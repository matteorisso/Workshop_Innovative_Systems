library verilog;
use verilog.vl_types.all;
entity test is
    generic(
        CLK             : integer := 2
    );
end test;
