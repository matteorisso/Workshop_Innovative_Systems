library ieee;
	use ieee.std_logic_1164.all;
	use ieee.numeric_std.all;

entity tb_conv_unit is

end tb_conv_unit;

architecture test of tb_conv_unit is

	component conv_unit is
		port(
			reset	:	in	std_logic;
			start	:	in	std_logic;
			done	:	in	std_logic;
			clk		:	in	std_logic;
			en_clk	:	in	std_logic;
			
			rf_in	:	in	std_logic_vector(83	downto 0);
			spw0_in	:	in	std_logic_vector(4	downto 0);
			spw1_in	:	in	std_logic_vector(4	downto 0);
			spw2_in	:	in	std_logic_vector(4	downto 0);
			spw3_in	:	in	std_logic_vector(4	downto 0);
			spw4_in	:	in	std_logic_vector(4	downto 0);
			spw5_in	:	in	std_logic_vector(4	downto 0);
			
			ofmap_0	:	out std_logic_vector(5	downto 0);
			ofmap_1	:	out std_logic_vector(5	downto 0);
			ofmap_2	:	out	std_logic_vector(5	downto 0);
			ofmap_3	:	out	std_logic_vector(5	downto 0);
			ofmap_4	:	out std_logic_vector(5	downto 0);
			ofmap_5	:	out std_logic_vector(5	downto 0)
		);
	end component;

	signal tb_reset		:	std_logic;
	signal tb_clk		:	std_logic;
	signal tb_start		:	std_logic;
	signal tb_done		:	std_logic;
	signal tb_en_clk	:	std_logic;
	
	signal tb_rf_in		:	std_logic_vector(0	to		83);
	signal tb_spw0_in	:	std_logic_vector(4	downto	0);
	signal tb_spw1_in	:	std_logic_vector(4	downto	0);
	signal tb_spw2_in	:	std_logic_vector(4	downto	0);
	signal tb_spw3_in	:	std_logic_vector(4	downto	0);
	signal tb_spw4_in	:	std_logic_vector(4	downto	0);
	signal tb_spw5_in	:	std_logic_vector(4	downto	0);
	
	signal tb_ofmap_0	:	std_logic_vector(5	downto	0);
	signal tb_ofmap_1	:	std_logic_vector(5	downto 	0);
	signal tb_ofmap_2	:	std_logic_vector(5	downto 	0);
	signal tb_ofmap_3	:	std_logic_vector(5	downto 	0);
	signal tb_ofmap_4	:	std_logic_vector(5	downto 	0);
	signal tb_ofmap_5	:	std_logic_vector(5	downto 	0);

begin

	dut : conv_unit
		port map(
			reset	=>	tb_reset,
			clk		=>	tb_clk,
			start	=>	tb_start,
			done	=>	tb_done,
			en_clk	=>	tb_en_clk,
			
			rf_in	=>	tb_rf_in,
			spw0_in	=>	tb_spw0_in,
			spw1_in	=>	tb_spw1_in,
			spw2_in	=>	tb_spw2_in,
			spw3_in	=>	tb_spw3_in,
			spw4_in	=>	tb_spw4_in,
			spw5_in	=>	tb_spw5_in,
			
			ofmap_0	=>	tb_ofmap_0,
			ofmap_1	=>	tb_ofmap_1,
			ofmap_2	=>	tb_ofmap_2,
			ofmap_3	=>	tb_ofmap_3,
			ofmap_4	=>	tb_ofmap_4,
			ofmap_5	=>	tb_ofmap_5
		);
	
	process -- clock generation at 500mhz.
	begin
		tb_clk <= '1';
		wait for 1 ns;
		tb_clk <= '0';
		wait for 1 ns;
	end process;
	
	process -- reset generation 
	begin
		tb_reset <= '0';
		wait for 4 ns;
		tb_reset <= '1';
		wait;
	end process;
	
	process 
	begin
		tb_start	<=	'0';
		tb_done		<=	'0';
		tb_en_clk	<=	'1';
		tb_rf_in	<=	(others	=> '1');
		tb_spw0_in	<=	(others	=> '1');
		tb_spw1_in	<=	(others	=> '1');
		tb_spw2_in	<=	(others	=> '1');
		tb_spw3_in	<=	(others	=> '1');
		tb_spw4_in	<=	(others	=> '1');
		tb_spw5_in	<=	(others	=> '1');
		
		wait for 6 ns;
		
		tb_start	<=	'1';
		
		wait for 2 ns;
		
		tb_start	<=	'0';
		
		wait for 2 ns;
		
		--load I5+I0 and row 0 of each filters.
		tb_rf_in(52	to		83)	<=	(others	=> '0'); --I0
		--tb_rf_in(52	to		83)	<=	"10101010111111000001100110000100";
		tb_rf_in(20	to		51)	<=	(others	=> '0'); --I5
		tb_rf_in(0	to		19)	<=	(others	=> '0'); 
		tb_spw0_in				<=	"01111";
		tb_spw1_in				<=	"11111";
		tb_spw2_in				<=	"10111";
		tb_spw3_in				<=	"11110";
		tb_spw4_in				<=	"11111";
		tb_spw5_in				<=	"11100";
		
		wait for 2 ns;
		--load I6+I1 and row 1 of each filters.
		tb_rf_in(52	to		83)	<=	(others	=> '0'); --I1
		tb_rf_in(20	to		51)	<=	(others	=> '0'); --I6
		tb_rf_in(0	to		19)	<=	(others	=> '0'); 
		tb_spw0_in				<=	"11111";
		tb_spw1_in				<=	"01011";
		tb_spw2_in				<=	"01111";
		tb_spw3_in				<=	"11111";
		tb_spw4_in				<=	"10000";
		tb_spw5_in				<=	"11110";
		
		wait for 2 ns;
		--load I7+I2 and row 2 of each filters.
		tb_rf_in(52	to		83)	<=	(others	=> '0'); --I2
		tb_rf_in(20	to		51)	<=	(others	=> '0'); --I7
		tb_rf_in(0	to		19)	<=	(others	=> '0'); 
		tb_spw0_in				<=	"01111";
		tb_spw1_in				<=	"00001";
		tb_spw2_in				<=	"11111";
		tb_spw3_in				<=	"11111";
		tb_spw4_in				<=	"10000";
		tb_spw5_in				<=	"01110";
		
		wait for 2 ns;
		--load I8+I3 and row 3 of each filters.
		tb_rf_in(52	to		83)	<=	(others	=> '0'); --I3
		tb_rf_in(20	to		51)	<=	(others	=> '0'); --I8
		tb_rf_in(0	to		19)	<=	(others	=> '0'); 
		tb_spw0_in				<=	"00000";
		tb_spw1_in				<=	"00000";
		tb_spw2_in				<=	"11000";
		tb_spw3_in				<=	"11111";
		tb_spw4_in				<=	"10000";
		tb_spw5_in				<=	"01110";
		
		wait for 2 ns;
		--load I9+I4 and row 4 of each filters.
		tb_rf_in(52	to		83)	<=	(others	=> '0'); --I4
		tb_rf_in(20	to		51)	<=	"00000000111111000000000000000000"; --I9
		tb_rf_in(0	to		19)	<=	(others	=> '0'); 
		tb_spw0_in				<=	"00000";
		tb_spw1_in				<=	"00001";
		tb_spw2_in				<=	"10000";
		tb_spw3_in				<=	"10000";
		tb_spw4_in				<=	"10000";
		tb_spw5_in				<=	"01111";
		
		wait for 384 ns;
		--load I15+I10.
		tb_rf_in(52	to		83)	<=	"00000000111111111111111100000000"; --I10
		tb_rf_in(20	to		51)	<=	"00000000000000000001111000000000"; --I15
		tb_rf_in(0	to		19)	<=	(others	=> '0'); 
		
		
		wait;
	end process;
	
end test;








