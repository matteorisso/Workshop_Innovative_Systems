library verilog;
use verilog.vl_types.all;
entity tb_fc is
end tb_fc;
