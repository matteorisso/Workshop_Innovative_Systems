library IEEE;
use IEEE.std_logic_1164.ALL;

entity wallace is
	port(
		in0,in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,in30,in31,in32,in33,in34,in35,in36,in37,in38,in39,in40,in41,in42,in43,in44,in45,in46,in47,in48,in49,in50,in51,in52,in53,in54,in55,in56,in57,in58,in59,in60,in61,in62,in63,in64,in65,in66,in67,in68,in69,in70,in71,in72,in73,in74,in75,in76,in77,in78,in79,in80,in81,in82,in83,in84,in85,in86,in87,in88,in89,in90,in91,in92,in93,in94,in95,in96,in97,in98,in99,in100,in101,in102,in103,in104,in105,in106,in107,in108,in109,in110,in111,in112,in113,in114,in115,in116,in117,in118,in119,in120,in121,in122,in123,in124,in125,in126,in127:IN std_logic_vector (127 downto 0);
clock,reset: IN std_logic;
		add1:OUT std_logic_vector(132 downto 0);
		add2:OUT std_logic_vector(132 downto 0);
		res:OUT std_logic_vector(1 downto 0));
end wallace;

architecture behavioural of wallace is
component HAff is
	 port(
		x,y,clock,reset:IN std_logic;
		s,c:OUT std_logic
	);
end component;
component FAff is
	port(
		cin,x,y,clock,reset:IN std_logic;
		s,cout:OUT std_logic
	);
end component;
component HA is
	 port(
		x,y:IN std_logic;
		s,c:OUT std_logic
	);
end component;
component FA is
	port(
		cin,x,y:IN std_logic;
		s,cout:OUT std_logic
	);
end component;

type bidimensional is array (0 to 389) of std_logic_vector(134 downto 0);
signal p:bidimensional;
begin
	p(0)(127 downto 0)<=in0;
	p(1)(127 downto 0)<=in1;
	p(2)(127 downto 0)<=in2;
	p(3)(127 downto 0)<=in3;
	p(4)(127 downto 0)<=in4;
	p(5)(127 downto 0)<=in5;
	p(6)(127 downto 0)<=in6;
	p(7)(127 downto 0)<=in7;
	p(8)(127 downto 0)<=in8;
	p(9)(127 downto 0)<=in9;
	p(10)(127 downto 0)<=in10;
	p(11)(127 downto 0)<=in11;
	p(12)(127 downto 0)<=in12;
	p(13)(127 downto 0)<=in13;
	p(14)(127 downto 0)<=in14;
	p(15)(127 downto 0)<=in15;
	p(16)(127 downto 0)<=in16;
	p(17)(127 downto 0)<=in17;
	p(18)(127 downto 0)<=in18;
	p(19)(127 downto 0)<=in19;
	p(20)(127 downto 0)<=in20;
	p(21)(127 downto 0)<=in21;
	p(22)(127 downto 0)<=in22;
	p(23)(127 downto 0)<=in23;
	p(24)(127 downto 0)<=in24;
	p(25)(127 downto 0)<=in25;
	p(26)(127 downto 0)<=in26;
	p(27)(127 downto 0)<=in27;
	p(28)(127 downto 0)<=in28;
	p(29)(127 downto 0)<=in29;
	p(30)(127 downto 0)<=in30;
	p(31)(127 downto 0)<=in31;
	p(32)(127 downto 0)<=in32;
	p(33)(127 downto 0)<=in33;
	p(34)(127 downto 0)<=in34;
	p(35)(127 downto 0)<=in35;
	p(36)(127 downto 0)<=in36;
	p(37)(127 downto 0)<=in37;
	p(38)(127 downto 0)<=in38;
	p(39)(127 downto 0)<=in39;
	p(40)(127 downto 0)<=in40;
	p(41)(127 downto 0)<=in41;
	p(42)(127 downto 0)<=in42;
	p(43)(127 downto 0)<=in43;
	p(44)(127 downto 0)<=in44;
	p(45)(127 downto 0)<=in45;
	p(46)(127 downto 0)<=in46;
	p(47)(127 downto 0)<=in47;
	p(48)(127 downto 0)<=in48;
	p(49)(127 downto 0)<=in49;
	p(50)(127 downto 0)<=in50;
	p(51)(127 downto 0)<=in51;
	p(52)(127 downto 0)<=in52;
	p(53)(127 downto 0)<=in53;
	p(54)(127 downto 0)<=in54;
	p(55)(127 downto 0)<=in55;
	p(56)(127 downto 0)<=in56;
	p(57)(127 downto 0)<=in57;
	p(58)(127 downto 0)<=in58;
	p(59)(127 downto 0)<=in59;
	p(60)(127 downto 0)<=in60;
	p(61)(127 downto 0)<=in61;
	p(62)(127 downto 0)<=in62;
	p(63)(127 downto 0)<=in63;
	p(64)(127 downto 0)<=in64;
	p(65)(127 downto 0)<=in65;
	p(66)(127 downto 0)<=in66;
	p(67)(127 downto 0)<=in67;
	p(68)(127 downto 0)<=in68;
	p(69)(127 downto 0)<=in69;
	p(70)(127 downto 0)<=in70;
	p(71)(127 downto 0)<=in71;
	p(72)(127 downto 0)<=in72;
	p(73)(127 downto 0)<=in73;
	p(74)(127 downto 0)<=in74;
	p(75)(127 downto 0)<=in75;
	p(76)(127 downto 0)<=in76;
	p(77)(127 downto 0)<=in77;
	p(78)(127 downto 0)<=in78;
	p(79)(127 downto 0)<=in79;
	p(80)(127 downto 0)<=in80;
	p(81)(127 downto 0)<=in81;
	p(82)(127 downto 0)<=in82;
	p(83)(127 downto 0)<=in83;
	p(84)(127 downto 0)<=in84;
	p(85)(127 downto 0)<=in85;
	p(86)(127 downto 0)<=in86;
	p(87)(127 downto 0)<=in87;
	p(88)(127 downto 0)<=in88;
	p(89)(127 downto 0)<=in89;
	p(90)(127 downto 0)<=in90;
	p(91)(127 downto 0)<=in91;
	p(92)(127 downto 0)<=in92;
	p(93)(127 downto 0)<=in93;
	p(94)(127 downto 0)<=in94;
	p(95)(127 downto 0)<=in95;
	p(96)(127 downto 0)<=in96;
	p(97)(127 downto 0)<=in97;
	p(98)(127 downto 0)<=in98;
	p(99)(127 downto 0)<=in99;
	p(100)(127 downto 0)<=in100;
	p(101)(127 downto 0)<=in101;
	p(102)(127 downto 0)<=in102;
	p(103)(127 downto 0)<=in103;
	p(104)(127 downto 0)<=in104;
	p(105)(127 downto 0)<=in105;
	p(106)(127 downto 0)<=in106;
	p(107)(127 downto 0)<=in107;
	p(108)(127 downto 0)<=in108;
	p(109)(127 downto 0)<=in109;
	p(110)(127 downto 0)<=in110;
	p(111)(127 downto 0)<=in111;
	p(112)(127 downto 0)<=in112;
	p(113)(127 downto 0)<=in113;
	p(114)(127 downto 0)<=in114;
	p(115)(127 downto 0)<=in115;
	p(116)(127 downto 0)<=in116;
	p(117)(127 downto 0)<=in117;
	p(118)(127 downto 0)<=in118;
	p(119)(127 downto 0)<=in119;
	p(120)(127 downto 0)<=in120;
	p(121)(127 downto 0)<=in121;
	p(122)(127 downto 0)<=in122;
	p(123)(127 downto 0)<=in123;
	p(124)(127 downto 0)<=in124;
	p(125)(127 downto 0)<=in125;
	p(126)(127 downto 0)<=in126;
	p(127)(127 downto 0)<=in127;
FA_ff_0:FAff port map(x=>p(0)(0),y=>p(1)(0),Cin=>p(2)(0),clock=>clock,reset=>reset,s=>p(128)(0),cout=>p(129)(1));
FA_ff_1:FAff port map(x=>p(0)(1),y=>p(1)(1),Cin=>p(2)(1),clock=>clock,reset=>reset,s=>p(128)(1),cout=>p(129)(2));
FA_ff_2:FAff port map(x=>p(0)(2),y=>p(1)(2),Cin=>p(2)(2),clock=>clock,reset=>reset,s=>p(128)(2),cout=>p(129)(3));
FA_ff_3:FAff port map(x=>p(0)(3),y=>p(1)(3),Cin=>p(2)(3),clock=>clock,reset=>reset,s=>p(128)(3),cout=>p(129)(4));
FA_ff_4:FAff port map(x=>p(0)(4),y=>p(1)(4),Cin=>p(2)(4),clock=>clock,reset=>reset,s=>p(128)(4),cout=>p(129)(5));
FA_ff_5:FAff port map(x=>p(0)(5),y=>p(1)(5),Cin=>p(2)(5),clock=>clock,reset=>reset,s=>p(128)(5),cout=>p(129)(6));
FA_ff_6:FAff port map(x=>p(0)(6),y=>p(1)(6),Cin=>p(2)(6),clock=>clock,reset=>reset,s=>p(128)(6),cout=>p(129)(7));
FA_ff_7:FAff port map(x=>p(0)(7),y=>p(1)(7),Cin=>p(2)(7),clock=>clock,reset=>reset,s=>p(128)(7),cout=>p(129)(8));
FA_ff_8:FAff port map(x=>p(0)(8),y=>p(1)(8),Cin=>p(2)(8),clock=>clock,reset=>reset,s=>p(128)(8),cout=>p(129)(9));
FA_ff_9:FAff port map(x=>p(0)(9),y=>p(1)(9),Cin=>p(2)(9),clock=>clock,reset=>reset,s=>p(128)(9),cout=>p(129)(10));
FA_ff_10:FAff port map(x=>p(0)(10),y=>p(1)(10),Cin=>p(2)(10),clock=>clock,reset=>reset,s=>p(128)(10),cout=>p(129)(11));
FA_ff_11:FAff port map(x=>p(0)(11),y=>p(1)(11),Cin=>p(2)(11),clock=>clock,reset=>reset,s=>p(128)(11),cout=>p(129)(12));
FA_ff_12:FAff port map(x=>p(0)(12),y=>p(1)(12),Cin=>p(2)(12),clock=>clock,reset=>reset,s=>p(128)(12),cout=>p(129)(13));
FA_ff_13:FAff port map(x=>p(0)(13),y=>p(1)(13),Cin=>p(2)(13),clock=>clock,reset=>reset,s=>p(128)(13),cout=>p(129)(14));
FA_ff_14:FAff port map(x=>p(0)(14),y=>p(1)(14),Cin=>p(2)(14),clock=>clock,reset=>reset,s=>p(128)(14),cout=>p(129)(15));
FA_ff_15:FAff port map(x=>p(0)(15),y=>p(1)(15),Cin=>p(2)(15),clock=>clock,reset=>reset,s=>p(128)(15),cout=>p(129)(16));
FA_ff_16:FAff port map(x=>p(0)(16),y=>p(1)(16),Cin=>p(2)(16),clock=>clock,reset=>reset,s=>p(128)(16),cout=>p(129)(17));
FA_ff_17:FAff port map(x=>p(0)(17),y=>p(1)(17),Cin=>p(2)(17),clock=>clock,reset=>reset,s=>p(128)(17),cout=>p(129)(18));
FA_ff_18:FAff port map(x=>p(0)(18),y=>p(1)(18),Cin=>p(2)(18),clock=>clock,reset=>reset,s=>p(128)(18),cout=>p(129)(19));
FA_ff_19:FAff port map(x=>p(0)(19),y=>p(1)(19),Cin=>p(2)(19),clock=>clock,reset=>reset,s=>p(128)(19),cout=>p(129)(20));
FA_ff_20:FAff port map(x=>p(0)(20),y=>p(1)(20),Cin=>p(2)(20),clock=>clock,reset=>reset,s=>p(128)(20),cout=>p(129)(21));
FA_ff_21:FAff port map(x=>p(0)(21),y=>p(1)(21),Cin=>p(2)(21),clock=>clock,reset=>reset,s=>p(128)(21),cout=>p(129)(22));
FA_ff_22:FAff port map(x=>p(0)(22),y=>p(1)(22),Cin=>p(2)(22),clock=>clock,reset=>reset,s=>p(128)(22),cout=>p(129)(23));
FA_ff_23:FAff port map(x=>p(0)(23),y=>p(1)(23),Cin=>p(2)(23),clock=>clock,reset=>reset,s=>p(128)(23),cout=>p(129)(24));
FA_ff_24:FAff port map(x=>p(0)(24),y=>p(1)(24),Cin=>p(2)(24),clock=>clock,reset=>reset,s=>p(128)(24),cout=>p(129)(25));
FA_ff_25:FAff port map(x=>p(0)(25),y=>p(1)(25),Cin=>p(2)(25),clock=>clock,reset=>reset,s=>p(128)(25),cout=>p(129)(26));
FA_ff_26:FAff port map(x=>p(0)(26),y=>p(1)(26),Cin=>p(2)(26),clock=>clock,reset=>reset,s=>p(128)(26),cout=>p(129)(27));
FA_ff_27:FAff port map(x=>p(0)(27),y=>p(1)(27),Cin=>p(2)(27),clock=>clock,reset=>reset,s=>p(128)(27),cout=>p(129)(28));
FA_ff_28:FAff port map(x=>p(0)(28),y=>p(1)(28),Cin=>p(2)(28),clock=>clock,reset=>reset,s=>p(128)(28),cout=>p(129)(29));
FA_ff_29:FAff port map(x=>p(0)(29),y=>p(1)(29),Cin=>p(2)(29),clock=>clock,reset=>reset,s=>p(128)(29),cout=>p(129)(30));
FA_ff_30:FAff port map(x=>p(0)(30),y=>p(1)(30),Cin=>p(2)(30),clock=>clock,reset=>reset,s=>p(128)(30),cout=>p(129)(31));
FA_ff_31:FAff port map(x=>p(0)(31),y=>p(1)(31),Cin=>p(2)(31),clock=>clock,reset=>reset,s=>p(128)(31),cout=>p(129)(32));
FA_ff_32:FAff port map(x=>p(0)(32),y=>p(1)(32),Cin=>p(2)(32),clock=>clock,reset=>reset,s=>p(128)(32),cout=>p(129)(33));
FA_ff_33:FAff port map(x=>p(0)(33),y=>p(1)(33),Cin=>p(2)(33),clock=>clock,reset=>reset,s=>p(128)(33),cout=>p(129)(34));
FA_ff_34:FAff port map(x=>p(0)(34),y=>p(1)(34),Cin=>p(2)(34),clock=>clock,reset=>reset,s=>p(128)(34),cout=>p(129)(35));
FA_ff_35:FAff port map(x=>p(0)(35),y=>p(1)(35),Cin=>p(2)(35),clock=>clock,reset=>reset,s=>p(128)(35),cout=>p(129)(36));
FA_ff_36:FAff port map(x=>p(0)(36),y=>p(1)(36),Cin=>p(2)(36),clock=>clock,reset=>reset,s=>p(128)(36),cout=>p(129)(37));
FA_ff_37:FAff port map(x=>p(0)(37),y=>p(1)(37),Cin=>p(2)(37),clock=>clock,reset=>reset,s=>p(128)(37),cout=>p(129)(38));
FA_ff_38:FAff port map(x=>p(0)(38),y=>p(1)(38),Cin=>p(2)(38),clock=>clock,reset=>reset,s=>p(128)(38),cout=>p(129)(39));
FA_ff_39:FAff port map(x=>p(0)(39),y=>p(1)(39),Cin=>p(2)(39),clock=>clock,reset=>reset,s=>p(128)(39),cout=>p(129)(40));
FA_ff_40:FAff port map(x=>p(0)(40),y=>p(1)(40),Cin=>p(2)(40),clock=>clock,reset=>reset,s=>p(128)(40),cout=>p(129)(41));
FA_ff_41:FAff port map(x=>p(0)(41),y=>p(1)(41),Cin=>p(2)(41),clock=>clock,reset=>reset,s=>p(128)(41),cout=>p(129)(42));
FA_ff_42:FAff port map(x=>p(0)(42),y=>p(1)(42),Cin=>p(2)(42),clock=>clock,reset=>reset,s=>p(128)(42),cout=>p(129)(43));
FA_ff_43:FAff port map(x=>p(0)(43),y=>p(1)(43),Cin=>p(2)(43),clock=>clock,reset=>reset,s=>p(128)(43),cout=>p(129)(44));
FA_ff_44:FAff port map(x=>p(0)(44),y=>p(1)(44),Cin=>p(2)(44),clock=>clock,reset=>reset,s=>p(128)(44),cout=>p(129)(45));
FA_ff_45:FAff port map(x=>p(0)(45),y=>p(1)(45),Cin=>p(2)(45),clock=>clock,reset=>reset,s=>p(128)(45),cout=>p(129)(46));
FA_ff_46:FAff port map(x=>p(0)(46),y=>p(1)(46),Cin=>p(2)(46),clock=>clock,reset=>reset,s=>p(128)(46),cout=>p(129)(47));
FA_ff_47:FAff port map(x=>p(0)(47),y=>p(1)(47),Cin=>p(2)(47),clock=>clock,reset=>reset,s=>p(128)(47),cout=>p(129)(48));
FA_ff_48:FAff port map(x=>p(0)(48),y=>p(1)(48),Cin=>p(2)(48),clock=>clock,reset=>reset,s=>p(128)(48),cout=>p(129)(49));
FA_ff_49:FAff port map(x=>p(0)(49),y=>p(1)(49),Cin=>p(2)(49),clock=>clock,reset=>reset,s=>p(128)(49),cout=>p(129)(50));
FA_ff_50:FAff port map(x=>p(0)(50),y=>p(1)(50),Cin=>p(2)(50),clock=>clock,reset=>reset,s=>p(128)(50),cout=>p(129)(51));
FA_ff_51:FAff port map(x=>p(0)(51),y=>p(1)(51),Cin=>p(2)(51),clock=>clock,reset=>reset,s=>p(128)(51),cout=>p(129)(52));
FA_ff_52:FAff port map(x=>p(0)(52),y=>p(1)(52),Cin=>p(2)(52),clock=>clock,reset=>reset,s=>p(128)(52),cout=>p(129)(53));
FA_ff_53:FAff port map(x=>p(0)(53),y=>p(1)(53),Cin=>p(2)(53),clock=>clock,reset=>reset,s=>p(128)(53),cout=>p(129)(54));
FA_ff_54:FAff port map(x=>p(0)(54),y=>p(1)(54),Cin=>p(2)(54),clock=>clock,reset=>reset,s=>p(128)(54),cout=>p(129)(55));
FA_ff_55:FAff port map(x=>p(0)(55),y=>p(1)(55),Cin=>p(2)(55),clock=>clock,reset=>reset,s=>p(128)(55),cout=>p(129)(56));
FA_ff_56:FAff port map(x=>p(0)(56),y=>p(1)(56),Cin=>p(2)(56),clock=>clock,reset=>reset,s=>p(128)(56),cout=>p(129)(57));
FA_ff_57:FAff port map(x=>p(0)(57),y=>p(1)(57),Cin=>p(2)(57),clock=>clock,reset=>reset,s=>p(128)(57),cout=>p(129)(58));
FA_ff_58:FAff port map(x=>p(0)(58),y=>p(1)(58),Cin=>p(2)(58),clock=>clock,reset=>reset,s=>p(128)(58),cout=>p(129)(59));
FA_ff_59:FAff port map(x=>p(0)(59),y=>p(1)(59),Cin=>p(2)(59),clock=>clock,reset=>reset,s=>p(128)(59),cout=>p(129)(60));
FA_ff_60:FAff port map(x=>p(0)(60),y=>p(1)(60),Cin=>p(2)(60),clock=>clock,reset=>reset,s=>p(128)(60),cout=>p(129)(61));
FA_ff_61:FAff port map(x=>p(0)(61),y=>p(1)(61),Cin=>p(2)(61),clock=>clock,reset=>reset,s=>p(128)(61),cout=>p(129)(62));
FA_ff_62:FAff port map(x=>p(0)(62),y=>p(1)(62),Cin=>p(2)(62),clock=>clock,reset=>reset,s=>p(128)(62),cout=>p(129)(63));
FA_ff_63:FAff port map(x=>p(0)(63),y=>p(1)(63),Cin=>p(2)(63),clock=>clock,reset=>reset,s=>p(128)(63),cout=>p(129)(64));
FA_ff_64:FAff port map(x=>p(0)(64),y=>p(1)(64),Cin=>p(2)(64),clock=>clock,reset=>reset,s=>p(128)(64),cout=>p(129)(65));
FA_ff_65:FAff port map(x=>p(0)(65),y=>p(1)(65),Cin=>p(2)(65),clock=>clock,reset=>reset,s=>p(128)(65),cout=>p(129)(66));
FA_ff_66:FAff port map(x=>p(0)(66),y=>p(1)(66),Cin=>p(2)(66),clock=>clock,reset=>reset,s=>p(128)(66),cout=>p(129)(67));
FA_ff_67:FAff port map(x=>p(0)(67),y=>p(1)(67),Cin=>p(2)(67),clock=>clock,reset=>reset,s=>p(128)(67),cout=>p(129)(68));
FA_ff_68:FAff port map(x=>p(0)(68),y=>p(1)(68),Cin=>p(2)(68),clock=>clock,reset=>reset,s=>p(128)(68),cout=>p(129)(69));
FA_ff_69:FAff port map(x=>p(0)(69),y=>p(1)(69),Cin=>p(2)(69),clock=>clock,reset=>reset,s=>p(128)(69),cout=>p(129)(70));
FA_ff_70:FAff port map(x=>p(0)(70),y=>p(1)(70),Cin=>p(2)(70),clock=>clock,reset=>reset,s=>p(128)(70),cout=>p(129)(71));
FA_ff_71:FAff port map(x=>p(0)(71),y=>p(1)(71),Cin=>p(2)(71),clock=>clock,reset=>reset,s=>p(128)(71),cout=>p(129)(72));
FA_ff_72:FAff port map(x=>p(0)(72),y=>p(1)(72),Cin=>p(2)(72),clock=>clock,reset=>reset,s=>p(128)(72),cout=>p(129)(73));
FA_ff_73:FAff port map(x=>p(0)(73),y=>p(1)(73),Cin=>p(2)(73),clock=>clock,reset=>reset,s=>p(128)(73),cout=>p(129)(74));
FA_ff_74:FAff port map(x=>p(0)(74),y=>p(1)(74),Cin=>p(2)(74),clock=>clock,reset=>reset,s=>p(128)(74),cout=>p(129)(75));
FA_ff_75:FAff port map(x=>p(0)(75),y=>p(1)(75),Cin=>p(2)(75),clock=>clock,reset=>reset,s=>p(128)(75),cout=>p(129)(76));
FA_ff_76:FAff port map(x=>p(0)(76),y=>p(1)(76),Cin=>p(2)(76),clock=>clock,reset=>reset,s=>p(128)(76),cout=>p(129)(77));
FA_ff_77:FAff port map(x=>p(0)(77),y=>p(1)(77),Cin=>p(2)(77),clock=>clock,reset=>reset,s=>p(128)(77),cout=>p(129)(78));
FA_ff_78:FAff port map(x=>p(0)(78),y=>p(1)(78),Cin=>p(2)(78),clock=>clock,reset=>reset,s=>p(128)(78),cout=>p(129)(79));
FA_ff_79:FAff port map(x=>p(0)(79),y=>p(1)(79),Cin=>p(2)(79),clock=>clock,reset=>reset,s=>p(128)(79),cout=>p(129)(80));
FA_ff_80:FAff port map(x=>p(0)(80),y=>p(1)(80),Cin=>p(2)(80),clock=>clock,reset=>reset,s=>p(128)(80),cout=>p(129)(81));
FA_ff_81:FAff port map(x=>p(0)(81),y=>p(1)(81),Cin=>p(2)(81),clock=>clock,reset=>reset,s=>p(128)(81),cout=>p(129)(82));
FA_ff_82:FAff port map(x=>p(0)(82),y=>p(1)(82),Cin=>p(2)(82),clock=>clock,reset=>reset,s=>p(128)(82),cout=>p(129)(83));
FA_ff_83:FAff port map(x=>p(0)(83),y=>p(1)(83),Cin=>p(2)(83),clock=>clock,reset=>reset,s=>p(128)(83),cout=>p(129)(84));
FA_ff_84:FAff port map(x=>p(0)(84),y=>p(1)(84),Cin=>p(2)(84),clock=>clock,reset=>reset,s=>p(128)(84),cout=>p(129)(85));
FA_ff_85:FAff port map(x=>p(0)(85),y=>p(1)(85),Cin=>p(2)(85),clock=>clock,reset=>reset,s=>p(128)(85),cout=>p(129)(86));
FA_ff_86:FAff port map(x=>p(0)(86),y=>p(1)(86),Cin=>p(2)(86),clock=>clock,reset=>reset,s=>p(128)(86),cout=>p(129)(87));
FA_ff_87:FAff port map(x=>p(0)(87),y=>p(1)(87),Cin=>p(2)(87),clock=>clock,reset=>reset,s=>p(128)(87),cout=>p(129)(88));
FA_ff_88:FAff port map(x=>p(0)(88),y=>p(1)(88),Cin=>p(2)(88),clock=>clock,reset=>reset,s=>p(128)(88),cout=>p(129)(89));
FA_ff_89:FAff port map(x=>p(0)(89),y=>p(1)(89),Cin=>p(2)(89),clock=>clock,reset=>reset,s=>p(128)(89),cout=>p(129)(90));
FA_ff_90:FAff port map(x=>p(0)(90),y=>p(1)(90),Cin=>p(2)(90),clock=>clock,reset=>reset,s=>p(128)(90),cout=>p(129)(91));
FA_ff_91:FAff port map(x=>p(0)(91),y=>p(1)(91),Cin=>p(2)(91),clock=>clock,reset=>reset,s=>p(128)(91),cout=>p(129)(92));
FA_ff_92:FAff port map(x=>p(0)(92),y=>p(1)(92),Cin=>p(2)(92),clock=>clock,reset=>reset,s=>p(128)(92),cout=>p(129)(93));
FA_ff_93:FAff port map(x=>p(0)(93),y=>p(1)(93),Cin=>p(2)(93),clock=>clock,reset=>reset,s=>p(128)(93),cout=>p(129)(94));
FA_ff_94:FAff port map(x=>p(0)(94),y=>p(1)(94),Cin=>p(2)(94),clock=>clock,reset=>reset,s=>p(128)(94),cout=>p(129)(95));
FA_ff_95:FAff port map(x=>p(0)(95),y=>p(1)(95),Cin=>p(2)(95),clock=>clock,reset=>reset,s=>p(128)(95),cout=>p(129)(96));
FA_ff_96:FAff port map(x=>p(0)(96),y=>p(1)(96),Cin=>p(2)(96),clock=>clock,reset=>reset,s=>p(128)(96),cout=>p(129)(97));
FA_ff_97:FAff port map(x=>p(0)(97),y=>p(1)(97),Cin=>p(2)(97),clock=>clock,reset=>reset,s=>p(128)(97),cout=>p(129)(98));
FA_ff_98:FAff port map(x=>p(0)(98),y=>p(1)(98),Cin=>p(2)(98),clock=>clock,reset=>reset,s=>p(128)(98),cout=>p(129)(99));
FA_ff_99:FAff port map(x=>p(0)(99),y=>p(1)(99),Cin=>p(2)(99),clock=>clock,reset=>reset,s=>p(128)(99),cout=>p(129)(100));
FA_ff_100:FAff port map(x=>p(0)(100),y=>p(1)(100),Cin=>p(2)(100),clock=>clock,reset=>reset,s=>p(128)(100),cout=>p(129)(101));
FA_ff_101:FAff port map(x=>p(0)(101),y=>p(1)(101),Cin=>p(2)(101),clock=>clock,reset=>reset,s=>p(128)(101),cout=>p(129)(102));
FA_ff_102:FAff port map(x=>p(0)(102),y=>p(1)(102),Cin=>p(2)(102),clock=>clock,reset=>reset,s=>p(128)(102),cout=>p(129)(103));
FA_ff_103:FAff port map(x=>p(0)(103),y=>p(1)(103),Cin=>p(2)(103),clock=>clock,reset=>reset,s=>p(128)(103),cout=>p(129)(104));
FA_ff_104:FAff port map(x=>p(0)(104),y=>p(1)(104),Cin=>p(2)(104),clock=>clock,reset=>reset,s=>p(128)(104),cout=>p(129)(105));
FA_ff_105:FAff port map(x=>p(0)(105),y=>p(1)(105),Cin=>p(2)(105),clock=>clock,reset=>reset,s=>p(128)(105),cout=>p(129)(106));
FA_ff_106:FAff port map(x=>p(0)(106),y=>p(1)(106),Cin=>p(2)(106),clock=>clock,reset=>reset,s=>p(128)(106),cout=>p(129)(107));
FA_ff_107:FAff port map(x=>p(0)(107),y=>p(1)(107),Cin=>p(2)(107),clock=>clock,reset=>reset,s=>p(128)(107),cout=>p(129)(108));
FA_ff_108:FAff port map(x=>p(0)(108),y=>p(1)(108),Cin=>p(2)(108),clock=>clock,reset=>reset,s=>p(128)(108),cout=>p(129)(109));
FA_ff_109:FAff port map(x=>p(0)(109),y=>p(1)(109),Cin=>p(2)(109),clock=>clock,reset=>reset,s=>p(128)(109),cout=>p(129)(110));
FA_ff_110:FAff port map(x=>p(0)(110),y=>p(1)(110),Cin=>p(2)(110),clock=>clock,reset=>reset,s=>p(128)(110),cout=>p(129)(111));
FA_ff_111:FAff port map(x=>p(0)(111),y=>p(1)(111),Cin=>p(2)(111),clock=>clock,reset=>reset,s=>p(128)(111),cout=>p(129)(112));
FA_ff_112:FAff port map(x=>p(0)(112),y=>p(1)(112),Cin=>p(2)(112),clock=>clock,reset=>reset,s=>p(128)(112),cout=>p(129)(113));
FA_ff_113:FAff port map(x=>p(0)(113),y=>p(1)(113),Cin=>p(2)(113),clock=>clock,reset=>reset,s=>p(128)(113),cout=>p(129)(114));
FA_ff_114:FAff port map(x=>p(0)(114),y=>p(1)(114),Cin=>p(2)(114),clock=>clock,reset=>reset,s=>p(128)(114),cout=>p(129)(115));
FA_ff_115:FAff port map(x=>p(0)(115),y=>p(1)(115),Cin=>p(2)(115),clock=>clock,reset=>reset,s=>p(128)(115),cout=>p(129)(116));
FA_ff_116:FAff port map(x=>p(0)(116),y=>p(1)(116),Cin=>p(2)(116),clock=>clock,reset=>reset,s=>p(128)(116),cout=>p(129)(117));
FA_ff_117:FAff port map(x=>p(0)(117),y=>p(1)(117),Cin=>p(2)(117),clock=>clock,reset=>reset,s=>p(128)(117),cout=>p(129)(118));
FA_ff_118:FAff port map(x=>p(0)(118),y=>p(1)(118),Cin=>p(2)(118),clock=>clock,reset=>reset,s=>p(128)(118),cout=>p(129)(119));
FA_ff_119:FAff port map(x=>p(0)(119),y=>p(1)(119),Cin=>p(2)(119),clock=>clock,reset=>reset,s=>p(128)(119),cout=>p(129)(120));
FA_ff_120:FAff port map(x=>p(0)(120),y=>p(1)(120),Cin=>p(2)(120),clock=>clock,reset=>reset,s=>p(128)(120),cout=>p(129)(121));
FA_ff_121:FAff port map(x=>p(0)(121),y=>p(1)(121),Cin=>p(2)(121),clock=>clock,reset=>reset,s=>p(128)(121),cout=>p(129)(122));
FA_ff_122:FAff port map(x=>p(0)(122),y=>p(1)(122),Cin=>p(2)(122),clock=>clock,reset=>reset,s=>p(128)(122),cout=>p(129)(123));
FA_ff_123:FAff port map(x=>p(0)(123),y=>p(1)(123),Cin=>p(2)(123),clock=>clock,reset=>reset,s=>p(128)(123),cout=>p(129)(124));
FA_ff_124:FAff port map(x=>p(0)(124),y=>p(1)(124),Cin=>p(2)(124),clock=>clock,reset=>reset,s=>p(128)(124),cout=>p(129)(125));
FA_ff_125:FAff port map(x=>p(0)(125),y=>p(1)(125),Cin=>p(2)(125),clock=>clock,reset=>reset,s=>p(128)(125),cout=>p(129)(126));
FA_ff_126:FAff port map(x=>p(0)(126),y=>p(1)(126),Cin=>p(2)(126),clock=>clock,reset=>reset,s=>p(128)(126),cout=>p(129)(127));
FA_ff_127:FAff port map(x=>p(0)(127),y=>p(1)(127),Cin=>p(2)(127),clock=>clock,reset=>reset,s=>p(128)(127),cout=>p(129)(128));
FA_ff_128:FAff port map(x=>p(3)(0),y=>p(4)(0),Cin=>p(5)(0),clock=>clock,reset=>reset,s=>p(130)(0),cout=>p(131)(1));
FA_ff_129:FAff port map(x=>p(3)(1),y=>p(4)(1),Cin=>p(5)(1),clock=>clock,reset=>reset,s=>p(130)(1),cout=>p(131)(2));
FA_ff_130:FAff port map(x=>p(3)(2),y=>p(4)(2),Cin=>p(5)(2),clock=>clock,reset=>reset,s=>p(130)(2),cout=>p(131)(3));
FA_ff_131:FAff port map(x=>p(3)(3),y=>p(4)(3),Cin=>p(5)(3),clock=>clock,reset=>reset,s=>p(130)(3),cout=>p(131)(4));
FA_ff_132:FAff port map(x=>p(3)(4),y=>p(4)(4),Cin=>p(5)(4),clock=>clock,reset=>reset,s=>p(130)(4),cout=>p(131)(5));
FA_ff_133:FAff port map(x=>p(3)(5),y=>p(4)(5),Cin=>p(5)(5),clock=>clock,reset=>reset,s=>p(130)(5),cout=>p(131)(6));
FA_ff_134:FAff port map(x=>p(3)(6),y=>p(4)(6),Cin=>p(5)(6),clock=>clock,reset=>reset,s=>p(130)(6),cout=>p(131)(7));
FA_ff_135:FAff port map(x=>p(3)(7),y=>p(4)(7),Cin=>p(5)(7),clock=>clock,reset=>reset,s=>p(130)(7),cout=>p(131)(8));
FA_ff_136:FAff port map(x=>p(3)(8),y=>p(4)(8),Cin=>p(5)(8),clock=>clock,reset=>reset,s=>p(130)(8),cout=>p(131)(9));
FA_ff_137:FAff port map(x=>p(3)(9),y=>p(4)(9),Cin=>p(5)(9),clock=>clock,reset=>reset,s=>p(130)(9),cout=>p(131)(10));
FA_ff_138:FAff port map(x=>p(3)(10),y=>p(4)(10),Cin=>p(5)(10),clock=>clock,reset=>reset,s=>p(130)(10),cout=>p(131)(11));
FA_ff_139:FAff port map(x=>p(3)(11),y=>p(4)(11),Cin=>p(5)(11),clock=>clock,reset=>reset,s=>p(130)(11),cout=>p(131)(12));
FA_ff_140:FAff port map(x=>p(3)(12),y=>p(4)(12),Cin=>p(5)(12),clock=>clock,reset=>reset,s=>p(130)(12),cout=>p(131)(13));
FA_ff_141:FAff port map(x=>p(3)(13),y=>p(4)(13),Cin=>p(5)(13),clock=>clock,reset=>reset,s=>p(130)(13),cout=>p(131)(14));
FA_ff_142:FAff port map(x=>p(3)(14),y=>p(4)(14),Cin=>p(5)(14),clock=>clock,reset=>reset,s=>p(130)(14),cout=>p(131)(15));
FA_ff_143:FAff port map(x=>p(3)(15),y=>p(4)(15),Cin=>p(5)(15),clock=>clock,reset=>reset,s=>p(130)(15),cout=>p(131)(16));
FA_ff_144:FAff port map(x=>p(3)(16),y=>p(4)(16),Cin=>p(5)(16),clock=>clock,reset=>reset,s=>p(130)(16),cout=>p(131)(17));
FA_ff_145:FAff port map(x=>p(3)(17),y=>p(4)(17),Cin=>p(5)(17),clock=>clock,reset=>reset,s=>p(130)(17),cout=>p(131)(18));
FA_ff_146:FAff port map(x=>p(3)(18),y=>p(4)(18),Cin=>p(5)(18),clock=>clock,reset=>reset,s=>p(130)(18),cout=>p(131)(19));
FA_ff_147:FAff port map(x=>p(3)(19),y=>p(4)(19),Cin=>p(5)(19),clock=>clock,reset=>reset,s=>p(130)(19),cout=>p(131)(20));
FA_ff_148:FAff port map(x=>p(3)(20),y=>p(4)(20),Cin=>p(5)(20),clock=>clock,reset=>reset,s=>p(130)(20),cout=>p(131)(21));
FA_ff_149:FAff port map(x=>p(3)(21),y=>p(4)(21),Cin=>p(5)(21),clock=>clock,reset=>reset,s=>p(130)(21),cout=>p(131)(22));
FA_ff_150:FAff port map(x=>p(3)(22),y=>p(4)(22),Cin=>p(5)(22),clock=>clock,reset=>reset,s=>p(130)(22),cout=>p(131)(23));
FA_ff_151:FAff port map(x=>p(3)(23),y=>p(4)(23),Cin=>p(5)(23),clock=>clock,reset=>reset,s=>p(130)(23),cout=>p(131)(24));
FA_ff_152:FAff port map(x=>p(3)(24),y=>p(4)(24),Cin=>p(5)(24),clock=>clock,reset=>reset,s=>p(130)(24),cout=>p(131)(25));
FA_ff_153:FAff port map(x=>p(3)(25),y=>p(4)(25),Cin=>p(5)(25),clock=>clock,reset=>reset,s=>p(130)(25),cout=>p(131)(26));
FA_ff_154:FAff port map(x=>p(3)(26),y=>p(4)(26),Cin=>p(5)(26),clock=>clock,reset=>reset,s=>p(130)(26),cout=>p(131)(27));
FA_ff_155:FAff port map(x=>p(3)(27),y=>p(4)(27),Cin=>p(5)(27),clock=>clock,reset=>reset,s=>p(130)(27),cout=>p(131)(28));
FA_ff_156:FAff port map(x=>p(3)(28),y=>p(4)(28),Cin=>p(5)(28),clock=>clock,reset=>reset,s=>p(130)(28),cout=>p(131)(29));
FA_ff_157:FAff port map(x=>p(3)(29),y=>p(4)(29),Cin=>p(5)(29),clock=>clock,reset=>reset,s=>p(130)(29),cout=>p(131)(30));
FA_ff_158:FAff port map(x=>p(3)(30),y=>p(4)(30),Cin=>p(5)(30),clock=>clock,reset=>reset,s=>p(130)(30),cout=>p(131)(31));
FA_ff_159:FAff port map(x=>p(3)(31),y=>p(4)(31),Cin=>p(5)(31),clock=>clock,reset=>reset,s=>p(130)(31),cout=>p(131)(32));
FA_ff_160:FAff port map(x=>p(3)(32),y=>p(4)(32),Cin=>p(5)(32),clock=>clock,reset=>reset,s=>p(130)(32),cout=>p(131)(33));
FA_ff_161:FAff port map(x=>p(3)(33),y=>p(4)(33),Cin=>p(5)(33),clock=>clock,reset=>reset,s=>p(130)(33),cout=>p(131)(34));
FA_ff_162:FAff port map(x=>p(3)(34),y=>p(4)(34),Cin=>p(5)(34),clock=>clock,reset=>reset,s=>p(130)(34),cout=>p(131)(35));
FA_ff_163:FAff port map(x=>p(3)(35),y=>p(4)(35),Cin=>p(5)(35),clock=>clock,reset=>reset,s=>p(130)(35),cout=>p(131)(36));
FA_ff_164:FAff port map(x=>p(3)(36),y=>p(4)(36),Cin=>p(5)(36),clock=>clock,reset=>reset,s=>p(130)(36),cout=>p(131)(37));
FA_ff_165:FAff port map(x=>p(3)(37),y=>p(4)(37),Cin=>p(5)(37),clock=>clock,reset=>reset,s=>p(130)(37),cout=>p(131)(38));
FA_ff_166:FAff port map(x=>p(3)(38),y=>p(4)(38),Cin=>p(5)(38),clock=>clock,reset=>reset,s=>p(130)(38),cout=>p(131)(39));
FA_ff_167:FAff port map(x=>p(3)(39),y=>p(4)(39),Cin=>p(5)(39),clock=>clock,reset=>reset,s=>p(130)(39),cout=>p(131)(40));
FA_ff_168:FAff port map(x=>p(3)(40),y=>p(4)(40),Cin=>p(5)(40),clock=>clock,reset=>reset,s=>p(130)(40),cout=>p(131)(41));
FA_ff_169:FAff port map(x=>p(3)(41),y=>p(4)(41),Cin=>p(5)(41),clock=>clock,reset=>reset,s=>p(130)(41),cout=>p(131)(42));
FA_ff_170:FAff port map(x=>p(3)(42),y=>p(4)(42),Cin=>p(5)(42),clock=>clock,reset=>reset,s=>p(130)(42),cout=>p(131)(43));
FA_ff_171:FAff port map(x=>p(3)(43),y=>p(4)(43),Cin=>p(5)(43),clock=>clock,reset=>reset,s=>p(130)(43),cout=>p(131)(44));
FA_ff_172:FAff port map(x=>p(3)(44),y=>p(4)(44),Cin=>p(5)(44),clock=>clock,reset=>reset,s=>p(130)(44),cout=>p(131)(45));
FA_ff_173:FAff port map(x=>p(3)(45),y=>p(4)(45),Cin=>p(5)(45),clock=>clock,reset=>reset,s=>p(130)(45),cout=>p(131)(46));
FA_ff_174:FAff port map(x=>p(3)(46),y=>p(4)(46),Cin=>p(5)(46),clock=>clock,reset=>reset,s=>p(130)(46),cout=>p(131)(47));
FA_ff_175:FAff port map(x=>p(3)(47),y=>p(4)(47),Cin=>p(5)(47),clock=>clock,reset=>reset,s=>p(130)(47),cout=>p(131)(48));
FA_ff_176:FAff port map(x=>p(3)(48),y=>p(4)(48),Cin=>p(5)(48),clock=>clock,reset=>reset,s=>p(130)(48),cout=>p(131)(49));
FA_ff_177:FAff port map(x=>p(3)(49),y=>p(4)(49),Cin=>p(5)(49),clock=>clock,reset=>reset,s=>p(130)(49),cout=>p(131)(50));
FA_ff_178:FAff port map(x=>p(3)(50),y=>p(4)(50),Cin=>p(5)(50),clock=>clock,reset=>reset,s=>p(130)(50),cout=>p(131)(51));
FA_ff_179:FAff port map(x=>p(3)(51),y=>p(4)(51),Cin=>p(5)(51),clock=>clock,reset=>reset,s=>p(130)(51),cout=>p(131)(52));
FA_ff_180:FAff port map(x=>p(3)(52),y=>p(4)(52),Cin=>p(5)(52),clock=>clock,reset=>reset,s=>p(130)(52),cout=>p(131)(53));
FA_ff_181:FAff port map(x=>p(3)(53),y=>p(4)(53),Cin=>p(5)(53),clock=>clock,reset=>reset,s=>p(130)(53),cout=>p(131)(54));
FA_ff_182:FAff port map(x=>p(3)(54),y=>p(4)(54),Cin=>p(5)(54),clock=>clock,reset=>reset,s=>p(130)(54),cout=>p(131)(55));
FA_ff_183:FAff port map(x=>p(3)(55),y=>p(4)(55),Cin=>p(5)(55),clock=>clock,reset=>reset,s=>p(130)(55),cout=>p(131)(56));
FA_ff_184:FAff port map(x=>p(3)(56),y=>p(4)(56),Cin=>p(5)(56),clock=>clock,reset=>reset,s=>p(130)(56),cout=>p(131)(57));
FA_ff_185:FAff port map(x=>p(3)(57),y=>p(4)(57),Cin=>p(5)(57),clock=>clock,reset=>reset,s=>p(130)(57),cout=>p(131)(58));
FA_ff_186:FAff port map(x=>p(3)(58),y=>p(4)(58),Cin=>p(5)(58),clock=>clock,reset=>reset,s=>p(130)(58),cout=>p(131)(59));
FA_ff_187:FAff port map(x=>p(3)(59),y=>p(4)(59),Cin=>p(5)(59),clock=>clock,reset=>reset,s=>p(130)(59),cout=>p(131)(60));
FA_ff_188:FAff port map(x=>p(3)(60),y=>p(4)(60),Cin=>p(5)(60),clock=>clock,reset=>reset,s=>p(130)(60),cout=>p(131)(61));
FA_ff_189:FAff port map(x=>p(3)(61),y=>p(4)(61),Cin=>p(5)(61),clock=>clock,reset=>reset,s=>p(130)(61),cout=>p(131)(62));
FA_ff_190:FAff port map(x=>p(3)(62),y=>p(4)(62),Cin=>p(5)(62),clock=>clock,reset=>reset,s=>p(130)(62),cout=>p(131)(63));
FA_ff_191:FAff port map(x=>p(3)(63),y=>p(4)(63),Cin=>p(5)(63),clock=>clock,reset=>reset,s=>p(130)(63),cout=>p(131)(64));
FA_ff_192:FAff port map(x=>p(3)(64),y=>p(4)(64),Cin=>p(5)(64),clock=>clock,reset=>reset,s=>p(130)(64),cout=>p(131)(65));
FA_ff_193:FAff port map(x=>p(3)(65),y=>p(4)(65),Cin=>p(5)(65),clock=>clock,reset=>reset,s=>p(130)(65),cout=>p(131)(66));
FA_ff_194:FAff port map(x=>p(3)(66),y=>p(4)(66),Cin=>p(5)(66),clock=>clock,reset=>reset,s=>p(130)(66),cout=>p(131)(67));
FA_ff_195:FAff port map(x=>p(3)(67),y=>p(4)(67),Cin=>p(5)(67),clock=>clock,reset=>reset,s=>p(130)(67),cout=>p(131)(68));
FA_ff_196:FAff port map(x=>p(3)(68),y=>p(4)(68),Cin=>p(5)(68),clock=>clock,reset=>reset,s=>p(130)(68),cout=>p(131)(69));
FA_ff_197:FAff port map(x=>p(3)(69),y=>p(4)(69),Cin=>p(5)(69),clock=>clock,reset=>reset,s=>p(130)(69),cout=>p(131)(70));
FA_ff_198:FAff port map(x=>p(3)(70),y=>p(4)(70),Cin=>p(5)(70),clock=>clock,reset=>reset,s=>p(130)(70),cout=>p(131)(71));
FA_ff_199:FAff port map(x=>p(3)(71),y=>p(4)(71),Cin=>p(5)(71),clock=>clock,reset=>reset,s=>p(130)(71),cout=>p(131)(72));
FA_ff_200:FAff port map(x=>p(3)(72),y=>p(4)(72),Cin=>p(5)(72),clock=>clock,reset=>reset,s=>p(130)(72),cout=>p(131)(73));
FA_ff_201:FAff port map(x=>p(3)(73),y=>p(4)(73),Cin=>p(5)(73),clock=>clock,reset=>reset,s=>p(130)(73),cout=>p(131)(74));
FA_ff_202:FAff port map(x=>p(3)(74),y=>p(4)(74),Cin=>p(5)(74),clock=>clock,reset=>reset,s=>p(130)(74),cout=>p(131)(75));
FA_ff_203:FAff port map(x=>p(3)(75),y=>p(4)(75),Cin=>p(5)(75),clock=>clock,reset=>reset,s=>p(130)(75),cout=>p(131)(76));
FA_ff_204:FAff port map(x=>p(3)(76),y=>p(4)(76),Cin=>p(5)(76),clock=>clock,reset=>reset,s=>p(130)(76),cout=>p(131)(77));
FA_ff_205:FAff port map(x=>p(3)(77),y=>p(4)(77),Cin=>p(5)(77),clock=>clock,reset=>reset,s=>p(130)(77),cout=>p(131)(78));
FA_ff_206:FAff port map(x=>p(3)(78),y=>p(4)(78),Cin=>p(5)(78),clock=>clock,reset=>reset,s=>p(130)(78),cout=>p(131)(79));
FA_ff_207:FAff port map(x=>p(3)(79),y=>p(4)(79),Cin=>p(5)(79),clock=>clock,reset=>reset,s=>p(130)(79),cout=>p(131)(80));
FA_ff_208:FAff port map(x=>p(3)(80),y=>p(4)(80),Cin=>p(5)(80),clock=>clock,reset=>reset,s=>p(130)(80),cout=>p(131)(81));
FA_ff_209:FAff port map(x=>p(3)(81),y=>p(4)(81),Cin=>p(5)(81),clock=>clock,reset=>reset,s=>p(130)(81),cout=>p(131)(82));
FA_ff_210:FAff port map(x=>p(3)(82),y=>p(4)(82),Cin=>p(5)(82),clock=>clock,reset=>reset,s=>p(130)(82),cout=>p(131)(83));
FA_ff_211:FAff port map(x=>p(3)(83),y=>p(4)(83),Cin=>p(5)(83),clock=>clock,reset=>reset,s=>p(130)(83),cout=>p(131)(84));
FA_ff_212:FAff port map(x=>p(3)(84),y=>p(4)(84),Cin=>p(5)(84),clock=>clock,reset=>reset,s=>p(130)(84),cout=>p(131)(85));
FA_ff_213:FAff port map(x=>p(3)(85),y=>p(4)(85),Cin=>p(5)(85),clock=>clock,reset=>reset,s=>p(130)(85),cout=>p(131)(86));
FA_ff_214:FAff port map(x=>p(3)(86),y=>p(4)(86),Cin=>p(5)(86),clock=>clock,reset=>reset,s=>p(130)(86),cout=>p(131)(87));
FA_ff_215:FAff port map(x=>p(3)(87),y=>p(4)(87),Cin=>p(5)(87),clock=>clock,reset=>reset,s=>p(130)(87),cout=>p(131)(88));
FA_ff_216:FAff port map(x=>p(3)(88),y=>p(4)(88),Cin=>p(5)(88),clock=>clock,reset=>reset,s=>p(130)(88),cout=>p(131)(89));
FA_ff_217:FAff port map(x=>p(3)(89),y=>p(4)(89),Cin=>p(5)(89),clock=>clock,reset=>reset,s=>p(130)(89),cout=>p(131)(90));
FA_ff_218:FAff port map(x=>p(3)(90),y=>p(4)(90),Cin=>p(5)(90),clock=>clock,reset=>reset,s=>p(130)(90),cout=>p(131)(91));
FA_ff_219:FAff port map(x=>p(3)(91),y=>p(4)(91),Cin=>p(5)(91),clock=>clock,reset=>reset,s=>p(130)(91),cout=>p(131)(92));
FA_ff_220:FAff port map(x=>p(3)(92),y=>p(4)(92),Cin=>p(5)(92),clock=>clock,reset=>reset,s=>p(130)(92),cout=>p(131)(93));
FA_ff_221:FAff port map(x=>p(3)(93),y=>p(4)(93),Cin=>p(5)(93),clock=>clock,reset=>reset,s=>p(130)(93),cout=>p(131)(94));
FA_ff_222:FAff port map(x=>p(3)(94),y=>p(4)(94),Cin=>p(5)(94),clock=>clock,reset=>reset,s=>p(130)(94),cout=>p(131)(95));
FA_ff_223:FAff port map(x=>p(3)(95),y=>p(4)(95),Cin=>p(5)(95),clock=>clock,reset=>reset,s=>p(130)(95),cout=>p(131)(96));
FA_ff_224:FAff port map(x=>p(3)(96),y=>p(4)(96),Cin=>p(5)(96),clock=>clock,reset=>reset,s=>p(130)(96),cout=>p(131)(97));
FA_ff_225:FAff port map(x=>p(3)(97),y=>p(4)(97),Cin=>p(5)(97),clock=>clock,reset=>reset,s=>p(130)(97),cout=>p(131)(98));
FA_ff_226:FAff port map(x=>p(3)(98),y=>p(4)(98),Cin=>p(5)(98),clock=>clock,reset=>reset,s=>p(130)(98),cout=>p(131)(99));
FA_ff_227:FAff port map(x=>p(3)(99),y=>p(4)(99),Cin=>p(5)(99),clock=>clock,reset=>reset,s=>p(130)(99),cout=>p(131)(100));
FA_ff_228:FAff port map(x=>p(3)(100),y=>p(4)(100),Cin=>p(5)(100),clock=>clock,reset=>reset,s=>p(130)(100),cout=>p(131)(101));
FA_ff_229:FAff port map(x=>p(3)(101),y=>p(4)(101),Cin=>p(5)(101),clock=>clock,reset=>reset,s=>p(130)(101),cout=>p(131)(102));
FA_ff_230:FAff port map(x=>p(3)(102),y=>p(4)(102),Cin=>p(5)(102),clock=>clock,reset=>reset,s=>p(130)(102),cout=>p(131)(103));
FA_ff_231:FAff port map(x=>p(3)(103),y=>p(4)(103),Cin=>p(5)(103),clock=>clock,reset=>reset,s=>p(130)(103),cout=>p(131)(104));
FA_ff_232:FAff port map(x=>p(3)(104),y=>p(4)(104),Cin=>p(5)(104),clock=>clock,reset=>reset,s=>p(130)(104),cout=>p(131)(105));
FA_ff_233:FAff port map(x=>p(3)(105),y=>p(4)(105),Cin=>p(5)(105),clock=>clock,reset=>reset,s=>p(130)(105),cout=>p(131)(106));
FA_ff_234:FAff port map(x=>p(3)(106),y=>p(4)(106),Cin=>p(5)(106),clock=>clock,reset=>reset,s=>p(130)(106),cout=>p(131)(107));
FA_ff_235:FAff port map(x=>p(3)(107),y=>p(4)(107),Cin=>p(5)(107),clock=>clock,reset=>reset,s=>p(130)(107),cout=>p(131)(108));
FA_ff_236:FAff port map(x=>p(3)(108),y=>p(4)(108),Cin=>p(5)(108),clock=>clock,reset=>reset,s=>p(130)(108),cout=>p(131)(109));
FA_ff_237:FAff port map(x=>p(3)(109),y=>p(4)(109),Cin=>p(5)(109),clock=>clock,reset=>reset,s=>p(130)(109),cout=>p(131)(110));
FA_ff_238:FAff port map(x=>p(3)(110),y=>p(4)(110),Cin=>p(5)(110),clock=>clock,reset=>reset,s=>p(130)(110),cout=>p(131)(111));
FA_ff_239:FAff port map(x=>p(3)(111),y=>p(4)(111),Cin=>p(5)(111),clock=>clock,reset=>reset,s=>p(130)(111),cout=>p(131)(112));
FA_ff_240:FAff port map(x=>p(3)(112),y=>p(4)(112),Cin=>p(5)(112),clock=>clock,reset=>reset,s=>p(130)(112),cout=>p(131)(113));
FA_ff_241:FAff port map(x=>p(3)(113),y=>p(4)(113),Cin=>p(5)(113),clock=>clock,reset=>reset,s=>p(130)(113),cout=>p(131)(114));
FA_ff_242:FAff port map(x=>p(3)(114),y=>p(4)(114),Cin=>p(5)(114),clock=>clock,reset=>reset,s=>p(130)(114),cout=>p(131)(115));
FA_ff_243:FAff port map(x=>p(3)(115),y=>p(4)(115),Cin=>p(5)(115),clock=>clock,reset=>reset,s=>p(130)(115),cout=>p(131)(116));
FA_ff_244:FAff port map(x=>p(3)(116),y=>p(4)(116),Cin=>p(5)(116),clock=>clock,reset=>reset,s=>p(130)(116),cout=>p(131)(117));
FA_ff_245:FAff port map(x=>p(3)(117),y=>p(4)(117),Cin=>p(5)(117),clock=>clock,reset=>reset,s=>p(130)(117),cout=>p(131)(118));
FA_ff_246:FAff port map(x=>p(3)(118),y=>p(4)(118),Cin=>p(5)(118),clock=>clock,reset=>reset,s=>p(130)(118),cout=>p(131)(119));
FA_ff_247:FAff port map(x=>p(3)(119),y=>p(4)(119),Cin=>p(5)(119),clock=>clock,reset=>reset,s=>p(130)(119),cout=>p(131)(120));
FA_ff_248:FAff port map(x=>p(3)(120),y=>p(4)(120),Cin=>p(5)(120),clock=>clock,reset=>reset,s=>p(130)(120),cout=>p(131)(121));
FA_ff_249:FAff port map(x=>p(3)(121),y=>p(4)(121),Cin=>p(5)(121),clock=>clock,reset=>reset,s=>p(130)(121),cout=>p(131)(122));
FA_ff_250:FAff port map(x=>p(3)(122),y=>p(4)(122),Cin=>p(5)(122),clock=>clock,reset=>reset,s=>p(130)(122),cout=>p(131)(123));
FA_ff_251:FAff port map(x=>p(3)(123),y=>p(4)(123),Cin=>p(5)(123),clock=>clock,reset=>reset,s=>p(130)(123),cout=>p(131)(124));
FA_ff_252:FAff port map(x=>p(3)(124),y=>p(4)(124),Cin=>p(5)(124),clock=>clock,reset=>reset,s=>p(130)(124),cout=>p(131)(125));
FA_ff_253:FAff port map(x=>p(3)(125),y=>p(4)(125),Cin=>p(5)(125),clock=>clock,reset=>reset,s=>p(130)(125),cout=>p(131)(126));
FA_ff_254:FAff port map(x=>p(3)(126),y=>p(4)(126),Cin=>p(5)(126),clock=>clock,reset=>reset,s=>p(130)(126),cout=>p(131)(127));
FA_ff_255:FAff port map(x=>p(3)(127),y=>p(4)(127),Cin=>p(5)(127),clock=>clock,reset=>reset,s=>p(130)(127),cout=>p(131)(128));
FA_ff_256:FAff port map(x=>p(6)(0),y=>p(7)(0),Cin=>p(8)(0),clock=>clock,reset=>reset,s=>p(132)(0),cout=>p(133)(1));
FA_ff_257:FAff port map(x=>p(6)(1),y=>p(7)(1),Cin=>p(8)(1),clock=>clock,reset=>reset,s=>p(132)(1),cout=>p(133)(2));
FA_ff_258:FAff port map(x=>p(6)(2),y=>p(7)(2),Cin=>p(8)(2),clock=>clock,reset=>reset,s=>p(132)(2),cout=>p(133)(3));
FA_ff_259:FAff port map(x=>p(6)(3),y=>p(7)(3),Cin=>p(8)(3),clock=>clock,reset=>reset,s=>p(132)(3),cout=>p(133)(4));
FA_ff_260:FAff port map(x=>p(6)(4),y=>p(7)(4),Cin=>p(8)(4),clock=>clock,reset=>reset,s=>p(132)(4),cout=>p(133)(5));
FA_ff_261:FAff port map(x=>p(6)(5),y=>p(7)(5),Cin=>p(8)(5),clock=>clock,reset=>reset,s=>p(132)(5),cout=>p(133)(6));
FA_ff_262:FAff port map(x=>p(6)(6),y=>p(7)(6),Cin=>p(8)(6),clock=>clock,reset=>reset,s=>p(132)(6),cout=>p(133)(7));
FA_ff_263:FAff port map(x=>p(6)(7),y=>p(7)(7),Cin=>p(8)(7),clock=>clock,reset=>reset,s=>p(132)(7),cout=>p(133)(8));
FA_ff_264:FAff port map(x=>p(6)(8),y=>p(7)(8),Cin=>p(8)(8),clock=>clock,reset=>reset,s=>p(132)(8),cout=>p(133)(9));
FA_ff_265:FAff port map(x=>p(6)(9),y=>p(7)(9),Cin=>p(8)(9),clock=>clock,reset=>reset,s=>p(132)(9),cout=>p(133)(10));
FA_ff_266:FAff port map(x=>p(6)(10),y=>p(7)(10),Cin=>p(8)(10),clock=>clock,reset=>reset,s=>p(132)(10),cout=>p(133)(11));
FA_ff_267:FAff port map(x=>p(6)(11),y=>p(7)(11),Cin=>p(8)(11),clock=>clock,reset=>reset,s=>p(132)(11),cout=>p(133)(12));
FA_ff_268:FAff port map(x=>p(6)(12),y=>p(7)(12),Cin=>p(8)(12),clock=>clock,reset=>reset,s=>p(132)(12),cout=>p(133)(13));
FA_ff_269:FAff port map(x=>p(6)(13),y=>p(7)(13),Cin=>p(8)(13),clock=>clock,reset=>reset,s=>p(132)(13),cout=>p(133)(14));
FA_ff_270:FAff port map(x=>p(6)(14),y=>p(7)(14),Cin=>p(8)(14),clock=>clock,reset=>reset,s=>p(132)(14),cout=>p(133)(15));
FA_ff_271:FAff port map(x=>p(6)(15),y=>p(7)(15),Cin=>p(8)(15),clock=>clock,reset=>reset,s=>p(132)(15),cout=>p(133)(16));
FA_ff_272:FAff port map(x=>p(6)(16),y=>p(7)(16),Cin=>p(8)(16),clock=>clock,reset=>reset,s=>p(132)(16),cout=>p(133)(17));
FA_ff_273:FAff port map(x=>p(6)(17),y=>p(7)(17),Cin=>p(8)(17),clock=>clock,reset=>reset,s=>p(132)(17),cout=>p(133)(18));
FA_ff_274:FAff port map(x=>p(6)(18),y=>p(7)(18),Cin=>p(8)(18),clock=>clock,reset=>reset,s=>p(132)(18),cout=>p(133)(19));
FA_ff_275:FAff port map(x=>p(6)(19),y=>p(7)(19),Cin=>p(8)(19),clock=>clock,reset=>reset,s=>p(132)(19),cout=>p(133)(20));
FA_ff_276:FAff port map(x=>p(6)(20),y=>p(7)(20),Cin=>p(8)(20),clock=>clock,reset=>reset,s=>p(132)(20),cout=>p(133)(21));
FA_ff_277:FAff port map(x=>p(6)(21),y=>p(7)(21),Cin=>p(8)(21),clock=>clock,reset=>reset,s=>p(132)(21),cout=>p(133)(22));
FA_ff_278:FAff port map(x=>p(6)(22),y=>p(7)(22),Cin=>p(8)(22),clock=>clock,reset=>reset,s=>p(132)(22),cout=>p(133)(23));
FA_ff_279:FAff port map(x=>p(6)(23),y=>p(7)(23),Cin=>p(8)(23),clock=>clock,reset=>reset,s=>p(132)(23),cout=>p(133)(24));
FA_ff_280:FAff port map(x=>p(6)(24),y=>p(7)(24),Cin=>p(8)(24),clock=>clock,reset=>reset,s=>p(132)(24),cout=>p(133)(25));
FA_ff_281:FAff port map(x=>p(6)(25),y=>p(7)(25),Cin=>p(8)(25),clock=>clock,reset=>reset,s=>p(132)(25),cout=>p(133)(26));
FA_ff_282:FAff port map(x=>p(6)(26),y=>p(7)(26),Cin=>p(8)(26),clock=>clock,reset=>reset,s=>p(132)(26),cout=>p(133)(27));
FA_ff_283:FAff port map(x=>p(6)(27),y=>p(7)(27),Cin=>p(8)(27),clock=>clock,reset=>reset,s=>p(132)(27),cout=>p(133)(28));
FA_ff_284:FAff port map(x=>p(6)(28),y=>p(7)(28),Cin=>p(8)(28),clock=>clock,reset=>reset,s=>p(132)(28),cout=>p(133)(29));
FA_ff_285:FAff port map(x=>p(6)(29),y=>p(7)(29),Cin=>p(8)(29),clock=>clock,reset=>reset,s=>p(132)(29),cout=>p(133)(30));
FA_ff_286:FAff port map(x=>p(6)(30),y=>p(7)(30),Cin=>p(8)(30),clock=>clock,reset=>reset,s=>p(132)(30),cout=>p(133)(31));
FA_ff_287:FAff port map(x=>p(6)(31),y=>p(7)(31),Cin=>p(8)(31),clock=>clock,reset=>reset,s=>p(132)(31),cout=>p(133)(32));
FA_ff_288:FAff port map(x=>p(6)(32),y=>p(7)(32),Cin=>p(8)(32),clock=>clock,reset=>reset,s=>p(132)(32),cout=>p(133)(33));
FA_ff_289:FAff port map(x=>p(6)(33),y=>p(7)(33),Cin=>p(8)(33),clock=>clock,reset=>reset,s=>p(132)(33),cout=>p(133)(34));
FA_ff_290:FAff port map(x=>p(6)(34),y=>p(7)(34),Cin=>p(8)(34),clock=>clock,reset=>reset,s=>p(132)(34),cout=>p(133)(35));
FA_ff_291:FAff port map(x=>p(6)(35),y=>p(7)(35),Cin=>p(8)(35),clock=>clock,reset=>reset,s=>p(132)(35),cout=>p(133)(36));
FA_ff_292:FAff port map(x=>p(6)(36),y=>p(7)(36),Cin=>p(8)(36),clock=>clock,reset=>reset,s=>p(132)(36),cout=>p(133)(37));
FA_ff_293:FAff port map(x=>p(6)(37),y=>p(7)(37),Cin=>p(8)(37),clock=>clock,reset=>reset,s=>p(132)(37),cout=>p(133)(38));
FA_ff_294:FAff port map(x=>p(6)(38),y=>p(7)(38),Cin=>p(8)(38),clock=>clock,reset=>reset,s=>p(132)(38),cout=>p(133)(39));
FA_ff_295:FAff port map(x=>p(6)(39),y=>p(7)(39),Cin=>p(8)(39),clock=>clock,reset=>reset,s=>p(132)(39),cout=>p(133)(40));
FA_ff_296:FAff port map(x=>p(6)(40),y=>p(7)(40),Cin=>p(8)(40),clock=>clock,reset=>reset,s=>p(132)(40),cout=>p(133)(41));
FA_ff_297:FAff port map(x=>p(6)(41),y=>p(7)(41),Cin=>p(8)(41),clock=>clock,reset=>reset,s=>p(132)(41),cout=>p(133)(42));
FA_ff_298:FAff port map(x=>p(6)(42),y=>p(7)(42),Cin=>p(8)(42),clock=>clock,reset=>reset,s=>p(132)(42),cout=>p(133)(43));
FA_ff_299:FAff port map(x=>p(6)(43),y=>p(7)(43),Cin=>p(8)(43),clock=>clock,reset=>reset,s=>p(132)(43),cout=>p(133)(44));
FA_ff_300:FAff port map(x=>p(6)(44),y=>p(7)(44),Cin=>p(8)(44),clock=>clock,reset=>reset,s=>p(132)(44),cout=>p(133)(45));
FA_ff_301:FAff port map(x=>p(6)(45),y=>p(7)(45),Cin=>p(8)(45),clock=>clock,reset=>reset,s=>p(132)(45),cout=>p(133)(46));
FA_ff_302:FAff port map(x=>p(6)(46),y=>p(7)(46),Cin=>p(8)(46),clock=>clock,reset=>reset,s=>p(132)(46),cout=>p(133)(47));
FA_ff_303:FAff port map(x=>p(6)(47),y=>p(7)(47),Cin=>p(8)(47),clock=>clock,reset=>reset,s=>p(132)(47),cout=>p(133)(48));
FA_ff_304:FAff port map(x=>p(6)(48),y=>p(7)(48),Cin=>p(8)(48),clock=>clock,reset=>reset,s=>p(132)(48),cout=>p(133)(49));
FA_ff_305:FAff port map(x=>p(6)(49),y=>p(7)(49),Cin=>p(8)(49),clock=>clock,reset=>reset,s=>p(132)(49),cout=>p(133)(50));
FA_ff_306:FAff port map(x=>p(6)(50),y=>p(7)(50),Cin=>p(8)(50),clock=>clock,reset=>reset,s=>p(132)(50),cout=>p(133)(51));
FA_ff_307:FAff port map(x=>p(6)(51),y=>p(7)(51),Cin=>p(8)(51),clock=>clock,reset=>reset,s=>p(132)(51),cout=>p(133)(52));
FA_ff_308:FAff port map(x=>p(6)(52),y=>p(7)(52),Cin=>p(8)(52),clock=>clock,reset=>reset,s=>p(132)(52),cout=>p(133)(53));
FA_ff_309:FAff port map(x=>p(6)(53),y=>p(7)(53),Cin=>p(8)(53),clock=>clock,reset=>reset,s=>p(132)(53),cout=>p(133)(54));
FA_ff_310:FAff port map(x=>p(6)(54),y=>p(7)(54),Cin=>p(8)(54),clock=>clock,reset=>reset,s=>p(132)(54),cout=>p(133)(55));
FA_ff_311:FAff port map(x=>p(6)(55),y=>p(7)(55),Cin=>p(8)(55),clock=>clock,reset=>reset,s=>p(132)(55),cout=>p(133)(56));
FA_ff_312:FAff port map(x=>p(6)(56),y=>p(7)(56),Cin=>p(8)(56),clock=>clock,reset=>reset,s=>p(132)(56),cout=>p(133)(57));
FA_ff_313:FAff port map(x=>p(6)(57),y=>p(7)(57),Cin=>p(8)(57),clock=>clock,reset=>reset,s=>p(132)(57),cout=>p(133)(58));
FA_ff_314:FAff port map(x=>p(6)(58),y=>p(7)(58),Cin=>p(8)(58),clock=>clock,reset=>reset,s=>p(132)(58),cout=>p(133)(59));
FA_ff_315:FAff port map(x=>p(6)(59),y=>p(7)(59),Cin=>p(8)(59),clock=>clock,reset=>reset,s=>p(132)(59),cout=>p(133)(60));
FA_ff_316:FAff port map(x=>p(6)(60),y=>p(7)(60),Cin=>p(8)(60),clock=>clock,reset=>reset,s=>p(132)(60),cout=>p(133)(61));
FA_ff_317:FAff port map(x=>p(6)(61),y=>p(7)(61),Cin=>p(8)(61),clock=>clock,reset=>reset,s=>p(132)(61),cout=>p(133)(62));
FA_ff_318:FAff port map(x=>p(6)(62),y=>p(7)(62),Cin=>p(8)(62),clock=>clock,reset=>reset,s=>p(132)(62),cout=>p(133)(63));
FA_ff_319:FAff port map(x=>p(6)(63),y=>p(7)(63),Cin=>p(8)(63),clock=>clock,reset=>reset,s=>p(132)(63),cout=>p(133)(64));
FA_ff_320:FAff port map(x=>p(6)(64),y=>p(7)(64),Cin=>p(8)(64),clock=>clock,reset=>reset,s=>p(132)(64),cout=>p(133)(65));
FA_ff_321:FAff port map(x=>p(6)(65),y=>p(7)(65),Cin=>p(8)(65),clock=>clock,reset=>reset,s=>p(132)(65),cout=>p(133)(66));
FA_ff_322:FAff port map(x=>p(6)(66),y=>p(7)(66),Cin=>p(8)(66),clock=>clock,reset=>reset,s=>p(132)(66),cout=>p(133)(67));
FA_ff_323:FAff port map(x=>p(6)(67),y=>p(7)(67),Cin=>p(8)(67),clock=>clock,reset=>reset,s=>p(132)(67),cout=>p(133)(68));
FA_ff_324:FAff port map(x=>p(6)(68),y=>p(7)(68),Cin=>p(8)(68),clock=>clock,reset=>reset,s=>p(132)(68),cout=>p(133)(69));
FA_ff_325:FAff port map(x=>p(6)(69),y=>p(7)(69),Cin=>p(8)(69),clock=>clock,reset=>reset,s=>p(132)(69),cout=>p(133)(70));
FA_ff_326:FAff port map(x=>p(6)(70),y=>p(7)(70),Cin=>p(8)(70),clock=>clock,reset=>reset,s=>p(132)(70),cout=>p(133)(71));
FA_ff_327:FAff port map(x=>p(6)(71),y=>p(7)(71),Cin=>p(8)(71),clock=>clock,reset=>reset,s=>p(132)(71),cout=>p(133)(72));
FA_ff_328:FAff port map(x=>p(6)(72),y=>p(7)(72),Cin=>p(8)(72),clock=>clock,reset=>reset,s=>p(132)(72),cout=>p(133)(73));
FA_ff_329:FAff port map(x=>p(6)(73),y=>p(7)(73),Cin=>p(8)(73),clock=>clock,reset=>reset,s=>p(132)(73),cout=>p(133)(74));
FA_ff_330:FAff port map(x=>p(6)(74),y=>p(7)(74),Cin=>p(8)(74),clock=>clock,reset=>reset,s=>p(132)(74),cout=>p(133)(75));
FA_ff_331:FAff port map(x=>p(6)(75),y=>p(7)(75),Cin=>p(8)(75),clock=>clock,reset=>reset,s=>p(132)(75),cout=>p(133)(76));
FA_ff_332:FAff port map(x=>p(6)(76),y=>p(7)(76),Cin=>p(8)(76),clock=>clock,reset=>reset,s=>p(132)(76),cout=>p(133)(77));
FA_ff_333:FAff port map(x=>p(6)(77),y=>p(7)(77),Cin=>p(8)(77),clock=>clock,reset=>reset,s=>p(132)(77),cout=>p(133)(78));
FA_ff_334:FAff port map(x=>p(6)(78),y=>p(7)(78),Cin=>p(8)(78),clock=>clock,reset=>reset,s=>p(132)(78),cout=>p(133)(79));
FA_ff_335:FAff port map(x=>p(6)(79),y=>p(7)(79),Cin=>p(8)(79),clock=>clock,reset=>reset,s=>p(132)(79),cout=>p(133)(80));
FA_ff_336:FAff port map(x=>p(6)(80),y=>p(7)(80),Cin=>p(8)(80),clock=>clock,reset=>reset,s=>p(132)(80),cout=>p(133)(81));
FA_ff_337:FAff port map(x=>p(6)(81),y=>p(7)(81),Cin=>p(8)(81),clock=>clock,reset=>reset,s=>p(132)(81),cout=>p(133)(82));
FA_ff_338:FAff port map(x=>p(6)(82),y=>p(7)(82),Cin=>p(8)(82),clock=>clock,reset=>reset,s=>p(132)(82),cout=>p(133)(83));
FA_ff_339:FAff port map(x=>p(6)(83),y=>p(7)(83),Cin=>p(8)(83),clock=>clock,reset=>reset,s=>p(132)(83),cout=>p(133)(84));
FA_ff_340:FAff port map(x=>p(6)(84),y=>p(7)(84),Cin=>p(8)(84),clock=>clock,reset=>reset,s=>p(132)(84),cout=>p(133)(85));
FA_ff_341:FAff port map(x=>p(6)(85),y=>p(7)(85),Cin=>p(8)(85),clock=>clock,reset=>reset,s=>p(132)(85),cout=>p(133)(86));
FA_ff_342:FAff port map(x=>p(6)(86),y=>p(7)(86),Cin=>p(8)(86),clock=>clock,reset=>reset,s=>p(132)(86),cout=>p(133)(87));
FA_ff_343:FAff port map(x=>p(6)(87),y=>p(7)(87),Cin=>p(8)(87),clock=>clock,reset=>reset,s=>p(132)(87),cout=>p(133)(88));
FA_ff_344:FAff port map(x=>p(6)(88),y=>p(7)(88),Cin=>p(8)(88),clock=>clock,reset=>reset,s=>p(132)(88),cout=>p(133)(89));
FA_ff_345:FAff port map(x=>p(6)(89),y=>p(7)(89),Cin=>p(8)(89),clock=>clock,reset=>reset,s=>p(132)(89),cout=>p(133)(90));
FA_ff_346:FAff port map(x=>p(6)(90),y=>p(7)(90),Cin=>p(8)(90),clock=>clock,reset=>reset,s=>p(132)(90),cout=>p(133)(91));
FA_ff_347:FAff port map(x=>p(6)(91),y=>p(7)(91),Cin=>p(8)(91),clock=>clock,reset=>reset,s=>p(132)(91),cout=>p(133)(92));
FA_ff_348:FAff port map(x=>p(6)(92),y=>p(7)(92),Cin=>p(8)(92),clock=>clock,reset=>reset,s=>p(132)(92),cout=>p(133)(93));
FA_ff_349:FAff port map(x=>p(6)(93),y=>p(7)(93),Cin=>p(8)(93),clock=>clock,reset=>reset,s=>p(132)(93),cout=>p(133)(94));
FA_ff_350:FAff port map(x=>p(6)(94),y=>p(7)(94),Cin=>p(8)(94),clock=>clock,reset=>reset,s=>p(132)(94),cout=>p(133)(95));
FA_ff_351:FAff port map(x=>p(6)(95),y=>p(7)(95),Cin=>p(8)(95),clock=>clock,reset=>reset,s=>p(132)(95),cout=>p(133)(96));
FA_ff_352:FAff port map(x=>p(6)(96),y=>p(7)(96),Cin=>p(8)(96),clock=>clock,reset=>reset,s=>p(132)(96),cout=>p(133)(97));
FA_ff_353:FAff port map(x=>p(6)(97),y=>p(7)(97),Cin=>p(8)(97),clock=>clock,reset=>reset,s=>p(132)(97),cout=>p(133)(98));
FA_ff_354:FAff port map(x=>p(6)(98),y=>p(7)(98),Cin=>p(8)(98),clock=>clock,reset=>reset,s=>p(132)(98),cout=>p(133)(99));
FA_ff_355:FAff port map(x=>p(6)(99),y=>p(7)(99),Cin=>p(8)(99),clock=>clock,reset=>reset,s=>p(132)(99),cout=>p(133)(100));
FA_ff_356:FAff port map(x=>p(6)(100),y=>p(7)(100),Cin=>p(8)(100),clock=>clock,reset=>reset,s=>p(132)(100),cout=>p(133)(101));
FA_ff_357:FAff port map(x=>p(6)(101),y=>p(7)(101),Cin=>p(8)(101),clock=>clock,reset=>reset,s=>p(132)(101),cout=>p(133)(102));
FA_ff_358:FAff port map(x=>p(6)(102),y=>p(7)(102),Cin=>p(8)(102),clock=>clock,reset=>reset,s=>p(132)(102),cout=>p(133)(103));
FA_ff_359:FAff port map(x=>p(6)(103),y=>p(7)(103),Cin=>p(8)(103),clock=>clock,reset=>reset,s=>p(132)(103),cout=>p(133)(104));
FA_ff_360:FAff port map(x=>p(6)(104),y=>p(7)(104),Cin=>p(8)(104),clock=>clock,reset=>reset,s=>p(132)(104),cout=>p(133)(105));
FA_ff_361:FAff port map(x=>p(6)(105),y=>p(7)(105),Cin=>p(8)(105),clock=>clock,reset=>reset,s=>p(132)(105),cout=>p(133)(106));
FA_ff_362:FAff port map(x=>p(6)(106),y=>p(7)(106),Cin=>p(8)(106),clock=>clock,reset=>reset,s=>p(132)(106),cout=>p(133)(107));
FA_ff_363:FAff port map(x=>p(6)(107),y=>p(7)(107),Cin=>p(8)(107),clock=>clock,reset=>reset,s=>p(132)(107),cout=>p(133)(108));
FA_ff_364:FAff port map(x=>p(6)(108),y=>p(7)(108),Cin=>p(8)(108),clock=>clock,reset=>reset,s=>p(132)(108),cout=>p(133)(109));
FA_ff_365:FAff port map(x=>p(6)(109),y=>p(7)(109),Cin=>p(8)(109),clock=>clock,reset=>reset,s=>p(132)(109),cout=>p(133)(110));
FA_ff_366:FAff port map(x=>p(6)(110),y=>p(7)(110),Cin=>p(8)(110),clock=>clock,reset=>reset,s=>p(132)(110),cout=>p(133)(111));
FA_ff_367:FAff port map(x=>p(6)(111),y=>p(7)(111),Cin=>p(8)(111),clock=>clock,reset=>reset,s=>p(132)(111),cout=>p(133)(112));
FA_ff_368:FAff port map(x=>p(6)(112),y=>p(7)(112),Cin=>p(8)(112),clock=>clock,reset=>reset,s=>p(132)(112),cout=>p(133)(113));
FA_ff_369:FAff port map(x=>p(6)(113),y=>p(7)(113),Cin=>p(8)(113),clock=>clock,reset=>reset,s=>p(132)(113),cout=>p(133)(114));
FA_ff_370:FAff port map(x=>p(6)(114),y=>p(7)(114),Cin=>p(8)(114),clock=>clock,reset=>reset,s=>p(132)(114),cout=>p(133)(115));
FA_ff_371:FAff port map(x=>p(6)(115),y=>p(7)(115),Cin=>p(8)(115),clock=>clock,reset=>reset,s=>p(132)(115),cout=>p(133)(116));
FA_ff_372:FAff port map(x=>p(6)(116),y=>p(7)(116),Cin=>p(8)(116),clock=>clock,reset=>reset,s=>p(132)(116),cout=>p(133)(117));
FA_ff_373:FAff port map(x=>p(6)(117),y=>p(7)(117),Cin=>p(8)(117),clock=>clock,reset=>reset,s=>p(132)(117),cout=>p(133)(118));
FA_ff_374:FAff port map(x=>p(6)(118),y=>p(7)(118),Cin=>p(8)(118),clock=>clock,reset=>reset,s=>p(132)(118),cout=>p(133)(119));
FA_ff_375:FAff port map(x=>p(6)(119),y=>p(7)(119),Cin=>p(8)(119),clock=>clock,reset=>reset,s=>p(132)(119),cout=>p(133)(120));
FA_ff_376:FAff port map(x=>p(6)(120),y=>p(7)(120),Cin=>p(8)(120),clock=>clock,reset=>reset,s=>p(132)(120),cout=>p(133)(121));
FA_ff_377:FAff port map(x=>p(6)(121),y=>p(7)(121),Cin=>p(8)(121),clock=>clock,reset=>reset,s=>p(132)(121),cout=>p(133)(122));
FA_ff_378:FAff port map(x=>p(6)(122),y=>p(7)(122),Cin=>p(8)(122),clock=>clock,reset=>reset,s=>p(132)(122),cout=>p(133)(123));
FA_ff_379:FAff port map(x=>p(6)(123),y=>p(7)(123),Cin=>p(8)(123),clock=>clock,reset=>reset,s=>p(132)(123),cout=>p(133)(124));
FA_ff_380:FAff port map(x=>p(6)(124),y=>p(7)(124),Cin=>p(8)(124),clock=>clock,reset=>reset,s=>p(132)(124),cout=>p(133)(125));
FA_ff_381:FAff port map(x=>p(6)(125),y=>p(7)(125),Cin=>p(8)(125),clock=>clock,reset=>reset,s=>p(132)(125),cout=>p(133)(126));
FA_ff_382:FAff port map(x=>p(6)(126),y=>p(7)(126),Cin=>p(8)(126),clock=>clock,reset=>reset,s=>p(132)(126),cout=>p(133)(127));
FA_ff_383:FAff port map(x=>p(6)(127),y=>p(7)(127),Cin=>p(8)(127),clock=>clock,reset=>reset,s=>p(132)(127),cout=>p(133)(128));
FA_ff_384:FAff port map(x=>p(9)(0),y=>p(10)(0),Cin=>p(11)(0),clock=>clock,reset=>reset,s=>p(134)(0),cout=>p(135)(1));
FA_ff_385:FAff port map(x=>p(9)(1),y=>p(10)(1),Cin=>p(11)(1),clock=>clock,reset=>reset,s=>p(134)(1),cout=>p(135)(2));
FA_ff_386:FAff port map(x=>p(9)(2),y=>p(10)(2),Cin=>p(11)(2),clock=>clock,reset=>reset,s=>p(134)(2),cout=>p(135)(3));
FA_ff_387:FAff port map(x=>p(9)(3),y=>p(10)(3),Cin=>p(11)(3),clock=>clock,reset=>reset,s=>p(134)(3),cout=>p(135)(4));
FA_ff_388:FAff port map(x=>p(9)(4),y=>p(10)(4),Cin=>p(11)(4),clock=>clock,reset=>reset,s=>p(134)(4),cout=>p(135)(5));
FA_ff_389:FAff port map(x=>p(9)(5),y=>p(10)(5),Cin=>p(11)(5),clock=>clock,reset=>reset,s=>p(134)(5),cout=>p(135)(6));
FA_ff_390:FAff port map(x=>p(9)(6),y=>p(10)(6),Cin=>p(11)(6),clock=>clock,reset=>reset,s=>p(134)(6),cout=>p(135)(7));
FA_ff_391:FAff port map(x=>p(9)(7),y=>p(10)(7),Cin=>p(11)(7),clock=>clock,reset=>reset,s=>p(134)(7),cout=>p(135)(8));
FA_ff_392:FAff port map(x=>p(9)(8),y=>p(10)(8),Cin=>p(11)(8),clock=>clock,reset=>reset,s=>p(134)(8),cout=>p(135)(9));
FA_ff_393:FAff port map(x=>p(9)(9),y=>p(10)(9),Cin=>p(11)(9),clock=>clock,reset=>reset,s=>p(134)(9),cout=>p(135)(10));
FA_ff_394:FAff port map(x=>p(9)(10),y=>p(10)(10),Cin=>p(11)(10),clock=>clock,reset=>reset,s=>p(134)(10),cout=>p(135)(11));
FA_ff_395:FAff port map(x=>p(9)(11),y=>p(10)(11),Cin=>p(11)(11),clock=>clock,reset=>reset,s=>p(134)(11),cout=>p(135)(12));
FA_ff_396:FAff port map(x=>p(9)(12),y=>p(10)(12),Cin=>p(11)(12),clock=>clock,reset=>reset,s=>p(134)(12),cout=>p(135)(13));
FA_ff_397:FAff port map(x=>p(9)(13),y=>p(10)(13),Cin=>p(11)(13),clock=>clock,reset=>reset,s=>p(134)(13),cout=>p(135)(14));
FA_ff_398:FAff port map(x=>p(9)(14),y=>p(10)(14),Cin=>p(11)(14),clock=>clock,reset=>reset,s=>p(134)(14),cout=>p(135)(15));
FA_ff_399:FAff port map(x=>p(9)(15),y=>p(10)(15),Cin=>p(11)(15),clock=>clock,reset=>reset,s=>p(134)(15),cout=>p(135)(16));
FA_ff_400:FAff port map(x=>p(9)(16),y=>p(10)(16),Cin=>p(11)(16),clock=>clock,reset=>reset,s=>p(134)(16),cout=>p(135)(17));
FA_ff_401:FAff port map(x=>p(9)(17),y=>p(10)(17),Cin=>p(11)(17),clock=>clock,reset=>reset,s=>p(134)(17),cout=>p(135)(18));
FA_ff_402:FAff port map(x=>p(9)(18),y=>p(10)(18),Cin=>p(11)(18),clock=>clock,reset=>reset,s=>p(134)(18),cout=>p(135)(19));
FA_ff_403:FAff port map(x=>p(9)(19),y=>p(10)(19),Cin=>p(11)(19),clock=>clock,reset=>reset,s=>p(134)(19),cout=>p(135)(20));
FA_ff_404:FAff port map(x=>p(9)(20),y=>p(10)(20),Cin=>p(11)(20),clock=>clock,reset=>reset,s=>p(134)(20),cout=>p(135)(21));
FA_ff_405:FAff port map(x=>p(9)(21),y=>p(10)(21),Cin=>p(11)(21),clock=>clock,reset=>reset,s=>p(134)(21),cout=>p(135)(22));
FA_ff_406:FAff port map(x=>p(9)(22),y=>p(10)(22),Cin=>p(11)(22),clock=>clock,reset=>reset,s=>p(134)(22),cout=>p(135)(23));
FA_ff_407:FAff port map(x=>p(9)(23),y=>p(10)(23),Cin=>p(11)(23),clock=>clock,reset=>reset,s=>p(134)(23),cout=>p(135)(24));
FA_ff_408:FAff port map(x=>p(9)(24),y=>p(10)(24),Cin=>p(11)(24),clock=>clock,reset=>reset,s=>p(134)(24),cout=>p(135)(25));
FA_ff_409:FAff port map(x=>p(9)(25),y=>p(10)(25),Cin=>p(11)(25),clock=>clock,reset=>reset,s=>p(134)(25),cout=>p(135)(26));
FA_ff_410:FAff port map(x=>p(9)(26),y=>p(10)(26),Cin=>p(11)(26),clock=>clock,reset=>reset,s=>p(134)(26),cout=>p(135)(27));
FA_ff_411:FAff port map(x=>p(9)(27),y=>p(10)(27),Cin=>p(11)(27),clock=>clock,reset=>reset,s=>p(134)(27),cout=>p(135)(28));
FA_ff_412:FAff port map(x=>p(9)(28),y=>p(10)(28),Cin=>p(11)(28),clock=>clock,reset=>reset,s=>p(134)(28),cout=>p(135)(29));
FA_ff_413:FAff port map(x=>p(9)(29),y=>p(10)(29),Cin=>p(11)(29),clock=>clock,reset=>reset,s=>p(134)(29),cout=>p(135)(30));
FA_ff_414:FAff port map(x=>p(9)(30),y=>p(10)(30),Cin=>p(11)(30),clock=>clock,reset=>reset,s=>p(134)(30),cout=>p(135)(31));
FA_ff_415:FAff port map(x=>p(9)(31),y=>p(10)(31),Cin=>p(11)(31),clock=>clock,reset=>reset,s=>p(134)(31),cout=>p(135)(32));
FA_ff_416:FAff port map(x=>p(9)(32),y=>p(10)(32),Cin=>p(11)(32),clock=>clock,reset=>reset,s=>p(134)(32),cout=>p(135)(33));
FA_ff_417:FAff port map(x=>p(9)(33),y=>p(10)(33),Cin=>p(11)(33),clock=>clock,reset=>reset,s=>p(134)(33),cout=>p(135)(34));
FA_ff_418:FAff port map(x=>p(9)(34),y=>p(10)(34),Cin=>p(11)(34),clock=>clock,reset=>reset,s=>p(134)(34),cout=>p(135)(35));
FA_ff_419:FAff port map(x=>p(9)(35),y=>p(10)(35),Cin=>p(11)(35),clock=>clock,reset=>reset,s=>p(134)(35),cout=>p(135)(36));
FA_ff_420:FAff port map(x=>p(9)(36),y=>p(10)(36),Cin=>p(11)(36),clock=>clock,reset=>reset,s=>p(134)(36),cout=>p(135)(37));
FA_ff_421:FAff port map(x=>p(9)(37),y=>p(10)(37),Cin=>p(11)(37),clock=>clock,reset=>reset,s=>p(134)(37),cout=>p(135)(38));
FA_ff_422:FAff port map(x=>p(9)(38),y=>p(10)(38),Cin=>p(11)(38),clock=>clock,reset=>reset,s=>p(134)(38),cout=>p(135)(39));
FA_ff_423:FAff port map(x=>p(9)(39),y=>p(10)(39),Cin=>p(11)(39),clock=>clock,reset=>reset,s=>p(134)(39),cout=>p(135)(40));
FA_ff_424:FAff port map(x=>p(9)(40),y=>p(10)(40),Cin=>p(11)(40),clock=>clock,reset=>reset,s=>p(134)(40),cout=>p(135)(41));
FA_ff_425:FAff port map(x=>p(9)(41),y=>p(10)(41),Cin=>p(11)(41),clock=>clock,reset=>reset,s=>p(134)(41),cout=>p(135)(42));
FA_ff_426:FAff port map(x=>p(9)(42),y=>p(10)(42),Cin=>p(11)(42),clock=>clock,reset=>reset,s=>p(134)(42),cout=>p(135)(43));
FA_ff_427:FAff port map(x=>p(9)(43),y=>p(10)(43),Cin=>p(11)(43),clock=>clock,reset=>reset,s=>p(134)(43),cout=>p(135)(44));
FA_ff_428:FAff port map(x=>p(9)(44),y=>p(10)(44),Cin=>p(11)(44),clock=>clock,reset=>reset,s=>p(134)(44),cout=>p(135)(45));
FA_ff_429:FAff port map(x=>p(9)(45),y=>p(10)(45),Cin=>p(11)(45),clock=>clock,reset=>reset,s=>p(134)(45),cout=>p(135)(46));
FA_ff_430:FAff port map(x=>p(9)(46),y=>p(10)(46),Cin=>p(11)(46),clock=>clock,reset=>reset,s=>p(134)(46),cout=>p(135)(47));
FA_ff_431:FAff port map(x=>p(9)(47),y=>p(10)(47),Cin=>p(11)(47),clock=>clock,reset=>reset,s=>p(134)(47),cout=>p(135)(48));
FA_ff_432:FAff port map(x=>p(9)(48),y=>p(10)(48),Cin=>p(11)(48),clock=>clock,reset=>reset,s=>p(134)(48),cout=>p(135)(49));
FA_ff_433:FAff port map(x=>p(9)(49),y=>p(10)(49),Cin=>p(11)(49),clock=>clock,reset=>reset,s=>p(134)(49),cout=>p(135)(50));
FA_ff_434:FAff port map(x=>p(9)(50),y=>p(10)(50),Cin=>p(11)(50),clock=>clock,reset=>reset,s=>p(134)(50),cout=>p(135)(51));
FA_ff_435:FAff port map(x=>p(9)(51),y=>p(10)(51),Cin=>p(11)(51),clock=>clock,reset=>reset,s=>p(134)(51),cout=>p(135)(52));
FA_ff_436:FAff port map(x=>p(9)(52),y=>p(10)(52),Cin=>p(11)(52),clock=>clock,reset=>reset,s=>p(134)(52),cout=>p(135)(53));
FA_ff_437:FAff port map(x=>p(9)(53),y=>p(10)(53),Cin=>p(11)(53),clock=>clock,reset=>reset,s=>p(134)(53),cout=>p(135)(54));
FA_ff_438:FAff port map(x=>p(9)(54),y=>p(10)(54),Cin=>p(11)(54),clock=>clock,reset=>reset,s=>p(134)(54),cout=>p(135)(55));
FA_ff_439:FAff port map(x=>p(9)(55),y=>p(10)(55),Cin=>p(11)(55),clock=>clock,reset=>reset,s=>p(134)(55),cout=>p(135)(56));
FA_ff_440:FAff port map(x=>p(9)(56),y=>p(10)(56),Cin=>p(11)(56),clock=>clock,reset=>reset,s=>p(134)(56),cout=>p(135)(57));
FA_ff_441:FAff port map(x=>p(9)(57),y=>p(10)(57),Cin=>p(11)(57),clock=>clock,reset=>reset,s=>p(134)(57),cout=>p(135)(58));
FA_ff_442:FAff port map(x=>p(9)(58),y=>p(10)(58),Cin=>p(11)(58),clock=>clock,reset=>reset,s=>p(134)(58),cout=>p(135)(59));
FA_ff_443:FAff port map(x=>p(9)(59),y=>p(10)(59),Cin=>p(11)(59),clock=>clock,reset=>reset,s=>p(134)(59),cout=>p(135)(60));
FA_ff_444:FAff port map(x=>p(9)(60),y=>p(10)(60),Cin=>p(11)(60),clock=>clock,reset=>reset,s=>p(134)(60),cout=>p(135)(61));
FA_ff_445:FAff port map(x=>p(9)(61),y=>p(10)(61),Cin=>p(11)(61),clock=>clock,reset=>reset,s=>p(134)(61),cout=>p(135)(62));
FA_ff_446:FAff port map(x=>p(9)(62),y=>p(10)(62),Cin=>p(11)(62),clock=>clock,reset=>reset,s=>p(134)(62),cout=>p(135)(63));
FA_ff_447:FAff port map(x=>p(9)(63),y=>p(10)(63),Cin=>p(11)(63),clock=>clock,reset=>reset,s=>p(134)(63),cout=>p(135)(64));
FA_ff_448:FAff port map(x=>p(9)(64),y=>p(10)(64),Cin=>p(11)(64),clock=>clock,reset=>reset,s=>p(134)(64),cout=>p(135)(65));
FA_ff_449:FAff port map(x=>p(9)(65),y=>p(10)(65),Cin=>p(11)(65),clock=>clock,reset=>reset,s=>p(134)(65),cout=>p(135)(66));
FA_ff_450:FAff port map(x=>p(9)(66),y=>p(10)(66),Cin=>p(11)(66),clock=>clock,reset=>reset,s=>p(134)(66),cout=>p(135)(67));
FA_ff_451:FAff port map(x=>p(9)(67),y=>p(10)(67),Cin=>p(11)(67),clock=>clock,reset=>reset,s=>p(134)(67),cout=>p(135)(68));
FA_ff_452:FAff port map(x=>p(9)(68),y=>p(10)(68),Cin=>p(11)(68),clock=>clock,reset=>reset,s=>p(134)(68),cout=>p(135)(69));
FA_ff_453:FAff port map(x=>p(9)(69),y=>p(10)(69),Cin=>p(11)(69),clock=>clock,reset=>reset,s=>p(134)(69),cout=>p(135)(70));
FA_ff_454:FAff port map(x=>p(9)(70),y=>p(10)(70),Cin=>p(11)(70),clock=>clock,reset=>reset,s=>p(134)(70),cout=>p(135)(71));
FA_ff_455:FAff port map(x=>p(9)(71),y=>p(10)(71),Cin=>p(11)(71),clock=>clock,reset=>reset,s=>p(134)(71),cout=>p(135)(72));
FA_ff_456:FAff port map(x=>p(9)(72),y=>p(10)(72),Cin=>p(11)(72),clock=>clock,reset=>reset,s=>p(134)(72),cout=>p(135)(73));
FA_ff_457:FAff port map(x=>p(9)(73),y=>p(10)(73),Cin=>p(11)(73),clock=>clock,reset=>reset,s=>p(134)(73),cout=>p(135)(74));
FA_ff_458:FAff port map(x=>p(9)(74),y=>p(10)(74),Cin=>p(11)(74),clock=>clock,reset=>reset,s=>p(134)(74),cout=>p(135)(75));
FA_ff_459:FAff port map(x=>p(9)(75),y=>p(10)(75),Cin=>p(11)(75),clock=>clock,reset=>reset,s=>p(134)(75),cout=>p(135)(76));
FA_ff_460:FAff port map(x=>p(9)(76),y=>p(10)(76),Cin=>p(11)(76),clock=>clock,reset=>reset,s=>p(134)(76),cout=>p(135)(77));
FA_ff_461:FAff port map(x=>p(9)(77),y=>p(10)(77),Cin=>p(11)(77),clock=>clock,reset=>reset,s=>p(134)(77),cout=>p(135)(78));
FA_ff_462:FAff port map(x=>p(9)(78),y=>p(10)(78),Cin=>p(11)(78),clock=>clock,reset=>reset,s=>p(134)(78),cout=>p(135)(79));
FA_ff_463:FAff port map(x=>p(9)(79),y=>p(10)(79),Cin=>p(11)(79),clock=>clock,reset=>reset,s=>p(134)(79),cout=>p(135)(80));
FA_ff_464:FAff port map(x=>p(9)(80),y=>p(10)(80),Cin=>p(11)(80),clock=>clock,reset=>reset,s=>p(134)(80),cout=>p(135)(81));
FA_ff_465:FAff port map(x=>p(9)(81),y=>p(10)(81),Cin=>p(11)(81),clock=>clock,reset=>reset,s=>p(134)(81),cout=>p(135)(82));
FA_ff_466:FAff port map(x=>p(9)(82),y=>p(10)(82),Cin=>p(11)(82),clock=>clock,reset=>reset,s=>p(134)(82),cout=>p(135)(83));
FA_ff_467:FAff port map(x=>p(9)(83),y=>p(10)(83),Cin=>p(11)(83),clock=>clock,reset=>reset,s=>p(134)(83),cout=>p(135)(84));
FA_ff_468:FAff port map(x=>p(9)(84),y=>p(10)(84),Cin=>p(11)(84),clock=>clock,reset=>reset,s=>p(134)(84),cout=>p(135)(85));
FA_ff_469:FAff port map(x=>p(9)(85),y=>p(10)(85),Cin=>p(11)(85),clock=>clock,reset=>reset,s=>p(134)(85),cout=>p(135)(86));
FA_ff_470:FAff port map(x=>p(9)(86),y=>p(10)(86),Cin=>p(11)(86),clock=>clock,reset=>reset,s=>p(134)(86),cout=>p(135)(87));
FA_ff_471:FAff port map(x=>p(9)(87),y=>p(10)(87),Cin=>p(11)(87),clock=>clock,reset=>reset,s=>p(134)(87),cout=>p(135)(88));
FA_ff_472:FAff port map(x=>p(9)(88),y=>p(10)(88),Cin=>p(11)(88),clock=>clock,reset=>reset,s=>p(134)(88),cout=>p(135)(89));
FA_ff_473:FAff port map(x=>p(9)(89),y=>p(10)(89),Cin=>p(11)(89),clock=>clock,reset=>reset,s=>p(134)(89),cout=>p(135)(90));
FA_ff_474:FAff port map(x=>p(9)(90),y=>p(10)(90),Cin=>p(11)(90),clock=>clock,reset=>reset,s=>p(134)(90),cout=>p(135)(91));
FA_ff_475:FAff port map(x=>p(9)(91),y=>p(10)(91),Cin=>p(11)(91),clock=>clock,reset=>reset,s=>p(134)(91),cout=>p(135)(92));
FA_ff_476:FAff port map(x=>p(9)(92),y=>p(10)(92),Cin=>p(11)(92),clock=>clock,reset=>reset,s=>p(134)(92),cout=>p(135)(93));
FA_ff_477:FAff port map(x=>p(9)(93),y=>p(10)(93),Cin=>p(11)(93),clock=>clock,reset=>reset,s=>p(134)(93),cout=>p(135)(94));
FA_ff_478:FAff port map(x=>p(9)(94),y=>p(10)(94),Cin=>p(11)(94),clock=>clock,reset=>reset,s=>p(134)(94),cout=>p(135)(95));
FA_ff_479:FAff port map(x=>p(9)(95),y=>p(10)(95),Cin=>p(11)(95),clock=>clock,reset=>reset,s=>p(134)(95),cout=>p(135)(96));
FA_ff_480:FAff port map(x=>p(9)(96),y=>p(10)(96),Cin=>p(11)(96),clock=>clock,reset=>reset,s=>p(134)(96),cout=>p(135)(97));
FA_ff_481:FAff port map(x=>p(9)(97),y=>p(10)(97),Cin=>p(11)(97),clock=>clock,reset=>reset,s=>p(134)(97),cout=>p(135)(98));
FA_ff_482:FAff port map(x=>p(9)(98),y=>p(10)(98),Cin=>p(11)(98),clock=>clock,reset=>reset,s=>p(134)(98),cout=>p(135)(99));
FA_ff_483:FAff port map(x=>p(9)(99),y=>p(10)(99),Cin=>p(11)(99),clock=>clock,reset=>reset,s=>p(134)(99),cout=>p(135)(100));
FA_ff_484:FAff port map(x=>p(9)(100),y=>p(10)(100),Cin=>p(11)(100),clock=>clock,reset=>reset,s=>p(134)(100),cout=>p(135)(101));
FA_ff_485:FAff port map(x=>p(9)(101),y=>p(10)(101),Cin=>p(11)(101),clock=>clock,reset=>reset,s=>p(134)(101),cout=>p(135)(102));
FA_ff_486:FAff port map(x=>p(9)(102),y=>p(10)(102),Cin=>p(11)(102),clock=>clock,reset=>reset,s=>p(134)(102),cout=>p(135)(103));
FA_ff_487:FAff port map(x=>p(9)(103),y=>p(10)(103),Cin=>p(11)(103),clock=>clock,reset=>reset,s=>p(134)(103),cout=>p(135)(104));
FA_ff_488:FAff port map(x=>p(9)(104),y=>p(10)(104),Cin=>p(11)(104),clock=>clock,reset=>reset,s=>p(134)(104),cout=>p(135)(105));
FA_ff_489:FAff port map(x=>p(9)(105),y=>p(10)(105),Cin=>p(11)(105),clock=>clock,reset=>reset,s=>p(134)(105),cout=>p(135)(106));
FA_ff_490:FAff port map(x=>p(9)(106),y=>p(10)(106),Cin=>p(11)(106),clock=>clock,reset=>reset,s=>p(134)(106),cout=>p(135)(107));
FA_ff_491:FAff port map(x=>p(9)(107),y=>p(10)(107),Cin=>p(11)(107),clock=>clock,reset=>reset,s=>p(134)(107),cout=>p(135)(108));
FA_ff_492:FAff port map(x=>p(9)(108),y=>p(10)(108),Cin=>p(11)(108),clock=>clock,reset=>reset,s=>p(134)(108),cout=>p(135)(109));
FA_ff_493:FAff port map(x=>p(9)(109),y=>p(10)(109),Cin=>p(11)(109),clock=>clock,reset=>reset,s=>p(134)(109),cout=>p(135)(110));
FA_ff_494:FAff port map(x=>p(9)(110),y=>p(10)(110),Cin=>p(11)(110),clock=>clock,reset=>reset,s=>p(134)(110),cout=>p(135)(111));
FA_ff_495:FAff port map(x=>p(9)(111),y=>p(10)(111),Cin=>p(11)(111),clock=>clock,reset=>reset,s=>p(134)(111),cout=>p(135)(112));
FA_ff_496:FAff port map(x=>p(9)(112),y=>p(10)(112),Cin=>p(11)(112),clock=>clock,reset=>reset,s=>p(134)(112),cout=>p(135)(113));
FA_ff_497:FAff port map(x=>p(9)(113),y=>p(10)(113),Cin=>p(11)(113),clock=>clock,reset=>reset,s=>p(134)(113),cout=>p(135)(114));
FA_ff_498:FAff port map(x=>p(9)(114),y=>p(10)(114),Cin=>p(11)(114),clock=>clock,reset=>reset,s=>p(134)(114),cout=>p(135)(115));
FA_ff_499:FAff port map(x=>p(9)(115),y=>p(10)(115),Cin=>p(11)(115),clock=>clock,reset=>reset,s=>p(134)(115),cout=>p(135)(116));
FA_ff_500:FAff port map(x=>p(9)(116),y=>p(10)(116),Cin=>p(11)(116),clock=>clock,reset=>reset,s=>p(134)(116),cout=>p(135)(117));
FA_ff_501:FAff port map(x=>p(9)(117),y=>p(10)(117),Cin=>p(11)(117),clock=>clock,reset=>reset,s=>p(134)(117),cout=>p(135)(118));
FA_ff_502:FAff port map(x=>p(9)(118),y=>p(10)(118),Cin=>p(11)(118),clock=>clock,reset=>reset,s=>p(134)(118),cout=>p(135)(119));
FA_ff_503:FAff port map(x=>p(9)(119),y=>p(10)(119),Cin=>p(11)(119),clock=>clock,reset=>reset,s=>p(134)(119),cout=>p(135)(120));
FA_ff_504:FAff port map(x=>p(9)(120),y=>p(10)(120),Cin=>p(11)(120),clock=>clock,reset=>reset,s=>p(134)(120),cout=>p(135)(121));
FA_ff_505:FAff port map(x=>p(9)(121),y=>p(10)(121),Cin=>p(11)(121),clock=>clock,reset=>reset,s=>p(134)(121),cout=>p(135)(122));
FA_ff_506:FAff port map(x=>p(9)(122),y=>p(10)(122),Cin=>p(11)(122),clock=>clock,reset=>reset,s=>p(134)(122),cout=>p(135)(123));
FA_ff_507:FAff port map(x=>p(9)(123),y=>p(10)(123),Cin=>p(11)(123),clock=>clock,reset=>reset,s=>p(134)(123),cout=>p(135)(124));
FA_ff_508:FAff port map(x=>p(9)(124),y=>p(10)(124),Cin=>p(11)(124),clock=>clock,reset=>reset,s=>p(134)(124),cout=>p(135)(125));
FA_ff_509:FAff port map(x=>p(9)(125),y=>p(10)(125),Cin=>p(11)(125),clock=>clock,reset=>reset,s=>p(134)(125),cout=>p(135)(126));
FA_ff_510:FAff port map(x=>p(9)(126),y=>p(10)(126),Cin=>p(11)(126),clock=>clock,reset=>reset,s=>p(134)(126),cout=>p(135)(127));
FA_ff_511:FAff port map(x=>p(9)(127),y=>p(10)(127),Cin=>p(11)(127),clock=>clock,reset=>reset,s=>p(134)(127),cout=>p(135)(128));
FA_ff_512:FAff port map(x=>p(12)(0),y=>p(13)(0),Cin=>p(14)(0),clock=>clock,reset=>reset,s=>p(136)(0),cout=>p(137)(1));
FA_ff_513:FAff port map(x=>p(12)(1),y=>p(13)(1),Cin=>p(14)(1),clock=>clock,reset=>reset,s=>p(136)(1),cout=>p(137)(2));
FA_ff_514:FAff port map(x=>p(12)(2),y=>p(13)(2),Cin=>p(14)(2),clock=>clock,reset=>reset,s=>p(136)(2),cout=>p(137)(3));
FA_ff_515:FAff port map(x=>p(12)(3),y=>p(13)(3),Cin=>p(14)(3),clock=>clock,reset=>reset,s=>p(136)(3),cout=>p(137)(4));
FA_ff_516:FAff port map(x=>p(12)(4),y=>p(13)(4),Cin=>p(14)(4),clock=>clock,reset=>reset,s=>p(136)(4),cout=>p(137)(5));
FA_ff_517:FAff port map(x=>p(12)(5),y=>p(13)(5),Cin=>p(14)(5),clock=>clock,reset=>reset,s=>p(136)(5),cout=>p(137)(6));
FA_ff_518:FAff port map(x=>p(12)(6),y=>p(13)(6),Cin=>p(14)(6),clock=>clock,reset=>reset,s=>p(136)(6),cout=>p(137)(7));
FA_ff_519:FAff port map(x=>p(12)(7),y=>p(13)(7),Cin=>p(14)(7),clock=>clock,reset=>reset,s=>p(136)(7),cout=>p(137)(8));
FA_ff_520:FAff port map(x=>p(12)(8),y=>p(13)(8),Cin=>p(14)(8),clock=>clock,reset=>reset,s=>p(136)(8),cout=>p(137)(9));
FA_ff_521:FAff port map(x=>p(12)(9),y=>p(13)(9),Cin=>p(14)(9),clock=>clock,reset=>reset,s=>p(136)(9),cout=>p(137)(10));
FA_ff_522:FAff port map(x=>p(12)(10),y=>p(13)(10),Cin=>p(14)(10),clock=>clock,reset=>reset,s=>p(136)(10),cout=>p(137)(11));
FA_ff_523:FAff port map(x=>p(12)(11),y=>p(13)(11),Cin=>p(14)(11),clock=>clock,reset=>reset,s=>p(136)(11),cout=>p(137)(12));
FA_ff_524:FAff port map(x=>p(12)(12),y=>p(13)(12),Cin=>p(14)(12),clock=>clock,reset=>reset,s=>p(136)(12),cout=>p(137)(13));
FA_ff_525:FAff port map(x=>p(12)(13),y=>p(13)(13),Cin=>p(14)(13),clock=>clock,reset=>reset,s=>p(136)(13),cout=>p(137)(14));
FA_ff_526:FAff port map(x=>p(12)(14),y=>p(13)(14),Cin=>p(14)(14),clock=>clock,reset=>reset,s=>p(136)(14),cout=>p(137)(15));
FA_ff_527:FAff port map(x=>p(12)(15),y=>p(13)(15),Cin=>p(14)(15),clock=>clock,reset=>reset,s=>p(136)(15),cout=>p(137)(16));
FA_ff_528:FAff port map(x=>p(12)(16),y=>p(13)(16),Cin=>p(14)(16),clock=>clock,reset=>reset,s=>p(136)(16),cout=>p(137)(17));
FA_ff_529:FAff port map(x=>p(12)(17),y=>p(13)(17),Cin=>p(14)(17),clock=>clock,reset=>reset,s=>p(136)(17),cout=>p(137)(18));
FA_ff_530:FAff port map(x=>p(12)(18),y=>p(13)(18),Cin=>p(14)(18),clock=>clock,reset=>reset,s=>p(136)(18),cout=>p(137)(19));
FA_ff_531:FAff port map(x=>p(12)(19),y=>p(13)(19),Cin=>p(14)(19),clock=>clock,reset=>reset,s=>p(136)(19),cout=>p(137)(20));
FA_ff_532:FAff port map(x=>p(12)(20),y=>p(13)(20),Cin=>p(14)(20),clock=>clock,reset=>reset,s=>p(136)(20),cout=>p(137)(21));
FA_ff_533:FAff port map(x=>p(12)(21),y=>p(13)(21),Cin=>p(14)(21),clock=>clock,reset=>reset,s=>p(136)(21),cout=>p(137)(22));
FA_ff_534:FAff port map(x=>p(12)(22),y=>p(13)(22),Cin=>p(14)(22),clock=>clock,reset=>reset,s=>p(136)(22),cout=>p(137)(23));
FA_ff_535:FAff port map(x=>p(12)(23),y=>p(13)(23),Cin=>p(14)(23),clock=>clock,reset=>reset,s=>p(136)(23),cout=>p(137)(24));
FA_ff_536:FAff port map(x=>p(12)(24),y=>p(13)(24),Cin=>p(14)(24),clock=>clock,reset=>reset,s=>p(136)(24),cout=>p(137)(25));
FA_ff_537:FAff port map(x=>p(12)(25),y=>p(13)(25),Cin=>p(14)(25),clock=>clock,reset=>reset,s=>p(136)(25),cout=>p(137)(26));
FA_ff_538:FAff port map(x=>p(12)(26),y=>p(13)(26),Cin=>p(14)(26),clock=>clock,reset=>reset,s=>p(136)(26),cout=>p(137)(27));
FA_ff_539:FAff port map(x=>p(12)(27),y=>p(13)(27),Cin=>p(14)(27),clock=>clock,reset=>reset,s=>p(136)(27),cout=>p(137)(28));
FA_ff_540:FAff port map(x=>p(12)(28),y=>p(13)(28),Cin=>p(14)(28),clock=>clock,reset=>reset,s=>p(136)(28),cout=>p(137)(29));
FA_ff_541:FAff port map(x=>p(12)(29),y=>p(13)(29),Cin=>p(14)(29),clock=>clock,reset=>reset,s=>p(136)(29),cout=>p(137)(30));
FA_ff_542:FAff port map(x=>p(12)(30),y=>p(13)(30),Cin=>p(14)(30),clock=>clock,reset=>reset,s=>p(136)(30),cout=>p(137)(31));
FA_ff_543:FAff port map(x=>p(12)(31),y=>p(13)(31),Cin=>p(14)(31),clock=>clock,reset=>reset,s=>p(136)(31),cout=>p(137)(32));
FA_ff_544:FAff port map(x=>p(12)(32),y=>p(13)(32),Cin=>p(14)(32),clock=>clock,reset=>reset,s=>p(136)(32),cout=>p(137)(33));
FA_ff_545:FAff port map(x=>p(12)(33),y=>p(13)(33),Cin=>p(14)(33),clock=>clock,reset=>reset,s=>p(136)(33),cout=>p(137)(34));
FA_ff_546:FAff port map(x=>p(12)(34),y=>p(13)(34),Cin=>p(14)(34),clock=>clock,reset=>reset,s=>p(136)(34),cout=>p(137)(35));
FA_ff_547:FAff port map(x=>p(12)(35),y=>p(13)(35),Cin=>p(14)(35),clock=>clock,reset=>reset,s=>p(136)(35),cout=>p(137)(36));
FA_ff_548:FAff port map(x=>p(12)(36),y=>p(13)(36),Cin=>p(14)(36),clock=>clock,reset=>reset,s=>p(136)(36),cout=>p(137)(37));
FA_ff_549:FAff port map(x=>p(12)(37),y=>p(13)(37),Cin=>p(14)(37),clock=>clock,reset=>reset,s=>p(136)(37),cout=>p(137)(38));
FA_ff_550:FAff port map(x=>p(12)(38),y=>p(13)(38),Cin=>p(14)(38),clock=>clock,reset=>reset,s=>p(136)(38),cout=>p(137)(39));
FA_ff_551:FAff port map(x=>p(12)(39),y=>p(13)(39),Cin=>p(14)(39),clock=>clock,reset=>reset,s=>p(136)(39),cout=>p(137)(40));
FA_ff_552:FAff port map(x=>p(12)(40),y=>p(13)(40),Cin=>p(14)(40),clock=>clock,reset=>reset,s=>p(136)(40),cout=>p(137)(41));
FA_ff_553:FAff port map(x=>p(12)(41),y=>p(13)(41),Cin=>p(14)(41),clock=>clock,reset=>reset,s=>p(136)(41),cout=>p(137)(42));
FA_ff_554:FAff port map(x=>p(12)(42),y=>p(13)(42),Cin=>p(14)(42),clock=>clock,reset=>reset,s=>p(136)(42),cout=>p(137)(43));
FA_ff_555:FAff port map(x=>p(12)(43),y=>p(13)(43),Cin=>p(14)(43),clock=>clock,reset=>reset,s=>p(136)(43),cout=>p(137)(44));
FA_ff_556:FAff port map(x=>p(12)(44),y=>p(13)(44),Cin=>p(14)(44),clock=>clock,reset=>reset,s=>p(136)(44),cout=>p(137)(45));
FA_ff_557:FAff port map(x=>p(12)(45),y=>p(13)(45),Cin=>p(14)(45),clock=>clock,reset=>reset,s=>p(136)(45),cout=>p(137)(46));
FA_ff_558:FAff port map(x=>p(12)(46),y=>p(13)(46),Cin=>p(14)(46),clock=>clock,reset=>reset,s=>p(136)(46),cout=>p(137)(47));
FA_ff_559:FAff port map(x=>p(12)(47),y=>p(13)(47),Cin=>p(14)(47),clock=>clock,reset=>reset,s=>p(136)(47),cout=>p(137)(48));
FA_ff_560:FAff port map(x=>p(12)(48),y=>p(13)(48),Cin=>p(14)(48),clock=>clock,reset=>reset,s=>p(136)(48),cout=>p(137)(49));
FA_ff_561:FAff port map(x=>p(12)(49),y=>p(13)(49),Cin=>p(14)(49),clock=>clock,reset=>reset,s=>p(136)(49),cout=>p(137)(50));
FA_ff_562:FAff port map(x=>p(12)(50),y=>p(13)(50),Cin=>p(14)(50),clock=>clock,reset=>reset,s=>p(136)(50),cout=>p(137)(51));
FA_ff_563:FAff port map(x=>p(12)(51),y=>p(13)(51),Cin=>p(14)(51),clock=>clock,reset=>reset,s=>p(136)(51),cout=>p(137)(52));
FA_ff_564:FAff port map(x=>p(12)(52),y=>p(13)(52),Cin=>p(14)(52),clock=>clock,reset=>reset,s=>p(136)(52),cout=>p(137)(53));
FA_ff_565:FAff port map(x=>p(12)(53),y=>p(13)(53),Cin=>p(14)(53),clock=>clock,reset=>reset,s=>p(136)(53),cout=>p(137)(54));
FA_ff_566:FAff port map(x=>p(12)(54),y=>p(13)(54),Cin=>p(14)(54),clock=>clock,reset=>reset,s=>p(136)(54),cout=>p(137)(55));
FA_ff_567:FAff port map(x=>p(12)(55),y=>p(13)(55),Cin=>p(14)(55),clock=>clock,reset=>reset,s=>p(136)(55),cout=>p(137)(56));
FA_ff_568:FAff port map(x=>p(12)(56),y=>p(13)(56),Cin=>p(14)(56),clock=>clock,reset=>reset,s=>p(136)(56),cout=>p(137)(57));
FA_ff_569:FAff port map(x=>p(12)(57),y=>p(13)(57),Cin=>p(14)(57),clock=>clock,reset=>reset,s=>p(136)(57),cout=>p(137)(58));
FA_ff_570:FAff port map(x=>p(12)(58),y=>p(13)(58),Cin=>p(14)(58),clock=>clock,reset=>reset,s=>p(136)(58),cout=>p(137)(59));
FA_ff_571:FAff port map(x=>p(12)(59),y=>p(13)(59),Cin=>p(14)(59),clock=>clock,reset=>reset,s=>p(136)(59),cout=>p(137)(60));
FA_ff_572:FAff port map(x=>p(12)(60),y=>p(13)(60),Cin=>p(14)(60),clock=>clock,reset=>reset,s=>p(136)(60),cout=>p(137)(61));
FA_ff_573:FAff port map(x=>p(12)(61),y=>p(13)(61),Cin=>p(14)(61),clock=>clock,reset=>reset,s=>p(136)(61),cout=>p(137)(62));
FA_ff_574:FAff port map(x=>p(12)(62),y=>p(13)(62),Cin=>p(14)(62),clock=>clock,reset=>reset,s=>p(136)(62),cout=>p(137)(63));
FA_ff_575:FAff port map(x=>p(12)(63),y=>p(13)(63),Cin=>p(14)(63),clock=>clock,reset=>reset,s=>p(136)(63),cout=>p(137)(64));
FA_ff_576:FAff port map(x=>p(12)(64),y=>p(13)(64),Cin=>p(14)(64),clock=>clock,reset=>reset,s=>p(136)(64),cout=>p(137)(65));
FA_ff_577:FAff port map(x=>p(12)(65),y=>p(13)(65),Cin=>p(14)(65),clock=>clock,reset=>reset,s=>p(136)(65),cout=>p(137)(66));
FA_ff_578:FAff port map(x=>p(12)(66),y=>p(13)(66),Cin=>p(14)(66),clock=>clock,reset=>reset,s=>p(136)(66),cout=>p(137)(67));
FA_ff_579:FAff port map(x=>p(12)(67),y=>p(13)(67),Cin=>p(14)(67),clock=>clock,reset=>reset,s=>p(136)(67),cout=>p(137)(68));
FA_ff_580:FAff port map(x=>p(12)(68),y=>p(13)(68),Cin=>p(14)(68),clock=>clock,reset=>reset,s=>p(136)(68),cout=>p(137)(69));
FA_ff_581:FAff port map(x=>p(12)(69),y=>p(13)(69),Cin=>p(14)(69),clock=>clock,reset=>reset,s=>p(136)(69),cout=>p(137)(70));
FA_ff_582:FAff port map(x=>p(12)(70),y=>p(13)(70),Cin=>p(14)(70),clock=>clock,reset=>reset,s=>p(136)(70),cout=>p(137)(71));
FA_ff_583:FAff port map(x=>p(12)(71),y=>p(13)(71),Cin=>p(14)(71),clock=>clock,reset=>reset,s=>p(136)(71),cout=>p(137)(72));
FA_ff_584:FAff port map(x=>p(12)(72),y=>p(13)(72),Cin=>p(14)(72),clock=>clock,reset=>reset,s=>p(136)(72),cout=>p(137)(73));
FA_ff_585:FAff port map(x=>p(12)(73),y=>p(13)(73),Cin=>p(14)(73),clock=>clock,reset=>reset,s=>p(136)(73),cout=>p(137)(74));
FA_ff_586:FAff port map(x=>p(12)(74),y=>p(13)(74),Cin=>p(14)(74),clock=>clock,reset=>reset,s=>p(136)(74),cout=>p(137)(75));
FA_ff_587:FAff port map(x=>p(12)(75),y=>p(13)(75),Cin=>p(14)(75),clock=>clock,reset=>reset,s=>p(136)(75),cout=>p(137)(76));
FA_ff_588:FAff port map(x=>p(12)(76),y=>p(13)(76),Cin=>p(14)(76),clock=>clock,reset=>reset,s=>p(136)(76),cout=>p(137)(77));
FA_ff_589:FAff port map(x=>p(12)(77),y=>p(13)(77),Cin=>p(14)(77),clock=>clock,reset=>reset,s=>p(136)(77),cout=>p(137)(78));
FA_ff_590:FAff port map(x=>p(12)(78),y=>p(13)(78),Cin=>p(14)(78),clock=>clock,reset=>reset,s=>p(136)(78),cout=>p(137)(79));
FA_ff_591:FAff port map(x=>p(12)(79),y=>p(13)(79),Cin=>p(14)(79),clock=>clock,reset=>reset,s=>p(136)(79),cout=>p(137)(80));
FA_ff_592:FAff port map(x=>p(12)(80),y=>p(13)(80),Cin=>p(14)(80),clock=>clock,reset=>reset,s=>p(136)(80),cout=>p(137)(81));
FA_ff_593:FAff port map(x=>p(12)(81),y=>p(13)(81),Cin=>p(14)(81),clock=>clock,reset=>reset,s=>p(136)(81),cout=>p(137)(82));
FA_ff_594:FAff port map(x=>p(12)(82),y=>p(13)(82),Cin=>p(14)(82),clock=>clock,reset=>reset,s=>p(136)(82),cout=>p(137)(83));
FA_ff_595:FAff port map(x=>p(12)(83),y=>p(13)(83),Cin=>p(14)(83),clock=>clock,reset=>reset,s=>p(136)(83),cout=>p(137)(84));
FA_ff_596:FAff port map(x=>p(12)(84),y=>p(13)(84),Cin=>p(14)(84),clock=>clock,reset=>reset,s=>p(136)(84),cout=>p(137)(85));
FA_ff_597:FAff port map(x=>p(12)(85),y=>p(13)(85),Cin=>p(14)(85),clock=>clock,reset=>reset,s=>p(136)(85),cout=>p(137)(86));
FA_ff_598:FAff port map(x=>p(12)(86),y=>p(13)(86),Cin=>p(14)(86),clock=>clock,reset=>reset,s=>p(136)(86),cout=>p(137)(87));
FA_ff_599:FAff port map(x=>p(12)(87),y=>p(13)(87),Cin=>p(14)(87),clock=>clock,reset=>reset,s=>p(136)(87),cout=>p(137)(88));
FA_ff_600:FAff port map(x=>p(12)(88),y=>p(13)(88),Cin=>p(14)(88),clock=>clock,reset=>reset,s=>p(136)(88),cout=>p(137)(89));
FA_ff_601:FAff port map(x=>p(12)(89),y=>p(13)(89),Cin=>p(14)(89),clock=>clock,reset=>reset,s=>p(136)(89),cout=>p(137)(90));
FA_ff_602:FAff port map(x=>p(12)(90),y=>p(13)(90),Cin=>p(14)(90),clock=>clock,reset=>reset,s=>p(136)(90),cout=>p(137)(91));
FA_ff_603:FAff port map(x=>p(12)(91),y=>p(13)(91),Cin=>p(14)(91),clock=>clock,reset=>reset,s=>p(136)(91),cout=>p(137)(92));
FA_ff_604:FAff port map(x=>p(12)(92),y=>p(13)(92),Cin=>p(14)(92),clock=>clock,reset=>reset,s=>p(136)(92),cout=>p(137)(93));
FA_ff_605:FAff port map(x=>p(12)(93),y=>p(13)(93),Cin=>p(14)(93),clock=>clock,reset=>reset,s=>p(136)(93),cout=>p(137)(94));
FA_ff_606:FAff port map(x=>p(12)(94),y=>p(13)(94),Cin=>p(14)(94),clock=>clock,reset=>reset,s=>p(136)(94),cout=>p(137)(95));
FA_ff_607:FAff port map(x=>p(12)(95),y=>p(13)(95),Cin=>p(14)(95),clock=>clock,reset=>reset,s=>p(136)(95),cout=>p(137)(96));
FA_ff_608:FAff port map(x=>p(12)(96),y=>p(13)(96),Cin=>p(14)(96),clock=>clock,reset=>reset,s=>p(136)(96),cout=>p(137)(97));
FA_ff_609:FAff port map(x=>p(12)(97),y=>p(13)(97),Cin=>p(14)(97),clock=>clock,reset=>reset,s=>p(136)(97),cout=>p(137)(98));
FA_ff_610:FAff port map(x=>p(12)(98),y=>p(13)(98),Cin=>p(14)(98),clock=>clock,reset=>reset,s=>p(136)(98),cout=>p(137)(99));
FA_ff_611:FAff port map(x=>p(12)(99),y=>p(13)(99),Cin=>p(14)(99),clock=>clock,reset=>reset,s=>p(136)(99),cout=>p(137)(100));
FA_ff_612:FAff port map(x=>p(12)(100),y=>p(13)(100),Cin=>p(14)(100),clock=>clock,reset=>reset,s=>p(136)(100),cout=>p(137)(101));
FA_ff_613:FAff port map(x=>p(12)(101),y=>p(13)(101),Cin=>p(14)(101),clock=>clock,reset=>reset,s=>p(136)(101),cout=>p(137)(102));
FA_ff_614:FAff port map(x=>p(12)(102),y=>p(13)(102),Cin=>p(14)(102),clock=>clock,reset=>reset,s=>p(136)(102),cout=>p(137)(103));
FA_ff_615:FAff port map(x=>p(12)(103),y=>p(13)(103),Cin=>p(14)(103),clock=>clock,reset=>reset,s=>p(136)(103),cout=>p(137)(104));
FA_ff_616:FAff port map(x=>p(12)(104),y=>p(13)(104),Cin=>p(14)(104),clock=>clock,reset=>reset,s=>p(136)(104),cout=>p(137)(105));
FA_ff_617:FAff port map(x=>p(12)(105),y=>p(13)(105),Cin=>p(14)(105),clock=>clock,reset=>reset,s=>p(136)(105),cout=>p(137)(106));
FA_ff_618:FAff port map(x=>p(12)(106),y=>p(13)(106),Cin=>p(14)(106),clock=>clock,reset=>reset,s=>p(136)(106),cout=>p(137)(107));
FA_ff_619:FAff port map(x=>p(12)(107),y=>p(13)(107),Cin=>p(14)(107),clock=>clock,reset=>reset,s=>p(136)(107),cout=>p(137)(108));
FA_ff_620:FAff port map(x=>p(12)(108),y=>p(13)(108),Cin=>p(14)(108),clock=>clock,reset=>reset,s=>p(136)(108),cout=>p(137)(109));
FA_ff_621:FAff port map(x=>p(12)(109),y=>p(13)(109),Cin=>p(14)(109),clock=>clock,reset=>reset,s=>p(136)(109),cout=>p(137)(110));
FA_ff_622:FAff port map(x=>p(12)(110),y=>p(13)(110),Cin=>p(14)(110),clock=>clock,reset=>reset,s=>p(136)(110),cout=>p(137)(111));
FA_ff_623:FAff port map(x=>p(12)(111),y=>p(13)(111),Cin=>p(14)(111),clock=>clock,reset=>reset,s=>p(136)(111),cout=>p(137)(112));
FA_ff_624:FAff port map(x=>p(12)(112),y=>p(13)(112),Cin=>p(14)(112),clock=>clock,reset=>reset,s=>p(136)(112),cout=>p(137)(113));
FA_ff_625:FAff port map(x=>p(12)(113),y=>p(13)(113),Cin=>p(14)(113),clock=>clock,reset=>reset,s=>p(136)(113),cout=>p(137)(114));
FA_ff_626:FAff port map(x=>p(12)(114),y=>p(13)(114),Cin=>p(14)(114),clock=>clock,reset=>reset,s=>p(136)(114),cout=>p(137)(115));
FA_ff_627:FAff port map(x=>p(12)(115),y=>p(13)(115),Cin=>p(14)(115),clock=>clock,reset=>reset,s=>p(136)(115),cout=>p(137)(116));
FA_ff_628:FAff port map(x=>p(12)(116),y=>p(13)(116),Cin=>p(14)(116),clock=>clock,reset=>reset,s=>p(136)(116),cout=>p(137)(117));
FA_ff_629:FAff port map(x=>p(12)(117),y=>p(13)(117),Cin=>p(14)(117),clock=>clock,reset=>reset,s=>p(136)(117),cout=>p(137)(118));
FA_ff_630:FAff port map(x=>p(12)(118),y=>p(13)(118),Cin=>p(14)(118),clock=>clock,reset=>reset,s=>p(136)(118),cout=>p(137)(119));
FA_ff_631:FAff port map(x=>p(12)(119),y=>p(13)(119),Cin=>p(14)(119),clock=>clock,reset=>reset,s=>p(136)(119),cout=>p(137)(120));
FA_ff_632:FAff port map(x=>p(12)(120),y=>p(13)(120),Cin=>p(14)(120),clock=>clock,reset=>reset,s=>p(136)(120),cout=>p(137)(121));
FA_ff_633:FAff port map(x=>p(12)(121),y=>p(13)(121),Cin=>p(14)(121),clock=>clock,reset=>reset,s=>p(136)(121),cout=>p(137)(122));
FA_ff_634:FAff port map(x=>p(12)(122),y=>p(13)(122),Cin=>p(14)(122),clock=>clock,reset=>reset,s=>p(136)(122),cout=>p(137)(123));
FA_ff_635:FAff port map(x=>p(12)(123),y=>p(13)(123),Cin=>p(14)(123),clock=>clock,reset=>reset,s=>p(136)(123),cout=>p(137)(124));
FA_ff_636:FAff port map(x=>p(12)(124),y=>p(13)(124),Cin=>p(14)(124),clock=>clock,reset=>reset,s=>p(136)(124),cout=>p(137)(125));
FA_ff_637:FAff port map(x=>p(12)(125),y=>p(13)(125),Cin=>p(14)(125),clock=>clock,reset=>reset,s=>p(136)(125),cout=>p(137)(126));
FA_ff_638:FAff port map(x=>p(12)(126),y=>p(13)(126),Cin=>p(14)(126),clock=>clock,reset=>reset,s=>p(136)(126),cout=>p(137)(127));
FA_ff_639:FAff port map(x=>p(12)(127),y=>p(13)(127),Cin=>p(14)(127),clock=>clock,reset=>reset,s=>p(136)(127),cout=>p(137)(128));
FA_ff_640:FAff port map(x=>p(15)(0),y=>p(16)(0),Cin=>p(17)(0),clock=>clock,reset=>reset,s=>p(138)(0),cout=>p(139)(1));
FA_ff_641:FAff port map(x=>p(15)(1),y=>p(16)(1),Cin=>p(17)(1),clock=>clock,reset=>reset,s=>p(138)(1),cout=>p(139)(2));
FA_ff_642:FAff port map(x=>p(15)(2),y=>p(16)(2),Cin=>p(17)(2),clock=>clock,reset=>reset,s=>p(138)(2),cout=>p(139)(3));
FA_ff_643:FAff port map(x=>p(15)(3),y=>p(16)(3),Cin=>p(17)(3),clock=>clock,reset=>reset,s=>p(138)(3),cout=>p(139)(4));
FA_ff_644:FAff port map(x=>p(15)(4),y=>p(16)(4),Cin=>p(17)(4),clock=>clock,reset=>reset,s=>p(138)(4),cout=>p(139)(5));
FA_ff_645:FAff port map(x=>p(15)(5),y=>p(16)(5),Cin=>p(17)(5),clock=>clock,reset=>reset,s=>p(138)(5),cout=>p(139)(6));
FA_ff_646:FAff port map(x=>p(15)(6),y=>p(16)(6),Cin=>p(17)(6),clock=>clock,reset=>reset,s=>p(138)(6),cout=>p(139)(7));
FA_ff_647:FAff port map(x=>p(15)(7),y=>p(16)(7),Cin=>p(17)(7),clock=>clock,reset=>reset,s=>p(138)(7),cout=>p(139)(8));
FA_ff_648:FAff port map(x=>p(15)(8),y=>p(16)(8),Cin=>p(17)(8),clock=>clock,reset=>reset,s=>p(138)(8),cout=>p(139)(9));
FA_ff_649:FAff port map(x=>p(15)(9),y=>p(16)(9),Cin=>p(17)(9),clock=>clock,reset=>reset,s=>p(138)(9),cout=>p(139)(10));
FA_ff_650:FAff port map(x=>p(15)(10),y=>p(16)(10),Cin=>p(17)(10),clock=>clock,reset=>reset,s=>p(138)(10),cout=>p(139)(11));
FA_ff_651:FAff port map(x=>p(15)(11),y=>p(16)(11),Cin=>p(17)(11),clock=>clock,reset=>reset,s=>p(138)(11),cout=>p(139)(12));
FA_ff_652:FAff port map(x=>p(15)(12),y=>p(16)(12),Cin=>p(17)(12),clock=>clock,reset=>reset,s=>p(138)(12),cout=>p(139)(13));
FA_ff_653:FAff port map(x=>p(15)(13),y=>p(16)(13),Cin=>p(17)(13),clock=>clock,reset=>reset,s=>p(138)(13),cout=>p(139)(14));
FA_ff_654:FAff port map(x=>p(15)(14),y=>p(16)(14),Cin=>p(17)(14),clock=>clock,reset=>reset,s=>p(138)(14),cout=>p(139)(15));
FA_ff_655:FAff port map(x=>p(15)(15),y=>p(16)(15),Cin=>p(17)(15),clock=>clock,reset=>reset,s=>p(138)(15),cout=>p(139)(16));
FA_ff_656:FAff port map(x=>p(15)(16),y=>p(16)(16),Cin=>p(17)(16),clock=>clock,reset=>reset,s=>p(138)(16),cout=>p(139)(17));
FA_ff_657:FAff port map(x=>p(15)(17),y=>p(16)(17),Cin=>p(17)(17),clock=>clock,reset=>reset,s=>p(138)(17),cout=>p(139)(18));
FA_ff_658:FAff port map(x=>p(15)(18),y=>p(16)(18),Cin=>p(17)(18),clock=>clock,reset=>reset,s=>p(138)(18),cout=>p(139)(19));
FA_ff_659:FAff port map(x=>p(15)(19),y=>p(16)(19),Cin=>p(17)(19),clock=>clock,reset=>reset,s=>p(138)(19),cout=>p(139)(20));
FA_ff_660:FAff port map(x=>p(15)(20),y=>p(16)(20),Cin=>p(17)(20),clock=>clock,reset=>reset,s=>p(138)(20),cout=>p(139)(21));
FA_ff_661:FAff port map(x=>p(15)(21),y=>p(16)(21),Cin=>p(17)(21),clock=>clock,reset=>reset,s=>p(138)(21),cout=>p(139)(22));
FA_ff_662:FAff port map(x=>p(15)(22),y=>p(16)(22),Cin=>p(17)(22),clock=>clock,reset=>reset,s=>p(138)(22),cout=>p(139)(23));
FA_ff_663:FAff port map(x=>p(15)(23),y=>p(16)(23),Cin=>p(17)(23),clock=>clock,reset=>reset,s=>p(138)(23),cout=>p(139)(24));
FA_ff_664:FAff port map(x=>p(15)(24),y=>p(16)(24),Cin=>p(17)(24),clock=>clock,reset=>reset,s=>p(138)(24),cout=>p(139)(25));
FA_ff_665:FAff port map(x=>p(15)(25),y=>p(16)(25),Cin=>p(17)(25),clock=>clock,reset=>reset,s=>p(138)(25),cout=>p(139)(26));
FA_ff_666:FAff port map(x=>p(15)(26),y=>p(16)(26),Cin=>p(17)(26),clock=>clock,reset=>reset,s=>p(138)(26),cout=>p(139)(27));
FA_ff_667:FAff port map(x=>p(15)(27),y=>p(16)(27),Cin=>p(17)(27),clock=>clock,reset=>reset,s=>p(138)(27),cout=>p(139)(28));
FA_ff_668:FAff port map(x=>p(15)(28),y=>p(16)(28),Cin=>p(17)(28),clock=>clock,reset=>reset,s=>p(138)(28),cout=>p(139)(29));
FA_ff_669:FAff port map(x=>p(15)(29),y=>p(16)(29),Cin=>p(17)(29),clock=>clock,reset=>reset,s=>p(138)(29),cout=>p(139)(30));
FA_ff_670:FAff port map(x=>p(15)(30),y=>p(16)(30),Cin=>p(17)(30),clock=>clock,reset=>reset,s=>p(138)(30),cout=>p(139)(31));
FA_ff_671:FAff port map(x=>p(15)(31),y=>p(16)(31),Cin=>p(17)(31),clock=>clock,reset=>reset,s=>p(138)(31),cout=>p(139)(32));
FA_ff_672:FAff port map(x=>p(15)(32),y=>p(16)(32),Cin=>p(17)(32),clock=>clock,reset=>reset,s=>p(138)(32),cout=>p(139)(33));
FA_ff_673:FAff port map(x=>p(15)(33),y=>p(16)(33),Cin=>p(17)(33),clock=>clock,reset=>reset,s=>p(138)(33),cout=>p(139)(34));
FA_ff_674:FAff port map(x=>p(15)(34),y=>p(16)(34),Cin=>p(17)(34),clock=>clock,reset=>reset,s=>p(138)(34),cout=>p(139)(35));
FA_ff_675:FAff port map(x=>p(15)(35),y=>p(16)(35),Cin=>p(17)(35),clock=>clock,reset=>reset,s=>p(138)(35),cout=>p(139)(36));
FA_ff_676:FAff port map(x=>p(15)(36),y=>p(16)(36),Cin=>p(17)(36),clock=>clock,reset=>reset,s=>p(138)(36),cout=>p(139)(37));
FA_ff_677:FAff port map(x=>p(15)(37),y=>p(16)(37),Cin=>p(17)(37),clock=>clock,reset=>reset,s=>p(138)(37),cout=>p(139)(38));
FA_ff_678:FAff port map(x=>p(15)(38),y=>p(16)(38),Cin=>p(17)(38),clock=>clock,reset=>reset,s=>p(138)(38),cout=>p(139)(39));
FA_ff_679:FAff port map(x=>p(15)(39),y=>p(16)(39),Cin=>p(17)(39),clock=>clock,reset=>reset,s=>p(138)(39),cout=>p(139)(40));
FA_ff_680:FAff port map(x=>p(15)(40),y=>p(16)(40),Cin=>p(17)(40),clock=>clock,reset=>reset,s=>p(138)(40),cout=>p(139)(41));
FA_ff_681:FAff port map(x=>p(15)(41),y=>p(16)(41),Cin=>p(17)(41),clock=>clock,reset=>reset,s=>p(138)(41),cout=>p(139)(42));
FA_ff_682:FAff port map(x=>p(15)(42),y=>p(16)(42),Cin=>p(17)(42),clock=>clock,reset=>reset,s=>p(138)(42),cout=>p(139)(43));
FA_ff_683:FAff port map(x=>p(15)(43),y=>p(16)(43),Cin=>p(17)(43),clock=>clock,reset=>reset,s=>p(138)(43),cout=>p(139)(44));
FA_ff_684:FAff port map(x=>p(15)(44),y=>p(16)(44),Cin=>p(17)(44),clock=>clock,reset=>reset,s=>p(138)(44),cout=>p(139)(45));
FA_ff_685:FAff port map(x=>p(15)(45),y=>p(16)(45),Cin=>p(17)(45),clock=>clock,reset=>reset,s=>p(138)(45),cout=>p(139)(46));
FA_ff_686:FAff port map(x=>p(15)(46),y=>p(16)(46),Cin=>p(17)(46),clock=>clock,reset=>reset,s=>p(138)(46),cout=>p(139)(47));
FA_ff_687:FAff port map(x=>p(15)(47),y=>p(16)(47),Cin=>p(17)(47),clock=>clock,reset=>reset,s=>p(138)(47),cout=>p(139)(48));
FA_ff_688:FAff port map(x=>p(15)(48),y=>p(16)(48),Cin=>p(17)(48),clock=>clock,reset=>reset,s=>p(138)(48),cout=>p(139)(49));
FA_ff_689:FAff port map(x=>p(15)(49),y=>p(16)(49),Cin=>p(17)(49),clock=>clock,reset=>reset,s=>p(138)(49),cout=>p(139)(50));
FA_ff_690:FAff port map(x=>p(15)(50),y=>p(16)(50),Cin=>p(17)(50),clock=>clock,reset=>reset,s=>p(138)(50),cout=>p(139)(51));
FA_ff_691:FAff port map(x=>p(15)(51),y=>p(16)(51),Cin=>p(17)(51),clock=>clock,reset=>reset,s=>p(138)(51),cout=>p(139)(52));
FA_ff_692:FAff port map(x=>p(15)(52),y=>p(16)(52),Cin=>p(17)(52),clock=>clock,reset=>reset,s=>p(138)(52),cout=>p(139)(53));
FA_ff_693:FAff port map(x=>p(15)(53),y=>p(16)(53),Cin=>p(17)(53),clock=>clock,reset=>reset,s=>p(138)(53),cout=>p(139)(54));
FA_ff_694:FAff port map(x=>p(15)(54),y=>p(16)(54),Cin=>p(17)(54),clock=>clock,reset=>reset,s=>p(138)(54),cout=>p(139)(55));
FA_ff_695:FAff port map(x=>p(15)(55),y=>p(16)(55),Cin=>p(17)(55),clock=>clock,reset=>reset,s=>p(138)(55),cout=>p(139)(56));
FA_ff_696:FAff port map(x=>p(15)(56),y=>p(16)(56),Cin=>p(17)(56),clock=>clock,reset=>reset,s=>p(138)(56),cout=>p(139)(57));
FA_ff_697:FAff port map(x=>p(15)(57),y=>p(16)(57),Cin=>p(17)(57),clock=>clock,reset=>reset,s=>p(138)(57),cout=>p(139)(58));
FA_ff_698:FAff port map(x=>p(15)(58),y=>p(16)(58),Cin=>p(17)(58),clock=>clock,reset=>reset,s=>p(138)(58),cout=>p(139)(59));
FA_ff_699:FAff port map(x=>p(15)(59),y=>p(16)(59),Cin=>p(17)(59),clock=>clock,reset=>reset,s=>p(138)(59),cout=>p(139)(60));
FA_ff_700:FAff port map(x=>p(15)(60),y=>p(16)(60),Cin=>p(17)(60),clock=>clock,reset=>reset,s=>p(138)(60),cout=>p(139)(61));
FA_ff_701:FAff port map(x=>p(15)(61),y=>p(16)(61),Cin=>p(17)(61),clock=>clock,reset=>reset,s=>p(138)(61),cout=>p(139)(62));
FA_ff_702:FAff port map(x=>p(15)(62),y=>p(16)(62),Cin=>p(17)(62),clock=>clock,reset=>reset,s=>p(138)(62),cout=>p(139)(63));
FA_ff_703:FAff port map(x=>p(15)(63),y=>p(16)(63),Cin=>p(17)(63),clock=>clock,reset=>reset,s=>p(138)(63),cout=>p(139)(64));
FA_ff_704:FAff port map(x=>p(15)(64),y=>p(16)(64),Cin=>p(17)(64),clock=>clock,reset=>reset,s=>p(138)(64),cout=>p(139)(65));
FA_ff_705:FAff port map(x=>p(15)(65),y=>p(16)(65),Cin=>p(17)(65),clock=>clock,reset=>reset,s=>p(138)(65),cout=>p(139)(66));
FA_ff_706:FAff port map(x=>p(15)(66),y=>p(16)(66),Cin=>p(17)(66),clock=>clock,reset=>reset,s=>p(138)(66),cout=>p(139)(67));
FA_ff_707:FAff port map(x=>p(15)(67),y=>p(16)(67),Cin=>p(17)(67),clock=>clock,reset=>reset,s=>p(138)(67),cout=>p(139)(68));
FA_ff_708:FAff port map(x=>p(15)(68),y=>p(16)(68),Cin=>p(17)(68),clock=>clock,reset=>reset,s=>p(138)(68),cout=>p(139)(69));
FA_ff_709:FAff port map(x=>p(15)(69),y=>p(16)(69),Cin=>p(17)(69),clock=>clock,reset=>reset,s=>p(138)(69),cout=>p(139)(70));
FA_ff_710:FAff port map(x=>p(15)(70),y=>p(16)(70),Cin=>p(17)(70),clock=>clock,reset=>reset,s=>p(138)(70),cout=>p(139)(71));
FA_ff_711:FAff port map(x=>p(15)(71),y=>p(16)(71),Cin=>p(17)(71),clock=>clock,reset=>reset,s=>p(138)(71),cout=>p(139)(72));
FA_ff_712:FAff port map(x=>p(15)(72),y=>p(16)(72),Cin=>p(17)(72),clock=>clock,reset=>reset,s=>p(138)(72),cout=>p(139)(73));
FA_ff_713:FAff port map(x=>p(15)(73),y=>p(16)(73),Cin=>p(17)(73),clock=>clock,reset=>reset,s=>p(138)(73),cout=>p(139)(74));
FA_ff_714:FAff port map(x=>p(15)(74),y=>p(16)(74),Cin=>p(17)(74),clock=>clock,reset=>reset,s=>p(138)(74),cout=>p(139)(75));
FA_ff_715:FAff port map(x=>p(15)(75),y=>p(16)(75),Cin=>p(17)(75),clock=>clock,reset=>reset,s=>p(138)(75),cout=>p(139)(76));
FA_ff_716:FAff port map(x=>p(15)(76),y=>p(16)(76),Cin=>p(17)(76),clock=>clock,reset=>reset,s=>p(138)(76),cout=>p(139)(77));
FA_ff_717:FAff port map(x=>p(15)(77),y=>p(16)(77),Cin=>p(17)(77),clock=>clock,reset=>reset,s=>p(138)(77),cout=>p(139)(78));
FA_ff_718:FAff port map(x=>p(15)(78),y=>p(16)(78),Cin=>p(17)(78),clock=>clock,reset=>reset,s=>p(138)(78),cout=>p(139)(79));
FA_ff_719:FAff port map(x=>p(15)(79),y=>p(16)(79),Cin=>p(17)(79),clock=>clock,reset=>reset,s=>p(138)(79),cout=>p(139)(80));
FA_ff_720:FAff port map(x=>p(15)(80),y=>p(16)(80),Cin=>p(17)(80),clock=>clock,reset=>reset,s=>p(138)(80),cout=>p(139)(81));
FA_ff_721:FAff port map(x=>p(15)(81),y=>p(16)(81),Cin=>p(17)(81),clock=>clock,reset=>reset,s=>p(138)(81),cout=>p(139)(82));
FA_ff_722:FAff port map(x=>p(15)(82),y=>p(16)(82),Cin=>p(17)(82),clock=>clock,reset=>reset,s=>p(138)(82),cout=>p(139)(83));
FA_ff_723:FAff port map(x=>p(15)(83),y=>p(16)(83),Cin=>p(17)(83),clock=>clock,reset=>reset,s=>p(138)(83),cout=>p(139)(84));
FA_ff_724:FAff port map(x=>p(15)(84),y=>p(16)(84),Cin=>p(17)(84),clock=>clock,reset=>reset,s=>p(138)(84),cout=>p(139)(85));
FA_ff_725:FAff port map(x=>p(15)(85),y=>p(16)(85),Cin=>p(17)(85),clock=>clock,reset=>reset,s=>p(138)(85),cout=>p(139)(86));
FA_ff_726:FAff port map(x=>p(15)(86),y=>p(16)(86),Cin=>p(17)(86),clock=>clock,reset=>reset,s=>p(138)(86),cout=>p(139)(87));
FA_ff_727:FAff port map(x=>p(15)(87),y=>p(16)(87),Cin=>p(17)(87),clock=>clock,reset=>reset,s=>p(138)(87),cout=>p(139)(88));
FA_ff_728:FAff port map(x=>p(15)(88),y=>p(16)(88),Cin=>p(17)(88),clock=>clock,reset=>reset,s=>p(138)(88),cout=>p(139)(89));
FA_ff_729:FAff port map(x=>p(15)(89),y=>p(16)(89),Cin=>p(17)(89),clock=>clock,reset=>reset,s=>p(138)(89),cout=>p(139)(90));
FA_ff_730:FAff port map(x=>p(15)(90),y=>p(16)(90),Cin=>p(17)(90),clock=>clock,reset=>reset,s=>p(138)(90),cout=>p(139)(91));
FA_ff_731:FAff port map(x=>p(15)(91),y=>p(16)(91),Cin=>p(17)(91),clock=>clock,reset=>reset,s=>p(138)(91),cout=>p(139)(92));
FA_ff_732:FAff port map(x=>p(15)(92),y=>p(16)(92),Cin=>p(17)(92),clock=>clock,reset=>reset,s=>p(138)(92),cout=>p(139)(93));
FA_ff_733:FAff port map(x=>p(15)(93),y=>p(16)(93),Cin=>p(17)(93),clock=>clock,reset=>reset,s=>p(138)(93),cout=>p(139)(94));
FA_ff_734:FAff port map(x=>p(15)(94),y=>p(16)(94),Cin=>p(17)(94),clock=>clock,reset=>reset,s=>p(138)(94),cout=>p(139)(95));
FA_ff_735:FAff port map(x=>p(15)(95),y=>p(16)(95),Cin=>p(17)(95),clock=>clock,reset=>reset,s=>p(138)(95),cout=>p(139)(96));
FA_ff_736:FAff port map(x=>p(15)(96),y=>p(16)(96),Cin=>p(17)(96),clock=>clock,reset=>reset,s=>p(138)(96),cout=>p(139)(97));
FA_ff_737:FAff port map(x=>p(15)(97),y=>p(16)(97),Cin=>p(17)(97),clock=>clock,reset=>reset,s=>p(138)(97),cout=>p(139)(98));
FA_ff_738:FAff port map(x=>p(15)(98),y=>p(16)(98),Cin=>p(17)(98),clock=>clock,reset=>reset,s=>p(138)(98),cout=>p(139)(99));
FA_ff_739:FAff port map(x=>p(15)(99),y=>p(16)(99),Cin=>p(17)(99),clock=>clock,reset=>reset,s=>p(138)(99),cout=>p(139)(100));
FA_ff_740:FAff port map(x=>p(15)(100),y=>p(16)(100),Cin=>p(17)(100),clock=>clock,reset=>reset,s=>p(138)(100),cout=>p(139)(101));
FA_ff_741:FAff port map(x=>p(15)(101),y=>p(16)(101),Cin=>p(17)(101),clock=>clock,reset=>reset,s=>p(138)(101),cout=>p(139)(102));
FA_ff_742:FAff port map(x=>p(15)(102),y=>p(16)(102),Cin=>p(17)(102),clock=>clock,reset=>reset,s=>p(138)(102),cout=>p(139)(103));
FA_ff_743:FAff port map(x=>p(15)(103),y=>p(16)(103),Cin=>p(17)(103),clock=>clock,reset=>reset,s=>p(138)(103),cout=>p(139)(104));
FA_ff_744:FAff port map(x=>p(15)(104),y=>p(16)(104),Cin=>p(17)(104),clock=>clock,reset=>reset,s=>p(138)(104),cout=>p(139)(105));
FA_ff_745:FAff port map(x=>p(15)(105),y=>p(16)(105),Cin=>p(17)(105),clock=>clock,reset=>reset,s=>p(138)(105),cout=>p(139)(106));
FA_ff_746:FAff port map(x=>p(15)(106),y=>p(16)(106),Cin=>p(17)(106),clock=>clock,reset=>reset,s=>p(138)(106),cout=>p(139)(107));
FA_ff_747:FAff port map(x=>p(15)(107),y=>p(16)(107),Cin=>p(17)(107),clock=>clock,reset=>reset,s=>p(138)(107),cout=>p(139)(108));
FA_ff_748:FAff port map(x=>p(15)(108),y=>p(16)(108),Cin=>p(17)(108),clock=>clock,reset=>reset,s=>p(138)(108),cout=>p(139)(109));
FA_ff_749:FAff port map(x=>p(15)(109),y=>p(16)(109),Cin=>p(17)(109),clock=>clock,reset=>reset,s=>p(138)(109),cout=>p(139)(110));
FA_ff_750:FAff port map(x=>p(15)(110),y=>p(16)(110),Cin=>p(17)(110),clock=>clock,reset=>reset,s=>p(138)(110),cout=>p(139)(111));
FA_ff_751:FAff port map(x=>p(15)(111),y=>p(16)(111),Cin=>p(17)(111),clock=>clock,reset=>reset,s=>p(138)(111),cout=>p(139)(112));
FA_ff_752:FAff port map(x=>p(15)(112),y=>p(16)(112),Cin=>p(17)(112),clock=>clock,reset=>reset,s=>p(138)(112),cout=>p(139)(113));
FA_ff_753:FAff port map(x=>p(15)(113),y=>p(16)(113),Cin=>p(17)(113),clock=>clock,reset=>reset,s=>p(138)(113),cout=>p(139)(114));
FA_ff_754:FAff port map(x=>p(15)(114),y=>p(16)(114),Cin=>p(17)(114),clock=>clock,reset=>reset,s=>p(138)(114),cout=>p(139)(115));
FA_ff_755:FAff port map(x=>p(15)(115),y=>p(16)(115),Cin=>p(17)(115),clock=>clock,reset=>reset,s=>p(138)(115),cout=>p(139)(116));
FA_ff_756:FAff port map(x=>p(15)(116),y=>p(16)(116),Cin=>p(17)(116),clock=>clock,reset=>reset,s=>p(138)(116),cout=>p(139)(117));
FA_ff_757:FAff port map(x=>p(15)(117),y=>p(16)(117),Cin=>p(17)(117),clock=>clock,reset=>reset,s=>p(138)(117),cout=>p(139)(118));
FA_ff_758:FAff port map(x=>p(15)(118),y=>p(16)(118),Cin=>p(17)(118),clock=>clock,reset=>reset,s=>p(138)(118),cout=>p(139)(119));
FA_ff_759:FAff port map(x=>p(15)(119),y=>p(16)(119),Cin=>p(17)(119),clock=>clock,reset=>reset,s=>p(138)(119),cout=>p(139)(120));
FA_ff_760:FAff port map(x=>p(15)(120),y=>p(16)(120),Cin=>p(17)(120),clock=>clock,reset=>reset,s=>p(138)(120),cout=>p(139)(121));
FA_ff_761:FAff port map(x=>p(15)(121),y=>p(16)(121),Cin=>p(17)(121),clock=>clock,reset=>reset,s=>p(138)(121),cout=>p(139)(122));
FA_ff_762:FAff port map(x=>p(15)(122),y=>p(16)(122),Cin=>p(17)(122),clock=>clock,reset=>reset,s=>p(138)(122),cout=>p(139)(123));
FA_ff_763:FAff port map(x=>p(15)(123),y=>p(16)(123),Cin=>p(17)(123),clock=>clock,reset=>reset,s=>p(138)(123),cout=>p(139)(124));
FA_ff_764:FAff port map(x=>p(15)(124),y=>p(16)(124),Cin=>p(17)(124),clock=>clock,reset=>reset,s=>p(138)(124),cout=>p(139)(125));
FA_ff_765:FAff port map(x=>p(15)(125),y=>p(16)(125),Cin=>p(17)(125),clock=>clock,reset=>reset,s=>p(138)(125),cout=>p(139)(126));
FA_ff_766:FAff port map(x=>p(15)(126),y=>p(16)(126),Cin=>p(17)(126),clock=>clock,reset=>reset,s=>p(138)(126),cout=>p(139)(127));
FA_ff_767:FAff port map(x=>p(15)(127),y=>p(16)(127),Cin=>p(17)(127),clock=>clock,reset=>reset,s=>p(138)(127),cout=>p(139)(128));
FA_ff_768:FAff port map(x=>p(18)(0),y=>p(19)(0),Cin=>p(20)(0),clock=>clock,reset=>reset,s=>p(140)(0),cout=>p(141)(1));
FA_ff_769:FAff port map(x=>p(18)(1),y=>p(19)(1),Cin=>p(20)(1),clock=>clock,reset=>reset,s=>p(140)(1),cout=>p(141)(2));
FA_ff_770:FAff port map(x=>p(18)(2),y=>p(19)(2),Cin=>p(20)(2),clock=>clock,reset=>reset,s=>p(140)(2),cout=>p(141)(3));
FA_ff_771:FAff port map(x=>p(18)(3),y=>p(19)(3),Cin=>p(20)(3),clock=>clock,reset=>reset,s=>p(140)(3),cout=>p(141)(4));
FA_ff_772:FAff port map(x=>p(18)(4),y=>p(19)(4),Cin=>p(20)(4),clock=>clock,reset=>reset,s=>p(140)(4),cout=>p(141)(5));
FA_ff_773:FAff port map(x=>p(18)(5),y=>p(19)(5),Cin=>p(20)(5),clock=>clock,reset=>reset,s=>p(140)(5),cout=>p(141)(6));
FA_ff_774:FAff port map(x=>p(18)(6),y=>p(19)(6),Cin=>p(20)(6),clock=>clock,reset=>reset,s=>p(140)(6),cout=>p(141)(7));
FA_ff_775:FAff port map(x=>p(18)(7),y=>p(19)(7),Cin=>p(20)(7),clock=>clock,reset=>reset,s=>p(140)(7),cout=>p(141)(8));
FA_ff_776:FAff port map(x=>p(18)(8),y=>p(19)(8),Cin=>p(20)(8),clock=>clock,reset=>reset,s=>p(140)(8),cout=>p(141)(9));
FA_ff_777:FAff port map(x=>p(18)(9),y=>p(19)(9),Cin=>p(20)(9),clock=>clock,reset=>reset,s=>p(140)(9),cout=>p(141)(10));
FA_ff_778:FAff port map(x=>p(18)(10),y=>p(19)(10),Cin=>p(20)(10),clock=>clock,reset=>reset,s=>p(140)(10),cout=>p(141)(11));
FA_ff_779:FAff port map(x=>p(18)(11),y=>p(19)(11),Cin=>p(20)(11),clock=>clock,reset=>reset,s=>p(140)(11),cout=>p(141)(12));
FA_ff_780:FAff port map(x=>p(18)(12),y=>p(19)(12),Cin=>p(20)(12),clock=>clock,reset=>reset,s=>p(140)(12),cout=>p(141)(13));
FA_ff_781:FAff port map(x=>p(18)(13),y=>p(19)(13),Cin=>p(20)(13),clock=>clock,reset=>reset,s=>p(140)(13),cout=>p(141)(14));
FA_ff_782:FAff port map(x=>p(18)(14),y=>p(19)(14),Cin=>p(20)(14),clock=>clock,reset=>reset,s=>p(140)(14),cout=>p(141)(15));
FA_ff_783:FAff port map(x=>p(18)(15),y=>p(19)(15),Cin=>p(20)(15),clock=>clock,reset=>reset,s=>p(140)(15),cout=>p(141)(16));
FA_ff_784:FAff port map(x=>p(18)(16),y=>p(19)(16),Cin=>p(20)(16),clock=>clock,reset=>reset,s=>p(140)(16),cout=>p(141)(17));
FA_ff_785:FAff port map(x=>p(18)(17),y=>p(19)(17),Cin=>p(20)(17),clock=>clock,reset=>reset,s=>p(140)(17),cout=>p(141)(18));
FA_ff_786:FAff port map(x=>p(18)(18),y=>p(19)(18),Cin=>p(20)(18),clock=>clock,reset=>reset,s=>p(140)(18),cout=>p(141)(19));
FA_ff_787:FAff port map(x=>p(18)(19),y=>p(19)(19),Cin=>p(20)(19),clock=>clock,reset=>reset,s=>p(140)(19),cout=>p(141)(20));
FA_ff_788:FAff port map(x=>p(18)(20),y=>p(19)(20),Cin=>p(20)(20),clock=>clock,reset=>reset,s=>p(140)(20),cout=>p(141)(21));
FA_ff_789:FAff port map(x=>p(18)(21),y=>p(19)(21),Cin=>p(20)(21),clock=>clock,reset=>reset,s=>p(140)(21),cout=>p(141)(22));
FA_ff_790:FAff port map(x=>p(18)(22),y=>p(19)(22),Cin=>p(20)(22),clock=>clock,reset=>reset,s=>p(140)(22),cout=>p(141)(23));
FA_ff_791:FAff port map(x=>p(18)(23),y=>p(19)(23),Cin=>p(20)(23),clock=>clock,reset=>reset,s=>p(140)(23),cout=>p(141)(24));
FA_ff_792:FAff port map(x=>p(18)(24),y=>p(19)(24),Cin=>p(20)(24),clock=>clock,reset=>reset,s=>p(140)(24),cout=>p(141)(25));
FA_ff_793:FAff port map(x=>p(18)(25),y=>p(19)(25),Cin=>p(20)(25),clock=>clock,reset=>reset,s=>p(140)(25),cout=>p(141)(26));
FA_ff_794:FAff port map(x=>p(18)(26),y=>p(19)(26),Cin=>p(20)(26),clock=>clock,reset=>reset,s=>p(140)(26),cout=>p(141)(27));
FA_ff_795:FAff port map(x=>p(18)(27),y=>p(19)(27),Cin=>p(20)(27),clock=>clock,reset=>reset,s=>p(140)(27),cout=>p(141)(28));
FA_ff_796:FAff port map(x=>p(18)(28),y=>p(19)(28),Cin=>p(20)(28),clock=>clock,reset=>reset,s=>p(140)(28),cout=>p(141)(29));
FA_ff_797:FAff port map(x=>p(18)(29),y=>p(19)(29),Cin=>p(20)(29),clock=>clock,reset=>reset,s=>p(140)(29),cout=>p(141)(30));
FA_ff_798:FAff port map(x=>p(18)(30),y=>p(19)(30),Cin=>p(20)(30),clock=>clock,reset=>reset,s=>p(140)(30),cout=>p(141)(31));
FA_ff_799:FAff port map(x=>p(18)(31),y=>p(19)(31),Cin=>p(20)(31),clock=>clock,reset=>reset,s=>p(140)(31),cout=>p(141)(32));
FA_ff_800:FAff port map(x=>p(18)(32),y=>p(19)(32),Cin=>p(20)(32),clock=>clock,reset=>reset,s=>p(140)(32),cout=>p(141)(33));
FA_ff_801:FAff port map(x=>p(18)(33),y=>p(19)(33),Cin=>p(20)(33),clock=>clock,reset=>reset,s=>p(140)(33),cout=>p(141)(34));
FA_ff_802:FAff port map(x=>p(18)(34),y=>p(19)(34),Cin=>p(20)(34),clock=>clock,reset=>reset,s=>p(140)(34),cout=>p(141)(35));
FA_ff_803:FAff port map(x=>p(18)(35),y=>p(19)(35),Cin=>p(20)(35),clock=>clock,reset=>reset,s=>p(140)(35),cout=>p(141)(36));
FA_ff_804:FAff port map(x=>p(18)(36),y=>p(19)(36),Cin=>p(20)(36),clock=>clock,reset=>reset,s=>p(140)(36),cout=>p(141)(37));
FA_ff_805:FAff port map(x=>p(18)(37),y=>p(19)(37),Cin=>p(20)(37),clock=>clock,reset=>reset,s=>p(140)(37),cout=>p(141)(38));
FA_ff_806:FAff port map(x=>p(18)(38),y=>p(19)(38),Cin=>p(20)(38),clock=>clock,reset=>reset,s=>p(140)(38),cout=>p(141)(39));
FA_ff_807:FAff port map(x=>p(18)(39),y=>p(19)(39),Cin=>p(20)(39),clock=>clock,reset=>reset,s=>p(140)(39),cout=>p(141)(40));
FA_ff_808:FAff port map(x=>p(18)(40),y=>p(19)(40),Cin=>p(20)(40),clock=>clock,reset=>reset,s=>p(140)(40),cout=>p(141)(41));
FA_ff_809:FAff port map(x=>p(18)(41),y=>p(19)(41),Cin=>p(20)(41),clock=>clock,reset=>reset,s=>p(140)(41),cout=>p(141)(42));
FA_ff_810:FAff port map(x=>p(18)(42),y=>p(19)(42),Cin=>p(20)(42),clock=>clock,reset=>reset,s=>p(140)(42),cout=>p(141)(43));
FA_ff_811:FAff port map(x=>p(18)(43),y=>p(19)(43),Cin=>p(20)(43),clock=>clock,reset=>reset,s=>p(140)(43),cout=>p(141)(44));
FA_ff_812:FAff port map(x=>p(18)(44),y=>p(19)(44),Cin=>p(20)(44),clock=>clock,reset=>reset,s=>p(140)(44),cout=>p(141)(45));
FA_ff_813:FAff port map(x=>p(18)(45),y=>p(19)(45),Cin=>p(20)(45),clock=>clock,reset=>reset,s=>p(140)(45),cout=>p(141)(46));
FA_ff_814:FAff port map(x=>p(18)(46),y=>p(19)(46),Cin=>p(20)(46),clock=>clock,reset=>reset,s=>p(140)(46),cout=>p(141)(47));
FA_ff_815:FAff port map(x=>p(18)(47),y=>p(19)(47),Cin=>p(20)(47),clock=>clock,reset=>reset,s=>p(140)(47),cout=>p(141)(48));
FA_ff_816:FAff port map(x=>p(18)(48),y=>p(19)(48),Cin=>p(20)(48),clock=>clock,reset=>reset,s=>p(140)(48),cout=>p(141)(49));
FA_ff_817:FAff port map(x=>p(18)(49),y=>p(19)(49),Cin=>p(20)(49),clock=>clock,reset=>reset,s=>p(140)(49),cout=>p(141)(50));
FA_ff_818:FAff port map(x=>p(18)(50),y=>p(19)(50),Cin=>p(20)(50),clock=>clock,reset=>reset,s=>p(140)(50),cout=>p(141)(51));
FA_ff_819:FAff port map(x=>p(18)(51),y=>p(19)(51),Cin=>p(20)(51),clock=>clock,reset=>reset,s=>p(140)(51),cout=>p(141)(52));
FA_ff_820:FAff port map(x=>p(18)(52),y=>p(19)(52),Cin=>p(20)(52),clock=>clock,reset=>reset,s=>p(140)(52),cout=>p(141)(53));
FA_ff_821:FAff port map(x=>p(18)(53),y=>p(19)(53),Cin=>p(20)(53),clock=>clock,reset=>reset,s=>p(140)(53),cout=>p(141)(54));
FA_ff_822:FAff port map(x=>p(18)(54),y=>p(19)(54),Cin=>p(20)(54),clock=>clock,reset=>reset,s=>p(140)(54),cout=>p(141)(55));
FA_ff_823:FAff port map(x=>p(18)(55),y=>p(19)(55),Cin=>p(20)(55),clock=>clock,reset=>reset,s=>p(140)(55),cout=>p(141)(56));
FA_ff_824:FAff port map(x=>p(18)(56),y=>p(19)(56),Cin=>p(20)(56),clock=>clock,reset=>reset,s=>p(140)(56),cout=>p(141)(57));
FA_ff_825:FAff port map(x=>p(18)(57),y=>p(19)(57),Cin=>p(20)(57),clock=>clock,reset=>reset,s=>p(140)(57),cout=>p(141)(58));
FA_ff_826:FAff port map(x=>p(18)(58),y=>p(19)(58),Cin=>p(20)(58),clock=>clock,reset=>reset,s=>p(140)(58),cout=>p(141)(59));
FA_ff_827:FAff port map(x=>p(18)(59),y=>p(19)(59),Cin=>p(20)(59),clock=>clock,reset=>reset,s=>p(140)(59),cout=>p(141)(60));
FA_ff_828:FAff port map(x=>p(18)(60),y=>p(19)(60),Cin=>p(20)(60),clock=>clock,reset=>reset,s=>p(140)(60),cout=>p(141)(61));
FA_ff_829:FAff port map(x=>p(18)(61),y=>p(19)(61),Cin=>p(20)(61),clock=>clock,reset=>reset,s=>p(140)(61),cout=>p(141)(62));
FA_ff_830:FAff port map(x=>p(18)(62),y=>p(19)(62),Cin=>p(20)(62),clock=>clock,reset=>reset,s=>p(140)(62),cout=>p(141)(63));
FA_ff_831:FAff port map(x=>p(18)(63),y=>p(19)(63),Cin=>p(20)(63),clock=>clock,reset=>reset,s=>p(140)(63),cout=>p(141)(64));
FA_ff_832:FAff port map(x=>p(18)(64),y=>p(19)(64),Cin=>p(20)(64),clock=>clock,reset=>reset,s=>p(140)(64),cout=>p(141)(65));
FA_ff_833:FAff port map(x=>p(18)(65),y=>p(19)(65),Cin=>p(20)(65),clock=>clock,reset=>reset,s=>p(140)(65),cout=>p(141)(66));
FA_ff_834:FAff port map(x=>p(18)(66),y=>p(19)(66),Cin=>p(20)(66),clock=>clock,reset=>reset,s=>p(140)(66),cout=>p(141)(67));
FA_ff_835:FAff port map(x=>p(18)(67),y=>p(19)(67),Cin=>p(20)(67),clock=>clock,reset=>reset,s=>p(140)(67),cout=>p(141)(68));
FA_ff_836:FAff port map(x=>p(18)(68),y=>p(19)(68),Cin=>p(20)(68),clock=>clock,reset=>reset,s=>p(140)(68),cout=>p(141)(69));
FA_ff_837:FAff port map(x=>p(18)(69),y=>p(19)(69),Cin=>p(20)(69),clock=>clock,reset=>reset,s=>p(140)(69),cout=>p(141)(70));
FA_ff_838:FAff port map(x=>p(18)(70),y=>p(19)(70),Cin=>p(20)(70),clock=>clock,reset=>reset,s=>p(140)(70),cout=>p(141)(71));
FA_ff_839:FAff port map(x=>p(18)(71),y=>p(19)(71),Cin=>p(20)(71),clock=>clock,reset=>reset,s=>p(140)(71),cout=>p(141)(72));
FA_ff_840:FAff port map(x=>p(18)(72),y=>p(19)(72),Cin=>p(20)(72),clock=>clock,reset=>reset,s=>p(140)(72),cout=>p(141)(73));
FA_ff_841:FAff port map(x=>p(18)(73),y=>p(19)(73),Cin=>p(20)(73),clock=>clock,reset=>reset,s=>p(140)(73),cout=>p(141)(74));
FA_ff_842:FAff port map(x=>p(18)(74),y=>p(19)(74),Cin=>p(20)(74),clock=>clock,reset=>reset,s=>p(140)(74),cout=>p(141)(75));
FA_ff_843:FAff port map(x=>p(18)(75),y=>p(19)(75),Cin=>p(20)(75),clock=>clock,reset=>reset,s=>p(140)(75),cout=>p(141)(76));
FA_ff_844:FAff port map(x=>p(18)(76),y=>p(19)(76),Cin=>p(20)(76),clock=>clock,reset=>reset,s=>p(140)(76),cout=>p(141)(77));
FA_ff_845:FAff port map(x=>p(18)(77),y=>p(19)(77),Cin=>p(20)(77),clock=>clock,reset=>reset,s=>p(140)(77),cout=>p(141)(78));
FA_ff_846:FAff port map(x=>p(18)(78),y=>p(19)(78),Cin=>p(20)(78),clock=>clock,reset=>reset,s=>p(140)(78),cout=>p(141)(79));
FA_ff_847:FAff port map(x=>p(18)(79),y=>p(19)(79),Cin=>p(20)(79),clock=>clock,reset=>reset,s=>p(140)(79),cout=>p(141)(80));
FA_ff_848:FAff port map(x=>p(18)(80),y=>p(19)(80),Cin=>p(20)(80),clock=>clock,reset=>reset,s=>p(140)(80),cout=>p(141)(81));
FA_ff_849:FAff port map(x=>p(18)(81),y=>p(19)(81),Cin=>p(20)(81),clock=>clock,reset=>reset,s=>p(140)(81),cout=>p(141)(82));
FA_ff_850:FAff port map(x=>p(18)(82),y=>p(19)(82),Cin=>p(20)(82),clock=>clock,reset=>reset,s=>p(140)(82),cout=>p(141)(83));
FA_ff_851:FAff port map(x=>p(18)(83),y=>p(19)(83),Cin=>p(20)(83),clock=>clock,reset=>reset,s=>p(140)(83),cout=>p(141)(84));
FA_ff_852:FAff port map(x=>p(18)(84),y=>p(19)(84),Cin=>p(20)(84),clock=>clock,reset=>reset,s=>p(140)(84),cout=>p(141)(85));
FA_ff_853:FAff port map(x=>p(18)(85),y=>p(19)(85),Cin=>p(20)(85),clock=>clock,reset=>reset,s=>p(140)(85),cout=>p(141)(86));
FA_ff_854:FAff port map(x=>p(18)(86),y=>p(19)(86),Cin=>p(20)(86),clock=>clock,reset=>reset,s=>p(140)(86),cout=>p(141)(87));
FA_ff_855:FAff port map(x=>p(18)(87),y=>p(19)(87),Cin=>p(20)(87),clock=>clock,reset=>reset,s=>p(140)(87),cout=>p(141)(88));
FA_ff_856:FAff port map(x=>p(18)(88),y=>p(19)(88),Cin=>p(20)(88),clock=>clock,reset=>reset,s=>p(140)(88),cout=>p(141)(89));
FA_ff_857:FAff port map(x=>p(18)(89),y=>p(19)(89),Cin=>p(20)(89),clock=>clock,reset=>reset,s=>p(140)(89),cout=>p(141)(90));
FA_ff_858:FAff port map(x=>p(18)(90),y=>p(19)(90),Cin=>p(20)(90),clock=>clock,reset=>reset,s=>p(140)(90),cout=>p(141)(91));
FA_ff_859:FAff port map(x=>p(18)(91),y=>p(19)(91),Cin=>p(20)(91),clock=>clock,reset=>reset,s=>p(140)(91),cout=>p(141)(92));
FA_ff_860:FAff port map(x=>p(18)(92),y=>p(19)(92),Cin=>p(20)(92),clock=>clock,reset=>reset,s=>p(140)(92),cout=>p(141)(93));
FA_ff_861:FAff port map(x=>p(18)(93),y=>p(19)(93),Cin=>p(20)(93),clock=>clock,reset=>reset,s=>p(140)(93),cout=>p(141)(94));
FA_ff_862:FAff port map(x=>p(18)(94),y=>p(19)(94),Cin=>p(20)(94),clock=>clock,reset=>reset,s=>p(140)(94),cout=>p(141)(95));
FA_ff_863:FAff port map(x=>p(18)(95),y=>p(19)(95),Cin=>p(20)(95),clock=>clock,reset=>reset,s=>p(140)(95),cout=>p(141)(96));
FA_ff_864:FAff port map(x=>p(18)(96),y=>p(19)(96),Cin=>p(20)(96),clock=>clock,reset=>reset,s=>p(140)(96),cout=>p(141)(97));
FA_ff_865:FAff port map(x=>p(18)(97),y=>p(19)(97),Cin=>p(20)(97),clock=>clock,reset=>reset,s=>p(140)(97),cout=>p(141)(98));
FA_ff_866:FAff port map(x=>p(18)(98),y=>p(19)(98),Cin=>p(20)(98),clock=>clock,reset=>reset,s=>p(140)(98),cout=>p(141)(99));
FA_ff_867:FAff port map(x=>p(18)(99),y=>p(19)(99),Cin=>p(20)(99),clock=>clock,reset=>reset,s=>p(140)(99),cout=>p(141)(100));
FA_ff_868:FAff port map(x=>p(18)(100),y=>p(19)(100),Cin=>p(20)(100),clock=>clock,reset=>reset,s=>p(140)(100),cout=>p(141)(101));
FA_ff_869:FAff port map(x=>p(18)(101),y=>p(19)(101),Cin=>p(20)(101),clock=>clock,reset=>reset,s=>p(140)(101),cout=>p(141)(102));
FA_ff_870:FAff port map(x=>p(18)(102),y=>p(19)(102),Cin=>p(20)(102),clock=>clock,reset=>reset,s=>p(140)(102),cout=>p(141)(103));
FA_ff_871:FAff port map(x=>p(18)(103),y=>p(19)(103),Cin=>p(20)(103),clock=>clock,reset=>reset,s=>p(140)(103),cout=>p(141)(104));
FA_ff_872:FAff port map(x=>p(18)(104),y=>p(19)(104),Cin=>p(20)(104),clock=>clock,reset=>reset,s=>p(140)(104),cout=>p(141)(105));
FA_ff_873:FAff port map(x=>p(18)(105),y=>p(19)(105),Cin=>p(20)(105),clock=>clock,reset=>reset,s=>p(140)(105),cout=>p(141)(106));
FA_ff_874:FAff port map(x=>p(18)(106),y=>p(19)(106),Cin=>p(20)(106),clock=>clock,reset=>reset,s=>p(140)(106),cout=>p(141)(107));
FA_ff_875:FAff port map(x=>p(18)(107),y=>p(19)(107),Cin=>p(20)(107),clock=>clock,reset=>reset,s=>p(140)(107),cout=>p(141)(108));
FA_ff_876:FAff port map(x=>p(18)(108),y=>p(19)(108),Cin=>p(20)(108),clock=>clock,reset=>reset,s=>p(140)(108),cout=>p(141)(109));
FA_ff_877:FAff port map(x=>p(18)(109),y=>p(19)(109),Cin=>p(20)(109),clock=>clock,reset=>reset,s=>p(140)(109),cout=>p(141)(110));
FA_ff_878:FAff port map(x=>p(18)(110),y=>p(19)(110),Cin=>p(20)(110),clock=>clock,reset=>reset,s=>p(140)(110),cout=>p(141)(111));
FA_ff_879:FAff port map(x=>p(18)(111),y=>p(19)(111),Cin=>p(20)(111),clock=>clock,reset=>reset,s=>p(140)(111),cout=>p(141)(112));
FA_ff_880:FAff port map(x=>p(18)(112),y=>p(19)(112),Cin=>p(20)(112),clock=>clock,reset=>reset,s=>p(140)(112),cout=>p(141)(113));
FA_ff_881:FAff port map(x=>p(18)(113),y=>p(19)(113),Cin=>p(20)(113),clock=>clock,reset=>reset,s=>p(140)(113),cout=>p(141)(114));
FA_ff_882:FAff port map(x=>p(18)(114),y=>p(19)(114),Cin=>p(20)(114),clock=>clock,reset=>reset,s=>p(140)(114),cout=>p(141)(115));
FA_ff_883:FAff port map(x=>p(18)(115),y=>p(19)(115),Cin=>p(20)(115),clock=>clock,reset=>reset,s=>p(140)(115),cout=>p(141)(116));
FA_ff_884:FAff port map(x=>p(18)(116),y=>p(19)(116),Cin=>p(20)(116),clock=>clock,reset=>reset,s=>p(140)(116),cout=>p(141)(117));
FA_ff_885:FAff port map(x=>p(18)(117),y=>p(19)(117),Cin=>p(20)(117),clock=>clock,reset=>reset,s=>p(140)(117),cout=>p(141)(118));
FA_ff_886:FAff port map(x=>p(18)(118),y=>p(19)(118),Cin=>p(20)(118),clock=>clock,reset=>reset,s=>p(140)(118),cout=>p(141)(119));
FA_ff_887:FAff port map(x=>p(18)(119),y=>p(19)(119),Cin=>p(20)(119),clock=>clock,reset=>reset,s=>p(140)(119),cout=>p(141)(120));
FA_ff_888:FAff port map(x=>p(18)(120),y=>p(19)(120),Cin=>p(20)(120),clock=>clock,reset=>reset,s=>p(140)(120),cout=>p(141)(121));
FA_ff_889:FAff port map(x=>p(18)(121),y=>p(19)(121),Cin=>p(20)(121),clock=>clock,reset=>reset,s=>p(140)(121),cout=>p(141)(122));
FA_ff_890:FAff port map(x=>p(18)(122),y=>p(19)(122),Cin=>p(20)(122),clock=>clock,reset=>reset,s=>p(140)(122),cout=>p(141)(123));
FA_ff_891:FAff port map(x=>p(18)(123),y=>p(19)(123),Cin=>p(20)(123),clock=>clock,reset=>reset,s=>p(140)(123),cout=>p(141)(124));
FA_ff_892:FAff port map(x=>p(18)(124),y=>p(19)(124),Cin=>p(20)(124),clock=>clock,reset=>reset,s=>p(140)(124),cout=>p(141)(125));
FA_ff_893:FAff port map(x=>p(18)(125),y=>p(19)(125),Cin=>p(20)(125),clock=>clock,reset=>reset,s=>p(140)(125),cout=>p(141)(126));
FA_ff_894:FAff port map(x=>p(18)(126),y=>p(19)(126),Cin=>p(20)(126),clock=>clock,reset=>reset,s=>p(140)(126),cout=>p(141)(127));
FA_ff_895:FAff port map(x=>p(18)(127),y=>p(19)(127),Cin=>p(20)(127),clock=>clock,reset=>reset,s=>p(140)(127),cout=>p(141)(128));
FA_ff_896:FAff port map(x=>p(21)(0),y=>p(22)(0),Cin=>p(23)(0),clock=>clock,reset=>reset,s=>p(142)(0),cout=>p(143)(1));
FA_ff_897:FAff port map(x=>p(21)(1),y=>p(22)(1),Cin=>p(23)(1),clock=>clock,reset=>reset,s=>p(142)(1),cout=>p(143)(2));
FA_ff_898:FAff port map(x=>p(21)(2),y=>p(22)(2),Cin=>p(23)(2),clock=>clock,reset=>reset,s=>p(142)(2),cout=>p(143)(3));
FA_ff_899:FAff port map(x=>p(21)(3),y=>p(22)(3),Cin=>p(23)(3),clock=>clock,reset=>reset,s=>p(142)(3),cout=>p(143)(4));
FA_ff_900:FAff port map(x=>p(21)(4),y=>p(22)(4),Cin=>p(23)(4),clock=>clock,reset=>reset,s=>p(142)(4),cout=>p(143)(5));
FA_ff_901:FAff port map(x=>p(21)(5),y=>p(22)(5),Cin=>p(23)(5),clock=>clock,reset=>reset,s=>p(142)(5),cout=>p(143)(6));
FA_ff_902:FAff port map(x=>p(21)(6),y=>p(22)(6),Cin=>p(23)(6),clock=>clock,reset=>reset,s=>p(142)(6),cout=>p(143)(7));
FA_ff_903:FAff port map(x=>p(21)(7),y=>p(22)(7),Cin=>p(23)(7),clock=>clock,reset=>reset,s=>p(142)(7),cout=>p(143)(8));
FA_ff_904:FAff port map(x=>p(21)(8),y=>p(22)(8),Cin=>p(23)(8),clock=>clock,reset=>reset,s=>p(142)(8),cout=>p(143)(9));
FA_ff_905:FAff port map(x=>p(21)(9),y=>p(22)(9),Cin=>p(23)(9),clock=>clock,reset=>reset,s=>p(142)(9),cout=>p(143)(10));
FA_ff_906:FAff port map(x=>p(21)(10),y=>p(22)(10),Cin=>p(23)(10),clock=>clock,reset=>reset,s=>p(142)(10),cout=>p(143)(11));
FA_ff_907:FAff port map(x=>p(21)(11),y=>p(22)(11),Cin=>p(23)(11),clock=>clock,reset=>reset,s=>p(142)(11),cout=>p(143)(12));
FA_ff_908:FAff port map(x=>p(21)(12),y=>p(22)(12),Cin=>p(23)(12),clock=>clock,reset=>reset,s=>p(142)(12),cout=>p(143)(13));
FA_ff_909:FAff port map(x=>p(21)(13),y=>p(22)(13),Cin=>p(23)(13),clock=>clock,reset=>reset,s=>p(142)(13),cout=>p(143)(14));
FA_ff_910:FAff port map(x=>p(21)(14),y=>p(22)(14),Cin=>p(23)(14),clock=>clock,reset=>reset,s=>p(142)(14),cout=>p(143)(15));
FA_ff_911:FAff port map(x=>p(21)(15),y=>p(22)(15),Cin=>p(23)(15),clock=>clock,reset=>reset,s=>p(142)(15),cout=>p(143)(16));
FA_ff_912:FAff port map(x=>p(21)(16),y=>p(22)(16),Cin=>p(23)(16),clock=>clock,reset=>reset,s=>p(142)(16),cout=>p(143)(17));
FA_ff_913:FAff port map(x=>p(21)(17),y=>p(22)(17),Cin=>p(23)(17),clock=>clock,reset=>reset,s=>p(142)(17),cout=>p(143)(18));
FA_ff_914:FAff port map(x=>p(21)(18),y=>p(22)(18),Cin=>p(23)(18),clock=>clock,reset=>reset,s=>p(142)(18),cout=>p(143)(19));
FA_ff_915:FAff port map(x=>p(21)(19),y=>p(22)(19),Cin=>p(23)(19),clock=>clock,reset=>reset,s=>p(142)(19),cout=>p(143)(20));
FA_ff_916:FAff port map(x=>p(21)(20),y=>p(22)(20),Cin=>p(23)(20),clock=>clock,reset=>reset,s=>p(142)(20),cout=>p(143)(21));
FA_ff_917:FAff port map(x=>p(21)(21),y=>p(22)(21),Cin=>p(23)(21),clock=>clock,reset=>reset,s=>p(142)(21),cout=>p(143)(22));
FA_ff_918:FAff port map(x=>p(21)(22),y=>p(22)(22),Cin=>p(23)(22),clock=>clock,reset=>reset,s=>p(142)(22),cout=>p(143)(23));
FA_ff_919:FAff port map(x=>p(21)(23),y=>p(22)(23),Cin=>p(23)(23),clock=>clock,reset=>reset,s=>p(142)(23),cout=>p(143)(24));
FA_ff_920:FAff port map(x=>p(21)(24),y=>p(22)(24),Cin=>p(23)(24),clock=>clock,reset=>reset,s=>p(142)(24),cout=>p(143)(25));
FA_ff_921:FAff port map(x=>p(21)(25),y=>p(22)(25),Cin=>p(23)(25),clock=>clock,reset=>reset,s=>p(142)(25),cout=>p(143)(26));
FA_ff_922:FAff port map(x=>p(21)(26),y=>p(22)(26),Cin=>p(23)(26),clock=>clock,reset=>reset,s=>p(142)(26),cout=>p(143)(27));
FA_ff_923:FAff port map(x=>p(21)(27),y=>p(22)(27),Cin=>p(23)(27),clock=>clock,reset=>reset,s=>p(142)(27),cout=>p(143)(28));
FA_ff_924:FAff port map(x=>p(21)(28),y=>p(22)(28),Cin=>p(23)(28),clock=>clock,reset=>reset,s=>p(142)(28),cout=>p(143)(29));
FA_ff_925:FAff port map(x=>p(21)(29),y=>p(22)(29),Cin=>p(23)(29),clock=>clock,reset=>reset,s=>p(142)(29),cout=>p(143)(30));
FA_ff_926:FAff port map(x=>p(21)(30),y=>p(22)(30),Cin=>p(23)(30),clock=>clock,reset=>reset,s=>p(142)(30),cout=>p(143)(31));
FA_ff_927:FAff port map(x=>p(21)(31),y=>p(22)(31),Cin=>p(23)(31),clock=>clock,reset=>reset,s=>p(142)(31),cout=>p(143)(32));
FA_ff_928:FAff port map(x=>p(21)(32),y=>p(22)(32),Cin=>p(23)(32),clock=>clock,reset=>reset,s=>p(142)(32),cout=>p(143)(33));
FA_ff_929:FAff port map(x=>p(21)(33),y=>p(22)(33),Cin=>p(23)(33),clock=>clock,reset=>reset,s=>p(142)(33),cout=>p(143)(34));
FA_ff_930:FAff port map(x=>p(21)(34),y=>p(22)(34),Cin=>p(23)(34),clock=>clock,reset=>reset,s=>p(142)(34),cout=>p(143)(35));
FA_ff_931:FAff port map(x=>p(21)(35),y=>p(22)(35),Cin=>p(23)(35),clock=>clock,reset=>reset,s=>p(142)(35),cout=>p(143)(36));
FA_ff_932:FAff port map(x=>p(21)(36),y=>p(22)(36),Cin=>p(23)(36),clock=>clock,reset=>reset,s=>p(142)(36),cout=>p(143)(37));
FA_ff_933:FAff port map(x=>p(21)(37),y=>p(22)(37),Cin=>p(23)(37),clock=>clock,reset=>reset,s=>p(142)(37),cout=>p(143)(38));
FA_ff_934:FAff port map(x=>p(21)(38),y=>p(22)(38),Cin=>p(23)(38),clock=>clock,reset=>reset,s=>p(142)(38),cout=>p(143)(39));
FA_ff_935:FAff port map(x=>p(21)(39),y=>p(22)(39),Cin=>p(23)(39),clock=>clock,reset=>reset,s=>p(142)(39),cout=>p(143)(40));
FA_ff_936:FAff port map(x=>p(21)(40),y=>p(22)(40),Cin=>p(23)(40),clock=>clock,reset=>reset,s=>p(142)(40),cout=>p(143)(41));
FA_ff_937:FAff port map(x=>p(21)(41),y=>p(22)(41),Cin=>p(23)(41),clock=>clock,reset=>reset,s=>p(142)(41),cout=>p(143)(42));
FA_ff_938:FAff port map(x=>p(21)(42),y=>p(22)(42),Cin=>p(23)(42),clock=>clock,reset=>reset,s=>p(142)(42),cout=>p(143)(43));
FA_ff_939:FAff port map(x=>p(21)(43),y=>p(22)(43),Cin=>p(23)(43),clock=>clock,reset=>reset,s=>p(142)(43),cout=>p(143)(44));
FA_ff_940:FAff port map(x=>p(21)(44),y=>p(22)(44),Cin=>p(23)(44),clock=>clock,reset=>reset,s=>p(142)(44),cout=>p(143)(45));
FA_ff_941:FAff port map(x=>p(21)(45),y=>p(22)(45),Cin=>p(23)(45),clock=>clock,reset=>reset,s=>p(142)(45),cout=>p(143)(46));
FA_ff_942:FAff port map(x=>p(21)(46),y=>p(22)(46),Cin=>p(23)(46),clock=>clock,reset=>reset,s=>p(142)(46),cout=>p(143)(47));
FA_ff_943:FAff port map(x=>p(21)(47),y=>p(22)(47),Cin=>p(23)(47),clock=>clock,reset=>reset,s=>p(142)(47),cout=>p(143)(48));
FA_ff_944:FAff port map(x=>p(21)(48),y=>p(22)(48),Cin=>p(23)(48),clock=>clock,reset=>reset,s=>p(142)(48),cout=>p(143)(49));
FA_ff_945:FAff port map(x=>p(21)(49),y=>p(22)(49),Cin=>p(23)(49),clock=>clock,reset=>reset,s=>p(142)(49),cout=>p(143)(50));
FA_ff_946:FAff port map(x=>p(21)(50),y=>p(22)(50),Cin=>p(23)(50),clock=>clock,reset=>reset,s=>p(142)(50),cout=>p(143)(51));
FA_ff_947:FAff port map(x=>p(21)(51),y=>p(22)(51),Cin=>p(23)(51),clock=>clock,reset=>reset,s=>p(142)(51),cout=>p(143)(52));
FA_ff_948:FAff port map(x=>p(21)(52),y=>p(22)(52),Cin=>p(23)(52),clock=>clock,reset=>reset,s=>p(142)(52),cout=>p(143)(53));
FA_ff_949:FAff port map(x=>p(21)(53),y=>p(22)(53),Cin=>p(23)(53),clock=>clock,reset=>reset,s=>p(142)(53),cout=>p(143)(54));
FA_ff_950:FAff port map(x=>p(21)(54),y=>p(22)(54),Cin=>p(23)(54),clock=>clock,reset=>reset,s=>p(142)(54),cout=>p(143)(55));
FA_ff_951:FAff port map(x=>p(21)(55),y=>p(22)(55),Cin=>p(23)(55),clock=>clock,reset=>reset,s=>p(142)(55),cout=>p(143)(56));
FA_ff_952:FAff port map(x=>p(21)(56),y=>p(22)(56),Cin=>p(23)(56),clock=>clock,reset=>reset,s=>p(142)(56),cout=>p(143)(57));
FA_ff_953:FAff port map(x=>p(21)(57),y=>p(22)(57),Cin=>p(23)(57),clock=>clock,reset=>reset,s=>p(142)(57),cout=>p(143)(58));
FA_ff_954:FAff port map(x=>p(21)(58),y=>p(22)(58),Cin=>p(23)(58),clock=>clock,reset=>reset,s=>p(142)(58),cout=>p(143)(59));
FA_ff_955:FAff port map(x=>p(21)(59),y=>p(22)(59),Cin=>p(23)(59),clock=>clock,reset=>reset,s=>p(142)(59),cout=>p(143)(60));
FA_ff_956:FAff port map(x=>p(21)(60),y=>p(22)(60),Cin=>p(23)(60),clock=>clock,reset=>reset,s=>p(142)(60),cout=>p(143)(61));
FA_ff_957:FAff port map(x=>p(21)(61),y=>p(22)(61),Cin=>p(23)(61),clock=>clock,reset=>reset,s=>p(142)(61),cout=>p(143)(62));
FA_ff_958:FAff port map(x=>p(21)(62),y=>p(22)(62),Cin=>p(23)(62),clock=>clock,reset=>reset,s=>p(142)(62),cout=>p(143)(63));
FA_ff_959:FAff port map(x=>p(21)(63),y=>p(22)(63),Cin=>p(23)(63),clock=>clock,reset=>reset,s=>p(142)(63),cout=>p(143)(64));
FA_ff_960:FAff port map(x=>p(21)(64),y=>p(22)(64),Cin=>p(23)(64),clock=>clock,reset=>reset,s=>p(142)(64),cout=>p(143)(65));
FA_ff_961:FAff port map(x=>p(21)(65),y=>p(22)(65),Cin=>p(23)(65),clock=>clock,reset=>reset,s=>p(142)(65),cout=>p(143)(66));
FA_ff_962:FAff port map(x=>p(21)(66),y=>p(22)(66),Cin=>p(23)(66),clock=>clock,reset=>reset,s=>p(142)(66),cout=>p(143)(67));
FA_ff_963:FAff port map(x=>p(21)(67),y=>p(22)(67),Cin=>p(23)(67),clock=>clock,reset=>reset,s=>p(142)(67),cout=>p(143)(68));
FA_ff_964:FAff port map(x=>p(21)(68),y=>p(22)(68),Cin=>p(23)(68),clock=>clock,reset=>reset,s=>p(142)(68),cout=>p(143)(69));
FA_ff_965:FAff port map(x=>p(21)(69),y=>p(22)(69),Cin=>p(23)(69),clock=>clock,reset=>reset,s=>p(142)(69),cout=>p(143)(70));
FA_ff_966:FAff port map(x=>p(21)(70),y=>p(22)(70),Cin=>p(23)(70),clock=>clock,reset=>reset,s=>p(142)(70),cout=>p(143)(71));
FA_ff_967:FAff port map(x=>p(21)(71),y=>p(22)(71),Cin=>p(23)(71),clock=>clock,reset=>reset,s=>p(142)(71),cout=>p(143)(72));
FA_ff_968:FAff port map(x=>p(21)(72),y=>p(22)(72),Cin=>p(23)(72),clock=>clock,reset=>reset,s=>p(142)(72),cout=>p(143)(73));
FA_ff_969:FAff port map(x=>p(21)(73),y=>p(22)(73),Cin=>p(23)(73),clock=>clock,reset=>reset,s=>p(142)(73),cout=>p(143)(74));
FA_ff_970:FAff port map(x=>p(21)(74),y=>p(22)(74),Cin=>p(23)(74),clock=>clock,reset=>reset,s=>p(142)(74),cout=>p(143)(75));
FA_ff_971:FAff port map(x=>p(21)(75),y=>p(22)(75),Cin=>p(23)(75),clock=>clock,reset=>reset,s=>p(142)(75),cout=>p(143)(76));
FA_ff_972:FAff port map(x=>p(21)(76),y=>p(22)(76),Cin=>p(23)(76),clock=>clock,reset=>reset,s=>p(142)(76),cout=>p(143)(77));
FA_ff_973:FAff port map(x=>p(21)(77),y=>p(22)(77),Cin=>p(23)(77),clock=>clock,reset=>reset,s=>p(142)(77),cout=>p(143)(78));
FA_ff_974:FAff port map(x=>p(21)(78),y=>p(22)(78),Cin=>p(23)(78),clock=>clock,reset=>reset,s=>p(142)(78),cout=>p(143)(79));
FA_ff_975:FAff port map(x=>p(21)(79),y=>p(22)(79),Cin=>p(23)(79),clock=>clock,reset=>reset,s=>p(142)(79),cout=>p(143)(80));
FA_ff_976:FAff port map(x=>p(21)(80),y=>p(22)(80),Cin=>p(23)(80),clock=>clock,reset=>reset,s=>p(142)(80),cout=>p(143)(81));
FA_ff_977:FAff port map(x=>p(21)(81),y=>p(22)(81),Cin=>p(23)(81),clock=>clock,reset=>reset,s=>p(142)(81),cout=>p(143)(82));
FA_ff_978:FAff port map(x=>p(21)(82),y=>p(22)(82),Cin=>p(23)(82),clock=>clock,reset=>reset,s=>p(142)(82),cout=>p(143)(83));
FA_ff_979:FAff port map(x=>p(21)(83),y=>p(22)(83),Cin=>p(23)(83),clock=>clock,reset=>reset,s=>p(142)(83),cout=>p(143)(84));
FA_ff_980:FAff port map(x=>p(21)(84),y=>p(22)(84),Cin=>p(23)(84),clock=>clock,reset=>reset,s=>p(142)(84),cout=>p(143)(85));
FA_ff_981:FAff port map(x=>p(21)(85),y=>p(22)(85),Cin=>p(23)(85),clock=>clock,reset=>reset,s=>p(142)(85),cout=>p(143)(86));
FA_ff_982:FAff port map(x=>p(21)(86),y=>p(22)(86),Cin=>p(23)(86),clock=>clock,reset=>reset,s=>p(142)(86),cout=>p(143)(87));
FA_ff_983:FAff port map(x=>p(21)(87),y=>p(22)(87),Cin=>p(23)(87),clock=>clock,reset=>reset,s=>p(142)(87),cout=>p(143)(88));
FA_ff_984:FAff port map(x=>p(21)(88),y=>p(22)(88),Cin=>p(23)(88),clock=>clock,reset=>reset,s=>p(142)(88),cout=>p(143)(89));
FA_ff_985:FAff port map(x=>p(21)(89),y=>p(22)(89),Cin=>p(23)(89),clock=>clock,reset=>reset,s=>p(142)(89),cout=>p(143)(90));
FA_ff_986:FAff port map(x=>p(21)(90),y=>p(22)(90),Cin=>p(23)(90),clock=>clock,reset=>reset,s=>p(142)(90),cout=>p(143)(91));
FA_ff_987:FAff port map(x=>p(21)(91),y=>p(22)(91),Cin=>p(23)(91),clock=>clock,reset=>reset,s=>p(142)(91),cout=>p(143)(92));
FA_ff_988:FAff port map(x=>p(21)(92),y=>p(22)(92),Cin=>p(23)(92),clock=>clock,reset=>reset,s=>p(142)(92),cout=>p(143)(93));
FA_ff_989:FAff port map(x=>p(21)(93),y=>p(22)(93),Cin=>p(23)(93),clock=>clock,reset=>reset,s=>p(142)(93),cout=>p(143)(94));
FA_ff_990:FAff port map(x=>p(21)(94),y=>p(22)(94),Cin=>p(23)(94),clock=>clock,reset=>reset,s=>p(142)(94),cout=>p(143)(95));
FA_ff_991:FAff port map(x=>p(21)(95),y=>p(22)(95),Cin=>p(23)(95),clock=>clock,reset=>reset,s=>p(142)(95),cout=>p(143)(96));
FA_ff_992:FAff port map(x=>p(21)(96),y=>p(22)(96),Cin=>p(23)(96),clock=>clock,reset=>reset,s=>p(142)(96),cout=>p(143)(97));
FA_ff_993:FAff port map(x=>p(21)(97),y=>p(22)(97),Cin=>p(23)(97),clock=>clock,reset=>reset,s=>p(142)(97),cout=>p(143)(98));
FA_ff_994:FAff port map(x=>p(21)(98),y=>p(22)(98),Cin=>p(23)(98),clock=>clock,reset=>reset,s=>p(142)(98),cout=>p(143)(99));
FA_ff_995:FAff port map(x=>p(21)(99),y=>p(22)(99),Cin=>p(23)(99),clock=>clock,reset=>reset,s=>p(142)(99),cout=>p(143)(100));
FA_ff_996:FAff port map(x=>p(21)(100),y=>p(22)(100),Cin=>p(23)(100),clock=>clock,reset=>reset,s=>p(142)(100),cout=>p(143)(101));
FA_ff_997:FAff port map(x=>p(21)(101),y=>p(22)(101),Cin=>p(23)(101),clock=>clock,reset=>reset,s=>p(142)(101),cout=>p(143)(102));
FA_ff_998:FAff port map(x=>p(21)(102),y=>p(22)(102),Cin=>p(23)(102),clock=>clock,reset=>reset,s=>p(142)(102),cout=>p(143)(103));
FA_ff_999:FAff port map(x=>p(21)(103),y=>p(22)(103),Cin=>p(23)(103),clock=>clock,reset=>reset,s=>p(142)(103),cout=>p(143)(104));
FA_ff_1000:FAff port map(x=>p(21)(104),y=>p(22)(104),Cin=>p(23)(104),clock=>clock,reset=>reset,s=>p(142)(104),cout=>p(143)(105));
FA_ff_1001:FAff port map(x=>p(21)(105),y=>p(22)(105),Cin=>p(23)(105),clock=>clock,reset=>reset,s=>p(142)(105),cout=>p(143)(106));
FA_ff_1002:FAff port map(x=>p(21)(106),y=>p(22)(106),Cin=>p(23)(106),clock=>clock,reset=>reset,s=>p(142)(106),cout=>p(143)(107));
FA_ff_1003:FAff port map(x=>p(21)(107),y=>p(22)(107),Cin=>p(23)(107),clock=>clock,reset=>reset,s=>p(142)(107),cout=>p(143)(108));
FA_ff_1004:FAff port map(x=>p(21)(108),y=>p(22)(108),Cin=>p(23)(108),clock=>clock,reset=>reset,s=>p(142)(108),cout=>p(143)(109));
FA_ff_1005:FAff port map(x=>p(21)(109),y=>p(22)(109),Cin=>p(23)(109),clock=>clock,reset=>reset,s=>p(142)(109),cout=>p(143)(110));
FA_ff_1006:FAff port map(x=>p(21)(110),y=>p(22)(110),Cin=>p(23)(110),clock=>clock,reset=>reset,s=>p(142)(110),cout=>p(143)(111));
FA_ff_1007:FAff port map(x=>p(21)(111),y=>p(22)(111),Cin=>p(23)(111),clock=>clock,reset=>reset,s=>p(142)(111),cout=>p(143)(112));
FA_ff_1008:FAff port map(x=>p(21)(112),y=>p(22)(112),Cin=>p(23)(112),clock=>clock,reset=>reset,s=>p(142)(112),cout=>p(143)(113));
FA_ff_1009:FAff port map(x=>p(21)(113),y=>p(22)(113),Cin=>p(23)(113),clock=>clock,reset=>reset,s=>p(142)(113),cout=>p(143)(114));
FA_ff_1010:FAff port map(x=>p(21)(114),y=>p(22)(114),Cin=>p(23)(114),clock=>clock,reset=>reset,s=>p(142)(114),cout=>p(143)(115));
FA_ff_1011:FAff port map(x=>p(21)(115),y=>p(22)(115),Cin=>p(23)(115),clock=>clock,reset=>reset,s=>p(142)(115),cout=>p(143)(116));
FA_ff_1012:FAff port map(x=>p(21)(116),y=>p(22)(116),Cin=>p(23)(116),clock=>clock,reset=>reset,s=>p(142)(116),cout=>p(143)(117));
FA_ff_1013:FAff port map(x=>p(21)(117),y=>p(22)(117),Cin=>p(23)(117),clock=>clock,reset=>reset,s=>p(142)(117),cout=>p(143)(118));
FA_ff_1014:FAff port map(x=>p(21)(118),y=>p(22)(118),Cin=>p(23)(118),clock=>clock,reset=>reset,s=>p(142)(118),cout=>p(143)(119));
FA_ff_1015:FAff port map(x=>p(21)(119),y=>p(22)(119),Cin=>p(23)(119),clock=>clock,reset=>reset,s=>p(142)(119),cout=>p(143)(120));
FA_ff_1016:FAff port map(x=>p(21)(120),y=>p(22)(120),Cin=>p(23)(120),clock=>clock,reset=>reset,s=>p(142)(120),cout=>p(143)(121));
FA_ff_1017:FAff port map(x=>p(21)(121),y=>p(22)(121),Cin=>p(23)(121),clock=>clock,reset=>reset,s=>p(142)(121),cout=>p(143)(122));
FA_ff_1018:FAff port map(x=>p(21)(122),y=>p(22)(122),Cin=>p(23)(122),clock=>clock,reset=>reset,s=>p(142)(122),cout=>p(143)(123));
FA_ff_1019:FAff port map(x=>p(21)(123),y=>p(22)(123),Cin=>p(23)(123),clock=>clock,reset=>reset,s=>p(142)(123),cout=>p(143)(124));
FA_ff_1020:FAff port map(x=>p(21)(124),y=>p(22)(124),Cin=>p(23)(124),clock=>clock,reset=>reset,s=>p(142)(124),cout=>p(143)(125));
FA_ff_1021:FAff port map(x=>p(21)(125),y=>p(22)(125),Cin=>p(23)(125),clock=>clock,reset=>reset,s=>p(142)(125),cout=>p(143)(126));
FA_ff_1022:FAff port map(x=>p(21)(126),y=>p(22)(126),Cin=>p(23)(126),clock=>clock,reset=>reset,s=>p(142)(126),cout=>p(143)(127));
FA_ff_1023:FAff port map(x=>p(21)(127),y=>p(22)(127),Cin=>p(23)(127),clock=>clock,reset=>reset,s=>p(142)(127),cout=>p(143)(128));
FA_ff_1024:FAff port map(x=>p(24)(0),y=>p(25)(0),Cin=>p(26)(0),clock=>clock,reset=>reset,s=>p(144)(0),cout=>p(145)(1));
FA_ff_1025:FAff port map(x=>p(24)(1),y=>p(25)(1),Cin=>p(26)(1),clock=>clock,reset=>reset,s=>p(144)(1),cout=>p(145)(2));
FA_ff_1026:FAff port map(x=>p(24)(2),y=>p(25)(2),Cin=>p(26)(2),clock=>clock,reset=>reset,s=>p(144)(2),cout=>p(145)(3));
FA_ff_1027:FAff port map(x=>p(24)(3),y=>p(25)(3),Cin=>p(26)(3),clock=>clock,reset=>reset,s=>p(144)(3),cout=>p(145)(4));
FA_ff_1028:FAff port map(x=>p(24)(4),y=>p(25)(4),Cin=>p(26)(4),clock=>clock,reset=>reset,s=>p(144)(4),cout=>p(145)(5));
FA_ff_1029:FAff port map(x=>p(24)(5),y=>p(25)(5),Cin=>p(26)(5),clock=>clock,reset=>reset,s=>p(144)(5),cout=>p(145)(6));
FA_ff_1030:FAff port map(x=>p(24)(6),y=>p(25)(6),Cin=>p(26)(6),clock=>clock,reset=>reset,s=>p(144)(6),cout=>p(145)(7));
FA_ff_1031:FAff port map(x=>p(24)(7),y=>p(25)(7),Cin=>p(26)(7),clock=>clock,reset=>reset,s=>p(144)(7),cout=>p(145)(8));
FA_ff_1032:FAff port map(x=>p(24)(8),y=>p(25)(8),Cin=>p(26)(8),clock=>clock,reset=>reset,s=>p(144)(8),cout=>p(145)(9));
FA_ff_1033:FAff port map(x=>p(24)(9),y=>p(25)(9),Cin=>p(26)(9),clock=>clock,reset=>reset,s=>p(144)(9),cout=>p(145)(10));
FA_ff_1034:FAff port map(x=>p(24)(10),y=>p(25)(10),Cin=>p(26)(10),clock=>clock,reset=>reset,s=>p(144)(10),cout=>p(145)(11));
FA_ff_1035:FAff port map(x=>p(24)(11),y=>p(25)(11),Cin=>p(26)(11),clock=>clock,reset=>reset,s=>p(144)(11),cout=>p(145)(12));
FA_ff_1036:FAff port map(x=>p(24)(12),y=>p(25)(12),Cin=>p(26)(12),clock=>clock,reset=>reset,s=>p(144)(12),cout=>p(145)(13));
FA_ff_1037:FAff port map(x=>p(24)(13),y=>p(25)(13),Cin=>p(26)(13),clock=>clock,reset=>reset,s=>p(144)(13),cout=>p(145)(14));
FA_ff_1038:FAff port map(x=>p(24)(14),y=>p(25)(14),Cin=>p(26)(14),clock=>clock,reset=>reset,s=>p(144)(14),cout=>p(145)(15));
FA_ff_1039:FAff port map(x=>p(24)(15),y=>p(25)(15),Cin=>p(26)(15),clock=>clock,reset=>reset,s=>p(144)(15),cout=>p(145)(16));
FA_ff_1040:FAff port map(x=>p(24)(16),y=>p(25)(16),Cin=>p(26)(16),clock=>clock,reset=>reset,s=>p(144)(16),cout=>p(145)(17));
FA_ff_1041:FAff port map(x=>p(24)(17),y=>p(25)(17),Cin=>p(26)(17),clock=>clock,reset=>reset,s=>p(144)(17),cout=>p(145)(18));
FA_ff_1042:FAff port map(x=>p(24)(18),y=>p(25)(18),Cin=>p(26)(18),clock=>clock,reset=>reset,s=>p(144)(18),cout=>p(145)(19));
FA_ff_1043:FAff port map(x=>p(24)(19),y=>p(25)(19),Cin=>p(26)(19),clock=>clock,reset=>reset,s=>p(144)(19),cout=>p(145)(20));
FA_ff_1044:FAff port map(x=>p(24)(20),y=>p(25)(20),Cin=>p(26)(20),clock=>clock,reset=>reset,s=>p(144)(20),cout=>p(145)(21));
FA_ff_1045:FAff port map(x=>p(24)(21),y=>p(25)(21),Cin=>p(26)(21),clock=>clock,reset=>reset,s=>p(144)(21),cout=>p(145)(22));
FA_ff_1046:FAff port map(x=>p(24)(22),y=>p(25)(22),Cin=>p(26)(22),clock=>clock,reset=>reset,s=>p(144)(22),cout=>p(145)(23));
FA_ff_1047:FAff port map(x=>p(24)(23),y=>p(25)(23),Cin=>p(26)(23),clock=>clock,reset=>reset,s=>p(144)(23),cout=>p(145)(24));
FA_ff_1048:FAff port map(x=>p(24)(24),y=>p(25)(24),Cin=>p(26)(24),clock=>clock,reset=>reset,s=>p(144)(24),cout=>p(145)(25));
FA_ff_1049:FAff port map(x=>p(24)(25),y=>p(25)(25),Cin=>p(26)(25),clock=>clock,reset=>reset,s=>p(144)(25),cout=>p(145)(26));
FA_ff_1050:FAff port map(x=>p(24)(26),y=>p(25)(26),Cin=>p(26)(26),clock=>clock,reset=>reset,s=>p(144)(26),cout=>p(145)(27));
FA_ff_1051:FAff port map(x=>p(24)(27),y=>p(25)(27),Cin=>p(26)(27),clock=>clock,reset=>reset,s=>p(144)(27),cout=>p(145)(28));
FA_ff_1052:FAff port map(x=>p(24)(28),y=>p(25)(28),Cin=>p(26)(28),clock=>clock,reset=>reset,s=>p(144)(28),cout=>p(145)(29));
FA_ff_1053:FAff port map(x=>p(24)(29),y=>p(25)(29),Cin=>p(26)(29),clock=>clock,reset=>reset,s=>p(144)(29),cout=>p(145)(30));
FA_ff_1054:FAff port map(x=>p(24)(30),y=>p(25)(30),Cin=>p(26)(30),clock=>clock,reset=>reset,s=>p(144)(30),cout=>p(145)(31));
FA_ff_1055:FAff port map(x=>p(24)(31),y=>p(25)(31),Cin=>p(26)(31),clock=>clock,reset=>reset,s=>p(144)(31),cout=>p(145)(32));
FA_ff_1056:FAff port map(x=>p(24)(32),y=>p(25)(32),Cin=>p(26)(32),clock=>clock,reset=>reset,s=>p(144)(32),cout=>p(145)(33));
FA_ff_1057:FAff port map(x=>p(24)(33),y=>p(25)(33),Cin=>p(26)(33),clock=>clock,reset=>reset,s=>p(144)(33),cout=>p(145)(34));
FA_ff_1058:FAff port map(x=>p(24)(34),y=>p(25)(34),Cin=>p(26)(34),clock=>clock,reset=>reset,s=>p(144)(34),cout=>p(145)(35));
FA_ff_1059:FAff port map(x=>p(24)(35),y=>p(25)(35),Cin=>p(26)(35),clock=>clock,reset=>reset,s=>p(144)(35),cout=>p(145)(36));
FA_ff_1060:FAff port map(x=>p(24)(36),y=>p(25)(36),Cin=>p(26)(36),clock=>clock,reset=>reset,s=>p(144)(36),cout=>p(145)(37));
FA_ff_1061:FAff port map(x=>p(24)(37),y=>p(25)(37),Cin=>p(26)(37),clock=>clock,reset=>reset,s=>p(144)(37),cout=>p(145)(38));
FA_ff_1062:FAff port map(x=>p(24)(38),y=>p(25)(38),Cin=>p(26)(38),clock=>clock,reset=>reset,s=>p(144)(38),cout=>p(145)(39));
FA_ff_1063:FAff port map(x=>p(24)(39),y=>p(25)(39),Cin=>p(26)(39),clock=>clock,reset=>reset,s=>p(144)(39),cout=>p(145)(40));
FA_ff_1064:FAff port map(x=>p(24)(40),y=>p(25)(40),Cin=>p(26)(40),clock=>clock,reset=>reset,s=>p(144)(40),cout=>p(145)(41));
FA_ff_1065:FAff port map(x=>p(24)(41),y=>p(25)(41),Cin=>p(26)(41),clock=>clock,reset=>reset,s=>p(144)(41),cout=>p(145)(42));
FA_ff_1066:FAff port map(x=>p(24)(42),y=>p(25)(42),Cin=>p(26)(42),clock=>clock,reset=>reset,s=>p(144)(42),cout=>p(145)(43));
FA_ff_1067:FAff port map(x=>p(24)(43),y=>p(25)(43),Cin=>p(26)(43),clock=>clock,reset=>reset,s=>p(144)(43),cout=>p(145)(44));
FA_ff_1068:FAff port map(x=>p(24)(44),y=>p(25)(44),Cin=>p(26)(44),clock=>clock,reset=>reset,s=>p(144)(44),cout=>p(145)(45));
FA_ff_1069:FAff port map(x=>p(24)(45),y=>p(25)(45),Cin=>p(26)(45),clock=>clock,reset=>reset,s=>p(144)(45),cout=>p(145)(46));
FA_ff_1070:FAff port map(x=>p(24)(46),y=>p(25)(46),Cin=>p(26)(46),clock=>clock,reset=>reset,s=>p(144)(46),cout=>p(145)(47));
FA_ff_1071:FAff port map(x=>p(24)(47),y=>p(25)(47),Cin=>p(26)(47),clock=>clock,reset=>reset,s=>p(144)(47),cout=>p(145)(48));
FA_ff_1072:FAff port map(x=>p(24)(48),y=>p(25)(48),Cin=>p(26)(48),clock=>clock,reset=>reset,s=>p(144)(48),cout=>p(145)(49));
FA_ff_1073:FAff port map(x=>p(24)(49),y=>p(25)(49),Cin=>p(26)(49),clock=>clock,reset=>reset,s=>p(144)(49),cout=>p(145)(50));
FA_ff_1074:FAff port map(x=>p(24)(50),y=>p(25)(50),Cin=>p(26)(50),clock=>clock,reset=>reset,s=>p(144)(50),cout=>p(145)(51));
FA_ff_1075:FAff port map(x=>p(24)(51),y=>p(25)(51),Cin=>p(26)(51),clock=>clock,reset=>reset,s=>p(144)(51),cout=>p(145)(52));
FA_ff_1076:FAff port map(x=>p(24)(52),y=>p(25)(52),Cin=>p(26)(52),clock=>clock,reset=>reset,s=>p(144)(52),cout=>p(145)(53));
FA_ff_1077:FAff port map(x=>p(24)(53),y=>p(25)(53),Cin=>p(26)(53),clock=>clock,reset=>reset,s=>p(144)(53),cout=>p(145)(54));
FA_ff_1078:FAff port map(x=>p(24)(54),y=>p(25)(54),Cin=>p(26)(54),clock=>clock,reset=>reset,s=>p(144)(54),cout=>p(145)(55));
FA_ff_1079:FAff port map(x=>p(24)(55),y=>p(25)(55),Cin=>p(26)(55),clock=>clock,reset=>reset,s=>p(144)(55),cout=>p(145)(56));
FA_ff_1080:FAff port map(x=>p(24)(56),y=>p(25)(56),Cin=>p(26)(56),clock=>clock,reset=>reset,s=>p(144)(56),cout=>p(145)(57));
FA_ff_1081:FAff port map(x=>p(24)(57),y=>p(25)(57),Cin=>p(26)(57),clock=>clock,reset=>reset,s=>p(144)(57),cout=>p(145)(58));
FA_ff_1082:FAff port map(x=>p(24)(58),y=>p(25)(58),Cin=>p(26)(58),clock=>clock,reset=>reset,s=>p(144)(58),cout=>p(145)(59));
FA_ff_1083:FAff port map(x=>p(24)(59),y=>p(25)(59),Cin=>p(26)(59),clock=>clock,reset=>reset,s=>p(144)(59),cout=>p(145)(60));
FA_ff_1084:FAff port map(x=>p(24)(60),y=>p(25)(60),Cin=>p(26)(60),clock=>clock,reset=>reset,s=>p(144)(60),cout=>p(145)(61));
FA_ff_1085:FAff port map(x=>p(24)(61),y=>p(25)(61),Cin=>p(26)(61),clock=>clock,reset=>reset,s=>p(144)(61),cout=>p(145)(62));
FA_ff_1086:FAff port map(x=>p(24)(62),y=>p(25)(62),Cin=>p(26)(62),clock=>clock,reset=>reset,s=>p(144)(62),cout=>p(145)(63));
FA_ff_1087:FAff port map(x=>p(24)(63),y=>p(25)(63),Cin=>p(26)(63),clock=>clock,reset=>reset,s=>p(144)(63),cout=>p(145)(64));
FA_ff_1088:FAff port map(x=>p(24)(64),y=>p(25)(64),Cin=>p(26)(64),clock=>clock,reset=>reset,s=>p(144)(64),cout=>p(145)(65));
FA_ff_1089:FAff port map(x=>p(24)(65),y=>p(25)(65),Cin=>p(26)(65),clock=>clock,reset=>reset,s=>p(144)(65),cout=>p(145)(66));
FA_ff_1090:FAff port map(x=>p(24)(66),y=>p(25)(66),Cin=>p(26)(66),clock=>clock,reset=>reset,s=>p(144)(66),cout=>p(145)(67));
FA_ff_1091:FAff port map(x=>p(24)(67),y=>p(25)(67),Cin=>p(26)(67),clock=>clock,reset=>reset,s=>p(144)(67),cout=>p(145)(68));
FA_ff_1092:FAff port map(x=>p(24)(68),y=>p(25)(68),Cin=>p(26)(68),clock=>clock,reset=>reset,s=>p(144)(68),cout=>p(145)(69));
FA_ff_1093:FAff port map(x=>p(24)(69),y=>p(25)(69),Cin=>p(26)(69),clock=>clock,reset=>reset,s=>p(144)(69),cout=>p(145)(70));
FA_ff_1094:FAff port map(x=>p(24)(70),y=>p(25)(70),Cin=>p(26)(70),clock=>clock,reset=>reset,s=>p(144)(70),cout=>p(145)(71));
FA_ff_1095:FAff port map(x=>p(24)(71),y=>p(25)(71),Cin=>p(26)(71),clock=>clock,reset=>reset,s=>p(144)(71),cout=>p(145)(72));
FA_ff_1096:FAff port map(x=>p(24)(72),y=>p(25)(72),Cin=>p(26)(72),clock=>clock,reset=>reset,s=>p(144)(72),cout=>p(145)(73));
FA_ff_1097:FAff port map(x=>p(24)(73),y=>p(25)(73),Cin=>p(26)(73),clock=>clock,reset=>reset,s=>p(144)(73),cout=>p(145)(74));
FA_ff_1098:FAff port map(x=>p(24)(74),y=>p(25)(74),Cin=>p(26)(74),clock=>clock,reset=>reset,s=>p(144)(74),cout=>p(145)(75));
FA_ff_1099:FAff port map(x=>p(24)(75),y=>p(25)(75),Cin=>p(26)(75),clock=>clock,reset=>reset,s=>p(144)(75),cout=>p(145)(76));
FA_ff_1100:FAff port map(x=>p(24)(76),y=>p(25)(76),Cin=>p(26)(76),clock=>clock,reset=>reset,s=>p(144)(76),cout=>p(145)(77));
FA_ff_1101:FAff port map(x=>p(24)(77),y=>p(25)(77),Cin=>p(26)(77),clock=>clock,reset=>reset,s=>p(144)(77),cout=>p(145)(78));
FA_ff_1102:FAff port map(x=>p(24)(78),y=>p(25)(78),Cin=>p(26)(78),clock=>clock,reset=>reset,s=>p(144)(78),cout=>p(145)(79));
FA_ff_1103:FAff port map(x=>p(24)(79),y=>p(25)(79),Cin=>p(26)(79),clock=>clock,reset=>reset,s=>p(144)(79),cout=>p(145)(80));
FA_ff_1104:FAff port map(x=>p(24)(80),y=>p(25)(80),Cin=>p(26)(80),clock=>clock,reset=>reset,s=>p(144)(80),cout=>p(145)(81));
FA_ff_1105:FAff port map(x=>p(24)(81),y=>p(25)(81),Cin=>p(26)(81),clock=>clock,reset=>reset,s=>p(144)(81),cout=>p(145)(82));
FA_ff_1106:FAff port map(x=>p(24)(82),y=>p(25)(82),Cin=>p(26)(82),clock=>clock,reset=>reset,s=>p(144)(82),cout=>p(145)(83));
FA_ff_1107:FAff port map(x=>p(24)(83),y=>p(25)(83),Cin=>p(26)(83),clock=>clock,reset=>reset,s=>p(144)(83),cout=>p(145)(84));
FA_ff_1108:FAff port map(x=>p(24)(84),y=>p(25)(84),Cin=>p(26)(84),clock=>clock,reset=>reset,s=>p(144)(84),cout=>p(145)(85));
FA_ff_1109:FAff port map(x=>p(24)(85),y=>p(25)(85),Cin=>p(26)(85),clock=>clock,reset=>reset,s=>p(144)(85),cout=>p(145)(86));
FA_ff_1110:FAff port map(x=>p(24)(86),y=>p(25)(86),Cin=>p(26)(86),clock=>clock,reset=>reset,s=>p(144)(86),cout=>p(145)(87));
FA_ff_1111:FAff port map(x=>p(24)(87),y=>p(25)(87),Cin=>p(26)(87),clock=>clock,reset=>reset,s=>p(144)(87),cout=>p(145)(88));
FA_ff_1112:FAff port map(x=>p(24)(88),y=>p(25)(88),Cin=>p(26)(88),clock=>clock,reset=>reset,s=>p(144)(88),cout=>p(145)(89));
FA_ff_1113:FAff port map(x=>p(24)(89),y=>p(25)(89),Cin=>p(26)(89),clock=>clock,reset=>reset,s=>p(144)(89),cout=>p(145)(90));
FA_ff_1114:FAff port map(x=>p(24)(90),y=>p(25)(90),Cin=>p(26)(90),clock=>clock,reset=>reset,s=>p(144)(90),cout=>p(145)(91));
FA_ff_1115:FAff port map(x=>p(24)(91),y=>p(25)(91),Cin=>p(26)(91),clock=>clock,reset=>reset,s=>p(144)(91),cout=>p(145)(92));
FA_ff_1116:FAff port map(x=>p(24)(92),y=>p(25)(92),Cin=>p(26)(92),clock=>clock,reset=>reset,s=>p(144)(92),cout=>p(145)(93));
FA_ff_1117:FAff port map(x=>p(24)(93),y=>p(25)(93),Cin=>p(26)(93),clock=>clock,reset=>reset,s=>p(144)(93),cout=>p(145)(94));
FA_ff_1118:FAff port map(x=>p(24)(94),y=>p(25)(94),Cin=>p(26)(94),clock=>clock,reset=>reset,s=>p(144)(94),cout=>p(145)(95));
FA_ff_1119:FAff port map(x=>p(24)(95),y=>p(25)(95),Cin=>p(26)(95),clock=>clock,reset=>reset,s=>p(144)(95),cout=>p(145)(96));
FA_ff_1120:FAff port map(x=>p(24)(96),y=>p(25)(96),Cin=>p(26)(96),clock=>clock,reset=>reset,s=>p(144)(96),cout=>p(145)(97));
FA_ff_1121:FAff port map(x=>p(24)(97),y=>p(25)(97),Cin=>p(26)(97),clock=>clock,reset=>reset,s=>p(144)(97),cout=>p(145)(98));
FA_ff_1122:FAff port map(x=>p(24)(98),y=>p(25)(98),Cin=>p(26)(98),clock=>clock,reset=>reset,s=>p(144)(98),cout=>p(145)(99));
FA_ff_1123:FAff port map(x=>p(24)(99),y=>p(25)(99),Cin=>p(26)(99),clock=>clock,reset=>reset,s=>p(144)(99),cout=>p(145)(100));
FA_ff_1124:FAff port map(x=>p(24)(100),y=>p(25)(100),Cin=>p(26)(100),clock=>clock,reset=>reset,s=>p(144)(100),cout=>p(145)(101));
FA_ff_1125:FAff port map(x=>p(24)(101),y=>p(25)(101),Cin=>p(26)(101),clock=>clock,reset=>reset,s=>p(144)(101),cout=>p(145)(102));
FA_ff_1126:FAff port map(x=>p(24)(102),y=>p(25)(102),Cin=>p(26)(102),clock=>clock,reset=>reset,s=>p(144)(102),cout=>p(145)(103));
FA_ff_1127:FAff port map(x=>p(24)(103),y=>p(25)(103),Cin=>p(26)(103),clock=>clock,reset=>reset,s=>p(144)(103),cout=>p(145)(104));
FA_ff_1128:FAff port map(x=>p(24)(104),y=>p(25)(104),Cin=>p(26)(104),clock=>clock,reset=>reset,s=>p(144)(104),cout=>p(145)(105));
FA_ff_1129:FAff port map(x=>p(24)(105),y=>p(25)(105),Cin=>p(26)(105),clock=>clock,reset=>reset,s=>p(144)(105),cout=>p(145)(106));
FA_ff_1130:FAff port map(x=>p(24)(106),y=>p(25)(106),Cin=>p(26)(106),clock=>clock,reset=>reset,s=>p(144)(106),cout=>p(145)(107));
FA_ff_1131:FAff port map(x=>p(24)(107),y=>p(25)(107),Cin=>p(26)(107),clock=>clock,reset=>reset,s=>p(144)(107),cout=>p(145)(108));
FA_ff_1132:FAff port map(x=>p(24)(108),y=>p(25)(108),Cin=>p(26)(108),clock=>clock,reset=>reset,s=>p(144)(108),cout=>p(145)(109));
FA_ff_1133:FAff port map(x=>p(24)(109),y=>p(25)(109),Cin=>p(26)(109),clock=>clock,reset=>reset,s=>p(144)(109),cout=>p(145)(110));
FA_ff_1134:FAff port map(x=>p(24)(110),y=>p(25)(110),Cin=>p(26)(110),clock=>clock,reset=>reset,s=>p(144)(110),cout=>p(145)(111));
FA_ff_1135:FAff port map(x=>p(24)(111),y=>p(25)(111),Cin=>p(26)(111),clock=>clock,reset=>reset,s=>p(144)(111),cout=>p(145)(112));
FA_ff_1136:FAff port map(x=>p(24)(112),y=>p(25)(112),Cin=>p(26)(112),clock=>clock,reset=>reset,s=>p(144)(112),cout=>p(145)(113));
FA_ff_1137:FAff port map(x=>p(24)(113),y=>p(25)(113),Cin=>p(26)(113),clock=>clock,reset=>reset,s=>p(144)(113),cout=>p(145)(114));
FA_ff_1138:FAff port map(x=>p(24)(114),y=>p(25)(114),Cin=>p(26)(114),clock=>clock,reset=>reset,s=>p(144)(114),cout=>p(145)(115));
FA_ff_1139:FAff port map(x=>p(24)(115),y=>p(25)(115),Cin=>p(26)(115),clock=>clock,reset=>reset,s=>p(144)(115),cout=>p(145)(116));
FA_ff_1140:FAff port map(x=>p(24)(116),y=>p(25)(116),Cin=>p(26)(116),clock=>clock,reset=>reset,s=>p(144)(116),cout=>p(145)(117));
FA_ff_1141:FAff port map(x=>p(24)(117),y=>p(25)(117),Cin=>p(26)(117),clock=>clock,reset=>reset,s=>p(144)(117),cout=>p(145)(118));
FA_ff_1142:FAff port map(x=>p(24)(118),y=>p(25)(118),Cin=>p(26)(118),clock=>clock,reset=>reset,s=>p(144)(118),cout=>p(145)(119));
FA_ff_1143:FAff port map(x=>p(24)(119),y=>p(25)(119),Cin=>p(26)(119),clock=>clock,reset=>reset,s=>p(144)(119),cout=>p(145)(120));
FA_ff_1144:FAff port map(x=>p(24)(120),y=>p(25)(120),Cin=>p(26)(120),clock=>clock,reset=>reset,s=>p(144)(120),cout=>p(145)(121));
FA_ff_1145:FAff port map(x=>p(24)(121),y=>p(25)(121),Cin=>p(26)(121),clock=>clock,reset=>reset,s=>p(144)(121),cout=>p(145)(122));
FA_ff_1146:FAff port map(x=>p(24)(122),y=>p(25)(122),Cin=>p(26)(122),clock=>clock,reset=>reset,s=>p(144)(122),cout=>p(145)(123));
FA_ff_1147:FAff port map(x=>p(24)(123),y=>p(25)(123),Cin=>p(26)(123),clock=>clock,reset=>reset,s=>p(144)(123),cout=>p(145)(124));
FA_ff_1148:FAff port map(x=>p(24)(124),y=>p(25)(124),Cin=>p(26)(124),clock=>clock,reset=>reset,s=>p(144)(124),cout=>p(145)(125));
FA_ff_1149:FAff port map(x=>p(24)(125),y=>p(25)(125),Cin=>p(26)(125),clock=>clock,reset=>reset,s=>p(144)(125),cout=>p(145)(126));
FA_ff_1150:FAff port map(x=>p(24)(126),y=>p(25)(126),Cin=>p(26)(126),clock=>clock,reset=>reset,s=>p(144)(126),cout=>p(145)(127));
FA_ff_1151:FAff port map(x=>p(24)(127),y=>p(25)(127),Cin=>p(26)(127),clock=>clock,reset=>reset,s=>p(144)(127),cout=>p(145)(128));
FA_ff_1152:FAff port map(x=>p(27)(0),y=>p(28)(0),Cin=>p(29)(0),clock=>clock,reset=>reset,s=>p(146)(0),cout=>p(147)(1));
FA_ff_1153:FAff port map(x=>p(27)(1),y=>p(28)(1),Cin=>p(29)(1),clock=>clock,reset=>reset,s=>p(146)(1),cout=>p(147)(2));
FA_ff_1154:FAff port map(x=>p(27)(2),y=>p(28)(2),Cin=>p(29)(2),clock=>clock,reset=>reset,s=>p(146)(2),cout=>p(147)(3));
FA_ff_1155:FAff port map(x=>p(27)(3),y=>p(28)(3),Cin=>p(29)(3),clock=>clock,reset=>reset,s=>p(146)(3),cout=>p(147)(4));
FA_ff_1156:FAff port map(x=>p(27)(4),y=>p(28)(4),Cin=>p(29)(4),clock=>clock,reset=>reset,s=>p(146)(4),cout=>p(147)(5));
FA_ff_1157:FAff port map(x=>p(27)(5),y=>p(28)(5),Cin=>p(29)(5),clock=>clock,reset=>reset,s=>p(146)(5),cout=>p(147)(6));
FA_ff_1158:FAff port map(x=>p(27)(6),y=>p(28)(6),Cin=>p(29)(6),clock=>clock,reset=>reset,s=>p(146)(6),cout=>p(147)(7));
FA_ff_1159:FAff port map(x=>p(27)(7),y=>p(28)(7),Cin=>p(29)(7),clock=>clock,reset=>reset,s=>p(146)(7),cout=>p(147)(8));
FA_ff_1160:FAff port map(x=>p(27)(8),y=>p(28)(8),Cin=>p(29)(8),clock=>clock,reset=>reset,s=>p(146)(8),cout=>p(147)(9));
FA_ff_1161:FAff port map(x=>p(27)(9),y=>p(28)(9),Cin=>p(29)(9),clock=>clock,reset=>reset,s=>p(146)(9),cout=>p(147)(10));
FA_ff_1162:FAff port map(x=>p(27)(10),y=>p(28)(10),Cin=>p(29)(10),clock=>clock,reset=>reset,s=>p(146)(10),cout=>p(147)(11));
FA_ff_1163:FAff port map(x=>p(27)(11),y=>p(28)(11),Cin=>p(29)(11),clock=>clock,reset=>reset,s=>p(146)(11),cout=>p(147)(12));
FA_ff_1164:FAff port map(x=>p(27)(12),y=>p(28)(12),Cin=>p(29)(12),clock=>clock,reset=>reset,s=>p(146)(12),cout=>p(147)(13));
FA_ff_1165:FAff port map(x=>p(27)(13),y=>p(28)(13),Cin=>p(29)(13),clock=>clock,reset=>reset,s=>p(146)(13),cout=>p(147)(14));
FA_ff_1166:FAff port map(x=>p(27)(14),y=>p(28)(14),Cin=>p(29)(14),clock=>clock,reset=>reset,s=>p(146)(14),cout=>p(147)(15));
FA_ff_1167:FAff port map(x=>p(27)(15),y=>p(28)(15),Cin=>p(29)(15),clock=>clock,reset=>reset,s=>p(146)(15),cout=>p(147)(16));
FA_ff_1168:FAff port map(x=>p(27)(16),y=>p(28)(16),Cin=>p(29)(16),clock=>clock,reset=>reset,s=>p(146)(16),cout=>p(147)(17));
FA_ff_1169:FAff port map(x=>p(27)(17),y=>p(28)(17),Cin=>p(29)(17),clock=>clock,reset=>reset,s=>p(146)(17),cout=>p(147)(18));
FA_ff_1170:FAff port map(x=>p(27)(18),y=>p(28)(18),Cin=>p(29)(18),clock=>clock,reset=>reset,s=>p(146)(18),cout=>p(147)(19));
FA_ff_1171:FAff port map(x=>p(27)(19),y=>p(28)(19),Cin=>p(29)(19),clock=>clock,reset=>reset,s=>p(146)(19),cout=>p(147)(20));
FA_ff_1172:FAff port map(x=>p(27)(20),y=>p(28)(20),Cin=>p(29)(20),clock=>clock,reset=>reset,s=>p(146)(20),cout=>p(147)(21));
FA_ff_1173:FAff port map(x=>p(27)(21),y=>p(28)(21),Cin=>p(29)(21),clock=>clock,reset=>reset,s=>p(146)(21),cout=>p(147)(22));
FA_ff_1174:FAff port map(x=>p(27)(22),y=>p(28)(22),Cin=>p(29)(22),clock=>clock,reset=>reset,s=>p(146)(22),cout=>p(147)(23));
FA_ff_1175:FAff port map(x=>p(27)(23),y=>p(28)(23),Cin=>p(29)(23),clock=>clock,reset=>reset,s=>p(146)(23),cout=>p(147)(24));
FA_ff_1176:FAff port map(x=>p(27)(24),y=>p(28)(24),Cin=>p(29)(24),clock=>clock,reset=>reset,s=>p(146)(24),cout=>p(147)(25));
FA_ff_1177:FAff port map(x=>p(27)(25),y=>p(28)(25),Cin=>p(29)(25),clock=>clock,reset=>reset,s=>p(146)(25),cout=>p(147)(26));
FA_ff_1178:FAff port map(x=>p(27)(26),y=>p(28)(26),Cin=>p(29)(26),clock=>clock,reset=>reset,s=>p(146)(26),cout=>p(147)(27));
FA_ff_1179:FAff port map(x=>p(27)(27),y=>p(28)(27),Cin=>p(29)(27),clock=>clock,reset=>reset,s=>p(146)(27),cout=>p(147)(28));
FA_ff_1180:FAff port map(x=>p(27)(28),y=>p(28)(28),Cin=>p(29)(28),clock=>clock,reset=>reset,s=>p(146)(28),cout=>p(147)(29));
FA_ff_1181:FAff port map(x=>p(27)(29),y=>p(28)(29),Cin=>p(29)(29),clock=>clock,reset=>reset,s=>p(146)(29),cout=>p(147)(30));
FA_ff_1182:FAff port map(x=>p(27)(30),y=>p(28)(30),Cin=>p(29)(30),clock=>clock,reset=>reset,s=>p(146)(30),cout=>p(147)(31));
FA_ff_1183:FAff port map(x=>p(27)(31),y=>p(28)(31),Cin=>p(29)(31),clock=>clock,reset=>reset,s=>p(146)(31),cout=>p(147)(32));
FA_ff_1184:FAff port map(x=>p(27)(32),y=>p(28)(32),Cin=>p(29)(32),clock=>clock,reset=>reset,s=>p(146)(32),cout=>p(147)(33));
FA_ff_1185:FAff port map(x=>p(27)(33),y=>p(28)(33),Cin=>p(29)(33),clock=>clock,reset=>reset,s=>p(146)(33),cout=>p(147)(34));
FA_ff_1186:FAff port map(x=>p(27)(34),y=>p(28)(34),Cin=>p(29)(34),clock=>clock,reset=>reset,s=>p(146)(34),cout=>p(147)(35));
FA_ff_1187:FAff port map(x=>p(27)(35),y=>p(28)(35),Cin=>p(29)(35),clock=>clock,reset=>reset,s=>p(146)(35),cout=>p(147)(36));
FA_ff_1188:FAff port map(x=>p(27)(36),y=>p(28)(36),Cin=>p(29)(36),clock=>clock,reset=>reset,s=>p(146)(36),cout=>p(147)(37));
FA_ff_1189:FAff port map(x=>p(27)(37),y=>p(28)(37),Cin=>p(29)(37),clock=>clock,reset=>reset,s=>p(146)(37),cout=>p(147)(38));
FA_ff_1190:FAff port map(x=>p(27)(38),y=>p(28)(38),Cin=>p(29)(38),clock=>clock,reset=>reset,s=>p(146)(38),cout=>p(147)(39));
FA_ff_1191:FAff port map(x=>p(27)(39),y=>p(28)(39),Cin=>p(29)(39),clock=>clock,reset=>reset,s=>p(146)(39),cout=>p(147)(40));
FA_ff_1192:FAff port map(x=>p(27)(40),y=>p(28)(40),Cin=>p(29)(40),clock=>clock,reset=>reset,s=>p(146)(40),cout=>p(147)(41));
FA_ff_1193:FAff port map(x=>p(27)(41),y=>p(28)(41),Cin=>p(29)(41),clock=>clock,reset=>reset,s=>p(146)(41),cout=>p(147)(42));
FA_ff_1194:FAff port map(x=>p(27)(42),y=>p(28)(42),Cin=>p(29)(42),clock=>clock,reset=>reset,s=>p(146)(42),cout=>p(147)(43));
FA_ff_1195:FAff port map(x=>p(27)(43),y=>p(28)(43),Cin=>p(29)(43),clock=>clock,reset=>reset,s=>p(146)(43),cout=>p(147)(44));
FA_ff_1196:FAff port map(x=>p(27)(44),y=>p(28)(44),Cin=>p(29)(44),clock=>clock,reset=>reset,s=>p(146)(44),cout=>p(147)(45));
FA_ff_1197:FAff port map(x=>p(27)(45),y=>p(28)(45),Cin=>p(29)(45),clock=>clock,reset=>reset,s=>p(146)(45),cout=>p(147)(46));
FA_ff_1198:FAff port map(x=>p(27)(46),y=>p(28)(46),Cin=>p(29)(46),clock=>clock,reset=>reset,s=>p(146)(46),cout=>p(147)(47));
FA_ff_1199:FAff port map(x=>p(27)(47),y=>p(28)(47),Cin=>p(29)(47),clock=>clock,reset=>reset,s=>p(146)(47),cout=>p(147)(48));
FA_ff_1200:FAff port map(x=>p(27)(48),y=>p(28)(48),Cin=>p(29)(48),clock=>clock,reset=>reset,s=>p(146)(48),cout=>p(147)(49));
FA_ff_1201:FAff port map(x=>p(27)(49),y=>p(28)(49),Cin=>p(29)(49),clock=>clock,reset=>reset,s=>p(146)(49),cout=>p(147)(50));
FA_ff_1202:FAff port map(x=>p(27)(50),y=>p(28)(50),Cin=>p(29)(50),clock=>clock,reset=>reset,s=>p(146)(50),cout=>p(147)(51));
FA_ff_1203:FAff port map(x=>p(27)(51),y=>p(28)(51),Cin=>p(29)(51),clock=>clock,reset=>reset,s=>p(146)(51),cout=>p(147)(52));
FA_ff_1204:FAff port map(x=>p(27)(52),y=>p(28)(52),Cin=>p(29)(52),clock=>clock,reset=>reset,s=>p(146)(52),cout=>p(147)(53));
FA_ff_1205:FAff port map(x=>p(27)(53),y=>p(28)(53),Cin=>p(29)(53),clock=>clock,reset=>reset,s=>p(146)(53),cout=>p(147)(54));
FA_ff_1206:FAff port map(x=>p(27)(54),y=>p(28)(54),Cin=>p(29)(54),clock=>clock,reset=>reset,s=>p(146)(54),cout=>p(147)(55));
FA_ff_1207:FAff port map(x=>p(27)(55),y=>p(28)(55),Cin=>p(29)(55),clock=>clock,reset=>reset,s=>p(146)(55),cout=>p(147)(56));
FA_ff_1208:FAff port map(x=>p(27)(56),y=>p(28)(56),Cin=>p(29)(56),clock=>clock,reset=>reset,s=>p(146)(56),cout=>p(147)(57));
FA_ff_1209:FAff port map(x=>p(27)(57),y=>p(28)(57),Cin=>p(29)(57),clock=>clock,reset=>reset,s=>p(146)(57),cout=>p(147)(58));
FA_ff_1210:FAff port map(x=>p(27)(58),y=>p(28)(58),Cin=>p(29)(58),clock=>clock,reset=>reset,s=>p(146)(58),cout=>p(147)(59));
FA_ff_1211:FAff port map(x=>p(27)(59),y=>p(28)(59),Cin=>p(29)(59),clock=>clock,reset=>reset,s=>p(146)(59),cout=>p(147)(60));
FA_ff_1212:FAff port map(x=>p(27)(60),y=>p(28)(60),Cin=>p(29)(60),clock=>clock,reset=>reset,s=>p(146)(60),cout=>p(147)(61));
FA_ff_1213:FAff port map(x=>p(27)(61),y=>p(28)(61),Cin=>p(29)(61),clock=>clock,reset=>reset,s=>p(146)(61),cout=>p(147)(62));
FA_ff_1214:FAff port map(x=>p(27)(62),y=>p(28)(62),Cin=>p(29)(62),clock=>clock,reset=>reset,s=>p(146)(62),cout=>p(147)(63));
FA_ff_1215:FAff port map(x=>p(27)(63),y=>p(28)(63),Cin=>p(29)(63),clock=>clock,reset=>reset,s=>p(146)(63),cout=>p(147)(64));
FA_ff_1216:FAff port map(x=>p(27)(64),y=>p(28)(64),Cin=>p(29)(64),clock=>clock,reset=>reset,s=>p(146)(64),cout=>p(147)(65));
FA_ff_1217:FAff port map(x=>p(27)(65),y=>p(28)(65),Cin=>p(29)(65),clock=>clock,reset=>reset,s=>p(146)(65),cout=>p(147)(66));
FA_ff_1218:FAff port map(x=>p(27)(66),y=>p(28)(66),Cin=>p(29)(66),clock=>clock,reset=>reset,s=>p(146)(66),cout=>p(147)(67));
FA_ff_1219:FAff port map(x=>p(27)(67),y=>p(28)(67),Cin=>p(29)(67),clock=>clock,reset=>reset,s=>p(146)(67),cout=>p(147)(68));
FA_ff_1220:FAff port map(x=>p(27)(68),y=>p(28)(68),Cin=>p(29)(68),clock=>clock,reset=>reset,s=>p(146)(68),cout=>p(147)(69));
FA_ff_1221:FAff port map(x=>p(27)(69),y=>p(28)(69),Cin=>p(29)(69),clock=>clock,reset=>reset,s=>p(146)(69),cout=>p(147)(70));
FA_ff_1222:FAff port map(x=>p(27)(70),y=>p(28)(70),Cin=>p(29)(70),clock=>clock,reset=>reset,s=>p(146)(70),cout=>p(147)(71));
FA_ff_1223:FAff port map(x=>p(27)(71),y=>p(28)(71),Cin=>p(29)(71),clock=>clock,reset=>reset,s=>p(146)(71),cout=>p(147)(72));
FA_ff_1224:FAff port map(x=>p(27)(72),y=>p(28)(72),Cin=>p(29)(72),clock=>clock,reset=>reset,s=>p(146)(72),cout=>p(147)(73));
FA_ff_1225:FAff port map(x=>p(27)(73),y=>p(28)(73),Cin=>p(29)(73),clock=>clock,reset=>reset,s=>p(146)(73),cout=>p(147)(74));
FA_ff_1226:FAff port map(x=>p(27)(74),y=>p(28)(74),Cin=>p(29)(74),clock=>clock,reset=>reset,s=>p(146)(74),cout=>p(147)(75));
FA_ff_1227:FAff port map(x=>p(27)(75),y=>p(28)(75),Cin=>p(29)(75),clock=>clock,reset=>reset,s=>p(146)(75),cout=>p(147)(76));
FA_ff_1228:FAff port map(x=>p(27)(76),y=>p(28)(76),Cin=>p(29)(76),clock=>clock,reset=>reset,s=>p(146)(76),cout=>p(147)(77));
FA_ff_1229:FAff port map(x=>p(27)(77),y=>p(28)(77),Cin=>p(29)(77),clock=>clock,reset=>reset,s=>p(146)(77),cout=>p(147)(78));
FA_ff_1230:FAff port map(x=>p(27)(78),y=>p(28)(78),Cin=>p(29)(78),clock=>clock,reset=>reset,s=>p(146)(78),cout=>p(147)(79));
FA_ff_1231:FAff port map(x=>p(27)(79),y=>p(28)(79),Cin=>p(29)(79),clock=>clock,reset=>reset,s=>p(146)(79),cout=>p(147)(80));
FA_ff_1232:FAff port map(x=>p(27)(80),y=>p(28)(80),Cin=>p(29)(80),clock=>clock,reset=>reset,s=>p(146)(80),cout=>p(147)(81));
FA_ff_1233:FAff port map(x=>p(27)(81),y=>p(28)(81),Cin=>p(29)(81),clock=>clock,reset=>reset,s=>p(146)(81),cout=>p(147)(82));
FA_ff_1234:FAff port map(x=>p(27)(82),y=>p(28)(82),Cin=>p(29)(82),clock=>clock,reset=>reset,s=>p(146)(82),cout=>p(147)(83));
FA_ff_1235:FAff port map(x=>p(27)(83),y=>p(28)(83),Cin=>p(29)(83),clock=>clock,reset=>reset,s=>p(146)(83),cout=>p(147)(84));
FA_ff_1236:FAff port map(x=>p(27)(84),y=>p(28)(84),Cin=>p(29)(84),clock=>clock,reset=>reset,s=>p(146)(84),cout=>p(147)(85));
FA_ff_1237:FAff port map(x=>p(27)(85),y=>p(28)(85),Cin=>p(29)(85),clock=>clock,reset=>reset,s=>p(146)(85),cout=>p(147)(86));
FA_ff_1238:FAff port map(x=>p(27)(86),y=>p(28)(86),Cin=>p(29)(86),clock=>clock,reset=>reset,s=>p(146)(86),cout=>p(147)(87));
FA_ff_1239:FAff port map(x=>p(27)(87),y=>p(28)(87),Cin=>p(29)(87),clock=>clock,reset=>reset,s=>p(146)(87),cout=>p(147)(88));
FA_ff_1240:FAff port map(x=>p(27)(88),y=>p(28)(88),Cin=>p(29)(88),clock=>clock,reset=>reset,s=>p(146)(88),cout=>p(147)(89));
FA_ff_1241:FAff port map(x=>p(27)(89),y=>p(28)(89),Cin=>p(29)(89),clock=>clock,reset=>reset,s=>p(146)(89),cout=>p(147)(90));
FA_ff_1242:FAff port map(x=>p(27)(90),y=>p(28)(90),Cin=>p(29)(90),clock=>clock,reset=>reset,s=>p(146)(90),cout=>p(147)(91));
FA_ff_1243:FAff port map(x=>p(27)(91),y=>p(28)(91),Cin=>p(29)(91),clock=>clock,reset=>reset,s=>p(146)(91),cout=>p(147)(92));
FA_ff_1244:FAff port map(x=>p(27)(92),y=>p(28)(92),Cin=>p(29)(92),clock=>clock,reset=>reset,s=>p(146)(92),cout=>p(147)(93));
FA_ff_1245:FAff port map(x=>p(27)(93),y=>p(28)(93),Cin=>p(29)(93),clock=>clock,reset=>reset,s=>p(146)(93),cout=>p(147)(94));
FA_ff_1246:FAff port map(x=>p(27)(94),y=>p(28)(94),Cin=>p(29)(94),clock=>clock,reset=>reset,s=>p(146)(94),cout=>p(147)(95));
FA_ff_1247:FAff port map(x=>p(27)(95),y=>p(28)(95),Cin=>p(29)(95),clock=>clock,reset=>reset,s=>p(146)(95),cout=>p(147)(96));
FA_ff_1248:FAff port map(x=>p(27)(96),y=>p(28)(96),Cin=>p(29)(96),clock=>clock,reset=>reset,s=>p(146)(96),cout=>p(147)(97));
FA_ff_1249:FAff port map(x=>p(27)(97),y=>p(28)(97),Cin=>p(29)(97),clock=>clock,reset=>reset,s=>p(146)(97),cout=>p(147)(98));
FA_ff_1250:FAff port map(x=>p(27)(98),y=>p(28)(98),Cin=>p(29)(98),clock=>clock,reset=>reset,s=>p(146)(98),cout=>p(147)(99));
FA_ff_1251:FAff port map(x=>p(27)(99),y=>p(28)(99),Cin=>p(29)(99),clock=>clock,reset=>reset,s=>p(146)(99),cout=>p(147)(100));
FA_ff_1252:FAff port map(x=>p(27)(100),y=>p(28)(100),Cin=>p(29)(100),clock=>clock,reset=>reset,s=>p(146)(100),cout=>p(147)(101));
FA_ff_1253:FAff port map(x=>p(27)(101),y=>p(28)(101),Cin=>p(29)(101),clock=>clock,reset=>reset,s=>p(146)(101),cout=>p(147)(102));
FA_ff_1254:FAff port map(x=>p(27)(102),y=>p(28)(102),Cin=>p(29)(102),clock=>clock,reset=>reset,s=>p(146)(102),cout=>p(147)(103));
FA_ff_1255:FAff port map(x=>p(27)(103),y=>p(28)(103),Cin=>p(29)(103),clock=>clock,reset=>reset,s=>p(146)(103),cout=>p(147)(104));
FA_ff_1256:FAff port map(x=>p(27)(104),y=>p(28)(104),Cin=>p(29)(104),clock=>clock,reset=>reset,s=>p(146)(104),cout=>p(147)(105));
FA_ff_1257:FAff port map(x=>p(27)(105),y=>p(28)(105),Cin=>p(29)(105),clock=>clock,reset=>reset,s=>p(146)(105),cout=>p(147)(106));
FA_ff_1258:FAff port map(x=>p(27)(106),y=>p(28)(106),Cin=>p(29)(106),clock=>clock,reset=>reset,s=>p(146)(106),cout=>p(147)(107));
FA_ff_1259:FAff port map(x=>p(27)(107),y=>p(28)(107),Cin=>p(29)(107),clock=>clock,reset=>reset,s=>p(146)(107),cout=>p(147)(108));
FA_ff_1260:FAff port map(x=>p(27)(108),y=>p(28)(108),Cin=>p(29)(108),clock=>clock,reset=>reset,s=>p(146)(108),cout=>p(147)(109));
FA_ff_1261:FAff port map(x=>p(27)(109),y=>p(28)(109),Cin=>p(29)(109),clock=>clock,reset=>reset,s=>p(146)(109),cout=>p(147)(110));
FA_ff_1262:FAff port map(x=>p(27)(110),y=>p(28)(110),Cin=>p(29)(110),clock=>clock,reset=>reset,s=>p(146)(110),cout=>p(147)(111));
FA_ff_1263:FAff port map(x=>p(27)(111),y=>p(28)(111),Cin=>p(29)(111),clock=>clock,reset=>reset,s=>p(146)(111),cout=>p(147)(112));
FA_ff_1264:FAff port map(x=>p(27)(112),y=>p(28)(112),Cin=>p(29)(112),clock=>clock,reset=>reset,s=>p(146)(112),cout=>p(147)(113));
FA_ff_1265:FAff port map(x=>p(27)(113),y=>p(28)(113),Cin=>p(29)(113),clock=>clock,reset=>reset,s=>p(146)(113),cout=>p(147)(114));
FA_ff_1266:FAff port map(x=>p(27)(114),y=>p(28)(114),Cin=>p(29)(114),clock=>clock,reset=>reset,s=>p(146)(114),cout=>p(147)(115));
FA_ff_1267:FAff port map(x=>p(27)(115),y=>p(28)(115),Cin=>p(29)(115),clock=>clock,reset=>reset,s=>p(146)(115),cout=>p(147)(116));
FA_ff_1268:FAff port map(x=>p(27)(116),y=>p(28)(116),Cin=>p(29)(116),clock=>clock,reset=>reset,s=>p(146)(116),cout=>p(147)(117));
FA_ff_1269:FAff port map(x=>p(27)(117),y=>p(28)(117),Cin=>p(29)(117),clock=>clock,reset=>reset,s=>p(146)(117),cout=>p(147)(118));
FA_ff_1270:FAff port map(x=>p(27)(118),y=>p(28)(118),Cin=>p(29)(118),clock=>clock,reset=>reset,s=>p(146)(118),cout=>p(147)(119));
FA_ff_1271:FAff port map(x=>p(27)(119),y=>p(28)(119),Cin=>p(29)(119),clock=>clock,reset=>reset,s=>p(146)(119),cout=>p(147)(120));
FA_ff_1272:FAff port map(x=>p(27)(120),y=>p(28)(120),Cin=>p(29)(120),clock=>clock,reset=>reset,s=>p(146)(120),cout=>p(147)(121));
FA_ff_1273:FAff port map(x=>p(27)(121),y=>p(28)(121),Cin=>p(29)(121),clock=>clock,reset=>reset,s=>p(146)(121),cout=>p(147)(122));
FA_ff_1274:FAff port map(x=>p(27)(122),y=>p(28)(122),Cin=>p(29)(122),clock=>clock,reset=>reset,s=>p(146)(122),cout=>p(147)(123));
FA_ff_1275:FAff port map(x=>p(27)(123),y=>p(28)(123),Cin=>p(29)(123),clock=>clock,reset=>reset,s=>p(146)(123),cout=>p(147)(124));
FA_ff_1276:FAff port map(x=>p(27)(124),y=>p(28)(124),Cin=>p(29)(124),clock=>clock,reset=>reset,s=>p(146)(124),cout=>p(147)(125));
FA_ff_1277:FAff port map(x=>p(27)(125),y=>p(28)(125),Cin=>p(29)(125),clock=>clock,reset=>reset,s=>p(146)(125),cout=>p(147)(126));
FA_ff_1278:FAff port map(x=>p(27)(126),y=>p(28)(126),Cin=>p(29)(126),clock=>clock,reset=>reset,s=>p(146)(126),cout=>p(147)(127));
FA_ff_1279:FAff port map(x=>p(27)(127),y=>p(28)(127),Cin=>p(29)(127),clock=>clock,reset=>reset,s=>p(146)(127),cout=>p(147)(128));
FA_ff_1280:FAff port map(x=>p(30)(0),y=>p(31)(0),Cin=>p(32)(0),clock=>clock,reset=>reset,s=>p(148)(0),cout=>p(149)(1));
FA_ff_1281:FAff port map(x=>p(30)(1),y=>p(31)(1),Cin=>p(32)(1),clock=>clock,reset=>reset,s=>p(148)(1),cout=>p(149)(2));
FA_ff_1282:FAff port map(x=>p(30)(2),y=>p(31)(2),Cin=>p(32)(2),clock=>clock,reset=>reset,s=>p(148)(2),cout=>p(149)(3));
FA_ff_1283:FAff port map(x=>p(30)(3),y=>p(31)(3),Cin=>p(32)(3),clock=>clock,reset=>reset,s=>p(148)(3),cout=>p(149)(4));
FA_ff_1284:FAff port map(x=>p(30)(4),y=>p(31)(4),Cin=>p(32)(4),clock=>clock,reset=>reset,s=>p(148)(4),cout=>p(149)(5));
FA_ff_1285:FAff port map(x=>p(30)(5),y=>p(31)(5),Cin=>p(32)(5),clock=>clock,reset=>reset,s=>p(148)(5),cout=>p(149)(6));
FA_ff_1286:FAff port map(x=>p(30)(6),y=>p(31)(6),Cin=>p(32)(6),clock=>clock,reset=>reset,s=>p(148)(6),cout=>p(149)(7));
FA_ff_1287:FAff port map(x=>p(30)(7),y=>p(31)(7),Cin=>p(32)(7),clock=>clock,reset=>reset,s=>p(148)(7),cout=>p(149)(8));
FA_ff_1288:FAff port map(x=>p(30)(8),y=>p(31)(8),Cin=>p(32)(8),clock=>clock,reset=>reset,s=>p(148)(8),cout=>p(149)(9));
FA_ff_1289:FAff port map(x=>p(30)(9),y=>p(31)(9),Cin=>p(32)(9),clock=>clock,reset=>reset,s=>p(148)(9),cout=>p(149)(10));
FA_ff_1290:FAff port map(x=>p(30)(10),y=>p(31)(10),Cin=>p(32)(10),clock=>clock,reset=>reset,s=>p(148)(10),cout=>p(149)(11));
FA_ff_1291:FAff port map(x=>p(30)(11),y=>p(31)(11),Cin=>p(32)(11),clock=>clock,reset=>reset,s=>p(148)(11),cout=>p(149)(12));
FA_ff_1292:FAff port map(x=>p(30)(12),y=>p(31)(12),Cin=>p(32)(12),clock=>clock,reset=>reset,s=>p(148)(12),cout=>p(149)(13));
FA_ff_1293:FAff port map(x=>p(30)(13),y=>p(31)(13),Cin=>p(32)(13),clock=>clock,reset=>reset,s=>p(148)(13),cout=>p(149)(14));
FA_ff_1294:FAff port map(x=>p(30)(14),y=>p(31)(14),Cin=>p(32)(14),clock=>clock,reset=>reset,s=>p(148)(14),cout=>p(149)(15));
FA_ff_1295:FAff port map(x=>p(30)(15),y=>p(31)(15),Cin=>p(32)(15),clock=>clock,reset=>reset,s=>p(148)(15),cout=>p(149)(16));
FA_ff_1296:FAff port map(x=>p(30)(16),y=>p(31)(16),Cin=>p(32)(16),clock=>clock,reset=>reset,s=>p(148)(16),cout=>p(149)(17));
FA_ff_1297:FAff port map(x=>p(30)(17),y=>p(31)(17),Cin=>p(32)(17),clock=>clock,reset=>reset,s=>p(148)(17),cout=>p(149)(18));
FA_ff_1298:FAff port map(x=>p(30)(18),y=>p(31)(18),Cin=>p(32)(18),clock=>clock,reset=>reset,s=>p(148)(18),cout=>p(149)(19));
FA_ff_1299:FAff port map(x=>p(30)(19),y=>p(31)(19),Cin=>p(32)(19),clock=>clock,reset=>reset,s=>p(148)(19),cout=>p(149)(20));
FA_ff_1300:FAff port map(x=>p(30)(20),y=>p(31)(20),Cin=>p(32)(20),clock=>clock,reset=>reset,s=>p(148)(20),cout=>p(149)(21));
FA_ff_1301:FAff port map(x=>p(30)(21),y=>p(31)(21),Cin=>p(32)(21),clock=>clock,reset=>reset,s=>p(148)(21),cout=>p(149)(22));
FA_ff_1302:FAff port map(x=>p(30)(22),y=>p(31)(22),Cin=>p(32)(22),clock=>clock,reset=>reset,s=>p(148)(22),cout=>p(149)(23));
FA_ff_1303:FAff port map(x=>p(30)(23),y=>p(31)(23),Cin=>p(32)(23),clock=>clock,reset=>reset,s=>p(148)(23),cout=>p(149)(24));
FA_ff_1304:FAff port map(x=>p(30)(24),y=>p(31)(24),Cin=>p(32)(24),clock=>clock,reset=>reset,s=>p(148)(24),cout=>p(149)(25));
FA_ff_1305:FAff port map(x=>p(30)(25),y=>p(31)(25),Cin=>p(32)(25),clock=>clock,reset=>reset,s=>p(148)(25),cout=>p(149)(26));
FA_ff_1306:FAff port map(x=>p(30)(26),y=>p(31)(26),Cin=>p(32)(26),clock=>clock,reset=>reset,s=>p(148)(26),cout=>p(149)(27));
FA_ff_1307:FAff port map(x=>p(30)(27),y=>p(31)(27),Cin=>p(32)(27),clock=>clock,reset=>reset,s=>p(148)(27),cout=>p(149)(28));
FA_ff_1308:FAff port map(x=>p(30)(28),y=>p(31)(28),Cin=>p(32)(28),clock=>clock,reset=>reset,s=>p(148)(28),cout=>p(149)(29));
FA_ff_1309:FAff port map(x=>p(30)(29),y=>p(31)(29),Cin=>p(32)(29),clock=>clock,reset=>reset,s=>p(148)(29),cout=>p(149)(30));
FA_ff_1310:FAff port map(x=>p(30)(30),y=>p(31)(30),Cin=>p(32)(30),clock=>clock,reset=>reset,s=>p(148)(30),cout=>p(149)(31));
FA_ff_1311:FAff port map(x=>p(30)(31),y=>p(31)(31),Cin=>p(32)(31),clock=>clock,reset=>reset,s=>p(148)(31),cout=>p(149)(32));
FA_ff_1312:FAff port map(x=>p(30)(32),y=>p(31)(32),Cin=>p(32)(32),clock=>clock,reset=>reset,s=>p(148)(32),cout=>p(149)(33));
FA_ff_1313:FAff port map(x=>p(30)(33),y=>p(31)(33),Cin=>p(32)(33),clock=>clock,reset=>reset,s=>p(148)(33),cout=>p(149)(34));
FA_ff_1314:FAff port map(x=>p(30)(34),y=>p(31)(34),Cin=>p(32)(34),clock=>clock,reset=>reset,s=>p(148)(34),cout=>p(149)(35));
FA_ff_1315:FAff port map(x=>p(30)(35),y=>p(31)(35),Cin=>p(32)(35),clock=>clock,reset=>reset,s=>p(148)(35),cout=>p(149)(36));
FA_ff_1316:FAff port map(x=>p(30)(36),y=>p(31)(36),Cin=>p(32)(36),clock=>clock,reset=>reset,s=>p(148)(36),cout=>p(149)(37));
FA_ff_1317:FAff port map(x=>p(30)(37),y=>p(31)(37),Cin=>p(32)(37),clock=>clock,reset=>reset,s=>p(148)(37),cout=>p(149)(38));
FA_ff_1318:FAff port map(x=>p(30)(38),y=>p(31)(38),Cin=>p(32)(38),clock=>clock,reset=>reset,s=>p(148)(38),cout=>p(149)(39));
FA_ff_1319:FAff port map(x=>p(30)(39),y=>p(31)(39),Cin=>p(32)(39),clock=>clock,reset=>reset,s=>p(148)(39),cout=>p(149)(40));
FA_ff_1320:FAff port map(x=>p(30)(40),y=>p(31)(40),Cin=>p(32)(40),clock=>clock,reset=>reset,s=>p(148)(40),cout=>p(149)(41));
FA_ff_1321:FAff port map(x=>p(30)(41),y=>p(31)(41),Cin=>p(32)(41),clock=>clock,reset=>reset,s=>p(148)(41),cout=>p(149)(42));
FA_ff_1322:FAff port map(x=>p(30)(42),y=>p(31)(42),Cin=>p(32)(42),clock=>clock,reset=>reset,s=>p(148)(42),cout=>p(149)(43));
FA_ff_1323:FAff port map(x=>p(30)(43),y=>p(31)(43),Cin=>p(32)(43),clock=>clock,reset=>reset,s=>p(148)(43),cout=>p(149)(44));
FA_ff_1324:FAff port map(x=>p(30)(44),y=>p(31)(44),Cin=>p(32)(44),clock=>clock,reset=>reset,s=>p(148)(44),cout=>p(149)(45));
FA_ff_1325:FAff port map(x=>p(30)(45),y=>p(31)(45),Cin=>p(32)(45),clock=>clock,reset=>reset,s=>p(148)(45),cout=>p(149)(46));
FA_ff_1326:FAff port map(x=>p(30)(46),y=>p(31)(46),Cin=>p(32)(46),clock=>clock,reset=>reset,s=>p(148)(46),cout=>p(149)(47));
FA_ff_1327:FAff port map(x=>p(30)(47),y=>p(31)(47),Cin=>p(32)(47),clock=>clock,reset=>reset,s=>p(148)(47),cout=>p(149)(48));
FA_ff_1328:FAff port map(x=>p(30)(48),y=>p(31)(48),Cin=>p(32)(48),clock=>clock,reset=>reset,s=>p(148)(48),cout=>p(149)(49));
FA_ff_1329:FAff port map(x=>p(30)(49),y=>p(31)(49),Cin=>p(32)(49),clock=>clock,reset=>reset,s=>p(148)(49),cout=>p(149)(50));
FA_ff_1330:FAff port map(x=>p(30)(50),y=>p(31)(50),Cin=>p(32)(50),clock=>clock,reset=>reset,s=>p(148)(50),cout=>p(149)(51));
FA_ff_1331:FAff port map(x=>p(30)(51),y=>p(31)(51),Cin=>p(32)(51),clock=>clock,reset=>reset,s=>p(148)(51),cout=>p(149)(52));
FA_ff_1332:FAff port map(x=>p(30)(52),y=>p(31)(52),Cin=>p(32)(52),clock=>clock,reset=>reset,s=>p(148)(52),cout=>p(149)(53));
FA_ff_1333:FAff port map(x=>p(30)(53),y=>p(31)(53),Cin=>p(32)(53),clock=>clock,reset=>reset,s=>p(148)(53),cout=>p(149)(54));
FA_ff_1334:FAff port map(x=>p(30)(54),y=>p(31)(54),Cin=>p(32)(54),clock=>clock,reset=>reset,s=>p(148)(54),cout=>p(149)(55));
FA_ff_1335:FAff port map(x=>p(30)(55),y=>p(31)(55),Cin=>p(32)(55),clock=>clock,reset=>reset,s=>p(148)(55),cout=>p(149)(56));
FA_ff_1336:FAff port map(x=>p(30)(56),y=>p(31)(56),Cin=>p(32)(56),clock=>clock,reset=>reset,s=>p(148)(56),cout=>p(149)(57));
FA_ff_1337:FAff port map(x=>p(30)(57),y=>p(31)(57),Cin=>p(32)(57),clock=>clock,reset=>reset,s=>p(148)(57),cout=>p(149)(58));
FA_ff_1338:FAff port map(x=>p(30)(58),y=>p(31)(58),Cin=>p(32)(58),clock=>clock,reset=>reset,s=>p(148)(58),cout=>p(149)(59));
FA_ff_1339:FAff port map(x=>p(30)(59),y=>p(31)(59),Cin=>p(32)(59),clock=>clock,reset=>reset,s=>p(148)(59),cout=>p(149)(60));
FA_ff_1340:FAff port map(x=>p(30)(60),y=>p(31)(60),Cin=>p(32)(60),clock=>clock,reset=>reset,s=>p(148)(60),cout=>p(149)(61));
FA_ff_1341:FAff port map(x=>p(30)(61),y=>p(31)(61),Cin=>p(32)(61),clock=>clock,reset=>reset,s=>p(148)(61),cout=>p(149)(62));
FA_ff_1342:FAff port map(x=>p(30)(62),y=>p(31)(62),Cin=>p(32)(62),clock=>clock,reset=>reset,s=>p(148)(62),cout=>p(149)(63));
FA_ff_1343:FAff port map(x=>p(30)(63),y=>p(31)(63),Cin=>p(32)(63),clock=>clock,reset=>reset,s=>p(148)(63),cout=>p(149)(64));
FA_ff_1344:FAff port map(x=>p(30)(64),y=>p(31)(64),Cin=>p(32)(64),clock=>clock,reset=>reset,s=>p(148)(64),cout=>p(149)(65));
FA_ff_1345:FAff port map(x=>p(30)(65),y=>p(31)(65),Cin=>p(32)(65),clock=>clock,reset=>reset,s=>p(148)(65),cout=>p(149)(66));
FA_ff_1346:FAff port map(x=>p(30)(66),y=>p(31)(66),Cin=>p(32)(66),clock=>clock,reset=>reset,s=>p(148)(66),cout=>p(149)(67));
FA_ff_1347:FAff port map(x=>p(30)(67),y=>p(31)(67),Cin=>p(32)(67),clock=>clock,reset=>reset,s=>p(148)(67),cout=>p(149)(68));
FA_ff_1348:FAff port map(x=>p(30)(68),y=>p(31)(68),Cin=>p(32)(68),clock=>clock,reset=>reset,s=>p(148)(68),cout=>p(149)(69));
FA_ff_1349:FAff port map(x=>p(30)(69),y=>p(31)(69),Cin=>p(32)(69),clock=>clock,reset=>reset,s=>p(148)(69),cout=>p(149)(70));
FA_ff_1350:FAff port map(x=>p(30)(70),y=>p(31)(70),Cin=>p(32)(70),clock=>clock,reset=>reset,s=>p(148)(70),cout=>p(149)(71));
FA_ff_1351:FAff port map(x=>p(30)(71),y=>p(31)(71),Cin=>p(32)(71),clock=>clock,reset=>reset,s=>p(148)(71),cout=>p(149)(72));
FA_ff_1352:FAff port map(x=>p(30)(72),y=>p(31)(72),Cin=>p(32)(72),clock=>clock,reset=>reset,s=>p(148)(72),cout=>p(149)(73));
FA_ff_1353:FAff port map(x=>p(30)(73),y=>p(31)(73),Cin=>p(32)(73),clock=>clock,reset=>reset,s=>p(148)(73),cout=>p(149)(74));
FA_ff_1354:FAff port map(x=>p(30)(74),y=>p(31)(74),Cin=>p(32)(74),clock=>clock,reset=>reset,s=>p(148)(74),cout=>p(149)(75));
FA_ff_1355:FAff port map(x=>p(30)(75),y=>p(31)(75),Cin=>p(32)(75),clock=>clock,reset=>reset,s=>p(148)(75),cout=>p(149)(76));
FA_ff_1356:FAff port map(x=>p(30)(76),y=>p(31)(76),Cin=>p(32)(76),clock=>clock,reset=>reset,s=>p(148)(76),cout=>p(149)(77));
FA_ff_1357:FAff port map(x=>p(30)(77),y=>p(31)(77),Cin=>p(32)(77),clock=>clock,reset=>reset,s=>p(148)(77),cout=>p(149)(78));
FA_ff_1358:FAff port map(x=>p(30)(78),y=>p(31)(78),Cin=>p(32)(78),clock=>clock,reset=>reset,s=>p(148)(78),cout=>p(149)(79));
FA_ff_1359:FAff port map(x=>p(30)(79),y=>p(31)(79),Cin=>p(32)(79),clock=>clock,reset=>reset,s=>p(148)(79),cout=>p(149)(80));
FA_ff_1360:FAff port map(x=>p(30)(80),y=>p(31)(80),Cin=>p(32)(80),clock=>clock,reset=>reset,s=>p(148)(80),cout=>p(149)(81));
FA_ff_1361:FAff port map(x=>p(30)(81),y=>p(31)(81),Cin=>p(32)(81),clock=>clock,reset=>reset,s=>p(148)(81),cout=>p(149)(82));
FA_ff_1362:FAff port map(x=>p(30)(82),y=>p(31)(82),Cin=>p(32)(82),clock=>clock,reset=>reset,s=>p(148)(82),cout=>p(149)(83));
FA_ff_1363:FAff port map(x=>p(30)(83),y=>p(31)(83),Cin=>p(32)(83),clock=>clock,reset=>reset,s=>p(148)(83),cout=>p(149)(84));
FA_ff_1364:FAff port map(x=>p(30)(84),y=>p(31)(84),Cin=>p(32)(84),clock=>clock,reset=>reset,s=>p(148)(84),cout=>p(149)(85));
FA_ff_1365:FAff port map(x=>p(30)(85),y=>p(31)(85),Cin=>p(32)(85),clock=>clock,reset=>reset,s=>p(148)(85),cout=>p(149)(86));
FA_ff_1366:FAff port map(x=>p(30)(86),y=>p(31)(86),Cin=>p(32)(86),clock=>clock,reset=>reset,s=>p(148)(86),cout=>p(149)(87));
FA_ff_1367:FAff port map(x=>p(30)(87),y=>p(31)(87),Cin=>p(32)(87),clock=>clock,reset=>reset,s=>p(148)(87),cout=>p(149)(88));
FA_ff_1368:FAff port map(x=>p(30)(88),y=>p(31)(88),Cin=>p(32)(88),clock=>clock,reset=>reset,s=>p(148)(88),cout=>p(149)(89));
FA_ff_1369:FAff port map(x=>p(30)(89),y=>p(31)(89),Cin=>p(32)(89),clock=>clock,reset=>reset,s=>p(148)(89),cout=>p(149)(90));
FA_ff_1370:FAff port map(x=>p(30)(90),y=>p(31)(90),Cin=>p(32)(90),clock=>clock,reset=>reset,s=>p(148)(90),cout=>p(149)(91));
FA_ff_1371:FAff port map(x=>p(30)(91),y=>p(31)(91),Cin=>p(32)(91),clock=>clock,reset=>reset,s=>p(148)(91),cout=>p(149)(92));
FA_ff_1372:FAff port map(x=>p(30)(92),y=>p(31)(92),Cin=>p(32)(92),clock=>clock,reset=>reset,s=>p(148)(92),cout=>p(149)(93));
FA_ff_1373:FAff port map(x=>p(30)(93),y=>p(31)(93),Cin=>p(32)(93),clock=>clock,reset=>reset,s=>p(148)(93),cout=>p(149)(94));
FA_ff_1374:FAff port map(x=>p(30)(94),y=>p(31)(94),Cin=>p(32)(94),clock=>clock,reset=>reset,s=>p(148)(94),cout=>p(149)(95));
FA_ff_1375:FAff port map(x=>p(30)(95),y=>p(31)(95),Cin=>p(32)(95),clock=>clock,reset=>reset,s=>p(148)(95),cout=>p(149)(96));
FA_ff_1376:FAff port map(x=>p(30)(96),y=>p(31)(96),Cin=>p(32)(96),clock=>clock,reset=>reset,s=>p(148)(96),cout=>p(149)(97));
FA_ff_1377:FAff port map(x=>p(30)(97),y=>p(31)(97),Cin=>p(32)(97),clock=>clock,reset=>reset,s=>p(148)(97),cout=>p(149)(98));
FA_ff_1378:FAff port map(x=>p(30)(98),y=>p(31)(98),Cin=>p(32)(98),clock=>clock,reset=>reset,s=>p(148)(98),cout=>p(149)(99));
FA_ff_1379:FAff port map(x=>p(30)(99),y=>p(31)(99),Cin=>p(32)(99),clock=>clock,reset=>reset,s=>p(148)(99),cout=>p(149)(100));
FA_ff_1380:FAff port map(x=>p(30)(100),y=>p(31)(100),Cin=>p(32)(100),clock=>clock,reset=>reset,s=>p(148)(100),cout=>p(149)(101));
FA_ff_1381:FAff port map(x=>p(30)(101),y=>p(31)(101),Cin=>p(32)(101),clock=>clock,reset=>reset,s=>p(148)(101),cout=>p(149)(102));
FA_ff_1382:FAff port map(x=>p(30)(102),y=>p(31)(102),Cin=>p(32)(102),clock=>clock,reset=>reset,s=>p(148)(102),cout=>p(149)(103));
FA_ff_1383:FAff port map(x=>p(30)(103),y=>p(31)(103),Cin=>p(32)(103),clock=>clock,reset=>reset,s=>p(148)(103),cout=>p(149)(104));
FA_ff_1384:FAff port map(x=>p(30)(104),y=>p(31)(104),Cin=>p(32)(104),clock=>clock,reset=>reset,s=>p(148)(104),cout=>p(149)(105));
FA_ff_1385:FAff port map(x=>p(30)(105),y=>p(31)(105),Cin=>p(32)(105),clock=>clock,reset=>reset,s=>p(148)(105),cout=>p(149)(106));
FA_ff_1386:FAff port map(x=>p(30)(106),y=>p(31)(106),Cin=>p(32)(106),clock=>clock,reset=>reset,s=>p(148)(106),cout=>p(149)(107));
FA_ff_1387:FAff port map(x=>p(30)(107),y=>p(31)(107),Cin=>p(32)(107),clock=>clock,reset=>reset,s=>p(148)(107),cout=>p(149)(108));
FA_ff_1388:FAff port map(x=>p(30)(108),y=>p(31)(108),Cin=>p(32)(108),clock=>clock,reset=>reset,s=>p(148)(108),cout=>p(149)(109));
FA_ff_1389:FAff port map(x=>p(30)(109),y=>p(31)(109),Cin=>p(32)(109),clock=>clock,reset=>reset,s=>p(148)(109),cout=>p(149)(110));
FA_ff_1390:FAff port map(x=>p(30)(110),y=>p(31)(110),Cin=>p(32)(110),clock=>clock,reset=>reset,s=>p(148)(110),cout=>p(149)(111));
FA_ff_1391:FAff port map(x=>p(30)(111),y=>p(31)(111),Cin=>p(32)(111),clock=>clock,reset=>reset,s=>p(148)(111),cout=>p(149)(112));
FA_ff_1392:FAff port map(x=>p(30)(112),y=>p(31)(112),Cin=>p(32)(112),clock=>clock,reset=>reset,s=>p(148)(112),cout=>p(149)(113));
FA_ff_1393:FAff port map(x=>p(30)(113),y=>p(31)(113),Cin=>p(32)(113),clock=>clock,reset=>reset,s=>p(148)(113),cout=>p(149)(114));
FA_ff_1394:FAff port map(x=>p(30)(114),y=>p(31)(114),Cin=>p(32)(114),clock=>clock,reset=>reset,s=>p(148)(114),cout=>p(149)(115));
FA_ff_1395:FAff port map(x=>p(30)(115),y=>p(31)(115),Cin=>p(32)(115),clock=>clock,reset=>reset,s=>p(148)(115),cout=>p(149)(116));
FA_ff_1396:FAff port map(x=>p(30)(116),y=>p(31)(116),Cin=>p(32)(116),clock=>clock,reset=>reset,s=>p(148)(116),cout=>p(149)(117));
FA_ff_1397:FAff port map(x=>p(30)(117),y=>p(31)(117),Cin=>p(32)(117),clock=>clock,reset=>reset,s=>p(148)(117),cout=>p(149)(118));
FA_ff_1398:FAff port map(x=>p(30)(118),y=>p(31)(118),Cin=>p(32)(118),clock=>clock,reset=>reset,s=>p(148)(118),cout=>p(149)(119));
FA_ff_1399:FAff port map(x=>p(30)(119),y=>p(31)(119),Cin=>p(32)(119),clock=>clock,reset=>reset,s=>p(148)(119),cout=>p(149)(120));
FA_ff_1400:FAff port map(x=>p(30)(120),y=>p(31)(120),Cin=>p(32)(120),clock=>clock,reset=>reset,s=>p(148)(120),cout=>p(149)(121));
FA_ff_1401:FAff port map(x=>p(30)(121),y=>p(31)(121),Cin=>p(32)(121),clock=>clock,reset=>reset,s=>p(148)(121),cout=>p(149)(122));
FA_ff_1402:FAff port map(x=>p(30)(122),y=>p(31)(122),Cin=>p(32)(122),clock=>clock,reset=>reset,s=>p(148)(122),cout=>p(149)(123));
FA_ff_1403:FAff port map(x=>p(30)(123),y=>p(31)(123),Cin=>p(32)(123),clock=>clock,reset=>reset,s=>p(148)(123),cout=>p(149)(124));
FA_ff_1404:FAff port map(x=>p(30)(124),y=>p(31)(124),Cin=>p(32)(124),clock=>clock,reset=>reset,s=>p(148)(124),cout=>p(149)(125));
FA_ff_1405:FAff port map(x=>p(30)(125),y=>p(31)(125),Cin=>p(32)(125),clock=>clock,reset=>reset,s=>p(148)(125),cout=>p(149)(126));
FA_ff_1406:FAff port map(x=>p(30)(126),y=>p(31)(126),Cin=>p(32)(126),clock=>clock,reset=>reset,s=>p(148)(126),cout=>p(149)(127));
FA_ff_1407:FAff port map(x=>p(30)(127),y=>p(31)(127),Cin=>p(32)(127),clock=>clock,reset=>reset,s=>p(148)(127),cout=>p(149)(128));
FA_ff_1408:FAff port map(x=>p(33)(0),y=>p(34)(0),Cin=>p(35)(0),clock=>clock,reset=>reset,s=>p(150)(0),cout=>p(151)(1));
FA_ff_1409:FAff port map(x=>p(33)(1),y=>p(34)(1),Cin=>p(35)(1),clock=>clock,reset=>reset,s=>p(150)(1),cout=>p(151)(2));
FA_ff_1410:FAff port map(x=>p(33)(2),y=>p(34)(2),Cin=>p(35)(2),clock=>clock,reset=>reset,s=>p(150)(2),cout=>p(151)(3));
FA_ff_1411:FAff port map(x=>p(33)(3),y=>p(34)(3),Cin=>p(35)(3),clock=>clock,reset=>reset,s=>p(150)(3),cout=>p(151)(4));
FA_ff_1412:FAff port map(x=>p(33)(4),y=>p(34)(4),Cin=>p(35)(4),clock=>clock,reset=>reset,s=>p(150)(4),cout=>p(151)(5));
FA_ff_1413:FAff port map(x=>p(33)(5),y=>p(34)(5),Cin=>p(35)(5),clock=>clock,reset=>reset,s=>p(150)(5),cout=>p(151)(6));
FA_ff_1414:FAff port map(x=>p(33)(6),y=>p(34)(6),Cin=>p(35)(6),clock=>clock,reset=>reset,s=>p(150)(6),cout=>p(151)(7));
FA_ff_1415:FAff port map(x=>p(33)(7),y=>p(34)(7),Cin=>p(35)(7),clock=>clock,reset=>reset,s=>p(150)(7),cout=>p(151)(8));
FA_ff_1416:FAff port map(x=>p(33)(8),y=>p(34)(8),Cin=>p(35)(8),clock=>clock,reset=>reset,s=>p(150)(8),cout=>p(151)(9));
FA_ff_1417:FAff port map(x=>p(33)(9),y=>p(34)(9),Cin=>p(35)(9),clock=>clock,reset=>reset,s=>p(150)(9),cout=>p(151)(10));
FA_ff_1418:FAff port map(x=>p(33)(10),y=>p(34)(10),Cin=>p(35)(10),clock=>clock,reset=>reset,s=>p(150)(10),cout=>p(151)(11));
FA_ff_1419:FAff port map(x=>p(33)(11),y=>p(34)(11),Cin=>p(35)(11),clock=>clock,reset=>reset,s=>p(150)(11),cout=>p(151)(12));
FA_ff_1420:FAff port map(x=>p(33)(12),y=>p(34)(12),Cin=>p(35)(12),clock=>clock,reset=>reset,s=>p(150)(12),cout=>p(151)(13));
FA_ff_1421:FAff port map(x=>p(33)(13),y=>p(34)(13),Cin=>p(35)(13),clock=>clock,reset=>reset,s=>p(150)(13),cout=>p(151)(14));
FA_ff_1422:FAff port map(x=>p(33)(14),y=>p(34)(14),Cin=>p(35)(14),clock=>clock,reset=>reset,s=>p(150)(14),cout=>p(151)(15));
FA_ff_1423:FAff port map(x=>p(33)(15),y=>p(34)(15),Cin=>p(35)(15),clock=>clock,reset=>reset,s=>p(150)(15),cout=>p(151)(16));
FA_ff_1424:FAff port map(x=>p(33)(16),y=>p(34)(16),Cin=>p(35)(16),clock=>clock,reset=>reset,s=>p(150)(16),cout=>p(151)(17));
FA_ff_1425:FAff port map(x=>p(33)(17),y=>p(34)(17),Cin=>p(35)(17),clock=>clock,reset=>reset,s=>p(150)(17),cout=>p(151)(18));
FA_ff_1426:FAff port map(x=>p(33)(18),y=>p(34)(18),Cin=>p(35)(18),clock=>clock,reset=>reset,s=>p(150)(18),cout=>p(151)(19));
FA_ff_1427:FAff port map(x=>p(33)(19),y=>p(34)(19),Cin=>p(35)(19),clock=>clock,reset=>reset,s=>p(150)(19),cout=>p(151)(20));
FA_ff_1428:FAff port map(x=>p(33)(20),y=>p(34)(20),Cin=>p(35)(20),clock=>clock,reset=>reset,s=>p(150)(20),cout=>p(151)(21));
FA_ff_1429:FAff port map(x=>p(33)(21),y=>p(34)(21),Cin=>p(35)(21),clock=>clock,reset=>reset,s=>p(150)(21),cout=>p(151)(22));
FA_ff_1430:FAff port map(x=>p(33)(22),y=>p(34)(22),Cin=>p(35)(22),clock=>clock,reset=>reset,s=>p(150)(22),cout=>p(151)(23));
FA_ff_1431:FAff port map(x=>p(33)(23),y=>p(34)(23),Cin=>p(35)(23),clock=>clock,reset=>reset,s=>p(150)(23),cout=>p(151)(24));
FA_ff_1432:FAff port map(x=>p(33)(24),y=>p(34)(24),Cin=>p(35)(24),clock=>clock,reset=>reset,s=>p(150)(24),cout=>p(151)(25));
FA_ff_1433:FAff port map(x=>p(33)(25),y=>p(34)(25),Cin=>p(35)(25),clock=>clock,reset=>reset,s=>p(150)(25),cout=>p(151)(26));
FA_ff_1434:FAff port map(x=>p(33)(26),y=>p(34)(26),Cin=>p(35)(26),clock=>clock,reset=>reset,s=>p(150)(26),cout=>p(151)(27));
FA_ff_1435:FAff port map(x=>p(33)(27),y=>p(34)(27),Cin=>p(35)(27),clock=>clock,reset=>reset,s=>p(150)(27),cout=>p(151)(28));
FA_ff_1436:FAff port map(x=>p(33)(28),y=>p(34)(28),Cin=>p(35)(28),clock=>clock,reset=>reset,s=>p(150)(28),cout=>p(151)(29));
FA_ff_1437:FAff port map(x=>p(33)(29),y=>p(34)(29),Cin=>p(35)(29),clock=>clock,reset=>reset,s=>p(150)(29),cout=>p(151)(30));
FA_ff_1438:FAff port map(x=>p(33)(30),y=>p(34)(30),Cin=>p(35)(30),clock=>clock,reset=>reset,s=>p(150)(30),cout=>p(151)(31));
FA_ff_1439:FAff port map(x=>p(33)(31),y=>p(34)(31),Cin=>p(35)(31),clock=>clock,reset=>reset,s=>p(150)(31),cout=>p(151)(32));
FA_ff_1440:FAff port map(x=>p(33)(32),y=>p(34)(32),Cin=>p(35)(32),clock=>clock,reset=>reset,s=>p(150)(32),cout=>p(151)(33));
FA_ff_1441:FAff port map(x=>p(33)(33),y=>p(34)(33),Cin=>p(35)(33),clock=>clock,reset=>reset,s=>p(150)(33),cout=>p(151)(34));
FA_ff_1442:FAff port map(x=>p(33)(34),y=>p(34)(34),Cin=>p(35)(34),clock=>clock,reset=>reset,s=>p(150)(34),cout=>p(151)(35));
FA_ff_1443:FAff port map(x=>p(33)(35),y=>p(34)(35),Cin=>p(35)(35),clock=>clock,reset=>reset,s=>p(150)(35),cout=>p(151)(36));
FA_ff_1444:FAff port map(x=>p(33)(36),y=>p(34)(36),Cin=>p(35)(36),clock=>clock,reset=>reset,s=>p(150)(36),cout=>p(151)(37));
FA_ff_1445:FAff port map(x=>p(33)(37),y=>p(34)(37),Cin=>p(35)(37),clock=>clock,reset=>reset,s=>p(150)(37),cout=>p(151)(38));
FA_ff_1446:FAff port map(x=>p(33)(38),y=>p(34)(38),Cin=>p(35)(38),clock=>clock,reset=>reset,s=>p(150)(38),cout=>p(151)(39));
FA_ff_1447:FAff port map(x=>p(33)(39),y=>p(34)(39),Cin=>p(35)(39),clock=>clock,reset=>reset,s=>p(150)(39),cout=>p(151)(40));
FA_ff_1448:FAff port map(x=>p(33)(40),y=>p(34)(40),Cin=>p(35)(40),clock=>clock,reset=>reset,s=>p(150)(40),cout=>p(151)(41));
FA_ff_1449:FAff port map(x=>p(33)(41),y=>p(34)(41),Cin=>p(35)(41),clock=>clock,reset=>reset,s=>p(150)(41),cout=>p(151)(42));
FA_ff_1450:FAff port map(x=>p(33)(42),y=>p(34)(42),Cin=>p(35)(42),clock=>clock,reset=>reset,s=>p(150)(42),cout=>p(151)(43));
FA_ff_1451:FAff port map(x=>p(33)(43),y=>p(34)(43),Cin=>p(35)(43),clock=>clock,reset=>reset,s=>p(150)(43),cout=>p(151)(44));
FA_ff_1452:FAff port map(x=>p(33)(44),y=>p(34)(44),Cin=>p(35)(44),clock=>clock,reset=>reset,s=>p(150)(44),cout=>p(151)(45));
FA_ff_1453:FAff port map(x=>p(33)(45),y=>p(34)(45),Cin=>p(35)(45),clock=>clock,reset=>reset,s=>p(150)(45),cout=>p(151)(46));
FA_ff_1454:FAff port map(x=>p(33)(46),y=>p(34)(46),Cin=>p(35)(46),clock=>clock,reset=>reset,s=>p(150)(46),cout=>p(151)(47));
FA_ff_1455:FAff port map(x=>p(33)(47),y=>p(34)(47),Cin=>p(35)(47),clock=>clock,reset=>reset,s=>p(150)(47),cout=>p(151)(48));
FA_ff_1456:FAff port map(x=>p(33)(48),y=>p(34)(48),Cin=>p(35)(48),clock=>clock,reset=>reset,s=>p(150)(48),cout=>p(151)(49));
FA_ff_1457:FAff port map(x=>p(33)(49),y=>p(34)(49),Cin=>p(35)(49),clock=>clock,reset=>reset,s=>p(150)(49),cout=>p(151)(50));
FA_ff_1458:FAff port map(x=>p(33)(50),y=>p(34)(50),Cin=>p(35)(50),clock=>clock,reset=>reset,s=>p(150)(50),cout=>p(151)(51));
FA_ff_1459:FAff port map(x=>p(33)(51),y=>p(34)(51),Cin=>p(35)(51),clock=>clock,reset=>reset,s=>p(150)(51),cout=>p(151)(52));
FA_ff_1460:FAff port map(x=>p(33)(52),y=>p(34)(52),Cin=>p(35)(52),clock=>clock,reset=>reset,s=>p(150)(52),cout=>p(151)(53));
FA_ff_1461:FAff port map(x=>p(33)(53),y=>p(34)(53),Cin=>p(35)(53),clock=>clock,reset=>reset,s=>p(150)(53),cout=>p(151)(54));
FA_ff_1462:FAff port map(x=>p(33)(54),y=>p(34)(54),Cin=>p(35)(54),clock=>clock,reset=>reset,s=>p(150)(54),cout=>p(151)(55));
FA_ff_1463:FAff port map(x=>p(33)(55),y=>p(34)(55),Cin=>p(35)(55),clock=>clock,reset=>reset,s=>p(150)(55),cout=>p(151)(56));
FA_ff_1464:FAff port map(x=>p(33)(56),y=>p(34)(56),Cin=>p(35)(56),clock=>clock,reset=>reset,s=>p(150)(56),cout=>p(151)(57));
FA_ff_1465:FAff port map(x=>p(33)(57),y=>p(34)(57),Cin=>p(35)(57),clock=>clock,reset=>reset,s=>p(150)(57),cout=>p(151)(58));
FA_ff_1466:FAff port map(x=>p(33)(58),y=>p(34)(58),Cin=>p(35)(58),clock=>clock,reset=>reset,s=>p(150)(58),cout=>p(151)(59));
FA_ff_1467:FAff port map(x=>p(33)(59),y=>p(34)(59),Cin=>p(35)(59),clock=>clock,reset=>reset,s=>p(150)(59),cout=>p(151)(60));
FA_ff_1468:FAff port map(x=>p(33)(60),y=>p(34)(60),Cin=>p(35)(60),clock=>clock,reset=>reset,s=>p(150)(60),cout=>p(151)(61));
FA_ff_1469:FAff port map(x=>p(33)(61),y=>p(34)(61),Cin=>p(35)(61),clock=>clock,reset=>reset,s=>p(150)(61),cout=>p(151)(62));
FA_ff_1470:FAff port map(x=>p(33)(62),y=>p(34)(62),Cin=>p(35)(62),clock=>clock,reset=>reset,s=>p(150)(62),cout=>p(151)(63));
FA_ff_1471:FAff port map(x=>p(33)(63),y=>p(34)(63),Cin=>p(35)(63),clock=>clock,reset=>reset,s=>p(150)(63),cout=>p(151)(64));
FA_ff_1472:FAff port map(x=>p(33)(64),y=>p(34)(64),Cin=>p(35)(64),clock=>clock,reset=>reset,s=>p(150)(64),cout=>p(151)(65));
FA_ff_1473:FAff port map(x=>p(33)(65),y=>p(34)(65),Cin=>p(35)(65),clock=>clock,reset=>reset,s=>p(150)(65),cout=>p(151)(66));
FA_ff_1474:FAff port map(x=>p(33)(66),y=>p(34)(66),Cin=>p(35)(66),clock=>clock,reset=>reset,s=>p(150)(66),cout=>p(151)(67));
FA_ff_1475:FAff port map(x=>p(33)(67),y=>p(34)(67),Cin=>p(35)(67),clock=>clock,reset=>reset,s=>p(150)(67),cout=>p(151)(68));
FA_ff_1476:FAff port map(x=>p(33)(68),y=>p(34)(68),Cin=>p(35)(68),clock=>clock,reset=>reset,s=>p(150)(68),cout=>p(151)(69));
FA_ff_1477:FAff port map(x=>p(33)(69),y=>p(34)(69),Cin=>p(35)(69),clock=>clock,reset=>reset,s=>p(150)(69),cout=>p(151)(70));
FA_ff_1478:FAff port map(x=>p(33)(70),y=>p(34)(70),Cin=>p(35)(70),clock=>clock,reset=>reset,s=>p(150)(70),cout=>p(151)(71));
FA_ff_1479:FAff port map(x=>p(33)(71),y=>p(34)(71),Cin=>p(35)(71),clock=>clock,reset=>reset,s=>p(150)(71),cout=>p(151)(72));
FA_ff_1480:FAff port map(x=>p(33)(72),y=>p(34)(72),Cin=>p(35)(72),clock=>clock,reset=>reset,s=>p(150)(72),cout=>p(151)(73));
FA_ff_1481:FAff port map(x=>p(33)(73),y=>p(34)(73),Cin=>p(35)(73),clock=>clock,reset=>reset,s=>p(150)(73),cout=>p(151)(74));
FA_ff_1482:FAff port map(x=>p(33)(74),y=>p(34)(74),Cin=>p(35)(74),clock=>clock,reset=>reset,s=>p(150)(74),cout=>p(151)(75));
FA_ff_1483:FAff port map(x=>p(33)(75),y=>p(34)(75),Cin=>p(35)(75),clock=>clock,reset=>reset,s=>p(150)(75),cout=>p(151)(76));
FA_ff_1484:FAff port map(x=>p(33)(76),y=>p(34)(76),Cin=>p(35)(76),clock=>clock,reset=>reset,s=>p(150)(76),cout=>p(151)(77));
FA_ff_1485:FAff port map(x=>p(33)(77),y=>p(34)(77),Cin=>p(35)(77),clock=>clock,reset=>reset,s=>p(150)(77),cout=>p(151)(78));
FA_ff_1486:FAff port map(x=>p(33)(78),y=>p(34)(78),Cin=>p(35)(78),clock=>clock,reset=>reset,s=>p(150)(78),cout=>p(151)(79));
FA_ff_1487:FAff port map(x=>p(33)(79),y=>p(34)(79),Cin=>p(35)(79),clock=>clock,reset=>reset,s=>p(150)(79),cout=>p(151)(80));
FA_ff_1488:FAff port map(x=>p(33)(80),y=>p(34)(80),Cin=>p(35)(80),clock=>clock,reset=>reset,s=>p(150)(80),cout=>p(151)(81));
FA_ff_1489:FAff port map(x=>p(33)(81),y=>p(34)(81),Cin=>p(35)(81),clock=>clock,reset=>reset,s=>p(150)(81),cout=>p(151)(82));
FA_ff_1490:FAff port map(x=>p(33)(82),y=>p(34)(82),Cin=>p(35)(82),clock=>clock,reset=>reset,s=>p(150)(82),cout=>p(151)(83));
FA_ff_1491:FAff port map(x=>p(33)(83),y=>p(34)(83),Cin=>p(35)(83),clock=>clock,reset=>reset,s=>p(150)(83),cout=>p(151)(84));
FA_ff_1492:FAff port map(x=>p(33)(84),y=>p(34)(84),Cin=>p(35)(84),clock=>clock,reset=>reset,s=>p(150)(84),cout=>p(151)(85));
FA_ff_1493:FAff port map(x=>p(33)(85),y=>p(34)(85),Cin=>p(35)(85),clock=>clock,reset=>reset,s=>p(150)(85),cout=>p(151)(86));
FA_ff_1494:FAff port map(x=>p(33)(86),y=>p(34)(86),Cin=>p(35)(86),clock=>clock,reset=>reset,s=>p(150)(86),cout=>p(151)(87));
FA_ff_1495:FAff port map(x=>p(33)(87),y=>p(34)(87),Cin=>p(35)(87),clock=>clock,reset=>reset,s=>p(150)(87),cout=>p(151)(88));
FA_ff_1496:FAff port map(x=>p(33)(88),y=>p(34)(88),Cin=>p(35)(88),clock=>clock,reset=>reset,s=>p(150)(88),cout=>p(151)(89));
FA_ff_1497:FAff port map(x=>p(33)(89),y=>p(34)(89),Cin=>p(35)(89),clock=>clock,reset=>reset,s=>p(150)(89),cout=>p(151)(90));
FA_ff_1498:FAff port map(x=>p(33)(90),y=>p(34)(90),Cin=>p(35)(90),clock=>clock,reset=>reset,s=>p(150)(90),cout=>p(151)(91));
FA_ff_1499:FAff port map(x=>p(33)(91),y=>p(34)(91),Cin=>p(35)(91),clock=>clock,reset=>reset,s=>p(150)(91),cout=>p(151)(92));
FA_ff_1500:FAff port map(x=>p(33)(92),y=>p(34)(92),Cin=>p(35)(92),clock=>clock,reset=>reset,s=>p(150)(92),cout=>p(151)(93));
FA_ff_1501:FAff port map(x=>p(33)(93),y=>p(34)(93),Cin=>p(35)(93),clock=>clock,reset=>reset,s=>p(150)(93),cout=>p(151)(94));
FA_ff_1502:FAff port map(x=>p(33)(94),y=>p(34)(94),Cin=>p(35)(94),clock=>clock,reset=>reset,s=>p(150)(94),cout=>p(151)(95));
FA_ff_1503:FAff port map(x=>p(33)(95),y=>p(34)(95),Cin=>p(35)(95),clock=>clock,reset=>reset,s=>p(150)(95),cout=>p(151)(96));
FA_ff_1504:FAff port map(x=>p(33)(96),y=>p(34)(96),Cin=>p(35)(96),clock=>clock,reset=>reset,s=>p(150)(96),cout=>p(151)(97));
FA_ff_1505:FAff port map(x=>p(33)(97),y=>p(34)(97),Cin=>p(35)(97),clock=>clock,reset=>reset,s=>p(150)(97),cout=>p(151)(98));
FA_ff_1506:FAff port map(x=>p(33)(98),y=>p(34)(98),Cin=>p(35)(98),clock=>clock,reset=>reset,s=>p(150)(98),cout=>p(151)(99));
FA_ff_1507:FAff port map(x=>p(33)(99),y=>p(34)(99),Cin=>p(35)(99),clock=>clock,reset=>reset,s=>p(150)(99),cout=>p(151)(100));
FA_ff_1508:FAff port map(x=>p(33)(100),y=>p(34)(100),Cin=>p(35)(100),clock=>clock,reset=>reset,s=>p(150)(100),cout=>p(151)(101));
FA_ff_1509:FAff port map(x=>p(33)(101),y=>p(34)(101),Cin=>p(35)(101),clock=>clock,reset=>reset,s=>p(150)(101),cout=>p(151)(102));
FA_ff_1510:FAff port map(x=>p(33)(102),y=>p(34)(102),Cin=>p(35)(102),clock=>clock,reset=>reset,s=>p(150)(102),cout=>p(151)(103));
FA_ff_1511:FAff port map(x=>p(33)(103),y=>p(34)(103),Cin=>p(35)(103),clock=>clock,reset=>reset,s=>p(150)(103),cout=>p(151)(104));
FA_ff_1512:FAff port map(x=>p(33)(104),y=>p(34)(104),Cin=>p(35)(104),clock=>clock,reset=>reset,s=>p(150)(104),cout=>p(151)(105));
FA_ff_1513:FAff port map(x=>p(33)(105),y=>p(34)(105),Cin=>p(35)(105),clock=>clock,reset=>reset,s=>p(150)(105),cout=>p(151)(106));
FA_ff_1514:FAff port map(x=>p(33)(106),y=>p(34)(106),Cin=>p(35)(106),clock=>clock,reset=>reset,s=>p(150)(106),cout=>p(151)(107));
FA_ff_1515:FAff port map(x=>p(33)(107),y=>p(34)(107),Cin=>p(35)(107),clock=>clock,reset=>reset,s=>p(150)(107),cout=>p(151)(108));
FA_ff_1516:FAff port map(x=>p(33)(108),y=>p(34)(108),Cin=>p(35)(108),clock=>clock,reset=>reset,s=>p(150)(108),cout=>p(151)(109));
FA_ff_1517:FAff port map(x=>p(33)(109),y=>p(34)(109),Cin=>p(35)(109),clock=>clock,reset=>reset,s=>p(150)(109),cout=>p(151)(110));
FA_ff_1518:FAff port map(x=>p(33)(110),y=>p(34)(110),Cin=>p(35)(110),clock=>clock,reset=>reset,s=>p(150)(110),cout=>p(151)(111));
FA_ff_1519:FAff port map(x=>p(33)(111),y=>p(34)(111),Cin=>p(35)(111),clock=>clock,reset=>reset,s=>p(150)(111),cout=>p(151)(112));
FA_ff_1520:FAff port map(x=>p(33)(112),y=>p(34)(112),Cin=>p(35)(112),clock=>clock,reset=>reset,s=>p(150)(112),cout=>p(151)(113));
FA_ff_1521:FAff port map(x=>p(33)(113),y=>p(34)(113),Cin=>p(35)(113),clock=>clock,reset=>reset,s=>p(150)(113),cout=>p(151)(114));
FA_ff_1522:FAff port map(x=>p(33)(114),y=>p(34)(114),Cin=>p(35)(114),clock=>clock,reset=>reset,s=>p(150)(114),cout=>p(151)(115));
FA_ff_1523:FAff port map(x=>p(33)(115),y=>p(34)(115),Cin=>p(35)(115),clock=>clock,reset=>reset,s=>p(150)(115),cout=>p(151)(116));
FA_ff_1524:FAff port map(x=>p(33)(116),y=>p(34)(116),Cin=>p(35)(116),clock=>clock,reset=>reset,s=>p(150)(116),cout=>p(151)(117));
FA_ff_1525:FAff port map(x=>p(33)(117),y=>p(34)(117),Cin=>p(35)(117),clock=>clock,reset=>reset,s=>p(150)(117),cout=>p(151)(118));
FA_ff_1526:FAff port map(x=>p(33)(118),y=>p(34)(118),Cin=>p(35)(118),clock=>clock,reset=>reset,s=>p(150)(118),cout=>p(151)(119));
FA_ff_1527:FAff port map(x=>p(33)(119),y=>p(34)(119),Cin=>p(35)(119),clock=>clock,reset=>reset,s=>p(150)(119),cout=>p(151)(120));
FA_ff_1528:FAff port map(x=>p(33)(120),y=>p(34)(120),Cin=>p(35)(120),clock=>clock,reset=>reset,s=>p(150)(120),cout=>p(151)(121));
FA_ff_1529:FAff port map(x=>p(33)(121),y=>p(34)(121),Cin=>p(35)(121),clock=>clock,reset=>reset,s=>p(150)(121),cout=>p(151)(122));
FA_ff_1530:FAff port map(x=>p(33)(122),y=>p(34)(122),Cin=>p(35)(122),clock=>clock,reset=>reset,s=>p(150)(122),cout=>p(151)(123));
FA_ff_1531:FAff port map(x=>p(33)(123),y=>p(34)(123),Cin=>p(35)(123),clock=>clock,reset=>reset,s=>p(150)(123),cout=>p(151)(124));
FA_ff_1532:FAff port map(x=>p(33)(124),y=>p(34)(124),Cin=>p(35)(124),clock=>clock,reset=>reset,s=>p(150)(124),cout=>p(151)(125));
FA_ff_1533:FAff port map(x=>p(33)(125),y=>p(34)(125),Cin=>p(35)(125),clock=>clock,reset=>reset,s=>p(150)(125),cout=>p(151)(126));
FA_ff_1534:FAff port map(x=>p(33)(126),y=>p(34)(126),Cin=>p(35)(126),clock=>clock,reset=>reset,s=>p(150)(126),cout=>p(151)(127));
FA_ff_1535:FAff port map(x=>p(33)(127),y=>p(34)(127),Cin=>p(35)(127),clock=>clock,reset=>reset,s=>p(150)(127),cout=>p(151)(128));
FA_ff_1536:FAff port map(x=>p(36)(0),y=>p(37)(0),Cin=>p(38)(0),clock=>clock,reset=>reset,s=>p(152)(0),cout=>p(153)(1));
FA_ff_1537:FAff port map(x=>p(36)(1),y=>p(37)(1),Cin=>p(38)(1),clock=>clock,reset=>reset,s=>p(152)(1),cout=>p(153)(2));
FA_ff_1538:FAff port map(x=>p(36)(2),y=>p(37)(2),Cin=>p(38)(2),clock=>clock,reset=>reset,s=>p(152)(2),cout=>p(153)(3));
FA_ff_1539:FAff port map(x=>p(36)(3),y=>p(37)(3),Cin=>p(38)(3),clock=>clock,reset=>reset,s=>p(152)(3),cout=>p(153)(4));
FA_ff_1540:FAff port map(x=>p(36)(4),y=>p(37)(4),Cin=>p(38)(4),clock=>clock,reset=>reset,s=>p(152)(4),cout=>p(153)(5));
FA_ff_1541:FAff port map(x=>p(36)(5),y=>p(37)(5),Cin=>p(38)(5),clock=>clock,reset=>reset,s=>p(152)(5),cout=>p(153)(6));
FA_ff_1542:FAff port map(x=>p(36)(6),y=>p(37)(6),Cin=>p(38)(6),clock=>clock,reset=>reset,s=>p(152)(6),cout=>p(153)(7));
FA_ff_1543:FAff port map(x=>p(36)(7),y=>p(37)(7),Cin=>p(38)(7),clock=>clock,reset=>reset,s=>p(152)(7),cout=>p(153)(8));
FA_ff_1544:FAff port map(x=>p(36)(8),y=>p(37)(8),Cin=>p(38)(8),clock=>clock,reset=>reset,s=>p(152)(8),cout=>p(153)(9));
FA_ff_1545:FAff port map(x=>p(36)(9),y=>p(37)(9),Cin=>p(38)(9),clock=>clock,reset=>reset,s=>p(152)(9),cout=>p(153)(10));
FA_ff_1546:FAff port map(x=>p(36)(10),y=>p(37)(10),Cin=>p(38)(10),clock=>clock,reset=>reset,s=>p(152)(10),cout=>p(153)(11));
FA_ff_1547:FAff port map(x=>p(36)(11),y=>p(37)(11),Cin=>p(38)(11),clock=>clock,reset=>reset,s=>p(152)(11),cout=>p(153)(12));
FA_ff_1548:FAff port map(x=>p(36)(12),y=>p(37)(12),Cin=>p(38)(12),clock=>clock,reset=>reset,s=>p(152)(12),cout=>p(153)(13));
FA_ff_1549:FAff port map(x=>p(36)(13),y=>p(37)(13),Cin=>p(38)(13),clock=>clock,reset=>reset,s=>p(152)(13),cout=>p(153)(14));
FA_ff_1550:FAff port map(x=>p(36)(14),y=>p(37)(14),Cin=>p(38)(14),clock=>clock,reset=>reset,s=>p(152)(14),cout=>p(153)(15));
FA_ff_1551:FAff port map(x=>p(36)(15),y=>p(37)(15),Cin=>p(38)(15),clock=>clock,reset=>reset,s=>p(152)(15),cout=>p(153)(16));
FA_ff_1552:FAff port map(x=>p(36)(16),y=>p(37)(16),Cin=>p(38)(16),clock=>clock,reset=>reset,s=>p(152)(16),cout=>p(153)(17));
FA_ff_1553:FAff port map(x=>p(36)(17),y=>p(37)(17),Cin=>p(38)(17),clock=>clock,reset=>reset,s=>p(152)(17),cout=>p(153)(18));
FA_ff_1554:FAff port map(x=>p(36)(18),y=>p(37)(18),Cin=>p(38)(18),clock=>clock,reset=>reset,s=>p(152)(18),cout=>p(153)(19));
FA_ff_1555:FAff port map(x=>p(36)(19),y=>p(37)(19),Cin=>p(38)(19),clock=>clock,reset=>reset,s=>p(152)(19),cout=>p(153)(20));
FA_ff_1556:FAff port map(x=>p(36)(20),y=>p(37)(20),Cin=>p(38)(20),clock=>clock,reset=>reset,s=>p(152)(20),cout=>p(153)(21));
FA_ff_1557:FAff port map(x=>p(36)(21),y=>p(37)(21),Cin=>p(38)(21),clock=>clock,reset=>reset,s=>p(152)(21),cout=>p(153)(22));
FA_ff_1558:FAff port map(x=>p(36)(22),y=>p(37)(22),Cin=>p(38)(22),clock=>clock,reset=>reset,s=>p(152)(22),cout=>p(153)(23));
FA_ff_1559:FAff port map(x=>p(36)(23),y=>p(37)(23),Cin=>p(38)(23),clock=>clock,reset=>reset,s=>p(152)(23),cout=>p(153)(24));
FA_ff_1560:FAff port map(x=>p(36)(24),y=>p(37)(24),Cin=>p(38)(24),clock=>clock,reset=>reset,s=>p(152)(24),cout=>p(153)(25));
FA_ff_1561:FAff port map(x=>p(36)(25),y=>p(37)(25),Cin=>p(38)(25),clock=>clock,reset=>reset,s=>p(152)(25),cout=>p(153)(26));
FA_ff_1562:FAff port map(x=>p(36)(26),y=>p(37)(26),Cin=>p(38)(26),clock=>clock,reset=>reset,s=>p(152)(26),cout=>p(153)(27));
FA_ff_1563:FAff port map(x=>p(36)(27),y=>p(37)(27),Cin=>p(38)(27),clock=>clock,reset=>reset,s=>p(152)(27),cout=>p(153)(28));
FA_ff_1564:FAff port map(x=>p(36)(28),y=>p(37)(28),Cin=>p(38)(28),clock=>clock,reset=>reset,s=>p(152)(28),cout=>p(153)(29));
FA_ff_1565:FAff port map(x=>p(36)(29),y=>p(37)(29),Cin=>p(38)(29),clock=>clock,reset=>reset,s=>p(152)(29),cout=>p(153)(30));
FA_ff_1566:FAff port map(x=>p(36)(30),y=>p(37)(30),Cin=>p(38)(30),clock=>clock,reset=>reset,s=>p(152)(30),cout=>p(153)(31));
FA_ff_1567:FAff port map(x=>p(36)(31),y=>p(37)(31),Cin=>p(38)(31),clock=>clock,reset=>reset,s=>p(152)(31),cout=>p(153)(32));
FA_ff_1568:FAff port map(x=>p(36)(32),y=>p(37)(32),Cin=>p(38)(32),clock=>clock,reset=>reset,s=>p(152)(32),cout=>p(153)(33));
FA_ff_1569:FAff port map(x=>p(36)(33),y=>p(37)(33),Cin=>p(38)(33),clock=>clock,reset=>reset,s=>p(152)(33),cout=>p(153)(34));
FA_ff_1570:FAff port map(x=>p(36)(34),y=>p(37)(34),Cin=>p(38)(34),clock=>clock,reset=>reset,s=>p(152)(34),cout=>p(153)(35));
FA_ff_1571:FAff port map(x=>p(36)(35),y=>p(37)(35),Cin=>p(38)(35),clock=>clock,reset=>reset,s=>p(152)(35),cout=>p(153)(36));
FA_ff_1572:FAff port map(x=>p(36)(36),y=>p(37)(36),Cin=>p(38)(36),clock=>clock,reset=>reset,s=>p(152)(36),cout=>p(153)(37));
FA_ff_1573:FAff port map(x=>p(36)(37),y=>p(37)(37),Cin=>p(38)(37),clock=>clock,reset=>reset,s=>p(152)(37),cout=>p(153)(38));
FA_ff_1574:FAff port map(x=>p(36)(38),y=>p(37)(38),Cin=>p(38)(38),clock=>clock,reset=>reset,s=>p(152)(38),cout=>p(153)(39));
FA_ff_1575:FAff port map(x=>p(36)(39),y=>p(37)(39),Cin=>p(38)(39),clock=>clock,reset=>reset,s=>p(152)(39),cout=>p(153)(40));
FA_ff_1576:FAff port map(x=>p(36)(40),y=>p(37)(40),Cin=>p(38)(40),clock=>clock,reset=>reset,s=>p(152)(40),cout=>p(153)(41));
FA_ff_1577:FAff port map(x=>p(36)(41),y=>p(37)(41),Cin=>p(38)(41),clock=>clock,reset=>reset,s=>p(152)(41),cout=>p(153)(42));
FA_ff_1578:FAff port map(x=>p(36)(42),y=>p(37)(42),Cin=>p(38)(42),clock=>clock,reset=>reset,s=>p(152)(42),cout=>p(153)(43));
FA_ff_1579:FAff port map(x=>p(36)(43),y=>p(37)(43),Cin=>p(38)(43),clock=>clock,reset=>reset,s=>p(152)(43),cout=>p(153)(44));
FA_ff_1580:FAff port map(x=>p(36)(44),y=>p(37)(44),Cin=>p(38)(44),clock=>clock,reset=>reset,s=>p(152)(44),cout=>p(153)(45));
FA_ff_1581:FAff port map(x=>p(36)(45),y=>p(37)(45),Cin=>p(38)(45),clock=>clock,reset=>reset,s=>p(152)(45),cout=>p(153)(46));
FA_ff_1582:FAff port map(x=>p(36)(46),y=>p(37)(46),Cin=>p(38)(46),clock=>clock,reset=>reset,s=>p(152)(46),cout=>p(153)(47));
FA_ff_1583:FAff port map(x=>p(36)(47),y=>p(37)(47),Cin=>p(38)(47),clock=>clock,reset=>reset,s=>p(152)(47),cout=>p(153)(48));
FA_ff_1584:FAff port map(x=>p(36)(48),y=>p(37)(48),Cin=>p(38)(48),clock=>clock,reset=>reset,s=>p(152)(48),cout=>p(153)(49));
FA_ff_1585:FAff port map(x=>p(36)(49),y=>p(37)(49),Cin=>p(38)(49),clock=>clock,reset=>reset,s=>p(152)(49),cout=>p(153)(50));
FA_ff_1586:FAff port map(x=>p(36)(50),y=>p(37)(50),Cin=>p(38)(50),clock=>clock,reset=>reset,s=>p(152)(50),cout=>p(153)(51));
FA_ff_1587:FAff port map(x=>p(36)(51),y=>p(37)(51),Cin=>p(38)(51),clock=>clock,reset=>reset,s=>p(152)(51),cout=>p(153)(52));
FA_ff_1588:FAff port map(x=>p(36)(52),y=>p(37)(52),Cin=>p(38)(52),clock=>clock,reset=>reset,s=>p(152)(52),cout=>p(153)(53));
FA_ff_1589:FAff port map(x=>p(36)(53),y=>p(37)(53),Cin=>p(38)(53),clock=>clock,reset=>reset,s=>p(152)(53),cout=>p(153)(54));
FA_ff_1590:FAff port map(x=>p(36)(54),y=>p(37)(54),Cin=>p(38)(54),clock=>clock,reset=>reset,s=>p(152)(54),cout=>p(153)(55));
FA_ff_1591:FAff port map(x=>p(36)(55),y=>p(37)(55),Cin=>p(38)(55),clock=>clock,reset=>reset,s=>p(152)(55),cout=>p(153)(56));
FA_ff_1592:FAff port map(x=>p(36)(56),y=>p(37)(56),Cin=>p(38)(56),clock=>clock,reset=>reset,s=>p(152)(56),cout=>p(153)(57));
FA_ff_1593:FAff port map(x=>p(36)(57),y=>p(37)(57),Cin=>p(38)(57),clock=>clock,reset=>reset,s=>p(152)(57),cout=>p(153)(58));
FA_ff_1594:FAff port map(x=>p(36)(58),y=>p(37)(58),Cin=>p(38)(58),clock=>clock,reset=>reset,s=>p(152)(58),cout=>p(153)(59));
FA_ff_1595:FAff port map(x=>p(36)(59),y=>p(37)(59),Cin=>p(38)(59),clock=>clock,reset=>reset,s=>p(152)(59),cout=>p(153)(60));
FA_ff_1596:FAff port map(x=>p(36)(60),y=>p(37)(60),Cin=>p(38)(60),clock=>clock,reset=>reset,s=>p(152)(60),cout=>p(153)(61));
FA_ff_1597:FAff port map(x=>p(36)(61),y=>p(37)(61),Cin=>p(38)(61),clock=>clock,reset=>reset,s=>p(152)(61),cout=>p(153)(62));
FA_ff_1598:FAff port map(x=>p(36)(62),y=>p(37)(62),Cin=>p(38)(62),clock=>clock,reset=>reset,s=>p(152)(62),cout=>p(153)(63));
FA_ff_1599:FAff port map(x=>p(36)(63),y=>p(37)(63),Cin=>p(38)(63),clock=>clock,reset=>reset,s=>p(152)(63),cout=>p(153)(64));
FA_ff_1600:FAff port map(x=>p(36)(64),y=>p(37)(64),Cin=>p(38)(64),clock=>clock,reset=>reset,s=>p(152)(64),cout=>p(153)(65));
FA_ff_1601:FAff port map(x=>p(36)(65),y=>p(37)(65),Cin=>p(38)(65),clock=>clock,reset=>reset,s=>p(152)(65),cout=>p(153)(66));
FA_ff_1602:FAff port map(x=>p(36)(66),y=>p(37)(66),Cin=>p(38)(66),clock=>clock,reset=>reset,s=>p(152)(66),cout=>p(153)(67));
FA_ff_1603:FAff port map(x=>p(36)(67),y=>p(37)(67),Cin=>p(38)(67),clock=>clock,reset=>reset,s=>p(152)(67),cout=>p(153)(68));
FA_ff_1604:FAff port map(x=>p(36)(68),y=>p(37)(68),Cin=>p(38)(68),clock=>clock,reset=>reset,s=>p(152)(68),cout=>p(153)(69));
FA_ff_1605:FAff port map(x=>p(36)(69),y=>p(37)(69),Cin=>p(38)(69),clock=>clock,reset=>reset,s=>p(152)(69),cout=>p(153)(70));
FA_ff_1606:FAff port map(x=>p(36)(70),y=>p(37)(70),Cin=>p(38)(70),clock=>clock,reset=>reset,s=>p(152)(70),cout=>p(153)(71));
FA_ff_1607:FAff port map(x=>p(36)(71),y=>p(37)(71),Cin=>p(38)(71),clock=>clock,reset=>reset,s=>p(152)(71),cout=>p(153)(72));
FA_ff_1608:FAff port map(x=>p(36)(72),y=>p(37)(72),Cin=>p(38)(72),clock=>clock,reset=>reset,s=>p(152)(72),cout=>p(153)(73));
FA_ff_1609:FAff port map(x=>p(36)(73),y=>p(37)(73),Cin=>p(38)(73),clock=>clock,reset=>reset,s=>p(152)(73),cout=>p(153)(74));
FA_ff_1610:FAff port map(x=>p(36)(74),y=>p(37)(74),Cin=>p(38)(74),clock=>clock,reset=>reset,s=>p(152)(74),cout=>p(153)(75));
FA_ff_1611:FAff port map(x=>p(36)(75),y=>p(37)(75),Cin=>p(38)(75),clock=>clock,reset=>reset,s=>p(152)(75),cout=>p(153)(76));
FA_ff_1612:FAff port map(x=>p(36)(76),y=>p(37)(76),Cin=>p(38)(76),clock=>clock,reset=>reset,s=>p(152)(76),cout=>p(153)(77));
FA_ff_1613:FAff port map(x=>p(36)(77),y=>p(37)(77),Cin=>p(38)(77),clock=>clock,reset=>reset,s=>p(152)(77),cout=>p(153)(78));
FA_ff_1614:FAff port map(x=>p(36)(78),y=>p(37)(78),Cin=>p(38)(78),clock=>clock,reset=>reset,s=>p(152)(78),cout=>p(153)(79));
FA_ff_1615:FAff port map(x=>p(36)(79),y=>p(37)(79),Cin=>p(38)(79),clock=>clock,reset=>reset,s=>p(152)(79),cout=>p(153)(80));
FA_ff_1616:FAff port map(x=>p(36)(80),y=>p(37)(80),Cin=>p(38)(80),clock=>clock,reset=>reset,s=>p(152)(80),cout=>p(153)(81));
FA_ff_1617:FAff port map(x=>p(36)(81),y=>p(37)(81),Cin=>p(38)(81),clock=>clock,reset=>reset,s=>p(152)(81),cout=>p(153)(82));
FA_ff_1618:FAff port map(x=>p(36)(82),y=>p(37)(82),Cin=>p(38)(82),clock=>clock,reset=>reset,s=>p(152)(82),cout=>p(153)(83));
FA_ff_1619:FAff port map(x=>p(36)(83),y=>p(37)(83),Cin=>p(38)(83),clock=>clock,reset=>reset,s=>p(152)(83),cout=>p(153)(84));
FA_ff_1620:FAff port map(x=>p(36)(84),y=>p(37)(84),Cin=>p(38)(84),clock=>clock,reset=>reset,s=>p(152)(84),cout=>p(153)(85));
FA_ff_1621:FAff port map(x=>p(36)(85),y=>p(37)(85),Cin=>p(38)(85),clock=>clock,reset=>reset,s=>p(152)(85),cout=>p(153)(86));
FA_ff_1622:FAff port map(x=>p(36)(86),y=>p(37)(86),Cin=>p(38)(86),clock=>clock,reset=>reset,s=>p(152)(86),cout=>p(153)(87));
FA_ff_1623:FAff port map(x=>p(36)(87),y=>p(37)(87),Cin=>p(38)(87),clock=>clock,reset=>reset,s=>p(152)(87),cout=>p(153)(88));
FA_ff_1624:FAff port map(x=>p(36)(88),y=>p(37)(88),Cin=>p(38)(88),clock=>clock,reset=>reset,s=>p(152)(88),cout=>p(153)(89));
FA_ff_1625:FAff port map(x=>p(36)(89),y=>p(37)(89),Cin=>p(38)(89),clock=>clock,reset=>reset,s=>p(152)(89),cout=>p(153)(90));
FA_ff_1626:FAff port map(x=>p(36)(90),y=>p(37)(90),Cin=>p(38)(90),clock=>clock,reset=>reset,s=>p(152)(90),cout=>p(153)(91));
FA_ff_1627:FAff port map(x=>p(36)(91),y=>p(37)(91),Cin=>p(38)(91),clock=>clock,reset=>reset,s=>p(152)(91),cout=>p(153)(92));
FA_ff_1628:FAff port map(x=>p(36)(92),y=>p(37)(92),Cin=>p(38)(92),clock=>clock,reset=>reset,s=>p(152)(92),cout=>p(153)(93));
FA_ff_1629:FAff port map(x=>p(36)(93),y=>p(37)(93),Cin=>p(38)(93),clock=>clock,reset=>reset,s=>p(152)(93),cout=>p(153)(94));
FA_ff_1630:FAff port map(x=>p(36)(94),y=>p(37)(94),Cin=>p(38)(94),clock=>clock,reset=>reset,s=>p(152)(94),cout=>p(153)(95));
FA_ff_1631:FAff port map(x=>p(36)(95),y=>p(37)(95),Cin=>p(38)(95),clock=>clock,reset=>reset,s=>p(152)(95),cout=>p(153)(96));
FA_ff_1632:FAff port map(x=>p(36)(96),y=>p(37)(96),Cin=>p(38)(96),clock=>clock,reset=>reset,s=>p(152)(96),cout=>p(153)(97));
FA_ff_1633:FAff port map(x=>p(36)(97),y=>p(37)(97),Cin=>p(38)(97),clock=>clock,reset=>reset,s=>p(152)(97),cout=>p(153)(98));
FA_ff_1634:FAff port map(x=>p(36)(98),y=>p(37)(98),Cin=>p(38)(98),clock=>clock,reset=>reset,s=>p(152)(98),cout=>p(153)(99));
FA_ff_1635:FAff port map(x=>p(36)(99),y=>p(37)(99),Cin=>p(38)(99),clock=>clock,reset=>reset,s=>p(152)(99),cout=>p(153)(100));
FA_ff_1636:FAff port map(x=>p(36)(100),y=>p(37)(100),Cin=>p(38)(100),clock=>clock,reset=>reset,s=>p(152)(100),cout=>p(153)(101));
FA_ff_1637:FAff port map(x=>p(36)(101),y=>p(37)(101),Cin=>p(38)(101),clock=>clock,reset=>reset,s=>p(152)(101),cout=>p(153)(102));
FA_ff_1638:FAff port map(x=>p(36)(102),y=>p(37)(102),Cin=>p(38)(102),clock=>clock,reset=>reset,s=>p(152)(102),cout=>p(153)(103));
FA_ff_1639:FAff port map(x=>p(36)(103),y=>p(37)(103),Cin=>p(38)(103),clock=>clock,reset=>reset,s=>p(152)(103),cout=>p(153)(104));
FA_ff_1640:FAff port map(x=>p(36)(104),y=>p(37)(104),Cin=>p(38)(104),clock=>clock,reset=>reset,s=>p(152)(104),cout=>p(153)(105));
FA_ff_1641:FAff port map(x=>p(36)(105),y=>p(37)(105),Cin=>p(38)(105),clock=>clock,reset=>reset,s=>p(152)(105),cout=>p(153)(106));
FA_ff_1642:FAff port map(x=>p(36)(106),y=>p(37)(106),Cin=>p(38)(106),clock=>clock,reset=>reset,s=>p(152)(106),cout=>p(153)(107));
FA_ff_1643:FAff port map(x=>p(36)(107),y=>p(37)(107),Cin=>p(38)(107),clock=>clock,reset=>reset,s=>p(152)(107),cout=>p(153)(108));
FA_ff_1644:FAff port map(x=>p(36)(108),y=>p(37)(108),Cin=>p(38)(108),clock=>clock,reset=>reset,s=>p(152)(108),cout=>p(153)(109));
FA_ff_1645:FAff port map(x=>p(36)(109),y=>p(37)(109),Cin=>p(38)(109),clock=>clock,reset=>reset,s=>p(152)(109),cout=>p(153)(110));
FA_ff_1646:FAff port map(x=>p(36)(110),y=>p(37)(110),Cin=>p(38)(110),clock=>clock,reset=>reset,s=>p(152)(110),cout=>p(153)(111));
FA_ff_1647:FAff port map(x=>p(36)(111),y=>p(37)(111),Cin=>p(38)(111),clock=>clock,reset=>reset,s=>p(152)(111),cout=>p(153)(112));
FA_ff_1648:FAff port map(x=>p(36)(112),y=>p(37)(112),Cin=>p(38)(112),clock=>clock,reset=>reset,s=>p(152)(112),cout=>p(153)(113));
FA_ff_1649:FAff port map(x=>p(36)(113),y=>p(37)(113),Cin=>p(38)(113),clock=>clock,reset=>reset,s=>p(152)(113),cout=>p(153)(114));
FA_ff_1650:FAff port map(x=>p(36)(114),y=>p(37)(114),Cin=>p(38)(114),clock=>clock,reset=>reset,s=>p(152)(114),cout=>p(153)(115));
FA_ff_1651:FAff port map(x=>p(36)(115),y=>p(37)(115),Cin=>p(38)(115),clock=>clock,reset=>reset,s=>p(152)(115),cout=>p(153)(116));
FA_ff_1652:FAff port map(x=>p(36)(116),y=>p(37)(116),Cin=>p(38)(116),clock=>clock,reset=>reset,s=>p(152)(116),cout=>p(153)(117));
FA_ff_1653:FAff port map(x=>p(36)(117),y=>p(37)(117),Cin=>p(38)(117),clock=>clock,reset=>reset,s=>p(152)(117),cout=>p(153)(118));
FA_ff_1654:FAff port map(x=>p(36)(118),y=>p(37)(118),Cin=>p(38)(118),clock=>clock,reset=>reset,s=>p(152)(118),cout=>p(153)(119));
FA_ff_1655:FAff port map(x=>p(36)(119),y=>p(37)(119),Cin=>p(38)(119),clock=>clock,reset=>reset,s=>p(152)(119),cout=>p(153)(120));
FA_ff_1656:FAff port map(x=>p(36)(120),y=>p(37)(120),Cin=>p(38)(120),clock=>clock,reset=>reset,s=>p(152)(120),cout=>p(153)(121));
FA_ff_1657:FAff port map(x=>p(36)(121),y=>p(37)(121),Cin=>p(38)(121),clock=>clock,reset=>reset,s=>p(152)(121),cout=>p(153)(122));
FA_ff_1658:FAff port map(x=>p(36)(122),y=>p(37)(122),Cin=>p(38)(122),clock=>clock,reset=>reset,s=>p(152)(122),cout=>p(153)(123));
FA_ff_1659:FAff port map(x=>p(36)(123),y=>p(37)(123),Cin=>p(38)(123),clock=>clock,reset=>reset,s=>p(152)(123),cout=>p(153)(124));
FA_ff_1660:FAff port map(x=>p(36)(124),y=>p(37)(124),Cin=>p(38)(124),clock=>clock,reset=>reset,s=>p(152)(124),cout=>p(153)(125));
FA_ff_1661:FAff port map(x=>p(36)(125),y=>p(37)(125),Cin=>p(38)(125),clock=>clock,reset=>reset,s=>p(152)(125),cout=>p(153)(126));
FA_ff_1662:FAff port map(x=>p(36)(126),y=>p(37)(126),Cin=>p(38)(126),clock=>clock,reset=>reset,s=>p(152)(126),cout=>p(153)(127));
FA_ff_1663:FAff port map(x=>p(36)(127),y=>p(37)(127),Cin=>p(38)(127),clock=>clock,reset=>reset,s=>p(152)(127),cout=>p(153)(128));
FA_ff_1664:FAff port map(x=>p(39)(0),y=>p(40)(0),Cin=>p(41)(0),clock=>clock,reset=>reset,s=>p(154)(0),cout=>p(155)(1));
FA_ff_1665:FAff port map(x=>p(39)(1),y=>p(40)(1),Cin=>p(41)(1),clock=>clock,reset=>reset,s=>p(154)(1),cout=>p(155)(2));
FA_ff_1666:FAff port map(x=>p(39)(2),y=>p(40)(2),Cin=>p(41)(2),clock=>clock,reset=>reset,s=>p(154)(2),cout=>p(155)(3));
FA_ff_1667:FAff port map(x=>p(39)(3),y=>p(40)(3),Cin=>p(41)(3),clock=>clock,reset=>reset,s=>p(154)(3),cout=>p(155)(4));
FA_ff_1668:FAff port map(x=>p(39)(4),y=>p(40)(4),Cin=>p(41)(4),clock=>clock,reset=>reset,s=>p(154)(4),cout=>p(155)(5));
FA_ff_1669:FAff port map(x=>p(39)(5),y=>p(40)(5),Cin=>p(41)(5),clock=>clock,reset=>reset,s=>p(154)(5),cout=>p(155)(6));
FA_ff_1670:FAff port map(x=>p(39)(6),y=>p(40)(6),Cin=>p(41)(6),clock=>clock,reset=>reset,s=>p(154)(6),cout=>p(155)(7));
FA_ff_1671:FAff port map(x=>p(39)(7),y=>p(40)(7),Cin=>p(41)(7),clock=>clock,reset=>reset,s=>p(154)(7),cout=>p(155)(8));
FA_ff_1672:FAff port map(x=>p(39)(8),y=>p(40)(8),Cin=>p(41)(8),clock=>clock,reset=>reset,s=>p(154)(8),cout=>p(155)(9));
FA_ff_1673:FAff port map(x=>p(39)(9),y=>p(40)(9),Cin=>p(41)(9),clock=>clock,reset=>reset,s=>p(154)(9),cout=>p(155)(10));
FA_ff_1674:FAff port map(x=>p(39)(10),y=>p(40)(10),Cin=>p(41)(10),clock=>clock,reset=>reset,s=>p(154)(10),cout=>p(155)(11));
FA_ff_1675:FAff port map(x=>p(39)(11),y=>p(40)(11),Cin=>p(41)(11),clock=>clock,reset=>reset,s=>p(154)(11),cout=>p(155)(12));
FA_ff_1676:FAff port map(x=>p(39)(12),y=>p(40)(12),Cin=>p(41)(12),clock=>clock,reset=>reset,s=>p(154)(12),cout=>p(155)(13));
FA_ff_1677:FAff port map(x=>p(39)(13),y=>p(40)(13),Cin=>p(41)(13),clock=>clock,reset=>reset,s=>p(154)(13),cout=>p(155)(14));
FA_ff_1678:FAff port map(x=>p(39)(14),y=>p(40)(14),Cin=>p(41)(14),clock=>clock,reset=>reset,s=>p(154)(14),cout=>p(155)(15));
FA_ff_1679:FAff port map(x=>p(39)(15),y=>p(40)(15),Cin=>p(41)(15),clock=>clock,reset=>reset,s=>p(154)(15),cout=>p(155)(16));
FA_ff_1680:FAff port map(x=>p(39)(16),y=>p(40)(16),Cin=>p(41)(16),clock=>clock,reset=>reset,s=>p(154)(16),cout=>p(155)(17));
FA_ff_1681:FAff port map(x=>p(39)(17),y=>p(40)(17),Cin=>p(41)(17),clock=>clock,reset=>reset,s=>p(154)(17),cout=>p(155)(18));
FA_ff_1682:FAff port map(x=>p(39)(18),y=>p(40)(18),Cin=>p(41)(18),clock=>clock,reset=>reset,s=>p(154)(18),cout=>p(155)(19));
FA_ff_1683:FAff port map(x=>p(39)(19),y=>p(40)(19),Cin=>p(41)(19),clock=>clock,reset=>reset,s=>p(154)(19),cout=>p(155)(20));
FA_ff_1684:FAff port map(x=>p(39)(20),y=>p(40)(20),Cin=>p(41)(20),clock=>clock,reset=>reset,s=>p(154)(20),cout=>p(155)(21));
FA_ff_1685:FAff port map(x=>p(39)(21),y=>p(40)(21),Cin=>p(41)(21),clock=>clock,reset=>reset,s=>p(154)(21),cout=>p(155)(22));
FA_ff_1686:FAff port map(x=>p(39)(22),y=>p(40)(22),Cin=>p(41)(22),clock=>clock,reset=>reset,s=>p(154)(22),cout=>p(155)(23));
FA_ff_1687:FAff port map(x=>p(39)(23),y=>p(40)(23),Cin=>p(41)(23),clock=>clock,reset=>reset,s=>p(154)(23),cout=>p(155)(24));
FA_ff_1688:FAff port map(x=>p(39)(24),y=>p(40)(24),Cin=>p(41)(24),clock=>clock,reset=>reset,s=>p(154)(24),cout=>p(155)(25));
FA_ff_1689:FAff port map(x=>p(39)(25),y=>p(40)(25),Cin=>p(41)(25),clock=>clock,reset=>reset,s=>p(154)(25),cout=>p(155)(26));
FA_ff_1690:FAff port map(x=>p(39)(26),y=>p(40)(26),Cin=>p(41)(26),clock=>clock,reset=>reset,s=>p(154)(26),cout=>p(155)(27));
FA_ff_1691:FAff port map(x=>p(39)(27),y=>p(40)(27),Cin=>p(41)(27),clock=>clock,reset=>reset,s=>p(154)(27),cout=>p(155)(28));
FA_ff_1692:FAff port map(x=>p(39)(28),y=>p(40)(28),Cin=>p(41)(28),clock=>clock,reset=>reset,s=>p(154)(28),cout=>p(155)(29));
FA_ff_1693:FAff port map(x=>p(39)(29),y=>p(40)(29),Cin=>p(41)(29),clock=>clock,reset=>reset,s=>p(154)(29),cout=>p(155)(30));
FA_ff_1694:FAff port map(x=>p(39)(30),y=>p(40)(30),Cin=>p(41)(30),clock=>clock,reset=>reset,s=>p(154)(30),cout=>p(155)(31));
FA_ff_1695:FAff port map(x=>p(39)(31),y=>p(40)(31),Cin=>p(41)(31),clock=>clock,reset=>reset,s=>p(154)(31),cout=>p(155)(32));
FA_ff_1696:FAff port map(x=>p(39)(32),y=>p(40)(32),Cin=>p(41)(32),clock=>clock,reset=>reset,s=>p(154)(32),cout=>p(155)(33));
FA_ff_1697:FAff port map(x=>p(39)(33),y=>p(40)(33),Cin=>p(41)(33),clock=>clock,reset=>reset,s=>p(154)(33),cout=>p(155)(34));
FA_ff_1698:FAff port map(x=>p(39)(34),y=>p(40)(34),Cin=>p(41)(34),clock=>clock,reset=>reset,s=>p(154)(34),cout=>p(155)(35));
FA_ff_1699:FAff port map(x=>p(39)(35),y=>p(40)(35),Cin=>p(41)(35),clock=>clock,reset=>reset,s=>p(154)(35),cout=>p(155)(36));
FA_ff_1700:FAff port map(x=>p(39)(36),y=>p(40)(36),Cin=>p(41)(36),clock=>clock,reset=>reset,s=>p(154)(36),cout=>p(155)(37));
FA_ff_1701:FAff port map(x=>p(39)(37),y=>p(40)(37),Cin=>p(41)(37),clock=>clock,reset=>reset,s=>p(154)(37),cout=>p(155)(38));
FA_ff_1702:FAff port map(x=>p(39)(38),y=>p(40)(38),Cin=>p(41)(38),clock=>clock,reset=>reset,s=>p(154)(38),cout=>p(155)(39));
FA_ff_1703:FAff port map(x=>p(39)(39),y=>p(40)(39),Cin=>p(41)(39),clock=>clock,reset=>reset,s=>p(154)(39),cout=>p(155)(40));
FA_ff_1704:FAff port map(x=>p(39)(40),y=>p(40)(40),Cin=>p(41)(40),clock=>clock,reset=>reset,s=>p(154)(40),cout=>p(155)(41));
FA_ff_1705:FAff port map(x=>p(39)(41),y=>p(40)(41),Cin=>p(41)(41),clock=>clock,reset=>reset,s=>p(154)(41),cout=>p(155)(42));
FA_ff_1706:FAff port map(x=>p(39)(42),y=>p(40)(42),Cin=>p(41)(42),clock=>clock,reset=>reset,s=>p(154)(42),cout=>p(155)(43));
FA_ff_1707:FAff port map(x=>p(39)(43),y=>p(40)(43),Cin=>p(41)(43),clock=>clock,reset=>reset,s=>p(154)(43),cout=>p(155)(44));
FA_ff_1708:FAff port map(x=>p(39)(44),y=>p(40)(44),Cin=>p(41)(44),clock=>clock,reset=>reset,s=>p(154)(44),cout=>p(155)(45));
FA_ff_1709:FAff port map(x=>p(39)(45),y=>p(40)(45),Cin=>p(41)(45),clock=>clock,reset=>reset,s=>p(154)(45),cout=>p(155)(46));
FA_ff_1710:FAff port map(x=>p(39)(46),y=>p(40)(46),Cin=>p(41)(46),clock=>clock,reset=>reset,s=>p(154)(46),cout=>p(155)(47));
FA_ff_1711:FAff port map(x=>p(39)(47),y=>p(40)(47),Cin=>p(41)(47),clock=>clock,reset=>reset,s=>p(154)(47),cout=>p(155)(48));
FA_ff_1712:FAff port map(x=>p(39)(48),y=>p(40)(48),Cin=>p(41)(48),clock=>clock,reset=>reset,s=>p(154)(48),cout=>p(155)(49));
FA_ff_1713:FAff port map(x=>p(39)(49),y=>p(40)(49),Cin=>p(41)(49),clock=>clock,reset=>reset,s=>p(154)(49),cout=>p(155)(50));
FA_ff_1714:FAff port map(x=>p(39)(50),y=>p(40)(50),Cin=>p(41)(50),clock=>clock,reset=>reset,s=>p(154)(50),cout=>p(155)(51));
FA_ff_1715:FAff port map(x=>p(39)(51),y=>p(40)(51),Cin=>p(41)(51),clock=>clock,reset=>reset,s=>p(154)(51),cout=>p(155)(52));
FA_ff_1716:FAff port map(x=>p(39)(52),y=>p(40)(52),Cin=>p(41)(52),clock=>clock,reset=>reset,s=>p(154)(52),cout=>p(155)(53));
FA_ff_1717:FAff port map(x=>p(39)(53),y=>p(40)(53),Cin=>p(41)(53),clock=>clock,reset=>reset,s=>p(154)(53),cout=>p(155)(54));
FA_ff_1718:FAff port map(x=>p(39)(54),y=>p(40)(54),Cin=>p(41)(54),clock=>clock,reset=>reset,s=>p(154)(54),cout=>p(155)(55));
FA_ff_1719:FAff port map(x=>p(39)(55),y=>p(40)(55),Cin=>p(41)(55),clock=>clock,reset=>reset,s=>p(154)(55),cout=>p(155)(56));
FA_ff_1720:FAff port map(x=>p(39)(56),y=>p(40)(56),Cin=>p(41)(56),clock=>clock,reset=>reset,s=>p(154)(56),cout=>p(155)(57));
FA_ff_1721:FAff port map(x=>p(39)(57),y=>p(40)(57),Cin=>p(41)(57),clock=>clock,reset=>reset,s=>p(154)(57),cout=>p(155)(58));
FA_ff_1722:FAff port map(x=>p(39)(58),y=>p(40)(58),Cin=>p(41)(58),clock=>clock,reset=>reset,s=>p(154)(58),cout=>p(155)(59));
FA_ff_1723:FAff port map(x=>p(39)(59),y=>p(40)(59),Cin=>p(41)(59),clock=>clock,reset=>reset,s=>p(154)(59),cout=>p(155)(60));
FA_ff_1724:FAff port map(x=>p(39)(60),y=>p(40)(60),Cin=>p(41)(60),clock=>clock,reset=>reset,s=>p(154)(60),cout=>p(155)(61));
FA_ff_1725:FAff port map(x=>p(39)(61),y=>p(40)(61),Cin=>p(41)(61),clock=>clock,reset=>reset,s=>p(154)(61),cout=>p(155)(62));
FA_ff_1726:FAff port map(x=>p(39)(62),y=>p(40)(62),Cin=>p(41)(62),clock=>clock,reset=>reset,s=>p(154)(62),cout=>p(155)(63));
FA_ff_1727:FAff port map(x=>p(39)(63),y=>p(40)(63),Cin=>p(41)(63),clock=>clock,reset=>reset,s=>p(154)(63),cout=>p(155)(64));
FA_ff_1728:FAff port map(x=>p(39)(64),y=>p(40)(64),Cin=>p(41)(64),clock=>clock,reset=>reset,s=>p(154)(64),cout=>p(155)(65));
FA_ff_1729:FAff port map(x=>p(39)(65),y=>p(40)(65),Cin=>p(41)(65),clock=>clock,reset=>reset,s=>p(154)(65),cout=>p(155)(66));
FA_ff_1730:FAff port map(x=>p(39)(66),y=>p(40)(66),Cin=>p(41)(66),clock=>clock,reset=>reset,s=>p(154)(66),cout=>p(155)(67));
FA_ff_1731:FAff port map(x=>p(39)(67),y=>p(40)(67),Cin=>p(41)(67),clock=>clock,reset=>reset,s=>p(154)(67),cout=>p(155)(68));
FA_ff_1732:FAff port map(x=>p(39)(68),y=>p(40)(68),Cin=>p(41)(68),clock=>clock,reset=>reset,s=>p(154)(68),cout=>p(155)(69));
FA_ff_1733:FAff port map(x=>p(39)(69),y=>p(40)(69),Cin=>p(41)(69),clock=>clock,reset=>reset,s=>p(154)(69),cout=>p(155)(70));
FA_ff_1734:FAff port map(x=>p(39)(70),y=>p(40)(70),Cin=>p(41)(70),clock=>clock,reset=>reset,s=>p(154)(70),cout=>p(155)(71));
FA_ff_1735:FAff port map(x=>p(39)(71),y=>p(40)(71),Cin=>p(41)(71),clock=>clock,reset=>reset,s=>p(154)(71),cout=>p(155)(72));
FA_ff_1736:FAff port map(x=>p(39)(72),y=>p(40)(72),Cin=>p(41)(72),clock=>clock,reset=>reset,s=>p(154)(72),cout=>p(155)(73));
FA_ff_1737:FAff port map(x=>p(39)(73),y=>p(40)(73),Cin=>p(41)(73),clock=>clock,reset=>reset,s=>p(154)(73),cout=>p(155)(74));
FA_ff_1738:FAff port map(x=>p(39)(74),y=>p(40)(74),Cin=>p(41)(74),clock=>clock,reset=>reset,s=>p(154)(74),cout=>p(155)(75));
FA_ff_1739:FAff port map(x=>p(39)(75),y=>p(40)(75),Cin=>p(41)(75),clock=>clock,reset=>reset,s=>p(154)(75),cout=>p(155)(76));
FA_ff_1740:FAff port map(x=>p(39)(76),y=>p(40)(76),Cin=>p(41)(76),clock=>clock,reset=>reset,s=>p(154)(76),cout=>p(155)(77));
FA_ff_1741:FAff port map(x=>p(39)(77),y=>p(40)(77),Cin=>p(41)(77),clock=>clock,reset=>reset,s=>p(154)(77),cout=>p(155)(78));
FA_ff_1742:FAff port map(x=>p(39)(78),y=>p(40)(78),Cin=>p(41)(78),clock=>clock,reset=>reset,s=>p(154)(78),cout=>p(155)(79));
FA_ff_1743:FAff port map(x=>p(39)(79),y=>p(40)(79),Cin=>p(41)(79),clock=>clock,reset=>reset,s=>p(154)(79),cout=>p(155)(80));
FA_ff_1744:FAff port map(x=>p(39)(80),y=>p(40)(80),Cin=>p(41)(80),clock=>clock,reset=>reset,s=>p(154)(80),cout=>p(155)(81));
FA_ff_1745:FAff port map(x=>p(39)(81),y=>p(40)(81),Cin=>p(41)(81),clock=>clock,reset=>reset,s=>p(154)(81),cout=>p(155)(82));
FA_ff_1746:FAff port map(x=>p(39)(82),y=>p(40)(82),Cin=>p(41)(82),clock=>clock,reset=>reset,s=>p(154)(82),cout=>p(155)(83));
FA_ff_1747:FAff port map(x=>p(39)(83),y=>p(40)(83),Cin=>p(41)(83),clock=>clock,reset=>reset,s=>p(154)(83),cout=>p(155)(84));
FA_ff_1748:FAff port map(x=>p(39)(84),y=>p(40)(84),Cin=>p(41)(84),clock=>clock,reset=>reset,s=>p(154)(84),cout=>p(155)(85));
FA_ff_1749:FAff port map(x=>p(39)(85),y=>p(40)(85),Cin=>p(41)(85),clock=>clock,reset=>reset,s=>p(154)(85),cout=>p(155)(86));
FA_ff_1750:FAff port map(x=>p(39)(86),y=>p(40)(86),Cin=>p(41)(86),clock=>clock,reset=>reset,s=>p(154)(86),cout=>p(155)(87));
FA_ff_1751:FAff port map(x=>p(39)(87),y=>p(40)(87),Cin=>p(41)(87),clock=>clock,reset=>reset,s=>p(154)(87),cout=>p(155)(88));
FA_ff_1752:FAff port map(x=>p(39)(88),y=>p(40)(88),Cin=>p(41)(88),clock=>clock,reset=>reset,s=>p(154)(88),cout=>p(155)(89));
FA_ff_1753:FAff port map(x=>p(39)(89),y=>p(40)(89),Cin=>p(41)(89),clock=>clock,reset=>reset,s=>p(154)(89),cout=>p(155)(90));
FA_ff_1754:FAff port map(x=>p(39)(90),y=>p(40)(90),Cin=>p(41)(90),clock=>clock,reset=>reset,s=>p(154)(90),cout=>p(155)(91));
FA_ff_1755:FAff port map(x=>p(39)(91),y=>p(40)(91),Cin=>p(41)(91),clock=>clock,reset=>reset,s=>p(154)(91),cout=>p(155)(92));
FA_ff_1756:FAff port map(x=>p(39)(92),y=>p(40)(92),Cin=>p(41)(92),clock=>clock,reset=>reset,s=>p(154)(92),cout=>p(155)(93));
FA_ff_1757:FAff port map(x=>p(39)(93),y=>p(40)(93),Cin=>p(41)(93),clock=>clock,reset=>reset,s=>p(154)(93),cout=>p(155)(94));
FA_ff_1758:FAff port map(x=>p(39)(94),y=>p(40)(94),Cin=>p(41)(94),clock=>clock,reset=>reset,s=>p(154)(94),cout=>p(155)(95));
FA_ff_1759:FAff port map(x=>p(39)(95),y=>p(40)(95),Cin=>p(41)(95),clock=>clock,reset=>reset,s=>p(154)(95),cout=>p(155)(96));
FA_ff_1760:FAff port map(x=>p(39)(96),y=>p(40)(96),Cin=>p(41)(96),clock=>clock,reset=>reset,s=>p(154)(96),cout=>p(155)(97));
FA_ff_1761:FAff port map(x=>p(39)(97),y=>p(40)(97),Cin=>p(41)(97),clock=>clock,reset=>reset,s=>p(154)(97),cout=>p(155)(98));
FA_ff_1762:FAff port map(x=>p(39)(98),y=>p(40)(98),Cin=>p(41)(98),clock=>clock,reset=>reset,s=>p(154)(98),cout=>p(155)(99));
FA_ff_1763:FAff port map(x=>p(39)(99),y=>p(40)(99),Cin=>p(41)(99),clock=>clock,reset=>reset,s=>p(154)(99),cout=>p(155)(100));
FA_ff_1764:FAff port map(x=>p(39)(100),y=>p(40)(100),Cin=>p(41)(100),clock=>clock,reset=>reset,s=>p(154)(100),cout=>p(155)(101));
FA_ff_1765:FAff port map(x=>p(39)(101),y=>p(40)(101),Cin=>p(41)(101),clock=>clock,reset=>reset,s=>p(154)(101),cout=>p(155)(102));
FA_ff_1766:FAff port map(x=>p(39)(102),y=>p(40)(102),Cin=>p(41)(102),clock=>clock,reset=>reset,s=>p(154)(102),cout=>p(155)(103));
FA_ff_1767:FAff port map(x=>p(39)(103),y=>p(40)(103),Cin=>p(41)(103),clock=>clock,reset=>reset,s=>p(154)(103),cout=>p(155)(104));
FA_ff_1768:FAff port map(x=>p(39)(104),y=>p(40)(104),Cin=>p(41)(104),clock=>clock,reset=>reset,s=>p(154)(104),cout=>p(155)(105));
FA_ff_1769:FAff port map(x=>p(39)(105),y=>p(40)(105),Cin=>p(41)(105),clock=>clock,reset=>reset,s=>p(154)(105),cout=>p(155)(106));
FA_ff_1770:FAff port map(x=>p(39)(106),y=>p(40)(106),Cin=>p(41)(106),clock=>clock,reset=>reset,s=>p(154)(106),cout=>p(155)(107));
FA_ff_1771:FAff port map(x=>p(39)(107),y=>p(40)(107),Cin=>p(41)(107),clock=>clock,reset=>reset,s=>p(154)(107),cout=>p(155)(108));
FA_ff_1772:FAff port map(x=>p(39)(108),y=>p(40)(108),Cin=>p(41)(108),clock=>clock,reset=>reset,s=>p(154)(108),cout=>p(155)(109));
FA_ff_1773:FAff port map(x=>p(39)(109),y=>p(40)(109),Cin=>p(41)(109),clock=>clock,reset=>reset,s=>p(154)(109),cout=>p(155)(110));
FA_ff_1774:FAff port map(x=>p(39)(110),y=>p(40)(110),Cin=>p(41)(110),clock=>clock,reset=>reset,s=>p(154)(110),cout=>p(155)(111));
FA_ff_1775:FAff port map(x=>p(39)(111),y=>p(40)(111),Cin=>p(41)(111),clock=>clock,reset=>reset,s=>p(154)(111),cout=>p(155)(112));
FA_ff_1776:FAff port map(x=>p(39)(112),y=>p(40)(112),Cin=>p(41)(112),clock=>clock,reset=>reset,s=>p(154)(112),cout=>p(155)(113));
FA_ff_1777:FAff port map(x=>p(39)(113),y=>p(40)(113),Cin=>p(41)(113),clock=>clock,reset=>reset,s=>p(154)(113),cout=>p(155)(114));
FA_ff_1778:FAff port map(x=>p(39)(114),y=>p(40)(114),Cin=>p(41)(114),clock=>clock,reset=>reset,s=>p(154)(114),cout=>p(155)(115));
FA_ff_1779:FAff port map(x=>p(39)(115),y=>p(40)(115),Cin=>p(41)(115),clock=>clock,reset=>reset,s=>p(154)(115),cout=>p(155)(116));
FA_ff_1780:FAff port map(x=>p(39)(116),y=>p(40)(116),Cin=>p(41)(116),clock=>clock,reset=>reset,s=>p(154)(116),cout=>p(155)(117));
FA_ff_1781:FAff port map(x=>p(39)(117),y=>p(40)(117),Cin=>p(41)(117),clock=>clock,reset=>reset,s=>p(154)(117),cout=>p(155)(118));
FA_ff_1782:FAff port map(x=>p(39)(118),y=>p(40)(118),Cin=>p(41)(118),clock=>clock,reset=>reset,s=>p(154)(118),cout=>p(155)(119));
FA_ff_1783:FAff port map(x=>p(39)(119),y=>p(40)(119),Cin=>p(41)(119),clock=>clock,reset=>reset,s=>p(154)(119),cout=>p(155)(120));
FA_ff_1784:FAff port map(x=>p(39)(120),y=>p(40)(120),Cin=>p(41)(120),clock=>clock,reset=>reset,s=>p(154)(120),cout=>p(155)(121));
FA_ff_1785:FAff port map(x=>p(39)(121),y=>p(40)(121),Cin=>p(41)(121),clock=>clock,reset=>reset,s=>p(154)(121),cout=>p(155)(122));
FA_ff_1786:FAff port map(x=>p(39)(122),y=>p(40)(122),Cin=>p(41)(122),clock=>clock,reset=>reset,s=>p(154)(122),cout=>p(155)(123));
FA_ff_1787:FAff port map(x=>p(39)(123),y=>p(40)(123),Cin=>p(41)(123),clock=>clock,reset=>reset,s=>p(154)(123),cout=>p(155)(124));
FA_ff_1788:FAff port map(x=>p(39)(124),y=>p(40)(124),Cin=>p(41)(124),clock=>clock,reset=>reset,s=>p(154)(124),cout=>p(155)(125));
FA_ff_1789:FAff port map(x=>p(39)(125),y=>p(40)(125),Cin=>p(41)(125),clock=>clock,reset=>reset,s=>p(154)(125),cout=>p(155)(126));
FA_ff_1790:FAff port map(x=>p(39)(126),y=>p(40)(126),Cin=>p(41)(126),clock=>clock,reset=>reset,s=>p(154)(126),cout=>p(155)(127));
FA_ff_1791:FAff port map(x=>p(39)(127),y=>p(40)(127),Cin=>p(41)(127),clock=>clock,reset=>reset,s=>p(154)(127),cout=>p(155)(128));
FA_ff_1792:FAff port map(x=>p(42)(0),y=>p(43)(0),Cin=>p(44)(0),clock=>clock,reset=>reset,s=>p(156)(0),cout=>p(157)(1));
FA_ff_1793:FAff port map(x=>p(42)(1),y=>p(43)(1),Cin=>p(44)(1),clock=>clock,reset=>reset,s=>p(156)(1),cout=>p(157)(2));
FA_ff_1794:FAff port map(x=>p(42)(2),y=>p(43)(2),Cin=>p(44)(2),clock=>clock,reset=>reset,s=>p(156)(2),cout=>p(157)(3));
FA_ff_1795:FAff port map(x=>p(42)(3),y=>p(43)(3),Cin=>p(44)(3),clock=>clock,reset=>reset,s=>p(156)(3),cout=>p(157)(4));
FA_ff_1796:FAff port map(x=>p(42)(4),y=>p(43)(4),Cin=>p(44)(4),clock=>clock,reset=>reset,s=>p(156)(4),cout=>p(157)(5));
FA_ff_1797:FAff port map(x=>p(42)(5),y=>p(43)(5),Cin=>p(44)(5),clock=>clock,reset=>reset,s=>p(156)(5),cout=>p(157)(6));
FA_ff_1798:FAff port map(x=>p(42)(6),y=>p(43)(6),Cin=>p(44)(6),clock=>clock,reset=>reset,s=>p(156)(6),cout=>p(157)(7));
FA_ff_1799:FAff port map(x=>p(42)(7),y=>p(43)(7),Cin=>p(44)(7),clock=>clock,reset=>reset,s=>p(156)(7),cout=>p(157)(8));
FA_ff_1800:FAff port map(x=>p(42)(8),y=>p(43)(8),Cin=>p(44)(8),clock=>clock,reset=>reset,s=>p(156)(8),cout=>p(157)(9));
FA_ff_1801:FAff port map(x=>p(42)(9),y=>p(43)(9),Cin=>p(44)(9),clock=>clock,reset=>reset,s=>p(156)(9),cout=>p(157)(10));
FA_ff_1802:FAff port map(x=>p(42)(10),y=>p(43)(10),Cin=>p(44)(10),clock=>clock,reset=>reset,s=>p(156)(10),cout=>p(157)(11));
FA_ff_1803:FAff port map(x=>p(42)(11),y=>p(43)(11),Cin=>p(44)(11),clock=>clock,reset=>reset,s=>p(156)(11),cout=>p(157)(12));
FA_ff_1804:FAff port map(x=>p(42)(12),y=>p(43)(12),Cin=>p(44)(12),clock=>clock,reset=>reset,s=>p(156)(12),cout=>p(157)(13));
FA_ff_1805:FAff port map(x=>p(42)(13),y=>p(43)(13),Cin=>p(44)(13),clock=>clock,reset=>reset,s=>p(156)(13),cout=>p(157)(14));
FA_ff_1806:FAff port map(x=>p(42)(14),y=>p(43)(14),Cin=>p(44)(14),clock=>clock,reset=>reset,s=>p(156)(14),cout=>p(157)(15));
FA_ff_1807:FAff port map(x=>p(42)(15),y=>p(43)(15),Cin=>p(44)(15),clock=>clock,reset=>reset,s=>p(156)(15),cout=>p(157)(16));
FA_ff_1808:FAff port map(x=>p(42)(16),y=>p(43)(16),Cin=>p(44)(16),clock=>clock,reset=>reset,s=>p(156)(16),cout=>p(157)(17));
FA_ff_1809:FAff port map(x=>p(42)(17),y=>p(43)(17),Cin=>p(44)(17),clock=>clock,reset=>reset,s=>p(156)(17),cout=>p(157)(18));
FA_ff_1810:FAff port map(x=>p(42)(18),y=>p(43)(18),Cin=>p(44)(18),clock=>clock,reset=>reset,s=>p(156)(18),cout=>p(157)(19));
FA_ff_1811:FAff port map(x=>p(42)(19),y=>p(43)(19),Cin=>p(44)(19),clock=>clock,reset=>reset,s=>p(156)(19),cout=>p(157)(20));
FA_ff_1812:FAff port map(x=>p(42)(20),y=>p(43)(20),Cin=>p(44)(20),clock=>clock,reset=>reset,s=>p(156)(20),cout=>p(157)(21));
FA_ff_1813:FAff port map(x=>p(42)(21),y=>p(43)(21),Cin=>p(44)(21),clock=>clock,reset=>reset,s=>p(156)(21),cout=>p(157)(22));
FA_ff_1814:FAff port map(x=>p(42)(22),y=>p(43)(22),Cin=>p(44)(22),clock=>clock,reset=>reset,s=>p(156)(22),cout=>p(157)(23));
FA_ff_1815:FAff port map(x=>p(42)(23),y=>p(43)(23),Cin=>p(44)(23),clock=>clock,reset=>reset,s=>p(156)(23),cout=>p(157)(24));
FA_ff_1816:FAff port map(x=>p(42)(24),y=>p(43)(24),Cin=>p(44)(24),clock=>clock,reset=>reset,s=>p(156)(24),cout=>p(157)(25));
FA_ff_1817:FAff port map(x=>p(42)(25),y=>p(43)(25),Cin=>p(44)(25),clock=>clock,reset=>reset,s=>p(156)(25),cout=>p(157)(26));
FA_ff_1818:FAff port map(x=>p(42)(26),y=>p(43)(26),Cin=>p(44)(26),clock=>clock,reset=>reset,s=>p(156)(26),cout=>p(157)(27));
FA_ff_1819:FAff port map(x=>p(42)(27),y=>p(43)(27),Cin=>p(44)(27),clock=>clock,reset=>reset,s=>p(156)(27),cout=>p(157)(28));
FA_ff_1820:FAff port map(x=>p(42)(28),y=>p(43)(28),Cin=>p(44)(28),clock=>clock,reset=>reset,s=>p(156)(28),cout=>p(157)(29));
FA_ff_1821:FAff port map(x=>p(42)(29),y=>p(43)(29),Cin=>p(44)(29),clock=>clock,reset=>reset,s=>p(156)(29),cout=>p(157)(30));
FA_ff_1822:FAff port map(x=>p(42)(30),y=>p(43)(30),Cin=>p(44)(30),clock=>clock,reset=>reset,s=>p(156)(30),cout=>p(157)(31));
FA_ff_1823:FAff port map(x=>p(42)(31),y=>p(43)(31),Cin=>p(44)(31),clock=>clock,reset=>reset,s=>p(156)(31),cout=>p(157)(32));
FA_ff_1824:FAff port map(x=>p(42)(32),y=>p(43)(32),Cin=>p(44)(32),clock=>clock,reset=>reset,s=>p(156)(32),cout=>p(157)(33));
FA_ff_1825:FAff port map(x=>p(42)(33),y=>p(43)(33),Cin=>p(44)(33),clock=>clock,reset=>reset,s=>p(156)(33),cout=>p(157)(34));
FA_ff_1826:FAff port map(x=>p(42)(34),y=>p(43)(34),Cin=>p(44)(34),clock=>clock,reset=>reset,s=>p(156)(34),cout=>p(157)(35));
FA_ff_1827:FAff port map(x=>p(42)(35),y=>p(43)(35),Cin=>p(44)(35),clock=>clock,reset=>reset,s=>p(156)(35),cout=>p(157)(36));
FA_ff_1828:FAff port map(x=>p(42)(36),y=>p(43)(36),Cin=>p(44)(36),clock=>clock,reset=>reset,s=>p(156)(36),cout=>p(157)(37));
FA_ff_1829:FAff port map(x=>p(42)(37),y=>p(43)(37),Cin=>p(44)(37),clock=>clock,reset=>reset,s=>p(156)(37),cout=>p(157)(38));
FA_ff_1830:FAff port map(x=>p(42)(38),y=>p(43)(38),Cin=>p(44)(38),clock=>clock,reset=>reset,s=>p(156)(38),cout=>p(157)(39));
FA_ff_1831:FAff port map(x=>p(42)(39),y=>p(43)(39),Cin=>p(44)(39),clock=>clock,reset=>reset,s=>p(156)(39),cout=>p(157)(40));
FA_ff_1832:FAff port map(x=>p(42)(40),y=>p(43)(40),Cin=>p(44)(40),clock=>clock,reset=>reset,s=>p(156)(40),cout=>p(157)(41));
FA_ff_1833:FAff port map(x=>p(42)(41),y=>p(43)(41),Cin=>p(44)(41),clock=>clock,reset=>reset,s=>p(156)(41),cout=>p(157)(42));
FA_ff_1834:FAff port map(x=>p(42)(42),y=>p(43)(42),Cin=>p(44)(42),clock=>clock,reset=>reset,s=>p(156)(42),cout=>p(157)(43));
FA_ff_1835:FAff port map(x=>p(42)(43),y=>p(43)(43),Cin=>p(44)(43),clock=>clock,reset=>reset,s=>p(156)(43),cout=>p(157)(44));
FA_ff_1836:FAff port map(x=>p(42)(44),y=>p(43)(44),Cin=>p(44)(44),clock=>clock,reset=>reset,s=>p(156)(44),cout=>p(157)(45));
FA_ff_1837:FAff port map(x=>p(42)(45),y=>p(43)(45),Cin=>p(44)(45),clock=>clock,reset=>reset,s=>p(156)(45),cout=>p(157)(46));
FA_ff_1838:FAff port map(x=>p(42)(46),y=>p(43)(46),Cin=>p(44)(46),clock=>clock,reset=>reset,s=>p(156)(46),cout=>p(157)(47));
FA_ff_1839:FAff port map(x=>p(42)(47),y=>p(43)(47),Cin=>p(44)(47),clock=>clock,reset=>reset,s=>p(156)(47),cout=>p(157)(48));
FA_ff_1840:FAff port map(x=>p(42)(48),y=>p(43)(48),Cin=>p(44)(48),clock=>clock,reset=>reset,s=>p(156)(48),cout=>p(157)(49));
FA_ff_1841:FAff port map(x=>p(42)(49),y=>p(43)(49),Cin=>p(44)(49),clock=>clock,reset=>reset,s=>p(156)(49),cout=>p(157)(50));
FA_ff_1842:FAff port map(x=>p(42)(50),y=>p(43)(50),Cin=>p(44)(50),clock=>clock,reset=>reset,s=>p(156)(50),cout=>p(157)(51));
FA_ff_1843:FAff port map(x=>p(42)(51),y=>p(43)(51),Cin=>p(44)(51),clock=>clock,reset=>reset,s=>p(156)(51),cout=>p(157)(52));
FA_ff_1844:FAff port map(x=>p(42)(52),y=>p(43)(52),Cin=>p(44)(52),clock=>clock,reset=>reset,s=>p(156)(52),cout=>p(157)(53));
FA_ff_1845:FAff port map(x=>p(42)(53),y=>p(43)(53),Cin=>p(44)(53),clock=>clock,reset=>reset,s=>p(156)(53),cout=>p(157)(54));
FA_ff_1846:FAff port map(x=>p(42)(54),y=>p(43)(54),Cin=>p(44)(54),clock=>clock,reset=>reset,s=>p(156)(54),cout=>p(157)(55));
FA_ff_1847:FAff port map(x=>p(42)(55),y=>p(43)(55),Cin=>p(44)(55),clock=>clock,reset=>reset,s=>p(156)(55),cout=>p(157)(56));
FA_ff_1848:FAff port map(x=>p(42)(56),y=>p(43)(56),Cin=>p(44)(56),clock=>clock,reset=>reset,s=>p(156)(56),cout=>p(157)(57));
FA_ff_1849:FAff port map(x=>p(42)(57),y=>p(43)(57),Cin=>p(44)(57),clock=>clock,reset=>reset,s=>p(156)(57),cout=>p(157)(58));
FA_ff_1850:FAff port map(x=>p(42)(58),y=>p(43)(58),Cin=>p(44)(58),clock=>clock,reset=>reset,s=>p(156)(58),cout=>p(157)(59));
FA_ff_1851:FAff port map(x=>p(42)(59),y=>p(43)(59),Cin=>p(44)(59),clock=>clock,reset=>reset,s=>p(156)(59),cout=>p(157)(60));
FA_ff_1852:FAff port map(x=>p(42)(60),y=>p(43)(60),Cin=>p(44)(60),clock=>clock,reset=>reset,s=>p(156)(60),cout=>p(157)(61));
FA_ff_1853:FAff port map(x=>p(42)(61),y=>p(43)(61),Cin=>p(44)(61),clock=>clock,reset=>reset,s=>p(156)(61),cout=>p(157)(62));
FA_ff_1854:FAff port map(x=>p(42)(62),y=>p(43)(62),Cin=>p(44)(62),clock=>clock,reset=>reset,s=>p(156)(62),cout=>p(157)(63));
FA_ff_1855:FAff port map(x=>p(42)(63),y=>p(43)(63),Cin=>p(44)(63),clock=>clock,reset=>reset,s=>p(156)(63),cout=>p(157)(64));
FA_ff_1856:FAff port map(x=>p(42)(64),y=>p(43)(64),Cin=>p(44)(64),clock=>clock,reset=>reset,s=>p(156)(64),cout=>p(157)(65));
FA_ff_1857:FAff port map(x=>p(42)(65),y=>p(43)(65),Cin=>p(44)(65),clock=>clock,reset=>reset,s=>p(156)(65),cout=>p(157)(66));
FA_ff_1858:FAff port map(x=>p(42)(66),y=>p(43)(66),Cin=>p(44)(66),clock=>clock,reset=>reset,s=>p(156)(66),cout=>p(157)(67));
FA_ff_1859:FAff port map(x=>p(42)(67),y=>p(43)(67),Cin=>p(44)(67),clock=>clock,reset=>reset,s=>p(156)(67),cout=>p(157)(68));
FA_ff_1860:FAff port map(x=>p(42)(68),y=>p(43)(68),Cin=>p(44)(68),clock=>clock,reset=>reset,s=>p(156)(68),cout=>p(157)(69));
FA_ff_1861:FAff port map(x=>p(42)(69),y=>p(43)(69),Cin=>p(44)(69),clock=>clock,reset=>reset,s=>p(156)(69),cout=>p(157)(70));
FA_ff_1862:FAff port map(x=>p(42)(70),y=>p(43)(70),Cin=>p(44)(70),clock=>clock,reset=>reset,s=>p(156)(70),cout=>p(157)(71));
FA_ff_1863:FAff port map(x=>p(42)(71),y=>p(43)(71),Cin=>p(44)(71),clock=>clock,reset=>reset,s=>p(156)(71),cout=>p(157)(72));
FA_ff_1864:FAff port map(x=>p(42)(72),y=>p(43)(72),Cin=>p(44)(72),clock=>clock,reset=>reset,s=>p(156)(72),cout=>p(157)(73));
FA_ff_1865:FAff port map(x=>p(42)(73),y=>p(43)(73),Cin=>p(44)(73),clock=>clock,reset=>reset,s=>p(156)(73),cout=>p(157)(74));
FA_ff_1866:FAff port map(x=>p(42)(74),y=>p(43)(74),Cin=>p(44)(74),clock=>clock,reset=>reset,s=>p(156)(74),cout=>p(157)(75));
FA_ff_1867:FAff port map(x=>p(42)(75),y=>p(43)(75),Cin=>p(44)(75),clock=>clock,reset=>reset,s=>p(156)(75),cout=>p(157)(76));
FA_ff_1868:FAff port map(x=>p(42)(76),y=>p(43)(76),Cin=>p(44)(76),clock=>clock,reset=>reset,s=>p(156)(76),cout=>p(157)(77));
FA_ff_1869:FAff port map(x=>p(42)(77),y=>p(43)(77),Cin=>p(44)(77),clock=>clock,reset=>reset,s=>p(156)(77),cout=>p(157)(78));
FA_ff_1870:FAff port map(x=>p(42)(78),y=>p(43)(78),Cin=>p(44)(78),clock=>clock,reset=>reset,s=>p(156)(78),cout=>p(157)(79));
FA_ff_1871:FAff port map(x=>p(42)(79),y=>p(43)(79),Cin=>p(44)(79),clock=>clock,reset=>reset,s=>p(156)(79),cout=>p(157)(80));
FA_ff_1872:FAff port map(x=>p(42)(80),y=>p(43)(80),Cin=>p(44)(80),clock=>clock,reset=>reset,s=>p(156)(80),cout=>p(157)(81));
FA_ff_1873:FAff port map(x=>p(42)(81),y=>p(43)(81),Cin=>p(44)(81),clock=>clock,reset=>reset,s=>p(156)(81),cout=>p(157)(82));
FA_ff_1874:FAff port map(x=>p(42)(82),y=>p(43)(82),Cin=>p(44)(82),clock=>clock,reset=>reset,s=>p(156)(82),cout=>p(157)(83));
FA_ff_1875:FAff port map(x=>p(42)(83),y=>p(43)(83),Cin=>p(44)(83),clock=>clock,reset=>reset,s=>p(156)(83),cout=>p(157)(84));
FA_ff_1876:FAff port map(x=>p(42)(84),y=>p(43)(84),Cin=>p(44)(84),clock=>clock,reset=>reset,s=>p(156)(84),cout=>p(157)(85));
FA_ff_1877:FAff port map(x=>p(42)(85),y=>p(43)(85),Cin=>p(44)(85),clock=>clock,reset=>reset,s=>p(156)(85),cout=>p(157)(86));
FA_ff_1878:FAff port map(x=>p(42)(86),y=>p(43)(86),Cin=>p(44)(86),clock=>clock,reset=>reset,s=>p(156)(86),cout=>p(157)(87));
FA_ff_1879:FAff port map(x=>p(42)(87),y=>p(43)(87),Cin=>p(44)(87),clock=>clock,reset=>reset,s=>p(156)(87),cout=>p(157)(88));
FA_ff_1880:FAff port map(x=>p(42)(88),y=>p(43)(88),Cin=>p(44)(88),clock=>clock,reset=>reset,s=>p(156)(88),cout=>p(157)(89));
FA_ff_1881:FAff port map(x=>p(42)(89),y=>p(43)(89),Cin=>p(44)(89),clock=>clock,reset=>reset,s=>p(156)(89),cout=>p(157)(90));
FA_ff_1882:FAff port map(x=>p(42)(90),y=>p(43)(90),Cin=>p(44)(90),clock=>clock,reset=>reset,s=>p(156)(90),cout=>p(157)(91));
FA_ff_1883:FAff port map(x=>p(42)(91),y=>p(43)(91),Cin=>p(44)(91),clock=>clock,reset=>reset,s=>p(156)(91),cout=>p(157)(92));
FA_ff_1884:FAff port map(x=>p(42)(92),y=>p(43)(92),Cin=>p(44)(92),clock=>clock,reset=>reset,s=>p(156)(92),cout=>p(157)(93));
FA_ff_1885:FAff port map(x=>p(42)(93),y=>p(43)(93),Cin=>p(44)(93),clock=>clock,reset=>reset,s=>p(156)(93),cout=>p(157)(94));
FA_ff_1886:FAff port map(x=>p(42)(94),y=>p(43)(94),Cin=>p(44)(94),clock=>clock,reset=>reset,s=>p(156)(94),cout=>p(157)(95));
FA_ff_1887:FAff port map(x=>p(42)(95),y=>p(43)(95),Cin=>p(44)(95),clock=>clock,reset=>reset,s=>p(156)(95),cout=>p(157)(96));
FA_ff_1888:FAff port map(x=>p(42)(96),y=>p(43)(96),Cin=>p(44)(96),clock=>clock,reset=>reset,s=>p(156)(96),cout=>p(157)(97));
FA_ff_1889:FAff port map(x=>p(42)(97),y=>p(43)(97),Cin=>p(44)(97),clock=>clock,reset=>reset,s=>p(156)(97),cout=>p(157)(98));
FA_ff_1890:FAff port map(x=>p(42)(98),y=>p(43)(98),Cin=>p(44)(98),clock=>clock,reset=>reset,s=>p(156)(98),cout=>p(157)(99));
FA_ff_1891:FAff port map(x=>p(42)(99),y=>p(43)(99),Cin=>p(44)(99),clock=>clock,reset=>reset,s=>p(156)(99),cout=>p(157)(100));
FA_ff_1892:FAff port map(x=>p(42)(100),y=>p(43)(100),Cin=>p(44)(100),clock=>clock,reset=>reset,s=>p(156)(100),cout=>p(157)(101));
FA_ff_1893:FAff port map(x=>p(42)(101),y=>p(43)(101),Cin=>p(44)(101),clock=>clock,reset=>reset,s=>p(156)(101),cout=>p(157)(102));
FA_ff_1894:FAff port map(x=>p(42)(102),y=>p(43)(102),Cin=>p(44)(102),clock=>clock,reset=>reset,s=>p(156)(102),cout=>p(157)(103));
FA_ff_1895:FAff port map(x=>p(42)(103),y=>p(43)(103),Cin=>p(44)(103),clock=>clock,reset=>reset,s=>p(156)(103),cout=>p(157)(104));
FA_ff_1896:FAff port map(x=>p(42)(104),y=>p(43)(104),Cin=>p(44)(104),clock=>clock,reset=>reset,s=>p(156)(104),cout=>p(157)(105));
FA_ff_1897:FAff port map(x=>p(42)(105),y=>p(43)(105),Cin=>p(44)(105),clock=>clock,reset=>reset,s=>p(156)(105),cout=>p(157)(106));
FA_ff_1898:FAff port map(x=>p(42)(106),y=>p(43)(106),Cin=>p(44)(106),clock=>clock,reset=>reset,s=>p(156)(106),cout=>p(157)(107));
FA_ff_1899:FAff port map(x=>p(42)(107),y=>p(43)(107),Cin=>p(44)(107),clock=>clock,reset=>reset,s=>p(156)(107),cout=>p(157)(108));
FA_ff_1900:FAff port map(x=>p(42)(108),y=>p(43)(108),Cin=>p(44)(108),clock=>clock,reset=>reset,s=>p(156)(108),cout=>p(157)(109));
FA_ff_1901:FAff port map(x=>p(42)(109),y=>p(43)(109),Cin=>p(44)(109),clock=>clock,reset=>reset,s=>p(156)(109),cout=>p(157)(110));
FA_ff_1902:FAff port map(x=>p(42)(110),y=>p(43)(110),Cin=>p(44)(110),clock=>clock,reset=>reset,s=>p(156)(110),cout=>p(157)(111));
FA_ff_1903:FAff port map(x=>p(42)(111),y=>p(43)(111),Cin=>p(44)(111),clock=>clock,reset=>reset,s=>p(156)(111),cout=>p(157)(112));
FA_ff_1904:FAff port map(x=>p(42)(112),y=>p(43)(112),Cin=>p(44)(112),clock=>clock,reset=>reset,s=>p(156)(112),cout=>p(157)(113));
FA_ff_1905:FAff port map(x=>p(42)(113),y=>p(43)(113),Cin=>p(44)(113),clock=>clock,reset=>reset,s=>p(156)(113),cout=>p(157)(114));
FA_ff_1906:FAff port map(x=>p(42)(114),y=>p(43)(114),Cin=>p(44)(114),clock=>clock,reset=>reset,s=>p(156)(114),cout=>p(157)(115));
FA_ff_1907:FAff port map(x=>p(42)(115),y=>p(43)(115),Cin=>p(44)(115),clock=>clock,reset=>reset,s=>p(156)(115),cout=>p(157)(116));
FA_ff_1908:FAff port map(x=>p(42)(116),y=>p(43)(116),Cin=>p(44)(116),clock=>clock,reset=>reset,s=>p(156)(116),cout=>p(157)(117));
FA_ff_1909:FAff port map(x=>p(42)(117),y=>p(43)(117),Cin=>p(44)(117),clock=>clock,reset=>reset,s=>p(156)(117),cout=>p(157)(118));
FA_ff_1910:FAff port map(x=>p(42)(118),y=>p(43)(118),Cin=>p(44)(118),clock=>clock,reset=>reset,s=>p(156)(118),cout=>p(157)(119));
FA_ff_1911:FAff port map(x=>p(42)(119),y=>p(43)(119),Cin=>p(44)(119),clock=>clock,reset=>reset,s=>p(156)(119),cout=>p(157)(120));
FA_ff_1912:FAff port map(x=>p(42)(120),y=>p(43)(120),Cin=>p(44)(120),clock=>clock,reset=>reset,s=>p(156)(120),cout=>p(157)(121));
FA_ff_1913:FAff port map(x=>p(42)(121),y=>p(43)(121),Cin=>p(44)(121),clock=>clock,reset=>reset,s=>p(156)(121),cout=>p(157)(122));
FA_ff_1914:FAff port map(x=>p(42)(122),y=>p(43)(122),Cin=>p(44)(122),clock=>clock,reset=>reset,s=>p(156)(122),cout=>p(157)(123));
FA_ff_1915:FAff port map(x=>p(42)(123),y=>p(43)(123),Cin=>p(44)(123),clock=>clock,reset=>reset,s=>p(156)(123),cout=>p(157)(124));
FA_ff_1916:FAff port map(x=>p(42)(124),y=>p(43)(124),Cin=>p(44)(124),clock=>clock,reset=>reset,s=>p(156)(124),cout=>p(157)(125));
FA_ff_1917:FAff port map(x=>p(42)(125),y=>p(43)(125),Cin=>p(44)(125),clock=>clock,reset=>reset,s=>p(156)(125),cout=>p(157)(126));
FA_ff_1918:FAff port map(x=>p(42)(126),y=>p(43)(126),Cin=>p(44)(126),clock=>clock,reset=>reset,s=>p(156)(126),cout=>p(157)(127));
FA_ff_1919:FAff port map(x=>p(42)(127),y=>p(43)(127),Cin=>p(44)(127),clock=>clock,reset=>reset,s=>p(156)(127),cout=>p(157)(128));
FA_ff_1920:FAff port map(x=>p(45)(0),y=>p(46)(0),Cin=>p(47)(0),clock=>clock,reset=>reset,s=>p(158)(0),cout=>p(159)(1));
FA_ff_1921:FAff port map(x=>p(45)(1),y=>p(46)(1),Cin=>p(47)(1),clock=>clock,reset=>reset,s=>p(158)(1),cout=>p(159)(2));
FA_ff_1922:FAff port map(x=>p(45)(2),y=>p(46)(2),Cin=>p(47)(2),clock=>clock,reset=>reset,s=>p(158)(2),cout=>p(159)(3));
FA_ff_1923:FAff port map(x=>p(45)(3),y=>p(46)(3),Cin=>p(47)(3),clock=>clock,reset=>reset,s=>p(158)(3),cout=>p(159)(4));
FA_ff_1924:FAff port map(x=>p(45)(4),y=>p(46)(4),Cin=>p(47)(4),clock=>clock,reset=>reset,s=>p(158)(4),cout=>p(159)(5));
FA_ff_1925:FAff port map(x=>p(45)(5),y=>p(46)(5),Cin=>p(47)(5),clock=>clock,reset=>reset,s=>p(158)(5),cout=>p(159)(6));
FA_ff_1926:FAff port map(x=>p(45)(6),y=>p(46)(6),Cin=>p(47)(6),clock=>clock,reset=>reset,s=>p(158)(6),cout=>p(159)(7));
FA_ff_1927:FAff port map(x=>p(45)(7),y=>p(46)(7),Cin=>p(47)(7),clock=>clock,reset=>reset,s=>p(158)(7),cout=>p(159)(8));
FA_ff_1928:FAff port map(x=>p(45)(8),y=>p(46)(8),Cin=>p(47)(8),clock=>clock,reset=>reset,s=>p(158)(8),cout=>p(159)(9));
FA_ff_1929:FAff port map(x=>p(45)(9),y=>p(46)(9),Cin=>p(47)(9),clock=>clock,reset=>reset,s=>p(158)(9),cout=>p(159)(10));
FA_ff_1930:FAff port map(x=>p(45)(10),y=>p(46)(10),Cin=>p(47)(10),clock=>clock,reset=>reset,s=>p(158)(10),cout=>p(159)(11));
FA_ff_1931:FAff port map(x=>p(45)(11),y=>p(46)(11),Cin=>p(47)(11),clock=>clock,reset=>reset,s=>p(158)(11),cout=>p(159)(12));
FA_ff_1932:FAff port map(x=>p(45)(12),y=>p(46)(12),Cin=>p(47)(12),clock=>clock,reset=>reset,s=>p(158)(12),cout=>p(159)(13));
FA_ff_1933:FAff port map(x=>p(45)(13),y=>p(46)(13),Cin=>p(47)(13),clock=>clock,reset=>reset,s=>p(158)(13),cout=>p(159)(14));
FA_ff_1934:FAff port map(x=>p(45)(14),y=>p(46)(14),Cin=>p(47)(14),clock=>clock,reset=>reset,s=>p(158)(14),cout=>p(159)(15));
FA_ff_1935:FAff port map(x=>p(45)(15),y=>p(46)(15),Cin=>p(47)(15),clock=>clock,reset=>reset,s=>p(158)(15),cout=>p(159)(16));
FA_ff_1936:FAff port map(x=>p(45)(16),y=>p(46)(16),Cin=>p(47)(16),clock=>clock,reset=>reset,s=>p(158)(16),cout=>p(159)(17));
FA_ff_1937:FAff port map(x=>p(45)(17),y=>p(46)(17),Cin=>p(47)(17),clock=>clock,reset=>reset,s=>p(158)(17),cout=>p(159)(18));
FA_ff_1938:FAff port map(x=>p(45)(18),y=>p(46)(18),Cin=>p(47)(18),clock=>clock,reset=>reset,s=>p(158)(18),cout=>p(159)(19));
FA_ff_1939:FAff port map(x=>p(45)(19),y=>p(46)(19),Cin=>p(47)(19),clock=>clock,reset=>reset,s=>p(158)(19),cout=>p(159)(20));
FA_ff_1940:FAff port map(x=>p(45)(20),y=>p(46)(20),Cin=>p(47)(20),clock=>clock,reset=>reset,s=>p(158)(20),cout=>p(159)(21));
FA_ff_1941:FAff port map(x=>p(45)(21),y=>p(46)(21),Cin=>p(47)(21),clock=>clock,reset=>reset,s=>p(158)(21),cout=>p(159)(22));
FA_ff_1942:FAff port map(x=>p(45)(22),y=>p(46)(22),Cin=>p(47)(22),clock=>clock,reset=>reset,s=>p(158)(22),cout=>p(159)(23));
FA_ff_1943:FAff port map(x=>p(45)(23),y=>p(46)(23),Cin=>p(47)(23),clock=>clock,reset=>reset,s=>p(158)(23),cout=>p(159)(24));
FA_ff_1944:FAff port map(x=>p(45)(24),y=>p(46)(24),Cin=>p(47)(24),clock=>clock,reset=>reset,s=>p(158)(24),cout=>p(159)(25));
FA_ff_1945:FAff port map(x=>p(45)(25),y=>p(46)(25),Cin=>p(47)(25),clock=>clock,reset=>reset,s=>p(158)(25),cout=>p(159)(26));
FA_ff_1946:FAff port map(x=>p(45)(26),y=>p(46)(26),Cin=>p(47)(26),clock=>clock,reset=>reset,s=>p(158)(26),cout=>p(159)(27));
FA_ff_1947:FAff port map(x=>p(45)(27),y=>p(46)(27),Cin=>p(47)(27),clock=>clock,reset=>reset,s=>p(158)(27),cout=>p(159)(28));
FA_ff_1948:FAff port map(x=>p(45)(28),y=>p(46)(28),Cin=>p(47)(28),clock=>clock,reset=>reset,s=>p(158)(28),cout=>p(159)(29));
FA_ff_1949:FAff port map(x=>p(45)(29),y=>p(46)(29),Cin=>p(47)(29),clock=>clock,reset=>reset,s=>p(158)(29),cout=>p(159)(30));
FA_ff_1950:FAff port map(x=>p(45)(30),y=>p(46)(30),Cin=>p(47)(30),clock=>clock,reset=>reset,s=>p(158)(30),cout=>p(159)(31));
FA_ff_1951:FAff port map(x=>p(45)(31),y=>p(46)(31),Cin=>p(47)(31),clock=>clock,reset=>reset,s=>p(158)(31),cout=>p(159)(32));
FA_ff_1952:FAff port map(x=>p(45)(32),y=>p(46)(32),Cin=>p(47)(32),clock=>clock,reset=>reset,s=>p(158)(32),cout=>p(159)(33));
FA_ff_1953:FAff port map(x=>p(45)(33),y=>p(46)(33),Cin=>p(47)(33),clock=>clock,reset=>reset,s=>p(158)(33),cout=>p(159)(34));
FA_ff_1954:FAff port map(x=>p(45)(34),y=>p(46)(34),Cin=>p(47)(34),clock=>clock,reset=>reset,s=>p(158)(34),cout=>p(159)(35));
FA_ff_1955:FAff port map(x=>p(45)(35),y=>p(46)(35),Cin=>p(47)(35),clock=>clock,reset=>reset,s=>p(158)(35),cout=>p(159)(36));
FA_ff_1956:FAff port map(x=>p(45)(36),y=>p(46)(36),Cin=>p(47)(36),clock=>clock,reset=>reset,s=>p(158)(36),cout=>p(159)(37));
FA_ff_1957:FAff port map(x=>p(45)(37),y=>p(46)(37),Cin=>p(47)(37),clock=>clock,reset=>reset,s=>p(158)(37),cout=>p(159)(38));
FA_ff_1958:FAff port map(x=>p(45)(38),y=>p(46)(38),Cin=>p(47)(38),clock=>clock,reset=>reset,s=>p(158)(38),cout=>p(159)(39));
FA_ff_1959:FAff port map(x=>p(45)(39),y=>p(46)(39),Cin=>p(47)(39),clock=>clock,reset=>reset,s=>p(158)(39),cout=>p(159)(40));
FA_ff_1960:FAff port map(x=>p(45)(40),y=>p(46)(40),Cin=>p(47)(40),clock=>clock,reset=>reset,s=>p(158)(40),cout=>p(159)(41));
FA_ff_1961:FAff port map(x=>p(45)(41),y=>p(46)(41),Cin=>p(47)(41),clock=>clock,reset=>reset,s=>p(158)(41),cout=>p(159)(42));
FA_ff_1962:FAff port map(x=>p(45)(42),y=>p(46)(42),Cin=>p(47)(42),clock=>clock,reset=>reset,s=>p(158)(42),cout=>p(159)(43));
FA_ff_1963:FAff port map(x=>p(45)(43),y=>p(46)(43),Cin=>p(47)(43),clock=>clock,reset=>reset,s=>p(158)(43),cout=>p(159)(44));
FA_ff_1964:FAff port map(x=>p(45)(44),y=>p(46)(44),Cin=>p(47)(44),clock=>clock,reset=>reset,s=>p(158)(44),cout=>p(159)(45));
FA_ff_1965:FAff port map(x=>p(45)(45),y=>p(46)(45),Cin=>p(47)(45),clock=>clock,reset=>reset,s=>p(158)(45),cout=>p(159)(46));
FA_ff_1966:FAff port map(x=>p(45)(46),y=>p(46)(46),Cin=>p(47)(46),clock=>clock,reset=>reset,s=>p(158)(46),cout=>p(159)(47));
FA_ff_1967:FAff port map(x=>p(45)(47),y=>p(46)(47),Cin=>p(47)(47),clock=>clock,reset=>reset,s=>p(158)(47),cout=>p(159)(48));
FA_ff_1968:FAff port map(x=>p(45)(48),y=>p(46)(48),Cin=>p(47)(48),clock=>clock,reset=>reset,s=>p(158)(48),cout=>p(159)(49));
FA_ff_1969:FAff port map(x=>p(45)(49),y=>p(46)(49),Cin=>p(47)(49),clock=>clock,reset=>reset,s=>p(158)(49),cout=>p(159)(50));
FA_ff_1970:FAff port map(x=>p(45)(50),y=>p(46)(50),Cin=>p(47)(50),clock=>clock,reset=>reset,s=>p(158)(50),cout=>p(159)(51));
FA_ff_1971:FAff port map(x=>p(45)(51),y=>p(46)(51),Cin=>p(47)(51),clock=>clock,reset=>reset,s=>p(158)(51),cout=>p(159)(52));
FA_ff_1972:FAff port map(x=>p(45)(52),y=>p(46)(52),Cin=>p(47)(52),clock=>clock,reset=>reset,s=>p(158)(52),cout=>p(159)(53));
FA_ff_1973:FAff port map(x=>p(45)(53),y=>p(46)(53),Cin=>p(47)(53),clock=>clock,reset=>reset,s=>p(158)(53),cout=>p(159)(54));
FA_ff_1974:FAff port map(x=>p(45)(54),y=>p(46)(54),Cin=>p(47)(54),clock=>clock,reset=>reset,s=>p(158)(54),cout=>p(159)(55));
FA_ff_1975:FAff port map(x=>p(45)(55),y=>p(46)(55),Cin=>p(47)(55),clock=>clock,reset=>reset,s=>p(158)(55),cout=>p(159)(56));
FA_ff_1976:FAff port map(x=>p(45)(56),y=>p(46)(56),Cin=>p(47)(56),clock=>clock,reset=>reset,s=>p(158)(56),cout=>p(159)(57));
FA_ff_1977:FAff port map(x=>p(45)(57),y=>p(46)(57),Cin=>p(47)(57),clock=>clock,reset=>reset,s=>p(158)(57),cout=>p(159)(58));
FA_ff_1978:FAff port map(x=>p(45)(58),y=>p(46)(58),Cin=>p(47)(58),clock=>clock,reset=>reset,s=>p(158)(58),cout=>p(159)(59));
FA_ff_1979:FAff port map(x=>p(45)(59),y=>p(46)(59),Cin=>p(47)(59),clock=>clock,reset=>reset,s=>p(158)(59),cout=>p(159)(60));
FA_ff_1980:FAff port map(x=>p(45)(60),y=>p(46)(60),Cin=>p(47)(60),clock=>clock,reset=>reset,s=>p(158)(60),cout=>p(159)(61));
FA_ff_1981:FAff port map(x=>p(45)(61),y=>p(46)(61),Cin=>p(47)(61),clock=>clock,reset=>reset,s=>p(158)(61),cout=>p(159)(62));
FA_ff_1982:FAff port map(x=>p(45)(62),y=>p(46)(62),Cin=>p(47)(62),clock=>clock,reset=>reset,s=>p(158)(62),cout=>p(159)(63));
FA_ff_1983:FAff port map(x=>p(45)(63),y=>p(46)(63),Cin=>p(47)(63),clock=>clock,reset=>reset,s=>p(158)(63),cout=>p(159)(64));
FA_ff_1984:FAff port map(x=>p(45)(64),y=>p(46)(64),Cin=>p(47)(64),clock=>clock,reset=>reset,s=>p(158)(64),cout=>p(159)(65));
FA_ff_1985:FAff port map(x=>p(45)(65),y=>p(46)(65),Cin=>p(47)(65),clock=>clock,reset=>reset,s=>p(158)(65),cout=>p(159)(66));
FA_ff_1986:FAff port map(x=>p(45)(66),y=>p(46)(66),Cin=>p(47)(66),clock=>clock,reset=>reset,s=>p(158)(66),cout=>p(159)(67));
FA_ff_1987:FAff port map(x=>p(45)(67),y=>p(46)(67),Cin=>p(47)(67),clock=>clock,reset=>reset,s=>p(158)(67),cout=>p(159)(68));
FA_ff_1988:FAff port map(x=>p(45)(68),y=>p(46)(68),Cin=>p(47)(68),clock=>clock,reset=>reset,s=>p(158)(68),cout=>p(159)(69));
FA_ff_1989:FAff port map(x=>p(45)(69),y=>p(46)(69),Cin=>p(47)(69),clock=>clock,reset=>reset,s=>p(158)(69),cout=>p(159)(70));
FA_ff_1990:FAff port map(x=>p(45)(70),y=>p(46)(70),Cin=>p(47)(70),clock=>clock,reset=>reset,s=>p(158)(70),cout=>p(159)(71));
FA_ff_1991:FAff port map(x=>p(45)(71),y=>p(46)(71),Cin=>p(47)(71),clock=>clock,reset=>reset,s=>p(158)(71),cout=>p(159)(72));
FA_ff_1992:FAff port map(x=>p(45)(72),y=>p(46)(72),Cin=>p(47)(72),clock=>clock,reset=>reset,s=>p(158)(72),cout=>p(159)(73));
FA_ff_1993:FAff port map(x=>p(45)(73),y=>p(46)(73),Cin=>p(47)(73),clock=>clock,reset=>reset,s=>p(158)(73),cout=>p(159)(74));
FA_ff_1994:FAff port map(x=>p(45)(74),y=>p(46)(74),Cin=>p(47)(74),clock=>clock,reset=>reset,s=>p(158)(74),cout=>p(159)(75));
FA_ff_1995:FAff port map(x=>p(45)(75),y=>p(46)(75),Cin=>p(47)(75),clock=>clock,reset=>reset,s=>p(158)(75),cout=>p(159)(76));
FA_ff_1996:FAff port map(x=>p(45)(76),y=>p(46)(76),Cin=>p(47)(76),clock=>clock,reset=>reset,s=>p(158)(76),cout=>p(159)(77));
FA_ff_1997:FAff port map(x=>p(45)(77),y=>p(46)(77),Cin=>p(47)(77),clock=>clock,reset=>reset,s=>p(158)(77),cout=>p(159)(78));
FA_ff_1998:FAff port map(x=>p(45)(78),y=>p(46)(78),Cin=>p(47)(78),clock=>clock,reset=>reset,s=>p(158)(78),cout=>p(159)(79));
FA_ff_1999:FAff port map(x=>p(45)(79),y=>p(46)(79),Cin=>p(47)(79),clock=>clock,reset=>reset,s=>p(158)(79),cout=>p(159)(80));
FA_ff_2000:FAff port map(x=>p(45)(80),y=>p(46)(80),Cin=>p(47)(80),clock=>clock,reset=>reset,s=>p(158)(80),cout=>p(159)(81));
FA_ff_2001:FAff port map(x=>p(45)(81),y=>p(46)(81),Cin=>p(47)(81),clock=>clock,reset=>reset,s=>p(158)(81),cout=>p(159)(82));
FA_ff_2002:FAff port map(x=>p(45)(82),y=>p(46)(82),Cin=>p(47)(82),clock=>clock,reset=>reset,s=>p(158)(82),cout=>p(159)(83));
FA_ff_2003:FAff port map(x=>p(45)(83),y=>p(46)(83),Cin=>p(47)(83),clock=>clock,reset=>reset,s=>p(158)(83),cout=>p(159)(84));
FA_ff_2004:FAff port map(x=>p(45)(84),y=>p(46)(84),Cin=>p(47)(84),clock=>clock,reset=>reset,s=>p(158)(84),cout=>p(159)(85));
FA_ff_2005:FAff port map(x=>p(45)(85),y=>p(46)(85),Cin=>p(47)(85),clock=>clock,reset=>reset,s=>p(158)(85),cout=>p(159)(86));
FA_ff_2006:FAff port map(x=>p(45)(86),y=>p(46)(86),Cin=>p(47)(86),clock=>clock,reset=>reset,s=>p(158)(86),cout=>p(159)(87));
FA_ff_2007:FAff port map(x=>p(45)(87),y=>p(46)(87),Cin=>p(47)(87),clock=>clock,reset=>reset,s=>p(158)(87),cout=>p(159)(88));
FA_ff_2008:FAff port map(x=>p(45)(88),y=>p(46)(88),Cin=>p(47)(88),clock=>clock,reset=>reset,s=>p(158)(88),cout=>p(159)(89));
FA_ff_2009:FAff port map(x=>p(45)(89),y=>p(46)(89),Cin=>p(47)(89),clock=>clock,reset=>reset,s=>p(158)(89),cout=>p(159)(90));
FA_ff_2010:FAff port map(x=>p(45)(90),y=>p(46)(90),Cin=>p(47)(90),clock=>clock,reset=>reset,s=>p(158)(90),cout=>p(159)(91));
FA_ff_2011:FAff port map(x=>p(45)(91),y=>p(46)(91),Cin=>p(47)(91),clock=>clock,reset=>reset,s=>p(158)(91),cout=>p(159)(92));
FA_ff_2012:FAff port map(x=>p(45)(92),y=>p(46)(92),Cin=>p(47)(92),clock=>clock,reset=>reset,s=>p(158)(92),cout=>p(159)(93));
FA_ff_2013:FAff port map(x=>p(45)(93),y=>p(46)(93),Cin=>p(47)(93),clock=>clock,reset=>reset,s=>p(158)(93),cout=>p(159)(94));
FA_ff_2014:FAff port map(x=>p(45)(94),y=>p(46)(94),Cin=>p(47)(94),clock=>clock,reset=>reset,s=>p(158)(94),cout=>p(159)(95));
FA_ff_2015:FAff port map(x=>p(45)(95),y=>p(46)(95),Cin=>p(47)(95),clock=>clock,reset=>reset,s=>p(158)(95),cout=>p(159)(96));
FA_ff_2016:FAff port map(x=>p(45)(96),y=>p(46)(96),Cin=>p(47)(96),clock=>clock,reset=>reset,s=>p(158)(96),cout=>p(159)(97));
FA_ff_2017:FAff port map(x=>p(45)(97),y=>p(46)(97),Cin=>p(47)(97),clock=>clock,reset=>reset,s=>p(158)(97),cout=>p(159)(98));
FA_ff_2018:FAff port map(x=>p(45)(98),y=>p(46)(98),Cin=>p(47)(98),clock=>clock,reset=>reset,s=>p(158)(98),cout=>p(159)(99));
FA_ff_2019:FAff port map(x=>p(45)(99),y=>p(46)(99),Cin=>p(47)(99),clock=>clock,reset=>reset,s=>p(158)(99),cout=>p(159)(100));
FA_ff_2020:FAff port map(x=>p(45)(100),y=>p(46)(100),Cin=>p(47)(100),clock=>clock,reset=>reset,s=>p(158)(100),cout=>p(159)(101));
FA_ff_2021:FAff port map(x=>p(45)(101),y=>p(46)(101),Cin=>p(47)(101),clock=>clock,reset=>reset,s=>p(158)(101),cout=>p(159)(102));
FA_ff_2022:FAff port map(x=>p(45)(102),y=>p(46)(102),Cin=>p(47)(102),clock=>clock,reset=>reset,s=>p(158)(102),cout=>p(159)(103));
FA_ff_2023:FAff port map(x=>p(45)(103),y=>p(46)(103),Cin=>p(47)(103),clock=>clock,reset=>reset,s=>p(158)(103),cout=>p(159)(104));
FA_ff_2024:FAff port map(x=>p(45)(104),y=>p(46)(104),Cin=>p(47)(104),clock=>clock,reset=>reset,s=>p(158)(104),cout=>p(159)(105));
FA_ff_2025:FAff port map(x=>p(45)(105),y=>p(46)(105),Cin=>p(47)(105),clock=>clock,reset=>reset,s=>p(158)(105),cout=>p(159)(106));
FA_ff_2026:FAff port map(x=>p(45)(106),y=>p(46)(106),Cin=>p(47)(106),clock=>clock,reset=>reset,s=>p(158)(106),cout=>p(159)(107));
FA_ff_2027:FAff port map(x=>p(45)(107),y=>p(46)(107),Cin=>p(47)(107),clock=>clock,reset=>reset,s=>p(158)(107),cout=>p(159)(108));
FA_ff_2028:FAff port map(x=>p(45)(108),y=>p(46)(108),Cin=>p(47)(108),clock=>clock,reset=>reset,s=>p(158)(108),cout=>p(159)(109));
FA_ff_2029:FAff port map(x=>p(45)(109),y=>p(46)(109),Cin=>p(47)(109),clock=>clock,reset=>reset,s=>p(158)(109),cout=>p(159)(110));
FA_ff_2030:FAff port map(x=>p(45)(110),y=>p(46)(110),Cin=>p(47)(110),clock=>clock,reset=>reset,s=>p(158)(110),cout=>p(159)(111));
FA_ff_2031:FAff port map(x=>p(45)(111),y=>p(46)(111),Cin=>p(47)(111),clock=>clock,reset=>reset,s=>p(158)(111),cout=>p(159)(112));
FA_ff_2032:FAff port map(x=>p(45)(112),y=>p(46)(112),Cin=>p(47)(112),clock=>clock,reset=>reset,s=>p(158)(112),cout=>p(159)(113));
FA_ff_2033:FAff port map(x=>p(45)(113),y=>p(46)(113),Cin=>p(47)(113),clock=>clock,reset=>reset,s=>p(158)(113),cout=>p(159)(114));
FA_ff_2034:FAff port map(x=>p(45)(114),y=>p(46)(114),Cin=>p(47)(114),clock=>clock,reset=>reset,s=>p(158)(114),cout=>p(159)(115));
FA_ff_2035:FAff port map(x=>p(45)(115),y=>p(46)(115),Cin=>p(47)(115),clock=>clock,reset=>reset,s=>p(158)(115),cout=>p(159)(116));
FA_ff_2036:FAff port map(x=>p(45)(116),y=>p(46)(116),Cin=>p(47)(116),clock=>clock,reset=>reset,s=>p(158)(116),cout=>p(159)(117));
FA_ff_2037:FAff port map(x=>p(45)(117),y=>p(46)(117),Cin=>p(47)(117),clock=>clock,reset=>reset,s=>p(158)(117),cout=>p(159)(118));
FA_ff_2038:FAff port map(x=>p(45)(118),y=>p(46)(118),Cin=>p(47)(118),clock=>clock,reset=>reset,s=>p(158)(118),cout=>p(159)(119));
FA_ff_2039:FAff port map(x=>p(45)(119),y=>p(46)(119),Cin=>p(47)(119),clock=>clock,reset=>reset,s=>p(158)(119),cout=>p(159)(120));
FA_ff_2040:FAff port map(x=>p(45)(120),y=>p(46)(120),Cin=>p(47)(120),clock=>clock,reset=>reset,s=>p(158)(120),cout=>p(159)(121));
FA_ff_2041:FAff port map(x=>p(45)(121),y=>p(46)(121),Cin=>p(47)(121),clock=>clock,reset=>reset,s=>p(158)(121),cout=>p(159)(122));
FA_ff_2042:FAff port map(x=>p(45)(122),y=>p(46)(122),Cin=>p(47)(122),clock=>clock,reset=>reset,s=>p(158)(122),cout=>p(159)(123));
FA_ff_2043:FAff port map(x=>p(45)(123),y=>p(46)(123),Cin=>p(47)(123),clock=>clock,reset=>reset,s=>p(158)(123),cout=>p(159)(124));
FA_ff_2044:FAff port map(x=>p(45)(124),y=>p(46)(124),Cin=>p(47)(124),clock=>clock,reset=>reset,s=>p(158)(124),cout=>p(159)(125));
FA_ff_2045:FAff port map(x=>p(45)(125),y=>p(46)(125),Cin=>p(47)(125),clock=>clock,reset=>reset,s=>p(158)(125),cout=>p(159)(126));
FA_ff_2046:FAff port map(x=>p(45)(126),y=>p(46)(126),Cin=>p(47)(126),clock=>clock,reset=>reset,s=>p(158)(126),cout=>p(159)(127));
FA_ff_2047:FAff port map(x=>p(45)(127),y=>p(46)(127),Cin=>p(47)(127),clock=>clock,reset=>reset,s=>p(158)(127),cout=>p(159)(128));
FA_ff_2048:FAff port map(x=>p(48)(0),y=>p(49)(0),Cin=>p(50)(0),clock=>clock,reset=>reset,s=>p(160)(0),cout=>p(161)(1));
FA_ff_2049:FAff port map(x=>p(48)(1),y=>p(49)(1),Cin=>p(50)(1),clock=>clock,reset=>reset,s=>p(160)(1),cout=>p(161)(2));
FA_ff_2050:FAff port map(x=>p(48)(2),y=>p(49)(2),Cin=>p(50)(2),clock=>clock,reset=>reset,s=>p(160)(2),cout=>p(161)(3));
FA_ff_2051:FAff port map(x=>p(48)(3),y=>p(49)(3),Cin=>p(50)(3),clock=>clock,reset=>reset,s=>p(160)(3),cout=>p(161)(4));
FA_ff_2052:FAff port map(x=>p(48)(4),y=>p(49)(4),Cin=>p(50)(4),clock=>clock,reset=>reset,s=>p(160)(4),cout=>p(161)(5));
FA_ff_2053:FAff port map(x=>p(48)(5),y=>p(49)(5),Cin=>p(50)(5),clock=>clock,reset=>reset,s=>p(160)(5),cout=>p(161)(6));
FA_ff_2054:FAff port map(x=>p(48)(6),y=>p(49)(6),Cin=>p(50)(6),clock=>clock,reset=>reset,s=>p(160)(6),cout=>p(161)(7));
FA_ff_2055:FAff port map(x=>p(48)(7),y=>p(49)(7),Cin=>p(50)(7),clock=>clock,reset=>reset,s=>p(160)(7),cout=>p(161)(8));
FA_ff_2056:FAff port map(x=>p(48)(8),y=>p(49)(8),Cin=>p(50)(8),clock=>clock,reset=>reset,s=>p(160)(8),cout=>p(161)(9));
FA_ff_2057:FAff port map(x=>p(48)(9),y=>p(49)(9),Cin=>p(50)(9),clock=>clock,reset=>reset,s=>p(160)(9),cout=>p(161)(10));
FA_ff_2058:FAff port map(x=>p(48)(10),y=>p(49)(10),Cin=>p(50)(10),clock=>clock,reset=>reset,s=>p(160)(10),cout=>p(161)(11));
FA_ff_2059:FAff port map(x=>p(48)(11),y=>p(49)(11),Cin=>p(50)(11),clock=>clock,reset=>reset,s=>p(160)(11),cout=>p(161)(12));
FA_ff_2060:FAff port map(x=>p(48)(12),y=>p(49)(12),Cin=>p(50)(12),clock=>clock,reset=>reset,s=>p(160)(12),cout=>p(161)(13));
FA_ff_2061:FAff port map(x=>p(48)(13),y=>p(49)(13),Cin=>p(50)(13),clock=>clock,reset=>reset,s=>p(160)(13),cout=>p(161)(14));
FA_ff_2062:FAff port map(x=>p(48)(14),y=>p(49)(14),Cin=>p(50)(14),clock=>clock,reset=>reset,s=>p(160)(14),cout=>p(161)(15));
FA_ff_2063:FAff port map(x=>p(48)(15),y=>p(49)(15),Cin=>p(50)(15),clock=>clock,reset=>reset,s=>p(160)(15),cout=>p(161)(16));
FA_ff_2064:FAff port map(x=>p(48)(16),y=>p(49)(16),Cin=>p(50)(16),clock=>clock,reset=>reset,s=>p(160)(16),cout=>p(161)(17));
FA_ff_2065:FAff port map(x=>p(48)(17),y=>p(49)(17),Cin=>p(50)(17),clock=>clock,reset=>reset,s=>p(160)(17),cout=>p(161)(18));
FA_ff_2066:FAff port map(x=>p(48)(18),y=>p(49)(18),Cin=>p(50)(18),clock=>clock,reset=>reset,s=>p(160)(18),cout=>p(161)(19));
FA_ff_2067:FAff port map(x=>p(48)(19),y=>p(49)(19),Cin=>p(50)(19),clock=>clock,reset=>reset,s=>p(160)(19),cout=>p(161)(20));
FA_ff_2068:FAff port map(x=>p(48)(20),y=>p(49)(20),Cin=>p(50)(20),clock=>clock,reset=>reset,s=>p(160)(20),cout=>p(161)(21));
FA_ff_2069:FAff port map(x=>p(48)(21),y=>p(49)(21),Cin=>p(50)(21),clock=>clock,reset=>reset,s=>p(160)(21),cout=>p(161)(22));
FA_ff_2070:FAff port map(x=>p(48)(22),y=>p(49)(22),Cin=>p(50)(22),clock=>clock,reset=>reset,s=>p(160)(22),cout=>p(161)(23));
FA_ff_2071:FAff port map(x=>p(48)(23),y=>p(49)(23),Cin=>p(50)(23),clock=>clock,reset=>reset,s=>p(160)(23),cout=>p(161)(24));
FA_ff_2072:FAff port map(x=>p(48)(24),y=>p(49)(24),Cin=>p(50)(24),clock=>clock,reset=>reset,s=>p(160)(24),cout=>p(161)(25));
FA_ff_2073:FAff port map(x=>p(48)(25),y=>p(49)(25),Cin=>p(50)(25),clock=>clock,reset=>reset,s=>p(160)(25),cout=>p(161)(26));
FA_ff_2074:FAff port map(x=>p(48)(26),y=>p(49)(26),Cin=>p(50)(26),clock=>clock,reset=>reset,s=>p(160)(26),cout=>p(161)(27));
FA_ff_2075:FAff port map(x=>p(48)(27),y=>p(49)(27),Cin=>p(50)(27),clock=>clock,reset=>reset,s=>p(160)(27),cout=>p(161)(28));
FA_ff_2076:FAff port map(x=>p(48)(28),y=>p(49)(28),Cin=>p(50)(28),clock=>clock,reset=>reset,s=>p(160)(28),cout=>p(161)(29));
FA_ff_2077:FAff port map(x=>p(48)(29),y=>p(49)(29),Cin=>p(50)(29),clock=>clock,reset=>reset,s=>p(160)(29),cout=>p(161)(30));
FA_ff_2078:FAff port map(x=>p(48)(30),y=>p(49)(30),Cin=>p(50)(30),clock=>clock,reset=>reset,s=>p(160)(30),cout=>p(161)(31));
FA_ff_2079:FAff port map(x=>p(48)(31),y=>p(49)(31),Cin=>p(50)(31),clock=>clock,reset=>reset,s=>p(160)(31),cout=>p(161)(32));
FA_ff_2080:FAff port map(x=>p(48)(32),y=>p(49)(32),Cin=>p(50)(32),clock=>clock,reset=>reset,s=>p(160)(32),cout=>p(161)(33));
FA_ff_2081:FAff port map(x=>p(48)(33),y=>p(49)(33),Cin=>p(50)(33),clock=>clock,reset=>reset,s=>p(160)(33),cout=>p(161)(34));
FA_ff_2082:FAff port map(x=>p(48)(34),y=>p(49)(34),Cin=>p(50)(34),clock=>clock,reset=>reset,s=>p(160)(34),cout=>p(161)(35));
FA_ff_2083:FAff port map(x=>p(48)(35),y=>p(49)(35),Cin=>p(50)(35),clock=>clock,reset=>reset,s=>p(160)(35),cout=>p(161)(36));
FA_ff_2084:FAff port map(x=>p(48)(36),y=>p(49)(36),Cin=>p(50)(36),clock=>clock,reset=>reset,s=>p(160)(36),cout=>p(161)(37));
FA_ff_2085:FAff port map(x=>p(48)(37),y=>p(49)(37),Cin=>p(50)(37),clock=>clock,reset=>reset,s=>p(160)(37),cout=>p(161)(38));
FA_ff_2086:FAff port map(x=>p(48)(38),y=>p(49)(38),Cin=>p(50)(38),clock=>clock,reset=>reset,s=>p(160)(38),cout=>p(161)(39));
FA_ff_2087:FAff port map(x=>p(48)(39),y=>p(49)(39),Cin=>p(50)(39),clock=>clock,reset=>reset,s=>p(160)(39),cout=>p(161)(40));
FA_ff_2088:FAff port map(x=>p(48)(40),y=>p(49)(40),Cin=>p(50)(40),clock=>clock,reset=>reset,s=>p(160)(40),cout=>p(161)(41));
FA_ff_2089:FAff port map(x=>p(48)(41),y=>p(49)(41),Cin=>p(50)(41),clock=>clock,reset=>reset,s=>p(160)(41),cout=>p(161)(42));
FA_ff_2090:FAff port map(x=>p(48)(42),y=>p(49)(42),Cin=>p(50)(42),clock=>clock,reset=>reset,s=>p(160)(42),cout=>p(161)(43));
FA_ff_2091:FAff port map(x=>p(48)(43),y=>p(49)(43),Cin=>p(50)(43),clock=>clock,reset=>reset,s=>p(160)(43),cout=>p(161)(44));
FA_ff_2092:FAff port map(x=>p(48)(44),y=>p(49)(44),Cin=>p(50)(44),clock=>clock,reset=>reset,s=>p(160)(44),cout=>p(161)(45));
FA_ff_2093:FAff port map(x=>p(48)(45),y=>p(49)(45),Cin=>p(50)(45),clock=>clock,reset=>reset,s=>p(160)(45),cout=>p(161)(46));
FA_ff_2094:FAff port map(x=>p(48)(46),y=>p(49)(46),Cin=>p(50)(46),clock=>clock,reset=>reset,s=>p(160)(46),cout=>p(161)(47));
FA_ff_2095:FAff port map(x=>p(48)(47),y=>p(49)(47),Cin=>p(50)(47),clock=>clock,reset=>reset,s=>p(160)(47),cout=>p(161)(48));
FA_ff_2096:FAff port map(x=>p(48)(48),y=>p(49)(48),Cin=>p(50)(48),clock=>clock,reset=>reset,s=>p(160)(48),cout=>p(161)(49));
FA_ff_2097:FAff port map(x=>p(48)(49),y=>p(49)(49),Cin=>p(50)(49),clock=>clock,reset=>reset,s=>p(160)(49),cout=>p(161)(50));
FA_ff_2098:FAff port map(x=>p(48)(50),y=>p(49)(50),Cin=>p(50)(50),clock=>clock,reset=>reset,s=>p(160)(50),cout=>p(161)(51));
FA_ff_2099:FAff port map(x=>p(48)(51),y=>p(49)(51),Cin=>p(50)(51),clock=>clock,reset=>reset,s=>p(160)(51),cout=>p(161)(52));
FA_ff_2100:FAff port map(x=>p(48)(52),y=>p(49)(52),Cin=>p(50)(52),clock=>clock,reset=>reset,s=>p(160)(52),cout=>p(161)(53));
FA_ff_2101:FAff port map(x=>p(48)(53),y=>p(49)(53),Cin=>p(50)(53),clock=>clock,reset=>reset,s=>p(160)(53),cout=>p(161)(54));
FA_ff_2102:FAff port map(x=>p(48)(54),y=>p(49)(54),Cin=>p(50)(54),clock=>clock,reset=>reset,s=>p(160)(54),cout=>p(161)(55));
FA_ff_2103:FAff port map(x=>p(48)(55),y=>p(49)(55),Cin=>p(50)(55),clock=>clock,reset=>reset,s=>p(160)(55),cout=>p(161)(56));
FA_ff_2104:FAff port map(x=>p(48)(56),y=>p(49)(56),Cin=>p(50)(56),clock=>clock,reset=>reset,s=>p(160)(56),cout=>p(161)(57));
FA_ff_2105:FAff port map(x=>p(48)(57),y=>p(49)(57),Cin=>p(50)(57),clock=>clock,reset=>reset,s=>p(160)(57),cout=>p(161)(58));
FA_ff_2106:FAff port map(x=>p(48)(58),y=>p(49)(58),Cin=>p(50)(58),clock=>clock,reset=>reset,s=>p(160)(58),cout=>p(161)(59));
FA_ff_2107:FAff port map(x=>p(48)(59),y=>p(49)(59),Cin=>p(50)(59),clock=>clock,reset=>reset,s=>p(160)(59),cout=>p(161)(60));
FA_ff_2108:FAff port map(x=>p(48)(60),y=>p(49)(60),Cin=>p(50)(60),clock=>clock,reset=>reset,s=>p(160)(60),cout=>p(161)(61));
FA_ff_2109:FAff port map(x=>p(48)(61),y=>p(49)(61),Cin=>p(50)(61),clock=>clock,reset=>reset,s=>p(160)(61),cout=>p(161)(62));
FA_ff_2110:FAff port map(x=>p(48)(62),y=>p(49)(62),Cin=>p(50)(62),clock=>clock,reset=>reset,s=>p(160)(62),cout=>p(161)(63));
FA_ff_2111:FAff port map(x=>p(48)(63),y=>p(49)(63),Cin=>p(50)(63),clock=>clock,reset=>reset,s=>p(160)(63),cout=>p(161)(64));
FA_ff_2112:FAff port map(x=>p(48)(64),y=>p(49)(64),Cin=>p(50)(64),clock=>clock,reset=>reset,s=>p(160)(64),cout=>p(161)(65));
FA_ff_2113:FAff port map(x=>p(48)(65),y=>p(49)(65),Cin=>p(50)(65),clock=>clock,reset=>reset,s=>p(160)(65),cout=>p(161)(66));
FA_ff_2114:FAff port map(x=>p(48)(66),y=>p(49)(66),Cin=>p(50)(66),clock=>clock,reset=>reset,s=>p(160)(66),cout=>p(161)(67));
FA_ff_2115:FAff port map(x=>p(48)(67),y=>p(49)(67),Cin=>p(50)(67),clock=>clock,reset=>reset,s=>p(160)(67),cout=>p(161)(68));
FA_ff_2116:FAff port map(x=>p(48)(68),y=>p(49)(68),Cin=>p(50)(68),clock=>clock,reset=>reset,s=>p(160)(68),cout=>p(161)(69));
FA_ff_2117:FAff port map(x=>p(48)(69),y=>p(49)(69),Cin=>p(50)(69),clock=>clock,reset=>reset,s=>p(160)(69),cout=>p(161)(70));
FA_ff_2118:FAff port map(x=>p(48)(70),y=>p(49)(70),Cin=>p(50)(70),clock=>clock,reset=>reset,s=>p(160)(70),cout=>p(161)(71));
FA_ff_2119:FAff port map(x=>p(48)(71),y=>p(49)(71),Cin=>p(50)(71),clock=>clock,reset=>reset,s=>p(160)(71),cout=>p(161)(72));
FA_ff_2120:FAff port map(x=>p(48)(72),y=>p(49)(72),Cin=>p(50)(72),clock=>clock,reset=>reset,s=>p(160)(72),cout=>p(161)(73));
FA_ff_2121:FAff port map(x=>p(48)(73),y=>p(49)(73),Cin=>p(50)(73),clock=>clock,reset=>reset,s=>p(160)(73),cout=>p(161)(74));
FA_ff_2122:FAff port map(x=>p(48)(74),y=>p(49)(74),Cin=>p(50)(74),clock=>clock,reset=>reset,s=>p(160)(74),cout=>p(161)(75));
FA_ff_2123:FAff port map(x=>p(48)(75),y=>p(49)(75),Cin=>p(50)(75),clock=>clock,reset=>reset,s=>p(160)(75),cout=>p(161)(76));
FA_ff_2124:FAff port map(x=>p(48)(76),y=>p(49)(76),Cin=>p(50)(76),clock=>clock,reset=>reset,s=>p(160)(76),cout=>p(161)(77));
FA_ff_2125:FAff port map(x=>p(48)(77),y=>p(49)(77),Cin=>p(50)(77),clock=>clock,reset=>reset,s=>p(160)(77),cout=>p(161)(78));
FA_ff_2126:FAff port map(x=>p(48)(78),y=>p(49)(78),Cin=>p(50)(78),clock=>clock,reset=>reset,s=>p(160)(78),cout=>p(161)(79));
FA_ff_2127:FAff port map(x=>p(48)(79),y=>p(49)(79),Cin=>p(50)(79),clock=>clock,reset=>reset,s=>p(160)(79),cout=>p(161)(80));
FA_ff_2128:FAff port map(x=>p(48)(80),y=>p(49)(80),Cin=>p(50)(80),clock=>clock,reset=>reset,s=>p(160)(80),cout=>p(161)(81));
FA_ff_2129:FAff port map(x=>p(48)(81),y=>p(49)(81),Cin=>p(50)(81),clock=>clock,reset=>reset,s=>p(160)(81),cout=>p(161)(82));
FA_ff_2130:FAff port map(x=>p(48)(82),y=>p(49)(82),Cin=>p(50)(82),clock=>clock,reset=>reset,s=>p(160)(82),cout=>p(161)(83));
FA_ff_2131:FAff port map(x=>p(48)(83),y=>p(49)(83),Cin=>p(50)(83),clock=>clock,reset=>reset,s=>p(160)(83),cout=>p(161)(84));
FA_ff_2132:FAff port map(x=>p(48)(84),y=>p(49)(84),Cin=>p(50)(84),clock=>clock,reset=>reset,s=>p(160)(84),cout=>p(161)(85));
FA_ff_2133:FAff port map(x=>p(48)(85),y=>p(49)(85),Cin=>p(50)(85),clock=>clock,reset=>reset,s=>p(160)(85),cout=>p(161)(86));
FA_ff_2134:FAff port map(x=>p(48)(86),y=>p(49)(86),Cin=>p(50)(86),clock=>clock,reset=>reset,s=>p(160)(86),cout=>p(161)(87));
FA_ff_2135:FAff port map(x=>p(48)(87),y=>p(49)(87),Cin=>p(50)(87),clock=>clock,reset=>reset,s=>p(160)(87),cout=>p(161)(88));
FA_ff_2136:FAff port map(x=>p(48)(88),y=>p(49)(88),Cin=>p(50)(88),clock=>clock,reset=>reset,s=>p(160)(88),cout=>p(161)(89));
FA_ff_2137:FAff port map(x=>p(48)(89),y=>p(49)(89),Cin=>p(50)(89),clock=>clock,reset=>reset,s=>p(160)(89),cout=>p(161)(90));
FA_ff_2138:FAff port map(x=>p(48)(90),y=>p(49)(90),Cin=>p(50)(90),clock=>clock,reset=>reset,s=>p(160)(90),cout=>p(161)(91));
FA_ff_2139:FAff port map(x=>p(48)(91),y=>p(49)(91),Cin=>p(50)(91),clock=>clock,reset=>reset,s=>p(160)(91),cout=>p(161)(92));
FA_ff_2140:FAff port map(x=>p(48)(92),y=>p(49)(92),Cin=>p(50)(92),clock=>clock,reset=>reset,s=>p(160)(92),cout=>p(161)(93));
FA_ff_2141:FAff port map(x=>p(48)(93),y=>p(49)(93),Cin=>p(50)(93),clock=>clock,reset=>reset,s=>p(160)(93),cout=>p(161)(94));
FA_ff_2142:FAff port map(x=>p(48)(94),y=>p(49)(94),Cin=>p(50)(94),clock=>clock,reset=>reset,s=>p(160)(94),cout=>p(161)(95));
FA_ff_2143:FAff port map(x=>p(48)(95),y=>p(49)(95),Cin=>p(50)(95),clock=>clock,reset=>reset,s=>p(160)(95),cout=>p(161)(96));
FA_ff_2144:FAff port map(x=>p(48)(96),y=>p(49)(96),Cin=>p(50)(96),clock=>clock,reset=>reset,s=>p(160)(96),cout=>p(161)(97));
FA_ff_2145:FAff port map(x=>p(48)(97),y=>p(49)(97),Cin=>p(50)(97),clock=>clock,reset=>reset,s=>p(160)(97),cout=>p(161)(98));
FA_ff_2146:FAff port map(x=>p(48)(98),y=>p(49)(98),Cin=>p(50)(98),clock=>clock,reset=>reset,s=>p(160)(98),cout=>p(161)(99));
FA_ff_2147:FAff port map(x=>p(48)(99),y=>p(49)(99),Cin=>p(50)(99),clock=>clock,reset=>reset,s=>p(160)(99),cout=>p(161)(100));
FA_ff_2148:FAff port map(x=>p(48)(100),y=>p(49)(100),Cin=>p(50)(100),clock=>clock,reset=>reset,s=>p(160)(100),cout=>p(161)(101));
FA_ff_2149:FAff port map(x=>p(48)(101),y=>p(49)(101),Cin=>p(50)(101),clock=>clock,reset=>reset,s=>p(160)(101),cout=>p(161)(102));
FA_ff_2150:FAff port map(x=>p(48)(102),y=>p(49)(102),Cin=>p(50)(102),clock=>clock,reset=>reset,s=>p(160)(102),cout=>p(161)(103));
FA_ff_2151:FAff port map(x=>p(48)(103),y=>p(49)(103),Cin=>p(50)(103),clock=>clock,reset=>reset,s=>p(160)(103),cout=>p(161)(104));
FA_ff_2152:FAff port map(x=>p(48)(104),y=>p(49)(104),Cin=>p(50)(104),clock=>clock,reset=>reset,s=>p(160)(104),cout=>p(161)(105));
FA_ff_2153:FAff port map(x=>p(48)(105),y=>p(49)(105),Cin=>p(50)(105),clock=>clock,reset=>reset,s=>p(160)(105),cout=>p(161)(106));
FA_ff_2154:FAff port map(x=>p(48)(106),y=>p(49)(106),Cin=>p(50)(106),clock=>clock,reset=>reset,s=>p(160)(106),cout=>p(161)(107));
FA_ff_2155:FAff port map(x=>p(48)(107),y=>p(49)(107),Cin=>p(50)(107),clock=>clock,reset=>reset,s=>p(160)(107),cout=>p(161)(108));
FA_ff_2156:FAff port map(x=>p(48)(108),y=>p(49)(108),Cin=>p(50)(108),clock=>clock,reset=>reset,s=>p(160)(108),cout=>p(161)(109));
FA_ff_2157:FAff port map(x=>p(48)(109),y=>p(49)(109),Cin=>p(50)(109),clock=>clock,reset=>reset,s=>p(160)(109),cout=>p(161)(110));
FA_ff_2158:FAff port map(x=>p(48)(110),y=>p(49)(110),Cin=>p(50)(110),clock=>clock,reset=>reset,s=>p(160)(110),cout=>p(161)(111));
FA_ff_2159:FAff port map(x=>p(48)(111),y=>p(49)(111),Cin=>p(50)(111),clock=>clock,reset=>reset,s=>p(160)(111),cout=>p(161)(112));
FA_ff_2160:FAff port map(x=>p(48)(112),y=>p(49)(112),Cin=>p(50)(112),clock=>clock,reset=>reset,s=>p(160)(112),cout=>p(161)(113));
FA_ff_2161:FAff port map(x=>p(48)(113),y=>p(49)(113),Cin=>p(50)(113),clock=>clock,reset=>reset,s=>p(160)(113),cout=>p(161)(114));
FA_ff_2162:FAff port map(x=>p(48)(114),y=>p(49)(114),Cin=>p(50)(114),clock=>clock,reset=>reset,s=>p(160)(114),cout=>p(161)(115));
FA_ff_2163:FAff port map(x=>p(48)(115),y=>p(49)(115),Cin=>p(50)(115),clock=>clock,reset=>reset,s=>p(160)(115),cout=>p(161)(116));
FA_ff_2164:FAff port map(x=>p(48)(116),y=>p(49)(116),Cin=>p(50)(116),clock=>clock,reset=>reset,s=>p(160)(116),cout=>p(161)(117));
FA_ff_2165:FAff port map(x=>p(48)(117),y=>p(49)(117),Cin=>p(50)(117),clock=>clock,reset=>reset,s=>p(160)(117),cout=>p(161)(118));
FA_ff_2166:FAff port map(x=>p(48)(118),y=>p(49)(118),Cin=>p(50)(118),clock=>clock,reset=>reset,s=>p(160)(118),cout=>p(161)(119));
FA_ff_2167:FAff port map(x=>p(48)(119),y=>p(49)(119),Cin=>p(50)(119),clock=>clock,reset=>reset,s=>p(160)(119),cout=>p(161)(120));
FA_ff_2168:FAff port map(x=>p(48)(120),y=>p(49)(120),Cin=>p(50)(120),clock=>clock,reset=>reset,s=>p(160)(120),cout=>p(161)(121));
FA_ff_2169:FAff port map(x=>p(48)(121),y=>p(49)(121),Cin=>p(50)(121),clock=>clock,reset=>reset,s=>p(160)(121),cout=>p(161)(122));
FA_ff_2170:FAff port map(x=>p(48)(122),y=>p(49)(122),Cin=>p(50)(122),clock=>clock,reset=>reset,s=>p(160)(122),cout=>p(161)(123));
FA_ff_2171:FAff port map(x=>p(48)(123),y=>p(49)(123),Cin=>p(50)(123),clock=>clock,reset=>reset,s=>p(160)(123),cout=>p(161)(124));
FA_ff_2172:FAff port map(x=>p(48)(124),y=>p(49)(124),Cin=>p(50)(124),clock=>clock,reset=>reset,s=>p(160)(124),cout=>p(161)(125));
FA_ff_2173:FAff port map(x=>p(48)(125),y=>p(49)(125),Cin=>p(50)(125),clock=>clock,reset=>reset,s=>p(160)(125),cout=>p(161)(126));
FA_ff_2174:FAff port map(x=>p(48)(126),y=>p(49)(126),Cin=>p(50)(126),clock=>clock,reset=>reset,s=>p(160)(126),cout=>p(161)(127));
FA_ff_2175:FAff port map(x=>p(48)(127),y=>p(49)(127),Cin=>p(50)(127),clock=>clock,reset=>reset,s=>p(160)(127),cout=>p(161)(128));
FA_ff_2176:FAff port map(x=>p(51)(0),y=>p(52)(0),Cin=>p(53)(0),clock=>clock,reset=>reset,s=>p(162)(0),cout=>p(163)(1));
FA_ff_2177:FAff port map(x=>p(51)(1),y=>p(52)(1),Cin=>p(53)(1),clock=>clock,reset=>reset,s=>p(162)(1),cout=>p(163)(2));
FA_ff_2178:FAff port map(x=>p(51)(2),y=>p(52)(2),Cin=>p(53)(2),clock=>clock,reset=>reset,s=>p(162)(2),cout=>p(163)(3));
FA_ff_2179:FAff port map(x=>p(51)(3),y=>p(52)(3),Cin=>p(53)(3),clock=>clock,reset=>reset,s=>p(162)(3),cout=>p(163)(4));
FA_ff_2180:FAff port map(x=>p(51)(4),y=>p(52)(4),Cin=>p(53)(4),clock=>clock,reset=>reset,s=>p(162)(4),cout=>p(163)(5));
FA_ff_2181:FAff port map(x=>p(51)(5),y=>p(52)(5),Cin=>p(53)(5),clock=>clock,reset=>reset,s=>p(162)(5),cout=>p(163)(6));
FA_ff_2182:FAff port map(x=>p(51)(6),y=>p(52)(6),Cin=>p(53)(6),clock=>clock,reset=>reset,s=>p(162)(6),cout=>p(163)(7));
FA_ff_2183:FAff port map(x=>p(51)(7),y=>p(52)(7),Cin=>p(53)(7),clock=>clock,reset=>reset,s=>p(162)(7),cout=>p(163)(8));
FA_ff_2184:FAff port map(x=>p(51)(8),y=>p(52)(8),Cin=>p(53)(8),clock=>clock,reset=>reset,s=>p(162)(8),cout=>p(163)(9));
FA_ff_2185:FAff port map(x=>p(51)(9),y=>p(52)(9),Cin=>p(53)(9),clock=>clock,reset=>reset,s=>p(162)(9),cout=>p(163)(10));
FA_ff_2186:FAff port map(x=>p(51)(10),y=>p(52)(10),Cin=>p(53)(10),clock=>clock,reset=>reset,s=>p(162)(10),cout=>p(163)(11));
FA_ff_2187:FAff port map(x=>p(51)(11),y=>p(52)(11),Cin=>p(53)(11),clock=>clock,reset=>reset,s=>p(162)(11),cout=>p(163)(12));
FA_ff_2188:FAff port map(x=>p(51)(12),y=>p(52)(12),Cin=>p(53)(12),clock=>clock,reset=>reset,s=>p(162)(12),cout=>p(163)(13));
FA_ff_2189:FAff port map(x=>p(51)(13),y=>p(52)(13),Cin=>p(53)(13),clock=>clock,reset=>reset,s=>p(162)(13),cout=>p(163)(14));
FA_ff_2190:FAff port map(x=>p(51)(14),y=>p(52)(14),Cin=>p(53)(14),clock=>clock,reset=>reset,s=>p(162)(14),cout=>p(163)(15));
FA_ff_2191:FAff port map(x=>p(51)(15),y=>p(52)(15),Cin=>p(53)(15),clock=>clock,reset=>reset,s=>p(162)(15),cout=>p(163)(16));
FA_ff_2192:FAff port map(x=>p(51)(16),y=>p(52)(16),Cin=>p(53)(16),clock=>clock,reset=>reset,s=>p(162)(16),cout=>p(163)(17));
FA_ff_2193:FAff port map(x=>p(51)(17),y=>p(52)(17),Cin=>p(53)(17),clock=>clock,reset=>reset,s=>p(162)(17),cout=>p(163)(18));
FA_ff_2194:FAff port map(x=>p(51)(18),y=>p(52)(18),Cin=>p(53)(18),clock=>clock,reset=>reset,s=>p(162)(18),cout=>p(163)(19));
FA_ff_2195:FAff port map(x=>p(51)(19),y=>p(52)(19),Cin=>p(53)(19),clock=>clock,reset=>reset,s=>p(162)(19),cout=>p(163)(20));
FA_ff_2196:FAff port map(x=>p(51)(20),y=>p(52)(20),Cin=>p(53)(20),clock=>clock,reset=>reset,s=>p(162)(20),cout=>p(163)(21));
FA_ff_2197:FAff port map(x=>p(51)(21),y=>p(52)(21),Cin=>p(53)(21),clock=>clock,reset=>reset,s=>p(162)(21),cout=>p(163)(22));
FA_ff_2198:FAff port map(x=>p(51)(22),y=>p(52)(22),Cin=>p(53)(22),clock=>clock,reset=>reset,s=>p(162)(22),cout=>p(163)(23));
FA_ff_2199:FAff port map(x=>p(51)(23),y=>p(52)(23),Cin=>p(53)(23),clock=>clock,reset=>reset,s=>p(162)(23),cout=>p(163)(24));
FA_ff_2200:FAff port map(x=>p(51)(24),y=>p(52)(24),Cin=>p(53)(24),clock=>clock,reset=>reset,s=>p(162)(24),cout=>p(163)(25));
FA_ff_2201:FAff port map(x=>p(51)(25),y=>p(52)(25),Cin=>p(53)(25),clock=>clock,reset=>reset,s=>p(162)(25),cout=>p(163)(26));
FA_ff_2202:FAff port map(x=>p(51)(26),y=>p(52)(26),Cin=>p(53)(26),clock=>clock,reset=>reset,s=>p(162)(26),cout=>p(163)(27));
FA_ff_2203:FAff port map(x=>p(51)(27),y=>p(52)(27),Cin=>p(53)(27),clock=>clock,reset=>reset,s=>p(162)(27),cout=>p(163)(28));
FA_ff_2204:FAff port map(x=>p(51)(28),y=>p(52)(28),Cin=>p(53)(28),clock=>clock,reset=>reset,s=>p(162)(28),cout=>p(163)(29));
FA_ff_2205:FAff port map(x=>p(51)(29),y=>p(52)(29),Cin=>p(53)(29),clock=>clock,reset=>reset,s=>p(162)(29),cout=>p(163)(30));
FA_ff_2206:FAff port map(x=>p(51)(30),y=>p(52)(30),Cin=>p(53)(30),clock=>clock,reset=>reset,s=>p(162)(30),cout=>p(163)(31));
FA_ff_2207:FAff port map(x=>p(51)(31),y=>p(52)(31),Cin=>p(53)(31),clock=>clock,reset=>reset,s=>p(162)(31),cout=>p(163)(32));
FA_ff_2208:FAff port map(x=>p(51)(32),y=>p(52)(32),Cin=>p(53)(32),clock=>clock,reset=>reset,s=>p(162)(32),cout=>p(163)(33));
FA_ff_2209:FAff port map(x=>p(51)(33),y=>p(52)(33),Cin=>p(53)(33),clock=>clock,reset=>reset,s=>p(162)(33),cout=>p(163)(34));
FA_ff_2210:FAff port map(x=>p(51)(34),y=>p(52)(34),Cin=>p(53)(34),clock=>clock,reset=>reset,s=>p(162)(34),cout=>p(163)(35));
FA_ff_2211:FAff port map(x=>p(51)(35),y=>p(52)(35),Cin=>p(53)(35),clock=>clock,reset=>reset,s=>p(162)(35),cout=>p(163)(36));
FA_ff_2212:FAff port map(x=>p(51)(36),y=>p(52)(36),Cin=>p(53)(36),clock=>clock,reset=>reset,s=>p(162)(36),cout=>p(163)(37));
FA_ff_2213:FAff port map(x=>p(51)(37),y=>p(52)(37),Cin=>p(53)(37),clock=>clock,reset=>reset,s=>p(162)(37),cout=>p(163)(38));
FA_ff_2214:FAff port map(x=>p(51)(38),y=>p(52)(38),Cin=>p(53)(38),clock=>clock,reset=>reset,s=>p(162)(38),cout=>p(163)(39));
FA_ff_2215:FAff port map(x=>p(51)(39),y=>p(52)(39),Cin=>p(53)(39),clock=>clock,reset=>reset,s=>p(162)(39),cout=>p(163)(40));
FA_ff_2216:FAff port map(x=>p(51)(40),y=>p(52)(40),Cin=>p(53)(40),clock=>clock,reset=>reset,s=>p(162)(40),cout=>p(163)(41));
FA_ff_2217:FAff port map(x=>p(51)(41),y=>p(52)(41),Cin=>p(53)(41),clock=>clock,reset=>reset,s=>p(162)(41),cout=>p(163)(42));
FA_ff_2218:FAff port map(x=>p(51)(42),y=>p(52)(42),Cin=>p(53)(42),clock=>clock,reset=>reset,s=>p(162)(42),cout=>p(163)(43));
FA_ff_2219:FAff port map(x=>p(51)(43),y=>p(52)(43),Cin=>p(53)(43),clock=>clock,reset=>reset,s=>p(162)(43),cout=>p(163)(44));
FA_ff_2220:FAff port map(x=>p(51)(44),y=>p(52)(44),Cin=>p(53)(44),clock=>clock,reset=>reset,s=>p(162)(44),cout=>p(163)(45));
FA_ff_2221:FAff port map(x=>p(51)(45),y=>p(52)(45),Cin=>p(53)(45),clock=>clock,reset=>reset,s=>p(162)(45),cout=>p(163)(46));
FA_ff_2222:FAff port map(x=>p(51)(46),y=>p(52)(46),Cin=>p(53)(46),clock=>clock,reset=>reset,s=>p(162)(46),cout=>p(163)(47));
FA_ff_2223:FAff port map(x=>p(51)(47),y=>p(52)(47),Cin=>p(53)(47),clock=>clock,reset=>reset,s=>p(162)(47),cout=>p(163)(48));
FA_ff_2224:FAff port map(x=>p(51)(48),y=>p(52)(48),Cin=>p(53)(48),clock=>clock,reset=>reset,s=>p(162)(48),cout=>p(163)(49));
FA_ff_2225:FAff port map(x=>p(51)(49),y=>p(52)(49),Cin=>p(53)(49),clock=>clock,reset=>reset,s=>p(162)(49),cout=>p(163)(50));
FA_ff_2226:FAff port map(x=>p(51)(50),y=>p(52)(50),Cin=>p(53)(50),clock=>clock,reset=>reset,s=>p(162)(50),cout=>p(163)(51));
FA_ff_2227:FAff port map(x=>p(51)(51),y=>p(52)(51),Cin=>p(53)(51),clock=>clock,reset=>reset,s=>p(162)(51),cout=>p(163)(52));
FA_ff_2228:FAff port map(x=>p(51)(52),y=>p(52)(52),Cin=>p(53)(52),clock=>clock,reset=>reset,s=>p(162)(52),cout=>p(163)(53));
FA_ff_2229:FAff port map(x=>p(51)(53),y=>p(52)(53),Cin=>p(53)(53),clock=>clock,reset=>reset,s=>p(162)(53),cout=>p(163)(54));
FA_ff_2230:FAff port map(x=>p(51)(54),y=>p(52)(54),Cin=>p(53)(54),clock=>clock,reset=>reset,s=>p(162)(54),cout=>p(163)(55));
FA_ff_2231:FAff port map(x=>p(51)(55),y=>p(52)(55),Cin=>p(53)(55),clock=>clock,reset=>reset,s=>p(162)(55),cout=>p(163)(56));
FA_ff_2232:FAff port map(x=>p(51)(56),y=>p(52)(56),Cin=>p(53)(56),clock=>clock,reset=>reset,s=>p(162)(56),cout=>p(163)(57));
FA_ff_2233:FAff port map(x=>p(51)(57),y=>p(52)(57),Cin=>p(53)(57),clock=>clock,reset=>reset,s=>p(162)(57),cout=>p(163)(58));
FA_ff_2234:FAff port map(x=>p(51)(58),y=>p(52)(58),Cin=>p(53)(58),clock=>clock,reset=>reset,s=>p(162)(58),cout=>p(163)(59));
FA_ff_2235:FAff port map(x=>p(51)(59),y=>p(52)(59),Cin=>p(53)(59),clock=>clock,reset=>reset,s=>p(162)(59),cout=>p(163)(60));
FA_ff_2236:FAff port map(x=>p(51)(60),y=>p(52)(60),Cin=>p(53)(60),clock=>clock,reset=>reset,s=>p(162)(60),cout=>p(163)(61));
FA_ff_2237:FAff port map(x=>p(51)(61),y=>p(52)(61),Cin=>p(53)(61),clock=>clock,reset=>reset,s=>p(162)(61),cout=>p(163)(62));
FA_ff_2238:FAff port map(x=>p(51)(62),y=>p(52)(62),Cin=>p(53)(62),clock=>clock,reset=>reset,s=>p(162)(62),cout=>p(163)(63));
FA_ff_2239:FAff port map(x=>p(51)(63),y=>p(52)(63),Cin=>p(53)(63),clock=>clock,reset=>reset,s=>p(162)(63),cout=>p(163)(64));
FA_ff_2240:FAff port map(x=>p(51)(64),y=>p(52)(64),Cin=>p(53)(64),clock=>clock,reset=>reset,s=>p(162)(64),cout=>p(163)(65));
FA_ff_2241:FAff port map(x=>p(51)(65),y=>p(52)(65),Cin=>p(53)(65),clock=>clock,reset=>reset,s=>p(162)(65),cout=>p(163)(66));
FA_ff_2242:FAff port map(x=>p(51)(66),y=>p(52)(66),Cin=>p(53)(66),clock=>clock,reset=>reset,s=>p(162)(66),cout=>p(163)(67));
FA_ff_2243:FAff port map(x=>p(51)(67),y=>p(52)(67),Cin=>p(53)(67),clock=>clock,reset=>reset,s=>p(162)(67),cout=>p(163)(68));
FA_ff_2244:FAff port map(x=>p(51)(68),y=>p(52)(68),Cin=>p(53)(68),clock=>clock,reset=>reset,s=>p(162)(68),cout=>p(163)(69));
FA_ff_2245:FAff port map(x=>p(51)(69),y=>p(52)(69),Cin=>p(53)(69),clock=>clock,reset=>reset,s=>p(162)(69),cout=>p(163)(70));
FA_ff_2246:FAff port map(x=>p(51)(70),y=>p(52)(70),Cin=>p(53)(70),clock=>clock,reset=>reset,s=>p(162)(70),cout=>p(163)(71));
FA_ff_2247:FAff port map(x=>p(51)(71),y=>p(52)(71),Cin=>p(53)(71),clock=>clock,reset=>reset,s=>p(162)(71),cout=>p(163)(72));
FA_ff_2248:FAff port map(x=>p(51)(72),y=>p(52)(72),Cin=>p(53)(72),clock=>clock,reset=>reset,s=>p(162)(72),cout=>p(163)(73));
FA_ff_2249:FAff port map(x=>p(51)(73),y=>p(52)(73),Cin=>p(53)(73),clock=>clock,reset=>reset,s=>p(162)(73),cout=>p(163)(74));
FA_ff_2250:FAff port map(x=>p(51)(74),y=>p(52)(74),Cin=>p(53)(74),clock=>clock,reset=>reset,s=>p(162)(74),cout=>p(163)(75));
FA_ff_2251:FAff port map(x=>p(51)(75),y=>p(52)(75),Cin=>p(53)(75),clock=>clock,reset=>reset,s=>p(162)(75),cout=>p(163)(76));
FA_ff_2252:FAff port map(x=>p(51)(76),y=>p(52)(76),Cin=>p(53)(76),clock=>clock,reset=>reset,s=>p(162)(76),cout=>p(163)(77));
FA_ff_2253:FAff port map(x=>p(51)(77),y=>p(52)(77),Cin=>p(53)(77),clock=>clock,reset=>reset,s=>p(162)(77),cout=>p(163)(78));
FA_ff_2254:FAff port map(x=>p(51)(78),y=>p(52)(78),Cin=>p(53)(78),clock=>clock,reset=>reset,s=>p(162)(78),cout=>p(163)(79));
FA_ff_2255:FAff port map(x=>p(51)(79),y=>p(52)(79),Cin=>p(53)(79),clock=>clock,reset=>reset,s=>p(162)(79),cout=>p(163)(80));
FA_ff_2256:FAff port map(x=>p(51)(80),y=>p(52)(80),Cin=>p(53)(80),clock=>clock,reset=>reset,s=>p(162)(80),cout=>p(163)(81));
FA_ff_2257:FAff port map(x=>p(51)(81),y=>p(52)(81),Cin=>p(53)(81),clock=>clock,reset=>reset,s=>p(162)(81),cout=>p(163)(82));
FA_ff_2258:FAff port map(x=>p(51)(82),y=>p(52)(82),Cin=>p(53)(82),clock=>clock,reset=>reset,s=>p(162)(82),cout=>p(163)(83));
FA_ff_2259:FAff port map(x=>p(51)(83),y=>p(52)(83),Cin=>p(53)(83),clock=>clock,reset=>reset,s=>p(162)(83),cout=>p(163)(84));
FA_ff_2260:FAff port map(x=>p(51)(84),y=>p(52)(84),Cin=>p(53)(84),clock=>clock,reset=>reset,s=>p(162)(84),cout=>p(163)(85));
FA_ff_2261:FAff port map(x=>p(51)(85),y=>p(52)(85),Cin=>p(53)(85),clock=>clock,reset=>reset,s=>p(162)(85),cout=>p(163)(86));
FA_ff_2262:FAff port map(x=>p(51)(86),y=>p(52)(86),Cin=>p(53)(86),clock=>clock,reset=>reset,s=>p(162)(86),cout=>p(163)(87));
FA_ff_2263:FAff port map(x=>p(51)(87),y=>p(52)(87),Cin=>p(53)(87),clock=>clock,reset=>reset,s=>p(162)(87),cout=>p(163)(88));
FA_ff_2264:FAff port map(x=>p(51)(88),y=>p(52)(88),Cin=>p(53)(88),clock=>clock,reset=>reset,s=>p(162)(88),cout=>p(163)(89));
FA_ff_2265:FAff port map(x=>p(51)(89),y=>p(52)(89),Cin=>p(53)(89),clock=>clock,reset=>reset,s=>p(162)(89),cout=>p(163)(90));
FA_ff_2266:FAff port map(x=>p(51)(90),y=>p(52)(90),Cin=>p(53)(90),clock=>clock,reset=>reset,s=>p(162)(90),cout=>p(163)(91));
FA_ff_2267:FAff port map(x=>p(51)(91),y=>p(52)(91),Cin=>p(53)(91),clock=>clock,reset=>reset,s=>p(162)(91),cout=>p(163)(92));
FA_ff_2268:FAff port map(x=>p(51)(92),y=>p(52)(92),Cin=>p(53)(92),clock=>clock,reset=>reset,s=>p(162)(92),cout=>p(163)(93));
FA_ff_2269:FAff port map(x=>p(51)(93),y=>p(52)(93),Cin=>p(53)(93),clock=>clock,reset=>reset,s=>p(162)(93),cout=>p(163)(94));
FA_ff_2270:FAff port map(x=>p(51)(94),y=>p(52)(94),Cin=>p(53)(94),clock=>clock,reset=>reset,s=>p(162)(94),cout=>p(163)(95));
FA_ff_2271:FAff port map(x=>p(51)(95),y=>p(52)(95),Cin=>p(53)(95),clock=>clock,reset=>reset,s=>p(162)(95),cout=>p(163)(96));
FA_ff_2272:FAff port map(x=>p(51)(96),y=>p(52)(96),Cin=>p(53)(96),clock=>clock,reset=>reset,s=>p(162)(96),cout=>p(163)(97));
FA_ff_2273:FAff port map(x=>p(51)(97),y=>p(52)(97),Cin=>p(53)(97),clock=>clock,reset=>reset,s=>p(162)(97),cout=>p(163)(98));
FA_ff_2274:FAff port map(x=>p(51)(98),y=>p(52)(98),Cin=>p(53)(98),clock=>clock,reset=>reset,s=>p(162)(98),cout=>p(163)(99));
FA_ff_2275:FAff port map(x=>p(51)(99),y=>p(52)(99),Cin=>p(53)(99),clock=>clock,reset=>reset,s=>p(162)(99),cout=>p(163)(100));
FA_ff_2276:FAff port map(x=>p(51)(100),y=>p(52)(100),Cin=>p(53)(100),clock=>clock,reset=>reset,s=>p(162)(100),cout=>p(163)(101));
FA_ff_2277:FAff port map(x=>p(51)(101),y=>p(52)(101),Cin=>p(53)(101),clock=>clock,reset=>reset,s=>p(162)(101),cout=>p(163)(102));
FA_ff_2278:FAff port map(x=>p(51)(102),y=>p(52)(102),Cin=>p(53)(102),clock=>clock,reset=>reset,s=>p(162)(102),cout=>p(163)(103));
FA_ff_2279:FAff port map(x=>p(51)(103),y=>p(52)(103),Cin=>p(53)(103),clock=>clock,reset=>reset,s=>p(162)(103),cout=>p(163)(104));
FA_ff_2280:FAff port map(x=>p(51)(104),y=>p(52)(104),Cin=>p(53)(104),clock=>clock,reset=>reset,s=>p(162)(104),cout=>p(163)(105));
FA_ff_2281:FAff port map(x=>p(51)(105),y=>p(52)(105),Cin=>p(53)(105),clock=>clock,reset=>reset,s=>p(162)(105),cout=>p(163)(106));
FA_ff_2282:FAff port map(x=>p(51)(106),y=>p(52)(106),Cin=>p(53)(106),clock=>clock,reset=>reset,s=>p(162)(106),cout=>p(163)(107));
FA_ff_2283:FAff port map(x=>p(51)(107),y=>p(52)(107),Cin=>p(53)(107),clock=>clock,reset=>reset,s=>p(162)(107),cout=>p(163)(108));
FA_ff_2284:FAff port map(x=>p(51)(108),y=>p(52)(108),Cin=>p(53)(108),clock=>clock,reset=>reset,s=>p(162)(108),cout=>p(163)(109));
FA_ff_2285:FAff port map(x=>p(51)(109),y=>p(52)(109),Cin=>p(53)(109),clock=>clock,reset=>reset,s=>p(162)(109),cout=>p(163)(110));
FA_ff_2286:FAff port map(x=>p(51)(110),y=>p(52)(110),Cin=>p(53)(110),clock=>clock,reset=>reset,s=>p(162)(110),cout=>p(163)(111));
FA_ff_2287:FAff port map(x=>p(51)(111),y=>p(52)(111),Cin=>p(53)(111),clock=>clock,reset=>reset,s=>p(162)(111),cout=>p(163)(112));
FA_ff_2288:FAff port map(x=>p(51)(112),y=>p(52)(112),Cin=>p(53)(112),clock=>clock,reset=>reset,s=>p(162)(112),cout=>p(163)(113));
FA_ff_2289:FAff port map(x=>p(51)(113),y=>p(52)(113),Cin=>p(53)(113),clock=>clock,reset=>reset,s=>p(162)(113),cout=>p(163)(114));
FA_ff_2290:FAff port map(x=>p(51)(114),y=>p(52)(114),Cin=>p(53)(114),clock=>clock,reset=>reset,s=>p(162)(114),cout=>p(163)(115));
FA_ff_2291:FAff port map(x=>p(51)(115),y=>p(52)(115),Cin=>p(53)(115),clock=>clock,reset=>reset,s=>p(162)(115),cout=>p(163)(116));
FA_ff_2292:FAff port map(x=>p(51)(116),y=>p(52)(116),Cin=>p(53)(116),clock=>clock,reset=>reset,s=>p(162)(116),cout=>p(163)(117));
FA_ff_2293:FAff port map(x=>p(51)(117),y=>p(52)(117),Cin=>p(53)(117),clock=>clock,reset=>reset,s=>p(162)(117),cout=>p(163)(118));
FA_ff_2294:FAff port map(x=>p(51)(118),y=>p(52)(118),Cin=>p(53)(118),clock=>clock,reset=>reset,s=>p(162)(118),cout=>p(163)(119));
FA_ff_2295:FAff port map(x=>p(51)(119),y=>p(52)(119),Cin=>p(53)(119),clock=>clock,reset=>reset,s=>p(162)(119),cout=>p(163)(120));
FA_ff_2296:FAff port map(x=>p(51)(120),y=>p(52)(120),Cin=>p(53)(120),clock=>clock,reset=>reset,s=>p(162)(120),cout=>p(163)(121));
FA_ff_2297:FAff port map(x=>p(51)(121),y=>p(52)(121),Cin=>p(53)(121),clock=>clock,reset=>reset,s=>p(162)(121),cout=>p(163)(122));
FA_ff_2298:FAff port map(x=>p(51)(122),y=>p(52)(122),Cin=>p(53)(122),clock=>clock,reset=>reset,s=>p(162)(122),cout=>p(163)(123));
FA_ff_2299:FAff port map(x=>p(51)(123),y=>p(52)(123),Cin=>p(53)(123),clock=>clock,reset=>reset,s=>p(162)(123),cout=>p(163)(124));
FA_ff_2300:FAff port map(x=>p(51)(124),y=>p(52)(124),Cin=>p(53)(124),clock=>clock,reset=>reset,s=>p(162)(124),cout=>p(163)(125));
FA_ff_2301:FAff port map(x=>p(51)(125),y=>p(52)(125),Cin=>p(53)(125),clock=>clock,reset=>reset,s=>p(162)(125),cout=>p(163)(126));
FA_ff_2302:FAff port map(x=>p(51)(126),y=>p(52)(126),Cin=>p(53)(126),clock=>clock,reset=>reset,s=>p(162)(126),cout=>p(163)(127));
FA_ff_2303:FAff port map(x=>p(51)(127),y=>p(52)(127),Cin=>p(53)(127),clock=>clock,reset=>reset,s=>p(162)(127),cout=>p(163)(128));
FA_ff_2304:FAff port map(x=>p(54)(0),y=>p(55)(0),Cin=>p(56)(0),clock=>clock,reset=>reset,s=>p(164)(0),cout=>p(165)(1));
FA_ff_2305:FAff port map(x=>p(54)(1),y=>p(55)(1),Cin=>p(56)(1),clock=>clock,reset=>reset,s=>p(164)(1),cout=>p(165)(2));
FA_ff_2306:FAff port map(x=>p(54)(2),y=>p(55)(2),Cin=>p(56)(2),clock=>clock,reset=>reset,s=>p(164)(2),cout=>p(165)(3));
FA_ff_2307:FAff port map(x=>p(54)(3),y=>p(55)(3),Cin=>p(56)(3),clock=>clock,reset=>reset,s=>p(164)(3),cout=>p(165)(4));
FA_ff_2308:FAff port map(x=>p(54)(4),y=>p(55)(4),Cin=>p(56)(4),clock=>clock,reset=>reset,s=>p(164)(4),cout=>p(165)(5));
FA_ff_2309:FAff port map(x=>p(54)(5),y=>p(55)(5),Cin=>p(56)(5),clock=>clock,reset=>reset,s=>p(164)(5),cout=>p(165)(6));
FA_ff_2310:FAff port map(x=>p(54)(6),y=>p(55)(6),Cin=>p(56)(6),clock=>clock,reset=>reset,s=>p(164)(6),cout=>p(165)(7));
FA_ff_2311:FAff port map(x=>p(54)(7),y=>p(55)(7),Cin=>p(56)(7),clock=>clock,reset=>reset,s=>p(164)(7),cout=>p(165)(8));
FA_ff_2312:FAff port map(x=>p(54)(8),y=>p(55)(8),Cin=>p(56)(8),clock=>clock,reset=>reset,s=>p(164)(8),cout=>p(165)(9));
FA_ff_2313:FAff port map(x=>p(54)(9),y=>p(55)(9),Cin=>p(56)(9),clock=>clock,reset=>reset,s=>p(164)(9),cout=>p(165)(10));
FA_ff_2314:FAff port map(x=>p(54)(10),y=>p(55)(10),Cin=>p(56)(10),clock=>clock,reset=>reset,s=>p(164)(10),cout=>p(165)(11));
FA_ff_2315:FAff port map(x=>p(54)(11),y=>p(55)(11),Cin=>p(56)(11),clock=>clock,reset=>reset,s=>p(164)(11),cout=>p(165)(12));
FA_ff_2316:FAff port map(x=>p(54)(12),y=>p(55)(12),Cin=>p(56)(12),clock=>clock,reset=>reset,s=>p(164)(12),cout=>p(165)(13));
FA_ff_2317:FAff port map(x=>p(54)(13),y=>p(55)(13),Cin=>p(56)(13),clock=>clock,reset=>reset,s=>p(164)(13),cout=>p(165)(14));
FA_ff_2318:FAff port map(x=>p(54)(14),y=>p(55)(14),Cin=>p(56)(14),clock=>clock,reset=>reset,s=>p(164)(14),cout=>p(165)(15));
FA_ff_2319:FAff port map(x=>p(54)(15),y=>p(55)(15),Cin=>p(56)(15),clock=>clock,reset=>reset,s=>p(164)(15),cout=>p(165)(16));
FA_ff_2320:FAff port map(x=>p(54)(16),y=>p(55)(16),Cin=>p(56)(16),clock=>clock,reset=>reset,s=>p(164)(16),cout=>p(165)(17));
FA_ff_2321:FAff port map(x=>p(54)(17),y=>p(55)(17),Cin=>p(56)(17),clock=>clock,reset=>reset,s=>p(164)(17),cout=>p(165)(18));
FA_ff_2322:FAff port map(x=>p(54)(18),y=>p(55)(18),Cin=>p(56)(18),clock=>clock,reset=>reset,s=>p(164)(18),cout=>p(165)(19));
FA_ff_2323:FAff port map(x=>p(54)(19),y=>p(55)(19),Cin=>p(56)(19),clock=>clock,reset=>reset,s=>p(164)(19),cout=>p(165)(20));
FA_ff_2324:FAff port map(x=>p(54)(20),y=>p(55)(20),Cin=>p(56)(20),clock=>clock,reset=>reset,s=>p(164)(20),cout=>p(165)(21));
FA_ff_2325:FAff port map(x=>p(54)(21),y=>p(55)(21),Cin=>p(56)(21),clock=>clock,reset=>reset,s=>p(164)(21),cout=>p(165)(22));
FA_ff_2326:FAff port map(x=>p(54)(22),y=>p(55)(22),Cin=>p(56)(22),clock=>clock,reset=>reset,s=>p(164)(22),cout=>p(165)(23));
FA_ff_2327:FAff port map(x=>p(54)(23),y=>p(55)(23),Cin=>p(56)(23),clock=>clock,reset=>reset,s=>p(164)(23),cout=>p(165)(24));
FA_ff_2328:FAff port map(x=>p(54)(24),y=>p(55)(24),Cin=>p(56)(24),clock=>clock,reset=>reset,s=>p(164)(24),cout=>p(165)(25));
FA_ff_2329:FAff port map(x=>p(54)(25),y=>p(55)(25),Cin=>p(56)(25),clock=>clock,reset=>reset,s=>p(164)(25),cout=>p(165)(26));
FA_ff_2330:FAff port map(x=>p(54)(26),y=>p(55)(26),Cin=>p(56)(26),clock=>clock,reset=>reset,s=>p(164)(26),cout=>p(165)(27));
FA_ff_2331:FAff port map(x=>p(54)(27),y=>p(55)(27),Cin=>p(56)(27),clock=>clock,reset=>reset,s=>p(164)(27),cout=>p(165)(28));
FA_ff_2332:FAff port map(x=>p(54)(28),y=>p(55)(28),Cin=>p(56)(28),clock=>clock,reset=>reset,s=>p(164)(28),cout=>p(165)(29));
FA_ff_2333:FAff port map(x=>p(54)(29),y=>p(55)(29),Cin=>p(56)(29),clock=>clock,reset=>reset,s=>p(164)(29),cout=>p(165)(30));
FA_ff_2334:FAff port map(x=>p(54)(30),y=>p(55)(30),Cin=>p(56)(30),clock=>clock,reset=>reset,s=>p(164)(30),cout=>p(165)(31));
FA_ff_2335:FAff port map(x=>p(54)(31),y=>p(55)(31),Cin=>p(56)(31),clock=>clock,reset=>reset,s=>p(164)(31),cout=>p(165)(32));
FA_ff_2336:FAff port map(x=>p(54)(32),y=>p(55)(32),Cin=>p(56)(32),clock=>clock,reset=>reset,s=>p(164)(32),cout=>p(165)(33));
FA_ff_2337:FAff port map(x=>p(54)(33),y=>p(55)(33),Cin=>p(56)(33),clock=>clock,reset=>reset,s=>p(164)(33),cout=>p(165)(34));
FA_ff_2338:FAff port map(x=>p(54)(34),y=>p(55)(34),Cin=>p(56)(34),clock=>clock,reset=>reset,s=>p(164)(34),cout=>p(165)(35));
FA_ff_2339:FAff port map(x=>p(54)(35),y=>p(55)(35),Cin=>p(56)(35),clock=>clock,reset=>reset,s=>p(164)(35),cout=>p(165)(36));
FA_ff_2340:FAff port map(x=>p(54)(36),y=>p(55)(36),Cin=>p(56)(36),clock=>clock,reset=>reset,s=>p(164)(36),cout=>p(165)(37));
FA_ff_2341:FAff port map(x=>p(54)(37),y=>p(55)(37),Cin=>p(56)(37),clock=>clock,reset=>reset,s=>p(164)(37),cout=>p(165)(38));
FA_ff_2342:FAff port map(x=>p(54)(38),y=>p(55)(38),Cin=>p(56)(38),clock=>clock,reset=>reset,s=>p(164)(38),cout=>p(165)(39));
FA_ff_2343:FAff port map(x=>p(54)(39),y=>p(55)(39),Cin=>p(56)(39),clock=>clock,reset=>reset,s=>p(164)(39),cout=>p(165)(40));
FA_ff_2344:FAff port map(x=>p(54)(40),y=>p(55)(40),Cin=>p(56)(40),clock=>clock,reset=>reset,s=>p(164)(40),cout=>p(165)(41));
FA_ff_2345:FAff port map(x=>p(54)(41),y=>p(55)(41),Cin=>p(56)(41),clock=>clock,reset=>reset,s=>p(164)(41),cout=>p(165)(42));
FA_ff_2346:FAff port map(x=>p(54)(42),y=>p(55)(42),Cin=>p(56)(42),clock=>clock,reset=>reset,s=>p(164)(42),cout=>p(165)(43));
FA_ff_2347:FAff port map(x=>p(54)(43),y=>p(55)(43),Cin=>p(56)(43),clock=>clock,reset=>reset,s=>p(164)(43),cout=>p(165)(44));
FA_ff_2348:FAff port map(x=>p(54)(44),y=>p(55)(44),Cin=>p(56)(44),clock=>clock,reset=>reset,s=>p(164)(44),cout=>p(165)(45));
FA_ff_2349:FAff port map(x=>p(54)(45),y=>p(55)(45),Cin=>p(56)(45),clock=>clock,reset=>reset,s=>p(164)(45),cout=>p(165)(46));
FA_ff_2350:FAff port map(x=>p(54)(46),y=>p(55)(46),Cin=>p(56)(46),clock=>clock,reset=>reset,s=>p(164)(46),cout=>p(165)(47));
FA_ff_2351:FAff port map(x=>p(54)(47),y=>p(55)(47),Cin=>p(56)(47),clock=>clock,reset=>reset,s=>p(164)(47),cout=>p(165)(48));
FA_ff_2352:FAff port map(x=>p(54)(48),y=>p(55)(48),Cin=>p(56)(48),clock=>clock,reset=>reset,s=>p(164)(48),cout=>p(165)(49));
FA_ff_2353:FAff port map(x=>p(54)(49),y=>p(55)(49),Cin=>p(56)(49),clock=>clock,reset=>reset,s=>p(164)(49),cout=>p(165)(50));
FA_ff_2354:FAff port map(x=>p(54)(50),y=>p(55)(50),Cin=>p(56)(50),clock=>clock,reset=>reset,s=>p(164)(50),cout=>p(165)(51));
FA_ff_2355:FAff port map(x=>p(54)(51),y=>p(55)(51),Cin=>p(56)(51),clock=>clock,reset=>reset,s=>p(164)(51),cout=>p(165)(52));
FA_ff_2356:FAff port map(x=>p(54)(52),y=>p(55)(52),Cin=>p(56)(52),clock=>clock,reset=>reset,s=>p(164)(52),cout=>p(165)(53));
FA_ff_2357:FAff port map(x=>p(54)(53),y=>p(55)(53),Cin=>p(56)(53),clock=>clock,reset=>reset,s=>p(164)(53),cout=>p(165)(54));
FA_ff_2358:FAff port map(x=>p(54)(54),y=>p(55)(54),Cin=>p(56)(54),clock=>clock,reset=>reset,s=>p(164)(54),cout=>p(165)(55));
FA_ff_2359:FAff port map(x=>p(54)(55),y=>p(55)(55),Cin=>p(56)(55),clock=>clock,reset=>reset,s=>p(164)(55),cout=>p(165)(56));
FA_ff_2360:FAff port map(x=>p(54)(56),y=>p(55)(56),Cin=>p(56)(56),clock=>clock,reset=>reset,s=>p(164)(56),cout=>p(165)(57));
FA_ff_2361:FAff port map(x=>p(54)(57),y=>p(55)(57),Cin=>p(56)(57),clock=>clock,reset=>reset,s=>p(164)(57),cout=>p(165)(58));
FA_ff_2362:FAff port map(x=>p(54)(58),y=>p(55)(58),Cin=>p(56)(58),clock=>clock,reset=>reset,s=>p(164)(58),cout=>p(165)(59));
FA_ff_2363:FAff port map(x=>p(54)(59),y=>p(55)(59),Cin=>p(56)(59),clock=>clock,reset=>reset,s=>p(164)(59),cout=>p(165)(60));
FA_ff_2364:FAff port map(x=>p(54)(60),y=>p(55)(60),Cin=>p(56)(60),clock=>clock,reset=>reset,s=>p(164)(60),cout=>p(165)(61));
FA_ff_2365:FAff port map(x=>p(54)(61),y=>p(55)(61),Cin=>p(56)(61),clock=>clock,reset=>reset,s=>p(164)(61),cout=>p(165)(62));
FA_ff_2366:FAff port map(x=>p(54)(62),y=>p(55)(62),Cin=>p(56)(62),clock=>clock,reset=>reset,s=>p(164)(62),cout=>p(165)(63));
FA_ff_2367:FAff port map(x=>p(54)(63),y=>p(55)(63),Cin=>p(56)(63),clock=>clock,reset=>reset,s=>p(164)(63),cout=>p(165)(64));
FA_ff_2368:FAff port map(x=>p(54)(64),y=>p(55)(64),Cin=>p(56)(64),clock=>clock,reset=>reset,s=>p(164)(64),cout=>p(165)(65));
FA_ff_2369:FAff port map(x=>p(54)(65),y=>p(55)(65),Cin=>p(56)(65),clock=>clock,reset=>reset,s=>p(164)(65),cout=>p(165)(66));
FA_ff_2370:FAff port map(x=>p(54)(66),y=>p(55)(66),Cin=>p(56)(66),clock=>clock,reset=>reset,s=>p(164)(66),cout=>p(165)(67));
FA_ff_2371:FAff port map(x=>p(54)(67),y=>p(55)(67),Cin=>p(56)(67),clock=>clock,reset=>reset,s=>p(164)(67),cout=>p(165)(68));
FA_ff_2372:FAff port map(x=>p(54)(68),y=>p(55)(68),Cin=>p(56)(68),clock=>clock,reset=>reset,s=>p(164)(68),cout=>p(165)(69));
FA_ff_2373:FAff port map(x=>p(54)(69),y=>p(55)(69),Cin=>p(56)(69),clock=>clock,reset=>reset,s=>p(164)(69),cout=>p(165)(70));
FA_ff_2374:FAff port map(x=>p(54)(70),y=>p(55)(70),Cin=>p(56)(70),clock=>clock,reset=>reset,s=>p(164)(70),cout=>p(165)(71));
FA_ff_2375:FAff port map(x=>p(54)(71),y=>p(55)(71),Cin=>p(56)(71),clock=>clock,reset=>reset,s=>p(164)(71),cout=>p(165)(72));
FA_ff_2376:FAff port map(x=>p(54)(72),y=>p(55)(72),Cin=>p(56)(72),clock=>clock,reset=>reset,s=>p(164)(72),cout=>p(165)(73));
FA_ff_2377:FAff port map(x=>p(54)(73),y=>p(55)(73),Cin=>p(56)(73),clock=>clock,reset=>reset,s=>p(164)(73),cout=>p(165)(74));
FA_ff_2378:FAff port map(x=>p(54)(74),y=>p(55)(74),Cin=>p(56)(74),clock=>clock,reset=>reset,s=>p(164)(74),cout=>p(165)(75));
FA_ff_2379:FAff port map(x=>p(54)(75),y=>p(55)(75),Cin=>p(56)(75),clock=>clock,reset=>reset,s=>p(164)(75),cout=>p(165)(76));
FA_ff_2380:FAff port map(x=>p(54)(76),y=>p(55)(76),Cin=>p(56)(76),clock=>clock,reset=>reset,s=>p(164)(76),cout=>p(165)(77));
FA_ff_2381:FAff port map(x=>p(54)(77),y=>p(55)(77),Cin=>p(56)(77),clock=>clock,reset=>reset,s=>p(164)(77),cout=>p(165)(78));
FA_ff_2382:FAff port map(x=>p(54)(78),y=>p(55)(78),Cin=>p(56)(78),clock=>clock,reset=>reset,s=>p(164)(78),cout=>p(165)(79));
FA_ff_2383:FAff port map(x=>p(54)(79),y=>p(55)(79),Cin=>p(56)(79),clock=>clock,reset=>reset,s=>p(164)(79),cout=>p(165)(80));
FA_ff_2384:FAff port map(x=>p(54)(80),y=>p(55)(80),Cin=>p(56)(80),clock=>clock,reset=>reset,s=>p(164)(80),cout=>p(165)(81));
FA_ff_2385:FAff port map(x=>p(54)(81),y=>p(55)(81),Cin=>p(56)(81),clock=>clock,reset=>reset,s=>p(164)(81),cout=>p(165)(82));
FA_ff_2386:FAff port map(x=>p(54)(82),y=>p(55)(82),Cin=>p(56)(82),clock=>clock,reset=>reset,s=>p(164)(82),cout=>p(165)(83));
FA_ff_2387:FAff port map(x=>p(54)(83),y=>p(55)(83),Cin=>p(56)(83),clock=>clock,reset=>reset,s=>p(164)(83),cout=>p(165)(84));
FA_ff_2388:FAff port map(x=>p(54)(84),y=>p(55)(84),Cin=>p(56)(84),clock=>clock,reset=>reset,s=>p(164)(84),cout=>p(165)(85));
FA_ff_2389:FAff port map(x=>p(54)(85),y=>p(55)(85),Cin=>p(56)(85),clock=>clock,reset=>reset,s=>p(164)(85),cout=>p(165)(86));
FA_ff_2390:FAff port map(x=>p(54)(86),y=>p(55)(86),Cin=>p(56)(86),clock=>clock,reset=>reset,s=>p(164)(86),cout=>p(165)(87));
FA_ff_2391:FAff port map(x=>p(54)(87),y=>p(55)(87),Cin=>p(56)(87),clock=>clock,reset=>reset,s=>p(164)(87),cout=>p(165)(88));
FA_ff_2392:FAff port map(x=>p(54)(88),y=>p(55)(88),Cin=>p(56)(88),clock=>clock,reset=>reset,s=>p(164)(88),cout=>p(165)(89));
FA_ff_2393:FAff port map(x=>p(54)(89),y=>p(55)(89),Cin=>p(56)(89),clock=>clock,reset=>reset,s=>p(164)(89),cout=>p(165)(90));
FA_ff_2394:FAff port map(x=>p(54)(90),y=>p(55)(90),Cin=>p(56)(90),clock=>clock,reset=>reset,s=>p(164)(90),cout=>p(165)(91));
FA_ff_2395:FAff port map(x=>p(54)(91),y=>p(55)(91),Cin=>p(56)(91),clock=>clock,reset=>reset,s=>p(164)(91),cout=>p(165)(92));
FA_ff_2396:FAff port map(x=>p(54)(92),y=>p(55)(92),Cin=>p(56)(92),clock=>clock,reset=>reset,s=>p(164)(92),cout=>p(165)(93));
FA_ff_2397:FAff port map(x=>p(54)(93),y=>p(55)(93),Cin=>p(56)(93),clock=>clock,reset=>reset,s=>p(164)(93),cout=>p(165)(94));
FA_ff_2398:FAff port map(x=>p(54)(94),y=>p(55)(94),Cin=>p(56)(94),clock=>clock,reset=>reset,s=>p(164)(94),cout=>p(165)(95));
FA_ff_2399:FAff port map(x=>p(54)(95),y=>p(55)(95),Cin=>p(56)(95),clock=>clock,reset=>reset,s=>p(164)(95),cout=>p(165)(96));
FA_ff_2400:FAff port map(x=>p(54)(96),y=>p(55)(96),Cin=>p(56)(96),clock=>clock,reset=>reset,s=>p(164)(96),cout=>p(165)(97));
FA_ff_2401:FAff port map(x=>p(54)(97),y=>p(55)(97),Cin=>p(56)(97),clock=>clock,reset=>reset,s=>p(164)(97),cout=>p(165)(98));
FA_ff_2402:FAff port map(x=>p(54)(98),y=>p(55)(98),Cin=>p(56)(98),clock=>clock,reset=>reset,s=>p(164)(98),cout=>p(165)(99));
FA_ff_2403:FAff port map(x=>p(54)(99),y=>p(55)(99),Cin=>p(56)(99),clock=>clock,reset=>reset,s=>p(164)(99),cout=>p(165)(100));
FA_ff_2404:FAff port map(x=>p(54)(100),y=>p(55)(100),Cin=>p(56)(100),clock=>clock,reset=>reset,s=>p(164)(100),cout=>p(165)(101));
FA_ff_2405:FAff port map(x=>p(54)(101),y=>p(55)(101),Cin=>p(56)(101),clock=>clock,reset=>reset,s=>p(164)(101),cout=>p(165)(102));
FA_ff_2406:FAff port map(x=>p(54)(102),y=>p(55)(102),Cin=>p(56)(102),clock=>clock,reset=>reset,s=>p(164)(102),cout=>p(165)(103));
FA_ff_2407:FAff port map(x=>p(54)(103),y=>p(55)(103),Cin=>p(56)(103),clock=>clock,reset=>reset,s=>p(164)(103),cout=>p(165)(104));
FA_ff_2408:FAff port map(x=>p(54)(104),y=>p(55)(104),Cin=>p(56)(104),clock=>clock,reset=>reset,s=>p(164)(104),cout=>p(165)(105));
FA_ff_2409:FAff port map(x=>p(54)(105),y=>p(55)(105),Cin=>p(56)(105),clock=>clock,reset=>reset,s=>p(164)(105),cout=>p(165)(106));
FA_ff_2410:FAff port map(x=>p(54)(106),y=>p(55)(106),Cin=>p(56)(106),clock=>clock,reset=>reset,s=>p(164)(106),cout=>p(165)(107));
FA_ff_2411:FAff port map(x=>p(54)(107),y=>p(55)(107),Cin=>p(56)(107),clock=>clock,reset=>reset,s=>p(164)(107),cout=>p(165)(108));
FA_ff_2412:FAff port map(x=>p(54)(108),y=>p(55)(108),Cin=>p(56)(108),clock=>clock,reset=>reset,s=>p(164)(108),cout=>p(165)(109));
FA_ff_2413:FAff port map(x=>p(54)(109),y=>p(55)(109),Cin=>p(56)(109),clock=>clock,reset=>reset,s=>p(164)(109),cout=>p(165)(110));
FA_ff_2414:FAff port map(x=>p(54)(110),y=>p(55)(110),Cin=>p(56)(110),clock=>clock,reset=>reset,s=>p(164)(110),cout=>p(165)(111));
FA_ff_2415:FAff port map(x=>p(54)(111),y=>p(55)(111),Cin=>p(56)(111),clock=>clock,reset=>reset,s=>p(164)(111),cout=>p(165)(112));
FA_ff_2416:FAff port map(x=>p(54)(112),y=>p(55)(112),Cin=>p(56)(112),clock=>clock,reset=>reset,s=>p(164)(112),cout=>p(165)(113));
FA_ff_2417:FAff port map(x=>p(54)(113),y=>p(55)(113),Cin=>p(56)(113),clock=>clock,reset=>reset,s=>p(164)(113),cout=>p(165)(114));
FA_ff_2418:FAff port map(x=>p(54)(114),y=>p(55)(114),Cin=>p(56)(114),clock=>clock,reset=>reset,s=>p(164)(114),cout=>p(165)(115));
FA_ff_2419:FAff port map(x=>p(54)(115),y=>p(55)(115),Cin=>p(56)(115),clock=>clock,reset=>reset,s=>p(164)(115),cout=>p(165)(116));
FA_ff_2420:FAff port map(x=>p(54)(116),y=>p(55)(116),Cin=>p(56)(116),clock=>clock,reset=>reset,s=>p(164)(116),cout=>p(165)(117));
FA_ff_2421:FAff port map(x=>p(54)(117),y=>p(55)(117),Cin=>p(56)(117),clock=>clock,reset=>reset,s=>p(164)(117),cout=>p(165)(118));
FA_ff_2422:FAff port map(x=>p(54)(118),y=>p(55)(118),Cin=>p(56)(118),clock=>clock,reset=>reset,s=>p(164)(118),cout=>p(165)(119));
FA_ff_2423:FAff port map(x=>p(54)(119),y=>p(55)(119),Cin=>p(56)(119),clock=>clock,reset=>reset,s=>p(164)(119),cout=>p(165)(120));
FA_ff_2424:FAff port map(x=>p(54)(120),y=>p(55)(120),Cin=>p(56)(120),clock=>clock,reset=>reset,s=>p(164)(120),cout=>p(165)(121));
FA_ff_2425:FAff port map(x=>p(54)(121),y=>p(55)(121),Cin=>p(56)(121),clock=>clock,reset=>reset,s=>p(164)(121),cout=>p(165)(122));
FA_ff_2426:FAff port map(x=>p(54)(122),y=>p(55)(122),Cin=>p(56)(122),clock=>clock,reset=>reset,s=>p(164)(122),cout=>p(165)(123));
FA_ff_2427:FAff port map(x=>p(54)(123),y=>p(55)(123),Cin=>p(56)(123),clock=>clock,reset=>reset,s=>p(164)(123),cout=>p(165)(124));
FA_ff_2428:FAff port map(x=>p(54)(124),y=>p(55)(124),Cin=>p(56)(124),clock=>clock,reset=>reset,s=>p(164)(124),cout=>p(165)(125));
FA_ff_2429:FAff port map(x=>p(54)(125),y=>p(55)(125),Cin=>p(56)(125),clock=>clock,reset=>reset,s=>p(164)(125),cout=>p(165)(126));
FA_ff_2430:FAff port map(x=>p(54)(126),y=>p(55)(126),Cin=>p(56)(126),clock=>clock,reset=>reset,s=>p(164)(126),cout=>p(165)(127));
FA_ff_2431:FAff port map(x=>p(54)(127),y=>p(55)(127),Cin=>p(56)(127),clock=>clock,reset=>reset,s=>p(164)(127),cout=>p(165)(128));
FA_ff_2432:FAff port map(x=>p(57)(0),y=>p(58)(0),Cin=>p(59)(0),clock=>clock,reset=>reset,s=>p(166)(0),cout=>p(167)(1));
FA_ff_2433:FAff port map(x=>p(57)(1),y=>p(58)(1),Cin=>p(59)(1),clock=>clock,reset=>reset,s=>p(166)(1),cout=>p(167)(2));
FA_ff_2434:FAff port map(x=>p(57)(2),y=>p(58)(2),Cin=>p(59)(2),clock=>clock,reset=>reset,s=>p(166)(2),cout=>p(167)(3));
FA_ff_2435:FAff port map(x=>p(57)(3),y=>p(58)(3),Cin=>p(59)(3),clock=>clock,reset=>reset,s=>p(166)(3),cout=>p(167)(4));
FA_ff_2436:FAff port map(x=>p(57)(4),y=>p(58)(4),Cin=>p(59)(4),clock=>clock,reset=>reset,s=>p(166)(4),cout=>p(167)(5));
FA_ff_2437:FAff port map(x=>p(57)(5),y=>p(58)(5),Cin=>p(59)(5),clock=>clock,reset=>reset,s=>p(166)(5),cout=>p(167)(6));
FA_ff_2438:FAff port map(x=>p(57)(6),y=>p(58)(6),Cin=>p(59)(6),clock=>clock,reset=>reset,s=>p(166)(6),cout=>p(167)(7));
FA_ff_2439:FAff port map(x=>p(57)(7),y=>p(58)(7),Cin=>p(59)(7),clock=>clock,reset=>reset,s=>p(166)(7),cout=>p(167)(8));
FA_ff_2440:FAff port map(x=>p(57)(8),y=>p(58)(8),Cin=>p(59)(8),clock=>clock,reset=>reset,s=>p(166)(8),cout=>p(167)(9));
FA_ff_2441:FAff port map(x=>p(57)(9),y=>p(58)(9),Cin=>p(59)(9),clock=>clock,reset=>reset,s=>p(166)(9),cout=>p(167)(10));
FA_ff_2442:FAff port map(x=>p(57)(10),y=>p(58)(10),Cin=>p(59)(10),clock=>clock,reset=>reset,s=>p(166)(10),cout=>p(167)(11));
FA_ff_2443:FAff port map(x=>p(57)(11),y=>p(58)(11),Cin=>p(59)(11),clock=>clock,reset=>reset,s=>p(166)(11),cout=>p(167)(12));
FA_ff_2444:FAff port map(x=>p(57)(12),y=>p(58)(12),Cin=>p(59)(12),clock=>clock,reset=>reset,s=>p(166)(12),cout=>p(167)(13));
FA_ff_2445:FAff port map(x=>p(57)(13),y=>p(58)(13),Cin=>p(59)(13),clock=>clock,reset=>reset,s=>p(166)(13),cout=>p(167)(14));
FA_ff_2446:FAff port map(x=>p(57)(14),y=>p(58)(14),Cin=>p(59)(14),clock=>clock,reset=>reset,s=>p(166)(14),cout=>p(167)(15));
FA_ff_2447:FAff port map(x=>p(57)(15),y=>p(58)(15),Cin=>p(59)(15),clock=>clock,reset=>reset,s=>p(166)(15),cout=>p(167)(16));
FA_ff_2448:FAff port map(x=>p(57)(16),y=>p(58)(16),Cin=>p(59)(16),clock=>clock,reset=>reset,s=>p(166)(16),cout=>p(167)(17));
FA_ff_2449:FAff port map(x=>p(57)(17),y=>p(58)(17),Cin=>p(59)(17),clock=>clock,reset=>reset,s=>p(166)(17),cout=>p(167)(18));
FA_ff_2450:FAff port map(x=>p(57)(18),y=>p(58)(18),Cin=>p(59)(18),clock=>clock,reset=>reset,s=>p(166)(18),cout=>p(167)(19));
FA_ff_2451:FAff port map(x=>p(57)(19),y=>p(58)(19),Cin=>p(59)(19),clock=>clock,reset=>reset,s=>p(166)(19),cout=>p(167)(20));
FA_ff_2452:FAff port map(x=>p(57)(20),y=>p(58)(20),Cin=>p(59)(20),clock=>clock,reset=>reset,s=>p(166)(20),cout=>p(167)(21));
FA_ff_2453:FAff port map(x=>p(57)(21),y=>p(58)(21),Cin=>p(59)(21),clock=>clock,reset=>reset,s=>p(166)(21),cout=>p(167)(22));
FA_ff_2454:FAff port map(x=>p(57)(22),y=>p(58)(22),Cin=>p(59)(22),clock=>clock,reset=>reset,s=>p(166)(22),cout=>p(167)(23));
FA_ff_2455:FAff port map(x=>p(57)(23),y=>p(58)(23),Cin=>p(59)(23),clock=>clock,reset=>reset,s=>p(166)(23),cout=>p(167)(24));
FA_ff_2456:FAff port map(x=>p(57)(24),y=>p(58)(24),Cin=>p(59)(24),clock=>clock,reset=>reset,s=>p(166)(24),cout=>p(167)(25));
FA_ff_2457:FAff port map(x=>p(57)(25),y=>p(58)(25),Cin=>p(59)(25),clock=>clock,reset=>reset,s=>p(166)(25),cout=>p(167)(26));
FA_ff_2458:FAff port map(x=>p(57)(26),y=>p(58)(26),Cin=>p(59)(26),clock=>clock,reset=>reset,s=>p(166)(26),cout=>p(167)(27));
FA_ff_2459:FAff port map(x=>p(57)(27),y=>p(58)(27),Cin=>p(59)(27),clock=>clock,reset=>reset,s=>p(166)(27),cout=>p(167)(28));
FA_ff_2460:FAff port map(x=>p(57)(28),y=>p(58)(28),Cin=>p(59)(28),clock=>clock,reset=>reset,s=>p(166)(28),cout=>p(167)(29));
FA_ff_2461:FAff port map(x=>p(57)(29),y=>p(58)(29),Cin=>p(59)(29),clock=>clock,reset=>reset,s=>p(166)(29),cout=>p(167)(30));
FA_ff_2462:FAff port map(x=>p(57)(30),y=>p(58)(30),Cin=>p(59)(30),clock=>clock,reset=>reset,s=>p(166)(30),cout=>p(167)(31));
FA_ff_2463:FAff port map(x=>p(57)(31),y=>p(58)(31),Cin=>p(59)(31),clock=>clock,reset=>reset,s=>p(166)(31),cout=>p(167)(32));
FA_ff_2464:FAff port map(x=>p(57)(32),y=>p(58)(32),Cin=>p(59)(32),clock=>clock,reset=>reset,s=>p(166)(32),cout=>p(167)(33));
FA_ff_2465:FAff port map(x=>p(57)(33),y=>p(58)(33),Cin=>p(59)(33),clock=>clock,reset=>reset,s=>p(166)(33),cout=>p(167)(34));
FA_ff_2466:FAff port map(x=>p(57)(34),y=>p(58)(34),Cin=>p(59)(34),clock=>clock,reset=>reset,s=>p(166)(34),cout=>p(167)(35));
FA_ff_2467:FAff port map(x=>p(57)(35),y=>p(58)(35),Cin=>p(59)(35),clock=>clock,reset=>reset,s=>p(166)(35),cout=>p(167)(36));
FA_ff_2468:FAff port map(x=>p(57)(36),y=>p(58)(36),Cin=>p(59)(36),clock=>clock,reset=>reset,s=>p(166)(36),cout=>p(167)(37));
FA_ff_2469:FAff port map(x=>p(57)(37),y=>p(58)(37),Cin=>p(59)(37),clock=>clock,reset=>reset,s=>p(166)(37),cout=>p(167)(38));
FA_ff_2470:FAff port map(x=>p(57)(38),y=>p(58)(38),Cin=>p(59)(38),clock=>clock,reset=>reset,s=>p(166)(38),cout=>p(167)(39));
FA_ff_2471:FAff port map(x=>p(57)(39),y=>p(58)(39),Cin=>p(59)(39),clock=>clock,reset=>reset,s=>p(166)(39),cout=>p(167)(40));
FA_ff_2472:FAff port map(x=>p(57)(40),y=>p(58)(40),Cin=>p(59)(40),clock=>clock,reset=>reset,s=>p(166)(40),cout=>p(167)(41));
FA_ff_2473:FAff port map(x=>p(57)(41),y=>p(58)(41),Cin=>p(59)(41),clock=>clock,reset=>reset,s=>p(166)(41),cout=>p(167)(42));
FA_ff_2474:FAff port map(x=>p(57)(42),y=>p(58)(42),Cin=>p(59)(42),clock=>clock,reset=>reset,s=>p(166)(42),cout=>p(167)(43));
FA_ff_2475:FAff port map(x=>p(57)(43),y=>p(58)(43),Cin=>p(59)(43),clock=>clock,reset=>reset,s=>p(166)(43),cout=>p(167)(44));
FA_ff_2476:FAff port map(x=>p(57)(44),y=>p(58)(44),Cin=>p(59)(44),clock=>clock,reset=>reset,s=>p(166)(44),cout=>p(167)(45));
FA_ff_2477:FAff port map(x=>p(57)(45),y=>p(58)(45),Cin=>p(59)(45),clock=>clock,reset=>reset,s=>p(166)(45),cout=>p(167)(46));
FA_ff_2478:FAff port map(x=>p(57)(46),y=>p(58)(46),Cin=>p(59)(46),clock=>clock,reset=>reset,s=>p(166)(46),cout=>p(167)(47));
FA_ff_2479:FAff port map(x=>p(57)(47),y=>p(58)(47),Cin=>p(59)(47),clock=>clock,reset=>reset,s=>p(166)(47),cout=>p(167)(48));
FA_ff_2480:FAff port map(x=>p(57)(48),y=>p(58)(48),Cin=>p(59)(48),clock=>clock,reset=>reset,s=>p(166)(48),cout=>p(167)(49));
FA_ff_2481:FAff port map(x=>p(57)(49),y=>p(58)(49),Cin=>p(59)(49),clock=>clock,reset=>reset,s=>p(166)(49),cout=>p(167)(50));
FA_ff_2482:FAff port map(x=>p(57)(50),y=>p(58)(50),Cin=>p(59)(50),clock=>clock,reset=>reset,s=>p(166)(50),cout=>p(167)(51));
FA_ff_2483:FAff port map(x=>p(57)(51),y=>p(58)(51),Cin=>p(59)(51),clock=>clock,reset=>reset,s=>p(166)(51),cout=>p(167)(52));
FA_ff_2484:FAff port map(x=>p(57)(52),y=>p(58)(52),Cin=>p(59)(52),clock=>clock,reset=>reset,s=>p(166)(52),cout=>p(167)(53));
FA_ff_2485:FAff port map(x=>p(57)(53),y=>p(58)(53),Cin=>p(59)(53),clock=>clock,reset=>reset,s=>p(166)(53),cout=>p(167)(54));
FA_ff_2486:FAff port map(x=>p(57)(54),y=>p(58)(54),Cin=>p(59)(54),clock=>clock,reset=>reset,s=>p(166)(54),cout=>p(167)(55));
FA_ff_2487:FAff port map(x=>p(57)(55),y=>p(58)(55),Cin=>p(59)(55),clock=>clock,reset=>reset,s=>p(166)(55),cout=>p(167)(56));
FA_ff_2488:FAff port map(x=>p(57)(56),y=>p(58)(56),Cin=>p(59)(56),clock=>clock,reset=>reset,s=>p(166)(56),cout=>p(167)(57));
FA_ff_2489:FAff port map(x=>p(57)(57),y=>p(58)(57),Cin=>p(59)(57),clock=>clock,reset=>reset,s=>p(166)(57),cout=>p(167)(58));
FA_ff_2490:FAff port map(x=>p(57)(58),y=>p(58)(58),Cin=>p(59)(58),clock=>clock,reset=>reset,s=>p(166)(58),cout=>p(167)(59));
FA_ff_2491:FAff port map(x=>p(57)(59),y=>p(58)(59),Cin=>p(59)(59),clock=>clock,reset=>reset,s=>p(166)(59),cout=>p(167)(60));
FA_ff_2492:FAff port map(x=>p(57)(60),y=>p(58)(60),Cin=>p(59)(60),clock=>clock,reset=>reset,s=>p(166)(60),cout=>p(167)(61));
FA_ff_2493:FAff port map(x=>p(57)(61),y=>p(58)(61),Cin=>p(59)(61),clock=>clock,reset=>reset,s=>p(166)(61),cout=>p(167)(62));
FA_ff_2494:FAff port map(x=>p(57)(62),y=>p(58)(62),Cin=>p(59)(62),clock=>clock,reset=>reset,s=>p(166)(62),cout=>p(167)(63));
FA_ff_2495:FAff port map(x=>p(57)(63),y=>p(58)(63),Cin=>p(59)(63),clock=>clock,reset=>reset,s=>p(166)(63),cout=>p(167)(64));
FA_ff_2496:FAff port map(x=>p(57)(64),y=>p(58)(64),Cin=>p(59)(64),clock=>clock,reset=>reset,s=>p(166)(64),cout=>p(167)(65));
FA_ff_2497:FAff port map(x=>p(57)(65),y=>p(58)(65),Cin=>p(59)(65),clock=>clock,reset=>reset,s=>p(166)(65),cout=>p(167)(66));
FA_ff_2498:FAff port map(x=>p(57)(66),y=>p(58)(66),Cin=>p(59)(66),clock=>clock,reset=>reset,s=>p(166)(66),cout=>p(167)(67));
FA_ff_2499:FAff port map(x=>p(57)(67),y=>p(58)(67),Cin=>p(59)(67),clock=>clock,reset=>reset,s=>p(166)(67),cout=>p(167)(68));
FA_ff_2500:FAff port map(x=>p(57)(68),y=>p(58)(68),Cin=>p(59)(68),clock=>clock,reset=>reset,s=>p(166)(68),cout=>p(167)(69));
FA_ff_2501:FAff port map(x=>p(57)(69),y=>p(58)(69),Cin=>p(59)(69),clock=>clock,reset=>reset,s=>p(166)(69),cout=>p(167)(70));
FA_ff_2502:FAff port map(x=>p(57)(70),y=>p(58)(70),Cin=>p(59)(70),clock=>clock,reset=>reset,s=>p(166)(70),cout=>p(167)(71));
FA_ff_2503:FAff port map(x=>p(57)(71),y=>p(58)(71),Cin=>p(59)(71),clock=>clock,reset=>reset,s=>p(166)(71),cout=>p(167)(72));
FA_ff_2504:FAff port map(x=>p(57)(72),y=>p(58)(72),Cin=>p(59)(72),clock=>clock,reset=>reset,s=>p(166)(72),cout=>p(167)(73));
FA_ff_2505:FAff port map(x=>p(57)(73),y=>p(58)(73),Cin=>p(59)(73),clock=>clock,reset=>reset,s=>p(166)(73),cout=>p(167)(74));
FA_ff_2506:FAff port map(x=>p(57)(74),y=>p(58)(74),Cin=>p(59)(74),clock=>clock,reset=>reset,s=>p(166)(74),cout=>p(167)(75));
FA_ff_2507:FAff port map(x=>p(57)(75),y=>p(58)(75),Cin=>p(59)(75),clock=>clock,reset=>reset,s=>p(166)(75),cout=>p(167)(76));
FA_ff_2508:FAff port map(x=>p(57)(76),y=>p(58)(76),Cin=>p(59)(76),clock=>clock,reset=>reset,s=>p(166)(76),cout=>p(167)(77));
FA_ff_2509:FAff port map(x=>p(57)(77),y=>p(58)(77),Cin=>p(59)(77),clock=>clock,reset=>reset,s=>p(166)(77),cout=>p(167)(78));
FA_ff_2510:FAff port map(x=>p(57)(78),y=>p(58)(78),Cin=>p(59)(78),clock=>clock,reset=>reset,s=>p(166)(78),cout=>p(167)(79));
FA_ff_2511:FAff port map(x=>p(57)(79),y=>p(58)(79),Cin=>p(59)(79),clock=>clock,reset=>reset,s=>p(166)(79),cout=>p(167)(80));
FA_ff_2512:FAff port map(x=>p(57)(80),y=>p(58)(80),Cin=>p(59)(80),clock=>clock,reset=>reset,s=>p(166)(80),cout=>p(167)(81));
FA_ff_2513:FAff port map(x=>p(57)(81),y=>p(58)(81),Cin=>p(59)(81),clock=>clock,reset=>reset,s=>p(166)(81),cout=>p(167)(82));
FA_ff_2514:FAff port map(x=>p(57)(82),y=>p(58)(82),Cin=>p(59)(82),clock=>clock,reset=>reset,s=>p(166)(82),cout=>p(167)(83));
FA_ff_2515:FAff port map(x=>p(57)(83),y=>p(58)(83),Cin=>p(59)(83),clock=>clock,reset=>reset,s=>p(166)(83),cout=>p(167)(84));
FA_ff_2516:FAff port map(x=>p(57)(84),y=>p(58)(84),Cin=>p(59)(84),clock=>clock,reset=>reset,s=>p(166)(84),cout=>p(167)(85));
FA_ff_2517:FAff port map(x=>p(57)(85),y=>p(58)(85),Cin=>p(59)(85),clock=>clock,reset=>reset,s=>p(166)(85),cout=>p(167)(86));
FA_ff_2518:FAff port map(x=>p(57)(86),y=>p(58)(86),Cin=>p(59)(86),clock=>clock,reset=>reset,s=>p(166)(86),cout=>p(167)(87));
FA_ff_2519:FAff port map(x=>p(57)(87),y=>p(58)(87),Cin=>p(59)(87),clock=>clock,reset=>reset,s=>p(166)(87),cout=>p(167)(88));
FA_ff_2520:FAff port map(x=>p(57)(88),y=>p(58)(88),Cin=>p(59)(88),clock=>clock,reset=>reset,s=>p(166)(88),cout=>p(167)(89));
FA_ff_2521:FAff port map(x=>p(57)(89),y=>p(58)(89),Cin=>p(59)(89),clock=>clock,reset=>reset,s=>p(166)(89),cout=>p(167)(90));
FA_ff_2522:FAff port map(x=>p(57)(90),y=>p(58)(90),Cin=>p(59)(90),clock=>clock,reset=>reset,s=>p(166)(90),cout=>p(167)(91));
FA_ff_2523:FAff port map(x=>p(57)(91),y=>p(58)(91),Cin=>p(59)(91),clock=>clock,reset=>reset,s=>p(166)(91),cout=>p(167)(92));
FA_ff_2524:FAff port map(x=>p(57)(92),y=>p(58)(92),Cin=>p(59)(92),clock=>clock,reset=>reset,s=>p(166)(92),cout=>p(167)(93));
FA_ff_2525:FAff port map(x=>p(57)(93),y=>p(58)(93),Cin=>p(59)(93),clock=>clock,reset=>reset,s=>p(166)(93),cout=>p(167)(94));
FA_ff_2526:FAff port map(x=>p(57)(94),y=>p(58)(94),Cin=>p(59)(94),clock=>clock,reset=>reset,s=>p(166)(94),cout=>p(167)(95));
FA_ff_2527:FAff port map(x=>p(57)(95),y=>p(58)(95),Cin=>p(59)(95),clock=>clock,reset=>reset,s=>p(166)(95),cout=>p(167)(96));
FA_ff_2528:FAff port map(x=>p(57)(96),y=>p(58)(96),Cin=>p(59)(96),clock=>clock,reset=>reset,s=>p(166)(96),cout=>p(167)(97));
FA_ff_2529:FAff port map(x=>p(57)(97),y=>p(58)(97),Cin=>p(59)(97),clock=>clock,reset=>reset,s=>p(166)(97),cout=>p(167)(98));
FA_ff_2530:FAff port map(x=>p(57)(98),y=>p(58)(98),Cin=>p(59)(98),clock=>clock,reset=>reset,s=>p(166)(98),cout=>p(167)(99));
FA_ff_2531:FAff port map(x=>p(57)(99),y=>p(58)(99),Cin=>p(59)(99),clock=>clock,reset=>reset,s=>p(166)(99),cout=>p(167)(100));
FA_ff_2532:FAff port map(x=>p(57)(100),y=>p(58)(100),Cin=>p(59)(100),clock=>clock,reset=>reset,s=>p(166)(100),cout=>p(167)(101));
FA_ff_2533:FAff port map(x=>p(57)(101),y=>p(58)(101),Cin=>p(59)(101),clock=>clock,reset=>reset,s=>p(166)(101),cout=>p(167)(102));
FA_ff_2534:FAff port map(x=>p(57)(102),y=>p(58)(102),Cin=>p(59)(102),clock=>clock,reset=>reset,s=>p(166)(102),cout=>p(167)(103));
FA_ff_2535:FAff port map(x=>p(57)(103),y=>p(58)(103),Cin=>p(59)(103),clock=>clock,reset=>reset,s=>p(166)(103),cout=>p(167)(104));
FA_ff_2536:FAff port map(x=>p(57)(104),y=>p(58)(104),Cin=>p(59)(104),clock=>clock,reset=>reset,s=>p(166)(104),cout=>p(167)(105));
FA_ff_2537:FAff port map(x=>p(57)(105),y=>p(58)(105),Cin=>p(59)(105),clock=>clock,reset=>reset,s=>p(166)(105),cout=>p(167)(106));
FA_ff_2538:FAff port map(x=>p(57)(106),y=>p(58)(106),Cin=>p(59)(106),clock=>clock,reset=>reset,s=>p(166)(106),cout=>p(167)(107));
FA_ff_2539:FAff port map(x=>p(57)(107),y=>p(58)(107),Cin=>p(59)(107),clock=>clock,reset=>reset,s=>p(166)(107),cout=>p(167)(108));
FA_ff_2540:FAff port map(x=>p(57)(108),y=>p(58)(108),Cin=>p(59)(108),clock=>clock,reset=>reset,s=>p(166)(108),cout=>p(167)(109));
FA_ff_2541:FAff port map(x=>p(57)(109),y=>p(58)(109),Cin=>p(59)(109),clock=>clock,reset=>reset,s=>p(166)(109),cout=>p(167)(110));
FA_ff_2542:FAff port map(x=>p(57)(110),y=>p(58)(110),Cin=>p(59)(110),clock=>clock,reset=>reset,s=>p(166)(110),cout=>p(167)(111));
FA_ff_2543:FAff port map(x=>p(57)(111),y=>p(58)(111),Cin=>p(59)(111),clock=>clock,reset=>reset,s=>p(166)(111),cout=>p(167)(112));
FA_ff_2544:FAff port map(x=>p(57)(112),y=>p(58)(112),Cin=>p(59)(112),clock=>clock,reset=>reset,s=>p(166)(112),cout=>p(167)(113));
FA_ff_2545:FAff port map(x=>p(57)(113),y=>p(58)(113),Cin=>p(59)(113),clock=>clock,reset=>reset,s=>p(166)(113),cout=>p(167)(114));
FA_ff_2546:FAff port map(x=>p(57)(114),y=>p(58)(114),Cin=>p(59)(114),clock=>clock,reset=>reset,s=>p(166)(114),cout=>p(167)(115));
FA_ff_2547:FAff port map(x=>p(57)(115),y=>p(58)(115),Cin=>p(59)(115),clock=>clock,reset=>reset,s=>p(166)(115),cout=>p(167)(116));
FA_ff_2548:FAff port map(x=>p(57)(116),y=>p(58)(116),Cin=>p(59)(116),clock=>clock,reset=>reset,s=>p(166)(116),cout=>p(167)(117));
FA_ff_2549:FAff port map(x=>p(57)(117),y=>p(58)(117),Cin=>p(59)(117),clock=>clock,reset=>reset,s=>p(166)(117),cout=>p(167)(118));
FA_ff_2550:FAff port map(x=>p(57)(118),y=>p(58)(118),Cin=>p(59)(118),clock=>clock,reset=>reset,s=>p(166)(118),cout=>p(167)(119));
FA_ff_2551:FAff port map(x=>p(57)(119),y=>p(58)(119),Cin=>p(59)(119),clock=>clock,reset=>reset,s=>p(166)(119),cout=>p(167)(120));
FA_ff_2552:FAff port map(x=>p(57)(120),y=>p(58)(120),Cin=>p(59)(120),clock=>clock,reset=>reset,s=>p(166)(120),cout=>p(167)(121));
FA_ff_2553:FAff port map(x=>p(57)(121),y=>p(58)(121),Cin=>p(59)(121),clock=>clock,reset=>reset,s=>p(166)(121),cout=>p(167)(122));
FA_ff_2554:FAff port map(x=>p(57)(122),y=>p(58)(122),Cin=>p(59)(122),clock=>clock,reset=>reset,s=>p(166)(122),cout=>p(167)(123));
FA_ff_2555:FAff port map(x=>p(57)(123),y=>p(58)(123),Cin=>p(59)(123),clock=>clock,reset=>reset,s=>p(166)(123),cout=>p(167)(124));
FA_ff_2556:FAff port map(x=>p(57)(124),y=>p(58)(124),Cin=>p(59)(124),clock=>clock,reset=>reset,s=>p(166)(124),cout=>p(167)(125));
FA_ff_2557:FAff port map(x=>p(57)(125),y=>p(58)(125),Cin=>p(59)(125),clock=>clock,reset=>reset,s=>p(166)(125),cout=>p(167)(126));
FA_ff_2558:FAff port map(x=>p(57)(126),y=>p(58)(126),Cin=>p(59)(126),clock=>clock,reset=>reset,s=>p(166)(126),cout=>p(167)(127));
FA_ff_2559:FAff port map(x=>p(57)(127),y=>p(58)(127),Cin=>p(59)(127),clock=>clock,reset=>reset,s=>p(166)(127),cout=>p(167)(128));
FA_ff_2560:FAff port map(x=>p(60)(0),y=>p(61)(0),Cin=>p(62)(0),clock=>clock,reset=>reset,s=>p(168)(0),cout=>p(169)(1));
FA_ff_2561:FAff port map(x=>p(60)(1),y=>p(61)(1),Cin=>p(62)(1),clock=>clock,reset=>reset,s=>p(168)(1),cout=>p(169)(2));
FA_ff_2562:FAff port map(x=>p(60)(2),y=>p(61)(2),Cin=>p(62)(2),clock=>clock,reset=>reset,s=>p(168)(2),cout=>p(169)(3));
FA_ff_2563:FAff port map(x=>p(60)(3),y=>p(61)(3),Cin=>p(62)(3),clock=>clock,reset=>reset,s=>p(168)(3),cout=>p(169)(4));
FA_ff_2564:FAff port map(x=>p(60)(4),y=>p(61)(4),Cin=>p(62)(4),clock=>clock,reset=>reset,s=>p(168)(4),cout=>p(169)(5));
FA_ff_2565:FAff port map(x=>p(60)(5),y=>p(61)(5),Cin=>p(62)(5),clock=>clock,reset=>reset,s=>p(168)(5),cout=>p(169)(6));
FA_ff_2566:FAff port map(x=>p(60)(6),y=>p(61)(6),Cin=>p(62)(6),clock=>clock,reset=>reset,s=>p(168)(6),cout=>p(169)(7));
FA_ff_2567:FAff port map(x=>p(60)(7),y=>p(61)(7),Cin=>p(62)(7),clock=>clock,reset=>reset,s=>p(168)(7),cout=>p(169)(8));
FA_ff_2568:FAff port map(x=>p(60)(8),y=>p(61)(8),Cin=>p(62)(8),clock=>clock,reset=>reset,s=>p(168)(8),cout=>p(169)(9));
FA_ff_2569:FAff port map(x=>p(60)(9),y=>p(61)(9),Cin=>p(62)(9),clock=>clock,reset=>reset,s=>p(168)(9),cout=>p(169)(10));
FA_ff_2570:FAff port map(x=>p(60)(10),y=>p(61)(10),Cin=>p(62)(10),clock=>clock,reset=>reset,s=>p(168)(10),cout=>p(169)(11));
FA_ff_2571:FAff port map(x=>p(60)(11),y=>p(61)(11),Cin=>p(62)(11),clock=>clock,reset=>reset,s=>p(168)(11),cout=>p(169)(12));
FA_ff_2572:FAff port map(x=>p(60)(12),y=>p(61)(12),Cin=>p(62)(12),clock=>clock,reset=>reset,s=>p(168)(12),cout=>p(169)(13));
FA_ff_2573:FAff port map(x=>p(60)(13),y=>p(61)(13),Cin=>p(62)(13),clock=>clock,reset=>reset,s=>p(168)(13),cout=>p(169)(14));
FA_ff_2574:FAff port map(x=>p(60)(14),y=>p(61)(14),Cin=>p(62)(14),clock=>clock,reset=>reset,s=>p(168)(14),cout=>p(169)(15));
FA_ff_2575:FAff port map(x=>p(60)(15),y=>p(61)(15),Cin=>p(62)(15),clock=>clock,reset=>reset,s=>p(168)(15),cout=>p(169)(16));
FA_ff_2576:FAff port map(x=>p(60)(16),y=>p(61)(16),Cin=>p(62)(16),clock=>clock,reset=>reset,s=>p(168)(16),cout=>p(169)(17));
FA_ff_2577:FAff port map(x=>p(60)(17),y=>p(61)(17),Cin=>p(62)(17),clock=>clock,reset=>reset,s=>p(168)(17),cout=>p(169)(18));
FA_ff_2578:FAff port map(x=>p(60)(18),y=>p(61)(18),Cin=>p(62)(18),clock=>clock,reset=>reset,s=>p(168)(18),cout=>p(169)(19));
FA_ff_2579:FAff port map(x=>p(60)(19),y=>p(61)(19),Cin=>p(62)(19),clock=>clock,reset=>reset,s=>p(168)(19),cout=>p(169)(20));
FA_ff_2580:FAff port map(x=>p(60)(20),y=>p(61)(20),Cin=>p(62)(20),clock=>clock,reset=>reset,s=>p(168)(20),cout=>p(169)(21));
FA_ff_2581:FAff port map(x=>p(60)(21),y=>p(61)(21),Cin=>p(62)(21),clock=>clock,reset=>reset,s=>p(168)(21),cout=>p(169)(22));
FA_ff_2582:FAff port map(x=>p(60)(22),y=>p(61)(22),Cin=>p(62)(22),clock=>clock,reset=>reset,s=>p(168)(22),cout=>p(169)(23));
FA_ff_2583:FAff port map(x=>p(60)(23),y=>p(61)(23),Cin=>p(62)(23),clock=>clock,reset=>reset,s=>p(168)(23),cout=>p(169)(24));
FA_ff_2584:FAff port map(x=>p(60)(24),y=>p(61)(24),Cin=>p(62)(24),clock=>clock,reset=>reset,s=>p(168)(24),cout=>p(169)(25));
FA_ff_2585:FAff port map(x=>p(60)(25),y=>p(61)(25),Cin=>p(62)(25),clock=>clock,reset=>reset,s=>p(168)(25),cout=>p(169)(26));
FA_ff_2586:FAff port map(x=>p(60)(26),y=>p(61)(26),Cin=>p(62)(26),clock=>clock,reset=>reset,s=>p(168)(26),cout=>p(169)(27));
FA_ff_2587:FAff port map(x=>p(60)(27),y=>p(61)(27),Cin=>p(62)(27),clock=>clock,reset=>reset,s=>p(168)(27),cout=>p(169)(28));
FA_ff_2588:FAff port map(x=>p(60)(28),y=>p(61)(28),Cin=>p(62)(28),clock=>clock,reset=>reset,s=>p(168)(28),cout=>p(169)(29));
FA_ff_2589:FAff port map(x=>p(60)(29),y=>p(61)(29),Cin=>p(62)(29),clock=>clock,reset=>reset,s=>p(168)(29),cout=>p(169)(30));
FA_ff_2590:FAff port map(x=>p(60)(30),y=>p(61)(30),Cin=>p(62)(30),clock=>clock,reset=>reset,s=>p(168)(30),cout=>p(169)(31));
FA_ff_2591:FAff port map(x=>p(60)(31),y=>p(61)(31),Cin=>p(62)(31),clock=>clock,reset=>reset,s=>p(168)(31),cout=>p(169)(32));
FA_ff_2592:FAff port map(x=>p(60)(32),y=>p(61)(32),Cin=>p(62)(32),clock=>clock,reset=>reset,s=>p(168)(32),cout=>p(169)(33));
FA_ff_2593:FAff port map(x=>p(60)(33),y=>p(61)(33),Cin=>p(62)(33),clock=>clock,reset=>reset,s=>p(168)(33),cout=>p(169)(34));
FA_ff_2594:FAff port map(x=>p(60)(34),y=>p(61)(34),Cin=>p(62)(34),clock=>clock,reset=>reset,s=>p(168)(34),cout=>p(169)(35));
FA_ff_2595:FAff port map(x=>p(60)(35),y=>p(61)(35),Cin=>p(62)(35),clock=>clock,reset=>reset,s=>p(168)(35),cout=>p(169)(36));
FA_ff_2596:FAff port map(x=>p(60)(36),y=>p(61)(36),Cin=>p(62)(36),clock=>clock,reset=>reset,s=>p(168)(36),cout=>p(169)(37));
FA_ff_2597:FAff port map(x=>p(60)(37),y=>p(61)(37),Cin=>p(62)(37),clock=>clock,reset=>reset,s=>p(168)(37),cout=>p(169)(38));
FA_ff_2598:FAff port map(x=>p(60)(38),y=>p(61)(38),Cin=>p(62)(38),clock=>clock,reset=>reset,s=>p(168)(38),cout=>p(169)(39));
FA_ff_2599:FAff port map(x=>p(60)(39),y=>p(61)(39),Cin=>p(62)(39),clock=>clock,reset=>reset,s=>p(168)(39),cout=>p(169)(40));
FA_ff_2600:FAff port map(x=>p(60)(40),y=>p(61)(40),Cin=>p(62)(40),clock=>clock,reset=>reset,s=>p(168)(40),cout=>p(169)(41));
FA_ff_2601:FAff port map(x=>p(60)(41),y=>p(61)(41),Cin=>p(62)(41),clock=>clock,reset=>reset,s=>p(168)(41),cout=>p(169)(42));
FA_ff_2602:FAff port map(x=>p(60)(42),y=>p(61)(42),Cin=>p(62)(42),clock=>clock,reset=>reset,s=>p(168)(42),cout=>p(169)(43));
FA_ff_2603:FAff port map(x=>p(60)(43),y=>p(61)(43),Cin=>p(62)(43),clock=>clock,reset=>reset,s=>p(168)(43),cout=>p(169)(44));
FA_ff_2604:FAff port map(x=>p(60)(44),y=>p(61)(44),Cin=>p(62)(44),clock=>clock,reset=>reset,s=>p(168)(44),cout=>p(169)(45));
FA_ff_2605:FAff port map(x=>p(60)(45),y=>p(61)(45),Cin=>p(62)(45),clock=>clock,reset=>reset,s=>p(168)(45),cout=>p(169)(46));
FA_ff_2606:FAff port map(x=>p(60)(46),y=>p(61)(46),Cin=>p(62)(46),clock=>clock,reset=>reset,s=>p(168)(46),cout=>p(169)(47));
FA_ff_2607:FAff port map(x=>p(60)(47),y=>p(61)(47),Cin=>p(62)(47),clock=>clock,reset=>reset,s=>p(168)(47),cout=>p(169)(48));
FA_ff_2608:FAff port map(x=>p(60)(48),y=>p(61)(48),Cin=>p(62)(48),clock=>clock,reset=>reset,s=>p(168)(48),cout=>p(169)(49));
FA_ff_2609:FAff port map(x=>p(60)(49),y=>p(61)(49),Cin=>p(62)(49),clock=>clock,reset=>reset,s=>p(168)(49),cout=>p(169)(50));
FA_ff_2610:FAff port map(x=>p(60)(50),y=>p(61)(50),Cin=>p(62)(50),clock=>clock,reset=>reset,s=>p(168)(50),cout=>p(169)(51));
FA_ff_2611:FAff port map(x=>p(60)(51),y=>p(61)(51),Cin=>p(62)(51),clock=>clock,reset=>reset,s=>p(168)(51),cout=>p(169)(52));
FA_ff_2612:FAff port map(x=>p(60)(52),y=>p(61)(52),Cin=>p(62)(52),clock=>clock,reset=>reset,s=>p(168)(52),cout=>p(169)(53));
FA_ff_2613:FAff port map(x=>p(60)(53),y=>p(61)(53),Cin=>p(62)(53),clock=>clock,reset=>reset,s=>p(168)(53),cout=>p(169)(54));
FA_ff_2614:FAff port map(x=>p(60)(54),y=>p(61)(54),Cin=>p(62)(54),clock=>clock,reset=>reset,s=>p(168)(54),cout=>p(169)(55));
FA_ff_2615:FAff port map(x=>p(60)(55),y=>p(61)(55),Cin=>p(62)(55),clock=>clock,reset=>reset,s=>p(168)(55),cout=>p(169)(56));
FA_ff_2616:FAff port map(x=>p(60)(56),y=>p(61)(56),Cin=>p(62)(56),clock=>clock,reset=>reset,s=>p(168)(56),cout=>p(169)(57));
FA_ff_2617:FAff port map(x=>p(60)(57),y=>p(61)(57),Cin=>p(62)(57),clock=>clock,reset=>reset,s=>p(168)(57),cout=>p(169)(58));
FA_ff_2618:FAff port map(x=>p(60)(58),y=>p(61)(58),Cin=>p(62)(58),clock=>clock,reset=>reset,s=>p(168)(58),cout=>p(169)(59));
FA_ff_2619:FAff port map(x=>p(60)(59),y=>p(61)(59),Cin=>p(62)(59),clock=>clock,reset=>reset,s=>p(168)(59),cout=>p(169)(60));
FA_ff_2620:FAff port map(x=>p(60)(60),y=>p(61)(60),Cin=>p(62)(60),clock=>clock,reset=>reset,s=>p(168)(60),cout=>p(169)(61));
FA_ff_2621:FAff port map(x=>p(60)(61),y=>p(61)(61),Cin=>p(62)(61),clock=>clock,reset=>reset,s=>p(168)(61),cout=>p(169)(62));
FA_ff_2622:FAff port map(x=>p(60)(62),y=>p(61)(62),Cin=>p(62)(62),clock=>clock,reset=>reset,s=>p(168)(62),cout=>p(169)(63));
FA_ff_2623:FAff port map(x=>p(60)(63),y=>p(61)(63),Cin=>p(62)(63),clock=>clock,reset=>reset,s=>p(168)(63),cout=>p(169)(64));
FA_ff_2624:FAff port map(x=>p(60)(64),y=>p(61)(64),Cin=>p(62)(64),clock=>clock,reset=>reset,s=>p(168)(64),cout=>p(169)(65));
FA_ff_2625:FAff port map(x=>p(60)(65),y=>p(61)(65),Cin=>p(62)(65),clock=>clock,reset=>reset,s=>p(168)(65),cout=>p(169)(66));
FA_ff_2626:FAff port map(x=>p(60)(66),y=>p(61)(66),Cin=>p(62)(66),clock=>clock,reset=>reset,s=>p(168)(66),cout=>p(169)(67));
FA_ff_2627:FAff port map(x=>p(60)(67),y=>p(61)(67),Cin=>p(62)(67),clock=>clock,reset=>reset,s=>p(168)(67),cout=>p(169)(68));
FA_ff_2628:FAff port map(x=>p(60)(68),y=>p(61)(68),Cin=>p(62)(68),clock=>clock,reset=>reset,s=>p(168)(68),cout=>p(169)(69));
FA_ff_2629:FAff port map(x=>p(60)(69),y=>p(61)(69),Cin=>p(62)(69),clock=>clock,reset=>reset,s=>p(168)(69),cout=>p(169)(70));
FA_ff_2630:FAff port map(x=>p(60)(70),y=>p(61)(70),Cin=>p(62)(70),clock=>clock,reset=>reset,s=>p(168)(70),cout=>p(169)(71));
FA_ff_2631:FAff port map(x=>p(60)(71),y=>p(61)(71),Cin=>p(62)(71),clock=>clock,reset=>reset,s=>p(168)(71),cout=>p(169)(72));
FA_ff_2632:FAff port map(x=>p(60)(72),y=>p(61)(72),Cin=>p(62)(72),clock=>clock,reset=>reset,s=>p(168)(72),cout=>p(169)(73));
FA_ff_2633:FAff port map(x=>p(60)(73),y=>p(61)(73),Cin=>p(62)(73),clock=>clock,reset=>reset,s=>p(168)(73),cout=>p(169)(74));
FA_ff_2634:FAff port map(x=>p(60)(74),y=>p(61)(74),Cin=>p(62)(74),clock=>clock,reset=>reset,s=>p(168)(74),cout=>p(169)(75));
FA_ff_2635:FAff port map(x=>p(60)(75),y=>p(61)(75),Cin=>p(62)(75),clock=>clock,reset=>reset,s=>p(168)(75),cout=>p(169)(76));
FA_ff_2636:FAff port map(x=>p(60)(76),y=>p(61)(76),Cin=>p(62)(76),clock=>clock,reset=>reset,s=>p(168)(76),cout=>p(169)(77));
FA_ff_2637:FAff port map(x=>p(60)(77),y=>p(61)(77),Cin=>p(62)(77),clock=>clock,reset=>reset,s=>p(168)(77),cout=>p(169)(78));
FA_ff_2638:FAff port map(x=>p(60)(78),y=>p(61)(78),Cin=>p(62)(78),clock=>clock,reset=>reset,s=>p(168)(78),cout=>p(169)(79));
FA_ff_2639:FAff port map(x=>p(60)(79),y=>p(61)(79),Cin=>p(62)(79),clock=>clock,reset=>reset,s=>p(168)(79),cout=>p(169)(80));
FA_ff_2640:FAff port map(x=>p(60)(80),y=>p(61)(80),Cin=>p(62)(80),clock=>clock,reset=>reset,s=>p(168)(80),cout=>p(169)(81));
FA_ff_2641:FAff port map(x=>p(60)(81),y=>p(61)(81),Cin=>p(62)(81),clock=>clock,reset=>reset,s=>p(168)(81),cout=>p(169)(82));
FA_ff_2642:FAff port map(x=>p(60)(82),y=>p(61)(82),Cin=>p(62)(82),clock=>clock,reset=>reset,s=>p(168)(82),cout=>p(169)(83));
FA_ff_2643:FAff port map(x=>p(60)(83),y=>p(61)(83),Cin=>p(62)(83),clock=>clock,reset=>reset,s=>p(168)(83),cout=>p(169)(84));
FA_ff_2644:FAff port map(x=>p(60)(84),y=>p(61)(84),Cin=>p(62)(84),clock=>clock,reset=>reset,s=>p(168)(84),cout=>p(169)(85));
FA_ff_2645:FAff port map(x=>p(60)(85),y=>p(61)(85),Cin=>p(62)(85),clock=>clock,reset=>reset,s=>p(168)(85),cout=>p(169)(86));
FA_ff_2646:FAff port map(x=>p(60)(86),y=>p(61)(86),Cin=>p(62)(86),clock=>clock,reset=>reset,s=>p(168)(86),cout=>p(169)(87));
FA_ff_2647:FAff port map(x=>p(60)(87),y=>p(61)(87),Cin=>p(62)(87),clock=>clock,reset=>reset,s=>p(168)(87),cout=>p(169)(88));
FA_ff_2648:FAff port map(x=>p(60)(88),y=>p(61)(88),Cin=>p(62)(88),clock=>clock,reset=>reset,s=>p(168)(88),cout=>p(169)(89));
FA_ff_2649:FAff port map(x=>p(60)(89),y=>p(61)(89),Cin=>p(62)(89),clock=>clock,reset=>reset,s=>p(168)(89),cout=>p(169)(90));
FA_ff_2650:FAff port map(x=>p(60)(90),y=>p(61)(90),Cin=>p(62)(90),clock=>clock,reset=>reset,s=>p(168)(90),cout=>p(169)(91));
FA_ff_2651:FAff port map(x=>p(60)(91),y=>p(61)(91),Cin=>p(62)(91),clock=>clock,reset=>reset,s=>p(168)(91),cout=>p(169)(92));
FA_ff_2652:FAff port map(x=>p(60)(92),y=>p(61)(92),Cin=>p(62)(92),clock=>clock,reset=>reset,s=>p(168)(92),cout=>p(169)(93));
FA_ff_2653:FAff port map(x=>p(60)(93),y=>p(61)(93),Cin=>p(62)(93),clock=>clock,reset=>reset,s=>p(168)(93),cout=>p(169)(94));
FA_ff_2654:FAff port map(x=>p(60)(94),y=>p(61)(94),Cin=>p(62)(94),clock=>clock,reset=>reset,s=>p(168)(94),cout=>p(169)(95));
FA_ff_2655:FAff port map(x=>p(60)(95),y=>p(61)(95),Cin=>p(62)(95),clock=>clock,reset=>reset,s=>p(168)(95),cout=>p(169)(96));
FA_ff_2656:FAff port map(x=>p(60)(96),y=>p(61)(96),Cin=>p(62)(96),clock=>clock,reset=>reset,s=>p(168)(96),cout=>p(169)(97));
FA_ff_2657:FAff port map(x=>p(60)(97),y=>p(61)(97),Cin=>p(62)(97),clock=>clock,reset=>reset,s=>p(168)(97),cout=>p(169)(98));
FA_ff_2658:FAff port map(x=>p(60)(98),y=>p(61)(98),Cin=>p(62)(98),clock=>clock,reset=>reset,s=>p(168)(98),cout=>p(169)(99));
FA_ff_2659:FAff port map(x=>p(60)(99),y=>p(61)(99),Cin=>p(62)(99),clock=>clock,reset=>reset,s=>p(168)(99),cout=>p(169)(100));
FA_ff_2660:FAff port map(x=>p(60)(100),y=>p(61)(100),Cin=>p(62)(100),clock=>clock,reset=>reset,s=>p(168)(100),cout=>p(169)(101));
FA_ff_2661:FAff port map(x=>p(60)(101),y=>p(61)(101),Cin=>p(62)(101),clock=>clock,reset=>reset,s=>p(168)(101),cout=>p(169)(102));
FA_ff_2662:FAff port map(x=>p(60)(102),y=>p(61)(102),Cin=>p(62)(102),clock=>clock,reset=>reset,s=>p(168)(102),cout=>p(169)(103));
FA_ff_2663:FAff port map(x=>p(60)(103),y=>p(61)(103),Cin=>p(62)(103),clock=>clock,reset=>reset,s=>p(168)(103),cout=>p(169)(104));
FA_ff_2664:FAff port map(x=>p(60)(104),y=>p(61)(104),Cin=>p(62)(104),clock=>clock,reset=>reset,s=>p(168)(104),cout=>p(169)(105));
FA_ff_2665:FAff port map(x=>p(60)(105),y=>p(61)(105),Cin=>p(62)(105),clock=>clock,reset=>reset,s=>p(168)(105),cout=>p(169)(106));
FA_ff_2666:FAff port map(x=>p(60)(106),y=>p(61)(106),Cin=>p(62)(106),clock=>clock,reset=>reset,s=>p(168)(106),cout=>p(169)(107));
FA_ff_2667:FAff port map(x=>p(60)(107),y=>p(61)(107),Cin=>p(62)(107),clock=>clock,reset=>reset,s=>p(168)(107),cout=>p(169)(108));
FA_ff_2668:FAff port map(x=>p(60)(108),y=>p(61)(108),Cin=>p(62)(108),clock=>clock,reset=>reset,s=>p(168)(108),cout=>p(169)(109));
FA_ff_2669:FAff port map(x=>p(60)(109),y=>p(61)(109),Cin=>p(62)(109),clock=>clock,reset=>reset,s=>p(168)(109),cout=>p(169)(110));
FA_ff_2670:FAff port map(x=>p(60)(110),y=>p(61)(110),Cin=>p(62)(110),clock=>clock,reset=>reset,s=>p(168)(110),cout=>p(169)(111));
FA_ff_2671:FAff port map(x=>p(60)(111),y=>p(61)(111),Cin=>p(62)(111),clock=>clock,reset=>reset,s=>p(168)(111),cout=>p(169)(112));
FA_ff_2672:FAff port map(x=>p(60)(112),y=>p(61)(112),Cin=>p(62)(112),clock=>clock,reset=>reset,s=>p(168)(112),cout=>p(169)(113));
FA_ff_2673:FAff port map(x=>p(60)(113),y=>p(61)(113),Cin=>p(62)(113),clock=>clock,reset=>reset,s=>p(168)(113),cout=>p(169)(114));
FA_ff_2674:FAff port map(x=>p(60)(114),y=>p(61)(114),Cin=>p(62)(114),clock=>clock,reset=>reset,s=>p(168)(114),cout=>p(169)(115));
FA_ff_2675:FAff port map(x=>p(60)(115),y=>p(61)(115),Cin=>p(62)(115),clock=>clock,reset=>reset,s=>p(168)(115),cout=>p(169)(116));
FA_ff_2676:FAff port map(x=>p(60)(116),y=>p(61)(116),Cin=>p(62)(116),clock=>clock,reset=>reset,s=>p(168)(116),cout=>p(169)(117));
FA_ff_2677:FAff port map(x=>p(60)(117),y=>p(61)(117),Cin=>p(62)(117),clock=>clock,reset=>reset,s=>p(168)(117),cout=>p(169)(118));
FA_ff_2678:FAff port map(x=>p(60)(118),y=>p(61)(118),Cin=>p(62)(118),clock=>clock,reset=>reset,s=>p(168)(118),cout=>p(169)(119));
FA_ff_2679:FAff port map(x=>p(60)(119),y=>p(61)(119),Cin=>p(62)(119),clock=>clock,reset=>reset,s=>p(168)(119),cout=>p(169)(120));
FA_ff_2680:FAff port map(x=>p(60)(120),y=>p(61)(120),Cin=>p(62)(120),clock=>clock,reset=>reset,s=>p(168)(120),cout=>p(169)(121));
FA_ff_2681:FAff port map(x=>p(60)(121),y=>p(61)(121),Cin=>p(62)(121),clock=>clock,reset=>reset,s=>p(168)(121),cout=>p(169)(122));
FA_ff_2682:FAff port map(x=>p(60)(122),y=>p(61)(122),Cin=>p(62)(122),clock=>clock,reset=>reset,s=>p(168)(122),cout=>p(169)(123));
FA_ff_2683:FAff port map(x=>p(60)(123),y=>p(61)(123),Cin=>p(62)(123),clock=>clock,reset=>reset,s=>p(168)(123),cout=>p(169)(124));
FA_ff_2684:FAff port map(x=>p(60)(124),y=>p(61)(124),Cin=>p(62)(124),clock=>clock,reset=>reset,s=>p(168)(124),cout=>p(169)(125));
FA_ff_2685:FAff port map(x=>p(60)(125),y=>p(61)(125),Cin=>p(62)(125),clock=>clock,reset=>reset,s=>p(168)(125),cout=>p(169)(126));
FA_ff_2686:FAff port map(x=>p(60)(126),y=>p(61)(126),Cin=>p(62)(126),clock=>clock,reset=>reset,s=>p(168)(126),cout=>p(169)(127));
FA_ff_2687:FAff port map(x=>p(60)(127),y=>p(61)(127),Cin=>p(62)(127),clock=>clock,reset=>reset,s=>p(168)(127),cout=>p(169)(128));
FA_ff_2688:FAff port map(x=>p(63)(0),y=>p(64)(0),Cin=>p(65)(0),clock=>clock,reset=>reset,s=>p(170)(0),cout=>p(171)(1));
FA_ff_2689:FAff port map(x=>p(63)(1),y=>p(64)(1),Cin=>p(65)(1),clock=>clock,reset=>reset,s=>p(170)(1),cout=>p(171)(2));
FA_ff_2690:FAff port map(x=>p(63)(2),y=>p(64)(2),Cin=>p(65)(2),clock=>clock,reset=>reset,s=>p(170)(2),cout=>p(171)(3));
FA_ff_2691:FAff port map(x=>p(63)(3),y=>p(64)(3),Cin=>p(65)(3),clock=>clock,reset=>reset,s=>p(170)(3),cout=>p(171)(4));
FA_ff_2692:FAff port map(x=>p(63)(4),y=>p(64)(4),Cin=>p(65)(4),clock=>clock,reset=>reset,s=>p(170)(4),cout=>p(171)(5));
FA_ff_2693:FAff port map(x=>p(63)(5),y=>p(64)(5),Cin=>p(65)(5),clock=>clock,reset=>reset,s=>p(170)(5),cout=>p(171)(6));
FA_ff_2694:FAff port map(x=>p(63)(6),y=>p(64)(6),Cin=>p(65)(6),clock=>clock,reset=>reset,s=>p(170)(6),cout=>p(171)(7));
FA_ff_2695:FAff port map(x=>p(63)(7),y=>p(64)(7),Cin=>p(65)(7),clock=>clock,reset=>reset,s=>p(170)(7),cout=>p(171)(8));
FA_ff_2696:FAff port map(x=>p(63)(8),y=>p(64)(8),Cin=>p(65)(8),clock=>clock,reset=>reset,s=>p(170)(8),cout=>p(171)(9));
FA_ff_2697:FAff port map(x=>p(63)(9),y=>p(64)(9),Cin=>p(65)(9),clock=>clock,reset=>reset,s=>p(170)(9),cout=>p(171)(10));
FA_ff_2698:FAff port map(x=>p(63)(10),y=>p(64)(10),Cin=>p(65)(10),clock=>clock,reset=>reset,s=>p(170)(10),cout=>p(171)(11));
FA_ff_2699:FAff port map(x=>p(63)(11),y=>p(64)(11),Cin=>p(65)(11),clock=>clock,reset=>reset,s=>p(170)(11),cout=>p(171)(12));
FA_ff_2700:FAff port map(x=>p(63)(12),y=>p(64)(12),Cin=>p(65)(12),clock=>clock,reset=>reset,s=>p(170)(12),cout=>p(171)(13));
FA_ff_2701:FAff port map(x=>p(63)(13),y=>p(64)(13),Cin=>p(65)(13),clock=>clock,reset=>reset,s=>p(170)(13),cout=>p(171)(14));
FA_ff_2702:FAff port map(x=>p(63)(14),y=>p(64)(14),Cin=>p(65)(14),clock=>clock,reset=>reset,s=>p(170)(14),cout=>p(171)(15));
FA_ff_2703:FAff port map(x=>p(63)(15),y=>p(64)(15),Cin=>p(65)(15),clock=>clock,reset=>reset,s=>p(170)(15),cout=>p(171)(16));
FA_ff_2704:FAff port map(x=>p(63)(16),y=>p(64)(16),Cin=>p(65)(16),clock=>clock,reset=>reset,s=>p(170)(16),cout=>p(171)(17));
FA_ff_2705:FAff port map(x=>p(63)(17),y=>p(64)(17),Cin=>p(65)(17),clock=>clock,reset=>reset,s=>p(170)(17),cout=>p(171)(18));
FA_ff_2706:FAff port map(x=>p(63)(18),y=>p(64)(18),Cin=>p(65)(18),clock=>clock,reset=>reset,s=>p(170)(18),cout=>p(171)(19));
FA_ff_2707:FAff port map(x=>p(63)(19),y=>p(64)(19),Cin=>p(65)(19),clock=>clock,reset=>reset,s=>p(170)(19),cout=>p(171)(20));
FA_ff_2708:FAff port map(x=>p(63)(20),y=>p(64)(20),Cin=>p(65)(20),clock=>clock,reset=>reset,s=>p(170)(20),cout=>p(171)(21));
FA_ff_2709:FAff port map(x=>p(63)(21),y=>p(64)(21),Cin=>p(65)(21),clock=>clock,reset=>reset,s=>p(170)(21),cout=>p(171)(22));
FA_ff_2710:FAff port map(x=>p(63)(22),y=>p(64)(22),Cin=>p(65)(22),clock=>clock,reset=>reset,s=>p(170)(22),cout=>p(171)(23));
FA_ff_2711:FAff port map(x=>p(63)(23),y=>p(64)(23),Cin=>p(65)(23),clock=>clock,reset=>reset,s=>p(170)(23),cout=>p(171)(24));
FA_ff_2712:FAff port map(x=>p(63)(24),y=>p(64)(24),Cin=>p(65)(24),clock=>clock,reset=>reset,s=>p(170)(24),cout=>p(171)(25));
FA_ff_2713:FAff port map(x=>p(63)(25),y=>p(64)(25),Cin=>p(65)(25),clock=>clock,reset=>reset,s=>p(170)(25),cout=>p(171)(26));
FA_ff_2714:FAff port map(x=>p(63)(26),y=>p(64)(26),Cin=>p(65)(26),clock=>clock,reset=>reset,s=>p(170)(26),cout=>p(171)(27));
FA_ff_2715:FAff port map(x=>p(63)(27),y=>p(64)(27),Cin=>p(65)(27),clock=>clock,reset=>reset,s=>p(170)(27),cout=>p(171)(28));
FA_ff_2716:FAff port map(x=>p(63)(28),y=>p(64)(28),Cin=>p(65)(28),clock=>clock,reset=>reset,s=>p(170)(28),cout=>p(171)(29));
FA_ff_2717:FAff port map(x=>p(63)(29),y=>p(64)(29),Cin=>p(65)(29),clock=>clock,reset=>reset,s=>p(170)(29),cout=>p(171)(30));
FA_ff_2718:FAff port map(x=>p(63)(30),y=>p(64)(30),Cin=>p(65)(30),clock=>clock,reset=>reset,s=>p(170)(30),cout=>p(171)(31));
FA_ff_2719:FAff port map(x=>p(63)(31),y=>p(64)(31),Cin=>p(65)(31),clock=>clock,reset=>reset,s=>p(170)(31),cout=>p(171)(32));
FA_ff_2720:FAff port map(x=>p(63)(32),y=>p(64)(32),Cin=>p(65)(32),clock=>clock,reset=>reset,s=>p(170)(32),cout=>p(171)(33));
FA_ff_2721:FAff port map(x=>p(63)(33),y=>p(64)(33),Cin=>p(65)(33),clock=>clock,reset=>reset,s=>p(170)(33),cout=>p(171)(34));
FA_ff_2722:FAff port map(x=>p(63)(34),y=>p(64)(34),Cin=>p(65)(34),clock=>clock,reset=>reset,s=>p(170)(34),cout=>p(171)(35));
FA_ff_2723:FAff port map(x=>p(63)(35),y=>p(64)(35),Cin=>p(65)(35),clock=>clock,reset=>reset,s=>p(170)(35),cout=>p(171)(36));
FA_ff_2724:FAff port map(x=>p(63)(36),y=>p(64)(36),Cin=>p(65)(36),clock=>clock,reset=>reset,s=>p(170)(36),cout=>p(171)(37));
FA_ff_2725:FAff port map(x=>p(63)(37),y=>p(64)(37),Cin=>p(65)(37),clock=>clock,reset=>reset,s=>p(170)(37),cout=>p(171)(38));
FA_ff_2726:FAff port map(x=>p(63)(38),y=>p(64)(38),Cin=>p(65)(38),clock=>clock,reset=>reset,s=>p(170)(38),cout=>p(171)(39));
FA_ff_2727:FAff port map(x=>p(63)(39),y=>p(64)(39),Cin=>p(65)(39),clock=>clock,reset=>reset,s=>p(170)(39),cout=>p(171)(40));
FA_ff_2728:FAff port map(x=>p(63)(40),y=>p(64)(40),Cin=>p(65)(40),clock=>clock,reset=>reset,s=>p(170)(40),cout=>p(171)(41));
FA_ff_2729:FAff port map(x=>p(63)(41),y=>p(64)(41),Cin=>p(65)(41),clock=>clock,reset=>reset,s=>p(170)(41),cout=>p(171)(42));
FA_ff_2730:FAff port map(x=>p(63)(42),y=>p(64)(42),Cin=>p(65)(42),clock=>clock,reset=>reset,s=>p(170)(42),cout=>p(171)(43));
FA_ff_2731:FAff port map(x=>p(63)(43),y=>p(64)(43),Cin=>p(65)(43),clock=>clock,reset=>reset,s=>p(170)(43),cout=>p(171)(44));
FA_ff_2732:FAff port map(x=>p(63)(44),y=>p(64)(44),Cin=>p(65)(44),clock=>clock,reset=>reset,s=>p(170)(44),cout=>p(171)(45));
FA_ff_2733:FAff port map(x=>p(63)(45),y=>p(64)(45),Cin=>p(65)(45),clock=>clock,reset=>reset,s=>p(170)(45),cout=>p(171)(46));
FA_ff_2734:FAff port map(x=>p(63)(46),y=>p(64)(46),Cin=>p(65)(46),clock=>clock,reset=>reset,s=>p(170)(46),cout=>p(171)(47));
FA_ff_2735:FAff port map(x=>p(63)(47),y=>p(64)(47),Cin=>p(65)(47),clock=>clock,reset=>reset,s=>p(170)(47),cout=>p(171)(48));
FA_ff_2736:FAff port map(x=>p(63)(48),y=>p(64)(48),Cin=>p(65)(48),clock=>clock,reset=>reset,s=>p(170)(48),cout=>p(171)(49));
FA_ff_2737:FAff port map(x=>p(63)(49),y=>p(64)(49),Cin=>p(65)(49),clock=>clock,reset=>reset,s=>p(170)(49),cout=>p(171)(50));
FA_ff_2738:FAff port map(x=>p(63)(50),y=>p(64)(50),Cin=>p(65)(50),clock=>clock,reset=>reset,s=>p(170)(50),cout=>p(171)(51));
FA_ff_2739:FAff port map(x=>p(63)(51),y=>p(64)(51),Cin=>p(65)(51),clock=>clock,reset=>reset,s=>p(170)(51),cout=>p(171)(52));
FA_ff_2740:FAff port map(x=>p(63)(52),y=>p(64)(52),Cin=>p(65)(52),clock=>clock,reset=>reset,s=>p(170)(52),cout=>p(171)(53));
FA_ff_2741:FAff port map(x=>p(63)(53),y=>p(64)(53),Cin=>p(65)(53),clock=>clock,reset=>reset,s=>p(170)(53),cout=>p(171)(54));
FA_ff_2742:FAff port map(x=>p(63)(54),y=>p(64)(54),Cin=>p(65)(54),clock=>clock,reset=>reset,s=>p(170)(54),cout=>p(171)(55));
FA_ff_2743:FAff port map(x=>p(63)(55),y=>p(64)(55),Cin=>p(65)(55),clock=>clock,reset=>reset,s=>p(170)(55),cout=>p(171)(56));
FA_ff_2744:FAff port map(x=>p(63)(56),y=>p(64)(56),Cin=>p(65)(56),clock=>clock,reset=>reset,s=>p(170)(56),cout=>p(171)(57));
FA_ff_2745:FAff port map(x=>p(63)(57),y=>p(64)(57),Cin=>p(65)(57),clock=>clock,reset=>reset,s=>p(170)(57),cout=>p(171)(58));
FA_ff_2746:FAff port map(x=>p(63)(58),y=>p(64)(58),Cin=>p(65)(58),clock=>clock,reset=>reset,s=>p(170)(58),cout=>p(171)(59));
FA_ff_2747:FAff port map(x=>p(63)(59),y=>p(64)(59),Cin=>p(65)(59),clock=>clock,reset=>reset,s=>p(170)(59),cout=>p(171)(60));
FA_ff_2748:FAff port map(x=>p(63)(60),y=>p(64)(60),Cin=>p(65)(60),clock=>clock,reset=>reset,s=>p(170)(60),cout=>p(171)(61));
FA_ff_2749:FAff port map(x=>p(63)(61),y=>p(64)(61),Cin=>p(65)(61),clock=>clock,reset=>reset,s=>p(170)(61),cout=>p(171)(62));
FA_ff_2750:FAff port map(x=>p(63)(62),y=>p(64)(62),Cin=>p(65)(62),clock=>clock,reset=>reset,s=>p(170)(62),cout=>p(171)(63));
FA_ff_2751:FAff port map(x=>p(63)(63),y=>p(64)(63),Cin=>p(65)(63),clock=>clock,reset=>reset,s=>p(170)(63),cout=>p(171)(64));
FA_ff_2752:FAff port map(x=>p(63)(64),y=>p(64)(64),Cin=>p(65)(64),clock=>clock,reset=>reset,s=>p(170)(64),cout=>p(171)(65));
FA_ff_2753:FAff port map(x=>p(63)(65),y=>p(64)(65),Cin=>p(65)(65),clock=>clock,reset=>reset,s=>p(170)(65),cout=>p(171)(66));
FA_ff_2754:FAff port map(x=>p(63)(66),y=>p(64)(66),Cin=>p(65)(66),clock=>clock,reset=>reset,s=>p(170)(66),cout=>p(171)(67));
FA_ff_2755:FAff port map(x=>p(63)(67),y=>p(64)(67),Cin=>p(65)(67),clock=>clock,reset=>reset,s=>p(170)(67),cout=>p(171)(68));
FA_ff_2756:FAff port map(x=>p(63)(68),y=>p(64)(68),Cin=>p(65)(68),clock=>clock,reset=>reset,s=>p(170)(68),cout=>p(171)(69));
FA_ff_2757:FAff port map(x=>p(63)(69),y=>p(64)(69),Cin=>p(65)(69),clock=>clock,reset=>reset,s=>p(170)(69),cout=>p(171)(70));
FA_ff_2758:FAff port map(x=>p(63)(70),y=>p(64)(70),Cin=>p(65)(70),clock=>clock,reset=>reset,s=>p(170)(70),cout=>p(171)(71));
FA_ff_2759:FAff port map(x=>p(63)(71),y=>p(64)(71),Cin=>p(65)(71),clock=>clock,reset=>reset,s=>p(170)(71),cout=>p(171)(72));
FA_ff_2760:FAff port map(x=>p(63)(72),y=>p(64)(72),Cin=>p(65)(72),clock=>clock,reset=>reset,s=>p(170)(72),cout=>p(171)(73));
FA_ff_2761:FAff port map(x=>p(63)(73),y=>p(64)(73),Cin=>p(65)(73),clock=>clock,reset=>reset,s=>p(170)(73),cout=>p(171)(74));
FA_ff_2762:FAff port map(x=>p(63)(74),y=>p(64)(74),Cin=>p(65)(74),clock=>clock,reset=>reset,s=>p(170)(74),cout=>p(171)(75));
FA_ff_2763:FAff port map(x=>p(63)(75),y=>p(64)(75),Cin=>p(65)(75),clock=>clock,reset=>reset,s=>p(170)(75),cout=>p(171)(76));
FA_ff_2764:FAff port map(x=>p(63)(76),y=>p(64)(76),Cin=>p(65)(76),clock=>clock,reset=>reset,s=>p(170)(76),cout=>p(171)(77));
FA_ff_2765:FAff port map(x=>p(63)(77),y=>p(64)(77),Cin=>p(65)(77),clock=>clock,reset=>reset,s=>p(170)(77),cout=>p(171)(78));
FA_ff_2766:FAff port map(x=>p(63)(78),y=>p(64)(78),Cin=>p(65)(78),clock=>clock,reset=>reset,s=>p(170)(78),cout=>p(171)(79));
FA_ff_2767:FAff port map(x=>p(63)(79),y=>p(64)(79),Cin=>p(65)(79),clock=>clock,reset=>reset,s=>p(170)(79),cout=>p(171)(80));
FA_ff_2768:FAff port map(x=>p(63)(80),y=>p(64)(80),Cin=>p(65)(80),clock=>clock,reset=>reset,s=>p(170)(80),cout=>p(171)(81));
FA_ff_2769:FAff port map(x=>p(63)(81),y=>p(64)(81),Cin=>p(65)(81),clock=>clock,reset=>reset,s=>p(170)(81),cout=>p(171)(82));
FA_ff_2770:FAff port map(x=>p(63)(82),y=>p(64)(82),Cin=>p(65)(82),clock=>clock,reset=>reset,s=>p(170)(82),cout=>p(171)(83));
FA_ff_2771:FAff port map(x=>p(63)(83),y=>p(64)(83),Cin=>p(65)(83),clock=>clock,reset=>reset,s=>p(170)(83),cout=>p(171)(84));
FA_ff_2772:FAff port map(x=>p(63)(84),y=>p(64)(84),Cin=>p(65)(84),clock=>clock,reset=>reset,s=>p(170)(84),cout=>p(171)(85));
FA_ff_2773:FAff port map(x=>p(63)(85),y=>p(64)(85),Cin=>p(65)(85),clock=>clock,reset=>reset,s=>p(170)(85),cout=>p(171)(86));
FA_ff_2774:FAff port map(x=>p(63)(86),y=>p(64)(86),Cin=>p(65)(86),clock=>clock,reset=>reset,s=>p(170)(86),cout=>p(171)(87));
FA_ff_2775:FAff port map(x=>p(63)(87),y=>p(64)(87),Cin=>p(65)(87),clock=>clock,reset=>reset,s=>p(170)(87),cout=>p(171)(88));
FA_ff_2776:FAff port map(x=>p(63)(88),y=>p(64)(88),Cin=>p(65)(88),clock=>clock,reset=>reset,s=>p(170)(88),cout=>p(171)(89));
FA_ff_2777:FAff port map(x=>p(63)(89),y=>p(64)(89),Cin=>p(65)(89),clock=>clock,reset=>reset,s=>p(170)(89),cout=>p(171)(90));
FA_ff_2778:FAff port map(x=>p(63)(90),y=>p(64)(90),Cin=>p(65)(90),clock=>clock,reset=>reset,s=>p(170)(90),cout=>p(171)(91));
FA_ff_2779:FAff port map(x=>p(63)(91),y=>p(64)(91),Cin=>p(65)(91),clock=>clock,reset=>reset,s=>p(170)(91),cout=>p(171)(92));
FA_ff_2780:FAff port map(x=>p(63)(92),y=>p(64)(92),Cin=>p(65)(92),clock=>clock,reset=>reset,s=>p(170)(92),cout=>p(171)(93));
FA_ff_2781:FAff port map(x=>p(63)(93),y=>p(64)(93),Cin=>p(65)(93),clock=>clock,reset=>reset,s=>p(170)(93),cout=>p(171)(94));
FA_ff_2782:FAff port map(x=>p(63)(94),y=>p(64)(94),Cin=>p(65)(94),clock=>clock,reset=>reset,s=>p(170)(94),cout=>p(171)(95));
FA_ff_2783:FAff port map(x=>p(63)(95),y=>p(64)(95),Cin=>p(65)(95),clock=>clock,reset=>reset,s=>p(170)(95),cout=>p(171)(96));
FA_ff_2784:FAff port map(x=>p(63)(96),y=>p(64)(96),Cin=>p(65)(96),clock=>clock,reset=>reset,s=>p(170)(96),cout=>p(171)(97));
FA_ff_2785:FAff port map(x=>p(63)(97),y=>p(64)(97),Cin=>p(65)(97),clock=>clock,reset=>reset,s=>p(170)(97),cout=>p(171)(98));
FA_ff_2786:FAff port map(x=>p(63)(98),y=>p(64)(98),Cin=>p(65)(98),clock=>clock,reset=>reset,s=>p(170)(98),cout=>p(171)(99));
FA_ff_2787:FAff port map(x=>p(63)(99),y=>p(64)(99),Cin=>p(65)(99),clock=>clock,reset=>reset,s=>p(170)(99),cout=>p(171)(100));
FA_ff_2788:FAff port map(x=>p(63)(100),y=>p(64)(100),Cin=>p(65)(100),clock=>clock,reset=>reset,s=>p(170)(100),cout=>p(171)(101));
FA_ff_2789:FAff port map(x=>p(63)(101),y=>p(64)(101),Cin=>p(65)(101),clock=>clock,reset=>reset,s=>p(170)(101),cout=>p(171)(102));
FA_ff_2790:FAff port map(x=>p(63)(102),y=>p(64)(102),Cin=>p(65)(102),clock=>clock,reset=>reset,s=>p(170)(102),cout=>p(171)(103));
FA_ff_2791:FAff port map(x=>p(63)(103),y=>p(64)(103),Cin=>p(65)(103),clock=>clock,reset=>reset,s=>p(170)(103),cout=>p(171)(104));
FA_ff_2792:FAff port map(x=>p(63)(104),y=>p(64)(104),Cin=>p(65)(104),clock=>clock,reset=>reset,s=>p(170)(104),cout=>p(171)(105));
FA_ff_2793:FAff port map(x=>p(63)(105),y=>p(64)(105),Cin=>p(65)(105),clock=>clock,reset=>reset,s=>p(170)(105),cout=>p(171)(106));
FA_ff_2794:FAff port map(x=>p(63)(106),y=>p(64)(106),Cin=>p(65)(106),clock=>clock,reset=>reset,s=>p(170)(106),cout=>p(171)(107));
FA_ff_2795:FAff port map(x=>p(63)(107),y=>p(64)(107),Cin=>p(65)(107),clock=>clock,reset=>reset,s=>p(170)(107),cout=>p(171)(108));
FA_ff_2796:FAff port map(x=>p(63)(108),y=>p(64)(108),Cin=>p(65)(108),clock=>clock,reset=>reset,s=>p(170)(108),cout=>p(171)(109));
FA_ff_2797:FAff port map(x=>p(63)(109),y=>p(64)(109),Cin=>p(65)(109),clock=>clock,reset=>reset,s=>p(170)(109),cout=>p(171)(110));
FA_ff_2798:FAff port map(x=>p(63)(110),y=>p(64)(110),Cin=>p(65)(110),clock=>clock,reset=>reset,s=>p(170)(110),cout=>p(171)(111));
FA_ff_2799:FAff port map(x=>p(63)(111),y=>p(64)(111),Cin=>p(65)(111),clock=>clock,reset=>reset,s=>p(170)(111),cout=>p(171)(112));
FA_ff_2800:FAff port map(x=>p(63)(112),y=>p(64)(112),Cin=>p(65)(112),clock=>clock,reset=>reset,s=>p(170)(112),cout=>p(171)(113));
FA_ff_2801:FAff port map(x=>p(63)(113),y=>p(64)(113),Cin=>p(65)(113),clock=>clock,reset=>reset,s=>p(170)(113),cout=>p(171)(114));
FA_ff_2802:FAff port map(x=>p(63)(114),y=>p(64)(114),Cin=>p(65)(114),clock=>clock,reset=>reset,s=>p(170)(114),cout=>p(171)(115));
FA_ff_2803:FAff port map(x=>p(63)(115),y=>p(64)(115),Cin=>p(65)(115),clock=>clock,reset=>reset,s=>p(170)(115),cout=>p(171)(116));
FA_ff_2804:FAff port map(x=>p(63)(116),y=>p(64)(116),Cin=>p(65)(116),clock=>clock,reset=>reset,s=>p(170)(116),cout=>p(171)(117));
FA_ff_2805:FAff port map(x=>p(63)(117),y=>p(64)(117),Cin=>p(65)(117),clock=>clock,reset=>reset,s=>p(170)(117),cout=>p(171)(118));
FA_ff_2806:FAff port map(x=>p(63)(118),y=>p(64)(118),Cin=>p(65)(118),clock=>clock,reset=>reset,s=>p(170)(118),cout=>p(171)(119));
FA_ff_2807:FAff port map(x=>p(63)(119),y=>p(64)(119),Cin=>p(65)(119),clock=>clock,reset=>reset,s=>p(170)(119),cout=>p(171)(120));
FA_ff_2808:FAff port map(x=>p(63)(120),y=>p(64)(120),Cin=>p(65)(120),clock=>clock,reset=>reset,s=>p(170)(120),cout=>p(171)(121));
FA_ff_2809:FAff port map(x=>p(63)(121),y=>p(64)(121),Cin=>p(65)(121),clock=>clock,reset=>reset,s=>p(170)(121),cout=>p(171)(122));
FA_ff_2810:FAff port map(x=>p(63)(122),y=>p(64)(122),Cin=>p(65)(122),clock=>clock,reset=>reset,s=>p(170)(122),cout=>p(171)(123));
FA_ff_2811:FAff port map(x=>p(63)(123),y=>p(64)(123),Cin=>p(65)(123),clock=>clock,reset=>reset,s=>p(170)(123),cout=>p(171)(124));
FA_ff_2812:FAff port map(x=>p(63)(124),y=>p(64)(124),Cin=>p(65)(124),clock=>clock,reset=>reset,s=>p(170)(124),cout=>p(171)(125));
FA_ff_2813:FAff port map(x=>p(63)(125),y=>p(64)(125),Cin=>p(65)(125),clock=>clock,reset=>reset,s=>p(170)(125),cout=>p(171)(126));
FA_ff_2814:FAff port map(x=>p(63)(126),y=>p(64)(126),Cin=>p(65)(126),clock=>clock,reset=>reset,s=>p(170)(126),cout=>p(171)(127));
FA_ff_2815:FAff port map(x=>p(63)(127),y=>p(64)(127),Cin=>p(65)(127),clock=>clock,reset=>reset,s=>p(170)(127),cout=>p(171)(128));
FA_ff_2816:FAff port map(x=>p(66)(0),y=>p(67)(0),Cin=>p(68)(0),clock=>clock,reset=>reset,s=>p(172)(0),cout=>p(173)(1));
FA_ff_2817:FAff port map(x=>p(66)(1),y=>p(67)(1),Cin=>p(68)(1),clock=>clock,reset=>reset,s=>p(172)(1),cout=>p(173)(2));
FA_ff_2818:FAff port map(x=>p(66)(2),y=>p(67)(2),Cin=>p(68)(2),clock=>clock,reset=>reset,s=>p(172)(2),cout=>p(173)(3));
FA_ff_2819:FAff port map(x=>p(66)(3),y=>p(67)(3),Cin=>p(68)(3),clock=>clock,reset=>reset,s=>p(172)(3),cout=>p(173)(4));
FA_ff_2820:FAff port map(x=>p(66)(4),y=>p(67)(4),Cin=>p(68)(4),clock=>clock,reset=>reset,s=>p(172)(4),cout=>p(173)(5));
FA_ff_2821:FAff port map(x=>p(66)(5),y=>p(67)(5),Cin=>p(68)(5),clock=>clock,reset=>reset,s=>p(172)(5),cout=>p(173)(6));
FA_ff_2822:FAff port map(x=>p(66)(6),y=>p(67)(6),Cin=>p(68)(6),clock=>clock,reset=>reset,s=>p(172)(6),cout=>p(173)(7));
FA_ff_2823:FAff port map(x=>p(66)(7),y=>p(67)(7),Cin=>p(68)(7),clock=>clock,reset=>reset,s=>p(172)(7),cout=>p(173)(8));
FA_ff_2824:FAff port map(x=>p(66)(8),y=>p(67)(8),Cin=>p(68)(8),clock=>clock,reset=>reset,s=>p(172)(8),cout=>p(173)(9));
FA_ff_2825:FAff port map(x=>p(66)(9),y=>p(67)(9),Cin=>p(68)(9),clock=>clock,reset=>reset,s=>p(172)(9),cout=>p(173)(10));
FA_ff_2826:FAff port map(x=>p(66)(10),y=>p(67)(10),Cin=>p(68)(10),clock=>clock,reset=>reset,s=>p(172)(10),cout=>p(173)(11));
FA_ff_2827:FAff port map(x=>p(66)(11),y=>p(67)(11),Cin=>p(68)(11),clock=>clock,reset=>reset,s=>p(172)(11),cout=>p(173)(12));
FA_ff_2828:FAff port map(x=>p(66)(12),y=>p(67)(12),Cin=>p(68)(12),clock=>clock,reset=>reset,s=>p(172)(12),cout=>p(173)(13));
FA_ff_2829:FAff port map(x=>p(66)(13),y=>p(67)(13),Cin=>p(68)(13),clock=>clock,reset=>reset,s=>p(172)(13),cout=>p(173)(14));
FA_ff_2830:FAff port map(x=>p(66)(14),y=>p(67)(14),Cin=>p(68)(14),clock=>clock,reset=>reset,s=>p(172)(14),cout=>p(173)(15));
FA_ff_2831:FAff port map(x=>p(66)(15),y=>p(67)(15),Cin=>p(68)(15),clock=>clock,reset=>reset,s=>p(172)(15),cout=>p(173)(16));
FA_ff_2832:FAff port map(x=>p(66)(16),y=>p(67)(16),Cin=>p(68)(16),clock=>clock,reset=>reset,s=>p(172)(16),cout=>p(173)(17));
FA_ff_2833:FAff port map(x=>p(66)(17),y=>p(67)(17),Cin=>p(68)(17),clock=>clock,reset=>reset,s=>p(172)(17),cout=>p(173)(18));
FA_ff_2834:FAff port map(x=>p(66)(18),y=>p(67)(18),Cin=>p(68)(18),clock=>clock,reset=>reset,s=>p(172)(18),cout=>p(173)(19));
FA_ff_2835:FAff port map(x=>p(66)(19),y=>p(67)(19),Cin=>p(68)(19),clock=>clock,reset=>reset,s=>p(172)(19),cout=>p(173)(20));
FA_ff_2836:FAff port map(x=>p(66)(20),y=>p(67)(20),Cin=>p(68)(20),clock=>clock,reset=>reset,s=>p(172)(20),cout=>p(173)(21));
FA_ff_2837:FAff port map(x=>p(66)(21),y=>p(67)(21),Cin=>p(68)(21),clock=>clock,reset=>reset,s=>p(172)(21),cout=>p(173)(22));
FA_ff_2838:FAff port map(x=>p(66)(22),y=>p(67)(22),Cin=>p(68)(22),clock=>clock,reset=>reset,s=>p(172)(22),cout=>p(173)(23));
FA_ff_2839:FAff port map(x=>p(66)(23),y=>p(67)(23),Cin=>p(68)(23),clock=>clock,reset=>reset,s=>p(172)(23),cout=>p(173)(24));
FA_ff_2840:FAff port map(x=>p(66)(24),y=>p(67)(24),Cin=>p(68)(24),clock=>clock,reset=>reset,s=>p(172)(24),cout=>p(173)(25));
FA_ff_2841:FAff port map(x=>p(66)(25),y=>p(67)(25),Cin=>p(68)(25),clock=>clock,reset=>reset,s=>p(172)(25),cout=>p(173)(26));
FA_ff_2842:FAff port map(x=>p(66)(26),y=>p(67)(26),Cin=>p(68)(26),clock=>clock,reset=>reset,s=>p(172)(26),cout=>p(173)(27));
FA_ff_2843:FAff port map(x=>p(66)(27),y=>p(67)(27),Cin=>p(68)(27),clock=>clock,reset=>reset,s=>p(172)(27),cout=>p(173)(28));
FA_ff_2844:FAff port map(x=>p(66)(28),y=>p(67)(28),Cin=>p(68)(28),clock=>clock,reset=>reset,s=>p(172)(28),cout=>p(173)(29));
FA_ff_2845:FAff port map(x=>p(66)(29),y=>p(67)(29),Cin=>p(68)(29),clock=>clock,reset=>reset,s=>p(172)(29),cout=>p(173)(30));
FA_ff_2846:FAff port map(x=>p(66)(30),y=>p(67)(30),Cin=>p(68)(30),clock=>clock,reset=>reset,s=>p(172)(30),cout=>p(173)(31));
FA_ff_2847:FAff port map(x=>p(66)(31),y=>p(67)(31),Cin=>p(68)(31),clock=>clock,reset=>reset,s=>p(172)(31),cout=>p(173)(32));
FA_ff_2848:FAff port map(x=>p(66)(32),y=>p(67)(32),Cin=>p(68)(32),clock=>clock,reset=>reset,s=>p(172)(32),cout=>p(173)(33));
FA_ff_2849:FAff port map(x=>p(66)(33),y=>p(67)(33),Cin=>p(68)(33),clock=>clock,reset=>reset,s=>p(172)(33),cout=>p(173)(34));
FA_ff_2850:FAff port map(x=>p(66)(34),y=>p(67)(34),Cin=>p(68)(34),clock=>clock,reset=>reset,s=>p(172)(34),cout=>p(173)(35));
FA_ff_2851:FAff port map(x=>p(66)(35),y=>p(67)(35),Cin=>p(68)(35),clock=>clock,reset=>reset,s=>p(172)(35),cout=>p(173)(36));
FA_ff_2852:FAff port map(x=>p(66)(36),y=>p(67)(36),Cin=>p(68)(36),clock=>clock,reset=>reset,s=>p(172)(36),cout=>p(173)(37));
FA_ff_2853:FAff port map(x=>p(66)(37),y=>p(67)(37),Cin=>p(68)(37),clock=>clock,reset=>reset,s=>p(172)(37),cout=>p(173)(38));
FA_ff_2854:FAff port map(x=>p(66)(38),y=>p(67)(38),Cin=>p(68)(38),clock=>clock,reset=>reset,s=>p(172)(38),cout=>p(173)(39));
FA_ff_2855:FAff port map(x=>p(66)(39),y=>p(67)(39),Cin=>p(68)(39),clock=>clock,reset=>reset,s=>p(172)(39),cout=>p(173)(40));
FA_ff_2856:FAff port map(x=>p(66)(40),y=>p(67)(40),Cin=>p(68)(40),clock=>clock,reset=>reset,s=>p(172)(40),cout=>p(173)(41));
FA_ff_2857:FAff port map(x=>p(66)(41),y=>p(67)(41),Cin=>p(68)(41),clock=>clock,reset=>reset,s=>p(172)(41),cout=>p(173)(42));
FA_ff_2858:FAff port map(x=>p(66)(42),y=>p(67)(42),Cin=>p(68)(42),clock=>clock,reset=>reset,s=>p(172)(42),cout=>p(173)(43));
FA_ff_2859:FAff port map(x=>p(66)(43),y=>p(67)(43),Cin=>p(68)(43),clock=>clock,reset=>reset,s=>p(172)(43),cout=>p(173)(44));
FA_ff_2860:FAff port map(x=>p(66)(44),y=>p(67)(44),Cin=>p(68)(44),clock=>clock,reset=>reset,s=>p(172)(44),cout=>p(173)(45));
FA_ff_2861:FAff port map(x=>p(66)(45),y=>p(67)(45),Cin=>p(68)(45),clock=>clock,reset=>reset,s=>p(172)(45),cout=>p(173)(46));
FA_ff_2862:FAff port map(x=>p(66)(46),y=>p(67)(46),Cin=>p(68)(46),clock=>clock,reset=>reset,s=>p(172)(46),cout=>p(173)(47));
FA_ff_2863:FAff port map(x=>p(66)(47),y=>p(67)(47),Cin=>p(68)(47),clock=>clock,reset=>reset,s=>p(172)(47),cout=>p(173)(48));
FA_ff_2864:FAff port map(x=>p(66)(48),y=>p(67)(48),Cin=>p(68)(48),clock=>clock,reset=>reset,s=>p(172)(48),cout=>p(173)(49));
FA_ff_2865:FAff port map(x=>p(66)(49),y=>p(67)(49),Cin=>p(68)(49),clock=>clock,reset=>reset,s=>p(172)(49),cout=>p(173)(50));
FA_ff_2866:FAff port map(x=>p(66)(50),y=>p(67)(50),Cin=>p(68)(50),clock=>clock,reset=>reset,s=>p(172)(50),cout=>p(173)(51));
FA_ff_2867:FAff port map(x=>p(66)(51),y=>p(67)(51),Cin=>p(68)(51),clock=>clock,reset=>reset,s=>p(172)(51),cout=>p(173)(52));
FA_ff_2868:FAff port map(x=>p(66)(52),y=>p(67)(52),Cin=>p(68)(52),clock=>clock,reset=>reset,s=>p(172)(52),cout=>p(173)(53));
FA_ff_2869:FAff port map(x=>p(66)(53),y=>p(67)(53),Cin=>p(68)(53),clock=>clock,reset=>reset,s=>p(172)(53),cout=>p(173)(54));
FA_ff_2870:FAff port map(x=>p(66)(54),y=>p(67)(54),Cin=>p(68)(54),clock=>clock,reset=>reset,s=>p(172)(54),cout=>p(173)(55));
FA_ff_2871:FAff port map(x=>p(66)(55),y=>p(67)(55),Cin=>p(68)(55),clock=>clock,reset=>reset,s=>p(172)(55),cout=>p(173)(56));
FA_ff_2872:FAff port map(x=>p(66)(56),y=>p(67)(56),Cin=>p(68)(56),clock=>clock,reset=>reset,s=>p(172)(56),cout=>p(173)(57));
FA_ff_2873:FAff port map(x=>p(66)(57),y=>p(67)(57),Cin=>p(68)(57),clock=>clock,reset=>reset,s=>p(172)(57),cout=>p(173)(58));
FA_ff_2874:FAff port map(x=>p(66)(58),y=>p(67)(58),Cin=>p(68)(58),clock=>clock,reset=>reset,s=>p(172)(58),cout=>p(173)(59));
FA_ff_2875:FAff port map(x=>p(66)(59),y=>p(67)(59),Cin=>p(68)(59),clock=>clock,reset=>reset,s=>p(172)(59),cout=>p(173)(60));
FA_ff_2876:FAff port map(x=>p(66)(60),y=>p(67)(60),Cin=>p(68)(60),clock=>clock,reset=>reset,s=>p(172)(60),cout=>p(173)(61));
FA_ff_2877:FAff port map(x=>p(66)(61),y=>p(67)(61),Cin=>p(68)(61),clock=>clock,reset=>reset,s=>p(172)(61),cout=>p(173)(62));
FA_ff_2878:FAff port map(x=>p(66)(62),y=>p(67)(62),Cin=>p(68)(62),clock=>clock,reset=>reset,s=>p(172)(62),cout=>p(173)(63));
FA_ff_2879:FAff port map(x=>p(66)(63),y=>p(67)(63),Cin=>p(68)(63),clock=>clock,reset=>reset,s=>p(172)(63),cout=>p(173)(64));
FA_ff_2880:FAff port map(x=>p(66)(64),y=>p(67)(64),Cin=>p(68)(64),clock=>clock,reset=>reset,s=>p(172)(64),cout=>p(173)(65));
FA_ff_2881:FAff port map(x=>p(66)(65),y=>p(67)(65),Cin=>p(68)(65),clock=>clock,reset=>reset,s=>p(172)(65),cout=>p(173)(66));
FA_ff_2882:FAff port map(x=>p(66)(66),y=>p(67)(66),Cin=>p(68)(66),clock=>clock,reset=>reset,s=>p(172)(66),cout=>p(173)(67));
FA_ff_2883:FAff port map(x=>p(66)(67),y=>p(67)(67),Cin=>p(68)(67),clock=>clock,reset=>reset,s=>p(172)(67),cout=>p(173)(68));
FA_ff_2884:FAff port map(x=>p(66)(68),y=>p(67)(68),Cin=>p(68)(68),clock=>clock,reset=>reset,s=>p(172)(68),cout=>p(173)(69));
FA_ff_2885:FAff port map(x=>p(66)(69),y=>p(67)(69),Cin=>p(68)(69),clock=>clock,reset=>reset,s=>p(172)(69),cout=>p(173)(70));
FA_ff_2886:FAff port map(x=>p(66)(70),y=>p(67)(70),Cin=>p(68)(70),clock=>clock,reset=>reset,s=>p(172)(70),cout=>p(173)(71));
FA_ff_2887:FAff port map(x=>p(66)(71),y=>p(67)(71),Cin=>p(68)(71),clock=>clock,reset=>reset,s=>p(172)(71),cout=>p(173)(72));
FA_ff_2888:FAff port map(x=>p(66)(72),y=>p(67)(72),Cin=>p(68)(72),clock=>clock,reset=>reset,s=>p(172)(72),cout=>p(173)(73));
FA_ff_2889:FAff port map(x=>p(66)(73),y=>p(67)(73),Cin=>p(68)(73),clock=>clock,reset=>reset,s=>p(172)(73),cout=>p(173)(74));
FA_ff_2890:FAff port map(x=>p(66)(74),y=>p(67)(74),Cin=>p(68)(74),clock=>clock,reset=>reset,s=>p(172)(74),cout=>p(173)(75));
FA_ff_2891:FAff port map(x=>p(66)(75),y=>p(67)(75),Cin=>p(68)(75),clock=>clock,reset=>reset,s=>p(172)(75),cout=>p(173)(76));
FA_ff_2892:FAff port map(x=>p(66)(76),y=>p(67)(76),Cin=>p(68)(76),clock=>clock,reset=>reset,s=>p(172)(76),cout=>p(173)(77));
FA_ff_2893:FAff port map(x=>p(66)(77),y=>p(67)(77),Cin=>p(68)(77),clock=>clock,reset=>reset,s=>p(172)(77),cout=>p(173)(78));
FA_ff_2894:FAff port map(x=>p(66)(78),y=>p(67)(78),Cin=>p(68)(78),clock=>clock,reset=>reset,s=>p(172)(78),cout=>p(173)(79));
FA_ff_2895:FAff port map(x=>p(66)(79),y=>p(67)(79),Cin=>p(68)(79),clock=>clock,reset=>reset,s=>p(172)(79),cout=>p(173)(80));
FA_ff_2896:FAff port map(x=>p(66)(80),y=>p(67)(80),Cin=>p(68)(80),clock=>clock,reset=>reset,s=>p(172)(80),cout=>p(173)(81));
FA_ff_2897:FAff port map(x=>p(66)(81),y=>p(67)(81),Cin=>p(68)(81),clock=>clock,reset=>reset,s=>p(172)(81),cout=>p(173)(82));
FA_ff_2898:FAff port map(x=>p(66)(82),y=>p(67)(82),Cin=>p(68)(82),clock=>clock,reset=>reset,s=>p(172)(82),cout=>p(173)(83));
FA_ff_2899:FAff port map(x=>p(66)(83),y=>p(67)(83),Cin=>p(68)(83),clock=>clock,reset=>reset,s=>p(172)(83),cout=>p(173)(84));
FA_ff_2900:FAff port map(x=>p(66)(84),y=>p(67)(84),Cin=>p(68)(84),clock=>clock,reset=>reset,s=>p(172)(84),cout=>p(173)(85));
FA_ff_2901:FAff port map(x=>p(66)(85),y=>p(67)(85),Cin=>p(68)(85),clock=>clock,reset=>reset,s=>p(172)(85),cout=>p(173)(86));
FA_ff_2902:FAff port map(x=>p(66)(86),y=>p(67)(86),Cin=>p(68)(86),clock=>clock,reset=>reset,s=>p(172)(86),cout=>p(173)(87));
FA_ff_2903:FAff port map(x=>p(66)(87),y=>p(67)(87),Cin=>p(68)(87),clock=>clock,reset=>reset,s=>p(172)(87),cout=>p(173)(88));
FA_ff_2904:FAff port map(x=>p(66)(88),y=>p(67)(88),Cin=>p(68)(88),clock=>clock,reset=>reset,s=>p(172)(88),cout=>p(173)(89));
FA_ff_2905:FAff port map(x=>p(66)(89),y=>p(67)(89),Cin=>p(68)(89),clock=>clock,reset=>reset,s=>p(172)(89),cout=>p(173)(90));
FA_ff_2906:FAff port map(x=>p(66)(90),y=>p(67)(90),Cin=>p(68)(90),clock=>clock,reset=>reset,s=>p(172)(90),cout=>p(173)(91));
FA_ff_2907:FAff port map(x=>p(66)(91),y=>p(67)(91),Cin=>p(68)(91),clock=>clock,reset=>reset,s=>p(172)(91),cout=>p(173)(92));
FA_ff_2908:FAff port map(x=>p(66)(92),y=>p(67)(92),Cin=>p(68)(92),clock=>clock,reset=>reset,s=>p(172)(92),cout=>p(173)(93));
FA_ff_2909:FAff port map(x=>p(66)(93),y=>p(67)(93),Cin=>p(68)(93),clock=>clock,reset=>reset,s=>p(172)(93),cout=>p(173)(94));
FA_ff_2910:FAff port map(x=>p(66)(94),y=>p(67)(94),Cin=>p(68)(94),clock=>clock,reset=>reset,s=>p(172)(94),cout=>p(173)(95));
FA_ff_2911:FAff port map(x=>p(66)(95),y=>p(67)(95),Cin=>p(68)(95),clock=>clock,reset=>reset,s=>p(172)(95),cout=>p(173)(96));
FA_ff_2912:FAff port map(x=>p(66)(96),y=>p(67)(96),Cin=>p(68)(96),clock=>clock,reset=>reset,s=>p(172)(96),cout=>p(173)(97));
FA_ff_2913:FAff port map(x=>p(66)(97),y=>p(67)(97),Cin=>p(68)(97),clock=>clock,reset=>reset,s=>p(172)(97),cout=>p(173)(98));
FA_ff_2914:FAff port map(x=>p(66)(98),y=>p(67)(98),Cin=>p(68)(98),clock=>clock,reset=>reset,s=>p(172)(98),cout=>p(173)(99));
FA_ff_2915:FAff port map(x=>p(66)(99),y=>p(67)(99),Cin=>p(68)(99),clock=>clock,reset=>reset,s=>p(172)(99),cout=>p(173)(100));
FA_ff_2916:FAff port map(x=>p(66)(100),y=>p(67)(100),Cin=>p(68)(100),clock=>clock,reset=>reset,s=>p(172)(100),cout=>p(173)(101));
FA_ff_2917:FAff port map(x=>p(66)(101),y=>p(67)(101),Cin=>p(68)(101),clock=>clock,reset=>reset,s=>p(172)(101),cout=>p(173)(102));
FA_ff_2918:FAff port map(x=>p(66)(102),y=>p(67)(102),Cin=>p(68)(102),clock=>clock,reset=>reset,s=>p(172)(102),cout=>p(173)(103));
FA_ff_2919:FAff port map(x=>p(66)(103),y=>p(67)(103),Cin=>p(68)(103),clock=>clock,reset=>reset,s=>p(172)(103),cout=>p(173)(104));
FA_ff_2920:FAff port map(x=>p(66)(104),y=>p(67)(104),Cin=>p(68)(104),clock=>clock,reset=>reset,s=>p(172)(104),cout=>p(173)(105));
FA_ff_2921:FAff port map(x=>p(66)(105),y=>p(67)(105),Cin=>p(68)(105),clock=>clock,reset=>reset,s=>p(172)(105),cout=>p(173)(106));
FA_ff_2922:FAff port map(x=>p(66)(106),y=>p(67)(106),Cin=>p(68)(106),clock=>clock,reset=>reset,s=>p(172)(106),cout=>p(173)(107));
FA_ff_2923:FAff port map(x=>p(66)(107),y=>p(67)(107),Cin=>p(68)(107),clock=>clock,reset=>reset,s=>p(172)(107),cout=>p(173)(108));
FA_ff_2924:FAff port map(x=>p(66)(108),y=>p(67)(108),Cin=>p(68)(108),clock=>clock,reset=>reset,s=>p(172)(108),cout=>p(173)(109));
FA_ff_2925:FAff port map(x=>p(66)(109),y=>p(67)(109),Cin=>p(68)(109),clock=>clock,reset=>reset,s=>p(172)(109),cout=>p(173)(110));
FA_ff_2926:FAff port map(x=>p(66)(110),y=>p(67)(110),Cin=>p(68)(110),clock=>clock,reset=>reset,s=>p(172)(110),cout=>p(173)(111));
FA_ff_2927:FAff port map(x=>p(66)(111),y=>p(67)(111),Cin=>p(68)(111),clock=>clock,reset=>reset,s=>p(172)(111),cout=>p(173)(112));
FA_ff_2928:FAff port map(x=>p(66)(112),y=>p(67)(112),Cin=>p(68)(112),clock=>clock,reset=>reset,s=>p(172)(112),cout=>p(173)(113));
FA_ff_2929:FAff port map(x=>p(66)(113),y=>p(67)(113),Cin=>p(68)(113),clock=>clock,reset=>reset,s=>p(172)(113),cout=>p(173)(114));
FA_ff_2930:FAff port map(x=>p(66)(114),y=>p(67)(114),Cin=>p(68)(114),clock=>clock,reset=>reset,s=>p(172)(114),cout=>p(173)(115));
FA_ff_2931:FAff port map(x=>p(66)(115),y=>p(67)(115),Cin=>p(68)(115),clock=>clock,reset=>reset,s=>p(172)(115),cout=>p(173)(116));
FA_ff_2932:FAff port map(x=>p(66)(116),y=>p(67)(116),Cin=>p(68)(116),clock=>clock,reset=>reset,s=>p(172)(116),cout=>p(173)(117));
FA_ff_2933:FAff port map(x=>p(66)(117),y=>p(67)(117),Cin=>p(68)(117),clock=>clock,reset=>reset,s=>p(172)(117),cout=>p(173)(118));
FA_ff_2934:FAff port map(x=>p(66)(118),y=>p(67)(118),Cin=>p(68)(118),clock=>clock,reset=>reset,s=>p(172)(118),cout=>p(173)(119));
FA_ff_2935:FAff port map(x=>p(66)(119),y=>p(67)(119),Cin=>p(68)(119),clock=>clock,reset=>reset,s=>p(172)(119),cout=>p(173)(120));
FA_ff_2936:FAff port map(x=>p(66)(120),y=>p(67)(120),Cin=>p(68)(120),clock=>clock,reset=>reset,s=>p(172)(120),cout=>p(173)(121));
FA_ff_2937:FAff port map(x=>p(66)(121),y=>p(67)(121),Cin=>p(68)(121),clock=>clock,reset=>reset,s=>p(172)(121),cout=>p(173)(122));
FA_ff_2938:FAff port map(x=>p(66)(122),y=>p(67)(122),Cin=>p(68)(122),clock=>clock,reset=>reset,s=>p(172)(122),cout=>p(173)(123));
FA_ff_2939:FAff port map(x=>p(66)(123),y=>p(67)(123),Cin=>p(68)(123),clock=>clock,reset=>reset,s=>p(172)(123),cout=>p(173)(124));
FA_ff_2940:FAff port map(x=>p(66)(124),y=>p(67)(124),Cin=>p(68)(124),clock=>clock,reset=>reset,s=>p(172)(124),cout=>p(173)(125));
FA_ff_2941:FAff port map(x=>p(66)(125),y=>p(67)(125),Cin=>p(68)(125),clock=>clock,reset=>reset,s=>p(172)(125),cout=>p(173)(126));
FA_ff_2942:FAff port map(x=>p(66)(126),y=>p(67)(126),Cin=>p(68)(126),clock=>clock,reset=>reset,s=>p(172)(126),cout=>p(173)(127));
FA_ff_2943:FAff port map(x=>p(66)(127),y=>p(67)(127),Cin=>p(68)(127),clock=>clock,reset=>reset,s=>p(172)(127),cout=>p(173)(128));
FA_ff_2944:FAff port map(x=>p(69)(0),y=>p(70)(0),Cin=>p(71)(0),clock=>clock,reset=>reset,s=>p(174)(0),cout=>p(175)(1));
FA_ff_2945:FAff port map(x=>p(69)(1),y=>p(70)(1),Cin=>p(71)(1),clock=>clock,reset=>reset,s=>p(174)(1),cout=>p(175)(2));
FA_ff_2946:FAff port map(x=>p(69)(2),y=>p(70)(2),Cin=>p(71)(2),clock=>clock,reset=>reset,s=>p(174)(2),cout=>p(175)(3));
FA_ff_2947:FAff port map(x=>p(69)(3),y=>p(70)(3),Cin=>p(71)(3),clock=>clock,reset=>reset,s=>p(174)(3),cout=>p(175)(4));
FA_ff_2948:FAff port map(x=>p(69)(4),y=>p(70)(4),Cin=>p(71)(4),clock=>clock,reset=>reset,s=>p(174)(4),cout=>p(175)(5));
FA_ff_2949:FAff port map(x=>p(69)(5),y=>p(70)(5),Cin=>p(71)(5),clock=>clock,reset=>reset,s=>p(174)(5),cout=>p(175)(6));
FA_ff_2950:FAff port map(x=>p(69)(6),y=>p(70)(6),Cin=>p(71)(6),clock=>clock,reset=>reset,s=>p(174)(6),cout=>p(175)(7));
FA_ff_2951:FAff port map(x=>p(69)(7),y=>p(70)(7),Cin=>p(71)(7),clock=>clock,reset=>reset,s=>p(174)(7),cout=>p(175)(8));
FA_ff_2952:FAff port map(x=>p(69)(8),y=>p(70)(8),Cin=>p(71)(8),clock=>clock,reset=>reset,s=>p(174)(8),cout=>p(175)(9));
FA_ff_2953:FAff port map(x=>p(69)(9),y=>p(70)(9),Cin=>p(71)(9),clock=>clock,reset=>reset,s=>p(174)(9),cout=>p(175)(10));
FA_ff_2954:FAff port map(x=>p(69)(10),y=>p(70)(10),Cin=>p(71)(10),clock=>clock,reset=>reset,s=>p(174)(10),cout=>p(175)(11));
FA_ff_2955:FAff port map(x=>p(69)(11),y=>p(70)(11),Cin=>p(71)(11),clock=>clock,reset=>reset,s=>p(174)(11),cout=>p(175)(12));
FA_ff_2956:FAff port map(x=>p(69)(12),y=>p(70)(12),Cin=>p(71)(12),clock=>clock,reset=>reset,s=>p(174)(12),cout=>p(175)(13));
FA_ff_2957:FAff port map(x=>p(69)(13),y=>p(70)(13),Cin=>p(71)(13),clock=>clock,reset=>reset,s=>p(174)(13),cout=>p(175)(14));
FA_ff_2958:FAff port map(x=>p(69)(14),y=>p(70)(14),Cin=>p(71)(14),clock=>clock,reset=>reset,s=>p(174)(14),cout=>p(175)(15));
FA_ff_2959:FAff port map(x=>p(69)(15),y=>p(70)(15),Cin=>p(71)(15),clock=>clock,reset=>reset,s=>p(174)(15),cout=>p(175)(16));
FA_ff_2960:FAff port map(x=>p(69)(16),y=>p(70)(16),Cin=>p(71)(16),clock=>clock,reset=>reset,s=>p(174)(16),cout=>p(175)(17));
FA_ff_2961:FAff port map(x=>p(69)(17),y=>p(70)(17),Cin=>p(71)(17),clock=>clock,reset=>reset,s=>p(174)(17),cout=>p(175)(18));
FA_ff_2962:FAff port map(x=>p(69)(18),y=>p(70)(18),Cin=>p(71)(18),clock=>clock,reset=>reset,s=>p(174)(18),cout=>p(175)(19));
FA_ff_2963:FAff port map(x=>p(69)(19),y=>p(70)(19),Cin=>p(71)(19),clock=>clock,reset=>reset,s=>p(174)(19),cout=>p(175)(20));
FA_ff_2964:FAff port map(x=>p(69)(20),y=>p(70)(20),Cin=>p(71)(20),clock=>clock,reset=>reset,s=>p(174)(20),cout=>p(175)(21));
FA_ff_2965:FAff port map(x=>p(69)(21),y=>p(70)(21),Cin=>p(71)(21),clock=>clock,reset=>reset,s=>p(174)(21),cout=>p(175)(22));
FA_ff_2966:FAff port map(x=>p(69)(22),y=>p(70)(22),Cin=>p(71)(22),clock=>clock,reset=>reset,s=>p(174)(22),cout=>p(175)(23));
FA_ff_2967:FAff port map(x=>p(69)(23),y=>p(70)(23),Cin=>p(71)(23),clock=>clock,reset=>reset,s=>p(174)(23),cout=>p(175)(24));
FA_ff_2968:FAff port map(x=>p(69)(24),y=>p(70)(24),Cin=>p(71)(24),clock=>clock,reset=>reset,s=>p(174)(24),cout=>p(175)(25));
FA_ff_2969:FAff port map(x=>p(69)(25),y=>p(70)(25),Cin=>p(71)(25),clock=>clock,reset=>reset,s=>p(174)(25),cout=>p(175)(26));
FA_ff_2970:FAff port map(x=>p(69)(26),y=>p(70)(26),Cin=>p(71)(26),clock=>clock,reset=>reset,s=>p(174)(26),cout=>p(175)(27));
FA_ff_2971:FAff port map(x=>p(69)(27),y=>p(70)(27),Cin=>p(71)(27),clock=>clock,reset=>reset,s=>p(174)(27),cout=>p(175)(28));
FA_ff_2972:FAff port map(x=>p(69)(28),y=>p(70)(28),Cin=>p(71)(28),clock=>clock,reset=>reset,s=>p(174)(28),cout=>p(175)(29));
FA_ff_2973:FAff port map(x=>p(69)(29),y=>p(70)(29),Cin=>p(71)(29),clock=>clock,reset=>reset,s=>p(174)(29),cout=>p(175)(30));
FA_ff_2974:FAff port map(x=>p(69)(30),y=>p(70)(30),Cin=>p(71)(30),clock=>clock,reset=>reset,s=>p(174)(30),cout=>p(175)(31));
FA_ff_2975:FAff port map(x=>p(69)(31),y=>p(70)(31),Cin=>p(71)(31),clock=>clock,reset=>reset,s=>p(174)(31),cout=>p(175)(32));
FA_ff_2976:FAff port map(x=>p(69)(32),y=>p(70)(32),Cin=>p(71)(32),clock=>clock,reset=>reset,s=>p(174)(32),cout=>p(175)(33));
FA_ff_2977:FAff port map(x=>p(69)(33),y=>p(70)(33),Cin=>p(71)(33),clock=>clock,reset=>reset,s=>p(174)(33),cout=>p(175)(34));
FA_ff_2978:FAff port map(x=>p(69)(34),y=>p(70)(34),Cin=>p(71)(34),clock=>clock,reset=>reset,s=>p(174)(34),cout=>p(175)(35));
FA_ff_2979:FAff port map(x=>p(69)(35),y=>p(70)(35),Cin=>p(71)(35),clock=>clock,reset=>reset,s=>p(174)(35),cout=>p(175)(36));
FA_ff_2980:FAff port map(x=>p(69)(36),y=>p(70)(36),Cin=>p(71)(36),clock=>clock,reset=>reset,s=>p(174)(36),cout=>p(175)(37));
FA_ff_2981:FAff port map(x=>p(69)(37),y=>p(70)(37),Cin=>p(71)(37),clock=>clock,reset=>reset,s=>p(174)(37),cout=>p(175)(38));
FA_ff_2982:FAff port map(x=>p(69)(38),y=>p(70)(38),Cin=>p(71)(38),clock=>clock,reset=>reset,s=>p(174)(38),cout=>p(175)(39));
FA_ff_2983:FAff port map(x=>p(69)(39),y=>p(70)(39),Cin=>p(71)(39),clock=>clock,reset=>reset,s=>p(174)(39),cout=>p(175)(40));
FA_ff_2984:FAff port map(x=>p(69)(40),y=>p(70)(40),Cin=>p(71)(40),clock=>clock,reset=>reset,s=>p(174)(40),cout=>p(175)(41));
FA_ff_2985:FAff port map(x=>p(69)(41),y=>p(70)(41),Cin=>p(71)(41),clock=>clock,reset=>reset,s=>p(174)(41),cout=>p(175)(42));
FA_ff_2986:FAff port map(x=>p(69)(42),y=>p(70)(42),Cin=>p(71)(42),clock=>clock,reset=>reset,s=>p(174)(42),cout=>p(175)(43));
FA_ff_2987:FAff port map(x=>p(69)(43),y=>p(70)(43),Cin=>p(71)(43),clock=>clock,reset=>reset,s=>p(174)(43),cout=>p(175)(44));
FA_ff_2988:FAff port map(x=>p(69)(44),y=>p(70)(44),Cin=>p(71)(44),clock=>clock,reset=>reset,s=>p(174)(44),cout=>p(175)(45));
FA_ff_2989:FAff port map(x=>p(69)(45),y=>p(70)(45),Cin=>p(71)(45),clock=>clock,reset=>reset,s=>p(174)(45),cout=>p(175)(46));
FA_ff_2990:FAff port map(x=>p(69)(46),y=>p(70)(46),Cin=>p(71)(46),clock=>clock,reset=>reset,s=>p(174)(46),cout=>p(175)(47));
FA_ff_2991:FAff port map(x=>p(69)(47),y=>p(70)(47),Cin=>p(71)(47),clock=>clock,reset=>reset,s=>p(174)(47),cout=>p(175)(48));
FA_ff_2992:FAff port map(x=>p(69)(48),y=>p(70)(48),Cin=>p(71)(48),clock=>clock,reset=>reset,s=>p(174)(48),cout=>p(175)(49));
FA_ff_2993:FAff port map(x=>p(69)(49),y=>p(70)(49),Cin=>p(71)(49),clock=>clock,reset=>reset,s=>p(174)(49),cout=>p(175)(50));
FA_ff_2994:FAff port map(x=>p(69)(50),y=>p(70)(50),Cin=>p(71)(50),clock=>clock,reset=>reset,s=>p(174)(50),cout=>p(175)(51));
FA_ff_2995:FAff port map(x=>p(69)(51),y=>p(70)(51),Cin=>p(71)(51),clock=>clock,reset=>reset,s=>p(174)(51),cout=>p(175)(52));
FA_ff_2996:FAff port map(x=>p(69)(52),y=>p(70)(52),Cin=>p(71)(52),clock=>clock,reset=>reset,s=>p(174)(52),cout=>p(175)(53));
FA_ff_2997:FAff port map(x=>p(69)(53),y=>p(70)(53),Cin=>p(71)(53),clock=>clock,reset=>reset,s=>p(174)(53),cout=>p(175)(54));
FA_ff_2998:FAff port map(x=>p(69)(54),y=>p(70)(54),Cin=>p(71)(54),clock=>clock,reset=>reset,s=>p(174)(54),cout=>p(175)(55));
FA_ff_2999:FAff port map(x=>p(69)(55),y=>p(70)(55),Cin=>p(71)(55),clock=>clock,reset=>reset,s=>p(174)(55),cout=>p(175)(56));
FA_ff_3000:FAff port map(x=>p(69)(56),y=>p(70)(56),Cin=>p(71)(56),clock=>clock,reset=>reset,s=>p(174)(56),cout=>p(175)(57));
FA_ff_3001:FAff port map(x=>p(69)(57),y=>p(70)(57),Cin=>p(71)(57),clock=>clock,reset=>reset,s=>p(174)(57),cout=>p(175)(58));
FA_ff_3002:FAff port map(x=>p(69)(58),y=>p(70)(58),Cin=>p(71)(58),clock=>clock,reset=>reset,s=>p(174)(58),cout=>p(175)(59));
FA_ff_3003:FAff port map(x=>p(69)(59),y=>p(70)(59),Cin=>p(71)(59),clock=>clock,reset=>reset,s=>p(174)(59),cout=>p(175)(60));
FA_ff_3004:FAff port map(x=>p(69)(60),y=>p(70)(60),Cin=>p(71)(60),clock=>clock,reset=>reset,s=>p(174)(60),cout=>p(175)(61));
FA_ff_3005:FAff port map(x=>p(69)(61),y=>p(70)(61),Cin=>p(71)(61),clock=>clock,reset=>reset,s=>p(174)(61),cout=>p(175)(62));
FA_ff_3006:FAff port map(x=>p(69)(62),y=>p(70)(62),Cin=>p(71)(62),clock=>clock,reset=>reset,s=>p(174)(62),cout=>p(175)(63));
FA_ff_3007:FAff port map(x=>p(69)(63),y=>p(70)(63),Cin=>p(71)(63),clock=>clock,reset=>reset,s=>p(174)(63),cout=>p(175)(64));
FA_ff_3008:FAff port map(x=>p(69)(64),y=>p(70)(64),Cin=>p(71)(64),clock=>clock,reset=>reset,s=>p(174)(64),cout=>p(175)(65));
FA_ff_3009:FAff port map(x=>p(69)(65),y=>p(70)(65),Cin=>p(71)(65),clock=>clock,reset=>reset,s=>p(174)(65),cout=>p(175)(66));
FA_ff_3010:FAff port map(x=>p(69)(66),y=>p(70)(66),Cin=>p(71)(66),clock=>clock,reset=>reset,s=>p(174)(66),cout=>p(175)(67));
FA_ff_3011:FAff port map(x=>p(69)(67),y=>p(70)(67),Cin=>p(71)(67),clock=>clock,reset=>reset,s=>p(174)(67),cout=>p(175)(68));
FA_ff_3012:FAff port map(x=>p(69)(68),y=>p(70)(68),Cin=>p(71)(68),clock=>clock,reset=>reset,s=>p(174)(68),cout=>p(175)(69));
FA_ff_3013:FAff port map(x=>p(69)(69),y=>p(70)(69),Cin=>p(71)(69),clock=>clock,reset=>reset,s=>p(174)(69),cout=>p(175)(70));
FA_ff_3014:FAff port map(x=>p(69)(70),y=>p(70)(70),Cin=>p(71)(70),clock=>clock,reset=>reset,s=>p(174)(70),cout=>p(175)(71));
FA_ff_3015:FAff port map(x=>p(69)(71),y=>p(70)(71),Cin=>p(71)(71),clock=>clock,reset=>reset,s=>p(174)(71),cout=>p(175)(72));
FA_ff_3016:FAff port map(x=>p(69)(72),y=>p(70)(72),Cin=>p(71)(72),clock=>clock,reset=>reset,s=>p(174)(72),cout=>p(175)(73));
FA_ff_3017:FAff port map(x=>p(69)(73),y=>p(70)(73),Cin=>p(71)(73),clock=>clock,reset=>reset,s=>p(174)(73),cout=>p(175)(74));
FA_ff_3018:FAff port map(x=>p(69)(74),y=>p(70)(74),Cin=>p(71)(74),clock=>clock,reset=>reset,s=>p(174)(74),cout=>p(175)(75));
FA_ff_3019:FAff port map(x=>p(69)(75),y=>p(70)(75),Cin=>p(71)(75),clock=>clock,reset=>reset,s=>p(174)(75),cout=>p(175)(76));
FA_ff_3020:FAff port map(x=>p(69)(76),y=>p(70)(76),Cin=>p(71)(76),clock=>clock,reset=>reset,s=>p(174)(76),cout=>p(175)(77));
FA_ff_3021:FAff port map(x=>p(69)(77),y=>p(70)(77),Cin=>p(71)(77),clock=>clock,reset=>reset,s=>p(174)(77),cout=>p(175)(78));
FA_ff_3022:FAff port map(x=>p(69)(78),y=>p(70)(78),Cin=>p(71)(78),clock=>clock,reset=>reset,s=>p(174)(78),cout=>p(175)(79));
FA_ff_3023:FAff port map(x=>p(69)(79),y=>p(70)(79),Cin=>p(71)(79),clock=>clock,reset=>reset,s=>p(174)(79),cout=>p(175)(80));
FA_ff_3024:FAff port map(x=>p(69)(80),y=>p(70)(80),Cin=>p(71)(80),clock=>clock,reset=>reset,s=>p(174)(80),cout=>p(175)(81));
FA_ff_3025:FAff port map(x=>p(69)(81),y=>p(70)(81),Cin=>p(71)(81),clock=>clock,reset=>reset,s=>p(174)(81),cout=>p(175)(82));
FA_ff_3026:FAff port map(x=>p(69)(82),y=>p(70)(82),Cin=>p(71)(82),clock=>clock,reset=>reset,s=>p(174)(82),cout=>p(175)(83));
FA_ff_3027:FAff port map(x=>p(69)(83),y=>p(70)(83),Cin=>p(71)(83),clock=>clock,reset=>reset,s=>p(174)(83),cout=>p(175)(84));
FA_ff_3028:FAff port map(x=>p(69)(84),y=>p(70)(84),Cin=>p(71)(84),clock=>clock,reset=>reset,s=>p(174)(84),cout=>p(175)(85));
FA_ff_3029:FAff port map(x=>p(69)(85),y=>p(70)(85),Cin=>p(71)(85),clock=>clock,reset=>reset,s=>p(174)(85),cout=>p(175)(86));
FA_ff_3030:FAff port map(x=>p(69)(86),y=>p(70)(86),Cin=>p(71)(86),clock=>clock,reset=>reset,s=>p(174)(86),cout=>p(175)(87));
FA_ff_3031:FAff port map(x=>p(69)(87),y=>p(70)(87),Cin=>p(71)(87),clock=>clock,reset=>reset,s=>p(174)(87),cout=>p(175)(88));
FA_ff_3032:FAff port map(x=>p(69)(88),y=>p(70)(88),Cin=>p(71)(88),clock=>clock,reset=>reset,s=>p(174)(88),cout=>p(175)(89));
FA_ff_3033:FAff port map(x=>p(69)(89),y=>p(70)(89),Cin=>p(71)(89),clock=>clock,reset=>reset,s=>p(174)(89),cout=>p(175)(90));
FA_ff_3034:FAff port map(x=>p(69)(90),y=>p(70)(90),Cin=>p(71)(90),clock=>clock,reset=>reset,s=>p(174)(90),cout=>p(175)(91));
FA_ff_3035:FAff port map(x=>p(69)(91),y=>p(70)(91),Cin=>p(71)(91),clock=>clock,reset=>reset,s=>p(174)(91),cout=>p(175)(92));
FA_ff_3036:FAff port map(x=>p(69)(92),y=>p(70)(92),Cin=>p(71)(92),clock=>clock,reset=>reset,s=>p(174)(92),cout=>p(175)(93));
FA_ff_3037:FAff port map(x=>p(69)(93),y=>p(70)(93),Cin=>p(71)(93),clock=>clock,reset=>reset,s=>p(174)(93),cout=>p(175)(94));
FA_ff_3038:FAff port map(x=>p(69)(94),y=>p(70)(94),Cin=>p(71)(94),clock=>clock,reset=>reset,s=>p(174)(94),cout=>p(175)(95));
FA_ff_3039:FAff port map(x=>p(69)(95),y=>p(70)(95),Cin=>p(71)(95),clock=>clock,reset=>reset,s=>p(174)(95),cout=>p(175)(96));
FA_ff_3040:FAff port map(x=>p(69)(96),y=>p(70)(96),Cin=>p(71)(96),clock=>clock,reset=>reset,s=>p(174)(96),cout=>p(175)(97));
FA_ff_3041:FAff port map(x=>p(69)(97),y=>p(70)(97),Cin=>p(71)(97),clock=>clock,reset=>reset,s=>p(174)(97),cout=>p(175)(98));
FA_ff_3042:FAff port map(x=>p(69)(98),y=>p(70)(98),Cin=>p(71)(98),clock=>clock,reset=>reset,s=>p(174)(98),cout=>p(175)(99));
FA_ff_3043:FAff port map(x=>p(69)(99),y=>p(70)(99),Cin=>p(71)(99),clock=>clock,reset=>reset,s=>p(174)(99),cout=>p(175)(100));
FA_ff_3044:FAff port map(x=>p(69)(100),y=>p(70)(100),Cin=>p(71)(100),clock=>clock,reset=>reset,s=>p(174)(100),cout=>p(175)(101));
FA_ff_3045:FAff port map(x=>p(69)(101),y=>p(70)(101),Cin=>p(71)(101),clock=>clock,reset=>reset,s=>p(174)(101),cout=>p(175)(102));
FA_ff_3046:FAff port map(x=>p(69)(102),y=>p(70)(102),Cin=>p(71)(102),clock=>clock,reset=>reset,s=>p(174)(102),cout=>p(175)(103));
FA_ff_3047:FAff port map(x=>p(69)(103),y=>p(70)(103),Cin=>p(71)(103),clock=>clock,reset=>reset,s=>p(174)(103),cout=>p(175)(104));
FA_ff_3048:FAff port map(x=>p(69)(104),y=>p(70)(104),Cin=>p(71)(104),clock=>clock,reset=>reset,s=>p(174)(104),cout=>p(175)(105));
FA_ff_3049:FAff port map(x=>p(69)(105),y=>p(70)(105),Cin=>p(71)(105),clock=>clock,reset=>reset,s=>p(174)(105),cout=>p(175)(106));
FA_ff_3050:FAff port map(x=>p(69)(106),y=>p(70)(106),Cin=>p(71)(106),clock=>clock,reset=>reset,s=>p(174)(106),cout=>p(175)(107));
FA_ff_3051:FAff port map(x=>p(69)(107),y=>p(70)(107),Cin=>p(71)(107),clock=>clock,reset=>reset,s=>p(174)(107),cout=>p(175)(108));
FA_ff_3052:FAff port map(x=>p(69)(108),y=>p(70)(108),Cin=>p(71)(108),clock=>clock,reset=>reset,s=>p(174)(108),cout=>p(175)(109));
FA_ff_3053:FAff port map(x=>p(69)(109),y=>p(70)(109),Cin=>p(71)(109),clock=>clock,reset=>reset,s=>p(174)(109),cout=>p(175)(110));
FA_ff_3054:FAff port map(x=>p(69)(110),y=>p(70)(110),Cin=>p(71)(110),clock=>clock,reset=>reset,s=>p(174)(110),cout=>p(175)(111));
FA_ff_3055:FAff port map(x=>p(69)(111),y=>p(70)(111),Cin=>p(71)(111),clock=>clock,reset=>reset,s=>p(174)(111),cout=>p(175)(112));
FA_ff_3056:FAff port map(x=>p(69)(112),y=>p(70)(112),Cin=>p(71)(112),clock=>clock,reset=>reset,s=>p(174)(112),cout=>p(175)(113));
FA_ff_3057:FAff port map(x=>p(69)(113),y=>p(70)(113),Cin=>p(71)(113),clock=>clock,reset=>reset,s=>p(174)(113),cout=>p(175)(114));
FA_ff_3058:FAff port map(x=>p(69)(114),y=>p(70)(114),Cin=>p(71)(114),clock=>clock,reset=>reset,s=>p(174)(114),cout=>p(175)(115));
FA_ff_3059:FAff port map(x=>p(69)(115),y=>p(70)(115),Cin=>p(71)(115),clock=>clock,reset=>reset,s=>p(174)(115),cout=>p(175)(116));
FA_ff_3060:FAff port map(x=>p(69)(116),y=>p(70)(116),Cin=>p(71)(116),clock=>clock,reset=>reset,s=>p(174)(116),cout=>p(175)(117));
FA_ff_3061:FAff port map(x=>p(69)(117),y=>p(70)(117),Cin=>p(71)(117),clock=>clock,reset=>reset,s=>p(174)(117),cout=>p(175)(118));
FA_ff_3062:FAff port map(x=>p(69)(118),y=>p(70)(118),Cin=>p(71)(118),clock=>clock,reset=>reset,s=>p(174)(118),cout=>p(175)(119));
FA_ff_3063:FAff port map(x=>p(69)(119),y=>p(70)(119),Cin=>p(71)(119),clock=>clock,reset=>reset,s=>p(174)(119),cout=>p(175)(120));
FA_ff_3064:FAff port map(x=>p(69)(120),y=>p(70)(120),Cin=>p(71)(120),clock=>clock,reset=>reset,s=>p(174)(120),cout=>p(175)(121));
FA_ff_3065:FAff port map(x=>p(69)(121),y=>p(70)(121),Cin=>p(71)(121),clock=>clock,reset=>reset,s=>p(174)(121),cout=>p(175)(122));
FA_ff_3066:FAff port map(x=>p(69)(122),y=>p(70)(122),Cin=>p(71)(122),clock=>clock,reset=>reset,s=>p(174)(122),cout=>p(175)(123));
FA_ff_3067:FAff port map(x=>p(69)(123),y=>p(70)(123),Cin=>p(71)(123),clock=>clock,reset=>reset,s=>p(174)(123),cout=>p(175)(124));
FA_ff_3068:FAff port map(x=>p(69)(124),y=>p(70)(124),Cin=>p(71)(124),clock=>clock,reset=>reset,s=>p(174)(124),cout=>p(175)(125));
FA_ff_3069:FAff port map(x=>p(69)(125),y=>p(70)(125),Cin=>p(71)(125),clock=>clock,reset=>reset,s=>p(174)(125),cout=>p(175)(126));
FA_ff_3070:FAff port map(x=>p(69)(126),y=>p(70)(126),Cin=>p(71)(126),clock=>clock,reset=>reset,s=>p(174)(126),cout=>p(175)(127));
FA_ff_3071:FAff port map(x=>p(69)(127),y=>p(70)(127),Cin=>p(71)(127),clock=>clock,reset=>reset,s=>p(174)(127),cout=>p(175)(128));
FA_ff_3072:FAff port map(x=>p(72)(0),y=>p(73)(0),Cin=>p(74)(0),clock=>clock,reset=>reset,s=>p(176)(0),cout=>p(177)(1));
FA_ff_3073:FAff port map(x=>p(72)(1),y=>p(73)(1),Cin=>p(74)(1),clock=>clock,reset=>reset,s=>p(176)(1),cout=>p(177)(2));
FA_ff_3074:FAff port map(x=>p(72)(2),y=>p(73)(2),Cin=>p(74)(2),clock=>clock,reset=>reset,s=>p(176)(2),cout=>p(177)(3));
FA_ff_3075:FAff port map(x=>p(72)(3),y=>p(73)(3),Cin=>p(74)(3),clock=>clock,reset=>reset,s=>p(176)(3),cout=>p(177)(4));
FA_ff_3076:FAff port map(x=>p(72)(4),y=>p(73)(4),Cin=>p(74)(4),clock=>clock,reset=>reset,s=>p(176)(4),cout=>p(177)(5));
FA_ff_3077:FAff port map(x=>p(72)(5),y=>p(73)(5),Cin=>p(74)(5),clock=>clock,reset=>reset,s=>p(176)(5),cout=>p(177)(6));
FA_ff_3078:FAff port map(x=>p(72)(6),y=>p(73)(6),Cin=>p(74)(6),clock=>clock,reset=>reset,s=>p(176)(6),cout=>p(177)(7));
FA_ff_3079:FAff port map(x=>p(72)(7),y=>p(73)(7),Cin=>p(74)(7),clock=>clock,reset=>reset,s=>p(176)(7),cout=>p(177)(8));
FA_ff_3080:FAff port map(x=>p(72)(8),y=>p(73)(8),Cin=>p(74)(8),clock=>clock,reset=>reset,s=>p(176)(8),cout=>p(177)(9));
FA_ff_3081:FAff port map(x=>p(72)(9),y=>p(73)(9),Cin=>p(74)(9),clock=>clock,reset=>reset,s=>p(176)(9),cout=>p(177)(10));
FA_ff_3082:FAff port map(x=>p(72)(10),y=>p(73)(10),Cin=>p(74)(10),clock=>clock,reset=>reset,s=>p(176)(10),cout=>p(177)(11));
FA_ff_3083:FAff port map(x=>p(72)(11),y=>p(73)(11),Cin=>p(74)(11),clock=>clock,reset=>reset,s=>p(176)(11),cout=>p(177)(12));
FA_ff_3084:FAff port map(x=>p(72)(12),y=>p(73)(12),Cin=>p(74)(12),clock=>clock,reset=>reset,s=>p(176)(12),cout=>p(177)(13));
FA_ff_3085:FAff port map(x=>p(72)(13),y=>p(73)(13),Cin=>p(74)(13),clock=>clock,reset=>reset,s=>p(176)(13),cout=>p(177)(14));
FA_ff_3086:FAff port map(x=>p(72)(14),y=>p(73)(14),Cin=>p(74)(14),clock=>clock,reset=>reset,s=>p(176)(14),cout=>p(177)(15));
FA_ff_3087:FAff port map(x=>p(72)(15),y=>p(73)(15),Cin=>p(74)(15),clock=>clock,reset=>reset,s=>p(176)(15),cout=>p(177)(16));
FA_ff_3088:FAff port map(x=>p(72)(16),y=>p(73)(16),Cin=>p(74)(16),clock=>clock,reset=>reset,s=>p(176)(16),cout=>p(177)(17));
FA_ff_3089:FAff port map(x=>p(72)(17),y=>p(73)(17),Cin=>p(74)(17),clock=>clock,reset=>reset,s=>p(176)(17),cout=>p(177)(18));
FA_ff_3090:FAff port map(x=>p(72)(18),y=>p(73)(18),Cin=>p(74)(18),clock=>clock,reset=>reset,s=>p(176)(18),cout=>p(177)(19));
FA_ff_3091:FAff port map(x=>p(72)(19),y=>p(73)(19),Cin=>p(74)(19),clock=>clock,reset=>reset,s=>p(176)(19),cout=>p(177)(20));
FA_ff_3092:FAff port map(x=>p(72)(20),y=>p(73)(20),Cin=>p(74)(20),clock=>clock,reset=>reset,s=>p(176)(20),cout=>p(177)(21));
FA_ff_3093:FAff port map(x=>p(72)(21),y=>p(73)(21),Cin=>p(74)(21),clock=>clock,reset=>reset,s=>p(176)(21),cout=>p(177)(22));
FA_ff_3094:FAff port map(x=>p(72)(22),y=>p(73)(22),Cin=>p(74)(22),clock=>clock,reset=>reset,s=>p(176)(22),cout=>p(177)(23));
FA_ff_3095:FAff port map(x=>p(72)(23),y=>p(73)(23),Cin=>p(74)(23),clock=>clock,reset=>reset,s=>p(176)(23),cout=>p(177)(24));
FA_ff_3096:FAff port map(x=>p(72)(24),y=>p(73)(24),Cin=>p(74)(24),clock=>clock,reset=>reset,s=>p(176)(24),cout=>p(177)(25));
FA_ff_3097:FAff port map(x=>p(72)(25),y=>p(73)(25),Cin=>p(74)(25),clock=>clock,reset=>reset,s=>p(176)(25),cout=>p(177)(26));
FA_ff_3098:FAff port map(x=>p(72)(26),y=>p(73)(26),Cin=>p(74)(26),clock=>clock,reset=>reset,s=>p(176)(26),cout=>p(177)(27));
FA_ff_3099:FAff port map(x=>p(72)(27),y=>p(73)(27),Cin=>p(74)(27),clock=>clock,reset=>reset,s=>p(176)(27),cout=>p(177)(28));
FA_ff_3100:FAff port map(x=>p(72)(28),y=>p(73)(28),Cin=>p(74)(28),clock=>clock,reset=>reset,s=>p(176)(28),cout=>p(177)(29));
FA_ff_3101:FAff port map(x=>p(72)(29),y=>p(73)(29),Cin=>p(74)(29),clock=>clock,reset=>reset,s=>p(176)(29),cout=>p(177)(30));
FA_ff_3102:FAff port map(x=>p(72)(30),y=>p(73)(30),Cin=>p(74)(30),clock=>clock,reset=>reset,s=>p(176)(30),cout=>p(177)(31));
FA_ff_3103:FAff port map(x=>p(72)(31),y=>p(73)(31),Cin=>p(74)(31),clock=>clock,reset=>reset,s=>p(176)(31),cout=>p(177)(32));
FA_ff_3104:FAff port map(x=>p(72)(32),y=>p(73)(32),Cin=>p(74)(32),clock=>clock,reset=>reset,s=>p(176)(32),cout=>p(177)(33));
FA_ff_3105:FAff port map(x=>p(72)(33),y=>p(73)(33),Cin=>p(74)(33),clock=>clock,reset=>reset,s=>p(176)(33),cout=>p(177)(34));
FA_ff_3106:FAff port map(x=>p(72)(34),y=>p(73)(34),Cin=>p(74)(34),clock=>clock,reset=>reset,s=>p(176)(34),cout=>p(177)(35));
FA_ff_3107:FAff port map(x=>p(72)(35),y=>p(73)(35),Cin=>p(74)(35),clock=>clock,reset=>reset,s=>p(176)(35),cout=>p(177)(36));
FA_ff_3108:FAff port map(x=>p(72)(36),y=>p(73)(36),Cin=>p(74)(36),clock=>clock,reset=>reset,s=>p(176)(36),cout=>p(177)(37));
FA_ff_3109:FAff port map(x=>p(72)(37),y=>p(73)(37),Cin=>p(74)(37),clock=>clock,reset=>reset,s=>p(176)(37),cout=>p(177)(38));
FA_ff_3110:FAff port map(x=>p(72)(38),y=>p(73)(38),Cin=>p(74)(38),clock=>clock,reset=>reset,s=>p(176)(38),cout=>p(177)(39));
FA_ff_3111:FAff port map(x=>p(72)(39),y=>p(73)(39),Cin=>p(74)(39),clock=>clock,reset=>reset,s=>p(176)(39),cout=>p(177)(40));
FA_ff_3112:FAff port map(x=>p(72)(40),y=>p(73)(40),Cin=>p(74)(40),clock=>clock,reset=>reset,s=>p(176)(40),cout=>p(177)(41));
FA_ff_3113:FAff port map(x=>p(72)(41),y=>p(73)(41),Cin=>p(74)(41),clock=>clock,reset=>reset,s=>p(176)(41),cout=>p(177)(42));
FA_ff_3114:FAff port map(x=>p(72)(42),y=>p(73)(42),Cin=>p(74)(42),clock=>clock,reset=>reset,s=>p(176)(42),cout=>p(177)(43));
FA_ff_3115:FAff port map(x=>p(72)(43),y=>p(73)(43),Cin=>p(74)(43),clock=>clock,reset=>reset,s=>p(176)(43),cout=>p(177)(44));
FA_ff_3116:FAff port map(x=>p(72)(44),y=>p(73)(44),Cin=>p(74)(44),clock=>clock,reset=>reset,s=>p(176)(44),cout=>p(177)(45));
FA_ff_3117:FAff port map(x=>p(72)(45),y=>p(73)(45),Cin=>p(74)(45),clock=>clock,reset=>reset,s=>p(176)(45),cout=>p(177)(46));
FA_ff_3118:FAff port map(x=>p(72)(46),y=>p(73)(46),Cin=>p(74)(46),clock=>clock,reset=>reset,s=>p(176)(46),cout=>p(177)(47));
FA_ff_3119:FAff port map(x=>p(72)(47),y=>p(73)(47),Cin=>p(74)(47),clock=>clock,reset=>reset,s=>p(176)(47),cout=>p(177)(48));
FA_ff_3120:FAff port map(x=>p(72)(48),y=>p(73)(48),Cin=>p(74)(48),clock=>clock,reset=>reset,s=>p(176)(48),cout=>p(177)(49));
FA_ff_3121:FAff port map(x=>p(72)(49),y=>p(73)(49),Cin=>p(74)(49),clock=>clock,reset=>reset,s=>p(176)(49),cout=>p(177)(50));
FA_ff_3122:FAff port map(x=>p(72)(50),y=>p(73)(50),Cin=>p(74)(50),clock=>clock,reset=>reset,s=>p(176)(50),cout=>p(177)(51));
FA_ff_3123:FAff port map(x=>p(72)(51),y=>p(73)(51),Cin=>p(74)(51),clock=>clock,reset=>reset,s=>p(176)(51),cout=>p(177)(52));
FA_ff_3124:FAff port map(x=>p(72)(52),y=>p(73)(52),Cin=>p(74)(52),clock=>clock,reset=>reset,s=>p(176)(52),cout=>p(177)(53));
FA_ff_3125:FAff port map(x=>p(72)(53),y=>p(73)(53),Cin=>p(74)(53),clock=>clock,reset=>reset,s=>p(176)(53),cout=>p(177)(54));
FA_ff_3126:FAff port map(x=>p(72)(54),y=>p(73)(54),Cin=>p(74)(54),clock=>clock,reset=>reset,s=>p(176)(54),cout=>p(177)(55));
FA_ff_3127:FAff port map(x=>p(72)(55),y=>p(73)(55),Cin=>p(74)(55),clock=>clock,reset=>reset,s=>p(176)(55),cout=>p(177)(56));
FA_ff_3128:FAff port map(x=>p(72)(56),y=>p(73)(56),Cin=>p(74)(56),clock=>clock,reset=>reset,s=>p(176)(56),cout=>p(177)(57));
FA_ff_3129:FAff port map(x=>p(72)(57),y=>p(73)(57),Cin=>p(74)(57),clock=>clock,reset=>reset,s=>p(176)(57),cout=>p(177)(58));
FA_ff_3130:FAff port map(x=>p(72)(58),y=>p(73)(58),Cin=>p(74)(58),clock=>clock,reset=>reset,s=>p(176)(58),cout=>p(177)(59));
FA_ff_3131:FAff port map(x=>p(72)(59),y=>p(73)(59),Cin=>p(74)(59),clock=>clock,reset=>reset,s=>p(176)(59),cout=>p(177)(60));
FA_ff_3132:FAff port map(x=>p(72)(60),y=>p(73)(60),Cin=>p(74)(60),clock=>clock,reset=>reset,s=>p(176)(60),cout=>p(177)(61));
FA_ff_3133:FAff port map(x=>p(72)(61),y=>p(73)(61),Cin=>p(74)(61),clock=>clock,reset=>reset,s=>p(176)(61),cout=>p(177)(62));
FA_ff_3134:FAff port map(x=>p(72)(62),y=>p(73)(62),Cin=>p(74)(62),clock=>clock,reset=>reset,s=>p(176)(62),cout=>p(177)(63));
FA_ff_3135:FAff port map(x=>p(72)(63),y=>p(73)(63),Cin=>p(74)(63),clock=>clock,reset=>reset,s=>p(176)(63),cout=>p(177)(64));
FA_ff_3136:FAff port map(x=>p(72)(64),y=>p(73)(64),Cin=>p(74)(64),clock=>clock,reset=>reset,s=>p(176)(64),cout=>p(177)(65));
FA_ff_3137:FAff port map(x=>p(72)(65),y=>p(73)(65),Cin=>p(74)(65),clock=>clock,reset=>reset,s=>p(176)(65),cout=>p(177)(66));
FA_ff_3138:FAff port map(x=>p(72)(66),y=>p(73)(66),Cin=>p(74)(66),clock=>clock,reset=>reset,s=>p(176)(66),cout=>p(177)(67));
FA_ff_3139:FAff port map(x=>p(72)(67),y=>p(73)(67),Cin=>p(74)(67),clock=>clock,reset=>reset,s=>p(176)(67),cout=>p(177)(68));
FA_ff_3140:FAff port map(x=>p(72)(68),y=>p(73)(68),Cin=>p(74)(68),clock=>clock,reset=>reset,s=>p(176)(68),cout=>p(177)(69));
FA_ff_3141:FAff port map(x=>p(72)(69),y=>p(73)(69),Cin=>p(74)(69),clock=>clock,reset=>reset,s=>p(176)(69),cout=>p(177)(70));
FA_ff_3142:FAff port map(x=>p(72)(70),y=>p(73)(70),Cin=>p(74)(70),clock=>clock,reset=>reset,s=>p(176)(70),cout=>p(177)(71));
FA_ff_3143:FAff port map(x=>p(72)(71),y=>p(73)(71),Cin=>p(74)(71),clock=>clock,reset=>reset,s=>p(176)(71),cout=>p(177)(72));
FA_ff_3144:FAff port map(x=>p(72)(72),y=>p(73)(72),Cin=>p(74)(72),clock=>clock,reset=>reset,s=>p(176)(72),cout=>p(177)(73));
FA_ff_3145:FAff port map(x=>p(72)(73),y=>p(73)(73),Cin=>p(74)(73),clock=>clock,reset=>reset,s=>p(176)(73),cout=>p(177)(74));
FA_ff_3146:FAff port map(x=>p(72)(74),y=>p(73)(74),Cin=>p(74)(74),clock=>clock,reset=>reset,s=>p(176)(74),cout=>p(177)(75));
FA_ff_3147:FAff port map(x=>p(72)(75),y=>p(73)(75),Cin=>p(74)(75),clock=>clock,reset=>reset,s=>p(176)(75),cout=>p(177)(76));
FA_ff_3148:FAff port map(x=>p(72)(76),y=>p(73)(76),Cin=>p(74)(76),clock=>clock,reset=>reset,s=>p(176)(76),cout=>p(177)(77));
FA_ff_3149:FAff port map(x=>p(72)(77),y=>p(73)(77),Cin=>p(74)(77),clock=>clock,reset=>reset,s=>p(176)(77),cout=>p(177)(78));
FA_ff_3150:FAff port map(x=>p(72)(78),y=>p(73)(78),Cin=>p(74)(78),clock=>clock,reset=>reset,s=>p(176)(78),cout=>p(177)(79));
FA_ff_3151:FAff port map(x=>p(72)(79),y=>p(73)(79),Cin=>p(74)(79),clock=>clock,reset=>reset,s=>p(176)(79),cout=>p(177)(80));
FA_ff_3152:FAff port map(x=>p(72)(80),y=>p(73)(80),Cin=>p(74)(80),clock=>clock,reset=>reset,s=>p(176)(80),cout=>p(177)(81));
FA_ff_3153:FAff port map(x=>p(72)(81),y=>p(73)(81),Cin=>p(74)(81),clock=>clock,reset=>reset,s=>p(176)(81),cout=>p(177)(82));
FA_ff_3154:FAff port map(x=>p(72)(82),y=>p(73)(82),Cin=>p(74)(82),clock=>clock,reset=>reset,s=>p(176)(82),cout=>p(177)(83));
FA_ff_3155:FAff port map(x=>p(72)(83),y=>p(73)(83),Cin=>p(74)(83),clock=>clock,reset=>reset,s=>p(176)(83),cout=>p(177)(84));
FA_ff_3156:FAff port map(x=>p(72)(84),y=>p(73)(84),Cin=>p(74)(84),clock=>clock,reset=>reset,s=>p(176)(84),cout=>p(177)(85));
FA_ff_3157:FAff port map(x=>p(72)(85),y=>p(73)(85),Cin=>p(74)(85),clock=>clock,reset=>reset,s=>p(176)(85),cout=>p(177)(86));
FA_ff_3158:FAff port map(x=>p(72)(86),y=>p(73)(86),Cin=>p(74)(86),clock=>clock,reset=>reset,s=>p(176)(86),cout=>p(177)(87));
FA_ff_3159:FAff port map(x=>p(72)(87),y=>p(73)(87),Cin=>p(74)(87),clock=>clock,reset=>reset,s=>p(176)(87),cout=>p(177)(88));
FA_ff_3160:FAff port map(x=>p(72)(88),y=>p(73)(88),Cin=>p(74)(88),clock=>clock,reset=>reset,s=>p(176)(88),cout=>p(177)(89));
FA_ff_3161:FAff port map(x=>p(72)(89),y=>p(73)(89),Cin=>p(74)(89),clock=>clock,reset=>reset,s=>p(176)(89),cout=>p(177)(90));
FA_ff_3162:FAff port map(x=>p(72)(90),y=>p(73)(90),Cin=>p(74)(90),clock=>clock,reset=>reset,s=>p(176)(90),cout=>p(177)(91));
FA_ff_3163:FAff port map(x=>p(72)(91),y=>p(73)(91),Cin=>p(74)(91),clock=>clock,reset=>reset,s=>p(176)(91),cout=>p(177)(92));
FA_ff_3164:FAff port map(x=>p(72)(92),y=>p(73)(92),Cin=>p(74)(92),clock=>clock,reset=>reset,s=>p(176)(92),cout=>p(177)(93));
FA_ff_3165:FAff port map(x=>p(72)(93),y=>p(73)(93),Cin=>p(74)(93),clock=>clock,reset=>reset,s=>p(176)(93),cout=>p(177)(94));
FA_ff_3166:FAff port map(x=>p(72)(94),y=>p(73)(94),Cin=>p(74)(94),clock=>clock,reset=>reset,s=>p(176)(94),cout=>p(177)(95));
FA_ff_3167:FAff port map(x=>p(72)(95),y=>p(73)(95),Cin=>p(74)(95),clock=>clock,reset=>reset,s=>p(176)(95),cout=>p(177)(96));
FA_ff_3168:FAff port map(x=>p(72)(96),y=>p(73)(96),Cin=>p(74)(96),clock=>clock,reset=>reset,s=>p(176)(96),cout=>p(177)(97));
FA_ff_3169:FAff port map(x=>p(72)(97),y=>p(73)(97),Cin=>p(74)(97),clock=>clock,reset=>reset,s=>p(176)(97),cout=>p(177)(98));
FA_ff_3170:FAff port map(x=>p(72)(98),y=>p(73)(98),Cin=>p(74)(98),clock=>clock,reset=>reset,s=>p(176)(98),cout=>p(177)(99));
FA_ff_3171:FAff port map(x=>p(72)(99),y=>p(73)(99),Cin=>p(74)(99),clock=>clock,reset=>reset,s=>p(176)(99),cout=>p(177)(100));
FA_ff_3172:FAff port map(x=>p(72)(100),y=>p(73)(100),Cin=>p(74)(100),clock=>clock,reset=>reset,s=>p(176)(100),cout=>p(177)(101));
FA_ff_3173:FAff port map(x=>p(72)(101),y=>p(73)(101),Cin=>p(74)(101),clock=>clock,reset=>reset,s=>p(176)(101),cout=>p(177)(102));
FA_ff_3174:FAff port map(x=>p(72)(102),y=>p(73)(102),Cin=>p(74)(102),clock=>clock,reset=>reset,s=>p(176)(102),cout=>p(177)(103));
FA_ff_3175:FAff port map(x=>p(72)(103),y=>p(73)(103),Cin=>p(74)(103),clock=>clock,reset=>reset,s=>p(176)(103),cout=>p(177)(104));
FA_ff_3176:FAff port map(x=>p(72)(104),y=>p(73)(104),Cin=>p(74)(104),clock=>clock,reset=>reset,s=>p(176)(104),cout=>p(177)(105));
FA_ff_3177:FAff port map(x=>p(72)(105),y=>p(73)(105),Cin=>p(74)(105),clock=>clock,reset=>reset,s=>p(176)(105),cout=>p(177)(106));
FA_ff_3178:FAff port map(x=>p(72)(106),y=>p(73)(106),Cin=>p(74)(106),clock=>clock,reset=>reset,s=>p(176)(106),cout=>p(177)(107));
FA_ff_3179:FAff port map(x=>p(72)(107),y=>p(73)(107),Cin=>p(74)(107),clock=>clock,reset=>reset,s=>p(176)(107),cout=>p(177)(108));
FA_ff_3180:FAff port map(x=>p(72)(108),y=>p(73)(108),Cin=>p(74)(108),clock=>clock,reset=>reset,s=>p(176)(108),cout=>p(177)(109));
FA_ff_3181:FAff port map(x=>p(72)(109),y=>p(73)(109),Cin=>p(74)(109),clock=>clock,reset=>reset,s=>p(176)(109),cout=>p(177)(110));
FA_ff_3182:FAff port map(x=>p(72)(110),y=>p(73)(110),Cin=>p(74)(110),clock=>clock,reset=>reset,s=>p(176)(110),cout=>p(177)(111));
FA_ff_3183:FAff port map(x=>p(72)(111),y=>p(73)(111),Cin=>p(74)(111),clock=>clock,reset=>reset,s=>p(176)(111),cout=>p(177)(112));
FA_ff_3184:FAff port map(x=>p(72)(112),y=>p(73)(112),Cin=>p(74)(112),clock=>clock,reset=>reset,s=>p(176)(112),cout=>p(177)(113));
FA_ff_3185:FAff port map(x=>p(72)(113),y=>p(73)(113),Cin=>p(74)(113),clock=>clock,reset=>reset,s=>p(176)(113),cout=>p(177)(114));
FA_ff_3186:FAff port map(x=>p(72)(114),y=>p(73)(114),Cin=>p(74)(114),clock=>clock,reset=>reset,s=>p(176)(114),cout=>p(177)(115));
FA_ff_3187:FAff port map(x=>p(72)(115),y=>p(73)(115),Cin=>p(74)(115),clock=>clock,reset=>reset,s=>p(176)(115),cout=>p(177)(116));
FA_ff_3188:FAff port map(x=>p(72)(116),y=>p(73)(116),Cin=>p(74)(116),clock=>clock,reset=>reset,s=>p(176)(116),cout=>p(177)(117));
FA_ff_3189:FAff port map(x=>p(72)(117),y=>p(73)(117),Cin=>p(74)(117),clock=>clock,reset=>reset,s=>p(176)(117),cout=>p(177)(118));
FA_ff_3190:FAff port map(x=>p(72)(118),y=>p(73)(118),Cin=>p(74)(118),clock=>clock,reset=>reset,s=>p(176)(118),cout=>p(177)(119));
FA_ff_3191:FAff port map(x=>p(72)(119),y=>p(73)(119),Cin=>p(74)(119),clock=>clock,reset=>reset,s=>p(176)(119),cout=>p(177)(120));
FA_ff_3192:FAff port map(x=>p(72)(120),y=>p(73)(120),Cin=>p(74)(120),clock=>clock,reset=>reset,s=>p(176)(120),cout=>p(177)(121));
FA_ff_3193:FAff port map(x=>p(72)(121),y=>p(73)(121),Cin=>p(74)(121),clock=>clock,reset=>reset,s=>p(176)(121),cout=>p(177)(122));
FA_ff_3194:FAff port map(x=>p(72)(122),y=>p(73)(122),Cin=>p(74)(122),clock=>clock,reset=>reset,s=>p(176)(122),cout=>p(177)(123));
FA_ff_3195:FAff port map(x=>p(72)(123),y=>p(73)(123),Cin=>p(74)(123),clock=>clock,reset=>reset,s=>p(176)(123),cout=>p(177)(124));
FA_ff_3196:FAff port map(x=>p(72)(124),y=>p(73)(124),Cin=>p(74)(124),clock=>clock,reset=>reset,s=>p(176)(124),cout=>p(177)(125));
FA_ff_3197:FAff port map(x=>p(72)(125),y=>p(73)(125),Cin=>p(74)(125),clock=>clock,reset=>reset,s=>p(176)(125),cout=>p(177)(126));
FA_ff_3198:FAff port map(x=>p(72)(126),y=>p(73)(126),Cin=>p(74)(126),clock=>clock,reset=>reset,s=>p(176)(126),cout=>p(177)(127));
FA_ff_3199:FAff port map(x=>p(72)(127),y=>p(73)(127),Cin=>p(74)(127),clock=>clock,reset=>reset,s=>p(176)(127),cout=>p(177)(128));
FA_ff_3200:FAff port map(x=>p(75)(0),y=>p(76)(0),Cin=>p(77)(0),clock=>clock,reset=>reset,s=>p(178)(0),cout=>p(179)(1));
FA_ff_3201:FAff port map(x=>p(75)(1),y=>p(76)(1),Cin=>p(77)(1),clock=>clock,reset=>reset,s=>p(178)(1),cout=>p(179)(2));
FA_ff_3202:FAff port map(x=>p(75)(2),y=>p(76)(2),Cin=>p(77)(2),clock=>clock,reset=>reset,s=>p(178)(2),cout=>p(179)(3));
FA_ff_3203:FAff port map(x=>p(75)(3),y=>p(76)(3),Cin=>p(77)(3),clock=>clock,reset=>reset,s=>p(178)(3),cout=>p(179)(4));
FA_ff_3204:FAff port map(x=>p(75)(4),y=>p(76)(4),Cin=>p(77)(4),clock=>clock,reset=>reset,s=>p(178)(4),cout=>p(179)(5));
FA_ff_3205:FAff port map(x=>p(75)(5),y=>p(76)(5),Cin=>p(77)(5),clock=>clock,reset=>reset,s=>p(178)(5),cout=>p(179)(6));
FA_ff_3206:FAff port map(x=>p(75)(6),y=>p(76)(6),Cin=>p(77)(6),clock=>clock,reset=>reset,s=>p(178)(6),cout=>p(179)(7));
FA_ff_3207:FAff port map(x=>p(75)(7),y=>p(76)(7),Cin=>p(77)(7),clock=>clock,reset=>reset,s=>p(178)(7),cout=>p(179)(8));
FA_ff_3208:FAff port map(x=>p(75)(8),y=>p(76)(8),Cin=>p(77)(8),clock=>clock,reset=>reset,s=>p(178)(8),cout=>p(179)(9));
FA_ff_3209:FAff port map(x=>p(75)(9),y=>p(76)(9),Cin=>p(77)(9),clock=>clock,reset=>reset,s=>p(178)(9),cout=>p(179)(10));
FA_ff_3210:FAff port map(x=>p(75)(10),y=>p(76)(10),Cin=>p(77)(10),clock=>clock,reset=>reset,s=>p(178)(10),cout=>p(179)(11));
FA_ff_3211:FAff port map(x=>p(75)(11),y=>p(76)(11),Cin=>p(77)(11),clock=>clock,reset=>reset,s=>p(178)(11),cout=>p(179)(12));
FA_ff_3212:FAff port map(x=>p(75)(12),y=>p(76)(12),Cin=>p(77)(12),clock=>clock,reset=>reset,s=>p(178)(12),cout=>p(179)(13));
FA_ff_3213:FAff port map(x=>p(75)(13),y=>p(76)(13),Cin=>p(77)(13),clock=>clock,reset=>reset,s=>p(178)(13),cout=>p(179)(14));
FA_ff_3214:FAff port map(x=>p(75)(14),y=>p(76)(14),Cin=>p(77)(14),clock=>clock,reset=>reset,s=>p(178)(14),cout=>p(179)(15));
FA_ff_3215:FAff port map(x=>p(75)(15),y=>p(76)(15),Cin=>p(77)(15),clock=>clock,reset=>reset,s=>p(178)(15),cout=>p(179)(16));
FA_ff_3216:FAff port map(x=>p(75)(16),y=>p(76)(16),Cin=>p(77)(16),clock=>clock,reset=>reset,s=>p(178)(16),cout=>p(179)(17));
FA_ff_3217:FAff port map(x=>p(75)(17),y=>p(76)(17),Cin=>p(77)(17),clock=>clock,reset=>reset,s=>p(178)(17),cout=>p(179)(18));
FA_ff_3218:FAff port map(x=>p(75)(18),y=>p(76)(18),Cin=>p(77)(18),clock=>clock,reset=>reset,s=>p(178)(18),cout=>p(179)(19));
FA_ff_3219:FAff port map(x=>p(75)(19),y=>p(76)(19),Cin=>p(77)(19),clock=>clock,reset=>reset,s=>p(178)(19),cout=>p(179)(20));
FA_ff_3220:FAff port map(x=>p(75)(20),y=>p(76)(20),Cin=>p(77)(20),clock=>clock,reset=>reset,s=>p(178)(20),cout=>p(179)(21));
FA_ff_3221:FAff port map(x=>p(75)(21),y=>p(76)(21),Cin=>p(77)(21),clock=>clock,reset=>reset,s=>p(178)(21),cout=>p(179)(22));
FA_ff_3222:FAff port map(x=>p(75)(22),y=>p(76)(22),Cin=>p(77)(22),clock=>clock,reset=>reset,s=>p(178)(22),cout=>p(179)(23));
FA_ff_3223:FAff port map(x=>p(75)(23),y=>p(76)(23),Cin=>p(77)(23),clock=>clock,reset=>reset,s=>p(178)(23),cout=>p(179)(24));
FA_ff_3224:FAff port map(x=>p(75)(24),y=>p(76)(24),Cin=>p(77)(24),clock=>clock,reset=>reset,s=>p(178)(24),cout=>p(179)(25));
FA_ff_3225:FAff port map(x=>p(75)(25),y=>p(76)(25),Cin=>p(77)(25),clock=>clock,reset=>reset,s=>p(178)(25),cout=>p(179)(26));
FA_ff_3226:FAff port map(x=>p(75)(26),y=>p(76)(26),Cin=>p(77)(26),clock=>clock,reset=>reset,s=>p(178)(26),cout=>p(179)(27));
FA_ff_3227:FAff port map(x=>p(75)(27),y=>p(76)(27),Cin=>p(77)(27),clock=>clock,reset=>reset,s=>p(178)(27),cout=>p(179)(28));
FA_ff_3228:FAff port map(x=>p(75)(28),y=>p(76)(28),Cin=>p(77)(28),clock=>clock,reset=>reset,s=>p(178)(28),cout=>p(179)(29));
FA_ff_3229:FAff port map(x=>p(75)(29),y=>p(76)(29),Cin=>p(77)(29),clock=>clock,reset=>reset,s=>p(178)(29),cout=>p(179)(30));
FA_ff_3230:FAff port map(x=>p(75)(30),y=>p(76)(30),Cin=>p(77)(30),clock=>clock,reset=>reset,s=>p(178)(30),cout=>p(179)(31));
FA_ff_3231:FAff port map(x=>p(75)(31),y=>p(76)(31),Cin=>p(77)(31),clock=>clock,reset=>reset,s=>p(178)(31),cout=>p(179)(32));
FA_ff_3232:FAff port map(x=>p(75)(32),y=>p(76)(32),Cin=>p(77)(32),clock=>clock,reset=>reset,s=>p(178)(32),cout=>p(179)(33));
FA_ff_3233:FAff port map(x=>p(75)(33),y=>p(76)(33),Cin=>p(77)(33),clock=>clock,reset=>reset,s=>p(178)(33),cout=>p(179)(34));
FA_ff_3234:FAff port map(x=>p(75)(34),y=>p(76)(34),Cin=>p(77)(34),clock=>clock,reset=>reset,s=>p(178)(34),cout=>p(179)(35));
FA_ff_3235:FAff port map(x=>p(75)(35),y=>p(76)(35),Cin=>p(77)(35),clock=>clock,reset=>reset,s=>p(178)(35),cout=>p(179)(36));
FA_ff_3236:FAff port map(x=>p(75)(36),y=>p(76)(36),Cin=>p(77)(36),clock=>clock,reset=>reset,s=>p(178)(36),cout=>p(179)(37));
FA_ff_3237:FAff port map(x=>p(75)(37),y=>p(76)(37),Cin=>p(77)(37),clock=>clock,reset=>reset,s=>p(178)(37),cout=>p(179)(38));
FA_ff_3238:FAff port map(x=>p(75)(38),y=>p(76)(38),Cin=>p(77)(38),clock=>clock,reset=>reset,s=>p(178)(38),cout=>p(179)(39));
FA_ff_3239:FAff port map(x=>p(75)(39),y=>p(76)(39),Cin=>p(77)(39),clock=>clock,reset=>reset,s=>p(178)(39),cout=>p(179)(40));
FA_ff_3240:FAff port map(x=>p(75)(40),y=>p(76)(40),Cin=>p(77)(40),clock=>clock,reset=>reset,s=>p(178)(40),cout=>p(179)(41));
FA_ff_3241:FAff port map(x=>p(75)(41),y=>p(76)(41),Cin=>p(77)(41),clock=>clock,reset=>reset,s=>p(178)(41),cout=>p(179)(42));
FA_ff_3242:FAff port map(x=>p(75)(42),y=>p(76)(42),Cin=>p(77)(42),clock=>clock,reset=>reset,s=>p(178)(42),cout=>p(179)(43));
FA_ff_3243:FAff port map(x=>p(75)(43),y=>p(76)(43),Cin=>p(77)(43),clock=>clock,reset=>reset,s=>p(178)(43),cout=>p(179)(44));
FA_ff_3244:FAff port map(x=>p(75)(44),y=>p(76)(44),Cin=>p(77)(44),clock=>clock,reset=>reset,s=>p(178)(44),cout=>p(179)(45));
FA_ff_3245:FAff port map(x=>p(75)(45),y=>p(76)(45),Cin=>p(77)(45),clock=>clock,reset=>reset,s=>p(178)(45),cout=>p(179)(46));
FA_ff_3246:FAff port map(x=>p(75)(46),y=>p(76)(46),Cin=>p(77)(46),clock=>clock,reset=>reset,s=>p(178)(46),cout=>p(179)(47));
FA_ff_3247:FAff port map(x=>p(75)(47),y=>p(76)(47),Cin=>p(77)(47),clock=>clock,reset=>reset,s=>p(178)(47),cout=>p(179)(48));
FA_ff_3248:FAff port map(x=>p(75)(48),y=>p(76)(48),Cin=>p(77)(48),clock=>clock,reset=>reset,s=>p(178)(48),cout=>p(179)(49));
FA_ff_3249:FAff port map(x=>p(75)(49),y=>p(76)(49),Cin=>p(77)(49),clock=>clock,reset=>reset,s=>p(178)(49),cout=>p(179)(50));
FA_ff_3250:FAff port map(x=>p(75)(50),y=>p(76)(50),Cin=>p(77)(50),clock=>clock,reset=>reset,s=>p(178)(50),cout=>p(179)(51));
FA_ff_3251:FAff port map(x=>p(75)(51),y=>p(76)(51),Cin=>p(77)(51),clock=>clock,reset=>reset,s=>p(178)(51),cout=>p(179)(52));
FA_ff_3252:FAff port map(x=>p(75)(52),y=>p(76)(52),Cin=>p(77)(52),clock=>clock,reset=>reset,s=>p(178)(52),cout=>p(179)(53));
FA_ff_3253:FAff port map(x=>p(75)(53),y=>p(76)(53),Cin=>p(77)(53),clock=>clock,reset=>reset,s=>p(178)(53),cout=>p(179)(54));
FA_ff_3254:FAff port map(x=>p(75)(54),y=>p(76)(54),Cin=>p(77)(54),clock=>clock,reset=>reset,s=>p(178)(54),cout=>p(179)(55));
FA_ff_3255:FAff port map(x=>p(75)(55),y=>p(76)(55),Cin=>p(77)(55),clock=>clock,reset=>reset,s=>p(178)(55),cout=>p(179)(56));
FA_ff_3256:FAff port map(x=>p(75)(56),y=>p(76)(56),Cin=>p(77)(56),clock=>clock,reset=>reset,s=>p(178)(56),cout=>p(179)(57));
FA_ff_3257:FAff port map(x=>p(75)(57),y=>p(76)(57),Cin=>p(77)(57),clock=>clock,reset=>reset,s=>p(178)(57),cout=>p(179)(58));
FA_ff_3258:FAff port map(x=>p(75)(58),y=>p(76)(58),Cin=>p(77)(58),clock=>clock,reset=>reset,s=>p(178)(58),cout=>p(179)(59));
FA_ff_3259:FAff port map(x=>p(75)(59),y=>p(76)(59),Cin=>p(77)(59),clock=>clock,reset=>reset,s=>p(178)(59),cout=>p(179)(60));
FA_ff_3260:FAff port map(x=>p(75)(60),y=>p(76)(60),Cin=>p(77)(60),clock=>clock,reset=>reset,s=>p(178)(60),cout=>p(179)(61));
FA_ff_3261:FAff port map(x=>p(75)(61),y=>p(76)(61),Cin=>p(77)(61),clock=>clock,reset=>reset,s=>p(178)(61),cout=>p(179)(62));
FA_ff_3262:FAff port map(x=>p(75)(62),y=>p(76)(62),Cin=>p(77)(62),clock=>clock,reset=>reset,s=>p(178)(62),cout=>p(179)(63));
FA_ff_3263:FAff port map(x=>p(75)(63),y=>p(76)(63),Cin=>p(77)(63),clock=>clock,reset=>reset,s=>p(178)(63),cout=>p(179)(64));
FA_ff_3264:FAff port map(x=>p(75)(64),y=>p(76)(64),Cin=>p(77)(64),clock=>clock,reset=>reset,s=>p(178)(64),cout=>p(179)(65));
FA_ff_3265:FAff port map(x=>p(75)(65),y=>p(76)(65),Cin=>p(77)(65),clock=>clock,reset=>reset,s=>p(178)(65),cout=>p(179)(66));
FA_ff_3266:FAff port map(x=>p(75)(66),y=>p(76)(66),Cin=>p(77)(66),clock=>clock,reset=>reset,s=>p(178)(66),cout=>p(179)(67));
FA_ff_3267:FAff port map(x=>p(75)(67),y=>p(76)(67),Cin=>p(77)(67),clock=>clock,reset=>reset,s=>p(178)(67),cout=>p(179)(68));
FA_ff_3268:FAff port map(x=>p(75)(68),y=>p(76)(68),Cin=>p(77)(68),clock=>clock,reset=>reset,s=>p(178)(68),cout=>p(179)(69));
FA_ff_3269:FAff port map(x=>p(75)(69),y=>p(76)(69),Cin=>p(77)(69),clock=>clock,reset=>reset,s=>p(178)(69),cout=>p(179)(70));
FA_ff_3270:FAff port map(x=>p(75)(70),y=>p(76)(70),Cin=>p(77)(70),clock=>clock,reset=>reset,s=>p(178)(70),cout=>p(179)(71));
FA_ff_3271:FAff port map(x=>p(75)(71),y=>p(76)(71),Cin=>p(77)(71),clock=>clock,reset=>reset,s=>p(178)(71),cout=>p(179)(72));
FA_ff_3272:FAff port map(x=>p(75)(72),y=>p(76)(72),Cin=>p(77)(72),clock=>clock,reset=>reset,s=>p(178)(72),cout=>p(179)(73));
FA_ff_3273:FAff port map(x=>p(75)(73),y=>p(76)(73),Cin=>p(77)(73),clock=>clock,reset=>reset,s=>p(178)(73),cout=>p(179)(74));
FA_ff_3274:FAff port map(x=>p(75)(74),y=>p(76)(74),Cin=>p(77)(74),clock=>clock,reset=>reset,s=>p(178)(74),cout=>p(179)(75));
FA_ff_3275:FAff port map(x=>p(75)(75),y=>p(76)(75),Cin=>p(77)(75),clock=>clock,reset=>reset,s=>p(178)(75),cout=>p(179)(76));
FA_ff_3276:FAff port map(x=>p(75)(76),y=>p(76)(76),Cin=>p(77)(76),clock=>clock,reset=>reset,s=>p(178)(76),cout=>p(179)(77));
FA_ff_3277:FAff port map(x=>p(75)(77),y=>p(76)(77),Cin=>p(77)(77),clock=>clock,reset=>reset,s=>p(178)(77),cout=>p(179)(78));
FA_ff_3278:FAff port map(x=>p(75)(78),y=>p(76)(78),Cin=>p(77)(78),clock=>clock,reset=>reset,s=>p(178)(78),cout=>p(179)(79));
FA_ff_3279:FAff port map(x=>p(75)(79),y=>p(76)(79),Cin=>p(77)(79),clock=>clock,reset=>reset,s=>p(178)(79),cout=>p(179)(80));
FA_ff_3280:FAff port map(x=>p(75)(80),y=>p(76)(80),Cin=>p(77)(80),clock=>clock,reset=>reset,s=>p(178)(80),cout=>p(179)(81));
FA_ff_3281:FAff port map(x=>p(75)(81),y=>p(76)(81),Cin=>p(77)(81),clock=>clock,reset=>reset,s=>p(178)(81),cout=>p(179)(82));
FA_ff_3282:FAff port map(x=>p(75)(82),y=>p(76)(82),Cin=>p(77)(82),clock=>clock,reset=>reset,s=>p(178)(82),cout=>p(179)(83));
FA_ff_3283:FAff port map(x=>p(75)(83),y=>p(76)(83),Cin=>p(77)(83),clock=>clock,reset=>reset,s=>p(178)(83),cout=>p(179)(84));
FA_ff_3284:FAff port map(x=>p(75)(84),y=>p(76)(84),Cin=>p(77)(84),clock=>clock,reset=>reset,s=>p(178)(84),cout=>p(179)(85));
FA_ff_3285:FAff port map(x=>p(75)(85),y=>p(76)(85),Cin=>p(77)(85),clock=>clock,reset=>reset,s=>p(178)(85),cout=>p(179)(86));
FA_ff_3286:FAff port map(x=>p(75)(86),y=>p(76)(86),Cin=>p(77)(86),clock=>clock,reset=>reset,s=>p(178)(86),cout=>p(179)(87));
FA_ff_3287:FAff port map(x=>p(75)(87),y=>p(76)(87),Cin=>p(77)(87),clock=>clock,reset=>reset,s=>p(178)(87),cout=>p(179)(88));
FA_ff_3288:FAff port map(x=>p(75)(88),y=>p(76)(88),Cin=>p(77)(88),clock=>clock,reset=>reset,s=>p(178)(88),cout=>p(179)(89));
FA_ff_3289:FAff port map(x=>p(75)(89),y=>p(76)(89),Cin=>p(77)(89),clock=>clock,reset=>reset,s=>p(178)(89),cout=>p(179)(90));
FA_ff_3290:FAff port map(x=>p(75)(90),y=>p(76)(90),Cin=>p(77)(90),clock=>clock,reset=>reset,s=>p(178)(90),cout=>p(179)(91));
FA_ff_3291:FAff port map(x=>p(75)(91),y=>p(76)(91),Cin=>p(77)(91),clock=>clock,reset=>reset,s=>p(178)(91),cout=>p(179)(92));
FA_ff_3292:FAff port map(x=>p(75)(92),y=>p(76)(92),Cin=>p(77)(92),clock=>clock,reset=>reset,s=>p(178)(92),cout=>p(179)(93));
FA_ff_3293:FAff port map(x=>p(75)(93),y=>p(76)(93),Cin=>p(77)(93),clock=>clock,reset=>reset,s=>p(178)(93),cout=>p(179)(94));
FA_ff_3294:FAff port map(x=>p(75)(94),y=>p(76)(94),Cin=>p(77)(94),clock=>clock,reset=>reset,s=>p(178)(94),cout=>p(179)(95));
FA_ff_3295:FAff port map(x=>p(75)(95),y=>p(76)(95),Cin=>p(77)(95),clock=>clock,reset=>reset,s=>p(178)(95),cout=>p(179)(96));
FA_ff_3296:FAff port map(x=>p(75)(96),y=>p(76)(96),Cin=>p(77)(96),clock=>clock,reset=>reset,s=>p(178)(96),cout=>p(179)(97));
FA_ff_3297:FAff port map(x=>p(75)(97),y=>p(76)(97),Cin=>p(77)(97),clock=>clock,reset=>reset,s=>p(178)(97),cout=>p(179)(98));
FA_ff_3298:FAff port map(x=>p(75)(98),y=>p(76)(98),Cin=>p(77)(98),clock=>clock,reset=>reset,s=>p(178)(98),cout=>p(179)(99));
FA_ff_3299:FAff port map(x=>p(75)(99),y=>p(76)(99),Cin=>p(77)(99),clock=>clock,reset=>reset,s=>p(178)(99),cout=>p(179)(100));
FA_ff_3300:FAff port map(x=>p(75)(100),y=>p(76)(100),Cin=>p(77)(100),clock=>clock,reset=>reset,s=>p(178)(100),cout=>p(179)(101));
FA_ff_3301:FAff port map(x=>p(75)(101),y=>p(76)(101),Cin=>p(77)(101),clock=>clock,reset=>reset,s=>p(178)(101),cout=>p(179)(102));
FA_ff_3302:FAff port map(x=>p(75)(102),y=>p(76)(102),Cin=>p(77)(102),clock=>clock,reset=>reset,s=>p(178)(102),cout=>p(179)(103));
FA_ff_3303:FAff port map(x=>p(75)(103),y=>p(76)(103),Cin=>p(77)(103),clock=>clock,reset=>reset,s=>p(178)(103),cout=>p(179)(104));
FA_ff_3304:FAff port map(x=>p(75)(104),y=>p(76)(104),Cin=>p(77)(104),clock=>clock,reset=>reset,s=>p(178)(104),cout=>p(179)(105));
FA_ff_3305:FAff port map(x=>p(75)(105),y=>p(76)(105),Cin=>p(77)(105),clock=>clock,reset=>reset,s=>p(178)(105),cout=>p(179)(106));
FA_ff_3306:FAff port map(x=>p(75)(106),y=>p(76)(106),Cin=>p(77)(106),clock=>clock,reset=>reset,s=>p(178)(106),cout=>p(179)(107));
FA_ff_3307:FAff port map(x=>p(75)(107),y=>p(76)(107),Cin=>p(77)(107),clock=>clock,reset=>reset,s=>p(178)(107),cout=>p(179)(108));
FA_ff_3308:FAff port map(x=>p(75)(108),y=>p(76)(108),Cin=>p(77)(108),clock=>clock,reset=>reset,s=>p(178)(108),cout=>p(179)(109));
FA_ff_3309:FAff port map(x=>p(75)(109),y=>p(76)(109),Cin=>p(77)(109),clock=>clock,reset=>reset,s=>p(178)(109),cout=>p(179)(110));
FA_ff_3310:FAff port map(x=>p(75)(110),y=>p(76)(110),Cin=>p(77)(110),clock=>clock,reset=>reset,s=>p(178)(110),cout=>p(179)(111));
FA_ff_3311:FAff port map(x=>p(75)(111),y=>p(76)(111),Cin=>p(77)(111),clock=>clock,reset=>reset,s=>p(178)(111),cout=>p(179)(112));
FA_ff_3312:FAff port map(x=>p(75)(112),y=>p(76)(112),Cin=>p(77)(112),clock=>clock,reset=>reset,s=>p(178)(112),cout=>p(179)(113));
FA_ff_3313:FAff port map(x=>p(75)(113),y=>p(76)(113),Cin=>p(77)(113),clock=>clock,reset=>reset,s=>p(178)(113),cout=>p(179)(114));
FA_ff_3314:FAff port map(x=>p(75)(114),y=>p(76)(114),Cin=>p(77)(114),clock=>clock,reset=>reset,s=>p(178)(114),cout=>p(179)(115));
FA_ff_3315:FAff port map(x=>p(75)(115),y=>p(76)(115),Cin=>p(77)(115),clock=>clock,reset=>reset,s=>p(178)(115),cout=>p(179)(116));
FA_ff_3316:FAff port map(x=>p(75)(116),y=>p(76)(116),Cin=>p(77)(116),clock=>clock,reset=>reset,s=>p(178)(116),cout=>p(179)(117));
FA_ff_3317:FAff port map(x=>p(75)(117),y=>p(76)(117),Cin=>p(77)(117),clock=>clock,reset=>reset,s=>p(178)(117),cout=>p(179)(118));
FA_ff_3318:FAff port map(x=>p(75)(118),y=>p(76)(118),Cin=>p(77)(118),clock=>clock,reset=>reset,s=>p(178)(118),cout=>p(179)(119));
FA_ff_3319:FAff port map(x=>p(75)(119),y=>p(76)(119),Cin=>p(77)(119),clock=>clock,reset=>reset,s=>p(178)(119),cout=>p(179)(120));
FA_ff_3320:FAff port map(x=>p(75)(120),y=>p(76)(120),Cin=>p(77)(120),clock=>clock,reset=>reset,s=>p(178)(120),cout=>p(179)(121));
FA_ff_3321:FAff port map(x=>p(75)(121),y=>p(76)(121),Cin=>p(77)(121),clock=>clock,reset=>reset,s=>p(178)(121),cout=>p(179)(122));
FA_ff_3322:FAff port map(x=>p(75)(122),y=>p(76)(122),Cin=>p(77)(122),clock=>clock,reset=>reset,s=>p(178)(122),cout=>p(179)(123));
FA_ff_3323:FAff port map(x=>p(75)(123),y=>p(76)(123),Cin=>p(77)(123),clock=>clock,reset=>reset,s=>p(178)(123),cout=>p(179)(124));
FA_ff_3324:FAff port map(x=>p(75)(124),y=>p(76)(124),Cin=>p(77)(124),clock=>clock,reset=>reset,s=>p(178)(124),cout=>p(179)(125));
FA_ff_3325:FAff port map(x=>p(75)(125),y=>p(76)(125),Cin=>p(77)(125),clock=>clock,reset=>reset,s=>p(178)(125),cout=>p(179)(126));
FA_ff_3326:FAff port map(x=>p(75)(126),y=>p(76)(126),Cin=>p(77)(126),clock=>clock,reset=>reset,s=>p(178)(126),cout=>p(179)(127));
FA_ff_3327:FAff port map(x=>p(75)(127),y=>p(76)(127),Cin=>p(77)(127),clock=>clock,reset=>reset,s=>p(178)(127),cout=>p(179)(128));
FA_ff_3328:FAff port map(x=>p(78)(0),y=>p(79)(0),Cin=>p(80)(0),clock=>clock,reset=>reset,s=>p(180)(0),cout=>p(181)(1));
FA_ff_3329:FAff port map(x=>p(78)(1),y=>p(79)(1),Cin=>p(80)(1),clock=>clock,reset=>reset,s=>p(180)(1),cout=>p(181)(2));
FA_ff_3330:FAff port map(x=>p(78)(2),y=>p(79)(2),Cin=>p(80)(2),clock=>clock,reset=>reset,s=>p(180)(2),cout=>p(181)(3));
FA_ff_3331:FAff port map(x=>p(78)(3),y=>p(79)(3),Cin=>p(80)(3),clock=>clock,reset=>reset,s=>p(180)(3),cout=>p(181)(4));
FA_ff_3332:FAff port map(x=>p(78)(4),y=>p(79)(4),Cin=>p(80)(4),clock=>clock,reset=>reset,s=>p(180)(4),cout=>p(181)(5));
FA_ff_3333:FAff port map(x=>p(78)(5),y=>p(79)(5),Cin=>p(80)(5),clock=>clock,reset=>reset,s=>p(180)(5),cout=>p(181)(6));
FA_ff_3334:FAff port map(x=>p(78)(6),y=>p(79)(6),Cin=>p(80)(6),clock=>clock,reset=>reset,s=>p(180)(6),cout=>p(181)(7));
FA_ff_3335:FAff port map(x=>p(78)(7),y=>p(79)(7),Cin=>p(80)(7),clock=>clock,reset=>reset,s=>p(180)(7),cout=>p(181)(8));
FA_ff_3336:FAff port map(x=>p(78)(8),y=>p(79)(8),Cin=>p(80)(8),clock=>clock,reset=>reset,s=>p(180)(8),cout=>p(181)(9));
FA_ff_3337:FAff port map(x=>p(78)(9),y=>p(79)(9),Cin=>p(80)(9),clock=>clock,reset=>reset,s=>p(180)(9),cout=>p(181)(10));
FA_ff_3338:FAff port map(x=>p(78)(10),y=>p(79)(10),Cin=>p(80)(10),clock=>clock,reset=>reset,s=>p(180)(10),cout=>p(181)(11));
FA_ff_3339:FAff port map(x=>p(78)(11),y=>p(79)(11),Cin=>p(80)(11),clock=>clock,reset=>reset,s=>p(180)(11),cout=>p(181)(12));
FA_ff_3340:FAff port map(x=>p(78)(12),y=>p(79)(12),Cin=>p(80)(12),clock=>clock,reset=>reset,s=>p(180)(12),cout=>p(181)(13));
FA_ff_3341:FAff port map(x=>p(78)(13),y=>p(79)(13),Cin=>p(80)(13),clock=>clock,reset=>reset,s=>p(180)(13),cout=>p(181)(14));
FA_ff_3342:FAff port map(x=>p(78)(14),y=>p(79)(14),Cin=>p(80)(14),clock=>clock,reset=>reset,s=>p(180)(14),cout=>p(181)(15));
FA_ff_3343:FAff port map(x=>p(78)(15),y=>p(79)(15),Cin=>p(80)(15),clock=>clock,reset=>reset,s=>p(180)(15),cout=>p(181)(16));
FA_ff_3344:FAff port map(x=>p(78)(16),y=>p(79)(16),Cin=>p(80)(16),clock=>clock,reset=>reset,s=>p(180)(16),cout=>p(181)(17));
FA_ff_3345:FAff port map(x=>p(78)(17),y=>p(79)(17),Cin=>p(80)(17),clock=>clock,reset=>reset,s=>p(180)(17),cout=>p(181)(18));
FA_ff_3346:FAff port map(x=>p(78)(18),y=>p(79)(18),Cin=>p(80)(18),clock=>clock,reset=>reset,s=>p(180)(18),cout=>p(181)(19));
FA_ff_3347:FAff port map(x=>p(78)(19),y=>p(79)(19),Cin=>p(80)(19),clock=>clock,reset=>reset,s=>p(180)(19),cout=>p(181)(20));
FA_ff_3348:FAff port map(x=>p(78)(20),y=>p(79)(20),Cin=>p(80)(20),clock=>clock,reset=>reset,s=>p(180)(20),cout=>p(181)(21));
FA_ff_3349:FAff port map(x=>p(78)(21),y=>p(79)(21),Cin=>p(80)(21),clock=>clock,reset=>reset,s=>p(180)(21),cout=>p(181)(22));
FA_ff_3350:FAff port map(x=>p(78)(22),y=>p(79)(22),Cin=>p(80)(22),clock=>clock,reset=>reset,s=>p(180)(22),cout=>p(181)(23));
FA_ff_3351:FAff port map(x=>p(78)(23),y=>p(79)(23),Cin=>p(80)(23),clock=>clock,reset=>reset,s=>p(180)(23),cout=>p(181)(24));
FA_ff_3352:FAff port map(x=>p(78)(24),y=>p(79)(24),Cin=>p(80)(24),clock=>clock,reset=>reset,s=>p(180)(24),cout=>p(181)(25));
FA_ff_3353:FAff port map(x=>p(78)(25),y=>p(79)(25),Cin=>p(80)(25),clock=>clock,reset=>reset,s=>p(180)(25),cout=>p(181)(26));
FA_ff_3354:FAff port map(x=>p(78)(26),y=>p(79)(26),Cin=>p(80)(26),clock=>clock,reset=>reset,s=>p(180)(26),cout=>p(181)(27));
FA_ff_3355:FAff port map(x=>p(78)(27),y=>p(79)(27),Cin=>p(80)(27),clock=>clock,reset=>reset,s=>p(180)(27),cout=>p(181)(28));
FA_ff_3356:FAff port map(x=>p(78)(28),y=>p(79)(28),Cin=>p(80)(28),clock=>clock,reset=>reset,s=>p(180)(28),cout=>p(181)(29));
FA_ff_3357:FAff port map(x=>p(78)(29),y=>p(79)(29),Cin=>p(80)(29),clock=>clock,reset=>reset,s=>p(180)(29),cout=>p(181)(30));
FA_ff_3358:FAff port map(x=>p(78)(30),y=>p(79)(30),Cin=>p(80)(30),clock=>clock,reset=>reset,s=>p(180)(30),cout=>p(181)(31));
FA_ff_3359:FAff port map(x=>p(78)(31),y=>p(79)(31),Cin=>p(80)(31),clock=>clock,reset=>reset,s=>p(180)(31),cout=>p(181)(32));
FA_ff_3360:FAff port map(x=>p(78)(32),y=>p(79)(32),Cin=>p(80)(32),clock=>clock,reset=>reset,s=>p(180)(32),cout=>p(181)(33));
FA_ff_3361:FAff port map(x=>p(78)(33),y=>p(79)(33),Cin=>p(80)(33),clock=>clock,reset=>reset,s=>p(180)(33),cout=>p(181)(34));
FA_ff_3362:FAff port map(x=>p(78)(34),y=>p(79)(34),Cin=>p(80)(34),clock=>clock,reset=>reset,s=>p(180)(34),cout=>p(181)(35));
FA_ff_3363:FAff port map(x=>p(78)(35),y=>p(79)(35),Cin=>p(80)(35),clock=>clock,reset=>reset,s=>p(180)(35),cout=>p(181)(36));
FA_ff_3364:FAff port map(x=>p(78)(36),y=>p(79)(36),Cin=>p(80)(36),clock=>clock,reset=>reset,s=>p(180)(36),cout=>p(181)(37));
FA_ff_3365:FAff port map(x=>p(78)(37),y=>p(79)(37),Cin=>p(80)(37),clock=>clock,reset=>reset,s=>p(180)(37),cout=>p(181)(38));
FA_ff_3366:FAff port map(x=>p(78)(38),y=>p(79)(38),Cin=>p(80)(38),clock=>clock,reset=>reset,s=>p(180)(38),cout=>p(181)(39));
FA_ff_3367:FAff port map(x=>p(78)(39),y=>p(79)(39),Cin=>p(80)(39),clock=>clock,reset=>reset,s=>p(180)(39),cout=>p(181)(40));
FA_ff_3368:FAff port map(x=>p(78)(40),y=>p(79)(40),Cin=>p(80)(40),clock=>clock,reset=>reset,s=>p(180)(40),cout=>p(181)(41));
FA_ff_3369:FAff port map(x=>p(78)(41),y=>p(79)(41),Cin=>p(80)(41),clock=>clock,reset=>reset,s=>p(180)(41),cout=>p(181)(42));
FA_ff_3370:FAff port map(x=>p(78)(42),y=>p(79)(42),Cin=>p(80)(42),clock=>clock,reset=>reset,s=>p(180)(42),cout=>p(181)(43));
FA_ff_3371:FAff port map(x=>p(78)(43),y=>p(79)(43),Cin=>p(80)(43),clock=>clock,reset=>reset,s=>p(180)(43),cout=>p(181)(44));
FA_ff_3372:FAff port map(x=>p(78)(44),y=>p(79)(44),Cin=>p(80)(44),clock=>clock,reset=>reset,s=>p(180)(44),cout=>p(181)(45));
FA_ff_3373:FAff port map(x=>p(78)(45),y=>p(79)(45),Cin=>p(80)(45),clock=>clock,reset=>reset,s=>p(180)(45),cout=>p(181)(46));
FA_ff_3374:FAff port map(x=>p(78)(46),y=>p(79)(46),Cin=>p(80)(46),clock=>clock,reset=>reset,s=>p(180)(46),cout=>p(181)(47));
FA_ff_3375:FAff port map(x=>p(78)(47),y=>p(79)(47),Cin=>p(80)(47),clock=>clock,reset=>reset,s=>p(180)(47),cout=>p(181)(48));
FA_ff_3376:FAff port map(x=>p(78)(48),y=>p(79)(48),Cin=>p(80)(48),clock=>clock,reset=>reset,s=>p(180)(48),cout=>p(181)(49));
FA_ff_3377:FAff port map(x=>p(78)(49),y=>p(79)(49),Cin=>p(80)(49),clock=>clock,reset=>reset,s=>p(180)(49),cout=>p(181)(50));
FA_ff_3378:FAff port map(x=>p(78)(50),y=>p(79)(50),Cin=>p(80)(50),clock=>clock,reset=>reset,s=>p(180)(50),cout=>p(181)(51));
FA_ff_3379:FAff port map(x=>p(78)(51),y=>p(79)(51),Cin=>p(80)(51),clock=>clock,reset=>reset,s=>p(180)(51),cout=>p(181)(52));
FA_ff_3380:FAff port map(x=>p(78)(52),y=>p(79)(52),Cin=>p(80)(52),clock=>clock,reset=>reset,s=>p(180)(52),cout=>p(181)(53));
FA_ff_3381:FAff port map(x=>p(78)(53),y=>p(79)(53),Cin=>p(80)(53),clock=>clock,reset=>reset,s=>p(180)(53),cout=>p(181)(54));
FA_ff_3382:FAff port map(x=>p(78)(54),y=>p(79)(54),Cin=>p(80)(54),clock=>clock,reset=>reset,s=>p(180)(54),cout=>p(181)(55));
FA_ff_3383:FAff port map(x=>p(78)(55),y=>p(79)(55),Cin=>p(80)(55),clock=>clock,reset=>reset,s=>p(180)(55),cout=>p(181)(56));
FA_ff_3384:FAff port map(x=>p(78)(56),y=>p(79)(56),Cin=>p(80)(56),clock=>clock,reset=>reset,s=>p(180)(56),cout=>p(181)(57));
FA_ff_3385:FAff port map(x=>p(78)(57),y=>p(79)(57),Cin=>p(80)(57),clock=>clock,reset=>reset,s=>p(180)(57),cout=>p(181)(58));
FA_ff_3386:FAff port map(x=>p(78)(58),y=>p(79)(58),Cin=>p(80)(58),clock=>clock,reset=>reset,s=>p(180)(58),cout=>p(181)(59));
FA_ff_3387:FAff port map(x=>p(78)(59),y=>p(79)(59),Cin=>p(80)(59),clock=>clock,reset=>reset,s=>p(180)(59),cout=>p(181)(60));
FA_ff_3388:FAff port map(x=>p(78)(60),y=>p(79)(60),Cin=>p(80)(60),clock=>clock,reset=>reset,s=>p(180)(60),cout=>p(181)(61));
FA_ff_3389:FAff port map(x=>p(78)(61),y=>p(79)(61),Cin=>p(80)(61),clock=>clock,reset=>reset,s=>p(180)(61),cout=>p(181)(62));
FA_ff_3390:FAff port map(x=>p(78)(62),y=>p(79)(62),Cin=>p(80)(62),clock=>clock,reset=>reset,s=>p(180)(62),cout=>p(181)(63));
FA_ff_3391:FAff port map(x=>p(78)(63),y=>p(79)(63),Cin=>p(80)(63),clock=>clock,reset=>reset,s=>p(180)(63),cout=>p(181)(64));
FA_ff_3392:FAff port map(x=>p(78)(64),y=>p(79)(64),Cin=>p(80)(64),clock=>clock,reset=>reset,s=>p(180)(64),cout=>p(181)(65));
FA_ff_3393:FAff port map(x=>p(78)(65),y=>p(79)(65),Cin=>p(80)(65),clock=>clock,reset=>reset,s=>p(180)(65),cout=>p(181)(66));
FA_ff_3394:FAff port map(x=>p(78)(66),y=>p(79)(66),Cin=>p(80)(66),clock=>clock,reset=>reset,s=>p(180)(66),cout=>p(181)(67));
FA_ff_3395:FAff port map(x=>p(78)(67),y=>p(79)(67),Cin=>p(80)(67),clock=>clock,reset=>reset,s=>p(180)(67),cout=>p(181)(68));
FA_ff_3396:FAff port map(x=>p(78)(68),y=>p(79)(68),Cin=>p(80)(68),clock=>clock,reset=>reset,s=>p(180)(68),cout=>p(181)(69));
FA_ff_3397:FAff port map(x=>p(78)(69),y=>p(79)(69),Cin=>p(80)(69),clock=>clock,reset=>reset,s=>p(180)(69),cout=>p(181)(70));
FA_ff_3398:FAff port map(x=>p(78)(70),y=>p(79)(70),Cin=>p(80)(70),clock=>clock,reset=>reset,s=>p(180)(70),cout=>p(181)(71));
FA_ff_3399:FAff port map(x=>p(78)(71),y=>p(79)(71),Cin=>p(80)(71),clock=>clock,reset=>reset,s=>p(180)(71),cout=>p(181)(72));
FA_ff_3400:FAff port map(x=>p(78)(72),y=>p(79)(72),Cin=>p(80)(72),clock=>clock,reset=>reset,s=>p(180)(72),cout=>p(181)(73));
FA_ff_3401:FAff port map(x=>p(78)(73),y=>p(79)(73),Cin=>p(80)(73),clock=>clock,reset=>reset,s=>p(180)(73),cout=>p(181)(74));
FA_ff_3402:FAff port map(x=>p(78)(74),y=>p(79)(74),Cin=>p(80)(74),clock=>clock,reset=>reset,s=>p(180)(74),cout=>p(181)(75));
FA_ff_3403:FAff port map(x=>p(78)(75),y=>p(79)(75),Cin=>p(80)(75),clock=>clock,reset=>reset,s=>p(180)(75),cout=>p(181)(76));
FA_ff_3404:FAff port map(x=>p(78)(76),y=>p(79)(76),Cin=>p(80)(76),clock=>clock,reset=>reset,s=>p(180)(76),cout=>p(181)(77));
FA_ff_3405:FAff port map(x=>p(78)(77),y=>p(79)(77),Cin=>p(80)(77),clock=>clock,reset=>reset,s=>p(180)(77),cout=>p(181)(78));
FA_ff_3406:FAff port map(x=>p(78)(78),y=>p(79)(78),Cin=>p(80)(78),clock=>clock,reset=>reset,s=>p(180)(78),cout=>p(181)(79));
FA_ff_3407:FAff port map(x=>p(78)(79),y=>p(79)(79),Cin=>p(80)(79),clock=>clock,reset=>reset,s=>p(180)(79),cout=>p(181)(80));
FA_ff_3408:FAff port map(x=>p(78)(80),y=>p(79)(80),Cin=>p(80)(80),clock=>clock,reset=>reset,s=>p(180)(80),cout=>p(181)(81));
FA_ff_3409:FAff port map(x=>p(78)(81),y=>p(79)(81),Cin=>p(80)(81),clock=>clock,reset=>reset,s=>p(180)(81),cout=>p(181)(82));
FA_ff_3410:FAff port map(x=>p(78)(82),y=>p(79)(82),Cin=>p(80)(82),clock=>clock,reset=>reset,s=>p(180)(82),cout=>p(181)(83));
FA_ff_3411:FAff port map(x=>p(78)(83),y=>p(79)(83),Cin=>p(80)(83),clock=>clock,reset=>reset,s=>p(180)(83),cout=>p(181)(84));
FA_ff_3412:FAff port map(x=>p(78)(84),y=>p(79)(84),Cin=>p(80)(84),clock=>clock,reset=>reset,s=>p(180)(84),cout=>p(181)(85));
FA_ff_3413:FAff port map(x=>p(78)(85),y=>p(79)(85),Cin=>p(80)(85),clock=>clock,reset=>reset,s=>p(180)(85),cout=>p(181)(86));
FA_ff_3414:FAff port map(x=>p(78)(86),y=>p(79)(86),Cin=>p(80)(86),clock=>clock,reset=>reset,s=>p(180)(86),cout=>p(181)(87));
FA_ff_3415:FAff port map(x=>p(78)(87),y=>p(79)(87),Cin=>p(80)(87),clock=>clock,reset=>reset,s=>p(180)(87),cout=>p(181)(88));
FA_ff_3416:FAff port map(x=>p(78)(88),y=>p(79)(88),Cin=>p(80)(88),clock=>clock,reset=>reset,s=>p(180)(88),cout=>p(181)(89));
FA_ff_3417:FAff port map(x=>p(78)(89),y=>p(79)(89),Cin=>p(80)(89),clock=>clock,reset=>reset,s=>p(180)(89),cout=>p(181)(90));
FA_ff_3418:FAff port map(x=>p(78)(90),y=>p(79)(90),Cin=>p(80)(90),clock=>clock,reset=>reset,s=>p(180)(90),cout=>p(181)(91));
FA_ff_3419:FAff port map(x=>p(78)(91),y=>p(79)(91),Cin=>p(80)(91),clock=>clock,reset=>reset,s=>p(180)(91),cout=>p(181)(92));
FA_ff_3420:FAff port map(x=>p(78)(92),y=>p(79)(92),Cin=>p(80)(92),clock=>clock,reset=>reset,s=>p(180)(92),cout=>p(181)(93));
FA_ff_3421:FAff port map(x=>p(78)(93),y=>p(79)(93),Cin=>p(80)(93),clock=>clock,reset=>reset,s=>p(180)(93),cout=>p(181)(94));
FA_ff_3422:FAff port map(x=>p(78)(94),y=>p(79)(94),Cin=>p(80)(94),clock=>clock,reset=>reset,s=>p(180)(94),cout=>p(181)(95));
FA_ff_3423:FAff port map(x=>p(78)(95),y=>p(79)(95),Cin=>p(80)(95),clock=>clock,reset=>reset,s=>p(180)(95),cout=>p(181)(96));
FA_ff_3424:FAff port map(x=>p(78)(96),y=>p(79)(96),Cin=>p(80)(96),clock=>clock,reset=>reset,s=>p(180)(96),cout=>p(181)(97));
FA_ff_3425:FAff port map(x=>p(78)(97),y=>p(79)(97),Cin=>p(80)(97),clock=>clock,reset=>reset,s=>p(180)(97),cout=>p(181)(98));
FA_ff_3426:FAff port map(x=>p(78)(98),y=>p(79)(98),Cin=>p(80)(98),clock=>clock,reset=>reset,s=>p(180)(98),cout=>p(181)(99));
FA_ff_3427:FAff port map(x=>p(78)(99),y=>p(79)(99),Cin=>p(80)(99),clock=>clock,reset=>reset,s=>p(180)(99),cout=>p(181)(100));
FA_ff_3428:FAff port map(x=>p(78)(100),y=>p(79)(100),Cin=>p(80)(100),clock=>clock,reset=>reset,s=>p(180)(100),cout=>p(181)(101));
FA_ff_3429:FAff port map(x=>p(78)(101),y=>p(79)(101),Cin=>p(80)(101),clock=>clock,reset=>reset,s=>p(180)(101),cout=>p(181)(102));
FA_ff_3430:FAff port map(x=>p(78)(102),y=>p(79)(102),Cin=>p(80)(102),clock=>clock,reset=>reset,s=>p(180)(102),cout=>p(181)(103));
FA_ff_3431:FAff port map(x=>p(78)(103),y=>p(79)(103),Cin=>p(80)(103),clock=>clock,reset=>reset,s=>p(180)(103),cout=>p(181)(104));
FA_ff_3432:FAff port map(x=>p(78)(104),y=>p(79)(104),Cin=>p(80)(104),clock=>clock,reset=>reset,s=>p(180)(104),cout=>p(181)(105));
FA_ff_3433:FAff port map(x=>p(78)(105),y=>p(79)(105),Cin=>p(80)(105),clock=>clock,reset=>reset,s=>p(180)(105),cout=>p(181)(106));
FA_ff_3434:FAff port map(x=>p(78)(106),y=>p(79)(106),Cin=>p(80)(106),clock=>clock,reset=>reset,s=>p(180)(106),cout=>p(181)(107));
FA_ff_3435:FAff port map(x=>p(78)(107),y=>p(79)(107),Cin=>p(80)(107),clock=>clock,reset=>reset,s=>p(180)(107),cout=>p(181)(108));
FA_ff_3436:FAff port map(x=>p(78)(108),y=>p(79)(108),Cin=>p(80)(108),clock=>clock,reset=>reset,s=>p(180)(108),cout=>p(181)(109));
FA_ff_3437:FAff port map(x=>p(78)(109),y=>p(79)(109),Cin=>p(80)(109),clock=>clock,reset=>reset,s=>p(180)(109),cout=>p(181)(110));
FA_ff_3438:FAff port map(x=>p(78)(110),y=>p(79)(110),Cin=>p(80)(110),clock=>clock,reset=>reset,s=>p(180)(110),cout=>p(181)(111));
FA_ff_3439:FAff port map(x=>p(78)(111),y=>p(79)(111),Cin=>p(80)(111),clock=>clock,reset=>reset,s=>p(180)(111),cout=>p(181)(112));
FA_ff_3440:FAff port map(x=>p(78)(112),y=>p(79)(112),Cin=>p(80)(112),clock=>clock,reset=>reset,s=>p(180)(112),cout=>p(181)(113));
FA_ff_3441:FAff port map(x=>p(78)(113),y=>p(79)(113),Cin=>p(80)(113),clock=>clock,reset=>reset,s=>p(180)(113),cout=>p(181)(114));
FA_ff_3442:FAff port map(x=>p(78)(114),y=>p(79)(114),Cin=>p(80)(114),clock=>clock,reset=>reset,s=>p(180)(114),cout=>p(181)(115));
FA_ff_3443:FAff port map(x=>p(78)(115),y=>p(79)(115),Cin=>p(80)(115),clock=>clock,reset=>reset,s=>p(180)(115),cout=>p(181)(116));
FA_ff_3444:FAff port map(x=>p(78)(116),y=>p(79)(116),Cin=>p(80)(116),clock=>clock,reset=>reset,s=>p(180)(116),cout=>p(181)(117));
FA_ff_3445:FAff port map(x=>p(78)(117),y=>p(79)(117),Cin=>p(80)(117),clock=>clock,reset=>reset,s=>p(180)(117),cout=>p(181)(118));
FA_ff_3446:FAff port map(x=>p(78)(118),y=>p(79)(118),Cin=>p(80)(118),clock=>clock,reset=>reset,s=>p(180)(118),cout=>p(181)(119));
FA_ff_3447:FAff port map(x=>p(78)(119),y=>p(79)(119),Cin=>p(80)(119),clock=>clock,reset=>reset,s=>p(180)(119),cout=>p(181)(120));
FA_ff_3448:FAff port map(x=>p(78)(120),y=>p(79)(120),Cin=>p(80)(120),clock=>clock,reset=>reset,s=>p(180)(120),cout=>p(181)(121));
FA_ff_3449:FAff port map(x=>p(78)(121),y=>p(79)(121),Cin=>p(80)(121),clock=>clock,reset=>reset,s=>p(180)(121),cout=>p(181)(122));
FA_ff_3450:FAff port map(x=>p(78)(122),y=>p(79)(122),Cin=>p(80)(122),clock=>clock,reset=>reset,s=>p(180)(122),cout=>p(181)(123));
FA_ff_3451:FAff port map(x=>p(78)(123),y=>p(79)(123),Cin=>p(80)(123),clock=>clock,reset=>reset,s=>p(180)(123),cout=>p(181)(124));
FA_ff_3452:FAff port map(x=>p(78)(124),y=>p(79)(124),Cin=>p(80)(124),clock=>clock,reset=>reset,s=>p(180)(124),cout=>p(181)(125));
FA_ff_3453:FAff port map(x=>p(78)(125),y=>p(79)(125),Cin=>p(80)(125),clock=>clock,reset=>reset,s=>p(180)(125),cout=>p(181)(126));
FA_ff_3454:FAff port map(x=>p(78)(126),y=>p(79)(126),Cin=>p(80)(126),clock=>clock,reset=>reset,s=>p(180)(126),cout=>p(181)(127));
FA_ff_3455:FAff port map(x=>p(78)(127),y=>p(79)(127),Cin=>p(80)(127),clock=>clock,reset=>reset,s=>p(180)(127),cout=>p(181)(128));
FA_ff_3456:FAff port map(x=>p(81)(0),y=>p(82)(0),Cin=>p(83)(0),clock=>clock,reset=>reset,s=>p(182)(0),cout=>p(183)(1));
FA_ff_3457:FAff port map(x=>p(81)(1),y=>p(82)(1),Cin=>p(83)(1),clock=>clock,reset=>reset,s=>p(182)(1),cout=>p(183)(2));
FA_ff_3458:FAff port map(x=>p(81)(2),y=>p(82)(2),Cin=>p(83)(2),clock=>clock,reset=>reset,s=>p(182)(2),cout=>p(183)(3));
FA_ff_3459:FAff port map(x=>p(81)(3),y=>p(82)(3),Cin=>p(83)(3),clock=>clock,reset=>reset,s=>p(182)(3),cout=>p(183)(4));
FA_ff_3460:FAff port map(x=>p(81)(4),y=>p(82)(4),Cin=>p(83)(4),clock=>clock,reset=>reset,s=>p(182)(4),cout=>p(183)(5));
FA_ff_3461:FAff port map(x=>p(81)(5),y=>p(82)(5),Cin=>p(83)(5),clock=>clock,reset=>reset,s=>p(182)(5),cout=>p(183)(6));
FA_ff_3462:FAff port map(x=>p(81)(6),y=>p(82)(6),Cin=>p(83)(6),clock=>clock,reset=>reset,s=>p(182)(6),cout=>p(183)(7));
FA_ff_3463:FAff port map(x=>p(81)(7),y=>p(82)(7),Cin=>p(83)(7),clock=>clock,reset=>reset,s=>p(182)(7),cout=>p(183)(8));
FA_ff_3464:FAff port map(x=>p(81)(8),y=>p(82)(8),Cin=>p(83)(8),clock=>clock,reset=>reset,s=>p(182)(8),cout=>p(183)(9));
FA_ff_3465:FAff port map(x=>p(81)(9),y=>p(82)(9),Cin=>p(83)(9),clock=>clock,reset=>reset,s=>p(182)(9),cout=>p(183)(10));
FA_ff_3466:FAff port map(x=>p(81)(10),y=>p(82)(10),Cin=>p(83)(10),clock=>clock,reset=>reset,s=>p(182)(10),cout=>p(183)(11));
FA_ff_3467:FAff port map(x=>p(81)(11),y=>p(82)(11),Cin=>p(83)(11),clock=>clock,reset=>reset,s=>p(182)(11),cout=>p(183)(12));
FA_ff_3468:FAff port map(x=>p(81)(12),y=>p(82)(12),Cin=>p(83)(12),clock=>clock,reset=>reset,s=>p(182)(12),cout=>p(183)(13));
FA_ff_3469:FAff port map(x=>p(81)(13),y=>p(82)(13),Cin=>p(83)(13),clock=>clock,reset=>reset,s=>p(182)(13),cout=>p(183)(14));
FA_ff_3470:FAff port map(x=>p(81)(14),y=>p(82)(14),Cin=>p(83)(14),clock=>clock,reset=>reset,s=>p(182)(14),cout=>p(183)(15));
FA_ff_3471:FAff port map(x=>p(81)(15),y=>p(82)(15),Cin=>p(83)(15),clock=>clock,reset=>reset,s=>p(182)(15),cout=>p(183)(16));
FA_ff_3472:FAff port map(x=>p(81)(16),y=>p(82)(16),Cin=>p(83)(16),clock=>clock,reset=>reset,s=>p(182)(16),cout=>p(183)(17));
FA_ff_3473:FAff port map(x=>p(81)(17),y=>p(82)(17),Cin=>p(83)(17),clock=>clock,reset=>reset,s=>p(182)(17),cout=>p(183)(18));
FA_ff_3474:FAff port map(x=>p(81)(18),y=>p(82)(18),Cin=>p(83)(18),clock=>clock,reset=>reset,s=>p(182)(18),cout=>p(183)(19));
FA_ff_3475:FAff port map(x=>p(81)(19),y=>p(82)(19),Cin=>p(83)(19),clock=>clock,reset=>reset,s=>p(182)(19),cout=>p(183)(20));
FA_ff_3476:FAff port map(x=>p(81)(20),y=>p(82)(20),Cin=>p(83)(20),clock=>clock,reset=>reset,s=>p(182)(20),cout=>p(183)(21));
FA_ff_3477:FAff port map(x=>p(81)(21),y=>p(82)(21),Cin=>p(83)(21),clock=>clock,reset=>reset,s=>p(182)(21),cout=>p(183)(22));
FA_ff_3478:FAff port map(x=>p(81)(22),y=>p(82)(22),Cin=>p(83)(22),clock=>clock,reset=>reset,s=>p(182)(22),cout=>p(183)(23));
FA_ff_3479:FAff port map(x=>p(81)(23),y=>p(82)(23),Cin=>p(83)(23),clock=>clock,reset=>reset,s=>p(182)(23),cout=>p(183)(24));
FA_ff_3480:FAff port map(x=>p(81)(24),y=>p(82)(24),Cin=>p(83)(24),clock=>clock,reset=>reset,s=>p(182)(24),cout=>p(183)(25));
FA_ff_3481:FAff port map(x=>p(81)(25),y=>p(82)(25),Cin=>p(83)(25),clock=>clock,reset=>reset,s=>p(182)(25),cout=>p(183)(26));
FA_ff_3482:FAff port map(x=>p(81)(26),y=>p(82)(26),Cin=>p(83)(26),clock=>clock,reset=>reset,s=>p(182)(26),cout=>p(183)(27));
FA_ff_3483:FAff port map(x=>p(81)(27),y=>p(82)(27),Cin=>p(83)(27),clock=>clock,reset=>reset,s=>p(182)(27),cout=>p(183)(28));
FA_ff_3484:FAff port map(x=>p(81)(28),y=>p(82)(28),Cin=>p(83)(28),clock=>clock,reset=>reset,s=>p(182)(28),cout=>p(183)(29));
FA_ff_3485:FAff port map(x=>p(81)(29),y=>p(82)(29),Cin=>p(83)(29),clock=>clock,reset=>reset,s=>p(182)(29),cout=>p(183)(30));
FA_ff_3486:FAff port map(x=>p(81)(30),y=>p(82)(30),Cin=>p(83)(30),clock=>clock,reset=>reset,s=>p(182)(30),cout=>p(183)(31));
FA_ff_3487:FAff port map(x=>p(81)(31),y=>p(82)(31),Cin=>p(83)(31),clock=>clock,reset=>reset,s=>p(182)(31),cout=>p(183)(32));
FA_ff_3488:FAff port map(x=>p(81)(32),y=>p(82)(32),Cin=>p(83)(32),clock=>clock,reset=>reset,s=>p(182)(32),cout=>p(183)(33));
FA_ff_3489:FAff port map(x=>p(81)(33),y=>p(82)(33),Cin=>p(83)(33),clock=>clock,reset=>reset,s=>p(182)(33),cout=>p(183)(34));
FA_ff_3490:FAff port map(x=>p(81)(34),y=>p(82)(34),Cin=>p(83)(34),clock=>clock,reset=>reset,s=>p(182)(34),cout=>p(183)(35));
FA_ff_3491:FAff port map(x=>p(81)(35),y=>p(82)(35),Cin=>p(83)(35),clock=>clock,reset=>reset,s=>p(182)(35),cout=>p(183)(36));
FA_ff_3492:FAff port map(x=>p(81)(36),y=>p(82)(36),Cin=>p(83)(36),clock=>clock,reset=>reset,s=>p(182)(36),cout=>p(183)(37));
FA_ff_3493:FAff port map(x=>p(81)(37),y=>p(82)(37),Cin=>p(83)(37),clock=>clock,reset=>reset,s=>p(182)(37),cout=>p(183)(38));
FA_ff_3494:FAff port map(x=>p(81)(38),y=>p(82)(38),Cin=>p(83)(38),clock=>clock,reset=>reset,s=>p(182)(38),cout=>p(183)(39));
FA_ff_3495:FAff port map(x=>p(81)(39),y=>p(82)(39),Cin=>p(83)(39),clock=>clock,reset=>reset,s=>p(182)(39),cout=>p(183)(40));
FA_ff_3496:FAff port map(x=>p(81)(40),y=>p(82)(40),Cin=>p(83)(40),clock=>clock,reset=>reset,s=>p(182)(40),cout=>p(183)(41));
FA_ff_3497:FAff port map(x=>p(81)(41),y=>p(82)(41),Cin=>p(83)(41),clock=>clock,reset=>reset,s=>p(182)(41),cout=>p(183)(42));
FA_ff_3498:FAff port map(x=>p(81)(42),y=>p(82)(42),Cin=>p(83)(42),clock=>clock,reset=>reset,s=>p(182)(42),cout=>p(183)(43));
FA_ff_3499:FAff port map(x=>p(81)(43),y=>p(82)(43),Cin=>p(83)(43),clock=>clock,reset=>reset,s=>p(182)(43),cout=>p(183)(44));
FA_ff_3500:FAff port map(x=>p(81)(44),y=>p(82)(44),Cin=>p(83)(44),clock=>clock,reset=>reset,s=>p(182)(44),cout=>p(183)(45));
FA_ff_3501:FAff port map(x=>p(81)(45),y=>p(82)(45),Cin=>p(83)(45),clock=>clock,reset=>reset,s=>p(182)(45),cout=>p(183)(46));
FA_ff_3502:FAff port map(x=>p(81)(46),y=>p(82)(46),Cin=>p(83)(46),clock=>clock,reset=>reset,s=>p(182)(46),cout=>p(183)(47));
FA_ff_3503:FAff port map(x=>p(81)(47),y=>p(82)(47),Cin=>p(83)(47),clock=>clock,reset=>reset,s=>p(182)(47),cout=>p(183)(48));
FA_ff_3504:FAff port map(x=>p(81)(48),y=>p(82)(48),Cin=>p(83)(48),clock=>clock,reset=>reset,s=>p(182)(48),cout=>p(183)(49));
FA_ff_3505:FAff port map(x=>p(81)(49),y=>p(82)(49),Cin=>p(83)(49),clock=>clock,reset=>reset,s=>p(182)(49),cout=>p(183)(50));
FA_ff_3506:FAff port map(x=>p(81)(50),y=>p(82)(50),Cin=>p(83)(50),clock=>clock,reset=>reset,s=>p(182)(50),cout=>p(183)(51));
FA_ff_3507:FAff port map(x=>p(81)(51),y=>p(82)(51),Cin=>p(83)(51),clock=>clock,reset=>reset,s=>p(182)(51),cout=>p(183)(52));
FA_ff_3508:FAff port map(x=>p(81)(52),y=>p(82)(52),Cin=>p(83)(52),clock=>clock,reset=>reset,s=>p(182)(52),cout=>p(183)(53));
FA_ff_3509:FAff port map(x=>p(81)(53),y=>p(82)(53),Cin=>p(83)(53),clock=>clock,reset=>reset,s=>p(182)(53),cout=>p(183)(54));
FA_ff_3510:FAff port map(x=>p(81)(54),y=>p(82)(54),Cin=>p(83)(54),clock=>clock,reset=>reset,s=>p(182)(54),cout=>p(183)(55));
FA_ff_3511:FAff port map(x=>p(81)(55),y=>p(82)(55),Cin=>p(83)(55),clock=>clock,reset=>reset,s=>p(182)(55),cout=>p(183)(56));
FA_ff_3512:FAff port map(x=>p(81)(56),y=>p(82)(56),Cin=>p(83)(56),clock=>clock,reset=>reset,s=>p(182)(56),cout=>p(183)(57));
FA_ff_3513:FAff port map(x=>p(81)(57),y=>p(82)(57),Cin=>p(83)(57),clock=>clock,reset=>reset,s=>p(182)(57),cout=>p(183)(58));
FA_ff_3514:FAff port map(x=>p(81)(58),y=>p(82)(58),Cin=>p(83)(58),clock=>clock,reset=>reset,s=>p(182)(58),cout=>p(183)(59));
FA_ff_3515:FAff port map(x=>p(81)(59),y=>p(82)(59),Cin=>p(83)(59),clock=>clock,reset=>reset,s=>p(182)(59),cout=>p(183)(60));
FA_ff_3516:FAff port map(x=>p(81)(60),y=>p(82)(60),Cin=>p(83)(60),clock=>clock,reset=>reset,s=>p(182)(60),cout=>p(183)(61));
FA_ff_3517:FAff port map(x=>p(81)(61),y=>p(82)(61),Cin=>p(83)(61),clock=>clock,reset=>reset,s=>p(182)(61),cout=>p(183)(62));
FA_ff_3518:FAff port map(x=>p(81)(62),y=>p(82)(62),Cin=>p(83)(62),clock=>clock,reset=>reset,s=>p(182)(62),cout=>p(183)(63));
FA_ff_3519:FAff port map(x=>p(81)(63),y=>p(82)(63),Cin=>p(83)(63),clock=>clock,reset=>reset,s=>p(182)(63),cout=>p(183)(64));
FA_ff_3520:FAff port map(x=>p(81)(64),y=>p(82)(64),Cin=>p(83)(64),clock=>clock,reset=>reset,s=>p(182)(64),cout=>p(183)(65));
FA_ff_3521:FAff port map(x=>p(81)(65),y=>p(82)(65),Cin=>p(83)(65),clock=>clock,reset=>reset,s=>p(182)(65),cout=>p(183)(66));
FA_ff_3522:FAff port map(x=>p(81)(66),y=>p(82)(66),Cin=>p(83)(66),clock=>clock,reset=>reset,s=>p(182)(66),cout=>p(183)(67));
FA_ff_3523:FAff port map(x=>p(81)(67),y=>p(82)(67),Cin=>p(83)(67),clock=>clock,reset=>reset,s=>p(182)(67),cout=>p(183)(68));
FA_ff_3524:FAff port map(x=>p(81)(68),y=>p(82)(68),Cin=>p(83)(68),clock=>clock,reset=>reset,s=>p(182)(68),cout=>p(183)(69));
FA_ff_3525:FAff port map(x=>p(81)(69),y=>p(82)(69),Cin=>p(83)(69),clock=>clock,reset=>reset,s=>p(182)(69),cout=>p(183)(70));
FA_ff_3526:FAff port map(x=>p(81)(70),y=>p(82)(70),Cin=>p(83)(70),clock=>clock,reset=>reset,s=>p(182)(70),cout=>p(183)(71));
FA_ff_3527:FAff port map(x=>p(81)(71),y=>p(82)(71),Cin=>p(83)(71),clock=>clock,reset=>reset,s=>p(182)(71),cout=>p(183)(72));
FA_ff_3528:FAff port map(x=>p(81)(72),y=>p(82)(72),Cin=>p(83)(72),clock=>clock,reset=>reset,s=>p(182)(72),cout=>p(183)(73));
FA_ff_3529:FAff port map(x=>p(81)(73),y=>p(82)(73),Cin=>p(83)(73),clock=>clock,reset=>reset,s=>p(182)(73),cout=>p(183)(74));
FA_ff_3530:FAff port map(x=>p(81)(74),y=>p(82)(74),Cin=>p(83)(74),clock=>clock,reset=>reset,s=>p(182)(74),cout=>p(183)(75));
FA_ff_3531:FAff port map(x=>p(81)(75),y=>p(82)(75),Cin=>p(83)(75),clock=>clock,reset=>reset,s=>p(182)(75),cout=>p(183)(76));
FA_ff_3532:FAff port map(x=>p(81)(76),y=>p(82)(76),Cin=>p(83)(76),clock=>clock,reset=>reset,s=>p(182)(76),cout=>p(183)(77));
FA_ff_3533:FAff port map(x=>p(81)(77),y=>p(82)(77),Cin=>p(83)(77),clock=>clock,reset=>reset,s=>p(182)(77),cout=>p(183)(78));
FA_ff_3534:FAff port map(x=>p(81)(78),y=>p(82)(78),Cin=>p(83)(78),clock=>clock,reset=>reset,s=>p(182)(78),cout=>p(183)(79));
FA_ff_3535:FAff port map(x=>p(81)(79),y=>p(82)(79),Cin=>p(83)(79),clock=>clock,reset=>reset,s=>p(182)(79),cout=>p(183)(80));
FA_ff_3536:FAff port map(x=>p(81)(80),y=>p(82)(80),Cin=>p(83)(80),clock=>clock,reset=>reset,s=>p(182)(80),cout=>p(183)(81));
FA_ff_3537:FAff port map(x=>p(81)(81),y=>p(82)(81),Cin=>p(83)(81),clock=>clock,reset=>reset,s=>p(182)(81),cout=>p(183)(82));
FA_ff_3538:FAff port map(x=>p(81)(82),y=>p(82)(82),Cin=>p(83)(82),clock=>clock,reset=>reset,s=>p(182)(82),cout=>p(183)(83));
FA_ff_3539:FAff port map(x=>p(81)(83),y=>p(82)(83),Cin=>p(83)(83),clock=>clock,reset=>reset,s=>p(182)(83),cout=>p(183)(84));
FA_ff_3540:FAff port map(x=>p(81)(84),y=>p(82)(84),Cin=>p(83)(84),clock=>clock,reset=>reset,s=>p(182)(84),cout=>p(183)(85));
FA_ff_3541:FAff port map(x=>p(81)(85),y=>p(82)(85),Cin=>p(83)(85),clock=>clock,reset=>reset,s=>p(182)(85),cout=>p(183)(86));
FA_ff_3542:FAff port map(x=>p(81)(86),y=>p(82)(86),Cin=>p(83)(86),clock=>clock,reset=>reset,s=>p(182)(86),cout=>p(183)(87));
FA_ff_3543:FAff port map(x=>p(81)(87),y=>p(82)(87),Cin=>p(83)(87),clock=>clock,reset=>reset,s=>p(182)(87),cout=>p(183)(88));
FA_ff_3544:FAff port map(x=>p(81)(88),y=>p(82)(88),Cin=>p(83)(88),clock=>clock,reset=>reset,s=>p(182)(88),cout=>p(183)(89));
FA_ff_3545:FAff port map(x=>p(81)(89),y=>p(82)(89),Cin=>p(83)(89),clock=>clock,reset=>reset,s=>p(182)(89),cout=>p(183)(90));
FA_ff_3546:FAff port map(x=>p(81)(90),y=>p(82)(90),Cin=>p(83)(90),clock=>clock,reset=>reset,s=>p(182)(90),cout=>p(183)(91));
FA_ff_3547:FAff port map(x=>p(81)(91),y=>p(82)(91),Cin=>p(83)(91),clock=>clock,reset=>reset,s=>p(182)(91),cout=>p(183)(92));
FA_ff_3548:FAff port map(x=>p(81)(92),y=>p(82)(92),Cin=>p(83)(92),clock=>clock,reset=>reset,s=>p(182)(92),cout=>p(183)(93));
FA_ff_3549:FAff port map(x=>p(81)(93),y=>p(82)(93),Cin=>p(83)(93),clock=>clock,reset=>reset,s=>p(182)(93),cout=>p(183)(94));
FA_ff_3550:FAff port map(x=>p(81)(94),y=>p(82)(94),Cin=>p(83)(94),clock=>clock,reset=>reset,s=>p(182)(94),cout=>p(183)(95));
FA_ff_3551:FAff port map(x=>p(81)(95),y=>p(82)(95),Cin=>p(83)(95),clock=>clock,reset=>reset,s=>p(182)(95),cout=>p(183)(96));
FA_ff_3552:FAff port map(x=>p(81)(96),y=>p(82)(96),Cin=>p(83)(96),clock=>clock,reset=>reset,s=>p(182)(96),cout=>p(183)(97));
FA_ff_3553:FAff port map(x=>p(81)(97),y=>p(82)(97),Cin=>p(83)(97),clock=>clock,reset=>reset,s=>p(182)(97),cout=>p(183)(98));
FA_ff_3554:FAff port map(x=>p(81)(98),y=>p(82)(98),Cin=>p(83)(98),clock=>clock,reset=>reset,s=>p(182)(98),cout=>p(183)(99));
FA_ff_3555:FAff port map(x=>p(81)(99),y=>p(82)(99),Cin=>p(83)(99),clock=>clock,reset=>reset,s=>p(182)(99),cout=>p(183)(100));
FA_ff_3556:FAff port map(x=>p(81)(100),y=>p(82)(100),Cin=>p(83)(100),clock=>clock,reset=>reset,s=>p(182)(100),cout=>p(183)(101));
FA_ff_3557:FAff port map(x=>p(81)(101),y=>p(82)(101),Cin=>p(83)(101),clock=>clock,reset=>reset,s=>p(182)(101),cout=>p(183)(102));
FA_ff_3558:FAff port map(x=>p(81)(102),y=>p(82)(102),Cin=>p(83)(102),clock=>clock,reset=>reset,s=>p(182)(102),cout=>p(183)(103));
FA_ff_3559:FAff port map(x=>p(81)(103),y=>p(82)(103),Cin=>p(83)(103),clock=>clock,reset=>reset,s=>p(182)(103),cout=>p(183)(104));
FA_ff_3560:FAff port map(x=>p(81)(104),y=>p(82)(104),Cin=>p(83)(104),clock=>clock,reset=>reset,s=>p(182)(104),cout=>p(183)(105));
FA_ff_3561:FAff port map(x=>p(81)(105),y=>p(82)(105),Cin=>p(83)(105),clock=>clock,reset=>reset,s=>p(182)(105),cout=>p(183)(106));
FA_ff_3562:FAff port map(x=>p(81)(106),y=>p(82)(106),Cin=>p(83)(106),clock=>clock,reset=>reset,s=>p(182)(106),cout=>p(183)(107));
FA_ff_3563:FAff port map(x=>p(81)(107),y=>p(82)(107),Cin=>p(83)(107),clock=>clock,reset=>reset,s=>p(182)(107),cout=>p(183)(108));
FA_ff_3564:FAff port map(x=>p(81)(108),y=>p(82)(108),Cin=>p(83)(108),clock=>clock,reset=>reset,s=>p(182)(108),cout=>p(183)(109));
FA_ff_3565:FAff port map(x=>p(81)(109),y=>p(82)(109),Cin=>p(83)(109),clock=>clock,reset=>reset,s=>p(182)(109),cout=>p(183)(110));
FA_ff_3566:FAff port map(x=>p(81)(110),y=>p(82)(110),Cin=>p(83)(110),clock=>clock,reset=>reset,s=>p(182)(110),cout=>p(183)(111));
FA_ff_3567:FAff port map(x=>p(81)(111),y=>p(82)(111),Cin=>p(83)(111),clock=>clock,reset=>reset,s=>p(182)(111),cout=>p(183)(112));
FA_ff_3568:FAff port map(x=>p(81)(112),y=>p(82)(112),Cin=>p(83)(112),clock=>clock,reset=>reset,s=>p(182)(112),cout=>p(183)(113));
FA_ff_3569:FAff port map(x=>p(81)(113),y=>p(82)(113),Cin=>p(83)(113),clock=>clock,reset=>reset,s=>p(182)(113),cout=>p(183)(114));
FA_ff_3570:FAff port map(x=>p(81)(114),y=>p(82)(114),Cin=>p(83)(114),clock=>clock,reset=>reset,s=>p(182)(114),cout=>p(183)(115));
FA_ff_3571:FAff port map(x=>p(81)(115),y=>p(82)(115),Cin=>p(83)(115),clock=>clock,reset=>reset,s=>p(182)(115),cout=>p(183)(116));
FA_ff_3572:FAff port map(x=>p(81)(116),y=>p(82)(116),Cin=>p(83)(116),clock=>clock,reset=>reset,s=>p(182)(116),cout=>p(183)(117));
FA_ff_3573:FAff port map(x=>p(81)(117),y=>p(82)(117),Cin=>p(83)(117),clock=>clock,reset=>reset,s=>p(182)(117),cout=>p(183)(118));
FA_ff_3574:FAff port map(x=>p(81)(118),y=>p(82)(118),Cin=>p(83)(118),clock=>clock,reset=>reset,s=>p(182)(118),cout=>p(183)(119));
FA_ff_3575:FAff port map(x=>p(81)(119),y=>p(82)(119),Cin=>p(83)(119),clock=>clock,reset=>reset,s=>p(182)(119),cout=>p(183)(120));
FA_ff_3576:FAff port map(x=>p(81)(120),y=>p(82)(120),Cin=>p(83)(120),clock=>clock,reset=>reset,s=>p(182)(120),cout=>p(183)(121));
FA_ff_3577:FAff port map(x=>p(81)(121),y=>p(82)(121),Cin=>p(83)(121),clock=>clock,reset=>reset,s=>p(182)(121),cout=>p(183)(122));
FA_ff_3578:FAff port map(x=>p(81)(122),y=>p(82)(122),Cin=>p(83)(122),clock=>clock,reset=>reset,s=>p(182)(122),cout=>p(183)(123));
FA_ff_3579:FAff port map(x=>p(81)(123),y=>p(82)(123),Cin=>p(83)(123),clock=>clock,reset=>reset,s=>p(182)(123),cout=>p(183)(124));
FA_ff_3580:FAff port map(x=>p(81)(124),y=>p(82)(124),Cin=>p(83)(124),clock=>clock,reset=>reset,s=>p(182)(124),cout=>p(183)(125));
FA_ff_3581:FAff port map(x=>p(81)(125),y=>p(82)(125),Cin=>p(83)(125),clock=>clock,reset=>reset,s=>p(182)(125),cout=>p(183)(126));
FA_ff_3582:FAff port map(x=>p(81)(126),y=>p(82)(126),Cin=>p(83)(126),clock=>clock,reset=>reset,s=>p(182)(126),cout=>p(183)(127));
FA_ff_3583:FAff port map(x=>p(81)(127),y=>p(82)(127),Cin=>p(83)(127),clock=>clock,reset=>reset,s=>p(182)(127),cout=>p(183)(128));
FA_ff_3584:FAff port map(x=>p(84)(0),y=>p(85)(0),Cin=>p(86)(0),clock=>clock,reset=>reset,s=>p(184)(0),cout=>p(185)(1));
FA_ff_3585:FAff port map(x=>p(84)(1),y=>p(85)(1),Cin=>p(86)(1),clock=>clock,reset=>reset,s=>p(184)(1),cout=>p(185)(2));
FA_ff_3586:FAff port map(x=>p(84)(2),y=>p(85)(2),Cin=>p(86)(2),clock=>clock,reset=>reset,s=>p(184)(2),cout=>p(185)(3));
FA_ff_3587:FAff port map(x=>p(84)(3),y=>p(85)(3),Cin=>p(86)(3),clock=>clock,reset=>reset,s=>p(184)(3),cout=>p(185)(4));
FA_ff_3588:FAff port map(x=>p(84)(4),y=>p(85)(4),Cin=>p(86)(4),clock=>clock,reset=>reset,s=>p(184)(4),cout=>p(185)(5));
FA_ff_3589:FAff port map(x=>p(84)(5),y=>p(85)(5),Cin=>p(86)(5),clock=>clock,reset=>reset,s=>p(184)(5),cout=>p(185)(6));
FA_ff_3590:FAff port map(x=>p(84)(6),y=>p(85)(6),Cin=>p(86)(6),clock=>clock,reset=>reset,s=>p(184)(6),cout=>p(185)(7));
FA_ff_3591:FAff port map(x=>p(84)(7),y=>p(85)(7),Cin=>p(86)(7),clock=>clock,reset=>reset,s=>p(184)(7),cout=>p(185)(8));
FA_ff_3592:FAff port map(x=>p(84)(8),y=>p(85)(8),Cin=>p(86)(8),clock=>clock,reset=>reset,s=>p(184)(8),cout=>p(185)(9));
FA_ff_3593:FAff port map(x=>p(84)(9),y=>p(85)(9),Cin=>p(86)(9),clock=>clock,reset=>reset,s=>p(184)(9),cout=>p(185)(10));
FA_ff_3594:FAff port map(x=>p(84)(10),y=>p(85)(10),Cin=>p(86)(10),clock=>clock,reset=>reset,s=>p(184)(10),cout=>p(185)(11));
FA_ff_3595:FAff port map(x=>p(84)(11),y=>p(85)(11),Cin=>p(86)(11),clock=>clock,reset=>reset,s=>p(184)(11),cout=>p(185)(12));
FA_ff_3596:FAff port map(x=>p(84)(12),y=>p(85)(12),Cin=>p(86)(12),clock=>clock,reset=>reset,s=>p(184)(12),cout=>p(185)(13));
FA_ff_3597:FAff port map(x=>p(84)(13),y=>p(85)(13),Cin=>p(86)(13),clock=>clock,reset=>reset,s=>p(184)(13),cout=>p(185)(14));
FA_ff_3598:FAff port map(x=>p(84)(14),y=>p(85)(14),Cin=>p(86)(14),clock=>clock,reset=>reset,s=>p(184)(14),cout=>p(185)(15));
FA_ff_3599:FAff port map(x=>p(84)(15),y=>p(85)(15),Cin=>p(86)(15),clock=>clock,reset=>reset,s=>p(184)(15),cout=>p(185)(16));
FA_ff_3600:FAff port map(x=>p(84)(16),y=>p(85)(16),Cin=>p(86)(16),clock=>clock,reset=>reset,s=>p(184)(16),cout=>p(185)(17));
FA_ff_3601:FAff port map(x=>p(84)(17),y=>p(85)(17),Cin=>p(86)(17),clock=>clock,reset=>reset,s=>p(184)(17),cout=>p(185)(18));
FA_ff_3602:FAff port map(x=>p(84)(18),y=>p(85)(18),Cin=>p(86)(18),clock=>clock,reset=>reset,s=>p(184)(18),cout=>p(185)(19));
FA_ff_3603:FAff port map(x=>p(84)(19),y=>p(85)(19),Cin=>p(86)(19),clock=>clock,reset=>reset,s=>p(184)(19),cout=>p(185)(20));
FA_ff_3604:FAff port map(x=>p(84)(20),y=>p(85)(20),Cin=>p(86)(20),clock=>clock,reset=>reset,s=>p(184)(20),cout=>p(185)(21));
FA_ff_3605:FAff port map(x=>p(84)(21),y=>p(85)(21),Cin=>p(86)(21),clock=>clock,reset=>reset,s=>p(184)(21),cout=>p(185)(22));
FA_ff_3606:FAff port map(x=>p(84)(22),y=>p(85)(22),Cin=>p(86)(22),clock=>clock,reset=>reset,s=>p(184)(22),cout=>p(185)(23));
FA_ff_3607:FAff port map(x=>p(84)(23),y=>p(85)(23),Cin=>p(86)(23),clock=>clock,reset=>reset,s=>p(184)(23),cout=>p(185)(24));
FA_ff_3608:FAff port map(x=>p(84)(24),y=>p(85)(24),Cin=>p(86)(24),clock=>clock,reset=>reset,s=>p(184)(24),cout=>p(185)(25));
FA_ff_3609:FAff port map(x=>p(84)(25),y=>p(85)(25),Cin=>p(86)(25),clock=>clock,reset=>reset,s=>p(184)(25),cout=>p(185)(26));
FA_ff_3610:FAff port map(x=>p(84)(26),y=>p(85)(26),Cin=>p(86)(26),clock=>clock,reset=>reset,s=>p(184)(26),cout=>p(185)(27));
FA_ff_3611:FAff port map(x=>p(84)(27),y=>p(85)(27),Cin=>p(86)(27),clock=>clock,reset=>reset,s=>p(184)(27),cout=>p(185)(28));
FA_ff_3612:FAff port map(x=>p(84)(28),y=>p(85)(28),Cin=>p(86)(28),clock=>clock,reset=>reset,s=>p(184)(28),cout=>p(185)(29));
FA_ff_3613:FAff port map(x=>p(84)(29),y=>p(85)(29),Cin=>p(86)(29),clock=>clock,reset=>reset,s=>p(184)(29),cout=>p(185)(30));
FA_ff_3614:FAff port map(x=>p(84)(30),y=>p(85)(30),Cin=>p(86)(30),clock=>clock,reset=>reset,s=>p(184)(30),cout=>p(185)(31));
FA_ff_3615:FAff port map(x=>p(84)(31),y=>p(85)(31),Cin=>p(86)(31),clock=>clock,reset=>reset,s=>p(184)(31),cout=>p(185)(32));
FA_ff_3616:FAff port map(x=>p(84)(32),y=>p(85)(32),Cin=>p(86)(32),clock=>clock,reset=>reset,s=>p(184)(32),cout=>p(185)(33));
FA_ff_3617:FAff port map(x=>p(84)(33),y=>p(85)(33),Cin=>p(86)(33),clock=>clock,reset=>reset,s=>p(184)(33),cout=>p(185)(34));
FA_ff_3618:FAff port map(x=>p(84)(34),y=>p(85)(34),Cin=>p(86)(34),clock=>clock,reset=>reset,s=>p(184)(34),cout=>p(185)(35));
FA_ff_3619:FAff port map(x=>p(84)(35),y=>p(85)(35),Cin=>p(86)(35),clock=>clock,reset=>reset,s=>p(184)(35),cout=>p(185)(36));
FA_ff_3620:FAff port map(x=>p(84)(36),y=>p(85)(36),Cin=>p(86)(36),clock=>clock,reset=>reset,s=>p(184)(36),cout=>p(185)(37));
FA_ff_3621:FAff port map(x=>p(84)(37),y=>p(85)(37),Cin=>p(86)(37),clock=>clock,reset=>reset,s=>p(184)(37),cout=>p(185)(38));
FA_ff_3622:FAff port map(x=>p(84)(38),y=>p(85)(38),Cin=>p(86)(38),clock=>clock,reset=>reset,s=>p(184)(38),cout=>p(185)(39));
FA_ff_3623:FAff port map(x=>p(84)(39),y=>p(85)(39),Cin=>p(86)(39),clock=>clock,reset=>reset,s=>p(184)(39),cout=>p(185)(40));
FA_ff_3624:FAff port map(x=>p(84)(40),y=>p(85)(40),Cin=>p(86)(40),clock=>clock,reset=>reset,s=>p(184)(40),cout=>p(185)(41));
FA_ff_3625:FAff port map(x=>p(84)(41),y=>p(85)(41),Cin=>p(86)(41),clock=>clock,reset=>reset,s=>p(184)(41),cout=>p(185)(42));
FA_ff_3626:FAff port map(x=>p(84)(42),y=>p(85)(42),Cin=>p(86)(42),clock=>clock,reset=>reset,s=>p(184)(42),cout=>p(185)(43));
FA_ff_3627:FAff port map(x=>p(84)(43),y=>p(85)(43),Cin=>p(86)(43),clock=>clock,reset=>reset,s=>p(184)(43),cout=>p(185)(44));
FA_ff_3628:FAff port map(x=>p(84)(44),y=>p(85)(44),Cin=>p(86)(44),clock=>clock,reset=>reset,s=>p(184)(44),cout=>p(185)(45));
FA_ff_3629:FAff port map(x=>p(84)(45),y=>p(85)(45),Cin=>p(86)(45),clock=>clock,reset=>reset,s=>p(184)(45),cout=>p(185)(46));
FA_ff_3630:FAff port map(x=>p(84)(46),y=>p(85)(46),Cin=>p(86)(46),clock=>clock,reset=>reset,s=>p(184)(46),cout=>p(185)(47));
FA_ff_3631:FAff port map(x=>p(84)(47),y=>p(85)(47),Cin=>p(86)(47),clock=>clock,reset=>reset,s=>p(184)(47),cout=>p(185)(48));
FA_ff_3632:FAff port map(x=>p(84)(48),y=>p(85)(48),Cin=>p(86)(48),clock=>clock,reset=>reset,s=>p(184)(48),cout=>p(185)(49));
FA_ff_3633:FAff port map(x=>p(84)(49),y=>p(85)(49),Cin=>p(86)(49),clock=>clock,reset=>reset,s=>p(184)(49),cout=>p(185)(50));
FA_ff_3634:FAff port map(x=>p(84)(50),y=>p(85)(50),Cin=>p(86)(50),clock=>clock,reset=>reset,s=>p(184)(50),cout=>p(185)(51));
FA_ff_3635:FAff port map(x=>p(84)(51),y=>p(85)(51),Cin=>p(86)(51),clock=>clock,reset=>reset,s=>p(184)(51),cout=>p(185)(52));
FA_ff_3636:FAff port map(x=>p(84)(52),y=>p(85)(52),Cin=>p(86)(52),clock=>clock,reset=>reset,s=>p(184)(52),cout=>p(185)(53));
FA_ff_3637:FAff port map(x=>p(84)(53),y=>p(85)(53),Cin=>p(86)(53),clock=>clock,reset=>reset,s=>p(184)(53),cout=>p(185)(54));
FA_ff_3638:FAff port map(x=>p(84)(54),y=>p(85)(54),Cin=>p(86)(54),clock=>clock,reset=>reset,s=>p(184)(54),cout=>p(185)(55));
FA_ff_3639:FAff port map(x=>p(84)(55),y=>p(85)(55),Cin=>p(86)(55),clock=>clock,reset=>reset,s=>p(184)(55),cout=>p(185)(56));
FA_ff_3640:FAff port map(x=>p(84)(56),y=>p(85)(56),Cin=>p(86)(56),clock=>clock,reset=>reset,s=>p(184)(56),cout=>p(185)(57));
FA_ff_3641:FAff port map(x=>p(84)(57),y=>p(85)(57),Cin=>p(86)(57),clock=>clock,reset=>reset,s=>p(184)(57),cout=>p(185)(58));
FA_ff_3642:FAff port map(x=>p(84)(58),y=>p(85)(58),Cin=>p(86)(58),clock=>clock,reset=>reset,s=>p(184)(58),cout=>p(185)(59));
FA_ff_3643:FAff port map(x=>p(84)(59),y=>p(85)(59),Cin=>p(86)(59),clock=>clock,reset=>reset,s=>p(184)(59),cout=>p(185)(60));
FA_ff_3644:FAff port map(x=>p(84)(60),y=>p(85)(60),Cin=>p(86)(60),clock=>clock,reset=>reset,s=>p(184)(60),cout=>p(185)(61));
FA_ff_3645:FAff port map(x=>p(84)(61),y=>p(85)(61),Cin=>p(86)(61),clock=>clock,reset=>reset,s=>p(184)(61),cout=>p(185)(62));
FA_ff_3646:FAff port map(x=>p(84)(62),y=>p(85)(62),Cin=>p(86)(62),clock=>clock,reset=>reset,s=>p(184)(62),cout=>p(185)(63));
FA_ff_3647:FAff port map(x=>p(84)(63),y=>p(85)(63),Cin=>p(86)(63),clock=>clock,reset=>reset,s=>p(184)(63),cout=>p(185)(64));
FA_ff_3648:FAff port map(x=>p(84)(64),y=>p(85)(64),Cin=>p(86)(64),clock=>clock,reset=>reset,s=>p(184)(64),cout=>p(185)(65));
FA_ff_3649:FAff port map(x=>p(84)(65),y=>p(85)(65),Cin=>p(86)(65),clock=>clock,reset=>reset,s=>p(184)(65),cout=>p(185)(66));
FA_ff_3650:FAff port map(x=>p(84)(66),y=>p(85)(66),Cin=>p(86)(66),clock=>clock,reset=>reset,s=>p(184)(66),cout=>p(185)(67));
FA_ff_3651:FAff port map(x=>p(84)(67),y=>p(85)(67),Cin=>p(86)(67),clock=>clock,reset=>reset,s=>p(184)(67),cout=>p(185)(68));
FA_ff_3652:FAff port map(x=>p(84)(68),y=>p(85)(68),Cin=>p(86)(68),clock=>clock,reset=>reset,s=>p(184)(68),cout=>p(185)(69));
FA_ff_3653:FAff port map(x=>p(84)(69),y=>p(85)(69),Cin=>p(86)(69),clock=>clock,reset=>reset,s=>p(184)(69),cout=>p(185)(70));
FA_ff_3654:FAff port map(x=>p(84)(70),y=>p(85)(70),Cin=>p(86)(70),clock=>clock,reset=>reset,s=>p(184)(70),cout=>p(185)(71));
FA_ff_3655:FAff port map(x=>p(84)(71),y=>p(85)(71),Cin=>p(86)(71),clock=>clock,reset=>reset,s=>p(184)(71),cout=>p(185)(72));
FA_ff_3656:FAff port map(x=>p(84)(72),y=>p(85)(72),Cin=>p(86)(72),clock=>clock,reset=>reset,s=>p(184)(72),cout=>p(185)(73));
FA_ff_3657:FAff port map(x=>p(84)(73),y=>p(85)(73),Cin=>p(86)(73),clock=>clock,reset=>reset,s=>p(184)(73),cout=>p(185)(74));
FA_ff_3658:FAff port map(x=>p(84)(74),y=>p(85)(74),Cin=>p(86)(74),clock=>clock,reset=>reset,s=>p(184)(74),cout=>p(185)(75));
FA_ff_3659:FAff port map(x=>p(84)(75),y=>p(85)(75),Cin=>p(86)(75),clock=>clock,reset=>reset,s=>p(184)(75),cout=>p(185)(76));
FA_ff_3660:FAff port map(x=>p(84)(76),y=>p(85)(76),Cin=>p(86)(76),clock=>clock,reset=>reset,s=>p(184)(76),cout=>p(185)(77));
FA_ff_3661:FAff port map(x=>p(84)(77),y=>p(85)(77),Cin=>p(86)(77),clock=>clock,reset=>reset,s=>p(184)(77),cout=>p(185)(78));
FA_ff_3662:FAff port map(x=>p(84)(78),y=>p(85)(78),Cin=>p(86)(78),clock=>clock,reset=>reset,s=>p(184)(78),cout=>p(185)(79));
FA_ff_3663:FAff port map(x=>p(84)(79),y=>p(85)(79),Cin=>p(86)(79),clock=>clock,reset=>reset,s=>p(184)(79),cout=>p(185)(80));
FA_ff_3664:FAff port map(x=>p(84)(80),y=>p(85)(80),Cin=>p(86)(80),clock=>clock,reset=>reset,s=>p(184)(80),cout=>p(185)(81));
FA_ff_3665:FAff port map(x=>p(84)(81),y=>p(85)(81),Cin=>p(86)(81),clock=>clock,reset=>reset,s=>p(184)(81),cout=>p(185)(82));
FA_ff_3666:FAff port map(x=>p(84)(82),y=>p(85)(82),Cin=>p(86)(82),clock=>clock,reset=>reset,s=>p(184)(82),cout=>p(185)(83));
FA_ff_3667:FAff port map(x=>p(84)(83),y=>p(85)(83),Cin=>p(86)(83),clock=>clock,reset=>reset,s=>p(184)(83),cout=>p(185)(84));
FA_ff_3668:FAff port map(x=>p(84)(84),y=>p(85)(84),Cin=>p(86)(84),clock=>clock,reset=>reset,s=>p(184)(84),cout=>p(185)(85));
FA_ff_3669:FAff port map(x=>p(84)(85),y=>p(85)(85),Cin=>p(86)(85),clock=>clock,reset=>reset,s=>p(184)(85),cout=>p(185)(86));
FA_ff_3670:FAff port map(x=>p(84)(86),y=>p(85)(86),Cin=>p(86)(86),clock=>clock,reset=>reset,s=>p(184)(86),cout=>p(185)(87));
FA_ff_3671:FAff port map(x=>p(84)(87),y=>p(85)(87),Cin=>p(86)(87),clock=>clock,reset=>reset,s=>p(184)(87),cout=>p(185)(88));
FA_ff_3672:FAff port map(x=>p(84)(88),y=>p(85)(88),Cin=>p(86)(88),clock=>clock,reset=>reset,s=>p(184)(88),cout=>p(185)(89));
FA_ff_3673:FAff port map(x=>p(84)(89),y=>p(85)(89),Cin=>p(86)(89),clock=>clock,reset=>reset,s=>p(184)(89),cout=>p(185)(90));
FA_ff_3674:FAff port map(x=>p(84)(90),y=>p(85)(90),Cin=>p(86)(90),clock=>clock,reset=>reset,s=>p(184)(90),cout=>p(185)(91));
FA_ff_3675:FAff port map(x=>p(84)(91),y=>p(85)(91),Cin=>p(86)(91),clock=>clock,reset=>reset,s=>p(184)(91),cout=>p(185)(92));
FA_ff_3676:FAff port map(x=>p(84)(92),y=>p(85)(92),Cin=>p(86)(92),clock=>clock,reset=>reset,s=>p(184)(92),cout=>p(185)(93));
FA_ff_3677:FAff port map(x=>p(84)(93),y=>p(85)(93),Cin=>p(86)(93),clock=>clock,reset=>reset,s=>p(184)(93),cout=>p(185)(94));
FA_ff_3678:FAff port map(x=>p(84)(94),y=>p(85)(94),Cin=>p(86)(94),clock=>clock,reset=>reset,s=>p(184)(94),cout=>p(185)(95));
FA_ff_3679:FAff port map(x=>p(84)(95),y=>p(85)(95),Cin=>p(86)(95),clock=>clock,reset=>reset,s=>p(184)(95),cout=>p(185)(96));
FA_ff_3680:FAff port map(x=>p(84)(96),y=>p(85)(96),Cin=>p(86)(96),clock=>clock,reset=>reset,s=>p(184)(96),cout=>p(185)(97));
FA_ff_3681:FAff port map(x=>p(84)(97),y=>p(85)(97),Cin=>p(86)(97),clock=>clock,reset=>reset,s=>p(184)(97),cout=>p(185)(98));
FA_ff_3682:FAff port map(x=>p(84)(98),y=>p(85)(98),Cin=>p(86)(98),clock=>clock,reset=>reset,s=>p(184)(98),cout=>p(185)(99));
FA_ff_3683:FAff port map(x=>p(84)(99),y=>p(85)(99),Cin=>p(86)(99),clock=>clock,reset=>reset,s=>p(184)(99),cout=>p(185)(100));
FA_ff_3684:FAff port map(x=>p(84)(100),y=>p(85)(100),Cin=>p(86)(100),clock=>clock,reset=>reset,s=>p(184)(100),cout=>p(185)(101));
FA_ff_3685:FAff port map(x=>p(84)(101),y=>p(85)(101),Cin=>p(86)(101),clock=>clock,reset=>reset,s=>p(184)(101),cout=>p(185)(102));
FA_ff_3686:FAff port map(x=>p(84)(102),y=>p(85)(102),Cin=>p(86)(102),clock=>clock,reset=>reset,s=>p(184)(102),cout=>p(185)(103));
FA_ff_3687:FAff port map(x=>p(84)(103),y=>p(85)(103),Cin=>p(86)(103),clock=>clock,reset=>reset,s=>p(184)(103),cout=>p(185)(104));
FA_ff_3688:FAff port map(x=>p(84)(104),y=>p(85)(104),Cin=>p(86)(104),clock=>clock,reset=>reset,s=>p(184)(104),cout=>p(185)(105));
FA_ff_3689:FAff port map(x=>p(84)(105),y=>p(85)(105),Cin=>p(86)(105),clock=>clock,reset=>reset,s=>p(184)(105),cout=>p(185)(106));
FA_ff_3690:FAff port map(x=>p(84)(106),y=>p(85)(106),Cin=>p(86)(106),clock=>clock,reset=>reset,s=>p(184)(106),cout=>p(185)(107));
FA_ff_3691:FAff port map(x=>p(84)(107),y=>p(85)(107),Cin=>p(86)(107),clock=>clock,reset=>reset,s=>p(184)(107),cout=>p(185)(108));
FA_ff_3692:FAff port map(x=>p(84)(108),y=>p(85)(108),Cin=>p(86)(108),clock=>clock,reset=>reset,s=>p(184)(108),cout=>p(185)(109));
FA_ff_3693:FAff port map(x=>p(84)(109),y=>p(85)(109),Cin=>p(86)(109),clock=>clock,reset=>reset,s=>p(184)(109),cout=>p(185)(110));
FA_ff_3694:FAff port map(x=>p(84)(110),y=>p(85)(110),Cin=>p(86)(110),clock=>clock,reset=>reset,s=>p(184)(110),cout=>p(185)(111));
FA_ff_3695:FAff port map(x=>p(84)(111),y=>p(85)(111),Cin=>p(86)(111),clock=>clock,reset=>reset,s=>p(184)(111),cout=>p(185)(112));
FA_ff_3696:FAff port map(x=>p(84)(112),y=>p(85)(112),Cin=>p(86)(112),clock=>clock,reset=>reset,s=>p(184)(112),cout=>p(185)(113));
FA_ff_3697:FAff port map(x=>p(84)(113),y=>p(85)(113),Cin=>p(86)(113),clock=>clock,reset=>reset,s=>p(184)(113),cout=>p(185)(114));
FA_ff_3698:FAff port map(x=>p(84)(114),y=>p(85)(114),Cin=>p(86)(114),clock=>clock,reset=>reset,s=>p(184)(114),cout=>p(185)(115));
FA_ff_3699:FAff port map(x=>p(84)(115),y=>p(85)(115),Cin=>p(86)(115),clock=>clock,reset=>reset,s=>p(184)(115),cout=>p(185)(116));
FA_ff_3700:FAff port map(x=>p(84)(116),y=>p(85)(116),Cin=>p(86)(116),clock=>clock,reset=>reset,s=>p(184)(116),cout=>p(185)(117));
FA_ff_3701:FAff port map(x=>p(84)(117),y=>p(85)(117),Cin=>p(86)(117),clock=>clock,reset=>reset,s=>p(184)(117),cout=>p(185)(118));
FA_ff_3702:FAff port map(x=>p(84)(118),y=>p(85)(118),Cin=>p(86)(118),clock=>clock,reset=>reset,s=>p(184)(118),cout=>p(185)(119));
FA_ff_3703:FAff port map(x=>p(84)(119),y=>p(85)(119),Cin=>p(86)(119),clock=>clock,reset=>reset,s=>p(184)(119),cout=>p(185)(120));
FA_ff_3704:FAff port map(x=>p(84)(120),y=>p(85)(120),Cin=>p(86)(120),clock=>clock,reset=>reset,s=>p(184)(120),cout=>p(185)(121));
FA_ff_3705:FAff port map(x=>p(84)(121),y=>p(85)(121),Cin=>p(86)(121),clock=>clock,reset=>reset,s=>p(184)(121),cout=>p(185)(122));
FA_ff_3706:FAff port map(x=>p(84)(122),y=>p(85)(122),Cin=>p(86)(122),clock=>clock,reset=>reset,s=>p(184)(122),cout=>p(185)(123));
FA_ff_3707:FAff port map(x=>p(84)(123),y=>p(85)(123),Cin=>p(86)(123),clock=>clock,reset=>reset,s=>p(184)(123),cout=>p(185)(124));
FA_ff_3708:FAff port map(x=>p(84)(124),y=>p(85)(124),Cin=>p(86)(124),clock=>clock,reset=>reset,s=>p(184)(124),cout=>p(185)(125));
FA_ff_3709:FAff port map(x=>p(84)(125),y=>p(85)(125),Cin=>p(86)(125),clock=>clock,reset=>reset,s=>p(184)(125),cout=>p(185)(126));
FA_ff_3710:FAff port map(x=>p(84)(126),y=>p(85)(126),Cin=>p(86)(126),clock=>clock,reset=>reset,s=>p(184)(126),cout=>p(185)(127));
FA_ff_3711:FAff port map(x=>p(84)(127),y=>p(85)(127),Cin=>p(86)(127),clock=>clock,reset=>reset,s=>p(184)(127),cout=>p(185)(128));
FA_ff_3712:FAff port map(x=>p(87)(0),y=>p(88)(0),Cin=>p(89)(0),clock=>clock,reset=>reset,s=>p(186)(0),cout=>p(187)(1));
FA_ff_3713:FAff port map(x=>p(87)(1),y=>p(88)(1),Cin=>p(89)(1),clock=>clock,reset=>reset,s=>p(186)(1),cout=>p(187)(2));
FA_ff_3714:FAff port map(x=>p(87)(2),y=>p(88)(2),Cin=>p(89)(2),clock=>clock,reset=>reset,s=>p(186)(2),cout=>p(187)(3));
FA_ff_3715:FAff port map(x=>p(87)(3),y=>p(88)(3),Cin=>p(89)(3),clock=>clock,reset=>reset,s=>p(186)(3),cout=>p(187)(4));
FA_ff_3716:FAff port map(x=>p(87)(4),y=>p(88)(4),Cin=>p(89)(4),clock=>clock,reset=>reset,s=>p(186)(4),cout=>p(187)(5));
FA_ff_3717:FAff port map(x=>p(87)(5),y=>p(88)(5),Cin=>p(89)(5),clock=>clock,reset=>reset,s=>p(186)(5),cout=>p(187)(6));
FA_ff_3718:FAff port map(x=>p(87)(6),y=>p(88)(6),Cin=>p(89)(6),clock=>clock,reset=>reset,s=>p(186)(6),cout=>p(187)(7));
FA_ff_3719:FAff port map(x=>p(87)(7),y=>p(88)(7),Cin=>p(89)(7),clock=>clock,reset=>reset,s=>p(186)(7),cout=>p(187)(8));
FA_ff_3720:FAff port map(x=>p(87)(8),y=>p(88)(8),Cin=>p(89)(8),clock=>clock,reset=>reset,s=>p(186)(8),cout=>p(187)(9));
FA_ff_3721:FAff port map(x=>p(87)(9),y=>p(88)(9),Cin=>p(89)(9),clock=>clock,reset=>reset,s=>p(186)(9),cout=>p(187)(10));
FA_ff_3722:FAff port map(x=>p(87)(10),y=>p(88)(10),Cin=>p(89)(10),clock=>clock,reset=>reset,s=>p(186)(10),cout=>p(187)(11));
FA_ff_3723:FAff port map(x=>p(87)(11),y=>p(88)(11),Cin=>p(89)(11),clock=>clock,reset=>reset,s=>p(186)(11),cout=>p(187)(12));
FA_ff_3724:FAff port map(x=>p(87)(12),y=>p(88)(12),Cin=>p(89)(12),clock=>clock,reset=>reset,s=>p(186)(12),cout=>p(187)(13));
FA_ff_3725:FAff port map(x=>p(87)(13),y=>p(88)(13),Cin=>p(89)(13),clock=>clock,reset=>reset,s=>p(186)(13),cout=>p(187)(14));
FA_ff_3726:FAff port map(x=>p(87)(14),y=>p(88)(14),Cin=>p(89)(14),clock=>clock,reset=>reset,s=>p(186)(14),cout=>p(187)(15));
FA_ff_3727:FAff port map(x=>p(87)(15),y=>p(88)(15),Cin=>p(89)(15),clock=>clock,reset=>reset,s=>p(186)(15),cout=>p(187)(16));
FA_ff_3728:FAff port map(x=>p(87)(16),y=>p(88)(16),Cin=>p(89)(16),clock=>clock,reset=>reset,s=>p(186)(16),cout=>p(187)(17));
FA_ff_3729:FAff port map(x=>p(87)(17),y=>p(88)(17),Cin=>p(89)(17),clock=>clock,reset=>reset,s=>p(186)(17),cout=>p(187)(18));
FA_ff_3730:FAff port map(x=>p(87)(18),y=>p(88)(18),Cin=>p(89)(18),clock=>clock,reset=>reset,s=>p(186)(18),cout=>p(187)(19));
FA_ff_3731:FAff port map(x=>p(87)(19),y=>p(88)(19),Cin=>p(89)(19),clock=>clock,reset=>reset,s=>p(186)(19),cout=>p(187)(20));
FA_ff_3732:FAff port map(x=>p(87)(20),y=>p(88)(20),Cin=>p(89)(20),clock=>clock,reset=>reset,s=>p(186)(20),cout=>p(187)(21));
FA_ff_3733:FAff port map(x=>p(87)(21),y=>p(88)(21),Cin=>p(89)(21),clock=>clock,reset=>reset,s=>p(186)(21),cout=>p(187)(22));
FA_ff_3734:FAff port map(x=>p(87)(22),y=>p(88)(22),Cin=>p(89)(22),clock=>clock,reset=>reset,s=>p(186)(22),cout=>p(187)(23));
FA_ff_3735:FAff port map(x=>p(87)(23),y=>p(88)(23),Cin=>p(89)(23),clock=>clock,reset=>reset,s=>p(186)(23),cout=>p(187)(24));
FA_ff_3736:FAff port map(x=>p(87)(24),y=>p(88)(24),Cin=>p(89)(24),clock=>clock,reset=>reset,s=>p(186)(24),cout=>p(187)(25));
FA_ff_3737:FAff port map(x=>p(87)(25),y=>p(88)(25),Cin=>p(89)(25),clock=>clock,reset=>reset,s=>p(186)(25),cout=>p(187)(26));
FA_ff_3738:FAff port map(x=>p(87)(26),y=>p(88)(26),Cin=>p(89)(26),clock=>clock,reset=>reset,s=>p(186)(26),cout=>p(187)(27));
FA_ff_3739:FAff port map(x=>p(87)(27),y=>p(88)(27),Cin=>p(89)(27),clock=>clock,reset=>reset,s=>p(186)(27),cout=>p(187)(28));
FA_ff_3740:FAff port map(x=>p(87)(28),y=>p(88)(28),Cin=>p(89)(28),clock=>clock,reset=>reset,s=>p(186)(28),cout=>p(187)(29));
FA_ff_3741:FAff port map(x=>p(87)(29),y=>p(88)(29),Cin=>p(89)(29),clock=>clock,reset=>reset,s=>p(186)(29),cout=>p(187)(30));
FA_ff_3742:FAff port map(x=>p(87)(30),y=>p(88)(30),Cin=>p(89)(30),clock=>clock,reset=>reset,s=>p(186)(30),cout=>p(187)(31));
FA_ff_3743:FAff port map(x=>p(87)(31),y=>p(88)(31),Cin=>p(89)(31),clock=>clock,reset=>reset,s=>p(186)(31),cout=>p(187)(32));
FA_ff_3744:FAff port map(x=>p(87)(32),y=>p(88)(32),Cin=>p(89)(32),clock=>clock,reset=>reset,s=>p(186)(32),cout=>p(187)(33));
FA_ff_3745:FAff port map(x=>p(87)(33),y=>p(88)(33),Cin=>p(89)(33),clock=>clock,reset=>reset,s=>p(186)(33),cout=>p(187)(34));
FA_ff_3746:FAff port map(x=>p(87)(34),y=>p(88)(34),Cin=>p(89)(34),clock=>clock,reset=>reset,s=>p(186)(34),cout=>p(187)(35));
FA_ff_3747:FAff port map(x=>p(87)(35),y=>p(88)(35),Cin=>p(89)(35),clock=>clock,reset=>reset,s=>p(186)(35),cout=>p(187)(36));
FA_ff_3748:FAff port map(x=>p(87)(36),y=>p(88)(36),Cin=>p(89)(36),clock=>clock,reset=>reset,s=>p(186)(36),cout=>p(187)(37));
FA_ff_3749:FAff port map(x=>p(87)(37),y=>p(88)(37),Cin=>p(89)(37),clock=>clock,reset=>reset,s=>p(186)(37),cout=>p(187)(38));
FA_ff_3750:FAff port map(x=>p(87)(38),y=>p(88)(38),Cin=>p(89)(38),clock=>clock,reset=>reset,s=>p(186)(38),cout=>p(187)(39));
FA_ff_3751:FAff port map(x=>p(87)(39),y=>p(88)(39),Cin=>p(89)(39),clock=>clock,reset=>reset,s=>p(186)(39),cout=>p(187)(40));
FA_ff_3752:FAff port map(x=>p(87)(40),y=>p(88)(40),Cin=>p(89)(40),clock=>clock,reset=>reset,s=>p(186)(40),cout=>p(187)(41));
FA_ff_3753:FAff port map(x=>p(87)(41),y=>p(88)(41),Cin=>p(89)(41),clock=>clock,reset=>reset,s=>p(186)(41),cout=>p(187)(42));
FA_ff_3754:FAff port map(x=>p(87)(42),y=>p(88)(42),Cin=>p(89)(42),clock=>clock,reset=>reset,s=>p(186)(42),cout=>p(187)(43));
FA_ff_3755:FAff port map(x=>p(87)(43),y=>p(88)(43),Cin=>p(89)(43),clock=>clock,reset=>reset,s=>p(186)(43),cout=>p(187)(44));
FA_ff_3756:FAff port map(x=>p(87)(44),y=>p(88)(44),Cin=>p(89)(44),clock=>clock,reset=>reset,s=>p(186)(44),cout=>p(187)(45));
FA_ff_3757:FAff port map(x=>p(87)(45),y=>p(88)(45),Cin=>p(89)(45),clock=>clock,reset=>reset,s=>p(186)(45),cout=>p(187)(46));
FA_ff_3758:FAff port map(x=>p(87)(46),y=>p(88)(46),Cin=>p(89)(46),clock=>clock,reset=>reset,s=>p(186)(46),cout=>p(187)(47));
FA_ff_3759:FAff port map(x=>p(87)(47),y=>p(88)(47),Cin=>p(89)(47),clock=>clock,reset=>reset,s=>p(186)(47),cout=>p(187)(48));
FA_ff_3760:FAff port map(x=>p(87)(48),y=>p(88)(48),Cin=>p(89)(48),clock=>clock,reset=>reset,s=>p(186)(48),cout=>p(187)(49));
FA_ff_3761:FAff port map(x=>p(87)(49),y=>p(88)(49),Cin=>p(89)(49),clock=>clock,reset=>reset,s=>p(186)(49),cout=>p(187)(50));
FA_ff_3762:FAff port map(x=>p(87)(50),y=>p(88)(50),Cin=>p(89)(50),clock=>clock,reset=>reset,s=>p(186)(50),cout=>p(187)(51));
FA_ff_3763:FAff port map(x=>p(87)(51),y=>p(88)(51),Cin=>p(89)(51),clock=>clock,reset=>reset,s=>p(186)(51),cout=>p(187)(52));
FA_ff_3764:FAff port map(x=>p(87)(52),y=>p(88)(52),Cin=>p(89)(52),clock=>clock,reset=>reset,s=>p(186)(52),cout=>p(187)(53));
FA_ff_3765:FAff port map(x=>p(87)(53),y=>p(88)(53),Cin=>p(89)(53),clock=>clock,reset=>reset,s=>p(186)(53),cout=>p(187)(54));
FA_ff_3766:FAff port map(x=>p(87)(54),y=>p(88)(54),Cin=>p(89)(54),clock=>clock,reset=>reset,s=>p(186)(54),cout=>p(187)(55));
FA_ff_3767:FAff port map(x=>p(87)(55),y=>p(88)(55),Cin=>p(89)(55),clock=>clock,reset=>reset,s=>p(186)(55),cout=>p(187)(56));
FA_ff_3768:FAff port map(x=>p(87)(56),y=>p(88)(56),Cin=>p(89)(56),clock=>clock,reset=>reset,s=>p(186)(56),cout=>p(187)(57));
FA_ff_3769:FAff port map(x=>p(87)(57),y=>p(88)(57),Cin=>p(89)(57),clock=>clock,reset=>reset,s=>p(186)(57),cout=>p(187)(58));
FA_ff_3770:FAff port map(x=>p(87)(58),y=>p(88)(58),Cin=>p(89)(58),clock=>clock,reset=>reset,s=>p(186)(58),cout=>p(187)(59));
FA_ff_3771:FAff port map(x=>p(87)(59),y=>p(88)(59),Cin=>p(89)(59),clock=>clock,reset=>reset,s=>p(186)(59),cout=>p(187)(60));
FA_ff_3772:FAff port map(x=>p(87)(60),y=>p(88)(60),Cin=>p(89)(60),clock=>clock,reset=>reset,s=>p(186)(60),cout=>p(187)(61));
FA_ff_3773:FAff port map(x=>p(87)(61),y=>p(88)(61),Cin=>p(89)(61),clock=>clock,reset=>reset,s=>p(186)(61),cout=>p(187)(62));
FA_ff_3774:FAff port map(x=>p(87)(62),y=>p(88)(62),Cin=>p(89)(62),clock=>clock,reset=>reset,s=>p(186)(62),cout=>p(187)(63));
FA_ff_3775:FAff port map(x=>p(87)(63),y=>p(88)(63),Cin=>p(89)(63),clock=>clock,reset=>reset,s=>p(186)(63),cout=>p(187)(64));
FA_ff_3776:FAff port map(x=>p(87)(64),y=>p(88)(64),Cin=>p(89)(64),clock=>clock,reset=>reset,s=>p(186)(64),cout=>p(187)(65));
FA_ff_3777:FAff port map(x=>p(87)(65),y=>p(88)(65),Cin=>p(89)(65),clock=>clock,reset=>reset,s=>p(186)(65),cout=>p(187)(66));
FA_ff_3778:FAff port map(x=>p(87)(66),y=>p(88)(66),Cin=>p(89)(66),clock=>clock,reset=>reset,s=>p(186)(66),cout=>p(187)(67));
FA_ff_3779:FAff port map(x=>p(87)(67),y=>p(88)(67),Cin=>p(89)(67),clock=>clock,reset=>reset,s=>p(186)(67),cout=>p(187)(68));
FA_ff_3780:FAff port map(x=>p(87)(68),y=>p(88)(68),Cin=>p(89)(68),clock=>clock,reset=>reset,s=>p(186)(68),cout=>p(187)(69));
FA_ff_3781:FAff port map(x=>p(87)(69),y=>p(88)(69),Cin=>p(89)(69),clock=>clock,reset=>reset,s=>p(186)(69),cout=>p(187)(70));
FA_ff_3782:FAff port map(x=>p(87)(70),y=>p(88)(70),Cin=>p(89)(70),clock=>clock,reset=>reset,s=>p(186)(70),cout=>p(187)(71));
FA_ff_3783:FAff port map(x=>p(87)(71),y=>p(88)(71),Cin=>p(89)(71),clock=>clock,reset=>reset,s=>p(186)(71),cout=>p(187)(72));
FA_ff_3784:FAff port map(x=>p(87)(72),y=>p(88)(72),Cin=>p(89)(72),clock=>clock,reset=>reset,s=>p(186)(72),cout=>p(187)(73));
FA_ff_3785:FAff port map(x=>p(87)(73),y=>p(88)(73),Cin=>p(89)(73),clock=>clock,reset=>reset,s=>p(186)(73),cout=>p(187)(74));
FA_ff_3786:FAff port map(x=>p(87)(74),y=>p(88)(74),Cin=>p(89)(74),clock=>clock,reset=>reset,s=>p(186)(74),cout=>p(187)(75));
FA_ff_3787:FAff port map(x=>p(87)(75),y=>p(88)(75),Cin=>p(89)(75),clock=>clock,reset=>reset,s=>p(186)(75),cout=>p(187)(76));
FA_ff_3788:FAff port map(x=>p(87)(76),y=>p(88)(76),Cin=>p(89)(76),clock=>clock,reset=>reset,s=>p(186)(76),cout=>p(187)(77));
FA_ff_3789:FAff port map(x=>p(87)(77),y=>p(88)(77),Cin=>p(89)(77),clock=>clock,reset=>reset,s=>p(186)(77),cout=>p(187)(78));
FA_ff_3790:FAff port map(x=>p(87)(78),y=>p(88)(78),Cin=>p(89)(78),clock=>clock,reset=>reset,s=>p(186)(78),cout=>p(187)(79));
FA_ff_3791:FAff port map(x=>p(87)(79),y=>p(88)(79),Cin=>p(89)(79),clock=>clock,reset=>reset,s=>p(186)(79),cout=>p(187)(80));
FA_ff_3792:FAff port map(x=>p(87)(80),y=>p(88)(80),Cin=>p(89)(80),clock=>clock,reset=>reset,s=>p(186)(80),cout=>p(187)(81));
FA_ff_3793:FAff port map(x=>p(87)(81),y=>p(88)(81),Cin=>p(89)(81),clock=>clock,reset=>reset,s=>p(186)(81),cout=>p(187)(82));
FA_ff_3794:FAff port map(x=>p(87)(82),y=>p(88)(82),Cin=>p(89)(82),clock=>clock,reset=>reset,s=>p(186)(82),cout=>p(187)(83));
FA_ff_3795:FAff port map(x=>p(87)(83),y=>p(88)(83),Cin=>p(89)(83),clock=>clock,reset=>reset,s=>p(186)(83),cout=>p(187)(84));
FA_ff_3796:FAff port map(x=>p(87)(84),y=>p(88)(84),Cin=>p(89)(84),clock=>clock,reset=>reset,s=>p(186)(84),cout=>p(187)(85));
FA_ff_3797:FAff port map(x=>p(87)(85),y=>p(88)(85),Cin=>p(89)(85),clock=>clock,reset=>reset,s=>p(186)(85),cout=>p(187)(86));
FA_ff_3798:FAff port map(x=>p(87)(86),y=>p(88)(86),Cin=>p(89)(86),clock=>clock,reset=>reset,s=>p(186)(86),cout=>p(187)(87));
FA_ff_3799:FAff port map(x=>p(87)(87),y=>p(88)(87),Cin=>p(89)(87),clock=>clock,reset=>reset,s=>p(186)(87),cout=>p(187)(88));
FA_ff_3800:FAff port map(x=>p(87)(88),y=>p(88)(88),Cin=>p(89)(88),clock=>clock,reset=>reset,s=>p(186)(88),cout=>p(187)(89));
FA_ff_3801:FAff port map(x=>p(87)(89),y=>p(88)(89),Cin=>p(89)(89),clock=>clock,reset=>reset,s=>p(186)(89),cout=>p(187)(90));
FA_ff_3802:FAff port map(x=>p(87)(90),y=>p(88)(90),Cin=>p(89)(90),clock=>clock,reset=>reset,s=>p(186)(90),cout=>p(187)(91));
FA_ff_3803:FAff port map(x=>p(87)(91),y=>p(88)(91),Cin=>p(89)(91),clock=>clock,reset=>reset,s=>p(186)(91),cout=>p(187)(92));
FA_ff_3804:FAff port map(x=>p(87)(92),y=>p(88)(92),Cin=>p(89)(92),clock=>clock,reset=>reset,s=>p(186)(92),cout=>p(187)(93));
FA_ff_3805:FAff port map(x=>p(87)(93),y=>p(88)(93),Cin=>p(89)(93),clock=>clock,reset=>reset,s=>p(186)(93),cout=>p(187)(94));
FA_ff_3806:FAff port map(x=>p(87)(94),y=>p(88)(94),Cin=>p(89)(94),clock=>clock,reset=>reset,s=>p(186)(94),cout=>p(187)(95));
FA_ff_3807:FAff port map(x=>p(87)(95),y=>p(88)(95),Cin=>p(89)(95),clock=>clock,reset=>reset,s=>p(186)(95),cout=>p(187)(96));
FA_ff_3808:FAff port map(x=>p(87)(96),y=>p(88)(96),Cin=>p(89)(96),clock=>clock,reset=>reset,s=>p(186)(96),cout=>p(187)(97));
FA_ff_3809:FAff port map(x=>p(87)(97),y=>p(88)(97),Cin=>p(89)(97),clock=>clock,reset=>reset,s=>p(186)(97),cout=>p(187)(98));
FA_ff_3810:FAff port map(x=>p(87)(98),y=>p(88)(98),Cin=>p(89)(98),clock=>clock,reset=>reset,s=>p(186)(98),cout=>p(187)(99));
FA_ff_3811:FAff port map(x=>p(87)(99),y=>p(88)(99),Cin=>p(89)(99),clock=>clock,reset=>reset,s=>p(186)(99),cout=>p(187)(100));
FA_ff_3812:FAff port map(x=>p(87)(100),y=>p(88)(100),Cin=>p(89)(100),clock=>clock,reset=>reset,s=>p(186)(100),cout=>p(187)(101));
FA_ff_3813:FAff port map(x=>p(87)(101),y=>p(88)(101),Cin=>p(89)(101),clock=>clock,reset=>reset,s=>p(186)(101),cout=>p(187)(102));
FA_ff_3814:FAff port map(x=>p(87)(102),y=>p(88)(102),Cin=>p(89)(102),clock=>clock,reset=>reset,s=>p(186)(102),cout=>p(187)(103));
FA_ff_3815:FAff port map(x=>p(87)(103),y=>p(88)(103),Cin=>p(89)(103),clock=>clock,reset=>reset,s=>p(186)(103),cout=>p(187)(104));
FA_ff_3816:FAff port map(x=>p(87)(104),y=>p(88)(104),Cin=>p(89)(104),clock=>clock,reset=>reset,s=>p(186)(104),cout=>p(187)(105));
FA_ff_3817:FAff port map(x=>p(87)(105),y=>p(88)(105),Cin=>p(89)(105),clock=>clock,reset=>reset,s=>p(186)(105),cout=>p(187)(106));
FA_ff_3818:FAff port map(x=>p(87)(106),y=>p(88)(106),Cin=>p(89)(106),clock=>clock,reset=>reset,s=>p(186)(106),cout=>p(187)(107));
FA_ff_3819:FAff port map(x=>p(87)(107),y=>p(88)(107),Cin=>p(89)(107),clock=>clock,reset=>reset,s=>p(186)(107),cout=>p(187)(108));
FA_ff_3820:FAff port map(x=>p(87)(108),y=>p(88)(108),Cin=>p(89)(108),clock=>clock,reset=>reset,s=>p(186)(108),cout=>p(187)(109));
FA_ff_3821:FAff port map(x=>p(87)(109),y=>p(88)(109),Cin=>p(89)(109),clock=>clock,reset=>reset,s=>p(186)(109),cout=>p(187)(110));
FA_ff_3822:FAff port map(x=>p(87)(110),y=>p(88)(110),Cin=>p(89)(110),clock=>clock,reset=>reset,s=>p(186)(110),cout=>p(187)(111));
FA_ff_3823:FAff port map(x=>p(87)(111),y=>p(88)(111),Cin=>p(89)(111),clock=>clock,reset=>reset,s=>p(186)(111),cout=>p(187)(112));
FA_ff_3824:FAff port map(x=>p(87)(112),y=>p(88)(112),Cin=>p(89)(112),clock=>clock,reset=>reset,s=>p(186)(112),cout=>p(187)(113));
FA_ff_3825:FAff port map(x=>p(87)(113),y=>p(88)(113),Cin=>p(89)(113),clock=>clock,reset=>reset,s=>p(186)(113),cout=>p(187)(114));
FA_ff_3826:FAff port map(x=>p(87)(114),y=>p(88)(114),Cin=>p(89)(114),clock=>clock,reset=>reset,s=>p(186)(114),cout=>p(187)(115));
FA_ff_3827:FAff port map(x=>p(87)(115),y=>p(88)(115),Cin=>p(89)(115),clock=>clock,reset=>reset,s=>p(186)(115),cout=>p(187)(116));
FA_ff_3828:FAff port map(x=>p(87)(116),y=>p(88)(116),Cin=>p(89)(116),clock=>clock,reset=>reset,s=>p(186)(116),cout=>p(187)(117));
FA_ff_3829:FAff port map(x=>p(87)(117),y=>p(88)(117),Cin=>p(89)(117),clock=>clock,reset=>reset,s=>p(186)(117),cout=>p(187)(118));
FA_ff_3830:FAff port map(x=>p(87)(118),y=>p(88)(118),Cin=>p(89)(118),clock=>clock,reset=>reset,s=>p(186)(118),cout=>p(187)(119));
FA_ff_3831:FAff port map(x=>p(87)(119),y=>p(88)(119),Cin=>p(89)(119),clock=>clock,reset=>reset,s=>p(186)(119),cout=>p(187)(120));
FA_ff_3832:FAff port map(x=>p(87)(120),y=>p(88)(120),Cin=>p(89)(120),clock=>clock,reset=>reset,s=>p(186)(120),cout=>p(187)(121));
FA_ff_3833:FAff port map(x=>p(87)(121),y=>p(88)(121),Cin=>p(89)(121),clock=>clock,reset=>reset,s=>p(186)(121),cout=>p(187)(122));
FA_ff_3834:FAff port map(x=>p(87)(122),y=>p(88)(122),Cin=>p(89)(122),clock=>clock,reset=>reset,s=>p(186)(122),cout=>p(187)(123));
FA_ff_3835:FAff port map(x=>p(87)(123),y=>p(88)(123),Cin=>p(89)(123),clock=>clock,reset=>reset,s=>p(186)(123),cout=>p(187)(124));
FA_ff_3836:FAff port map(x=>p(87)(124),y=>p(88)(124),Cin=>p(89)(124),clock=>clock,reset=>reset,s=>p(186)(124),cout=>p(187)(125));
FA_ff_3837:FAff port map(x=>p(87)(125),y=>p(88)(125),Cin=>p(89)(125),clock=>clock,reset=>reset,s=>p(186)(125),cout=>p(187)(126));
FA_ff_3838:FAff port map(x=>p(87)(126),y=>p(88)(126),Cin=>p(89)(126),clock=>clock,reset=>reset,s=>p(186)(126),cout=>p(187)(127));
FA_ff_3839:FAff port map(x=>p(87)(127),y=>p(88)(127),Cin=>p(89)(127),clock=>clock,reset=>reset,s=>p(186)(127),cout=>p(187)(128));
FA_ff_3840:FAff port map(x=>p(90)(0),y=>p(91)(0),Cin=>p(92)(0),clock=>clock,reset=>reset,s=>p(188)(0),cout=>p(189)(1));
FA_ff_3841:FAff port map(x=>p(90)(1),y=>p(91)(1),Cin=>p(92)(1),clock=>clock,reset=>reset,s=>p(188)(1),cout=>p(189)(2));
FA_ff_3842:FAff port map(x=>p(90)(2),y=>p(91)(2),Cin=>p(92)(2),clock=>clock,reset=>reset,s=>p(188)(2),cout=>p(189)(3));
FA_ff_3843:FAff port map(x=>p(90)(3),y=>p(91)(3),Cin=>p(92)(3),clock=>clock,reset=>reset,s=>p(188)(3),cout=>p(189)(4));
FA_ff_3844:FAff port map(x=>p(90)(4),y=>p(91)(4),Cin=>p(92)(4),clock=>clock,reset=>reset,s=>p(188)(4),cout=>p(189)(5));
FA_ff_3845:FAff port map(x=>p(90)(5),y=>p(91)(5),Cin=>p(92)(5),clock=>clock,reset=>reset,s=>p(188)(5),cout=>p(189)(6));
FA_ff_3846:FAff port map(x=>p(90)(6),y=>p(91)(6),Cin=>p(92)(6),clock=>clock,reset=>reset,s=>p(188)(6),cout=>p(189)(7));
FA_ff_3847:FAff port map(x=>p(90)(7),y=>p(91)(7),Cin=>p(92)(7),clock=>clock,reset=>reset,s=>p(188)(7),cout=>p(189)(8));
FA_ff_3848:FAff port map(x=>p(90)(8),y=>p(91)(8),Cin=>p(92)(8),clock=>clock,reset=>reset,s=>p(188)(8),cout=>p(189)(9));
FA_ff_3849:FAff port map(x=>p(90)(9),y=>p(91)(9),Cin=>p(92)(9),clock=>clock,reset=>reset,s=>p(188)(9),cout=>p(189)(10));
FA_ff_3850:FAff port map(x=>p(90)(10),y=>p(91)(10),Cin=>p(92)(10),clock=>clock,reset=>reset,s=>p(188)(10),cout=>p(189)(11));
FA_ff_3851:FAff port map(x=>p(90)(11),y=>p(91)(11),Cin=>p(92)(11),clock=>clock,reset=>reset,s=>p(188)(11),cout=>p(189)(12));
FA_ff_3852:FAff port map(x=>p(90)(12),y=>p(91)(12),Cin=>p(92)(12),clock=>clock,reset=>reset,s=>p(188)(12),cout=>p(189)(13));
FA_ff_3853:FAff port map(x=>p(90)(13),y=>p(91)(13),Cin=>p(92)(13),clock=>clock,reset=>reset,s=>p(188)(13),cout=>p(189)(14));
FA_ff_3854:FAff port map(x=>p(90)(14),y=>p(91)(14),Cin=>p(92)(14),clock=>clock,reset=>reset,s=>p(188)(14),cout=>p(189)(15));
FA_ff_3855:FAff port map(x=>p(90)(15),y=>p(91)(15),Cin=>p(92)(15),clock=>clock,reset=>reset,s=>p(188)(15),cout=>p(189)(16));
FA_ff_3856:FAff port map(x=>p(90)(16),y=>p(91)(16),Cin=>p(92)(16),clock=>clock,reset=>reset,s=>p(188)(16),cout=>p(189)(17));
FA_ff_3857:FAff port map(x=>p(90)(17),y=>p(91)(17),Cin=>p(92)(17),clock=>clock,reset=>reset,s=>p(188)(17),cout=>p(189)(18));
FA_ff_3858:FAff port map(x=>p(90)(18),y=>p(91)(18),Cin=>p(92)(18),clock=>clock,reset=>reset,s=>p(188)(18),cout=>p(189)(19));
FA_ff_3859:FAff port map(x=>p(90)(19),y=>p(91)(19),Cin=>p(92)(19),clock=>clock,reset=>reset,s=>p(188)(19),cout=>p(189)(20));
FA_ff_3860:FAff port map(x=>p(90)(20),y=>p(91)(20),Cin=>p(92)(20),clock=>clock,reset=>reset,s=>p(188)(20),cout=>p(189)(21));
FA_ff_3861:FAff port map(x=>p(90)(21),y=>p(91)(21),Cin=>p(92)(21),clock=>clock,reset=>reset,s=>p(188)(21),cout=>p(189)(22));
FA_ff_3862:FAff port map(x=>p(90)(22),y=>p(91)(22),Cin=>p(92)(22),clock=>clock,reset=>reset,s=>p(188)(22),cout=>p(189)(23));
FA_ff_3863:FAff port map(x=>p(90)(23),y=>p(91)(23),Cin=>p(92)(23),clock=>clock,reset=>reset,s=>p(188)(23),cout=>p(189)(24));
FA_ff_3864:FAff port map(x=>p(90)(24),y=>p(91)(24),Cin=>p(92)(24),clock=>clock,reset=>reset,s=>p(188)(24),cout=>p(189)(25));
FA_ff_3865:FAff port map(x=>p(90)(25),y=>p(91)(25),Cin=>p(92)(25),clock=>clock,reset=>reset,s=>p(188)(25),cout=>p(189)(26));
FA_ff_3866:FAff port map(x=>p(90)(26),y=>p(91)(26),Cin=>p(92)(26),clock=>clock,reset=>reset,s=>p(188)(26),cout=>p(189)(27));
FA_ff_3867:FAff port map(x=>p(90)(27),y=>p(91)(27),Cin=>p(92)(27),clock=>clock,reset=>reset,s=>p(188)(27),cout=>p(189)(28));
FA_ff_3868:FAff port map(x=>p(90)(28),y=>p(91)(28),Cin=>p(92)(28),clock=>clock,reset=>reset,s=>p(188)(28),cout=>p(189)(29));
FA_ff_3869:FAff port map(x=>p(90)(29),y=>p(91)(29),Cin=>p(92)(29),clock=>clock,reset=>reset,s=>p(188)(29),cout=>p(189)(30));
FA_ff_3870:FAff port map(x=>p(90)(30),y=>p(91)(30),Cin=>p(92)(30),clock=>clock,reset=>reset,s=>p(188)(30),cout=>p(189)(31));
FA_ff_3871:FAff port map(x=>p(90)(31),y=>p(91)(31),Cin=>p(92)(31),clock=>clock,reset=>reset,s=>p(188)(31),cout=>p(189)(32));
FA_ff_3872:FAff port map(x=>p(90)(32),y=>p(91)(32),Cin=>p(92)(32),clock=>clock,reset=>reset,s=>p(188)(32),cout=>p(189)(33));
FA_ff_3873:FAff port map(x=>p(90)(33),y=>p(91)(33),Cin=>p(92)(33),clock=>clock,reset=>reset,s=>p(188)(33),cout=>p(189)(34));
FA_ff_3874:FAff port map(x=>p(90)(34),y=>p(91)(34),Cin=>p(92)(34),clock=>clock,reset=>reset,s=>p(188)(34),cout=>p(189)(35));
FA_ff_3875:FAff port map(x=>p(90)(35),y=>p(91)(35),Cin=>p(92)(35),clock=>clock,reset=>reset,s=>p(188)(35),cout=>p(189)(36));
FA_ff_3876:FAff port map(x=>p(90)(36),y=>p(91)(36),Cin=>p(92)(36),clock=>clock,reset=>reset,s=>p(188)(36),cout=>p(189)(37));
FA_ff_3877:FAff port map(x=>p(90)(37),y=>p(91)(37),Cin=>p(92)(37),clock=>clock,reset=>reset,s=>p(188)(37),cout=>p(189)(38));
FA_ff_3878:FAff port map(x=>p(90)(38),y=>p(91)(38),Cin=>p(92)(38),clock=>clock,reset=>reset,s=>p(188)(38),cout=>p(189)(39));
FA_ff_3879:FAff port map(x=>p(90)(39),y=>p(91)(39),Cin=>p(92)(39),clock=>clock,reset=>reset,s=>p(188)(39),cout=>p(189)(40));
FA_ff_3880:FAff port map(x=>p(90)(40),y=>p(91)(40),Cin=>p(92)(40),clock=>clock,reset=>reset,s=>p(188)(40),cout=>p(189)(41));
FA_ff_3881:FAff port map(x=>p(90)(41),y=>p(91)(41),Cin=>p(92)(41),clock=>clock,reset=>reset,s=>p(188)(41),cout=>p(189)(42));
FA_ff_3882:FAff port map(x=>p(90)(42),y=>p(91)(42),Cin=>p(92)(42),clock=>clock,reset=>reset,s=>p(188)(42),cout=>p(189)(43));
FA_ff_3883:FAff port map(x=>p(90)(43),y=>p(91)(43),Cin=>p(92)(43),clock=>clock,reset=>reset,s=>p(188)(43),cout=>p(189)(44));
FA_ff_3884:FAff port map(x=>p(90)(44),y=>p(91)(44),Cin=>p(92)(44),clock=>clock,reset=>reset,s=>p(188)(44),cout=>p(189)(45));
FA_ff_3885:FAff port map(x=>p(90)(45),y=>p(91)(45),Cin=>p(92)(45),clock=>clock,reset=>reset,s=>p(188)(45),cout=>p(189)(46));
FA_ff_3886:FAff port map(x=>p(90)(46),y=>p(91)(46),Cin=>p(92)(46),clock=>clock,reset=>reset,s=>p(188)(46),cout=>p(189)(47));
FA_ff_3887:FAff port map(x=>p(90)(47),y=>p(91)(47),Cin=>p(92)(47),clock=>clock,reset=>reset,s=>p(188)(47),cout=>p(189)(48));
FA_ff_3888:FAff port map(x=>p(90)(48),y=>p(91)(48),Cin=>p(92)(48),clock=>clock,reset=>reset,s=>p(188)(48),cout=>p(189)(49));
FA_ff_3889:FAff port map(x=>p(90)(49),y=>p(91)(49),Cin=>p(92)(49),clock=>clock,reset=>reset,s=>p(188)(49),cout=>p(189)(50));
FA_ff_3890:FAff port map(x=>p(90)(50),y=>p(91)(50),Cin=>p(92)(50),clock=>clock,reset=>reset,s=>p(188)(50),cout=>p(189)(51));
FA_ff_3891:FAff port map(x=>p(90)(51),y=>p(91)(51),Cin=>p(92)(51),clock=>clock,reset=>reset,s=>p(188)(51),cout=>p(189)(52));
FA_ff_3892:FAff port map(x=>p(90)(52),y=>p(91)(52),Cin=>p(92)(52),clock=>clock,reset=>reset,s=>p(188)(52),cout=>p(189)(53));
FA_ff_3893:FAff port map(x=>p(90)(53),y=>p(91)(53),Cin=>p(92)(53),clock=>clock,reset=>reset,s=>p(188)(53),cout=>p(189)(54));
FA_ff_3894:FAff port map(x=>p(90)(54),y=>p(91)(54),Cin=>p(92)(54),clock=>clock,reset=>reset,s=>p(188)(54),cout=>p(189)(55));
FA_ff_3895:FAff port map(x=>p(90)(55),y=>p(91)(55),Cin=>p(92)(55),clock=>clock,reset=>reset,s=>p(188)(55),cout=>p(189)(56));
FA_ff_3896:FAff port map(x=>p(90)(56),y=>p(91)(56),Cin=>p(92)(56),clock=>clock,reset=>reset,s=>p(188)(56),cout=>p(189)(57));
FA_ff_3897:FAff port map(x=>p(90)(57),y=>p(91)(57),Cin=>p(92)(57),clock=>clock,reset=>reset,s=>p(188)(57),cout=>p(189)(58));
FA_ff_3898:FAff port map(x=>p(90)(58),y=>p(91)(58),Cin=>p(92)(58),clock=>clock,reset=>reset,s=>p(188)(58),cout=>p(189)(59));
FA_ff_3899:FAff port map(x=>p(90)(59),y=>p(91)(59),Cin=>p(92)(59),clock=>clock,reset=>reset,s=>p(188)(59),cout=>p(189)(60));
FA_ff_3900:FAff port map(x=>p(90)(60),y=>p(91)(60),Cin=>p(92)(60),clock=>clock,reset=>reset,s=>p(188)(60),cout=>p(189)(61));
FA_ff_3901:FAff port map(x=>p(90)(61),y=>p(91)(61),Cin=>p(92)(61),clock=>clock,reset=>reset,s=>p(188)(61),cout=>p(189)(62));
FA_ff_3902:FAff port map(x=>p(90)(62),y=>p(91)(62),Cin=>p(92)(62),clock=>clock,reset=>reset,s=>p(188)(62),cout=>p(189)(63));
FA_ff_3903:FAff port map(x=>p(90)(63),y=>p(91)(63),Cin=>p(92)(63),clock=>clock,reset=>reset,s=>p(188)(63),cout=>p(189)(64));
FA_ff_3904:FAff port map(x=>p(90)(64),y=>p(91)(64),Cin=>p(92)(64),clock=>clock,reset=>reset,s=>p(188)(64),cout=>p(189)(65));
FA_ff_3905:FAff port map(x=>p(90)(65),y=>p(91)(65),Cin=>p(92)(65),clock=>clock,reset=>reset,s=>p(188)(65),cout=>p(189)(66));
FA_ff_3906:FAff port map(x=>p(90)(66),y=>p(91)(66),Cin=>p(92)(66),clock=>clock,reset=>reset,s=>p(188)(66),cout=>p(189)(67));
FA_ff_3907:FAff port map(x=>p(90)(67),y=>p(91)(67),Cin=>p(92)(67),clock=>clock,reset=>reset,s=>p(188)(67),cout=>p(189)(68));
FA_ff_3908:FAff port map(x=>p(90)(68),y=>p(91)(68),Cin=>p(92)(68),clock=>clock,reset=>reset,s=>p(188)(68),cout=>p(189)(69));
FA_ff_3909:FAff port map(x=>p(90)(69),y=>p(91)(69),Cin=>p(92)(69),clock=>clock,reset=>reset,s=>p(188)(69),cout=>p(189)(70));
FA_ff_3910:FAff port map(x=>p(90)(70),y=>p(91)(70),Cin=>p(92)(70),clock=>clock,reset=>reset,s=>p(188)(70),cout=>p(189)(71));
FA_ff_3911:FAff port map(x=>p(90)(71),y=>p(91)(71),Cin=>p(92)(71),clock=>clock,reset=>reset,s=>p(188)(71),cout=>p(189)(72));
FA_ff_3912:FAff port map(x=>p(90)(72),y=>p(91)(72),Cin=>p(92)(72),clock=>clock,reset=>reset,s=>p(188)(72),cout=>p(189)(73));
FA_ff_3913:FAff port map(x=>p(90)(73),y=>p(91)(73),Cin=>p(92)(73),clock=>clock,reset=>reset,s=>p(188)(73),cout=>p(189)(74));
FA_ff_3914:FAff port map(x=>p(90)(74),y=>p(91)(74),Cin=>p(92)(74),clock=>clock,reset=>reset,s=>p(188)(74),cout=>p(189)(75));
FA_ff_3915:FAff port map(x=>p(90)(75),y=>p(91)(75),Cin=>p(92)(75),clock=>clock,reset=>reset,s=>p(188)(75),cout=>p(189)(76));
FA_ff_3916:FAff port map(x=>p(90)(76),y=>p(91)(76),Cin=>p(92)(76),clock=>clock,reset=>reset,s=>p(188)(76),cout=>p(189)(77));
FA_ff_3917:FAff port map(x=>p(90)(77),y=>p(91)(77),Cin=>p(92)(77),clock=>clock,reset=>reset,s=>p(188)(77),cout=>p(189)(78));
FA_ff_3918:FAff port map(x=>p(90)(78),y=>p(91)(78),Cin=>p(92)(78),clock=>clock,reset=>reset,s=>p(188)(78),cout=>p(189)(79));
FA_ff_3919:FAff port map(x=>p(90)(79),y=>p(91)(79),Cin=>p(92)(79),clock=>clock,reset=>reset,s=>p(188)(79),cout=>p(189)(80));
FA_ff_3920:FAff port map(x=>p(90)(80),y=>p(91)(80),Cin=>p(92)(80),clock=>clock,reset=>reset,s=>p(188)(80),cout=>p(189)(81));
FA_ff_3921:FAff port map(x=>p(90)(81),y=>p(91)(81),Cin=>p(92)(81),clock=>clock,reset=>reset,s=>p(188)(81),cout=>p(189)(82));
FA_ff_3922:FAff port map(x=>p(90)(82),y=>p(91)(82),Cin=>p(92)(82),clock=>clock,reset=>reset,s=>p(188)(82),cout=>p(189)(83));
FA_ff_3923:FAff port map(x=>p(90)(83),y=>p(91)(83),Cin=>p(92)(83),clock=>clock,reset=>reset,s=>p(188)(83),cout=>p(189)(84));
FA_ff_3924:FAff port map(x=>p(90)(84),y=>p(91)(84),Cin=>p(92)(84),clock=>clock,reset=>reset,s=>p(188)(84),cout=>p(189)(85));
FA_ff_3925:FAff port map(x=>p(90)(85),y=>p(91)(85),Cin=>p(92)(85),clock=>clock,reset=>reset,s=>p(188)(85),cout=>p(189)(86));
FA_ff_3926:FAff port map(x=>p(90)(86),y=>p(91)(86),Cin=>p(92)(86),clock=>clock,reset=>reset,s=>p(188)(86),cout=>p(189)(87));
FA_ff_3927:FAff port map(x=>p(90)(87),y=>p(91)(87),Cin=>p(92)(87),clock=>clock,reset=>reset,s=>p(188)(87),cout=>p(189)(88));
FA_ff_3928:FAff port map(x=>p(90)(88),y=>p(91)(88),Cin=>p(92)(88),clock=>clock,reset=>reset,s=>p(188)(88),cout=>p(189)(89));
FA_ff_3929:FAff port map(x=>p(90)(89),y=>p(91)(89),Cin=>p(92)(89),clock=>clock,reset=>reset,s=>p(188)(89),cout=>p(189)(90));
FA_ff_3930:FAff port map(x=>p(90)(90),y=>p(91)(90),Cin=>p(92)(90),clock=>clock,reset=>reset,s=>p(188)(90),cout=>p(189)(91));
FA_ff_3931:FAff port map(x=>p(90)(91),y=>p(91)(91),Cin=>p(92)(91),clock=>clock,reset=>reset,s=>p(188)(91),cout=>p(189)(92));
FA_ff_3932:FAff port map(x=>p(90)(92),y=>p(91)(92),Cin=>p(92)(92),clock=>clock,reset=>reset,s=>p(188)(92),cout=>p(189)(93));
FA_ff_3933:FAff port map(x=>p(90)(93),y=>p(91)(93),Cin=>p(92)(93),clock=>clock,reset=>reset,s=>p(188)(93),cout=>p(189)(94));
FA_ff_3934:FAff port map(x=>p(90)(94),y=>p(91)(94),Cin=>p(92)(94),clock=>clock,reset=>reset,s=>p(188)(94),cout=>p(189)(95));
FA_ff_3935:FAff port map(x=>p(90)(95),y=>p(91)(95),Cin=>p(92)(95),clock=>clock,reset=>reset,s=>p(188)(95),cout=>p(189)(96));
FA_ff_3936:FAff port map(x=>p(90)(96),y=>p(91)(96),Cin=>p(92)(96),clock=>clock,reset=>reset,s=>p(188)(96),cout=>p(189)(97));
FA_ff_3937:FAff port map(x=>p(90)(97),y=>p(91)(97),Cin=>p(92)(97),clock=>clock,reset=>reset,s=>p(188)(97),cout=>p(189)(98));
FA_ff_3938:FAff port map(x=>p(90)(98),y=>p(91)(98),Cin=>p(92)(98),clock=>clock,reset=>reset,s=>p(188)(98),cout=>p(189)(99));
FA_ff_3939:FAff port map(x=>p(90)(99),y=>p(91)(99),Cin=>p(92)(99),clock=>clock,reset=>reset,s=>p(188)(99),cout=>p(189)(100));
FA_ff_3940:FAff port map(x=>p(90)(100),y=>p(91)(100),Cin=>p(92)(100),clock=>clock,reset=>reset,s=>p(188)(100),cout=>p(189)(101));
FA_ff_3941:FAff port map(x=>p(90)(101),y=>p(91)(101),Cin=>p(92)(101),clock=>clock,reset=>reset,s=>p(188)(101),cout=>p(189)(102));
FA_ff_3942:FAff port map(x=>p(90)(102),y=>p(91)(102),Cin=>p(92)(102),clock=>clock,reset=>reset,s=>p(188)(102),cout=>p(189)(103));
FA_ff_3943:FAff port map(x=>p(90)(103),y=>p(91)(103),Cin=>p(92)(103),clock=>clock,reset=>reset,s=>p(188)(103),cout=>p(189)(104));
FA_ff_3944:FAff port map(x=>p(90)(104),y=>p(91)(104),Cin=>p(92)(104),clock=>clock,reset=>reset,s=>p(188)(104),cout=>p(189)(105));
FA_ff_3945:FAff port map(x=>p(90)(105),y=>p(91)(105),Cin=>p(92)(105),clock=>clock,reset=>reset,s=>p(188)(105),cout=>p(189)(106));
FA_ff_3946:FAff port map(x=>p(90)(106),y=>p(91)(106),Cin=>p(92)(106),clock=>clock,reset=>reset,s=>p(188)(106),cout=>p(189)(107));
FA_ff_3947:FAff port map(x=>p(90)(107),y=>p(91)(107),Cin=>p(92)(107),clock=>clock,reset=>reset,s=>p(188)(107),cout=>p(189)(108));
FA_ff_3948:FAff port map(x=>p(90)(108),y=>p(91)(108),Cin=>p(92)(108),clock=>clock,reset=>reset,s=>p(188)(108),cout=>p(189)(109));
FA_ff_3949:FAff port map(x=>p(90)(109),y=>p(91)(109),Cin=>p(92)(109),clock=>clock,reset=>reset,s=>p(188)(109),cout=>p(189)(110));
FA_ff_3950:FAff port map(x=>p(90)(110),y=>p(91)(110),Cin=>p(92)(110),clock=>clock,reset=>reset,s=>p(188)(110),cout=>p(189)(111));
FA_ff_3951:FAff port map(x=>p(90)(111),y=>p(91)(111),Cin=>p(92)(111),clock=>clock,reset=>reset,s=>p(188)(111),cout=>p(189)(112));
FA_ff_3952:FAff port map(x=>p(90)(112),y=>p(91)(112),Cin=>p(92)(112),clock=>clock,reset=>reset,s=>p(188)(112),cout=>p(189)(113));
FA_ff_3953:FAff port map(x=>p(90)(113),y=>p(91)(113),Cin=>p(92)(113),clock=>clock,reset=>reset,s=>p(188)(113),cout=>p(189)(114));
FA_ff_3954:FAff port map(x=>p(90)(114),y=>p(91)(114),Cin=>p(92)(114),clock=>clock,reset=>reset,s=>p(188)(114),cout=>p(189)(115));
FA_ff_3955:FAff port map(x=>p(90)(115),y=>p(91)(115),Cin=>p(92)(115),clock=>clock,reset=>reset,s=>p(188)(115),cout=>p(189)(116));
FA_ff_3956:FAff port map(x=>p(90)(116),y=>p(91)(116),Cin=>p(92)(116),clock=>clock,reset=>reset,s=>p(188)(116),cout=>p(189)(117));
FA_ff_3957:FAff port map(x=>p(90)(117),y=>p(91)(117),Cin=>p(92)(117),clock=>clock,reset=>reset,s=>p(188)(117),cout=>p(189)(118));
FA_ff_3958:FAff port map(x=>p(90)(118),y=>p(91)(118),Cin=>p(92)(118),clock=>clock,reset=>reset,s=>p(188)(118),cout=>p(189)(119));
FA_ff_3959:FAff port map(x=>p(90)(119),y=>p(91)(119),Cin=>p(92)(119),clock=>clock,reset=>reset,s=>p(188)(119),cout=>p(189)(120));
FA_ff_3960:FAff port map(x=>p(90)(120),y=>p(91)(120),Cin=>p(92)(120),clock=>clock,reset=>reset,s=>p(188)(120),cout=>p(189)(121));
FA_ff_3961:FAff port map(x=>p(90)(121),y=>p(91)(121),Cin=>p(92)(121),clock=>clock,reset=>reset,s=>p(188)(121),cout=>p(189)(122));
FA_ff_3962:FAff port map(x=>p(90)(122),y=>p(91)(122),Cin=>p(92)(122),clock=>clock,reset=>reset,s=>p(188)(122),cout=>p(189)(123));
FA_ff_3963:FAff port map(x=>p(90)(123),y=>p(91)(123),Cin=>p(92)(123),clock=>clock,reset=>reset,s=>p(188)(123),cout=>p(189)(124));
FA_ff_3964:FAff port map(x=>p(90)(124),y=>p(91)(124),Cin=>p(92)(124),clock=>clock,reset=>reset,s=>p(188)(124),cout=>p(189)(125));
FA_ff_3965:FAff port map(x=>p(90)(125),y=>p(91)(125),Cin=>p(92)(125),clock=>clock,reset=>reset,s=>p(188)(125),cout=>p(189)(126));
FA_ff_3966:FAff port map(x=>p(90)(126),y=>p(91)(126),Cin=>p(92)(126),clock=>clock,reset=>reset,s=>p(188)(126),cout=>p(189)(127));
FA_ff_3967:FAff port map(x=>p(90)(127),y=>p(91)(127),Cin=>p(92)(127),clock=>clock,reset=>reset,s=>p(188)(127),cout=>p(189)(128));
FA_ff_3968:FAff port map(x=>p(93)(0),y=>p(94)(0),Cin=>p(95)(0),clock=>clock,reset=>reset,s=>p(190)(0),cout=>p(191)(1));
FA_ff_3969:FAff port map(x=>p(93)(1),y=>p(94)(1),Cin=>p(95)(1),clock=>clock,reset=>reset,s=>p(190)(1),cout=>p(191)(2));
FA_ff_3970:FAff port map(x=>p(93)(2),y=>p(94)(2),Cin=>p(95)(2),clock=>clock,reset=>reset,s=>p(190)(2),cout=>p(191)(3));
FA_ff_3971:FAff port map(x=>p(93)(3),y=>p(94)(3),Cin=>p(95)(3),clock=>clock,reset=>reset,s=>p(190)(3),cout=>p(191)(4));
FA_ff_3972:FAff port map(x=>p(93)(4),y=>p(94)(4),Cin=>p(95)(4),clock=>clock,reset=>reset,s=>p(190)(4),cout=>p(191)(5));
FA_ff_3973:FAff port map(x=>p(93)(5),y=>p(94)(5),Cin=>p(95)(5),clock=>clock,reset=>reset,s=>p(190)(5),cout=>p(191)(6));
FA_ff_3974:FAff port map(x=>p(93)(6),y=>p(94)(6),Cin=>p(95)(6),clock=>clock,reset=>reset,s=>p(190)(6),cout=>p(191)(7));
FA_ff_3975:FAff port map(x=>p(93)(7),y=>p(94)(7),Cin=>p(95)(7),clock=>clock,reset=>reset,s=>p(190)(7),cout=>p(191)(8));
FA_ff_3976:FAff port map(x=>p(93)(8),y=>p(94)(8),Cin=>p(95)(8),clock=>clock,reset=>reset,s=>p(190)(8),cout=>p(191)(9));
FA_ff_3977:FAff port map(x=>p(93)(9),y=>p(94)(9),Cin=>p(95)(9),clock=>clock,reset=>reset,s=>p(190)(9),cout=>p(191)(10));
FA_ff_3978:FAff port map(x=>p(93)(10),y=>p(94)(10),Cin=>p(95)(10),clock=>clock,reset=>reset,s=>p(190)(10),cout=>p(191)(11));
FA_ff_3979:FAff port map(x=>p(93)(11),y=>p(94)(11),Cin=>p(95)(11),clock=>clock,reset=>reset,s=>p(190)(11),cout=>p(191)(12));
FA_ff_3980:FAff port map(x=>p(93)(12),y=>p(94)(12),Cin=>p(95)(12),clock=>clock,reset=>reset,s=>p(190)(12),cout=>p(191)(13));
FA_ff_3981:FAff port map(x=>p(93)(13),y=>p(94)(13),Cin=>p(95)(13),clock=>clock,reset=>reset,s=>p(190)(13),cout=>p(191)(14));
FA_ff_3982:FAff port map(x=>p(93)(14),y=>p(94)(14),Cin=>p(95)(14),clock=>clock,reset=>reset,s=>p(190)(14),cout=>p(191)(15));
FA_ff_3983:FAff port map(x=>p(93)(15),y=>p(94)(15),Cin=>p(95)(15),clock=>clock,reset=>reset,s=>p(190)(15),cout=>p(191)(16));
FA_ff_3984:FAff port map(x=>p(93)(16),y=>p(94)(16),Cin=>p(95)(16),clock=>clock,reset=>reset,s=>p(190)(16),cout=>p(191)(17));
FA_ff_3985:FAff port map(x=>p(93)(17),y=>p(94)(17),Cin=>p(95)(17),clock=>clock,reset=>reset,s=>p(190)(17),cout=>p(191)(18));
FA_ff_3986:FAff port map(x=>p(93)(18),y=>p(94)(18),Cin=>p(95)(18),clock=>clock,reset=>reset,s=>p(190)(18),cout=>p(191)(19));
FA_ff_3987:FAff port map(x=>p(93)(19),y=>p(94)(19),Cin=>p(95)(19),clock=>clock,reset=>reset,s=>p(190)(19),cout=>p(191)(20));
FA_ff_3988:FAff port map(x=>p(93)(20),y=>p(94)(20),Cin=>p(95)(20),clock=>clock,reset=>reset,s=>p(190)(20),cout=>p(191)(21));
FA_ff_3989:FAff port map(x=>p(93)(21),y=>p(94)(21),Cin=>p(95)(21),clock=>clock,reset=>reset,s=>p(190)(21),cout=>p(191)(22));
FA_ff_3990:FAff port map(x=>p(93)(22),y=>p(94)(22),Cin=>p(95)(22),clock=>clock,reset=>reset,s=>p(190)(22),cout=>p(191)(23));
FA_ff_3991:FAff port map(x=>p(93)(23),y=>p(94)(23),Cin=>p(95)(23),clock=>clock,reset=>reset,s=>p(190)(23),cout=>p(191)(24));
FA_ff_3992:FAff port map(x=>p(93)(24),y=>p(94)(24),Cin=>p(95)(24),clock=>clock,reset=>reset,s=>p(190)(24),cout=>p(191)(25));
FA_ff_3993:FAff port map(x=>p(93)(25),y=>p(94)(25),Cin=>p(95)(25),clock=>clock,reset=>reset,s=>p(190)(25),cout=>p(191)(26));
FA_ff_3994:FAff port map(x=>p(93)(26),y=>p(94)(26),Cin=>p(95)(26),clock=>clock,reset=>reset,s=>p(190)(26),cout=>p(191)(27));
FA_ff_3995:FAff port map(x=>p(93)(27),y=>p(94)(27),Cin=>p(95)(27),clock=>clock,reset=>reset,s=>p(190)(27),cout=>p(191)(28));
FA_ff_3996:FAff port map(x=>p(93)(28),y=>p(94)(28),Cin=>p(95)(28),clock=>clock,reset=>reset,s=>p(190)(28),cout=>p(191)(29));
FA_ff_3997:FAff port map(x=>p(93)(29),y=>p(94)(29),Cin=>p(95)(29),clock=>clock,reset=>reset,s=>p(190)(29),cout=>p(191)(30));
FA_ff_3998:FAff port map(x=>p(93)(30),y=>p(94)(30),Cin=>p(95)(30),clock=>clock,reset=>reset,s=>p(190)(30),cout=>p(191)(31));
FA_ff_3999:FAff port map(x=>p(93)(31),y=>p(94)(31),Cin=>p(95)(31),clock=>clock,reset=>reset,s=>p(190)(31),cout=>p(191)(32));
FA_ff_4000:FAff port map(x=>p(93)(32),y=>p(94)(32),Cin=>p(95)(32),clock=>clock,reset=>reset,s=>p(190)(32),cout=>p(191)(33));
FA_ff_4001:FAff port map(x=>p(93)(33),y=>p(94)(33),Cin=>p(95)(33),clock=>clock,reset=>reset,s=>p(190)(33),cout=>p(191)(34));
FA_ff_4002:FAff port map(x=>p(93)(34),y=>p(94)(34),Cin=>p(95)(34),clock=>clock,reset=>reset,s=>p(190)(34),cout=>p(191)(35));
FA_ff_4003:FAff port map(x=>p(93)(35),y=>p(94)(35),Cin=>p(95)(35),clock=>clock,reset=>reset,s=>p(190)(35),cout=>p(191)(36));
FA_ff_4004:FAff port map(x=>p(93)(36),y=>p(94)(36),Cin=>p(95)(36),clock=>clock,reset=>reset,s=>p(190)(36),cout=>p(191)(37));
FA_ff_4005:FAff port map(x=>p(93)(37),y=>p(94)(37),Cin=>p(95)(37),clock=>clock,reset=>reset,s=>p(190)(37),cout=>p(191)(38));
FA_ff_4006:FAff port map(x=>p(93)(38),y=>p(94)(38),Cin=>p(95)(38),clock=>clock,reset=>reset,s=>p(190)(38),cout=>p(191)(39));
FA_ff_4007:FAff port map(x=>p(93)(39),y=>p(94)(39),Cin=>p(95)(39),clock=>clock,reset=>reset,s=>p(190)(39),cout=>p(191)(40));
FA_ff_4008:FAff port map(x=>p(93)(40),y=>p(94)(40),Cin=>p(95)(40),clock=>clock,reset=>reset,s=>p(190)(40),cout=>p(191)(41));
FA_ff_4009:FAff port map(x=>p(93)(41),y=>p(94)(41),Cin=>p(95)(41),clock=>clock,reset=>reset,s=>p(190)(41),cout=>p(191)(42));
FA_ff_4010:FAff port map(x=>p(93)(42),y=>p(94)(42),Cin=>p(95)(42),clock=>clock,reset=>reset,s=>p(190)(42),cout=>p(191)(43));
FA_ff_4011:FAff port map(x=>p(93)(43),y=>p(94)(43),Cin=>p(95)(43),clock=>clock,reset=>reset,s=>p(190)(43),cout=>p(191)(44));
FA_ff_4012:FAff port map(x=>p(93)(44),y=>p(94)(44),Cin=>p(95)(44),clock=>clock,reset=>reset,s=>p(190)(44),cout=>p(191)(45));
FA_ff_4013:FAff port map(x=>p(93)(45),y=>p(94)(45),Cin=>p(95)(45),clock=>clock,reset=>reset,s=>p(190)(45),cout=>p(191)(46));
FA_ff_4014:FAff port map(x=>p(93)(46),y=>p(94)(46),Cin=>p(95)(46),clock=>clock,reset=>reset,s=>p(190)(46),cout=>p(191)(47));
FA_ff_4015:FAff port map(x=>p(93)(47),y=>p(94)(47),Cin=>p(95)(47),clock=>clock,reset=>reset,s=>p(190)(47),cout=>p(191)(48));
FA_ff_4016:FAff port map(x=>p(93)(48),y=>p(94)(48),Cin=>p(95)(48),clock=>clock,reset=>reset,s=>p(190)(48),cout=>p(191)(49));
FA_ff_4017:FAff port map(x=>p(93)(49),y=>p(94)(49),Cin=>p(95)(49),clock=>clock,reset=>reset,s=>p(190)(49),cout=>p(191)(50));
FA_ff_4018:FAff port map(x=>p(93)(50),y=>p(94)(50),Cin=>p(95)(50),clock=>clock,reset=>reset,s=>p(190)(50),cout=>p(191)(51));
FA_ff_4019:FAff port map(x=>p(93)(51),y=>p(94)(51),Cin=>p(95)(51),clock=>clock,reset=>reset,s=>p(190)(51),cout=>p(191)(52));
FA_ff_4020:FAff port map(x=>p(93)(52),y=>p(94)(52),Cin=>p(95)(52),clock=>clock,reset=>reset,s=>p(190)(52),cout=>p(191)(53));
FA_ff_4021:FAff port map(x=>p(93)(53),y=>p(94)(53),Cin=>p(95)(53),clock=>clock,reset=>reset,s=>p(190)(53),cout=>p(191)(54));
FA_ff_4022:FAff port map(x=>p(93)(54),y=>p(94)(54),Cin=>p(95)(54),clock=>clock,reset=>reset,s=>p(190)(54),cout=>p(191)(55));
FA_ff_4023:FAff port map(x=>p(93)(55),y=>p(94)(55),Cin=>p(95)(55),clock=>clock,reset=>reset,s=>p(190)(55),cout=>p(191)(56));
FA_ff_4024:FAff port map(x=>p(93)(56),y=>p(94)(56),Cin=>p(95)(56),clock=>clock,reset=>reset,s=>p(190)(56),cout=>p(191)(57));
FA_ff_4025:FAff port map(x=>p(93)(57),y=>p(94)(57),Cin=>p(95)(57),clock=>clock,reset=>reset,s=>p(190)(57),cout=>p(191)(58));
FA_ff_4026:FAff port map(x=>p(93)(58),y=>p(94)(58),Cin=>p(95)(58),clock=>clock,reset=>reset,s=>p(190)(58),cout=>p(191)(59));
FA_ff_4027:FAff port map(x=>p(93)(59),y=>p(94)(59),Cin=>p(95)(59),clock=>clock,reset=>reset,s=>p(190)(59),cout=>p(191)(60));
FA_ff_4028:FAff port map(x=>p(93)(60),y=>p(94)(60),Cin=>p(95)(60),clock=>clock,reset=>reset,s=>p(190)(60),cout=>p(191)(61));
FA_ff_4029:FAff port map(x=>p(93)(61),y=>p(94)(61),Cin=>p(95)(61),clock=>clock,reset=>reset,s=>p(190)(61),cout=>p(191)(62));
FA_ff_4030:FAff port map(x=>p(93)(62),y=>p(94)(62),Cin=>p(95)(62),clock=>clock,reset=>reset,s=>p(190)(62),cout=>p(191)(63));
FA_ff_4031:FAff port map(x=>p(93)(63),y=>p(94)(63),Cin=>p(95)(63),clock=>clock,reset=>reset,s=>p(190)(63),cout=>p(191)(64));
FA_ff_4032:FAff port map(x=>p(93)(64),y=>p(94)(64),Cin=>p(95)(64),clock=>clock,reset=>reset,s=>p(190)(64),cout=>p(191)(65));
FA_ff_4033:FAff port map(x=>p(93)(65),y=>p(94)(65),Cin=>p(95)(65),clock=>clock,reset=>reset,s=>p(190)(65),cout=>p(191)(66));
FA_ff_4034:FAff port map(x=>p(93)(66),y=>p(94)(66),Cin=>p(95)(66),clock=>clock,reset=>reset,s=>p(190)(66),cout=>p(191)(67));
FA_ff_4035:FAff port map(x=>p(93)(67),y=>p(94)(67),Cin=>p(95)(67),clock=>clock,reset=>reset,s=>p(190)(67),cout=>p(191)(68));
FA_ff_4036:FAff port map(x=>p(93)(68),y=>p(94)(68),Cin=>p(95)(68),clock=>clock,reset=>reset,s=>p(190)(68),cout=>p(191)(69));
FA_ff_4037:FAff port map(x=>p(93)(69),y=>p(94)(69),Cin=>p(95)(69),clock=>clock,reset=>reset,s=>p(190)(69),cout=>p(191)(70));
FA_ff_4038:FAff port map(x=>p(93)(70),y=>p(94)(70),Cin=>p(95)(70),clock=>clock,reset=>reset,s=>p(190)(70),cout=>p(191)(71));
FA_ff_4039:FAff port map(x=>p(93)(71),y=>p(94)(71),Cin=>p(95)(71),clock=>clock,reset=>reset,s=>p(190)(71),cout=>p(191)(72));
FA_ff_4040:FAff port map(x=>p(93)(72),y=>p(94)(72),Cin=>p(95)(72),clock=>clock,reset=>reset,s=>p(190)(72),cout=>p(191)(73));
FA_ff_4041:FAff port map(x=>p(93)(73),y=>p(94)(73),Cin=>p(95)(73),clock=>clock,reset=>reset,s=>p(190)(73),cout=>p(191)(74));
FA_ff_4042:FAff port map(x=>p(93)(74),y=>p(94)(74),Cin=>p(95)(74),clock=>clock,reset=>reset,s=>p(190)(74),cout=>p(191)(75));
FA_ff_4043:FAff port map(x=>p(93)(75),y=>p(94)(75),Cin=>p(95)(75),clock=>clock,reset=>reset,s=>p(190)(75),cout=>p(191)(76));
FA_ff_4044:FAff port map(x=>p(93)(76),y=>p(94)(76),Cin=>p(95)(76),clock=>clock,reset=>reset,s=>p(190)(76),cout=>p(191)(77));
FA_ff_4045:FAff port map(x=>p(93)(77),y=>p(94)(77),Cin=>p(95)(77),clock=>clock,reset=>reset,s=>p(190)(77),cout=>p(191)(78));
FA_ff_4046:FAff port map(x=>p(93)(78),y=>p(94)(78),Cin=>p(95)(78),clock=>clock,reset=>reset,s=>p(190)(78),cout=>p(191)(79));
FA_ff_4047:FAff port map(x=>p(93)(79),y=>p(94)(79),Cin=>p(95)(79),clock=>clock,reset=>reset,s=>p(190)(79),cout=>p(191)(80));
FA_ff_4048:FAff port map(x=>p(93)(80),y=>p(94)(80),Cin=>p(95)(80),clock=>clock,reset=>reset,s=>p(190)(80),cout=>p(191)(81));
FA_ff_4049:FAff port map(x=>p(93)(81),y=>p(94)(81),Cin=>p(95)(81),clock=>clock,reset=>reset,s=>p(190)(81),cout=>p(191)(82));
FA_ff_4050:FAff port map(x=>p(93)(82),y=>p(94)(82),Cin=>p(95)(82),clock=>clock,reset=>reset,s=>p(190)(82),cout=>p(191)(83));
FA_ff_4051:FAff port map(x=>p(93)(83),y=>p(94)(83),Cin=>p(95)(83),clock=>clock,reset=>reset,s=>p(190)(83),cout=>p(191)(84));
FA_ff_4052:FAff port map(x=>p(93)(84),y=>p(94)(84),Cin=>p(95)(84),clock=>clock,reset=>reset,s=>p(190)(84),cout=>p(191)(85));
FA_ff_4053:FAff port map(x=>p(93)(85),y=>p(94)(85),Cin=>p(95)(85),clock=>clock,reset=>reset,s=>p(190)(85),cout=>p(191)(86));
FA_ff_4054:FAff port map(x=>p(93)(86),y=>p(94)(86),Cin=>p(95)(86),clock=>clock,reset=>reset,s=>p(190)(86),cout=>p(191)(87));
FA_ff_4055:FAff port map(x=>p(93)(87),y=>p(94)(87),Cin=>p(95)(87),clock=>clock,reset=>reset,s=>p(190)(87),cout=>p(191)(88));
FA_ff_4056:FAff port map(x=>p(93)(88),y=>p(94)(88),Cin=>p(95)(88),clock=>clock,reset=>reset,s=>p(190)(88),cout=>p(191)(89));
FA_ff_4057:FAff port map(x=>p(93)(89),y=>p(94)(89),Cin=>p(95)(89),clock=>clock,reset=>reset,s=>p(190)(89),cout=>p(191)(90));
FA_ff_4058:FAff port map(x=>p(93)(90),y=>p(94)(90),Cin=>p(95)(90),clock=>clock,reset=>reset,s=>p(190)(90),cout=>p(191)(91));
FA_ff_4059:FAff port map(x=>p(93)(91),y=>p(94)(91),Cin=>p(95)(91),clock=>clock,reset=>reset,s=>p(190)(91),cout=>p(191)(92));
FA_ff_4060:FAff port map(x=>p(93)(92),y=>p(94)(92),Cin=>p(95)(92),clock=>clock,reset=>reset,s=>p(190)(92),cout=>p(191)(93));
FA_ff_4061:FAff port map(x=>p(93)(93),y=>p(94)(93),Cin=>p(95)(93),clock=>clock,reset=>reset,s=>p(190)(93),cout=>p(191)(94));
FA_ff_4062:FAff port map(x=>p(93)(94),y=>p(94)(94),Cin=>p(95)(94),clock=>clock,reset=>reset,s=>p(190)(94),cout=>p(191)(95));
FA_ff_4063:FAff port map(x=>p(93)(95),y=>p(94)(95),Cin=>p(95)(95),clock=>clock,reset=>reset,s=>p(190)(95),cout=>p(191)(96));
FA_ff_4064:FAff port map(x=>p(93)(96),y=>p(94)(96),Cin=>p(95)(96),clock=>clock,reset=>reset,s=>p(190)(96),cout=>p(191)(97));
FA_ff_4065:FAff port map(x=>p(93)(97),y=>p(94)(97),Cin=>p(95)(97),clock=>clock,reset=>reset,s=>p(190)(97),cout=>p(191)(98));
FA_ff_4066:FAff port map(x=>p(93)(98),y=>p(94)(98),Cin=>p(95)(98),clock=>clock,reset=>reset,s=>p(190)(98),cout=>p(191)(99));
FA_ff_4067:FAff port map(x=>p(93)(99),y=>p(94)(99),Cin=>p(95)(99),clock=>clock,reset=>reset,s=>p(190)(99),cout=>p(191)(100));
FA_ff_4068:FAff port map(x=>p(93)(100),y=>p(94)(100),Cin=>p(95)(100),clock=>clock,reset=>reset,s=>p(190)(100),cout=>p(191)(101));
FA_ff_4069:FAff port map(x=>p(93)(101),y=>p(94)(101),Cin=>p(95)(101),clock=>clock,reset=>reset,s=>p(190)(101),cout=>p(191)(102));
FA_ff_4070:FAff port map(x=>p(93)(102),y=>p(94)(102),Cin=>p(95)(102),clock=>clock,reset=>reset,s=>p(190)(102),cout=>p(191)(103));
FA_ff_4071:FAff port map(x=>p(93)(103),y=>p(94)(103),Cin=>p(95)(103),clock=>clock,reset=>reset,s=>p(190)(103),cout=>p(191)(104));
FA_ff_4072:FAff port map(x=>p(93)(104),y=>p(94)(104),Cin=>p(95)(104),clock=>clock,reset=>reset,s=>p(190)(104),cout=>p(191)(105));
FA_ff_4073:FAff port map(x=>p(93)(105),y=>p(94)(105),Cin=>p(95)(105),clock=>clock,reset=>reset,s=>p(190)(105),cout=>p(191)(106));
FA_ff_4074:FAff port map(x=>p(93)(106),y=>p(94)(106),Cin=>p(95)(106),clock=>clock,reset=>reset,s=>p(190)(106),cout=>p(191)(107));
FA_ff_4075:FAff port map(x=>p(93)(107),y=>p(94)(107),Cin=>p(95)(107),clock=>clock,reset=>reset,s=>p(190)(107),cout=>p(191)(108));
FA_ff_4076:FAff port map(x=>p(93)(108),y=>p(94)(108),Cin=>p(95)(108),clock=>clock,reset=>reset,s=>p(190)(108),cout=>p(191)(109));
FA_ff_4077:FAff port map(x=>p(93)(109),y=>p(94)(109),Cin=>p(95)(109),clock=>clock,reset=>reset,s=>p(190)(109),cout=>p(191)(110));
FA_ff_4078:FAff port map(x=>p(93)(110),y=>p(94)(110),Cin=>p(95)(110),clock=>clock,reset=>reset,s=>p(190)(110),cout=>p(191)(111));
FA_ff_4079:FAff port map(x=>p(93)(111),y=>p(94)(111),Cin=>p(95)(111),clock=>clock,reset=>reset,s=>p(190)(111),cout=>p(191)(112));
FA_ff_4080:FAff port map(x=>p(93)(112),y=>p(94)(112),Cin=>p(95)(112),clock=>clock,reset=>reset,s=>p(190)(112),cout=>p(191)(113));
FA_ff_4081:FAff port map(x=>p(93)(113),y=>p(94)(113),Cin=>p(95)(113),clock=>clock,reset=>reset,s=>p(190)(113),cout=>p(191)(114));
FA_ff_4082:FAff port map(x=>p(93)(114),y=>p(94)(114),Cin=>p(95)(114),clock=>clock,reset=>reset,s=>p(190)(114),cout=>p(191)(115));
FA_ff_4083:FAff port map(x=>p(93)(115),y=>p(94)(115),Cin=>p(95)(115),clock=>clock,reset=>reset,s=>p(190)(115),cout=>p(191)(116));
FA_ff_4084:FAff port map(x=>p(93)(116),y=>p(94)(116),Cin=>p(95)(116),clock=>clock,reset=>reset,s=>p(190)(116),cout=>p(191)(117));
FA_ff_4085:FAff port map(x=>p(93)(117),y=>p(94)(117),Cin=>p(95)(117),clock=>clock,reset=>reset,s=>p(190)(117),cout=>p(191)(118));
FA_ff_4086:FAff port map(x=>p(93)(118),y=>p(94)(118),Cin=>p(95)(118),clock=>clock,reset=>reset,s=>p(190)(118),cout=>p(191)(119));
FA_ff_4087:FAff port map(x=>p(93)(119),y=>p(94)(119),Cin=>p(95)(119),clock=>clock,reset=>reset,s=>p(190)(119),cout=>p(191)(120));
FA_ff_4088:FAff port map(x=>p(93)(120),y=>p(94)(120),Cin=>p(95)(120),clock=>clock,reset=>reset,s=>p(190)(120),cout=>p(191)(121));
FA_ff_4089:FAff port map(x=>p(93)(121),y=>p(94)(121),Cin=>p(95)(121),clock=>clock,reset=>reset,s=>p(190)(121),cout=>p(191)(122));
FA_ff_4090:FAff port map(x=>p(93)(122),y=>p(94)(122),Cin=>p(95)(122),clock=>clock,reset=>reset,s=>p(190)(122),cout=>p(191)(123));
FA_ff_4091:FAff port map(x=>p(93)(123),y=>p(94)(123),Cin=>p(95)(123),clock=>clock,reset=>reset,s=>p(190)(123),cout=>p(191)(124));
FA_ff_4092:FAff port map(x=>p(93)(124),y=>p(94)(124),Cin=>p(95)(124),clock=>clock,reset=>reset,s=>p(190)(124),cout=>p(191)(125));
FA_ff_4093:FAff port map(x=>p(93)(125),y=>p(94)(125),Cin=>p(95)(125),clock=>clock,reset=>reset,s=>p(190)(125),cout=>p(191)(126));
FA_ff_4094:FAff port map(x=>p(93)(126),y=>p(94)(126),Cin=>p(95)(126),clock=>clock,reset=>reset,s=>p(190)(126),cout=>p(191)(127));
FA_ff_4095:FAff port map(x=>p(93)(127),y=>p(94)(127),Cin=>p(95)(127),clock=>clock,reset=>reset,s=>p(190)(127),cout=>p(191)(128));
FA_ff_4096:FAff port map(x=>p(96)(0),y=>p(97)(0),Cin=>p(98)(0),clock=>clock,reset=>reset,s=>p(192)(0),cout=>p(193)(1));
FA_ff_4097:FAff port map(x=>p(96)(1),y=>p(97)(1),Cin=>p(98)(1),clock=>clock,reset=>reset,s=>p(192)(1),cout=>p(193)(2));
FA_ff_4098:FAff port map(x=>p(96)(2),y=>p(97)(2),Cin=>p(98)(2),clock=>clock,reset=>reset,s=>p(192)(2),cout=>p(193)(3));
FA_ff_4099:FAff port map(x=>p(96)(3),y=>p(97)(3),Cin=>p(98)(3),clock=>clock,reset=>reset,s=>p(192)(3),cout=>p(193)(4));
FA_ff_4100:FAff port map(x=>p(96)(4),y=>p(97)(4),Cin=>p(98)(4),clock=>clock,reset=>reset,s=>p(192)(4),cout=>p(193)(5));
FA_ff_4101:FAff port map(x=>p(96)(5),y=>p(97)(5),Cin=>p(98)(5),clock=>clock,reset=>reset,s=>p(192)(5),cout=>p(193)(6));
FA_ff_4102:FAff port map(x=>p(96)(6),y=>p(97)(6),Cin=>p(98)(6),clock=>clock,reset=>reset,s=>p(192)(6),cout=>p(193)(7));
FA_ff_4103:FAff port map(x=>p(96)(7),y=>p(97)(7),Cin=>p(98)(7),clock=>clock,reset=>reset,s=>p(192)(7),cout=>p(193)(8));
FA_ff_4104:FAff port map(x=>p(96)(8),y=>p(97)(8),Cin=>p(98)(8),clock=>clock,reset=>reset,s=>p(192)(8),cout=>p(193)(9));
FA_ff_4105:FAff port map(x=>p(96)(9),y=>p(97)(9),Cin=>p(98)(9),clock=>clock,reset=>reset,s=>p(192)(9),cout=>p(193)(10));
FA_ff_4106:FAff port map(x=>p(96)(10),y=>p(97)(10),Cin=>p(98)(10),clock=>clock,reset=>reset,s=>p(192)(10),cout=>p(193)(11));
FA_ff_4107:FAff port map(x=>p(96)(11),y=>p(97)(11),Cin=>p(98)(11),clock=>clock,reset=>reset,s=>p(192)(11),cout=>p(193)(12));
FA_ff_4108:FAff port map(x=>p(96)(12),y=>p(97)(12),Cin=>p(98)(12),clock=>clock,reset=>reset,s=>p(192)(12),cout=>p(193)(13));
FA_ff_4109:FAff port map(x=>p(96)(13),y=>p(97)(13),Cin=>p(98)(13),clock=>clock,reset=>reset,s=>p(192)(13),cout=>p(193)(14));
FA_ff_4110:FAff port map(x=>p(96)(14),y=>p(97)(14),Cin=>p(98)(14),clock=>clock,reset=>reset,s=>p(192)(14),cout=>p(193)(15));
FA_ff_4111:FAff port map(x=>p(96)(15),y=>p(97)(15),Cin=>p(98)(15),clock=>clock,reset=>reset,s=>p(192)(15),cout=>p(193)(16));
FA_ff_4112:FAff port map(x=>p(96)(16),y=>p(97)(16),Cin=>p(98)(16),clock=>clock,reset=>reset,s=>p(192)(16),cout=>p(193)(17));
FA_ff_4113:FAff port map(x=>p(96)(17),y=>p(97)(17),Cin=>p(98)(17),clock=>clock,reset=>reset,s=>p(192)(17),cout=>p(193)(18));
FA_ff_4114:FAff port map(x=>p(96)(18),y=>p(97)(18),Cin=>p(98)(18),clock=>clock,reset=>reset,s=>p(192)(18),cout=>p(193)(19));
FA_ff_4115:FAff port map(x=>p(96)(19),y=>p(97)(19),Cin=>p(98)(19),clock=>clock,reset=>reset,s=>p(192)(19),cout=>p(193)(20));
FA_ff_4116:FAff port map(x=>p(96)(20),y=>p(97)(20),Cin=>p(98)(20),clock=>clock,reset=>reset,s=>p(192)(20),cout=>p(193)(21));
FA_ff_4117:FAff port map(x=>p(96)(21),y=>p(97)(21),Cin=>p(98)(21),clock=>clock,reset=>reset,s=>p(192)(21),cout=>p(193)(22));
FA_ff_4118:FAff port map(x=>p(96)(22),y=>p(97)(22),Cin=>p(98)(22),clock=>clock,reset=>reset,s=>p(192)(22),cout=>p(193)(23));
FA_ff_4119:FAff port map(x=>p(96)(23),y=>p(97)(23),Cin=>p(98)(23),clock=>clock,reset=>reset,s=>p(192)(23),cout=>p(193)(24));
FA_ff_4120:FAff port map(x=>p(96)(24),y=>p(97)(24),Cin=>p(98)(24),clock=>clock,reset=>reset,s=>p(192)(24),cout=>p(193)(25));
FA_ff_4121:FAff port map(x=>p(96)(25),y=>p(97)(25),Cin=>p(98)(25),clock=>clock,reset=>reset,s=>p(192)(25),cout=>p(193)(26));
FA_ff_4122:FAff port map(x=>p(96)(26),y=>p(97)(26),Cin=>p(98)(26),clock=>clock,reset=>reset,s=>p(192)(26),cout=>p(193)(27));
FA_ff_4123:FAff port map(x=>p(96)(27),y=>p(97)(27),Cin=>p(98)(27),clock=>clock,reset=>reset,s=>p(192)(27),cout=>p(193)(28));
FA_ff_4124:FAff port map(x=>p(96)(28),y=>p(97)(28),Cin=>p(98)(28),clock=>clock,reset=>reset,s=>p(192)(28),cout=>p(193)(29));
FA_ff_4125:FAff port map(x=>p(96)(29),y=>p(97)(29),Cin=>p(98)(29),clock=>clock,reset=>reset,s=>p(192)(29),cout=>p(193)(30));
FA_ff_4126:FAff port map(x=>p(96)(30),y=>p(97)(30),Cin=>p(98)(30),clock=>clock,reset=>reset,s=>p(192)(30),cout=>p(193)(31));
FA_ff_4127:FAff port map(x=>p(96)(31),y=>p(97)(31),Cin=>p(98)(31),clock=>clock,reset=>reset,s=>p(192)(31),cout=>p(193)(32));
FA_ff_4128:FAff port map(x=>p(96)(32),y=>p(97)(32),Cin=>p(98)(32),clock=>clock,reset=>reset,s=>p(192)(32),cout=>p(193)(33));
FA_ff_4129:FAff port map(x=>p(96)(33),y=>p(97)(33),Cin=>p(98)(33),clock=>clock,reset=>reset,s=>p(192)(33),cout=>p(193)(34));
FA_ff_4130:FAff port map(x=>p(96)(34),y=>p(97)(34),Cin=>p(98)(34),clock=>clock,reset=>reset,s=>p(192)(34),cout=>p(193)(35));
FA_ff_4131:FAff port map(x=>p(96)(35),y=>p(97)(35),Cin=>p(98)(35),clock=>clock,reset=>reset,s=>p(192)(35),cout=>p(193)(36));
FA_ff_4132:FAff port map(x=>p(96)(36),y=>p(97)(36),Cin=>p(98)(36),clock=>clock,reset=>reset,s=>p(192)(36),cout=>p(193)(37));
FA_ff_4133:FAff port map(x=>p(96)(37),y=>p(97)(37),Cin=>p(98)(37),clock=>clock,reset=>reset,s=>p(192)(37),cout=>p(193)(38));
FA_ff_4134:FAff port map(x=>p(96)(38),y=>p(97)(38),Cin=>p(98)(38),clock=>clock,reset=>reset,s=>p(192)(38),cout=>p(193)(39));
FA_ff_4135:FAff port map(x=>p(96)(39),y=>p(97)(39),Cin=>p(98)(39),clock=>clock,reset=>reset,s=>p(192)(39),cout=>p(193)(40));
FA_ff_4136:FAff port map(x=>p(96)(40),y=>p(97)(40),Cin=>p(98)(40),clock=>clock,reset=>reset,s=>p(192)(40),cout=>p(193)(41));
FA_ff_4137:FAff port map(x=>p(96)(41),y=>p(97)(41),Cin=>p(98)(41),clock=>clock,reset=>reset,s=>p(192)(41),cout=>p(193)(42));
FA_ff_4138:FAff port map(x=>p(96)(42),y=>p(97)(42),Cin=>p(98)(42),clock=>clock,reset=>reset,s=>p(192)(42),cout=>p(193)(43));
FA_ff_4139:FAff port map(x=>p(96)(43),y=>p(97)(43),Cin=>p(98)(43),clock=>clock,reset=>reset,s=>p(192)(43),cout=>p(193)(44));
FA_ff_4140:FAff port map(x=>p(96)(44),y=>p(97)(44),Cin=>p(98)(44),clock=>clock,reset=>reset,s=>p(192)(44),cout=>p(193)(45));
FA_ff_4141:FAff port map(x=>p(96)(45),y=>p(97)(45),Cin=>p(98)(45),clock=>clock,reset=>reset,s=>p(192)(45),cout=>p(193)(46));
FA_ff_4142:FAff port map(x=>p(96)(46),y=>p(97)(46),Cin=>p(98)(46),clock=>clock,reset=>reset,s=>p(192)(46),cout=>p(193)(47));
FA_ff_4143:FAff port map(x=>p(96)(47),y=>p(97)(47),Cin=>p(98)(47),clock=>clock,reset=>reset,s=>p(192)(47),cout=>p(193)(48));
FA_ff_4144:FAff port map(x=>p(96)(48),y=>p(97)(48),Cin=>p(98)(48),clock=>clock,reset=>reset,s=>p(192)(48),cout=>p(193)(49));
FA_ff_4145:FAff port map(x=>p(96)(49),y=>p(97)(49),Cin=>p(98)(49),clock=>clock,reset=>reset,s=>p(192)(49),cout=>p(193)(50));
FA_ff_4146:FAff port map(x=>p(96)(50),y=>p(97)(50),Cin=>p(98)(50),clock=>clock,reset=>reset,s=>p(192)(50),cout=>p(193)(51));
FA_ff_4147:FAff port map(x=>p(96)(51),y=>p(97)(51),Cin=>p(98)(51),clock=>clock,reset=>reset,s=>p(192)(51),cout=>p(193)(52));
FA_ff_4148:FAff port map(x=>p(96)(52),y=>p(97)(52),Cin=>p(98)(52),clock=>clock,reset=>reset,s=>p(192)(52),cout=>p(193)(53));
FA_ff_4149:FAff port map(x=>p(96)(53),y=>p(97)(53),Cin=>p(98)(53),clock=>clock,reset=>reset,s=>p(192)(53),cout=>p(193)(54));
FA_ff_4150:FAff port map(x=>p(96)(54),y=>p(97)(54),Cin=>p(98)(54),clock=>clock,reset=>reset,s=>p(192)(54),cout=>p(193)(55));
FA_ff_4151:FAff port map(x=>p(96)(55),y=>p(97)(55),Cin=>p(98)(55),clock=>clock,reset=>reset,s=>p(192)(55),cout=>p(193)(56));
FA_ff_4152:FAff port map(x=>p(96)(56),y=>p(97)(56),Cin=>p(98)(56),clock=>clock,reset=>reset,s=>p(192)(56),cout=>p(193)(57));
FA_ff_4153:FAff port map(x=>p(96)(57),y=>p(97)(57),Cin=>p(98)(57),clock=>clock,reset=>reset,s=>p(192)(57),cout=>p(193)(58));
FA_ff_4154:FAff port map(x=>p(96)(58),y=>p(97)(58),Cin=>p(98)(58),clock=>clock,reset=>reset,s=>p(192)(58),cout=>p(193)(59));
FA_ff_4155:FAff port map(x=>p(96)(59),y=>p(97)(59),Cin=>p(98)(59),clock=>clock,reset=>reset,s=>p(192)(59),cout=>p(193)(60));
FA_ff_4156:FAff port map(x=>p(96)(60),y=>p(97)(60),Cin=>p(98)(60),clock=>clock,reset=>reset,s=>p(192)(60),cout=>p(193)(61));
FA_ff_4157:FAff port map(x=>p(96)(61),y=>p(97)(61),Cin=>p(98)(61),clock=>clock,reset=>reset,s=>p(192)(61),cout=>p(193)(62));
FA_ff_4158:FAff port map(x=>p(96)(62),y=>p(97)(62),Cin=>p(98)(62),clock=>clock,reset=>reset,s=>p(192)(62),cout=>p(193)(63));
FA_ff_4159:FAff port map(x=>p(96)(63),y=>p(97)(63),Cin=>p(98)(63),clock=>clock,reset=>reset,s=>p(192)(63),cout=>p(193)(64));
FA_ff_4160:FAff port map(x=>p(96)(64),y=>p(97)(64),Cin=>p(98)(64),clock=>clock,reset=>reset,s=>p(192)(64),cout=>p(193)(65));
FA_ff_4161:FAff port map(x=>p(96)(65),y=>p(97)(65),Cin=>p(98)(65),clock=>clock,reset=>reset,s=>p(192)(65),cout=>p(193)(66));
FA_ff_4162:FAff port map(x=>p(96)(66),y=>p(97)(66),Cin=>p(98)(66),clock=>clock,reset=>reset,s=>p(192)(66),cout=>p(193)(67));
FA_ff_4163:FAff port map(x=>p(96)(67),y=>p(97)(67),Cin=>p(98)(67),clock=>clock,reset=>reset,s=>p(192)(67),cout=>p(193)(68));
FA_ff_4164:FAff port map(x=>p(96)(68),y=>p(97)(68),Cin=>p(98)(68),clock=>clock,reset=>reset,s=>p(192)(68),cout=>p(193)(69));
FA_ff_4165:FAff port map(x=>p(96)(69),y=>p(97)(69),Cin=>p(98)(69),clock=>clock,reset=>reset,s=>p(192)(69),cout=>p(193)(70));
FA_ff_4166:FAff port map(x=>p(96)(70),y=>p(97)(70),Cin=>p(98)(70),clock=>clock,reset=>reset,s=>p(192)(70),cout=>p(193)(71));
FA_ff_4167:FAff port map(x=>p(96)(71),y=>p(97)(71),Cin=>p(98)(71),clock=>clock,reset=>reset,s=>p(192)(71),cout=>p(193)(72));
FA_ff_4168:FAff port map(x=>p(96)(72),y=>p(97)(72),Cin=>p(98)(72),clock=>clock,reset=>reset,s=>p(192)(72),cout=>p(193)(73));
FA_ff_4169:FAff port map(x=>p(96)(73),y=>p(97)(73),Cin=>p(98)(73),clock=>clock,reset=>reset,s=>p(192)(73),cout=>p(193)(74));
FA_ff_4170:FAff port map(x=>p(96)(74),y=>p(97)(74),Cin=>p(98)(74),clock=>clock,reset=>reset,s=>p(192)(74),cout=>p(193)(75));
FA_ff_4171:FAff port map(x=>p(96)(75),y=>p(97)(75),Cin=>p(98)(75),clock=>clock,reset=>reset,s=>p(192)(75),cout=>p(193)(76));
FA_ff_4172:FAff port map(x=>p(96)(76),y=>p(97)(76),Cin=>p(98)(76),clock=>clock,reset=>reset,s=>p(192)(76),cout=>p(193)(77));
FA_ff_4173:FAff port map(x=>p(96)(77),y=>p(97)(77),Cin=>p(98)(77),clock=>clock,reset=>reset,s=>p(192)(77),cout=>p(193)(78));
FA_ff_4174:FAff port map(x=>p(96)(78),y=>p(97)(78),Cin=>p(98)(78),clock=>clock,reset=>reset,s=>p(192)(78),cout=>p(193)(79));
FA_ff_4175:FAff port map(x=>p(96)(79),y=>p(97)(79),Cin=>p(98)(79),clock=>clock,reset=>reset,s=>p(192)(79),cout=>p(193)(80));
FA_ff_4176:FAff port map(x=>p(96)(80),y=>p(97)(80),Cin=>p(98)(80),clock=>clock,reset=>reset,s=>p(192)(80),cout=>p(193)(81));
FA_ff_4177:FAff port map(x=>p(96)(81),y=>p(97)(81),Cin=>p(98)(81),clock=>clock,reset=>reset,s=>p(192)(81),cout=>p(193)(82));
FA_ff_4178:FAff port map(x=>p(96)(82),y=>p(97)(82),Cin=>p(98)(82),clock=>clock,reset=>reset,s=>p(192)(82),cout=>p(193)(83));
FA_ff_4179:FAff port map(x=>p(96)(83),y=>p(97)(83),Cin=>p(98)(83),clock=>clock,reset=>reset,s=>p(192)(83),cout=>p(193)(84));
FA_ff_4180:FAff port map(x=>p(96)(84),y=>p(97)(84),Cin=>p(98)(84),clock=>clock,reset=>reset,s=>p(192)(84),cout=>p(193)(85));
FA_ff_4181:FAff port map(x=>p(96)(85),y=>p(97)(85),Cin=>p(98)(85),clock=>clock,reset=>reset,s=>p(192)(85),cout=>p(193)(86));
FA_ff_4182:FAff port map(x=>p(96)(86),y=>p(97)(86),Cin=>p(98)(86),clock=>clock,reset=>reset,s=>p(192)(86),cout=>p(193)(87));
FA_ff_4183:FAff port map(x=>p(96)(87),y=>p(97)(87),Cin=>p(98)(87),clock=>clock,reset=>reset,s=>p(192)(87),cout=>p(193)(88));
FA_ff_4184:FAff port map(x=>p(96)(88),y=>p(97)(88),Cin=>p(98)(88),clock=>clock,reset=>reset,s=>p(192)(88),cout=>p(193)(89));
FA_ff_4185:FAff port map(x=>p(96)(89),y=>p(97)(89),Cin=>p(98)(89),clock=>clock,reset=>reset,s=>p(192)(89),cout=>p(193)(90));
FA_ff_4186:FAff port map(x=>p(96)(90),y=>p(97)(90),Cin=>p(98)(90),clock=>clock,reset=>reset,s=>p(192)(90),cout=>p(193)(91));
FA_ff_4187:FAff port map(x=>p(96)(91),y=>p(97)(91),Cin=>p(98)(91),clock=>clock,reset=>reset,s=>p(192)(91),cout=>p(193)(92));
FA_ff_4188:FAff port map(x=>p(96)(92),y=>p(97)(92),Cin=>p(98)(92),clock=>clock,reset=>reset,s=>p(192)(92),cout=>p(193)(93));
FA_ff_4189:FAff port map(x=>p(96)(93),y=>p(97)(93),Cin=>p(98)(93),clock=>clock,reset=>reset,s=>p(192)(93),cout=>p(193)(94));
FA_ff_4190:FAff port map(x=>p(96)(94),y=>p(97)(94),Cin=>p(98)(94),clock=>clock,reset=>reset,s=>p(192)(94),cout=>p(193)(95));
FA_ff_4191:FAff port map(x=>p(96)(95),y=>p(97)(95),Cin=>p(98)(95),clock=>clock,reset=>reset,s=>p(192)(95),cout=>p(193)(96));
FA_ff_4192:FAff port map(x=>p(96)(96),y=>p(97)(96),Cin=>p(98)(96),clock=>clock,reset=>reset,s=>p(192)(96),cout=>p(193)(97));
FA_ff_4193:FAff port map(x=>p(96)(97),y=>p(97)(97),Cin=>p(98)(97),clock=>clock,reset=>reset,s=>p(192)(97),cout=>p(193)(98));
FA_ff_4194:FAff port map(x=>p(96)(98),y=>p(97)(98),Cin=>p(98)(98),clock=>clock,reset=>reset,s=>p(192)(98),cout=>p(193)(99));
FA_ff_4195:FAff port map(x=>p(96)(99),y=>p(97)(99),Cin=>p(98)(99),clock=>clock,reset=>reset,s=>p(192)(99),cout=>p(193)(100));
FA_ff_4196:FAff port map(x=>p(96)(100),y=>p(97)(100),Cin=>p(98)(100),clock=>clock,reset=>reset,s=>p(192)(100),cout=>p(193)(101));
FA_ff_4197:FAff port map(x=>p(96)(101),y=>p(97)(101),Cin=>p(98)(101),clock=>clock,reset=>reset,s=>p(192)(101),cout=>p(193)(102));
FA_ff_4198:FAff port map(x=>p(96)(102),y=>p(97)(102),Cin=>p(98)(102),clock=>clock,reset=>reset,s=>p(192)(102),cout=>p(193)(103));
FA_ff_4199:FAff port map(x=>p(96)(103),y=>p(97)(103),Cin=>p(98)(103),clock=>clock,reset=>reset,s=>p(192)(103),cout=>p(193)(104));
FA_ff_4200:FAff port map(x=>p(96)(104),y=>p(97)(104),Cin=>p(98)(104),clock=>clock,reset=>reset,s=>p(192)(104),cout=>p(193)(105));
FA_ff_4201:FAff port map(x=>p(96)(105),y=>p(97)(105),Cin=>p(98)(105),clock=>clock,reset=>reset,s=>p(192)(105),cout=>p(193)(106));
FA_ff_4202:FAff port map(x=>p(96)(106),y=>p(97)(106),Cin=>p(98)(106),clock=>clock,reset=>reset,s=>p(192)(106),cout=>p(193)(107));
FA_ff_4203:FAff port map(x=>p(96)(107),y=>p(97)(107),Cin=>p(98)(107),clock=>clock,reset=>reset,s=>p(192)(107),cout=>p(193)(108));
FA_ff_4204:FAff port map(x=>p(96)(108),y=>p(97)(108),Cin=>p(98)(108),clock=>clock,reset=>reset,s=>p(192)(108),cout=>p(193)(109));
FA_ff_4205:FAff port map(x=>p(96)(109),y=>p(97)(109),Cin=>p(98)(109),clock=>clock,reset=>reset,s=>p(192)(109),cout=>p(193)(110));
FA_ff_4206:FAff port map(x=>p(96)(110),y=>p(97)(110),Cin=>p(98)(110),clock=>clock,reset=>reset,s=>p(192)(110),cout=>p(193)(111));
FA_ff_4207:FAff port map(x=>p(96)(111),y=>p(97)(111),Cin=>p(98)(111),clock=>clock,reset=>reset,s=>p(192)(111),cout=>p(193)(112));
FA_ff_4208:FAff port map(x=>p(96)(112),y=>p(97)(112),Cin=>p(98)(112),clock=>clock,reset=>reset,s=>p(192)(112),cout=>p(193)(113));
FA_ff_4209:FAff port map(x=>p(96)(113),y=>p(97)(113),Cin=>p(98)(113),clock=>clock,reset=>reset,s=>p(192)(113),cout=>p(193)(114));
FA_ff_4210:FAff port map(x=>p(96)(114),y=>p(97)(114),Cin=>p(98)(114),clock=>clock,reset=>reset,s=>p(192)(114),cout=>p(193)(115));
FA_ff_4211:FAff port map(x=>p(96)(115),y=>p(97)(115),Cin=>p(98)(115),clock=>clock,reset=>reset,s=>p(192)(115),cout=>p(193)(116));
FA_ff_4212:FAff port map(x=>p(96)(116),y=>p(97)(116),Cin=>p(98)(116),clock=>clock,reset=>reset,s=>p(192)(116),cout=>p(193)(117));
FA_ff_4213:FAff port map(x=>p(96)(117),y=>p(97)(117),Cin=>p(98)(117),clock=>clock,reset=>reset,s=>p(192)(117),cout=>p(193)(118));
FA_ff_4214:FAff port map(x=>p(96)(118),y=>p(97)(118),Cin=>p(98)(118),clock=>clock,reset=>reset,s=>p(192)(118),cout=>p(193)(119));
FA_ff_4215:FAff port map(x=>p(96)(119),y=>p(97)(119),Cin=>p(98)(119),clock=>clock,reset=>reset,s=>p(192)(119),cout=>p(193)(120));
FA_ff_4216:FAff port map(x=>p(96)(120),y=>p(97)(120),Cin=>p(98)(120),clock=>clock,reset=>reset,s=>p(192)(120),cout=>p(193)(121));
FA_ff_4217:FAff port map(x=>p(96)(121),y=>p(97)(121),Cin=>p(98)(121),clock=>clock,reset=>reset,s=>p(192)(121),cout=>p(193)(122));
FA_ff_4218:FAff port map(x=>p(96)(122),y=>p(97)(122),Cin=>p(98)(122),clock=>clock,reset=>reset,s=>p(192)(122),cout=>p(193)(123));
FA_ff_4219:FAff port map(x=>p(96)(123),y=>p(97)(123),Cin=>p(98)(123),clock=>clock,reset=>reset,s=>p(192)(123),cout=>p(193)(124));
FA_ff_4220:FAff port map(x=>p(96)(124),y=>p(97)(124),Cin=>p(98)(124),clock=>clock,reset=>reset,s=>p(192)(124),cout=>p(193)(125));
FA_ff_4221:FAff port map(x=>p(96)(125),y=>p(97)(125),Cin=>p(98)(125),clock=>clock,reset=>reset,s=>p(192)(125),cout=>p(193)(126));
FA_ff_4222:FAff port map(x=>p(96)(126),y=>p(97)(126),Cin=>p(98)(126),clock=>clock,reset=>reset,s=>p(192)(126),cout=>p(193)(127));
FA_ff_4223:FAff port map(x=>p(96)(127),y=>p(97)(127),Cin=>p(98)(127),clock=>clock,reset=>reset,s=>p(192)(127),cout=>p(193)(128));
FA_ff_4224:FAff port map(x=>p(99)(0),y=>p(100)(0),Cin=>p(101)(0),clock=>clock,reset=>reset,s=>p(194)(0),cout=>p(195)(1));
FA_ff_4225:FAff port map(x=>p(99)(1),y=>p(100)(1),Cin=>p(101)(1),clock=>clock,reset=>reset,s=>p(194)(1),cout=>p(195)(2));
FA_ff_4226:FAff port map(x=>p(99)(2),y=>p(100)(2),Cin=>p(101)(2),clock=>clock,reset=>reset,s=>p(194)(2),cout=>p(195)(3));
FA_ff_4227:FAff port map(x=>p(99)(3),y=>p(100)(3),Cin=>p(101)(3),clock=>clock,reset=>reset,s=>p(194)(3),cout=>p(195)(4));
FA_ff_4228:FAff port map(x=>p(99)(4),y=>p(100)(4),Cin=>p(101)(4),clock=>clock,reset=>reset,s=>p(194)(4),cout=>p(195)(5));
FA_ff_4229:FAff port map(x=>p(99)(5),y=>p(100)(5),Cin=>p(101)(5),clock=>clock,reset=>reset,s=>p(194)(5),cout=>p(195)(6));
FA_ff_4230:FAff port map(x=>p(99)(6),y=>p(100)(6),Cin=>p(101)(6),clock=>clock,reset=>reset,s=>p(194)(6),cout=>p(195)(7));
FA_ff_4231:FAff port map(x=>p(99)(7),y=>p(100)(7),Cin=>p(101)(7),clock=>clock,reset=>reset,s=>p(194)(7),cout=>p(195)(8));
FA_ff_4232:FAff port map(x=>p(99)(8),y=>p(100)(8),Cin=>p(101)(8),clock=>clock,reset=>reset,s=>p(194)(8),cout=>p(195)(9));
FA_ff_4233:FAff port map(x=>p(99)(9),y=>p(100)(9),Cin=>p(101)(9),clock=>clock,reset=>reset,s=>p(194)(9),cout=>p(195)(10));
FA_ff_4234:FAff port map(x=>p(99)(10),y=>p(100)(10),Cin=>p(101)(10),clock=>clock,reset=>reset,s=>p(194)(10),cout=>p(195)(11));
FA_ff_4235:FAff port map(x=>p(99)(11),y=>p(100)(11),Cin=>p(101)(11),clock=>clock,reset=>reset,s=>p(194)(11),cout=>p(195)(12));
FA_ff_4236:FAff port map(x=>p(99)(12),y=>p(100)(12),Cin=>p(101)(12),clock=>clock,reset=>reset,s=>p(194)(12),cout=>p(195)(13));
FA_ff_4237:FAff port map(x=>p(99)(13),y=>p(100)(13),Cin=>p(101)(13),clock=>clock,reset=>reset,s=>p(194)(13),cout=>p(195)(14));
FA_ff_4238:FAff port map(x=>p(99)(14),y=>p(100)(14),Cin=>p(101)(14),clock=>clock,reset=>reset,s=>p(194)(14),cout=>p(195)(15));
FA_ff_4239:FAff port map(x=>p(99)(15),y=>p(100)(15),Cin=>p(101)(15),clock=>clock,reset=>reset,s=>p(194)(15),cout=>p(195)(16));
FA_ff_4240:FAff port map(x=>p(99)(16),y=>p(100)(16),Cin=>p(101)(16),clock=>clock,reset=>reset,s=>p(194)(16),cout=>p(195)(17));
FA_ff_4241:FAff port map(x=>p(99)(17),y=>p(100)(17),Cin=>p(101)(17),clock=>clock,reset=>reset,s=>p(194)(17),cout=>p(195)(18));
FA_ff_4242:FAff port map(x=>p(99)(18),y=>p(100)(18),Cin=>p(101)(18),clock=>clock,reset=>reset,s=>p(194)(18),cout=>p(195)(19));
FA_ff_4243:FAff port map(x=>p(99)(19),y=>p(100)(19),Cin=>p(101)(19),clock=>clock,reset=>reset,s=>p(194)(19),cout=>p(195)(20));
FA_ff_4244:FAff port map(x=>p(99)(20),y=>p(100)(20),Cin=>p(101)(20),clock=>clock,reset=>reset,s=>p(194)(20),cout=>p(195)(21));
FA_ff_4245:FAff port map(x=>p(99)(21),y=>p(100)(21),Cin=>p(101)(21),clock=>clock,reset=>reset,s=>p(194)(21),cout=>p(195)(22));
FA_ff_4246:FAff port map(x=>p(99)(22),y=>p(100)(22),Cin=>p(101)(22),clock=>clock,reset=>reset,s=>p(194)(22),cout=>p(195)(23));
FA_ff_4247:FAff port map(x=>p(99)(23),y=>p(100)(23),Cin=>p(101)(23),clock=>clock,reset=>reset,s=>p(194)(23),cout=>p(195)(24));
FA_ff_4248:FAff port map(x=>p(99)(24),y=>p(100)(24),Cin=>p(101)(24),clock=>clock,reset=>reset,s=>p(194)(24),cout=>p(195)(25));
FA_ff_4249:FAff port map(x=>p(99)(25),y=>p(100)(25),Cin=>p(101)(25),clock=>clock,reset=>reset,s=>p(194)(25),cout=>p(195)(26));
FA_ff_4250:FAff port map(x=>p(99)(26),y=>p(100)(26),Cin=>p(101)(26),clock=>clock,reset=>reset,s=>p(194)(26),cout=>p(195)(27));
FA_ff_4251:FAff port map(x=>p(99)(27),y=>p(100)(27),Cin=>p(101)(27),clock=>clock,reset=>reset,s=>p(194)(27),cout=>p(195)(28));
FA_ff_4252:FAff port map(x=>p(99)(28),y=>p(100)(28),Cin=>p(101)(28),clock=>clock,reset=>reset,s=>p(194)(28),cout=>p(195)(29));
FA_ff_4253:FAff port map(x=>p(99)(29),y=>p(100)(29),Cin=>p(101)(29),clock=>clock,reset=>reset,s=>p(194)(29),cout=>p(195)(30));
FA_ff_4254:FAff port map(x=>p(99)(30),y=>p(100)(30),Cin=>p(101)(30),clock=>clock,reset=>reset,s=>p(194)(30),cout=>p(195)(31));
FA_ff_4255:FAff port map(x=>p(99)(31),y=>p(100)(31),Cin=>p(101)(31),clock=>clock,reset=>reset,s=>p(194)(31),cout=>p(195)(32));
FA_ff_4256:FAff port map(x=>p(99)(32),y=>p(100)(32),Cin=>p(101)(32),clock=>clock,reset=>reset,s=>p(194)(32),cout=>p(195)(33));
FA_ff_4257:FAff port map(x=>p(99)(33),y=>p(100)(33),Cin=>p(101)(33),clock=>clock,reset=>reset,s=>p(194)(33),cout=>p(195)(34));
FA_ff_4258:FAff port map(x=>p(99)(34),y=>p(100)(34),Cin=>p(101)(34),clock=>clock,reset=>reset,s=>p(194)(34),cout=>p(195)(35));
FA_ff_4259:FAff port map(x=>p(99)(35),y=>p(100)(35),Cin=>p(101)(35),clock=>clock,reset=>reset,s=>p(194)(35),cout=>p(195)(36));
FA_ff_4260:FAff port map(x=>p(99)(36),y=>p(100)(36),Cin=>p(101)(36),clock=>clock,reset=>reset,s=>p(194)(36),cout=>p(195)(37));
FA_ff_4261:FAff port map(x=>p(99)(37),y=>p(100)(37),Cin=>p(101)(37),clock=>clock,reset=>reset,s=>p(194)(37),cout=>p(195)(38));
FA_ff_4262:FAff port map(x=>p(99)(38),y=>p(100)(38),Cin=>p(101)(38),clock=>clock,reset=>reset,s=>p(194)(38),cout=>p(195)(39));
FA_ff_4263:FAff port map(x=>p(99)(39),y=>p(100)(39),Cin=>p(101)(39),clock=>clock,reset=>reset,s=>p(194)(39),cout=>p(195)(40));
FA_ff_4264:FAff port map(x=>p(99)(40),y=>p(100)(40),Cin=>p(101)(40),clock=>clock,reset=>reset,s=>p(194)(40),cout=>p(195)(41));
FA_ff_4265:FAff port map(x=>p(99)(41),y=>p(100)(41),Cin=>p(101)(41),clock=>clock,reset=>reset,s=>p(194)(41),cout=>p(195)(42));
FA_ff_4266:FAff port map(x=>p(99)(42),y=>p(100)(42),Cin=>p(101)(42),clock=>clock,reset=>reset,s=>p(194)(42),cout=>p(195)(43));
FA_ff_4267:FAff port map(x=>p(99)(43),y=>p(100)(43),Cin=>p(101)(43),clock=>clock,reset=>reset,s=>p(194)(43),cout=>p(195)(44));
FA_ff_4268:FAff port map(x=>p(99)(44),y=>p(100)(44),Cin=>p(101)(44),clock=>clock,reset=>reset,s=>p(194)(44),cout=>p(195)(45));
FA_ff_4269:FAff port map(x=>p(99)(45),y=>p(100)(45),Cin=>p(101)(45),clock=>clock,reset=>reset,s=>p(194)(45),cout=>p(195)(46));
FA_ff_4270:FAff port map(x=>p(99)(46),y=>p(100)(46),Cin=>p(101)(46),clock=>clock,reset=>reset,s=>p(194)(46),cout=>p(195)(47));
FA_ff_4271:FAff port map(x=>p(99)(47),y=>p(100)(47),Cin=>p(101)(47),clock=>clock,reset=>reset,s=>p(194)(47),cout=>p(195)(48));
FA_ff_4272:FAff port map(x=>p(99)(48),y=>p(100)(48),Cin=>p(101)(48),clock=>clock,reset=>reset,s=>p(194)(48),cout=>p(195)(49));
FA_ff_4273:FAff port map(x=>p(99)(49),y=>p(100)(49),Cin=>p(101)(49),clock=>clock,reset=>reset,s=>p(194)(49),cout=>p(195)(50));
FA_ff_4274:FAff port map(x=>p(99)(50),y=>p(100)(50),Cin=>p(101)(50),clock=>clock,reset=>reset,s=>p(194)(50),cout=>p(195)(51));
FA_ff_4275:FAff port map(x=>p(99)(51),y=>p(100)(51),Cin=>p(101)(51),clock=>clock,reset=>reset,s=>p(194)(51),cout=>p(195)(52));
FA_ff_4276:FAff port map(x=>p(99)(52),y=>p(100)(52),Cin=>p(101)(52),clock=>clock,reset=>reset,s=>p(194)(52),cout=>p(195)(53));
FA_ff_4277:FAff port map(x=>p(99)(53),y=>p(100)(53),Cin=>p(101)(53),clock=>clock,reset=>reset,s=>p(194)(53),cout=>p(195)(54));
FA_ff_4278:FAff port map(x=>p(99)(54),y=>p(100)(54),Cin=>p(101)(54),clock=>clock,reset=>reset,s=>p(194)(54),cout=>p(195)(55));
FA_ff_4279:FAff port map(x=>p(99)(55),y=>p(100)(55),Cin=>p(101)(55),clock=>clock,reset=>reset,s=>p(194)(55),cout=>p(195)(56));
FA_ff_4280:FAff port map(x=>p(99)(56),y=>p(100)(56),Cin=>p(101)(56),clock=>clock,reset=>reset,s=>p(194)(56),cout=>p(195)(57));
FA_ff_4281:FAff port map(x=>p(99)(57),y=>p(100)(57),Cin=>p(101)(57),clock=>clock,reset=>reset,s=>p(194)(57),cout=>p(195)(58));
FA_ff_4282:FAff port map(x=>p(99)(58),y=>p(100)(58),Cin=>p(101)(58),clock=>clock,reset=>reset,s=>p(194)(58),cout=>p(195)(59));
FA_ff_4283:FAff port map(x=>p(99)(59),y=>p(100)(59),Cin=>p(101)(59),clock=>clock,reset=>reset,s=>p(194)(59),cout=>p(195)(60));
FA_ff_4284:FAff port map(x=>p(99)(60),y=>p(100)(60),Cin=>p(101)(60),clock=>clock,reset=>reset,s=>p(194)(60),cout=>p(195)(61));
FA_ff_4285:FAff port map(x=>p(99)(61),y=>p(100)(61),Cin=>p(101)(61),clock=>clock,reset=>reset,s=>p(194)(61),cout=>p(195)(62));
FA_ff_4286:FAff port map(x=>p(99)(62),y=>p(100)(62),Cin=>p(101)(62),clock=>clock,reset=>reset,s=>p(194)(62),cout=>p(195)(63));
FA_ff_4287:FAff port map(x=>p(99)(63),y=>p(100)(63),Cin=>p(101)(63),clock=>clock,reset=>reset,s=>p(194)(63),cout=>p(195)(64));
FA_ff_4288:FAff port map(x=>p(99)(64),y=>p(100)(64),Cin=>p(101)(64),clock=>clock,reset=>reset,s=>p(194)(64),cout=>p(195)(65));
FA_ff_4289:FAff port map(x=>p(99)(65),y=>p(100)(65),Cin=>p(101)(65),clock=>clock,reset=>reset,s=>p(194)(65),cout=>p(195)(66));
FA_ff_4290:FAff port map(x=>p(99)(66),y=>p(100)(66),Cin=>p(101)(66),clock=>clock,reset=>reset,s=>p(194)(66),cout=>p(195)(67));
FA_ff_4291:FAff port map(x=>p(99)(67),y=>p(100)(67),Cin=>p(101)(67),clock=>clock,reset=>reset,s=>p(194)(67),cout=>p(195)(68));
FA_ff_4292:FAff port map(x=>p(99)(68),y=>p(100)(68),Cin=>p(101)(68),clock=>clock,reset=>reset,s=>p(194)(68),cout=>p(195)(69));
FA_ff_4293:FAff port map(x=>p(99)(69),y=>p(100)(69),Cin=>p(101)(69),clock=>clock,reset=>reset,s=>p(194)(69),cout=>p(195)(70));
FA_ff_4294:FAff port map(x=>p(99)(70),y=>p(100)(70),Cin=>p(101)(70),clock=>clock,reset=>reset,s=>p(194)(70),cout=>p(195)(71));
FA_ff_4295:FAff port map(x=>p(99)(71),y=>p(100)(71),Cin=>p(101)(71),clock=>clock,reset=>reset,s=>p(194)(71),cout=>p(195)(72));
FA_ff_4296:FAff port map(x=>p(99)(72),y=>p(100)(72),Cin=>p(101)(72),clock=>clock,reset=>reset,s=>p(194)(72),cout=>p(195)(73));
FA_ff_4297:FAff port map(x=>p(99)(73),y=>p(100)(73),Cin=>p(101)(73),clock=>clock,reset=>reset,s=>p(194)(73),cout=>p(195)(74));
FA_ff_4298:FAff port map(x=>p(99)(74),y=>p(100)(74),Cin=>p(101)(74),clock=>clock,reset=>reset,s=>p(194)(74),cout=>p(195)(75));
FA_ff_4299:FAff port map(x=>p(99)(75),y=>p(100)(75),Cin=>p(101)(75),clock=>clock,reset=>reset,s=>p(194)(75),cout=>p(195)(76));
FA_ff_4300:FAff port map(x=>p(99)(76),y=>p(100)(76),Cin=>p(101)(76),clock=>clock,reset=>reset,s=>p(194)(76),cout=>p(195)(77));
FA_ff_4301:FAff port map(x=>p(99)(77),y=>p(100)(77),Cin=>p(101)(77),clock=>clock,reset=>reset,s=>p(194)(77),cout=>p(195)(78));
FA_ff_4302:FAff port map(x=>p(99)(78),y=>p(100)(78),Cin=>p(101)(78),clock=>clock,reset=>reset,s=>p(194)(78),cout=>p(195)(79));
FA_ff_4303:FAff port map(x=>p(99)(79),y=>p(100)(79),Cin=>p(101)(79),clock=>clock,reset=>reset,s=>p(194)(79),cout=>p(195)(80));
FA_ff_4304:FAff port map(x=>p(99)(80),y=>p(100)(80),Cin=>p(101)(80),clock=>clock,reset=>reset,s=>p(194)(80),cout=>p(195)(81));
FA_ff_4305:FAff port map(x=>p(99)(81),y=>p(100)(81),Cin=>p(101)(81),clock=>clock,reset=>reset,s=>p(194)(81),cout=>p(195)(82));
FA_ff_4306:FAff port map(x=>p(99)(82),y=>p(100)(82),Cin=>p(101)(82),clock=>clock,reset=>reset,s=>p(194)(82),cout=>p(195)(83));
FA_ff_4307:FAff port map(x=>p(99)(83),y=>p(100)(83),Cin=>p(101)(83),clock=>clock,reset=>reset,s=>p(194)(83),cout=>p(195)(84));
FA_ff_4308:FAff port map(x=>p(99)(84),y=>p(100)(84),Cin=>p(101)(84),clock=>clock,reset=>reset,s=>p(194)(84),cout=>p(195)(85));
FA_ff_4309:FAff port map(x=>p(99)(85),y=>p(100)(85),Cin=>p(101)(85),clock=>clock,reset=>reset,s=>p(194)(85),cout=>p(195)(86));
FA_ff_4310:FAff port map(x=>p(99)(86),y=>p(100)(86),Cin=>p(101)(86),clock=>clock,reset=>reset,s=>p(194)(86),cout=>p(195)(87));
FA_ff_4311:FAff port map(x=>p(99)(87),y=>p(100)(87),Cin=>p(101)(87),clock=>clock,reset=>reset,s=>p(194)(87),cout=>p(195)(88));
FA_ff_4312:FAff port map(x=>p(99)(88),y=>p(100)(88),Cin=>p(101)(88),clock=>clock,reset=>reset,s=>p(194)(88),cout=>p(195)(89));
FA_ff_4313:FAff port map(x=>p(99)(89),y=>p(100)(89),Cin=>p(101)(89),clock=>clock,reset=>reset,s=>p(194)(89),cout=>p(195)(90));
FA_ff_4314:FAff port map(x=>p(99)(90),y=>p(100)(90),Cin=>p(101)(90),clock=>clock,reset=>reset,s=>p(194)(90),cout=>p(195)(91));
FA_ff_4315:FAff port map(x=>p(99)(91),y=>p(100)(91),Cin=>p(101)(91),clock=>clock,reset=>reset,s=>p(194)(91),cout=>p(195)(92));
FA_ff_4316:FAff port map(x=>p(99)(92),y=>p(100)(92),Cin=>p(101)(92),clock=>clock,reset=>reset,s=>p(194)(92),cout=>p(195)(93));
FA_ff_4317:FAff port map(x=>p(99)(93),y=>p(100)(93),Cin=>p(101)(93),clock=>clock,reset=>reset,s=>p(194)(93),cout=>p(195)(94));
FA_ff_4318:FAff port map(x=>p(99)(94),y=>p(100)(94),Cin=>p(101)(94),clock=>clock,reset=>reset,s=>p(194)(94),cout=>p(195)(95));
FA_ff_4319:FAff port map(x=>p(99)(95),y=>p(100)(95),Cin=>p(101)(95),clock=>clock,reset=>reset,s=>p(194)(95),cout=>p(195)(96));
FA_ff_4320:FAff port map(x=>p(99)(96),y=>p(100)(96),Cin=>p(101)(96),clock=>clock,reset=>reset,s=>p(194)(96),cout=>p(195)(97));
FA_ff_4321:FAff port map(x=>p(99)(97),y=>p(100)(97),Cin=>p(101)(97),clock=>clock,reset=>reset,s=>p(194)(97),cout=>p(195)(98));
FA_ff_4322:FAff port map(x=>p(99)(98),y=>p(100)(98),Cin=>p(101)(98),clock=>clock,reset=>reset,s=>p(194)(98),cout=>p(195)(99));
FA_ff_4323:FAff port map(x=>p(99)(99),y=>p(100)(99),Cin=>p(101)(99),clock=>clock,reset=>reset,s=>p(194)(99),cout=>p(195)(100));
FA_ff_4324:FAff port map(x=>p(99)(100),y=>p(100)(100),Cin=>p(101)(100),clock=>clock,reset=>reset,s=>p(194)(100),cout=>p(195)(101));
FA_ff_4325:FAff port map(x=>p(99)(101),y=>p(100)(101),Cin=>p(101)(101),clock=>clock,reset=>reset,s=>p(194)(101),cout=>p(195)(102));
FA_ff_4326:FAff port map(x=>p(99)(102),y=>p(100)(102),Cin=>p(101)(102),clock=>clock,reset=>reset,s=>p(194)(102),cout=>p(195)(103));
FA_ff_4327:FAff port map(x=>p(99)(103),y=>p(100)(103),Cin=>p(101)(103),clock=>clock,reset=>reset,s=>p(194)(103),cout=>p(195)(104));
FA_ff_4328:FAff port map(x=>p(99)(104),y=>p(100)(104),Cin=>p(101)(104),clock=>clock,reset=>reset,s=>p(194)(104),cout=>p(195)(105));
FA_ff_4329:FAff port map(x=>p(99)(105),y=>p(100)(105),Cin=>p(101)(105),clock=>clock,reset=>reset,s=>p(194)(105),cout=>p(195)(106));
FA_ff_4330:FAff port map(x=>p(99)(106),y=>p(100)(106),Cin=>p(101)(106),clock=>clock,reset=>reset,s=>p(194)(106),cout=>p(195)(107));
FA_ff_4331:FAff port map(x=>p(99)(107),y=>p(100)(107),Cin=>p(101)(107),clock=>clock,reset=>reset,s=>p(194)(107),cout=>p(195)(108));
FA_ff_4332:FAff port map(x=>p(99)(108),y=>p(100)(108),Cin=>p(101)(108),clock=>clock,reset=>reset,s=>p(194)(108),cout=>p(195)(109));
FA_ff_4333:FAff port map(x=>p(99)(109),y=>p(100)(109),Cin=>p(101)(109),clock=>clock,reset=>reset,s=>p(194)(109),cout=>p(195)(110));
FA_ff_4334:FAff port map(x=>p(99)(110),y=>p(100)(110),Cin=>p(101)(110),clock=>clock,reset=>reset,s=>p(194)(110),cout=>p(195)(111));
FA_ff_4335:FAff port map(x=>p(99)(111),y=>p(100)(111),Cin=>p(101)(111),clock=>clock,reset=>reset,s=>p(194)(111),cout=>p(195)(112));
FA_ff_4336:FAff port map(x=>p(99)(112),y=>p(100)(112),Cin=>p(101)(112),clock=>clock,reset=>reset,s=>p(194)(112),cout=>p(195)(113));
FA_ff_4337:FAff port map(x=>p(99)(113),y=>p(100)(113),Cin=>p(101)(113),clock=>clock,reset=>reset,s=>p(194)(113),cout=>p(195)(114));
FA_ff_4338:FAff port map(x=>p(99)(114),y=>p(100)(114),Cin=>p(101)(114),clock=>clock,reset=>reset,s=>p(194)(114),cout=>p(195)(115));
FA_ff_4339:FAff port map(x=>p(99)(115),y=>p(100)(115),Cin=>p(101)(115),clock=>clock,reset=>reset,s=>p(194)(115),cout=>p(195)(116));
FA_ff_4340:FAff port map(x=>p(99)(116),y=>p(100)(116),Cin=>p(101)(116),clock=>clock,reset=>reset,s=>p(194)(116),cout=>p(195)(117));
FA_ff_4341:FAff port map(x=>p(99)(117),y=>p(100)(117),Cin=>p(101)(117),clock=>clock,reset=>reset,s=>p(194)(117),cout=>p(195)(118));
FA_ff_4342:FAff port map(x=>p(99)(118),y=>p(100)(118),Cin=>p(101)(118),clock=>clock,reset=>reset,s=>p(194)(118),cout=>p(195)(119));
FA_ff_4343:FAff port map(x=>p(99)(119),y=>p(100)(119),Cin=>p(101)(119),clock=>clock,reset=>reset,s=>p(194)(119),cout=>p(195)(120));
FA_ff_4344:FAff port map(x=>p(99)(120),y=>p(100)(120),Cin=>p(101)(120),clock=>clock,reset=>reset,s=>p(194)(120),cout=>p(195)(121));
FA_ff_4345:FAff port map(x=>p(99)(121),y=>p(100)(121),Cin=>p(101)(121),clock=>clock,reset=>reset,s=>p(194)(121),cout=>p(195)(122));
FA_ff_4346:FAff port map(x=>p(99)(122),y=>p(100)(122),Cin=>p(101)(122),clock=>clock,reset=>reset,s=>p(194)(122),cout=>p(195)(123));
FA_ff_4347:FAff port map(x=>p(99)(123),y=>p(100)(123),Cin=>p(101)(123),clock=>clock,reset=>reset,s=>p(194)(123),cout=>p(195)(124));
FA_ff_4348:FAff port map(x=>p(99)(124),y=>p(100)(124),Cin=>p(101)(124),clock=>clock,reset=>reset,s=>p(194)(124),cout=>p(195)(125));
FA_ff_4349:FAff port map(x=>p(99)(125),y=>p(100)(125),Cin=>p(101)(125),clock=>clock,reset=>reset,s=>p(194)(125),cout=>p(195)(126));
FA_ff_4350:FAff port map(x=>p(99)(126),y=>p(100)(126),Cin=>p(101)(126),clock=>clock,reset=>reset,s=>p(194)(126),cout=>p(195)(127));
FA_ff_4351:FAff port map(x=>p(99)(127),y=>p(100)(127),Cin=>p(101)(127),clock=>clock,reset=>reset,s=>p(194)(127),cout=>p(195)(128));
FA_ff_4352:FAff port map(x=>p(102)(0),y=>p(103)(0),Cin=>p(104)(0),clock=>clock,reset=>reset,s=>p(196)(0),cout=>p(197)(1));
FA_ff_4353:FAff port map(x=>p(102)(1),y=>p(103)(1),Cin=>p(104)(1),clock=>clock,reset=>reset,s=>p(196)(1),cout=>p(197)(2));
FA_ff_4354:FAff port map(x=>p(102)(2),y=>p(103)(2),Cin=>p(104)(2),clock=>clock,reset=>reset,s=>p(196)(2),cout=>p(197)(3));
FA_ff_4355:FAff port map(x=>p(102)(3),y=>p(103)(3),Cin=>p(104)(3),clock=>clock,reset=>reset,s=>p(196)(3),cout=>p(197)(4));
FA_ff_4356:FAff port map(x=>p(102)(4),y=>p(103)(4),Cin=>p(104)(4),clock=>clock,reset=>reset,s=>p(196)(4),cout=>p(197)(5));
FA_ff_4357:FAff port map(x=>p(102)(5),y=>p(103)(5),Cin=>p(104)(5),clock=>clock,reset=>reset,s=>p(196)(5),cout=>p(197)(6));
FA_ff_4358:FAff port map(x=>p(102)(6),y=>p(103)(6),Cin=>p(104)(6),clock=>clock,reset=>reset,s=>p(196)(6),cout=>p(197)(7));
FA_ff_4359:FAff port map(x=>p(102)(7),y=>p(103)(7),Cin=>p(104)(7),clock=>clock,reset=>reset,s=>p(196)(7),cout=>p(197)(8));
FA_ff_4360:FAff port map(x=>p(102)(8),y=>p(103)(8),Cin=>p(104)(8),clock=>clock,reset=>reset,s=>p(196)(8),cout=>p(197)(9));
FA_ff_4361:FAff port map(x=>p(102)(9),y=>p(103)(9),Cin=>p(104)(9),clock=>clock,reset=>reset,s=>p(196)(9),cout=>p(197)(10));
FA_ff_4362:FAff port map(x=>p(102)(10),y=>p(103)(10),Cin=>p(104)(10),clock=>clock,reset=>reset,s=>p(196)(10),cout=>p(197)(11));
FA_ff_4363:FAff port map(x=>p(102)(11),y=>p(103)(11),Cin=>p(104)(11),clock=>clock,reset=>reset,s=>p(196)(11),cout=>p(197)(12));
FA_ff_4364:FAff port map(x=>p(102)(12),y=>p(103)(12),Cin=>p(104)(12),clock=>clock,reset=>reset,s=>p(196)(12),cout=>p(197)(13));
FA_ff_4365:FAff port map(x=>p(102)(13),y=>p(103)(13),Cin=>p(104)(13),clock=>clock,reset=>reset,s=>p(196)(13),cout=>p(197)(14));
FA_ff_4366:FAff port map(x=>p(102)(14),y=>p(103)(14),Cin=>p(104)(14),clock=>clock,reset=>reset,s=>p(196)(14),cout=>p(197)(15));
FA_ff_4367:FAff port map(x=>p(102)(15),y=>p(103)(15),Cin=>p(104)(15),clock=>clock,reset=>reset,s=>p(196)(15),cout=>p(197)(16));
FA_ff_4368:FAff port map(x=>p(102)(16),y=>p(103)(16),Cin=>p(104)(16),clock=>clock,reset=>reset,s=>p(196)(16),cout=>p(197)(17));
FA_ff_4369:FAff port map(x=>p(102)(17),y=>p(103)(17),Cin=>p(104)(17),clock=>clock,reset=>reset,s=>p(196)(17),cout=>p(197)(18));
FA_ff_4370:FAff port map(x=>p(102)(18),y=>p(103)(18),Cin=>p(104)(18),clock=>clock,reset=>reset,s=>p(196)(18),cout=>p(197)(19));
FA_ff_4371:FAff port map(x=>p(102)(19),y=>p(103)(19),Cin=>p(104)(19),clock=>clock,reset=>reset,s=>p(196)(19),cout=>p(197)(20));
FA_ff_4372:FAff port map(x=>p(102)(20),y=>p(103)(20),Cin=>p(104)(20),clock=>clock,reset=>reset,s=>p(196)(20),cout=>p(197)(21));
FA_ff_4373:FAff port map(x=>p(102)(21),y=>p(103)(21),Cin=>p(104)(21),clock=>clock,reset=>reset,s=>p(196)(21),cout=>p(197)(22));
FA_ff_4374:FAff port map(x=>p(102)(22),y=>p(103)(22),Cin=>p(104)(22),clock=>clock,reset=>reset,s=>p(196)(22),cout=>p(197)(23));
FA_ff_4375:FAff port map(x=>p(102)(23),y=>p(103)(23),Cin=>p(104)(23),clock=>clock,reset=>reset,s=>p(196)(23),cout=>p(197)(24));
FA_ff_4376:FAff port map(x=>p(102)(24),y=>p(103)(24),Cin=>p(104)(24),clock=>clock,reset=>reset,s=>p(196)(24),cout=>p(197)(25));
FA_ff_4377:FAff port map(x=>p(102)(25),y=>p(103)(25),Cin=>p(104)(25),clock=>clock,reset=>reset,s=>p(196)(25),cout=>p(197)(26));
FA_ff_4378:FAff port map(x=>p(102)(26),y=>p(103)(26),Cin=>p(104)(26),clock=>clock,reset=>reset,s=>p(196)(26),cout=>p(197)(27));
FA_ff_4379:FAff port map(x=>p(102)(27),y=>p(103)(27),Cin=>p(104)(27),clock=>clock,reset=>reset,s=>p(196)(27),cout=>p(197)(28));
FA_ff_4380:FAff port map(x=>p(102)(28),y=>p(103)(28),Cin=>p(104)(28),clock=>clock,reset=>reset,s=>p(196)(28),cout=>p(197)(29));
FA_ff_4381:FAff port map(x=>p(102)(29),y=>p(103)(29),Cin=>p(104)(29),clock=>clock,reset=>reset,s=>p(196)(29),cout=>p(197)(30));
FA_ff_4382:FAff port map(x=>p(102)(30),y=>p(103)(30),Cin=>p(104)(30),clock=>clock,reset=>reset,s=>p(196)(30),cout=>p(197)(31));
FA_ff_4383:FAff port map(x=>p(102)(31),y=>p(103)(31),Cin=>p(104)(31),clock=>clock,reset=>reset,s=>p(196)(31),cout=>p(197)(32));
FA_ff_4384:FAff port map(x=>p(102)(32),y=>p(103)(32),Cin=>p(104)(32),clock=>clock,reset=>reset,s=>p(196)(32),cout=>p(197)(33));
FA_ff_4385:FAff port map(x=>p(102)(33),y=>p(103)(33),Cin=>p(104)(33),clock=>clock,reset=>reset,s=>p(196)(33),cout=>p(197)(34));
FA_ff_4386:FAff port map(x=>p(102)(34),y=>p(103)(34),Cin=>p(104)(34),clock=>clock,reset=>reset,s=>p(196)(34),cout=>p(197)(35));
FA_ff_4387:FAff port map(x=>p(102)(35),y=>p(103)(35),Cin=>p(104)(35),clock=>clock,reset=>reset,s=>p(196)(35),cout=>p(197)(36));
FA_ff_4388:FAff port map(x=>p(102)(36),y=>p(103)(36),Cin=>p(104)(36),clock=>clock,reset=>reset,s=>p(196)(36),cout=>p(197)(37));
FA_ff_4389:FAff port map(x=>p(102)(37),y=>p(103)(37),Cin=>p(104)(37),clock=>clock,reset=>reset,s=>p(196)(37),cout=>p(197)(38));
FA_ff_4390:FAff port map(x=>p(102)(38),y=>p(103)(38),Cin=>p(104)(38),clock=>clock,reset=>reset,s=>p(196)(38),cout=>p(197)(39));
FA_ff_4391:FAff port map(x=>p(102)(39),y=>p(103)(39),Cin=>p(104)(39),clock=>clock,reset=>reset,s=>p(196)(39),cout=>p(197)(40));
FA_ff_4392:FAff port map(x=>p(102)(40),y=>p(103)(40),Cin=>p(104)(40),clock=>clock,reset=>reset,s=>p(196)(40),cout=>p(197)(41));
FA_ff_4393:FAff port map(x=>p(102)(41),y=>p(103)(41),Cin=>p(104)(41),clock=>clock,reset=>reset,s=>p(196)(41),cout=>p(197)(42));
FA_ff_4394:FAff port map(x=>p(102)(42),y=>p(103)(42),Cin=>p(104)(42),clock=>clock,reset=>reset,s=>p(196)(42),cout=>p(197)(43));
FA_ff_4395:FAff port map(x=>p(102)(43),y=>p(103)(43),Cin=>p(104)(43),clock=>clock,reset=>reset,s=>p(196)(43),cout=>p(197)(44));
FA_ff_4396:FAff port map(x=>p(102)(44),y=>p(103)(44),Cin=>p(104)(44),clock=>clock,reset=>reset,s=>p(196)(44),cout=>p(197)(45));
FA_ff_4397:FAff port map(x=>p(102)(45),y=>p(103)(45),Cin=>p(104)(45),clock=>clock,reset=>reset,s=>p(196)(45),cout=>p(197)(46));
FA_ff_4398:FAff port map(x=>p(102)(46),y=>p(103)(46),Cin=>p(104)(46),clock=>clock,reset=>reset,s=>p(196)(46),cout=>p(197)(47));
FA_ff_4399:FAff port map(x=>p(102)(47),y=>p(103)(47),Cin=>p(104)(47),clock=>clock,reset=>reset,s=>p(196)(47),cout=>p(197)(48));
FA_ff_4400:FAff port map(x=>p(102)(48),y=>p(103)(48),Cin=>p(104)(48),clock=>clock,reset=>reset,s=>p(196)(48),cout=>p(197)(49));
FA_ff_4401:FAff port map(x=>p(102)(49),y=>p(103)(49),Cin=>p(104)(49),clock=>clock,reset=>reset,s=>p(196)(49),cout=>p(197)(50));
FA_ff_4402:FAff port map(x=>p(102)(50),y=>p(103)(50),Cin=>p(104)(50),clock=>clock,reset=>reset,s=>p(196)(50),cout=>p(197)(51));
FA_ff_4403:FAff port map(x=>p(102)(51),y=>p(103)(51),Cin=>p(104)(51),clock=>clock,reset=>reset,s=>p(196)(51),cout=>p(197)(52));
FA_ff_4404:FAff port map(x=>p(102)(52),y=>p(103)(52),Cin=>p(104)(52),clock=>clock,reset=>reset,s=>p(196)(52),cout=>p(197)(53));
FA_ff_4405:FAff port map(x=>p(102)(53),y=>p(103)(53),Cin=>p(104)(53),clock=>clock,reset=>reset,s=>p(196)(53),cout=>p(197)(54));
FA_ff_4406:FAff port map(x=>p(102)(54),y=>p(103)(54),Cin=>p(104)(54),clock=>clock,reset=>reset,s=>p(196)(54),cout=>p(197)(55));
FA_ff_4407:FAff port map(x=>p(102)(55),y=>p(103)(55),Cin=>p(104)(55),clock=>clock,reset=>reset,s=>p(196)(55),cout=>p(197)(56));
FA_ff_4408:FAff port map(x=>p(102)(56),y=>p(103)(56),Cin=>p(104)(56),clock=>clock,reset=>reset,s=>p(196)(56),cout=>p(197)(57));
FA_ff_4409:FAff port map(x=>p(102)(57),y=>p(103)(57),Cin=>p(104)(57),clock=>clock,reset=>reset,s=>p(196)(57),cout=>p(197)(58));
FA_ff_4410:FAff port map(x=>p(102)(58),y=>p(103)(58),Cin=>p(104)(58),clock=>clock,reset=>reset,s=>p(196)(58),cout=>p(197)(59));
FA_ff_4411:FAff port map(x=>p(102)(59),y=>p(103)(59),Cin=>p(104)(59),clock=>clock,reset=>reset,s=>p(196)(59),cout=>p(197)(60));
FA_ff_4412:FAff port map(x=>p(102)(60),y=>p(103)(60),Cin=>p(104)(60),clock=>clock,reset=>reset,s=>p(196)(60),cout=>p(197)(61));
FA_ff_4413:FAff port map(x=>p(102)(61),y=>p(103)(61),Cin=>p(104)(61),clock=>clock,reset=>reset,s=>p(196)(61),cout=>p(197)(62));
FA_ff_4414:FAff port map(x=>p(102)(62),y=>p(103)(62),Cin=>p(104)(62),clock=>clock,reset=>reset,s=>p(196)(62),cout=>p(197)(63));
FA_ff_4415:FAff port map(x=>p(102)(63),y=>p(103)(63),Cin=>p(104)(63),clock=>clock,reset=>reset,s=>p(196)(63),cout=>p(197)(64));
FA_ff_4416:FAff port map(x=>p(102)(64),y=>p(103)(64),Cin=>p(104)(64),clock=>clock,reset=>reset,s=>p(196)(64),cout=>p(197)(65));
FA_ff_4417:FAff port map(x=>p(102)(65),y=>p(103)(65),Cin=>p(104)(65),clock=>clock,reset=>reset,s=>p(196)(65),cout=>p(197)(66));
FA_ff_4418:FAff port map(x=>p(102)(66),y=>p(103)(66),Cin=>p(104)(66),clock=>clock,reset=>reset,s=>p(196)(66),cout=>p(197)(67));
FA_ff_4419:FAff port map(x=>p(102)(67),y=>p(103)(67),Cin=>p(104)(67),clock=>clock,reset=>reset,s=>p(196)(67),cout=>p(197)(68));
FA_ff_4420:FAff port map(x=>p(102)(68),y=>p(103)(68),Cin=>p(104)(68),clock=>clock,reset=>reset,s=>p(196)(68),cout=>p(197)(69));
FA_ff_4421:FAff port map(x=>p(102)(69),y=>p(103)(69),Cin=>p(104)(69),clock=>clock,reset=>reset,s=>p(196)(69),cout=>p(197)(70));
FA_ff_4422:FAff port map(x=>p(102)(70),y=>p(103)(70),Cin=>p(104)(70),clock=>clock,reset=>reset,s=>p(196)(70),cout=>p(197)(71));
FA_ff_4423:FAff port map(x=>p(102)(71),y=>p(103)(71),Cin=>p(104)(71),clock=>clock,reset=>reset,s=>p(196)(71),cout=>p(197)(72));
FA_ff_4424:FAff port map(x=>p(102)(72),y=>p(103)(72),Cin=>p(104)(72),clock=>clock,reset=>reset,s=>p(196)(72),cout=>p(197)(73));
FA_ff_4425:FAff port map(x=>p(102)(73),y=>p(103)(73),Cin=>p(104)(73),clock=>clock,reset=>reset,s=>p(196)(73),cout=>p(197)(74));
FA_ff_4426:FAff port map(x=>p(102)(74),y=>p(103)(74),Cin=>p(104)(74),clock=>clock,reset=>reset,s=>p(196)(74),cout=>p(197)(75));
FA_ff_4427:FAff port map(x=>p(102)(75),y=>p(103)(75),Cin=>p(104)(75),clock=>clock,reset=>reset,s=>p(196)(75),cout=>p(197)(76));
FA_ff_4428:FAff port map(x=>p(102)(76),y=>p(103)(76),Cin=>p(104)(76),clock=>clock,reset=>reset,s=>p(196)(76),cout=>p(197)(77));
FA_ff_4429:FAff port map(x=>p(102)(77),y=>p(103)(77),Cin=>p(104)(77),clock=>clock,reset=>reset,s=>p(196)(77),cout=>p(197)(78));
FA_ff_4430:FAff port map(x=>p(102)(78),y=>p(103)(78),Cin=>p(104)(78),clock=>clock,reset=>reset,s=>p(196)(78),cout=>p(197)(79));
FA_ff_4431:FAff port map(x=>p(102)(79),y=>p(103)(79),Cin=>p(104)(79),clock=>clock,reset=>reset,s=>p(196)(79),cout=>p(197)(80));
FA_ff_4432:FAff port map(x=>p(102)(80),y=>p(103)(80),Cin=>p(104)(80),clock=>clock,reset=>reset,s=>p(196)(80),cout=>p(197)(81));
FA_ff_4433:FAff port map(x=>p(102)(81),y=>p(103)(81),Cin=>p(104)(81),clock=>clock,reset=>reset,s=>p(196)(81),cout=>p(197)(82));
FA_ff_4434:FAff port map(x=>p(102)(82),y=>p(103)(82),Cin=>p(104)(82),clock=>clock,reset=>reset,s=>p(196)(82),cout=>p(197)(83));
FA_ff_4435:FAff port map(x=>p(102)(83),y=>p(103)(83),Cin=>p(104)(83),clock=>clock,reset=>reset,s=>p(196)(83),cout=>p(197)(84));
FA_ff_4436:FAff port map(x=>p(102)(84),y=>p(103)(84),Cin=>p(104)(84),clock=>clock,reset=>reset,s=>p(196)(84),cout=>p(197)(85));
FA_ff_4437:FAff port map(x=>p(102)(85),y=>p(103)(85),Cin=>p(104)(85),clock=>clock,reset=>reset,s=>p(196)(85),cout=>p(197)(86));
FA_ff_4438:FAff port map(x=>p(102)(86),y=>p(103)(86),Cin=>p(104)(86),clock=>clock,reset=>reset,s=>p(196)(86),cout=>p(197)(87));
FA_ff_4439:FAff port map(x=>p(102)(87),y=>p(103)(87),Cin=>p(104)(87),clock=>clock,reset=>reset,s=>p(196)(87),cout=>p(197)(88));
FA_ff_4440:FAff port map(x=>p(102)(88),y=>p(103)(88),Cin=>p(104)(88),clock=>clock,reset=>reset,s=>p(196)(88),cout=>p(197)(89));
FA_ff_4441:FAff port map(x=>p(102)(89),y=>p(103)(89),Cin=>p(104)(89),clock=>clock,reset=>reset,s=>p(196)(89),cout=>p(197)(90));
FA_ff_4442:FAff port map(x=>p(102)(90),y=>p(103)(90),Cin=>p(104)(90),clock=>clock,reset=>reset,s=>p(196)(90),cout=>p(197)(91));
FA_ff_4443:FAff port map(x=>p(102)(91),y=>p(103)(91),Cin=>p(104)(91),clock=>clock,reset=>reset,s=>p(196)(91),cout=>p(197)(92));
FA_ff_4444:FAff port map(x=>p(102)(92),y=>p(103)(92),Cin=>p(104)(92),clock=>clock,reset=>reset,s=>p(196)(92),cout=>p(197)(93));
FA_ff_4445:FAff port map(x=>p(102)(93),y=>p(103)(93),Cin=>p(104)(93),clock=>clock,reset=>reset,s=>p(196)(93),cout=>p(197)(94));
FA_ff_4446:FAff port map(x=>p(102)(94),y=>p(103)(94),Cin=>p(104)(94),clock=>clock,reset=>reset,s=>p(196)(94),cout=>p(197)(95));
FA_ff_4447:FAff port map(x=>p(102)(95),y=>p(103)(95),Cin=>p(104)(95),clock=>clock,reset=>reset,s=>p(196)(95),cout=>p(197)(96));
FA_ff_4448:FAff port map(x=>p(102)(96),y=>p(103)(96),Cin=>p(104)(96),clock=>clock,reset=>reset,s=>p(196)(96),cout=>p(197)(97));
FA_ff_4449:FAff port map(x=>p(102)(97),y=>p(103)(97),Cin=>p(104)(97),clock=>clock,reset=>reset,s=>p(196)(97),cout=>p(197)(98));
FA_ff_4450:FAff port map(x=>p(102)(98),y=>p(103)(98),Cin=>p(104)(98),clock=>clock,reset=>reset,s=>p(196)(98),cout=>p(197)(99));
FA_ff_4451:FAff port map(x=>p(102)(99),y=>p(103)(99),Cin=>p(104)(99),clock=>clock,reset=>reset,s=>p(196)(99),cout=>p(197)(100));
FA_ff_4452:FAff port map(x=>p(102)(100),y=>p(103)(100),Cin=>p(104)(100),clock=>clock,reset=>reset,s=>p(196)(100),cout=>p(197)(101));
FA_ff_4453:FAff port map(x=>p(102)(101),y=>p(103)(101),Cin=>p(104)(101),clock=>clock,reset=>reset,s=>p(196)(101),cout=>p(197)(102));
FA_ff_4454:FAff port map(x=>p(102)(102),y=>p(103)(102),Cin=>p(104)(102),clock=>clock,reset=>reset,s=>p(196)(102),cout=>p(197)(103));
FA_ff_4455:FAff port map(x=>p(102)(103),y=>p(103)(103),Cin=>p(104)(103),clock=>clock,reset=>reset,s=>p(196)(103),cout=>p(197)(104));
FA_ff_4456:FAff port map(x=>p(102)(104),y=>p(103)(104),Cin=>p(104)(104),clock=>clock,reset=>reset,s=>p(196)(104),cout=>p(197)(105));
FA_ff_4457:FAff port map(x=>p(102)(105),y=>p(103)(105),Cin=>p(104)(105),clock=>clock,reset=>reset,s=>p(196)(105),cout=>p(197)(106));
FA_ff_4458:FAff port map(x=>p(102)(106),y=>p(103)(106),Cin=>p(104)(106),clock=>clock,reset=>reset,s=>p(196)(106),cout=>p(197)(107));
FA_ff_4459:FAff port map(x=>p(102)(107),y=>p(103)(107),Cin=>p(104)(107),clock=>clock,reset=>reset,s=>p(196)(107),cout=>p(197)(108));
FA_ff_4460:FAff port map(x=>p(102)(108),y=>p(103)(108),Cin=>p(104)(108),clock=>clock,reset=>reset,s=>p(196)(108),cout=>p(197)(109));
FA_ff_4461:FAff port map(x=>p(102)(109),y=>p(103)(109),Cin=>p(104)(109),clock=>clock,reset=>reset,s=>p(196)(109),cout=>p(197)(110));
FA_ff_4462:FAff port map(x=>p(102)(110),y=>p(103)(110),Cin=>p(104)(110),clock=>clock,reset=>reset,s=>p(196)(110),cout=>p(197)(111));
FA_ff_4463:FAff port map(x=>p(102)(111),y=>p(103)(111),Cin=>p(104)(111),clock=>clock,reset=>reset,s=>p(196)(111),cout=>p(197)(112));
FA_ff_4464:FAff port map(x=>p(102)(112),y=>p(103)(112),Cin=>p(104)(112),clock=>clock,reset=>reset,s=>p(196)(112),cout=>p(197)(113));
FA_ff_4465:FAff port map(x=>p(102)(113),y=>p(103)(113),Cin=>p(104)(113),clock=>clock,reset=>reset,s=>p(196)(113),cout=>p(197)(114));
FA_ff_4466:FAff port map(x=>p(102)(114),y=>p(103)(114),Cin=>p(104)(114),clock=>clock,reset=>reset,s=>p(196)(114),cout=>p(197)(115));
FA_ff_4467:FAff port map(x=>p(102)(115),y=>p(103)(115),Cin=>p(104)(115),clock=>clock,reset=>reset,s=>p(196)(115),cout=>p(197)(116));
FA_ff_4468:FAff port map(x=>p(102)(116),y=>p(103)(116),Cin=>p(104)(116),clock=>clock,reset=>reset,s=>p(196)(116),cout=>p(197)(117));
FA_ff_4469:FAff port map(x=>p(102)(117),y=>p(103)(117),Cin=>p(104)(117),clock=>clock,reset=>reset,s=>p(196)(117),cout=>p(197)(118));
FA_ff_4470:FAff port map(x=>p(102)(118),y=>p(103)(118),Cin=>p(104)(118),clock=>clock,reset=>reset,s=>p(196)(118),cout=>p(197)(119));
FA_ff_4471:FAff port map(x=>p(102)(119),y=>p(103)(119),Cin=>p(104)(119),clock=>clock,reset=>reset,s=>p(196)(119),cout=>p(197)(120));
FA_ff_4472:FAff port map(x=>p(102)(120),y=>p(103)(120),Cin=>p(104)(120),clock=>clock,reset=>reset,s=>p(196)(120),cout=>p(197)(121));
FA_ff_4473:FAff port map(x=>p(102)(121),y=>p(103)(121),Cin=>p(104)(121),clock=>clock,reset=>reset,s=>p(196)(121),cout=>p(197)(122));
FA_ff_4474:FAff port map(x=>p(102)(122),y=>p(103)(122),Cin=>p(104)(122),clock=>clock,reset=>reset,s=>p(196)(122),cout=>p(197)(123));
FA_ff_4475:FAff port map(x=>p(102)(123),y=>p(103)(123),Cin=>p(104)(123),clock=>clock,reset=>reset,s=>p(196)(123),cout=>p(197)(124));
FA_ff_4476:FAff port map(x=>p(102)(124),y=>p(103)(124),Cin=>p(104)(124),clock=>clock,reset=>reset,s=>p(196)(124),cout=>p(197)(125));
FA_ff_4477:FAff port map(x=>p(102)(125),y=>p(103)(125),Cin=>p(104)(125),clock=>clock,reset=>reset,s=>p(196)(125),cout=>p(197)(126));
FA_ff_4478:FAff port map(x=>p(102)(126),y=>p(103)(126),Cin=>p(104)(126),clock=>clock,reset=>reset,s=>p(196)(126),cout=>p(197)(127));
FA_ff_4479:FAff port map(x=>p(102)(127),y=>p(103)(127),Cin=>p(104)(127),clock=>clock,reset=>reset,s=>p(196)(127),cout=>p(197)(128));
FA_ff_4480:FAff port map(x=>p(105)(0),y=>p(106)(0),Cin=>p(107)(0),clock=>clock,reset=>reset,s=>p(198)(0),cout=>p(199)(1));
FA_ff_4481:FAff port map(x=>p(105)(1),y=>p(106)(1),Cin=>p(107)(1),clock=>clock,reset=>reset,s=>p(198)(1),cout=>p(199)(2));
FA_ff_4482:FAff port map(x=>p(105)(2),y=>p(106)(2),Cin=>p(107)(2),clock=>clock,reset=>reset,s=>p(198)(2),cout=>p(199)(3));
FA_ff_4483:FAff port map(x=>p(105)(3),y=>p(106)(3),Cin=>p(107)(3),clock=>clock,reset=>reset,s=>p(198)(3),cout=>p(199)(4));
FA_ff_4484:FAff port map(x=>p(105)(4),y=>p(106)(4),Cin=>p(107)(4),clock=>clock,reset=>reset,s=>p(198)(4),cout=>p(199)(5));
FA_ff_4485:FAff port map(x=>p(105)(5),y=>p(106)(5),Cin=>p(107)(5),clock=>clock,reset=>reset,s=>p(198)(5),cout=>p(199)(6));
FA_ff_4486:FAff port map(x=>p(105)(6),y=>p(106)(6),Cin=>p(107)(6),clock=>clock,reset=>reset,s=>p(198)(6),cout=>p(199)(7));
FA_ff_4487:FAff port map(x=>p(105)(7),y=>p(106)(7),Cin=>p(107)(7),clock=>clock,reset=>reset,s=>p(198)(7),cout=>p(199)(8));
FA_ff_4488:FAff port map(x=>p(105)(8),y=>p(106)(8),Cin=>p(107)(8),clock=>clock,reset=>reset,s=>p(198)(8),cout=>p(199)(9));
FA_ff_4489:FAff port map(x=>p(105)(9),y=>p(106)(9),Cin=>p(107)(9),clock=>clock,reset=>reset,s=>p(198)(9),cout=>p(199)(10));
FA_ff_4490:FAff port map(x=>p(105)(10),y=>p(106)(10),Cin=>p(107)(10),clock=>clock,reset=>reset,s=>p(198)(10),cout=>p(199)(11));
FA_ff_4491:FAff port map(x=>p(105)(11),y=>p(106)(11),Cin=>p(107)(11),clock=>clock,reset=>reset,s=>p(198)(11),cout=>p(199)(12));
FA_ff_4492:FAff port map(x=>p(105)(12),y=>p(106)(12),Cin=>p(107)(12),clock=>clock,reset=>reset,s=>p(198)(12),cout=>p(199)(13));
FA_ff_4493:FAff port map(x=>p(105)(13),y=>p(106)(13),Cin=>p(107)(13),clock=>clock,reset=>reset,s=>p(198)(13),cout=>p(199)(14));
FA_ff_4494:FAff port map(x=>p(105)(14),y=>p(106)(14),Cin=>p(107)(14),clock=>clock,reset=>reset,s=>p(198)(14),cout=>p(199)(15));
FA_ff_4495:FAff port map(x=>p(105)(15),y=>p(106)(15),Cin=>p(107)(15),clock=>clock,reset=>reset,s=>p(198)(15),cout=>p(199)(16));
FA_ff_4496:FAff port map(x=>p(105)(16),y=>p(106)(16),Cin=>p(107)(16),clock=>clock,reset=>reset,s=>p(198)(16),cout=>p(199)(17));
FA_ff_4497:FAff port map(x=>p(105)(17),y=>p(106)(17),Cin=>p(107)(17),clock=>clock,reset=>reset,s=>p(198)(17),cout=>p(199)(18));
FA_ff_4498:FAff port map(x=>p(105)(18),y=>p(106)(18),Cin=>p(107)(18),clock=>clock,reset=>reset,s=>p(198)(18),cout=>p(199)(19));
FA_ff_4499:FAff port map(x=>p(105)(19),y=>p(106)(19),Cin=>p(107)(19),clock=>clock,reset=>reset,s=>p(198)(19),cout=>p(199)(20));
FA_ff_4500:FAff port map(x=>p(105)(20),y=>p(106)(20),Cin=>p(107)(20),clock=>clock,reset=>reset,s=>p(198)(20),cout=>p(199)(21));
FA_ff_4501:FAff port map(x=>p(105)(21),y=>p(106)(21),Cin=>p(107)(21),clock=>clock,reset=>reset,s=>p(198)(21),cout=>p(199)(22));
FA_ff_4502:FAff port map(x=>p(105)(22),y=>p(106)(22),Cin=>p(107)(22),clock=>clock,reset=>reset,s=>p(198)(22),cout=>p(199)(23));
FA_ff_4503:FAff port map(x=>p(105)(23),y=>p(106)(23),Cin=>p(107)(23),clock=>clock,reset=>reset,s=>p(198)(23),cout=>p(199)(24));
FA_ff_4504:FAff port map(x=>p(105)(24),y=>p(106)(24),Cin=>p(107)(24),clock=>clock,reset=>reset,s=>p(198)(24),cout=>p(199)(25));
FA_ff_4505:FAff port map(x=>p(105)(25),y=>p(106)(25),Cin=>p(107)(25),clock=>clock,reset=>reset,s=>p(198)(25),cout=>p(199)(26));
FA_ff_4506:FAff port map(x=>p(105)(26),y=>p(106)(26),Cin=>p(107)(26),clock=>clock,reset=>reset,s=>p(198)(26),cout=>p(199)(27));
FA_ff_4507:FAff port map(x=>p(105)(27),y=>p(106)(27),Cin=>p(107)(27),clock=>clock,reset=>reset,s=>p(198)(27),cout=>p(199)(28));
FA_ff_4508:FAff port map(x=>p(105)(28),y=>p(106)(28),Cin=>p(107)(28),clock=>clock,reset=>reset,s=>p(198)(28),cout=>p(199)(29));
FA_ff_4509:FAff port map(x=>p(105)(29),y=>p(106)(29),Cin=>p(107)(29),clock=>clock,reset=>reset,s=>p(198)(29),cout=>p(199)(30));
FA_ff_4510:FAff port map(x=>p(105)(30),y=>p(106)(30),Cin=>p(107)(30),clock=>clock,reset=>reset,s=>p(198)(30),cout=>p(199)(31));
FA_ff_4511:FAff port map(x=>p(105)(31),y=>p(106)(31),Cin=>p(107)(31),clock=>clock,reset=>reset,s=>p(198)(31),cout=>p(199)(32));
FA_ff_4512:FAff port map(x=>p(105)(32),y=>p(106)(32),Cin=>p(107)(32),clock=>clock,reset=>reset,s=>p(198)(32),cout=>p(199)(33));
FA_ff_4513:FAff port map(x=>p(105)(33),y=>p(106)(33),Cin=>p(107)(33),clock=>clock,reset=>reset,s=>p(198)(33),cout=>p(199)(34));
FA_ff_4514:FAff port map(x=>p(105)(34),y=>p(106)(34),Cin=>p(107)(34),clock=>clock,reset=>reset,s=>p(198)(34),cout=>p(199)(35));
FA_ff_4515:FAff port map(x=>p(105)(35),y=>p(106)(35),Cin=>p(107)(35),clock=>clock,reset=>reset,s=>p(198)(35),cout=>p(199)(36));
FA_ff_4516:FAff port map(x=>p(105)(36),y=>p(106)(36),Cin=>p(107)(36),clock=>clock,reset=>reset,s=>p(198)(36),cout=>p(199)(37));
FA_ff_4517:FAff port map(x=>p(105)(37),y=>p(106)(37),Cin=>p(107)(37),clock=>clock,reset=>reset,s=>p(198)(37),cout=>p(199)(38));
FA_ff_4518:FAff port map(x=>p(105)(38),y=>p(106)(38),Cin=>p(107)(38),clock=>clock,reset=>reset,s=>p(198)(38),cout=>p(199)(39));
FA_ff_4519:FAff port map(x=>p(105)(39),y=>p(106)(39),Cin=>p(107)(39),clock=>clock,reset=>reset,s=>p(198)(39),cout=>p(199)(40));
FA_ff_4520:FAff port map(x=>p(105)(40),y=>p(106)(40),Cin=>p(107)(40),clock=>clock,reset=>reset,s=>p(198)(40),cout=>p(199)(41));
FA_ff_4521:FAff port map(x=>p(105)(41),y=>p(106)(41),Cin=>p(107)(41),clock=>clock,reset=>reset,s=>p(198)(41),cout=>p(199)(42));
FA_ff_4522:FAff port map(x=>p(105)(42),y=>p(106)(42),Cin=>p(107)(42),clock=>clock,reset=>reset,s=>p(198)(42),cout=>p(199)(43));
FA_ff_4523:FAff port map(x=>p(105)(43),y=>p(106)(43),Cin=>p(107)(43),clock=>clock,reset=>reset,s=>p(198)(43),cout=>p(199)(44));
FA_ff_4524:FAff port map(x=>p(105)(44),y=>p(106)(44),Cin=>p(107)(44),clock=>clock,reset=>reset,s=>p(198)(44),cout=>p(199)(45));
FA_ff_4525:FAff port map(x=>p(105)(45),y=>p(106)(45),Cin=>p(107)(45),clock=>clock,reset=>reset,s=>p(198)(45),cout=>p(199)(46));
FA_ff_4526:FAff port map(x=>p(105)(46),y=>p(106)(46),Cin=>p(107)(46),clock=>clock,reset=>reset,s=>p(198)(46),cout=>p(199)(47));
FA_ff_4527:FAff port map(x=>p(105)(47),y=>p(106)(47),Cin=>p(107)(47),clock=>clock,reset=>reset,s=>p(198)(47),cout=>p(199)(48));
FA_ff_4528:FAff port map(x=>p(105)(48),y=>p(106)(48),Cin=>p(107)(48),clock=>clock,reset=>reset,s=>p(198)(48),cout=>p(199)(49));
FA_ff_4529:FAff port map(x=>p(105)(49),y=>p(106)(49),Cin=>p(107)(49),clock=>clock,reset=>reset,s=>p(198)(49),cout=>p(199)(50));
FA_ff_4530:FAff port map(x=>p(105)(50),y=>p(106)(50),Cin=>p(107)(50),clock=>clock,reset=>reset,s=>p(198)(50),cout=>p(199)(51));
FA_ff_4531:FAff port map(x=>p(105)(51),y=>p(106)(51),Cin=>p(107)(51),clock=>clock,reset=>reset,s=>p(198)(51),cout=>p(199)(52));
FA_ff_4532:FAff port map(x=>p(105)(52),y=>p(106)(52),Cin=>p(107)(52),clock=>clock,reset=>reset,s=>p(198)(52),cout=>p(199)(53));
FA_ff_4533:FAff port map(x=>p(105)(53),y=>p(106)(53),Cin=>p(107)(53),clock=>clock,reset=>reset,s=>p(198)(53),cout=>p(199)(54));
FA_ff_4534:FAff port map(x=>p(105)(54),y=>p(106)(54),Cin=>p(107)(54),clock=>clock,reset=>reset,s=>p(198)(54),cout=>p(199)(55));
FA_ff_4535:FAff port map(x=>p(105)(55),y=>p(106)(55),Cin=>p(107)(55),clock=>clock,reset=>reset,s=>p(198)(55),cout=>p(199)(56));
FA_ff_4536:FAff port map(x=>p(105)(56),y=>p(106)(56),Cin=>p(107)(56),clock=>clock,reset=>reset,s=>p(198)(56),cout=>p(199)(57));
FA_ff_4537:FAff port map(x=>p(105)(57),y=>p(106)(57),Cin=>p(107)(57),clock=>clock,reset=>reset,s=>p(198)(57),cout=>p(199)(58));
FA_ff_4538:FAff port map(x=>p(105)(58),y=>p(106)(58),Cin=>p(107)(58),clock=>clock,reset=>reset,s=>p(198)(58),cout=>p(199)(59));
FA_ff_4539:FAff port map(x=>p(105)(59),y=>p(106)(59),Cin=>p(107)(59),clock=>clock,reset=>reset,s=>p(198)(59),cout=>p(199)(60));
FA_ff_4540:FAff port map(x=>p(105)(60),y=>p(106)(60),Cin=>p(107)(60),clock=>clock,reset=>reset,s=>p(198)(60),cout=>p(199)(61));
FA_ff_4541:FAff port map(x=>p(105)(61),y=>p(106)(61),Cin=>p(107)(61),clock=>clock,reset=>reset,s=>p(198)(61),cout=>p(199)(62));
FA_ff_4542:FAff port map(x=>p(105)(62),y=>p(106)(62),Cin=>p(107)(62),clock=>clock,reset=>reset,s=>p(198)(62),cout=>p(199)(63));
FA_ff_4543:FAff port map(x=>p(105)(63),y=>p(106)(63),Cin=>p(107)(63),clock=>clock,reset=>reset,s=>p(198)(63),cout=>p(199)(64));
FA_ff_4544:FAff port map(x=>p(105)(64),y=>p(106)(64),Cin=>p(107)(64),clock=>clock,reset=>reset,s=>p(198)(64),cout=>p(199)(65));
FA_ff_4545:FAff port map(x=>p(105)(65),y=>p(106)(65),Cin=>p(107)(65),clock=>clock,reset=>reset,s=>p(198)(65),cout=>p(199)(66));
FA_ff_4546:FAff port map(x=>p(105)(66),y=>p(106)(66),Cin=>p(107)(66),clock=>clock,reset=>reset,s=>p(198)(66),cout=>p(199)(67));
FA_ff_4547:FAff port map(x=>p(105)(67),y=>p(106)(67),Cin=>p(107)(67),clock=>clock,reset=>reset,s=>p(198)(67),cout=>p(199)(68));
FA_ff_4548:FAff port map(x=>p(105)(68),y=>p(106)(68),Cin=>p(107)(68),clock=>clock,reset=>reset,s=>p(198)(68),cout=>p(199)(69));
FA_ff_4549:FAff port map(x=>p(105)(69),y=>p(106)(69),Cin=>p(107)(69),clock=>clock,reset=>reset,s=>p(198)(69),cout=>p(199)(70));
FA_ff_4550:FAff port map(x=>p(105)(70),y=>p(106)(70),Cin=>p(107)(70),clock=>clock,reset=>reset,s=>p(198)(70),cout=>p(199)(71));
FA_ff_4551:FAff port map(x=>p(105)(71),y=>p(106)(71),Cin=>p(107)(71),clock=>clock,reset=>reset,s=>p(198)(71),cout=>p(199)(72));
FA_ff_4552:FAff port map(x=>p(105)(72),y=>p(106)(72),Cin=>p(107)(72),clock=>clock,reset=>reset,s=>p(198)(72),cout=>p(199)(73));
FA_ff_4553:FAff port map(x=>p(105)(73),y=>p(106)(73),Cin=>p(107)(73),clock=>clock,reset=>reset,s=>p(198)(73),cout=>p(199)(74));
FA_ff_4554:FAff port map(x=>p(105)(74),y=>p(106)(74),Cin=>p(107)(74),clock=>clock,reset=>reset,s=>p(198)(74),cout=>p(199)(75));
FA_ff_4555:FAff port map(x=>p(105)(75),y=>p(106)(75),Cin=>p(107)(75),clock=>clock,reset=>reset,s=>p(198)(75),cout=>p(199)(76));
FA_ff_4556:FAff port map(x=>p(105)(76),y=>p(106)(76),Cin=>p(107)(76),clock=>clock,reset=>reset,s=>p(198)(76),cout=>p(199)(77));
FA_ff_4557:FAff port map(x=>p(105)(77),y=>p(106)(77),Cin=>p(107)(77),clock=>clock,reset=>reset,s=>p(198)(77),cout=>p(199)(78));
FA_ff_4558:FAff port map(x=>p(105)(78),y=>p(106)(78),Cin=>p(107)(78),clock=>clock,reset=>reset,s=>p(198)(78),cout=>p(199)(79));
FA_ff_4559:FAff port map(x=>p(105)(79),y=>p(106)(79),Cin=>p(107)(79),clock=>clock,reset=>reset,s=>p(198)(79),cout=>p(199)(80));
FA_ff_4560:FAff port map(x=>p(105)(80),y=>p(106)(80),Cin=>p(107)(80),clock=>clock,reset=>reset,s=>p(198)(80),cout=>p(199)(81));
FA_ff_4561:FAff port map(x=>p(105)(81),y=>p(106)(81),Cin=>p(107)(81),clock=>clock,reset=>reset,s=>p(198)(81),cout=>p(199)(82));
FA_ff_4562:FAff port map(x=>p(105)(82),y=>p(106)(82),Cin=>p(107)(82),clock=>clock,reset=>reset,s=>p(198)(82),cout=>p(199)(83));
FA_ff_4563:FAff port map(x=>p(105)(83),y=>p(106)(83),Cin=>p(107)(83),clock=>clock,reset=>reset,s=>p(198)(83),cout=>p(199)(84));
FA_ff_4564:FAff port map(x=>p(105)(84),y=>p(106)(84),Cin=>p(107)(84),clock=>clock,reset=>reset,s=>p(198)(84),cout=>p(199)(85));
FA_ff_4565:FAff port map(x=>p(105)(85),y=>p(106)(85),Cin=>p(107)(85),clock=>clock,reset=>reset,s=>p(198)(85),cout=>p(199)(86));
FA_ff_4566:FAff port map(x=>p(105)(86),y=>p(106)(86),Cin=>p(107)(86),clock=>clock,reset=>reset,s=>p(198)(86),cout=>p(199)(87));
FA_ff_4567:FAff port map(x=>p(105)(87),y=>p(106)(87),Cin=>p(107)(87),clock=>clock,reset=>reset,s=>p(198)(87),cout=>p(199)(88));
FA_ff_4568:FAff port map(x=>p(105)(88),y=>p(106)(88),Cin=>p(107)(88),clock=>clock,reset=>reset,s=>p(198)(88),cout=>p(199)(89));
FA_ff_4569:FAff port map(x=>p(105)(89),y=>p(106)(89),Cin=>p(107)(89),clock=>clock,reset=>reset,s=>p(198)(89),cout=>p(199)(90));
FA_ff_4570:FAff port map(x=>p(105)(90),y=>p(106)(90),Cin=>p(107)(90),clock=>clock,reset=>reset,s=>p(198)(90),cout=>p(199)(91));
FA_ff_4571:FAff port map(x=>p(105)(91),y=>p(106)(91),Cin=>p(107)(91),clock=>clock,reset=>reset,s=>p(198)(91),cout=>p(199)(92));
FA_ff_4572:FAff port map(x=>p(105)(92),y=>p(106)(92),Cin=>p(107)(92),clock=>clock,reset=>reset,s=>p(198)(92),cout=>p(199)(93));
FA_ff_4573:FAff port map(x=>p(105)(93),y=>p(106)(93),Cin=>p(107)(93),clock=>clock,reset=>reset,s=>p(198)(93),cout=>p(199)(94));
FA_ff_4574:FAff port map(x=>p(105)(94),y=>p(106)(94),Cin=>p(107)(94),clock=>clock,reset=>reset,s=>p(198)(94),cout=>p(199)(95));
FA_ff_4575:FAff port map(x=>p(105)(95),y=>p(106)(95),Cin=>p(107)(95),clock=>clock,reset=>reset,s=>p(198)(95),cout=>p(199)(96));
FA_ff_4576:FAff port map(x=>p(105)(96),y=>p(106)(96),Cin=>p(107)(96),clock=>clock,reset=>reset,s=>p(198)(96),cout=>p(199)(97));
FA_ff_4577:FAff port map(x=>p(105)(97),y=>p(106)(97),Cin=>p(107)(97),clock=>clock,reset=>reset,s=>p(198)(97),cout=>p(199)(98));
FA_ff_4578:FAff port map(x=>p(105)(98),y=>p(106)(98),Cin=>p(107)(98),clock=>clock,reset=>reset,s=>p(198)(98),cout=>p(199)(99));
FA_ff_4579:FAff port map(x=>p(105)(99),y=>p(106)(99),Cin=>p(107)(99),clock=>clock,reset=>reset,s=>p(198)(99),cout=>p(199)(100));
FA_ff_4580:FAff port map(x=>p(105)(100),y=>p(106)(100),Cin=>p(107)(100),clock=>clock,reset=>reset,s=>p(198)(100),cout=>p(199)(101));
FA_ff_4581:FAff port map(x=>p(105)(101),y=>p(106)(101),Cin=>p(107)(101),clock=>clock,reset=>reset,s=>p(198)(101),cout=>p(199)(102));
FA_ff_4582:FAff port map(x=>p(105)(102),y=>p(106)(102),Cin=>p(107)(102),clock=>clock,reset=>reset,s=>p(198)(102),cout=>p(199)(103));
FA_ff_4583:FAff port map(x=>p(105)(103),y=>p(106)(103),Cin=>p(107)(103),clock=>clock,reset=>reset,s=>p(198)(103),cout=>p(199)(104));
FA_ff_4584:FAff port map(x=>p(105)(104),y=>p(106)(104),Cin=>p(107)(104),clock=>clock,reset=>reset,s=>p(198)(104),cout=>p(199)(105));
FA_ff_4585:FAff port map(x=>p(105)(105),y=>p(106)(105),Cin=>p(107)(105),clock=>clock,reset=>reset,s=>p(198)(105),cout=>p(199)(106));
FA_ff_4586:FAff port map(x=>p(105)(106),y=>p(106)(106),Cin=>p(107)(106),clock=>clock,reset=>reset,s=>p(198)(106),cout=>p(199)(107));
FA_ff_4587:FAff port map(x=>p(105)(107),y=>p(106)(107),Cin=>p(107)(107),clock=>clock,reset=>reset,s=>p(198)(107),cout=>p(199)(108));
FA_ff_4588:FAff port map(x=>p(105)(108),y=>p(106)(108),Cin=>p(107)(108),clock=>clock,reset=>reset,s=>p(198)(108),cout=>p(199)(109));
FA_ff_4589:FAff port map(x=>p(105)(109),y=>p(106)(109),Cin=>p(107)(109),clock=>clock,reset=>reset,s=>p(198)(109),cout=>p(199)(110));
FA_ff_4590:FAff port map(x=>p(105)(110),y=>p(106)(110),Cin=>p(107)(110),clock=>clock,reset=>reset,s=>p(198)(110),cout=>p(199)(111));
FA_ff_4591:FAff port map(x=>p(105)(111),y=>p(106)(111),Cin=>p(107)(111),clock=>clock,reset=>reset,s=>p(198)(111),cout=>p(199)(112));
FA_ff_4592:FAff port map(x=>p(105)(112),y=>p(106)(112),Cin=>p(107)(112),clock=>clock,reset=>reset,s=>p(198)(112),cout=>p(199)(113));
FA_ff_4593:FAff port map(x=>p(105)(113),y=>p(106)(113),Cin=>p(107)(113),clock=>clock,reset=>reset,s=>p(198)(113),cout=>p(199)(114));
FA_ff_4594:FAff port map(x=>p(105)(114),y=>p(106)(114),Cin=>p(107)(114),clock=>clock,reset=>reset,s=>p(198)(114),cout=>p(199)(115));
FA_ff_4595:FAff port map(x=>p(105)(115),y=>p(106)(115),Cin=>p(107)(115),clock=>clock,reset=>reset,s=>p(198)(115),cout=>p(199)(116));
FA_ff_4596:FAff port map(x=>p(105)(116),y=>p(106)(116),Cin=>p(107)(116),clock=>clock,reset=>reset,s=>p(198)(116),cout=>p(199)(117));
FA_ff_4597:FAff port map(x=>p(105)(117),y=>p(106)(117),Cin=>p(107)(117),clock=>clock,reset=>reset,s=>p(198)(117),cout=>p(199)(118));
FA_ff_4598:FAff port map(x=>p(105)(118),y=>p(106)(118),Cin=>p(107)(118),clock=>clock,reset=>reset,s=>p(198)(118),cout=>p(199)(119));
FA_ff_4599:FAff port map(x=>p(105)(119),y=>p(106)(119),Cin=>p(107)(119),clock=>clock,reset=>reset,s=>p(198)(119),cout=>p(199)(120));
FA_ff_4600:FAff port map(x=>p(105)(120),y=>p(106)(120),Cin=>p(107)(120),clock=>clock,reset=>reset,s=>p(198)(120),cout=>p(199)(121));
FA_ff_4601:FAff port map(x=>p(105)(121),y=>p(106)(121),Cin=>p(107)(121),clock=>clock,reset=>reset,s=>p(198)(121),cout=>p(199)(122));
FA_ff_4602:FAff port map(x=>p(105)(122),y=>p(106)(122),Cin=>p(107)(122),clock=>clock,reset=>reset,s=>p(198)(122),cout=>p(199)(123));
FA_ff_4603:FAff port map(x=>p(105)(123),y=>p(106)(123),Cin=>p(107)(123),clock=>clock,reset=>reset,s=>p(198)(123),cout=>p(199)(124));
FA_ff_4604:FAff port map(x=>p(105)(124),y=>p(106)(124),Cin=>p(107)(124),clock=>clock,reset=>reset,s=>p(198)(124),cout=>p(199)(125));
FA_ff_4605:FAff port map(x=>p(105)(125),y=>p(106)(125),Cin=>p(107)(125),clock=>clock,reset=>reset,s=>p(198)(125),cout=>p(199)(126));
FA_ff_4606:FAff port map(x=>p(105)(126),y=>p(106)(126),Cin=>p(107)(126),clock=>clock,reset=>reset,s=>p(198)(126),cout=>p(199)(127));
FA_ff_4607:FAff port map(x=>p(105)(127),y=>p(106)(127),Cin=>p(107)(127),clock=>clock,reset=>reset,s=>p(198)(127),cout=>p(199)(128));
FA_ff_4608:FAff port map(x=>p(108)(0),y=>p(109)(0),Cin=>p(110)(0),clock=>clock,reset=>reset,s=>p(200)(0),cout=>p(201)(1));
FA_ff_4609:FAff port map(x=>p(108)(1),y=>p(109)(1),Cin=>p(110)(1),clock=>clock,reset=>reset,s=>p(200)(1),cout=>p(201)(2));
FA_ff_4610:FAff port map(x=>p(108)(2),y=>p(109)(2),Cin=>p(110)(2),clock=>clock,reset=>reset,s=>p(200)(2),cout=>p(201)(3));
FA_ff_4611:FAff port map(x=>p(108)(3),y=>p(109)(3),Cin=>p(110)(3),clock=>clock,reset=>reset,s=>p(200)(3),cout=>p(201)(4));
FA_ff_4612:FAff port map(x=>p(108)(4),y=>p(109)(4),Cin=>p(110)(4),clock=>clock,reset=>reset,s=>p(200)(4),cout=>p(201)(5));
FA_ff_4613:FAff port map(x=>p(108)(5),y=>p(109)(5),Cin=>p(110)(5),clock=>clock,reset=>reset,s=>p(200)(5),cout=>p(201)(6));
FA_ff_4614:FAff port map(x=>p(108)(6),y=>p(109)(6),Cin=>p(110)(6),clock=>clock,reset=>reset,s=>p(200)(6),cout=>p(201)(7));
FA_ff_4615:FAff port map(x=>p(108)(7),y=>p(109)(7),Cin=>p(110)(7),clock=>clock,reset=>reset,s=>p(200)(7),cout=>p(201)(8));
FA_ff_4616:FAff port map(x=>p(108)(8),y=>p(109)(8),Cin=>p(110)(8),clock=>clock,reset=>reset,s=>p(200)(8),cout=>p(201)(9));
FA_ff_4617:FAff port map(x=>p(108)(9),y=>p(109)(9),Cin=>p(110)(9),clock=>clock,reset=>reset,s=>p(200)(9),cout=>p(201)(10));
FA_ff_4618:FAff port map(x=>p(108)(10),y=>p(109)(10),Cin=>p(110)(10),clock=>clock,reset=>reset,s=>p(200)(10),cout=>p(201)(11));
FA_ff_4619:FAff port map(x=>p(108)(11),y=>p(109)(11),Cin=>p(110)(11),clock=>clock,reset=>reset,s=>p(200)(11),cout=>p(201)(12));
FA_ff_4620:FAff port map(x=>p(108)(12),y=>p(109)(12),Cin=>p(110)(12),clock=>clock,reset=>reset,s=>p(200)(12),cout=>p(201)(13));
FA_ff_4621:FAff port map(x=>p(108)(13),y=>p(109)(13),Cin=>p(110)(13),clock=>clock,reset=>reset,s=>p(200)(13),cout=>p(201)(14));
FA_ff_4622:FAff port map(x=>p(108)(14),y=>p(109)(14),Cin=>p(110)(14),clock=>clock,reset=>reset,s=>p(200)(14),cout=>p(201)(15));
FA_ff_4623:FAff port map(x=>p(108)(15),y=>p(109)(15),Cin=>p(110)(15),clock=>clock,reset=>reset,s=>p(200)(15),cout=>p(201)(16));
FA_ff_4624:FAff port map(x=>p(108)(16),y=>p(109)(16),Cin=>p(110)(16),clock=>clock,reset=>reset,s=>p(200)(16),cout=>p(201)(17));
FA_ff_4625:FAff port map(x=>p(108)(17),y=>p(109)(17),Cin=>p(110)(17),clock=>clock,reset=>reset,s=>p(200)(17),cout=>p(201)(18));
FA_ff_4626:FAff port map(x=>p(108)(18),y=>p(109)(18),Cin=>p(110)(18),clock=>clock,reset=>reset,s=>p(200)(18),cout=>p(201)(19));
FA_ff_4627:FAff port map(x=>p(108)(19),y=>p(109)(19),Cin=>p(110)(19),clock=>clock,reset=>reset,s=>p(200)(19),cout=>p(201)(20));
FA_ff_4628:FAff port map(x=>p(108)(20),y=>p(109)(20),Cin=>p(110)(20),clock=>clock,reset=>reset,s=>p(200)(20),cout=>p(201)(21));
FA_ff_4629:FAff port map(x=>p(108)(21),y=>p(109)(21),Cin=>p(110)(21),clock=>clock,reset=>reset,s=>p(200)(21),cout=>p(201)(22));
FA_ff_4630:FAff port map(x=>p(108)(22),y=>p(109)(22),Cin=>p(110)(22),clock=>clock,reset=>reset,s=>p(200)(22),cout=>p(201)(23));
FA_ff_4631:FAff port map(x=>p(108)(23),y=>p(109)(23),Cin=>p(110)(23),clock=>clock,reset=>reset,s=>p(200)(23),cout=>p(201)(24));
FA_ff_4632:FAff port map(x=>p(108)(24),y=>p(109)(24),Cin=>p(110)(24),clock=>clock,reset=>reset,s=>p(200)(24),cout=>p(201)(25));
FA_ff_4633:FAff port map(x=>p(108)(25),y=>p(109)(25),Cin=>p(110)(25),clock=>clock,reset=>reset,s=>p(200)(25),cout=>p(201)(26));
FA_ff_4634:FAff port map(x=>p(108)(26),y=>p(109)(26),Cin=>p(110)(26),clock=>clock,reset=>reset,s=>p(200)(26),cout=>p(201)(27));
FA_ff_4635:FAff port map(x=>p(108)(27),y=>p(109)(27),Cin=>p(110)(27),clock=>clock,reset=>reset,s=>p(200)(27),cout=>p(201)(28));
FA_ff_4636:FAff port map(x=>p(108)(28),y=>p(109)(28),Cin=>p(110)(28),clock=>clock,reset=>reset,s=>p(200)(28),cout=>p(201)(29));
FA_ff_4637:FAff port map(x=>p(108)(29),y=>p(109)(29),Cin=>p(110)(29),clock=>clock,reset=>reset,s=>p(200)(29),cout=>p(201)(30));
FA_ff_4638:FAff port map(x=>p(108)(30),y=>p(109)(30),Cin=>p(110)(30),clock=>clock,reset=>reset,s=>p(200)(30),cout=>p(201)(31));
FA_ff_4639:FAff port map(x=>p(108)(31),y=>p(109)(31),Cin=>p(110)(31),clock=>clock,reset=>reset,s=>p(200)(31),cout=>p(201)(32));
FA_ff_4640:FAff port map(x=>p(108)(32),y=>p(109)(32),Cin=>p(110)(32),clock=>clock,reset=>reset,s=>p(200)(32),cout=>p(201)(33));
FA_ff_4641:FAff port map(x=>p(108)(33),y=>p(109)(33),Cin=>p(110)(33),clock=>clock,reset=>reset,s=>p(200)(33),cout=>p(201)(34));
FA_ff_4642:FAff port map(x=>p(108)(34),y=>p(109)(34),Cin=>p(110)(34),clock=>clock,reset=>reset,s=>p(200)(34),cout=>p(201)(35));
FA_ff_4643:FAff port map(x=>p(108)(35),y=>p(109)(35),Cin=>p(110)(35),clock=>clock,reset=>reset,s=>p(200)(35),cout=>p(201)(36));
FA_ff_4644:FAff port map(x=>p(108)(36),y=>p(109)(36),Cin=>p(110)(36),clock=>clock,reset=>reset,s=>p(200)(36),cout=>p(201)(37));
FA_ff_4645:FAff port map(x=>p(108)(37),y=>p(109)(37),Cin=>p(110)(37),clock=>clock,reset=>reset,s=>p(200)(37),cout=>p(201)(38));
FA_ff_4646:FAff port map(x=>p(108)(38),y=>p(109)(38),Cin=>p(110)(38),clock=>clock,reset=>reset,s=>p(200)(38),cout=>p(201)(39));
FA_ff_4647:FAff port map(x=>p(108)(39),y=>p(109)(39),Cin=>p(110)(39),clock=>clock,reset=>reset,s=>p(200)(39),cout=>p(201)(40));
FA_ff_4648:FAff port map(x=>p(108)(40),y=>p(109)(40),Cin=>p(110)(40),clock=>clock,reset=>reset,s=>p(200)(40),cout=>p(201)(41));
FA_ff_4649:FAff port map(x=>p(108)(41),y=>p(109)(41),Cin=>p(110)(41),clock=>clock,reset=>reset,s=>p(200)(41),cout=>p(201)(42));
FA_ff_4650:FAff port map(x=>p(108)(42),y=>p(109)(42),Cin=>p(110)(42),clock=>clock,reset=>reset,s=>p(200)(42),cout=>p(201)(43));
FA_ff_4651:FAff port map(x=>p(108)(43),y=>p(109)(43),Cin=>p(110)(43),clock=>clock,reset=>reset,s=>p(200)(43),cout=>p(201)(44));
FA_ff_4652:FAff port map(x=>p(108)(44),y=>p(109)(44),Cin=>p(110)(44),clock=>clock,reset=>reset,s=>p(200)(44),cout=>p(201)(45));
FA_ff_4653:FAff port map(x=>p(108)(45),y=>p(109)(45),Cin=>p(110)(45),clock=>clock,reset=>reset,s=>p(200)(45),cout=>p(201)(46));
FA_ff_4654:FAff port map(x=>p(108)(46),y=>p(109)(46),Cin=>p(110)(46),clock=>clock,reset=>reset,s=>p(200)(46),cout=>p(201)(47));
FA_ff_4655:FAff port map(x=>p(108)(47),y=>p(109)(47),Cin=>p(110)(47),clock=>clock,reset=>reset,s=>p(200)(47),cout=>p(201)(48));
FA_ff_4656:FAff port map(x=>p(108)(48),y=>p(109)(48),Cin=>p(110)(48),clock=>clock,reset=>reset,s=>p(200)(48),cout=>p(201)(49));
FA_ff_4657:FAff port map(x=>p(108)(49),y=>p(109)(49),Cin=>p(110)(49),clock=>clock,reset=>reset,s=>p(200)(49),cout=>p(201)(50));
FA_ff_4658:FAff port map(x=>p(108)(50),y=>p(109)(50),Cin=>p(110)(50),clock=>clock,reset=>reset,s=>p(200)(50),cout=>p(201)(51));
FA_ff_4659:FAff port map(x=>p(108)(51),y=>p(109)(51),Cin=>p(110)(51),clock=>clock,reset=>reset,s=>p(200)(51),cout=>p(201)(52));
FA_ff_4660:FAff port map(x=>p(108)(52),y=>p(109)(52),Cin=>p(110)(52),clock=>clock,reset=>reset,s=>p(200)(52),cout=>p(201)(53));
FA_ff_4661:FAff port map(x=>p(108)(53),y=>p(109)(53),Cin=>p(110)(53),clock=>clock,reset=>reset,s=>p(200)(53),cout=>p(201)(54));
FA_ff_4662:FAff port map(x=>p(108)(54),y=>p(109)(54),Cin=>p(110)(54),clock=>clock,reset=>reset,s=>p(200)(54),cout=>p(201)(55));
FA_ff_4663:FAff port map(x=>p(108)(55),y=>p(109)(55),Cin=>p(110)(55),clock=>clock,reset=>reset,s=>p(200)(55),cout=>p(201)(56));
FA_ff_4664:FAff port map(x=>p(108)(56),y=>p(109)(56),Cin=>p(110)(56),clock=>clock,reset=>reset,s=>p(200)(56),cout=>p(201)(57));
FA_ff_4665:FAff port map(x=>p(108)(57),y=>p(109)(57),Cin=>p(110)(57),clock=>clock,reset=>reset,s=>p(200)(57),cout=>p(201)(58));
FA_ff_4666:FAff port map(x=>p(108)(58),y=>p(109)(58),Cin=>p(110)(58),clock=>clock,reset=>reset,s=>p(200)(58),cout=>p(201)(59));
FA_ff_4667:FAff port map(x=>p(108)(59),y=>p(109)(59),Cin=>p(110)(59),clock=>clock,reset=>reset,s=>p(200)(59),cout=>p(201)(60));
FA_ff_4668:FAff port map(x=>p(108)(60),y=>p(109)(60),Cin=>p(110)(60),clock=>clock,reset=>reset,s=>p(200)(60),cout=>p(201)(61));
FA_ff_4669:FAff port map(x=>p(108)(61),y=>p(109)(61),Cin=>p(110)(61),clock=>clock,reset=>reset,s=>p(200)(61),cout=>p(201)(62));
FA_ff_4670:FAff port map(x=>p(108)(62),y=>p(109)(62),Cin=>p(110)(62),clock=>clock,reset=>reset,s=>p(200)(62),cout=>p(201)(63));
FA_ff_4671:FAff port map(x=>p(108)(63),y=>p(109)(63),Cin=>p(110)(63),clock=>clock,reset=>reset,s=>p(200)(63),cout=>p(201)(64));
FA_ff_4672:FAff port map(x=>p(108)(64),y=>p(109)(64),Cin=>p(110)(64),clock=>clock,reset=>reset,s=>p(200)(64),cout=>p(201)(65));
FA_ff_4673:FAff port map(x=>p(108)(65),y=>p(109)(65),Cin=>p(110)(65),clock=>clock,reset=>reset,s=>p(200)(65),cout=>p(201)(66));
FA_ff_4674:FAff port map(x=>p(108)(66),y=>p(109)(66),Cin=>p(110)(66),clock=>clock,reset=>reset,s=>p(200)(66),cout=>p(201)(67));
FA_ff_4675:FAff port map(x=>p(108)(67),y=>p(109)(67),Cin=>p(110)(67),clock=>clock,reset=>reset,s=>p(200)(67),cout=>p(201)(68));
FA_ff_4676:FAff port map(x=>p(108)(68),y=>p(109)(68),Cin=>p(110)(68),clock=>clock,reset=>reset,s=>p(200)(68),cout=>p(201)(69));
FA_ff_4677:FAff port map(x=>p(108)(69),y=>p(109)(69),Cin=>p(110)(69),clock=>clock,reset=>reset,s=>p(200)(69),cout=>p(201)(70));
FA_ff_4678:FAff port map(x=>p(108)(70),y=>p(109)(70),Cin=>p(110)(70),clock=>clock,reset=>reset,s=>p(200)(70),cout=>p(201)(71));
FA_ff_4679:FAff port map(x=>p(108)(71),y=>p(109)(71),Cin=>p(110)(71),clock=>clock,reset=>reset,s=>p(200)(71),cout=>p(201)(72));
FA_ff_4680:FAff port map(x=>p(108)(72),y=>p(109)(72),Cin=>p(110)(72),clock=>clock,reset=>reset,s=>p(200)(72),cout=>p(201)(73));
FA_ff_4681:FAff port map(x=>p(108)(73),y=>p(109)(73),Cin=>p(110)(73),clock=>clock,reset=>reset,s=>p(200)(73),cout=>p(201)(74));
FA_ff_4682:FAff port map(x=>p(108)(74),y=>p(109)(74),Cin=>p(110)(74),clock=>clock,reset=>reset,s=>p(200)(74),cout=>p(201)(75));
FA_ff_4683:FAff port map(x=>p(108)(75),y=>p(109)(75),Cin=>p(110)(75),clock=>clock,reset=>reset,s=>p(200)(75),cout=>p(201)(76));
FA_ff_4684:FAff port map(x=>p(108)(76),y=>p(109)(76),Cin=>p(110)(76),clock=>clock,reset=>reset,s=>p(200)(76),cout=>p(201)(77));
FA_ff_4685:FAff port map(x=>p(108)(77),y=>p(109)(77),Cin=>p(110)(77),clock=>clock,reset=>reset,s=>p(200)(77),cout=>p(201)(78));
FA_ff_4686:FAff port map(x=>p(108)(78),y=>p(109)(78),Cin=>p(110)(78),clock=>clock,reset=>reset,s=>p(200)(78),cout=>p(201)(79));
FA_ff_4687:FAff port map(x=>p(108)(79),y=>p(109)(79),Cin=>p(110)(79),clock=>clock,reset=>reset,s=>p(200)(79),cout=>p(201)(80));
FA_ff_4688:FAff port map(x=>p(108)(80),y=>p(109)(80),Cin=>p(110)(80),clock=>clock,reset=>reset,s=>p(200)(80),cout=>p(201)(81));
FA_ff_4689:FAff port map(x=>p(108)(81),y=>p(109)(81),Cin=>p(110)(81),clock=>clock,reset=>reset,s=>p(200)(81),cout=>p(201)(82));
FA_ff_4690:FAff port map(x=>p(108)(82),y=>p(109)(82),Cin=>p(110)(82),clock=>clock,reset=>reset,s=>p(200)(82),cout=>p(201)(83));
FA_ff_4691:FAff port map(x=>p(108)(83),y=>p(109)(83),Cin=>p(110)(83),clock=>clock,reset=>reset,s=>p(200)(83),cout=>p(201)(84));
FA_ff_4692:FAff port map(x=>p(108)(84),y=>p(109)(84),Cin=>p(110)(84),clock=>clock,reset=>reset,s=>p(200)(84),cout=>p(201)(85));
FA_ff_4693:FAff port map(x=>p(108)(85),y=>p(109)(85),Cin=>p(110)(85),clock=>clock,reset=>reset,s=>p(200)(85),cout=>p(201)(86));
FA_ff_4694:FAff port map(x=>p(108)(86),y=>p(109)(86),Cin=>p(110)(86),clock=>clock,reset=>reset,s=>p(200)(86),cout=>p(201)(87));
FA_ff_4695:FAff port map(x=>p(108)(87),y=>p(109)(87),Cin=>p(110)(87),clock=>clock,reset=>reset,s=>p(200)(87),cout=>p(201)(88));
FA_ff_4696:FAff port map(x=>p(108)(88),y=>p(109)(88),Cin=>p(110)(88),clock=>clock,reset=>reset,s=>p(200)(88),cout=>p(201)(89));
FA_ff_4697:FAff port map(x=>p(108)(89),y=>p(109)(89),Cin=>p(110)(89),clock=>clock,reset=>reset,s=>p(200)(89),cout=>p(201)(90));
FA_ff_4698:FAff port map(x=>p(108)(90),y=>p(109)(90),Cin=>p(110)(90),clock=>clock,reset=>reset,s=>p(200)(90),cout=>p(201)(91));
FA_ff_4699:FAff port map(x=>p(108)(91),y=>p(109)(91),Cin=>p(110)(91),clock=>clock,reset=>reset,s=>p(200)(91),cout=>p(201)(92));
FA_ff_4700:FAff port map(x=>p(108)(92),y=>p(109)(92),Cin=>p(110)(92),clock=>clock,reset=>reset,s=>p(200)(92),cout=>p(201)(93));
FA_ff_4701:FAff port map(x=>p(108)(93),y=>p(109)(93),Cin=>p(110)(93),clock=>clock,reset=>reset,s=>p(200)(93),cout=>p(201)(94));
FA_ff_4702:FAff port map(x=>p(108)(94),y=>p(109)(94),Cin=>p(110)(94),clock=>clock,reset=>reset,s=>p(200)(94),cout=>p(201)(95));
FA_ff_4703:FAff port map(x=>p(108)(95),y=>p(109)(95),Cin=>p(110)(95),clock=>clock,reset=>reset,s=>p(200)(95),cout=>p(201)(96));
FA_ff_4704:FAff port map(x=>p(108)(96),y=>p(109)(96),Cin=>p(110)(96),clock=>clock,reset=>reset,s=>p(200)(96),cout=>p(201)(97));
FA_ff_4705:FAff port map(x=>p(108)(97),y=>p(109)(97),Cin=>p(110)(97),clock=>clock,reset=>reset,s=>p(200)(97),cout=>p(201)(98));
FA_ff_4706:FAff port map(x=>p(108)(98),y=>p(109)(98),Cin=>p(110)(98),clock=>clock,reset=>reset,s=>p(200)(98),cout=>p(201)(99));
FA_ff_4707:FAff port map(x=>p(108)(99),y=>p(109)(99),Cin=>p(110)(99),clock=>clock,reset=>reset,s=>p(200)(99),cout=>p(201)(100));
FA_ff_4708:FAff port map(x=>p(108)(100),y=>p(109)(100),Cin=>p(110)(100),clock=>clock,reset=>reset,s=>p(200)(100),cout=>p(201)(101));
FA_ff_4709:FAff port map(x=>p(108)(101),y=>p(109)(101),Cin=>p(110)(101),clock=>clock,reset=>reset,s=>p(200)(101),cout=>p(201)(102));
FA_ff_4710:FAff port map(x=>p(108)(102),y=>p(109)(102),Cin=>p(110)(102),clock=>clock,reset=>reset,s=>p(200)(102),cout=>p(201)(103));
FA_ff_4711:FAff port map(x=>p(108)(103),y=>p(109)(103),Cin=>p(110)(103),clock=>clock,reset=>reset,s=>p(200)(103),cout=>p(201)(104));
FA_ff_4712:FAff port map(x=>p(108)(104),y=>p(109)(104),Cin=>p(110)(104),clock=>clock,reset=>reset,s=>p(200)(104),cout=>p(201)(105));
FA_ff_4713:FAff port map(x=>p(108)(105),y=>p(109)(105),Cin=>p(110)(105),clock=>clock,reset=>reset,s=>p(200)(105),cout=>p(201)(106));
FA_ff_4714:FAff port map(x=>p(108)(106),y=>p(109)(106),Cin=>p(110)(106),clock=>clock,reset=>reset,s=>p(200)(106),cout=>p(201)(107));
FA_ff_4715:FAff port map(x=>p(108)(107),y=>p(109)(107),Cin=>p(110)(107),clock=>clock,reset=>reset,s=>p(200)(107),cout=>p(201)(108));
FA_ff_4716:FAff port map(x=>p(108)(108),y=>p(109)(108),Cin=>p(110)(108),clock=>clock,reset=>reset,s=>p(200)(108),cout=>p(201)(109));
FA_ff_4717:FAff port map(x=>p(108)(109),y=>p(109)(109),Cin=>p(110)(109),clock=>clock,reset=>reset,s=>p(200)(109),cout=>p(201)(110));
FA_ff_4718:FAff port map(x=>p(108)(110),y=>p(109)(110),Cin=>p(110)(110),clock=>clock,reset=>reset,s=>p(200)(110),cout=>p(201)(111));
FA_ff_4719:FAff port map(x=>p(108)(111),y=>p(109)(111),Cin=>p(110)(111),clock=>clock,reset=>reset,s=>p(200)(111),cout=>p(201)(112));
FA_ff_4720:FAff port map(x=>p(108)(112),y=>p(109)(112),Cin=>p(110)(112),clock=>clock,reset=>reset,s=>p(200)(112),cout=>p(201)(113));
FA_ff_4721:FAff port map(x=>p(108)(113),y=>p(109)(113),Cin=>p(110)(113),clock=>clock,reset=>reset,s=>p(200)(113),cout=>p(201)(114));
FA_ff_4722:FAff port map(x=>p(108)(114),y=>p(109)(114),Cin=>p(110)(114),clock=>clock,reset=>reset,s=>p(200)(114),cout=>p(201)(115));
FA_ff_4723:FAff port map(x=>p(108)(115),y=>p(109)(115),Cin=>p(110)(115),clock=>clock,reset=>reset,s=>p(200)(115),cout=>p(201)(116));
FA_ff_4724:FAff port map(x=>p(108)(116),y=>p(109)(116),Cin=>p(110)(116),clock=>clock,reset=>reset,s=>p(200)(116),cout=>p(201)(117));
FA_ff_4725:FAff port map(x=>p(108)(117),y=>p(109)(117),Cin=>p(110)(117),clock=>clock,reset=>reset,s=>p(200)(117),cout=>p(201)(118));
FA_ff_4726:FAff port map(x=>p(108)(118),y=>p(109)(118),Cin=>p(110)(118),clock=>clock,reset=>reset,s=>p(200)(118),cout=>p(201)(119));
FA_ff_4727:FAff port map(x=>p(108)(119),y=>p(109)(119),Cin=>p(110)(119),clock=>clock,reset=>reset,s=>p(200)(119),cout=>p(201)(120));
FA_ff_4728:FAff port map(x=>p(108)(120),y=>p(109)(120),Cin=>p(110)(120),clock=>clock,reset=>reset,s=>p(200)(120),cout=>p(201)(121));
FA_ff_4729:FAff port map(x=>p(108)(121),y=>p(109)(121),Cin=>p(110)(121),clock=>clock,reset=>reset,s=>p(200)(121),cout=>p(201)(122));
FA_ff_4730:FAff port map(x=>p(108)(122),y=>p(109)(122),Cin=>p(110)(122),clock=>clock,reset=>reset,s=>p(200)(122),cout=>p(201)(123));
FA_ff_4731:FAff port map(x=>p(108)(123),y=>p(109)(123),Cin=>p(110)(123),clock=>clock,reset=>reset,s=>p(200)(123),cout=>p(201)(124));
FA_ff_4732:FAff port map(x=>p(108)(124),y=>p(109)(124),Cin=>p(110)(124),clock=>clock,reset=>reset,s=>p(200)(124),cout=>p(201)(125));
FA_ff_4733:FAff port map(x=>p(108)(125),y=>p(109)(125),Cin=>p(110)(125),clock=>clock,reset=>reset,s=>p(200)(125),cout=>p(201)(126));
FA_ff_4734:FAff port map(x=>p(108)(126),y=>p(109)(126),Cin=>p(110)(126),clock=>clock,reset=>reset,s=>p(200)(126),cout=>p(201)(127));
FA_ff_4735:FAff port map(x=>p(108)(127),y=>p(109)(127),Cin=>p(110)(127),clock=>clock,reset=>reset,s=>p(200)(127),cout=>p(201)(128));
FA_ff_4736:FAff port map(x=>p(111)(0),y=>p(112)(0),Cin=>p(113)(0),clock=>clock,reset=>reset,s=>p(202)(0),cout=>p(203)(1));
FA_ff_4737:FAff port map(x=>p(111)(1),y=>p(112)(1),Cin=>p(113)(1),clock=>clock,reset=>reset,s=>p(202)(1),cout=>p(203)(2));
FA_ff_4738:FAff port map(x=>p(111)(2),y=>p(112)(2),Cin=>p(113)(2),clock=>clock,reset=>reset,s=>p(202)(2),cout=>p(203)(3));
FA_ff_4739:FAff port map(x=>p(111)(3),y=>p(112)(3),Cin=>p(113)(3),clock=>clock,reset=>reset,s=>p(202)(3),cout=>p(203)(4));
FA_ff_4740:FAff port map(x=>p(111)(4),y=>p(112)(4),Cin=>p(113)(4),clock=>clock,reset=>reset,s=>p(202)(4),cout=>p(203)(5));
FA_ff_4741:FAff port map(x=>p(111)(5),y=>p(112)(5),Cin=>p(113)(5),clock=>clock,reset=>reset,s=>p(202)(5),cout=>p(203)(6));
FA_ff_4742:FAff port map(x=>p(111)(6),y=>p(112)(6),Cin=>p(113)(6),clock=>clock,reset=>reset,s=>p(202)(6),cout=>p(203)(7));
FA_ff_4743:FAff port map(x=>p(111)(7),y=>p(112)(7),Cin=>p(113)(7),clock=>clock,reset=>reset,s=>p(202)(7),cout=>p(203)(8));
FA_ff_4744:FAff port map(x=>p(111)(8),y=>p(112)(8),Cin=>p(113)(8),clock=>clock,reset=>reset,s=>p(202)(8),cout=>p(203)(9));
FA_ff_4745:FAff port map(x=>p(111)(9),y=>p(112)(9),Cin=>p(113)(9),clock=>clock,reset=>reset,s=>p(202)(9),cout=>p(203)(10));
FA_ff_4746:FAff port map(x=>p(111)(10),y=>p(112)(10),Cin=>p(113)(10),clock=>clock,reset=>reset,s=>p(202)(10),cout=>p(203)(11));
FA_ff_4747:FAff port map(x=>p(111)(11),y=>p(112)(11),Cin=>p(113)(11),clock=>clock,reset=>reset,s=>p(202)(11),cout=>p(203)(12));
FA_ff_4748:FAff port map(x=>p(111)(12),y=>p(112)(12),Cin=>p(113)(12),clock=>clock,reset=>reset,s=>p(202)(12),cout=>p(203)(13));
FA_ff_4749:FAff port map(x=>p(111)(13),y=>p(112)(13),Cin=>p(113)(13),clock=>clock,reset=>reset,s=>p(202)(13),cout=>p(203)(14));
FA_ff_4750:FAff port map(x=>p(111)(14),y=>p(112)(14),Cin=>p(113)(14),clock=>clock,reset=>reset,s=>p(202)(14),cout=>p(203)(15));
FA_ff_4751:FAff port map(x=>p(111)(15),y=>p(112)(15),Cin=>p(113)(15),clock=>clock,reset=>reset,s=>p(202)(15),cout=>p(203)(16));
FA_ff_4752:FAff port map(x=>p(111)(16),y=>p(112)(16),Cin=>p(113)(16),clock=>clock,reset=>reset,s=>p(202)(16),cout=>p(203)(17));
FA_ff_4753:FAff port map(x=>p(111)(17),y=>p(112)(17),Cin=>p(113)(17),clock=>clock,reset=>reset,s=>p(202)(17),cout=>p(203)(18));
FA_ff_4754:FAff port map(x=>p(111)(18),y=>p(112)(18),Cin=>p(113)(18),clock=>clock,reset=>reset,s=>p(202)(18),cout=>p(203)(19));
FA_ff_4755:FAff port map(x=>p(111)(19),y=>p(112)(19),Cin=>p(113)(19),clock=>clock,reset=>reset,s=>p(202)(19),cout=>p(203)(20));
FA_ff_4756:FAff port map(x=>p(111)(20),y=>p(112)(20),Cin=>p(113)(20),clock=>clock,reset=>reset,s=>p(202)(20),cout=>p(203)(21));
FA_ff_4757:FAff port map(x=>p(111)(21),y=>p(112)(21),Cin=>p(113)(21),clock=>clock,reset=>reset,s=>p(202)(21),cout=>p(203)(22));
FA_ff_4758:FAff port map(x=>p(111)(22),y=>p(112)(22),Cin=>p(113)(22),clock=>clock,reset=>reset,s=>p(202)(22),cout=>p(203)(23));
FA_ff_4759:FAff port map(x=>p(111)(23),y=>p(112)(23),Cin=>p(113)(23),clock=>clock,reset=>reset,s=>p(202)(23),cout=>p(203)(24));
FA_ff_4760:FAff port map(x=>p(111)(24),y=>p(112)(24),Cin=>p(113)(24),clock=>clock,reset=>reset,s=>p(202)(24),cout=>p(203)(25));
FA_ff_4761:FAff port map(x=>p(111)(25),y=>p(112)(25),Cin=>p(113)(25),clock=>clock,reset=>reset,s=>p(202)(25),cout=>p(203)(26));
FA_ff_4762:FAff port map(x=>p(111)(26),y=>p(112)(26),Cin=>p(113)(26),clock=>clock,reset=>reset,s=>p(202)(26),cout=>p(203)(27));
FA_ff_4763:FAff port map(x=>p(111)(27),y=>p(112)(27),Cin=>p(113)(27),clock=>clock,reset=>reset,s=>p(202)(27),cout=>p(203)(28));
FA_ff_4764:FAff port map(x=>p(111)(28),y=>p(112)(28),Cin=>p(113)(28),clock=>clock,reset=>reset,s=>p(202)(28),cout=>p(203)(29));
FA_ff_4765:FAff port map(x=>p(111)(29),y=>p(112)(29),Cin=>p(113)(29),clock=>clock,reset=>reset,s=>p(202)(29),cout=>p(203)(30));
FA_ff_4766:FAff port map(x=>p(111)(30),y=>p(112)(30),Cin=>p(113)(30),clock=>clock,reset=>reset,s=>p(202)(30),cout=>p(203)(31));
FA_ff_4767:FAff port map(x=>p(111)(31),y=>p(112)(31),Cin=>p(113)(31),clock=>clock,reset=>reset,s=>p(202)(31),cout=>p(203)(32));
FA_ff_4768:FAff port map(x=>p(111)(32),y=>p(112)(32),Cin=>p(113)(32),clock=>clock,reset=>reset,s=>p(202)(32),cout=>p(203)(33));
FA_ff_4769:FAff port map(x=>p(111)(33),y=>p(112)(33),Cin=>p(113)(33),clock=>clock,reset=>reset,s=>p(202)(33),cout=>p(203)(34));
FA_ff_4770:FAff port map(x=>p(111)(34),y=>p(112)(34),Cin=>p(113)(34),clock=>clock,reset=>reset,s=>p(202)(34),cout=>p(203)(35));
FA_ff_4771:FAff port map(x=>p(111)(35),y=>p(112)(35),Cin=>p(113)(35),clock=>clock,reset=>reset,s=>p(202)(35),cout=>p(203)(36));
FA_ff_4772:FAff port map(x=>p(111)(36),y=>p(112)(36),Cin=>p(113)(36),clock=>clock,reset=>reset,s=>p(202)(36),cout=>p(203)(37));
FA_ff_4773:FAff port map(x=>p(111)(37),y=>p(112)(37),Cin=>p(113)(37),clock=>clock,reset=>reset,s=>p(202)(37),cout=>p(203)(38));
FA_ff_4774:FAff port map(x=>p(111)(38),y=>p(112)(38),Cin=>p(113)(38),clock=>clock,reset=>reset,s=>p(202)(38),cout=>p(203)(39));
FA_ff_4775:FAff port map(x=>p(111)(39),y=>p(112)(39),Cin=>p(113)(39),clock=>clock,reset=>reset,s=>p(202)(39),cout=>p(203)(40));
FA_ff_4776:FAff port map(x=>p(111)(40),y=>p(112)(40),Cin=>p(113)(40),clock=>clock,reset=>reset,s=>p(202)(40),cout=>p(203)(41));
FA_ff_4777:FAff port map(x=>p(111)(41),y=>p(112)(41),Cin=>p(113)(41),clock=>clock,reset=>reset,s=>p(202)(41),cout=>p(203)(42));
FA_ff_4778:FAff port map(x=>p(111)(42),y=>p(112)(42),Cin=>p(113)(42),clock=>clock,reset=>reset,s=>p(202)(42),cout=>p(203)(43));
FA_ff_4779:FAff port map(x=>p(111)(43),y=>p(112)(43),Cin=>p(113)(43),clock=>clock,reset=>reset,s=>p(202)(43),cout=>p(203)(44));
FA_ff_4780:FAff port map(x=>p(111)(44),y=>p(112)(44),Cin=>p(113)(44),clock=>clock,reset=>reset,s=>p(202)(44),cout=>p(203)(45));
FA_ff_4781:FAff port map(x=>p(111)(45),y=>p(112)(45),Cin=>p(113)(45),clock=>clock,reset=>reset,s=>p(202)(45),cout=>p(203)(46));
FA_ff_4782:FAff port map(x=>p(111)(46),y=>p(112)(46),Cin=>p(113)(46),clock=>clock,reset=>reset,s=>p(202)(46),cout=>p(203)(47));
FA_ff_4783:FAff port map(x=>p(111)(47),y=>p(112)(47),Cin=>p(113)(47),clock=>clock,reset=>reset,s=>p(202)(47),cout=>p(203)(48));
FA_ff_4784:FAff port map(x=>p(111)(48),y=>p(112)(48),Cin=>p(113)(48),clock=>clock,reset=>reset,s=>p(202)(48),cout=>p(203)(49));
FA_ff_4785:FAff port map(x=>p(111)(49),y=>p(112)(49),Cin=>p(113)(49),clock=>clock,reset=>reset,s=>p(202)(49),cout=>p(203)(50));
FA_ff_4786:FAff port map(x=>p(111)(50),y=>p(112)(50),Cin=>p(113)(50),clock=>clock,reset=>reset,s=>p(202)(50),cout=>p(203)(51));
FA_ff_4787:FAff port map(x=>p(111)(51),y=>p(112)(51),Cin=>p(113)(51),clock=>clock,reset=>reset,s=>p(202)(51),cout=>p(203)(52));
FA_ff_4788:FAff port map(x=>p(111)(52),y=>p(112)(52),Cin=>p(113)(52),clock=>clock,reset=>reset,s=>p(202)(52),cout=>p(203)(53));
FA_ff_4789:FAff port map(x=>p(111)(53),y=>p(112)(53),Cin=>p(113)(53),clock=>clock,reset=>reset,s=>p(202)(53),cout=>p(203)(54));
FA_ff_4790:FAff port map(x=>p(111)(54),y=>p(112)(54),Cin=>p(113)(54),clock=>clock,reset=>reset,s=>p(202)(54),cout=>p(203)(55));
FA_ff_4791:FAff port map(x=>p(111)(55),y=>p(112)(55),Cin=>p(113)(55),clock=>clock,reset=>reset,s=>p(202)(55),cout=>p(203)(56));
FA_ff_4792:FAff port map(x=>p(111)(56),y=>p(112)(56),Cin=>p(113)(56),clock=>clock,reset=>reset,s=>p(202)(56),cout=>p(203)(57));
FA_ff_4793:FAff port map(x=>p(111)(57),y=>p(112)(57),Cin=>p(113)(57),clock=>clock,reset=>reset,s=>p(202)(57),cout=>p(203)(58));
FA_ff_4794:FAff port map(x=>p(111)(58),y=>p(112)(58),Cin=>p(113)(58),clock=>clock,reset=>reset,s=>p(202)(58),cout=>p(203)(59));
FA_ff_4795:FAff port map(x=>p(111)(59),y=>p(112)(59),Cin=>p(113)(59),clock=>clock,reset=>reset,s=>p(202)(59),cout=>p(203)(60));
FA_ff_4796:FAff port map(x=>p(111)(60),y=>p(112)(60),Cin=>p(113)(60),clock=>clock,reset=>reset,s=>p(202)(60),cout=>p(203)(61));
FA_ff_4797:FAff port map(x=>p(111)(61),y=>p(112)(61),Cin=>p(113)(61),clock=>clock,reset=>reset,s=>p(202)(61),cout=>p(203)(62));
FA_ff_4798:FAff port map(x=>p(111)(62),y=>p(112)(62),Cin=>p(113)(62),clock=>clock,reset=>reset,s=>p(202)(62),cout=>p(203)(63));
FA_ff_4799:FAff port map(x=>p(111)(63),y=>p(112)(63),Cin=>p(113)(63),clock=>clock,reset=>reset,s=>p(202)(63),cout=>p(203)(64));
FA_ff_4800:FAff port map(x=>p(111)(64),y=>p(112)(64),Cin=>p(113)(64),clock=>clock,reset=>reset,s=>p(202)(64),cout=>p(203)(65));
FA_ff_4801:FAff port map(x=>p(111)(65),y=>p(112)(65),Cin=>p(113)(65),clock=>clock,reset=>reset,s=>p(202)(65),cout=>p(203)(66));
FA_ff_4802:FAff port map(x=>p(111)(66),y=>p(112)(66),Cin=>p(113)(66),clock=>clock,reset=>reset,s=>p(202)(66),cout=>p(203)(67));
FA_ff_4803:FAff port map(x=>p(111)(67),y=>p(112)(67),Cin=>p(113)(67),clock=>clock,reset=>reset,s=>p(202)(67),cout=>p(203)(68));
FA_ff_4804:FAff port map(x=>p(111)(68),y=>p(112)(68),Cin=>p(113)(68),clock=>clock,reset=>reset,s=>p(202)(68),cout=>p(203)(69));
FA_ff_4805:FAff port map(x=>p(111)(69),y=>p(112)(69),Cin=>p(113)(69),clock=>clock,reset=>reset,s=>p(202)(69),cout=>p(203)(70));
FA_ff_4806:FAff port map(x=>p(111)(70),y=>p(112)(70),Cin=>p(113)(70),clock=>clock,reset=>reset,s=>p(202)(70),cout=>p(203)(71));
FA_ff_4807:FAff port map(x=>p(111)(71),y=>p(112)(71),Cin=>p(113)(71),clock=>clock,reset=>reset,s=>p(202)(71),cout=>p(203)(72));
FA_ff_4808:FAff port map(x=>p(111)(72),y=>p(112)(72),Cin=>p(113)(72),clock=>clock,reset=>reset,s=>p(202)(72),cout=>p(203)(73));
FA_ff_4809:FAff port map(x=>p(111)(73),y=>p(112)(73),Cin=>p(113)(73),clock=>clock,reset=>reset,s=>p(202)(73),cout=>p(203)(74));
FA_ff_4810:FAff port map(x=>p(111)(74),y=>p(112)(74),Cin=>p(113)(74),clock=>clock,reset=>reset,s=>p(202)(74),cout=>p(203)(75));
FA_ff_4811:FAff port map(x=>p(111)(75),y=>p(112)(75),Cin=>p(113)(75),clock=>clock,reset=>reset,s=>p(202)(75),cout=>p(203)(76));
FA_ff_4812:FAff port map(x=>p(111)(76),y=>p(112)(76),Cin=>p(113)(76),clock=>clock,reset=>reset,s=>p(202)(76),cout=>p(203)(77));
FA_ff_4813:FAff port map(x=>p(111)(77),y=>p(112)(77),Cin=>p(113)(77),clock=>clock,reset=>reset,s=>p(202)(77),cout=>p(203)(78));
FA_ff_4814:FAff port map(x=>p(111)(78),y=>p(112)(78),Cin=>p(113)(78),clock=>clock,reset=>reset,s=>p(202)(78),cout=>p(203)(79));
FA_ff_4815:FAff port map(x=>p(111)(79),y=>p(112)(79),Cin=>p(113)(79),clock=>clock,reset=>reset,s=>p(202)(79),cout=>p(203)(80));
FA_ff_4816:FAff port map(x=>p(111)(80),y=>p(112)(80),Cin=>p(113)(80),clock=>clock,reset=>reset,s=>p(202)(80),cout=>p(203)(81));
FA_ff_4817:FAff port map(x=>p(111)(81),y=>p(112)(81),Cin=>p(113)(81),clock=>clock,reset=>reset,s=>p(202)(81),cout=>p(203)(82));
FA_ff_4818:FAff port map(x=>p(111)(82),y=>p(112)(82),Cin=>p(113)(82),clock=>clock,reset=>reset,s=>p(202)(82),cout=>p(203)(83));
FA_ff_4819:FAff port map(x=>p(111)(83),y=>p(112)(83),Cin=>p(113)(83),clock=>clock,reset=>reset,s=>p(202)(83),cout=>p(203)(84));
FA_ff_4820:FAff port map(x=>p(111)(84),y=>p(112)(84),Cin=>p(113)(84),clock=>clock,reset=>reset,s=>p(202)(84),cout=>p(203)(85));
FA_ff_4821:FAff port map(x=>p(111)(85),y=>p(112)(85),Cin=>p(113)(85),clock=>clock,reset=>reset,s=>p(202)(85),cout=>p(203)(86));
FA_ff_4822:FAff port map(x=>p(111)(86),y=>p(112)(86),Cin=>p(113)(86),clock=>clock,reset=>reset,s=>p(202)(86),cout=>p(203)(87));
FA_ff_4823:FAff port map(x=>p(111)(87),y=>p(112)(87),Cin=>p(113)(87),clock=>clock,reset=>reset,s=>p(202)(87),cout=>p(203)(88));
FA_ff_4824:FAff port map(x=>p(111)(88),y=>p(112)(88),Cin=>p(113)(88),clock=>clock,reset=>reset,s=>p(202)(88),cout=>p(203)(89));
FA_ff_4825:FAff port map(x=>p(111)(89),y=>p(112)(89),Cin=>p(113)(89),clock=>clock,reset=>reset,s=>p(202)(89),cout=>p(203)(90));
FA_ff_4826:FAff port map(x=>p(111)(90),y=>p(112)(90),Cin=>p(113)(90),clock=>clock,reset=>reset,s=>p(202)(90),cout=>p(203)(91));
FA_ff_4827:FAff port map(x=>p(111)(91),y=>p(112)(91),Cin=>p(113)(91),clock=>clock,reset=>reset,s=>p(202)(91),cout=>p(203)(92));
FA_ff_4828:FAff port map(x=>p(111)(92),y=>p(112)(92),Cin=>p(113)(92),clock=>clock,reset=>reset,s=>p(202)(92),cout=>p(203)(93));
FA_ff_4829:FAff port map(x=>p(111)(93),y=>p(112)(93),Cin=>p(113)(93),clock=>clock,reset=>reset,s=>p(202)(93),cout=>p(203)(94));
FA_ff_4830:FAff port map(x=>p(111)(94),y=>p(112)(94),Cin=>p(113)(94),clock=>clock,reset=>reset,s=>p(202)(94),cout=>p(203)(95));
FA_ff_4831:FAff port map(x=>p(111)(95),y=>p(112)(95),Cin=>p(113)(95),clock=>clock,reset=>reset,s=>p(202)(95),cout=>p(203)(96));
FA_ff_4832:FAff port map(x=>p(111)(96),y=>p(112)(96),Cin=>p(113)(96),clock=>clock,reset=>reset,s=>p(202)(96),cout=>p(203)(97));
FA_ff_4833:FAff port map(x=>p(111)(97),y=>p(112)(97),Cin=>p(113)(97),clock=>clock,reset=>reset,s=>p(202)(97),cout=>p(203)(98));
FA_ff_4834:FAff port map(x=>p(111)(98),y=>p(112)(98),Cin=>p(113)(98),clock=>clock,reset=>reset,s=>p(202)(98),cout=>p(203)(99));
FA_ff_4835:FAff port map(x=>p(111)(99),y=>p(112)(99),Cin=>p(113)(99),clock=>clock,reset=>reset,s=>p(202)(99),cout=>p(203)(100));
FA_ff_4836:FAff port map(x=>p(111)(100),y=>p(112)(100),Cin=>p(113)(100),clock=>clock,reset=>reset,s=>p(202)(100),cout=>p(203)(101));
FA_ff_4837:FAff port map(x=>p(111)(101),y=>p(112)(101),Cin=>p(113)(101),clock=>clock,reset=>reset,s=>p(202)(101),cout=>p(203)(102));
FA_ff_4838:FAff port map(x=>p(111)(102),y=>p(112)(102),Cin=>p(113)(102),clock=>clock,reset=>reset,s=>p(202)(102),cout=>p(203)(103));
FA_ff_4839:FAff port map(x=>p(111)(103),y=>p(112)(103),Cin=>p(113)(103),clock=>clock,reset=>reset,s=>p(202)(103),cout=>p(203)(104));
FA_ff_4840:FAff port map(x=>p(111)(104),y=>p(112)(104),Cin=>p(113)(104),clock=>clock,reset=>reset,s=>p(202)(104),cout=>p(203)(105));
FA_ff_4841:FAff port map(x=>p(111)(105),y=>p(112)(105),Cin=>p(113)(105),clock=>clock,reset=>reset,s=>p(202)(105),cout=>p(203)(106));
FA_ff_4842:FAff port map(x=>p(111)(106),y=>p(112)(106),Cin=>p(113)(106),clock=>clock,reset=>reset,s=>p(202)(106),cout=>p(203)(107));
FA_ff_4843:FAff port map(x=>p(111)(107),y=>p(112)(107),Cin=>p(113)(107),clock=>clock,reset=>reset,s=>p(202)(107),cout=>p(203)(108));
FA_ff_4844:FAff port map(x=>p(111)(108),y=>p(112)(108),Cin=>p(113)(108),clock=>clock,reset=>reset,s=>p(202)(108),cout=>p(203)(109));
FA_ff_4845:FAff port map(x=>p(111)(109),y=>p(112)(109),Cin=>p(113)(109),clock=>clock,reset=>reset,s=>p(202)(109),cout=>p(203)(110));
FA_ff_4846:FAff port map(x=>p(111)(110),y=>p(112)(110),Cin=>p(113)(110),clock=>clock,reset=>reset,s=>p(202)(110),cout=>p(203)(111));
FA_ff_4847:FAff port map(x=>p(111)(111),y=>p(112)(111),Cin=>p(113)(111),clock=>clock,reset=>reset,s=>p(202)(111),cout=>p(203)(112));
FA_ff_4848:FAff port map(x=>p(111)(112),y=>p(112)(112),Cin=>p(113)(112),clock=>clock,reset=>reset,s=>p(202)(112),cout=>p(203)(113));
FA_ff_4849:FAff port map(x=>p(111)(113),y=>p(112)(113),Cin=>p(113)(113),clock=>clock,reset=>reset,s=>p(202)(113),cout=>p(203)(114));
FA_ff_4850:FAff port map(x=>p(111)(114),y=>p(112)(114),Cin=>p(113)(114),clock=>clock,reset=>reset,s=>p(202)(114),cout=>p(203)(115));
FA_ff_4851:FAff port map(x=>p(111)(115),y=>p(112)(115),Cin=>p(113)(115),clock=>clock,reset=>reset,s=>p(202)(115),cout=>p(203)(116));
FA_ff_4852:FAff port map(x=>p(111)(116),y=>p(112)(116),Cin=>p(113)(116),clock=>clock,reset=>reset,s=>p(202)(116),cout=>p(203)(117));
FA_ff_4853:FAff port map(x=>p(111)(117),y=>p(112)(117),Cin=>p(113)(117),clock=>clock,reset=>reset,s=>p(202)(117),cout=>p(203)(118));
FA_ff_4854:FAff port map(x=>p(111)(118),y=>p(112)(118),Cin=>p(113)(118),clock=>clock,reset=>reset,s=>p(202)(118),cout=>p(203)(119));
FA_ff_4855:FAff port map(x=>p(111)(119),y=>p(112)(119),Cin=>p(113)(119),clock=>clock,reset=>reset,s=>p(202)(119),cout=>p(203)(120));
FA_ff_4856:FAff port map(x=>p(111)(120),y=>p(112)(120),Cin=>p(113)(120),clock=>clock,reset=>reset,s=>p(202)(120),cout=>p(203)(121));
FA_ff_4857:FAff port map(x=>p(111)(121),y=>p(112)(121),Cin=>p(113)(121),clock=>clock,reset=>reset,s=>p(202)(121),cout=>p(203)(122));
FA_ff_4858:FAff port map(x=>p(111)(122),y=>p(112)(122),Cin=>p(113)(122),clock=>clock,reset=>reset,s=>p(202)(122),cout=>p(203)(123));
FA_ff_4859:FAff port map(x=>p(111)(123),y=>p(112)(123),Cin=>p(113)(123),clock=>clock,reset=>reset,s=>p(202)(123),cout=>p(203)(124));
FA_ff_4860:FAff port map(x=>p(111)(124),y=>p(112)(124),Cin=>p(113)(124),clock=>clock,reset=>reset,s=>p(202)(124),cout=>p(203)(125));
FA_ff_4861:FAff port map(x=>p(111)(125),y=>p(112)(125),Cin=>p(113)(125),clock=>clock,reset=>reset,s=>p(202)(125),cout=>p(203)(126));
FA_ff_4862:FAff port map(x=>p(111)(126),y=>p(112)(126),Cin=>p(113)(126),clock=>clock,reset=>reset,s=>p(202)(126),cout=>p(203)(127));
FA_ff_4863:FAff port map(x=>p(111)(127),y=>p(112)(127),Cin=>p(113)(127),clock=>clock,reset=>reset,s=>p(202)(127),cout=>p(203)(128));
FA_ff_4864:FAff port map(x=>p(114)(0),y=>p(115)(0),Cin=>p(116)(0),clock=>clock,reset=>reset,s=>p(204)(0),cout=>p(205)(1));
FA_ff_4865:FAff port map(x=>p(114)(1),y=>p(115)(1),Cin=>p(116)(1),clock=>clock,reset=>reset,s=>p(204)(1),cout=>p(205)(2));
FA_ff_4866:FAff port map(x=>p(114)(2),y=>p(115)(2),Cin=>p(116)(2),clock=>clock,reset=>reset,s=>p(204)(2),cout=>p(205)(3));
FA_ff_4867:FAff port map(x=>p(114)(3),y=>p(115)(3),Cin=>p(116)(3),clock=>clock,reset=>reset,s=>p(204)(3),cout=>p(205)(4));
FA_ff_4868:FAff port map(x=>p(114)(4),y=>p(115)(4),Cin=>p(116)(4),clock=>clock,reset=>reset,s=>p(204)(4),cout=>p(205)(5));
FA_ff_4869:FAff port map(x=>p(114)(5),y=>p(115)(5),Cin=>p(116)(5),clock=>clock,reset=>reset,s=>p(204)(5),cout=>p(205)(6));
FA_ff_4870:FAff port map(x=>p(114)(6),y=>p(115)(6),Cin=>p(116)(6),clock=>clock,reset=>reset,s=>p(204)(6),cout=>p(205)(7));
FA_ff_4871:FAff port map(x=>p(114)(7),y=>p(115)(7),Cin=>p(116)(7),clock=>clock,reset=>reset,s=>p(204)(7),cout=>p(205)(8));
FA_ff_4872:FAff port map(x=>p(114)(8),y=>p(115)(8),Cin=>p(116)(8),clock=>clock,reset=>reset,s=>p(204)(8),cout=>p(205)(9));
FA_ff_4873:FAff port map(x=>p(114)(9),y=>p(115)(9),Cin=>p(116)(9),clock=>clock,reset=>reset,s=>p(204)(9),cout=>p(205)(10));
FA_ff_4874:FAff port map(x=>p(114)(10),y=>p(115)(10),Cin=>p(116)(10),clock=>clock,reset=>reset,s=>p(204)(10),cout=>p(205)(11));
FA_ff_4875:FAff port map(x=>p(114)(11),y=>p(115)(11),Cin=>p(116)(11),clock=>clock,reset=>reset,s=>p(204)(11),cout=>p(205)(12));
FA_ff_4876:FAff port map(x=>p(114)(12),y=>p(115)(12),Cin=>p(116)(12),clock=>clock,reset=>reset,s=>p(204)(12),cout=>p(205)(13));
FA_ff_4877:FAff port map(x=>p(114)(13),y=>p(115)(13),Cin=>p(116)(13),clock=>clock,reset=>reset,s=>p(204)(13),cout=>p(205)(14));
FA_ff_4878:FAff port map(x=>p(114)(14),y=>p(115)(14),Cin=>p(116)(14),clock=>clock,reset=>reset,s=>p(204)(14),cout=>p(205)(15));
FA_ff_4879:FAff port map(x=>p(114)(15),y=>p(115)(15),Cin=>p(116)(15),clock=>clock,reset=>reset,s=>p(204)(15),cout=>p(205)(16));
FA_ff_4880:FAff port map(x=>p(114)(16),y=>p(115)(16),Cin=>p(116)(16),clock=>clock,reset=>reset,s=>p(204)(16),cout=>p(205)(17));
FA_ff_4881:FAff port map(x=>p(114)(17),y=>p(115)(17),Cin=>p(116)(17),clock=>clock,reset=>reset,s=>p(204)(17),cout=>p(205)(18));
FA_ff_4882:FAff port map(x=>p(114)(18),y=>p(115)(18),Cin=>p(116)(18),clock=>clock,reset=>reset,s=>p(204)(18),cout=>p(205)(19));
FA_ff_4883:FAff port map(x=>p(114)(19),y=>p(115)(19),Cin=>p(116)(19),clock=>clock,reset=>reset,s=>p(204)(19),cout=>p(205)(20));
FA_ff_4884:FAff port map(x=>p(114)(20),y=>p(115)(20),Cin=>p(116)(20),clock=>clock,reset=>reset,s=>p(204)(20),cout=>p(205)(21));
FA_ff_4885:FAff port map(x=>p(114)(21),y=>p(115)(21),Cin=>p(116)(21),clock=>clock,reset=>reset,s=>p(204)(21),cout=>p(205)(22));
FA_ff_4886:FAff port map(x=>p(114)(22),y=>p(115)(22),Cin=>p(116)(22),clock=>clock,reset=>reset,s=>p(204)(22),cout=>p(205)(23));
FA_ff_4887:FAff port map(x=>p(114)(23),y=>p(115)(23),Cin=>p(116)(23),clock=>clock,reset=>reset,s=>p(204)(23),cout=>p(205)(24));
FA_ff_4888:FAff port map(x=>p(114)(24),y=>p(115)(24),Cin=>p(116)(24),clock=>clock,reset=>reset,s=>p(204)(24),cout=>p(205)(25));
FA_ff_4889:FAff port map(x=>p(114)(25),y=>p(115)(25),Cin=>p(116)(25),clock=>clock,reset=>reset,s=>p(204)(25),cout=>p(205)(26));
FA_ff_4890:FAff port map(x=>p(114)(26),y=>p(115)(26),Cin=>p(116)(26),clock=>clock,reset=>reset,s=>p(204)(26),cout=>p(205)(27));
FA_ff_4891:FAff port map(x=>p(114)(27),y=>p(115)(27),Cin=>p(116)(27),clock=>clock,reset=>reset,s=>p(204)(27),cout=>p(205)(28));
FA_ff_4892:FAff port map(x=>p(114)(28),y=>p(115)(28),Cin=>p(116)(28),clock=>clock,reset=>reset,s=>p(204)(28),cout=>p(205)(29));
FA_ff_4893:FAff port map(x=>p(114)(29),y=>p(115)(29),Cin=>p(116)(29),clock=>clock,reset=>reset,s=>p(204)(29),cout=>p(205)(30));
FA_ff_4894:FAff port map(x=>p(114)(30),y=>p(115)(30),Cin=>p(116)(30),clock=>clock,reset=>reset,s=>p(204)(30),cout=>p(205)(31));
FA_ff_4895:FAff port map(x=>p(114)(31),y=>p(115)(31),Cin=>p(116)(31),clock=>clock,reset=>reset,s=>p(204)(31),cout=>p(205)(32));
FA_ff_4896:FAff port map(x=>p(114)(32),y=>p(115)(32),Cin=>p(116)(32),clock=>clock,reset=>reset,s=>p(204)(32),cout=>p(205)(33));
FA_ff_4897:FAff port map(x=>p(114)(33),y=>p(115)(33),Cin=>p(116)(33),clock=>clock,reset=>reset,s=>p(204)(33),cout=>p(205)(34));
FA_ff_4898:FAff port map(x=>p(114)(34),y=>p(115)(34),Cin=>p(116)(34),clock=>clock,reset=>reset,s=>p(204)(34),cout=>p(205)(35));
FA_ff_4899:FAff port map(x=>p(114)(35),y=>p(115)(35),Cin=>p(116)(35),clock=>clock,reset=>reset,s=>p(204)(35),cout=>p(205)(36));
FA_ff_4900:FAff port map(x=>p(114)(36),y=>p(115)(36),Cin=>p(116)(36),clock=>clock,reset=>reset,s=>p(204)(36),cout=>p(205)(37));
FA_ff_4901:FAff port map(x=>p(114)(37),y=>p(115)(37),Cin=>p(116)(37),clock=>clock,reset=>reset,s=>p(204)(37),cout=>p(205)(38));
FA_ff_4902:FAff port map(x=>p(114)(38),y=>p(115)(38),Cin=>p(116)(38),clock=>clock,reset=>reset,s=>p(204)(38),cout=>p(205)(39));
FA_ff_4903:FAff port map(x=>p(114)(39),y=>p(115)(39),Cin=>p(116)(39),clock=>clock,reset=>reset,s=>p(204)(39),cout=>p(205)(40));
FA_ff_4904:FAff port map(x=>p(114)(40),y=>p(115)(40),Cin=>p(116)(40),clock=>clock,reset=>reset,s=>p(204)(40),cout=>p(205)(41));
FA_ff_4905:FAff port map(x=>p(114)(41),y=>p(115)(41),Cin=>p(116)(41),clock=>clock,reset=>reset,s=>p(204)(41),cout=>p(205)(42));
FA_ff_4906:FAff port map(x=>p(114)(42),y=>p(115)(42),Cin=>p(116)(42),clock=>clock,reset=>reset,s=>p(204)(42),cout=>p(205)(43));
FA_ff_4907:FAff port map(x=>p(114)(43),y=>p(115)(43),Cin=>p(116)(43),clock=>clock,reset=>reset,s=>p(204)(43),cout=>p(205)(44));
FA_ff_4908:FAff port map(x=>p(114)(44),y=>p(115)(44),Cin=>p(116)(44),clock=>clock,reset=>reset,s=>p(204)(44),cout=>p(205)(45));
FA_ff_4909:FAff port map(x=>p(114)(45),y=>p(115)(45),Cin=>p(116)(45),clock=>clock,reset=>reset,s=>p(204)(45),cout=>p(205)(46));
FA_ff_4910:FAff port map(x=>p(114)(46),y=>p(115)(46),Cin=>p(116)(46),clock=>clock,reset=>reset,s=>p(204)(46),cout=>p(205)(47));
FA_ff_4911:FAff port map(x=>p(114)(47),y=>p(115)(47),Cin=>p(116)(47),clock=>clock,reset=>reset,s=>p(204)(47),cout=>p(205)(48));
FA_ff_4912:FAff port map(x=>p(114)(48),y=>p(115)(48),Cin=>p(116)(48),clock=>clock,reset=>reset,s=>p(204)(48),cout=>p(205)(49));
FA_ff_4913:FAff port map(x=>p(114)(49),y=>p(115)(49),Cin=>p(116)(49),clock=>clock,reset=>reset,s=>p(204)(49),cout=>p(205)(50));
FA_ff_4914:FAff port map(x=>p(114)(50),y=>p(115)(50),Cin=>p(116)(50),clock=>clock,reset=>reset,s=>p(204)(50),cout=>p(205)(51));
FA_ff_4915:FAff port map(x=>p(114)(51),y=>p(115)(51),Cin=>p(116)(51),clock=>clock,reset=>reset,s=>p(204)(51),cout=>p(205)(52));
FA_ff_4916:FAff port map(x=>p(114)(52),y=>p(115)(52),Cin=>p(116)(52),clock=>clock,reset=>reset,s=>p(204)(52),cout=>p(205)(53));
FA_ff_4917:FAff port map(x=>p(114)(53),y=>p(115)(53),Cin=>p(116)(53),clock=>clock,reset=>reset,s=>p(204)(53),cout=>p(205)(54));
FA_ff_4918:FAff port map(x=>p(114)(54),y=>p(115)(54),Cin=>p(116)(54),clock=>clock,reset=>reset,s=>p(204)(54),cout=>p(205)(55));
FA_ff_4919:FAff port map(x=>p(114)(55),y=>p(115)(55),Cin=>p(116)(55),clock=>clock,reset=>reset,s=>p(204)(55),cout=>p(205)(56));
FA_ff_4920:FAff port map(x=>p(114)(56),y=>p(115)(56),Cin=>p(116)(56),clock=>clock,reset=>reset,s=>p(204)(56),cout=>p(205)(57));
FA_ff_4921:FAff port map(x=>p(114)(57),y=>p(115)(57),Cin=>p(116)(57),clock=>clock,reset=>reset,s=>p(204)(57),cout=>p(205)(58));
FA_ff_4922:FAff port map(x=>p(114)(58),y=>p(115)(58),Cin=>p(116)(58),clock=>clock,reset=>reset,s=>p(204)(58),cout=>p(205)(59));
FA_ff_4923:FAff port map(x=>p(114)(59),y=>p(115)(59),Cin=>p(116)(59),clock=>clock,reset=>reset,s=>p(204)(59),cout=>p(205)(60));
FA_ff_4924:FAff port map(x=>p(114)(60),y=>p(115)(60),Cin=>p(116)(60),clock=>clock,reset=>reset,s=>p(204)(60),cout=>p(205)(61));
FA_ff_4925:FAff port map(x=>p(114)(61),y=>p(115)(61),Cin=>p(116)(61),clock=>clock,reset=>reset,s=>p(204)(61),cout=>p(205)(62));
FA_ff_4926:FAff port map(x=>p(114)(62),y=>p(115)(62),Cin=>p(116)(62),clock=>clock,reset=>reset,s=>p(204)(62),cout=>p(205)(63));
FA_ff_4927:FAff port map(x=>p(114)(63),y=>p(115)(63),Cin=>p(116)(63),clock=>clock,reset=>reset,s=>p(204)(63),cout=>p(205)(64));
FA_ff_4928:FAff port map(x=>p(114)(64),y=>p(115)(64),Cin=>p(116)(64),clock=>clock,reset=>reset,s=>p(204)(64),cout=>p(205)(65));
FA_ff_4929:FAff port map(x=>p(114)(65),y=>p(115)(65),Cin=>p(116)(65),clock=>clock,reset=>reset,s=>p(204)(65),cout=>p(205)(66));
FA_ff_4930:FAff port map(x=>p(114)(66),y=>p(115)(66),Cin=>p(116)(66),clock=>clock,reset=>reset,s=>p(204)(66),cout=>p(205)(67));
FA_ff_4931:FAff port map(x=>p(114)(67),y=>p(115)(67),Cin=>p(116)(67),clock=>clock,reset=>reset,s=>p(204)(67),cout=>p(205)(68));
FA_ff_4932:FAff port map(x=>p(114)(68),y=>p(115)(68),Cin=>p(116)(68),clock=>clock,reset=>reset,s=>p(204)(68),cout=>p(205)(69));
FA_ff_4933:FAff port map(x=>p(114)(69),y=>p(115)(69),Cin=>p(116)(69),clock=>clock,reset=>reset,s=>p(204)(69),cout=>p(205)(70));
FA_ff_4934:FAff port map(x=>p(114)(70),y=>p(115)(70),Cin=>p(116)(70),clock=>clock,reset=>reset,s=>p(204)(70),cout=>p(205)(71));
FA_ff_4935:FAff port map(x=>p(114)(71),y=>p(115)(71),Cin=>p(116)(71),clock=>clock,reset=>reset,s=>p(204)(71),cout=>p(205)(72));
FA_ff_4936:FAff port map(x=>p(114)(72),y=>p(115)(72),Cin=>p(116)(72),clock=>clock,reset=>reset,s=>p(204)(72),cout=>p(205)(73));
FA_ff_4937:FAff port map(x=>p(114)(73),y=>p(115)(73),Cin=>p(116)(73),clock=>clock,reset=>reset,s=>p(204)(73),cout=>p(205)(74));
FA_ff_4938:FAff port map(x=>p(114)(74),y=>p(115)(74),Cin=>p(116)(74),clock=>clock,reset=>reset,s=>p(204)(74),cout=>p(205)(75));
FA_ff_4939:FAff port map(x=>p(114)(75),y=>p(115)(75),Cin=>p(116)(75),clock=>clock,reset=>reset,s=>p(204)(75),cout=>p(205)(76));
FA_ff_4940:FAff port map(x=>p(114)(76),y=>p(115)(76),Cin=>p(116)(76),clock=>clock,reset=>reset,s=>p(204)(76),cout=>p(205)(77));
FA_ff_4941:FAff port map(x=>p(114)(77),y=>p(115)(77),Cin=>p(116)(77),clock=>clock,reset=>reset,s=>p(204)(77),cout=>p(205)(78));
FA_ff_4942:FAff port map(x=>p(114)(78),y=>p(115)(78),Cin=>p(116)(78),clock=>clock,reset=>reset,s=>p(204)(78),cout=>p(205)(79));
FA_ff_4943:FAff port map(x=>p(114)(79),y=>p(115)(79),Cin=>p(116)(79),clock=>clock,reset=>reset,s=>p(204)(79),cout=>p(205)(80));
FA_ff_4944:FAff port map(x=>p(114)(80),y=>p(115)(80),Cin=>p(116)(80),clock=>clock,reset=>reset,s=>p(204)(80),cout=>p(205)(81));
FA_ff_4945:FAff port map(x=>p(114)(81),y=>p(115)(81),Cin=>p(116)(81),clock=>clock,reset=>reset,s=>p(204)(81),cout=>p(205)(82));
FA_ff_4946:FAff port map(x=>p(114)(82),y=>p(115)(82),Cin=>p(116)(82),clock=>clock,reset=>reset,s=>p(204)(82),cout=>p(205)(83));
FA_ff_4947:FAff port map(x=>p(114)(83),y=>p(115)(83),Cin=>p(116)(83),clock=>clock,reset=>reset,s=>p(204)(83),cout=>p(205)(84));
FA_ff_4948:FAff port map(x=>p(114)(84),y=>p(115)(84),Cin=>p(116)(84),clock=>clock,reset=>reset,s=>p(204)(84),cout=>p(205)(85));
FA_ff_4949:FAff port map(x=>p(114)(85),y=>p(115)(85),Cin=>p(116)(85),clock=>clock,reset=>reset,s=>p(204)(85),cout=>p(205)(86));
FA_ff_4950:FAff port map(x=>p(114)(86),y=>p(115)(86),Cin=>p(116)(86),clock=>clock,reset=>reset,s=>p(204)(86),cout=>p(205)(87));
FA_ff_4951:FAff port map(x=>p(114)(87),y=>p(115)(87),Cin=>p(116)(87),clock=>clock,reset=>reset,s=>p(204)(87),cout=>p(205)(88));
FA_ff_4952:FAff port map(x=>p(114)(88),y=>p(115)(88),Cin=>p(116)(88),clock=>clock,reset=>reset,s=>p(204)(88),cout=>p(205)(89));
FA_ff_4953:FAff port map(x=>p(114)(89),y=>p(115)(89),Cin=>p(116)(89),clock=>clock,reset=>reset,s=>p(204)(89),cout=>p(205)(90));
FA_ff_4954:FAff port map(x=>p(114)(90),y=>p(115)(90),Cin=>p(116)(90),clock=>clock,reset=>reset,s=>p(204)(90),cout=>p(205)(91));
FA_ff_4955:FAff port map(x=>p(114)(91),y=>p(115)(91),Cin=>p(116)(91),clock=>clock,reset=>reset,s=>p(204)(91),cout=>p(205)(92));
FA_ff_4956:FAff port map(x=>p(114)(92),y=>p(115)(92),Cin=>p(116)(92),clock=>clock,reset=>reset,s=>p(204)(92),cout=>p(205)(93));
FA_ff_4957:FAff port map(x=>p(114)(93),y=>p(115)(93),Cin=>p(116)(93),clock=>clock,reset=>reset,s=>p(204)(93),cout=>p(205)(94));
FA_ff_4958:FAff port map(x=>p(114)(94),y=>p(115)(94),Cin=>p(116)(94),clock=>clock,reset=>reset,s=>p(204)(94),cout=>p(205)(95));
FA_ff_4959:FAff port map(x=>p(114)(95),y=>p(115)(95),Cin=>p(116)(95),clock=>clock,reset=>reset,s=>p(204)(95),cout=>p(205)(96));
FA_ff_4960:FAff port map(x=>p(114)(96),y=>p(115)(96),Cin=>p(116)(96),clock=>clock,reset=>reset,s=>p(204)(96),cout=>p(205)(97));
FA_ff_4961:FAff port map(x=>p(114)(97),y=>p(115)(97),Cin=>p(116)(97),clock=>clock,reset=>reset,s=>p(204)(97),cout=>p(205)(98));
FA_ff_4962:FAff port map(x=>p(114)(98),y=>p(115)(98),Cin=>p(116)(98),clock=>clock,reset=>reset,s=>p(204)(98),cout=>p(205)(99));
FA_ff_4963:FAff port map(x=>p(114)(99),y=>p(115)(99),Cin=>p(116)(99),clock=>clock,reset=>reset,s=>p(204)(99),cout=>p(205)(100));
FA_ff_4964:FAff port map(x=>p(114)(100),y=>p(115)(100),Cin=>p(116)(100),clock=>clock,reset=>reset,s=>p(204)(100),cout=>p(205)(101));
FA_ff_4965:FAff port map(x=>p(114)(101),y=>p(115)(101),Cin=>p(116)(101),clock=>clock,reset=>reset,s=>p(204)(101),cout=>p(205)(102));
FA_ff_4966:FAff port map(x=>p(114)(102),y=>p(115)(102),Cin=>p(116)(102),clock=>clock,reset=>reset,s=>p(204)(102),cout=>p(205)(103));
FA_ff_4967:FAff port map(x=>p(114)(103),y=>p(115)(103),Cin=>p(116)(103),clock=>clock,reset=>reset,s=>p(204)(103),cout=>p(205)(104));
FA_ff_4968:FAff port map(x=>p(114)(104),y=>p(115)(104),Cin=>p(116)(104),clock=>clock,reset=>reset,s=>p(204)(104),cout=>p(205)(105));
FA_ff_4969:FAff port map(x=>p(114)(105),y=>p(115)(105),Cin=>p(116)(105),clock=>clock,reset=>reset,s=>p(204)(105),cout=>p(205)(106));
FA_ff_4970:FAff port map(x=>p(114)(106),y=>p(115)(106),Cin=>p(116)(106),clock=>clock,reset=>reset,s=>p(204)(106),cout=>p(205)(107));
FA_ff_4971:FAff port map(x=>p(114)(107),y=>p(115)(107),Cin=>p(116)(107),clock=>clock,reset=>reset,s=>p(204)(107),cout=>p(205)(108));
FA_ff_4972:FAff port map(x=>p(114)(108),y=>p(115)(108),Cin=>p(116)(108),clock=>clock,reset=>reset,s=>p(204)(108),cout=>p(205)(109));
FA_ff_4973:FAff port map(x=>p(114)(109),y=>p(115)(109),Cin=>p(116)(109),clock=>clock,reset=>reset,s=>p(204)(109),cout=>p(205)(110));
FA_ff_4974:FAff port map(x=>p(114)(110),y=>p(115)(110),Cin=>p(116)(110),clock=>clock,reset=>reset,s=>p(204)(110),cout=>p(205)(111));
FA_ff_4975:FAff port map(x=>p(114)(111),y=>p(115)(111),Cin=>p(116)(111),clock=>clock,reset=>reset,s=>p(204)(111),cout=>p(205)(112));
FA_ff_4976:FAff port map(x=>p(114)(112),y=>p(115)(112),Cin=>p(116)(112),clock=>clock,reset=>reset,s=>p(204)(112),cout=>p(205)(113));
FA_ff_4977:FAff port map(x=>p(114)(113),y=>p(115)(113),Cin=>p(116)(113),clock=>clock,reset=>reset,s=>p(204)(113),cout=>p(205)(114));
FA_ff_4978:FAff port map(x=>p(114)(114),y=>p(115)(114),Cin=>p(116)(114),clock=>clock,reset=>reset,s=>p(204)(114),cout=>p(205)(115));
FA_ff_4979:FAff port map(x=>p(114)(115),y=>p(115)(115),Cin=>p(116)(115),clock=>clock,reset=>reset,s=>p(204)(115),cout=>p(205)(116));
FA_ff_4980:FAff port map(x=>p(114)(116),y=>p(115)(116),Cin=>p(116)(116),clock=>clock,reset=>reset,s=>p(204)(116),cout=>p(205)(117));
FA_ff_4981:FAff port map(x=>p(114)(117),y=>p(115)(117),Cin=>p(116)(117),clock=>clock,reset=>reset,s=>p(204)(117),cout=>p(205)(118));
FA_ff_4982:FAff port map(x=>p(114)(118),y=>p(115)(118),Cin=>p(116)(118),clock=>clock,reset=>reset,s=>p(204)(118),cout=>p(205)(119));
FA_ff_4983:FAff port map(x=>p(114)(119),y=>p(115)(119),Cin=>p(116)(119),clock=>clock,reset=>reset,s=>p(204)(119),cout=>p(205)(120));
FA_ff_4984:FAff port map(x=>p(114)(120),y=>p(115)(120),Cin=>p(116)(120),clock=>clock,reset=>reset,s=>p(204)(120),cout=>p(205)(121));
FA_ff_4985:FAff port map(x=>p(114)(121),y=>p(115)(121),Cin=>p(116)(121),clock=>clock,reset=>reset,s=>p(204)(121),cout=>p(205)(122));
FA_ff_4986:FAff port map(x=>p(114)(122),y=>p(115)(122),Cin=>p(116)(122),clock=>clock,reset=>reset,s=>p(204)(122),cout=>p(205)(123));
FA_ff_4987:FAff port map(x=>p(114)(123),y=>p(115)(123),Cin=>p(116)(123),clock=>clock,reset=>reset,s=>p(204)(123),cout=>p(205)(124));
FA_ff_4988:FAff port map(x=>p(114)(124),y=>p(115)(124),Cin=>p(116)(124),clock=>clock,reset=>reset,s=>p(204)(124),cout=>p(205)(125));
FA_ff_4989:FAff port map(x=>p(114)(125),y=>p(115)(125),Cin=>p(116)(125),clock=>clock,reset=>reset,s=>p(204)(125),cout=>p(205)(126));
FA_ff_4990:FAff port map(x=>p(114)(126),y=>p(115)(126),Cin=>p(116)(126),clock=>clock,reset=>reset,s=>p(204)(126),cout=>p(205)(127));
FA_ff_4991:FAff port map(x=>p(114)(127),y=>p(115)(127),Cin=>p(116)(127),clock=>clock,reset=>reset,s=>p(204)(127),cout=>p(205)(128));
FA_ff_4992:FAff port map(x=>p(117)(0),y=>p(118)(0),Cin=>p(119)(0),clock=>clock,reset=>reset,s=>p(206)(0),cout=>p(207)(1));
FA_ff_4993:FAff port map(x=>p(117)(1),y=>p(118)(1),Cin=>p(119)(1),clock=>clock,reset=>reset,s=>p(206)(1),cout=>p(207)(2));
FA_ff_4994:FAff port map(x=>p(117)(2),y=>p(118)(2),Cin=>p(119)(2),clock=>clock,reset=>reset,s=>p(206)(2),cout=>p(207)(3));
FA_ff_4995:FAff port map(x=>p(117)(3),y=>p(118)(3),Cin=>p(119)(3),clock=>clock,reset=>reset,s=>p(206)(3),cout=>p(207)(4));
FA_ff_4996:FAff port map(x=>p(117)(4),y=>p(118)(4),Cin=>p(119)(4),clock=>clock,reset=>reset,s=>p(206)(4),cout=>p(207)(5));
FA_ff_4997:FAff port map(x=>p(117)(5),y=>p(118)(5),Cin=>p(119)(5),clock=>clock,reset=>reset,s=>p(206)(5),cout=>p(207)(6));
FA_ff_4998:FAff port map(x=>p(117)(6),y=>p(118)(6),Cin=>p(119)(6),clock=>clock,reset=>reset,s=>p(206)(6),cout=>p(207)(7));
FA_ff_4999:FAff port map(x=>p(117)(7),y=>p(118)(7),Cin=>p(119)(7),clock=>clock,reset=>reset,s=>p(206)(7),cout=>p(207)(8));
FA_ff_5000:FAff port map(x=>p(117)(8),y=>p(118)(8),Cin=>p(119)(8),clock=>clock,reset=>reset,s=>p(206)(8),cout=>p(207)(9));
FA_ff_5001:FAff port map(x=>p(117)(9),y=>p(118)(9),Cin=>p(119)(9),clock=>clock,reset=>reset,s=>p(206)(9),cout=>p(207)(10));
FA_ff_5002:FAff port map(x=>p(117)(10),y=>p(118)(10),Cin=>p(119)(10),clock=>clock,reset=>reset,s=>p(206)(10),cout=>p(207)(11));
FA_ff_5003:FAff port map(x=>p(117)(11),y=>p(118)(11),Cin=>p(119)(11),clock=>clock,reset=>reset,s=>p(206)(11),cout=>p(207)(12));
FA_ff_5004:FAff port map(x=>p(117)(12),y=>p(118)(12),Cin=>p(119)(12),clock=>clock,reset=>reset,s=>p(206)(12),cout=>p(207)(13));
FA_ff_5005:FAff port map(x=>p(117)(13),y=>p(118)(13),Cin=>p(119)(13),clock=>clock,reset=>reset,s=>p(206)(13),cout=>p(207)(14));
FA_ff_5006:FAff port map(x=>p(117)(14),y=>p(118)(14),Cin=>p(119)(14),clock=>clock,reset=>reset,s=>p(206)(14),cout=>p(207)(15));
FA_ff_5007:FAff port map(x=>p(117)(15),y=>p(118)(15),Cin=>p(119)(15),clock=>clock,reset=>reset,s=>p(206)(15),cout=>p(207)(16));
FA_ff_5008:FAff port map(x=>p(117)(16),y=>p(118)(16),Cin=>p(119)(16),clock=>clock,reset=>reset,s=>p(206)(16),cout=>p(207)(17));
FA_ff_5009:FAff port map(x=>p(117)(17),y=>p(118)(17),Cin=>p(119)(17),clock=>clock,reset=>reset,s=>p(206)(17),cout=>p(207)(18));
FA_ff_5010:FAff port map(x=>p(117)(18),y=>p(118)(18),Cin=>p(119)(18),clock=>clock,reset=>reset,s=>p(206)(18),cout=>p(207)(19));
FA_ff_5011:FAff port map(x=>p(117)(19),y=>p(118)(19),Cin=>p(119)(19),clock=>clock,reset=>reset,s=>p(206)(19),cout=>p(207)(20));
FA_ff_5012:FAff port map(x=>p(117)(20),y=>p(118)(20),Cin=>p(119)(20),clock=>clock,reset=>reset,s=>p(206)(20),cout=>p(207)(21));
FA_ff_5013:FAff port map(x=>p(117)(21),y=>p(118)(21),Cin=>p(119)(21),clock=>clock,reset=>reset,s=>p(206)(21),cout=>p(207)(22));
FA_ff_5014:FAff port map(x=>p(117)(22),y=>p(118)(22),Cin=>p(119)(22),clock=>clock,reset=>reset,s=>p(206)(22),cout=>p(207)(23));
FA_ff_5015:FAff port map(x=>p(117)(23),y=>p(118)(23),Cin=>p(119)(23),clock=>clock,reset=>reset,s=>p(206)(23),cout=>p(207)(24));
FA_ff_5016:FAff port map(x=>p(117)(24),y=>p(118)(24),Cin=>p(119)(24),clock=>clock,reset=>reset,s=>p(206)(24),cout=>p(207)(25));
FA_ff_5017:FAff port map(x=>p(117)(25),y=>p(118)(25),Cin=>p(119)(25),clock=>clock,reset=>reset,s=>p(206)(25),cout=>p(207)(26));
FA_ff_5018:FAff port map(x=>p(117)(26),y=>p(118)(26),Cin=>p(119)(26),clock=>clock,reset=>reset,s=>p(206)(26),cout=>p(207)(27));
FA_ff_5019:FAff port map(x=>p(117)(27),y=>p(118)(27),Cin=>p(119)(27),clock=>clock,reset=>reset,s=>p(206)(27),cout=>p(207)(28));
FA_ff_5020:FAff port map(x=>p(117)(28),y=>p(118)(28),Cin=>p(119)(28),clock=>clock,reset=>reset,s=>p(206)(28),cout=>p(207)(29));
FA_ff_5021:FAff port map(x=>p(117)(29),y=>p(118)(29),Cin=>p(119)(29),clock=>clock,reset=>reset,s=>p(206)(29),cout=>p(207)(30));
FA_ff_5022:FAff port map(x=>p(117)(30),y=>p(118)(30),Cin=>p(119)(30),clock=>clock,reset=>reset,s=>p(206)(30),cout=>p(207)(31));
FA_ff_5023:FAff port map(x=>p(117)(31),y=>p(118)(31),Cin=>p(119)(31),clock=>clock,reset=>reset,s=>p(206)(31),cout=>p(207)(32));
FA_ff_5024:FAff port map(x=>p(117)(32),y=>p(118)(32),Cin=>p(119)(32),clock=>clock,reset=>reset,s=>p(206)(32),cout=>p(207)(33));
FA_ff_5025:FAff port map(x=>p(117)(33),y=>p(118)(33),Cin=>p(119)(33),clock=>clock,reset=>reset,s=>p(206)(33),cout=>p(207)(34));
FA_ff_5026:FAff port map(x=>p(117)(34),y=>p(118)(34),Cin=>p(119)(34),clock=>clock,reset=>reset,s=>p(206)(34),cout=>p(207)(35));
FA_ff_5027:FAff port map(x=>p(117)(35),y=>p(118)(35),Cin=>p(119)(35),clock=>clock,reset=>reset,s=>p(206)(35),cout=>p(207)(36));
FA_ff_5028:FAff port map(x=>p(117)(36),y=>p(118)(36),Cin=>p(119)(36),clock=>clock,reset=>reset,s=>p(206)(36),cout=>p(207)(37));
FA_ff_5029:FAff port map(x=>p(117)(37),y=>p(118)(37),Cin=>p(119)(37),clock=>clock,reset=>reset,s=>p(206)(37),cout=>p(207)(38));
FA_ff_5030:FAff port map(x=>p(117)(38),y=>p(118)(38),Cin=>p(119)(38),clock=>clock,reset=>reset,s=>p(206)(38),cout=>p(207)(39));
FA_ff_5031:FAff port map(x=>p(117)(39),y=>p(118)(39),Cin=>p(119)(39),clock=>clock,reset=>reset,s=>p(206)(39),cout=>p(207)(40));
FA_ff_5032:FAff port map(x=>p(117)(40),y=>p(118)(40),Cin=>p(119)(40),clock=>clock,reset=>reset,s=>p(206)(40),cout=>p(207)(41));
FA_ff_5033:FAff port map(x=>p(117)(41),y=>p(118)(41),Cin=>p(119)(41),clock=>clock,reset=>reset,s=>p(206)(41),cout=>p(207)(42));
FA_ff_5034:FAff port map(x=>p(117)(42),y=>p(118)(42),Cin=>p(119)(42),clock=>clock,reset=>reset,s=>p(206)(42),cout=>p(207)(43));
FA_ff_5035:FAff port map(x=>p(117)(43),y=>p(118)(43),Cin=>p(119)(43),clock=>clock,reset=>reset,s=>p(206)(43),cout=>p(207)(44));
FA_ff_5036:FAff port map(x=>p(117)(44),y=>p(118)(44),Cin=>p(119)(44),clock=>clock,reset=>reset,s=>p(206)(44),cout=>p(207)(45));
FA_ff_5037:FAff port map(x=>p(117)(45),y=>p(118)(45),Cin=>p(119)(45),clock=>clock,reset=>reset,s=>p(206)(45),cout=>p(207)(46));
FA_ff_5038:FAff port map(x=>p(117)(46),y=>p(118)(46),Cin=>p(119)(46),clock=>clock,reset=>reset,s=>p(206)(46),cout=>p(207)(47));
FA_ff_5039:FAff port map(x=>p(117)(47),y=>p(118)(47),Cin=>p(119)(47),clock=>clock,reset=>reset,s=>p(206)(47),cout=>p(207)(48));
FA_ff_5040:FAff port map(x=>p(117)(48),y=>p(118)(48),Cin=>p(119)(48),clock=>clock,reset=>reset,s=>p(206)(48),cout=>p(207)(49));
FA_ff_5041:FAff port map(x=>p(117)(49),y=>p(118)(49),Cin=>p(119)(49),clock=>clock,reset=>reset,s=>p(206)(49),cout=>p(207)(50));
FA_ff_5042:FAff port map(x=>p(117)(50),y=>p(118)(50),Cin=>p(119)(50),clock=>clock,reset=>reset,s=>p(206)(50),cout=>p(207)(51));
FA_ff_5043:FAff port map(x=>p(117)(51),y=>p(118)(51),Cin=>p(119)(51),clock=>clock,reset=>reset,s=>p(206)(51),cout=>p(207)(52));
FA_ff_5044:FAff port map(x=>p(117)(52),y=>p(118)(52),Cin=>p(119)(52),clock=>clock,reset=>reset,s=>p(206)(52),cout=>p(207)(53));
FA_ff_5045:FAff port map(x=>p(117)(53),y=>p(118)(53),Cin=>p(119)(53),clock=>clock,reset=>reset,s=>p(206)(53),cout=>p(207)(54));
FA_ff_5046:FAff port map(x=>p(117)(54),y=>p(118)(54),Cin=>p(119)(54),clock=>clock,reset=>reset,s=>p(206)(54),cout=>p(207)(55));
FA_ff_5047:FAff port map(x=>p(117)(55),y=>p(118)(55),Cin=>p(119)(55),clock=>clock,reset=>reset,s=>p(206)(55),cout=>p(207)(56));
FA_ff_5048:FAff port map(x=>p(117)(56),y=>p(118)(56),Cin=>p(119)(56),clock=>clock,reset=>reset,s=>p(206)(56),cout=>p(207)(57));
FA_ff_5049:FAff port map(x=>p(117)(57),y=>p(118)(57),Cin=>p(119)(57),clock=>clock,reset=>reset,s=>p(206)(57),cout=>p(207)(58));
FA_ff_5050:FAff port map(x=>p(117)(58),y=>p(118)(58),Cin=>p(119)(58),clock=>clock,reset=>reset,s=>p(206)(58),cout=>p(207)(59));
FA_ff_5051:FAff port map(x=>p(117)(59),y=>p(118)(59),Cin=>p(119)(59),clock=>clock,reset=>reset,s=>p(206)(59),cout=>p(207)(60));
FA_ff_5052:FAff port map(x=>p(117)(60),y=>p(118)(60),Cin=>p(119)(60),clock=>clock,reset=>reset,s=>p(206)(60),cout=>p(207)(61));
FA_ff_5053:FAff port map(x=>p(117)(61),y=>p(118)(61),Cin=>p(119)(61),clock=>clock,reset=>reset,s=>p(206)(61),cout=>p(207)(62));
FA_ff_5054:FAff port map(x=>p(117)(62),y=>p(118)(62),Cin=>p(119)(62),clock=>clock,reset=>reset,s=>p(206)(62),cout=>p(207)(63));
FA_ff_5055:FAff port map(x=>p(117)(63),y=>p(118)(63),Cin=>p(119)(63),clock=>clock,reset=>reset,s=>p(206)(63),cout=>p(207)(64));
FA_ff_5056:FAff port map(x=>p(117)(64),y=>p(118)(64),Cin=>p(119)(64),clock=>clock,reset=>reset,s=>p(206)(64),cout=>p(207)(65));
FA_ff_5057:FAff port map(x=>p(117)(65),y=>p(118)(65),Cin=>p(119)(65),clock=>clock,reset=>reset,s=>p(206)(65),cout=>p(207)(66));
FA_ff_5058:FAff port map(x=>p(117)(66),y=>p(118)(66),Cin=>p(119)(66),clock=>clock,reset=>reset,s=>p(206)(66),cout=>p(207)(67));
FA_ff_5059:FAff port map(x=>p(117)(67),y=>p(118)(67),Cin=>p(119)(67),clock=>clock,reset=>reset,s=>p(206)(67),cout=>p(207)(68));
FA_ff_5060:FAff port map(x=>p(117)(68),y=>p(118)(68),Cin=>p(119)(68),clock=>clock,reset=>reset,s=>p(206)(68),cout=>p(207)(69));
FA_ff_5061:FAff port map(x=>p(117)(69),y=>p(118)(69),Cin=>p(119)(69),clock=>clock,reset=>reset,s=>p(206)(69),cout=>p(207)(70));
FA_ff_5062:FAff port map(x=>p(117)(70),y=>p(118)(70),Cin=>p(119)(70),clock=>clock,reset=>reset,s=>p(206)(70),cout=>p(207)(71));
FA_ff_5063:FAff port map(x=>p(117)(71),y=>p(118)(71),Cin=>p(119)(71),clock=>clock,reset=>reset,s=>p(206)(71),cout=>p(207)(72));
FA_ff_5064:FAff port map(x=>p(117)(72),y=>p(118)(72),Cin=>p(119)(72),clock=>clock,reset=>reset,s=>p(206)(72),cout=>p(207)(73));
FA_ff_5065:FAff port map(x=>p(117)(73),y=>p(118)(73),Cin=>p(119)(73),clock=>clock,reset=>reset,s=>p(206)(73),cout=>p(207)(74));
FA_ff_5066:FAff port map(x=>p(117)(74),y=>p(118)(74),Cin=>p(119)(74),clock=>clock,reset=>reset,s=>p(206)(74),cout=>p(207)(75));
FA_ff_5067:FAff port map(x=>p(117)(75),y=>p(118)(75),Cin=>p(119)(75),clock=>clock,reset=>reset,s=>p(206)(75),cout=>p(207)(76));
FA_ff_5068:FAff port map(x=>p(117)(76),y=>p(118)(76),Cin=>p(119)(76),clock=>clock,reset=>reset,s=>p(206)(76),cout=>p(207)(77));
FA_ff_5069:FAff port map(x=>p(117)(77),y=>p(118)(77),Cin=>p(119)(77),clock=>clock,reset=>reset,s=>p(206)(77),cout=>p(207)(78));
FA_ff_5070:FAff port map(x=>p(117)(78),y=>p(118)(78),Cin=>p(119)(78),clock=>clock,reset=>reset,s=>p(206)(78),cout=>p(207)(79));
FA_ff_5071:FAff port map(x=>p(117)(79),y=>p(118)(79),Cin=>p(119)(79),clock=>clock,reset=>reset,s=>p(206)(79),cout=>p(207)(80));
FA_ff_5072:FAff port map(x=>p(117)(80),y=>p(118)(80),Cin=>p(119)(80),clock=>clock,reset=>reset,s=>p(206)(80),cout=>p(207)(81));
FA_ff_5073:FAff port map(x=>p(117)(81),y=>p(118)(81),Cin=>p(119)(81),clock=>clock,reset=>reset,s=>p(206)(81),cout=>p(207)(82));
FA_ff_5074:FAff port map(x=>p(117)(82),y=>p(118)(82),Cin=>p(119)(82),clock=>clock,reset=>reset,s=>p(206)(82),cout=>p(207)(83));
FA_ff_5075:FAff port map(x=>p(117)(83),y=>p(118)(83),Cin=>p(119)(83),clock=>clock,reset=>reset,s=>p(206)(83),cout=>p(207)(84));
FA_ff_5076:FAff port map(x=>p(117)(84),y=>p(118)(84),Cin=>p(119)(84),clock=>clock,reset=>reset,s=>p(206)(84),cout=>p(207)(85));
FA_ff_5077:FAff port map(x=>p(117)(85),y=>p(118)(85),Cin=>p(119)(85),clock=>clock,reset=>reset,s=>p(206)(85),cout=>p(207)(86));
FA_ff_5078:FAff port map(x=>p(117)(86),y=>p(118)(86),Cin=>p(119)(86),clock=>clock,reset=>reset,s=>p(206)(86),cout=>p(207)(87));
FA_ff_5079:FAff port map(x=>p(117)(87),y=>p(118)(87),Cin=>p(119)(87),clock=>clock,reset=>reset,s=>p(206)(87),cout=>p(207)(88));
FA_ff_5080:FAff port map(x=>p(117)(88),y=>p(118)(88),Cin=>p(119)(88),clock=>clock,reset=>reset,s=>p(206)(88),cout=>p(207)(89));
FA_ff_5081:FAff port map(x=>p(117)(89),y=>p(118)(89),Cin=>p(119)(89),clock=>clock,reset=>reset,s=>p(206)(89),cout=>p(207)(90));
FA_ff_5082:FAff port map(x=>p(117)(90),y=>p(118)(90),Cin=>p(119)(90),clock=>clock,reset=>reset,s=>p(206)(90),cout=>p(207)(91));
FA_ff_5083:FAff port map(x=>p(117)(91),y=>p(118)(91),Cin=>p(119)(91),clock=>clock,reset=>reset,s=>p(206)(91),cout=>p(207)(92));
FA_ff_5084:FAff port map(x=>p(117)(92),y=>p(118)(92),Cin=>p(119)(92),clock=>clock,reset=>reset,s=>p(206)(92),cout=>p(207)(93));
FA_ff_5085:FAff port map(x=>p(117)(93),y=>p(118)(93),Cin=>p(119)(93),clock=>clock,reset=>reset,s=>p(206)(93),cout=>p(207)(94));
FA_ff_5086:FAff port map(x=>p(117)(94),y=>p(118)(94),Cin=>p(119)(94),clock=>clock,reset=>reset,s=>p(206)(94),cout=>p(207)(95));
FA_ff_5087:FAff port map(x=>p(117)(95),y=>p(118)(95),Cin=>p(119)(95),clock=>clock,reset=>reset,s=>p(206)(95),cout=>p(207)(96));
FA_ff_5088:FAff port map(x=>p(117)(96),y=>p(118)(96),Cin=>p(119)(96),clock=>clock,reset=>reset,s=>p(206)(96),cout=>p(207)(97));
FA_ff_5089:FAff port map(x=>p(117)(97),y=>p(118)(97),Cin=>p(119)(97),clock=>clock,reset=>reset,s=>p(206)(97),cout=>p(207)(98));
FA_ff_5090:FAff port map(x=>p(117)(98),y=>p(118)(98),Cin=>p(119)(98),clock=>clock,reset=>reset,s=>p(206)(98),cout=>p(207)(99));
FA_ff_5091:FAff port map(x=>p(117)(99),y=>p(118)(99),Cin=>p(119)(99),clock=>clock,reset=>reset,s=>p(206)(99),cout=>p(207)(100));
FA_ff_5092:FAff port map(x=>p(117)(100),y=>p(118)(100),Cin=>p(119)(100),clock=>clock,reset=>reset,s=>p(206)(100),cout=>p(207)(101));
FA_ff_5093:FAff port map(x=>p(117)(101),y=>p(118)(101),Cin=>p(119)(101),clock=>clock,reset=>reset,s=>p(206)(101),cout=>p(207)(102));
FA_ff_5094:FAff port map(x=>p(117)(102),y=>p(118)(102),Cin=>p(119)(102),clock=>clock,reset=>reset,s=>p(206)(102),cout=>p(207)(103));
FA_ff_5095:FAff port map(x=>p(117)(103),y=>p(118)(103),Cin=>p(119)(103),clock=>clock,reset=>reset,s=>p(206)(103),cout=>p(207)(104));
FA_ff_5096:FAff port map(x=>p(117)(104),y=>p(118)(104),Cin=>p(119)(104),clock=>clock,reset=>reset,s=>p(206)(104),cout=>p(207)(105));
FA_ff_5097:FAff port map(x=>p(117)(105),y=>p(118)(105),Cin=>p(119)(105),clock=>clock,reset=>reset,s=>p(206)(105),cout=>p(207)(106));
FA_ff_5098:FAff port map(x=>p(117)(106),y=>p(118)(106),Cin=>p(119)(106),clock=>clock,reset=>reset,s=>p(206)(106),cout=>p(207)(107));
FA_ff_5099:FAff port map(x=>p(117)(107),y=>p(118)(107),Cin=>p(119)(107),clock=>clock,reset=>reset,s=>p(206)(107),cout=>p(207)(108));
FA_ff_5100:FAff port map(x=>p(117)(108),y=>p(118)(108),Cin=>p(119)(108),clock=>clock,reset=>reset,s=>p(206)(108),cout=>p(207)(109));
FA_ff_5101:FAff port map(x=>p(117)(109),y=>p(118)(109),Cin=>p(119)(109),clock=>clock,reset=>reset,s=>p(206)(109),cout=>p(207)(110));
FA_ff_5102:FAff port map(x=>p(117)(110),y=>p(118)(110),Cin=>p(119)(110),clock=>clock,reset=>reset,s=>p(206)(110),cout=>p(207)(111));
FA_ff_5103:FAff port map(x=>p(117)(111),y=>p(118)(111),Cin=>p(119)(111),clock=>clock,reset=>reset,s=>p(206)(111),cout=>p(207)(112));
FA_ff_5104:FAff port map(x=>p(117)(112),y=>p(118)(112),Cin=>p(119)(112),clock=>clock,reset=>reset,s=>p(206)(112),cout=>p(207)(113));
FA_ff_5105:FAff port map(x=>p(117)(113),y=>p(118)(113),Cin=>p(119)(113),clock=>clock,reset=>reset,s=>p(206)(113),cout=>p(207)(114));
FA_ff_5106:FAff port map(x=>p(117)(114),y=>p(118)(114),Cin=>p(119)(114),clock=>clock,reset=>reset,s=>p(206)(114),cout=>p(207)(115));
FA_ff_5107:FAff port map(x=>p(117)(115),y=>p(118)(115),Cin=>p(119)(115),clock=>clock,reset=>reset,s=>p(206)(115),cout=>p(207)(116));
FA_ff_5108:FAff port map(x=>p(117)(116),y=>p(118)(116),Cin=>p(119)(116),clock=>clock,reset=>reset,s=>p(206)(116),cout=>p(207)(117));
FA_ff_5109:FAff port map(x=>p(117)(117),y=>p(118)(117),Cin=>p(119)(117),clock=>clock,reset=>reset,s=>p(206)(117),cout=>p(207)(118));
FA_ff_5110:FAff port map(x=>p(117)(118),y=>p(118)(118),Cin=>p(119)(118),clock=>clock,reset=>reset,s=>p(206)(118),cout=>p(207)(119));
FA_ff_5111:FAff port map(x=>p(117)(119),y=>p(118)(119),Cin=>p(119)(119),clock=>clock,reset=>reset,s=>p(206)(119),cout=>p(207)(120));
FA_ff_5112:FAff port map(x=>p(117)(120),y=>p(118)(120),Cin=>p(119)(120),clock=>clock,reset=>reset,s=>p(206)(120),cout=>p(207)(121));
FA_ff_5113:FAff port map(x=>p(117)(121),y=>p(118)(121),Cin=>p(119)(121),clock=>clock,reset=>reset,s=>p(206)(121),cout=>p(207)(122));
FA_ff_5114:FAff port map(x=>p(117)(122),y=>p(118)(122),Cin=>p(119)(122),clock=>clock,reset=>reset,s=>p(206)(122),cout=>p(207)(123));
FA_ff_5115:FAff port map(x=>p(117)(123),y=>p(118)(123),Cin=>p(119)(123),clock=>clock,reset=>reset,s=>p(206)(123),cout=>p(207)(124));
FA_ff_5116:FAff port map(x=>p(117)(124),y=>p(118)(124),Cin=>p(119)(124),clock=>clock,reset=>reset,s=>p(206)(124),cout=>p(207)(125));
FA_ff_5117:FAff port map(x=>p(117)(125),y=>p(118)(125),Cin=>p(119)(125),clock=>clock,reset=>reset,s=>p(206)(125),cout=>p(207)(126));
FA_ff_5118:FAff port map(x=>p(117)(126),y=>p(118)(126),Cin=>p(119)(126),clock=>clock,reset=>reset,s=>p(206)(126),cout=>p(207)(127));
FA_ff_5119:FAff port map(x=>p(117)(127),y=>p(118)(127),Cin=>p(119)(127),clock=>clock,reset=>reset,s=>p(206)(127),cout=>p(207)(128));
FA_ff_5120:FAff port map(x=>p(120)(0),y=>p(121)(0),Cin=>p(122)(0),clock=>clock,reset=>reset,s=>p(208)(0),cout=>p(209)(1));
FA_ff_5121:FAff port map(x=>p(120)(1),y=>p(121)(1),Cin=>p(122)(1),clock=>clock,reset=>reset,s=>p(208)(1),cout=>p(209)(2));
FA_ff_5122:FAff port map(x=>p(120)(2),y=>p(121)(2),Cin=>p(122)(2),clock=>clock,reset=>reset,s=>p(208)(2),cout=>p(209)(3));
FA_ff_5123:FAff port map(x=>p(120)(3),y=>p(121)(3),Cin=>p(122)(3),clock=>clock,reset=>reset,s=>p(208)(3),cout=>p(209)(4));
FA_ff_5124:FAff port map(x=>p(120)(4),y=>p(121)(4),Cin=>p(122)(4),clock=>clock,reset=>reset,s=>p(208)(4),cout=>p(209)(5));
FA_ff_5125:FAff port map(x=>p(120)(5),y=>p(121)(5),Cin=>p(122)(5),clock=>clock,reset=>reset,s=>p(208)(5),cout=>p(209)(6));
FA_ff_5126:FAff port map(x=>p(120)(6),y=>p(121)(6),Cin=>p(122)(6),clock=>clock,reset=>reset,s=>p(208)(6),cout=>p(209)(7));
FA_ff_5127:FAff port map(x=>p(120)(7),y=>p(121)(7),Cin=>p(122)(7),clock=>clock,reset=>reset,s=>p(208)(7),cout=>p(209)(8));
FA_ff_5128:FAff port map(x=>p(120)(8),y=>p(121)(8),Cin=>p(122)(8),clock=>clock,reset=>reset,s=>p(208)(8),cout=>p(209)(9));
FA_ff_5129:FAff port map(x=>p(120)(9),y=>p(121)(9),Cin=>p(122)(9),clock=>clock,reset=>reset,s=>p(208)(9),cout=>p(209)(10));
FA_ff_5130:FAff port map(x=>p(120)(10),y=>p(121)(10),Cin=>p(122)(10),clock=>clock,reset=>reset,s=>p(208)(10),cout=>p(209)(11));
FA_ff_5131:FAff port map(x=>p(120)(11),y=>p(121)(11),Cin=>p(122)(11),clock=>clock,reset=>reset,s=>p(208)(11),cout=>p(209)(12));
FA_ff_5132:FAff port map(x=>p(120)(12),y=>p(121)(12),Cin=>p(122)(12),clock=>clock,reset=>reset,s=>p(208)(12),cout=>p(209)(13));
FA_ff_5133:FAff port map(x=>p(120)(13),y=>p(121)(13),Cin=>p(122)(13),clock=>clock,reset=>reset,s=>p(208)(13),cout=>p(209)(14));
FA_ff_5134:FAff port map(x=>p(120)(14),y=>p(121)(14),Cin=>p(122)(14),clock=>clock,reset=>reset,s=>p(208)(14),cout=>p(209)(15));
FA_ff_5135:FAff port map(x=>p(120)(15),y=>p(121)(15),Cin=>p(122)(15),clock=>clock,reset=>reset,s=>p(208)(15),cout=>p(209)(16));
FA_ff_5136:FAff port map(x=>p(120)(16),y=>p(121)(16),Cin=>p(122)(16),clock=>clock,reset=>reset,s=>p(208)(16),cout=>p(209)(17));
FA_ff_5137:FAff port map(x=>p(120)(17),y=>p(121)(17),Cin=>p(122)(17),clock=>clock,reset=>reset,s=>p(208)(17),cout=>p(209)(18));
FA_ff_5138:FAff port map(x=>p(120)(18),y=>p(121)(18),Cin=>p(122)(18),clock=>clock,reset=>reset,s=>p(208)(18),cout=>p(209)(19));
FA_ff_5139:FAff port map(x=>p(120)(19),y=>p(121)(19),Cin=>p(122)(19),clock=>clock,reset=>reset,s=>p(208)(19),cout=>p(209)(20));
FA_ff_5140:FAff port map(x=>p(120)(20),y=>p(121)(20),Cin=>p(122)(20),clock=>clock,reset=>reset,s=>p(208)(20),cout=>p(209)(21));
FA_ff_5141:FAff port map(x=>p(120)(21),y=>p(121)(21),Cin=>p(122)(21),clock=>clock,reset=>reset,s=>p(208)(21),cout=>p(209)(22));
FA_ff_5142:FAff port map(x=>p(120)(22),y=>p(121)(22),Cin=>p(122)(22),clock=>clock,reset=>reset,s=>p(208)(22),cout=>p(209)(23));
FA_ff_5143:FAff port map(x=>p(120)(23),y=>p(121)(23),Cin=>p(122)(23),clock=>clock,reset=>reset,s=>p(208)(23),cout=>p(209)(24));
FA_ff_5144:FAff port map(x=>p(120)(24),y=>p(121)(24),Cin=>p(122)(24),clock=>clock,reset=>reset,s=>p(208)(24),cout=>p(209)(25));
FA_ff_5145:FAff port map(x=>p(120)(25),y=>p(121)(25),Cin=>p(122)(25),clock=>clock,reset=>reset,s=>p(208)(25),cout=>p(209)(26));
FA_ff_5146:FAff port map(x=>p(120)(26),y=>p(121)(26),Cin=>p(122)(26),clock=>clock,reset=>reset,s=>p(208)(26),cout=>p(209)(27));
FA_ff_5147:FAff port map(x=>p(120)(27),y=>p(121)(27),Cin=>p(122)(27),clock=>clock,reset=>reset,s=>p(208)(27),cout=>p(209)(28));
FA_ff_5148:FAff port map(x=>p(120)(28),y=>p(121)(28),Cin=>p(122)(28),clock=>clock,reset=>reset,s=>p(208)(28),cout=>p(209)(29));
FA_ff_5149:FAff port map(x=>p(120)(29),y=>p(121)(29),Cin=>p(122)(29),clock=>clock,reset=>reset,s=>p(208)(29),cout=>p(209)(30));
FA_ff_5150:FAff port map(x=>p(120)(30),y=>p(121)(30),Cin=>p(122)(30),clock=>clock,reset=>reset,s=>p(208)(30),cout=>p(209)(31));
FA_ff_5151:FAff port map(x=>p(120)(31),y=>p(121)(31),Cin=>p(122)(31),clock=>clock,reset=>reset,s=>p(208)(31),cout=>p(209)(32));
FA_ff_5152:FAff port map(x=>p(120)(32),y=>p(121)(32),Cin=>p(122)(32),clock=>clock,reset=>reset,s=>p(208)(32),cout=>p(209)(33));
FA_ff_5153:FAff port map(x=>p(120)(33),y=>p(121)(33),Cin=>p(122)(33),clock=>clock,reset=>reset,s=>p(208)(33),cout=>p(209)(34));
FA_ff_5154:FAff port map(x=>p(120)(34),y=>p(121)(34),Cin=>p(122)(34),clock=>clock,reset=>reset,s=>p(208)(34),cout=>p(209)(35));
FA_ff_5155:FAff port map(x=>p(120)(35),y=>p(121)(35),Cin=>p(122)(35),clock=>clock,reset=>reset,s=>p(208)(35),cout=>p(209)(36));
FA_ff_5156:FAff port map(x=>p(120)(36),y=>p(121)(36),Cin=>p(122)(36),clock=>clock,reset=>reset,s=>p(208)(36),cout=>p(209)(37));
FA_ff_5157:FAff port map(x=>p(120)(37),y=>p(121)(37),Cin=>p(122)(37),clock=>clock,reset=>reset,s=>p(208)(37),cout=>p(209)(38));
FA_ff_5158:FAff port map(x=>p(120)(38),y=>p(121)(38),Cin=>p(122)(38),clock=>clock,reset=>reset,s=>p(208)(38),cout=>p(209)(39));
FA_ff_5159:FAff port map(x=>p(120)(39),y=>p(121)(39),Cin=>p(122)(39),clock=>clock,reset=>reset,s=>p(208)(39),cout=>p(209)(40));
FA_ff_5160:FAff port map(x=>p(120)(40),y=>p(121)(40),Cin=>p(122)(40),clock=>clock,reset=>reset,s=>p(208)(40),cout=>p(209)(41));
FA_ff_5161:FAff port map(x=>p(120)(41),y=>p(121)(41),Cin=>p(122)(41),clock=>clock,reset=>reset,s=>p(208)(41),cout=>p(209)(42));
FA_ff_5162:FAff port map(x=>p(120)(42),y=>p(121)(42),Cin=>p(122)(42),clock=>clock,reset=>reset,s=>p(208)(42),cout=>p(209)(43));
FA_ff_5163:FAff port map(x=>p(120)(43),y=>p(121)(43),Cin=>p(122)(43),clock=>clock,reset=>reset,s=>p(208)(43),cout=>p(209)(44));
FA_ff_5164:FAff port map(x=>p(120)(44),y=>p(121)(44),Cin=>p(122)(44),clock=>clock,reset=>reset,s=>p(208)(44),cout=>p(209)(45));
FA_ff_5165:FAff port map(x=>p(120)(45),y=>p(121)(45),Cin=>p(122)(45),clock=>clock,reset=>reset,s=>p(208)(45),cout=>p(209)(46));
FA_ff_5166:FAff port map(x=>p(120)(46),y=>p(121)(46),Cin=>p(122)(46),clock=>clock,reset=>reset,s=>p(208)(46),cout=>p(209)(47));
FA_ff_5167:FAff port map(x=>p(120)(47),y=>p(121)(47),Cin=>p(122)(47),clock=>clock,reset=>reset,s=>p(208)(47),cout=>p(209)(48));
FA_ff_5168:FAff port map(x=>p(120)(48),y=>p(121)(48),Cin=>p(122)(48),clock=>clock,reset=>reset,s=>p(208)(48),cout=>p(209)(49));
FA_ff_5169:FAff port map(x=>p(120)(49),y=>p(121)(49),Cin=>p(122)(49),clock=>clock,reset=>reset,s=>p(208)(49),cout=>p(209)(50));
FA_ff_5170:FAff port map(x=>p(120)(50),y=>p(121)(50),Cin=>p(122)(50),clock=>clock,reset=>reset,s=>p(208)(50),cout=>p(209)(51));
FA_ff_5171:FAff port map(x=>p(120)(51),y=>p(121)(51),Cin=>p(122)(51),clock=>clock,reset=>reset,s=>p(208)(51),cout=>p(209)(52));
FA_ff_5172:FAff port map(x=>p(120)(52),y=>p(121)(52),Cin=>p(122)(52),clock=>clock,reset=>reset,s=>p(208)(52),cout=>p(209)(53));
FA_ff_5173:FAff port map(x=>p(120)(53),y=>p(121)(53),Cin=>p(122)(53),clock=>clock,reset=>reset,s=>p(208)(53),cout=>p(209)(54));
FA_ff_5174:FAff port map(x=>p(120)(54),y=>p(121)(54),Cin=>p(122)(54),clock=>clock,reset=>reset,s=>p(208)(54),cout=>p(209)(55));
FA_ff_5175:FAff port map(x=>p(120)(55),y=>p(121)(55),Cin=>p(122)(55),clock=>clock,reset=>reset,s=>p(208)(55),cout=>p(209)(56));
FA_ff_5176:FAff port map(x=>p(120)(56),y=>p(121)(56),Cin=>p(122)(56),clock=>clock,reset=>reset,s=>p(208)(56),cout=>p(209)(57));
FA_ff_5177:FAff port map(x=>p(120)(57),y=>p(121)(57),Cin=>p(122)(57),clock=>clock,reset=>reset,s=>p(208)(57),cout=>p(209)(58));
FA_ff_5178:FAff port map(x=>p(120)(58),y=>p(121)(58),Cin=>p(122)(58),clock=>clock,reset=>reset,s=>p(208)(58),cout=>p(209)(59));
FA_ff_5179:FAff port map(x=>p(120)(59),y=>p(121)(59),Cin=>p(122)(59),clock=>clock,reset=>reset,s=>p(208)(59),cout=>p(209)(60));
FA_ff_5180:FAff port map(x=>p(120)(60),y=>p(121)(60),Cin=>p(122)(60),clock=>clock,reset=>reset,s=>p(208)(60),cout=>p(209)(61));
FA_ff_5181:FAff port map(x=>p(120)(61),y=>p(121)(61),Cin=>p(122)(61),clock=>clock,reset=>reset,s=>p(208)(61),cout=>p(209)(62));
FA_ff_5182:FAff port map(x=>p(120)(62),y=>p(121)(62),Cin=>p(122)(62),clock=>clock,reset=>reset,s=>p(208)(62),cout=>p(209)(63));
FA_ff_5183:FAff port map(x=>p(120)(63),y=>p(121)(63),Cin=>p(122)(63),clock=>clock,reset=>reset,s=>p(208)(63),cout=>p(209)(64));
FA_ff_5184:FAff port map(x=>p(120)(64),y=>p(121)(64),Cin=>p(122)(64),clock=>clock,reset=>reset,s=>p(208)(64),cout=>p(209)(65));
FA_ff_5185:FAff port map(x=>p(120)(65),y=>p(121)(65),Cin=>p(122)(65),clock=>clock,reset=>reset,s=>p(208)(65),cout=>p(209)(66));
FA_ff_5186:FAff port map(x=>p(120)(66),y=>p(121)(66),Cin=>p(122)(66),clock=>clock,reset=>reset,s=>p(208)(66),cout=>p(209)(67));
FA_ff_5187:FAff port map(x=>p(120)(67),y=>p(121)(67),Cin=>p(122)(67),clock=>clock,reset=>reset,s=>p(208)(67),cout=>p(209)(68));
FA_ff_5188:FAff port map(x=>p(120)(68),y=>p(121)(68),Cin=>p(122)(68),clock=>clock,reset=>reset,s=>p(208)(68),cout=>p(209)(69));
FA_ff_5189:FAff port map(x=>p(120)(69),y=>p(121)(69),Cin=>p(122)(69),clock=>clock,reset=>reset,s=>p(208)(69),cout=>p(209)(70));
FA_ff_5190:FAff port map(x=>p(120)(70),y=>p(121)(70),Cin=>p(122)(70),clock=>clock,reset=>reset,s=>p(208)(70),cout=>p(209)(71));
FA_ff_5191:FAff port map(x=>p(120)(71),y=>p(121)(71),Cin=>p(122)(71),clock=>clock,reset=>reset,s=>p(208)(71),cout=>p(209)(72));
FA_ff_5192:FAff port map(x=>p(120)(72),y=>p(121)(72),Cin=>p(122)(72),clock=>clock,reset=>reset,s=>p(208)(72),cout=>p(209)(73));
FA_ff_5193:FAff port map(x=>p(120)(73),y=>p(121)(73),Cin=>p(122)(73),clock=>clock,reset=>reset,s=>p(208)(73),cout=>p(209)(74));
FA_ff_5194:FAff port map(x=>p(120)(74),y=>p(121)(74),Cin=>p(122)(74),clock=>clock,reset=>reset,s=>p(208)(74),cout=>p(209)(75));
FA_ff_5195:FAff port map(x=>p(120)(75),y=>p(121)(75),Cin=>p(122)(75),clock=>clock,reset=>reset,s=>p(208)(75),cout=>p(209)(76));
FA_ff_5196:FAff port map(x=>p(120)(76),y=>p(121)(76),Cin=>p(122)(76),clock=>clock,reset=>reset,s=>p(208)(76),cout=>p(209)(77));
FA_ff_5197:FAff port map(x=>p(120)(77),y=>p(121)(77),Cin=>p(122)(77),clock=>clock,reset=>reset,s=>p(208)(77),cout=>p(209)(78));
FA_ff_5198:FAff port map(x=>p(120)(78),y=>p(121)(78),Cin=>p(122)(78),clock=>clock,reset=>reset,s=>p(208)(78),cout=>p(209)(79));
FA_ff_5199:FAff port map(x=>p(120)(79),y=>p(121)(79),Cin=>p(122)(79),clock=>clock,reset=>reset,s=>p(208)(79),cout=>p(209)(80));
FA_ff_5200:FAff port map(x=>p(120)(80),y=>p(121)(80),Cin=>p(122)(80),clock=>clock,reset=>reset,s=>p(208)(80),cout=>p(209)(81));
FA_ff_5201:FAff port map(x=>p(120)(81),y=>p(121)(81),Cin=>p(122)(81),clock=>clock,reset=>reset,s=>p(208)(81),cout=>p(209)(82));
FA_ff_5202:FAff port map(x=>p(120)(82),y=>p(121)(82),Cin=>p(122)(82),clock=>clock,reset=>reset,s=>p(208)(82),cout=>p(209)(83));
FA_ff_5203:FAff port map(x=>p(120)(83),y=>p(121)(83),Cin=>p(122)(83),clock=>clock,reset=>reset,s=>p(208)(83),cout=>p(209)(84));
FA_ff_5204:FAff port map(x=>p(120)(84),y=>p(121)(84),Cin=>p(122)(84),clock=>clock,reset=>reset,s=>p(208)(84),cout=>p(209)(85));
FA_ff_5205:FAff port map(x=>p(120)(85),y=>p(121)(85),Cin=>p(122)(85),clock=>clock,reset=>reset,s=>p(208)(85),cout=>p(209)(86));
FA_ff_5206:FAff port map(x=>p(120)(86),y=>p(121)(86),Cin=>p(122)(86),clock=>clock,reset=>reset,s=>p(208)(86),cout=>p(209)(87));
FA_ff_5207:FAff port map(x=>p(120)(87),y=>p(121)(87),Cin=>p(122)(87),clock=>clock,reset=>reset,s=>p(208)(87),cout=>p(209)(88));
FA_ff_5208:FAff port map(x=>p(120)(88),y=>p(121)(88),Cin=>p(122)(88),clock=>clock,reset=>reset,s=>p(208)(88),cout=>p(209)(89));
FA_ff_5209:FAff port map(x=>p(120)(89),y=>p(121)(89),Cin=>p(122)(89),clock=>clock,reset=>reset,s=>p(208)(89),cout=>p(209)(90));
FA_ff_5210:FAff port map(x=>p(120)(90),y=>p(121)(90),Cin=>p(122)(90),clock=>clock,reset=>reset,s=>p(208)(90),cout=>p(209)(91));
FA_ff_5211:FAff port map(x=>p(120)(91),y=>p(121)(91),Cin=>p(122)(91),clock=>clock,reset=>reset,s=>p(208)(91),cout=>p(209)(92));
FA_ff_5212:FAff port map(x=>p(120)(92),y=>p(121)(92),Cin=>p(122)(92),clock=>clock,reset=>reset,s=>p(208)(92),cout=>p(209)(93));
FA_ff_5213:FAff port map(x=>p(120)(93),y=>p(121)(93),Cin=>p(122)(93),clock=>clock,reset=>reset,s=>p(208)(93),cout=>p(209)(94));
FA_ff_5214:FAff port map(x=>p(120)(94),y=>p(121)(94),Cin=>p(122)(94),clock=>clock,reset=>reset,s=>p(208)(94),cout=>p(209)(95));
FA_ff_5215:FAff port map(x=>p(120)(95),y=>p(121)(95),Cin=>p(122)(95),clock=>clock,reset=>reset,s=>p(208)(95),cout=>p(209)(96));
FA_ff_5216:FAff port map(x=>p(120)(96),y=>p(121)(96),Cin=>p(122)(96),clock=>clock,reset=>reset,s=>p(208)(96),cout=>p(209)(97));
FA_ff_5217:FAff port map(x=>p(120)(97),y=>p(121)(97),Cin=>p(122)(97),clock=>clock,reset=>reset,s=>p(208)(97),cout=>p(209)(98));
FA_ff_5218:FAff port map(x=>p(120)(98),y=>p(121)(98),Cin=>p(122)(98),clock=>clock,reset=>reset,s=>p(208)(98),cout=>p(209)(99));
FA_ff_5219:FAff port map(x=>p(120)(99),y=>p(121)(99),Cin=>p(122)(99),clock=>clock,reset=>reset,s=>p(208)(99),cout=>p(209)(100));
FA_ff_5220:FAff port map(x=>p(120)(100),y=>p(121)(100),Cin=>p(122)(100),clock=>clock,reset=>reset,s=>p(208)(100),cout=>p(209)(101));
FA_ff_5221:FAff port map(x=>p(120)(101),y=>p(121)(101),Cin=>p(122)(101),clock=>clock,reset=>reset,s=>p(208)(101),cout=>p(209)(102));
FA_ff_5222:FAff port map(x=>p(120)(102),y=>p(121)(102),Cin=>p(122)(102),clock=>clock,reset=>reset,s=>p(208)(102),cout=>p(209)(103));
FA_ff_5223:FAff port map(x=>p(120)(103),y=>p(121)(103),Cin=>p(122)(103),clock=>clock,reset=>reset,s=>p(208)(103),cout=>p(209)(104));
FA_ff_5224:FAff port map(x=>p(120)(104),y=>p(121)(104),Cin=>p(122)(104),clock=>clock,reset=>reset,s=>p(208)(104),cout=>p(209)(105));
FA_ff_5225:FAff port map(x=>p(120)(105),y=>p(121)(105),Cin=>p(122)(105),clock=>clock,reset=>reset,s=>p(208)(105),cout=>p(209)(106));
FA_ff_5226:FAff port map(x=>p(120)(106),y=>p(121)(106),Cin=>p(122)(106),clock=>clock,reset=>reset,s=>p(208)(106),cout=>p(209)(107));
FA_ff_5227:FAff port map(x=>p(120)(107),y=>p(121)(107),Cin=>p(122)(107),clock=>clock,reset=>reset,s=>p(208)(107),cout=>p(209)(108));
FA_ff_5228:FAff port map(x=>p(120)(108),y=>p(121)(108),Cin=>p(122)(108),clock=>clock,reset=>reset,s=>p(208)(108),cout=>p(209)(109));
FA_ff_5229:FAff port map(x=>p(120)(109),y=>p(121)(109),Cin=>p(122)(109),clock=>clock,reset=>reset,s=>p(208)(109),cout=>p(209)(110));
FA_ff_5230:FAff port map(x=>p(120)(110),y=>p(121)(110),Cin=>p(122)(110),clock=>clock,reset=>reset,s=>p(208)(110),cout=>p(209)(111));
FA_ff_5231:FAff port map(x=>p(120)(111),y=>p(121)(111),Cin=>p(122)(111),clock=>clock,reset=>reset,s=>p(208)(111),cout=>p(209)(112));
FA_ff_5232:FAff port map(x=>p(120)(112),y=>p(121)(112),Cin=>p(122)(112),clock=>clock,reset=>reset,s=>p(208)(112),cout=>p(209)(113));
FA_ff_5233:FAff port map(x=>p(120)(113),y=>p(121)(113),Cin=>p(122)(113),clock=>clock,reset=>reset,s=>p(208)(113),cout=>p(209)(114));
FA_ff_5234:FAff port map(x=>p(120)(114),y=>p(121)(114),Cin=>p(122)(114),clock=>clock,reset=>reset,s=>p(208)(114),cout=>p(209)(115));
FA_ff_5235:FAff port map(x=>p(120)(115),y=>p(121)(115),Cin=>p(122)(115),clock=>clock,reset=>reset,s=>p(208)(115),cout=>p(209)(116));
FA_ff_5236:FAff port map(x=>p(120)(116),y=>p(121)(116),Cin=>p(122)(116),clock=>clock,reset=>reset,s=>p(208)(116),cout=>p(209)(117));
FA_ff_5237:FAff port map(x=>p(120)(117),y=>p(121)(117),Cin=>p(122)(117),clock=>clock,reset=>reset,s=>p(208)(117),cout=>p(209)(118));
FA_ff_5238:FAff port map(x=>p(120)(118),y=>p(121)(118),Cin=>p(122)(118),clock=>clock,reset=>reset,s=>p(208)(118),cout=>p(209)(119));
FA_ff_5239:FAff port map(x=>p(120)(119),y=>p(121)(119),Cin=>p(122)(119),clock=>clock,reset=>reset,s=>p(208)(119),cout=>p(209)(120));
FA_ff_5240:FAff port map(x=>p(120)(120),y=>p(121)(120),Cin=>p(122)(120),clock=>clock,reset=>reset,s=>p(208)(120),cout=>p(209)(121));
FA_ff_5241:FAff port map(x=>p(120)(121),y=>p(121)(121),Cin=>p(122)(121),clock=>clock,reset=>reset,s=>p(208)(121),cout=>p(209)(122));
FA_ff_5242:FAff port map(x=>p(120)(122),y=>p(121)(122),Cin=>p(122)(122),clock=>clock,reset=>reset,s=>p(208)(122),cout=>p(209)(123));
FA_ff_5243:FAff port map(x=>p(120)(123),y=>p(121)(123),Cin=>p(122)(123),clock=>clock,reset=>reset,s=>p(208)(123),cout=>p(209)(124));
FA_ff_5244:FAff port map(x=>p(120)(124),y=>p(121)(124),Cin=>p(122)(124),clock=>clock,reset=>reset,s=>p(208)(124),cout=>p(209)(125));
FA_ff_5245:FAff port map(x=>p(120)(125),y=>p(121)(125),Cin=>p(122)(125),clock=>clock,reset=>reset,s=>p(208)(125),cout=>p(209)(126));
FA_ff_5246:FAff port map(x=>p(120)(126),y=>p(121)(126),Cin=>p(122)(126),clock=>clock,reset=>reset,s=>p(208)(126),cout=>p(209)(127));
FA_ff_5247:FAff port map(x=>p(120)(127),y=>p(121)(127),Cin=>p(122)(127),clock=>clock,reset=>reset,s=>p(208)(127),cout=>p(209)(128));
FA_ff_5248:FAff port map(x=>p(123)(0),y=>p(124)(0),Cin=>p(125)(0),clock=>clock,reset=>reset,s=>p(210)(0),cout=>p(211)(1));
FA_ff_5249:FAff port map(x=>p(123)(1),y=>p(124)(1),Cin=>p(125)(1),clock=>clock,reset=>reset,s=>p(210)(1),cout=>p(211)(2));
FA_ff_5250:FAff port map(x=>p(123)(2),y=>p(124)(2),Cin=>p(125)(2),clock=>clock,reset=>reset,s=>p(210)(2),cout=>p(211)(3));
FA_ff_5251:FAff port map(x=>p(123)(3),y=>p(124)(3),Cin=>p(125)(3),clock=>clock,reset=>reset,s=>p(210)(3),cout=>p(211)(4));
FA_ff_5252:FAff port map(x=>p(123)(4),y=>p(124)(4),Cin=>p(125)(4),clock=>clock,reset=>reset,s=>p(210)(4),cout=>p(211)(5));
FA_ff_5253:FAff port map(x=>p(123)(5),y=>p(124)(5),Cin=>p(125)(5),clock=>clock,reset=>reset,s=>p(210)(5),cout=>p(211)(6));
FA_ff_5254:FAff port map(x=>p(123)(6),y=>p(124)(6),Cin=>p(125)(6),clock=>clock,reset=>reset,s=>p(210)(6),cout=>p(211)(7));
FA_ff_5255:FAff port map(x=>p(123)(7),y=>p(124)(7),Cin=>p(125)(7),clock=>clock,reset=>reset,s=>p(210)(7),cout=>p(211)(8));
FA_ff_5256:FAff port map(x=>p(123)(8),y=>p(124)(8),Cin=>p(125)(8),clock=>clock,reset=>reset,s=>p(210)(8),cout=>p(211)(9));
FA_ff_5257:FAff port map(x=>p(123)(9),y=>p(124)(9),Cin=>p(125)(9),clock=>clock,reset=>reset,s=>p(210)(9),cout=>p(211)(10));
FA_ff_5258:FAff port map(x=>p(123)(10),y=>p(124)(10),Cin=>p(125)(10),clock=>clock,reset=>reset,s=>p(210)(10),cout=>p(211)(11));
FA_ff_5259:FAff port map(x=>p(123)(11),y=>p(124)(11),Cin=>p(125)(11),clock=>clock,reset=>reset,s=>p(210)(11),cout=>p(211)(12));
FA_ff_5260:FAff port map(x=>p(123)(12),y=>p(124)(12),Cin=>p(125)(12),clock=>clock,reset=>reset,s=>p(210)(12),cout=>p(211)(13));
FA_ff_5261:FAff port map(x=>p(123)(13),y=>p(124)(13),Cin=>p(125)(13),clock=>clock,reset=>reset,s=>p(210)(13),cout=>p(211)(14));
FA_ff_5262:FAff port map(x=>p(123)(14),y=>p(124)(14),Cin=>p(125)(14),clock=>clock,reset=>reset,s=>p(210)(14),cout=>p(211)(15));
FA_ff_5263:FAff port map(x=>p(123)(15),y=>p(124)(15),Cin=>p(125)(15),clock=>clock,reset=>reset,s=>p(210)(15),cout=>p(211)(16));
FA_ff_5264:FAff port map(x=>p(123)(16),y=>p(124)(16),Cin=>p(125)(16),clock=>clock,reset=>reset,s=>p(210)(16),cout=>p(211)(17));
FA_ff_5265:FAff port map(x=>p(123)(17),y=>p(124)(17),Cin=>p(125)(17),clock=>clock,reset=>reset,s=>p(210)(17),cout=>p(211)(18));
FA_ff_5266:FAff port map(x=>p(123)(18),y=>p(124)(18),Cin=>p(125)(18),clock=>clock,reset=>reset,s=>p(210)(18),cout=>p(211)(19));
FA_ff_5267:FAff port map(x=>p(123)(19),y=>p(124)(19),Cin=>p(125)(19),clock=>clock,reset=>reset,s=>p(210)(19),cout=>p(211)(20));
FA_ff_5268:FAff port map(x=>p(123)(20),y=>p(124)(20),Cin=>p(125)(20),clock=>clock,reset=>reset,s=>p(210)(20),cout=>p(211)(21));
FA_ff_5269:FAff port map(x=>p(123)(21),y=>p(124)(21),Cin=>p(125)(21),clock=>clock,reset=>reset,s=>p(210)(21),cout=>p(211)(22));
FA_ff_5270:FAff port map(x=>p(123)(22),y=>p(124)(22),Cin=>p(125)(22),clock=>clock,reset=>reset,s=>p(210)(22),cout=>p(211)(23));
FA_ff_5271:FAff port map(x=>p(123)(23),y=>p(124)(23),Cin=>p(125)(23),clock=>clock,reset=>reset,s=>p(210)(23),cout=>p(211)(24));
FA_ff_5272:FAff port map(x=>p(123)(24),y=>p(124)(24),Cin=>p(125)(24),clock=>clock,reset=>reset,s=>p(210)(24),cout=>p(211)(25));
FA_ff_5273:FAff port map(x=>p(123)(25),y=>p(124)(25),Cin=>p(125)(25),clock=>clock,reset=>reset,s=>p(210)(25),cout=>p(211)(26));
FA_ff_5274:FAff port map(x=>p(123)(26),y=>p(124)(26),Cin=>p(125)(26),clock=>clock,reset=>reset,s=>p(210)(26),cout=>p(211)(27));
FA_ff_5275:FAff port map(x=>p(123)(27),y=>p(124)(27),Cin=>p(125)(27),clock=>clock,reset=>reset,s=>p(210)(27),cout=>p(211)(28));
FA_ff_5276:FAff port map(x=>p(123)(28),y=>p(124)(28),Cin=>p(125)(28),clock=>clock,reset=>reset,s=>p(210)(28),cout=>p(211)(29));
FA_ff_5277:FAff port map(x=>p(123)(29),y=>p(124)(29),Cin=>p(125)(29),clock=>clock,reset=>reset,s=>p(210)(29),cout=>p(211)(30));
FA_ff_5278:FAff port map(x=>p(123)(30),y=>p(124)(30),Cin=>p(125)(30),clock=>clock,reset=>reset,s=>p(210)(30),cout=>p(211)(31));
FA_ff_5279:FAff port map(x=>p(123)(31),y=>p(124)(31),Cin=>p(125)(31),clock=>clock,reset=>reset,s=>p(210)(31),cout=>p(211)(32));
FA_ff_5280:FAff port map(x=>p(123)(32),y=>p(124)(32),Cin=>p(125)(32),clock=>clock,reset=>reset,s=>p(210)(32),cout=>p(211)(33));
FA_ff_5281:FAff port map(x=>p(123)(33),y=>p(124)(33),Cin=>p(125)(33),clock=>clock,reset=>reset,s=>p(210)(33),cout=>p(211)(34));
FA_ff_5282:FAff port map(x=>p(123)(34),y=>p(124)(34),Cin=>p(125)(34),clock=>clock,reset=>reset,s=>p(210)(34),cout=>p(211)(35));
FA_ff_5283:FAff port map(x=>p(123)(35),y=>p(124)(35),Cin=>p(125)(35),clock=>clock,reset=>reset,s=>p(210)(35),cout=>p(211)(36));
FA_ff_5284:FAff port map(x=>p(123)(36),y=>p(124)(36),Cin=>p(125)(36),clock=>clock,reset=>reset,s=>p(210)(36),cout=>p(211)(37));
FA_ff_5285:FAff port map(x=>p(123)(37),y=>p(124)(37),Cin=>p(125)(37),clock=>clock,reset=>reset,s=>p(210)(37),cout=>p(211)(38));
FA_ff_5286:FAff port map(x=>p(123)(38),y=>p(124)(38),Cin=>p(125)(38),clock=>clock,reset=>reset,s=>p(210)(38),cout=>p(211)(39));
FA_ff_5287:FAff port map(x=>p(123)(39),y=>p(124)(39),Cin=>p(125)(39),clock=>clock,reset=>reset,s=>p(210)(39),cout=>p(211)(40));
FA_ff_5288:FAff port map(x=>p(123)(40),y=>p(124)(40),Cin=>p(125)(40),clock=>clock,reset=>reset,s=>p(210)(40),cout=>p(211)(41));
FA_ff_5289:FAff port map(x=>p(123)(41),y=>p(124)(41),Cin=>p(125)(41),clock=>clock,reset=>reset,s=>p(210)(41),cout=>p(211)(42));
FA_ff_5290:FAff port map(x=>p(123)(42),y=>p(124)(42),Cin=>p(125)(42),clock=>clock,reset=>reset,s=>p(210)(42),cout=>p(211)(43));
FA_ff_5291:FAff port map(x=>p(123)(43),y=>p(124)(43),Cin=>p(125)(43),clock=>clock,reset=>reset,s=>p(210)(43),cout=>p(211)(44));
FA_ff_5292:FAff port map(x=>p(123)(44),y=>p(124)(44),Cin=>p(125)(44),clock=>clock,reset=>reset,s=>p(210)(44),cout=>p(211)(45));
FA_ff_5293:FAff port map(x=>p(123)(45),y=>p(124)(45),Cin=>p(125)(45),clock=>clock,reset=>reset,s=>p(210)(45),cout=>p(211)(46));
FA_ff_5294:FAff port map(x=>p(123)(46),y=>p(124)(46),Cin=>p(125)(46),clock=>clock,reset=>reset,s=>p(210)(46),cout=>p(211)(47));
FA_ff_5295:FAff port map(x=>p(123)(47),y=>p(124)(47),Cin=>p(125)(47),clock=>clock,reset=>reset,s=>p(210)(47),cout=>p(211)(48));
FA_ff_5296:FAff port map(x=>p(123)(48),y=>p(124)(48),Cin=>p(125)(48),clock=>clock,reset=>reset,s=>p(210)(48),cout=>p(211)(49));
FA_ff_5297:FAff port map(x=>p(123)(49),y=>p(124)(49),Cin=>p(125)(49),clock=>clock,reset=>reset,s=>p(210)(49),cout=>p(211)(50));
FA_ff_5298:FAff port map(x=>p(123)(50),y=>p(124)(50),Cin=>p(125)(50),clock=>clock,reset=>reset,s=>p(210)(50),cout=>p(211)(51));
FA_ff_5299:FAff port map(x=>p(123)(51),y=>p(124)(51),Cin=>p(125)(51),clock=>clock,reset=>reset,s=>p(210)(51),cout=>p(211)(52));
FA_ff_5300:FAff port map(x=>p(123)(52),y=>p(124)(52),Cin=>p(125)(52),clock=>clock,reset=>reset,s=>p(210)(52),cout=>p(211)(53));
FA_ff_5301:FAff port map(x=>p(123)(53),y=>p(124)(53),Cin=>p(125)(53),clock=>clock,reset=>reset,s=>p(210)(53),cout=>p(211)(54));
FA_ff_5302:FAff port map(x=>p(123)(54),y=>p(124)(54),Cin=>p(125)(54),clock=>clock,reset=>reset,s=>p(210)(54),cout=>p(211)(55));
FA_ff_5303:FAff port map(x=>p(123)(55),y=>p(124)(55),Cin=>p(125)(55),clock=>clock,reset=>reset,s=>p(210)(55),cout=>p(211)(56));
FA_ff_5304:FAff port map(x=>p(123)(56),y=>p(124)(56),Cin=>p(125)(56),clock=>clock,reset=>reset,s=>p(210)(56),cout=>p(211)(57));
FA_ff_5305:FAff port map(x=>p(123)(57),y=>p(124)(57),Cin=>p(125)(57),clock=>clock,reset=>reset,s=>p(210)(57),cout=>p(211)(58));
FA_ff_5306:FAff port map(x=>p(123)(58),y=>p(124)(58),Cin=>p(125)(58),clock=>clock,reset=>reset,s=>p(210)(58),cout=>p(211)(59));
FA_ff_5307:FAff port map(x=>p(123)(59),y=>p(124)(59),Cin=>p(125)(59),clock=>clock,reset=>reset,s=>p(210)(59),cout=>p(211)(60));
FA_ff_5308:FAff port map(x=>p(123)(60),y=>p(124)(60),Cin=>p(125)(60),clock=>clock,reset=>reset,s=>p(210)(60),cout=>p(211)(61));
FA_ff_5309:FAff port map(x=>p(123)(61),y=>p(124)(61),Cin=>p(125)(61),clock=>clock,reset=>reset,s=>p(210)(61),cout=>p(211)(62));
FA_ff_5310:FAff port map(x=>p(123)(62),y=>p(124)(62),Cin=>p(125)(62),clock=>clock,reset=>reset,s=>p(210)(62),cout=>p(211)(63));
FA_ff_5311:FAff port map(x=>p(123)(63),y=>p(124)(63),Cin=>p(125)(63),clock=>clock,reset=>reset,s=>p(210)(63),cout=>p(211)(64));
FA_ff_5312:FAff port map(x=>p(123)(64),y=>p(124)(64),Cin=>p(125)(64),clock=>clock,reset=>reset,s=>p(210)(64),cout=>p(211)(65));
FA_ff_5313:FAff port map(x=>p(123)(65),y=>p(124)(65),Cin=>p(125)(65),clock=>clock,reset=>reset,s=>p(210)(65),cout=>p(211)(66));
FA_ff_5314:FAff port map(x=>p(123)(66),y=>p(124)(66),Cin=>p(125)(66),clock=>clock,reset=>reset,s=>p(210)(66),cout=>p(211)(67));
FA_ff_5315:FAff port map(x=>p(123)(67),y=>p(124)(67),Cin=>p(125)(67),clock=>clock,reset=>reset,s=>p(210)(67),cout=>p(211)(68));
FA_ff_5316:FAff port map(x=>p(123)(68),y=>p(124)(68),Cin=>p(125)(68),clock=>clock,reset=>reset,s=>p(210)(68),cout=>p(211)(69));
FA_ff_5317:FAff port map(x=>p(123)(69),y=>p(124)(69),Cin=>p(125)(69),clock=>clock,reset=>reset,s=>p(210)(69),cout=>p(211)(70));
FA_ff_5318:FAff port map(x=>p(123)(70),y=>p(124)(70),Cin=>p(125)(70),clock=>clock,reset=>reset,s=>p(210)(70),cout=>p(211)(71));
FA_ff_5319:FAff port map(x=>p(123)(71),y=>p(124)(71),Cin=>p(125)(71),clock=>clock,reset=>reset,s=>p(210)(71),cout=>p(211)(72));
FA_ff_5320:FAff port map(x=>p(123)(72),y=>p(124)(72),Cin=>p(125)(72),clock=>clock,reset=>reset,s=>p(210)(72),cout=>p(211)(73));
FA_ff_5321:FAff port map(x=>p(123)(73),y=>p(124)(73),Cin=>p(125)(73),clock=>clock,reset=>reset,s=>p(210)(73),cout=>p(211)(74));
FA_ff_5322:FAff port map(x=>p(123)(74),y=>p(124)(74),Cin=>p(125)(74),clock=>clock,reset=>reset,s=>p(210)(74),cout=>p(211)(75));
FA_ff_5323:FAff port map(x=>p(123)(75),y=>p(124)(75),Cin=>p(125)(75),clock=>clock,reset=>reset,s=>p(210)(75),cout=>p(211)(76));
FA_ff_5324:FAff port map(x=>p(123)(76),y=>p(124)(76),Cin=>p(125)(76),clock=>clock,reset=>reset,s=>p(210)(76),cout=>p(211)(77));
FA_ff_5325:FAff port map(x=>p(123)(77),y=>p(124)(77),Cin=>p(125)(77),clock=>clock,reset=>reset,s=>p(210)(77),cout=>p(211)(78));
FA_ff_5326:FAff port map(x=>p(123)(78),y=>p(124)(78),Cin=>p(125)(78),clock=>clock,reset=>reset,s=>p(210)(78),cout=>p(211)(79));
FA_ff_5327:FAff port map(x=>p(123)(79),y=>p(124)(79),Cin=>p(125)(79),clock=>clock,reset=>reset,s=>p(210)(79),cout=>p(211)(80));
FA_ff_5328:FAff port map(x=>p(123)(80),y=>p(124)(80),Cin=>p(125)(80),clock=>clock,reset=>reset,s=>p(210)(80),cout=>p(211)(81));
FA_ff_5329:FAff port map(x=>p(123)(81),y=>p(124)(81),Cin=>p(125)(81),clock=>clock,reset=>reset,s=>p(210)(81),cout=>p(211)(82));
FA_ff_5330:FAff port map(x=>p(123)(82),y=>p(124)(82),Cin=>p(125)(82),clock=>clock,reset=>reset,s=>p(210)(82),cout=>p(211)(83));
FA_ff_5331:FAff port map(x=>p(123)(83),y=>p(124)(83),Cin=>p(125)(83),clock=>clock,reset=>reset,s=>p(210)(83),cout=>p(211)(84));
FA_ff_5332:FAff port map(x=>p(123)(84),y=>p(124)(84),Cin=>p(125)(84),clock=>clock,reset=>reset,s=>p(210)(84),cout=>p(211)(85));
FA_ff_5333:FAff port map(x=>p(123)(85),y=>p(124)(85),Cin=>p(125)(85),clock=>clock,reset=>reset,s=>p(210)(85),cout=>p(211)(86));
FA_ff_5334:FAff port map(x=>p(123)(86),y=>p(124)(86),Cin=>p(125)(86),clock=>clock,reset=>reset,s=>p(210)(86),cout=>p(211)(87));
FA_ff_5335:FAff port map(x=>p(123)(87),y=>p(124)(87),Cin=>p(125)(87),clock=>clock,reset=>reset,s=>p(210)(87),cout=>p(211)(88));
FA_ff_5336:FAff port map(x=>p(123)(88),y=>p(124)(88),Cin=>p(125)(88),clock=>clock,reset=>reset,s=>p(210)(88),cout=>p(211)(89));
FA_ff_5337:FAff port map(x=>p(123)(89),y=>p(124)(89),Cin=>p(125)(89),clock=>clock,reset=>reset,s=>p(210)(89),cout=>p(211)(90));
FA_ff_5338:FAff port map(x=>p(123)(90),y=>p(124)(90),Cin=>p(125)(90),clock=>clock,reset=>reset,s=>p(210)(90),cout=>p(211)(91));
FA_ff_5339:FAff port map(x=>p(123)(91),y=>p(124)(91),Cin=>p(125)(91),clock=>clock,reset=>reset,s=>p(210)(91),cout=>p(211)(92));
FA_ff_5340:FAff port map(x=>p(123)(92),y=>p(124)(92),Cin=>p(125)(92),clock=>clock,reset=>reset,s=>p(210)(92),cout=>p(211)(93));
FA_ff_5341:FAff port map(x=>p(123)(93),y=>p(124)(93),Cin=>p(125)(93),clock=>clock,reset=>reset,s=>p(210)(93),cout=>p(211)(94));
FA_ff_5342:FAff port map(x=>p(123)(94),y=>p(124)(94),Cin=>p(125)(94),clock=>clock,reset=>reset,s=>p(210)(94),cout=>p(211)(95));
FA_ff_5343:FAff port map(x=>p(123)(95),y=>p(124)(95),Cin=>p(125)(95),clock=>clock,reset=>reset,s=>p(210)(95),cout=>p(211)(96));
FA_ff_5344:FAff port map(x=>p(123)(96),y=>p(124)(96),Cin=>p(125)(96),clock=>clock,reset=>reset,s=>p(210)(96),cout=>p(211)(97));
FA_ff_5345:FAff port map(x=>p(123)(97),y=>p(124)(97),Cin=>p(125)(97),clock=>clock,reset=>reset,s=>p(210)(97),cout=>p(211)(98));
FA_ff_5346:FAff port map(x=>p(123)(98),y=>p(124)(98),Cin=>p(125)(98),clock=>clock,reset=>reset,s=>p(210)(98),cout=>p(211)(99));
FA_ff_5347:FAff port map(x=>p(123)(99),y=>p(124)(99),Cin=>p(125)(99),clock=>clock,reset=>reset,s=>p(210)(99),cout=>p(211)(100));
FA_ff_5348:FAff port map(x=>p(123)(100),y=>p(124)(100),Cin=>p(125)(100),clock=>clock,reset=>reset,s=>p(210)(100),cout=>p(211)(101));
FA_ff_5349:FAff port map(x=>p(123)(101),y=>p(124)(101),Cin=>p(125)(101),clock=>clock,reset=>reset,s=>p(210)(101),cout=>p(211)(102));
FA_ff_5350:FAff port map(x=>p(123)(102),y=>p(124)(102),Cin=>p(125)(102),clock=>clock,reset=>reset,s=>p(210)(102),cout=>p(211)(103));
FA_ff_5351:FAff port map(x=>p(123)(103),y=>p(124)(103),Cin=>p(125)(103),clock=>clock,reset=>reset,s=>p(210)(103),cout=>p(211)(104));
FA_ff_5352:FAff port map(x=>p(123)(104),y=>p(124)(104),Cin=>p(125)(104),clock=>clock,reset=>reset,s=>p(210)(104),cout=>p(211)(105));
FA_ff_5353:FAff port map(x=>p(123)(105),y=>p(124)(105),Cin=>p(125)(105),clock=>clock,reset=>reset,s=>p(210)(105),cout=>p(211)(106));
FA_ff_5354:FAff port map(x=>p(123)(106),y=>p(124)(106),Cin=>p(125)(106),clock=>clock,reset=>reset,s=>p(210)(106),cout=>p(211)(107));
FA_ff_5355:FAff port map(x=>p(123)(107),y=>p(124)(107),Cin=>p(125)(107),clock=>clock,reset=>reset,s=>p(210)(107),cout=>p(211)(108));
FA_ff_5356:FAff port map(x=>p(123)(108),y=>p(124)(108),Cin=>p(125)(108),clock=>clock,reset=>reset,s=>p(210)(108),cout=>p(211)(109));
FA_ff_5357:FAff port map(x=>p(123)(109),y=>p(124)(109),Cin=>p(125)(109),clock=>clock,reset=>reset,s=>p(210)(109),cout=>p(211)(110));
FA_ff_5358:FAff port map(x=>p(123)(110),y=>p(124)(110),Cin=>p(125)(110),clock=>clock,reset=>reset,s=>p(210)(110),cout=>p(211)(111));
FA_ff_5359:FAff port map(x=>p(123)(111),y=>p(124)(111),Cin=>p(125)(111),clock=>clock,reset=>reset,s=>p(210)(111),cout=>p(211)(112));
FA_ff_5360:FAff port map(x=>p(123)(112),y=>p(124)(112),Cin=>p(125)(112),clock=>clock,reset=>reset,s=>p(210)(112),cout=>p(211)(113));
FA_ff_5361:FAff port map(x=>p(123)(113),y=>p(124)(113),Cin=>p(125)(113),clock=>clock,reset=>reset,s=>p(210)(113),cout=>p(211)(114));
FA_ff_5362:FAff port map(x=>p(123)(114),y=>p(124)(114),Cin=>p(125)(114),clock=>clock,reset=>reset,s=>p(210)(114),cout=>p(211)(115));
FA_ff_5363:FAff port map(x=>p(123)(115),y=>p(124)(115),Cin=>p(125)(115),clock=>clock,reset=>reset,s=>p(210)(115),cout=>p(211)(116));
FA_ff_5364:FAff port map(x=>p(123)(116),y=>p(124)(116),Cin=>p(125)(116),clock=>clock,reset=>reset,s=>p(210)(116),cout=>p(211)(117));
FA_ff_5365:FAff port map(x=>p(123)(117),y=>p(124)(117),Cin=>p(125)(117),clock=>clock,reset=>reset,s=>p(210)(117),cout=>p(211)(118));
FA_ff_5366:FAff port map(x=>p(123)(118),y=>p(124)(118),Cin=>p(125)(118),clock=>clock,reset=>reset,s=>p(210)(118),cout=>p(211)(119));
FA_ff_5367:FAff port map(x=>p(123)(119),y=>p(124)(119),Cin=>p(125)(119),clock=>clock,reset=>reset,s=>p(210)(119),cout=>p(211)(120));
FA_ff_5368:FAff port map(x=>p(123)(120),y=>p(124)(120),Cin=>p(125)(120),clock=>clock,reset=>reset,s=>p(210)(120),cout=>p(211)(121));
FA_ff_5369:FAff port map(x=>p(123)(121),y=>p(124)(121),Cin=>p(125)(121),clock=>clock,reset=>reset,s=>p(210)(121),cout=>p(211)(122));
FA_ff_5370:FAff port map(x=>p(123)(122),y=>p(124)(122),Cin=>p(125)(122),clock=>clock,reset=>reset,s=>p(210)(122),cout=>p(211)(123));
FA_ff_5371:FAff port map(x=>p(123)(123),y=>p(124)(123),Cin=>p(125)(123),clock=>clock,reset=>reset,s=>p(210)(123),cout=>p(211)(124));
FA_ff_5372:FAff port map(x=>p(123)(124),y=>p(124)(124),Cin=>p(125)(124),clock=>clock,reset=>reset,s=>p(210)(124),cout=>p(211)(125));
FA_ff_5373:FAff port map(x=>p(123)(125),y=>p(124)(125),Cin=>p(125)(125),clock=>clock,reset=>reset,s=>p(210)(125),cout=>p(211)(126));
FA_ff_5374:FAff port map(x=>p(123)(126),y=>p(124)(126),Cin=>p(125)(126),clock=>clock,reset=>reset,s=>p(210)(126),cout=>p(211)(127));
FA_ff_5375:FAff port map(x=>p(123)(127),y=>p(124)(127),Cin=>p(125)(127),clock=>clock,reset=>reset,s=>p(210)(127),cout=>p(211)(128));
p(212)(0)<=p(126)(0);
p(212)(1)<=p(126)(1);
p(212)(2)<=p(126)(2);
p(212)(3)<=p(126)(3);
p(212)(4)<=p(126)(4);
p(212)(5)<=p(126)(5);
p(212)(6)<=p(126)(6);
p(212)(7)<=p(126)(7);
p(212)(8)<=p(126)(8);
p(212)(9)<=p(126)(9);
p(212)(10)<=p(126)(10);
p(212)(11)<=p(126)(11);
p(212)(12)<=p(126)(12);
p(212)(13)<=p(126)(13);
p(212)(14)<=p(126)(14);
p(212)(15)<=p(126)(15);
p(212)(16)<=p(126)(16);
p(212)(17)<=p(126)(17);
p(212)(18)<=p(126)(18);
p(212)(19)<=p(126)(19);
p(212)(20)<=p(126)(20);
p(212)(21)<=p(126)(21);
p(212)(22)<=p(126)(22);
p(212)(23)<=p(126)(23);
p(212)(24)<=p(126)(24);
p(212)(25)<=p(126)(25);
p(212)(26)<=p(126)(26);
p(212)(27)<=p(126)(27);
p(212)(28)<=p(126)(28);
p(212)(29)<=p(126)(29);
p(212)(30)<=p(126)(30);
p(212)(31)<=p(126)(31);
p(212)(32)<=p(126)(32);
p(212)(33)<=p(126)(33);
p(212)(34)<=p(126)(34);
p(212)(35)<=p(126)(35);
p(212)(36)<=p(126)(36);
p(212)(37)<=p(126)(37);
p(212)(38)<=p(126)(38);
p(212)(39)<=p(126)(39);
p(212)(40)<=p(126)(40);
p(212)(41)<=p(126)(41);
p(212)(42)<=p(126)(42);
p(212)(43)<=p(126)(43);
p(212)(44)<=p(126)(44);
p(212)(45)<=p(126)(45);
p(212)(46)<=p(126)(46);
p(212)(47)<=p(126)(47);
p(212)(48)<=p(126)(48);
p(212)(49)<=p(126)(49);
p(212)(50)<=p(126)(50);
p(212)(51)<=p(126)(51);
p(212)(52)<=p(126)(52);
p(212)(53)<=p(126)(53);
p(212)(54)<=p(126)(54);
p(212)(55)<=p(126)(55);
p(212)(56)<=p(126)(56);
p(212)(57)<=p(126)(57);
p(212)(58)<=p(126)(58);
p(212)(59)<=p(126)(59);
p(212)(60)<=p(126)(60);
p(212)(61)<=p(126)(61);
p(212)(62)<=p(126)(62);
p(212)(63)<=p(126)(63);
p(212)(64)<=p(126)(64);
p(212)(65)<=p(126)(65);
p(212)(66)<=p(126)(66);
p(212)(67)<=p(126)(67);
p(212)(68)<=p(126)(68);
p(212)(69)<=p(126)(69);
p(212)(70)<=p(126)(70);
p(212)(71)<=p(126)(71);
p(212)(72)<=p(126)(72);
p(212)(73)<=p(126)(73);
p(212)(74)<=p(126)(74);
p(212)(75)<=p(126)(75);
p(212)(76)<=p(126)(76);
p(212)(77)<=p(126)(77);
p(212)(78)<=p(126)(78);
p(212)(79)<=p(126)(79);
p(212)(80)<=p(126)(80);
p(212)(81)<=p(126)(81);
p(212)(82)<=p(126)(82);
p(212)(83)<=p(126)(83);
p(212)(84)<=p(126)(84);
p(212)(85)<=p(126)(85);
p(212)(86)<=p(126)(86);
p(212)(87)<=p(126)(87);
p(212)(88)<=p(126)(88);
p(212)(89)<=p(126)(89);
p(212)(90)<=p(126)(90);
p(212)(91)<=p(126)(91);
p(212)(92)<=p(126)(92);
p(212)(93)<=p(126)(93);
p(212)(94)<=p(126)(94);
p(212)(95)<=p(126)(95);
p(212)(96)<=p(126)(96);
p(212)(97)<=p(126)(97);
p(212)(98)<=p(126)(98);
p(212)(99)<=p(126)(99);
p(212)(100)<=p(126)(100);
p(212)(101)<=p(126)(101);
p(212)(102)<=p(126)(102);
p(212)(103)<=p(126)(103);
p(212)(104)<=p(126)(104);
p(212)(105)<=p(126)(105);
p(212)(106)<=p(126)(106);
p(212)(107)<=p(126)(107);
p(212)(108)<=p(126)(108);
p(212)(109)<=p(126)(109);
p(212)(110)<=p(126)(110);
p(212)(111)<=p(126)(111);
p(212)(112)<=p(126)(112);
p(212)(113)<=p(126)(113);
p(212)(114)<=p(126)(114);
p(212)(115)<=p(126)(115);
p(212)(116)<=p(126)(116);
p(212)(117)<=p(126)(117);
p(212)(118)<=p(126)(118);
p(212)(119)<=p(126)(119);
p(212)(120)<=p(126)(120);
p(212)(121)<=p(126)(121);
p(212)(122)<=p(126)(122);
p(212)(123)<=p(126)(123);
p(212)(124)<=p(126)(124);
p(212)(125)<=p(126)(125);
p(212)(126)<=p(126)(126);
p(212)(127)<=p(126)(127);
p(212)(128)<=p(126)(128);
p(212)(129)<=p(126)(129);
p(212)(130)<=p(126)(130);
p(212)(131)<=p(126)(131);
p(212)(132)<=p(126)(132);
p(212)(133)<=p(126)(133);
p(212)(134)<=p(126)(134);
p(213)(0)<=p(127)(0);
p(213)(1)<=p(127)(1);
p(213)(2)<=p(127)(2);
p(213)(3)<=p(127)(3);
p(213)(4)<=p(127)(4);
p(213)(5)<=p(127)(5);
p(213)(6)<=p(127)(6);
p(213)(7)<=p(127)(7);
p(213)(8)<=p(127)(8);
p(213)(9)<=p(127)(9);
p(213)(10)<=p(127)(10);
p(213)(11)<=p(127)(11);
p(213)(12)<=p(127)(12);
p(213)(13)<=p(127)(13);
p(213)(14)<=p(127)(14);
p(213)(15)<=p(127)(15);
p(213)(16)<=p(127)(16);
p(213)(17)<=p(127)(17);
p(213)(18)<=p(127)(18);
p(213)(19)<=p(127)(19);
p(213)(20)<=p(127)(20);
p(213)(21)<=p(127)(21);
p(213)(22)<=p(127)(22);
p(213)(23)<=p(127)(23);
p(213)(24)<=p(127)(24);
p(213)(25)<=p(127)(25);
p(213)(26)<=p(127)(26);
p(213)(27)<=p(127)(27);
p(213)(28)<=p(127)(28);
p(213)(29)<=p(127)(29);
p(213)(30)<=p(127)(30);
p(213)(31)<=p(127)(31);
p(213)(32)<=p(127)(32);
p(213)(33)<=p(127)(33);
p(213)(34)<=p(127)(34);
p(213)(35)<=p(127)(35);
p(213)(36)<=p(127)(36);
p(213)(37)<=p(127)(37);
p(213)(38)<=p(127)(38);
p(213)(39)<=p(127)(39);
p(213)(40)<=p(127)(40);
p(213)(41)<=p(127)(41);
p(213)(42)<=p(127)(42);
p(213)(43)<=p(127)(43);
p(213)(44)<=p(127)(44);
p(213)(45)<=p(127)(45);
p(213)(46)<=p(127)(46);
p(213)(47)<=p(127)(47);
p(213)(48)<=p(127)(48);
p(213)(49)<=p(127)(49);
p(213)(50)<=p(127)(50);
p(213)(51)<=p(127)(51);
p(213)(52)<=p(127)(52);
p(213)(53)<=p(127)(53);
p(213)(54)<=p(127)(54);
p(213)(55)<=p(127)(55);
p(213)(56)<=p(127)(56);
p(213)(57)<=p(127)(57);
p(213)(58)<=p(127)(58);
p(213)(59)<=p(127)(59);
p(213)(60)<=p(127)(60);
p(213)(61)<=p(127)(61);
p(213)(62)<=p(127)(62);
p(213)(63)<=p(127)(63);
p(213)(64)<=p(127)(64);
p(213)(65)<=p(127)(65);
p(213)(66)<=p(127)(66);
p(213)(67)<=p(127)(67);
p(213)(68)<=p(127)(68);
p(213)(69)<=p(127)(69);
p(213)(70)<=p(127)(70);
p(213)(71)<=p(127)(71);
p(213)(72)<=p(127)(72);
p(213)(73)<=p(127)(73);
p(213)(74)<=p(127)(74);
p(213)(75)<=p(127)(75);
p(213)(76)<=p(127)(76);
p(213)(77)<=p(127)(77);
p(213)(78)<=p(127)(78);
p(213)(79)<=p(127)(79);
p(213)(80)<=p(127)(80);
p(213)(81)<=p(127)(81);
p(213)(82)<=p(127)(82);
p(213)(83)<=p(127)(83);
p(213)(84)<=p(127)(84);
p(213)(85)<=p(127)(85);
p(213)(86)<=p(127)(86);
p(213)(87)<=p(127)(87);
p(213)(88)<=p(127)(88);
p(213)(89)<=p(127)(89);
p(213)(90)<=p(127)(90);
p(213)(91)<=p(127)(91);
p(213)(92)<=p(127)(92);
p(213)(93)<=p(127)(93);
p(213)(94)<=p(127)(94);
p(213)(95)<=p(127)(95);
p(213)(96)<=p(127)(96);
p(213)(97)<=p(127)(97);
p(213)(98)<=p(127)(98);
p(213)(99)<=p(127)(99);
p(213)(100)<=p(127)(100);
p(213)(101)<=p(127)(101);
p(213)(102)<=p(127)(102);
p(213)(103)<=p(127)(103);
p(213)(104)<=p(127)(104);
p(213)(105)<=p(127)(105);
p(213)(106)<=p(127)(106);
p(213)(107)<=p(127)(107);
p(213)(108)<=p(127)(108);
p(213)(109)<=p(127)(109);
p(213)(110)<=p(127)(110);
p(213)(111)<=p(127)(111);
p(213)(112)<=p(127)(112);
p(213)(113)<=p(127)(113);
p(213)(114)<=p(127)(114);
p(213)(115)<=p(127)(115);
p(213)(116)<=p(127)(116);
p(213)(117)<=p(127)(117);
p(213)(118)<=p(127)(118);
p(213)(119)<=p(127)(119);
p(213)(120)<=p(127)(120);
p(213)(121)<=p(127)(121);
p(213)(122)<=p(127)(122);
p(213)(123)<=p(127)(123);
p(213)(124)<=p(127)(124);
p(213)(125)<=p(127)(125);
p(213)(126)<=p(127)(126);
p(213)(127)<=p(127)(127);
p(213)(128)<=p(127)(128);
p(213)(129)<=p(127)(129);
p(213)(130)<=p(127)(130);
p(213)(131)<=p(127)(131);
p(213)(132)<=p(127)(132);
p(213)(133)<=p(127)(133);
p(213)(134)<=p(127)(134);
HA_ff_0:HAff port map(x=>p(128)(0),y=>p(130)(0),clock=>clock,reset=>reset,s=>p(214)(0),c=>p(215)(1));
FA_ff_5376:FAff port map(x=>p(128)(1),y=>p(129)(1),Cin=>p(130)(1),clock=>clock,reset=>reset,s=>p(214)(1),cout=>p(215)(2));
FA_ff_5377:FAff port map(x=>p(128)(2),y=>p(129)(2),Cin=>p(130)(2),clock=>clock,reset=>reset,s=>p(214)(2),cout=>p(215)(3));
FA_ff_5378:FAff port map(x=>p(128)(3),y=>p(129)(3),Cin=>p(130)(3),clock=>clock,reset=>reset,s=>p(214)(3),cout=>p(215)(4));
FA_ff_5379:FAff port map(x=>p(128)(4),y=>p(129)(4),Cin=>p(130)(4),clock=>clock,reset=>reset,s=>p(214)(4),cout=>p(215)(5));
FA_ff_5380:FAff port map(x=>p(128)(5),y=>p(129)(5),Cin=>p(130)(5),clock=>clock,reset=>reset,s=>p(214)(5),cout=>p(215)(6));
FA_ff_5381:FAff port map(x=>p(128)(6),y=>p(129)(6),Cin=>p(130)(6),clock=>clock,reset=>reset,s=>p(214)(6),cout=>p(215)(7));
FA_ff_5382:FAff port map(x=>p(128)(7),y=>p(129)(7),Cin=>p(130)(7),clock=>clock,reset=>reset,s=>p(214)(7),cout=>p(215)(8));
FA_ff_5383:FAff port map(x=>p(128)(8),y=>p(129)(8),Cin=>p(130)(8),clock=>clock,reset=>reset,s=>p(214)(8),cout=>p(215)(9));
FA_ff_5384:FAff port map(x=>p(128)(9),y=>p(129)(9),Cin=>p(130)(9),clock=>clock,reset=>reset,s=>p(214)(9),cout=>p(215)(10));
FA_ff_5385:FAff port map(x=>p(128)(10),y=>p(129)(10),Cin=>p(130)(10),clock=>clock,reset=>reset,s=>p(214)(10),cout=>p(215)(11));
FA_ff_5386:FAff port map(x=>p(128)(11),y=>p(129)(11),Cin=>p(130)(11),clock=>clock,reset=>reset,s=>p(214)(11),cout=>p(215)(12));
FA_ff_5387:FAff port map(x=>p(128)(12),y=>p(129)(12),Cin=>p(130)(12),clock=>clock,reset=>reset,s=>p(214)(12),cout=>p(215)(13));
FA_ff_5388:FAff port map(x=>p(128)(13),y=>p(129)(13),Cin=>p(130)(13),clock=>clock,reset=>reset,s=>p(214)(13),cout=>p(215)(14));
FA_ff_5389:FAff port map(x=>p(128)(14),y=>p(129)(14),Cin=>p(130)(14),clock=>clock,reset=>reset,s=>p(214)(14),cout=>p(215)(15));
FA_ff_5390:FAff port map(x=>p(128)(15),y=>p(129)(15),Cin=>p(130)(15),clock=>clock,reset=>reset,s=>p(214)(15),cout=>p(215)(16));
FA_ff_5391:FAff port map(x=>p(128)(16),y=>p(129)(16),Cin=>p(130)(16),clock=>clock,reset=>reset,s=>p(214)(16),cout=>p(215)(17));
FA_ff_5392:FAff port map(x=>p(128)(17),y=>p(129)(17),Cin=>p(130)(17),clock=>clock,reset=>reset,s=>p(214)(17),cout=>p(215)(18));
FA_ff_5393:FAff port map(x=>p(128)(18),y=>p(129)(18),Cin=>p(130)(18),clock=>clock,reset=>reset,s=>p(214)(18),cout=>p(215)(19));
FA_ff_5394:FAff port map(x=>p(128)(19),y=>p(129)(19),Cin=>p(130)(19),clock=>clock,reset=>reset,s=>p(214)(19),cout=>p(215)(20));
FA_ff_5395:FAff port map(x=>p(128)(20),y=>p(129)(20),Cin=>p(130)(20),clock=>clock,reset=>reset,s=>p(214)(20),cout=>p(215)(21));
FA_ff_5396:FAff port map(x=>p(128)(21),y=>p(129)(21),Cin=>p(130)(21),clock=>clock,reset=>reset,s=>p(214)(21),cout=>p(215)(22));
FA_ff_5397:FAff port map(x=>p(128)(22),y=>p(129)(22),Cin=>p(130)(22),clock=>clock,reset=>reset,s=>p(214)(22),cout=>p(215)(23));
FA_ff_5398:FAff port map(x=>p(128)(23),y=>p(129)(23),Cin=>p(130)(23),clock=>clock,reset=>reset,s=>p(214)(23),cout=>p(215)(24));
FA_ff_5399:FAff port map(x=>p(128)(24),y=>p(129)(24),Cin=>p(130)(24),clock=>clock,reset=>reset,s=>p(214)(24),cout=>p(215)(25));
FA_ff_5400:FAff port map(x=>p(128)(25),y=>p(129)(25),Cin=>p(130)(25),clock=>clock,reset=>reset,s=>p(214)(25),cout=>p(215)(26));
FA_ff_5401:FAff port map(x=>p(128)(26),y=>p(129)(26),Cin=>p(130)(26),clock=>clock,reset=>reset,s=>p(214)(26),cout=>p(215)(27));
FA_ff_5402:FAff port map(x=>p(128)(27),y=>p(129)(27),Cin=>p(130)(27),clock=>clock,reset=>reset,s=>p(214)(27),cout=>p(215)(28));
FA_ff_5403:FAff port map(x=>p(128)(28),y=>p(129)(28),Cin=>p(130)(28),clock=>clock,reset=>reset,s=>p(214)(28),cout=>p(215)(29));
FA_ff_5404:FAff port map(x=>p(128)(29),y=>p(129)(29),Cin=>p(130)(29),clock=>clock,reset=>reset,s=>p(214)(29),cout=>p(215)(30));
FA_ff_5405:FAff port map(x=>p(128)(30),y=>p(129)(30),Cin=>p(130)(30),clock=>clock,reset=>reset,s=>p(214)(30),cout=>p(215)(31));
FA_ff_5406:FAff port map(x=>p(128)(31),y=>p(129)(31),Cin=>p(130)(31),clock=>clock,reset=>reset,s=>p(214)(31),cout=>p(215)(32));
FA_ff_5407:FAff port map(x=>p(128)(32),y=>p(129)(32),Cin=>p(130)(32),clock=>clock,reset=>reset,s=>p(214)(32),cout=>p(215)(33));
FA_ff_5408:FAff port map(x=>p(128)(33),y=>p(129)(33),Cin=>p(130)(33),clock=>clock,reset=>reset,s=>p(214)(33),cout=>p(215)(34));
FA_ff_5409:FAff port map(x=>p(128)(34),y=>p(129)(34),Cin=>p(130)(34),clock=>clock,reset=>reset,s=>p(214)(34),cout=>p(215)(35));
FA_ff_5410:FAff port map(x=>p(128)(35),y=>p(129)(35),Cin=>p(130)(35),clock=>clock,reset=>reset,s=>p(214)(35),cout=>p(215)(36));
FA_ff_5411:FAff port map(x=>p(128)(36),y=>p(129)(36),Cin=>p(130)(36),clock=>clock,reset=>reset,s=>p(214)(36),cout=>p(215)(37));
FA_ff_5412:FAff port map(x=>p(128)(37),y=>p(129)(37),Cin=>p(130)(37),clock=>clock,reset=>reset,s=>p(214)(37),cout=>p(215)(38));
FA_ff_5413:FAff port map(x=>p(128)(38),y=>p(129)(38),Cin=>p(130)(38),clock=>clock,reset=>reset,s=>p(214)(38),cout=>p(215)(39));
FA_ff_5414:FAff port map(x=>p(128)(39),y=>p(129)(39),Cin=>p(130)(39),clock=>clock,reset=>reset,s=>p(214)(39),cout=>p(215)(40));
FA_ff_5415:FAff port map(x=>p(128)(40),y=>p(129)(40),Cin=>p(130)(40),clock=>clock,reset=>reset,s=>p(214)(40),cout=>p(215)(41));
FA_ff_5416:FAff port map(x=>p(128)(41),y=>p(129)(41),Cin=>p(130)(41),clock=>clock,reset=>reset,s=>p(214)(41),cout=>p(215)(42));
FA_ff_5417:FAff port map(x=>p(128)(42),y=>p(129)(42),Cin=>p(130)(42),clock=>clock,reset=>reset,s=>p(214)(42),cout=>p(215)(43));
FA_ff_5418:FAff port map(x=>p(128)(43),y=>p(129)(43),Cin=>p(130)(43),clock=>clock,reset=>reset,s=>p(214)(43),cout=>p(215)(44));
FA_ff_5419:FAff port map(x=>p(128)(44),y=>p(129)(44),Cin=>p(130)(44),clock=>clock,reset=>reset,s=>p(214)(44),cout=>p(215)(45));
FA_ff_5420:FAff port map(x=>p(128)(45),y=>p(129)(45),Cin=>p(130)(45),clock=>clock,reset=>reset,s=>p(214)(45),cout=>p(215)(46));
FA_ff_5421:FAff port map(x=>p(128)(46),y=>p(129)(46),Cin=>p(130)(46),clock=>clock,reset=>reset,s=>p(214)(46),cout=>p(215)(47));
FA_ff_5422:FAff port map(x=>p(128)(47),y=>p(129)(47),Cin=>p(130)(47),clock=>clock,reset=>reset,s=>p(214)(47),cout=>p(215)(48));
FA_ff_5423:FAff port map(x=>p(128)(48),y=>p(129)(48),Cin=>p(130)(48),clock=>clock,reset=>reset,s=>p(214)(48),cout=>p(215)(49));
FA_ff_5424:FAff port map(x=>p(128)(49),y=>p(129)(49),Cin=>p(130)(49),clock=>clock,reset=>reset,s=>p(214)(49),cout=>p(215)(50));
FA_ff_5425:FAff port map(x=>p(128)(50),y=>p(129)(50),Cin=>p(130)(50),clock=>clock,reset=>reset,s=>p(214)(50),cout=>p(215)(51));
FA_ff_5426:FAff port map(x=>p(128)(51),y=>p(129)(51),Cin=>p(130)(51),clock=>clock,reset=>reset,s=>p(214)(51),cout=>p(215)(52));
FA_ff_5427:FAff port map(x=>p(128)(52),y=>p(129)(52),Cin=>p(130)(52),clock=>clock,reset=>reset,s=>p(214)(52),cout=>p(215)(53));
FA_ff_5428:FAff port map(x=>p(128)(53),y=>p(129)(53),Cin=>p(130)(53),clock=>clock,reset=>reset,s=>p(214)(53),cout=>p(215)(54));
FA_ff_5429:FAff port map(x=>p(128)(54),y=>p(129)(54),Cin=>p(130)(54),clock=>clock,reset=>reset,s=>p(214)(54),cout=>p(215)(55));
FA_ff_5430:FAff port map(x=>p(128)(55),y=>p(129)(55),Cin=>p(130)(55),clock=>clock,reset=>reset,s=>p(214)(55),cout=>p(215)(56));
FA_ff_5431:FAff port map(x=>p(128)(56),y=>p(129)(56),Cin=>p(130)(56),clock=>clock,reset=>reset,s=>p(214)(56),cout=>p(215)(57));
FA_ff_5432:FAff port map(x=>p(128)(57),y=>p(129)(57),Cin=>p(130)(57),clock=>clock,reset=>reset,s=>p(214)(57),cout=>p(215)(58));
FA_ff_5433:FAff port map(x=>p(128)(58),y=>p(129)(58),Cin=>p(130)(58),clock=>clock,reset=>reset,s=>p(214)(58),cout=>p(215)(59));
FA_ff_5434:FAff port map(x=>p(128)(59),y=>p(129)(59),Cin=>p(130)(59),clock=>clock,reset=>reset,s=>p(214)(59),cout=>p(215)(60));
FA_ff_5435:FAff port map(x=>p(128)(60),y=>p(129)(60),Cin=>p(130)(60),clock=>clock,reset=>reset,s=>p(214)(60),cout=>p(215)(61));
FA_ff_5436:FAff port map(x=>p(128)(61),y=>p(129)(61),Cin=>p(130)(61),clock=>clock,reset=>reset,s=>p(214)(61),cout=>p(215)(62));
FA_ff_5437:FAff port map(x=>p(128)(62),y=>p(129)(62),Cin=>p(130)(62),clock=>clock,reset=>reset,s=>p(214)(62),cout=>p(215)(63));
FA_ff_5438:FAff port map(x=>p(128)(63),y=>p(129)(63),Cin=>p(130)(63),clock=>clock,reset=>reset,s=>p(214)(63),cout=>p(215)(64));
FA_ff_5439:FAff port map(x=>p(128)(64),y=>p(129)(64),Cin=>p(130)(64),clock=>clock,reset=>reset,s=>p(214)(64),cout=>p(215)(65));
FA_ff_5440:FAff port map(x=>p(128)(65),y=>p(129)(65),Cin=>p(130)(65),clock=>clock,reset=>reset,s=>p(214)(65),cout=>p(215)(66));
FA_ff_5441:FAff port map(x=>p(128)(66),y=>p(129)(66),Cin=>p(130)(66),clock=>clock,reset=>reset,s=>p(214)(66),cout=>p(215)(67));
FA_ff_5442:FAff port map(x=>p(128)(67),y=>p(129)(67),Cin=>p(130)(67),clock=>clock,reset=>reset,s=>p(214)(67),cout=>p(215)(68));
FA_ff_5443:FAff port map(x=>p(128)(68),y=>p(129)(68),Cin=>p(130)(68),clock=>clock,reset=>reset,s=>p(214)(68),cout=>p(215)(69));
FA_ff_5444:FAff port map(x=>p(128)(69),y=>p(129)(69),Cin=>p(130)(69),clock=>clock,reset=>reset,s=>p(214)(69),cout=>p(215)(70));
FA_ff_5445:FAff port map(x=>p(128)(70),y=>p(129)(70),Cin=>p(130)(70),clock=>clock,reset=>reset,s=>p(214)(70),cout=>p(215)(71));
FA_ff_5446:FAff port map(x=>p(128)(71),y=>p(129)(71),Cin=>p(130)(71),clock=>clock,reset=>reset,s=>p(214)(71),cout=>p(215)(72));
FA_ff_5447:FAff port map(x=>p(128)(72),y=>p(129)(72),Cin=>p(130)(72),clock=>clock,reset=>reset,s=>p(214)(72),cout=>p(215)(73));
FA_ff_5448:FAff port map(x=>p(128)(73),y=>p(129)(73),Cin=>p(130)(73),clock=>clock,reset=>reset,s=>p(214)(73),cout=>p(215)(74));
FA_ff_5449:FAff port map(x=>p(128)(74),y=>p(129)(74),Cin=>p(130)(74),clock=>clock,reset=>reset,s=>p(214)(74),cout=>p(215)(75));
FA_ff_5450:FAff port map(x=>p(128)(75),y=>p(129)(75),Cin=>p(130)(75),clock=>clock,reset=>reset,s=>p(214)(75),cout=>p(215)(76));
FA_ff_5451:FAff port map(x=>p(128)(76),y=>p(129)(76),Cin=>p(130)(76),clock=>clock,reset=>reset,s=>p(214)(76),cout=>p(215)(77));
FA_ff_5452:FAff port map(x=>p(128)(77),y=>p(129)(77),Cin=>p(130)(77),clock=>clock,reset=>reset,s=>p(214)(77),cout=>p(215)(78));
FA_ff_5453:FAff port map(x=>p(128)(78),y=>p(129)(78),Cin=>p(130)(78),clock=>clock,reset=>reset,s=>p(214)(78),cout=>p(215)(79));
FA_ff_5454:FAff port map(x=>p(128)(79),y=>p(129)(79),Cin=>p(130)(79),clock=>clock,reset=>reset,s=>p(214)(79),cout=>p(215)(80));
FA_ff_5455:FAff port map(x=>p(128)(80),y=>p(129)(80),Cin=>p(130)(80),clock=>clock,reset=>reset,s=>p(214)(80),cout=>p(215)(81));
FA_ff_5456:FAff port map(x=>p(128)(81),y=>p(129)(81),Cin=>p(130)(81),clock=>clock,reset=>reset,s=>p(214)(81),cout=>p(215)(82));
FA_ff_5457:FAff port map(x=>p(128)(82),y=>p(129)(82),Cin=>p(130)(82),clock=>clock,reset=>reset,s=>p(214)(82),cout=>p(215)(83));
FA_ff_5458:FAff port map(x=>p(128)(83),y=>p(129)(83),Cin=>p(130)(83),clock=>clock,reset=>reset,s=>p(214)(83),cout=>p(215)(84));
FA_ff_5459:FAff port map(x=>p(128)(84),y=>p(129)(84),Cin=>p(130)(84),clock=>clock,reset=>reset,s=>p(214)(84),cout=>p(215)(85));
FA_ff_5460:FAff port map(x=>p(128)(85),y=>p(129)(85),Cin=>p(130)(85),clock=>clock,reset=>reset,s=>p(214)(85),cout=>p(215)(86));
FA_ff_5461:FAff port map(x=>p(128)(86),y=>p(129)(86),Cin=>p(130)(86),clock=>clock,reset=>reset,s=>p(214)(86),cout=>p(215)(87));
FA_ff_5462:FAff port map(x=>p(128)(87),y=>p(129)(87),Cin=>p(130)(87),clock=>clock,reset=>reset,s=>p(214)(87),cout=>p(215)(88));
FA_ff_5463:FAff port map(x=>p(128)(88),y=>p(129)(88),Cin=>p(130)(88),clock=>clock,reset=>reset,s=>p(214)(88),cout=>p(215)(89));
FA_ff_5464:FAff port map(x=>p(128)(89),y=>p(129)(89),Cin=>p(130)(89),clock=>clock,reset=>reset,s=>p(214)(89),cout=>p(215)(90));
FA_ff_5465:FAff port map(x=>p(128)(90),y=>p(129)(90),Cin=>p(130)(90),clock=>clock,reset=>reset,s=>p(214)(90),cout=>p(215)(91));
FA_ff_5466:FAff port map(x=>p(128)(91),y=>p(129)(91),Cin=>p(130)(91),clock=>clock,reset=>reset,s=>p(214)(91),cout=>p(215)(92));
FA_ff_5467:FAff port map(x=>p(128)(92),y=>p(129)(92),Cin=>p(130)(92),clock=>clock,reset=>reset,s=>p(214)(92),cout=>p(215)(93));
FA_ff_5468:FAff port map(x=>p(128)(93),y=>p(129)(93),Cin=>p(130)(93),clock=>clock,reset=>reset,s=>p(214)(93),cout=>p(215)(94));
FA_ff_5469:FAff port map(x=>p(128)(94),y=>p(129)(94),Cin=>p(130)(94),clock=>clock,reset=>reset,s=>p(214)(94),cout=>p(215)(95));
FA_ff_5470:FAff port map(x=>p(128)(95),y=>p(129)(95),Cin=>p(130)(95),clock=>clock,reset=>reset,s=>p(214)(95),cout=>p(215)(96));
FA_ff_5471:FAff port map(x=>p(128)(96),y=>p(129)(96),Cin=>p(130)(96),clock=>clock,reset=>reset,s=>p(214)(96),cout=>p(215)(97));
FA_ff_5472:FAff port map(x=>p(128)(97),y=>p(129)(97),Cin=>p(130)(97),clock=>clock,reset=>reset,s=>p(214)(97),cout=>p(215)(98));
FA_ff_5473:FAff port map(x=>p(128)(98),y=>p(129)(98),Cin=>p(130)(98),clock=>clock,reset=>reset,s=>p(214)(98),cout=>p(215)(99));
FA_ff_5474:FAff port map(x=>p(128)(99),y=>p(129)(99),Cin=>p(130)(99),clock=>clock,reset=>reset,s=>p(214)(99),cout=>p(215)(100));
FA_ff_5475:FAff port map(x=>p(128)(100),y=>p(129)(100),Cin=>p(130)(100),clock=>clock,reset=>reset,s=>p(214)(100),cout=>p(215)(101));
FA_ff_5476:FAff port map(x=>p(128)(101),y=>p(129)(101),Cin=>p(130)(101),clock=>clock,reset=>reset,s=>p(214)(101),cout=>p(215)(102));
FA_ff_5477:FAff port map(x=>p(128)(102),y=>p(129)(102),Cin=>p(130)(102),clock=>clock,reset=>reset,s=>p(214)(102),cout=>p(215)(103));
FA_ff_5478:FAff port map(x=>p(128)(103),y=>p(129)(103),Cin=>p(130)(103),clock=>clock,reset=>reset,s=>p(214)(103),cout=>p(215)(104));
FA_ff_5479:FAff port map(x=>p(128)(104),y=>p(129)(104),Cin=>p(130)(104),clock=>clock,reset=>reset,s=>p(214)(104),cout=>p(215)(105));
FA_ff_5480:FAff port map(x=>p(128)(105),y=>p(129)(105),Cin=>p(130)(105),clock=>clock,reset=>reset,s=>p(214)(105),cout=>p(215)(106));
FA_ff_5481:FAff port map(x=>p(128)(106),y=>p(129)(106),Cin=>p(130)(106),clock=>clock,reset=>reset,s=>p(214)(106),cout=>p(215)(107));
FA_ff_5482:FAff port map(x=>p(128)(107),y=>p(129)(107),Cin=>p(130)(107),clock=>clock,reset=>reset,s=>p(214)(107),cout=>p(215)(108));
FA_ff_5483:FAff port map(x=>p(128)(108),y=>p(129)(108),Cin=>p(130)(108),clock=>clock,reset=>reset,s=>p(214)(108),cout=>p(215)(109));
FA_ff_5484:FAff port map(x=>p(128)(109),y=>p(129)(109),Cin=>p(130)(109),clock=>clock,reset=>reset,s=>p(214)(109),cout=>p(215)(110));
FA_ff_5485:FAff port map(x=>p(128)(110),y=>p(129)(110),Cin=>p(130)(110),clock=>clock,reset=>reset,s=>p(214)(110),cout=>p(215)(111));
FA_ff_5486:FAff port map(x=>p(128)(111),y=>p(129)(111),Cin=>p(130)(111),clock=>clock,reset=>reset,s=>p(214)(111),cout=>p(215)(112));
FA_ff_5487:FAff port map(x=>p(128)(112),y=>p(129)(112),Cin=>p(130)(112),clock=>clock,reset=>reset,s=>p(214)(112),cout=>p(215)(113));
FA_ff_5488:FAff port map(x=>p(128)(113),y=>p(129)(113),Cin=>p(130)(113),clock=>clock,reset=>reset,s=>p(214)(113),cout=>p(215)(114));
FA_ff_5489:FAff port map(x=>p(128)(114),y=>p(129)(114),Cin=>p(130)(114),clock=>clock,reset=>reset,s=>p(214)(114),cout=>p(215)(115));
FA_ff_5490:FAff port map(x=>p(128)(115),y=>p(129)(115),Cin=>p(130)(115),clock=>clock,reset=>reset,s=>p(214)(115),cout=>p(215)(116));
FA_ff_5491:FAff port map(x=>p(128)(116),y=>p(129)(116),Cin=>p(130)(116),clock=>clock,reset=>reset,s=>p(214)(116),cout=>p(215)(117));
FA_ff_5492:FAff port map(x=>p(128)(117),y=>p(129)(117),Cin=>p(130)(117),clock=>clock,reset=>reset,s=>p(214)(117),cout=>p(215)(118));
FA_ff_5493:FAff port map(x=>p(128)(118),y=>p(129)(118),Cin=>p(130)(118),clock=>clock,reset=>reset,s=>p(214)(118),cout=>p(215)(119));
FA_ff_5494:FAff port map(x=>p(128)(119),y=>p(129)(119),Cin=>p(130)(119),clock=>clock,reset=>reset,s=>p(214)(119),cout=>p(215)(120));
FA_ff_5495:FAff port map(x=>p(128)(120),y=>p(129)(120),Cin=>p(130)(120),clock=>clock,reset=>reset,s=>p(214)(120),cout=>p(215)(121));
FA_ff_5496:FAff port map(x=>p(128)(121),y=>p(129)(121),Cin=>p(130)(121),clock=>clock,reset=>reset,s=>p(214)(121),cout=>p(215)(122));
FA_ff_5497:FAff port map(x=>p(128)(122),y=>p(129)(122),Cin=>p(130)(122),clock=>clock,reset=>reset,s=>p(214)(122),cout=>p(215)(123));
FA_ff_5498:FAff port map(x=>p(128)(123),y=>p(129)(123),Cin=>p(130)(123),clock=>clock,reset=>reset,s=>p(214)(123),cout=>p(215)(124));
FA_ff_5499:FAff port map(x=>p(128)(124),y=>p(129)(124),Cin=>p(130)(124),clock=>clock,reset=>reset,s=>p(214)(124),cout=>p(215)(125));
FA_ff_5500:FAff port map(x=>p(128)(125),y=>p(129)(125),Cin=>p(130)(125),clock=>clock,reset=>reset,s=>p(214)(125),cout=>p(215)(126));
FA_ff_5501:FAff port map(x=>p(128)(126),y=>p(129)(126),Cin=>p(130)(126),clock=>clock,reset=>reset,s=>p(214)(126),cout=>p(215)(127));
FA_ff_5502:FAff port map(x=>p(128)(127),y=>p(129)(127),Cin=>p(130)(127),clock=>clock,reset=>reset,s=>p(214)(127),cout=>p(215)(128));
p(214)(128)<=p(129)(128);
p(216)(0)<=p(132)(0);
FA_ff_5503:FAff port map(x=>p(131)(1),y=>p(132)(1),Cin=>p(133)(1),clock=>clock,reset=>reset,s=>p(216)(1),cout=>p(217)(2));
FA_ff_5504:FAff port map(x=>p(131)(2),y=>p(132)(2),Cin=>p(133)(2),clock=>clock,reset=>reset,s=>p(216)(2),cout=>p(217)(3));
FA_ff_5505:FAff port map(x=>p(131)(3),y=>p(132)(3),Cin=>p(133)(3),clock=>clock,reset=>reset,s=>p(216)(3),cout=>p(217)(4));
FA_ff_5506:FAff port map(x=>p(131)(4),y=>p(132)(4),Cin=>p(133)(4),clock=>clock,reset=>reset,s=>p(216)(4),cout=>p(217)(5));
FA_ff_5507:FAff port map(x=>p(131)(5),y=>p(132)(5),Cin=>p(133)(5),clock=>clock,reset=>reset,s=>p(216)(5),cout=>p(217)(6));
FA_ff_5508:FAff port map(x=>p(131)(6),y=>p(132)(6),Cin=>p(133)(6),clock=>clock,reset=>reset,s=>p(216)(6),cout=>p(217)(7));
FA_ff_5509:FAff port map(x=>p(131)(7),y=>p(132)(7),Cin=>p(133)(7),clock=>clock,reset=>reset,s=>p(216)(7),cout=>p(217)(8));
FA_ff_5510:FAff port map(x=>p(131)(8),y=>p(132)(8),Cin=>p(133)(8),clock=>clock,reset=>reset,s=>p(216)(8),cout=>p(217)(9));
FA_ff_5511:FAff port map(x=>p(131)(9),y=>p(132)(9),Cin=>p(133)(9),clock=>clock,reset=>reset,s=>p(216)(9),cout=>p(217)(10));
FA_ff_5512:FAff port map(x=>p(131)(10),y=>p(132)(10),Cin=>p(133)(10),clock=>clock,reset=>reset,s=>p(216)(10),cout=>p(217)(11));
FA_ff_5513:FAff port map(x=>p(131)(11),y=>p(132)(11),Cin=>p(133)(11),clock=>clock,reset=>reset,s=>p(216)(11),cout=>p(217)(12));
FA_ff_5514:FAff port map(x=>p(131)(12),y=>p(132)(12),Cin=>p(133)(12),clock=>clock,reset=>reset,s=>p(216)(12),cout=>p(217)(13));
FA_ff_5515:FAff port map(x=>p(131)(13),y=>p(132)(13),Cin=>p(133)(13),clock=>clock,reset=>reset,s=>p(216)(13),cout=>p(217)(14));
FA_ff_5516:FAff port map(x=>p(131)(14),y=>p(132)(14),Cin=>p(133)(14),clock=>clock,reset=>reset,s=>p(216)(14),cout=>p(217)(15));
FA_ff_5517:FAff port map(x=>p(131)(15),y=>p(132)(15),Cin=>p(133)(15),clock=>clock,reset=>reset,s=>p(216)(15),cout=>p(217)(16));
FA_ff_5518:FAff port map(x=>p(131)(16),y=>p(132)(16),Cin=>p(133)(16),clock=>clock,reset=>reset,s=>p(216)(16),cout=>p(217)(17));
FA_ff_5519:FAff port map(x=>p(131)(17),y=>p(132)(17),Cin=>p(133)(17),clock=>clock,reset=>reset,s=>p(216)(17),cout=>p(217)(18));
FA_ff_5520:FAff port map(x=>p(131)(18),y=>p(132)(18),Cin=>p(133)(18),clock=>clock,reset=>reset,s=>p(216)(18),cout=>p(217)(19));
FA_ff_5521:FAff port map(x=>p(131)(19),y=>p(132)(19),Cin=>p(133)(19),clock=>clock,reset=>reset,s=>p(216)(19),cout=>p(217)(20));
FA_ff_5522:FAff port map(x=>p(131)(20),y=>p(132)(20),Cin=>p(133)(20),clock=>clock,reset=>reset,s=>p(216)(20),cout=>p(217)(21));
FA_ff_5523:FAff port map(x=>p(131)(21),y=>p(132)(21),Cin=>p(133)(21),clock=>clock,reset=>reset,s=>p(216)(21),cout=>p(217)(22));
FA_ff_5524:FAff port map(x=>p(131)(22),y=>p(132)(22),Cin=>p(133)(22),clock=>clock,reset=>reset,s=>p(216)(22),cout=>p(217)(23));
FA_ff_5525:FAff port map(x=>p(131)(23),y=>p(132)(23),Cin=>p(133)(23),clock=>clock,reset=>reset,s=>p(216)(23),cout=>p(217)(24));
FA_ff_5526:FAff port map(x=>p(131)(24),y=>p(132)(24),Cin=>p(133)(24),clock=>clock,reset=>reset,s=>p(216)(24),cout=>p(217)(25));
FA_ff_5527:FAff port map(x=>p(131)(25),y=>p(132)(25),Cin=>p(133)(25),clock=>clock,reset=>reset,s=>p(216)(25),cout=>p(217)(26));
FA_ff_5528:FAff port map(x=>p(131)(26),y=>p(132)(26),Cin=>p(133)(26),clock=>clock,reset=>reset,s=>p(216)(26),cout=>p(217)(27));
FA_ff_5529:FAff port map(x=>p(131)(27),y=>p(132)(27),Cin=>p(133)(27),clock=>clock,reset=>reset,s=>p(216)(27),cout=>p(217)(28));
FA_ff_5530:FAff port map(x=>p(131)(28),y=>p(132)(28),Cin=>p(133)(28),clock=>clock,reset=>reset,s=>p(216)(28),cout=>p(217)(29));
FA_ff_5531:FAff port map(x=>p(131)(29),y=>p(132)(29),Cin=>p(133)(29),clock=>clock,reset=>reset,s=>p(216)(29),cout=>p(217)(30));
FA_ff_5532:FAff port map(x=>p(131)(30),y=>p(132)(30),Cin=>p(133)(30),clock=>clock,reset=>reset,s=>p(216)(30),cout=>p(217)(31));
FA_ff_5533:FAff port map(x=>p(131)(31),y=>p(132)(31),Cin=>p(133)(31),clock=>clock,reset=>reset,s=>p(216)(31),cout=>p(217)(32));
FA_ff_5534:FAff port map(x=>p(131)(32),y=>p(132)(32),Cin=>p(133)(32),clock=>clock,reset=>reset,s=>p(216)(32),cout=>p(217)(33));
FA_ff_5535:FAff port map(x=>p(131)(33),y=>p(132)(33),Cin=>p(133)(33),clock=>clock,reset=>reset,s=>p(216)(33),cout=>p(217)(34));
FA_ff_5536:FAff port map(x=>p(131)(34),y=>p(132)(34),Cin=>p(133)(34),clock=>clock,reset=>reset,s=>p(216)(34),cout=>p(217)(35));
FA_ff_5537:FAff port map(x=>p(131)(35),y=>p(132)(35),Cin=>p(133)(35),clock=>clock,reset=>reset,s=>p(216)(35),cout=>p(217)(36));
FA_ff_5538:FAff port map(x=>p(131)(36),y=>p(132)(36),Cin=>p(133)(36),clock=>clock,reset=>reset,s=>p(216)(36),cout=>p(217)(37));
FA_ff_5539:FAff port map(x=>p(131)(37),y=>p(132)(37),Cin=>p(133)(37),clock=>clock,reset=>reset,s=>p(216)(37),cout=>p(217)(38));
FA_ff_5540:FAff port map(x=>p(131)(38),y=>p(132)(38),Cin=>p(133)(38),clock=>clock,reset=>reset,s=>p(216)(38),cout=>p(217)(39));
FA_ff_5541:FAff port map(x=>p(131)(39),y=>p(132)(39),Cin=>p(133)(39),clock=>clock,reset=>reset,s=>p(216)(39),cout=>p(217)(40));
FA_ff_5542:FAff port map(x=>p(131)(40),y=>p(132)(40),Cin=>p(133)(40),clock=>clock,reset=>reset,s=>p(216)(40),cout=>p(217)(41));
FA_ff_5543:FAff port map(x=>p(131)(41),y=>p(132)(41),Cin=>p(133)(41),clock=>clock,reset=>reset,s=>p(216)(41),cout=>p(217)(42));
FA_ff_5544:FAff port map(x=>p(131)(42),y=>p(132)(42),Cin=>p(133)(42),clock=>clock,reset=>reset,s=>p(216)(42),cout=>p(217)(43));
FA_ff_5545:FAff port map(x=>p(131)(43),y=>p(132)(43),Cin=>p(133)(43),clock=>clock,reset=>reset,s=>p(216)(43),cout=>p(217)(44));
FA_ff_5546:FAff port map(x=>p(131)(44),y=>p(132)(44),Cin=>p(133)(44),clock=>clock,reset=>reset,s=>p(216)(44),cout=>p(217)(45));
FA_ff_5547:FAff port map(x=>p(131)(45),y=>p(132)(45),Cin=>p(133)(45),clock=>clock,reset=>reset,s=>p(216)(45),cout=>p(217)(46));
FA_ff_5548:FAff port map(x=>p(131)(46),y=>p(132)(46),Cin=>p(133)(46),clock=>clock,reset=>reset,s=>p(216)(46),cout=>p(217)(47));
FA_ff_5549:FAff port map(x=>p(131)(47),y=>p(132)(47),Cin=>p(133)(47),clock=>clock,reset=>reset,s=>p(216)(47),cout=>p(217)(48));
FA_ff_5550:FAff port map(x=>p(131)(48),y=>p(132)(48),Cin=>p(133)(48),clock=>clock,reset=>reset,s=>p(216)(48),cout=>p(217)(49));
FA_ff_5551:FAff port map(x=>p(131)(49),y=>p(132)(49),Cin=>p(133)(49),clock=>clock,reset=>reset,s=>p(216)(49),cout=>p(217)(50));
FA_ff_5552:FAff port map(x=>p(131)(50),y=>p(132)(50),Cin=>p(133)(50),clock=>clock,reset=>reset,s=>p(216)(50),cout=>p(217)(51));
FA_ff_5553:FAff port map(x=>p(131)(51),y=>p(132)(51),Cin=>p(133)(51),clock=>clock,reset=>reset,s=>p(216)(51),cout=>p(217)(52));
FA_ff_5554:FAff port map(x=>p(131)(52),y=>p(132)(52),Cin=>p(133)(52),clock=>clock,reset=>reset,s=>p(216)(52),cout=>p(217)(53));
FA_ff_5555:FAff port map(x=>p(131)(53),y=>p(132)(53),Cin=>p(133)(53),clock=>clock,reset=>reset,s=>p(216)(53),cout=>p(217)(54));
FA_ff_5556:FAff port map(x=>p(131)(54),y=>p(132)(54),Cin=>p(133)(54),clock=>clock,reset=>reset,s=>p(216)(54),cout=>p(217)(55));
FA_ff_5557:FAff port map(x=>p(131)(55),y=>p(132)(55),Cin=>p(133)(55),clock=>clock,reset=>reset,s=>p(216)(55),cout=>p(217)(56));
FA_ff_5558:FAff port map(x=>p(131)(56),y=>p(132)(56),Cin=>p(133)(56),clock=>clock,reset=>reset,s=>p(216)(56),cout=>p(217)(57));
FA_ff_5559:FAff port map(x=>p(131)(57),y=>p(132)(57),Cin=>p(133)(57),clock=>clock,reset=>reset,s=>p(216)(57),cout=>p(217)(58));
FA_ff_5560:FAff port map(x=>p(131)(58),y=>p(132)(58),Cin=>p(133)(58),clock=>clock,reset=>reset,s=>p(216)(58),cout=>p(217)(59));
FA_ff_5561:FAff port map(x=>p(131)(59),y=>p(132)(59),Cin=>p(133)(59),clock=>clock,reset=>reset,s=>p(216)(59),cout=>p(217)(60));
FA_ff_5562:FAff port map(x=>p(131)(60),y=>p(132)(60),Cin=>p(133)(60),clock=>clock,reset=>reset,s=>p(216)(60),cout=>p(217)(61));
FA_ff_5563:FAff port map(x=>p(131)(61),y=>p(132)(61),Cin=>p(133)(61),clock=>clock,reset=>reset,s=>p(216)(61),cout=>p(217)(62));
FA_ff_5564:FAff port map(x=>p(131)(62),y=>p(132)(62),Cin=>p(133)(62),clock=>clock,reset=>reset,s=>p(216)(62),cout=>p(217)(63));
FA_ff_5565:FAff port map(x=>p(131)(63),y=>p(132)(63),Cin=>p(133)(63),clock=>clock,reset=>reset,s=>p(216)(63),cout=>p(217)(64));
FA_ff_5566:FAff port map(x=>p(131)(64),y=>p(132)(64),Cin=>p(133)(64),clock=>clock,reset=>reset,s=>p(216)(64),cout=>p(217)(65));
FA_ff_5567:FAff port map(x=>p(131)(65),y=>p(132)(65),Cin=>p(133)(65),clock=>clock,reset=>reset,s=>p(216)(65),cout=>p(217)(66));
FA_ff_5568:FAff port map(x=>p(131)(66),y=>p(132)(66),Cin=>p(133)(66),clock=>clock,reset=>reset,s=>p(216)(66),cout=>p(217)(67));
FA_ff_5569:FAff port map(x=>p(131)(67),y=>p(132)(67),Cin=>p(133)(67),clock=>clock,reset=>reset,s=>p(216)(67),cout=>p(217)(68));
FA_ff_5570:FAff port map(x=>p(131)(68),y=>p(132)(68),Cin=>p(133)(68),clock=>clock,reset=>reset,s=>p(216)(68),cout=>p(217)(69));
FA_ff_5571:FAff port map(x=>p(131)(69),y=>p(132)(69),Cin=>p(133)(69),clock=>clock,reset=>reset,s=>p(216)(69),cout=>p(217)(70));
FA_ff_5572:FAff port map(x=>p(131)(70),y=>p(132)(70),Cin=>p(133)(70),clock=>clock,reset=>reset,s=>p(216)(70),cout=>p(217)(71));
FA_ff_5573:FAff port map(x=>p(131)(71),y=>p(132)(71),Cin=>p(133)(71),clock=>clock,reset=>reset,s=>p(216)(71),cout=>p(217)(72));
FA_ff_5574:FAff port map(x=>p(131)(72),y=>p(132)(72),Cin=>p(133)(72),clock=>clock,reset=>reset,s=>p(216)(72),cout=>p(217)(73));
FA_ff_5575:FAff port map(x=>p(131)(73),y=>p(132)(73),Cin=>p(133)(73),clock=>clock,reset=>reset,s=>p(216)(73),cout=>p(217)(74));
FA_ff_5576:FAff port map(x=>p(131)(74),y=>p(132)(74),Cin=>p(133)(74),clock=>clock,reset=>reset,s=>p(216)(74),cout=>p(217)(75));
FA_ff_5577:FAff port map(x=>p(131)(75),y=>p(132)(75),Cin=>p(133)(75),clock=>clock,reset=>reset,s=>p(216)(75),cout=>p(217)(76));
FA_ff_5578:FAff port map(x=>p(131)(76),y=>p(132)(76),Cin=>p(133)(76),clock=>clock,reset=>reset,s=>p(216)(76),cout=>p(217)(77));
FA_ff_5579:FAff port map(x=>p(131)(77),y=>p(132)(77),Cin=>p(133)(77),clock=>clock,reset=>reset,s=>p(216)(77),cout=>p(217)(78));
FA_ff_5580:FAff port map(x=>p(131)(78),y=>p(132)(78),Cin=>p(133)(78),clock=>clock,reset=>reset,s=>p(216)(78),cout=>p(217)(79));
FA_ff_5581:FAff port map(x=>p(131)(79),y=>p(132)(79),Cin=>p(133)(79),clock=>clock,reset=>reset,s=>p(216)(79),cout=>p(217)(80));
FA_ff_5582:FAff port map(x=>p(131)(80),y=>p(132)(80),Cin=>p(133)(80),clock=>clock,reset=>reset,s=>p(216)(80),cout=>p(217)(81));
FA_ff_5583:FAff port map(x=>p(131)(81),y=>p(132)(81),Cin=>p(133)(81),clock=>clock,reset=>reset,s=>p(216)(81),cout=>p(217)(82));
FA_ff_5584:FAff port map(x=>p(131)(82),y=>p(132)(82),Cin=>p(133)(82),clock=>clock,reset=>reset,s=>p(216)(82),cout=>p(217)(83));
FA_ff_5585:FAff port map(x=>p(131)(83),y=>p(132)(83),Cin=>p(133)(83),clock=>clock,reset=>reset,s=>p(216)(83),cout=>p(217)(84));
FA_ff_5586:FAff port map(x=>p(131)(84),y=>p(132)(84),Cin=>p(133)(84),clock=>clock,reset=>reset,s=>p(216)(84),cout=>p(217)(85));
FA_ff_5587:FAff port map(x=>p(131)(85),y=>p(132)(85),Cin=>p(133)(85),clock=>clock,reset=>reset,s=>p(216)(85),cout=>p(217)(86));
FA_ff_5588:FAff port map(x=>p(131)(86),y=>p(132)(86),Cin=>p(133)(86),clock=>clock,reset=>reset,s=>p(216)(86),cout=>p(217)(87));
FA_ff_5589:FAff port map(x=>p(131)(87),y=>p(132)(87),Cin=>p(133)(87),clock=>clock,reset=>reset,s=>p(216)(87),cout=>p(217)(88));
FA_ff_5590:FAff port map(x=>p(131)(88),y=>p(132)(88),Cin=>p(133)(88),clock=>clock,reset=>reset,s=>p(216)(88),cout=>p(217)(89));
FA_ff_5591:FAff port map(x=>p(131)(89),y=>p(132)(89),Cin=>p(133)(89),clock=>clock,reset=>reset,s=>p(216)(89),cout=>p(217)(90));
FA_ff_5592:FAff port map(x=>p(131)(90),y=>p(132)(90),Cin=>p(133)(90),clock=>clock,reset=>reset,s=>p(216)(90),cout=>p(217)(91));
FA_ff_5593:FAff port map(x=>p(131)(91),y=>p(132)(91),Cin=>p(133)(91),clock=>clock,reset=>reset,s=>p(216)(91),cout=>p(217)(92));
FA_ff_5594:FAff port map(x=>p(131)(92),y=>p(132)(92),Cin=>p(133)(92),clock=>clock,reset=>reset,s=>p(216)(92),cout=>p(217)(93));
FA_ff_5595:FAff port map(x=>p(131)(93),y=>p(132)(93),Cin=>p(133)(93),clock=>clock,reset=>reset,s=>p(216)(93),cout=>p(217)(94));
FA_ff_5596:FAff port map(x=>p(131)(94),y=>p(132)(94),Cin=>p(133)(94),clock=>clock,reset=>reset,s=>p(216)(94),cout=>p(217)(95));
FA_ff_5597:FAff port map(x=>p(131)(95),y=>p(132)(95),Cin=>p(133)(95),clock=>clock,reset=>reset,s=>p(216)(95),cout=>p(217)(96));
FA_ff_5598:FAff port map(x=>p(131)(96),y=>p(132)(96),Cin=>p(133)(96),clock=>clock,reset=>reset,s=>p(216)(96),cout=>p(217)(97));
FA_ff_5599:FAff port map(x=>p(131)(97),y=>p(132)(97),Cin=>p(133)(97),clock=>clock,reset=>reset,s=>p(216)(97),cout=>p(217)(98));
FA_ff_5600:FAff port map(x=>p(131)(98),y=>p(132)(98),Cin=>p(133)(98),clock=>clock,reset=>reset,s=>p(216)(98),cout=>p(217)(99));
FA_ff_5601:FAff port map(x=>p(131)(99),y=>p(132)(99),Cin=>p(133)(99),clock=>clock,reset=>reset,s=>p(216)(99),cout=>p(217)(100));
FA_ff_5602:FAff port map(x=>p(131)(100),y=>p(132)(100),Cin=>p(133)(100),clock=>clock,reset=>reset,s=>p(216)(100),cout=>p(217)(101));
FA_ff_5603:FAff port map(x=>p(131)(101),y=>p(132)(101),Cin=>p(133)(101),clock=>clock,reset=>reset,s=>p(216)(101),cout=>p(217)(102));
FA_ff_5604:FAff port map(x=>p(131)(102),y=>p(132)(102),Cin=>p(133)(102),clock=>clock,reset=>reset,s=>p(216)(102),cout=>p(217)(103));
FA_ff_5605:FAff port map(x=>p(131)(103),y=>p(132)(103),Cin=>p(133)(103),clock=>clock,reset=>reset,s=>p(216)(103),cout=>p(217)(104));
FA_ff_5606:FAff port map(x=>p(131)(104),y=>p(132)(104),Cin=>p(133)(104),clock=>clock,reset=>reset,s=>p(216)(104),cout=>p(217)(105));
FA_ff_5607:FAff port map(x=>p(131)(105),y=>p(132)(105),Cin=>p(133)(105),clock=>clock,reset=>reset,s=>p(216)(105),cout=>p(217)(106));
FA_ff_5608:FAff port map(x=>p(131)(106),y=>p(132)(106),Cin=>p(133)(106),clock=>clock,reset=>reset,s=>p(216)(106),cout=>p(217)(107));
FA_ff_5609:FAff port map(x=>p(131)(107),y=>p(132)(107),Cin=>p(133)(107),clock=>clock,reset=>reset,s=>p(216)(107),cout=>p(217)(108));
FA_ff_5610:FAff port map(x=>p(131)(108),y=>p(132)(108),Cin=>p(133)(108),clock=>clock,reset=>reset,s=>p(216)(108),cout=>p(217)(109));
FA_ff_5611:FAff port map(x=>p(131)(109),y=>p(132)(109),Cin=>p(133)(109),clock=>clock,reset=>reset,s=>p(216)(109),cout=>p(217)(110));
FA_ff_5612:FAff port map(x=>p(131)(110),y=>p(132)(110),Cin=>p(133)(110),clock=>clock,reset=>reset,s=>p(216)(110),cout=>p(217)(111));
FA_ff_5613:FAff port map(x=>p(131)(111),y=>p(132)(111),Cin=>p(133)(111),clock=>clock,reset=>reset,s=>p(216)(111),cout=>p(217)(112));
FA_ff_5614:FAff port map(x=>p(131)(112),y=>p(132)(112),Cin=>p(133)(112),clock=>clock,reset=>reset,s=>p(216)(112),cout=>p(217)(113));
FA_ff_5615:FAff port map(x=>p(131)(113),y=>p(132)(113),Cin=>p(133)(113),clock=>clock,reset=>reset,s=>p(216)(113),cout=>p(217)(114));
FA_ff_5616:FAff port map(x=>p(131)(114),y=>p(132)(114),Cin=>p(133)(114),clock=>clock,reset=>reset,s=>p(216)(114),cout=>p(217)(115));
FA_ff_5617:FAff port map(x=>p(131)(115),y=>p(132)(115),Cin=>p(133)(115),clock=>clock,reset=>reset,s=>p(216)(115),cout=>p(217)(116));
FA_ff_5618:FAff port map(x=>p(131)(116),y=>p(132)(116),Cin=>p(133)(116),clock=>clock,reset=>reset,s=>p(216)(116),cout=>p(217)(117));
FA_ff_5619:FAff port map(x=>p(131)(117),y=>p(132)(117),Cin=>p(133)(117),clock=>clock,reset=>reset,s=>p(216)(117),cout=>p(217)(118));
FA_ff_5620:FAff port map(x=>p(131)(118),y=>p(132)(118),Cin=>p(133)(118),clock=>clock,reset=>reset,s=>p(216)(118),cout=>p(217)(119));
FA_ff_5621:FAff port map(x=>p(131)(119),y=>p(132)(119),Cin=>p(133)(119),clock=>clock,reset=>reset,s=>p(216)(119),cout=>p(217)(120));
FA_ff_5622:FAff port map(x=>p(131)(120),y=>p(132)(120),Cin=>p(133)(120),clock=>clock,reset=>reset,s=>p(216)(120),cout=>p(217)(121));
FA_ff_5623:FAff port map(x=>p(131)(121),y=>p(132)(121),Cin=>p(133)(121),clock=>clock,reset=>reset,s=>p(216)(121),cout=>p(217)(122));
FA_ff_5624:FAff port map(x=>p(131)(122),y=>p(132)(122),Cin=>p(133)(122),clock=>clock,reset=>reset,s=>p(216)(122),cout=>p(217)(123));
FA_ff_5625:FAff port map(x=>p(131)(123),y=>p(132)(123),Cin=>p(133)(123),clock=>clock,reset=>reset,s=>p(216)(123),cout=>p(217)(124));
FA_ff_5626:FAff port map(x=>p(131)(124),y=>p(132)(124),Cin=>p(133)(124),clock=>clock,reset=>reset,s=>p(216)(124),cout=>p(217)(125));
FA_ff_5627:FAff port map(x=>p(131)(125),y=>p(132)(125),Cin=>p(133)(125),clock=>clock,reset=>reset,s=>p(216)(125),cout=>p(217)(126));
FA_ff_5628:FAff port map(x=>p(131)(126),y=>p(132)(126),Cin=>p(133)(126),clock=>clock,reset=>reset,s=>p(216)(126),cout=>p(217)(127));
FA_ff_5629:FAff port map(x=>p(131)(127),y=>p(132)(127),Cin=>p(133)(127),clock=>clock,reset=>reset,s=>p(216)(127),cout=>p(217)(128));
HA_ff_1:HAff port map(x=>p(131)(128),y=>p(133)(128),clock=>clock,reset=>reset,s=>p(216)(128),c=>p(217)(129));
HA_ff_2:HAff port map(x=>p(134)(0),y=>p(136)(0),clock=>clock,reset=>reset,s=>p(218)(0),c=>p(219)(1));
FA_ff_5630:FAff port map(x=>p(134)(1),y=>p(135)(1),Cin=>p(136)(1),clock=>clock,reset=>reset,s=>p(218)(1),cout=>p(219)(2));
FA_ff_5631:FAff port map(x=>p(134)(2),y=>p(135)(2),Cin=>p(136)(2),clock=>clock,reset=>reset,s=>p(218)(2),cout=>p(219)(3));
FA_ff_5632:FAff port map(x=>p(134)(3),y=>p(135)(3),Cin=>p(136)(3),clock=>clock,reset=>reset,s=>p(218)(3),cout=>p(219)(4));
FA_ff_5633:FAff port map(x=>p(134)(4),y=>p(135)(4),Cin=>p(136)(4),clock=>clock,reset=>reset,s=>p(218)(4),cout=>p(219)(5));
FA_ff_5634:FAff port map(x=>p(134)(5),y=>p(135)(5),Cin=>p(136)(5),clock=>clock,reset=>reset,s=>p(218)(5),cout=>p(219)(6));
FA_ff_5635:FAff port map(x=>p(134)(6),y=>p(135)(6),Cin=>p(136)(6),clock=>clock,reset=>reset,s=>p(218)(6),cout=>p(219)(7));
FA_ff_5636:FAff port map(x=>p(134)(7),y=>p(135)(7),Cin=>p(136)(7),clock=>clock,reset=>reset,s=>p(218)(7),cout=>p(219)(8));
FA_ff_5637:FAff port map(x=>p(134)(8),y=>p(135)(8),Cin=>p(136)(8),clock=>clock,reset=>reset,s=>p(218)(8),cout=>p(219)(9));
FA_ff_5638:FAff port map(x=>p(134)(9),y=>p(135)(9),Cin=>p(136)(9),clock=>clock,reset=>reset,s=>p(218)(9),cout=>p(219)(10));
FA_ff_5639:FAff port map(x=>p(134)(10),y=>p(135)(10),Cin=>p(136)(10),clock=>clock,reset=>reset,s=>p(218)(10),cout=>p(219)(11));
FA_ff_5640:FAff port map(x=>p(134)(11),y=>p(135)(11),Cin=>p(136)(11),clock=>clock,reset=>reset,s=>p(218)(11),cout=>p(219)(12));
FA_ff_5641:FAff port map(x=>p(134)(12),y=>p(135)(12),Cin=>p(136)(12),clock=>clock,reset=>reset,s=>p(218)(12),cout=>p(219)(13));
FA_ff_5642:FAff port map(x=>p(134)(13),y=>p(135)(13),Cin=>p(136)(13),clock=>clock,reset=>reset,s=>p(218)(13),cout=>p(219)(14));
FA_ff_5643:FAff port map(x=>p(134)(14),y=>p(135)(14),Cin=>p(136)(14),clock=>clock,reset=>reset,s=>p(218)(14),cout=>p(219)(15));
FA_ff_5644:FAff port map(x=>p(134)(15),y=>p(135)(15),Cin=>p(136)(15),clock=>clock,reset=>reset,s=>p(218)(15),cout=>p(219)(16));
FA_ff_5645:FAff port map(x=>p(134)(16),y=>p(135)(16),Cin=>p(136)(16),clock=>clock,reset=>reset,s=>p(218)(16),cout=>p(219)(17));
FA_ff_5646:FAff port map(x=>p(134)(17),y=>p(135)(17),Cin=>p(136)(17),clock=>clock,reset=>reset,s=>p(218)(17),cout=>p(219)(18));
FA_ff_5647:FAff port map(x=>p(134)(18),y=>p(135)(18),Cin=>p(136)(18),clock=>clock,reset=>reset,s=>p(218)(18),cout=>p(219)(19));
FA_ff_5648:FAff port map(x=>p(134)(19),y=>p(135)(19),Cin=>p(136)(19),clock=>clock,reset=>reset,s=>p(218)(19),cout=>p(219)(20));
FA_ff_5649:FAff port map(x=>p(134)(20),y=>p(135)(20),Cin=>p(136)(20),clock=>clock,reset=>reset,s=>p(218)(20),cout=>p(219)(21));
FA_ff_5650:FAff port map(x=>p(134)(21),y=>p(135)(21),Cin=>p(136)(21),clock=>clock,reset=>reset,s=>p(218)(21),cout=>p(219)(22));
FA_ff_5651:FAff port map(x=>p(134)(22),y=>p(135)(22),Cin=>p(136)(22),clock=>clock,reset=>reset,s=>p(218)(22),cout=>p(219)(23));
FA_ff_5652:FAff port map(x=>p(134)(23),y=>p(135)(23),Cin=>p(136)(23),clock=>clock,reset=>reset,s=>p(218)(23),cout=>p(219)(24));
FA_ff_5653:FAff port map(x=>p(134)(24),y=>p(135)(24),Cin=>p(136)(24),clock=>clock,reset=>reset,s=>p(218)(24),cout=>p(219)(25));
FA_ff_5654:FAff port map(x=>p(134)(25),y=>p(135)(25),Cin=>p(136)(25),clock=>clock,reset=>reset,s=>p(218)(25),cout=>p(219)(26));
FA_ff_5655:FAff port map(x=>p(134)(26),y=>p(135)(26),Cin=>p(136)(26),clock=>clock,reset=>reset,s=>p(218)(26),cout=>p(219)(27));
FA_ff_5656:FAff port map(x=>p(134)(27),y=>p(135)(27),Cin=>p(136)(27),clock=>clock,reset=>reset,s=>p(218)(27),cout=>p(219)(28));
FA_ff_5657:FAff port map(x=>p(134)(28),y=>p(135)(28),Cin=>p(136)(28),clock=>clock,reset=>reset,s=>p(218)(28),cout=>p(219)(29));
FA_ff_5658:FAff port map(x=>p(134)(29),y=>p(135)(29),Cin=>p(136)(29),clock=>clock,reset=>reset,s=>p(218)(29),cout=>p(219)(30));
FA_ff_5659:FAff port map(x=>p(134)(30),y=>p(135)(30),Cin=>p(136)(30),clock=>clock,reset=>reset,s=>p(218)(30),cout=>p(219)(31));
FA_ff_5660:FAff port map(x=>p(134)(31),y=>p(135)(31),Cin=>p(136)(31),clock=>clock,reset=>reset,s=>p(218)(31),cout=>p(219)(32));
FA_ff_5661:FAff port map(x=>p(134)(32),y=>p(135)(32),Cin=>p(136)(32),clock=>clock,reset=>reset,s=>p(218)(32),cout=>p(219)(33));
FA_ff_5662:FAff port map(x=>p(134)(33),y=>p(135)(33),Cin=>p(136)(33),clock=>clock,reset=>reset,s=>p(218)(33),cout=>p(219)(34));
FA_ff_5663:FAff port map(x=>p(134)(34),y=>p(135)(34),Cin=>p(136)(34),clock=>clock,reset=>reset,s=>p(218)(34),cout=>p(219)(35));
FA_ff_5664:FAff port map(x=>p(134)(35),y=>p(135)(35),Cin=>p(136)(35),clock=>clock,reset=>reset,s=>p(218)(35),cout=>p(219)(36));
FA_ff_5665:FAff port map(x=>p(134)(36),y=>p(135)(36),Cin=>p(136)(36),clock=>clock,reset=>reset,s=>p(218)(36),cout=>p(219)(37));
FA_ff_5666:FAff port map(x=>p(134)(37),y=>p(135)(37),Cin=>p(136)(37),clock=>clock,reset=>reset,s=>p(218)(37),cout=>p(219)(38));
FA_ff_5667:FAff port map(x=>p(134)(38),y=>p(135)(38),Cin=>p(136)(38),clock=>clock,reset=>reset,s=>p(218)(38),cout=>p(219)(39));
FA_ff_5668:FAff port map(x=>p(134)(39),y=>p(135)(39),Cin=>p(136)(39),clock=>clock,reset=>reset,s=>p(218)(39),cout=>p(219)(40));
FA_ff_5669:FAff port map(x=>p(134)(40),y=>p(135)(40),Cin=>p(136)(40),clock=>clock,reset=>reset,s=>p(218)(40),cout=>p(219)(41));
FA_ff_5670:FAff port map(x=>p(134)(41),y=>p(135)(41),Cin=>p(136)(41),clock=>clock,reset=>reset,s=>p(218)(41),cout=>p(219)(42));
FA_ff_5671:FAff port map(x=>p(134)(42),y=>p(135)(42),Cin=>p(136)(42),clock=>clock,reset=>reset,s=>p(218)(42),cout=>p(219)(43));
FA_ff_5672:FAff port map(x=>p(134)(43),y=>p(135)(43),Cin=>p(136)(43),clock=>clock,reset=>reset,s=>p(218)(43),cout=>p(219)(44));
FA_ff_5673:FAff port map(x=>p(134)(44),y=>p(135)(44),Cin=>p(136)(44),clock=>clock,reset=>reset,s=>p(218)(44),cout=>p(219)(45));
FA_ff_5674:FAff port map(x=>p(134)(45),y=>p(135)(45),Cin=>p(136)(45),clock=>clock,reset=>reset,s=>p(218)(45),cout=>p(219)(46));
FA_ff_5675:FAff port map(x=>p(134)(46),y=>p(135)(46),Cin=>p(136)(46),clock=>clock,reset=>reset,s=>p(218)(46),cout=>p(219)(47));
FA_ff_5676:FAff port map(x=>p(134)(47),y=>p(135)(47),Cin=>p(136)(47),clock=>clock,reset=>reset,s=>p(218)(47),cout=>p(219)(48));
FA_ff_5677:FAff port map(x=>p(134)(48),y=>p(135)(48),Cin=>p(136)(48),clock=>clock,reset=>reset,s=>p(218)(48),cout=>p(219)(49));
FA_ff_5678:FAff port map(x=>p(134)(49),y=>p(135)(49),Cin=>p(136)(49),clock=>clock,reset=>reset,s=>p(218)(49),cout=>p(219)(50));
FA_ff_5679:FAff port map(x=>p(134)(50),y=>p(135)(50),Cin=>p(136)(50),clock=>clock,reset=>reset,s=>p(218)(50),cout=>p(219)(51));
FA_ff_5680:FAff port map(x=>p(134)(51),y=>p(135)(51),Cin=>p(136)(51),clock=>clock,reset=>reset,s=>p(218)(51),cout=>p(219)(52));
FA_ff_5681:FAff port map(x=>p(134)(52),y=>p(135)(52),Cin=>p(136)(52),clock=>clock,reset=>reset,s=>p(218)(52),cout=>p(219)(53));
FA_ff_5682:FAff port map(x=>p(134)(53),y=>p(135)(53),Cin=>p(136)(53),clock=>clock,reset=>reset,s=>p(218)(53),cout=>p(219)(54));
FA_ff_5683:FAff port map(x=>p(134)(54),y=>p(135)(54),Cin=>p(136)(54),clock=>clock,reset=>reset,s=>p(218)(54),cout=>p(219)(55));
FA_ff_5684:FAff port map(x=>p(134)(55),y=>p(135)(55),Cin=>p(136)(55),clock=>clock,reset=>reset,s=>p(218)(55),cout=>p(219)(56));
FA_ff_5685:FAff port map(x=>p(134)(56),y=>p(135)(56),Cin=>p(136)(56),clock=>clock,reset=>reset,s=>p(218)(56),cout=>p(219)(57));
FA_ff_5686:FAff port map(x=>p(134)(57),y=>p(135)(57),Cin=>p(136)(57),clock=>clock,reset=>reset,s=>p(218)(57),cout=>p(219)(58));
FA_ff_5687:FAff port map(x=>p(134)(58),y=>p(135)(58),Cin=>p(136)(58),clock=>clock,reset=>reset,s=>p(218)(58),cout=>p(219)(59));
FA_ff_5688:FAff port map(x=>p(134)(59),y=>p(135)(59),Cin=>p(136)(59),clock=>clock,reset=>reset,s=>p(218)(59),cout=>p(219)(60));
FA_ff_5689:FAff port map(x=>p(134)(60),y=>p(135)(60),Cin=>p(136)(60),clock=>clock,reset=>reset,s=>p(218)(60),cout=>p(219)(61));
FA_ff_5690:FAff port map(x=>p(134)(61),y=>p(135)(61),Cin=>p(136)(61),clock=>clock,reset=>reset,s=>p(218)(61),cout=>p(219)(62));
FA_ff_5691:FAff port map(x=>p(134)(62),y=>p(135)(62),Cin=>p(136)(62),clock=>clock,reset=>reset,s=>p(218)(62),cout=>p(219)(63));
FA_ff_5692:FAff port map(x=>p(134)(63),y=>p(135)(63),Cin=>p(136)(63),clock=>clock,reset=>reset,s=>p(218)(63),cout=>p(219)(64));
FA_ff_5693:FAff port map(x=>p(134)(64),y=>p(135)(64),Cin=>p(136)(64),clock=>clock,reset=>reset,s=>p(218)(64),cout=>p(219)(65));
FA_ff_5694:FAff port map(x=>p(134)(65),y=>p(135)(65),Cin=>p(136)(65),clock=>clock,reset=>reset,s=>p(218)(65),cout=>p(219)(66));
FA_ff_5695:FAff port map(x=>p(134)(66),y=>p(135)(66),Cin=>p(136)(66),clock=>clock,reset=>reset,s=>p(218)(66),cout=>p(219)(67));
FA_ff_5696:FAff port map(x=>p(134)(67),y=>p(135)(67),Cin=>p(136)(67),clock=>clock,reset=>reset,s=>p(218)(67),cout=>p(219)(68));
FA_ff_5697:FAff port map(x=>p(134)(68),y=>p(135)(68),Cin=>p(136)(68),clock=>clock,reset=>reset,s=>p(218)(68),cout=>p(219)(69));
FA_ff_5698:FAff port map(x=>p(134)(69),y=>p(135)(69),Cin=>p(136)(69),clock=>clock,reset=>reset,s=>p(218)(69),cout=>p(219)(70));
FA_ff_5699:FAff port map(x=>p(134)(70),y=>p(135)(70),Cin=>p(136)(70),clock=>clock,reset=>reset,s=>p(218)(70),cout=>p(219)(71));
FA_ff_5700:FAff port map(x=>p(134)(71),y=>p(135)(71),Cin=>p(136)(71),clock=>clock,reset=>reset,s=>p(218)(71),cout=>p(219)(72));
FA_ff_5701:FAff port map(x=>p(134)(72),y=>p(135)(72),Cin=>p(136)(72),clock=>clock,reset=>reset,s=>p(218)(72),cout=>p(219)(73));
FA_ff_5702:FAff port map(x=>p(134)(73),y=>p(135)(73),Cin=>p(136)(73),clock=>clock,reset=>reset,s=>p(218)(73),cout=>p(219)(74));
FA_ff_5703:FAff port map(x=>p(134)(74),y=>p(135)(74),Cin=>p(136)(74),clock=>clock,reset=>reset,s=>p(218)(74),cout=>p(219)(75));
FA_ff_5704:FAff port map(x=>p(134)(75),y=>p(135)(75),Cin=>p(136)(75),clock=>clock,reset=>reset,s=>p(218)(75),cout=>p(219)(76));
FA_ff_5705:FAff port map(x=>p(134)(76),y=>p(135)(76),Cin=>p(136)(76),clock=>clock,reset=>reset,s=>p(218)(76),cout=>p(219)(77));
FA_ff_5706:FAff port map(x=>p(134)(77),y=>p(135)(77),Cin=>p(136)(77),clock=>clock,reset=>reset,s=>p(218)(77),cout=>p(219)(78));
FA_ff_5707:FAff port map(x=>p(134)(78),y=>p(135)(78),Cin=>p(136)(78),clock=>clock,reset=>reset,s=>p(218)(78),cout=>p(219)(79));
FA_ff_5708:FAff port map(x=>p(134)(79),y=>p(135)(79),Cin=>p(136)(79),clock=>clock,reset=>reset,s=>p(218)(79),cout=>p(219)(80));
FA_ff_5709:FAff port map(x=>p(134)(80),y=>p(135)(80),Cin=>p(136)(80),clock=>clock,reset=>reset,s=>p(218)(80),cout=>p(219)(81));
FA_ff_5710:FAff port map(x=>p(134)(81),y=>p(135)(81),Cin=>p(136)(81),clock=>clock,reset=>reset,s=>p(218)(81),cout=>p(219)(82));
FA_ff_5711:FAff port map(x=>p(134)(82),y=>p(135)(82),Cin=>p(136)(82),clock=>clock,reset=>reset,s=>p(218)(82),cout=>p(219)(83));
FA_ff_5712:FAff port map(x=>p(134)(83),y=>p(135)(83),Cin=>p(136)(83),clock=>clock,reset=>reset,s=>p(218)(83),cout=>p(219)(84));
FA_ff_5713:FAff port map(x=>p(134)(84),y=>p(135)(84),Cin=>p(136)(84),clock=>clock,reset=>reset,s=>p(218)(84),cout=>p(219)(85));
FA_ff_5714:FAff port map(x=>p(134)(85),y=>p(135)(85),Cin=>p(136)(85),clock=>clock,reset=>reset,s=>p(218)(85),cout=>p(219)(86));
FA_ff_5715:FAff port map(x=>p(134)(86),y=>p(135)(86),Cin=>p(136)(86),clock=>clock,reset=>reset,s=>p(218)(86),cout=>p(219)(87));
FA_ff_5716:FAff port map(x=>p(134)(87),y=>p(135)(87),Cin=>p(136)(87),clock=>clock,reset=>reset,s=>p(218)(87),cout=>p(219)(88));
FA_ff_5717:FAff port map(x=>p(134)(88),y=>p(135)(88),Cin=>p(136)(88),clock=>clock,reset=>reset,s=>p(218)(88),cout=>p(219)(89));
FA_ff_5718:FAff port map(x=>p(134)(89),y=>p(135)(89),Cin=>p(136)(89),clock=>clock,reset=>reset,s=>p(218)(89),cout=>p(219)(90));
FA_ff_5719:FAff port map(x=>p(134)(90),y=>p(135)(90),Cin=>p(136)(90),clock=>clock,reset=>reset,s=>p(218)(90),cout=>p(219)(91));
FA_ff_5720:FAff port map(x=>p(134)(91),y=>p(135)(91),Cin=>p(136)(91),clock=>clock,reset=>reset,s=>p(218)(91),cout=>p(219)(92));
FA_ff_5721:FAff port map(x=>p(134)(92),y=>p(135)(92),Cin=>p(136)(92),clock=>clock,reset=>reset,s=>p(218)(92),cout=>p(219)(93));
FA_ff_5722:FAff port map(x=>p(134)(93),y=>p(135)(93),Cin=>p(136)(93),clock=>clock,reset=>reset,s=>p(218)(93),cout=>p(219)(94));
FA_ff_5723:FAff port map(x=>p(134)(94),y=>p(135)(94),Cin=>p(136)(94),clock=>clock,reset=>reset,s=>p(218)(94),cout=>p(219)(95));
FA_ff_5724:FAff port map(x=>p(134)(95),y=>p(135)(95),Cin=>p(136)(95),clock=>clock,reset=>reset,s=>p(218)(95),cout=>p(219)(96));
FA_ff_5725:FAff port map(x=>p(134)(96),y=>p(135)(96),Cin=>p(136)(96),clock=>clock,reset=>reset,s=>p(218)(96),cout=>p(219)(97));
FA_ff_5726:FAff port map(x=>p(134)(97),y=>p(135)(97),Cin=>p(136)(97),clock=>clock,reset=>reset,s=>p(218)(97),cout=>p(219)(98));
FA_ff_5727:FAff port map(x=>p(134)(98),y=>p(135)(98),Cin=>p(136)(98),clock=>clock,reset=>reset,s=>p(218)(98),cout=>p(219)(99));
FA_ff_5728:FAff port map(x=>p(134)(99),y=>p(135)(99),Cin=>p(136)(99),clock=>clock,reset=>reset,s=>p(218)(99),cout=>p(219)(100));
FA_ff_5729:FAff port map(x=>p(134)(100),y=>p(135)(100),Cin=>p(136)(100),clock=>clock,reset=>reset,s=>p(218)(100),cout=>p(219)(101));
FA_ff_5730:FAff port map(x=>p(134)(101),y=>p(135)(101),Cin=>p(136)(101),clock=>clock,reset=>reset,s=>p(218)(101),cout=>p(219)(102));
FA_ff_5731:FAff port map(x=>p(134)(102),y=>p(135)(102),Cin=>p(136)(102),clock=>clock,reset=>reset,s=>p(218)(102),cout=>p(219)(103));
FA_ff_5732:FAff port map(x=>p(134)(103),y=>p(135)(103),Cin=>p(136)(103),clock=>clock,reset=>reset,s=>p(218)(103),cout=>p(219)(104));
FA_ff_5733:FAff port map(x=>p(134)(104),y=>p(135)(104),Cin=>p(136)(104),clock=>clock,reset=>reset,s=>p(218)(104),cout=>p(219)(105));
FA_ff_5734:FAff port map(x=>p(134)(105),y=>p(135)(105),Cin=>p(136)(105),clock=>clock,reset=>reset,s=>p(218)(105),cout=>p(219)(106));
FA_ff_5735:FAff port map(x=>p(134)(106),y=>p(135)(106),Cin=>p(136)(106),clock=>clock,reset=>reset,s=>p(218)(106),cout=>p(219)(107));
FA_ff_5736:FAff port map(x=>p(134)(107),y=>p(135)(107),Cin=>p(136)(107),clock=>clock,reset=>reset,s=>p(218)(107),cout=>p(219)(108));
FA_ff_5737:FAff port map(x=>p(134)(108),y=>p(135)(108),Cin=>p(136)(108),clock=>clock,reset=>reset,s=>p(218)(108),cout=>p(219)(109));
FA_ff_5738:FAff port map(x=>p(134)(109),y=>p(135)(109),Cin=>p(136)(109),clock=>clock,reset=>reset,s=>p(218)(109),cout=>p(219)(110));
FA_ff_5739:FAff port map(x=>p(134)(110),y=>p(135)(110),Cin=>p(136)(110),clock=>clock,reset=>reset,s=>p(218)(110),cout=>p(219)(111));
FA_ff_5740:FAff port map(x=>p(134)(111),y=>p(135)(111),Cin=>p(136)(111),clock=>clock,reset=>reset,s=>p(218)(111),cout=>p(219)(112));
FA_ff_5741:FAff port map(x=>p(134)(112),y=>p(135)(112),Cin=>p(136)(112),clock=>clock,reset=>reset,s=>p(218)(112),cout=>p(219)(113));
FA_ff_5742:FAff port map(x=>p(134)(113),y=>p(135)(113),Cin=>p(136)(113),clock=>clock,reset=>reset,s=>p(218)(113),cout=>p(219)(114));
FA_ff_5743:FAff port map(x=>p(134)(114),y=>p(135)(114),Cin=>p(136)(114),clock=>clock,reset=>reset,s=>p(218)(114),cout=>p(219)(115));
FA_ff_5744:FAff port map(x=>p(134)(115),y=>p(135)(115),Cin=>p(136)(115),clock=>clock,reset=>reset,s=>p(218)(115),cout=>p(219)(116));
FA_ff_5745:FAff port map(x=>p(134)(116),y=>p(135)(116),Cin=>p(136)(116),clock=>clock,reset=>reset,s=>p(218)(116),cout=>p(219)(117));
FA_ff_5746:FAff port map(x=>p(134)(117),y=>p(135)(117),Cin=>p(136)(117),clock=>clock,reset=>reset,s=>p(218)(117),cout=>p(219)(118));
FA_ff_5747:FAff port map(x=>p(134)(118),y=>p(135)(118),Cin=>p(136)(118),clock=>clock,reset=>reset,s=>p(218)(118),cout=>p(219)(119));
FA_ff_5748:FAff port map(x=>p(134)(119),y=>p(135)(119),Cin=>p(136)(119),clock=>clock,reset=>reset,s=>p(218)(119),cout=>p(219)(120));
FA_ff_5749:FAff port map(x=>p(134)(120),y=>p(135)(120),Cin=>p(136)(120),clock=>clock,reset=>reset,s=>p(218)(120),cout=>p(219)(121));
FA_ff_5750:FAff port map(x=>p(134)(121),y=>p(135)(121),Cin=>p(136)(121),clock=>clock,reset=>reset,s=>p(218)(121),cout=>p(219)(122));
FA_ff_5751:FAff port map(x=>p(134)(122),y=>p(135)(122),Cin=>p(136)(122),clock=>clock,reset=>reset,s=>p(218)(122),cout=>p(219)(123));
FA_ff_5752:FAff port map(x=>p(134)(123),y=>p(135)(123),Cin=>p(136)(123),clock=>clock,reset=>reset,s=>p(218)(123),cout=>p(219)(124));
FA_ff_5753:FAff port map(x=>p(134)(124),y=>p(135)(124),Cin=>p(136)(124),clock=>clock,reset=>reset,s=>p(218)(124),cout=>p(219)(125));
FA_ff_5754:FAff port map(x=>p(134)(125),y=>p(135)(125),Cin=>p(136)(125),clock=>clock,reset=>reset,s=>p(218)(125),cout=>p(219)(126));
FA_ff_5755:FAff port map(x=>p(134)(126),y=>p(135)(126),Cin=>p(136)(126),clock=>clock,reset=>reset,s=>p(218)(126),cout=>p(219)(127));
FA_ff_5756:FAff port map(x=>p(134)(127),y=>p(135)(127),Cin=>p(136)(127),clock=>clock,reset=>reset,s=>p(218)(127),cout=>p(219)(128));
p(218)(128)<=p(135)(128);
p(220)(0)<=p(138)(0);
FA_ff_5757:FAff port map(x=>p(137)(1),y=>p(138)(1),Cin=>p(139)(1),clock=>clock,reset=>reset,s=>p(220)(1),cout=>p(221)(2));
FA_ff_5758:FAff port map(x=>p(137)(2),y=>p(138)(2),Cin=>p(139)(2),clock=>clock,reset=>reset,s=>p(220)(2),cout=>p(221)(3));
FA_ff_5759:FAff port map(x=>p(137)(3),y=>p(138)(3),Cin=>p(139)(3),clock=>clock,reset=>reset,s=>p(220)(3),cout=>p(221)(4));
FA_ff_5760:FAff port map(x=>p(137)(4),y=>p(138)(4),Cin=>p(139)(4),clock=>clock,reset=>reset,s=>p(220)(4),cout=>p(221)(5));
FA_ff_5761:FAff port map(x=>p(137)(5),y=>p(138)(5),Cin=>p(139)(5),clock=>clock,reset=>reset,s=>p(220)(5),cout=>p(221)(6));
FA_ff_5762:FAff port map(x=>p(137)(6),y=>p(138)(6),Cin=>p(139)(6),clock=>clock,reset=>reset,s=>p(220)(6),cout=>p(221)(7));
FA_ff_5763:FAff port map(x=>p(137)(7),y=>p(138)(7),Cin=>p(139)(7),clock=>clock,reset=>reset,s=>p(220)(7),cout=>p(221)(8));
FA_ff_5764:FAff port map(x=>p(137)(8),y=>p(138)(8),Cin=>p(139)(8),clock=>clock,reset=>reset,s=>p(220)(8),cout=>p(221)(9));
FA_ff_5765:FAff port map(x=>p(137)(9),y=>p(138)(9),Cin=>p(139)(9),clock=>clock,reset=>reset,s=>p(220)(9),cout=>p(221)(10));
FA_ff_5766:FAff port map(x=>p(137)(10),y=>p(138)(10),Cin=>p(139)(10),clock=>clock,reset=>reset,s=>p(220)(10),cout=>p(221)(11));
FA_ff_5767:FAff port map(x=>p(137)(11),y=>p(138)(11),Cin=>p(139)(11),clock=>clock,reset=>reset,s=>p(220)(11),cout=>p(221)(12));
FA_ff_5768:FAff port map(x=>p(137)(12),y=>p(138)(12),Cin=>p(139)(12),clock=>clock,reset=>reset,s=>p(220)(12),cout=>p(221)(13));
FA_ff_5769:FAff port map(x=>p(137)(13),y=>p(138)(13),Cin=>p(139)(13),clock=>clock,reset=>reset,s=>p(220)(13),cout=>p(221)(14));
FA_ff_5770:FAff port map(x=>p(137)(14),y=>p(138)(14),Cin=>p(139)(14),clock=>clock,reset=>reset,s=>p(220)(14),cout=>p(221)(15));
FA_ff_5771:FAff port map(x=>p(137)(15),y=>p(138)(15),Cin=>p(139)(15),clock=>clock,reset=>reset,s=>p(220)(15),cout=>p(221)(16));
FA_ff_5772:FAff port map(x=>p(137)(16),y=>p(138)(16),Cin=>p(139)(16),clock=>clock,reset=>reset,s=>p(220)(16),cout=>p(221)(17));
FA_ff_5773:FAff port map(x=>p(137)(17),y=>p(138)(17),Cin=>p(139)(17),clock=>clock,reset=>reset,s=>p(220)(17),cout=>p(221)(18));
FA_ff_5774:FAff port map(x=>p(137)(18),y=>p(138)(18),Cin=>p(139)(18),clock=>clock,reset=>reset,s=>p(220)(18),cout=>p(221)(19));
FA_ff_5775:FAff port map(x=>p(137)(19),y=>p(138)(19),Cin=>p(139)(19),clock=>clock,reset=>reset,s=>p(220)(19),cout=>p(221)(20));
FA_ff_5776:FAff port map(x=>p(137)(20),y=>p(138)(20),Cin=>p(139)(20),clock=>clock,reset=>reset,s=>p(220)(20),cout=>p(221)(21));
FA_ff_5777:FAff port map(x=>p(137)(21),y=>p(138)(21),Cin=>p(139)(21),clock=>clock,reset=>reset,s=>p(220)(21),cout=>p(221)(22));
FA_ff_5778:FAff port map(x=>p(137)(22),y=>p(138)(22),Cin=>p(139)(22),clock=>clock,reset=>reset,s=>p(220)(22),cout=>p(221)(23));
FA_ff_5779:FAff port map(x=>p(137)(23),y=>p(138)(23),Cin=>p(139)(23),clock=>clock,reset=>reset,s=>p(220)(23),cout=>p(221)(24));
FA_ff_5780:FAff port map(x=>p(137)(24),y=>p(138)(24),Cin=>p(139)(24),clock=>clock,reset=>reset,s=>p(220)(24),cout=>p(221)(25));
FA_ff_5781:FAff port map(x=>p(137)(25),y=>p(138)(25),Cin=>p(139)(25),clock=>clock,reset=>reset,s=>p(220)(25),cout=>p(221)(26));
FA_ff_5782:FAff port map(x=>p(137)(26),y=>p(138)(26),Cin=>p(139)(26),clock=>clock,reset=>reset,s=>p(220)(26),cout=>p(221)(27));
FA_ff_5783:FAff port map(x=>p(137)(27),y=>p(138)(27),Cin=>p(139)(27),clock=>clock,reset=>reset,s=>p(220)(27),cout=>p(221)(28));
FA_ff_5784:FAff port map(x=>p(137)(28),y=>p(138)(28),Cin=>p(139)(28),clock=>clock,reset=>reset,s=>p(220)(28),cout=>p(221)(29));
FA_ff_5785:FAff port map(x=>p(137)(29),y=>p(138)(29),Cin=>p(139)(29),clock=>clock,reset=>reset,s=>p(220)(29),cout=>p(221)(30));
FA_ff_5786:FAff port map(x=>p(137)(30),y=>p(138)(30),Cin=>p(139)(30),clock=>clock,reset=>reset,s=>p(220)(30),cout=>p(221)(31));
FA_ff_5787:FAff port map(x=>p(137)(31),y=>p(138)(31),Cin=>p(139)(31),clock=>clock,reset=>reset,s=>p(220)(31),cout=>p(221)(32));
FA_ff_5788:FAff port map(x=>p(137)(32),y=>p(138)(32),Cin=>p(139)(32),clock=>clock,reset=>reset,s=>p(220)(32),cout=>p(221)(33));
FA_ff_5789:FAff port map(x=>p(137)(33),y=>p(138)(33),Cin=>p(139)(33),clock=>clock,reset=>reset,s=>p(220)(33),cout=>p(221)(34));
FA_ff_5790:FAff port map(x=>p(137)(34),y=>p(138)(34),Cin=>p(139)(34),clock=>clock,reset=>reset,s=>p(220)(34),cout=>p(221)(35));
FA_ff_5791:FAff port map(x=>p(137)(35),y=>p(138)(35),Cin=>p(139)(35),clock=>clock,reset=>reset,s=>p(220)(35),cout=>p(221)(36));
FA_ff_5792:FAff port map(x=>p(137)(36),y=>p(138)(36),Cin=>p(139)(36),clock=>clock,reset=>reset,s=>p(220)(36),cout=>p(221)(37));
FA_ff_5793:FAff port map(x=>p(137)(37),y=>p(138)(37),Cin=>p(139)(37),clock=>clock,reset=>reset,s=>p(220)(37),cout=>p(221)(38));
FA_ff_5794:FAff port map(x=>p(137)(38),y=>p(138)(38),Cin=>p(139)(38),clock=>clock,reset=>reset,s=>p(220)(38),cout=>p(221)(39));
FA_ff_5795:FAff port map(x=>p(137)(39),y=>p(138)(39),Cin=>p(139)(39),clock=>clock,reset=>reset,s=>p(220)(39),cout=>p(221)(40));
FA_ff_5796:FAff port map(x=>p(137)(40),y=>p(138)(40),Cin=>p(139)(40),clock=>clock,reset=>reset,s=>p(220)(40),cout=>p(221)(41));
FA_ff_5797:FAff port map(x=>p(137)(41),y=>p(138)(41),Cin=>p(139)(41),clock=>clock,reset=>reset,s=>p(220)(41),cout=>p(221)(42));
FA_ff_5798:FAff port map(x=>p(137)(42),y=>p(138)(42),Cin=>p(139)(42),clock=>clock,reset=>reset,s=>p(220)(42),cout=>p(221)(43));
FA_ff_5799:FAff port map(x=>p(137)(43),y=>p(138)(43),Cin=>p(139)(43),clock=>clock,reset=>reset,s=>p(220)(43),cout=>p(221)(44));
FA_ff_5800:FAff port map(x=>p(137)(44),y=>p(138)(44),Cin=>p(139)(44),clock=>clock,reset=>reset,s=>p(220)(44),cout=>p(221)(45));
FA_ff_5801:FAff port map(x=>p(137)(45),y=>p(138)(45),Cin=>p(139)(45),clock=>clock,reset=>reset,s=>p(220)(45),cout=>p(221)(46));
FA_ff_5802:FAff port map(x=>p(137)(46),y=>p(138)(46),Cin=>p(139)(46),clock=>clock,reset=>reset,s=>p(220)(46),cout=>p(221)(47));
FA_ff_5803:FAff port map(x=>p(137)(47),y=>p(138)(47),Cin=>p(139)(47),clock=>clock,reset=>reset,s=>p(220)(47),cout=>p(221)(48));
FA_ff_5804:FAff port map(x=>p(137)(48),y=>p(138)(48),Cin=>p(139)(48),clock=>clock,reset=>reset,s=>p(220)(48),cout=>p(221)(49));
FA_ff_5805:FAff port map(x=>p(137)(49),y=>p(138)(49),Cin=>p(139)(49),clock=>clock,reset=>reset,s=>p(220)(49),cout=>p(221)(50));
FA_ff_5806:FAff port map(x=>p(137)(50),y=>p(138)(50),Cin=>p(139)(50),clock=>clock,reset=>reset,s=>p(220)(50),cout=>p(221)(51));
FA_ff_5807:FAff port map(x=>p(137)(51),y=>p(138)(51),Cin=>p(139)(51),clock=>clock,reset=>reset,s=>p(220)(51),cout=>p(221)(52));
FA_ff_5808:FAff port map(x=>p(137)(52),y=>p(138)(52),Cin=>p(139)(52),clock=>clock,reset=>reset,s=>p(220)(52),cout=>p(221)(53));
FA_ff_5809:FAff port map(x=>p(137)(53),y=>p(138)(53),Cin=>p(139)(53),clock=>clock,reset=>reset,s=>p(220)(53),cout=>p(221)(54));
FA_ff_5810:FAff port map(x=>p(137)(54),y=>p(138)(54),Cin=>p(139)(54),clock=>clock,reset=>reset,s=>p(220)(54),cout=>p(221)(55));
FA_ff_5811:FAff port map(x=>p(137)(55),y=>p(138)(55),Cin=>p(139)(55),clock=>clock,reset=>reset,s=>p(220)(55),cout=>p(221)(56));
FA_ff_5812:FAff port map(x=>p(137)(56),y=>p(138)(56),Cin=>p(139)(56),clock=>clock,reset=>reset,s=>p(220)(56),cout=>p(221)(57));
FA_ff_5813:FAff port map(x=>p(137)(57),y=>p(138)(57),Cin=>p(139)(57),clock=>clock,reset=>reset,s=>p(220)(57),cout=>p(221)(58));
FA_ff_5814:FAff port map(x=>p(137)(58),y=>p(138)(58),Cin=>p(139)(58),clock=>clock,reset=>reset,s=>p(220)(58),cout=>p(221)(59));
FA_ff_5815:FAff port map(x=>p(137)(59),y=>p(138)(59),Cin=>p(139)(59),clock=>clock,reset=>reset,s=>p(220)(59),cout=>p(221)(60));
FA_ff_5816:FAff port map(x=>p(137)(60),y=>p(138)(60),Cin=>p(139)(60),clock=>clock,reset=>reset,s=>p(220)(60),cout=>p(221)(61));
FA_ff_5817:FAff port map(x=>p(137)(61),y=>p(138)(61),Cin=>p(139)(61),clock=>clock,reset=>reset,s=>p(220)(61),cout=>p(221)(62));
FA_ff_5818:FAff port map(x=>p(137)(62),y=>p(138)(62),Cin=>p(139)(62),clock=>clock,reset=>reset,s=>p(220)(62),cout=>p(221)(63));
FA_ff_5819:FAff port map(x=>p(137)(63),y=>p(138)(63),Cin=>p(139)(63),clock=>clock,reset=>reset,s=>p(220)(63),cout=>p(221)(64));
FA_ff_5820:FAff port map(x=>p(137)(64),y=>p(138)(64),Cin=>p(139)(64),clock=>clock,reset=>reset,s=>p(220)(64),cout=>p(221)(65));
FA_ff_5821:FAff port map(x=>p(137)(65),y=>p(138)(65),Cin=>p(139)(65),clock=>clock,reset=>reset,s=>p(220)(65),cout=>p(221)(66));
FA_ff_5822:FAff port map(x=>p(137)(66),y=>p(138)(66),Cin=>p(139)(66),clock=>clock,reset=>reset,s=>p(220)(66),cout=>p(221)(67));
FA_ff_5823:FAff port map(x=>p(137)(67),y=>p(138)(67),Cin=>p(139)(67),clock=>clock,reset=>reset,s=>p(220)(67),cout=>p(221)(68));
FA_ff_5824:FAff port map(x=>p(137)(68),y=>p(138)(68),Cin=>p(139)(68),clock=>clock,reset=>reset,s=>p(220)(68),cout=>p(221)(69));
FA_ff_5825:FAff port map(x=>p(137)(69),y=>p(138)(69),Cin=>p(139)(69),clock=>clock,reset=>reset,s=>p(220)(69),cout=>p(221)(70));
FA_ff_5826:FAff port map(x=>p(137)(70),y=>p(138)(70),Cin=>p(139)(70),clock=>clock,reset=>reset,s=>p(220)(70),cout=>p(221)(71));
FA_ff_5827:FAff port map(x=>p(137)(71),y=>p(138)(71),Cin=>p(139)(71),clock=>clock,reset=>reset,s=>p(220)(71),cout=>p(221)(72));
FA_ff_5828:FAff port map(x=>p(137)(72),y=>p(138)(72),Cin=>p(139)(72),clock=>clock,reset=>reset,s=>p(220)(72),cout=>p(221)(73));
FA_ff_5829:FAff port map(x=>p(137)(73),y=>p(138)(73),Cin=>p(139)(73),clock=>clock,reset=>reset,s=>p(220)(73),cout=>p(221)(74));
FA_ff_5830:FAff port map(x=>p(137)(74),y=>p(138)(74),Cin=>p(139)(74),clock=>clock,reset=>reset,s=>p(220)(74),cout=>p(221)(75));
FA_ff_5831:FAff port map(x=>p(137)(75),y=>p(138)(75),Cin=>p(139)(75),clock=>clock,reset=>reset,s=>p(220)(75),cout=>p(221)(76));
FA_ff_5832:FAff port map(x=>p(137)(76),y=>p(138)(76),Cin=>p(139)(76),clock=>clock,reset=>reset,s=>p(220)(76),cout=>p(221)(77));
FA_ff_5833:FAff port map(x=>p(137)(77),y=>p(138)(77),Cin=>p(139)(77),clock=>clock,reset=>reset,s=>p(220)(77),cout=>p(221)(78));
FA_ff_5834:FAff port map(x=>p(137)(78),y=>p(138)(78),Cin=>p(139)(78),clock=>clock,reset=>reset,s=>p(220)(78),cout=>p(221)(79));
FA_ff_5835:FAff port map(x=>p(137)(79),y=>p(138)(79),Cin=>p(139)(79),clock=>clock,reset=>reset,s=>p(220)(79),cout=>p(221)(80));
FA_ff_5836:FAff port map(x=>p(137)(80),y=>p(138)(80),Cin=>p(139)(80),clock=>clock,reset=>reset,s=>p(220)(80),cout=>p(221)(81));
FA_ff_5837:FAff port map(x=>p(137)(81),y=>p(138)(81),Cin=>p(139)(81),clock=>clock,reset=>reset,s=>p(220)(81),cout=>p(221)(82));
FA_ff_5838:FAff port map(x=>p(137)(82),y=>p(138)(82),Cin=>p(139)(82),clock=>clock,reset=>reset,s=>p(220)(82),cout=>p(221)(83));
FA_ff_5839:FAff port map(x=>p(137)(83),y=>p(138)(83),Cin=>p(139)(83),clock=>clock,reset=>reset,s=>p(220)(83),cout=>p(221)(84));
FA_ff_5840:FAff port map(x=>p(137)(84),y=>p(138)(84),Cin=>p(139)(84),clock=>clock,reset=>reset,s=>p(220)(84),cout=>p(221)(85));
FA_ff_5841:FAff port map(x=>p(137)(85),y=>p(138)(85),Cin=>p(139)(85),clock=>clock,reset=>reset,s=>p(220)(85),cout=>p(221)(86));
FA_ff_5842:FAff port map(x=>p(137)(86),y=>p(138)(86),Cin=>p(139)(86),clock=>clock,reset=>reset,s=>p(220)(86),cout=>p(221)(87));
FA_ff_5843:FAff port map(x=>p(137)(87),y=>p(138)(87),Cin=>p(139)(87),clock=>clock,reset=>reset,s=>p(220)(87),cout=>p(221)(88));
FA_ff_5844:FAff port map(x=>p(137)(88),y=>p(138)(88),Cin=>p(139)(88),clock=>clock,reset=>reset,s=>p(220)(88),cout=>p(221)(89));
FA_ff_5845:FAff port map(x=>p(137)(89),y=>p(138)(89),Cin=>p(139)(89),clock=>clock,reset=>reset,s=>p(220)(89),cout=>p(221)(90));
FA_ff_5846:FAff port map(x=>p(137)(90),y=>p(138)(90),Cin=>p(139)(90),clock=>clock,reset=>reset,s=>p(220)(90),cout=>p(221)(91));
FA_ff_5847:FAff port map(x=>p(137)(91),y=>p(138)(91),Cin=>p(139)(91),clock=>clock,reset=>reset,s=>p(220)(91),cout=>p(221)(92));
FA_ff_5848:FAff port map(x=>p(137)(92),y=>p(138)(92),Cin=>p(139)(92),clock=>clock,reset=>reset,s=>p(220)(92),cout=>p(221)(93));
FA_ff_5849:FAff port map(x=>p(137)(93),y=>p(138)(93),Cin=>p(139)(93),clock=>clock,reset=>reset,s=>p(220)(93),cout=>p(221)(94));
FA_ff_5850:FAff port map(x=>p(137)(94),y=>p(138)(94),Cin=>p(139)(94),clock=>clock,reset=>reset,s=>p(220)(94),cout=>p(221)(95));
FA_ff_5851:FAff port map(x=>p(137)(95),y=>p(138)(95),Cin=>p(139)(95),clock=>clock,reset=>reset,s=>p(220)(95),cout=>p(221)(96));
FA_ff_5852:FAff port map(x=>p(137)(96),y=>p(138)(96),Cin=>p(139)(96),clock=>clock,reset=>reset,s=>p(220)(96),cout=>p(221)(97));
FA_ff_5853:FAff port map(x=>p(137)(97),y=>p(138)(97),Cin=>p(139)(97),clock=>clock,reset=>reset,s=>p(220)(97),cout=>p(221)(98));
FA_ff_5854:FAff port map(x=>p(137)(98),y=>p(138)(98),Cin=>p(139)(98),clock=>clock,reset=>reset,s=>p(220)(98),cout=>p(221)(99));
FA_ff_5855:FAff port map(x=>p(137)(99),y=>p(138)(99),Cin=>p(139)(99),clock=>clock,reset=>reset,s=>p(220)(99),cout=>p(221)(100));
FA_ff_5856:FAff port map(x=>p(137)(100),y=>p(138)(100),Cin=>p(139)(100),clock=>clock,reset=>reset,s=>p(220)(100),cout=>p(221)(101));
FA_ff_5857:FAff port map(x=>p(137)(101),y=>p(138)(101),Cin=>p(139)(101),clock=>clock,reset=>reset,s=>p(220)(101),cout=>p(221)(102));
FA_ff_5858:FAff port map(x=>p(137)(102),y=>p(138)(102),Cin=>p(139)(102),clock=>clock,reset=>reset,s=>p(220)(102),cout=>p(221)(103));
FA_ff_5859:FAff port map(x=>p(137)(103),y=>p(138)(103),Cin=>p(139)(103),clock=>clock,reset=>reset,s=>p(220)(103),cout=>p(221)(104));
FA_ff_5860:FAff port map(x=>p(137)(104),y=>p(138)(104),Cin=>p(139)(104),clock=>clock,reset=>reset,s=>p(220)(104),cout=>p(221)(105));
FA_ff_5861:FAff port map(x=>p(137)(105),y=>p(138)(105),Cin=>p(139)(105),clock=>clock,reset=>reset,s=>p(220)(105),cout=>p(221)(106));
FA_ff_5862:FAff port map(x=>p(137)(106),y=>p(138)(106),Cin=>p(139)(106),clock=>clock,reset=>reset,s=>p(220)(106),cout=>p(221)(107));
FA_ff_5863:FAff port map(x=>p(137)(107),y=>p(138)(107),Cin=>p(139)(107),clock=>clock,reset=>reset,s=>p(220)(107),cout=>p(221)(108));
FA_ff_5864:FAff port map(x=>p(137)(108),y=>p(138)(108),Cin=>p(139)(108),clock=>clock,reset=>reset,s=>p(220)(108),cout=>p(221)(109));
FA_ff_5865:FAff port map(x=>p(137)(109),y=>p(138)(109),Cin=>p(139)(109),clock=>clock,reset=>reset,s=>p(220)(109),cout=>p(221)(110));
FA_ff_5866:FAff port map(x=>p(137)(110),y=>p(138)(110),Cin=>p(139)(110),clock=>clock,reset=>reset,s=>p(220)(110),cout=>p(221)(111));
FA_ff_5867:FAff port map(x=>p(137)(111),y=>p(138)(111),Cin=>p(139)(111),clock=>clock,reset=>reset,s=>p(220)(111),cout=>p(221)(112));
FA_ff_5868:FAff port map(x=>p(137)(112),y=>p(138)(112),Cin=>p(139)(112),clock=>clock,reset=>reset,s=>p(220)(112),cout=>p(221)(113));
FA_ff_5869:FAff port map(x=>p(137)(113),y=>p(138)(113),Cin=>p(139)(113),clock=>clock,reset=>reset,s=>p(220)(113),cout=>p(221)(114));
FA_ff_5870:FAff port map(x=>p(137)(114),y=>p(138)(114),Cin=>p(139)(114),clock=>clock,reset=>reset,s=>p(220)(114),cout=>p(221)(115));
FA_ff_5871:FAff port map(x=>p(137)(115),y=>p(138)(115),Cin=>p(139)(115),clock=>clock,reset=>reset,s=>p(220)(115),cout=>p(221)(116));
FA_ff_5872:FAff port map(x=>p(137)(116),y=>p(138)(116),Cin=>p(139)(116),clock=>clock,reset=>reset,s=>p(220)(116),cout=>p(221)(117));
FA_ff_5873:FAff port map(x=>p(137)(117),y=>p(138)(117),Cin=>p(139)(117),clock=>clock,reset=>reset,s=>p(220)(117),cout=>p(221)(118));
FA_ff_5874:FAff port map(x=>p(137)(118),y=>p(138)(118),Cin=>p(139)(118),clock=>clock,reset=>reset,s=>p(220)(118),cout=>p(221)(119));
FA_ff_5875:FAff port map(x=>p(137)(119),y=>p(138)(119),Cin=>p(139)(119),clock=>clock,reset=>reset,s=>p(220)(119),cout=>p(221)(120));
FA_ff_5876:FAff port map(x=>p(137)(120),y=>p(138)(120),Cin=>p(139)(120),clock=>clock,reset=>reset,s=>p(220)(120),cout=>p(221)(121));
FA_ff_5877:FAff port map(x=>p(137)(121),y=>p(138)(121),Cin=>p(139)(121),clock=>clock,reset=>reset,s=>p(220)(121),cout=>p(221)(122));
FA_ff_5878:FAff port map(x=>p(137)(122),y=>p(138)(122),Cin=>p(139)(122),clock=>clock,reset=>reset,s=>p(220)(122),cout=>p(221)(123));
FA_ff_5879:FAff port map(x=>p(137)(123),y=>p(138)(123),Cin=>p(139)(123),clock=>clock,reset=>reset,s=>p(220)(123),cout=>p(221)(124));
FA_ff_5880:FAff port map(x=>p(137)(124),y=>p(138)(124),Cin=>p(139)(124),clock=>clock,reset=>reset,s=>p(220)(124),cout=>p(221)(125));
FA_ff_5881:FAff port map(x=>p(137)(125),y=>p(138)(125),Cin=>p(139)(125),clock=>clock,reset=>reset,s=>p(220)(125),cout=>p(221)(126));
FA_ff_5882:FAff port map(x=>p(137)(126),y=>p(138)(126),Cin=>p(139)(126),clock=>clock,reset=>reset,s=>p(220)(126),cout=>p(221)(127));
FA_ff_5883:FAff port map(x=>p(137)(127),y=>p(138)(127),Cin=>p(139)(127),clock=>clock,reset=>reset,s=>p(220)(127),cout=>p(221)(128));
HA_ff_3:HAff port map(x=>p(137)(128),y=>p(139)(128),clock=>clock,reset=>reset,s=>p(220)(128),c=>p(221)(129));
HA_ff_4:HAff port map(x=>p(140)(0),y=>p(142)(0),clock=>clock,reset=>reset,s=>p(222)(0),c=>p(223)(1));
FA_ff_5884:FAff port map(x=>p(140)(1),y=>p(141)(1),Cin=>p(142)(1),clock=>clock,reset=>reset,s=>p(222)(1),cout=>p(223)(2));
FA_ff_5885:FAff port map(x=>p(140)(2),y=>p(141)(2),Cin=>p(142)(2),clock=>clock,reset=>reset,s=>p(222)(2),cout=>p(223)(3));
FA_ff_5886:FAff port map(x=>p(140)(3),y=>p(141)(3),Cin=>p(142)(3),clock=>clock,reset=>reset,s=>p(222)(3),cout=>p(223)(4));
FA_ff_5887:FAff port map(x=>p(140)(4),y=>p(141)(4),Cin=>p(142)(4),clock=>clock,reset=>reset,s=>p(222)(4),cout=>p(223)(5));
FA_ff_5888:FAff port map(x=>p(140)(5),y=>p(141)(5),Cin=>p(142)(5),clock=>clock,reset=>reset,s=>p(222)(5),cout=>p(223)(6));
FA_ff_5889:FAff port map(x=>p(140)(6),y=>p(141)(6),Cin=>p(142)(6),clock=>clock,reset=>reset,s=>p(222)(6),cout=>p(223)(7));
FA_ff_5890:FAff port map(x=>p(140)(7),y=>p(141)(7),Cin=>p(142)(7),clock=>clock,reset=>reset,s=>p(222)(7),cout=>p(223)(8));
FA_ff_5891:FAff port map(x=>p(140)(8),y=>p(141)(8),Cin=>p(142)(8),clock=>clock,reset=>reset,s=>p(222)(8),cout=>p(223)(9));
FA_ff_5892:FAff port map(x=>p(140)(9),y=>p(141)(9),Cin=>p(142)(9),clock=>clock,reset=>reset,s=>p(222)(9),cout=>p(223)(10));
FA_ff_5893:FAff port map(x=>p(140)(10),y=>p(141)(10),Cin=>p(142)(10),clock=>clock,reset=>reset,s=>p(222)(10),cout=>p(223)(11));
FA_ff_5894:FAff port map(x=>p(140)(11),y=>p(141)(11),Cin=>p(142)(11),clock=>clock,reset=>reset,s=>p(222)(11),cout=>p(223)(12));
FA_ff_5895:FAff port map(x=>p(140)(12),y=>p(141)(12),Cin=>p(142)(12),clock=>clock,reset=>reset,s=>p(222)(12),cout=>p(223)(13));
FA_ff_5896:FAff port map(x=>p(140)(13),y=>p(141)(13),Cin=>p(142)(13),clock=>clock,reset=>reset,s=>p(222)(13),cout=>p(223)(14));
FA_ff_5897:FAff port map(x=>p(140)(14),y=>p(141)(14),Cin=>p(142)(14),clock=>clock,reset=>reset,s=>p(222)(14),cout=>p(223)(15));
FA_ff_5898:FAff port map(x=>p(140)(15),y=>p(141)(15),Cin=>p(142)(15),clock=>clock,reset=>reset,s=>p(222)(15),cout=>p(223)(16));
FA_ff_5899:FAff port map(x=>p(140)(16),y=>p(141)(16),Cin=>p(142)(16),clock=>clock,reset=>reset,s=>p(222)(16),cout=>p(223)(17));
FA_ff_5900:FAff port map(x=>p(140)(17),y=>p(141)(17),Cin=>p(142)(17),clock=>clock,reset=>reset,s=>p(222)(17),cout=>p(223)(18));
FA_ff_5901:FAff port map(x=>p(140)(18),y=>p(141)(18),Cin=>p(142)(18),clock=>clock,reset=>reset,s=>p(222)(18),cout=>p(223)(19));
FA_ff_5902:FAff port map(x=>p(140)(19),y=>p(141)(19),Cin=>p(142)(19),clock=>clock,reset=>reset,s=>p(222)(19),cout=>p(223)(20));
FA_ff_5903:FAff port map(x=>p(140)(20),y=>p(141)(20),Cin=>p(142)(20),clock=>clock,reset=>reset,s=>p(222)(20),cout=>p(223)(21));
FA_ff_5904:FAff port map(x=>p(140)(21),y=>p(141)(21),Cin=>p(142)(21),clock=>clock,reset=>reset,s=>p(222)(21),cout=>p(223)(22));
FA_ff_5905:FAff port map(x=>p(140)(22),y=>p(141)(22),Cin=>p(142)(22),clock=>clock,reset=>reset,s=>p(222)(22),cout=>p(223)(23));
FA_ff_5906:FAff port map(x=>p(140)(23),y=>p(141)(23),Cin=>p(142)(23),clock=>clock,reset=>reset,s=>p(222)(23),cout=>p(223)(24));
FA_ff_5907:FAff port map(x=>p(140)(24),y=>p(141)(24),Cin=>p(142)(24),clock=>clock,reset=>reset,s=>p(222)(24),cout=>p(223)(25));
FA_ff_5908:FAff port map(x=>p(140)(25),y=>p(141)(25),Cin=>p(142)(25),clock=>clock,reset=>reset,s=>p(222)(25),cout=>p(223)(26));
FA_ff_5909:FAff port map(x=>p(140)(26),y=>p(141)(26),Cin=>p(142)(26),clock=>clock,reset=>reset,s=>p(222)(26),cout=>p(223)(27));
FA_ff_5910:FAff port map(x=>p(140)(27),y=>p(141)(27),Cin=>p(142)(27),clock=>clock,reset=>reset,s=>p(222)(27),cout=>p(223)(28));
FA_ff_5911:FAff port map(x=>p(140)(28),y=>p(141)(28),Cin=>p(142)(28),clock=>clock,reset=>reset,s=>p(222)(28),cout=>p(223)(29));
FA_ff_5912:FAff port map(x=>p(140)(29),y=>p(141)(29),Cin=>p(142)(29),clock=>clock,reset=>reset,s=>p(222)(29),cout=>p(223)(30));
FA_ff_5913:FAff port map(x=>p(140)(30),y=>p(141)(30),Cin=>p(142)(30),clock=>clock,reset=>reset,s=>p(222)(30),cout=>p(223)(31));
FA_ff_5914:FAff port map(x=>p(140)(31),y=>p(141)(31),Cin=>p(142)(31),clock=>clock,reset=>reset,s=>p(222)(31),cout=>p(223)(32));
FA_ff_5915:FAff port map(x=>p(140)(32),y=>p(141)(32),Cin=>p(142)(32),clock=>clock,reset=>reset,s=>p(222)(32),cout=>p(223)(33));
FA_ff_5916:FAff port map(x=>p(140)(33),y=>p(141)(33),Cin=>p(142)(33),clock=>clock,reset=>reset,s=>p(222)(33),cout=>p(223)(34));
FA_ff_5917:FAff port map(x=>p(140)(34),y=>p(141)(34),Cin=>p(142)(34),clock=>clock,reset=>reset,s=>p(222)(34),cout=>p(223)(35));
FA_ff_5918:FAff port map(x=>p(140)(35),y=>p(141)(35),Cin=>p(142)(35),clock=>clock,reset=>reset,s=>p(222)(35),cout=>p(223)(36));
FA_ff_5919:FAff port map(x=>p(140)(36),y=>p(141)(36),Cin=>p(142)(36),clock=>clock,reset=>reset,s=>p(222)(36),cout=>p(223)(37));
FA_ff_5920:FAff port map(x=>p(140)(37),y=>p(141)(37),Cin=>p(142)(37),clock=>clock,reset=>reset,s=>p(222)(37),cout=>p(223)(38));
FA_ff_5921:FAff port map(x=>p(140)(38),y=>p(141)(38),Cin=>p(142)(38),clock=>clock,reset=>reset,s=>p(222)(38),cout=>p(223)(39));
FA_ff_5922:FAff port map(x=>p(140)(39),y=>p(141)(39),Cin=>p(142)(39),clock=>clock,reset=>reset,s=>p(222)(39),cout=>p(223)(40));
FA_ff_5923:FAff port map(x=>p(140)(40),y=>p(141)(40),Cin=>p(142)(40),clock=>clock,reset=>reset,s=>p(222)(40),cout=>p(223)(41));
FA_ff_5924:FAff port map(x=>p(140)(41),y=>p(141)(41),Cin=>p(142)(41),clock=>clock,reset=>reset,s=>p(222)(41),cout=>p(223)(42));
FA_ff_5925:FAff port map(x=>p(140)(42),y=>p(141)(42),Cin=>p(142)(42),clock=>clock,reset=>reset,s=>p(222)(42),cout=>p(223)(43));
FA_ff_5926:FAff port map(x=>p(140)(43),y=>p(141)(43),Cin=>p(142)(43),clock=>clock,reset=>reset,s=>p(222)(43),cout=>p(223)(44));
FA_ff_5927:FAff port map(x=>p(140)(44),y=>p(141)(44),Cin=>p(142)(44),clock=>clock,reset=>reset,s=>p(222)(44),cout=>p(223)(45));
FA_ff_5928:FAff port map(x=>p(140)(45),y=>p(141)(45),Cin=>p(142)(45),clock=>clock,reset=>reset,s=>p(222)(45),cout=>p(223)(46));
FA_ff_5929:FAff port map(x=>p(140)(46),y=>p(141)(46),Cin=>p(142)(46),clock=>clock,reset=>reset,s=>p(222)(46),cout=>p(223)(47));
FA_ff_5930:FAff port map(x=>p(140)(47),y=>p(141)(47),Cin=>p(142)(47),clock=>clock,reset=>reset,s=>p(222)(47),cout=>p(223)(48));
FA_ff_5931:FAff port map(x=>p(140)(48),y=>p(141)(48),Cin=>p(142)(48),clock=>clock,reset=>reset,s=>p(222)(48),cout=>p(223)(49));
FA_ff_5932:FAff port map(x=>p(140)(49),y=>p(141)(49),Cin=>p(142)(49),clock=>clock,reset=>reset,s=>p(222)(49),cout=>p(223)(50));
FA_ff_5933:FAff port map(x=>p(140)(50),y=>p(141)(50),Cin=>p(142)(50),clock=>clock,reset=>reset,s=>p(222)(50),cout=>p(223)(51));
FA_ff_5934:FAff port map(x=>p(140)(51),y=>p(141)(51),Cin=>p(142)(51),clock=>clock,reset=>reset,s=>p(222)(51),cout=>p(223)(52));
FA_ff_5935:FAff port map(x=>p(140)(52),y=>p(141)(52),Cin=>p(142)(52),clock=>clock,reset=>reset,s=>p(222)(52),cout=>p(223)(53));
FA_ff_5936:FAff port map(x=>p(140)(53),y=>p(141)(53),Cin=>p(142)(53),clock=>clock,reset=>reset,s=>p(222)(53),cout=>p(223)(54));
FA_ff_5937:FAff port map(x=>p(140)(54),y=>p(141)(54),Cin=>p(142)(54),clock=>clock,reset=>reset,s=>p(222)(54),cout=>p(223)(55));
FA_ff_5938:FAff port map(x=>p(140)(55),y=>p(141)(55),Cin=>p(142)(55),clock=>clock,reset=>reset,s=>p(222)(55),cout=>p(223)(56));
FA_ff_5939:FAff port map(x=>p(140)(56),y=>p(141)(56),Cin=>p(142)(56),clock=>clock,reset=>reset,s=>p(222)(56),cout=>p(223)(57));
FA_ff_5940:FAff port map(x=>p(140)(57),y=>p(141)(57),Cin=>p(142)(57),clock=>clock,reset=>reset,s=>p(222)(57),cout=>p(223)(58));
FA_ff_5941:FAff port map(x=>p(140)(58),y=>p(141)(58),Cin=>p(142)(58),clock=>clock,reset=>reset,s=>p(222)(58),cout=>p(223)(59));
FA_ff_5942:FAff port map(x=>p(140)(59),y=>p(141)(59),Cin=>p(142)(59),clock=>clock,reset=>reset,s=>p(222)(59),cout=>p(223)(60));
FA_ff_5943:FAff port map(x=>p(140)(60),y=>p(141)(60),Cin=>p(142)(60),clock=>clock,reset=>reset,s=>p(222)(60),cout=>p(223)(61));
FA_ff_5944:FAff port map(x=>p(140)(61),y=>p(141)(61),Cin=>p(142)(61),clock=>clock,reset=>reset,s=>p(222)(61),cout=>p(223)(62));
FA_ff_5945:FAff port map(x=>p(140)(62),y=>p(141)(62),Cin=>p(142)(62),clock=>clock,reset=>reset,s=>p(222)(62),cout=>p(223)(63));
FA_ff_5946:FAff port map(x=>p(140)(63),y=>p(141)(63),Cin=>p(142)(63),clock=>clock,reset=>reset,s=>p(222)(63),cout=>p(223)(64));
FA_ff_5947:FAff port map(x=>p(140)(64),y=>p(141)(64),Cin=>p(142)(64),clock=>clock,reset=>reset,s=>p(222)(64),cout=>p(223)(65));
FA_ff_5948:FAff port map(x=>p(140)(65),y=>p(141)(65),Cin=>p(142)(65),clock=>clock,reset=>reset,s=>p(222)(65),cout=>p(223)(66));
FA_ff_5949:FAff port map(x=>p(140)(66),y=>p(141)(66),Cin=>p(142)(66),clock=>clock,reset=>reset,s=>p(222)(66),cout=>p(223)(67));
FA_ff_5950:FAff port map(x=>p(140)(67),y=>p(141)(67),Cin=>p(142)(67),clock=>clock,reset=>reset,s=>p(222)(67),cout=>p(223)(68));
FA_ff_5951:FAff port map(x=>p(140)(68),y=>p(141)(68),Cin=>p(142)(68),clock=>clock,reset=>reset,s=>p(222)(68),cout=>p(223)(69));
FA_ff_5952:FAff port map(x=>p(140)(69),y=>p(141)(69),Cin=>p(142)(69),clock=>clock,reset=>reset,s=>p(222)(69),cout=>p(223)(70));
FA_ff_5953:FAff port map(x=>p(140)(70),y=>p(141)(70),Cin=>p(142)(70),clock=>clock,reset=>reset,s=>p(222)(70),cout=>p(223)(71));
FA_ff_5954:FAff port map(x=>p(140)(71),y=>p(141)(71),Cin=>p(142)(71),clock=>clock,reset=>reset,s=>p(222)(71),cout=>p(223)(72));
FA_ff_5955:FAff port map(x=>p(140)(72),y=>p(141)(72),Cin=>p(142)(72),clock=>clock,reset=>reset,s=>p(222)(72),cout=>p(223)(73));
FA_ff_5956:FAff port map(x=>p(140)(73),y=>p(141)(73),Cin=>p(142)(73),clock=>clock,reset=>reset,s=>p(222)(73),cout=>p(223)(74));
FA_ff_5957:FAff port map(x=>p(140)(74),y=>p(141)(74),Cin=>p(142)(74),clock=>clock,reset=>reset,s=>p(222)(74),cout=>p(223)(75));
FA_ff_5958:FAff port map(x=>p(140)(75),y=>p(141)(75),Cin=>p(142)(75),clock=>clock,reset=>reset,s=>p(222)(75),cout=>p(223)(76));
FA_ff_5959:FAff port map(x=>p(140)(76),y=>p(141)(76),Cin=>p(142)(76),clock=>clock,reset=>reset,s=>p(222)(76),cout=>p(223)(77));
FA_ff_5960:FAff port map(x=>p(140)(77),y=>p(141)(77),Cin=>p(142)(77),clock=>clock,reset=>reset,s=>p(222)(77),cout=>p(223)(78));
FA_ff_5961:FAff port map(x=>p(140)(78),y=>p(141)(78),Cin=>p(142)(78),clock=>clock,reset=>reset,s=>p(222)(78),cout=>p(223)(79));
FA_ff_5962:FAff port map(x=>p(140)(79),y=>p(141)(79),Cin=>p(142)(79),clock=>clock,reset=>reset,s=>p(222)(79),cout=>p(223)(80));
FA_ff_5963:FAff port map(x=>p(140)(80),y=>p(141)(80),Cin=>p(142)(80),clock=>clock,reset=>reset,s=>p(222)(80),cout=>p(223)(81));
FA_ff_5964:FAff port map(x=>p(140)(81),y=>p(141)(81),Cin=>p(142)(81),clock=>clock,reset=>reset,s=>p(222)(81),cout=>p(223)(82));
FA_ff_5965:FAff port map(x=>p(140)(82),y=>p(141)(82),Cin=>p(142)(82),clock=>clock,reset=>reset,s=>p(222)(82),cout=>p(223)(83));
FA_ff_5966:FAff port map(x=>p(140)(83),y=>p(141)(83),Cin=>p(142)(83),clock=>clock,reset=>reset,s=>p(222)(83),cout=>p(223)(84));
FA_ff_5967:FAff port map(x=>p(140)(84),y=>p(141)(84),Cin=>p(142)(84),clock=>clock,reset=>reset,s=>p(222)(84),cout=>p(223)(85));
FA_ff_5968:FAff port map(x=>p(140)(85),y=>p(141)(85),Cin=>p(142)(85),clock=>clock,reset=>reset,s=>p(222)(85),cout=>p(223)(86));
FA_ff_5969:FAff port map(x=>p(140)(86),y=>p(141)(86),Cin=>p(142)(86),clock=>clock,reset=>reset,s=>p(222)(86),cout=>p(223)(87));
FA_ff_5970:FAff port map(x=>p(140)(87),y=>p(141)(87),Cin=>p(142)(87),clock=>clock,reset=>reset,s=>p(222)(87),cout=>p(223)(88));
FA_ff_5971:FAff port map(x=>p(140)(88),y=>p(141)(88),Cin=>p(142)(88),clock=>clock,reset=>reset,s=>p(222)(88),cout=>p(223)(89));
FA_ff_5972:FAff port map(x=>p(140)(89),y=>p(141)(89),Cin=>p(142)(89),clock=>clock,reset=>reset,s=>p(222)(89),cout=>p(223)(90));
FA_ff_5973:FAff port map(x=>p(140)(90),y=>p(141)(90),Cin=>p(142)(90),clock=>clock,reset=>reset,s=>p(222)(90),cout=>p(223)(91));
FA_ff_5974:FAff port map(x=>p(140)(91),y=>p(141)(91),Cin=>p(142)(91),clock=>clock,reset=>reset,s=>p(222)(91),cout=>p(223)(92));
FA_ff_5975:FAff port map(x=>p(140)(92),y=>p(141)(92),Cin=>p(142)(92),clock=>clock,reset=>reset,s=>p(222)(92),cout=>p(223)(93));
FA_ff_5976:FAff port map(x=>p(140)(93),y=>p(141)(93),Cin=>p(142)(93),clock=>clock,reset=>reset,s=>p(222)(93),cout=>p(223)(94));
FA_ff_5977:FAff port map(x=>p(140)(94),y=>p(141)(94),Cin=>p(142)(94),clock=>clock,reset=>reset,s=>p(222)(94),cout=>p(223)(95));
FA_ff_5978:FAff port map(x=>p(140)(95),y=>p(141)(95),Cin=>p(142)(95),clock=>clock,reset=>reset,s=>p(222)(95),cout=>p(223)(96));
FA_ff_5979:FAff port map(x=>p(140)(96),y=>p(141)(96),Cin=>p(142)(96),clock=>clock,reset=>reset,s=>p(222)(96),cout=>p(223)(97));
FA_ff_5980:FAff port map(x=>p(140)(97),y=>p(141)(97),Cin=>p(142)(97),clock=>clock,reset=>reset,s=>p(222)(97),cout=>p(223)(98));
FA_ff_5981:FAff port map(x=>p(140)(98),y=>p(141)(98),Cin=>p(142)(98),clock=>clock,reset=>reset,s=>p(222)(98),cout=>p(223)(99));
FA_ff_5982:FAff port map(x=>p(140)(99),y=>p(141)(99),Cin=>p(142)(99),clock=>clock,reset=>reset,s=>p(222)(99),cout=>p(223)(100));
FA_ff_5983:FAff port map(x=>p(140)(100),y=>p(141)(100),Cin=>p(142)(100),clock=>clock,reset=>reset,s=>p(222)(100),cout=>p(223)(101));
FA_ff_5984:FAff port map(x=>p(140)(101),y=>p(141)(101),Cin=>p(142)(101),clock=>clock,reset=>reset,s=>p(222)(101),cout=>p(223)(102));
FA_ff_5985:FAff port map(x=>p(140)(102),y=>p(141)(102),Cin=>p(142)(102),clock=>clock,reset=>reset,s=>p(222)(102),cout=>p(223)(103));
FA_ff_5986:FAff port map(x=>p(140)(103),y=>p(141)(103),Cin=>p(142)(103),clock=>clock,reset=>reset,s=>p(222)(103),cout=>p(223)(104));
FA_ff_5987:FAff port map(x=>p(140)(104),y=>p(141)(104),Cin=>p(142)(104),clock=>clock,reset=>reset,s=>p(222)(104),cout=>p(223)(105));
FA_ff_5988:FAff port map(x=>p(140)(105),y=>p(141)(105),Cin=>p(142)(105),clock=>clock,reset=>reset,s=>p(222)(105),cout=>p(223)(106));
FA_ff_5989:FAff port map(x=>p(140)(106),y=>p(141)(106),Cin=>p(142)(106),clock=>clock,reset=>reset,s=>p(222)(106),cout=>p(223)(107));
FA_ff_5990:FAff port map(x=>p(140)(107),y=>p(141)(107),Cin=>p(142)(107),clock=>clock,reset=>reset,s=>p(222)(107),cout=>p(223)(108));
FA_ff_5991:FAff port map(x=>p(140)(108),y=>p(141)(108),Cin=>p(142)(108),clock=>clock,reset=>reset,s=>p(222)(108),cout=>p(223)(109));
FA_ff_5992:FAff port map(x=>p(140)(109),y=>p(141)(109),Cin=>p(142)(109),clock=>clock,reset=>reset,s=>p(222)(109),cout=>p(223)(110));
FA_ff_5993:FAff port map(x=>p(140)(110),y=>p(141)(110),Cin=>p(142)(110),clock=>clock,reset=>reset,s=>p(222)(110),cout=>p(223)(111));
FA_ff_5994:FAff port map(x=>p(140)(111),y=>p(141)(111),Cin=>p(142)(111),clock=>clock,reset=>reset,s=>p(222)(111),cout=>p(223)(112));
FA_ff_5995:FAff port map(x=>p(140)(112),y=>p(141)(112),Cin=>p(142)(112),clock=>clock,reset=>reset,s=>p(222)(112),cout=>p(223)(113));
FA_ff_5996:FAff port map(x=>p(140)(113),y=>p(141)(113),Cin=>p(142)(113),clock=>clock,reset=>reset,s=>p(222)(113),cout=>p(223)(114));
FA_ff_5997:FAff port map(x=>p(140)(114),y=>p(141)(114),Cin=>p(142)(114),clock=>clock,reset=>reset,s=>p(222)(114),cout=>p(223)(115));
FA_ff_5998:FAff port map(x=>p(140)(115),y=>p(141)(115),Cin=>p(142)(115),clock=>clock,reset=>reset,s=>p(222)(115),cout=>p(223)(116));
FA_ff_5999:FAff port map(x=>p(140)(116),y=>p(141)(116),Cin=>p(142)(116),clock=>clock,reset=>reset,s=>p(222)(116),cout=>p(223)(117));
FA_ff_6000:FAff port map(x=>p(140)(117),y=>p(141)(117),Cin=>p(142)(117),clock=>clock,reset=>reset,s=>p(222)(117),cout=>p(223)(118));
FA_ff_6001:FAff port map(x=>p(140)(118),y=>p(141)(118),Cin=>p(142)(118),clock=>clock,reset=>reset,s=>p(222)(118),cout=>p(223)(119));
FA_ff_6002:FAff port map(x=>p(140)(119),y=>p(141)(119),Cin=>p(142)(119),clock=>clock,reset=>reset,s=>p(222)(119),cout=>p(223)(120));
FA_ff_6003:FAff port map(x=>p(140)(120),y=>p(141)(120),Cin=>p(142)(120),clock=>clock,reset=>reset,s=>p(222)(120),cout=>p(223)(121));
FA_ff_6004:FAff port map(x=>p(140)(121),y=>p(141)(121),Cin=>p(142)(121),clock=>clock,reset=>reset,s=>p(222)(121),cout=>p(223)(122));
FA_ff_6005:FAff port map(x=>p(140)(122),y=>p(141)(122),Cin=>p(142)(122),clock=>clock,reset=>reset,s=>p(222)(122),cout=>p(223)(123));
FA_ff_6006:FAff port map(x=>p(140)(123),y=>p(141)(123),Cin=>p(142)(123),clock=>clock,reset=>reset,s=>p(222)(123),cout=>p(223)(124));
FA_ff_6007:FAff port map(x=>p(140)(124),y=>p(141)(124),Cin=>p(142)(124),clock=>clock,reset=>reset,s=>p(222)(124),cout=>p(223)(125));
FA_ff_6008:FAff port map(x=>p(140)(125),y=>p(141)(125),Cin=>p(142)(125),clock=>clock,reset=>reset,s=>p(222)(125),cout=>p(223)(126));
FA_ff_6009:FAff port map(x=>p(140)(126),y=>p(141)(126),Cin=>p(142)(126),clock=>clock,reset=>reset,s=>p(222)(126),cout=>p(223)(127));
FA_ff_6010:FAff port map(x=>p(140)(127),y=>p(141)(127),Cin=>p(142)(127),clock=>clock,reset=>reset,s=>p(222)(127),cout=>p(223)(128));
p(222)(128)<=p(141)(128);
p(224)(0)<=p(144)(0);
FA_ff_6011:FAff port map(x=>p(143)(1),y=>p(144)(1),Cin=>p(145)(1),clock=>clock,reset=>reset,s=>p(224)(1),cout=>p(225)(2));
FA_ff_6012:FAff port map(x=>p(143)(2),y=>p(144)(2),Cin=>p(145)(2),clock=>clock,reset=>reset,s=>p(224)(2),cout=>p(225)(3));
FA_ff_6013:FAff port map(x=>p(143)(3),y=>p(144)(3),Cin=>p(145)(3),clock=>clock,reset=>reset,s=>p(224)(3),cout=>p(225)(4));
FA_ff_6014:FAff port map(x=>p(143)(4),y=>p(144)(4),Cin=>p(145)(4),clock=>clock,reset=>reset,s=>p(224)(4),cout=>p(225)(5));
FA_ff_6015:FAff port map(x=>p(143)(5),y=>p(144)(5),Cin=>p(145)(5),clock=>clock,reset=>reset,s=>p(224)(5),cout=>p(225)(6));
FA_ff_6016:FAff port map(x=>p(143)(6),y=>p(144)(6),Cin=>p(145)(6),clock=>clock,reset=>reset,s=>p(224)(6),cout=>p(225)(7));
FA_ff_6017:FAff port map(x=>p(143)(7),y=>p(144)(7),Cin=>p(145)(7),clock=>clock,reset=>reset,s=>p(224)(7),cout=>p(225)(8));
FA_ff_6018:FAff port map(x=>p(143)(8),y=>p(144)(8),Cin=>p(145)(8),clock=>clock,reset=>reset,s=>p(224)(8),cout=>p(225)(9));
FA_ff_6019:FAff port map(x=>p(143)(9),y=>p(144)(9),Cin=>p(145)(9),clock=>clock,reset=>reset,s=>p(224)(9),cout=>p(225)(10));
FA_ff_6020:FAff port map(x=>p(143)(10),y=>p(144)(10),Cin=>p(145)(10),clock=>clock,reset=>reset,s=>p(224)(10),cout=>p(225)(11));
FA_ff_6021:FAff port map(x=>p(143)(11),y=>p(144)(11),Cin=>p(145)(11),clock=>clock,reset=>reset,s=>p(224)(11),cout=>p(225)(12));
FA_ff_6022:FAff port map(x=>p(143)(12),y=>p(144)(12),Cin=>p(145)(12),clock=>clock,reset=>reset,s=>p(224)(12),cout=>p(225)(13));
FA_ff_6023:FAff port map(x=>p(143)(13),y=>p(144)(13),Cin=>p(145)(13),clock=>clock,reset=>reset,s=>p(224)(13),cout=>p(225)(14));
FA_ff_6024:FAff port map(x=>p(143)(14),y=>p(144)(14),Cin=>p(145)(14),clock=>clock,reset=>reset,s=>p(224)(14),cout=>p(225)(15));
FA_ff_6025:FAff port map(x=>p(143)(15),y=>p(144)(15),Cin=>p(145)(15),clock=>clock,reset=>reset,s=>p(224)(15),cout=>p(225)(16));
FA_ff_6026:FAff port map(x=>p(143)(16),y=>p(144)(16),Cin=>p(145)(16),clock=>clock,reset=>reset,s=>p(224)(16),cout=>p(225)(17));
FA_ff_6027:FAff port map(x=>p(143)(17),y=>p(144)(17),Cin=>p(145)(17),clock=>clock,reset=>reset,s=>p(224)(17),cout=>p(225)(18));
FA_ff_6028:FAff port map(x=>p(143)(18),y=>p(144)(18),Cin=>p(145)(18),clock=>clock,reset=>reset,s=>p(224)(18),cout=>p(225)(19));
FA_ff_6029:FAff port map(x=>p(143)(19),y=>p(144)(19),Cin=>p(145)(19),clock=>clock,reset=>reset,s=>p(224)(19),cout=>p(225)(20));
FA_ff_6030:FAff port map(x=>p(143)(20),y=>p(144)(20),Cin=>p(145)(20),clock=>clock,reset=>reset,s=>p(224)(20),cout=>p(225)(21));
FA_ff_6031:FAff port map(x=>p(143)(21),y=>p(144)(21),Cin=>p(145)(21),clock=>clock,reset=>reset,s=>p(224)(21),cout=>p(225)(22));
FA_ff_6032:FAff port map(x=>p(143)(22),y=>p(144)(22),Cin=>p(145)(22),clock=>clock,reset=>reset,s=>p(224)(22),cout=>p(225)(23));
FA_ff_6033:FAff port map(x=>p(143)(23),y=>p(144)(23),Cin=>p(145)(23),clock=>clock,reset=>reset,s=>p(224)(23),cout=>p(225)(24));
FA_ff_6034:FAff port map(x=>p(143)(24),y=>p(144)(24),Cin=>p(145)(24),clock=>clock,reset=>reset,s=>p(224)(24),cout=>p(225)(25));
FA_ff_6035:FAff port map(x=>p(143)(25),y=>p(144)(25),Cin=>p(145)(25),clock=>clock,reset=>reset,s=>p(224)(25),cout=>p(225)(26));
FA_ff_6036:FAff port map(x=>p(143)(26),y=>p(144)(26),Cin=>p(145)(26),clock=>clock,reset=>reset,s=>p(224)(26),cout=>p(225)(27));
FA_ff_6037:FAff port map(x=>p(143)(27),y=>p(144)(27),Cin=>p(145)(27),clock=>clock,reset=>reset,s=>p(224)(27),cout=>p(225)(28));
FA_ff_6038:FAff port map(x=>p(143)(28),y=>p(144)(28),Cin=>p(145)(28),clock=>clock,reset=>reset,s=>p(224)(28),cout=>p(225)(29));
FA_ff_6039:FAff port map(x=>p(143)(29),y=>p(144)(29),Cin=>p(145)(29),clock=>clock,reset=>reset,s=>p(224)(29),cout=>p(225)(30));
FA_ff_6040:FAff port map(x=>p(143)(30),y=>p(144)(30),Cin=>p(145)(30),clock=>clock,reset=>reset,s=>p(224)(30),cout=>p(225)(31));
FA_ff_6041:FAff port map(x=>p(143)(31),y=>p(144)(31),Cin=>p(145)(31),clock=>clock,reset=>reset,s=>p(224)(31),cout=>p(225)(32));
FA_ff_6042:FAff port map(x=>p(143)(32),y=>p(144)(32),Cin=>p(145)(32),clock=>clock,reset=>reset,s=>p(224)(32),cout=>p(225)(33));
FA_ff_6043:FAff port map(x=>p(143)(33),y=>p(144)(33),Cin=>p(145)(33),clock=>clock,reset=>reset,s=>p(224)(33),cout=>p(225)(34));
FA_ff_6044:FAff port map(x=>p(143)(34),y=>p(144)(34),Cin=>p(145)(34),clock=>clock,reset=>reset,s=>p(224)(34),cout=>p(225)(35));
FA_ff_6045:FAff port map(x=>p(143)(35),y=>p(144)(35),Cin=>p(145)(35),clock=>clock,reset=>reset,s=>p(224)(35),cout=>p(225)(36));
FA_ff_6046:FAff port map(x=>p(143)(36),y=>p(144)(36),Cin=>p(145)(36),clock=>clock,reset=>reset,s=>p(224)(36),cout=>p(225)(37));
FA_ff_6047:FAff port map(x=>p(143)(37),y=>p(144)(37),Cin=>p(145)(37),clock=>clock,reset=>reset,s=>p(224)(37),cout=>p(225)(38));
FA_ff_6048:FAff port map(x=>p(143)(38),y=>p(144)(38),Cin=>p(145)(38),clock=>clock,reset=>reset,s=>p(224)(38),cout=>p(225)(39));
FA_ff_6049:FAff port map(x=>p(143)(39),y=>p(144)(39),Cin=>p(145)(39),clock=>clock,reset=>reset,s=>p(224)(39),cout=>p(225)(40));
FA_ff_6050:FAff port map(x=>p(143)(40),y=>p(144)(40),Cin=>p(145)(40),clock=>clock,reset=>reset,s=>p(224)(40),cout=>p(225)(41));
FA_ff_6051:FAff port map(x=>p(143)(41),y=>p(144)(41),Cin=>p(145)(41),clock=>clock,reset=>reset,s=>p(224)(41),cout=>p(225)(42));
FA_ff_6052:FAff port map(x=>p(143)(42),y=>p(144)(42),Cin=>p(145)(42),clock=>clock,reset=>reset,s=>p(224)(42),cout=>p(225)(43));
FA_ff_6053:FAff port map(x=>p(143)(43),y=>p(144)(43),Cin=>p(145)(43),clock=>clock,reset=>reset,s=>p(224)(43),cout=>p(225)(44));
FA_ff_6054:FAff port map(x=>p(143)(44),y=>p(144)(44),Cin=>p(145)(44),clock=>clock,reset=>reset,s=>p(224)(44),cout=>p(225)(45));
FA_ff_6055:FAff port map(x=>p(143)(45),y=>p(144)(45),Cin=>p(145)(45),clock=>clock,reset=>reset,s=>p(224)(45),cout=>p(225)(46));
FA_ff_6056:FAff port map(x=>p(143)(46),y=>p(144)(46),Cin=>p(145)(46),clock=>clock,reset=>reset,s=>p(224)(46),cout=>p(225)(47));
FA_ff_6057:FAff port map(x=>p(143)(47),y=>p(144)(47),Cin=>p(145)(47),clock=>clock,reset=>reset,s=>p(224)(47),cout=>p(225)(48));
FA_ff_6058:FAff port map(x=>p(143)(48),y=>p(144)(48),Cin=>p(145)(48),clock=>clock,reset=>reset,s=>p(224)(48),cout=>p(225)(49));
FA_ff_6059:FAff port map(x=>p(143)(49),y=>p(144)(49),Cin=>p(145)(49),clock=>clock,reset=>reset,s=>p(224)(49),cout=>p(225)(50));
FA_ff_6060:FAff port map(x=>p(143)(50),y=>p(144)(50),Cin=>p(145)(50),clock=>clock,reset=>reset,s=>p(224)(50),cout=>p(225)(51));
FA_ff_6061:FAff port map(x=>p(143)(51),y=>p(144)(51),Cin=>p(145)(51),clock=>clock,reset=>reset,s=>p(224)(51),cout=>p(225)(52));
FA_ff_6062:FAff port map(x=>p(143)(52),y=>p(144)(52),Cin=>p(145)(52),clock=>clock,reset=>reset,s=>p(224)(52),cout=>p(225)(53));
FA_ff_6063:FAff port map(x=>p(143)(53),y=>p(144)(53),Cin=>p(145)(53),clock=>clock,reset=>reset,s=>p(224)(53),cout=>p(225)(54));
FA_ff_6064:FAff port map(x=>p(143)(54),y=>p(144)(54),Cin=>p(145)(54),clock=>clock,reset=>reset,s=>p(224)(54),cout=>p(225)(55));
FA_ff_6065:FAff port map(x=>p(143)(55),y=>p(144)(55),Cin=>p(145)(55),clock=>clock,reset=>reset,s=>p(224)(55),cout=>p(225)(56));
FA_ff_6066:FAff port map(x=>p(143)(56),y=>p(144)(56),Cin=>p(145)(56),clock=>clock,reset=>reset,s=>p(224)(56),cout=>p(225)(57));
FA_ff_6067:FAff port map(x=>p(143)(57),y=>p(144)(57),Cin=>p(145)(57),clock=>clock,reset=>reset,s=>p(224)(57),cout=>p(225)(58));
FA_ff_6068:FAff port map(x=>p(143)(58),y=>p(144)(58),Cin=>p(145)(58),clock=>clock,reset=>reset,s=>p(224)(58),cout=>p(225)(59));
FA_ff_6069:FAff port map(x=>p(143)(59),y=>p(144)(59),Cin=>p(145)(59),clock=>clock,reset=>reset,s=>p(224)(59),cout=>p(225)(60));
FA_ff_6070:FAff port map(x=>p(143)(60),y=>p(144)(60),Cin=>p(145)(60),clock=>clock,reset=>reset,s=>p(224)(60),cout=>p(225)(61));
FA_ff_6071:FAff port map(x=>p(143)(61),y=>p(144)(61),Cin=>p(145)(61),clock=>clock,reset=>reset,s=>p(224)(61),cout=>p(225)(62));
FA_ff_6072:FAff port map(x=>p(143)(62),y=>p(144)(62),Cin=>p(145)(62),clock=>clock,reset=>reset,s=>p(224)(62),cout=>p(225)(63));
FA_ff_6073:FAff port map(x=>p(143)(63),y=>p(144)(63),Cin=>p(145)(63),clock=>clock,reset=>reset,s=>p(224)(63),cout=>p(225)(64));
FA_ff_6074:FAff port map(x=>p(143)(64),y=>p(144)(64),Cin=>p(145)(64),clock=>clock,reset=>reset,s=>p(224)(64),cout=>p(225)(65));
FA_ff_6075:FAff port map(x=>p(143)(65),y=>p(144)(65),Cin=>p(145)(65),clock=>clock,reset=>reset,s=>p(224)(65),cout=>p(225)(66));
FA_ff_6076:FAff port map(x=>p(143)(66),y=>p(144)(66),Cin=>p(145)(66),clock=>clock,reset=>reset,s=>p(224)(66),cout=>p(225)(67));
FA_ff_6077:FAff port map(x=>p(143)(67),y=>p(144)(67),Cin=>p(145)(67),clock=>clock,reset=>reset,s=>p(224)(67),cout=>p(225)(68));
FA_ff_6078:FAff port map(x=>p(143)(68),y=>p(144)(68),Cin=>p(145)(68),clock=>clock,reset=>reset,s=>p(224)(68),cout=>p(225)(69));
FA_ff_6079:FAff port map(x=>p(143)(69),y=>p(144)(69),Cin=>p(145)(69),clock=>clock,reset=>reset,s=>p(224)(69),cout=>p(225)(70));
FA_ff_6080:FAff port map(x=>p(143)(70),y=>p(144)(70),Cin=>p(145)(70),clock=>clock,reset=>reset,s=>p(224)(70),cout=>p(225)(71));
FA_ff_6081:FAff port map(x=>p(143)(71),y=>p(144)(71),Cin=>p(145)(71),clock=>clock,reset=>reset,s=>p(224)(71),cout=>p(225)(72));
FA_ff_6082:FAff port map(x=>p(143)(72),y=>p(144)(72),Cin=>p(145)(72),clock=>clock,reset=>reset,s=>p(224)(72),cout=>p(225)(73));
FA_ff_6083:FAff port map(x=>p(143)(73),y=>p(144)(73),Cin=>p(145)(73),clock=>clock,reset=>reset,s=>p(224)(73),cout=>p(225)(74));
FA_ff_6084:FAff port map(x=>p(143)(74),y=>p(144)(74),Cin=>p(145)(74),clock=>clock,reset=>reset,s=>p(224)(74),cout=>p(225)(75));
FA_ff_6085:FAff port map(x=>p(143)(75),y=>p(144)(75),Cin=>p(145)(75),clock=>clock,reset=>reset,s=>p(224)(75),cout=>p(225)(76));
FA_ff_6086:FAff port map(x=>p(143)(76),y=>p(144)(76),Cin=>p(145)(76),clock=>clock,reset=>reset,s=>p(224)(76),cout=>p(225)(77));
FA_ff_6087:FAff port map(x=>p(143)(77),y=>p(144)(77),Cin=>p(145)(77),clock=>clock,reset=>reset,s=>p(224)(77),cout=>p(225)(78));
FA_ff_6088:FAff port map(x=>p(143)(78),y=>p(144)(78),Cin=>p(145)(78),clock=>clock,reset=>reset,s=>p(224)(78),cout=>p(225)(79));
FA_ff_6089:FAff port map(x=>p(143)(79),y=>p(144)(79),Cin=>p(145)(79),clock=>clock,reset=>reset,s=>p(224)(79),cout=>p(225)(80));
FA_ff_6090:FAff port map(x=>p(143)(80),y=>p(144)(80),Cin=>p(145)(80),clock=>clock,reset=>reset,s=>p(224)(80),cout=>p(225)(81));
FA_ff_6091:FAff port map(x=>p(143)(81),y=>p(144)(81),Cin=>p(145)(81),clock=>clock,reset=>reset,s=>p(224)(81),cout=>p(225)(82));
FA_ff_6092:FAff port map(x=>p(143)(82),y=>p(144)(82),Cin=>p(145)(82),clock=>clock,reset=>reset,s=>p(224)(82),cout=>p(225)(83));
FA_ff_6093:FAff port map(x=>p(143)(83),y=>p(144)(83),Cin=>p(145)(83),clock=>clock,reset=>reset,s=>p(224)(83),cout=>p(225)(84));
FA_ff_6094:FAff port map(x=>p(143)(84),y=>p(144)(84),Cin=>p(145)(84),clock=>clock,reset=>reset,s=>p(224)(84),cout=>p(225)(85));
FA_ff_6095:FAff port map(x=>p(143)(85),y=>p(144)(85),Cin=>p(145)(85),clock=>clock,reset=>reset,s=>p(224)(85),cout=>p(225)(86));
FA_ff_6096:FAff port map(x=>p(143)(86),y=>p(144)(86),Cin=>p(145)(86),clock=>clock,reset=>reset,s=>p(224)(86),cout=>p(225)(87));
FA_ff_6097:FAff port map(x=>p(143)(87),y=>p(144)(87),Cin=>p(145)(87),clock=>clock,reset=>reset,s=>p(224)(87),cout=>p(225)(88));
FA_ff_6098:FAff port map(x=>p(143)(88),y=>p(144)(88),Cin=>p(145)(88),clock=>clock,reset=>reset,s=>p(224)(88),cout=>p(225)(89));
FA_ff_6099:FAff port map(x=>p(143)(89),y=>p(144)(89),Cin=>p(145)(89),clock=>clock,reset=>reset,s=>p(224)(89),cout=>p(225)(90));
FA_ff_6100:FAff port map(x=>p(143)(90),y=>p(144)(90),Cin=>p(145)(90),clock=>clock,reset=>reset,s=>p(224)(90),cout=>p(225)(91));
FA_ff_6101:FAff port map(x=>p(143)(91),y=>p(144)(91),Cin=>p(145)(91),clock=>clock,reset=>reset,s=>p(224)(91),cout=>p(225)(92));
FA_ff_6102:FAff port map(x=>p(143)(92),y=>p(144)(92),Cin=>p(145)(92),clock=>clock,reset=>reset,s=>p(224)(92),cout=>p(225)(93));
FA_ff_6103:FAff port map(x=>p(143)(93),y=>p(144)(93),Cin=>p(145)(93),clock=>clock,reset=>reset,s=>p(224)(93),cout=>p(225)(94));
FA_ff_6104:FAff port map(x=>p(143)(94),y=>p(144)(94),Cin=>p(145)(94),clock=>clock,reset=>reset,s=>p(224)(94),cout=>p(225)(95));
FA_ff_6105:FAff port map(x=>p(143)(95),y=>p(144)(95),Cin=>p(145)(95),clock=>clock,reset=>reset,s=>p(224)(95),cout=>p(225)(96));
FA_ff_6106:FAff port map(x=>p(143)(96),y=>p(144)(96),Cin=>p(145)(96),clock=>clock,reset=>reset,s=>p(224)(96),cout=>p(225)(97));
FA_ff_6107:FAff port map(x=>p(143)(97),y=>p(144)(97),Cin=>p(145)(97),clock=>clock,reset=>reset,s=>p(224)(97),cout=>p(225)(98));
FA_ff_6108:FAff port map(x=>p(143)(98),y=>p(144)(98),Cin=>p(145)(98),clock=>clock,reset=>reset,s=>p(224)(98),cout=>p(225)(99));
FA_ff_6109:FAff port map(x=>p(143)(99),y=>p(144)(99),Cin=>p(145)(99),clock=>clock,reset=>reset,s=>p(224)(99),cout=>p(225)(100));
FA_ff_6110:FAff port map(x=>p(143)(100),y=>p(144)(100),Cin=>p(145)(100),clock=>clock,reset=>reset,s=>p(224)(100),cout=>p(225)(101));
FA_ff_6111:FAff port map(x=>p(143)(101),y=>p(144)(101),Cin=>p(145)(101),clock=>clock,reset=>reset,s=>p(224)(101),cout=>p(225)(102));
FA_ff_6112:FAff port map(x=>p(143)(102),y=>p(144)(102),Cin=>p(145)(102),clock=>clock,reset=>reset,s=>p(224)(102),cout=>p(225)(103));
FA_ff_6113:FAff port map(x=>p(143)(103),y=>p(144)(103),Cin=>p(145)(103),clock=>clock,reset=>reset,s=>p(224)(103),cout=>p(225)(104));
FA_ff_6114:FAff port map(x=>p(143)(104),y=>p(144)(104),Cin=>p(145)(104),clock=>clock,reset=>reset,s=>p(224)(104),cout=>p(225)(105));
FA_ff_6115:FAff port map(x=>p(143)(105),y=>p(144)(105),Cin=>p(145)(105),clock=>clock,reset=>reset,s=>p(224)(105),cout=>p(225)(106));
FA_ff_6116:FAff port map(x=>p(143)(106),y=>p(144)(106),Cin=>p(145)(106),clock=>clock,reset=>reset,s=>p(224)(106),cout=>p(225)(107));
FA_ff_6117:FAff port map(x=>p(143)(107),y=>p(144)(107),Cin=>p(145)(107),clock=>clock,reset=>reset,s=>p(224)(107),cout=>p(225)(108));
FA_ff_6118:FAff port map(x=>p(143)(108),y=>p(144)(108),Cin=>p(145)(108),clock=>clock,reset=>reset,s=>p(224)(108),cout=>p(225)(109));
FA_ff_6119:FAff port map(x=>p(143)(109),y=>p(144)(109),Cin=>p(145)(109),clock=>clock,reset=>reset,s=>p(224)(109),cout=>p(225)(110));
FA_ff_6120:FAff port map(x=>p(143)(110),y=>p(144)(110),Cin=>p(145)(110),clock=>clock,reset=>reset,s=>p(224)(110),cout=>p(225)(111));
FA_ff_6121:FAff port map(x=>p(143)(111),y=>p(144)(111),Cin=>p(145)(111),clock=>clock,reset=>reset,s=>p(224)(111),cout=>p(225)(112));
FA_ff_6122:FAff port map(x=>p(143)(112),y=>p(144)(112),Cin=>p(145)(112),clock=>clock,reset=>reset,s=>p(224)(112),cout=>p(225)(113));
FA_ff_6123:FAff port map(x=>p(143)(113),y=>p(144)(113),Cin=>p(145)(113),clock=>clock,reset=>reset,s=>p(224)(113),cout=>p(225)(114));
FA_ff_6124:FAff port map(x=>p(143)(114),y=>p(144)(114),Cin=>p(145)(114),clock=>clock,reset=>reset,s=>p(224)(114),cout=>p(225)(115));
FA_ff_6125:FAff port map(x=>p(143)(115),y=>p(144)(115),Cin=>p(145)(115),clock=>clock,reset=>reset,s=>p(224)(115),cout=>p(225)(116));
FA_ff_6126:FAff port map(x=>p(143)(116),y=>p(144)(116),Cin=>p(145)(116),clock=>clock,reset=>reset,s=>p(224)(116),cout=>p(225)(117));
FA_ff_6127:FAff port map(x=>p(143)(117),y=>p(144)(117),Cin=>p(145)(117),clock=>clock,reset=>reset,s=>p(224)(117),cout=>p(225)(118));
FA_ff_6128:FAff port map(x=>p(143)(118),y=>p(144)(118),Cin=>p(145)(118),clock=>clock,reset=>reset,s=>p(224)(118),cout=>p(225)(119));
FA_ff_6129:FAff port map(x=>p(143)(119),y=>p(144)(119),Cin=>p(145)(119),clock=>clock,reset=>reset,s=>p(224)(119),cout=>p(225)(120));
FA_ff_6130:FAff port map(x=>p(143)(120),y=>p(144)(120),Cin=>p(145)(120),clock=>clock,reset=>reset,s=>p(224)(120),cout=>p(225)(121));
FA_ff_6131:FAff port map(x=>p(143)(121),y=>p(144)(121),Cin=>p(145)(121),clock=>clock,reset=>reset,s=>p(224)(121),cout=>p(225)(122));
FA_ff_6132:FAff port map(x=>p(143)(122),y=>p(144)(122),Cin=>p(145)(122),clock=>clock,reset=>reset,s=>p(224)(122),cout=>p(225)(123));
FA_ff_6133:FAff port map(x=>p(143)(123),y=>p(144)(123),Cin=>p(145)(123),clock=>clock,reset=>reset,s=>p(224)(123),cout=>p(225)(124));
FA_ff_6134:FAff port map(x=>p(143)(124),y=>p(144)(124),Cin=>p(145)(124),clock=>clock,reset=>reset,s=>p(224)(124),cout=>p(225)(125));
FA_ff_6135:FAff port map(x=>p(143)(125),y=>p(144)(125),Cin=>p(145)(125),clock=>clock,reset=>reset,s=>p(224)(125),cout=>p(225)(126));
FA_ff_6136:FAff port map(x=>p(143)(126),y=>p(144)(126),Cin=>p(145)(126),clock=>clock,reset=>reset,s=>p(224)(126),cout=>p(225)(127));
FA_ff_6137:FAff port map(x=>p(143)(127),y=>p(144)(127),Cin=>p(145)(127),clock=>clock,reset=>reset,s=>p(224)(127),cout=>p(225)(128));
HA_ff_5:HAff port map(x=>p(143)(128),y=>p(145)(128),clock=>clock,reset=>reset,s=>p(224)(128),c=>p(225)(129));
HA_ff_6:HAff port map(x=>p(146)(0),y=>p(148)(0),clock=>clock,reset=>reset,s=>p(226)(0),c=>p(227)(1));
FA_ff_6138:FAff port map(x=>p(146)(1),y=>p(147)(1),Cin=>p(148)(1),clock=>clock,reset=>reset,s=>p(226)(1),cout=>p(227)(2));
FA_ff_6139:FAff port map(x=>p(146)(2),y=>p(147)(2),Cin=>p(148)(2),clock=>clock,reset=>reset,s=>p(226)(2),cout=>p(227)(3));
FA_ff_6140:FAff port map(x=>p(146)(3),y=>p(147)(3),Cin=>p(148)(3),clock=>clock,reset=>reset,s=>p(226)(3),cout=>p(227)(4));
FA_ff_6141:FAff port map(x=>p(146)(4),y=>p(147)(4),Cin=>p(148)(4),clock=>clock,reset=>reset,s=>p(226)(4),cout=>p(227)(5));
FA_ff_6142:FAff port map(x=>p(146)(5),y=>p(147)(5),Cin=>p(148)(5),clock=>clock,reset=>reset,s=>p(226)(5),cout=>p(227)(6));
FA_ff_6143:FAff port map(x=>p(146)(6),y=>p(147)(6),Cin=>p(148)(6),clock=>clock,reset=>reset,s=>p(226)(6),cout=>p(227)(7));
FA_ff_6144:FAff port map(x=>p(146)(7),y=>p(147)(7),Cin=>p(148)(7),clock=>clock,reset=>reset,s=>p(226)(7),cout=>p(227)(8));
FA_ff_6145:FAff port map(x=>p(146)(8),y=>p(147)(8),Cin=>p(148)(8),clock=>clock,reset=>reset,s=>p(226)(8),cout=>p(227)(9));
FA_ff_6146:FAff port map(x=>p(146)(9),y=>p(147)(9),Cin=>p(148)(9),clock=>clock,reset=>reset,s=>p(226)(9),cout=>p(227)(10));
FA_ff_6147:FAff port map(x=>p(146)(10),y=>p(147)(10),Cin=>p(148)(10),clock=>clock,reset=>reset,s=>p(226)(10),cout=>p(227)(11));
FA_ff_6148:FAff port map(x=>p(146)(11),y=>p(147)(11),Cin=>p(148)(11),clock=>clock,reset=>reset,s=>p(226)(11),cout=>p(227)(12));
FA_ff_6149:FAff port map(x=>p(146)(12),y=>p(147)(12),Cin=>p(148)(12),clock=>clock,reset=>reset,s=>p(226)(12),cout=>p(227)(13));
FA_ff_6150:FAff port map(x=>p(146)(13),y=>p(147)(13),Cin=>p(148)(13),clock=>clock,reset=>reset,s=>p(226)(13),cout=>p(227)(14));
FA_ff_6151:FAff port map(x=>p(146)(14),y=>p(147)(14),Cin=>p(148)(14),clock=>clock,reset=>reset,s=>p(226)(14),cout=>p(227)(15));
FA_ff_6152:FAff port map(x=>p(146)(15),y=>p(147)(15),Cin=>p(148)(15),clock=>clock,reset=>reset,s=>p(226)(15),cout=>p(227)(16));
FA_ff_6153:FAff port map(x=>p(146)(16),y=>p(147)(16),Cin=>p(148)(16),clock=>clock,reset=>reset,s=>p(226)(16),cout=>p(227)(17));
FA_ff_6154:FAff port map(x=>p(146)(17),y=>p(147)(17),Cin=>p(148)(17),clock=>clock,reset=>reset,s=>p(226)(17),cout=>p(227)(18));
FA_ff_6155:FAff port map(x=>p(146)(18),y=>p(147)(18),Cin=>p(148)(18),clock=>clock,reset=>reset,s=>p(226)(18),cout=>p(227)(19));
FA_ff_6156:FAff port map(x=>p(146)(19),y=>p(147)(19),Cin=>p(148)(19),clock=>clock,reset=>reset,s=>p(226)(19),cout=>p(227)(20));
FA_ff_6157:FAff port map(x=>p(146)(20),y=>p(147)(20),Cin=>p(148)(20),clock=>clock,reset=>reset,s=>p(226)(20),cout=>p(227)(21));
FA_ff_6158:FAff port map(x=>p(146)(21),y=>p(147)(21),Cin=>p(148)(21),clock=>clock,reset=>reset,s=>p(226)(21),cout=>p(227)(22));
FA_ff_6159:FAff port map(x=>p(146)(22),y=>p(147)(22),Cin=>p(148)(22),clock=>clock,reset=>reset,s=>p(226)(22),cout=>p(227)(23));
FA_ff_6160:FAff port map(x=>p(146)(23),y=>p(147)(23),Cin=>p(148)(23),clock=>clock,reset=>reset,s=>p(226)(23),cout=>p(227)(24));
FA_ff_6161:FAff port map(x=>p(146)(24),y=>p(147)(24),Cin=>p(148)(24),clock=>clock,reset=>reset,s=>p(226)(24),cout=>p(227)(25));
FA_ff_6162:FAff port map(x=>p(146)(25),y=>p(147)(25),Cin=>p(148)(25),clock=>clock,reset=>reset,s=>p(226)(25),cout=>p(227)(26));
FA_ff_6163:FAff port map(x=>p(146)(26),y=>p(147)(26),Cin=>p(148)(26),clock=>clock,reset=>reset,s=>p(226)(26),cout=>p(227)(27));
FA_ff_6164:FAff port map(x=>p(146)(27),y=>p(147)(27),Cin=>p(148)(27),clock=>clock,reset=>reset,s=>p(226)(27),cout=>p(227)(28));
FA_ff_6165:FAff port map(x=>p(146)(28),y=>p(147)(28),Cin=>p(148)(28),clock=>clock,reset=>reset,s=>p(226)(28),cout=>p(227)(29));
FA_ff_6166:FAff port map(x=>p(146)(29),y=>p(147)(29),Cin=>p(148)(29),clock=>clock,reset=>reset,s=>p(226)(29),cout=>p(227)(30));
FA_ff_6167:FAff port map(x=>p(146)(30),y=>p(147)(30),Cin=>p(148)(30),clock=>clock,reset=>reset,s=>p(226)(30),cout=>p(227)(31));
FA_ff_6168:FAff port map(x=>p(146)(31),y=>p(147)(31),Cin=>p(148)(31),clock=>clock,reset=>reset,s=>p(226)(31),cout=>p(227)(32));
FA_ff_6169:FAff port map(x=>p(146)(32),y=>p(147)(32),Cin=>p(148)(32),clock=>clock,reset=>reset,s=>p(226)(32),cout=>p(227)(33));
FA_ff_6170:FAff port map(x=>p(146)(33),y=>p(147)(33),Cin=>p(148)(33),clock=>clock,reset=>reset,s=>p(226)(33),cout=>p(227)(34));
FA_ff_6171:FAff port map(x=>p(146)(34),y=>p(147)(34),Cin=>p(148)(34),clock=>clock,reset=>reset,s=>p(226)(34),cout=>p(227)(35));
FA_ff_6172:FAff port map(x=>p(146)(35),y=>p(147)(35),Cin=>p(148)(35),clock=>clock,reset=>reset,s=>p(226)(35),cout=>p(227)(36));
FA_ff_6173:FAff port map(x=>p(146)(36),y=>p(147)(36),Cin=>p(148)(36),clock=>clock,reset=>reset,s=>p(226)(36),cout=>p(227)(37));
FA_ff_6174:FAff port map(x=>p(146)(37),y=>p(147)(37),Cin=>p(148)(37),clock=>clock,reset=>reset,s=>p(226)(37),cout=>p(227)(38));
FA_ff_6175:FAff port map(x=>p(146)(38),y=>p(147)(38),Cin=>p(148)(38),clock=>clock,reset=>reset,s=>p(226)(38),cout=>p(227)(39));
FA_ff_6176:FAff port map(x=>p(146)(39),y=>p(147)(39),Cin=>p(148)(39),clock=>clock,reset=>reset,s=>p(226)(39),cout=>p(227)(40));
FA_ff_6177:FAff port map(x=>p(146)(40),y=>p(147)(40),Cin=>p(148)(40),clock=>clock,reset=>reset,s=>p(226)(40),cout=>p(227)(41));
FA_ff_6178:FAff port map(x=>p(146)(41),y=>p(147)(41),Cin=>p(148)(41),clock=>clock,reset=>reset,s=>p(226)(41),cout=>p(227)(42));
FA_ff_6179:FAff port map(x=>p(146)(42),y=>p(147)(42),Cin=>p(148)(42),clock=>clock,reset=>reset,s=>p(226)(42),cout=>p(227)(43));
FA_ff_6180:FAff port map(x=>p(146)(43),y=>p(147)(43),Cin=>p(148)(43),clock=>clock,reset=>reset,s=>p(226)(43),cout=>p(227)(44));
FA_ff_6181:FAff port map(x=>p(146)(44),y=>p(147)(44),Cin=>p(148)(44),clock=>clock,reset=>reset,s=>p(226)(44),cout=>p(227)(45));
FA_ff_6182:FAff port map(x=>p(146)(45),y=>p(147)(45),Cin=>p(148)(45),clock=>clock,reset=>reset,s=>p(226)(45),cout=>p(227)(46));
FA_ff_6183:FAff port map(x=>p(146)(46),y=>p(147)(46),Cin=>p(148)(46),clock=>clock,reset=>reset,s=>p(226)(46),cout=>p(227)(47));
FA_ff_6184:FAff port map(x=>p(146)(47),y=>p(147)(47),Cin=>p(148)(47),clock=>clock,reset=>reset,s=>p(226)(47),cout=>p(227)(48));
FA_ff_6185:FAff port map(x=>p(146)(48),y=>p(147)(48),Cin=>p(148)(48),clock=>clock,reset=>reset,s=>p(226)(48),cout=>p(227)(49));
FA_ff_6186:FAff port map(x=>p(146)(49),y=>p(147)(49),Cin=>p(148)(49),clock=>clock,reset=>reset,s=>p(226)(49),cout=>p(227)(50));
FA_ff_6187:FAff port map(x=>p(146)(50),y=>p(147)(50),Cin=>p(148)(50),clock=>clock,reset=>reset,s=>p(226)(50),cout=>p(227)(51));
FA_ff_6188:FAff port map(x=>p(146)(51),y=>p(147)(51),Cin=>p(148)(51),clock=>clock,reset=>reset,s=>p(226)(51),cout=>p(227)(52));
FA_ff_6189:FAff port map(x=>p(146)(52),y=>p(147)(52),Cin=>p(148)(52),clock=>clock,reset=>reset,s=>p(226)(52),cout=>p(227)(53));
FA_ff_6190:FAff port map(x=>p(146)(53),y=>p(147)(53),Cin=>p(148)(53),clock=>clock,reset=>reset,s=>p(226)(53),cout=>p(227)(54));
FA_ff_6191:FAff port map(x=>p(146)(54),y=>p(147)(54),Cin=>p(148)(54),clock=>clock,reset=>reset,s=>p(226)(54),cout=>p(227)(55));
FA_ff_6192:FAff port map(x=>p(146)(55),y=>p(147)(55),Cin=>p(148)(55),clock=>clock,reset=>reset,s=>p(226)(55),cout=>p(227)(56));
FA_ff_6193:FAff port map(x=>p(146)(56),y=>p(147)(56),Cin=>p(148)(56),clock=>clock,reset=>reset,s=>p(226)(56),cout=>p(227)(57));
FA_ff_6194:FAff port map(x=>p(146)(57),y=>p(147)(57),Cin=>p(148)(57),clock=>clock,reset=>reset,s=>p(226)(57),cout=>p(227)(58));
FA_ff_6195:FAff port map(x=>p(146)(58),y=>p(147)(58),Cin=>p(148)(58),clock=>clock,reset=>reset,s=>p(226)(58),cout=>p(227)(59));
FA_ff_6196:FAff port map(x=>p(146)(59),y=>p(147)(59),Cin=>p(148)(59),clock=>clock,reset=>reset,s=>p(226)(59),cout=>p(227)(60));
FA_ff_6197:FAff port map(x=>p(146)(60),y=>p(147)(60),Cin=>p(148)(60),clock=>clock,reset=>reset,s=>p(226)(60),cout=>p(227)(61));
FA_ff_6198:FAff port map(x=>p(146)(61),y=>p(147)(61),Cin=>p(148)(61),clock=>clock,reset=>reset,s=>p(226)(61),cout=>p(227)(62));
FA_ff_6199:FAff port map(x=>p(146)(62),y=>p(147)(62),Cin=>p(148)(62),clock=>clock,reset=>reset,s=>p(226)(62),cout=>p(227)(63));
FA_ff_6200:FAff port map(x=>p(146)(63),y=>p(147)(63),Cin=>p(148)(63),clock=>clock,reset=>reset,s=>p(226)(63),cout=>p(227)(64));
FA_ff_6201:FAff port map(x=>p(146)(64),y=>p(147)(64),Cin=>p(148)(64),clock=>clock,reset=>reset,s=>p(226)(64),cout=>p(227)(65));
FA_ff_6202:FAff port map(x=>p(146)(65),y=>p(147)(65),Cin=>p(148)(65),clock=>clock,reset=>reset,s=>p(226)(65),cout=>p(227)(66));
FA_ff_6203:FAff port map(x=>p(146)(66),y=>p(147)(66),Cin=>p(148)(66),clock=>clock,reset=>reset,s=>p(226)(66),cout=>p(227)(67));
FA_ff_6204:FAff port map(x=>p(146)(67),y=>p(147)(67),Cin=>p(148)(67),clock=>clock,reset=>reset,s=>p(226)(67),cout=>p(227)(68));
FA_ff_6205:FAff port map(x=>p(146)(68),y=>p(147)(68),Cin=>p(148)(68),clock=>clock,reset=>reset,s=>p(226)(68),cout=>p(227)(69));
FA_ff_6206:FAff port map(x=>p(146)(69),y=>p(147)(69),Cin=>p(148)(69),clock=>clock,reset=>reset,s=>p(226)(69),cout=>p(227)(70));
FA_ff_6207:FAff port map(x=>p(146)(70),y=>p(147)(70),Cin=>p(148)(70),clock=>clock,reset=>reset,s=>p(226)(70),cout=>p(227)(71));
FA_ff_6208:FAff port map(x=>p(146)(71),y=>p(147)(71),Cin=>p(148)(71),clock=>clock,reset=>reset,s=>p(226)(71),cout=>p(227)(72));
FA_ff_6209:FAff port map(x=>p(146)(72),y=>p(147)(72),Cin=>p(148)(72),clock=>clock,reset=>reset,s=>p(226)(72),cout=>p(227)(73));
FA_ff_6210:FAff port map(x=>p(146)(73),y=>p(147)(73),Cin=>p(148)(73),clock=>clock,reset=>reset,s=>p(226)(73),cout=>p(227)(74));
FA_ff_6211:FAff port map(x=>p(146)(74),y=>p(147)(74),Cin=>p(148)(74),clock=>clock,reset=>reset,s=>p(226)(74),cout=>p(227)(75));
FA_ff_6212:FAff port map(x=>p(146)(75),y=>p(147)(75),Cin=>p(148)(75),clock=>clock,reset=>reset,s=>p(226)(75),cout=>p(227)(76));
FA_ff_6213:FAff port map(x=>p(146)(76),y=>p(147)(76),Cin=>p(148)(76),clock=>clock,reset=>reset,s=>p(226)(76),cout=>p(227)(77));
FA_ff_6214:FAff port map(x=>p(146)(77),y=>p(147)(77),Cin=>p(148)(77),clock=>clock,reset=>reset,s=>p(226)(77),cout=>p(227)(78));
FA_ff_6215:FAff port map(x=>p(146)(78),y=>p(147)(78),Cin=>p(148)(78),clock=>clock,reset=>reset,s=>p(226)(78),cout=>p(227)(79));
FA_ff_6216:FAff port map(x=>p(146)(79),y=>p(147)(79),Cin=>p(148)(79),clock=>clock,reset=>reset,s=>p(226)(79),cout=>p(227)(80));
FA_ff_6217:FAff port map(x=>p(146)(80),y=>p(147)(80),Cin=>p(148)(80),clock=>clock,reset=>reset,s=>p(226)(80),cout=>p(227)(81));
FA_ff_6218:FAff port map(x=>p(146)(81),y=>p(147)(81),Cin=>p(148)(81),clock=>clock,reset=>reset,s=>p(226)(81),cout=>p(227)(82));
FA_ff_6219:FAff port map(x=>p(146)(82),y=>p(147)(82),Cin=>p(148)(82),clock=>clock,reset=>reset,s=>p(226)(82),cout=>p(227)(83));
FA_ff_6220:FAff port map(x=>p(146)(83),y=>p(147)(83),Cin=>p(148)(83),clock=>clock,reset=>reset,s=>p(226)(83),cout=>p(227)(84));
FA_ff_6221:FAff port map(x=>p(146)(84),y=>p(147)(84),Cin=>p(148)(84),clock=>clock,reset=>reset,s=>p(226)(84),cout=>p(227)(85));
FA_ff_6222:FAff port map(x=>p(146)(85),y=>p(147)(85),Cin=>p(148)(85),clock=>clock,reset=>reset,s=>p(226)(85),cout=>p(227)(86));
FA_ff_6223:FAff port map(x=>p(146)(86),y=>p(147)(86),Cin=>p(148)(86),clock=>clock,reset=>reset,s=>p(226)(86),cout=>p(227)(87));
FA_ff_6224:FAff port map(x=>p(146)(87),y=>p(147)(87),Cin=>p(148)(87),clock=>clock,reset=>reset,s=>p(226)(87),cout=>p(227)(88));
FA_ff_6225:FAff port map(x=>p(146)(88),y=>p(147)(88),Cin=>p(148)(88),clock=>clock,reset=>reset,s=>p(226)(88),cout=>p(227)(89));
FA_ff_6226:FAff port map(x=>p(146)(89),y=>p(147)(89),Cin=>p(148)(89),clock=>clock,reset=>reset,s=>p(226)(89),cout=>p(227)(90));
FA_ff_6227:FAff port map(x=>p(146)(90),y=>p(147)(90),Cin=>p(148)(90),clock=>clock,reset=>reset,s=>p(226)(90),cout=>p(227)(91));
FA_ff_6228:FAff port map(x=>p(146)(91),y=>p(147)(91),Cin=>p(148)(91),clock=>clock,reset=>reset,s=>p(226)(91),cout=>p(227)(92));
FA_ff_6229:FAff port map(x=>p(146)(92),y=>p(147)(92),Cin=>p(148)(92),clock=>clock,reset=>reset,s=>p(226)(92),cout=>p(227)(93));
FA_ff_6230:FAff port map(x=>p(146)(93),y=>p(147)(93),Cin=>p(148)(93),clock=>clock,reset=>reset,s=>p(226)(93),cout=>p(227)(94));
FA_ff_6231:FAff port map(x=>p(146)(94),y=>p(147)(94),Cin=>p(148)(94),clock=>clock,reset=>reset,s=>p(226)(94),cout=>p(227)(95));
FA_ff_6232:FAff port map(x=>p(146)(95),y=>p(147)(95),Cin=>p(148)(95),clock=>clock,reset=>reset,s=>p(226)(95),cout=>p(227)(96));
FA_ff_6233:FAff port map(x=>p(146)(96),y=>p(147)(96),Cin=>p(148)(96),clock=>clock,reset=>reset,s=>p(226)(96),cout=>p(227)(97));
FA_ff_6234:FAff port map(x=>p(146)(97),y=>p(147)(97),Cin=>p(148)(97),clock=>clock,reset=>reset,s=>p(226)(97),cout=>p(227)(98));
FA_ff_6235:FAff port map(x=>p(146)(98),y=>p(147)(98),Cin=>p(148)(98),clock=>clock,reset=>reset,s=>p(226)(98),cout=>p(227)(99));
FA_ff_6236:FAff port map(x=>p(146)(99),y=>p(147)(99),Cin=>p(148)(99),clock=>clock,reset=>reset,s=>p(226)(99),cout=>p(227)(100));
FA_ff_6237:FAff port map(x=>p(146)(100),y=>p(147)(100),Cin=>p(148)(100),clock=>clock,reset=>reset,s=>p(226)(100),cout=>p(227)(101));
FA_ff_6238:FAff port map(x=>p(146)(101),y=>p(147)(101),Cin=>p(148)(101),clock=>clock,reset=>reset,s=>p(226)(101),cout=>p(227)(102));
FA_ff_6239:FAff port map(x=>p(146)(102),y=>p(147)(102),Cin=>p(148)(102),clock=>clock,reset=>reset,s=>p(226)(102),cout=>p(227)(103));
FA_ff_6240:FAff port map(x=>p(146)(103),y=>p(147)(103),Cin=>p(148)(103),clock=>clock,reset=>reset,s=>p(226)(103),cout=>p(227)(104));
FA_ff_6241:FAff port map(x=>p(146)(104),y=>p(147)(104),Cin=>p(148)(104),clock=>clock,reset=>reset,s=>p(226)(104),cout=>p(227)(105));
FA_ff_6242:FAff port map(x=>p(146)(105),y=>p(147)(105),Cin=>p(148)(105),clock=>clock,reset=>reset,s=>p(226)(105),cout=>p(227)(106));
FA_ff_6243:FAff port map(x=>p(146)(106),y=>p(147)(106),Cin=>p(148)(106),clock=>clock,reset=>reset,s=>p(226)(106),cout=>p(227)(107));
FA_ff_6244:FAff port map(x=>p(146)(107),y=>p(147)(107),Cin=>p(148)(107),clock=>clock,reset=>reset,s=>p(226)(107),cout=>p(227)(108));
FA_ff_6245:FAff port map(x=>p(146)(108),y=>p(147)(108),Cin=>p(148)(108),clock=>clock,reset=>reset,s=>p(226)(108),cout=>p(227)(109));
FA_ff_6246:FAff port map(x=>p(146)(109),y=>p(147)(109),Cin=>p(148)(109),clock=>clock,reset=>reset,s=>p(226)(109),cout=>p(227)(110));
FA_ff_6247:FAff port map(x=>p(146)(110),y=>p(147)(110),Cin=>p(148)(110),clock=>clock,reset=>reset,s=>p(226)(110),cout=>p(227)(111));
FA_ff_6248:FAff port map(x=>p(146)(111),y=>p(147)(111),Cin=>p(148)(111),clock=>clock,reset=>reset,s=>p(226)(111),cout=>p(227)(112));
FA_ff_6249:FAff port map(x=>p(146)(112),y=>p(147)(112),Cin=>p(148)(112),clock=>clock,reset=>reset,s=>p(226)(112),cout=>p(227)(113));
FA_ff_6250:FAff port map(x=>p(146)(113),y=>p(147)(113),Cin=>p(148)(113),clock=>clock,reset=>reset,s=>p(226)(113),cout=>p(227)(114));
FA_ff_6251:FAff port map(x=>p(146)(114),y=>p(147)(114),Cin=>p(148)(114),clock=>clock,reset=>reset,s=>p(226)(114),cout=>p(227)(115));
FA_ff_6252:FAff port map(x=>p(146)(115),y=>p(147)(115),Cin=>p(148)(115),clock=>clock,reset=>reset,s=>p(226)(115),cout=>p(227)(116));
FA_ff_6253:FAff port map(x=>p(146)(116),y=>p(147)(116),Cin=>p(148)(116),clock=>clock,reset=>reset,s=>p(226)(116),cout=>p(227)(117));
FA_ff_6254:FAff port map(x=>p(146)(117),y=>p(147)(117),Cin=>p(148)(117),clock=>clock,reset=>reset,s=>p(226)(117),cout=>p(227)(118));
FA_ff_6255:FAff port map(x=>p(146)(118),y=>p(147)(118),Cin=>p(148)(118),clock=>clock,reset=>reset,s=>p(226)(118),cout=>p(227)(119));
FA_ff_6256:FAff port map(x=>p(146)(119),y=>p(147)(119),Cin=>p(148)(119),clock=>clock,reset=>reset,s=>p(226)(119),cout=>p(227)(120));
FA_ff_6257:FAff port map(x=>p(146)(120),y=>p(147)(120),Cin=>p(148)(120),clock=>clock,reset=>reset,s=>p(226)(120),cout=>p(227)(121));
FA_ff_6258:FAff port map(x=>p(146)(121),y=>p(147)(121),Cin=>p(148)(121),clock=>clock,reset=>reset,s=>p(226)(121),cout=>p(227)(122));
FA_ff_6259:FAff port map(x=>p(146)(122),y=>p(147)(122),Cin=>p(148)(122),clock=>clock,reset=>reset,s=>p(226)(122),cout=>p(227)(123));
FA_ff_6260:FAff port map(x=>p(146)(123),y=>p(147)(123),Cin=>p(148)(123),clock=>clock,reset=>reset,s=>p(226)(123),cout=>p(227)(124));
FA_ff_6261:FAff port map(x=>p(146)(124),y=>p(147)(124),Cin=>p(148)(124),clock=>clock,reset=>reset,s=>p(226)(124),cout=>p(227)(125));
FA_ff_6262:FAff port map(x=>p(146)(125),y=>p(147)(125),Cin=>p(148)(125),clock=>clock,reset=>reset,s=>p(226)(125),cout=>p(227)(126));
FA_ff_6263:FAff port map(x=>p(146)(126),y=>p(147)(126),Cin=>p(148)(126),clock=>clock,reset=>reset,s=>p(226)(126),cout=>p(227)(127));
FA_ff_6264:FAff port map(x=>p(146)(127),y=>p(147)(127),Cin=>p(148)(127),clock=>clock,reset=>reset,s=>p(226)(127),cout=>p(227)(128));
p(226)(128)<=p(147)(128);
p(228)(0)<=p(150)(0);
FA_ff_6265:FAff port map(x=>p(149)(1),y=>p(150)(1),Cin=>p(151)(1),clock=>clock,reset=>reset,s=>p(228)(1),cout=>p(229)(2));
FA_ff_6266:FAff port map(x=>p(149)(2),y=>p(150)(2),Cin=>p(151)(2),clock=>clock,reset=>reset,s=>p(228)(2),cout=>p(229)(3));
FA_ff_6267:FAff port map(x=>p(149)(3),y=>p(150)(3),Cin=>p(151)(3),clock=>clock,reset=>reset,s=>p(228)(3),cout=>p(229)(4));
FA_ff_6268:FAff port map(x=>p(149)(4),y=>p(150)(4),Cin=>p(151)(4),clock=>clock,reset=>reset,s=>p(228)(4),cout=>p(229)(5));
FA_ff_6269:FAff port map(x=>p(149)(5),y=>p(150)(5),Cin=>p(151)(5),clock=>clock,reset=>reset,s=>p(228)(5),cout=>p(229)(6));
FA_ff_6270:FAff port map(x=>p(149)(6),y=>p(150)(6),Cin=>p(151)(6),clock=>clock,reset=>reset,s=>p(228)(6),cout=>p(229)(7));
FA_ff_6271:FAff port map(x=>p(149)(7),y=>p(150)(7),Cin=>p(151)(7),clock=>clock,reset=>reset,s=>p(228)(7),cout=>p(229)(8));
FA_ff_6272:FAff port map(x=>p(149)(8),y=>p(150)(8),Cin=>p(151)(8),clock=>clock,reset=>reset,s=>p(228)(8),cout=>p(229)(9));
FA_ff_6273:FAff port map(x=>p(149)(9),y=>p(150)(9),Cin=>p(151)(9),clock=>clock,reset=>reset,s=>p(228)(9),cout=>p(229)(10));
FA_ff_6274:FAff port map(x=>p(149)(10),y=>p(150)(10),Cin=>p(151)(10),clock=>clock,reset=>reset,s=>p(228)(10),cout=>p(229)(11));
FA_ff_6275:FAff port map(x=>p(149)(11),y=>p(150)(11),Cin=>p(151)(11),clock=>clock,reset=>reset,s=>p(228)(11),cout=>p(229)(12));
FA_ff_6276:FAff port map(x=>p(149)(12),y=>p(150)(12),Cin=>p(151)(12),clock=>clock,reset=>reset,s=>p(228)(12),cout=>p(229)(13));
FA_ff_6277:FAff port map(x=>p(149)(13),y=>p(150)(13),Cin=>p(151)(13),clock=>clock,reset=>reset,s=>p(228)(13),cout=>p(229)(14));
FA_ff_6278:FAff port map(x=>p(149)(14),y=>p(150)(14),Cin=>p(151)(14),clock=>clock,reset=>reset,s=>p(228)(14),cout=>p(229)(15));
FA_ff_6279:FAff port map(x=>p(149)(15),y=>p(150)(15),Cin=>p(151)(15),clock=>clock,reset=>reset,s=>p(228)(15),cout=>p(229)(16));
FA_ff_6280:FAff port map(x=>p(149)(16),y=>p(150)(16),Cin=>p(151)(16),clock=>clock,reset=>reset,s=>p(228)(16),cout=>p(229)(17));
FA_ff_6281:FAff port map(x=>p(149)(17),y=>p(150)(17),Cin=>p(151)(17),clock=>clock,reset=>reset,s=>p(228)(17),cout=>p(229)(18));
FA_ff_6282:FAff port map(x=>p(149)(18),y=>p(150)(18),Cin=>p(151)(18),clock=>clock,reset=>reset,s=>p(228)(18),cout=>p(229)(19));
FA_ff_6283:FAff port map(x=>p(149)(19),y=>p(150)(19),Cin=>p(151)(19),clock=>clock,reset=>reset,s=>p(228)(19),cout=>p(229)(20));
FA_ff_6284:FAff port map(x=>p(149)(20),y=>p(150)(20),Cin=>p(151)(20),clock=>clock,reset=>reset,s=>p(228)(20),cout=>p(229)(21));
FA_ff_6285:FAff port map(x=>p(149)(21),y=>p(150)(21),Cin=>p(151)(21),clock=>clock,reset=>reset,s=>p(228)(21),cout=>p(229)(22));
FA_ff_6286:FAff port map(x=>p(149)(22),y=>p(150)(22),Cin=>p(151)(22),clock=>clock,reset=>reset,s=>p(228)(22),cout=>p(229)(23));
FA_ff_6287:FAff port map(x=>p(149)(23),y=>p(150)(23),Cin=>p(151)(23),clock=>clock,reset=>reset,s=>p(228)(23),cout=>p(229)(24));
FA_ff_6288:FAff port map(x=>p(149)(24),y=>p(150)(24),Cin=>p(151)(24),clock=>clock,reset=>reset,s=>p(228)(24),cout=>p(229)(25));
FA_ff_6289:FAff port map(x=>p(149)(25),y=>p(150)(25),Cin=>p(151)(25),clock=>clock,reset=>reset,s=>p(228)(25),cout=>p(229)(26));
FA_ff_6290:FAff port map(x=>p(149)(26),y=>p(150)(26),Cin=>p(151)(26),clock=>clock,reset=>reset,s=>p(228)(26),cout=>p(229)(27));
FA_ff_6291:FAff port map(x=>p(149)(27),y=>p(150)(27),Cin=>p(151)(27),clock=>clock,reset=>reset,s=>p(228)(27),cout=>p(229)(28));
FA_ff_6292:FAff port map(x=>p(149)(28),y=>p(150)(28),Cin=>p(151)(28),clock=>clock,reset=>reset,s=>p(228)(28),cout=>p(229)(29));
FA_ff_6293:FAff port map(x=>p(149)(29),y=>p(150)(29),Cin=>p(151)(29),clock=>clock,reset=>reset,s=>p(228)(29),cout=>p(229)(30));
FA_ff_6294:FAff port map(x=>p(149)(30),y=>p(150)(30),Cin=>p(151)(30),clock=>clock,reset=>reset,s=>p(228)(30),cout=>p(229)(31));
FA_ff_6295:FAff port map(x=>p(149)(31),y=>p(150)(31),Cin=>p(151)(31),clock=>clock,reset=>reset,s=>p(228)(31),cout=>p(229)(32));
FA_ff_6296:FAff port map(x=>p(149)(32),y=>p(150)(32),Cin=>p(151)(32),clock=>clock,reset=>reset,s=>p(228)(32),cout=>p(229)(33));
FA_ff_6297:FAff port map(x=>p(149)(33),y=>p(150)(33),Cin=>p(151)(33),clock=>clock,reset=>reset,s=>p(228)(33),cout=>p(229)(34));
FA_ff_6298:FAff port map(x=>p(149)(34),y=>p(150)(34),Cin=>p(151)(34),clock=>clock,reset=>reset,s=>p(228)(34),cout=>p(229)(35));
FA_ff_6299:FAff port map(x=>p(149)(35),y=>p(150)(35),Cin=>p(151)(35),clock=>clock,reset=>reset,s=>p(228)(35),cout=>p(229)(36));
FA_ff_6300:FAff port map(x=>p(149)(36),y=>p(150)(36),Cin=>p(151)(36),clock=>clock,reset=>reset,s=>p(228)(36),cout=>p(229)(37));
FA_ff_6301:FAff port map(x=>p(149)(37),y=>p(150)(37),Cin=>p(151)(37),clock=>clock,reset=>reset,s=>p(228)(37),cout=>p(229)(38));
FA_ff_6302:FAff port map(x=>p(149)(38),y=>p(150)(38),Cin=>p(151)(38),clock=>clock,reset=>reset,s=>p(228)(38),cout=>p(229)(39));
FA_ff_6303:FAff port map(x=>p(149)(39),y=>p(150)(39),Cin=>p(151)(39),clock=>clock,reset=>reset,s=>p(228)(39),cout=>p(229)(40));
FA_ff_6304:FAff port map(x=>p(149)(40),y=>p(150)(40),Cin=>p(151)(40),clock=>clock,reset=>reset,s=>p(228)(40),cout=>p(229)(41));
FA_ff_6305:FAff port map(x=>p(149)(41),y=>p(150)(41),Cin=>p(151)(41),clock=>clock,reset=>reset,s=>p(228)(41),cout=>p(229)(42));
FA_ff_6306:FAff port map(x=>p(149)(42),y=>p(150)(42),Cin=>p(151)(42),clock=>clock,reset=>reset,s=>p(228)(42),cout=>p(229)(43));
FA_ff_6307:FAff port map(x=>p(149)(43),y=>p(150)(43),Cin=>p(151)(43),clock=>clock,reset=>reset,s=>p(228)(43),cout=>p(229)(44));
FA_ff_6308:FAff port map(x=>p(149)(44),y=>p(150)(44),Cin=>p(151)(44),clock=>clock,reset=>reset,s=>p(228)(44),cout=>p(229)(45));
FA_ff_6309:FAff port map(x=>p(149)(45),y=>p(150)(45),Cin=>p(151)(45),clock=>clock,reset=>reset,s=>p(228)(45),cout=>p(229)(46));
FA_ff_6310:FAff port map(x=>p(149)(46),y=>p(150)(46),Cin=>p(151)(46),clock=>clock,reset=>reset,s=>p(228)(46),cout=>p(229)(47));
FA_ff_6311:FAff port map(x=>p(149)(47),y=>p(150)(47),Cin=>p(151)(47),clock=>clock,reset=>reset,s=>p(228)(47),cout=>p(229)(48));
FA_ff_6312:FAff port map(x=>p(149)(48),y=>p(150)(48),Cin=>p(151)(48),clock=>clock,reset=>reset,s=>p(228)(48),cout=>p(229)(49));
FA_ff_6313:FAff port map(x=>p(149)(49),y=>p(150)(49),Cin=>p(151)(49),clock=>clock,reset=>reset,s=>p(228)(49),cout=>p(229)(50));
FA_ff_6314:FAff port map(x=>p(149)(50),y=>p(150)(50),Cin=>p(151)(50),clock=>clock,reset=>reset,s=>p(228)(50),cout=>p(229)(51));
FA_ff_6315:FAff port map(x=>p(149)(51),y=>p(150)(51),Cin=>p(151)(51),clock=>clock,reset=>reset,s=>p(228)(51),cout=>p(229)(52));
FA_ff_6316:FAff port map(x=>p(149)(52),y=>p(150)(52),Cin=>p(151)(52),clock=>clock,reset=>reset,s=>p(228)(52),cout=>p(229)(53));
FA_ff_6317:FAff port map(x=>p(149)(53),y=>p(150)(53),Cin=>p(151)(53),clock=>clock,reset=>reset,s=>p(228)(53),cout=>p(229)(54));
FA_ff_6318:FAff port map(x=>p(149)(54),y=>p(150)(54),Cin=>p(151)(54),clock=>clock,reset=>reset,s=>p(228)(54),cout=>p(229)(55));
FA_ff_6319:FAff port map(x=>p(149)(55),y=>p(150)(55),Cin=>p(151)(55),clock=>clock,reset=>reset,s=>p(228)(55),cout=>p(229)(56));
FA_ff_6320:FAff port map(x=>p(149)(56),y=>p(150)(56),Cin=>p(151)(56),clock=>clock,reset=>reset,s=>p(228)(56),cout=>p(229)(57));
FA_ff_6321:FAff port map(x=>p(149)(57),y=>p(150)(57),Cin=>p(151)(57),clock=>clock,reset=>reset,s=>p(228)(57),cout=>p(229)(58));
FA_ff_6322:FAff port map(x=>p(149)(58),y=>p(150)(58),Cin=>p(151)(58),clock=>clock,reset=>reset,s=>p(228)(58),cout=>p(229)(59));
FA_ff_6323:FAff port map(x=>p(149)(59),y=>p(150)(59),Cin=>p(151)(59),clock=>clock,reset=>reset,s=>p(228)(59),cout=>p(229)(60));
FA_ff_6324:FAff port map(x=>p(149)(60),y=>p(150)(60),Cin=>p(151)(60),clock=>clock,reset=>reset,s=>p(228)(60),cout=>p(229)(61));
FA_ff_6325:FAff port map(x=>p(149)(61),y=>p(150)(61),Cin=>p(151)(61),clock=>clock,reset=>reset,s=>p(228)(61),cout=>p(229)(62));
FA_ff_6326:FAff port map(x=>p(149)(62),y=>p(150)(62),Cin=>p(151)(62),clock=>clock,reset=>reset,s=>p(228)(62),cout=>p(229)(63));
FA_ff_6327:FAff port map(x=>p(149)(63),y=>p(150)(63),Cin=>p(151)(63),clock=>clock,reset=>reset,s=>p(228)(63),cout=>p(229)(64));
FA_ff_6328:FAff port map(x=>p(149)(64),y=>p(150)(64),Cin=>p(151)(64),clock=>clock,reset=>reset,s=>p(228)(64),cout=>p(229)(65));
FA_ff_6329:FAff port map(x=>p(149)(65),y=>p(150)(65),Cin=>p(151)(65),clock=>clock,reset=>reset,s=>p(228)(65),cout=>p(229)(66));
FA_ff_6330:FAff port map(x=>p(149)(66),y=>p(150)(66),Cin=>p(151)(66),clock=>clock,reset=>reset,s=>p(228)(66),cout=>p(229)(67));
FA_ff_6331:FAff port map(x=>p(149)(67),y=>p(150)(67),Cin=>p(151)(67),clock=>clock,reset=>reset,s=>p(228)(67),cout=>p(229)(68));
FA_ff_6332:FAff port map(x=>p(149)(68),y=>p(150)(68),Cin=>p(151)(68),clock=>clock,reset=>reset,s=>p(228)(68),cout=>p(229)(69));
FA_ff_6333:FAff port map(x=>p(149)(69),y=>p(150)(69),Cin=>p(151)(69),clock=>clock,reset=>reset,s=>p(228)(69),cout=>p(229)(70));
FA_ff_6334:FAff port map(x=>p(149)(70),y=>p(150)(70),Cin=>p(151)(70),clock=>clock,reset=>reset,s=>p(228)(70),cout=>p(229)(71));
FA_ff_6335:FAff port map(x=>p(149)(71),y=>p(150)(71),Cin=>p(151)(71),clock=>clock,reset=>reset,s=>p(228)(71),cout=>p(229)(72));
FA_ff_6336:FAff port map(x=>p(149)(72),y=>p(150)(72),Cin=>p(151)(72),clock=>clock,reset=>reset,s=>p(228)(72),cout=>p(229)(73));
FA_ff_6337:FAff port map(x=>p(149)(73),y=>p(150)(73),Cin=>p(151)(73),clock=>clock,reset=>reset,s=>p(228)(73),cout=>p(229)(74));
FA_ff_6338:FAff port map(x=>p(149)(74),y=>p(150)(74),Cin=>p(151)(74),clock=>clock,reset=>reset,s=>p(228)(74),cout=>p(229)(75));
FA_ff_6339:FAff port map(x=>p(149)(75),y=>p(150)(75),Cin=>p(151)(75),clock=>clock,reset=>reset,s=>p(228)(75),cout=>p(229)(76));
FA_ff_6340:FAff port map(x=>p(149)(76),y=>p(150)(76),Cin=>p(151)(76),clock=>clock,reset=>reset,s=>p(228)(76),cout=>p(229)(77));
FA_ff_6341:FAff port map(x=>p(149)(77),y=>p(150)(77),Cin=>p(151)(77),clock=>clock,reset=>reset,s=>p(228)(77),cout=>p(229)(78));
FA_ff_6342:FAff port map(x=>p(149)(78),y=>p(150)(78),Cin=>p(151)(78),clock=>clock,reset=>reset,s=>p(228)(78),cout=>p(229)(79));
FA_ff_6343:FAff port map(x=>p(149)(79),y=>p(150)(79),Cin=>p(151)(79),clock=>clock,reset=>reset,s=>p(228)(79),cout=>p(229)(80));
FA_ff_6344:FAff port map(x=>p(149)(80),y=>p(150)(80),Cin=>p(151)(80),clock=>clock,reset=>reset,s=>p(228)(80),cout=>p(229)(81));
FA_ff_6345:FAff port map(x=>p(149)(81),y=>p(150)(81),Cin=>p(151)(81),clock=>clock,reset=>reset,s=>p(228)(81),cout=>p(229)(82));
FA_ff_6346:FAff port map(x=>p(149)(82),y=>p(150)(82),Cin=>p(151)(82),clock=>clock,reset=>reset,s=>p(228)(82),cout=>p(229)(83));
FA_ff_6347:FAff port map(x=>p(149)(83),y=>p(150)(83),Cin=>p(151)(83),clock=>clock,reset=>reset,s=>p(228)(83),cout=>p(229)(84));
FA_ff_6348:FAff port map(x=>p(149)(84),y=>p(150)(84),Cin=>p(151)(84),clock=>clock,reset=>reset,s=>p(228)(84),cout=>p(229)(85));
FA_ff_6349:FAff port map(x=>p(149)(85),y=>p(150)(85),Cin=>p(151)(85),clock=>clock,reset=>reset,s=>p(228)(85),cout=>p(229)(86));
FA_ff_6350:FAff port map(x=>p(149)(86),y=>p(150)(86),Cin=>p(151)(86),clock=>clock,reset=>reset,s=>p(228)(86),cout=>p(229)(87));
FA_ff_6351:FAff port map(x=>p(149)(87),y=>p(150)(87),Cin=>p(151)(87),clock=>clock,reset=>reset,s=>p(228)(87),cout=>p(229)(88));
FA_ff_6352:FAff port map(x=>p(149)(88),y=>p(150)(88),Cin=>p(151)(88),clock=>clock,reset=>reset,s=>p(228)(88),cout=>p(229)(89));
FA_ff_6353:FAff port map(x=>p(149)(89),y=>p(150)(89),Cin=>p(151)(89),clock=>clock,reset=>reset,s=>p(228)(89),cout=>p(229)(90));
FA_ff_6354:FAff port map(x=>p(149)(90),y=>p(150)(90),Cin=>p(151)(90),clock=>clock,reset=>reset,s=>p(228)(90),cout=>p(229)(91));
FA_ff_6355:FAff port map(x=>p(149)(91),y=>p(150)(91),Cin=>p(151)(91),clock=>clock,reset=>reset,s=>p(228)(91),cout=>p(229)(92));
FA_ff_6356:FAff port map(x=>p(149)(92),y=>p(150)(92),Cin=>p(151)(92),clock=>clock,reset=>reset,s=>p(228)(92),cout=>p(229)(93));
FA_ff_6357:FAff port map(x=>p(149)(93),y=>p(150)(93),Cin=>p(151)(93),clock=>clock,reset=>reset,s=>p(228)(93),cout=>p(229)(94));
FA_ff_6358:FAff port map(x=>p(149)(94),y=>p(150)(94),Cin=>p(151)(94),clock=>clock,reset=>reset,s=>p(228)(94),cout=>p(229)(95));
FA_ff_6359:FAff port map(x=>p(149)(95),y=>p(150)(95),Cin=>p(151)(95),clock=>clock,reset=>reset,s=>p(228)(95),cout=>p(229)(96));
FA_ff_6360:FAff port map(x=>p(149)(96),y=>p(150)(96),Cin=>p(151)(96),clock=>clock,reset=>reset,s=>p(228)(96),cout=>p(229)(97));
FA_ff_6361:FAff port map(x=>p(149)(97),y=>p(150)(97),Cin=>p(151)(97),clock=>clock,reset=>reset,s=>p(228)(97),cout=>p(229)(98));
FA_ff_6362:FAff port map(x=>p(149)(98),y=>p(150)(98),Cin=>p(151)(98),clock=>clock,reset=>reset,s=>p(228)(98),cout=>p(229)(99));
FA_ff_6363:FAff port map(x=>p(149)(99),y=>p(150)(99),Cin=>p(151)(99),clock=>clock,reset=>reset,s=>p(228)(99),cout=>p(229)(100));
FA_ff_6364:FAff port map(x=>p(149)(100),y=>p(150)(100),Cin=>p(151)(100),clock=>clock,reset=>reset,s=>p(228)(100),cout=>p(229)(101));
FA_ff_6365:FAff port map(x=>p(149)(101),y=>p(150)(101),Cin=>p(151)(101),clock=>clock,reset=>reset,s=>p(228)(101),cout=>p(229)(102));
FA_ff_6366:FAff port map(x=>p(149)(102),y=>p(150)(102),Cin=>p(151)(102),clock=>clock,reset=>reset,s=>p(228)(102),cout=>p(229)(103));
FA_ff_6367:FAff port map(x=>p(149)(103),y=>p(150)(103),Cin=>p(151)(103),clock=>clock,reset=>reset,s=>p(228)(103),cout=>p(229)(104));
FA_ff_6368:FAff port map(x=>p(149)(104),y=>p(150)(104),Cin=>p(151)(104),clock=>clock,reset=>reset,s=>p(228)(104),cout=>p(229)(105));
FA_ff_6369:FAff port map(x=>p(149)(105),y=>p(150)(105),Cin=>p(151)(105),clock=>clock,reset=>reset,s=>p(228)(105),cout=>p(229)(106));
FA_ff_6370:FAff port map(x=>p(149)(106),y=>p(150)(106),Cin=>p(151)(106),clock=>clock,reset=>reset,s=>p(228)(106),cout=>p(229)(107));
FA_ff_6371:FAff port map(x=>p(149)(107),y=>p(150)(107),Cin=>p(151)(107),clock=>clock,reset=>reset,s=>p(228)(107),cout=>p(229)(108));
FA_ff_6372:FAff port map(x=>p(149)(108),y=>p(150)(108),Cin=>p(151)(108),clock=>clock,reset=>reset,s=>p(228)(108),cout=>p(229)(109));
FA_ff_6373:FAff port map(x=>p(149)(109),y=>p(150)(109),Cin=>p(151)(109),clock=>clock,reset=>reset,s=>p(228)(109),cout=>p(229)(110));
FA_ff_6374:FAff port map(x=>p(149)(110),y=>p(150)(110),Cin=>p(151)(110),clock=>clock,reset=>reset,s=>p(228)(110),cout=>p(229)(111));
FA_ff_6375:FAff port map(x=>p(149)(111),y=>p(150)(111),Cin=>p(151)(111),clock=>clock,reset=>reset,s=>p(228)(111),cout=>p(229)(112));
FA_ff_6376:FAff port map(x=>p(149)(112),y=>p(150)(112),Cin=>p(151)(112),clock=>clock,reset=>reset,s=>p(228)(112),cout=>p(229)(113));
FA_ff_6377:FAff port map(x=>p(149)(113),y=>p(150)(113),Cin=>p(151)(113),clock=>clock,reset=>reset,s=>p(228)(113),cout=>p(229)(114));
FA_ff_6378:FAff port map(x=>p(149)(114),y=>p(150)(114),Cin=>p(151)(114),clock=>clock,reset=>reset,s=>p(228)(114),cout=>p(229)(115));
FA_ff_6379:FAff port map(x=>p(149)(115),y=>p(150)(115),Cin=>p(151)(115),clock=>clock,reset=>reset,s=>p(228)(115),cout=>p(229)(116));
FA_ff_6380:FAff port map(x=>p(149)(116),y=>p(150)(116),Cin=>p(151)(116),clock=>clock,reset=>reset,s=>p(228)(116),cout=>p(229)(117));
FA_ff_6381:FAff port map(x=>p(149)(117),y=>p(150)(117),Cin=>p(151)(117),clock=>clock,reset=>reset,s=>p(228)(117),cout=>p(229)(118));
FA_ff_6382:FAff port map(x=>p(149)(118),y=>p(150)(118),Cin=>p(151)(118),clock=>clock,reset=>reset,s=>p(228)(118),cout=>p(229)(119));
FA_ff_6383:FAff port map(x=>p(149)(119),y=>p(150)(119),Cin=>p(151)(119),clock=>clock,reset=>reset,s=>p(228)(119),cout=>p(229)(120));
FA_ff_6384:FAff port map(x=>p(149)(120),y=>p(150)(120),Cin=>p(151)(120),clock=>clock,reset=>reset,s=>p(228)(120),cout=>p(229)(121));
FA_ff_6385:FAff port map(x=>p(149)(121),y=>p(150)(121),Cin=>p(151)(121),clock=>clock,reset=>reset,s=>p(228)(121),cout=>p(229)(122));
FA_ff_6386:FAff port map(x=>p(149)(122),y=>p(150)(122),Cin=>p(151)(122),clock=>clock,reset=>reset,s=>p(228)(122),cout=>p(229)(123));
FA_ff_6387:FAff port map(x=>p(149)(123),y=>p(150)(123),Cin=>p(151)(123),clock=>clock,reset=>reset,s=>p(228)(123),cout=>p(229)(124));
FA_ff_6388:FAff port map(x=>p(149)(124),y=>p(150)(124),Cin=>p(151)(124),clock=>clock,reset=>reset,s=>p(228)(124),cout=>p(229)(125));
FA_ff_6389:FAff port map(x=>p(149)(125),y=>p(150)(125),Cin=>p(151)(125),clock=>clock,reset=>reset,s=>p(228)(125),cout=>p(229)(126));
FA_ff_6390:FAff port map(x=>p(149)(126),y=>p(150)(126),Cin=>p(151)(126),clock=>clock,reset=>reset,s=>p(228)(126),cout=>p(229)(127));
FA_ff_6391:FAff port map(x=>p(149)(127),y=>p(150)(127),Cin=>p(151)(127),clock=>clock,reset=>reset,s=>p(228)(127),cout=>p(229)(128));
HA_ff_7:HAff port map(x=>p(149)(128),y=>p(151)(128),clock=>clock,reset=>reset,s=>p(228)(128),c=>p(229)(129));
HA_ff_8:HAff port map(x=>p(152)(0),y=>p(154)(0),clock=>clock,reset=>reset,s=>p(230)(0),c=>p(231)(1));
FA_ff_6392:FAff port map(x=>p(152)(1),y=>p(153)(1),Cin=>p(154)(1),clock=>clock,reset=>reset,s=>p(230)(1),cout=>p(231)(2));
FA_ff_6393:FAff port map(x=>p(152)(2),y=>p(153)(2),Cin=>p(154)(2),clock=>clock,reset=>reset,s=>p(230)(2),cout=>p(231)(3));
FA_ff_6394:FAff port map(x=>p(152)(3),y=>p(153)(3),Cin=>p(154)(3),clock=>clock,reset=>reset,s=>p(230)(3),cout=>p(231)(4));
FA_ff_6395:FAff port map(x=>p(152)(4),y=>p(153)(4),Cin=>p(154)(4),clock=>clock,reset=>reset,s=>p(230)(4),cout=>p(231)(5));
FA_ff_6396:FAff port map(x=>p(152)(5),y=>p(153)(5),Cin=>p(154)(5),clock=>clock,reset=>reset,s=>p(230)(5),cout=>p(231)(6));
FA_ff_6397:FAff port map(x=>p(152)(6),y=>p(153)(6),Cin=>p(154)(6),clock=>clock,reset=>reset,s=>p(230)(6),cout=>p(231)(7));
FA_ff_6398:FAff port map(x=>p(152)(7),y=>p(153)(7),Cin=>p(154)(7),clock=>clock,reset=>reset,s=>p(230)(7),cout=>p(231)(8));
FA_ff_6399:FAff port map(x=>p(152)(8),y=>p(153)(8),Cin=>p(154)(8),clock=>clock,reset=>reset,s=>p(230)(8),cout=>p(231)(9));
FA_ff_6400:FAff port map(x=>p(152)(9),y=>p(153)(9),Cin=>p(154)(9),clock=>clock,reset=>reset,s=>p(230)(9),cout=>p(231)(10));
FA_ff_6401:FAff port map(x=>p(152)(10),y=>p(153)(10),Cin=>p(154)(10),clock=>clock,reset=>reset,s=>p(230)(10),cout=>p(231)(11));
FA_ff_6402:FAff port map(x=>p(152)(11),y=>p(153)(11),Cin=>p(154)(11),clock=>clock,reset=>reset,s=>p(230)(11),cout=>p(231)(12));
FA_ff_6403:FAff port map(x=>p(152)(12),y=>p(153)(12),Cin=>p(154)(12),clock=>clock,reset=>reset,s=>p(230)(12),cout=>p(231)(13));
FA_ff_6404:FAff port map(x=>p(152)(13),y=>p(153)(13),Cin=>p(154)(13),clock=>clock,reset=>reset,s=>p(230)(13),cout=>p(231)(14));
FA_ff_6405:FAff port map(x=>p(152)(14),y=>p(153)(14),Cin=>p(154)(14),clock=>clock,reset=>reset,s=>p(230)(14),cout=>p(231)(15));
FA_ff_6406:FAff port map(x=>p(152)(15),y=>p(153)(15),Cin=>p(154)(15),clock=>clock,reset=>reset,s=>p(230)(15),cout=>p(231)(16));
FA_ff_6407:FAff port map(x=>p(152)(16),y=>p(153)(16),Cin=>p(154)(16),clock=>clock,reset=>reset,s=>p(230)(16),cout=>p(231)(17));
FA_ff_6408:FAff port map(x=>p(152)(17),y=>p(153)(17),Cin=>p(154)(17),clock=>clock,reset=>reset,s=>p(230)(17),cout=>p(231)(18));
FA_ff_6409:FAff port map(x=>p(152)(18),y=>p(153)(18),Cin=>p(154)(18),clock=>clock,reset=>reset,s=>p(230)(18),cout=>p(231)(19));
FA_ff_6410:FAff port map(x=>p(152)(19),y=>p(153)(19),Cin=>p(154)(19),clock=>clock,reset=>reset,s=>p(230)(19),cout=>p(231)(20));
FA_ff_6411:FAff port map(x=>p(152)(20),y=>p(153)(20),Cin=>p(154)(20),clock=>clock,reset=>reset,s=>p(230)(20),cout=>p(231)(21));
FA_ff_6412:FAff port map(x=>p(152)(21),y=>p(153)(21),Cin=>p(154)(21),clock=>clock,reset=>reset,s=>p(230)(21),cout=>p(231)(22));
FA_ff_6413:FAff port map(x=>p(152)(22),y=>p(153)(22),Cin=>p(154)(22),clock=>clock,reset=>reset,s=>p(230)(22),cout=>p(231)(23));
FA_ff_6414:FAff port map(x=>p(152)(23),y=>p(153)(23),Cin=>p(154)(23),clock=>clock,reset=>reset,s=>p(230)(23),cout=>p(231)(24));
FA_ff_6415:FAff port map(x=>p(152)(24),y=>p(153)(24),Cin=>p(154)(24),clock=>clock,reset=>reset,s=>p(230)(24),cout=>p(231)(25));
FA_ff_6416:FAff port map(x=>p(152)(25),y=>p(153)(25),Cin=>p(154)(25),clock=>clock,reset=>reset,s=>p(230)(25),cout=>p(231)(26));
FA_ff_6417:FAff port map(x=>p(152)(26),y=>p(153)(26),Cin=>p(154)(26),clock=>clock,reset=>reset,s=>p(230)(26),cout=>p(231)(27));
FA_ff_6418:FAff port map(x=>p(152)(27),y=>p(153)(27),Cin=>p(154)(27),clock=>clock,reset=>reset,s=>p(230)(27),cout=>p(231)(28));
FA_ff_6419:FAff port map(x=>p(152)(28),y=>p(153)(28),Cin=>p(154)(28),clock=>clock,reset=>reset,s=>p(230)(28),cout=>p(231)(29));
FA_ff_6420:FAff port map(x=>p(152)(29),y=>p(153)(29),Cin=>p(154)(29),clock=>clock,reset=>reset,s=>p(230)(29),cout=>p(231)(30));
FA_ff_6421:FAff port map(x=>p(152)(30),y=>p(153)(30),Cin=>p(154)(30),clock=>clock,reset=>reset,s=>p(230)(30),cout=>p(231)(31));
FA_ff_6422:FAff port map(x=>p(152)(31),y=>p(153)(31),Cin=>p(154)(31),clock=>clock,reset=>reset,s=>p(230)(31),cout=>p(231)(32));
FA_ff_6423:FAff port map(x=>p(152)(32),y=>p(153)(32),Cin=>p(154)(32),clock=>clock,reset=>reset,s=>p(230)(32),cout=>p(231)(33));
FA_ff_6424:FAff port map(x=>p(152)(33),y=>p(153)(33),Cin=>p(154)(33),clock=>clock,reset=>reset,s=>p(230)(33),cout=>p(231)(34));
FA_ff_6425:FAff port map(x=>p(152)(34),y=>p(153)(34),Cin=>p(154)(34),clock=>clock,reset=>reset,s=>p(230)(34),cout=>p(231)(35));
FA_ff_6426:FAff port map(x=>p(152)(35),y=>p(153)(35),Cin=>p(154)(35),clock=>clock,reset=>reset,s=>p(230)(35),cout=>p(231)(36));
FA_ff_6427:FAff port map(x=>p(152)(36),y=>p(153)(36),Cin=>p(154)(36),clock=>clock,reset=>reset,s=>p(230)(36),cout=>p(231)(37));
FA_ff_6428:FAff port map(x=>p(152)(37),y=>p(153)(37),Cin=>p(154)(37),clock=>clock,reset=>reset,s=>p(230)(37),cout=>p(231)(38));
FA_ff_6429:FAff port map(x=>p(152)(38),y=>p(153)(38),Cin=>p(154)(38),clock=>clock,reset=>reset,s=>p(230)(38),cout=>p(231)(39));
FA_ff_6430:FAff port map(x=>p(152)(39),y=>p(153)(39),Cin=>p(154)(39),clock=>clock,reset=>reset,s=>p(230)(39),cout=>p(231)(40));
FA_ff_6431:FAff port map(x=>p(152)(40),y=>p(153)(40),Cin=>p(154)(40),clock=>clock,reset=>reset,s=>p(230)(40),cout=>p(231)(41));
FA_ff_6432:FAff port map(x=>p(152)(41),y=>p(153)(41),Cin=>p(154)(41),clock=>clock,reset=>reset,s=>p(230)(41),cout=>p(231)(42));
FA_ff_6433:FAff port map(x=>p(152)(42),y=>p(153)(42),Cin=>p(154)(42),clock=>clock,reset=>reset,s=>p(230)(42),cout=>p(231)(43));
FA_ff_6434:FAff port map(x=>p(152)(43),y=>p(153)(43),Cin=>p(154)(43),clock=>clock,reset=>reset,s=>p(230)(43),cout=>p(231)(44));
FA_ff_6435:FAff port map(x=>p(152)(44),y=>p(153)(44),Cin=>p(154)(44),clock=>clock,reset=>reset,s=>p(230)(44),cout=>p(231)(45));
FA_ff_6436:FAff port map(x=>p(152)(45),y=>p(153)(45),Cin=>p(154)(45),clock=>clock,reset=>reset,s=>p(230)(45),cout=>p(231)(46));
FA_ff_6437:FAff port map(x=>p(152)(46),y=>p(153)(46),Cin=>p(154)(46),clock=>clock,reset=>reset,s=>p(230)(46),cout=>p(231)(47));
FA_ff_6438:FAff port map(x=>p(152)(47),y=>p(153)(47),Cin=>p(154)(47),clock=>clock,reset=>reset,s=>p(230)(47),cout=>p(231)(48));
FA_ff_6439:FAff port map(x=>p(152)(48),y=>p(153)(48),Cin=>p(154)(48),clock=>clock,reset=>reset,s=>p(230)(48),cout=>p(231)(49));
FA_ff_6440:FAff port map(x=>p(152)(49),y=>p(153)(49),Cin=>p(154)(49),clock=>clock,reset=>reset,s=>p(230)(49),cout=>p(231)(50));
FA_ff_6441:FAff port map(x=>p(152)(50),y=>p(153)(50),Cin=>p(154)(50),clock=>clock,reset=>reset,s=>p(230)(50),cout=>p(231)(51));
FA_ff_6442:FAff port map(x=>p(152)(51),y=>p(153)(51),Cin=>p(154)(51),clock=>clock,reset=>reset,s=>p(230)(51),cout=>p(231)(52));
FA_ff_6443:FAff port map(x=>p(152)(52),y=>p(153)(52),Cin=>p(154)(52),clock=>clock,reset=>reset,s=>p(230)(52),cout=>p(231)(53));
FA_ff_6444:FAff port map(x=>p(152)(53),y=>p(153)(53),Cin=>p(154)(53),clock=>clock,reset=>reset,s=>p(230)(53),cout=>p(231)(54));
FA_ff_6445:FAff port map(x=>p(152)(54),y=>p(153)(54),Cin=>p(154)(54),clock=>clock,reset=>reset,s=>p(230)(54),cout=>p(231)(55));
FA_ff_6446:FAff port map(x=>p(152)(55),y=>p(153)(55),Cin=>p(154)(55),clock=>clock,reset=>reset,s=>p(230)(55),cout=>p(231)(56));
FA_ff_6447:FAff port map(x=>p(152)(56),y=>p(153)(56),Cin=>p(154)(56),clock=>clock,reset=>reset,s=>p(230)(56),cout=>p(231)(57));
FA_ff_6448:FAff port map(x=>p(152)(57),y=>p(153)(57),Cin=>p(154)(57),clock=>clock,reset=>reset,s=>p(230)(57),cout=>p(231)(58));
FA_ff_6449:FAff port map(x=>p(152)(58),y=>p(153)(58),Cin=>p(154)(58),clock=>clock,reset=>reset,s=>p(230)(58),cout=>p(231)(59));
FA_ff_6450:FAff port map(x=>p(152)(59),y=>p(153)(59),Cin=>p(154)(59),clock=>clock,reset=>reset,s=>p(230)(59),cout=>p(231)(60));
FA_ff_6451:FAff port map(x=>p(152)(60),y=>p(153)(60),Cin=>p(154)(60),clock=>clock,reset=>reset,s=>p(230)(60),cout=>p(231)(61));
FA_ff_6452:FAff port map(x=>p(152)(61),y=>p(153)(61),Cin=>p(154)(61),clock=>clock,reset=>reset,s=>p(230)(61),cout=>p(231)(62));
FA_ff_6453:FAff port map(x=>p(152)(62),y=>p(153)(62),Cin=>p(154)(62),clock=>clock,reset=>reset,s=>p(230)(62),cout=>p(231)(63));
FA_ff_6454:FAff port map(x=>p(152)(63),y=>p(153)(63),Cin=>p(154)(63),clock=>clock,reset=>reset,s=>p(230)(63),cout=>p(231)(64));
FA_ff_6455:FAff port map(x=>p(152)(64),y=>p(153)(64),Cin=>p(154)(64),clock=>clock,reset=>reset,s=>p(230)(64),cout=>p(231)(65));
FA_ff_6456:FAff port map(x=>p(152)(65),y=>p(153)(65),Cin=>p(154)(65),clock=>clock,reset=>reset,s=>p(230)(65),cout=>p(231)(66));
FA_ff_6457:FAff port map(x=>p(152)(66),y=>p(153)(66),Cin=>p(154)(66),clock=>clock,reset=>reset,s=>p(230)(66),cout=>p(231)(67));
FA_ff_6458:FAff port map(x=>p(152)(67),y=>p(153)(67),Cin=>p(154)(67),clock=>clock,reset=>reset,s=>p(230)(67),cout=>p(231)(68));
FA_ff_6459:FAff port map(x=>p(152)(68),y=>p(153)(68),Cin=>p(154)(68),clock=>clock,reset=>reset,s=>p(230)(68),cout=>p(231)(69));
FA_ff_6460:FAff port map(x=>p(152)(69),y=>p(153)(69),Cin=>p(154)(69),clock=>clock,reset=>reset,s=>p(230)(69),cout=>p(231)(70));
FA_ff_6461:FAff port map(x=>p(152)(70),y=>p(153)(70),Cin=>p(154)(70),clock=>clock,reset=>reset,s=>p(230)(70),cout=>p(231)(71));
FA_ff_6462:FAff port map(x=>p(152)(71),y=>p(153)(71),Cin=>p(154)(71),clock=>clock,reset=>reset,s=>p(230)(71),cout=>p(231)(72));
FA_ff_6463:FAff port map(x=>p(152)(72),y=>p(153)(72),Cin=>p(154)(72),clock=>clock,reset=>reset,s=>p(230)(72),cout=>p(231)(73));
FA_ff_6464:FAff port map(x=>p(152)(73),y=>p(153)(73),Cin=>p(154)(73),clock=>clock,reset=>reset,s=>p(230)(73),cout=>p(231)(74));
FA_ff_6465:FAff port map(x=>p(152)(74),y=>p(153)(74),Cin=>p(154)(74),clock=>clock,reset=>reset,s=>p(230)(74),cout=>p(231)(75));
FA_ff_6466:FAff port map(x=>p(152)(75),y=>p(153)(75),Cin=>p(154)(75),clock=>clock,reset=>reset,s=>p(230)(75),cout=>p(231)(76));
FA_ff_6467:FAff port map(x=>p(152)(76),y=>p(153)(76),Cin=>p(154)(76),clock=>clock,reset=>reset,s=>p(230)(76),cout=>p(231)(77));
FA_ff_6468:FAff port map(x=>p(152)(77),y=>p(153)(77),Cin=>p(154)(77),clock=>clock,reset=>reset,s=>p(230)(77),cout=>p(231)(78));
FA_ff_6469:FAff port map(x=>p(152)(78),y=>p(153)(78),Cin=>p(154)(78),clock=>clock,reset=>reset,s=>p(230)(78),cout=>p(231)(79));
FA_ff_6470:FAff port map(x=>p(152)(79),y=>p(153)(79),Cin=>p(154)(79),clock=>clock,reset=>reset,s=>p(230)(79),cout=>p(231)(80));
FA_ff_6471:FAff port map(x=>p(152)(80),y=>p(153)(80),Cin=>p(154)(80),clock=>clock,reset=>reset,s=>p(230)(80),cout=>p(231)(81));
FA_ff_6472:FAff port map(x=>p(152)(81),y=>p(153)(81),Cin=>p(154)(81),clock=>clock,reset=>reset,s=>p(230)(81),cout=>p(231)(82));
FA_ff_6473:FAff port map(x=>p(152)(82),y=>p(153)(82),Cin=>p(154)(82),clock=>clock,reset=>reset,s=>p(230)(82),cout=>p(231)(83));
FA_ff_6474:FAff port map(x=>p(152)(83),y=>p(153)(83),Cin=>p(154)(83),clock=>clock,reset=>reset,s=>p(230)(83),cout=>p(231)(84));
FA_ff_6475:FAff port map(x=>p(152)(84),y=>p(153)(84),Cin=>p(154)(84),clock=>clock,reset=>reset,s=>p(230)(84),cout=>p(231)(85));
FA_ff_6476:FAff port map(x=>p(152)(85),y=>p(153)(85),Cin=>p(154)(85),clock=>clock,reset=>reset,s=>p(230)(85),cout=>p(231)(86));
FA_ff_6477:FAff port map(x=>p(152)(86),y=>p(153)(86),Cin=>p(154)(86),clock=>clock,reset=>reset,s=>p(230)(86),cout=>p(231)(87));
FA_ff_6478:FAff port map(x=>p(152)(87),y=>p(153)(87),Cin=>p(154)(87),clock=>clock,reset=>reset,s=>p(230)(87),cout=>p(231)(88));
FA_ff_6479:FAff port map(x=>p(152)(88),y=>p(153)(88),Cin=>p(154)(88),clock=>clock,reset=>reset,s=>p(230)(88),cout=>p(231)(89));
FA_ff_6480:FAff port map(x=>p(152)(89),y=>p(153)(89),Cin=>p(154)(89),clock=>clock,reset=>reset,s=>p(230)(89),cout=>p(231)(90));
FA_ff_6481:FAff port map(x=>p(152)(90),y=>p(153)(90),Cin=>p(154)(90),clock=>clock,reset=>reset,s=>p(230)(90),cout=>p(231)(91));
FA_ff_6482:FAff port map(x=>p(152)(91),y=>p(153)(91),Cin=>p(154)(91),clock=>clock,reset=>reset,s=>p(230)(91),cout=>p(231)(92));
FA_ff_6483:FAff port map(x=>p(152)(92),y=>p(153)(92),Cin=>p(154)(92),clock=>clock,reset=>reset,s=>p(230)(92),cout=>p(231)(93));
FA_ff_6484:FAff port map(x=>p(152)(93),y=>p(153)(93),Cin=>p(154)(93),clock=>clock,reset=>reset,s=>p(230)(93),cout=>p(231)(94));
FA_ff_6485:FAff port map(x=>p(152)(94),y=>p(153)(94),Cin=>p(154)(94),clock=>clock,reset=>reset,s=>p(230)(94),cout=>p(231)(95));
FA_ff_6486:FAff port map(x=>p(152)(95),y=>p(153)(95),Cin=>p(154)(95),clock=>clock,reset=>reset,s=>p(230)(95),cout=>p(231)(96));
FA_ff_6487:FAff port map(x=>p(152)(96),y=>p(153)(96),Cin=>p(154)(96),clock=>clock,reset=>reset,s=>p(230)(96),cout=>p(231)(97));
FA_ff_6488:FAff port map(x=>p(152)(97),y=>p(153)(97),Cin=>p(154)(97),clock=>clock,reset=>reset,s=>p(230)(97),cout=>p(231)(98));
FA_ff_6489:FAff port map(x=>p(152)(98),y=>p(153)(98),Cin=>p(154)(98),clock=>clock,reset=>reset,s=>p(230)(98),cout=>p(231)(99));
FA_ff_6490:FAff port map(x=>p(152)(99),y=>p(153)(99),Cin=>p(154)(99),clock=>clock,reset=>reset,s=>p(230)(99),cout=>p(231)(100));
FA_ff_6491:FAff port map(x=>p(152)(100),y=>p(153)(100),Cin=>p(154)(100),clock=>clock,reset=>reset,s=>p(230)(100),cout=>p(231)(101));
FA_ff_6492:FAff port map(x=>p(152)(101),y=>p(153)(101),Cin=>p(154)(101),clock=>clock,reset=>reset,s=>p(230)(101),cout=>p(231)(102));
FA_ff_6493:FAff port map(x=>p(152)(102),y=>p(153)(102),Cin=>p(154)(102),clock=>clock,reset=>reset,s=>p(230)(102),cout=>p(231)(103));
FA_ff_6494:FAff port map(x=>p(152)(103),y=>p(153)(103),Cin=>p(154)(103),clock=>clock,reset=>reset,s=>p(230)(103),cout=>p(231)(104));
FA_ff_6495:FAff port map(x=>p(152)(104),y=>p(153)(104),Cin=>p(154)(104),clock=>clock,reset=>reset,s=>p(230)(104),cout=>p(231)(105));
FA_ff_6496:FAff port map(x=>p(152)(105),y=>p(153)(105),Cin=>p(154)(105),clock=>clock,reset=>reset,s=>p(230)(105),cout=>p(231)(106));
FA_ff_6497:FAff port map(x=>p(152)(106),y=>p(153)(106),Cin=>p(154)(106),clock=>clock,reset=>reset,s=>p(230)(106),cout=>p(231)(107));
FA_ff_6498:FAff port map(x=>p(152)(107),y=>p(153)(107),Cin=>p(154)(107),clock=>clock,reset=>reset,s=>p(230)(107),cout=>p(231)(108));
FA_ff_6499:FAff port map(x=>p(152)(108),y=>p(153)(108),Cin=>p(154)(108),clock=>clock,reset=>reset,s=>p(230)(108),cout=>p(231)(109));
FA_ff_6500:FAff port map(x=>p(152)(109),y=>p(153)(109),Cin=>p(154)(109),clock=>clock,reset=>reset,s=>p(230)(109),cout=>p(231)(110));
FA_ff_6501:FAff port map(x=>p(152)(110),y=>p(153)(110),Cin=>p(154)(110),clock=>clock,reset=>reset,s=>p(230)(110),cout=>p(231)(111));
FA_ff_6502:FAff port map(x=>p(152)(111),y=>p(153)(111),Cin=>p(154)(111),clock=>clock,reset=>reset,s=>p(230)(111),cout=>p(231)(112));
FA_ff_6503:FAff port map(x=>p(152)(112),y=>p(153)(112),Cin=>p(154)(112),clock=>clock,reset=>reset,s=>p(230)(112),cout=>p(231)(113));
FA_ff_6504:FAff port map(x=>p(152)(113),y=>p(153)(113),Cin=>p(154)(113),clock=>clock,reset=>reset,s=>p(230)(113),cout=>p(231)(114));
FA_ff_6505:FAff port map(x=>p(152)(114),y=>p(153)(114),Cin=>p(154)(114),clock=>clock,reset=>reset,s=>p(230)(114),cout=>p(231)(115));
FA_ff_6506:FAff port map(x=>p(152)(115),y=>p(153)(115),Cin=>p(154)(115),clock=>clock,reset=>reset,s=>p(230)(115),cout=>p(231)(116));
FA_ff_6507:FAff port map(x=>p(152)(116),y=>p(153)(116),Cin=>p(154)(116),clock=>clock,reset=>reset,s=>p(230)(116),cout=>p(231)(117));
FA_ff_6508:FAff port map(x=>p(152)(117),y=>p(153)(117),Cin=>p(154)(117),clock=>clock,reset=>reset,s=>p(230)(117),cout=>p(231)(118));
FA_ff_6509:FAff port map(x=>p(152)(118),y=>p(153)(118),Cin=>p(154)(118),clock=>clock,reset=>reset,s=>p(230)(118),cout=>p(231)(119));
FA_ff_6510:FAff port map(x=>p(152)(119),y=>p(153)(119),Cin=>p(154)(119),clock=>clock,reset=>reset,s=>p(230)(119),cout=>p(231)(120));
FA_ff_6511:FAff port map(x=>p(152)(120),y=>p(153)(120),Cin=>p(154)(120),clock=>clock,reset=>reset,s=>p(230)(120),cout=>p(231)(121));
FA_ff_6512:FAff port map(x=>p(152)(121),y=>p(153)(121),Cin=>p(154)(121),clock=>clock,reset=>reset,s=>p(230)(121),cout=>p(231)(122));
FA_ff_6513:FAff port map(x=>p(152)(122),y=>p(153)(122),Cin=>p(154)(122),clock=>clock,reset=>reset,s=>p(230)(122),cout=>p(231)(123));
FA_ff_6514:FAff port map(x=>p(152)(123),y=>p(153)(123),Cin=>p(154)(123),clock=>clock,reset=>reset,s=>p(230)(123),cout=>p(231)(124));
FA_ff_6515:FAff port map(x=>p(152)(124),y=>p(153)(124),Cin=>p(154)(124),clock=>clock,reset=>reset,s=>p(230)(124),cout=>p(231)(125));
FA_ff_6516:FAff port map(x=>p(152)(125),y=>p(153)(125),Cin=>p(154)(125),clock=>clock,reset=>reset,s=>p(230)(125),cout=>p(231)(126));
FA_ff_6517:FAff port map(x=>p(152)(126),y=>p(153)(126),Cin=>p(154)(126),clock=>clock,reset=>reset,s=>p(230)(126),cout=>p(231)(127));
FA_ff_6518:FAff port map(x=>p(152)(127),y=>p(153)(127),Cin=>p(154)(127),clock=>clock,reset=>reset,s=>p(230)(127),cout=>p(231)(128));
p(230)(128)<=p(153)(128);
p(232)(0)<=p(156)(0);
FA_ff_6519:FAff port map(x=>p(155)(1),y=>p(156)(1),Cin=>p(157)(1),clock=>clock,reset=>reset,s=>p(232)(1),cout=>p(233)(2));
FA_ff_6520:FAff port map(x=>p(155)(2),y=>p(156)(2),Cin=>p(157)(2),clock=>clock,reset=>reset,s=>p(232)(2),cout=>p(233)(3));
FA_ff_6521:FAff port map(x=>p(155)(3),y=>p(156)(3),Cin=>p(157)(3),clock=>clock,reset=>reset,s=>p(232)(3),cout=>p(233)(4));
FA_ff_6522:FAff port map(x=>p(155)(4),y=>p(156)(4),Cin=>p(157)(4),clock=>clock,reset=>reset,s=>p(232)(4),cout=>p(233)(5));
FA_ff_6523:FAff port map(x=>p(155)(5),y=>p(156)(5),Cin=>p(157)(5),clock=>clock,reset=>reset,s=>p(232)(5),cout=>p(233)(6));
FA_ff_6524:FAff port map(x=>p(155)(6),y=>p(156)(6),Cin=>p(157)(6),clock=>clock,reset=>reset,s=>p(232)(6),cout=>p(233)(7));
FA_ff_6525:FAff port map(x=>p(155)(7),y=>p(156)(7),Cin=>p(157)(7),clock=>clock,reset=>reset,s=>p(232)(7),cout=>p(233)(8));
FA_ff_6526:FAff port map(x=>p(155)(8),y=>p(156)(8),Cin=>p(157)(8),clock=>clock,reset=>reset,s=>p(232)(8),cout=>p(233)(9));
FA_ff_6527:FAff port map(x=>p(155)(9),y=>p(156)(9),Cin=>p(157)(9),clock=>clock,reset=>reset,s=>p(232)(9),cout=>p(233)(10));
FA_ff_6528:FAff port map(x=>p(155)(10),y=>p(156)(10),Cin=>p(157)(10),clock=>clock,reset=>reset,s=>p(232)(10),cout=>p(233)(11));
FA_ff_6529:FAff port map(x=>p(155)(11),y=>p(156)(11),Cin=>p(157)(11),clock=>clock,reset=>reset,s=>p(232)(11),cout=>p(233)(12));
FA_ff_6530:FAff port map(x=>p(155)(12),y=>p(156)(12),Cin=>p(157)(12),clock=>clock,reset=>reset,s=>p(232)(12),cout=>p(233)(13));
FA_ff_6531:FAff port map(x=>p(155)(13),y=>p(156)(13),Cin=>p(157)(13),clock=>clock,reset=>reset,s=>p(232)(13),cout=>p(233)(14));
FA_ff_6532:FAff port map(x=>p(155)(14),y=>p(156)(14),Cin=>p(157)(14),clock=>clock,reset=>reset,s=>p(232)(14),cout=>p(233)(15));
FA_ff_6533:FAff port map(x=>p(155)(15),y=>p(156)(15),Cin=>p(157)(15),clock=>clock,reset=>reset,s=>p(232)(15),cout=>p(233)(16));
FA_ff_6534:FAff port map(x=>p(155)(16),y=>p(156)(16),Cin=>p(157)(16),clock=>clock,reset=>reset,s=>p(232)(16),cout=>p(233)(17));
FA_ff_6535:FAff port map(x=>p(155)(17),y=>p(156)(17),Cin=>p(157)(17),clock=>clock,reset=>reset,s=>p(232)(17),cout=>p(233)(18));
FA_ff_6536:FAff port map(x=>p(155)(18),y=>p(156)(18),Cin=>p(157)(18),clock=>clock,reset=>reset,s=>p(232)(18),cout=>p(233)(19));
FA_ff_6537:FAff port map(x=>p(155)(19),y=>p(156)(19),Cin=>p(157)(19),clock=>clock,reset=>reset,s=>p(232)(19),cout=>p(233)(20));
FA_ff_6538:FAff port map(x=>p(155)(20),y=>p(156)(20),Cin=>p(157)(20),clock=>clock,reset=>reset,s=>p(232)(20),cout=>p(233)(21));
FA_ff_6539:FAff port map(x=>p(155)(21),y=>p(156)(21),Cin=>p(157)(21),clock=>clock,reset=>reset,s=>p(232)(21),cout=>p(233)(22));
FA_ff_6540:FAff port map(x=>p(155)(22),y=>p(156)(22),Cin=>p(157)(22),clock=>clock,reset=>reset,s=>p(232)(22),cout=>p(233)(23));
FA_ff_6541:FAff port map(x=>p(155)(23),y=>p(156)(23),Cin=>p(157)(23),clock=>clock,reset=>reset,s=>p(232)(23),cout=>p(233)(24));
FA_ff_6542:FAff port map(x=>p(155)(24),y=>p(156)(24),Cin=>p(157)(24),clock=>clock,reset=>reset,s=>p(232)(24),cout=>p(233)(25));
FA_ff_6543:FAff port map(x=>p(155)(25),y=>p(156)(25),Cin=>p(157)(25),clock=>clock,reset=>reset,s=>p(232)(25),cout=>p(233)(26));
FA_ff_6544:FAff port map(x=>p(155)(26),y=>p(156)(26),Cin=>p(157)(26),clock=>clock,reset=>reset,s=>p(232)(26),cout=>p(233)(27));
FA_ff_6545:FAff port map(x=>p(155)(27),y=>p(156)(27),Cin=>p(157)(27),clock=>clock,reset=>reset,s=>p(232)(27),cout=>p(233)(28));
FA_ff_6546:FAff port map(x=>p(155)(28),y=>p(156)(28),Cin=>p(157)(28),clock=>clock,reset=>reset,s=>p(232)(28),cout=>p(233)(29));
FA_ff_6547:FAff port map(x=>p(155)(29),y=>p(156)(29),Cin=>p(157)(29),clock=>clock,reset=>reset,s=>p(232)(29),cout=>p(233)(30));
FA_ff_6548:FAff port map(x=>p(155)(30),y=>p(156)(30),Cin=>p(157)(30),clock=>clock,reset=>reset,s=>p(232)(30),cout=>p(233)(31));
FA_ff_6549:FAff port map(x=>p(155)(31),y=>p(156)(31),Cin=>p(157)(31),clock=>clock,reset=>reset,s=>p(232)(31),cout=>p(233)(32));
FA_ff_6550:FAff port map(x=>p(155)(32),y=>p(156)(32),Cin=>p(157)(32),clock=>clock,reset=>reset,s=>p(232)(32),cout=>p(233)(33));
FA_ff_6551:FAff port map(x=>p(155)(33),y=>p(156)(33),Cin=>p(157)(33),clock=>clock,reset=>reset,s=>p(232)(33),cout=>p(233)(34));
FA_ff_6552:FAff port map(x=>p(155)(34),y=>p(156)(34),Cin=>p(157)(34),clock=>clock,reset=>reset,s=>p(232)(34),cout=>p(233)(35));
FA_ff_6553:FAff port map(x=>p(155)(35),y=>p(156)(35),Cin=>p(157)(35),clock=>clock,reset=>reset,s=>p(232)(35),cout=>p(233)(36));
FA_ff_6554:FAff port map(x=>p(155)(36),y=>p(156)(36),Cin=>p(157)(36),clock=>clock,reset=>reset,s=>p(232)(36),cout=>p(233)(37));
FA_ff_6555:FAff port map(x=>p(155)(37),y=>p(156)(37),Cin=>p(157)(37),clock=>clock,reset=>reset,s=>p(232)(37),cout=>p(233)(38));
FA_ff_6556:FAff port map(x=>p(155)(38),y=>p(156)(38),Cin=>p(157)(38),clock=>clock,reset=>reset,s=>p(232)(38),cout=>p(233)(39));
FA_ff_6557:FAff port map(x=>p(155)(39),y=>p(156)(39),Cin=>p(157)(39),clock=>clock,reset=>reset,s=>p(232)(39),cout=>p(233)(40));
FA_ff_6558:FAff port map(x=>p(155)(40),y=>p(156)(40),Cin=>p(157)(40),clock=>clock,reset=>reset,s=>p(232)(40),cout=>p(233)(41));
FA_ff_6559:FAff port map(x=>p(155)(41),y=>p(156)(41),Cin=>p(157)(41),clock=>clock,reset=>reset,s=>p(232)(41),cout=>p(233)(42));
FA_ff_6560:FAff port map(x=>p(155)(42),y=>p(156)(42),Cin=>p(157)(42),clock=>clock,reset=>reset,s=>p(232)(42),cout=>p(233)(43));
FA_ff_6561:FAff port map(x=>p(155)(43),y=>p(156)(43),Cin=>p(157)(43),clock=>clock,reset=>reset,s=>p(232)(43),cout=>p(233)(44));
FA_ff_6562:FAff port map(x=>p(155)(44),y=>p(156)(44),Cin=>p(157)(44),clock=>clock,reset=>reset,s=>p(232)(44),cout=>p(233)(45));
FA_ff_6563:FAff port map(x=>p(155)(45),y=>p(156)(45),Cin=>p(157)(45),clock=>clock,reset=>reset,s=>p(232)(45),cout=>p(233)(46));
FA_ff_6564:FAff port map(x=>p(155)(46),y=>p(156)(46),Cin=>p(157)(46),clock=>clock,reset=>reset,s=>p(232)(46),cout=>p(233)(47));
FA_ff_6565:FAff port map(x=>p(155)(47),y=>p(156)(47),Cin=>p(157)(47),clock=>clock,reset=>reset,s=>p(232)(47),cout=>p(233)(48));
FA_ff_6566:FAff port map(x=>p(155)(48),y=>p(156)(48),Cin=>p(157)(48),clock=>clock,reset=>reset,s=>p(232)(48),cout=>p(233)(49));
FA_ff_6567:FAff port map(x=>p(155)(49),y=>p(156)(49),Cin=>p(157)(49),clock=>clock,reset=>reset,s=>p(232)(49),cout=>p(233)(50));
FA_ff_6568:FAff port map(x=>p(155)(50),y=>p(156)(50),Cin=>p(157)(50),clock=>clock,reset=>reset,s=>p(232)(50),cout=>p(233)(51));
FA_ff_6569:FAff port map(x=>p(155)(51),y=>p(156)(51),Cin=>p(157)(51),clock=>clock,reset=>reset,s=>p(232)(51),cout=>p(233)(52));
FA_ff_6570:FAff port map(x=>p(155)(52),y=>p(156)(52),Cin=>p(157)(52),clock=>clock,reset=>reset,s=>p(232)(52),cout=>p(233)(53));
FA_ff_6571:FAff port map(x=>p(155)(53),y=>p(156)(53),Cin=>p(157)(53),clock=>clock,reset=>reset,s=>p(232)(53),cout=>p(233)(54));
FA_ff_6572:FAff port map(x=>p(155)(54),y=>p(156)(54),Cin=>p(157)(54),clock=>clock,reset=>reset,s=>p(232)(54),cout=>p(233)(55));
FA_ff_6573:FAff port map(x=>p(155)(55),y=>p(156)(55),Cin=>p(157)(55),clock=>clock,reset=>reset,s=>p(232)(55),cout=>p(233)(56));
FA_ff_6574:FAff port map(x=>p(155)(56),y=>p(156)(56),Cin=>p(157)(56),clock=>clock,reset=>reset,s=>p(232)(56),cout=>p(233)(57));
FA_ff_6575:FAff port map(x=>p(155)(57),y=>p(156)(57),Cin=>p(157)(57),clock=>clock,reset=>reset,s=>p(232)(57),cout=>p(233)(58));
FA_ff_6576:FAff port map(x=>p(155)(58),y=>p(156)(58),Cin=>p(157)(58),clock=>clock,reset=>reset,s=>p(232)(58),cout=>p(233)(59));
FA_ff_6577:FAff port map(x=>p(155)(59),y=>p(156)(59),Cin=>p(157)(59),clock=>clock,reset=>reset,s=>p(232)(59),cout=>p(233)(60));
FA_ff_6578:FAff port map(x=>p(155)(60),y=>p(156)(60),Cin=>p(157)(60),clock=>clock,reset=>reset,s=>p(232)(60),cout=>p(233)(61));
FA_ff_6579:FAff port map(x=>p(155)(61),y=>p(156)(61),Cin=>p(157)(61),clock=>clock,reset=>reset,s=>p(232)(61),cout=>p(233)(62));
FA_ff_6580:FAff port map(x=>p(155)(62),y=>p(156)(62),Cin=>p(157)(62),clock=>clock,reset=>reset,s=>p(232)(62),cout=>p(233)(63));
FA_ff_6581:FAff port map(x=>p(155)(63),y=>p(156)(63),Cin=>p(157)(63),clock=>clock,reset=>reset,s=>p(232)(63),cout=>p(233)(64));
FA_ff_6582:FAff port map(x=>p(155)(64),y=>p(156)(64),Cin=>p(157)(64),clock=>clock,reset=>reset,s=>p(232)(64),cout=>p(233)(65));
FA_ff_6583:FAff port map(x=>p(155)(65),y=>p(156)(65),Cin=>p(157)(65),clock=>clock,reset=>reset,s=>p(232)(65),cout=>p(233)(66));
FA_ff_6584:FAff port map(x=>p(155)(66),y=>p(156)(66),Cin=>p(157)(66),clock=>clock,reset=>reset,s=>p(232)(66),cout=>p(233)(67));
FA_ff_6585:FAff port map(x=>p(155)(67),y=>p(156)(67),Cin=>p(157)(67),clock=>clock,reset=>reset,s=>p(232)(67),cout=>p(233)(68));
FA_ff_6586:FAff port map(x=>p(155)(68),y=>p(156)(68),Cin=>p(157)(68),clock=>clock,reset=>reset,s=>p(232)(68),cout=>p(233)(69));
FA_ff_6587:FAff port map(x=>p(155)(69),y=>p(156)(69),Cin=>p(157)(69),clock=>clock,reset=>reset,s=>p(232)(69),cout=>p(233)(70));
FA_ff_6588:FAff port map(x=>p(155)(70),y=>p(156)(70),Cin=>p(157)(70),clock=>clock,reset=>reset,s=>p(232)(70),cout=>p(233)(71));
FA_ff_6589:FAff port map(x=>p(155)(71),y=>p(156)(71),Cin=>p(157)(71),clock=>clock,reset=>reset,s=>p(232)(71),cout=>p(233)(72));
FA_ff_6590:FAff port map(x=>p(155)(72),y=>p(156)(72),Cin=>p(157)(72),clock=>clock,reset=>reset,s=>p(232)(72),cout=>p(233)(73));
FA_ff_6591:FAff port map(x=>p(155)(73),y=>p(156)(73),Cin=>p(157)(73),clock=>clock,reset=>reset,s=>p(232)(73),cout=>p(233)(74));
FA_ff_6592:FAff port map(x=>p(155)(74),y=>p(156)(74),Cin=>p(157)(74),clock=>clock,reset=>reset,s=>p(232)(74),cout=>p(233)(75));
FA_ff_6593:FAff port map(x=>p(155)(75),y=>p(156)(75),Cin=>p(157)(75),clock=>clock,reset=>reset,s=>p(232)(75),cout=>p(233)(76));
FA_ff_6594:FAff port map(x=>p(155)(76),y=>p(156)(76),Cin=>p(157)(76),clock=>clock,reset=>reset,s=>p(232)(76),cout=>p(233)(77));
FA_ff_6595:FAff port map(x=>p(155)(77),y=>p(156)(77),Cin=>p(157)(77),clock=>clock,reset=>reset,s=>p(232)(77),cout=>p(233)(78));
FA_ff_6596:FAff port map(x=>p(155)(78),y=>p(156)(78),Cin=>p(157)(78),clock=>clock,reset=>reset,s=>p(232)(78),cout=>p(233)(79));
FA_ff_6597:FAff port map(x=>p(155)(79),y=>p(156)(79),Cin=>p(157)(79),clock=>clock,reset=>reset,s=>p(232)(79),cout=>p(233)(80));
FA_ff_6598:FAff port map(x=>p(155)(80),y=>p(156)(80),Cin=>p(157)(80),clock=>clock,reset=>reset,s=>p(232)(80),cout=>p(233)(81));
FA_ff_6599:FAff port map(x=>p(155)(81),y=>p(156)(81),Cin=>p(157)(81),clock=>clock,reset=>reset,s=>p(232)(81),cout=>p(233)(82));
FA_ff_6600:FAff port map(x=>p(155)(82),y=>p(156)(82),Cin=>p(157)(82),clock=>clock,reset=>reset,s=>p(232)(82),cout=>p(233)(83));
FA_ff_6601:FAff port map(x=>p(155)(83),y=>p(156)(83),Cin=>p(157)(83),clock=>clock,reset=>reset,s=>p(232)(83),cout=>p(233)(84));
FA_ff_6602:FAff port map(x=>p(155)(84),y=>p(156)(84),Cin=>p(157)(84),clock=>clock,reset=>reset,s=>p(232)(84),cout=>p(233)(85));
FA_ff_6603:FAff port map(x=>p(155)(85),y=>p(156)(85),Cin=>p(157)(85),clock=>clock,reset=>reset,s=>p(232)(85),cout=>p(233)(86));
FA_ff_6604:FAff port map(x=>p(155)(86),y=>p(156)(86),Cin=>p(157)(86),clock=>clock,reset=>reset,s=>p(232)(86),cout=>p(233)(87));
FA_ff_6605:FAff port map(x=>p(155)(87),y=>p(156)(87),Cin=>p(157)(87),clock=>clock,reset=>reset,s=>p(232)(87),cout=>p(233)(88));
FA_ff_6606:FAff port map(x=>p(155)(88),y=>p(156)(88),Cin=>p(157)(88),clock=>clock,reset=>reset,s=>p(232)(88),cout=>p(233)(89));
FA_ff_6607:FAff port map(x=>p(155)(89),y=>p(156)(89),Cin=>p(157)(89),clock=>clock,reset=>reset,s=>p(232)(89),cout=>p(233)(90));
FA_ff_6608:FAff port map(x=>p(155)(90),y=>p(156)(90),Cin=>p(157)(90),clock=>clock,reset=>reset,s=>p(232)(90),cout=>p(233)(91));
FA_ff_6609:FAff port map(x=>p(155)(91),y=>p(156)(91),Cin=>p(157)(91),clock=>clock,reset=>reset,s=>p(232)(91),cout=>p(233)(92));
FA_ff_6610:FAff port map(x=>p(155)(92),y=>p(156)(92),Cin=>p(157)(92),clock=>clock,reset=>reset,s=>p(232)(92),cout=>p(233)(93));
FA_ff_6611:FAff port map(x=>p(155)(93),y=>p(156)(93),Cin=>p(157)(93),clock=>clock,reset=>reset,s=>p(232)(93),cout=>p(233)(94));
FA_ff_6612:FAff port map(x=>p(155)(94),y=>p(156)(94),Cin=>p(157)(94),clock=>clock,reset=>reset,s=>p(232)(94),cout=>p(233)(95));
FA_ff_6613:FAff port map(x=>p(155)(95),y=>p(156)(95),Cin=>p(157)(95),clock=>clock,reset=>reset,s=>p(232)(95),cout=>p(233)(96));
FA_ff_6614:FAff port map(x=>p(155)(96),y=>p(156)(96),Cin=>p(157)(96),clock=>clock,reset=>reset,s=>p(232)(96),cout=>p(233)(97));
FA_ff_6615:FAff port map(x=>p(155)(97),y=>p(156)(97),Cin=>p(157)(97),clock=>clock,reset=>reset,s=>p(232)(97),cout=>p(233)(98));
FA_ff_6616:FAff port map(x=>p(155)(98),y=>p(156)(98),Cin=>p(157)(98),clock=>clock,reset=>reset,s=>p(232)(98),cout=>p(233)(99));
FA_ff_6617:FAff port map(x=>p(155)(99),y=>p(156)(99),Cin=>p(157)(99),clock=>clock,reset=>reset,s=>p(232)(99),cout=>p(233)(100));
FA_ff_6618:FAff port map(x=>p(155)(100),y=>p(156)(100),Cin=>p(157)(100),clock=>clock,reset=>reset,s=>p(232)(100),cout=>p(233)(101));
FA_ff_6619:FAff port map(x=>p(155)(101),y=>p(156)(101),Cin=>p(157)(101),clock=>clock,reset=>reset,s=>p(232)(101),cout=>p(233)(102));
FA_ff_6620:FAff port map(x=>p(155)(102),y=>p(156)(102),Cin=>p(157)(102),clock=>clock,reset=>reset,s=>p(232)(102),cout=>p(233)(103));
FA_ff_6621:FAff port map(x=>p(155)(103),y=>p(156)(103),Cin=>p(157)(103),clock=>clock,reset=>reset,s=>p(232)(103),cout=>p(233)(104));
FA_ff_6622:FAff port map(x=>p(155)(104),y=>p(156)(104),Cin=>p(157)(104),clock=>clock,reset=>reset,s=>p(232)(104),cout=>p(233)(105));
FA_ff_6623:FAff port map(x=>p(155)(105),y=>p(156)(105),Cin=>p(157)(105),clock=>clock,reset=>reset,s=>p(232)(105),cout=>p(233)(106));
FA_ff_6624:FAff port map(x=>p(155)(106),y=>p(156)(106),Cin=>p(157)(106),clock=>clock,reset=>reset,s=>p(232)(106),cout=>p(233)(107));
FA_ff_6625:FAff port map(x=>p(155)(107),y=>p(156)(107),Cin=>p(157)(107),clock=>clock,reset=>reset,s=>p(232)(107),cout=>p(233)(108));
FA_ff_6626:FAff port map(x=>p(155)(108),y=>p(156)(108),Cin=>p(157)(108),clock=>clock,reset=>reset,s=>p(232)(108),cout=>p(233)(109));
FA_ff_6627:FAff port map(x=>p(155)(109),y=>p(156)(109),Cin=>p(157)(109),clock=>clock,reset=>reset,s=>p(232)(109),cout=>p(233)(110));
FA_ff_6628:FAff port map(x=>p(155)(110),y=>p(156)(110),Cin=>p(157)(110),clock=>clock,reset=>reset,s=>p(232)(110),cout=>p(233)(111));
FA_ff_6629:FAff port map(x=>p(155)(111),y=>p(156)(111),Cin=>p(157)(111),clock=>clock,reset=>reset,s=>p(232)(111),cout=>p(233)(112));
FA_ff_6630:FAff port map(x=>p(155)(112),y=>p(156)(112),Cin=>p(157)(112),clock=>clock,reset=>reset,s=>p(232)(112),cout=>p(233)(113));
FA_ff_6631:FAff port map(x=>p(155)(113),y=>p(156)(113),Cin=>p(157)(113),clock=>clock,reset=>reset,s=>p(232)(113),cout=>p(233)(114));
FA_ff_6632:FAff port map(x=>p(155)(114),y=>p(156)(114),Cin=>p(157)(114),clock=>clock,reset=>reset,s=>p(232)(114),cout=>p(233)(115));
FA_ff_6633:FAff port map(x=>p(155)(115),y=>p(156)(115),Cin=>p(157)(115),clock=>clock,reset=>reset,s=>p(232)(115),cout=>p(233)(116));
FA_ff_6634:FAff port map(x=>p(155)(116),y=>p(156)(116),Cin=>p(157)(116),clock=>clock,reset=>reset,s=>p(232)(116),cout=>p(233)(117));
FA_ff_6635:FAff port map(x=>p(155)(117),y=>p(156)(117),Cin=>p(157)(117),clock=>clock,reset=>reset,s=>p(232)(117),cout=>p(233)(118));
FA_ff_6636:FAff port map(x=>p(155)(118),y=>p(156)(118),Cin=>p(157)(118),clock=>clock,reset=>reset,s=>p(232)(118),cout=>p(233)(119));
FA_ff_6637:FAff port map(x=>p(155)(119),y=>p(156)(119),Cin=>p(157)(119),clock=>clock,reset=>reset,s=>p(232)(119),cout=>p(233)(120));
FA_ff_6638:FAff port map(x=>p(155)(120),y=>p(156)(120),Cin=>p(157)(120),clock=>clock,reset=>reset,s=>p(232)(120),cout=>p(233)(121));
FA_ff_6639:FAff port map(x=>p(155)(121),y=>p(156)(121),Cin=>p(157)(121),clock=>clock,reset=>reset,s=>p(232)(121),cout=>p(233)(122));
FA_ff_6640:FAff port map(x=>p(155)(122),y=>p(156)(122),Cin=>p(157)(122),clock=>clock,reset=>reset,s=>p(232)(122),cout=>p(233)(123));
FA_ff_6641:FAff port map(x=>p(155)(123),y=>p(156)(123),Cin=>p(157)(123),clock=>clock,reset=>reset,s=>p(232)(123),cout=>p(233)(124));
FA_ff_6642:FAff port map(x=>p(155)(124),y=>p(156)(124),Cin=>p(157)(124),clock=>clock,reset=>reset,s=>p(232)(124),cout=>p(233)(125));
FA_ff_6643:FAff port map(x=>p(155)(125),y=>p(156)(125),Cin=>p(157)(125),clock=>clock,reset=>reset,s=>p(232)(125),cout=>p(233)(126));
FA_ff_6644:FAff port map(x=>p(155)(126),y=>p(156)(126),Cin=>p(157)(126),clock=>clock,reset=>reset,s=>p(232)(126),cout=>p(233)(127));
FA_ff_6645:FAff port map(x=>p(155)(127),y=>p(156)(127),Cin=>p(157)(127),clock=>clock,reset=>reset,s=>p(232)(127),cout=>p(233)(128));
HA_ff_9:HAff port map(x=>p(155)(128),y=>p(157)(128),clock=>clock,reset=>reset,s=>p(232)(128),c=>p(233)(129));
HA_ff_10:HAff port map(x=>p(158)(0),y=>p(160)(0),clock=>clock,reset=>reset,s=>p(234)(0),c=>p(235)(1));
FA_ff_6646:FAff port map(x=>p(158)(1),y=>p(159)(1),Cin=>p(160)(1),clock=>clock,reset=>reset,s=>p(234)(1),cout=>p(235)(2));
FA_ff_6647:FAff port map(x=>p(158)(2),y=>p(159)(2),Cin=>p(160)(2),clock=>clock,reset=>reset,s=>p(234)(2),cout=>p(235)(3));
FA_ff_6648:FAff port map(x=>p(158)(3),y=>p(159)(3),Cin=>p(160)(3),clock=>clock,reset=>reset,s=>p(234)(3),cout=>p(235)(4));
FA_ff_6649:FAff port map(x=>p(158)(4),y=>p(159)(4),Cin=>p(160)(4),clock=>clock,reset=>reset,s=>p(234)(4),cout=>p(235)(5));
FA_ff_6650:FAff port map(x=>p(158)(5),y=>p(159)(5),Cin=>p(160)(5),clock=>clock,reset=>reset,s=>p(234)(5),cout=>p(235)(6));
FA_ff_6651:FAff port map(x=>p(158)(6),y=>p(159)(6),Cin=>p(160)(6),clock=>clock,reset=>reset,s=>p(234)(6),cout=>p(235)(7));
FA_ff_6652:FAff port map(x=>p(158)(7),y=>p(159)(7),Cin=>p(160)(7),clock=>clock,reset=>reset,s=>p(234)(7),cout=>p(235)(8));
FA_ff_6653:FAff port map(x=>p(158)(8),y=>p(159)(8),Cin=>p(160)(8),clock=>clock,reset=>reset,s=>p(234)(8),cout=>p(235)(9));
FA_ff_6654:FAff port map(x=>p(158)(9),y=>p(159)(9),Cin=>p(160)(9),clock=>clock,reset=>reset,s=>p(234)(9),cout=>p(235)(10));
FA_ff_6655:FAff port map(x=>p(158)(10),y=>p(159)(10),Cin=>p(160)(10),clock=>clock,reset=>reset,s=>p(234)(10),cout=>p(235)(11));
FA_ff_6656:FAff port map(x=>p(158)(11),y=>p(159)(11),Cin=>p(160)(11),clock=>clock,reset=>reset,s=>p(234)(11),cout=>p(235)(12));
FA_ff_6657:FAff port map(x=>p(158)(12),y=>p(159)(12),Cin=>p(160)(12),clock=>clock,reset=>reset,s=>p(234)(12),cout=>p(235)(13));
FA_ff_6658:FAff port map(x=>p(158)(13),y=>p(159)(13),Cin=>p(160)(13),clock=>clock,reset=>reset,s=>p(234)(13),cout=>p(235)(14));
FA_ff_6659:FAff port map(x=>p(158)(14),y=>p(159)(14),Cin=>p(160)(14),clock=>clock,reset=>reset,s=>p(234)(14),cout=>p(235)(15));
FA_ff_6660:FAff port map(x=>p(158)(15),y=>p(159)(15),Cin=>p(160)(15),clock=>clock,reset=>reset,s=>p(234)(15),cout=>p(235)(16));
FA_ff_6661:FAff port map(x=>p(158)(16),y=>p(159)(16),Cin=>p(160)(16),clock=>clock,reset=>reset,s=>p(234)(16),cout=>p(235)(17));
FA_ff_6662:FAff port map(x=>p(158)(17),y=>p(159)(17),Cin=>p(160)(17),clock=>clock,reset=>reset,s=>p(234)(17),cout=>p(235)(18));
FA_ff_6663:FAff port map(x=>p(158)(18),y=>p(159)(18),Cin=>p(160)(18),clock=>clock,reset=>reset,s=>p(234)(18),cout=>p(235)(19));
FA_ff_6664:FAff port map(x=>p(158)(19),y=>p(159)(19),Cin=>p(160)(19),clock=>clock,reset=>reset,s=>p(234)(19),cout=>p(235)(20));
FA_ff_6665:FAff port map(x=>p(158)(20),y=>p(159)(20),Cin=>p(160)(20),clock=>clock,reset=>reset,s=>p(234)(20),cout=>p(235)(21));
FA_ff_6666:FAff port map(x=>p(158)(21),y=>p(159)(21),Cin=>p(160)(21),clock=>clock,reset=>reset,s=>p(234)(21),cout=>p(235)(22));
FA_ff_6667:FAff port map(x=>p(158)(22),y=>p(159)(22),Cin=>p(160)(22),clock=>clock,reset=>reset,s=>p(234)(22),cout=>p(235)(23));
FA_ff_6668:FAff port map(x=>p(158)(23),y=>p(159)(23),Cin=>p(160)(23),clock=>clock,reset=>reset,s=>p(234)(23),cout=>p(235)(24));
FA_ff_6669:FAff port map(x=>p(158)(24),y=>p(159)(24),Cin=>p(160)(24),clock=>clock,reset=>reset,s=>p(234)(24),cout=>p(235)(25));
FA_ff_6670:FAff port map(x=>p(158)(25),y=>p(159)(25),Cin=>p(160)(25),clock=>clock,reset=>reset,s=>p(234)(25),cout=>p(235)(26));
FA_ff_6671:FAff port map(x=>p(158)(26),y=>p(159)(26),Cin=>p(160)(26),clock=>clock,reset=>reset,s=>p(234)(26),cout=>p(235)(27));
FA_ff_6672:FAff port map(x=>p(158)(27),y=>p(159)(27),Cin=>p(160)(27),clock=>clock,reset=>reset,s=>p(234)(27),cout=>p(235)(28));
FA_ff_6673:FAff port map(x=>p(158)(28),y=>p(159)(28),Cin=>p(160)(28),clock=>clock,reset=>reset,s=>p(234)(28),cout=>p(235)(29));
FA_ff_6674:FAff port map(x=>p(158)(29),y=>p(159)(29),Cin=>p(160)(29),clock=>clock,reset=>reset,s=>p(234)(29),cout=>p(235)(30));
FA_ff_6675:FAff port map(x=>p(158)(30),y=>p(159)(30),Cin=>p(160)(30),clock=>clock,reset=>reset,s=>p(234)(30),cout=>p(235)(31));
FA_ff_6676:FAff port map(x=>p(158)(31),y=>p(159)(31),Cin=>p(160)(31),clock=>clock,reset=>reset,s=>p(234)(31),cout=>p(235)(32));
FA_ff_6677:FAff port map(x=>p(158)(32),y=>p(159)(32),Cin=>p(160)(32),clock=>clock,reset=>reset,s=>p(234)(32),cout=>p(235)(33));
FA_ff_6678:FAff port map(x=>p(158)(33),y=>p(159)(33),Cin=>p(160)(33),clock=>clock,reset=>reset,s=>p(234)(33),cout=>p(235)(34));
FA_ff_6679:FAff port map(x=>p(158)(34),y=>p(159)(34),Cin=>p(160)(34),clock=>clock,reset=>reset,s=>p(234)(34),cout=>p(235)(35));
FA_ff_6680:FAff port map(x=>p(158)(35),y=>p(159)(35),Cin=>p(160)(35),clock=>clock,reset=>reset,s=>p(234)(35),cout=>p(235)(36));
FA_ff_6681:FAff port map(x=>p(158)(36),y=>p(159)(36),Cin=>p(160)(36),clock=>clock,reset=>reset,s=>p(234)(36),cout=>p(235)(37));
FA_ff_6682:FAff port map(x=>p(158)(37),y=>p(159)(37),Cin=>p(160)(37),clock=>clock,reset=>reset,s=>p(234)(37),cout=>p(235)(38));
FA_ff_6683:FAff port map(x=>p(158)(38),y=>p(159)(38),Cin=>p(160)(38),clock=>clock,reset=>reset,s=>p(234)(38),cout=>p(235)(39));
FA_ff_6684:FAff port map(x=>p(158)(39),y=>p(159)(39),Cin=>p(160)(39),clock=>clock,reset=>reset,s=>p(234)(39),cout=>p(235)(40));
FA_ff_6685:FAff port map(x=>p(158)(40),y=>p(159)(40),Cin=>p(160)(40),clock=>clock,reset=>reset,s=>p(234)(40),cout=>p(235)(41));
FA_ff_6686:FAff port map(x=>p(158)(41),y=>p(159)(41),Cin=>p(160)(41),clock=>clock,reset=>reset,s=>p(234)(41),cout=>p(235)(42));
FA_ff_6687:FAff port map(x=>p(158)(42),y=>p(159)(42),Cin=>p(160)(42),clock=>clock,reset=>reset,s=>p(234)(42),cout=>p(235)(43));
FA_ff_6688:FAff port map(x=>p(158)(43),y=>p(159)(43),Cin=>p(160)(43),clock=>clock,reset=>reset,s=>p(234)(43),cout=>p(235)(44));
FA_ff_6689:FAff port map(x=>p(158)(44),y=>p(159)(44),Cin=>p(160)(44),clock=>clock,reset=>reset,s=>p(234)(44),cout=>p(235)(45));
FA_ff_6690:FAff port map(x=>p(158)(45),y=>p(159)(45),Cin=>p(160)(45),clock=>clock,reset=>reset,s=>p(234)(45),cout=>p(235)(46));
FA_ff_6691:FAff port map(x=>p(158)(46),y=>p(159)(46),Cin=>p(160)(46),clock=>clock,reset=>reset,s=>p(234)(46),cout=>p(235)(47));
FA_ff_6692:FAff port map(x=>p(158)(47),y=>p(159)(47),Cin=>p(160)(47),clock=>clock,reset=>reset,s=>p(234)(47),cout=>p(235)(48));
FA_ff_6693:FAff port map(x=>p(158)(48),y=>p(159)(48),Cin=>p(160)(48),clock=>clock,reset=>reset,s=>p(234)(48),cout=>p(235)(49));
FA_ff_6694:FAff port map(x=>p(158)(49),y=>p(159)(49),Cin=>p(160)(49),clock=>clock,reset=>reset,s=>p(234)(49),cout=>p(235)(50));
FA_ff_6695:FAff port map(x=>p(158)(50),y=>p(159)(50),Cin=>p(160)(50),clock=>clock,reset=>reset,s=>p(234)(50),cout=>p(235)(51));
FA_ff_6696:FAff port map(x=>p(158)(51),y=>p(159)(51),Cin=>p(160)(51),clock=>clock,reset=>reset,s=>p(234)(51),cout=>p(235)(52));
FA_ff_6697:FAff port map(x=>p(158)(52),y=>p(159)(52),Cin=>p(160)(52),clock=>clock,reset=>reset,s=>p(234)(52),cout=>p(235)(53));
FA_ff_6698:FAff port map(x=>p(158)(53),y=>p(159)(53),Cin=>p(160)(53),clock=>clock,reset=>reset,s=>p(234)(53),cout=>p(235)(54));
FA_ff_6699:FAff port map(x=>p(158)(54),y=>p(159)(54),Cin=>p(160)(54),clock=>clock,reset=>reset,s=>p(234)(54),cout=>p(235)(55));
FA_ff_6700:FAff port map(x=>p(158)(55),y=>p(159)(55),Cin=>p(160)(55),clock=>clock,reset=>reset,s=>p(234)(55),cout=>p(235)(56));
FA_ff_6701:FAff port map(x=>p(158)(56),y=>p(159)(56),Cin=>p(160)(56),clock=>clock,reset=>reset,s=>p(234)(56),cout=>p(235)(57));
FA_ff_6702:FAff port map(x=>p(158)(57),y=>p(159)(57),Cin=>p(160)(57),clock=>clock,reset=>reset,s=>p(234)(57),cout=>p(235)(58));
FA_ff_6703:FAff port map(x=>p(158)(58),y=>p(159)(58),Cin=>p(160)(58),clock=>clock,reset=>reset,s=>p(234)(58),cout=>p(235)(59));
FA_ff_6704:FAff port map(x=>p(158)(59),y=>p(159)(59),Cin=>p(160)(59),clock=>clock,reset=>reset,s=>p(234)(59),cout=>p(235)(60));
FA_ff_6705:FAff port map(x=>p(158)(60),y=>p(159)(60),Cin=>p(160)(60),clock=>clock,reset=>reset,s=>p(234)(60),cout=>p(235)(61));
FA_ff_6706:FAff port map(x=>p(158)(61),y=>p(159)(61),Cin=>p(160)(61),clock=>clock,reset=>reset,s=>p(234)(61),cout=>p(235)(62));
FA_ff_6707:FAff port map(x=>p(158)(62),y=>p(159)(62),Cin=>p(160)(62),clock=>clock,reset=>reset,s=>p(234)(62),cout=>p(235)(63));
FA_ff_6708:FAff port map(x=>p(158)(63),y=>p(159)(63),Cin=>p(160)(63),clock=>clock,reset=>reset,s=>p(234)(63),cout=>p(235)(64));
FA_ff_6709:FAff port map(x=>p(158)(64),y=>p(159)(64),Cin=>p(160)(64),clock=>clock,reset=>reset,s=>p(234)(64),cout=>p(235)(65));
FA_ff_6710:FAff port map(x=>p(158)(65),y=>p(159)(65),Cin=>p(160)(65),clock=>clock,reset=>reset,s=>p(234)(65),cout=>p(235)(66));
FA_ff_6711:FAff port map(x=>p(158)(66),y=>p(159)(66),Cin=>p(160)(66),clock=>clock,reset=>reset,s=>p(234)(66),cout=>p(235)(67));
FA_ff_6712:FAff port map(x=>p(158)(67),y=>p(159)(67),Cin=>p(160)(67),clock=>clock,reset=>reset,s=>p(234)(67),cout=>p(235)(68));
FA_ff_6713:FAff port map(x=>p(158)(68),y=>p(159)(68),Cin=>p(160)(68),clock=>clock,reset=>reset,s=>p(234)(68),cout=>p(235)(69));
FA_ff_6714:FAff port map(x=>p(158)(69),y=>p(159)(69),Cin=>p(160)(69),clock=>clock,reset=>reset,s=>p(234)(69),cout=>p(235)(70));
FA_ff_6715:FAff port map(x=>p(158)(70),y=>p(159)(70),Cin=>p(160)(70),clock=>clock,reset=>reset,s=>p(234)(70),cout=>p(235)(71));
FA_ff_6716:FAff port map(x=>p(158)(71),y=>p(159)(71),Cin=>p(160)(71),clock=>clock,reset=>reset,s=>p(234)(71),cout=>p(235)(72));
FA_ff_6717:FAff port map(x=>p(158)(72),y=>p(159)(72),Cin=>p(160)(72),clock=>clock,reset=>reset,s=>p(234)(72),cout=>p(235)(73));
FA_ff_6718:FAff port map(x=>p(158)(73),y=>p(159)(73),Cin=>p(160)(73),clock=>clock,reset=>reset,s=>p(234)(73),cout=>p(235)(74));
FA_ff_6719:FAff port map(x=>p(158)(74),y=>p(159)(74),Cin=>p(160)(74),clock=>clock,reset=>reset,s=>p(234)(74),cout=>p(235)(75));
FA_ff_6720:FAff port map(x=>p(158)(75),y=>p(159)(75),Cin=>p(160)(75),clock=>clock,reset=>reset,s=>p(234)(75),cout=>p(235)(76));
FA_ff_6721:FAff port map(x=>p(158)(76),y=>p(159)(76),Cin=>p(160)(76),clock=>clock,reset=>reset,s=>p(234)(76),cout=>p(235)(77));
FA_ff_6722:FAff port map(x=>p(158)(77),y=>p(159)(77),Cin=>p(160)(77),clock=>clock,reset=>reset,s=>p(234)(77),cout=>p(235)(78));
FA_ff_6723:FAff port map(x=>p(158)(78),y=>p(159)(78),Cin=>p(160)(78),clock=>clock,reset=>reset,s=>p(234)(78),cout=>p(235)(79));
FA_ff_6724:FAff port map(x=>p(158)(79),y=>p(159)(79),Cin=>p(160)(79),clock=>clock,reset=>reset,s=>p(234)(79),cout=>p(235)(80));
FA_ff_6725:FAff port map(x=>p(158)(80),y=>p(159)(80),Cin=>p(160)(80),clock=>clock,reset=>reset,s=>p(234)(80),cout=>p(235)(81));
FA_ff_6726:FAff port map(x=>p(158)(81),y=>p(159)(81),Cin=>p(160)(81),clock=>clock,reset=>reset,s=>p(234)(81),cout=>p(235)(82));
FA_ff_6727:FAff port map(x=>p(158)(82),y=>p(159)(82),Cin=>p(160)(82),clock=>clock,reset=>reset,s=>p(234)(82),cout=>p(235)(83));
FA_ff_6728:FAff port map(x=>p(158)(83),y=>p(159)(83),Cin=>p(160)(83),clock=>clock,reset=>reset,s=>p(234)(83),cout=>p(235)(84));
FA_ff_6729:FAff port map(x=>p(158)(84),y=>p(159)(84),Cin=>p(160)(84),clock=>clock,reset=>reset,s=>p(234)(84),cout=>p(235)(85));
FA_ff_6730:FAff port map(x=>p(158)(85),y=>p(159)(85),Cin=>p(160)(85),clock=>clock,reset=>reset,s=>p(234)(85),cout=>p(235)(86));
FA_ff_6731:FAff port map(x=>p(158)(86),y=>p(159)(86),Cin=>p(160)(86),clock=>clock,reset=>reset,s=>p(234)(86),cout=>p(235)(87));
FA_ff_6732:FAff port map(x=>p(158)(87),y=>p(159)(87),Cin=>p(160)(87),clock=>clock,reset=>reset,s=>p(234)(87),cout=>p(235)(88));
FA_ff_6733:FAff port map(x=>p(158)(88),y=>p(159)(88),Cin=>p(160)(88),clock=>clock,reset=>reset,s=>p(234)(88),cout=>p(235)(89));
FA_ff_6734:FAff port map(x=>p(158)(89),y=>p(159)(89),Cin=>p(160)(89),clock=>clock,reset=>reset,s=>p(234)(89),cout=>p(235)(90));
FA_ff_6735:FAff port map(x=>p(158)(90),y=>p(159)(90),Cin=>p(160)(90),clock=>clock,reset=>reset,s=>p(234)(90),cout=>p(235)(91));
FA_ff_6736:FAff port map(x=>p(158)(91),y=>p(159)(91),Cin=>p(160)(91),clock=>clock,reset=>reset,s=>p(234)(91),cout=>p(235)(92));
FA_ff_6737:FAff port map(x=>p(158)(92),y=>p(159)(92),Cin=>p(160)(92),clock=>clock,reset=>reset,s=>p(234)(92),cout=>p(235)(93));
FA_ff_6738:FAff port map(x=>p(158)(93),y=>p(159)(93),Cin=>p(160)(93),clock=>clock,reset=>reset,s=>p(234)(93),cout=>p(235)(94));
FA_ff_6739:FAff port map(x=>p(158)(94),y=>p(159)(94),Cin=>p(160)(94),clock=>clock,reset=>reset,s=>p(234)(94),cout=>p(235)(95));
FA_ff_6740:FAff port map(x=>p(158)(95),y=>p(159)(95),Cin=>p(160)(95),clock=>clock,reset=>reset,s=>p(234)(95),cout=>p(235)(96));
FA_ff_6741:FAff port map(x=>p(158)(96),y=>p(159)(96),Cin=>p(160)(96),clock=>clock,reset=>reset,s=>p(234)(96),cout=>p(235)(97));
FA_ff_6742:FAff port map(x=>p(158)(97),y=>p(159)(97),Cin=>p(160)(97),clock=>clock,reset=>reset,s=>p(234)(97),cout=>p(235)(98));
FA_ff_6743:FAff port map(x=>p(158)(98),y=>p(159)(98),Cin=>p(160)(98),clock=>clock,reset=>reset,s=>p(234)(98),cout=>p(235)(99));
FA_ff_6744:FAff port map(x=>p(158)(99),y=>p(159)(99),Cin=>p(160)(99),clock=>clock,reset=>reset,s=>p(234)(99),cout=>p(235)(100));
FA_ff_6745:FAff port map(x=>p(158)(100),y=>p(159)(100),Cin=>p(160)(100),clock=>clock,reset=>reset,s=>p(234)(100),cout=>p(235)(101));
FA_ff_6746:FAff port map(x=>p(158)(101),y=>p(159)(101),Cin=>p(160)(101),clock=>clock,reset=>reset,s=>p(234)(101),cout=>p(235)(102));
FA_ff_6747:FAff port map(x=>p(158)(102),y=>p(159)(102),Cin=>p(160)(102),clock=>clock,reset=>reset,s=>p(234)(102),cout=>p(235)(103));
FA_ff_6748:FAff port map(x=>p(158)(103),y=>p(159)(103),Cin=>p(160)(103),clock=>clock,reset=>reset,s=>p(234)(103),cout=>p(235)(104));
FA_ff_6749:FAff port map(x=>p(158)(104),y=>p(159)(104),Cin=>p(160)(104),clock=>clock,reset=>reset,s=>p(234)(104),cout=>p(235)(105));
FA_ff_6750:FAff port map(x=>p(158)(105),y=>p(159)(105),Cin=>p(160)(105),clock=>clock,reset=>reset,s=>p(234)(105),cout=>p(235)(106));
FA_ff_6751:FAff port map(x=>p(158)(106),y=>p(159)(106),Cin=>p(160)(106),clock=>clock,reset=>reset,s=>p(234)(106),cout=>p(235)(107));
FA_ff_6752:FAff port map(x=>p(158)(107),y=>p(159)(107),Cin=>p(160)(107),clock=>clock,reset=>reset,s=>p(234)(107),cout=>p(235)(108));
FA_ff_6753:FAff port map(x=>p(158)(108),y=>p(159)(108),Cin=>p(160)(108),clock=>clock,reset=>reset,s=>p(234)(108),cout=>p(235)(109));
FA_ff_6754:FAff port map(x=>p(158)(109),y=>p(159)(109),Cin=>p(160)(109),clock=>clock,reset=>reset,s=>p(234)(109),cout=>p(235)(110));
FA_ff_6755:FAff port map(x=>p(158)(110),y=>p(159)(110),Cin=>p(160)(110),clock=>clock,reset=>reset,s=>p(234)(110),cout=>p(235)(111));
FA_ff_6756:FAff port map(x=>p(158)(111),y=>p(159)(111),Cin=>p(160)(111),clock=>clock,reset=>reset,s=>p(234)(111),cout=>p(235)(112));
FA_ff_6757:FAff port map(x=>p(158)(112),y=>p(159)(112),Cin=>p(160)(112),clock=>clock,reset=>reset,s=>p(234)(112),cout=>p(235)(113));
FA_ff_6758:FAff port map(x=>p(158)(113),y=>p(159)(113),Cin=>p(160)(113),clock=>clock,reset=>reset,s=>p(234)(113),cout=>p(235)(114));
FA_ff_6759:FAff port map(x=>p(158)(114),y=>p(159)(114),Cin=>p(160)(114),clock=>clock,reset=>reset,s=>p(234)(114),cout=>p(235)(115));
FA_ff_6760:FAff port map(x=>p(158)(115),y=>p(159)(115),Cin=>p(160)(115),clock=>clock,reset=>reset,s=>p(234)(115),cout=>p(235)(116));
FA_ff_6761:FAff port map(x=>p(158)(116),y=>p(159)(116),Cin=>p(160)(116),clock=>clock,reset=>reset,s=>p(234)(116),cout=>p(235)(117));
FA_ff_6762:FAff port map(x=>p(158)(117),y=>p(159)(117),Cin=>p(160)(117),clock=>clock,reset=>reset,s=>p(234)(117),cout=>p(235)(118));
FA_ff_6763:FAff port map(x=>p(158)(118),y=>p(159)(118),Cin=>p(160)(118),clock=>clock,reset=>reset,s=>p(234)(118),cout=>p(235)(119));
FA_ff_6764:FAff port map(x=>p(158)(119),y=>p(159)(119),Cin=>p(160)(119),clock=>clock,reset=>reset,s=>p(234)(119),cout=>p(235)(120));
FA_ff_6765:FAff port map(x=>p(158)(120),y=>p(159)(120),Cin=>p(160)(120),clock=>clock,reset=>reset,s=>p(234)(120),cout=>p(235)(121));
FA_ff_6766:FAff port map(x=>p(158)(121),y=>p(159)(121),Cin=>p(160)(121),clock=>clock,reset=>reset,s=>p(234)(121),cout=>p(235)(122));
FA_ff_6767:FAff port map(x=>p(158)(122),y=>p(159)(122),Cin=>p(160)(122),clock=>clock,reset=>reset,s=>p(234)(122),cout=>p(235)(123));
FA_ff_6768:FAff port map(x=>p(158)(123),y=>p(159)(123),Cin=>p(160)(123),clock=>clock,reset=>reset,s=>p(234)(123),cout=>p(235)(124));
FA_ff_6769:FAff port map(x=>p(158)(124),y=>p(159)(124),Cin=>p(160)(124),clock=>clock,reset=>reset,s=>p(234)(124),cout=>p(235)(125));
FA_ff_6770:FAff port map(x=>p(158)(125),y=>p(159)(125),Cin=>p(160)(125),clock=>clock,reset=>reset,s=>p(234)(125),cout=>p(235)(126));
FA_ff_6771:FAff port map(x=>p(158)(126),y=>p(159)(126),Cin=>p(160)(126),clock=>clock,reset=>reset,s=>p(234)(126),cout=>p(235)(127));
FA_ff_6772:FAff port map(x=>p(158)(127),y=>p(159)(127),Cin=>p(160)(127),clock=>clock,reset=>reset,s=>p(234)(127),cout=>p(235)(128));
p(234)(128)<=p(159)(128);
p(236)(0)<=p(162)(0);
FA_ff_6773:FAff port map(x=>p(161)(1),y=>p(162)(1),Cin=>p(163)(1),clock=>clock,reset=>reset,s=>p(236)(1),cout=>p(237)(2));
FA_ff_6774:FAff port map(x=>p(161)(2),y=>p(162)(2),Cin=>p(163)(2),clock=>clock,reset=>reset,s=>p(236)(2),cout=>p(237)(3));
FA_ff_6775:FAff port map(x=>p(161)(3),y=>p(162)(3),Cin=>p(163)(3),clock=>clock,reset=>reset,s=>p(236)(3),cout=>p(237)(4));
FA_ff_6776:FAff port map(x=>p(161)(4),y=>p(162)(4),Cin=>p(163)(4),clock=>clock,reset=>reset,s=>p(236)(4),cout=>p(237)(5));
FA_ff_6777:FAff port map(x=>p(161)(5),y=>p(162)(5),Cin=>p(163)(5),clock=>clock,reset=>reset,s=>p(236)(5),cout=>p(237)(6));
FA_ff_6778:FAff port map(x=>p(161)(6),y=>p(162)(6),Cin=>p(163)(6),clock=>clock,reset=>reset,s=>p(236)(6),cout=>p(237)(7));
FA_ff_6779:FAff port map(x=>p(161)(7),y=>p(162)(7),Cin=>p(163)(7),clock=>clock,reset=>reset,s=>p(236)(7),cout=>p(237)(8));
FA_ff_6780:FAff port map(x=>p(161)(8),y=>p(162)(8),Cin=>p(163)(8),clock=>clock,reset=>reset,s=>p(236)(8),cout=>p(237)(9));
FA_ff_6781:FAff port map(x=>p(161)(9),y=>p(162)(9),Cin=>p(163)(9),clock=>clock,reset=>reset,s=>p(236)(9),cout=>p(237)(10));
FA_ff_6782:FAff port map(x=>p(161)(10),y=>p(162)(10),Cin=>p(163)(10),clock=>clock,reset=>reset,s=>p(236)(10),cout=>p(237)(11));
FA_ff_6783:FAff port map(x=>p(161)(11),y=>p(162)(11),Cin=>p(163)(11),clock=>clock,reset=>reset,s=>p(236)(11),cout=>p(237)(12));
FA_ff_6784:FAff port map(x=>p(161)(12),y=>p(162)(12),Cin=>p(163)(12),clock=>clock,reset=>reset,s=>p(236)(12),cout=>p(237)(13));
FA_ff_6785:FAff port map(x=>p(161)(13),y=>p(162)(13),Cin=>p(163)(13),clock=>clock,reset=>reset,s=>p(236)(13),cout=>p(237)(14));
FA_ff_6786:FAff port map(x=>p(161)(14),y=>p(162)(14),Cin=>p(163)(14),clock=>clock,reset=>reset,s=>p(236)(14),cout=>p(237)(15));
FA_ff_6787:FAff port map(x=>p(161)(15),y=>p(162)(15),Cin=>p(163)(15),clock=>clock,reset=>reset,s=>p(236)(15),cout=>p(237)(16));
FA_ff_6788:FAff port map(x=>p(161)(16),y=>p(162)(16),Cin=>p(163)(16),clock=>clock,reset=>reset,s=>p(236)(16),cout=>p(237)(17));
FA_ff_6789:FAff port map(x=>p(161)(17),y=>p(162)(17),Cin=>p(163)(17),clock=>clock,reset=>reset,s=>p(236)(17),cout=>p(237)(18));
FA_ff_6790:FAff port map(x=>p(161)(18),y=>p(162)(18),Cin=>p(163)(18),clock=>clock,reset=>reset,s=>p(236)(18),cout=>p(237)(19));
FA_ff_6791:FAff port map(x=>p(161)(19),y=>p(162)(19),Cin=>p(163)(19),clock=>clock,reset=>reset,s=>p(236)(19),cout=>p(237)(20));
FA_ff_6792:FAff port map(x=>p(161)(20),y=>p(162)(20),Cin=>p(163)(20),clock=>clock,reset=>reset,s=>p(236)(20),cout=>p(237)(21));
FA_ff_6793:FAff port map(x=>p(161)(21),y=>p(162)(21),Cin=>p(163)(21),clock=>clock,reset=>reset,s=>p(236)(21),cout=>p(237)(22));
FA_ff_6794:FAff port map(x=>p(161)(22),y=>p(162)(22),Cin=>p(163)(22),clock=>clock,reset=>reset,s=>p(236)(22),cout=>p(237)(23));
FA_ff_6795:FAff port map(x=>p(161)(23),y=>p(162)(23),Cin=>p(163)(23),clock=>clock,reset=>reset,s=>p(236)(23),cout=>p(237)(24));
FA_ff_6796:FAff port map(x=>p(161)(24),y=>p(162)(24),Cin=>p(163)(24),clock=>clock,reset=>reset,s=>p(236)(24),cout=>p(237)(25));
FA_ff_6797:FAff port map(x=>p(161)(25),y=>p(162)(25),Cin=>p(163)(25),clock=>clock,reset=>reset,s=>p(236)(25),cout=>p(237)(26));
FA_ff_6798:FAff port map(x=>p(161)(26),y=>p(162)(26),Cin=>p(163)(26),clock=>clock,reset=>reset,s=>p(236)(26),cout=>p(237)(27));
FA_ff_6799:FAff port map(x=>p(161)(27),y=>p(162)(27),Cin=>p(163)(27),clock=>clock,reset=>reset,s=>p(236)(27),cout=>p(237)(28));
FA_ff_6800:FAff port map(x=>p(161)(28),y=>p(162)(28),Cin=>p(163)(28),clock=>clock,reset=>reset,s=>p(236)(28),cout=>p(237)(29));
FA_ff_6801:FAff port map(x=>p(161)(29),y=>p(162)(29),Cin=>p(163)(29),clock=>clock,reset=>reset,s=>p(236)(29),cout=>p(237)(30));
FA_ff_6802:FAff port map(x=>p(161)(30),y=>p(162)(30),Cin=>p(163)(30),clock=>clock,reset=>reset,s=>p(236)(30),cout=>p(237)(31));
FA_ff_6803:FAff port map(x=>p(161)(31),y=>p(162)(31),Cin=>p(163)(31),clock=>clock,reset=>reset,s=>p(236)(31),cout=>p(237)(32));
FA_ff_6804:FAff port map(x=>p(161)(32),y=>p(162)(32),Cin=>p(163)(32),clock=>clock,reset=>reset,s=>p(236)(32),cout=>p(237)(33));
FA_ff_6805:FAff port map(x=>p(161)(33),y=>p(162)(33),Cin=>p(163)(33),clock=>clock,reset=>reset,s=>p(236)(33),cout=>p(237)(34));
FA_ff_6806:FAff port map(x=>p(161)(34),y=>p(162)(34),Cin=>p(163)(34),clock=>clock,reset=>reset,s=>p(236)(34),cout=>p(237)(35));
FA_ff_6807:FAff port map(x=>p(161)(35),y=>p(162)(35),Cin=>p(163)(35),clock=>clock,reset=>reset,s=>p(236)(35),cout=>p(237)(36));
FA_ff_6808:FAff port map(x=>p(161)(36),y=>p(162)(36),Cin=>p(163)(36),clock=>clock,reset=>reset,s=>p(236)(36),cout=>p(237)(37));
FA_ff_6809:FAff port map(x=>p(161)(37),y=>p(162)(37),Cin=>p(163)(37),clock=>clock,reset=>reset,s=>p(236)(37),cout=>p(237)(38));
FA_ff_6810:FAff port map(x=>p(161)(38),y=>p(162)(38),Cin=>p(163)(38),clock=>clock,reset=>reset,s=>p(236)(38),cout=>p(237)(39));
FA_ff_6811:FAff port map(x=>p(161)(39),y=>p(162)(39),Cin=>p(163)(39),clock=>clock,reset=>reset,s=>p(236)(39),cout=>p(237)(40));
FA_ff_6812:FAff port map(x=>p(161)(40),y=>p(162)(40),Cin=>p(163)(40),clock=>clock,reset=>reset,s=>p(236)(40),cout=>p(237)(41));
FA_ff_6813:FAff port map(x=>p(161)(41),y=>p(162)(41),Cin=>p(163)(41),clock=>clock,reset=>reset,s=>p(236)(41),cout=>p(237)(42));
FA_ff_6814:FAff port map(x=>p(161)(42),y=>p(162)(42),Cin=>p(163)(42),clock=>clock,reset=>reset,s=>p(236)(42),cout=>p(237)(43));
FA_ff_6815:FAff port map(x=>p(161)(43),y=>p(162)(43),Cin=>p(163)(43),clock=>clock,reset=>reset,s=>p(236)(43),cout=>p(237)(44));
FA_ff_6816:FAff port map(x=>p(161)(44),y=>p(162)(44),Cin=>p(163)(44),clock=>clock,reset=>reset,s=>p(236)(44),cout=>p(237)(45));
FA_ff_6817:FAff port map(x=>p(161)(45),y=>p(162)(45),Cin=>p(163)(45),clock=>clock,reset=>reset,s=>p(236)(45),cout=>p(237)(46));
FA_ff_6818:FAff port map(x=>p(161)(46),y=>p(162)(46),Cin=>p(163)(46),clock=>clock,reset=>reset,s=>p(236)(46),cout=>p(237)(47));
FA_ff_6819:FAff port map(x=>p(161)(47),y=>p(162)(47),Cin=>p(163)(47),clock=>clock,reset=>reset,s=>p(236)(47),cout=>p(237)(48));
FA_ff_6820:FAff port map(x=>p(161)(48),y=>p(162)(48),Cin=>p(163)(48),clock=>clock,reset=>reset,s=>p(236)(48),cout=>p(237)(49));
FA_ff_6821:FAff port map(x=>p(161)(49),y=>p(162)(49),Cin=>p(163)(49),clock=>clock,reset=>reset,s=>p(236)(49),cout=>p(237)(50));
FA_ff_6822:FAff port map(x=>p(161)(50),y=>p(162)(50),Cin=>p(163)(50),clock=>clock,reset=>reset,s=>p(236)(50),cout=>p(237)(51));
FA_ff_6823:FAff port map(x=>p(161)(51),y=>p(162)(51),Cin=>p(163)(51),clock=>clock,reset=>reset,s=>p(236)(51),cout=>p(237)(52));
FA_ff_6824:FAff port map(x=>p(161)(52),y=>p(162)(52),Cin=>p(163)(52),clock=>clock,reset=>reset,s=>p(236)(52),cout=>p(237)(53));
FA_ff_6825:FAff port map(x=>p(161)(53),y=>p(162)(53),Cin=>p(163)(53),clock=>clock,reset=>reset,s=>p(236)(53),cout=>p(237)(54));
FA_ff_6826:FAff port map(x=>p(161)(54),y=>p(162)(54),Cin=>p(163)(54),clock=>clock,reset=>reset,s=>p(236)(54),cout=>p(237)(55));
FA_ff_6827:FAff port map(x=>p(161)(55),y=>p(162)(55),Cin=>p(163)(55),clock=>clock,reset=>reset,s=>p(236)(55),cout=>p(237)(56));
FA_ff_6828:FAff port map(x=>p(161)(56),y=>p(162)(56),Cin=>p(163)(56),clock=>clock,reset=>reset,s=>p(236)(56),cout=>p(237)(57));
FA_ff_6829:FAff port map(x=>p(161)(57),y=>p(162)(57),Cin=>p(163)(57),clock=>clock,reset=>reset,s=>p(236)(57),cout=>p(237)(58));
FA_ff_6830:FAff port map(x=>p(161)(58),y=>p(162)(58),Cin=>p(163)(58),clock=>clock,reset=>reset,s=>p(236)(58),cout=>p(237)(59));
FA_ff_6831:FAff port map(x=>p(161)(59),y=>p(162)(59),Cin=>p(163)(59),clock=>clock,reset=>reset,s=>p(236)(59),cout=>p(237)(60));
FA_ff_6832:FAff port map(x=>p(161)(60),y=>p(162)(60),Cin=>p(163)(60),clock=>clock,reset=>reset,s=>p(236)(60),cout=>p(237)(61));
FA_ff_6833:FAff port map(x=>p(161)(61),y=>p(162)(61),Cin=>p(163)(61),clock=>clock,reset=>reset,s=>p(236)(61),cout=>p(237)(62));
FA_ff_6834:FAff port map(x=>p(161)(62),y=>p(162)(62),Cin=>p(163)(62),clock=>clock,reset=>reset,s=>p(236)(62),cout=>p(237)(63));
FA_ff_6835:FAff port map(x=>p(161)(63),y=>p(162)(63),Cin=>p(163)(63),clock=>clock,reset=>reset,s=>p(236)(63),cout=>p(237)(64));
FA_ff_6836:FAff port map(x=>p(161)(64),y=>p(162)(64),Cin=>p(163)(64),clock=>clock,reset=>reset,s=>p(236)(64),cout=>p(237)(65));
FA_ff_6837:FAff port map(x=>p(161)(65),y=>p(162)(65),Cin=>p(163)(65),clock=>clock,reset=>reset,s=>p(236)(65),cout=>p(237)(66));
FA_ff_6838:FAff port map(x=>p(161)(66),y=>p(162)(66),Cin=>p(163)(66),clock=>clock,reset=>reset,s=>p(236)(66),cout=>p(237)(67));
FA_ff_6839:FAff port map(x=>p(161)(67),y=>p(162)(67),Cin=>p(163)(67),clock=>clock,reset=>reset,s=>p(236)(67),cout=>p(237)(68));
FA_ff_6840:FAff port map(x=>p(161)(68),y=>p(162)(68),Cin=>p(163)(68),clock=>clock,reset=>reset,s=>p(236)(68),cout=>p(237)(69));
FA_ff_6841:FAff port map(x=>p(161)(69),y=>p(162)(69),Cin=>p(163)(69),clock=>clock,reset=>reset,s=>p(236)(69),cout=>p(237)(70));
FA_ff_6842:FAff port map(x=>p(161)(70),y=>p(162)(70),Cin=>p(163)(70),clock=>clock,reset=>reset,s=>p(236)(70),cout=>p(237)(71));
FA_ff_6843:FAff port map(x=>p(161)(71),y=>p(162)(71),Cin=>p(163)(71),clock=>clock,reset=>reset,s=>p(236)(71),cout=>p(237)(72));
FA_ff_6844:FAff port map(x=>p(161)(72),y=>p(162)(72),Cin=>p(163)(72),clock=>clock,reset=>reset,s=>p(236)(72),cout=>p(237)(73));
FA_ff_6845:FAff port map(x=>p(161)(73),y=>p(162)(73),Cin=>p(163)(73),clock=>clock,reset=>reset,s=>p(236)(73),cout=>p(237)(74));
FA_ff_6846:FAff port map(x=>p(161)(74),y=>p(162)(74),Cin=>p(163)(74),clock=>clock,reset=>reset,s=>p(236)(74),cout=>p(237)(75));
FA_ff_6847:FAff port map(x=>p(161)(75),y=>p(162)(75),Cin=>p(163)(75),clock=>clock,reset=>reset,s=>p(236)(75),cout=>p(237)(76));
FA_ff_6848:FAff port map(x=>p(161)(76),y=>p(162)(76),Cin=>p(163)(76),clock=>clock,reset=>reset,s=>p(236)(76),cout=>p(237)(77));
FA_ff_6849:FAff port map(x=>p(161)(77),y=>p(162)(77),Cin=>p(163)(77),clock=>clock,reset=>reset,s=>p(236)(77),cout=>p(237)(78));
FA_ff_6850:FAff port map(x=>p(161)(78),y=>p(162)(78),Cin=>p(163)(78),clock=>clock,reset=>reset,s=>p(236)(78),cout=>p(237)(79));
FA_ff_6851:FAff port map(x=>p(161)(79),y=>p(162)(79),Cin=>p(163)(79),clock=>clock,reset=>reset,s=>p(236)(79),cout=>p(237)(80));
FA_ff_6852:FAff port map(x=>p(161)(80),y=>p(162)(80),Cin=>p(163)(80),clock=>clock,reset=>reset,s=>p(236)(80),cout=>p(237)(81));
FA_ff_6853:FAff port map(x=>p(161)(81),y=>p(162)(81),Cin=>p(163)(81),clock=>clock,reset=>reset,s=>p(236)(81),cout=>p(237)(82));
FA_ff_6854:FAff port map(x=>p(161)(82),y=>p(162)(82),Cin=>p(163)(82),clock=>clock,reset=>reset,s=>p(236)(82),cout=>p(237)(83));
FA_ff_6855:FAff port map(x=>p(161)(83),y=>p(162)(83),Cin=>p(163)(83),clock=>clock,reset=>reset,s=>p(236)(83),cout=>p(237)(84));
FA_ff_6856:FAff port map(x=>p(161)(84),y=>p(162)(84),Cin=>p(163)(84),clock=>clock,reset=>reset,s=>p(236)(84),cout=>p(237)(85));
FA_ff_6857:FAff port map(x=>p(161)(85),y=>p(162)(85),Cin=>p(163)(85),clock=>clock,reset=>reset,s=>p(236)(85),cout=>p(237)(86));
FA_ff_6858:FAff port map(x=>p(161)(86),y=>p(162)(86),Cin=>p(163)(86),clock=>clock,reset=>reset,s=>p(236)(86),cout=>p(237)(87));
FA_ff_6859:FAff port map(x=>p(161)(87),y=>p(162)(87),Cin=>p(163)(87),clock=>clock,reset=>reset,s=>p(236)(87),cout=>p(237)(88));
FA_ff_6860:FAff port map(x=>p(161)(88),y=>p(162)(88),Cin=>p(163)(88),clock=>clock,reset=>reset,s=>p(236)(88),cout=>p(237)(89));
FA_ff_6861:FAff port map(x=>p(161)(89),y=>p(162)(89),Cin=>p(163)(89),clock=>clock,reset=>reset,s=>p(236)(89),cout=>p(237)(90));
FA_ff_6862:FAff port map(x=>p(161)(90),y=>p(162)(90),Cin=>p(163)(90),clock=>clock,reset=>reset,s=>p(236)(90),cout=>p(237)(91));
FA_ff_6863:FAff port map(x=>p(161)(91),y=>p(162)(91),Cin=>p(163)(91),clock=>clock,reset=>reset,s=>p(236)(91),cout=>p(237)(92));
FA_ff_6864:FAff port map(x=>p(161)(92),y=>p(162)(92),Cin=>p(163)(92),clock=>clock,reset=>reset,s=>p(236)(92),cout=>p(237)(93));
FA_ff_6865:FAff port map(x=>p(161)(93),y=>p(162)(93),Cin=>p(163)(93),clock=>clock,reset=>reset,s=>p(236)(93),cout=>p(237)(94));
FA_ff_6866:FAff port map(x=>p(161)(94),y=>p(162)(94),Cin=>p(163)(94),clock=>clock,reset=>reset,s=>p(236)(94),cout=>p(237)(95));
FA_ff_6867:FAff port map(x=>p(161)(95),y=>p(162)(95),Cin=>p(163)(95),clock=>clock,reset=>reset,s=>p(236)(95),cout=>p(237)(96));
FA_ff_6868:FAff port map(x=>p(161)(96),y=>p(162)(96),Cin=>p(163)(96),clock=>clock,reset=>reset,s=>p(236)(96),cout=>p(237)(97));
FA_ff_6869:FAff port map(x=>p(161)(97),y=>p(162)(97),Cin=>p(163)(97),clock=>clock,reset=>reset,s=>p(236)(97),cout=>p(237)(98));
FA_ff_6870:FAff port map(x=>p(161)(98),y=>p(162)(98),Cin=>p(163)(98),clock=>clock,reset=>reset,s=>p(236)(98),cout=>p(237)(99));
FA_ff_6871:FAff port map(x=>p(161)(99),y=>p(162)(99),Cin=>p(163)(99),clock=>clock,reset=>reset,s=>p(236)(99),cout=>p(237)(100));
FA_ff_6872:FAff port map(x=>p(161)(100),y=>p(162)(100),Cin=>p(163)(100),clock=>clock,reset=>reset,s=>p(236)(100),cout=>p(237)(101));
FA_ff_6873:FAff port map(x=>p(161)(101),y=>p(162)(101),Cin=>p(163)(101),clock=>clock,reset=>reset,s=>p(236)(101),cout=>p(237)(102));
FA_ff_6874:FAff port map(x=>p(161)(102),y=>p(162)(102),Cin=>p(163)(102),clock=>clock,reset=>reset,s=>p(236)(102),cout=>p(237)(103));
FA_ff_6875:FAff port map(x=>p(161)(103),y=>p(162)(103),Cin=>p(163)(103),clock=>clock,reset=>reset,s=>p(236)(103),cout=>p(237)(104));
FA_ff_6876:FAff port map(x=>p(161)(104),y=>p(162)(104),Cin=>p(163)(104),clock=>clock,reset=>reset,s=>p(236)(104),cout=>p(237)(105));
FA_ff_6877:FAff port map(x=>p(161)(105),y=>p(162)(105),Cin=>p(163)(105),clock=>clock,reset=>reset,s=>p(236)(105),cout=>p(237)(106));
FA_ff_6878:FAff port map(x=>p(161)(106),y=>p(162)(106),Cin=>p(163)(106),clock=>clock,reset=>reset,s=>p(236)(106),cout=>p(237)(107));
FA_ff_6879:FAff port map(x=>p(161)(107),y=>p(162)(107),Cin=>p(163)(107),clock=>clock,reset=>reset,s=>p(236)(107),cout=>p(237)(108));
FA_ff_6880:FAff port map(x=>p(161)(108),y=>p(162)(108),Cin=>p(163)(108),clock=>clock,reset=>reset,s=>p(236)(108),cout=>p(237)(109));
FA_ff_6881:FAff port map(x=>p(161)(109),y=>p(162)(109),Cin=>p(163)(109),clock=>clock,reset=>reset,s=>p(236)(109),cout=>p(237)(110));
FA_ff_6882:FAff port map(x=>p(161)(110),y=>p(162)(110),Cin=>p(163)(110),clock=>clock,reset=>reset,s=>p(236)(110),cout=>p(237)(111));
FA_ff_6883:FAff port map(x=>p(161)(111),y=>p(162)(111),Cin=>p(163)(111),clock=>clock,reset=>reset,s=>p(236)(111),cout=>p(237)(112));
FA_ff_6884:FAff port map(x=>p(161)(112),y=>p(162)(112),Cin=>p(163)(112),clock=>clock,reset=>reset,s=>p(236)(112),cout=>p(237)(113));
FA_ff_6885:FAff port map(x=>p(161)(113),y=>p(162)(113),Cin=>p(163)(113),clock=>clock,reset=>reset,s=>p(236)(113),cout=>p(237)(114));
FA_ff_6886:FAff port map(x=>p(161)(114),y=>p(162)(114),Cin=>p(163)(114),clock=>clock,reset=>reset,s=>p(236)(114),cout=>p(237)(115));
FA_ff_6887:FAff port map(x=>p(161)(115),y=>p(162)(115),Cin=>p(163)(115),clock=>clock,reset=>reset,s=>p(236)(115),cout=>p(237)(116));
FA_ff_6888:FAff port map(x=>p(161)(116),y=>p(162)(116),Cin=>p(163)(116),clock=>clock,reset=>reset,s=>p(236)(116),cout=>p(237)(117));
FA_ff_6889:FAff port map(x=>p(161)(117),y=>p(162)(117),Cin=>p(163)(117),clock=>clock,reset=>reset,s=>p(236)(117),cout=>p(237)(118));
FA_ff_6890:FAff port map(x=>p(161)(118),y=>p(162)(118),Cin=>p(163)(118),clock=>clock,reset=>reset,s=>p(236)(118),cout=>p(237)(119));
FA_ff_6891:FAff port map(x=>p(161)(119),y=>p(162)(119),Cin=>p(163)(119),clock=>clock,reset=>reset,s=>p(236)(119),cout=>p(237)(120));
FA_ff_6892:FAff port map(x=>p(161)(120),y=>p(162)(120),Cin=>p(163)(120),clock=>clock,reset=>reset,s=>p(236)(120),cout=>p(237)(121));
FA_ff_6893:FAff port map(x=>p(161)(121),y=>p(162)(121),Cin=>p(163)(121),clock=>clock,reset=>reset,s=>p(236)(121),cout=>p(237)(122));
FA_ff_6894:FAff port map(x=>p(161)(122),y=>p(162)(122),Cin=>p(163)(122),clock=>clock,reset=>reset,s=>p(236)(122),cout=>p(237)(123));
FA_ff_6895:FAff port map(x=>p(161)(123),y=>p(162)(123),Cin=>p(163)(123),clock=>clock,reset=>reset,s=>p(236)(123),cout=>p(237)(124));
FA_ff_6896:FAff port map(x=>p(161)(124),y=>p(162)(124),Cin=>p(163)(124),clock=>clock,reset=>reset,s=>p(236)(124),cout=>p(237)(125));
FA_ff_6897:FAff port map(x=>p(161)(125),y=>p(162)(125),Cin=>p(163)(125),clock=>clock,reset=>reset,s=>p(236)(125),cout=>p(237)(126));
FA_ff_6898:FAff port map(x=>p(161)(126),y=>p(162)(126),Cin=>p(163)(126),clock=>clock,reset=>reset,s=>p(236)(126),cout=>p(237)(127));
FA_ff_6899:FAff port map(x=>p(161)(127),y=>p(162)(127),Cin=>p(163)(127),clock=>clock,reset=>reset,s=>p(236)(127),cout=>p(237)(128));
HA_ff_11:HAff port map(x=>p(161)(128),y=>p(163)(128),clock=>clock,reset=>reset,s=>p(236)(128),c=>p(237)(129));
HA_ff_12:HAff port map(x=>p(164)(0),y=>p(166)(0),clock=>clock,reset=>reset,s=>p(238)(0),c=>p(239)(1));
FA_ff_6900:FAff port map(x=>p(164)(1),y=>p(165)(1),Cin=>p(166)(1),clock=>clock,reset=>reset,s=>p(238)(1),cout=>p(239)(2));
FA_ff_6901:FAff port map(x=>p(164)(2),y=>p(165)(2),Cin=>p(166)(2),clock=>clock,reset=>reset,s=>p(238)(2),cout=>p(239)(3));
FA_ff_6902:FAff port map(x=>p(164)(3),y=>p(165)(3),Cin=>p(166)(3),clock=>clock,reset=>reset,s=>p(238)(3),cout=>p(239)(4));
FA_ff_6903:FAff port map(x=>p(164)(4),y=>p(165)(4),Cin=>p(166)(4),clock=>clock,reset=>reset,s=>p(238)(4),cout=>p(239)(5));
FA_ff_6904:FAff port map(x=>p(164)(5),y=>p(165)(5),Cin=>p(166)(5),clock=>clock,reset=>reset,s=>p(238)(5),cout=>p(239)(6));
FA_ff_6905:FAff port map(x=>p(164)(6),y=>p(165)(6),Cin=>p(166)(6),clock=>clock,reset=>reset,s=>p(238)(6),cout=>p(239)(7));
FA_ff_6906:FAff port map(x=>p(164)(7),y=>p(165)(7),Cin=>p(166)(7),clock=>clock,reset=>reset,s=>p(238)(7),cout=>p(239)(8));
FA_ff_6907:FAff port map(x=>p(164)(8),y=>p(165)(8),Cin=>p(166)(8),clock=>clock,reset=>reset,s=>p(238)(8),cout=>p(239)(9));
FA_ff_6908:FAff port map(x=>p(164)(9),y=>p(165)(9),Cin=>p(166)(9),clock=>clock,reset=>reset,s=>p(238)(9),cout=>p(239)(10));
FA_ff_6909:FAff port map(x=>p(164)(10),y=>p(165)(10),Cin=>p(166)(10),clock=>clock,reset=>reset,s=>p(238)(10),cout=>p(239)(11));
FA_ff_6910:FAff port map(x=>p(164)(11),y=>p(165)(11),Cin=>p(166)(11),clock=>clock,reset=>reset,s=>p(238)(11),cout=>p(239)(12));
FA_ff_6911:FAff port map(x=>p(164)(12),y=>p(165)(12),Cin=>p(166)(12),clock=>clock,reset=>reset,s=>p(238)(12),cout=>p(239)(13));
FA_ff_6912:FAff port map(x=>p(164)(13),y=>p(165)(13),Cin=>p(166)(13),clock=>clock,reset=>reset,s=>p(238)(13),cout=>p(239)(14));
FA_ff_6913:FAff port map(x=>p(164)(14),y=>p(165)(14),Cin=>p(166)(14),clock=>clock,reset=>reset,s=>p(238)(14),cout=>p(239)(15));
FA_ff_6914:FAff port map(x=>p(164)(15),y=>p(165)(15),Cin=>p(166)(15),clock=>clock,reset=>reset,s=>p(238)(15),cout=>p(239)(16));
FA_ff_6915:FAff port map(x=>p(164)(16),y=>p(165)(16),Cin=>p(166)(16),clock=>clock,reset=>reset,s=>p(238)(16),cout=>p(239)(17));
FA_ff_6916:FAff port map(x=>p(164)(17),y=>p(165)(17),Cin=>p(166)(17),clock=>clock,reset=>reset,s=>p(238)(17),cout=>p(239)(18));
FA_ff_6917:FAff port map(x=>p(164)(18),y=>p(165)(18),Cin=>p(166)(18),clock=>clock,reset=>reset,s=>p(238)(18),cout=>p(239)(19));
FA_ff_6918:FAff port map(x=>p(164)(19),y=>p(165)(19),Cin=>p(166)(19),clock=>clock,reset=>reset,s=>p(238)(19),cout=>p(239)(20));
FA_ff_6919:FAff port map(x=>p(164)(20),y=>p(165)(20),Cin=>p(166)(20),clock=>clock,reset=>reset,s=>p(238)(20),cout=>p(239)(21));
FA_ff_6920:FAff port map(x=>p(164)(21),y=>p(165)(21),Cin=>p(166)(21),clock=>clock,reset=>reset,s=>p(238)(21),cout=>p(239)(22));
FA_ff_6921:FAff port map(x=>p(164)(22),y=>p(165)(22),Cin=>p(166)(22),clock=>clock,reset=>reset,s=>p(238)(22),cout=>p(239)(23));
FA_ff_6922:FAff port map(x=>p(164)(23),y=>p(165)(23),Cin=>p(166)(23),clock=>clock,reset=>reset,s=>p(238)(23),cout=>p(239)(24));
FA_ff_6923:FAff port map(x=>p(164)(24),y=>p(165)(24),Cin=>p(166)(24),clock=>clock,reset=>reset,s=>p(238)(24),cout=>p(239)(25));
FA_ff_6924:FAff port map(x=>p(164)(25),y=>p(165)(25),Cin=>p(166)(25),clock=>clock,reset=>reset,s=>p(238)(25),cout=>p(239)(26));
FA_ff_6925:FAff port map(x=>p(164)(26),y=>p(165)(26),Cin=>p(166)(26),clock=>clock,reset=>reset,s=>p(238)(26),cout=>p(239)(27));
FA_ff_6926:FAff port map(x=>p(164)(27),y=>p(165)(27),Cin=>p(166)(27),clock=>clock,reset=>reset,s=>p(238)(27),cout=>p(239)(28));
FA_ff_6927:FAff port map(x=>p(164)(28),y=>p(165)(28),Cin=>p(166)(28),clock=>clock,reset=>reset,s=>p(238)(28),cout=>p(239)(29));
FA_ff_6928:FAff port map(x=>p(164)(29),y=>p(165)(29),Cin=>p(166)(29),clock=>clock,reset=>reset,s=>p(238)(29),cout=>p(239)(30));
FA_ff_6929:FAff port map(x=>p(164)(30),y=>p(165)(30),Cin=>p(166)(30),clock=>clock,reset=>reset,s=>p(238)(30),cout=>p(239)(31));
FA_ff_6930:FAff port map(x=>p(164)(31),y=>p(165)(31),Cin=>p(166)(31),clock=>clock,reset=>reset,s=>p(238)(31),cout=>p(239)(32));
FA_ff_6931:FAff port map(x=>p(164)(32),y=>p(165)(32),Cin=>p(166)(32),clock=>clock,reset=>reset,s=>p(238)(32),cout=>p(239)(33));
FA_ff_6932:FAff port map(x=>p(164)(33),y=>p(165)(33),Cin=>p(166)(33),clock=>clock,reset=>reset,s=>p(238)(33),cout=>p(239)(34));
FA_ff_6933:FAff port map(x=>p(164)(34),y=>p(165)(34),Cin=>p(166)(34),clock=>clock,reset=>reset,s=>p(238)(34),cout=>p(239)(35));
FA_ff_6934:FAff port map(x=>p(164)(35),y=>p(165)(35),Cin=>p(166)(35),clock=>clock,reset=>reset,s=>p(238)(35),cout=>p(239)(36));
FA_ff_6935:FAff port map(x=>p(164)(36),y=>p(165)(36),Cin=>p(166)(36),clock=>clock,reset=>reset,s=>p(238)(36),cout=>p(239)(37));
FA_ff_6936:FAff port map(x=>p(164)(37),y=>p(165)(37),Cin=>p(166)(37),clock=>clock,reset=>reset,s=>p(238)(37),cout=>p(239)(38));
FA_ff_6937:FAff port map(x=>p(164)(38),y=>p(165)(38),Cin=>p(166)(38),clock=>clock,reset=>reset,s=>p(238)(38),cout=>p(239)(39));
FA_ff_6938:FAff port map(x=>p(164)(39),y=>p(165)(39),Cin=>p(166)(39),clock=>clock,reset=>reset,s=>p(238)(39),cout=>p(239)(40));
FA_ff_6939:FAff port map(x=>p(164)(40),y=>p(165)(40),Cin=>p(166)(40),clock=>clock,reset=>reset,s=>p(238)(40),cout=>p(239)(41));
FA_ff_6940:FAff port map(x=>p(164)(41),y=>p(165)(41),Cin=>p(166)(41),clock=>clock,reset=>reset,s=>p(238)(41),cout=>p(239)(42));
FA_ff_6941:FAff port map(x=>p(164)(42),y=>p(165)(42),Cin=>p(166)(42),clock=>clock,reset=>reset,s=>p(238)(42),cout=>p(239)(43));
FA_ff_6942:FAff port map(x=>p(164)(43),y=>p(165)(43),Cin=>p(166)(43),clock=>clock,reset=>reset,s=>p(238)(43),cout=>p(239)(44));
FA_ff_6943:FAff port map(x=>p(164)(44),y=>p(165)(44),Cin=>p(166)(44),clock=>clock,reset=>reset,s=>p(238)(44),cout=>p(239)(45));
FA_ff_6944:FAff port map(x=>p(164)(45),y=>p(165)(45),Cin=>p(166)(45),clock=>clock,reset=>reset,s=>p(238)(45),cout=>p(239)(46));
FA_ff_6945:FAff port map(x=>p(164)(46),y=>p(165)(46),Cin=>p(166)(46),clock=>clock,reset=>reset,s=>p(238)(46),cout=>p(239)(47));
FA_ff_6946:FAff port map(x=>p(164)(47),y=>p(165)(47),Cin=>p(166)(47),clock=>clock,reset=>reset,s=>p(238)(47),cout=>p(239)(48));
FA_ff_6947:FAff port map(x=>p(164)(48),y=>p(165)(48),Cin=>p(166)(48),clock=>clock,reset=>reset,s=>p(238)(48),cout=>p(239)(49));
FA_ff_6948:FAff port map(x=>p(164)(49),y=>p(165)(49),Cin=>p(166)(49),clock=>clock,reset=>reset,s=>p(238)(49),cout=>p(239)(50));
FA_ff_6949:FAff port map(x=>p(164)(50),y=>p(165)(50),Cin=>p(166)(50),clock=>clock,reset=>reset,s=>p(238)(50),cout=>p(239)(51));
FA_ff_6950:FAff port map(x=>p(164)(51),y=>p(165)(51),Cin=>p(166)(51),clock=>clock,reset=>reset,s=>p(238)(51),cout=>p(239)(52));
FA_ff_6951:FAff port map(x=>p(164)(52),y=>p(165)(52),Cin=>p(166)(52),clock=>clock,reset=>reset,s=>p(238)(52),cout=>p(239)(53));
FA_ff_6952:FAff port map(x=>p(164)(53),y=>p(165)(53),Cin=>p(166)(53),clock=>clock,reset=>reset,s=>p(238)(53),cout=>p(239)(54));
FA_ff_6953:FAff port map(x=>p(164)(54),y=>p(165)(54),Cin=>p(166)(54),clock=>clock,reset=>reset,s=>p(238)(54),cout=>p(239)(55));
FA_ff_6954:FAff port map(x=>p(164)(55),y=>p(165)(55),Cin=>p(166)(55),clock=>clock,reset=>reset,s=>p(238)(55),cout=>p(239)(56));
FA_ff_6955:FAff port map(x=>p(164)(56),y=>p(165)(56),Cin=>p(166)(56),clock=>clock,reset=>reset,s=>p(238)(56),cout=>p(239)(57));
FA_ff_6956:FAff port map(x=>p(164)(57),y=>p(165)(57),Cin=>p(166)(57),clock=>clock,reset=>reset,s=>p(238)(57),cout=>p(239)(58));
FA_ff_6957:FAff port map(x=>p(164)(58),y=>p(165)(58),Cin=>p(166)(58),clock=>clock,reset=>reset,s=>p(238)(58),cout=>p(239)(59));
FA_ff_6958:FAff port map(x=>p(164)(59),y=>p(165)(59),Cin=>p(166)(59),clock=>clock,reset=>reset,s=>p(238)(59),cout=>p(239)(60));
FA_ff_6959:FAff port map(x=>p(164)(60),y=>p(165)(60),Cin=>p(166)(60),clock=>clock,reset=>reset,s=>p(238)(60),cout=>p(239)(61));
FA_ff_6960:FAff port map(x=>p(164)(61),y=>p(165)(61),Cin=>p(166)(61),clock=>clock,reset=>reset,s=>p(238)(61),cout=>p(239)(62));
FA_ff_6961:FAff port map(x=>p(164)(62),y=>p(165)(62),Cin=>p(166)(62),clock=>clock,reset=>reset,s=>p(238)(62),cout=>p(239)(63));
FA_ff_6962:FAff port map(x=>p(164)(63),y=>p(165)(63),Cin=>p(166)(63),clock=>clock,reset=>reset,s=>p(238)(63),cout=>p(239)(64));
FA_ff_6963:FAff port map(x=>p(164)(64),y=>p(165)(64),Cin=>p(166)(64),clock=>clock,reset=>reset,s=>p(238)(64),cout=>p(239)(65));
FA_ff_6964:FAff port map(x=>p(164)(65),y=>p(165)(65),Cin=>p(166)(65),clock=>clock,reset=>reset,s=>p(238)(65),cout=>p(239)(66));
FA_ff_6965:FAff port map(x=>p(164)(66),y=>p(165)(66),Cin=>p(166)(66),clock=>clock,reset=>reset,s=>p(238)(66),cout=>p(239)(67));
FA_ff_6966:FAff port map(x=>p(164)(67),y=>p(165)(67),Cin=>p(166)(67),clock=>clock,reset=>reset,s=>p(238)(67),cout=>p(239)(68));
FA_ff_6967:FAff port map(x=>p(164)(68),y=>p(165)(68),Cin=>p(166)(68),clock=>clock,reset=>reset,s=>p(238)(68),cout=>p(239)(69));
FA_ff_6968:FAff port map(x=>p(164)(69),y=>p(165)(69),Cin=>p(166)(69),clock=>clock,reset=>reset,s=>p(238)(69),cout=>p(239)(70));
FA_ff_6969:FAff port map(x=>p(164)(70),y=>p(165)(70),Cin=>p(166)(70),clock=>clock,reset=>reset,s=>p(238)(70),cout=>p(239)(71));
FA_ff_6970:FAff port map(x=>p(164)(71),y=>p(165)(71),Cin=>p(166)(71),clock=>clock,reset=>reset,s=>p(238)(71),cout=>p(239)(72));
FA_ff_6971:FAff port map(x=>p(164)(72),y=>p(165)(72),Cin=>p(166)(72),clock=>clock,reset=>reset,s=>p(238)(72),cout=>p(239)(73));
FA_ff_6972:FAff port map(x=>p(164)(73),y=>p(165)(73),Cin=>p(166)(73),clock=>clock,reset=>reset,s=>p(238)(73),cout=>p(239)(74));
FA_ff_6973:FAff port map(x=>p(164)(74),y=>p(165)(74),Cin=>p(166)(74),clock=>clock,reset=>reset,s=>p(238)(74),cout=>p(239)(75));
FA_ff_6974:FAff port map(x=>p(164)(75),y=>p(165)(75),Cin=>p(166)(75),clock=>clock,reset=>reset,s=>p(238)(75),cout=>p(239)(76));
FA_ff_6975:FAff port map(x=>p(164)(76),y=>p(165)(76),Cin=>p(166)(76),clock=>clock,reset=>reset,s=>p(238)(76),cout=>p(239)(77));
FA_ff_6976:FAff port map(x=>p(164)(77),y=>p(165)(77),Cin=>p(166)(77),clock=>clock,reset=>reset,s=>p(238)(77),cout=>p(239)(78));
FA_ff_6977:FAff port map(x=>p(164)(78),y=>p(165)(78),Cin=>p(166)(78),clock=>clock,reset=>reset,s=>p(238)(78),cout=>p(239)(79));
FA_ff_6978:FAff port map(x=>p(164)(79),y=>p(165)(79),Cin=>p(166)(79),clock=>clock,reset=>reset,s=>p(238)(79),cout=>p(239)(80));
FA_ff_6979:FAff port map(x=>p(164)(80),y=>p(165)(80),Cin=>p(166)(80),clock=>clock,reset=>reset,s=>p(238)(80),cout=>p(239)(81));
FA_ff_6980:FAff port map(x=>p(164)(81),y=>p(165)(81),Cin=>p(166)(81),clock=>clock,reset=>reset,s=>p(238)(81),cout=>p(239)(82));
FA_ff_6981:FAff port map(x=>p(164)(82),y=>p(165)(82),Cin=>p(166)(82),clock=>clock,reset=>reset,s=>p(238)(82),cout=>p(239)(83));
FA_ff_6982:FAff port map(x=>p(164)(83),y=>p(165)(83),Cin=>p(166)(83),clock=>clock,reset=>reset,s=>p(238)(83),cout=>p(239)(84));
FA_ff_6983:FAff port map(x=>p(164)(84),y=>p(165)(84),Cin=>p(166)(84),clock=>clock,reset=>reset,s=>p(238)(84),cout=>p(239)(85));
FA_ff_6984:FAff port map(x=>p(164)(85),y=>p(165)(85),Cin=>p(166)(85),clock=>clock,reset=>reset,s=>p(238)(85),cout=>p(239)(86));
FA_ff_6985:FAff port map(x=>p(164)(86),y=>p(165)(86),Cin=>p(166)(86),clock=>clock,reset=>reset,s=>p(238)(86),cout=>p(239)(87));
FA_ff_6986:FAff port map(x=>p(164)(87),y=>p(165)(87),Cin=>p(166)(87),clock=>clock,reset=>reset,s=>p(238)(87),cout=>p(239)(88));
FA_ff_6987:FAff port map(x=>p(164)(88),y=>p(165)(88),Cin=>p(166)(88),clock=>clock,reset=>reset,s=>p(238)(88),cout=>p(239)(89));
FA_ff_6988:FAff port map(x=>p(164)(89),y=>p(165)(89),Cin=>p(166)(89),clock=>clock,reset=>reset,s=>p(238)(89),cout=>p(239)(90));
FA_ff_6989:FAff port map(x=>p(164)(90),y=>p(165)(90),Cin=>p(166)(90),clock=>clock,reset=>reset,s=>p(238)(90),cout=>p(239)(91));
FA_ff_6990:FAff port map(x=>p(164)(91),y=>p(165)(91),Cin=>p(166)(91),clock=>clock,reset=>reset,s=>p(238)(91),cout=>p(239)(92));
FA_ff_6991:FAff port map(x=>p(164)(92),y=>p(165)(92),Cin=>p(166)(92),clock=>clock,reset=>reset,s=>p(238)(92),cout=>p(239)(93));
FA_ff_6992:FAff port map(x=>p(164)(93),y=>p(165)(93),Cin=>p(166)(93),clock=>clock,reset=>reset,s=>p(238)(93),cout=>p(239)(94));
FA_ff_6993:FAff port map(x=>p(164)(94),y=>p(165)(94),Cin=>p(166)(94),clock=>clock,reset=>reset,s=>p(238)(94),cout=>p(239)(95));
FA_ff_6994:FAff port map(x=>p(164)(95),y=>p(165)(95),Cin=>p(166)(95),clock=>clock,reset=>reset,s=>p(238)(95),cout=>p(239)(96));
FA_ff_6995:FAff port map(x=>p(164)(96),y=>p(165)(96),Cin=>p(166)(96),clock=>clock,reset=>reset,s=>p(238)(96),cout=>p(239)(97));
FA_ff_6996:FAff port map(x=>p(164)(97),y=>p(165)(97),Cin=>p(166)(97),clock=>clock,reset=>reset,s=>p(238)(97),cout=>p(239)(98));
FA_ff_6997:FAff port map(x=>p(164)(98),y=>p(165)(98),Cin=>p(166)(98),clock=>clock,reset=>reset,s=>p(238)(98),cout=>p(239)(99));
FA_ff_6998:FAff port map(x=>p(164)(99),y=>p(165)(99),Cin=>p(166)(99),clock=>clock,reset=>reset,s=>p(238)(99),cout=>p(239)(100));
FA_ff_6999:FAff port map(x=>p(164)(100),y=>p(165)(100),Cin=>p(166)(100),clock=>clock,reset=>reset,s=>p(238)(100),cout=>p(239)(101));
FA_ff_7000:FAff port map(x=>p(164)(101),y=>p(165)(101),Cin=>p(166)(101),clock=>clock,reset=>reset,s=>p(238)(101),cout=>p(239)(102));
FA_ff_7001:FAff port map(x=>p(164)(102),y=>p(165)(102),Cin=>p(166)(102),clock=>clock,reset=>reset,s=>p(238)(102),cout=>p(239)(103));
FA_ff_7002:FAff port map(x=>p(164)(103),y=>p(165)(103),Cin=>p(166)(103),clock=>clock,reset=>reset,s=>p(238)(103),cout=>p(239)(104));
FA_ff_7003:FAff port map(x=>p(164)(104),y=>p(165)(104),Cin=>p(166)(104),clock=>clock,reset=>reset,s=>p(238)(104),cout=>p(239)(105));
FA_ff_7004:FAff port map(x=>p(164)(105),y=>p(165)(105),Cin=>p(166)(105),clock=>clock,reset=>reset,s=>p(238)(105),cout=>p(239)(106));
FA_ff_7005:FAff port map(x=>p(164)(106),y=>p(165)(106),Cin=>p(166)(106),clock=>clock,reset=>reset,s=>p(238)(106),cout=>p(239)(107));
FA_ff_7006:FAff port map(x=>p(164)(107),y=>p(165)(107),Cin=>p(166)(107),clock=>clock,reset=>reset,s=>p(238)(107),cout=>p(239)(108));
FA_ff_7007:FAff port map(x=>p(164)(108),y=>p(165)(108),Cin=>p(166)(108),clock=>clock,reset=>reset,s=>p(238)(108),cout=>p(239)(109));
FA_ff_7008:FAff port map(x=>p(164)(109),y=>p(165)(109),Cin=>p(166)(109),clock=>clock,reset=>reset,s=>p(238)(109),cout=>p(239)(110));
FA_ff_7009:FAff port map(x=>p(164)(110),y=>p(165)(110),Cin=>p(166)(110),clock=>clock,reset=>reset,s=>p(238)(110),cout=>p(239)(111));
FA_ff_7010:FAff port map(x=>p(164)(111),y=>p(165)(111),Cin=>p(166)(111),clock=>clock,reset=>reset,s=>p(238)(111),cout=>p(239)(112));
FA_ff_7011:FAff port map(x=>p(164)(112),y=>p(165)(112),Cin=>p(166)(112),clock=>clock,reset=>reset,s=>p(238)(112),cout=>p(239)(113));
FA_ff_7012:FAff port map(x=>p(164)(113),y=>p(165)(113),Cin=>p(166)(113),clock=>clock,reset=>reset,s=>p(238)(113),cout=>p(239)(114));
FA_ff_7013:FAff port map(x=>p(164)(114),y=>p(165)(114),Cin=>p(166)(114),clock=>clock,reset=>reset,s=>p(238)(114),cout=>p(239)(115));
FA_ff_7014:FAff port map(x=>p(164)(115),y=>p(165)(115),Cin=>p(166)(115),clock=>clock,reset=>reset,s=>p(238)(115),cout=>p(239)(116));
FA_ff_7015:FAff port map(x=>p(164)(116),y=>p(165)(116),Cin=>p(166)(116),clock=>clock,reset=>reset,s=>p(238)(116),cout=>p(239)(117));
FA_ff_7016:FAff port map(x=>p(164)(117),y=>p(165)(117),Cin=>p(166)(117),clock=>clock,reset=>reset,s=>p(238)(117),cout=>p(239)(118));
FA_ff_7017:FAff port map(x=>p(164)(118),y=>p(165)(118),Cin=>p(166)(118),clock=>clock,reset=>reset,s=>p(238)(118),cout=>p(239)(119));
FA_ff_7018:FAff port map(x=>p(164)(119),y=>p(165)(119),Cin=>p(166)(119),clock=>clock,reset=>reset,s=>p(238)(119),cout=>p(239)(120));
FA_ff_7019:FAff port map(x=>p(164)(120),y=>p(165)(120),Cin=>p(166)(120),clock=>clock,reset=>reset,s=>p(238)(120),cout=>p(239)(121));
FA_ff_7020:FAff port map(x=>p(164)(121),y=>p(165)(121),Cin=>p(166)(121),clock=>clock,reset=>reset,s=>p(238)(121),cout=>p(239)(122));
FA_ff_7021:FAff port map(x=>p(164)(122),y=>p(165)(122),Cin=>p(166)(122),clock=>clock,reset=>reset,s=>p(238)(122),cout=>p(239)(123));
FA_ff_7022:FAff port map(x=>p(164)(123),y=>p(165)(123),Cin=>p(166)(123),clock=>clock,reset=>reset,s=>p(238)(123),cout=>p(239)(124));
FA_ff_7023:FAff port map(x=>p(164)(124),y=>p(165)(124),Cin=>p(166)(124),clock=>clock,reset=>reset,s=>p(238)(124),cout=>p(239)(125));
FA_ff_7024:FAff port map(x=>p(164)(125),y=>p(165)(125),Cin=>p(166)(125),clock=>clock,reset=>reset,s=>p(238)(125),cout=>p(239)(126));
FA_ff_7025:FAff port map(x=>p(164)(126),y=>p(165)(126),Cin=>p(166)(126),clock=>clock,reset=>reset,s=>p(238)(126),cout=>p(239)(127));
FA_ff_7026:FAff port map(x=>p(164)(127),y=>p(165)(127),Cin=>p(166)(127),clock=>clock,reset=>reset,s=>p(238)(127),cout=>p(239)(128));
p(238)(128)<=p(165)(128);
p(240)(0)<=p(168)(0);
FA_ff_7027:FAff port map(x=>p(167)(1),y=>p(168)(1),Cin=>p(169)(1),clock=>clock,reset=>reset,s=>p(240)(1),cout=>p(241)(2));
FA_ff_7028:FAff port map(x=>p(167)(2),y=>p(168)(2),Cin=>p(169)(2),clock=>clock,reset=>reset,s=>p(240)(2),cout=>p(241)(3));
FA_ff_7029:FAff port map(x=>p(167)(3),y=>p(168)(3),Cin=>p(169)(3),clock=>clock,reset=>reset,s=>p(240)(3),cout=>p(241)(4));
FA_ff_7030:FAff port map(x=>p(167)(4),y=>p(168)(4),Cin=>p(169)(4),clock=>clock,reset=>reset,s=>p(240)(4),cout=>p(241)(5));
FA_ff_7031:FAff port map(x=>p(167)(5),y=>p(168)(5),Cin=>p(169)(5),clock=>clock,reset=>reset,s=>p(240)(5),cout=>p(241)(6));
FA_ff_7032:FAff port map(x=>p(167)(6),y=>p(168)(6),Cin=>p(169)(6),clock=>clock,reset=>reset,s=>p(240)(6),cout=>p(241)(7));
FA_ff_7033:FAff port map(x=>p(167)(7),y=>p(168)(7),Cin=>p(169)(7),clock=>clock,reset=>reset,s=>p(240)(7),cout=>p(241)(8));
FA_ff_7034:FAff port map(x=>p(167)(8),y=>p(168)(8),Cin=>p(169)(8),clock=>clock,reset=>reset,s=>p(240)(8),cout=>p(241)(9));
FA_ff_7035:FAff port map(x=>p(167)(9),y=>p(168)(9),Cin=>p(169)(9),clock=>clock,reset=>reset,s=>p(240)(9),cout=>p(241)(10));
FA_ff_7036:FAff port map(x=>p(167)(10),y=>p(168)(10),Cin=>p(169)(10),clock=>clock,reset=>reset,s=>p(240)(10),cout=>p(241)(11));
FA_ff_7037:FAff port map(x=>p(167)(11),y=>p(168)(11),Cin=>p(169)(11),clock=>clock,reset=>reset,s=>p(240)(11),cout=>p(241)(12));
FA_ff_7038:FAff port map(x=>p(167)(12),y=>p(168)(12),Cin=>p(169)(12),clock=>clock,reset=>reset,s=>p(240)(12),cout=>p(241)(13));
FA_ff_7039:FAff port map(x=>p(167)(13),y=>p(168)(13),Cin=>p(169)(13),clock=>clock,reset=>reset,s=>p(240)(13),cout=>p(241)(14));
FA_ff_7040:FAff port map(x=>p(167)(14),y=>p(168)(14),Cin=>p(169)(14),clock=>clock,reset=>reset,s=>p(240)(14),cout=>p(241)(15));
FA_ff_7041:FAff port map(x=>p(167)(15),y=>p(168)(15),Cin=>p(169)(15),clock=>clock,reset=>reset,s=>p(240)(15),cout=>p(241)(16));
FA_ff_7042:FAff port map(x=>p(167)(16),y=>p(168)(16),Cin=>p(169)(16),clock=>clock,reset=>reset,s=>p(240)(16),cout=>p(241)(17));
FA_ff_7043:FAff port map(x=>p(167)(17),y=>p(168)(17),Cin=>p(169)(17),clock=>clock,reset=>reset,s=>p(240)(17),cout=>p(241)(18));
FA_ff_7044:FAff port map(x=>p(167)(18),y=>p(168)(18),Cin=>p(169)(18),clock=>clock,reset=>reset,s=>p(240)(18),cout=>p(241)(19));
FA_ff_7045:FAff port map(x=>p(167)(19),y=>p(168)(19),Cin=>p(169)(19),clock=>clock,reset=>reset,s=>p(240)(19),cout=>p(241)(20));
FA_ff_7046:FAff port map(x=>p(167)(20),y=>p(168)(20),Cin=>p(169)(20),clock=>clock,reset=>reset,s=>p(240)(20),cout=>p(241)(21));
FA_ff_7047:FAff port map(x=>p(167)(21),y=>p(168)(21),Cin=>p(169)(21),clock=>clock,reset=>reset,s=>p(240)(21),cout=>p(241)(22));
FA_ff_7048:FAff port map(x=>p(167)(22),y=>p(168)(22),Cin=>p(169)(22),clock=>clock,reset=>reset,s=>p(240)(22),cout=>p(241)(23));
FA_ff_7049:FAff port map(x=>p(167)(23),y=>p(168)(23),Cin=>p(169)(23),clock=>clock,reset=>reset,s=>p(240)(23),cout=>p(241)(24));
FA_ff_7050:FAff port map(x=>p(167)(24),y=>p(168)(24),Cin=>p(169)(24),clock=>clock,reset=>reset,s=>p(240)(24),cout=>p(241)(25));
FA_ff_7051:FAff port map(x=>p(167)(25),y=>p(168)(25),Cin=>p(169)(25),clock=>clock,reset=>reset,s=>p(240)(25),cout=>p(241)(26));
FA_ff_7052:FAff port map(x=>p(167)(26),y=>p(168)(26),Cin=>p(169)(26),clock=>clock,reset=>reset,s=>p(240)(26),cout=>p(241)(27));
FA_ff_7053:FAff port map(x=>p(167)(27),y=>p(168)(27),Cin=>p(169)(27),clock=>clock,reset=>reset,s=>p(240)(27),cout=>p(241)(28));
FA_ff_7054:FAff port map(x=>p(167)(28),y=>p(168)(28),Cin=>p(169)(28),clock=>clock,reset=>reset,s=>p(240)(28),cout=>p(241)(29));
FA_ff_7055:FAff port map(x=>p(167)(29),y=>p(168)(29),Cin=>p(169)(29),clock=>clock,reset=>reset,s=>p(240)(29),cout=>p(241)(30));
FA_ff_7056:FAff port map(x=>p(167)(30),y=>p(168)(30),Cin=>p(169)(30),clock=>clock,reset=>reset,s=>p(240)(30),cout=>p(241)(31));
FA_ff_7057:FAff port map(x=>p(167)(31),y=>p(168)(31),Cin=>p(169)(31),clock=>clock,reset=>reset,s=>p(240)(31),cout=>p(241)(32));
FA_ff_7058:FAff port map(x=>p(167)(32),y=>p(168)(32),Cin=>p(169)(32),clock=>clock,reset=>reset,s=>p(240)(32),cout=>p(241)(33));
FA_ff_7059:FAff port map(x=>p(167)(33),y=>p(168)(33),Cin=>p(169)(33),clock=>clock,reset=>reset,s=>p(240)(33),cout=>p(241)(34));
FA_ff_7060:FAff port map(x=>p(167)(34),y=>p(168)(34),Cin=>p(169)(34),clock=>clock,reset=>reset,s=>p(240)(34),cout=>p(241)(35));
FA_ff_7061:FAff port map(x=>p(167)(35),y=>p(168)(35),Cin=>p(169)(35),clock=>clock,reset=>reset,s=>p(240)(35),cout=>p(241)(36));
FA_ff_7062:FAff port map(x=>p(167)(36),y=>p(168)(36),Cin=>p(169)(36),clock=>clock,reset=>reset,s=>p(240)(36),cout=>p(241)(37));
FA_ff_7063:FAff port map(x=>p(167)(37),y=>p(168)(37),Cin=>p(169)(37),clock=>clock,reset=>reset,s=>p(240)(37),cout=>p(241)(38));
FA_ff_7064:FAff port map(x=>p(167)(38),y=>p(168)(38),Cin=>p(169)(38),clock=>clock,reset=>reset,s=>p(240)(38),cout=>p(241)(39));
FA_ff_7065:FAff port map(x=>p(167)(39),y=>p(168)(39),Cin=>p(169)(39),clock=>clock,reset=>reset,s=>p(240)(39),cout=>p(241)(40));
FA_ff_7066:FAff port map(x=>p(167)(40),y=>p(168)(40),Cin=>p(169)(40),clock=>clock,reset=>reset,s=>p(240)(40),cout=>p(241)(41));
FA_ff_7067:FAff port map(x=>p(167)(41),y=>p(168)(41),Cin=>p(169)(41),clock=>clock,reset=>reset,s=>p(240)(41),cout=>p(241)(42));
FA_ff_7068:FAff port map(x=>p(167)(42),y=>p(168)(42),Cin=>p(169)(42),clock=>clock,reset=>reset,s=>p(240)(42),cout=>p(241)(43));
FA_ff_7069:FAff port map(x=>p(167)(43),y=>p(168)(43),Cin=>p(169)(43),clock=>clock,reset=>reset,s=>p(240)(43),cout=>p(241)(44));
FA_ff_7070:FAff port map(x=>p(167)(44),y=>p(168)(44),Cin=>p(169)(44),clock=>clock,reset=>reset,s=>p(240)(44),cout=>p(241)(45));
FA_ff_7071:FAff port map(x=>p(167)(45),y=>p(168)(45),Cin=>p(169)(45),clock=>clock,reset=>reset,s=>p(240)(45),cout=>p(241)(46));
FA_ff_7072:FAff port map(x=>p(167)(46),y=>p(168)(46),Cin=>p(169)(46),clock=>clock,reset=>reset,s=>p(240)(46),cout=>p(241)(47));
FA_ff_7073:FAff port map(x=>p(167)(47),y=>p(168)(47),Cin=>p(169)(47),clock=>clock,reset=>reset,s=>p(240)(47),cout=>p(241)(48));
FA_ff_7074:FAff port map(x=>p(167)(48),y=>p(168)(48),Cin=>p(169)(48),clock=>clock,reset=>reset,s=>p(240)(48),cout=>p(241)(49));
FA_ff_7075:FAff port map(x=>p(167)(49),y=>p(168)(49),Cin=>p(169)(49),clock=>clock,reset=>reset,s=>p(240)(49),cout=>p(241)(50));
FA_ff_7076:FAff port map(x=>p(167)(50),y=>p(168)(50),Cin=>p(169)(50),clock=>clock,reset=>reset,s=>p(240)(50),cout=>p(241)(51));
FA_ff_7077:FAff port map(x=>p(167)(51),y=>p(168)(51),Cin=>p(169)(51),clock=>clock,reset=>reset,s=>p(240)(51),cout=>p(241)(52));
FA_ff_7078:FAff port map(x=>p(167)(52),y=>p(168)(52),Cin=>p(169)(52),clock=>clock,reset=>reset,s=>p(240)(52),cout=>p(241)(53));
FA_ff_7079:FAff port map(x=>p(167)(53),y=>p(168)(53),Cin=>p(169)(53),clock=>clock,reset=>reset,s=>p(240)(53),cout=>p(241)(54));
FA_ff_7080:FAff port map(x=>p(167)(54),y=>p(168)(54),Cin=>p(169)(54),clock=>clock,reset=>reset,s=>p(240)(54),cout=>p(241)(55));
FA_ff_7081:FAff port map(x=>p(167)(55),y=>p(168)(55),Cin=>p(169)(55),clock=>clock,reset=>reset,s=>p(240)(55),cout=>p(241)(56));
FA_ff_7082:FAff port map(x=>p(167)(56),y=>p(168)(56),Cin=>p(169)(56),clock=>clock,reset=>reset,s=>p(240)(56),cout=>p(241)(57));
FA_ff_7083:FAff port map(x=>p(167)(57),y=>p(168)(57),Cin=>p(169)(57),clock=>clock,reset=>reset,s=>p(240)(57),cout=>p(241)(58));
FA_ff_7084:FAff port map(x=>p(167)(58),y=>p(168)(58),Cin=>p(169)(58),clock=>clock,reset=>reset,s=>p(240)(58),cout=>p(241)(59));
FA_ff_7085:FAff port map(x=>p(167)(59),y=>p(168)(59),Cin=>p(169)(59),clock=>clock,reset=>reset,s=>p(240)(59),cout=>p(241)(60));
FA_ff_7086:FAff port map(x=>p(167)(60),y=>p(168)(60),Cin=>p(169)(60),clock=>clock,reset=>reset,s=>p(240)(60),cout=>p(241)(61));
FA_ff_7087:FAff port map(x=>p(167)(61),y=>p(168)(61),Cin=>p(169)(61),clock=>clock,reset=>reset,s=>p(240)(61),cout=>p(241)(62));
FA_ff_7088:FAff port map(x=>p(167)(62),y=>p(168)(62),Cin=>p(169)(62),clock=>clock,reset=>reset,s=>p(240)(62),cout=>p(241)(63));
FA_ff_7089:FAff port map(x=>p(167)(63),y=>p(168)(63),Cin=>p(169)(63),clock=>clock,reset=>reset,s=>p(240)(63),cout=>p(241)(64));
FA_ff_7090:FAff port map(x=>p(167)(64),y=>p(168)(64),Cin=>p(169)(64),clock=>clock,reset=>reset,s=>p(240)(64),cout=>p(241)(65));
FA_ff_7091:FAff port map(x=>p(167)(65),y=>p(168)(65),Cin=>p(169)(65),clock=>clock,reset=>reset,s=>p(240)(65),cout=>p(241)(66));
FA_ff_7092:FAff port map(x=>p(167)(66),y=>p(168)(66),Cin=>p(169)(66),clock=>clock,reset=>reset,s=>p(240)(66),cout=>p(241)(67));
FA_ff_7093:FAff port map(x=>p(167)(67),y=>p(168)(67),Cin=>p(169)(67),clock=>clock,reset=>reset,s=>p(240)(67),cout=>p(241)(68));
FA_ff_7094:FAff port map(x=>p(167)(68),y=>p(168)(68),Cin=>p(169)(68),clock=>clock,reset=>reset,s=>p(240)(68),cout=>p(241)(69));
FA_ff_7095:FAff port map(x=>p(167)(69),y=>p(168)(69),Cin=>p(169)(69),clock=>clock,reset=>reset,s=>p(240)(69),cout=>p(241)(70));
FA_ff_7096:FAff port map(x=>p(167)(70),y=>p(168)(70),Cin=>p(169)(70),clock=>clock,reset=>reset,s=>p(240)(70),cout=>p(241)(71));
FA_ff_7097:FAff port map(x=>p(167)(71),y=>p(168)(71),Cin=>p(169)(71),clock=>clock,reset=>reset,s=>p(240)(71),cout=>p(241)(72));
FA_ff_7098:FAff port map(x=>p(167)(72),y=>p(168)(72),Cin=>p(169)(72),clock=>clock,reset=>reset,s=>p(240)(72),cout=>p(241)(73));
FA_ff_7099:FAff port map(x=>p(167)(73),y=>p(168)(73),Cin=>p(169)(73),clock=>clock,reset=>reset,s=>p(240)(73),cout=>p(241)(74));
FA_ff_7100:FAff port map(x=>p(167)(74),y=>p(168)(74),Cin=>p(169)(74),clock=>clock,reset=>reset,s=>p(240)(74),cout=>p(241)(75));
FA_ff_7101:FAff port map(x=>p(167)(75),y=>p(168)(75),Cin=>p(169)(75),clock=>clock,reset=>reset,s=>p(240)(75),cout=>p(241)(76));
FA_ff_7102:FAff port map(x=>p(167)(76),y=>p(168)(76),Cin=>p(169)(76),clock=>clock,reset=>reset,s=>p(240)(76),cout=>p(241)(77));
FA_ff_7103:FAff port map(x=>p(167)(77),y=>p(168)(77),Cin=>p(169)(77),clock=>clock,reset=>reset,s=>p(240)(77),cout=>p(241)(78));
FA_ff_7104:FAff port map(x=>p(167)(78),y=>p(168)(78),Cin=>p(169)(78),clock=>clock,reset=>reset,s=>p(240)(78),cout=>p(241)(79));
FA_ff_7105:FAff port map(x=>p(167)(79),y=>p(168)(79),Cin=>p(169)(79),clock=>clock,reset=>reset,s=>p(240)(79),cout=>p(241)(80));
FA_ff_7106:FAff port map(x=>p(167)(80),y=>p(168)(80),Cin=>p(169)(80),clock=>clock,reset=>reset,s=>p(240)(80),cout=>p(241)(81));
FA_ff_7107:FAff port map(x=>p(167)(81),y=>p(168)(81),Cin=>p(169)(81),clock=>clock,reset=>reset,s=>p(240)(81),cout=>p(241)(82));
FA_ff_7108:FAff port map(x=>p(167)(82),y=>p(168)(82),Cin=>p(169)(82),clock=>clock,reset=>reset,s=>p(240)(82),cout=>p(241)(83));
FA_ff_7109:FAff port map(x=>p(167)(83),y=>p(168)(83),Cin=>p(169)(83),clock=>clock,reset=>reset,s=>p(240)(83),cout=>p(241)(84));
FA_ff_7110:FAff port map(x=>p(167)(84),y=>p(168)(84),Cin=>p(169)(84),clock=>clock,reset=>reset,s=>p(240)(84),cout=>p(241)(85));
FA_ff_7111:FAff port map(x=>p(167)(85),y=>p(168)(85),Cin=>p(169)(85),clock=>clock,reset=>reset,s=>p(240)(85),cout=>p(241)(86));
FA_ff_7112:FAff port map(x=>p(167)(86),y=>p(168)(86),Cin=>p(169)(86),clock=>clock,reset=>reset,s=>p(240)(86),cout=>p(241)(87));
FA_ff_7113:FAff port map(x=>p(167)(87),y=>p(168)(87),Cin=>p(169)(87),clock=>clock,reset=>reset,s=>p(240)(87),cout=>p(241)(88));
FA_ff_7114:FAff port map(x=>p(167)(88),y=>p(168)(88),Cin=>p(169)(88),clock=>clock,reset=>reset,s=>p(240)(88),cout=>p(241)(89));
FA_ff_7115:FAff port map(x=>p(167)(89),y=>p(168)(89),Cin=>p(169)(89),clock=>clock,reset=>reset,s=>p(240)(89),cout=>p(241)(90));
FA_ff_7116:FAff port map(x=>p(167)(90),y=>p(168)(90),Cin=>p(169)(90),clock=>clock,reset=>reset,s=>p(240)(90),cout=>p(241)(91));
FA_ff_7117:FAff port map(x=>p(167)(91),y=>p(168)(91),Cin=>p(169)(91),clock=>clock,reset=>reset,s=>p(240)(91),cout=>p(241)(92));
FA_ff_7118:FAff port map(x=>p(167)(92),y=>p(168)(92),Cin=>p(169)(92),clock=>clock,reset=>reset,s=>p(240)(92),cout=>p(241)(93));
FA_ff_7119:FAff port map(x=>p(167)(93),y=>p(168)(93),Cin=>p(169)(93),clock=>clock,reset=>reset,s=>p(240)(93),cout=>p(241)(94));
FA_ff_7120:FAff port map(x=>p(167)(94),y=>p(168)(94),Cin=>p(169)(94),clock=>clock,reset=>reset,s=>p(240)(94),cout=>p(241)(95));
FA_ff_7121:FAff port map(x=>p(167)(95),y=>p(168)(95),Cin=>p(169)(95),clock=>clock,reset=>reset,s=>p(240)(95),cout=>p(241)(96));
FA_ff_7122:FAff port map(x=>p(167)(96),y=>p(168)(96),Cin=>p(169)(96),clock=>clock,reset=>reset,s=>p(240)(96),cout=>p(241)(97));
FA_ff_7123:FAff port map(x=>p(167)(97),y=>p(168)(97),Cin=>p(169)(97),clock=>clock,reset=>reset,s=>p(240)(97),cout=>p(241)(98));
FA_ff_7124:FAff port map(x=>p(167)(98),y=>p(168)(98),Cin=>p(169)(98),clock=>clock,reset=>reset,s=>p(240)(98),cout=>p(241)(99));
FA_ff_7125:FAff port map(x=>p(167)(99),y=>p(168)(99),Cin=>p(169)(99),clock=>clock,reset=>reset,s=>p(240)(99),cout=>p(241)(100));
FA_ff_7126:FAff port map(x=>p(167)(100),y=>p(168)(100),Cin=>p(169)(100),clock=>clock,reset=>reset,s=>p(240)(100),cout=>p(241)(101));
FA_ff_7127:FAff port map(x=>p(167)(101),y=>p(168)(101),Cin=>p(169)(101),clock=>clock,reset=>reset,s=>p(240)(101),cout=>p(241)(102));
FA_ff_7128:FAff port map(x=>p(167)(102),y=>p(168)(102),Cin=>p(169)(102),clock=>clock,reset=>reset,s=>p(240)(102),cout=>p(241)(103));
FA_ff_7129:FAff port map(x=>p(167)(103),y=>p(168)(103),Cin=>p(169)(103),clock=>clock,reset=>reset,s=>p(240)(103),cout=>p(241)(104));
FA_ff_7130:FAff port map(x=>p(167)(104),y=>p(168)(104),Cin=>p(169)(104),clock=>clock,reset=>reset,s=>p(240)(104),cout=>p(241)(105));
FA_ff_7131:FAff port map(x=>p(167)(105),y=>p(168)(105),Cin=>p(169)(105),clock=>clock,reset=>reset,s=>p(240)(105),cout=>p(241)(106));
FA_ff_7132:FAff port map(x=>p(167)(106),y=>p(168)(106),Cin=>p(169)(106),clock=>clock,reset=>reset,s=>p(240)(106),cout=>p(241)(107));
FA_ff_7133:FAff port map(x=>p(167)(107),y=>p(168)(107),Cin=>p(169)(107),clock=>clock,reset=>reset,s=>p(240)(107),cout=>p(241)(108));
FA_ff_7134:FAff port map(x=>p(167)(108),y=>p(168)(108),Cin=>p(169)(108),clock=>clock,reset=>reset,s=>p(240)(108),cout=>p(241)(109));
FA_ff_7135:FAff port map(x=>p(167)(109),y=>p(168)(109),Cin=>p(169)(109),clock=>clock,reset=>reset,s=>p(240)(109),cout=>p(241)(110));
FA_ff_7136:FAff port map(x=>p(167)(110),y=>p(168)(110),Cin=>p(169)(110),clock=>clock,reset=>reset,s=>p(240)(110),cout=>p(241)(111));
FA_ff_7137:FAff port map(x=>p(167)(111),y=>p(168)(111),Cin=>p(169)(111),clock=>clock,reset=>reset,s=>p(240)(111),cout=>p(241)(112));
FA_ff_7138:FAff port map(x=>p(167)(112),y=>p(168)(112),Cin=>p(169)(112),clock=>clock,reset=>reset,s=>p(240)(112),cout=>p(241)(113));
FA_ff_7139:FAff port map(x=>p(167)(113),y=>p(168)(113),Cin=>p(169)(113),clock=>clock,reset=>reset,s=>p(240)(113),cout=>p(241)(114));
FA_ff_7140:FAff port map(x=>p(167)(114),y=>p(168)(114),Cin=>p(169)(114),clock=>clock,reset=>reset,s=>p(240)(114),cout=>p(241)(115));
FA_ff_7141:FAff port map(x=>p(167)(115),y=>p(168)(115),Cin=>p(169)(115),clock=>clock,reset=>reset,s=>p(240)(115),cout=>p(241)(116));
FA_ff_7142:FAff port map(x=>p(167)(116),y=>p(168)(116),Cin=>p(169)(116),clock=>clock,reset=>reset,s=>p(240)(116),cout=>p(241)(117));
FA_ff_7143:FAff port map(x=>p(167)(117),y=>p(168)(117),Cin=>p(169)(117),clock=>clock,reset=>reset,s=>p(240)(117),cout=>p(241)(118));
FA_ff_7144:FAff port map(x=>p(167)(118),y=>p(168)(118),Cin=>p(169)(118),clock=>clock,reset=>reset,s=>p(240)(118),cout=>p(241)(119));
FA_ff_7145:FAff port map(x=>p(167)(119),y=>p(168)(119),Cin=>p(169)(119),clock=>clock,reset=>reset,s=>p(240)(119),cout=>p(241)(120));
FA_ff_7146:FAff port map(x=>p(167)(120),y=>p(168)(120),Cin=>p(169)(120),clock=>clock,reset=>reset,s=>p(240)(120),cout=>p(241)(121));
FA_ff_7147:FAff port map(x=>p(167)(121),y=>p(168)(121),Cin=>p(169)(121),clock=>clock,reset=>reset,s=>p(240)(121),cout=>p(241)(122));
FA_ff_7148:FAff port map(x=>p(167)(122),y=>p(168)(122),Cin=>p(169)(122),clock=>clock,reset=>reset,s=>p(240)(122),cout=>p(241)(123));
FA_ff_7149:FAff port map(x=>p(167)(123),y=>p(168)(123),Cin=>p(169)(123),clock=>clock,reset=>reset,s=>p(240)(123),cout=>p(241)(124));
FA_ff_7150:FAff port map(x=>p(167)(124),y=>p(168)(124),Cin=>p(169)(124),clock=>clock,reset=>reset,s=>p(240)(124),cout=>p(241)(125));
FA_ff_7151:FAff port map(x=>p(167)(125),y=>p(168)(125),Cin=>p(169)(125),clock=>clock,reset=>reset,s=>p(240)(125),cout=>p(241)(126));
FA_ff_7152:FAff port map(x=>p(167)(126),y=>p(168)(126),Cin=>p(169)(126),clock=>clock,reset=>reset,s=>p(240)(126),cout=>p(241)(127));
FA_ff_7153:FAff port map(x=>p(167)(127),y=>p(168)(127),Cin=>p(169)(127),clock=>clock,reset=>reset,s=>p(240)(127),cout=>p(241)(128));
HA_ff_13:HAff port map(x=>p(167)(128),y=>p(169)(128),clock=>clock,reset=>reset,s=>p(240)(128),c=>p(241)(129));
HA_ff_14:HAff port map(x=>p(170)(0),y=>p(172)(0),clock=>clock,reset=>reset,s=>p(242)(0),c=>p(243)(1));
FA_ff_7154:FAff port map(x=>p(170)(1),y=>p(171)(1),Cin=>p(172)(1),clock=>clock,reset=>reset,s=>p(242)(1),cout=>p(243)(2));
FA_ff_7155:FAff port map(x=>p(170)(2),y=>p(171)(2),Cin=>p(172)(2),clock=>clock,reset=>reset,s=>p(242)(2),cout=>p(243)(3));
FA_ff_7156:FAff port map(x=>p(170)(3),y=>p(171)(3),Cin=>p(172)(3),clock=>clock,reset=>reset,s=>p(242)(3),cout=>p(243)(4));
FA_ff_7157:FAff port map(x=>p(170)(4),y=>p(171)(4),Cin=>p(172)(4),clock=>clock,reset=>reset,s=>p(242)(4),cout=>p(243)(5));
FA_ff_7158:FAff port map(x=>p(170)(5),y=>p(171)(5),Cin=>p(172)(5),clock=>clock,reset=>reset,s=>p(242)(5),cout=>p(243)(6));
FA_ff_7159:FAff port map(x=>p(170)(6),y=>p(171)(6),Cin=>p(172)(6),clock=>clock,reset=>reset,s=>p(242)(6),cout=>p(243)(7));
FA_ff_7160:FAff port map(x=>p(170)(7),y=>p(171)(7),Cin=>p(172)(7),clock=>clock,reset=>reset,s=>p(242)(7),cout=>p(243)(8));
FA_ff_7161:FAff port map(x=>p(170)(8),y=>p(171)(8),Cin=>p(172)(8),clock=>clock,reset=>reset,s=>p(242)(8),cout=>p(243)(9));
FA_ff_7162:FAff port map(x=>p(170)(9),y=>p(171)(9),Cin=>p(172)(9),clock=>clock,reset=>reset,s=>p(242)(9),cout=>p(243)(10));
FA_ff_7163:FAff port map(x=>p(170)(10),y=>p(171)(10),Cin=>p(172)(10),clock=>clock,reset=>reset,s=>p(242)(10),cout=>p(243)(11));
FA_ff_7164:FAff port map(x=>p(170)(11),y=>p(171)(11),Cin=>p(172)(11),clock=>clock,reset=>reset,s=>p(242)(11),cout=>p(243)(12));
FA_ff_7165:FAff port map(x=>p(170)(12),y=>p(171)(12),Cin=>p(172)(12),clock=>clock,reset=>reset,s=>p(242)(12),cout=>p(243)(13));
FA_ff_7166:FAff port map(x=>p(170)(13),y=>p(171)(13),Cin=>p(172)(13),clock=>clock,reset=>reset,s=>p(242)(13),cout=>p(243)(14));
FA_ff_7167:FAff port map(x=>p(170)(14),y=>p(171)(14),Cin=>p(172)(14),clock=>clock,reset=>reset,s=>p(242)(14),cout=>p(243)(15));
FA_ff_7168:FAff port map(x=>p(170)(15),y=>p(171)(15),Cin=>p(172)(15),clock=>clock,reset=>reset,s=>p(242)(15),cout=>p(243)(16));
FA_ff_7169:FAff port map(x=>p(170)(16),y=>p(171)(16),Cin=>p(172)(16),clock=>clock,reset=>reset,s=>p(242)(16),cout=>p(243)(17));
FA_ff_7170:FAff port map(x=>p(170)(17),y=>p(171)(17),Cin=>p(172)(17),clock=>clock,reset=>reset,s=>p(242)(17),cout=>p(243)(18));
FA_ff_7171:FAff port map(x=>p(170)(18),y=>p(171)(18),Cin=>p(172)(18),clock=>clock,reset=>reset,s=>p(242)(18),cout=>p(243)(19));
FA_ff_7172:FAff port map(x=>p(170)(19),y=>p(171)(19),Cin=>p(172)(19),clock=>clock,reset=>reset,s=>p(242)(19),cout=>p(243)(20));
FA_ff_7173:FAff port map(x=>p(170)(20),y=>p(171)(20),Cin=>p(172)(20),clock=>clock,reset=>reset,s=>p(242)(20),cout=>p(243)(21));
FA_ff_7174:FAff port map(x=>p(170)(21),y=>p(171)(21),Cin=>p(172)(21),clock=>clock,reset=>reset,s=>p(242)(21),cout=>p(243)(22));
FA_ff_7175:FAff port map(x=>p(170)(22),y=>p(171)(22),Cin=>p(172)(22),clock=>clock,reset=>reset,s=>p(242)(22),cout=>p(243)(23));
FA_ff_7176:FAff port map(x=>p(170)(23),y=>p(171)(23),Cin=>p(172)(23),clock=>clock,reset=>reset,s=>p(242)(23),cout=>p(243)(24));
FA_ff_7177:FAff port map(x=>p(170)(24),y=>p(171)(24),Cin=>p(172)(24),clock=>clock,reset=>reset,s=>p(242)(24),cout=>p(243)(25));
FA_ff_7178:FAff port map(x=>p(170)(25),y=>p(171)(25),Cin=>p(172)(25),clock=>clock,reset=>reset,s=>p(242)(25),cout=>p(243)(26));
FA_ff_7179:FAff port map(x=>p(170)(26),y=>p(171)(26),Cin=>p(172)(26),clock=>clock,reset=>reset,s=>p(242)(26),cout=>p(243)(27));
FA_ff_7180:FAff port map(x=>p(170)(27),y=>p(171)(27),Cin=>p(172)(27),clock=>clock,reset=>reset,s=>p(242)(27),cout=>p(243)(28));
FA_ff_7181:FAff port map(x=>p(170)(28),y=>p(171)(28),Cin=>p(172)(28),clock=>clock,reset=>reset,s=>p(242)(28),cout=>p(243)(29));
FA_ff_7182:FAff port map(x=>p(170)(29),y=>p(171)(29),Cin=>p(172)(29),clock=>clock,reset=>reset,s=>p(242)(29),cout=>p(243)(30));
FA_ff_7183:FAff port map(x=>p(170)(30),y=>p(171)(30),Cin=>p(172)(30),clock=>clock,reset=>reset,s=>p(242)(30),cout=>p(243)(31));
FA_ff_7184:FAff port map(x=>p(170)(31),y=>p(171)(31),Cin=>p(172)(31),clock=>clock,reset=>reset,s=>p(242)(31),cout=>p(243)(32));
FA_ff_7185:FAff port map(x=>p(170)(32),y=>p(171)(32),Cin=>p(172)(32),clock=>clock,reset=>reset,s=>p(242)(32),cout=>p(243)(33));
FA_ff_7186:FAff port map(x=>p(170)(33),y=>p(171)(33),Cin=>p(172)(33),clock=>clock,reset=>reset,s=>p(242)(33),cout=>p(243)(34));
FA_ff_7187:FAff port map(x=>p(170)(34),y=>p(171)(34),Cin=>p(172)(34),clock=>clock,reset=>reset,s=>p(242)(34),cout=>p(243)(35));
FA_ff_7188:FAff port map(x=>p(170)(35),y=>p(171)(35),Cin=>p(172)(35),clock=>clock,reset=>reset,s=>p(242)(35),cout=>p(243)(36));
FA_ff_7189:FAff port map(x=>p(170)(36),y=>p(171)(36),Cin=>p(172)(36),clock=>clock,reset=>reset,s=>p(242)(36),cout=>p(243)(37));
FA_ff_7190:FAff port map(x=>p(170)(37),y=>p(171)(37),Cin=>p(172)(37),clock=>clock,reset=>reset,s=>p(242)(37),cout=>p(243)(38));
FA_ff_7191:FAff port map(x=>p(170)(38),y=>p(171)(38),Cin=>p(172)(38),clock=>clock,reset=>reset,s=>p(242)(38),cout=>p(243)(39));
FA_ff_7192:FAff port map(x=>p(170)(39),y=>p(171)(39),Cin=>p(172)(39),clock=>clock,reset=>reset,s=>p(242)(39),cout=>p(243)(40));
FA_ff_7193:FAff port map(x=>p(170)(40),y=>p(171)(40),Cin=>p(172)(40),clock=>clock,reset=>reset,s=>p(242)(40),cout=>p(243)(41));
FA_ff_7194:FAff port map(x=>p(170)(41),y=>p(171)(41),Cin=>p(172)(41),clock=>clock,reset=>reset,s=>p(242)(41),cout=>p(243)(42));
FA_ff_7195:FAff port map(x=>p(170)(42),y=>p(171)(42),Cin=>p(172)(42),clock=>clock,reset=>reset,s=>p(242)(42),cout=>p(243)(43));
FA_ff_7196:FAff port map(x=>p(170)(43),y=>p(171)(43),Cin=>p(172)(43),clock=>clock,reset=>reset,s=>p(242)(43),cout=>p(243)(44));
FA_ff_7197:FAff port map(x=>p(170)(44),y=>p(171)(44),Cin=>p(172)(44),clock=>clock,reset=>reset,s=>p(242)(44),cout=>p(243)(45));
FA_ff_7198:FAff port map(x=>p(170)(45),y=>p(171)(45),Cin=>p(172)(45),clock=>clock,reset=>reset,s=>p(242)(45),cout=>p(243)(46));
FA_ff_7199:FAff port map(x=>p(170)(46),y=>p(171)(46),Cin=>p(172)(46),clock=>clock,reset=>reset,s=>p(242)(46),cout=>p(243)(47));
FA_ff_7200:FAff port map(x=>p(170)(47),y=>p(171)(47),Cin=>p(172)(47),clock=>clock,reset=>reset,s=>p(242)(47),cout=>p(243)(48));
FA_ff_7201:FAff port map(x=>p(170)(48),y=>p(171)(48),Cin=>p(172)(48),clock=>clock,reset=>reset,s=>p(242)(48),cout=>p(243)(49));
FA_ff_7202:FAff port map(x=>p(170)(49),y=>p(171)(49),Cin=>p(172)(49),clock=>clock,reset=>reset,s=>p(242)(49),cout=>p(243)(50));
FA_ff_7203:FAff port map(x=>p(170)(50),y=>p(171)(50),Cin=>p(172)(50),clock=>clock,reset=>reset,s=>p(242)(50),cout=>p(243)(51));
FA_ff_7204:FAff port map(x=>p(170)(51),y=>p(171)(51),Cin=>p(172)(51),clock=>clock,reset=>reset,s=>p(242)(51),cout=>p(243)(52));
FA_ff_7205:FAff port map(x=>p(170)(52),y=>p(171)(52),Cin=>p(172)(52),clock=>clock,reset=>reset,s=>p(242)(52),cout=>p(243)(53));
FA_ff_7206:FAff port map(x=>p(170)(53),y=>p(171)(53),Cin=>p(172)(53),clock=>clock,reset=>reset,s=>p(242)(53),cout=>p(243)(54));
FA_ff_7207:FAff port map(x=>p(170)(54),y=>p(171)(54),Cin=>p(172)(54),clock=>clock,reset=>reset,s=>p(242)(54),cout=>p(243)(55));
FA_ff_7208:FAff port map(x=>p(170)(55),y=>p(171)(55),Cin=>p(172)(55),clock=>clock,reset=>reset,s=>p(242)(55),cout=>p(243)(56));
FA_ff_7209:FAff port map(x=>p(170)(56),y=>p(171)(56),Cin=>p(172)(56),clock=>clock,reset=>reset,s=>p(242)(56),cout=>p(243)(57));
FA_ff_7210:FAff port map(x=>p(170)(57),y=>p(171)(57),Cin=>p(172)(57),clock=>clock,reset=>reset,s=>p(242)(57),cout=>p(243)(58));
FA_ff_7211:FAff port map(x=>p(170)(58),y=>p(171)(58),Cin=>p(172)(58),clock=>clock,reset=>reset,s=>p(242)(58),cout=>p(243)(59));
FA_ff_7212:FAff port map(x=>p(170)(59),y=>p(171)(59),Cin=>p(172)(59),clock=>clock,reset=>reset,s=>p(242)(59),cout=>p(243)(60));
FA_ff_7213:FAff port map(x=>p(170)(60),y=>p(171)(60),Cin=>p(172)(60),clock=>clock,reset=>reset,s=>p(242)(60),cout=>p(243)(61));
FA_ff_7214:FAff port map(x=>p(170)(61),y=>p(171)(61),Cin=>p(172)(61),clock=>clock,reset=>reset,s=>p(242)(61),cout=>p(243)(62));
FA_ff_7215:FAff port map(x=>p(170)(62),y=>p(171)(62),Cin=>p(172)(62),clock=>clock,reset=>reset,s=>p(242)(62),cout=>p(243)(63));
FA_ff_7216:FAff port map(x=>p(170)(63),y=>p(171)(63),Cin=>p(172)(63),clock=>clock,reset=>reset,s=>p(242)(63),cout=>p(243)(64));
FA_ff_7217:FAff port map(x=>p(170)(64),y=>p(171)(64),Cin=>p(172)(64),clock=>clock,reset=>reset,s=>p(242)(64),cout=>p(243)(65));
FA_ff_7218:FAff port map(x=>p(170)(65),y=>p(171)(65),Cin=>p(172)(65),clock=>clock,reset=>reset,s=>p(242)(65),cout=>p(243)(66));
FA_ff_7219:FAff port map(x=>p(170)(66),y=>p(171)(66),Cin=>p(172)(66),clock=>clock,reset=>reset,s=>p(242)(66),cout=>p(243)(67));
FA_ff_7220:FAff port map(x=>p(170)(67),y=>p(171)(67),Cin=>p(172)(67),clock=>clock,reset=>reset,s=>p(242)(67),cout=>p(243)(68));
FA_ff_7221:FAff port map(x=>p(170)(68),y=>p(171)(68),Cin=>p(172)(68),clock=>clock,reset=>reset,s=>p(242)(68),cout=>p(243)(69));
FA_ff_7222:FAff port map(x=>p(170)(69),y=>p(171)(69),Cin=>p(172)(69),clock=>clock,reset=>reset,s=>p(242)(69),cout=>p(243)(70));
FA_ff_7223:FAff port map(x=>p(170)(70),y=>p(171)(70),Cin=>p(172)(70),clock=>clock,reset=>reset,s=>p(242)(70),cout=>p(243)(71));
FA_ff_7224:FAff port map(x=>p(170)(71),y=>p(171)(71),Cin=>p(172)(71),clock=>clock,reset=>reset,s=>p(242)(71),cout=>p(243)(72));
FA_ff_7225:FAff port map(x=>p(170)(72),y=>p(171)(72),Cin=>p(172)(72),clock=>clock,reset=>reset,s=>p(242)(72),cout=>p(243)(73));
FA_ff_7226:FAff port map(x=>p(170)(73),y=>p(171)(73),Cin=>p(172)(73),clock=>clock,reset=>reset,s=>p(242)(73),cout=>p(243)(74));
FA_ff_7227:FAff port map(x=>p(170)(74),y=>p(171)(74),Cin=>p(172)(74),clock=>clock,reset=>reset,s=>p(242)(74),cout=>p(243)(75));
FA_ff_7228:FAff port map(x=>p(170)(75),y=>p(171)(75),Cin=>p(172)(75),clock=>clock,reset=>reset,s=>p(242)(75),cout=>p(243)(76));
FA_ff_7229:FAff port map(x=>p(170)(76),y=>p(171)(76),Cin=>p(172)(76),clock=>clock,reset=>reset,s=>p(242)(76),cout=>p(243)(77));
FA_ff_7230:FAff port map(x=>p(170)(77),y=>p(171)(77),Cin=>p(172)(77),clock=>clock,reset=>reset,s=>p(242)(77),cout=>p(243)(78));
FA_ff_7231:FAff port map(x=>p(170)(78),y=>p(171)(78),Cin=>p(172)(78),clock=>clock,reset=>reset,s=>p(242)(78),cout=>p(243)(79));
FA_ff_7232:FAff port map(x=>p(170)(79),y=>p(171)(79),Cin=>p(172)(79),clock=>clock,reset=>reset,s=>p(242)(79),cout=>p(243)(80));
FA_ff_7233:FAff port map(x=>p(170)(80),y=>p(171)(80),Cin=>p(172)(80),clock=>clock,reset=>reset,s=>p(242)(80),cout=>p(243)(81));
FA_ff_7234:FAff port map(x=>p(170)(81),y=>p(171)(81),Cin=>p(172)(81),clock=>clock,reset=>reset,s=>p(242)(81),cout=>p(243)(82));
FA_ff_7235:FAff port map(x=>p(170)(82),y=>p(171)(82),Cin=>p(172)(82),clock=>clock,reset=>reset,s=>p(242)(82),cout=>p(243)(83));
FA_ff_7236:FAff port map(x=>p(170)(83),y=>p(171)(83),Cin=>p(172)(83),clock=>clock,reset=>reset,s=>p(242)(83),cout=>p(243)(84));
FA_ff_7237:FAff port map(x=>p(170)(84),y=>p(171)(84),Cin=>p(172)(84),clock=>clock,reset=>reset,s=>p(242)(84),cout=>p(243)(85));
FA_ff_7238:FAff port map(x=>p(170)(85),y=>p(171)(85),Cin=>p(172)(85),clock=>clock,reset=>reset,s=>p(242)(85),cout=>p(243)(86));
FA_ff_7239:FAff port map(x=>p(170)(86),y=>p(171)(86),Cin=>p(172)(86),clock=>clock,reset=>reset,s=>p(242)(86),cout=>p(243)(87));
FA_ff_7240:FAff port map(x=>p(170)(87),y=>p(171)(87),Cin=>p(172)(87),clock=>clock,reset=>reset,s=>p(242)(87),cout=>p(243)(88));
FA_ff_7241:FAff port map(x=>p(170)(88),y=>p(171)(88),Cin=>p(172)(88),clock=>clock,reset=>reset,s=>p(242)(88),cout=>p(243)(89));
FA_ff_7242:FAff port map(x=>p(170)(89),y=>p(171)(89),Cin=>p(172)(89),clock=>clock,reset=>reset,s=>p(242)(89),cout=>p(243)(90));
FA_ff_7243:FAff port map(x=>p(170)(90),y=>p(171)(90),Cin=>p(172)(90),clock=>clock,reset=>reset,s=>p(242)(90),cout=>p(243)(91));
FA_ff_7244:FAff port map(x=>p(170)(91),y=>p(171)(91),Cin=>p(172)(91),clock=>clock,reset=>reset,s=>p(242)(91),cout=>p(243)(92));
FA_ff_7245:FAff port map(x=>p(170)(92),y=>p(171)(92),Cin=>p(172)(92),clock=>clock,reset=>reset,s=>p(242)(92),cout=>p(243)(93));
FA_ff_7246:FAff port map(x=>p(170)(93),y=>p(171)(93),Cin=>p(172)(93),clock=>clock,reset=>reset,s=>p(242)(93),cout=>p(243)(94));
FA_ff_7247:FAff port map(x=>p(170)(94),y=>p(171)(94),Cin=>p(172)(94),clock=>clock,reset=>reset,s=>p(242)(94),cout=>p(243)(95));
FA_ff_7248:FAff port map(x=>p(170)(95),y=>p(171)(95),Cin=>p(172)(95),clock=>clock,reset=>reset,s=>p(242)(95),cout=>p(243)(96));
FA_ff_7249:FAff port map(x=>p(170)(96),y=>p(171)(96),Cin=>p(172)(96),clock=>clock,reset=>reset,s=>p(242)(96),cout=>p(243)(97));
FA_ff_7250:FAff port map(x=>p(170)(97),y=>p(171)(97),Cin=>p(172)(97),clock=>clock,reset=>reset,s=>p(242)(97),cout=>p(243)(98));
FA_ff_7251:FAff port map(x=>p(170)(98),y=>p(171)(98),Cin=>p(172)(98),clock=>clock,reset=>reset,s=>p(242)(98),cout=>p(243)(99));
FA_ff_7252:FAff port map(x=>p(170)(99),y=>p(171)(99),Cin=>p(172)(99),clock=>clock,reset=>reset,s=>p(242)(99),cout=>p(243)(100));
FA_ff_7253:FAff port map(x=>p(170)(100),y=>p(171)(100),Cin=>p(172)(100),clock=>clock,reset=>reset,s=>p(242)(100),cout=>p(243)(101));
FA_ff_7254:FAff port map(x=>p(170)(101),y=>p(171)(101),Cin=>p(172)(101),clock=>clock,reset=>reset,s=>p(242)(101),cout=>p(243)(102));
FA_ff_7255:FAff port map(x=>p(170)(102),y=>p(171)(102),Cin=>p(172)(102),clock=>clock,reset=>reset,s=>p(242)(102),cout=>p(243)(103));
FA_ff_7256:FAff port map(x=>p(170)(103),y=>p(171)(103),Cin=>p(172)(103),clock=>clock,reset=>reset,s=>p(242)(103),cout=>p(243)(104));
FA_ff_7257:FAff port map(x=>p(170)(104),y=>p(171)(104),Cin=>p(172)(104),clock=>clock,reset=>reset,s=>p(242)(104),cout=>p(243)(105));
FA_ff_7258:FAff port map(x=>p(170)(105),y=>p(171)(105),Cin=>p(172)(105),clock=>clock,reset=>reset,s=>p(242)(105),cout=>p(243)(106));
FA_ff_7259:FAff port map(x=>p(170)(106),y=>p(171)(106),Cin=>p(172)(106),clock=>clock,reset=>reset,s=>p(242)(106),cout=>p(243)(107));
FA_ff_7260:FAff port map(x=>p(170)(107),y=>p(171)(107),Cin=>p(172)(107),clock=>clock,reset=>reset,s=>p(242)(107),cout=>p(243)(108));
FA_ff_7261:FAff port map(x=>p(170)(108),y=>p(171)(108),Cin=>p(172)(108),clock=>clock,reset=>reset,s=>p(242)(108),cout=>p(243)(109));
FA_ff_7262:FAff port map(x=>p(170)(109),y=>p(171)(109),Cin=>p(172)(109),clock=>clock,reset=>reset,s=>p(242)(109),cout=>p(243)(110));
FA_ff_7263:FAff port map(x=>p(170)(110),y=>p(171)(110),Cin=>p(172)(110),clock=>clock,reset=>reset,s=>p(242)(110),cout=>p(243)(111));
FA_ff_7264:FAff port map(x=>p(170)(111),y=>p(171)(111),Cin=>p(172)(111),clock=>clock,reset=>reset,s=>p(242)(111),cout=>p(243)(112));
FA_ff_7265:FAff port map(x=>p(170)(112),y=>p(171)(112),Cin=>p(172)(112),clock=>clock,reset=>reset,s=>p(242)(112),cout=>p(243)(113));
FA_ff_7266:FAff port map(x=>p(170)(113),y=>p(171)(113),Cin=>p(172)(113),clock=>clock,reset=>reset,s=>p(242)(113),cout=>p(243)(114));
FA_ff_7267:FAff port map(x=>p(170)(114),y=>p(171)(114),Cin=>p(172)(114),clock=>clock,reset=>reset,s=>p(242)(114),cout=>p(243)(115));
FA_ff_7268:FAff port map(x=>p(170)(115),y=>p(171)(115),Cin=>p(172)(115),clock=>clock,reset=>reset,s=>p(242)(115),cout=>p(243)(116));
FA_ff_7269:FAff port map(x=>p(170)(116),y=>p(171)(116),Cin=>p(172)(116),clock=>clock,reset=>reset,s=>p(242)(116),cout=>p(243)(117));
FA_ff_7270:FAff port map(x=>p(170)(117),y=>p(171)(117),Cin=>p(172)(117),clock=>clock,reset=>reset,s=>p(242)(117),cout=>p(243)(118));
FA_ff_7271:FAff port map(x=>p(170)(118),y=>p(171)(118),Cin=>p(172)(118),clock=>clock,reset=>reset,s=>p(242)(118),cout=>p(243)(119));
FA_ff_7272:FAff port map(x=>p(170)(119),y=>p(171)(119),Cin=>p(172)(119),clock=>clock,reset=>reset,s=>p(242)(119),cout=>p(243)(120));
FA_ff_7273:FAff port map(x=>p(170)(120),y=>p(171)(120),Cin=>p(172)(120),clock=>clock,reset=>reset,s=>p(242)(120),cout=>p(243)(121));
FA_ff_7274:FAff port map(x=>p(170)(121),y=>p(171)(121),Cin=>p(172)(121),clock=>clock,reset=>reset,s=>p(242)(121),cout=>p(243)(122));
FA_ff_7275:FAff port map(x=>p(170)(122),y=>p(171)(122),Cin=>p(172)(122),clock=>clock,reset=>reset,s=>p(242)(122),cout=>p(243)(123));
FA_ff_7276:FAff port map(x=>p(170)(123),y=>p(171)(123),Cin=>p(172)(123),clock=>clock,reset=>reset,s=>p(242)(123),cout=>p(243)(124));
FA_ff_7277:FAff port map(x=>p(170)(124),y=>p(171)(124),Cin=>p(172)(124),clock=>clock,reset=>reset,s=>p(242)(124),cout=>p(243)(125));
FA_ff_7278:FAff port map(x=>p(170)(125),y=>p(171)(125),Cin=>p(172)(125),clock=>clock,reset=>reset,s=>p(242)(125),cout=>p(243)(126));
FA_ff_7279:FAff port map(x=>p(170)(126),y=>p(171)(126),Cin=>p(172)(126),clock=>clock,reset=>reset,s=>p(242)(126),cout=>p(243)(127));
FA_ff_7280:FAff port map(x=>p(170)(127),y=>p(171)(127),Cin=>p(172)(127),clock=>clock,reset=>reset,s=>p(242)(127),cout=>p(243)(128));
p(242)(128)<=p(171)(128);
p(244)(0)<=p(174)(0);
FA_ff_7281:FAff port map(x=>p(173)(1),y=>p(174)(1),Cin=>p(175)(1),clock=>clock,reset=>reset,s=>p(244)(1),cout=>p(245)(2));
FA_ff_7282:FAff port map(x=>p(173)(2),y=>p(174)(2),Cin=>p(175)(2),clock=>clock,reset=>reset,s=>p(244)(2),cout=>p(245)(3));
FA_ff_7283:FAff port map(x=>p(173)(3),y=>p(174)(3),Cin=>p(175)(3),clock=>clock,reset=>reset,s=>p(244)(3),cout=>p(245)(4));
FA_ff_7284:FAff port map(x=>p(173)(4),y=>p(174)(4),Cin=>p(175)(4),clock=>clock,reset=>reset,s=>p(244)(4),cout=>p(245)(5));
FA_ff_7285:FAff port map(x=>p(173)(5),y=>p(174)(5),Cin=>p(175)(5),clock=>clock,reset=>reset,s=>p(244)(5),cout=>p(245)(6));
FA_ff_7286:FAff port map(x=>p(173)(6),y=>p(174)(6),Cin=>p(175)(6),clock=>clock,reset=>reset,s=>p(244)(6),cout=>p(245)(7));
FA_ff_7287:FAff port map(x=>p(173)(7),y=>p(174)(7),Cin=>p(175)(7),clock=>clock,reset=>reset,s=>p(244)(7),cout=>p(245)(8));
FA_ff_7288:FAff port map(x=>p(173)(8),y=>p(174)(8),Cin=>p(175)(8),clock=>clock,reset=>reset,s=>p(244)(8),cout=>p(245)(9));
FA_ff_7289:FAff port map(x=>p(173)(9),y=>p(174)(9),Cin=>p(175)(9),clock=>clock,reset=>reset,s=>p(244)(9),cout=>p(245)(10));
FA_ff_7290:FAff port map(x=>p(173)(10),y=>p(174)(10),Cin=>p(175)(10),clock=>clock,reset=>reset,s=>p(244)(10),cout=>p(245)(11));
FA_ff_7291:FAff port map(x=>p(173)(11),y=>p(174)(11),Cin=>p(175)(11),clock=>clock,reset=>reset,s=>p(244)(11),cout=>p(245)(12));
FA_ff_7292:FAff port map(x=>p(173)(12),y=>p(174)(12),Cin=>p(175)(12),clock=>clock,reset=>reset,s=>p(244)(12),cout=>p(245)(13));
FA_ff_7293:FAff port map(x=>p(173)(13),y=>p(174)(13),Cin=>p(175)(13),clock=>clock,reset=>reset,s=>p(244)(13),cout=>p(245)(14));
FA_ff_7294:FAff port map(x=>p(173)(14),y=>p(174)(14),Cin=>p(175)(14),clock=>clock,reset=>reset,s=>p(244)(14),cout=>p(245)(15));
FA_ff_7295:FAff port map(x=>p(173)(15),y=>p(174)(15),Cin=>p(175)(15),clock=>clock,reset=>reset,s=>p(244)(15),cout=>p(245)(16));
FA_ff_7296:FAff port map(x=>p(173)(16),y=>p(174)(16),Cin=>p(175)(16),clock=>clock,reset=>reset,s=>p(244)(16),cout=>p(245)(17));
FA_ff_7297:FAff port map(x=>p(173)(17),y=>p(174)(17),Cin=>p(175)(17),clock=>clock,reset=>reset,s=>p(244)(17),cout=>p(245)(18));
FA_ff_7298:FAff port map(x=>p(173)(18),y=>p(174)(18),Cin=>p(175)(18),clock=>clock,reset=>reset,s=>p(244)(18),cout=>p(245)(19));
FA_ff_7299:FAff port map(x=>p(173)(19),y=>p(174)(19),Cin=>p(175)(19),clock=>clock,reset=>reset,s=>p(244)(19),cout=>p(245)(20));
FA_ff_7300:FAff port map(x=>p(173)(20),y=>p(174)(20),Cin=>p(175)(20),clock=>clock,reset=>reset,s=>p(244)(20),cout=>p(245)(21));
FA_ff_7301:FAff port map(x=>p(173)(21),y=>p(174)(21),Cin=>p(175)(21),clock=>clock,reset=>reset,s=>p(244)(21),cout=>p(245)(22));
FA_ff_7302:FAff port map(x=>p(173)(22),y=>p(174)(22),Cin=>p(175)(22),clock=>clock,reset=>reset,s=>p(244)(22),cout=>p(245)(23));
FA_ff_7303:FAff port map(x=>p(173)(23),y=>p(174)(23),Cin=>p(175)(23),clock=>clock,reset=>reset,s=>p(244)(23),cout=>p(245)(24));
FA_ff_7304:FAff port map(x=>p(173)(24),y=>p(174)(24),Cin=>p(175)(24),clock=>clock,reset=>reset,s=>p(244)(24),cout=>p(245)(25));
FA_ff_7305:FAff port map(x=>p(173)(25),y=>p(174)(25),Cin=>p(175)(25),clock=>clock,reset=>reset,s=>p(244)(25),cout=>p(245)(26));
FA_ff_7306:FAff port map(x=>p(173)(26),y=>p(174)(26),Cin=>p(175)(26),clock=>clock,reset=>reset,s=>p(244)(26),cout=>p(245)(27));
FA_ff_7307:FAff port map(x=>p(173)(27),y=>p(174)(27),Cin=>p(175)(27),clock=>clock,reset=>reset,s=>p(244)(27),cout=>p(245)(28));
FA_ff_7308:FAff port map(x=>p(173)(28),y=>p(174)(28),Cin=>p(175)(28),clock=>clock,reset=>reset,s=>p(244)(28),cout=>p(245)(29));
FA_ff_7309:FAff port map(x=>p(173)(29),y=>p(174)(29),Cin=>p(175)(29),clock=>clock,reset=>reset,s=>p(244)(29),cout=>p(245)(30));
FA_ff_7310:FAff port map(x=>p(173)(30),y=>p(174)(30),Cin=>p(175)(30),clock=>clock,reset=>reset,s=>p(244)(30),cout=>p(245)(31));
FA_ff_7311:FAff port map(x=>p(173)(31),y=>p(174)(31),Cin=>p(175)(31),clock=>clock,reset=>reset,s=>p(244)(31),cout=>p(245)(32));
FA_ff_7312:FAff port map(x=>p(173)(32),y=>p(174)(32),Cin=>p(175)(32),clock=>clock,reset=>reset,s=>p(244)(32),cout=>p(245)(33));
FA_ff_7313:FAff port map(x=>p(173)(33),y=>p(174)(33),Cin=>p(175)(33),clock=>clock,reset=>reset,s=>p(244)(33),cout=>p(245)(34));
FA_ff_7314:FAff port map(x=>p(173)(34),y=>p(174)(34),Cin=>p(175)(34),clock=>clock,reset=>reset,s=>p(244)(34),cout=>p(245)(35));
FA_ff_7315:FAff port map(x=>p(173)(35),y=>p(174)(35),Cin=>p(175)(35),clock=>clock,reset=>reset,s=>p(244)(35),cout=>p(245)(36));
FA_ff_7316:FAff port map(x=>p(173)(36),y=>p(174)(36),Cin=>p(175)(36),clock=>clock,reset=>reset,s=>p(244)(36),cout=>p(245)(37));
FA_ff_7317:FAff port map(x=>p(173)(37),y=>p(174)(37),Cin=>p(175)(37),clock=>clock,reset=>reset,s=>p(244)(37),cout=>p(245)(38));
FA_ff_7318:FAff port map(x=>p(173)(38),y=>p(174)(38),Cin=>p(175)(38),clock=>clock,reset=>reset,s=>p(244)(38),cout=>p(245)(39));
FA_ff_7319:FAff port map(x=>p(173)(39),y=>p(174)(39),Cin=>p(175)(39),clock=>clock,reset=>reset,s=>p(244)(39),cout=>p(245)(40));
FA_ff_7320:FAff port map(x=>p(173)(40),y=>p(174)(40),Cin=>p(175)(40),clock=>clock,reset=>reset,s=>p(244)(40),cout=>p(245)(41));
FA_ff_7321:FAff port map(x=>p(173)(41),y=>p(174)(41),Cin=>p(175)(41),clock=>clock,reset=>reset,s=>p(244)(41),cout=>p(245)(42));
FA_ff_7322:FAff port map(x=>p(173)(42),y=>p(174)(42),Cin=>p(175)(42),clock=>clock,reset=>reset,s=>p(244)(42),cout=>p(245)(43));
FA_ff_7323:FAff port map(x=>p(173)(43),y=>p(174)(43),Cin=>p(175)(43),clock=>clock,reset=>reset,s=>p(244)(43),cout=>p(245)(44));
FA_ff_7324:FAff port map(x=>p(173)(44),y=>p(174)(44),Cin=>p(175)(44),clock=>clock,reset=>reset,s=>p(244)(44),cout=>p(245)(45));
FA_ff_7325:FAff port map(x=>p(173)(45),y=>p(174)(45),Cin=>p(175)(45),clock=>clock,reset=>reset,s=>p(244)(45),cout=>p(245)(46));
FA_ff_7326:FAff port map(x=>p(173)(46),y=>p(174)(46),Cin=>p(175)(46),clock=>clock,reset=>reset,s=>p(244)(46),cout=>p(245)(47));
FA_ff_7327:FAff port map(x=>p(173)(47),y=>p(174)(47),Cin=>p(175)(47),clock=>clock,reset=>reset,s=>p(244)(47),cout=>p(245)(48));
FA_ff_7328:FAff port map(x=>p(173)(48),y=>p(174)(48),Cin=>p(175)(48),clock=>clock,reset=>reset,s=>p(244)(48),cout=>p(245)(49));
FA_ff_7329:FAff port map(x=>p(173)(49),y=>p(174)(49),Cin=>p(175)(49),clock=>clock,reset=>reset,s=>p(244)(49),cout=>p(245)(50));
FA_ff_7330:FAff port map(x=>p(173)(50),y=>p(174)(50),Cin=>p(175)(50),clock=>clock,reset=>reset,s=>p(244)(50),cout=>p(245)(51));
FA_ff_7331:FAff port map(x=>p(173)(51),y=>p(174)(51),Cin=>p(175)(51),clock=>clock,reset=>reset,s=>p(244)(51),cout=>p(245)(52));
FA_ff_7332:FAff port map(x=>p(173)(52),y=>p(174)(52),Cin=>p(175)(52),clock=>clock,reset=>reset,s=>p(244)(52),cout=>p(245)(53));
FA_ff_7333:FAff port map(x=>p(173)(53),y=>p(174)(53),Cin=>p(175)(53),clock=>clock,reset=>reset,s=>p(244)(53),cout=>p(245)(54));
FA_ff_7334:FAff port map(x=>p(173)(54),y=>p(174)(54),Cin=>p(175)(54),clock=>clock,reset=>reset,s=>p(244)(54),cout=>p(245)(55));
FA_ff_7335:FAff port map(x=>p(173)(55),y=>p(174)(55),Cin=>p(175)(55),clock=>clock,reset=>reset,s=>p(244)(55),cout=>p(245)(56));
FA_ff_7336:FAff port map(x=>p(173)(56),y=>p(174)(56),Cin=>p(175)(56),clock=>clock,reset=>reset,s=>p(244)(56),cout=>p(245)(57));
FA_ff_7337:FAff port map(x=>p(173)(57),y=>p(174)(57),Cin=>p(175)(57),clock=>clock,reset=>reset,s=>p(244)(57),cout=>p(245)(58));
FA_ff_7338:FAff port map(x=>p(173)(58),y=>p(174)(58),Cin=>p(175)(58),clock=>clock,reset=>reset,s=>p(244)(58),cout=>p(245)(59));
FA_ff_7339:FAff port map(x=>p(173)(59),y=>p(174)(59),Cin=>p(175)(59),clock=>clock,reset=>reset,s=>p(244)(59),cout=>p(245)(60));
FA_ff_7340:FAff port map(x=>p(173)(60),y=>p(174)(60),Cin=>p(175)(60),clock=>clock,reset=>reset,s=>p(244)(60),cout=>p(245)(61));
FA_ff_7341:FAff port map(x=>p(173)(61),y=>p(174)(61),Cin=>p(175)(61),clock=>clock,reset=>reset,s=>p(244)(61),cout=>p(245)(62));
FA_ff_7342:FAff port map(x=>p(173)(62),y=>p(174)(62),Cin=>p(175)(62),clock=>clock,reset=>reset,s=>p(244)(62),cout=>p(245)(63));
FA_ff_7343:FAff port map(x=>p(173)(63),y=>p(174)(63),Cin=>p(175)(63),clock=>clock,reset=>reset,s=>p(244)(63),cout=>p(245)(64));
FA_ff_7344:FAff port map(x=>p(173)(64),y=>p(174)(64),Cin=>p(175)(64),clock=>clock,reset=>reset,s=>p(244)(64),cout=>p(245)(65));
FA_ff_7345:FAff port map(x=>p(173)(65),y=>p(174)(65),Cin=>p(175)(65),clock=>clock,reset=>reset,s=>p(244)(65),cout=>p(245)(66));
FA_ff_7346:FAff port map(x=>p(173)(66),y=>p(174)(66),Cin=>p(175)(66),clock=>clock,reset=>reset,s=>p(244)(66),cout=>p(245)(67));
FA_ff_7347:FAff port map(x=>p(173)(67),y=>p(174)(67),Cin=>p(175)(67),clock=>clock,reset=>reset,s=>p(244)(67),cout=>p(245)(68));
FA_ff_7348:FAff port map(x=>p(173)(68),y=>p(174)(68),Cin=>p(175)(68),clock=>clock,reset=>reset,s=>p(244)(68),cout=>p(245)(69));
FA_ff_7349:FAff port map(x=>p(173)(69),y=>p(174)(69),Cin=>p(175)(69),clock=>clock,reset=>reset,s=>p(244)(69),cout=>p(245)(70));
FA_ff_7350:FAff port map(x=>p(173)(70),y=>p(174)(70),Cin=>p(175)(70),clock=>clock,reset=>reset,s=>p(244)(70),cout=>p(245)(71));
FA_ff_7351:FAff port map(x=>p(173)(71),y=>p(174)(71),Cin=>p(175)(71),clock=>clock,reset=>reset,s=>p(244)(71),cout=>p(245)(72));
FA_ff_7352:FAff port map(x=>p(173)(72),y=>p(174)(72),Cin=>p(175)(72),clock=>clock,reset=>reset,s=>p(244)(72),cout=>p(245)(73));
FA_ff_7353:FAff port map(x=>p(173)(73),y=>p(174)(73),Cin=>p(175)(73),clock=>clock,reset=>reset,s=>p(244)(73),cout=>p(245)(74));
FA_ff_7354:FAff port map(x=>p(173)(74),y=>p(174)(74),Cin=>p(175)(74),clock=>clock,reset=>reset,s=>p(244)(74),cout=>p(245)(75));
FA_ff_7355:FAff port map(x=>p(173)(75),y=>p(174)(75),Cin=>p(175)(75),clock=>clock,reset=>reset,s=>p(244)(75),cout=>p(245)(76));
FA_ff_7356:FAff port map(x=>p(173)(76),y=>p(174)(76),Cin=>p(175)(76),clock=>clock,reset=>reset,s=>p(244)(76),cout=>p(245)(77));
FA_ff_7357:FAff port map(x=>p(173)(77),y=>p(174)(77),Cin=>p(175)(77),clock=>clock,reset=>reset,s=>p(244)(77),cout=>p(245)(78));
FA_ff_7358:FAff port map(x=>p(173)(78),y=>p(174)(78),Cin=>p(175)(78),clock=>clock,reset=>reset,s=>p(244)(78),cout=>p(245)(79));
FA_ff_7359:FAff port map(x=>p(173)(79),y=>p(174)(79),Cin=>p(175)(79),clock=>clock,reset=>reset,s=>p(244)(79),cout=>p(245)(80));
FA_ff_7360:FAff port map(x=>p(173)(80),y=>p(174)(80),Cin=>p(175)(80),clock=>clock,reset=>reset,s=>p(244)(80),cout=>p(245)(81));
FA_ff_7361:FAff port map(x=>p(173)(81),y=>p(174)(81),Cin=>p(175)(81),clock=>clock,reset=>reset,s=>p(244)(81),cout=>p(245)(82));
FA_ff_7362:FAff port map(x=>p(173)(82),y=>p(174)(82),Cin=>p(175)(82),clock=>clock,reset=>reset,s=>p(244)(82),cout=>p(245)(83));
FA_ff_7363:FAff port map(x=>p(173)(83),y=>p(174)(83),Cin=>p(175)(83),clock=>clock,reset=>reset,s=>p(244)(83),cout=>p(245)(84));
FA_ff_7364:FAff port map(x=>p(173)(84),y=>p(174)(84),Cin=>p(175)(84),clock=>clock,reset=>reset,s=>p(244)(84),cout=>p(245)(85));
FA_ff_7365:FAff port map(x=>p(173)(85),y=>p(174)(85),Cin=>p(175)(85),clock=>clock,reset=>reset,s=>p(244)(85),cout=>p(245)(86));
FA_ff_7366:FAff port map(x=>p(173)(86),y=>p(174)(86),Cin=>p(175)(86),clock=>clock,reset=>reset,s=>p(244)(86),cout=>p(245)(87));
FA_ff_7367:FAff port map(x=>p(173)(87),y=>p(174)(87),Cin=>p(175)(87),clock=>clock,reset=>reset,s=>p(244)(87),cout=>p(245)(88));
FA_ff_7368:FAff port map(x=>p(173)(88),y=>p(174)(88),Cin=>p(175)(88),clock=>clock,reset=>reset,s=>p(244)(88),cout=>p(245)(89));
FA_ff_7369:FAff port map(x=>p(173)(89),y=>p(174)(89),Cin=>p(175)(89),clock=>clock,reset=>reset,s=>p(244)(89),cout=>p(245)(90));
FA_ff_7370:FAff port map(x=>p(173)(90),y=>p(174)(90),Cin=>p(175)(90),clock=>clock,reset=>reset,s=>p(244)(90),cout=>p(245)(91));
FA_ff_7371:FAff port map(x=>p(173)(91),y=>p(174)(91),Cin=>p(175)(91),clock=>clock,reset=>reset,s=>p(244)(91),cout=>p(245)(92));
FA_ff_7372:FAff port map(x=>p(173)(92),y=>p(174)(92),Cin=>p(175)(92),clock=>clock,reset=>reset,s=>p(244)(92),cout=>p(245)(93));
FA_ff_7373:FAff port map(x=>p(173)(93),y=>p(174)(93),Cin=>p(175)(93),clock=>clock,reset=>reset,s=>p(244)(93),cout=>p(245)(94));
FA_ff_7374:FAff port map(x=>p(173)(94),y=>p(174)(94),Cin=>p(175)(94),clock=>clock,reset=>reset,s=>p(244)(94),cout=>p(245)(95));
FA_ff_7375:FAff port map(x=>p(173)(95),y=>p(174)(95),Cin=>p(175)(95),clock=>clock,reset=>reset,s=>p(244)(95),cout=>p(245)(96));
FA_ff_7376:FAff port map(x=>p(173)(96),y=>p(174)(96),Cin=>p(175)(96),clock=>clock,reset=>reset,s=>p(244)(96),cout=>p(245)(97));
FA_ff_7377:FAff port map(x=>p(173)(97),y=>p(174)(97),Cin=>p(175)(97),clock=>clock,reset=>reset,s=>p(244)(97),cout=>p(245)(98));
FA_ff_7378:FAff port map(x=>p(173)(98),y=>p(174)(98),Cin=>p(175)(98),clock=>clock,reset=>reset,s=>p(244)(98),cout=>p(245)(99));
FA_ff_7379:FAff port map(x=>p(173)(99),y=>p(174)(99),Cin=>p(175)(99),clock=>clock,reset=>reset,s=>p(244)(99),cout=>p(245)(100));
FA_ff_7380:FAff port map(x=>p(173)(100),y=>p(174)(100),Cin=>p(175)(100),clock=>clock,reset=>reset,s=>p(244)(100),cout=>p(245)(101));
FA_ff_7381:FAff port map(x=>p(173)(101),y=>p(174)(101),Cin=>p(175)(101),clock=>clock,reset=>reset,s=>p(244)(101),cout=>p(245)(102));
FA_ff_7382:FAff port map(x=>p(173)(102),y=>p(174)(102),Cin=>p(175)(102),clock=>clock,reset=>reset,s=>p(244)(102),cout=>p(245)(103));
FA_ff_7383:FAff port map(x=>p(173)(103),y=>p(174)(103),Cin=>p(175)(103),clock=>clock,reset=>reset,s=>p(244)(103),cout=>p(245)(104));
FA_ff_7384:FAff port map(x=>p(173)(104),y=>p(174)(104),Cin=>p(175)(104),clock=>clock,reset=>reset,s=>p(244)(104),cout=>p(245)(105));
FA_ff_7385:FAff port map(x=>p(173)(105),y=>p(174)(105),Cin=>p(175)(105),clock=>clock,reset=>reset,s=>p(244)(105),cout=>p(245)(106));
FA_ff_7386:FAff port map(x=>p(173)(106),y=>p(174)(106),Cin=>p(175)(106),clock=>clock,reset=>reset,s=>p(244)(106),cout=>p(245)(107));
FA_ff_7387:FAff port map(x=>p(173)(107),y=>p(174)(107),Cin=>p(175)(107),clock=>clock,reset=>reset,s=>p(244)(107),cout=>p(245)(108));
FA_ff_7388:FAff port map(x=>p(173)(108),y=>p(174)(108),Cin=>p(175)(108),clock=>clock,reset=>reset,s=>p(244)(108),cout=>p(245)(109));
FA_ff_7389:FAff port map(x=>p(173)(109),y=>p(174)(109),Cin=>p(175)(109),clock=>clock,reset=>reset,s=>p(244)(109),cout=>p(245)(110));
FA_ff_7390:FAff port map(x=>p(173)(110),y=>p(174)(110),Cin=>p(175)(110),clock=>clock,reset=>reset,s=>p(244)(110),cout=>p(245)(111));
FA_ff_7391:FAff port map(x=>p(173)(111),y=>p(174)(111),Cin=>p(175)(111),clock=>clock,reset=>reset,s=>p(244)(111),cout=>p(245)(112));
FA_ff_7392:FAff port map(x=>p(173)(112),y=>p(174)(112),Cin=>p(175)(112),clock=>clock,reset=>reset,s=>p(244)(112),cout=>p(245)(113));
FA_ff_7393:FAff port map(x=>p(173)(113),y=>p(174)(113),Cin=>p(175)(113),clock=>clock,reset=>reset,s=>p(244)(113),cout=>p(245)(114));
FA_ff_7394:FAff port map(x=>p(173)(114),y=>p(174)(114),Cin=>p(175)(114),clock=>clock,reset=>reset,s=>p(244)(114),cout=>p(245)(115));
FA_ff_7395:FAff port map(x=>p(173)(115),y=>p(174)(115),Cin=>p(175)(115),clock=>clock,reset=>reset,s=>p(244)(115),cout=>p(245)(116));
FA_ff_7396:FAff port map(x=>p(173)(116),y=>p(174)(116),Cin=>p(175)(116),clock=>clock,reset=>reset,s=>p(244)(116),cout=>p(245)(117));
FA_ff_7397:FAff port map(x=>p(173)(117),y=>p(174)(117),Cin=>p(175)(117),clock=>clock,reset=>reset,s=>p(244)(117),cout=>p(245)(118));
FA_ff_7398:FAff port map(x=>p(173)(118),y=>p(174)(118),Cin=>p(175)(118),clock=>clock,reset=>reset,s=>p(244)(118),cout=>p(245)(119));
FA_ff_7399:FAff port map(x=>p(173)(119),y=>p(174)(119),Cin=>p(175)(119),clock=>clock,reset=>reset,s=>p(244)(119),cout=>p(245)(120));
FA_ff_7400:FAff port map(x=>p(173)(120),y=>p(174)(120),Cin=>p(175)(120),clock=>clock,reset=>reset,s=>p(244)(120),cout=>p(245)(121));
FA_ff_7401:FAff port map(x=>p(173)(121),y=>p(174)(121),Cin=>p(175)(121),clock=>clock,reset=>reset,s=>p(244)(121),cout=>p(245)(122));
FA_ff_7402:FAff port map(x=>p(173)(122),y=>p(174)(122),Cin=>p(175)(122),clock=>clock,reset=>reset,s=>p(244)(122),cout=>p(245)(123));
FA_ff_7403:FAff port map(x=>p(173)(123),y=>p(174)(123),Cin=>p(175)(123),clock=>clock,reset=>reset,s=>p(244)(123),cout=>p(245)(124));
FA_ff_7404:FAff port map(x=>p(173)(124),y=>p(174)(124),Cin=>p(175)(124),clock=>clock,reset=>reset,s=>p(244)(124),cout=>p(245)(125));
FA_ff_7405:FAff port map(x=>p(173)(125),y=>p(174)(125),Cin=>p(175)(125),clock=>clock,reset=>reset,s=>p(244)(125),cout=>p(245)(126));
FA_ff_7406:FAff port map(x=>p(173)(126),y=>p(174)(126),Cin=>p(175)(126),clock=>clock,reset=>reset,s=>p(244)(126),cout=>p(245)(127));
FA_ff_7407:FAff port map(x=>p(173)(127),y=>p(174)(127),Cin=>p(175)(127),clock=>clock,reset=>reset,s=>p(244)(127),cout=>p(245)(128));
HA_ff_15:HAff port map(x=>p(173)(128),y=>p(175)(128),clock=>clock,reset=>reset,s=>p(244)(128),c=>p(245)(129));
HA_ff_16:HAff port map(x=>p(176)(0),y=>p(178)(0),clock=>clock,reset=>reset,s=>p(246)(0),c=>p(247)(1));
FA_ff_7408:FAff port map(x=>p(176)(1),y=>p(177)(1),Cin=>p(178)(1),clock=>clock,reset=>reset,s=>p(246)(1),cout=>p(247)(2));
FA_ff_7409:FAff port map(x=>p(176)(2),y=>p(177)(2),Cin=>p(178)(2),clock=>clock,reset=>reset,s=>p(246)(2),cout=>p(247)(3));
FA_ff_7410:FAff port map(x=>p(176)(3),y=>p(177)(3),Cin=>p(178)(3),clock=>clock,reset=>reset,s=>p(246)(3),cout=>p(247)(4));
FA_ff_7411:FAff port map(x=>p(176)(4),y=>p(177)(4),Cin=>p(178)(4),clock=>clock,reset=>reset,s=>p(246)(4),cout=>p(247)(5));
FA_ff_7412:FAff port map(x=>p(176)(5),y=>p(177)(5),Cin=>p(178)(5),clock=>clock,reset=>reset,s=>p(246)(5),cout=>p(247)(6));
FA_ff_7413:FAff port map(x=>p(176)(6),y=>p(177)(6),Cin=>p(178)(6),clock=>clock,reset=>reset,s=>p(246)(6),cout=>p(247)(7));
FA_ff_7414:FAff port map(x=>p(176)(7),y=>p(177)(7),Cin=>p(178)(7),clock=>clock,reset=>reset,s=>p(246)(7),cout=>p(247)(8));
FA_ff_7415:FAff port map(x=>p(176)(8),y=>p(177)(8),Cin=>p(178)(8),clock=>clock,reset=>reset,s=>p(246)(8),cout=>p(247)(9));
FA_ff_7416:FAff port map(x=>p(176)(9),y=>p(177)(9),Cin=>p(178)(9),clock=>clock,reset=>reset,s=>p(246)(9),cout=>p(247)(10));
FA_ff_7417:FAff port map(x=>p(176)(10),y=>p(177)(10),Cin=>p(178)(10),clock=>clock,reset=>reset,s=>p(246)(10),cout=>p(247)(11));
FA_ff_7418:FAff port map(x=>p(176)(11),y=>p(177)(11),Cin=>p(178)(11),clock=>clock,reset=>reset,s=>p(246)(11),cout=>p(247)(12));
FA_ff_7419:FAff port map(x=>p(176)(12),y=>p(177)(12),Cin=>p(178)(12),clock=>clock,reset=>reset,s=>p(246)(12),cout=>p(247)(13));
FA_ff_7420:FAff port map(x=>p(176)(13),y=>p(177)(13),Cin=>p(178)(13),clock=>clock,reset=>reset,s=>p(246)(13),cout=>p(247)(14));
FA_ff_7421:FAff port map(x=>p(176)(14),y=>p(177)(14),Cin=>p(178)(14),clock=>clock,reset=>reset,s=>p(246)(14),cout=>p(247)(15));
FA_ff_7422:FAff port map(x=>p(176)(15),y=>p(177)(15),Cin=>p(178)(15),clock=>clock,reset=>reset,s=>p(246)(15),cout=>p(247)(16));
FA_ff_7423:FAff port map(x=>p(176)(16),y=>p(177)(16),Cin=>p(178)(16),clock=>clock,reset=>reset,s=>p(246)(16),cout=>p(247)(17));
FA_ff_7424:FAff port map(x=>p(176)(17),y=>p(177)(17),Cin=>p(178)(17),clock=>clock,reset=>reset,s=>p(246)(17),cout=>p(247)(18));
FA_ff_7425:FAff port map(x=>p(176)(18),y=>p(177)(18),Cin=>p(178)(18),clock=>clock,reset=>reset,s=>p(246)(18),cout=>p(247)(19));
FA_ff_7426:FAff port map(x=>p(176)(19),y=>p(177)(19),Cin=>p(178)(19),clock=>clock,reset=>reset,s=>p(246)(19),cout=>p(247)(20));
FA_ff_7427:FAff port map(x=>p(176)(20),y=>p(177)(20),Cin=>p(178)(20),clock=>clock,reset=>reset,s=>p(246)(20),cout=>p(247)(21));
FA_ff_7428:FAff port map(x=>p(176)(21),y=>p(177)(21),Cin=>p(178)(21),clock=>clock,reset=>reset,s=>p(246)(21),cout=>p(247)(22));
FA_ff_7429:FAff port map(x=>p(176)(22),y=>p(177)(22),Cin=>p(178)(22),clock=>clock,reset=>reset,s=>p(246)(22),cout=>p(247)(23));
FA_ff_7430:FAff port map(x=>p(176)(23),y=>p(177)(23),Cin=>p(178)(23),clock=>clock,reset=>reset,s=>p(246)(23),cout=>p(247)(24));
FA_ff_7431:FAff port map(x=>p(176)(24),y=>p(177)(24),Cin=>p(178)(24),clock=>clock,reset=>reset,s=>p(246)(24),cout=>p(247)(25));
FA_ff_7432:FAff port map(x=>p(176)(25),y=>p(177)(25),Cin=>p(178)(25),clock=>clock,reset=>reset,s=>p(246)(25),cout=>p(247)(26));
FA_ff_7433:FAff port map(x=>p(176)(26),y=>p(177)(26),Cin=>p(178)(26),clock=>clock,reset=>reset,s=>p(246)(26),cout=>p(247)(27));
FA_ff_7434:FAff port map(x=>p(176)(27),y=>p(177)(27),Cin=>p(178)(27),clock=>clock,reset=>reset,s=>p(246)(27),cout=>p(247)(28));
FA_ff_7435:FAff port map(x=>p(176)(28),y=>p(177)(28),Cin=>p(178)(28),clock=>clock,reset=>reset,s=>p(246)(28),cout=>p(247)(29));
FA_ff_7436:FAff port map(x=>p(176)(29),y=>p(177)(29),Cin=>p(178)(29),clock=>clock,reset=>reset,s=>p(246)(29),cout=>p(247)(30));
FA_ff_7437:FAff port map(x=>p(176)(30),y=>p(177)(30),Cin=>p(178)(30),clock=>clock,reset=>reset,s=>p(246)(30),cout=>p(247)(31));
FA_ff_7438:FAff port map(x=>p(176)(31),y=>p(177)(31),Cin=>p(178)(31),clock=>clock,reset=>reset,s=>p(246)(31),cout=>p(247)(32));
FA_ff_7439:FAff port map(x=>p(176)(32),y=>p(177)(32),Cin=>p(178)(32),clock=>clock,reset=>reset,s=>p(246)(32),cout=>p(247)(33));
FA_ff_7440:FAff port map(x=>p(176)(33),y=>p(177)(33),Cin=>p(178)(33),clock=>clock,reset=>reset,s=>p(246)(33),cout=>p(247)(34));
FA_ff_7441:FAff port map(x=>p(176)(34),y=>p(177)(34),Cin=>p(178)(34),clock=>clock,reset=>reset,s=>p(246)(34),cout=>p(247)(35));
FA_ff_7442:FAff port map(x=>p(176)(35),y=>p(177)(35),Cin=>p(178)(35),clock=>clock,reset=>reset,s=>p(246)(35),cout=>p(247)(36));
FA_ff_7443:FAff port map(x=>p(176)(36),y=>p(177)(36),Cin=>p(178)(36),clock=>clock,reset=>reset,s=>p(246)(36),cout=>p(247)(37));
FA_ff_7444:FAff port map(x=>p(176)(37),y=>p(177)(37),Cin=>p(178)(37),clock=>clock,reset=>reset,s=>p(246)(37),cout=>p(247)(38));
FA_ff_7445:FAff port map(x=>p(176)(38),y=>p(177)(38),Cin=>p(178)(38),clock=>clock,reset=>reset,s=>p(246)(38),cout=>p(247)(39));
FA_ff_7446:FAff port map(x=>p(176)(39),y=>p(177)(39),Cin=>p(178)(39),clock=>clock,reset=>reset,s=>p(246)(39),cout=>p(247)(40));
FA_ff_7447:FAff port map(x=>p(176)(40),y=>p(177)(40),Cin=>p(178)(40),clock=>clock,reset=>reset,s=>p(246)(40),cout=>p(247)(41));
FA_ff_7448:FAff port map(x=>p(176)(41),y=>p(177)(41),Cin=>p(178)(41),clock=>clock,reset=>reset,s=>p(246)(41),cout=>p(247)(42));
FA_ff_7449:FAff port map(x=>p(176)(42),y=>p(177)(42),Cin=>p(178)(42),clock=>clock,reset=>reset,s=>p(246)(42),cout=>p(247)(43));
FA_ff_7450:FAff port map(x=>p(176)(43),y=>p(177)(43),Cin=>p(178)(43),clock=>clock,reset=>reset,s=>p(246)(43),cout=>p(247)(44));
FA_ff_7451:FAff port map(x=>p(176)(44),y=>p(177)(44),Cin=>p(178)(44),clock=>clock,reset=>reset,s=>p(246)(44),cout=>p(247)(45));
FA_ff_7452:FAff port map(x=>p(176)(45),y=>p(177)(45),Cin=>p(178)(45),clock=>clock,reset=>reset,s=>p(246)(45),cout=>p(247)(46));
FA_ff_7453:FAff port map(x=>p(176)(46),y=>p(177)(46),Cin=>p(178)(46),clock=>clock,reset=>reset,s=>p(246)(46),cout=>p(247)(47));
FA_ff_7454:FAff port map(x=>p(176)(47),y=>p(177)(47),Cin=>p(178)(47),clock=>clock,reset=>reset,s=>p(246)(47),cout=>p(247)(48));
FA_ff_7455:FAff port map(x=>p(176)(48),y=>p(177)(48),Cin=>p(178)(48),clock=>clock,reset=>reset,s=>p(246)(48),cout=>p(247)(49));
FA_ff_7456:FAff port map(x=>p(176)(49),y=>p(177)(49),Cin=>p(178)(49),clock=>clock,reset=>reset,s=>p(246)(49),cout=>p(247)(50));
FA_ff_7457:FAff port map(x=>p(176)(50),y=>p(177)(50),Cin=>p(178)(50),clock=>clock,reset=>reset,s=>p(246)(50),cout=>p(247)(51));
FA_ff_7458:FAff port map(x=>p(176)(51),y=>p(177)(51),Cin=>p(178)(51),clock=>clock,reset=>reset,s=>p(246)(51),cout=>p(247)(52));
FA_ff_7459:FAff port map(x=>p(176)(52),y=>p(177)(52),Cin=>p(178)(52),clock=>clock,reset=>reset,s=>p(246)(52),cout=>p(247)(53));
FA_ff_7460:FAff port map(x=>p(176)(53),y=>p(177)(53),Cin=>p(178)(53),clock=>clock,reset=>reset,s=>p(246)(53),cout=>p(247)(54));
FA_ff_7461:FAff port map(x=>p(176)(54),y=>p(177)(54),Cin=>p(178)(54),clock=>clock,reset=>reset,s=>p(246)(54),cout=>p(247)(55));
FA_ff_7462:FAff port map(x=>p(176)(55),y=>p(177)(55),Cin=>p(178)(55),clock=>clock,reset=>reset,s=>p(246)(55),cout=>p(247)(56));
FA_ff_7463:FAff port map(x=>p(176)(56),y=>p(177)(56),Cin=>p(178)(56),clock=>clock,reset=>reset,s=>p(246)(56),cout=>p(247)(57));
FA_ff_7464:FAff port map(x=>p(176)(57),y=>p(177)(57),Cin=>p(178)(57),clock=>clock,reset=>reset,s=>p(246)(57),cout=>p(247)(58));
FA_ff_7465:FAff port map(x=>p(176)(58),y=>p(177)(58),Cin=>p(178)(58),clock=>clock,reset=>reset,s=>p(246)(58),cout=>p(247)(59));
FA_ff_7466:FAff port map(x=>p(176)(59),y=>p(177)(59),Cin=>p(178)(59),clock=>clock,reset=>reset,s=>p(246)(59),cout=>p(247)(60));
FA_ff_7467:FAff port map(x=>p(176)(60),y=>p(177)(60),Cin=>p(178)(60),clock=>clock,reset=>reset,s=>p(246)(60),cout=>p(247)(61));
FA_ff_7468:FAff port map(x=>p(176)(61),y=>p(177)(61),Cin=>p(178)(61),clock=>clock,reset=>reset,s=>p(246)(61),cout=>p(247)(62));
FA_ff_7469:FAff port map(x=>p(176)(62),y=>p(177)(62),Cin=>p(178)(62),clock=>clock,reset=>reset,s=>p(246)(62),cout=>p(247)(63));
FA_ff_7470:FAff port map(x=>p(176)(63),y=>p(177)(63),Cin=>p(178)(63),clock=>clock,reset=>reset,s=>p(246)(63),cout=>p(247)(64));
FA_ff_7471:FAff port map(x=>p(176)(64),y=>p(177)(64),Cin=>p(178)(64),clock=>clock,reset=>reset,s=>p(246)(64),cout=>p(247)(65));
FA_ff_7472:FAff port map(x=>p(176)(65),y=>p(177)(65),Cin=>p(178)(65),clock=>clock,reset=>reset,s=>p(246)(65),cout=>p(247)(66));
FA_ff_7473:FAff port map(x=>p(176)(66),y=>p(177)(66),Cin=>p(178)(66),clock=>clock,reset=>reset,s=>p(246)(66),cout=>p(247)(67));
FA_ff_7474:FAff port map(x=>p(176)(67),y=>p(177)(67),Cin=>p(178)(67),clock=>clock,reset=>reset,s=>p(246)(67),cout=>p(247)(68));
FA_ff_7475:FAff port map(x=>p(176)(68),y=>p(177)(68),Cin=>p(178)(68),clock=>clock,reset=>reset,s=>p(246)(68),cout=>p(247)(69));
FA_ff_7476:FAff port map(x=>p(176)(69),y=>p(177)(69),Cin=>p(178)(69),clock=>clock,reset=>reset,s=>p(246)(69),cout=>p(247)(70));
FA_ff_7477:FAff port map(x=>p(176)(70),y=>p(177)(70),Cin=>p(178)(70),clock=>clock,reset=>reset,s=>p(246)(70),cout=>p(247)(71));
FA_ff_7478:FAff port map(x=>p(176)(71),y=>p(177)(71),Cin=>p(178)(71),clock=>clock,reset=>reset,s=>p(246)(71),cout=>p(247)(72));
FA_ff_7479:FAff port map(x=>p(176)(72),y=>p(177)(72),Cin=>p(178)(72),clock=>clock,reset=>reset,s=>p(246)(72),cout=>p(247)(73));
FA_ff_7480:FAff port map(x=>p(176)(73),y=>p(177)(73),Cin=>p(178)(73),clock=>clock,reset=>reset,s=>p(246)(73),cout=>p(247)(74));
FA_ff_7481:FAff port map(x=>p(176)(74),y=>p(177)(74),Cin=>p(178)(74),clock=>clock,reset=>reset,s=>p(246)(74),cout=>p(247)(75));
FA_ff_7482:FAff port map(x=>p(176)(75),y=>p(177)(75),Cin=>p(178)(75),clock=>clock,reset=>reset,s=>p(246)(75),cout=>p(247)(76));
FA_ff_7483:FAff port map(x=>p(176)(76),y=>p(177)(76),Cin=>p(178)(76),clock=>clock,reset=>reset,s=>p(246)(76),cout=>p(247)(77));
FA_ff_7484:FAff port map(x=>p(176)(77),y=>p(177)(77),Cin=>p(178)(77),clock=>clock,reset=>reset,s=>p(246)(77),cout=>p(247)(78));
FA_ff_7485:FAff port map(x=>p(176)(78),y=>p(177)(78),Cin=>p(178)(78),clock=>clock,reset=>reset,s=>p(246)(78),cout=>p(247)(79));
FA_ff_7486:FAff port map(x=>p(176)(79),y=>p(177)(79),Cin=>p(178)(79),clock=>clock,reset=>reset,s=>p(246)(79),cout=>p(247)(80));
FA_ff_7487:FAff port map(x=>p(176)(80),y=>p(177)(80),Cin=>p(178)(80),clock=>clock,reset=>reset,s=>p(246)(80),cout=>p(247)(81));
FA_ff_7488:FAff port map(x=>p(176)(81),y=>p(177)(81),Cin=>p(178)(81),clock=>clock,reset=>reset,s=>p(246)(81),cout=>p(247)(82));
FA_ff_7489:FAff port map(x=>p(176)(82),y=>p(177)(82),Cin=>p(178)(82),clock=>clock,reset=>reset,s=>p(246)(82),cout=>p(247)(83));
FA_ff_7490:FAff port map(x=>p(176)(83),y=>p(177)(83),Cin=>p(178)(83),clock=>clock,reset=>reset,s=>p(246)(83),cout=>p(247)(84));
FA_ff_7491:FAff port map(x=>p(176)(84),y=>p(177)(84),Cin=>p(178)(84),clock=>clock,reset=>reset,s=>p(246)(84),cout=>p(247)(85));
FA_ff_7492:FAff port map(x=>p(176)(85),y=>p(177)(85),Cin=>p(178)(85),clock=>clock,reset=>reset,s=>p(246)(85),cout=>p(247)(86));
FA_ff_7493:FAff port map(x=>p(176)(86),y=>p(177)(86),Cin=>p(178)(86),clock=>clock,reset=>reset,s=>p(246)(86),cout=>p(247)(87));
FA_ff_7494:FAff port map(x=>p(176)(87),y=>p(177)(87),Cin=>p(178)(87),clock=>clock,reset=>reset,s=>p(246)(87),cout=>p(247)(88));
FA_ff_7495:FAff port map(x=>p(176)(88),y=>p(177)(88),Cin=>p(178)(88),clock=>clock,reset=>reset,s=>p(246)(88),cout=>p(247)(89));
FA_ff_7496:FAff port map(x=>p(176)(89),y=>p(177)(89),Cin=>p(178)(89),clock=>clock,reset=>reset,s=>p(246)(89),cout=>p(247)(90));
FA_ff_7497:FAff port map(x=>p(176)(90),y=>p(177)(90),Cin=>p(178)(90),clock=>clock,reset=>reset,s=>p(246)(90),cout=>p(247)(91));
FA_ff_7498:FAff port map(x=>p(176)(91),y=>p(177)(91),Cin=>p(178)(91),clock=>clock,reset=>reset,s=>p(246)(91),cout=>p(247)(92));
FA_ff_7499:FAff port map(x=>p(176)(92),y=>p(177)(92),Cin=>p(178)(92),clock=>clock,reset=>reset,s=>p(246)(92),cout=>p(247)(93));
FA_ff_7500:FAff port map(x=>p(176)(93),y=>p(177)(93),Cin=>p(178)(93),clock=>clock,reset=>reset,s=>p(246)(93),cout=>p(247)(94));
FA_ff_7501:FAff port map(x=>p(176)(94),y=>p(177)(94),Cin=>p(178)(94),clock=>clock,reset=>reset,s=>p(246)(94),cout=>p(247)(95));
FA_ff_7502:FAff port map(x=>p(176)(95),y=>p(177)(95),Cin=>p(178)(95),clock=>clock,reset=>reset,s=>p(246)(95),cout=>p(247)(96));
FA_ff_7503:FAff port map(x=>p(176)(96),y=>p(177)(96),Cin=>p(178)(96),clock=>clock,reset=>reset,s=>p(246)(96),cout=>p(247)(97));
FA_ff_7504:FAff port map(x=>p(176)(97),y=>p(177)(97),Cin=>p(178)(97),clock=>clock,reset=>reset,s=>p(246)(97),cout=>p(247)(98));
FA_ff_7505:FAff port map(x=>p(176)(98),y=>p(177)(98),Cin=>p(178)(98),clock=>clock,reset=>reset,s=>p(246)(98),cout=>p(247)(99));
FA_ff_7506:FAff port map(x=>p(176)(99),y=>p(177)(99),Cin=>p(178)(99),clock=>clock,reset=>reset,s=>p(246)(99),cout=>p(247)(100));
FA_ff_7507:FAff port map(x=>p(176)(100),y=>p(177)(100),Cin=>p(178)(100),clock=>clock,reset=>reset,s=>p(246)(100),cout=>p(247)(101));
FA_ff_7508:FAff port map(x=>p(176)(101),y=>p(177)(101),Cin=>p(178)(101),clock=>clock,reset=>reset,s=>p(246)(101),cout=>p(247)(102));
FA_ff_7509:FAff port map(x=>p(176)(102),y=>p(177)(102),Cin=>p(178)(102),clock=>clock,reset=>reset,s=>p(246)(102),cout=>p(247)(103));
FA_ff_7510:FAff port map(x=>p(176)(103),y=>p(177)(103),Cin=>p(178)(103),clock=>clock,reset=>reset,s=>p(246)(103),cout=>p(247)(104));
FA_ff_7511:FAff port map(x=>p(176)(104),y=>p(177)(104),Cin=>p(178)(104),clock=>clock,reset=>reset,s=>p(246)(104),cout=>p(247)(105));
FA_ff_7512:FAff port map(x=>p(176)(105),y=>p(177)(105),Cin=>p(178)(105),clock=>clock,reset=>reset,s=>p(246)(105),cout=>p(247)(106));
FA_ff_7513:FAff port map(x=>p(176)(106),y=>p(177)(106),Cin=>p(178)(106),clock=>clock,reset=>reset,s=>p(246)(106),cout=>p(247)(107));
FA_ff_7514:FAff port map(x=>p(176)(107),y=>p(177)(107),Cin=>p(178)(107),clock=>clock,reset=>reset,s=>p(246)(107),cout=>p(247)(108));
FA_ff_7515:FAff port map(x=>p(176)(108),y=>p(177)(108),Cin=>p(178)(108),clock=>clock,reset=>reset,s=>p(246)(108),cout=>p(247)(109));
FA_ff_7516:FAff port map(x=>p(176)(109),y=>p(177)(109),Cin=>p(178)(109),clock=>clock,reset=>reset,s=>p(246)(109),cout=>p(247)(110));
FA_ff_7517:FAff port map(x=>p(176)(110),y=>p(177)(110),Cin=>p(178)(110),clock=>clock,reset=>reset,s=>p(246)(110),cout=>p(247)(111));
FA_ff_7518:FAff port map(x=>p(176)(111),y=>p(177)(111),Cin=>p(178)(111),clock=>clock,reset=>reset,s=>p(246)(111),cout=>p(247)(112));
FA_ff_7519:FAff port map(x=>p(176)(112),y=>p(177)(112),Cin=>p(178)(112),clock=>clock,reset=>reset,s=>p(246)(112),cout=>p(247)(113));
FA_ff_7520:FAff port map(x=>p(176)(113),y=>p(177)(113),Cin=>p(178)(113),clock=>clock,reset=>reset,s=>p(246)(113),cout=>p(247)(114));
FA_ff_7521:FAff port map(x=>p(176)(114),y=>p(177)(114),Cin=>p(178)(114),clock=>clock,reset=>reset,s=>p(246)(114),cout=>p(247)(115));
FA_ff_7522:FAff port map(x=>p(176)(115),y=>p(177)(115),Cin=>p(178)(115),clock=>clock,reset=>reset,s=>p(246)(115),cout=>p(247)(116));
FA_ff_7523:FAff port map(x=>p(176)(116),y=>p(177)(116),Cin=>p(178)(116),clock=>clock,reset=>reset,s=>p(246)(116),cout=>p(247)(117));
FA_ff_7524:FAff port map(x=>p(176)(117),y=>p(177)(117),Cin=>p(178)(117),clock=>clock,reset=>reset,s=>p(246)(117),cout=>p(247)(118));
FA_ff_7525:FAff port map(x=>p(176)(118),y=>p(177)(118),Cin=>p(178)(118),clock=>clock,reset=>reset,s=>p(246)(118),cout=>p(247)(119));
FA_ff_7526:FAff port map(x=>p(176)(119),y=>p(177)(119),Cin=>p(178)(119),clock=>clock,reset=>reset,s=>p(246)(119),cout=>p(247)(120));
FA_ff_7527:FAff port map(x=>p(176)(120),y=>p(177)(120),Cin=>p(178)(120),clock=>clock,reset=>reset,s=>p(246)(120),cout=>p(247)(121));
FA_ff_7528:FAff port map(x=>p(176)(121),y=>p(177)(121),Cin=>p(178)(121),clock=>clock,reset=>reset,s=>p(246)(121),cout=>p(247)(122));
FA_ff_7529:FAff port map(x=>p(176)(122),y=>p(177)(122),Cin=>p(178)(122),clock=>clock,reset=>reset,s=>p(246)(122),cout=>p(247)(123));
FA_ff_7530:FAff port map(x=>p(176)(123),y=>p(177)(123),Cin=>p(178)(123),clock=>clock,reset=>reset,s=>p(246)(123),cout=>p(247)(124));
FA_ff_7531:FAff port map(x=>p(176)(124),y=>p(177)(124),Cin=>p(178)(124),clock=>clock,reset=>reset,s=>p(246)(124),cout=>p(247)(125));
FA_ff_7532:FAff port map(x=>p(176)(125),y=>p(177)(125),Cin=>p(178)(125),clock=>clock,reset=>reset,s=>p(246)(125),cout=>p(247)(126));
FA_ff_7533:FAff port map(x=>p(176)(126),y=>p(177)(126),Cin=>p(178)(126),clock=>clock,reset=>reset,s=>p(246)(126),cout=>p(247)(127));
FA_ff_7534:FAff port map(x=>p(176)(127),y=>p(177)(127),Cin=>p(178)(127),clock=>clock,reset=>reset,s=>p(246)(127),cout=>p(247)(128));
p(246)(128)<=p(177)(128);
p(248)(0)<=p(180)(0);
FA_ff_7535:FAff port map(x=>p(179)(1),y=>p(180)(1),Cin=>p(181)(1),clock=>clock,reset=>reset,s=>p(248)(1),cout=>p(249)(2));
FA_ff_7536:FAff port map(x=>p(179)(2),y=>p(180)(2),Cin=>p(181)(2),clock=>clock,reset=>reset,s=>p(248)(2),cout=>p(249)(3));
FA_ff_7537:FAff port map(x=>p(179)(3),y=>p(180)(3),Cin=>p(181)(3),clock=>clock,reset=>reset,s=>p(248)(3),cout=>p(249)(4));
FA_ff_7538:FAff port map(x=>p(179)(4),y=>p(180)(4),Cin=>p(181)(4),clock=>clock,reset=>reset,s=>p(248)(4),cout=>p(249)(5));
FA_ff_7539:FAff port map(x=>p(179)(5),y=>p(180)(5),Cin=>p(181)(5),clock=>clock,reset=>reset,s=>p(248)(5),cout=>p(249)(6));
FA_ff_7540:FAff port map(x=>p(179)(6),y=>p(180)(6),Cin=>p(181)(6),clock=>clock,reset=>reset,s=>p(248)(6),cout=>p(249)(7));
FA_ff_7541:FAff port map(x=>p(179)(7),y=>p(180)(7),Cin=>p(181)(7),clock=>clock,reset=>reset,s=>p(248)(7),cout=>p(249)(8));
FA_ff_7542:FAff port map(x=>p(179)(8),y=>p(180)(8),Cin=>p(181)(8),clock=>clock,reset=>reset,s=>p(248)(8),cout=>p(249)(9));
FA_ff_7543:FAff port map(x=>p(179)(9),y=>p(180)(9),Cin=>p(181)(9),clock=>clock,reset=>reset,s=>p(248)(9),cout=>p(249)(10));
FA_ff_7544:FAff port map(x=>p(179)(10),y=>p(180)(10),Cin=>p(181)(10),clock=>clock,reset=>reset,s=>p(248)(10),cout=>p(249)(11));
FA_ff_7545:FAff port map(x=>p(179)(11),y=>p(180)(11),Cin=>p(181)(11),clock=>clock,reset=>reset,s=>p(248)(11),cout=>p(249)(12));
FA_ff_7546:FAff port map(x=>p(179)(12),y=>p(180)(12),Cin=>p(181)(12),clock=>clock,reset=>reset,s=>p(248)(12),cout=>p(249)(13));
FA_ff_7547:FAff port map(x=>p(179)(13),y=>p(180)(13),Cin=>p(181)(13),clock=>clock,reset=>reset,s=>p(248)(13),cout=>p(249)(14));
FA_ff_7548:FAff port map(x=>p(179)(14),y=>p(180)(14),Cin=>p(181)(14),clock=>clock,reset=>reset,s=>p(248)(14),cout=>p(249)(15));
FA_ff_7549:FAff port map(x=>p(179)(15),y=>p(180)(15),Cin=>p(181)(15),clock=>clock,reset=>reset,s=>p(248)(15),cout=>p(249)(16));
FA_ff_7550:FAff port map(x=>p(179)(16),y=>p(180)(16),Cin=>p(181)(16),clock=>clock,reset=>reset,s=>p(248)(16),cout=>p(249)(17));
FA_ff_7551:FAff port map(x=>p(179)(17),y=>p(180)(17),Cin=>p(181)(17),clock=>clock,reset=>reset,s=>p(248)(17),cout=>p(249)(18));
FA_ff_7552:FAff port map(x=>p(179)(18),y=>p(180)(18),Cin=>p(181)(18),clock=>clock,reset=>reset,s=>p(248)(18),cout=>p(249)(19));
FA_ff_7553:FAff port map(x=>p(179)(19),y=>p(180)(19),Cin=>p(181)(19),clock=>clock,reset=>reset,s=>p(248)(19),cout=>p(249)(20));
FA_ff_7554:FAff port map(x=>p(179)(20),y=>p(180)(20),Cin=>p(181)(20),clock=>clock,reset=>reset,s=>p(248)(20),cout=>p(249)(21));
FA_ff_7555:FAff port map(x=>p(179)(21),y=>p(180)(21),Cin=>p(181)(21),clock=>clock,reset=>reset,s=>p(248)(21),cout=>p(249)(22));
FA_ff_7556:FAff port map(x=>p(179)(22),y=>p(180)(22),Cin=>p(181)(22),clock=>clock,reset=>reset,s=>p(248)(22),cout=>p(249)(23));
FA_ff_7557:FAff port map(x=>p(179)(23),y=>p(180)(23),Cin=>p(181)(23),clock=>clock,reset=>reset,s=>p(248)(23),cout=>p(249)(24));
FA_ff_7558:FAff port map(x=>p(179)(24),y=>p(180)(24),Cin=>p(181)(24),clock=>clock,reset=>reset,s=>p(248)(24),cout=>p(249)(25));
FA_ff_7559:FAff port map(x=>p(179)(25),y=>p(180)(25),Cin=>p(181)(25),clock=>clock,reset=>reset,s=>p(248)(25),cout=>p(249)(26));
FA_ff_7560:FAff port map(x=>p(179)(26),y=>p(180)(26),Cin=>p(181)(26),clock=>clock,reset=>reset,s=>p(248)(26),cout=>p(249)(27));
FA_ff_7561:FAff port map(x=>p(179)(27),y=>p(180)(27),Cin=>p(181)(27),clock=>clock,reset=>reset,s=>p(248)(27),cout=>p(249)(28));
FA_ff_7562:FAff port map(x=>p(179)(28),y=>p(180)(28),Cin=>p(181)(28),clock=>clock,reset=>reset,s=>p(248)(28),cout=>p(249)(29));
FA_ff_7563:FAff port map(x=>p(179)(29),y=>p(180)(29),Cin=>p(181)(29),clock=>clock,reset=>reset,s=>p(248)(29),cout=>p(249)(30));
FA_ff_7564:FAff port map(x=>p(179)(30),y=>p(180)(30),Cin=>p(181)(30),clock=>clock,reset=>reset,s=>p(248)(30),cout=>p(249)(31));
FA_ff_7565:FAff port map(x=>p(179)(31),y=>p(180)(31),Cin=>p(181)(31),clock=>clock,reset=>reset,s=>p(248)(31),cout=>p(249)(32));
FA_ff_7566:FAff port map(x=>p(179)(32),y=>p(180)(32),Cin=>p(181)(32),clock=>clock,reset=>reset,s=>p(248)(32),cout=>p(249)(33));
FA_ff_7567:FAff port map(x=>p(179)(33),y=>p(180)(33),Cin=>p(181)(33),clock=>clock,reset=>reset,s=>p(248)(33),cout=>p(249)(34));
FA_ff_7568:FAff port map(x=>p(179)(34),y=>p(180)(34),Cin=>p(181)(34),clock=>clock,reset=>reset,s=>p(248)(34),cout=>p(249)(35));
FA_ff_7569:FAff port map(x=>p(179)(35),y=>p(180)(35),Cin=>p(181)(35),clock=>clock,reset=>reset,s=>p(248)(35),cout=>p(249)(36));
FA_ff_7570:FAff port map(x=>p(179)(36),y=>p(180)(36),Cin=>p(181)(36),clock=>clock,reset=>reset,s=>p(248)(36),cout=>p(249)(37));
FA_ff_7571:FAff port map(x=>p(179)(37),y=>p(180)(37),Cin=>p(181)(37),clock=>clock,reset=>reset,s=>p(248)(37),cout=>p(249)(38));
FA_ff_7572:FAff port map(x=>p(179)(38),y=>p(180)(38),Cin=>p(181)(38),clock=>clock,reset=>reset,s=>p(248)(38),cout=>p(249)(39));
FA_ff_7573:FAff port map(x=>p(179)(39),y=>p(180)(39),Cin=>p(181)(39),clock=>clock,reset=>reset,s=>p(248)(39),cout=>p(249)(40));
FA_ff_7574:FAff port map(x=>p(179)(40),y=>p(180)(40),Cin=>p(181)(40),clock=>clock,reset=>reset,s=>p(248)(40),cout=>p(249)(41));
FA_ff_7575:FAff port map(x=>p(179)(41),y=>p(180)(41),Cin=>p(181)(41),clock=>clock,reset=>reset,s=>p(248)(41),cout=>p(249)(42));
FA_ff_7576:FAff port map(x=>p(179)(42),y=>p(180)(42),Cin=>p(181)(42),clock=>clock,reset=>reset,s=>p(248)(42),cout=>p(249)(43));
FA_ff_7577:FAff port map(x=>p(179)(43),y=>p(180)(43),Cin=>p(181)(43),clock=>clock,reset=>reset,s=>p(248)(43),cout=>p(249)(44));
FA_ff_7578:FAff port map(x=>p(179)(44),y=>p(180)(44),Cin=>p(181)(44),clock=>clock,reset=>reset,s=>p(248)(44),cout=>p(249)(45));
FA_ff_7579:FAff port map(x=>p(179)(45),y=>p(180)(45),Cin=>p(181)(45),clock=>clock,reset=>reset,s=>p(248)(45),cout=>p(249)(46));
FA_ff_7580:FAff port map(x=>p(179)(46),y=>p(180)(46),Cin=>p(181)(46),clock=>clock,reset=>reset,s=>p(248)(46),cout=>p(249)(47));
FA_ff_7581:FAff port map(x=>p(179)(47),y=>p(180)(47),Cin=>p(181)(47),clock=>clock,reset=>reset,s=>p(248)(47),cout=>p(249)(48));
FA_ff_7582:FAff port map(x=>p(179)(48),y=>p(180)(48),Cin=>p(181)(48),clock=>clock,reset=>reset,s=>p(248)(48),cout=>p(249)(49));
FA_ff_7583:FAff port map(x=>p(179)(49),y=>p(180)(49),Cin=>p(181)(49),clock=>clock,reset=>reset,s=>p(248)(49),cout=>p(249)(50));
FA_ff_7584:FAff port map(x=>p(179)(50),y=>p(180)(50),Cin=>p(181)(50),clock=>clock,reset=>reset,s=>p(248)(50),cout=>p(249)(51));
FA_ff_7585:FAff port map(x=>p(179)(51),y=>p(180)(51),Cin=>p(181)(51),clock=>clock,reset=>reset,s=>p(248)(51),cout=>p(249)(52));
FA_ff_7586:FAff port map(x=>p(179)(52),y=>p(180)(52),Cin=>p(181)(52),clock=>clock,reset=>reset,s=>p(248)(52),cout=>p(249)(53));
FA_ff_7587:FAff port map(x=>p(179)(53),y=>p(180)(53),Cin=>p(181)(53),clock=>clock,reset=>reset,s=>p(248)(53),cout=>p(249)(54));
FA_ff_7588:FAff port map(x=>p(179)(54),y=>p(180)(54),Cin=>p(181)(54),clock=>clock,reset=>reset,s=>p(248)(54),cout=>p(249)(55));
FA_ff_7589:FAff port map(x=>p(179)(55),y=>p(180)(55),Cin=>p(181)(55),clock=>clock,reset=>reset,s=>p(248)(55),cout=>p(249)(56));
FA_ff_7590:FAff port map(x=>p(179)(56),y=>p(180)(56),Cin=>p(181)(56),clock=>clock,reset=>reset,s=>p(248)(56),cout=>p(249)(57));
FA_ff_7591:FAff port map(x=>p(179)(57),y=>p(180)(57),Cin=>p(181)(57),clock=>clock,reset=>reset,s=>p(248)(57),cout=>p(249)(58));
FA_ff_7592:FAff port map(x=>p(179)(58),y=>p(180)(58),Cin=>p(181)(58),clock=>clock,reset=>reset,s=>p(248)(58),cout=>p(249)(59));
FA_ff_7593:FAff port map(x=>p(179)(59),y=>p(180)(59),Cin=>p(181)(59),clock=>clock,reset=>reset,s=>p(248)(59),cout=>p(249)(60));
FA_ff_7594:FAff port map(x=>p(179)(60),y=>p(180)(60),Cin=>p(181)(60),clock=>clock,reset=>reset,s=>p(248)(60),cout=>p(249)(61));
FA_ff_7595:FAff port map(x=>p(179)(61),y=>p(180)(61),Cin=>p(181)(61),clock=>clock,reset=>reset,s=>p(248)(61),cout=>p(249)(62));
FA_ff_7596:FAff port map(x=>p(179)(62),y=>p(180)(62),Cin=>p(181)(62),clock=>clock,reset=>reset,s=>p(248)(62),cout=>p(249)(63));
FA_ff_7597:FAff port map(x=>p(179)(63),y=>p(180)(63),Cin=>p(181)(63),clock=>clock,reset=>reset,s=>p(248)(63),cout=>p(249)(64));
FA_ff_7598:FAff port map(x=>p(179)(64),y=>p(180)(64),Cin=>p(181)(64),clock=>clock,reset=>reset,s=>p(248)(64),cout=>p(249)(65));
FA_ff_7599:FAff port map(x=>p(179)(65),y=>p(180)(65),Cin=>p(181)(65),clock=>clock,reset=>reset,s=>p(248)(65),cout=>p(249)(66));
FA_ff_7600:FAff port map(x=>p(179)(66),y=>p(180)(66),Cin=>p(181)(66),clock=>clock,reset=>reset,s=>p(248)(66),cout=>p(249)(67));
FA_ff_7601:FAff port map(x=>p(179)(67),y=>p(180)(67),Cin=>p(181)(67),clock=>clock,reset=>reset,s=>p(248)(67),cout=>p(249)(68));
FA_ff_7602:FAff port map(x=>p(179)(68),y=>p(180)(68),Cin=>p(181)(68),clock=>clock,reset=>reset,s=>p(248)(68),cout=>p(249)(69));
FA_ff_7603:FAff port map(x=>p(179)(69),y=>p(180)(69),Cin=>p(181)(69),clock=>clock,reset=>reset,s=>p(248)(69),cout=>p(249)(70));
FA_ff_7604:FAff port map(x=>p(179)(70),y=>p(180)(70),Cin=>p(181)(70),clock=>clock,reset=>reset,s=>p(248)(70),cout=>p(249)(71));
FA_ff_7605:FAff port map(x=>p(179)(71),y=>p(180)(71),Cin=>p(181)(71),clock=>clock,reset=>reset,s=>p(248)(71),cout=>p(249)(72));
FA_ff_7606:FAff port map(x=>p(179)(72),y=>p(180)(72),Cin=>p(181)(72),clock=>clock,reset=>reset,s=>p(248)(72),cout=>p(249)(73));
FA_ff_7607:FAff port map(x=>p(179)(73),y=>p(180)(73),Cin=>p(181)(73),clock=>clock,reset=>reset,s=>p(248)(73),cout=>p(249)(74));
FA_ff_7608:FAff port map(x=>p(179)(74),y=>p(180)(74),Cin=>p(181)(74),clock=>clock,reset=>reset,s=>p(248)(74),cout=>p(249)(75));
FA_ff_7609:FAff port map(x=>p(179)(75),y=>p(180)(75),Cin=>p(181)(75),clock=>clock,reset=>reset,s=>p(248)(75),cout=>p(249)(76));
FA_ff_7610:FAff port map(x=>p(179)(76),y=>p(180)(76),Cin=>p(181)(76),clock=>clock,reset=>reset,s=>p(248)(76),cout=>p(249)(77));
FA_ff_7611:FAff port map(x=>p(179)(77),y=>p(180)(77),Cin=>p(181)(77),clock=>clock,reset=>reset,s=>p(248)(77),cout=>p(249)(78));
FA_ff_7612:FAff port map(x=>p(179)(78),y=>p(180)(78),Cin=>p(181)(78),clock=>clock,reset=>reset,s=>p(248)(78),cout=>p(249)(79));
FA_ff_7613:FAff port map(x=>p(179)(79),y=>p(180)(79),Cin=>p(181)(79),clock=>clock,reset=>reset,s=>p(248)(79),cout=>p(249)(80));
FA_ff_7614:FAff port map(x=>p(179)(80),y=>p(180)(80),Cin=>p(181)(80),clock=>clock,reset=>reset,s=>p(248)(80),cout=>p(249)(81));
FA_ff_7615:FAff port map(x=>p(179)(81),y=>p(180)(81),Cin=>p(181)(81),clock=>clock,reset=>reset,s=>p(248)(81),cout=>p(249)(82));
FA_ff_7616:FAff port map(x=>p(179)(82),y=>p(180)(82),Cin=>p(181)(82),clock=>clock,reset=>reset,s=>p(248)(82),cout=>p(249)(83));
FA_ff_7617:FAff port map(x=>p(179)(83),y=>p(180)(83),Cin=>p(181)(83),clock=>clock,reset=>reset,s=>p(248)(83),cout=>p(249)(84));
FA_ff_7618:FAff port map(x=>p(179)(84),y=>p(180)(84),Cin=>p(181)(84),clock=>clock,reset=>reset,s=>p(248)(84),cout=>p(249)(85));
FA_ff_7619:FAff port map(x=>p(179)(85),y=>p(180)(85),Cin=>p(181)(85),clock=>clock,reset=>reset,s=>p(248)(85),cout=>p(249)(86));
FA_ff_7620:FAff port map(x=>p(179)(86),y=>p(180)(86),Cin=>p(181)(86),clock=>clock,reset=>reset,s=>p(248)(86),cout=>p(249)(87));
FA_ff_7621:FAff port map(x=>p(179)(87),y=>p(180)(87),Cin=>p(181)(87),clock=>clock,reset=>reset,s=>p(248)(87),cout=>p(249)(88));
FA_ff_7622:FAff port map(x=>p(179)(88),y=>p(180)(88),Cin=>p(181)(88),clock=>clock,reset=>reset,s=>p(248)(88),cout=>p(249)(89));
FA_ff_7623:FAff port map(x=>p(179)(89),y=>p(180)(89),Cin=>p(181)(89),clock=>clock,reset=>reset,s=>p(248)(89),cout=>p(249)(90));
FA_ff_7624:FAff port map(x=>p(179)(90),y=>p(180)(90),Cin=>p(181)(90),clock=>clock,reset=>reset,s=>p(248)(90),cout=>p(249)(91));
FA_ff_7625:FAff port map(x=>p(179)(91),y=>p(180)(91),Cin=>p(181)(91),clock=>clock,reset=>reset,s=>p(248)(91),cout=>p(249)(92));
FA_ff_7626:FAff port map(x=>p(179)(92),y=>p(180)(92),Cin=>p(181)(92),clock=>clock,reset=>reset,s=>p(248)(92),cout=>p(249)(93));
FA_ff_7627:FAff port map(x=>p(179)(93),y=>p(180)(93),Cin=>p(181)(93),clock=>clock,reset=>reset,s=>p(248)(93),cout=>p(249)(94));
FA_ff_7628:FAff port map(x=>p(179)(94),y=>p(180)(94),Cin=>p(181)(94),clock=>clock,reset=>reset,s=>p(248)(94),cout=>p(249)(95));
FA_ff_7629:FAff port map(x=>p(179)(95),y=>p(180)(95),Cin=>p(181)(95),clock=>clock,reset=>reset,s=>p(248)(95),cout=>p(249)(96));
FA_ff_7630:FAff port map(x=>p(179)(96),y=>p(180)(96),Cin=>p(181)(96),clock=>clock,reset=>reset,s=>p(248)(96),cout=>p(249)(97));
FA_ff_7631:FAff port map(x=>p(179)(97),y=>p(180)(97),Cin=>p(181)(97),clock=>clock,reset=>reset,s=>p(248)(97),cout=>p(249)(98));
FA_ff_7632:FAff port map(x=>p(179)(98),y=>p(180)(98),Cin=>p(181)(98),clock=>clock,reset=>reset,s=>p(248)(98),cout=>p(249)(99));
FA_ff_7633:FAff port map(x=>p(179)(99),y=>p(180)(99),Cin=>p(181)(99),clock=>clock,reset=>reset,s=>p(248)(99),cout=>p(249)(100));
FA_ff_7634:FAff port map(x=>p(179)(100),y=>p(180)(100),Cin=>p(181)(100),clock=>clock,reset=>reset,s=>p(248)(100),cout=>p(249)(101));
FA_ff_7635:FAff port map(x=>p(179)(101),y=>p(180)(101),Cin=>p(181)(101),clock=>clock,reset=>reset,s=>p(248)(101),cout=>p(249)(102));
FA_ff_7636:FAff port map(x=>p(179)(102),y=>p(180)(102),Cin=>p(181)(102),clock=>clock,reset=>reset,s=>p(248)(102),cout=>p(249)(103));
FA_ff_7637:FAff port map(x=>p(179)(103),y=>p(180)(103),Cin=>p(181)(103),clock=>clock,reset=>reset,s=>p(248)(103),cout=>p(249)(104));
FA_ff_7638:FAff port map(x=>p(179)(104),y=>p(180)(104),Cin=>p(181)(104),clock=>clock,reset=>reset,s=>p(248)(104),cout=>p(249)(105));
FA_ff_7639:FAff port map(x=>p(179)(105),y=>p(180)(105),Cin=>p(181)(105),clock=>clock,reset=>reset,s=>p(248)(105),cout=>p(249)(106));
FA_ff_7640:FAff port map(x=>p(179)(106),y=>p(180)(106),Cin=>p(181)(106),clock=>clock,reset=>reset,s=>p(248)(106),cout=>p(249)(107));
FA_ff_7641:FAff port map(x=>p(179)(107),y=>p(180)(107),Cin=>p(181)(107),clock=>clock,reset=>reset,s=>p(248)(107),cout=>p(249)(108));
FA_ff_7642:FAff port map(x=>p(179)(108),y=>p(180)(108),Cin=>p(181)(108),clock=>clock,reset=>reset,s=>p(248)(108),cout=>p(249)(109));
FA_ff_7643:FAff port map(x=>p(179)(109),y=>p(180)(109),Cin=>p(181)(109),clock=>clock,reset=>reset,s=>p(248)(109),cout=>p(249)(110));
FA_ff_7644:FAff port map(x=>p(179)(110),y=>p(180)(110),Cin=>p(181)(110),clock=>clock,reset=>reset,s=>p(248)(110),cout=>p(249)(111));
FA_ff_7645:FAff port map(x=>p(179)(111),y=>p(180)(111),Cin=>p(181)(111),clock=>clock,reset=>reset,s=>p(248)(111),cout=>p(249)(112));
FA_ff_7646:FAff port map(x=>p(179)(112),y=>p(180)(112),Cin=>p(181)(112),clock=>clock,reset=>reset,s=>p(248)(112),cout=>p(249)(113));
FA_ff_7647:FAff port map(x=>p(179)(113),y=>p(180)(113),Cin=>p(181)(113),clock=>clock,reset=>reset,s=>p(248)(113),cout=>p(249)(114));
FA_ff_7648:FAff port map(x=>p(179)(114),y=>p(180)(114),Cin=>p(181)(114),clock=>clock,reset=>reset,s=>p(248)(114),cout=>p(249)(115));
FA_ff_7649:FAff port map(x=>p(179)(115),y=>p(180)(115),Cin=>p(181)(115),clock=>clock,reset=>reset,s=>p(248)(115),cout=>p(249)(116));
FA_ff_7650:FAff port map(x=>p(179)(116),y=>p(180)(116),Cin=>p(181)(116),clock=>clock,reset=>reset,s=>p(248)(116),cout=>p(249)(117));
FA_ff_7651:FAff port map(x=>p(179)(117),y=>p(180)(117),Cin=>p(181)(117),clock=>clock,reset=>reset,s=>p(248)(117),cout=>p(249)(118));
FA_ff_7652:FAff port map(x=>p(179)(118),y=>p(180)(118),Cin=>p(181)(118),clock=>clock,reset=>reset,s=>p(248)(118),cout=>p(249)(119));
FA_ff_7653:FAff port map(x=>p(179)(119),y=>p(180)(119),Cin=>p(181)(119),clock=>clock,reset=>reset,s=>p(248)(119),cout=>p(249)(120));
FA_ff_7654:FAff port map(x=>p(179)(120),y=>p(180)(120),Cin=>p(181)(120),clock=>clock,reset=>reset,s=>p(248)(120),cout=>p(249)(121));
FA_ff_7655:FAff port map(x=>p(179)(121),y=>p(180)(121),Cin=>p(181)(121),clock=>clock,reset=>reset,s=>p(248)(121),cout=>p(249)(122));
FA_ff_7656:FAff port map(x=>p(179)(122),y=>p(180)(122),Cin=>p(181)(122),clock=>clock,reset=>reset,s=>p(248)(122),cout=>p(249)(123));
FA_ff_7657:FAff port map(x=>p(179)(123),y=>p(180)(123),Cin=>p(181)(123),clock=>clock,reset=>reset,s=>p(248)(123),cout=>p(249)(124));
FA_ff_7658:FAff port map(x=>p(179)(124),y=>p(180)(124),Cin=>p(181)(124),clock=>clock,reset=>reset,s=>p(248)(124),cout=>p(249)(125));
FA_ff_7659:FAff port map(x=>p(179)(125),y=>p(180)(125),Cin=>p(181)(125),clock=>clock,reset=>reset,s=>p(248)(125),cout=>p(249)(126));
FA_ff_7660:FAff port map(x=>p(179)(126),y=>p(180)(126),Cin=>p(181)(126),clock=>clock,reset=>reset,s=>p(248)(126),cout=>p(249)(127));
FA_ff_7661:FAff port map(x=>p(179)(127),y=>p(180)(127),Cin=>p(181)(127),clock=>clock,reset=>reset,s=>p(248)(127),cout=>p(249)(128));
HA_ff_17:HAff port map(x=>p(179)(128),y=>p(181)(128),clock=>clock,reset=>reset,s=>p(248)(128),c=>p(249)(129));
HA_ff_18:HAff port map(x=>p(182)(0),y=>p(184)(0),clock=>clock,reset=>reset,s=>p(250)(0),c=>p(251)(1));
FA_ff_7662:FAff port map(x=>p(182)(1),y=>p(183)(1),Cin=>p(184)(1),clock=>clock,reset=>reset,s=>p(250)(1),cout=>p(251)(2));
FA_ff_7663:FAff port map(x=>p(182)(2),y=>p(183)(2),Cin=>p(184)(2),clock=>clock,reset=>reset,s=>p(250)(2),cout=>p(251)(3));
FA_ff_7664:FAff port map(x=>p(182)(3),y=>p(183)(3),Cin=>p(184)(3),clock=>clock,reset=>reset,s=>p(250)(3),cout=>p(251)(4));
FA_ff_7665:FAff port map(x=>p(182)(4),y=>p(183)(4),Cin=>p(184)(4),clock=>clock,reset=>reset,s=>p(250)(4),cout=>p(251)(5));
FA_ff_7666:FAff port map(x=>p(182)(5),y=>p(183)(5),Cin=>p(184)(5),clock=>clock,reset=>reset,s=>p(250)(5),cout=>p(251)(6));
FA_ff_7667:FAff port map(x=>p(182)(6),y=>p(183)(6),Cin=>p(184)(6),clock=>clock,reset=>reset,s=>p(250)(6),cout=>p(251)(7));
FA_ff_7668:FAff port map(x=>p(182)(7),y=>p(183)(7),Cin=>p(184)(7),clock=>clock,reset=>reset,s=>p(250)(7),cout=>p(251)(8));
FA_ff_7669:FAff port map(x=>p(182)(8),y=>p(183)(8),Cin=>p(184)(8),clock=>clock,reset=>reset,s=>p(250)(8),cout=>p(251)(9));
FA_ff_7670:FAff port map(x=>p(182)(9),y=>p(183)(9),Cin=>p(184)(9),clock=>clock,reset=>reset,s=>p(250)(9),cout=>p(251)(10));
FA_ff_7671:FAff port map(x=>p(182)(10),y=>p(183)(10),Cin=>p(184)(10),clock=>clock,reset=>reset,s=>p(250)(10),cout=>p(251)(11));
FA_ff_7672:FAff port map(x=>p(182)(11),y=>p(183)(11),Cin=>p(184)(11),clock=>clock,reset=>reset,s=>p(250)(11),cout=>p(251)(12));
FA_ff_7673:FAff port map(x=>p(182)(12),y=>p(183)(12),Cin=>p(184)(12),clock=>clock,reset=>reset,s=>p(250)(12),cout=>p(251)(13));
FA_ff_7674:FAff port map(x=>p(182)(13),y=>p(183)(13),Cin=>p(184)(13),clock=>clock,reset=>reset,s=>p(250)(13),cout=>p(251)(14));
FA_ff_7675:FAff port map(x=>p(182)(14),y=>p(183)(14),Cin=>p(184)(14),clock=>clock,reset=>reset,s=>p(250)(14),cout=>p(251)(15));
FA_ff_7676:FAff port map(x=>p(182)(15),y=>p(183)(15),Cin=>p(184)(15),clock=>clock,reset=>reset,s=>p(250)(15),cout=>p(251)(16));
FA_ff_7677:FAff port map(x=>p(182)(16),y=>p(183)(16),Cin=>p(184)(16),clock=>clock,reset=>reset,s=>p(250)(16),cout=>p(251)(17));
FA_ff_7678:FAff port map(x=>p(182)(17),y=>p(183)(17),Cin=>p(184)(17),clock=>clock,reset=>reset,s=>p(250)(17),cout=>p(251)(18));
FA_ff_7679:FAff port map(x=>p(182)(18),y=>p(183)(18),Cin=>p(184)(18),clock=>clock,reset=>reset,s=>p(250)(18),cout=>p(251)(19));
FA_ff_7680:FAff port map(x=>p(182)(19),y=>p(183)(19),Cin=>p(184)(19),clock=>clock,reset=>reset,s=>p(250)(19),cout=>p(251)(20));
FA_ff_7681:FAff port map(x=>p(182)(20),y=>p(183)(20),Cin=>p(184)(20),clock=>clock,reset=>reset,s=>p(250)(20),cout=>p(251)(21));
FA_ff_7682:FAff port map(x=>p(182)(21),y=>p(183)(21),Cin=>p(184)(21),clock=>clock,reset=>reset,s=>p(250)(21),cout=>p(251)(22));
FA_ff_7683:FAff port map(x=>p(182)(22),y=>p(183)(22),Cin=>p(184)(22),clock=>clock,reset=>reset,s=>p(250)(22),cout=>p(251)(23));
FA_ff_7684:FAff port map(x=>p(182)(23),y=>p(183)(23),Cin=>p(184)(23),clock=>clock,reset=>reset,s=>p(250)(23),cout=>p(251)(24));
FA_ff_7685:FAff port map(x=>p(182)(24),y=>p(183)(24),Cin=>p(184)(24),clock=>clock,reset=>reset,s=>p(250)(24),cout=>p(251)(25));
FA_ff_7686:FAff port map(x=>p(182)(25),y=>p(183)(25),Cin=>p(184)(25),clock=>clock,reset=>reset,s=>p(250)(25),cout=>p(251)(26));
FA_ff_7687:FAff port map(x=>p(182)(26),y=>p(183)(26),Cin=>p(184)(26),clock=>clock,reset=>reset,s=>p(250)(26),cout=>p(251)(27));
FA_ff_7688:FAff port map(x=>p(182)(27),y=>p(183)(27),Cin=>p(184)(27),clock=>clock,reset=>reset,s=>p(250)(27),cout=>p(251)(28));
FA_ff_7689:FAff port map(x=>p(182)(28),y=>p(183)(28),Cin=>p(184)(28),clock=>clock,reset=>reset,s=>p(250)(28),cout=>p(251)(29));
FA_ff_7690:FAff port map(x=>p(182)(29),y=>p(183)(29),Cin=>p(184)(29),clock=>clock,reset=>reset,s=>p(250)(29),cout=>p(251)(30));
FA_ff_7691:FAff port map(x=>p(182)(30),y=>p(183)(30),Cin=>p(184)(30),clock=>clock,reset=>reset,s=>p(250)(30),cout=>p(251)(31));
FA_ff_7692:FAff port map(x=>p(182)(31),y=>p(183)(31),Cin=>p(184)(31),clock=>clock,reset=>reset,s=>p(250)(31),cout=>p(251)(32));
FA_ff_7693:FAff port map(x=>p(182)(32),y=>p(183)(32),Cin=>p(184)(32),clock=>clock,reset=>reset,s=>p(250)(32),cout=>p(251)(33));
FA_ff_7694:FAff port map(x=>p(182)(33),y=>p(183)(33),Cin=>p(184)(33),clock=>clock,reset=>reset,s=>p(250)(33),cout=>p(251)(34));
FA_ff_7695:FAff port map(x=>p(182)(34),y=>p(183)(34),Cin=>p(184)(34),clock=>clock,reset=>reset,s=>p(250)(34),cout=>p(251)(35));
FA_ff_7696:FAff port map(x=>p(182)(35),y=>p(183)(35),Cin=>p(184)(35),clock=>clock,reset=>reset,s=>p(250)(35),cout=>p(251)(36));
FA_ff_7697:FAff port map(x=>p(182)(36),y=>p(183)(36),Cin=>p(184)(36),clock=>clock,reset=>reset,s=>p(250)(36),cout=>p(251)(37));
FA_ff_7698:FAff port map(x=>p(182)(37),y=>p(183)(37),Cin=>p(184)(37),clock=>clock,reset=>reset,s=>p(250)(37),cout=>p(251)(38));
FA_ff_7699:FAff port map(x=>p(182)(38),y=>p(183)(38),Cin=>p(184)(38),clock=>clock,reset=>reset,s=>p(250)(38),cout=>p(251)(39));
FA_ff_7700:FAff port map(x=>p(182)(39),y=>p(183)(39),Cin=>p(184)(39),clock=>clock,reset=>reset,s=>p(250)(39),cout=>p(251)(40));
FA_ff_7701:FAff port map(x=>p(182)(40),y=>p(183)(40),Cin=>p(184)(40),clock=>clock,reset=>reset,s=>p(250)(40),cout=>p(251)(41));
FA_ff_7702:FAff port map(x=>p(182)(41),y=>p(183)(41),Cin=>p(184)(41),clock=>clock,reset=>reset,s=>p(250)(41),cout=>p(251)(42));
FA_ff_7703:FAff port map(x=>p(182)(42),y=>p(183)(42),Cin=>p(184)(42),clock=>clock,reset=>reset,s=>p(250)(42),cout=>p(251)(43));
FA_ff_7704:FAff port map(x=>p(182)(43),y=>p(183)(43),Cin=>p(184)(43),clock=>clock,reset=>reset,s=>p(250)(43),cout=>p(251)(44));
FA_ff_7705:FAff port map(x=>p(182)(44),y=>p(183)(44),Cin=>p(184)(44),clock=>clock,reset=>reset,s=>p(250)(44),cout=>p(251)(45));
FA_ff_7706:FAff port map(x=>p(182)(45),y=>p(183)(45),Cin=>p(184)(45),clock=>clock,reset=>reset,s=>p(250)(45),cout=>p(251)(46));
FA_ff_7707:FAff port map(x=>p(182)(46),y=>p(183)(46),Cin=>p(184)(46),clock=>clock,reset=>reset,s=>p(250)(46),cout=>p(251)(47));
FA_ff_7708:FAff port map(x=>p(182)(47),y=>p(183)(47),Cin=>p(184)(47),clock=>clock,reset=>reset,s=>p(250)(47),cout=>p(251)(48));
FA_ff_7709:FAff port map(x=>p(182)(48),y=>p(183)(48),Cin=>p(184)(48),clock=>clock,reset=>reset,s=>p(250)(48),cout=>p(251)(49));
FA_ff_7710:FAff port map(x=>p(182)(49),y=>p(183)(49),Cin=>p(184)(49),clock=>clock,reset=>reset,s=>p(250)(49),cout=>p(251)(50));
FA_ff_7711:FAff port map(x=>p(182)(50),y=>p(183)(50),Cin=>p(184)(50),clock=>clock,reset=>reset,s=>p(250)(50),cout=>p(251)(51));
FA_ff_7712:FAff port map(x=>p(182)(51),y=>p(183)(51),Cin=>p(184)(51),clock=>clock,reset=>reset,s=>p(250)(51),cout=>p(251)(52));
FA_ff_7713:FAff port map(x=>p(182)(52),y=>p(183)(52),Cin=>p(184)(52),clock=>clock,reset=>reset,s=>p(250)(52),cout=>p(251)(53));
FA_ff_7714:FAff port map(x=>p(182)(53),y=>p(183)(53),Cin=>p(184)(53),clock=>clock,reset=>reset,s=>p(250)(53),cout=>p(251)(54));
FA_ff_7715:FAff port map(x=>p(182)(54),y=>p(183)(54),Cin=>p(184)(54),clock=>clock,reset=>reset,s=>p(250)(54),cout=>p(251)(55));
FA_ff_7716:FAff port map(x=>p(182)(55),y=>p(183)(55),Cin=>p(184)(55),clock=>clock,reset=>reset,s=>p(250)(55),cout=>p(251)(56));
FA_ff_7717:FAff port map(x=>p(182)(56),y=>p(183)(56),Cin=>p(184)(56),clock=>clock,reset=>reset,s=>p(250)(56),cout=>p(251)(57));
FA_ff_7718:FAff port map(x=>p(182)(57),y=>p(183)(57),Cin=>p(184)(57),clock=>clock,reset=>reset,s=>p(250)(57),cout=>p(251)(58));
FA_ff_7719:FAff port map(x=>p(182)(58),y=>p(183)(58),Cin=>p(184)(58),clock=>clock,reset=>reset,s=>p(250)(58),cout=>p(251)(59));
FA_ff_7720:FAff port map(x=>p(182)(59),y=>p(183)(59),Cin=>p(184)(59),clock=>clock,reset=>reset,s=>p(250)(59),cout=>p(251)(60));
FA_ff_7721:FAff port map(x=>p(182)(60),y=>p(183)(60),Cin=>p(184)(60),clock=>clock,reset=>reset,s=>p(250)(60),cout=>p(251)(61));
FA_ff_7722:FAff port map(x=>p(182)(61),y=>p(183)(61),Cin=>p(184)(61),clock=>clock,reset=>reset,s=>p(250)(61),cout=>p(251)(62));
FA_ff_7723:FAff port map(x=>p(182)(62),y=>p(183)(62),Cin=>p(184)(62),clock=>clock,reset=>reset,s=>p(250)(62),cout=>p(251)(63));
FA_ff_7724:FAff port map(x=>p(182)(63),y=>p(183)(63),Cin=>p(184)(63),clock=>clock,reset=>reset,s=>p(250)(63),cout=>p(251)(64));
FA_ff_7725:FAff port map(x=>p(182)(64),y=>p(183)(64),Cin=>p(184)(64),clock=>clock,reset=>reset,s=>p(250)(64),cout=>p(251)(65));
FA_ff_7726:FAff port map(x=>p(182)(65),y=>p(183)(65),Cin=>p(184)(65),clock=>clock,reset=>reset,s=>p(250)(65),cout=>p(251)(66));
FA_ff_7727:FAff port map(x=>p(182)(66),y=>p(183)(66),Cin=>p(184)(66),clock=>clock,reset=>reset,s=>p(250)(66),cout=>p(251)(67));
FA_ff_7728:FAff port map(x=>p(182)(67),y=>p(183)(67),Cin=>p(184)(67),clock=>clock,reset=>reset,s=>p(250)(67),cout=>p(251)(68));
FA_ff_7729:FAff port map(x=>p(182)(68),y=>p(183)(68),Cin=>p(184)(68),clock=>clock,reset=>reset,s=>p(250)(68),cout=>p(251)(69));
FA_ff_7730:FAff port map(x=>p(182)(69),y=>p(183)(69),Cin=>p(184)(69),clock=>clock,reset=>reset,s=>p(250)(69),cout=>p(251)(70));
FA_ff_7731:FAff port map(x=>p(182)(70),y=>p(183)(70),Cin=>p(184)(70),clock=>clock,reset=>reset,s=>p(250)(70),cout=>p(251)(71));
FA_ff_7732:FAff port map(x=>p(182)(71),y=>p(183)(71),Cin=>p(184)(71),clock=>clock,reset=>reset,s=>p(250)(71),cout=>p(251)(72));
FA_ff_7733:FAff port map(x=>p(182)(72),y=>p(183)(72),Cin=>p(184)(72),clock=>clock,reset=>reset,s=>p(250)(72),cout=>p(251)(73));
FA_ff_7734:FAff port map(x=>p(182)(73),y=>p(183)(73),Cin=>p(184)(73),clock=>clock,reset=>reset,s=>p(250)(73),cout=>p(251)(74));
FA_ff_7735:FAff port map(x=>p(182)(74),y=>p(183)(74),Cin=>p(184)(74),clock=>clock,reset=>reset,s=>p(250)(74),cout=>p(251)(75));
FA_ff_7736:FAff port map(x=>p(182)(75),y=>p(183)(75),Cin=>p(184)(75),clock=>clock,reset=>reset,s=>p(250)(75),cout=>p(251)(76));
FA_ff_7737:FAff port map(x=>p(182)(76),y=>p(183)(76),Cin=>p(184)(76),clock=>clock,reset=>reset,s=>p(250)(76),cout=>p(251)(77));
FA_ff_7738:FAff port map(x=>p(182)(77),y=>p(183)(77),Cin=>p(184)(77),clock=>clock,reset=>reset,s=>p(250)(77),cout=>p(251)(78));
FA_ff_7739:FAff port map(x=>p(182)(78),y=>p(183)(78),Cin=>p(184)(78),clock=>clock,reset=>reset,s=>p(250)(78),cout=>p(251)(79));
FA_ff_7740:FAff port map(x=>p(182)(79),y=>p(183)(79),Cin=>p(184)(79),clock=>clock,reset=>reset,s=>p(250)(79),cout=>p(251)(80));
FA_ff_7741:FAff port map(x=>p(182)(80),y=>p(183)(80),Cin=>p(184)(80),clock=>clock,reset=>reset,s=>p(250)(80),cout=>p(251)(81));
FA_ff_7742:FAff port map(x=>p(182)(81),y=>p(183)(81),Cin=>p(184)(81),clock=>clock,reset=>reset,s=>p(250)(81),cout=>p(251)(82));
FA_ff_7743:FAff port map(x=>p(182)(82),y=>p(183)(82),Cin=>p(184)(82),clock=>clock,reset=>reset,s=>p(250)(82),cout=>p(251)(83));
FA_ff_7744:FAff port map(x=>p(182)(83),y=>p(183)(83),Cin=>p(184)(83),clock=>clock,reset=>reset,s=>p(250)(83),cout=>p(251)(84));
FA_ff_7745:FAff port map(x=>p(182)(84),y=>p(183)(84),Cin=>p(184)(84),clock=>clock,reset=>reset,s=>p(250)(84),cout=>p(251)(85));
FA_ff_7746:FAff port map(x=>p(182)(85),y=>p(183)(85),Cin=>p(184)(85),clock=>clock,reset=>reset,s=>p(250)(85),cout=>p(251)(86));
FA_ff_7747:FAff port map(x=>p(182)(86),y=>p(183)(86),Cin=>p(184)(86),clock=>clock,reset=>reset,s=>p(250)(86),cout=>p(251)(87));
FA_ff_7748:FAff port map(x=>p(182)(87),y=>p(183)(87),Cin=>p(184)(87),clock=>clock,reset=>reset,s=>p(250)(87),cout=>p(251)(88));
FA_ff_7749:FAff port map(x=>p(182)(88),y=>p(183)(88),Cin=>p(184)(88),clock=>clock,reset=>reset,s=>p(250)(88),cout=>p(251)(89));
FA_ff_7750:FAff port map(x=>p(182)(89),y=>p(183)(89),Cin=>p(184)(89),clock=>clock,reset=>reset,s=>p(250)(89),cout=>p(251)(90));
FA_ff_7751:FAff port map(x=>p(182)(90),y=>p(183)(90),Cin=>p(184)(90),clock=>clock,reset=>reset,s=>p(250)(90),cout=>p(251)(91));
FA_ff_7752:FAff port map(x=>p(182)(91),y=>p(183)(91),Cin=>p(184)(91),clock=>clock,reset=>reset,s=>p(250)(91),cout=>p(251)(92));
FA_ff_7753:FAff port map(x=>p(182)(92),y=>p(183)(92),Cin=>p(184)(92),clock=>clock,reset=>reset,s=>p(250)(92),cout=>p(251)(93));
FA_ff_7754:FAff port map(x=>p(182)(93),y=>p(183)(93),Cin=>p(184)(93),clock=>clock,reset=>reset,s=>p(250)(93),cout=>p(251)(94));
FA_ff_7755:FAff port map(x=>p(182)(94),y=>p(183)(94),Cin=>p(184)(94),clock=>clock,reset=>reset,s=>p(250)(94),cout=>p(251)(95));
FA_ff_7756:FAff port map(x=>p(182)(95),y=>p(183)(95),Cin=>p(184)(95),clock=>clock,reset=>reset,s=>p(250)(95),cout=>p(251)(96));
FA_ff_7757:FAff port map(x=>p(182)(96),y=>p(183)(96),Cin=>p(184)(96),clock=>clock,reset=>reset,s=>p(250)(96),cout=>p(251)(97));
FA_ff_7758:FAff port map(x=>p(182)(97),y=>p(183)(97),Cin=>p(184)(97),clock=>clock,reset=>reset,s=>p(250)(97),cout=>p(251)(98));
FA_ff_7759:FAff port map(x=>p(182)(98),y=>p(183)(98),Cin=>p(184)(98),clock=>clock,reset=>reset,s=>p(250)(98),cout=>p(251)(99));
FA_ff_7760:FAff port map(x=>p(182)(99),y=>p(183)(99),Cin=>p(184)(99),clock=>clock,reset=>reset,s=>p(250)(99),cout=>p(251)(100));
FA_ff_7761:FAff port map(x=>p(182)(100),y=>p(183)(100),Cin=>p(184)(100),clock=>clock,reset=>reset,s=>p(250)(100),cout=>p(251)(101));
FA_ff_7762:FAff port map(x=>p(182)(101),y=>p(183)(101),Cin=>p(184)(101),clock=>clock,reset=>reset,s=>p(250)(101),cout=>p(251)(102));
FA_ff_7763:FAff port map(x=>p(182)(102),y=>p(183)(102),Cin=>p(184)(102),clock=>clock,reset=>reset,s=>p(250)(102),cout=>p(251)(103));
FA_ff_7764:FAff port map(x=>p(182)(103),y=>p(183)(103),Cin=>p(184)(103),clock=>clock,reset=>reset,s=>p(250)(103),cout=>p(251)(104));
FA_ff_7765:FAff port map(x=>p(182)(104),y=>p(183)(104),Cin=>p(184)(104),clock=>clock,reset=>reset,s=>p(250)(104),cout=>p(251)(105));
FA_ff_7766:FAff port map(x=>p(182)(105),y=>p(183)(105),Cin=>p(184)(105),clock=>clock,reset=>reset,s=>p(250)(105),cout=>p(251)(106));
FA_ff_7767:FAff port map(x=>p(182)(106),y=>p(183)(106),Cin=>p(184)(106),clock=>clock,reset=>reset,s=>p(250)(106),cout=>p(251)(107));
FA_ff_7768:FAff port map(x=>p(182)(107),y=>p(183)(107),Cin=>p(184)(107),clock=>clock,reset=>reset,s=>p(250)(107),cout=>p(251)(108));
FA_ff_7769:FAff port map(x=>p(182)(108),y=>p(183)(108),Cin=>p(184)(108),clock=>clock,reset=>reset,s=>p(250)(108),cout=>p(251)(109));
FA_ff_7770:FAff port map(x=>p(182)(109),y=>p(183)(109),Cin=>p(184)(109),clock=>clock,reset=>reset,s=>p(250)(109),cout=>p(251)(110));
FA_ff_7771:FAff port map(x=>p(182)(110),y=>p(183)(110),Cin=>p(184)(110),clock=>clock,reset=>reset,s=>p(250)(110),cout=>p(251)(111));
FA_ff_7772:FAff port map(x=>p(182)(111),y=>p(183)(111),Cin=>p(184)(111),clock=>clock,reset=>reset,s=>p(250)(111),cout=>p(251)(112));
FA_ff_7773:FAff port map(x=>p(182)(112),y=>p(183)(112),Cin=>p(184)(112),clock=>clock,reset=>reset,s=>p(250)(112),cout=>p(251)(113));
FA_ff_7774:FAff port map(x=>p(182)(113),y=>p(183)(113),Cin=>p(184)(113),clock=>clock,reset=>reset,s=>p(250)(113),cout=>p(251)(114));
FA_ff_7775:FAff port map(x=>p(182)(114),y=>p(183)(114),Cin=>p(184)(114),clock=>clock,reset=>reset,s=>p(250)(114),cout=>p(251)(115));
FA_ff_7776:FAff port map(x=>p(182)(115),y=>p(183)(115),Cin=>p(184)(115),clock=>clock,reset=>reset,s=>p(250)(115),cout=>p(251)(116));
FA_ff_7777:FAff port map(x=>p(182)(116),y=>p(183)(116),Cin=>p(184)(116),clock=>clock,reset=>reset,s=>p(250)(116),cout=>p(251)(117));
FA_ff_7778:FAff port map(x=>p(182)(117),y=>p(183)(117),Cin=>p(184)(117),clock=>clock,reset=>reset,s=>p(250)(117),cout=>p(251)(118));
FA_ff_7779:FAff port map(x=>p(182)(118),y=>p(183)(118),Cin=>p(184)(118),clock=>clock,reset=>reset,s=>p(250)(118),cout=>p(251)(119));
FA_ff_7780:FAff port map(x=>p(182)(119),y=>p(183)(119),Cin=>p(184)(119),clock=>clock,reset=>reset,s=>p(250)(119),cout=>p(251)(120));
FA_ff_7781:FAff port map(x=>p(182)(120),y=>p(183)(120),Cin=>p(184)(120),clock=>clock,reset=>reset,s=>p(250)(120),cout=>p(251)(121));
FA_ff_7782:FAff port map(x=>p(182)(121),y=>p(183)(121),Cin=>p(184)(121),clock=>clock,reset=>reset,s=>p(250)(121),cout=>p(251)(122));
FA_ff_7783:FAff port map(x=>p(182)(122),y=>p(183)(122),Cin=>p(184)(122),clock=>clock,reset=>reset,s=>p(250)(122),cout=>p(251)(123));
FA_ff_7784:FAff port map(x=>p(182)(123),y=>p(183)(123),Cin=>p(184)(123),clock=>clock,reset=>reset,s=>p(250)(123),cout=>p(251)(124));
FA_ff_7785:FAff port map(x=>p(182)(124),y=>p(183)(124),Cin=>p(184)(124),clock=>clock,reset=>reset,s=>p(250)(124),cout=>p(251)(125));
FA_ff_7786:FAff port map(x=>p(182)(125),y=>p(183)(125),Cin=>p(184)(125),clock=>clock,reset=>reset,s=>p(250)(125),cout=>p(251)(126));
FA_ff_7787:FAff port map(x=>p(182)(126),y=>p(183)(126),Cin=>p(184)(126),clock=>clock,reset=>reset,s=>p(250)(126),cout=>p(251)(127));
FA_ff_7788:FAff port map(x=>p(182)(127),y=>p(183)(127),Cin=>p(184)(127),clock=>clock,reset=>reset,s=>p(250)(127),cout=>p(251)(128));
p(250)(128)<=p(183)(128);
p(252)(0)<=p(186)(0);
FA_ff_7789:FAff port map(x=>p(185)(1),y=>p(186)(1),Cin=>p(187)(1),clock=>clock,reset=>reset,s=>p(252)(1),cout=>p(253)(2));
FA_ff_7790:FAff port map(x=>p(185)(2),y=>p(186)(2),Cin=>p(187)(2),clock=>clock,reset=>reset,s=>p(252)(2),cout=>p(253)(3));
FA_ff_7791:FAff port map(x=>p(185)(3),y=>p(186)(3),Cin=>p(187)(3),clock=>clock,reset=>reset,s=>p(252)(3),cout=>p(253)(4));
FA_ff_7792:FAff port map(x=>p(185)(4),y=>p(186)(4),Cin=>p(187)(4),clock=>clock,reset=>reset,s=>p(252)(4),cout=>p(253)(5));
FA_ff_7793:FAff port map(x=>p(185)(5),y=>p(186)(5),Cin=>p(187)(5),clock=>clock,reset=>reset,s=>p(252)(5),cout=>p(253)(6));
FA_ff_7794:FAff port map(x=>p(185)(6),y=>p(186)(6),Cin=>p(187)(6),clock=>clock,reset=>reset,s=>p(252)(6),cout=>p(253)(7));
FA_ff_7795:FAff port map(x=>p(185)(7),y=>p(186)(7),Cin=>p(187)(7),clock=>clock,reset=>reset,s=>p(252)(7),cout=>p(253)(8));
FA_ff_7796:FAff port map(x=>p(185)(8),y=>p(186)(8),Cin=>p(187)(8),clock=>clock,reset=>reset,s=>p(252)(8),cout=>p(253)(9));
FA_ff_7797:FAff port map(x=>p(185)(9),y=>p(186)(9),Cin=>p(187)(9),clock=>clock,reset=>reset,s=>p(252)(9),cout=>p(253)(10));
FA_ff_7798:FAff port map(x=>p(185)(10),y=>p(186)(10),Cin=>p(187)(10),clock=>clock,reset=>reset,s=>p(252)(10),cout=>p(253)(11));
FA_ff_7799:FAff port map(x=>p(185)(11),y=>p(186)(11),Cin=>p(187)(11),clock=>clock,reset=>reset,s=>p(252)(11),cout=>p(253)(12));
FA_ff_7800:FAff port map(x=>p(185)(12),y=>p(186)(12),Cin=>p(187)(12),clock=>clock,reset=>reset,s=>p(252)(12),cout=>p(253)(13));
FA_ff_7801:FAff port map(x=>p(185)(13),y=>p(186)(13),Cin=>p(187)(13),clock=>clock,reset=>reset,s=>p(252)(13),cout=>p(253)(14));
FA_ff_7802:FAff port map(x=>p(185)(14),y=>p(186)(14),Cin=>p(187)(14),clock=>clock,reset=>reset,s=>p(252)(14),cout=>p(253)(15));
FA_ff_7803:FAff port map(x=>p(185)(15),y=>p(186)(15),Cin=>p(187)(15),clock=>clock,reset=>reset,s=>p(252)(15),cout=>p(253)(16));
FA_ff_7804:FAff port map(x=>p(185)(16),y=>p(186)(16),Cin=>p(187)(16),clock=>clock,reset=>reset,s=>p(252)(16),cout=>p(253)(17));
FA_ff_7805:FAff port map(x=>p(185)(17),y=>p(186)(17),Cin=>p(187)(17),clock=>clock,reset=>reset,s=>p(252)(17),cout=>p(253)(18));
FA_ff_7806:FAff port map(x=>p(185)(18),y=>p(186)(18),Cin=>p(187)(18),clock=>clock,reset=>reset,s=>p(252)(18),cout=>p(253)(19));
FA_ff_7807:FAff port map(x=>p(185)(19),y=>p(186)(19),Cin=>p(187)(19),clock=>clock,reset=>reset,s=>p(252)(19),cout=>p(253)(20));
FA_ff_7808:FAff port map(x=>p(185)(20),y=>p(186)(20),Cin=>p(187)(20),clock=>clock,reset=>reset,s=>p(252)(20),cout=>p(253)(21));
FA_ff_7809:FAff port map(x=>p(185)(21),y=>p(186)(21),Cin=>p(187)(21),clock=>clock,reset=>reset,s=>p(252)(21),cout=>p(253)(22));
FA_ff_7810:FAff port map(x=>p(185)(22),y=>p(186)(22),Cin=>p(187)(22),clock=>clock,reset=>reset,s=>p(252)(22),cout=>p(253)(23));
FA_ff_7811:FAff port map(x=>p(185)(23),y=>p(186)(23),Cin=>p(187)(23),clock=>clock,reset=>reset,s=>p(252)(23),cout=>p(253)(24));
FA_ff_7812:FAff port map(x=>p(185)(24),y=>p(186)(24),Cin=>p(187)(24),clock=>clock,reset=>reset,s=>p(252)(24),cout=>p(253)(25));
FA_ff_7813:FAff port map(x=>p(185)(25),y=>p(186)(25),Cin=>p(187)(25),clock=>clock,reset=>reset,s=>p(252)(25),cout=>p(253)(26));
FA_ff_7814:FAff port map(x=>p(185)(26),y=>p(186)(26),Cin=>p(187)(26),clock=>clock,reset=>reset,s=>p(252)(26),cout=>p(253)(27));
FA_ff_7815:FAff port map(x=>p(185)(27),y=>p(186)(27),Cin=>p(187)(27),clock=>clock,reset=>reset,s=>p(252)(27),cout=>p(253)(28));
FA_ff_7816:FAff port map(x=>p(185)(28),y=>p(186)(28),Cin=>p(187)(28),clock=>clock,reset=>reset,s=>p(252)(28),cout=>p(253)(29));
FA_ff_7817:FAff port map(x=>p(185)(29),y=>p(186)(29),Cin=>p(187)(29),clock=>clock,reset=>reset,s=>p(252)(29),cout=>p(253)(30));
FA_ff_7818:FAff port map(x=>p(185)(30),y=>p(186)(30),Cin=>p(187)(30),clock=>clock,reset=>reset,s=>p(252)(30),cout=>p(253)(31));
FA_ff_7819:FAff port map(x=>p(185)(31),y=>p(186)(31),Cin=>p(187)(31),clock=>clock,reset=>reset,s=>p(252)(31),cout=>p(253)(32));
FA_ff_7820:FAff port map(x=>p(185)(32),y=>p(186)(32),Cin=>p(187)(32),clock=>clock,reset=>reset,s=>p(252)(32),cout=>p(253)(33));
FA_ff_7821:FAff port map(x=>p(185)(33),y=>p(186)(33),Cin=>p(187)(33),clock=>clock,reset=>reset,s=>p(252)(33),cout=>p(253)(34));
FA_ff_7822:FAff port map(x=>p(185)(34),y=>p(186)(34),Cin=>p(187)(34),clock=>clock,reset=>reset,s=>p(252)(34),cout=>p(253)(35));
FA_ff_7823:FAff port map(x=>p(185)(35),y=>p(186)(35),Cin=>p(187)(35),clock=>clock,reset=>reset,s=>p(252)(35),cout=>p(253)(36));
FA_ff_7824:FAff port map(x=>p(185)(36),y=>p(186)(36),Cin=>p(187)(36),clock=>clock,reset=>reset,s=>p(252)(36),cout=>p(253)(37));
FA_ff_7825:FAff port map(x=>p(185)(37),y=>p(186)(37),Cin=>p(187)(37),clock=>clock,reset=>reset,s=>p(252)(37),cout=>p(253)(38));
FA_ff_7826:FAff port map(x=>p(185)(38),y=>p(186)(38),Cin=>p(187)(38),clock=>clock,reset=>reset,s=>p(252)(38),cout=>p(253)(39));
FA_ff_7827:FAff port map(x=>p(185)(39),y=>p(186)(39),Cin=>p(187)(39),clock=>clock,reset=>reset,s=>p(252)(39),cout=>p(253)(40));
FA_ff_7828:FAff port map(x=>p(185)(40),y=>p(186)(40),Cin=>p(187)(40),clock=>clock,reset=>reset,s=>p(252)(40),cout=>p(253)(41));
FA_ff_7829:FAff port map(x=>p(185)(41),y=>p(186)(41),Cin=>p(187)(41),clock=>clock,reset=>reset,s=>p(252)(41),cout=>p(253)(42));
FA_ff_7830:FAff port map(x=>p(185)(42),y=>p(186)(42),Cin=>p(187)(42),clock=>clock,reset=>reset,s=>p(252)(42),cout=>p(253)(43));
FA_ff_7831:FAff port map(x=>p(185)(43),y=>p(186)(43),Cin=>p(187)(43),clock=>clock,reset=>reset,s=>p(252)(43),cout=>p(253)(44));
FA_ff_7832:FAff port map(x=>p(185)(44),y=>p(186)(44),Cin=>p(187)(44),clock=>clock,reset=>reset,s=>p(252)(44),cout=>p(253)(45));
FA_ff_7833:FAff port map(x=>p(185)(45),y=>p(186)(45),Cin=>p(187)(45),clock=>clock,reset=>reset,s=>p(252)(45),cout=>p(253)(46));
FA_ff_7834:FAff port map(x=>p(185)(46),y=>p(186)(46),Cin=>p(187)(46),clock=>clock,reset=>reset,s=>p(252)(46),cout=>p(253)(47));
FA_ff_7835:FAff port map(x=>p(185)(47),y=>p(186)(47),Cin=>p(187)(47),clock=>clock,reset=>reset,s=>p(252)(47),cout=>p(253)(48));
FA_ff_7836:FAff port map(x=>p(185)(48),y=>p(186)(48),Cin=>p(187)(48),clock=>clock,reset=>reset,s=>p(252)(48),cout=>p(253)(49));
FA_ff_7837:FAff port map(x=>p(185)(49),y=>p(186)(49),Cin=>p(187)(49),clock=>clock,reset=>reset,s=>p(252)(49),cout=>p(253)(50));
FA_ff_7838:FAff port map(x=>p(185)(50),y=>p(186)(50),Cin=>p(187)(50),clock=>clock,reset=>reset,s=>p(252)(50),cout=>p(253)(51));
FA_ff_7839:FAff port map(x=>p(185)(51),y=>p(186)(51),Cin=>p(187)(51),clock=>clock,reset=>reset,s=>p(252)(51),cout=>p(253)(52));
FA_ff_7840:FAff port map(x=>p(185)(52),y=>p(186)(52),Cin=>p(187)(52),clock=>clock,reset=>reset,s=>p(252)(52),cout=>p(253)(53));
FA_ff_7841:FAff port map(x=>p(185)(53),y=>p(186)(53),Cin=>p(187)(53),clock=>clock,reset=>reset,s=>p(252)(53),cout=>p(253)(54));
FA_ff_7842:FAff port map(x=>p(185)(54),y=>p(186)(54),Cin=>p(187)(54),clock=>clock,reset=>reset,s=>p(252)(54),cout=>p(253)(55));
FA_ff_7843:FAff port map(x=>p(185)(55),y=>p(186)(55),Cin=>p(187)(55),clock=>clock,reset=>reset,s=>p(252)(55),cout=>p(253)(56));
FA_ff_7844:FAff port map(x=>p(185)(56),y=>p(186)(56),Cin=>p(187)(56),clock=>clock,reset=>reset,s=>p(252)(56),cout=>p(253)(57));
FA_ff_7845:FAff port map(x=>p(185)(57),y=>p(186)(57),Cin=>p(187)(57),clock=>clock,reset=>reset,s=>p(252)(57),cout=>p(253)(58));
FA_ff_7846:FAff port map(x=>p(185)(58),y=>p(186)(58),Cin=>p(187)(58),clock=>clock,reset=>reset,s=>p(252)(58),cout=>p(253)(59));
FA_ff_7847:FAff port map(x=>p(185)(59),y=>p(186)(59),Cin=>p(187)(59),clock=>clock,reset=>reset,s=>p(252)(59),cout=>p(253)(60));
FA_ff_7848:FAff port map(x=>p(185)(60),y=>p(186)(60),Cin=>p(187)(60),clock=>clock,reset=>reset,s=>p(252)(60),cout=>p(253)(61));
FA_ff_7849:FAff port map(x=>p(185)(61),y=>p(186)(61),Cin=>p(187)(61),clock=>clock,reset=>reset,s=>p(252)(61),cout=>p(253)(62));
FA_ff_7850:FAff port map(x=>p(185)(62),y=>p(186)(62),Cin=>p(187)(62),clock=>clock,reset=>reset,s=>p(252)(62),cout=>p(253)(63));
FA_ff_7851:FAff port map(x=>p(185)(63),y=>p(186)(63),Cin=>p(187)(63),clock=>clock,reset=>reset,s=>p(252)(63),cout=>p(253)(64));
FA_ff_7852:FAff port map(x=>p(185)(64),y=>p(186)(64),Cin=>p(187)(64),clock=>clock,reset=>reset,s=>p(252)(64),cout=>p(253)(65));
FA_ff_7853:FAff port map(x=>p(185)(65),y=>p(186)(65),Cin=>p(187)(65),clock=>clock,reset=>reset,s=>p(252)(65),cout=>p(253)(66));
FA_ff_7854:FAff port map(x=>p(185)(66),y=>p(186)(66),Cin=>p(187)(66),clock=>clock,reset=>reset,s=>p(252)(66),cout=>p(253)(67));
FA_ff_7855:FAff port map(x=>p(185)(67),y=>p(186)(67),Cin=>p(187)(67),clock=>clock,reset=>reset,s=>p(252)(67),cout=>p(253)(68));
FA_ff_7856:FAff port map(x=>p(185)(68),y=>p(186)(68),Cin=>p(187)(68),clock=>clock,reset=>reset,s=>p(252)(68),cout=>p(253)(69));
FA_ff_7857:FAff port map(x=>p(185)(69),y=>p(186)(69),Cin=>p(187)(69),clock=>clock,reset=>reset,s=>p(252)(69),cout=>p(253)(70));
FA_ff_7858:FAff port map(x=>p(185)(70),y=>p(186)(70),Cin=>p(187)(70),clock=>clock,reset=>reset,s=>p(252)(70),cout=>p(253)(71));
FA_ff_7859:FAff port map(x=>p(185)(71),y=>p(186)(71),Cin=>p(187)(71),clock=>clock,reset=>reset,s=>p(252)(71),cout=>p(253)(72));
FA_ff_7860:FAff port map(x=>p(185)(72),y=>p(186)(72),Cin=>p(187)(72),clock=>clock,reset=>reset,s=>p(252)(72),cout=>p(253)(73));
FA_ff_7861:FAff port map(x=>p(185)(73),y=>p(186)(73),Cin=>p(187)(73),clock=>clock,reset=>reset,s=>p(252)(73),cout=>p(253)(74));
FA_ff_7862:FAff port map(x=>p(185)(74),y=>p(186)(74),Cin=>p(187)(74),clock=>clock,reset=>reset,s=>p(252)(74),cout=>p(253)(75));
FA_ff_7863:FAff port map(x=>p(185)(75),y=>p(186)(75),Cin=>p(187)(75),clock=>clock,reset=>reset,s=>p(252)(75),cout=>p(253)(76));
FA_ff_7864:FAff port map(x=>p(185)(76),y=>p(186)(76),Cin=>p(187)(76),clock=>clock,reset=>reset,s=>p(252)(76),cout=>p(253)(77));
FA_ff_7865:FAff port map(x=>p(185)(77),y=>p(186)(77),Cin=>p(187)(77),clock=>clock,reset=>reset,s=>p(252)(77),cout=>p(253)(78));
FA_ff_7866:FAff port map(x=>p(185)(78),y=>p(186)(78),Cin=>p(187)(78),clock=>clock,reset=>reset,s=>p(252)(78),cout=>p(253)(79));
FA_ff_7867:FAff port map(x=>p(185)(79),y=>p(186)(79),Cin=>p(187)(79),clock=>clock,reset=>reset,s=>p(252)(79),cout=>p(253)(80));
FA_ff_7868:FAff port map(x=>p(185)(80),y=>p(186)(80),Cin=>p(187)(80),clock=>clock,reset=>reset,s=>p(252)(80),cout=>p(253)(81));
FA_ff_7869:FAff port map(x=>p(185)(81),y=>p(186)(81),Cin=>p(187)(81),clock=>clock,reset=>reset,s=>p(252)(81),cout=>p(253)(82));
FA_ff_7870:FAff port map(x=>p(185)(82),y=>p(186)(82),Cin=>p(187)(82),clock=>clock,reset=>reset,s=>p(252)(82),cout=>p(253)(83));
FA_ff_7871:FAff port map(x=>p(185)(83),y=>p(186)(83),Cin=>p(187)(83),clock=>clock,reset=>reset,s=>p(252)(83),cout=>p(253)(84));
FA_ff_7872:FAff port map(x=>p(185)(84),y=>p(186)(84),Cin=>p(187)(84),clock=>clock,reset=>reset,s=>p(252)(84),cout=>p(253)(85));
FA_ff_7873:FAff port map(x=>p(185)(85),y=>p(186)(85),Cin=>p(187)(85),clock=>clock,reset=>reset,s=>p(252)(85),cout=>p(253)(86));
FA_ff_7874:FAff port map(x=>p(185)(86),y=>p(186)(86),Cin=>p(187)(86),clock=>clock,reset=>reset,s=>p(252)(86),cout=>p(253)(87));
FA_ff_7875:FAff port map(x=>p(185)(87),y=>p(186)(87),Cin=>p(187)(87),clock=>clock,reset=>reset,s=>p(252)(87),cout=>p(253)(88));
FA_ff_7876:FAff port map(x=>p(185)(88),y=>p(186)(88),Cin=>p(187)(88),clock=>clock,reset=>reset,s=>p(252)(88),cout=>p(253)(89));
FA_ff_7877:FAff port map(x=>p(185)(89),y=>p(186)(89),Cin=>p(187)(89),clock=>clock,reset=>reset,s=>p(252)(89),cout=>p(253)(90));
FA_ff_7878:FAff port map(x=>p(185)(90),y=>p(186)(90),Cin=>p(187)(90),clock=>clock,reset=>reset,s=>p(252)(90),cout=>p(253)(91));
FA_ff_7879:FAff port map(x=>p(185)(91),y=>p(186)(91),Cin=>p(187)(91),clock=>clock,reset=>reset,s=>p(252)(91),cout=>p(253)(92));
FA_ff_7880:FAff port map(x=>p(185)(92),y=>p(186)(92),Cin=>p(187)(92),clock=>clock,reset=>reset,s=>p(252)(92),cout=>p(253)(93));
FA_ff_7881:FAff port map(x=>p(185)(93),y=>p(186)(93),Cin=>p(187)(93),clock=>clock,reset=>reset,s=>p(252)(93),cout=>p(253)(94));
FA_ff_7882:FAff port map(x=>p(185)(94),y=>p(186)(94),Cin=>p(187)(94),clock=>clock,reset=>reset,s=>p(252)(94),cout=>p(253)(95));
FA_ff_7883:FAff port map(x=>p(185)(95),y=>p(186)(95),Cin=>p(187)(95),clock=>clock,reset=>reset,s=>p(252)(95),cout=>p(253)(96));
FA_ff_7884:FAff port map(x=>p(185)(96),y=>p(186)(96),Cin=>p(187)(96),clock=>clock,reset=>reset,s=>p(252)(96),cout=>p(253)(97));
FA_ff_7885:FAff port map(x=>p(185)(97),y=>p(186)(97),Cin=>p(187)(97),clock=>clock,reset=>reset,s=>p(252)(97),cout=>p(253)(98));
FA_ff_7886:FAff port map(x=>p(185)(98),y=>p(186)(98),Cin=>p(187)(98),clock=>clock,reset=>reset,s=>p(252)(98),cout=>p(253)(99));
FA_ff_7887:FAff port map(x=>p(185)(99),y=>p(186)(99),Cin=>p(187)(99),clock=>clock,reset=>reset,s=>p(252)(99),cout=>p(253)(100));
FA_ff_7888:FAff port map(x=>p(185)(100),y=>p(186)(100),Cin=>p(187)(100),clock=>clock,reset=>reset,s=>p(252)(100),cout=>p(253)(101));
FA_ff_7889:FAff port map(x=>p(185)(101),y=>p(186)(101),Cin=>p(187)(101),clock=>clock,reset=>reset,s=>p(252)(101),cout=>p(253)(102));
FA_ff_7890:FAff port map(x=>p(185)(102),y=>p(186)(102),Cin=>p(187)(102),clock=>clock,reset=>reset,s=>p(252)(102),cout=>p(253)(103));
FA_ff_7891:FAff port map(x=>p(185)(103),y=>p(186)(103),Cin=>p(187)(103),clock=>clock,reset=>reset,s=>p(252)(103),cout=>p(253)(104));
FA_ff_7892:FAff port map(x=>p(185)(104),y=>p(186)(104),Cin=>p(187)(104),clock=>clock,reset=>reset,s=>p(252)(104),cout=>p(253)(105));
FA_ff_7893:FAff port map(x=>p(185)(105),y=>p(186)(105),Cin=>p(187)(105),clock=>clock,reset=>reset,s=>p(252)(105),cout=>p(253)(106));
FA_ff_7894:FAff port map(x=>p(185)(106),y=>p(186)(106),Cin=>p(187)(106),clock=>clock,reset=>reset,s=>p(252)(106),cout=>p(253)(107));
FA_ff_7895:FAff port map(x=>p(185)(107),y=>p(186)(107),Cin=>p(187)(107),clock=>clock,reset=>reset,s=>p(252)(107),cout=>p(253)(108));
FA_ff_7896:FAff port map(x=>p(185)(108),y=>p(186)(108),Cin=>p(187)(108),clock=>clock,reset=>reset,s=>p(252)(108),cout=>p(253)(109));
FA_ff_7897:FAff port map(x=>p(185)(109),y=>p(186)(109),Cin=>p(187)(109),clock=>clock,reset=>reset,s=>p(252)(109),cout=>p(253)(110));
FA_ff_7898:FAff port map(x=>p(185)(110),y=>p(186)(110),Cin=>p(187)(110),clock=>clock,reset=>reset,s=>p(252)(110),cout=>p(253)(111));
FA_ff_7899:FAff port map(x=>p(185)(111),y=>p(186)(111),Cin=>p(187)(111),clock=>clock,reset=>reset,s=>p(252)(111),cout=>p(253)(112));
FA_ff_7900:FAff port map(x=>p(185)(112),y=>p(186)(112),Cin=>p(187)(112),clock=>clock,reset=>reset,s=>p(252)(112),cout=>p(253)(113));
FA_ff_7901:FAff port map(x=>p(185)(113),y=>p(186)(113),Cin=>p(187)(113),clock=>clock,reset=>reset,s=>p(252)(113),cout=>p(253)(114));
FA_ff_7902:FAff port map(x=>p(185)(114),y=>p(186)(114),Cin=>p(187)(114),clock=>clock,reset=>reset,s=>p(252)(114),cout=>p(253)(115));
FA_ff_7903:FAff port map(x=>p(185)(115),y=>p(186)(115),Cin=>p(187)(115),clock=>clock,reset=>reset,s=>p(252)(115),cout=>p(253)(116));
FA_ff_7904:FAff port map(x=>p(185)(116),y=>p(186)(116),Cin=>p(187)(116),clock=>clock,reset=>reset,s=>p(252)(116),cout=>p(253)(117));
FA_ff_7905:FAff port map(x=>p(185)(117),y=>p(186)(117),Cin=>p(187)(117),clock=>clock,reset=>reset,s=>p(252)(117),cout=>p(253)(118));
FA_ff_7906:FAff port map(x=>p(185)(118),y=>p(186)(118),Cin=>p(187)(118),clock=>clock,reset=>reset,s=>p(252)(118),cout=>p(253)(119));
FA_ff_7907:FAff port map(x=>p(185)(119),y=>p(186)(119),Cin=>p(187)(119),clock=>clock,reset=>reset,s=>p(252)(119),cout=>p(253)(120));
FA_ff_7908:FAff port map(x=>p(185)(120),y=>p(186)(120),Cin=>p(187)(120),clock=>clock,reset=>reset,s=>p(252)(120),cout=>p(253)(121));
FA_ff_7909:FAff port map(x=>p(185)(121),y=>p(186)(121),Cin=>p(187)(121),clock=>clock,reset=>reset,s=>p(252)(121),cout=>p(253)(122));
FA_ff_7910:FAff port map(x=>p(185)(122),y=>p(186)(122),Cin=>p(187)(122),clock=>clock,reset=>reset,s=>p(252)(122),cout=>p(253)(123));
FA_ff_7911:FAff port map(x=>p(185)(123),y=>p(186)(123),Cin=>p(187)(123),clock=>clock,reset=>reset,s=>p(252)(123),cout=>p(253)(124));
FA_ff_7912:FAff port map(x=>p(185)(124),y=>p(186)(124),Cin=>p(187)(124),clock=>clock,reset=>reset,s=>p(252)(124),cout=>p(253)(125));
FA_ff_7913:FAff port map(x=>p(185)(125),y=>p(186)(125),Cin=>p(187)(125),clock=>clock,reset=>reset,s=>p(252)(125),cout=>p(253)(126));
FA_ff_7914:FAff port map(x=>p(185)(126),y=>p(186)(126),Cin=>p(187)(126),clock=>clock,reset=>reset,s=>p(252)(126),cout=>p(253)(127));
FA_ff_7915:FAff port map(x=>p(185)(127),y=>p(186)(127),Cin=>p(187)(127),clock=>clock,reset=>reset,s=>p(252)(127),cout=>p(253)(128));
HA_ff_19:HAff port map(x=>p(185)(128),y=>p(187)(128),clock=>clock,reset=>reset,s=>p(252)(128),c=>p(253)(129));
HA_ff_20:HAff port map(x=>p(188)(0),y=>p(190)(0),clock=>clock,reset=>reset,s=>p(254)(0),c=>p(255)(1));
FA_ff_7916:FAff port map(x=>p(188)(1),y=>p(189)(1),Cin=>p(190)(1),clock=>clock,reset=>reset,s=>p(254)(1),cout=>p(255)(2));
FA_ff_7917:FAff port map(x=>p(188)(2),y=>p(189)(2),Cin=>p(190)(2),clock=>clock,reset=>reset,s=>p(254)(2),cout=>p(255)(3));
FA_ff_7918:FAff port map(x=>p(188)(3),y=>p(189)(3),Cin=>p(190)(3),clock=>clock,reset=>reset,s=>p(254)(3),cout=>p(255)(4));
FA_ff_7919:FAff port map(x=>p(188)(4),y=>p(189)(4),Cin=>p(190)(4),clock=>clock,reset=>reset,s=>p(254)(4),cout=>p(255)(5));
FA_ff_7920:FAff port map(x=>p(188)(5),y=>p(189)(5),Cin=>p(190)(5),clock=>clock,reset=>reset,s=>p(254)(5),cout=>p(255)(6));
FA_ff_7921:FAff port map(x=>p(188)(6),y=>p(189)(6),Cin=>p(190)(6),clock=>clock,reset=>reset,s=>p(254)(6),cout=>p(255)(7));
FA_ff_7922:FAff port map(x=>p(188)(7),y=>p(189)(7),Cin=>p(190)(7),clock=>clock,reset=>reset,s=>p(254)(7),cout=>p(255)(8));
FA_ff_7923:FAff port map(x=>p(188)(8),y=>p(189)(8),Cin=>p(190)(8),clock=>clock,reset=>reset,s=>p(254)(8),cout=>p(255)(9));
FA_ff_7924:FAff port map(x=>p(188)(9),y=>p(189)(9),Cin=>p(190)(9),clock=>clock,reset=>reset,s=>p(254)(9),cout=>p(255)(10));
FA_ff_7925:FAff port map(x=>p(188)(10),y=>p(189)(10),Cin=>p(190)(10),clock=>clock,reset=>reset,s=>p(254)(10),cout=>p(255)(11));
FA_ff_7926:FAff port map(x=>p(188)(11),y=>p(189)(11),Cin=>p(190)(11),clock=>clock,reset=>reset,s=>p(254)(11),cout=>p(255)(12));
FA_ff_7927:FAff port map(x=>p(188)(12),y=>p(189)(12),Cin=>p(190)(12),clock=>clock,reset=>reset,s=>p(254)(12),cout=>p(255)(13));
FA_ff_7928:FAff port map(x=>p(188)(13),y=>p(189)(13),Cin=>p(190)(13),clock=>clock,reset=>reset,s=>p(254)(13),cout=>p(255)(14));
FA_ff_7929:FAff port map(x=>p(188)(14),y=>p(189)(14),Cin=>p(190)(14),clock=>clock,reset=>reset,s=>p(254)(14),cout=>p(255)(15));
FA_ff_7930:FAff port map(x=>p(188)(15),y=>p(189)(15),Cin=>p(190)(15),clock=>clock,reset=>reset,s=>p(254)(15),cout=>p(255)(16));
FA_ff_7931:FAff port map(x=>p(188)(16),y=>p(189)(16),Cin=>p(190)(16),clock=>clock,reset=>reset,s=>p(254)(16),cout=>p(255)(17));
FA_ff_7932:FAff port map(x=>p(188)(17),y=>p(189)(17),Cin=>p(190)(17),clock=>clock,reset=>reset,s=>p(254)(17),cout=>p(255)(18));
FA_ff_7933:FAff port map(x=>p(188)(18),y=>p(189)(18),Cin=>p(190)(18),clock=>clock,reset=>reset,s=>p(254)(18),cout=>p(255)(19));
FA_ff_7934:FAff port map(x=>p(188)(19),y=>p(189)(19),Cin=>p(190)(19),clock=>clock,reset=>reset,s=>p(254)(19),cout=>p(255)(20));
FA_ff_7935:FAff port map(x=>p(188)(20),y=>p(189)(20),Cin=>p(190)(20),clock=>clock,reset=>reset,s=>p(254)(20),cout=>p(255)(21));
FA_ff_7936:FAff port map(x=>p(188)(21),y=>p(189)(21),Cin=>p(190)(21),clock=>clock,reset=>reset,s=>p(254)(21),cout=>p(255)(22));
FA_ff_7937:FAff port map(x=>p(188)(22),y=>p(189)(22),Cin=>p(190)(22),clock=>clock,reset=>reset,s=>p(254)(22),cout=>p(255)(23));
FA_ff_7938:FAff port map(x=>p(188)(23),y=>p(189)(23),Cin=>p(190)(23),clock=>clock,reset=>reset,s=>p(254)(23),cout=>p(255)(24));
FA_ff_7939:FAff port map(x=>p(188)(24),y=>p(189)(24),Cin=>p(190)(24),clock=>clock,reset=>reset,s=>p(254)(24),cout=>p(255)(25));
FA_ff_7940:FAff port map(x=>p(188)(25),y=>p(189)(25),Cin=>p(190)(25),clock=>clock,reset=>reset,s=>p(254)(25),cout=>p(255)(26));
FA_ff_7941:FAff port map(x=>p(188)(26),y=>p(189)(26),Cin=>p(190)(26),clock=>clock,reset=>reset,s=>p(254)(26),cout=>p(255)(27));
FA_ff_7942:FAff port map(x=>p(188)(27),y=>p(189)(27),Cin=>p(190)(27),clock=>clock,reset=>reset,s=>p(254)(27),cout=>p(255)(28));
FA_ff_7943:FAff port map(x=>p(188)(28),y=>p(189)(28),Cin=>p(190)(28),clock=>clock,reset=>reset,s=>p(254)(28),cout=>p(255)(29));
FA_ff_7944:FAff port map(x=>p(188)(29),y=>p(189)(29),Cin=>p(190)(29),clock=>clock,reset=>reset,s=>p(254)(29),cout=>p(255)(30));
FA_ff_7945:FAff port map(x=>p(188)(30),y=>p(189)(30),Cin=>p(190)(30),clock=>clock,reset=>reset,s=>p(254)(30),cout=>p(255)(31));
FA_ff_7946:FAff port map(x=>p(188)(31),y=>p(189)(31),Cin=>p(190)(31),clock=>clock,reset=>reset,s=>p(254)(31),cout=>p(255)(32));
FA_ff_7947:FAff port map(x=>p(188)(32),y=>p(189)(32),Cin=>p(190)(32),clock=>clock,reset=>reset,s=>p(254)(32),cout=>p(255)(33));
FA_ff_7948:FAff port map(x=>p(188)(33),y=>p(189)(33),Cin=>p(190)(33),clock=>clock,reset=>reset,s=>p(254)(33),cout=>p(255)(34));
FA_ff_7949:FAff port map(x=>p(188)(34),y=>p(189)(34),Cin=>p(190)(34),clock=>clock,reset=>reset,s=>p(254)(34),cout=>p(255)(35));
FA_ff_7950:FAff port map(x=>p(188)(35),y=>p(189)(35),Cin=>p(190)(35),clock=>clock,reset=>reset,s=>p(254)(35),cout=>p(255)(36));
FA_ff_7951:FAff port map(x=>p(188)(36),y=>p(189)(36),Cin=>p(190)(36),clock=>clock,reset=>reset,s=>p(254)(36),cout=>p(255)(37));
FA_ff_7952:FAff port map(x=>p(188)(37),y=>p(189)(37),Cin=>p(190)(37),clock=>clock,reset=>reset,s=>p(254)(37),cout=>p(255)(38));
FA_ff_7953:FAff port map(x=>p(188)(38),y=>p(189)(38),Cin=>p(190)(38),clock=>clock,reset=>reset,s=>p(254)(38),cout=>p(255)(39));
FA_ff_7954:FAff port map(x=>p(188)(39),y=>p(189)(39),Cin=>p(190)(39),clock=>clock,reset=>reset,s=>p(254)(39),cout=>p(255)(40));
FA_ff_7955:FAff port map(x=>p(188)(40),y=>p(189)(40),Cin=>p(190)(40),clock=>clock,reset=>reset,s=>p(254)(40),cout=>p(255)(41));
FA_ff_7956:FAff port map(x=>p(188)(41),y=>p(189)(41),Cin=>p(190)(41),clock=>clock,reset=>reset,s=>p(254)(41),cout=>p(255)(42));
FA_ff_7957:FAff port map(x=>p(188)(42),y=>p(189)(42),Cin=>p(190)(42),clock=>clock,reset=>reset,s=>p(254)(42),cout=>p(255)(43));
FA_ff_7958:FAff port map(x=>p(188)(43),y=>p(189)(43),Cin=>p(190)(43),clock=>clock,reset=>reset,s=>p(254)(43),cout=>p(255)(44));
FA_ff_7959:FAff port map(x=>p(188)(44),y=>p(189)(44),Cin=>p(190)(44),clock=>clock,reset=>reset,s=>p(254)(44),cout=>p(255)(45));
FA_ff_7960:FAff port map(x=>p(188)(45),y=>p(189)(45),Cin=>p(190)(45),clock=>clock,reset=>reset,s=>p(254)(45),cout=>p(255)(46));
FA_ff_7961:FAff port map(x=>p(188)(46),y=>p(189)(46),Cin=>p(190)(46),clock=>clock,reset=>reset,s=>p(254)(46),cout=>p(255)(47));
FA_ff_7962:FAff port map(x=>p(188)(47),y=>p(189)(47),Cin=>p(190)(47),clock=>clock,reset=>reset,s=>p(254)(47),cout=>p(255)(48));
FA_ff_7963:FAff port map(x=>p(188)(48),y=>p(189)(48),Cin=>p(190)(48),clock=>clock,reset=>reset,s=>p(254)(48),cout=>p(255)(49));
FA_ff_7964:FAff port map(x=>p(188)(49),y=>p(189)(49),Cin=>p(190)(49),clock=>clock,reset=>reset,s=>p(254)(49),cout=>p(255)(50));
FA_ff_7965:FAff port map(x=>p(188)(50),y=>p(189)(50),Cin=>p(190)(50),clock=>clock,reset=>reset,s=>p(254)(50),cout=>p(255)(51));
FA_ff_7966:FAff port map(x=>p(188)(51),y=>p(189)(51),Cin=>p(190)(51),clock=>clock,reset=>reset,s=>p(254)(51),cout=>p(255)(52));
FA_ff_7967:FAff port map(x=>p(188)(52),y=>p(189)(52),Cin=>p(190)(52),clock=>clock,reset=>reset,s=>p(254)(52),cout=>p(255)(53));
FA_ff_7968:FAff port map(x=>p(188)(53),y=>p(189)(53),Cin=>p(190)(53),clock=>clock,reset=>reset,s=>p(254)(53),cout=>p(255)(54));
FA_ff_7969:FAff port map(x=>p(188)(54),y=>p(189)(54),Cin=>p(190)(54),clock=>clock,reset=>reset,s=>p(254)(54),cout=>p(255)(55));
FA_ff_7970:FAff port map(x=>p(188)(55),y=>p(189)(55),Cin=>p(190)(55),clock=>clock,reset=>reset,s=>p(254)(55),cout=>p(255)(56));
FA_ff_7971:FAff port map(x=>p(188)(56),y=>p(189)(56),Cin=>p(190)(56),clock=>clock,reset=>reset,s=>p(254)(56),cout=>p(255)(57));
FA_ff_7972:FAff port map(x=>p(188)(57),y=>p(189)(57),Cin=>p(190)(57),clock=>clock,reset=>reset,s=>p(254)(57),cout=>p(255)(58));
FA_ff_7973:FAff port map(x=>p(188)(58),y=>p(189)(58),Cin=>p(190)(58),clock=>clock,reset=>reset,s=>p(254)(58),cout=>p(255)(59));
FA_ff_7974:FAff port map(x=>p(188)(59),y=>p(189)(59),Cin=>p(190)(59),clock=>clock,reset=>reset,s=>p(254)(59),cout=>p(255)(60));
FA_ff_7975:FAff port map(x=>p(188)(60),y=>p(189)(60),Cin=>p(190)(60),clock=>clock,reset=>reset,s=>p(254)(60),cout=>p(255)(61));
FA_ff_7976:FAff port map(x=>p(188)(61),y=>p(189)(61),Cin=>p(190)(61),clock=>clock,reset=>reset,s=>p(254)(61),cout=>p(255)(62));
FA_ff_7977:FAff port map(x=>p(188)(62),y=>p(189)(62),Cin=>p(190)(62),clock=>clock,reset=>reset,s=>p(254)(62),cout=>p(255)(63));
FA_ff_7978:FAff port map(x=>p(188)(63),y=>p(189)(63),Cin=>p(190)(63),clock=>clock,reset=>reset,s=>p(254)(63),cout=>p(255)(64));
FA_ff_7979:FAff port map(x=>p(188)(64),y=>p(189)(64),Cin=>p(190)(64),clock=>clock,reset=>reset,s=>p(254)(64),cout=>p(255)(65));
FA_ff_7980:FAff port map(x=>p(188)(65),y=>p(189)(65),Cin=>p(190)(65),clock=>clock,reset=>reset,s=>p(254)(65),cout=>p(255)(66));
FA_ff_7981:FAff port map(x=>p(188)(66),y=>p(189)(66),Cin=>p(190)(66),clock=>clock,reset=>reset,s=>p(254)(66),cout=>p(255)(67));
FA_ff_7982:FAff port map(x=>p(188)(67),y=>p(189)(67),Cin=>p(190)(67),clock=>clock,reset=>reset,s=>p(254)(67),cout=>p(255)(68));
FA_ff_7983:FAff port map(x=>p(188)(68),y=>p(189)(68),Cin=>p(190)(68),clock=>clock,reset=>reset,s=>p(254)(68),cout=>p(255)(69));
FA_ff_7984:FAff port map(x=>p(188)(69),y=>p(189)(69),Cin=>p(190)(69),clock=>clock,reset=>reset,s=>p(254)(69),cout=>p(255)(70));
FA_ff_7985:FAff port map(x=>p(188)(70),y=>p(189)(70),Cin=>p(190)(70),clock=>clock,reset=>reset,s=>p(254)(70),cout=>p(255)(71));
FA_ff_7986:FAff port map(x=>p(188)(71),y=>p(189)(71),Cin=>p(190)(71),clock=>clock,reset=>reset,s=>p(254)(71),cout=>p(255)(72));
FA_ff_7987:FAff port map(x=>p(188)(72),y=>p(189)(72),Cin=>p(190)(72),clock=>clock,reset=>reset,s=>p(254)(72),cout=>p(255)(73));
FA_ff_7988:FAff port map(x=>p(188)(73),y=>p(189)(73),Cin=>p(190)(73),clock=>clock,reset=>reset,s=>p(254)(73),cout=>p(255)(74));
FA_ff_7989:FAff port map(x=>p(188)(74),y=>p(189)(74),Cin=>p(190)(74),clock=>clock,reset=>reset,s=>p(254)(74),cout=>p(255)(75));
FA_ff_7990:FAff port map(x=>p(188)(75),y=>p(189)(75),Cin=>p(190)(75),clock=>clock,reset=>reset,s=>p(254)(75),cout=>p(255)(76));
FA_ff_7991:FAff port map(x=>p(188)(76),y=>p(189)(76),Cin=>p(190)(76),clock=>clock,reset=>reset,s=>p(254)(76),cout=>p(255)(77));
FA_ff_7992:FAff port map(x=>p(188)(77),y=>p(189)(77),Cin=>p(190)(77),clock=>clock,reset=>reset,s=>p(254)(77),cout=>p(255)(78));
FA_ff_7993:FAff port map(x=>p(188)(78),y=>p(189)(78),Cin=>p(190)(78),clock=>clock,reset=>reset,s=>p(254)(78),cout=>p(255)(79));
FA_ff_7994:FAff port map(x=>p(188)(79),y=>p(189)(79),Cin=>p(190)(79),clock=>clock,reset=>reset,s=>p(254)(79),cout=>p(255)(80));
FA_ff_7995:FAff port map(x=>p(188)(80),y=>p(189)(80),Cin=>p(190)(80),clock=>clock,reset=>reset,s=>p(254)(80),cout=>p(255)(81));
FA_ff_7996:FAff port map(x=>p(188)(81),y=>p(189)(81),Cin=>p(190)(81),clock=>clock,reset=>reset,s=>p(254)(81),cout=>p(255)(82));
FA_ff_7997:FAff port map(x=>p(188)(82),y=>p(189)(82),Cin=>p(190)(82),clock=>clock,reset=>reset,s=>p(254)(82),cout=>p(255)(83));
FA_ff_7998:FAff port map(x=>p(188)(83),y=>p(189)(83),Cin=>p(190)(83),clock=>clock,reset=>reset,s=>p(254)(83),cout=>p(255)(84));
FA_ff_7999:FAff port map(x=>p(188)(84),y=>p(189)(84),Cin=>p(190)(84),clock=>clock,reset=>reset,s=>p(254)(84),cout=>p(255)(85));
FA_ff_8000:FAff port map(x=>p(188)(85),y=>p(189)(85),Cin=>p(190)(85),clock=>clock,reset=>reset,s=>p(254)(85),cout=>p(255)(86));
FA_ff_8001:FAff port map(x=>p(188)(86),y=>p(189)(86),Cin=>p(190)(86),clock=>clock,reset=>reset,s=>p(254)(86),cout=>p(255)(87));
FA_ff_8002:FAff port map(x=>p(188)(87),y=>p(189)(87),Cin=>p(190)(87),clock=>clock,reset=>reset,s=>p(254)(87),cout=>p(255)(88));
FA_ff_8003:FAff port map(x=>p(188)(88),y=>p(189)(88),Cin=>p(190)(88),clock=>clock,reset=>reset,s=>p(254)(88),cout=>p(255)(89));
FA_ff_8004:FAff port map(x=>p(188)(89),y=>p(189)(89),Cin=>p(190)(89),clock=>clock,reset=>reset,s=>p(254)(89),cout=>p(255)(90));
FA_ff_8005:FAff port map(x=>p(188)(90),y=>p(189)(90),Cin=>p(190)(90),clock=>clock,reset=>reset,s=>p(254)(90),cout=>p(255)(91));
FA_ff_8006:FAff port map(x=>p(188)(91),y=>p(189)(91),Cin=>p(190)(91),clock=>clock,reset=>reset,s=>p(254)(91),cout=>p(255)(92));
FA_ff_8007:FAff port map(x=>p(188)(92),y=>p(189)(92),Cin=>p(190)(92),clock=>clock,reset=>reset,s=>p(254)(92),cout=>p(255)(93));
FA_ff_8008:FAff port map(x=>p(188)(93),y=>p(189)(93),Cin=>p(190)(93),clock=>clock,reset=>reset,s=>p(254)(93),cout=>p(255)(94));
FA_ff_8009:FAff port map(x=>p(188)(94),y=>p(189)(94),Cin=>p(190)(94),clock=>clock,reset=>reset,s=>p(254)(94),cout=>p(255)(95));
FA_ff_8010:FAff port map(x=>p(188)(95),y=>p(189)(95),Cin=>p(190)(95),clock=>clock,reset=>reset,s=>p(254)(95),cout=>p(255)(96));
FA_ff_8011:FAff port map(x=>p(188)(96),y=>p(189)(96),Cin=>p(190)(96),clock=>clock,reset=>reset,s=>p(254)(96),cout=>p(255)(97));
FA_ff_8012:FAff port map(x=>p(188)(97),y=>p(189)(97),Cin=>p(190)(97),clock=>clock,reset=>reset,s=>p(254)(97),cout=>p(255)(98));
FA_ff_8013:FAff port map(x=>p(188)(98),y=>p(189)(98),Cin=>p(190)(98),clock=>clock,reset=>reset,s=>p(254)(98),cout=>p(255)(99));
FA_ff_8014:FAff port map(x=>p(188)(99),y=>p(189)(99),Cin=>p(190)(99),clock=>clock,reset=>reset,s=>p(254)(99),cout=>p(255)(100));
FA_ff_8015:FAff port map(x=>p(188)(100),y=>p(189)(100),Cin=>p(190)(100),clock=>clock,reset=>reset,s=>p(254)(100),cout=>p(255)(101));
FA_ff_8016:FAff port map(x=>p(188)(101),y=>p(189)(101),Cin=>p(190)(101),clock=>clock,reset=>reset,s=>p(254)(101),cout=>p(255)(102));
FA_ff_8017:FAff port map(x=>p(188)(102),y=>p(189)(102),Cin=>p(190)(102),clock=>clock,reset=>reset,s=>p(254)(102),cout=>p(255)(103));
FA_ff_8018:FAff port map(x=>p(188)(103),y=>p(189)(103),Cin=>p(190)(103),clock=>clock,reset=>reset,s=>p(254)(103),cout=>p(255)(104));
FA_ff_8019:FAff port map(x=>p(188)(104),y=>p(189)(104),Cin=>p(190)(104),clock=>clock,reset=>reset,s=>p(254)(104),cout=>p(255)(105));
FA_ff_8020:FAff port map(x=>p(188)(105),y=>p(189)(105),Cin=>p(190)(105),clock=>clock,reset=>reset,s=>p(254)(105),cout=>p(255)(106));
FA_ff_8021:FAff port map(x=>p(188)(106),y=>p(189)(106),Cin=>p(190)(106),clock=>clock,reset=>reset,s=>p(254)(106),cout=>p(255)(107));
FA_ff_8022:FAff port map(x=>p(188)(107),y=>p(189)(107),Cin=>p(190)(107),clock=>clock,reset=>reset,s=>p(254)(107),cout=>p(255)(108));
FA_ff_8023:FAff port map(x=>p(188)(108),y=>p(189)(108),Cin=>p(190)(108),clock=>clock,reset=>reset,s=>p(254)(108),cout=>p(255)(109));
FA_ff_8024:FAff port map(x=>p(188)(109),y=>p(189)(109),Cin=>p(190)(109),clock=>clock,reset=>reset,s=>p(254)(109),cout=>p(255)(110));
FA_ff_8025:FAff port map(x=>p(188)(110),y=>p(189)(110),Cin=>p(190)(110),clock=>clock,reset=>reset,s=>p(254)(110),cout=>p(255)(111));
FA_ff_8026:FAff port map(x=>p(188)(111),y=>p(189)(111),Cin=>p(190)(111),clock=>clock,reset=>reset,s=>p(254)(111),cout=>p(255)(112));
FA_ff_8027:FAff port map(x=>p(188)(112),y=>p(189)(112),Cin=>p(190)(112),clock=>clock,reset=>reset,s=>p(254)(112),cout=>p(255)(113));
FA_ff_8028:FAff port map(x=>p(188)(113),y=>p(189)(113),Cin=>p(190)(113),clock=>clock,reset=>reset,s=>p(254)(113),cout=>p(255)(114));
FA_ff_8029:FAff port map(x=>p(188)(114),y=>p(189)(114),Cin=>p(190)(114),clock=>clock,reset=>reset,s=>p(254)(114),cout=>p(255)(115));
FA_ff_8030:FAff port map(x=>p(188)(115),y=>p(189)(115),Cin=>p(190)(115),clock=>clock,reset=>reset,s=>p(254)(115),cout=>p(255)(116));
FA_ff_8031:FAff port map(x=>p(188)(116),y=>p(189)(116),Cin=>p(190)(116),clock=>clock,reset=>reset,s=>p(254)(116),cout=>p(255)(117));
FA_ff_8032:FAff port map(x=>p(188)(117),y=>p(189)(117),Cin=>p(190)(117),clock=>clock,reset=>reset,s=>p(254)(117),cout=>p(255)(118));
FA_ff_8033:FAff port map(x=>p(188)(118),y=>p(189)(118),Cin=>p(190)(118),clock=>clock,reset=>reset,s=>p(254)(118),cout=>p(255)(119));
FA_ff_8034:FAff port map(x=>p(188)(119),y=>p(189)(119),Cin=>p(190)(119),clock=>clock,reset=>reset,s=>p(254)(119),cout=>p(255)(120));
FA_ff_8035:FAff port map(x=>p(188)(120),y=>p(189)(120),Cin=>p(190)(120),clock=>clock,reset=>reset,s=>p(254)(120),cout=>p(255)(121));
FA_ff_8036:FAff port map(x=>p(188)(121),y=>p(189)(121),Cin=>p(190)(121),clock=>clock,reset=>reset,s=>p(254)(121),cout=>p(255)(122));
FA_ff_8037:FAff port map(x=>p(188)(122),y=>p(189)(122),Cin=>p(190)(122),clock=>clock,reset=>reset,s=>p(254)(122),cout=>p(255)(123));
FA_ff_8038:FAff port map(x=>p(188)(123),y=>p(189)(123),Cin=>p(190)(123),clock=>clock,reset=>reset,s=>p(254)(123),cout=>p(255)(124));
FA_ff_8039:FAff port map(x=>p(188)(124),y=>p(189)(124),Cin=>p(190)(124),clock=>clock,reset=>reset,s=>p(254)(124),cout=>p(255)(125));
FA_ff_8040:FAff port map(x=>p(188)(125),y=>p(189)(125),Cin=>p(190)(125),clock=>clock,reset=>reset,s=>p(254)(125),cout=>p(255)(126));
FA_ff_8041:FAff port map(x=>p(188)(126),y=>p(189)(126),Cin=>p(190)(126),clock=>clock,reset=>reset,s=>p(254)(126),cout=>p(255)(127));
FA_ff_8042:FAff port map(x=>p(188)(127),y=>p(189)(127),Cin=>p(190)(127),clock=>clock,reset=>reset,s=>p(254)(127),cout=>p(255)(128));
p(254)(128)<=p(189)(128);
p(256)(0)<=p(192)(0);
FA_ff_8043:FAff port map(x=>p(191)(1),y=>p(192)(1),Cin=>p(193)(1),clock=>clock,reset=>reset,s=>p(256)(1),cout=>p(257)(2));
FA_ff_8044:FAff port map(x=>p(191)(2),y=>p(192)(2),Cin=>p(193)(2),clock=>clock,reset=>reset,s=>p(256)(2),cout=>p(257)(3));
FA_ff_8045:FAff port map(x=>p(191)(3),y=>p(192)(3),Cin=>p(193)(3),clock=>clock,reset=>reset,s=>p(256)(3),cout=>p(257)(4));
FA_ff_8046:FAff port map(x=>p(191)(4),y=>p(192)(4),Cin=>p(193)(4),clock=>clock,reset=>reset,s=>p(256)(4),cout=>p(257)(5));
FA_ff_8047:FAff port map(x=>p(191)(5),y=>p(192)(5),Cin=>p(193)(5),clock=>clock,reset=>reset,s=>p(256)(5),cout=>p(257)(6));
FA_ff_8048:FAff port map(x=>p(191)(6),y=>p(192)(6),Cin=>p(193)(6),clock=>clock,reset=>reset,s=>p(256)(6),cout=>p(257)(7));
FA_ff_8049:FAff port map(x=>p(191)(7),y=>p(192)(7),Cin=>p(193)(7),clock=>clock,reset=>reset,s=>p(256)(7),cout=>p(257)(8));
FA_ff_8050:FAff port map(x=>p(191)(8),y=>p(192)(8),Cin=>p(193)(8),clock=>clock,reset=>reset,s=>p(256)(8),cout=>p(257)(9));
FA_ff_8051:FAff port map(x=>p(191)(9),y=>p(192)(9),Cin=>p(193)(9),clock=>clock,reset=>reset,s=>p(256)(9),cout=>p(257)(10));
FA_ff_8052:FAff port map(x=>p(191)(10),y=>p(192)(10),Cin=>p(193)(10),clock=>clock,reset=>reset,s=>p(256)(10),cout=>p(257)(11));
FA_ff_8053:FAff port map(x=>p(191)(11),y=>p(192)(11),Cin=>p(193)(11),clock=>clock,reset=>reset,s=>p(256)(11),cout=>p(257)(12));
FA_ff_8054:FAff port map(x=>p(191)(12),y=>p(192)(12),Cin=>p(193)(12),clock=>clock,reset=>reset,s=>p(256)(12),cout=>p(257)(13));
FA_ff_8055:FAff port map(x=>p(191)(13),y=>p(192)(13),Cin=>p(193)(13),clock=>clock,reset=>reset,s=>p(256)(13),cout=>p(257)(14));
FA_ff_8056:FAff port map(x=>p(191)(14),y=>p(192)(14),Cin=>p(193)(14),clock=>clock,reset=>reset,s=>p(256)(14),cout=>p(257)(15));
FA_ff_8057:FAff port map(x=>p(191)(15),y=>p(192)(15),Cin=>p(193)(15),clock=>clock,reset=>reset,s=>p(256)(15),cout=>p(257)(16));
FA_ff_8058:FAff port map(x=>p(191)(16),y=>p(192)(16),Cin=>p(193)(16),clock=>clock,reset=>reset,s=>p(256)(16),cout=>p(257)(17));
FA_ff_8059:FAff port map(x=>p(191)(17),y=>p(192)(17),Cin=>p(193)(17),clock=>clock,reset=>reset,s=>p(256)(17),cout=>p(257)(18));
FA_ff_8060:FAff port map(x=>p(191)(18),y=>p(192)(18),Cin=>p(193)(18),clock=>clock,reset=>reset,s=>p(256)(18),cout=>p(257)(19));
FA_ff_8061:FAff port map(x=>p(191)(19),y=>p(192)(19),Cin=>p(193)(19),clock=>clock,reset=>reset,s=>p(256)(19),cout=>p(257)(20));
FA_ff_8062:FAff port map(x=>p(191)(20),y=>p(192)(20),Cin=>p(193)(20),clock=>clock,reset=>reset,s=>p(256)(20),cout=>p(257)(21));
FA_ff_8063:FAff port map(x=>p(191)(21),y=>p(192)(21),Cin=>p(193)(21),clock=>clock,reset=>reset,s=>p(256)(21),cout=>p(257)(22));
FA_ff_8064:FAff port map(x=>p(191)(22),y=>p(192)(22),Cin=>p(193)(22),clock=>clock,reset=>reset,s=>p(256)(22),cout=>p(257)(23));
FA_ff_8065:FAff port map(x=>p(191)(23),y=>p(192)(23),Cin=>p(193)(23),clock=>clock,reset=>reset,s=>p(256)(23),cout=>p(257)(24));
FA_ff_8066:FAff port map(x=>p(191)(24),y=>p(192)(24),Cin=>p(193)(24),clock=>clock,reset=>reset,s=>p(256)(24),cout=>p(257)(25));
FA_ff_8067:FAff port map(x=>p(191)(25),y=>p(192)(25),Cin=>p(193)(25),clock=>clock,reset=>reset,s=>p(256)(25),cout=>p(257)(26));
FA_ff_8068:FAff port map(x=>p(191)(26),y=>p(192)(26),Cin=>p(193)(26),clock=>clock,reset=>reset,s=>p(256)(26),cout=>p(257)(27));
FA_ff_8069:FAff port map(x=>p(191)(27),y=>p(192)(27),Cin=>p(193)(27),clock=>clock,reset=>reset,s=>p(256)(27),cout=>p(257)(28));
FA_ff_8070:FAff port map(x=>p(191)(28),y=>p(192)(28),Cin=>p(193)(28),clock=>clock,reset=>reset,s=>p(256)(28),cout=>p(257)(29));
FA_ff_8071:FAff port map(x=>p(191)(29),y=>p(192)(29),Cin=>p(193)(29),clock=>clock,reset=>reset,s=>p(256)(29),cout=>p(257)(30));
FA_ff_8072:FAff port map(x=>p(191)(30),y=>p(192)(30),Cin=>p(193)(30),clock=>clock,reset=>reset,s=>p(256)(30),cout=>p(257)(31));
FA_ff_8073:FAff port map(x=>p(191)(31),y=>p(192)(31),Cin=>p(193)(31),clock=>clock,reset=>reset,s=>p(256)(31),cout=>p(257)(32));
FA_ff_8074:FAff port map(x=>p(191)(32),y=>p(192)(32),Cin=>p(193)(32),clock=>clock,reset=>reset,s=>p(256)(32),cout=>p(257)(33));
FA_ff_8075:FAff port map(x=>p(191)(33),y=>p(192)(33),Cin=>p(193)(33),clock=>clock,reset=>reset,s=>p(256)(33),cout=>p(257)(34));
FA_ff_8076:FAff port map(x=>p(191)(34),y=>p(192)(34),Cin=>p(193)(34),clock=>clock,reset=>reset,s=>p(256)(34),cout=>p(257)(35));
FA_ff_8077:FAff port map(x=>p(191)(35),y=>p(192)(35),Cin=>p(193)(35),clock=>clock,reset=>reset,s=>p(256)(35),cout=>p(257)(36));
FA_ff_8078:FAff port map(x=>p(191)(36),y=>p(192)(36),Cin=>p(193)(36),clock=>clock,reset=>reset,s=>p(256)(36),cout=>p(257)(37));
FA_ff_8079:FAff port map(x=>p(191)(37),y=>p(192)(37),Cin=>p(193)(37),clock=>clock,reset=>reset,s=>p(256)(37),cout=>p(257)(38));
FA_ff_8080:FAff port map(x=>p(191)(38),y=>p(192)(38),Cin=>p(193)(38),clock=>clock,reset=>reset,s=>p(256)(38),cout=>p(257)(39));
FA_ff_8081:FAff port map(x=>p(191)(39),y=>p(192)(39),Cin=>p(193)(39),clock=>clock,reset=>reset,s=>p(256)(39),cout=>p(257)(40));
FA_ff_8082:FAff port map(x=>p(191)(40),y=>p(192)(40),Cin=>p(193)(40),clock=>clock,reset=>reset,s=>p(256)(40),cout=>p(257)(41));
FA_ff_8083:FAff port map(x=>p(191)(41),y=>p(192)(41),Cin=>p(193)(41),clock=>clock,reset=>reset,s=>p(256)(41),cout=>p(257)(42));
FA_ff_8084:FAff port map(x=>p(191)(42),y=>p(192)(42),Cin=>p(193)(42),clock=>clock,reset=>reset,s=>p(256)(42),cout=>p(257)(43));
FA_ff_8085:FAff port map(x=>p(191)(43),y=>p(192)(43),Cin=>p(193)(43),clock=>clock,reset=>reset,s=>p(256)(43),cout=>p(257)(44));
FA_ff_8086:FAff port map(x=>p(191)(44),y=>p(192)(44),Cin=>p(193)(44),clock=>clock,reset=>reset,s=>p(256)(44),cout=>p(257)(45));
FA_ff_8087:FAff port map(x=>p(191)(45),y=>p(192)(45),Cin=>p(193)(45),clock=>clock,reset=>reset,s=>p(256)(45),cout=>p(257)(46));
FA_ff_8088:FAff port map(x=>p(191)(46),y=>p(192)(46),Cin=>p(193)(46),clock=>clock,reset=>reset,s=>p(256)(46),cout=>p(257)(47));
FA_ff_8089:FAff port map(x=>p(191)(47),y=>p(192)(47),Cin=>p(193)(47),clock=>clock,reset=>reset,s=>p(256)(47),cout=>p(257)(48));
FA_ff_8090:FAff port map(x=>p(191)(48),y=>p(192)(48),Cin=>p(193)(48),clock=>clock,reset=>reset,s=>p(256)(48),cout=>p(257)(49));
FA_ff_8091:FAff port map(x=>p(191)(49),y=>p(192)(49),Cin=>p(193)(49),clock=>clock,reset=>reset,s=>p(256)(49),cout=>p(257)(50));
FA_ff_8092:FAff port map(x=>p(191)(50),y=>p(192)(50),Cin=>p(193)(50),clock=>clock,reset=>reset,s=>p(256)(50),cout=>p(257)(51));
FA_ff_8093:FAff port map(x=>p(191)(51),y=>p(192)(51),Cin=>p(193)(51),clock=>clock,reset=>reset,s=>p(256)(51),cout=>p(257)(52));
FA_ff_8094:FAff port map(x=>p(191)(52),y=>p(192)(52),Cin=>p(193)(52),clock=>clock,reset=>reset,s=>p(256)(52),cout=>p(257)(53));
FA_ff_8095:FAff port map(x=>p(191)(53),y=>p(192)(53),Cin=>p(193)(53),clock=>clock,reset=>reset,s=>p(256)(53),cout=>p(257)(54));
FA_ff_8096:FAff port map(x=>p(191)(54),y=>p(192)(54),Cin=>p(193)(54),clock=>clock,reset=>reset,s=>p(256)(54),cout=>p(257)(55));
FA_ff_8097:FAff port map(x=>p(191)(55),y=>p(192)(55),Cin=>p(193)(55),clock=>clock,reset=>reset,s=>p(256)(55),cout=>p(257)(56));
FA_ff_8098:FAff port map(x=>p(191)(56),y=>p(192)(56),Cin=>p(193)(56),clock=>clock,reset=>reset,s=>p(256)(56),cout=>p(257)(57));
FA_ff_8099:FAff port map(x=>p(191)(57),y=>p(192)(57),Cin=>p(193)(57),clock=>clock,reset=>reset,s=>p(256)(57),cout=>p(257)(58));
FA_ff_8100:FAff port map(x=>p(191)(58),y=>p(192)(58),Cin=>p(193)(58),clock=>clock,reset=>reset,s=>p(256)(58),cout=>p(257)(59));
FA_ff_8101:FAff port map(x=>p(191)(59),y=>p(192)(59),Cin=>p(193)(59),clock=>clock,reset=>reset,s=>p(256)(59),cout=>p(257)(60));
FA_ff_8102:FAff port map(x=>p(191)(60),y=>p(192)(60),Cin=>p(193)(60),clock=>clock,reset=>reset,s=>p(256)(60),cout=>p(257)(61));
FA_ff_8103:FAff port map(x=>p(191)(61),y=>p(192)(61),Cin=>p(193)(61),clock=>clock,reset=>reset,s=>p(256)(61),cout=>p(257)(62));
FA_ff_8104:FAff port map(x=>p(191)(62),y=>p(192)(62),Cin=>p(193)(62),clock=>clock,reset=>reset,s=>p(256)(62),cout=>p(257)(63));
FA_ff_8105:FAff port map(x=>p(191)(63),y=>p(192)(63),Cin=>p(193)(63),clock=>clock,reset=>reset,s=>p(256)(63),cout=>p(257)(64));
FA_ff_8106:FAff port map(x=>p(191)(64),y=>p(192)(64),Cin=>p(193)(64),clock=>clock,reset=>reset,s=>p(256)(64),cout=>p(257)(65));
FA_ff_8107:FAff port map(x=>p(191)(65),y=>p(192)(65),Cin=>p(193)(65),clock=>clock,reset=>reset,s=>p(256)(65),cout=>p(257)(66));
FA_ff_8108:FAff port map(x=>p(191)(66),y=>p(192)(66),Cin=>p(193)(66),clock=>clock,reset=>reset,s=>p(256)(66),cout=>p(257)(67));
FA_ff_8109:FAff port map(x=>p(191)(67),y=>p(192)(67),Cin=>p(193)(67),clock=>clock,reset=>reset,s=>p(256)(67),cout=>p(257)(68));
FA_ff_8110:FAff port map(x=>p(191)(68),y=>p(192)(68),Cin=>p(193)(68),clock=>clock,reset=>reset,s=>p(256)(68),cout=>p(257)(69));
FA_ff_8111:FAff port map(x=>p(191)(69),y=>p(192)(69),Cin=>p(193)(69),clock=>clock,reset=>reset,s=>p(256)(69),cout=>p(257)(70));
FA_ff_8112:FAff port map(x=>p(191)(70),y=>p(192)(70),Cin=>p(193)(70),clock=>clock,reset=>reset,s=>p(256)(70),cout=>p(257)(71));
FA_ff_8113:FAff port map(x=>p(191)(71),y=>p(192)(71),Cin=>p(193)(71),clock=>clock,reset=>reset,s=>p(256)(71),cout=>p(257)(72));
FA_ff_8114:FAff port map(x=>p(191)(72),y=>p(192)(72),Cin=>p(193)(72),clock=>clock,reset=>reset,s=>p(256)(72),cout=>p(257)(73));
FA_ff_8115:FAff port map(x=>p(191)(73),y=>p(192)(73),Cin=>p(193)(73),clock=>clock,reset=>reset,s=>p(256)(73),cout=>p(257)(74));
FA_ff_8116:FAff port map(x=>p(191)(74),y=>p(192)(74),Cin=>p(193)(74),clock=>clock,reset=>reset,s=>p(256)(74),cout=>p(257)(75));
FA_ff_8117:FAff port map(x=>p(191)(75),y=>p(192)(75),Cin=>p(193)(75),clock=>clock,reset=>reset,s=>p(256)(75),cout=>p(257)(76));
FA_ff_8118:FAff port map(x=>p(191)(76),y=>p(192)(76),Cin=>p(193)(76),clock=>clock,reset=>reset,s=>p(256)(76),cout=>p(257)(77));
FA_ff_8119:FAff port map(x=>p(191)(77),y=>p(192)(77),Cin=>p(193)(77),clock=>clock,reset=>reset,s=>p(256)(77),cout=>p(257)(78));
FA_ff_8120:FAff port map(x=>p(191)(78),y=>p(192)(78),Cin=>p(193)(78),clock=>clock,reset=>reset,s=>p(256)(78),cout=>p(257)(79));
FA_ff_8121:FAff port map(x=>p(191)(79),y=>p(192)(79),Cin=>p(193)(79),clock=>clock,reset=>reset,s=>p(256)(79),cout=>p(257)(80));
FA_ff_8122:FAff port map(x=>p(191)(80),y=>p(192)(80),Cin=>p(193)(80),clock=>clock,reset=>reset,s=>p(256)(80),cout=>p(257)(81));
FA_ff_8123:FAff port map(x=>p(191)(81),y=>p(192)(81),Cin=>p(193)(81),clock=>clock,reset=>reset,s=>p(256)(81),cout=>p(257)(82));
FA_ff_8124:FAff port map(x=>p(191)(82),y=>p(192)(82),Cin=>p(193)(82),clock=>clock,reset=>reset,s=>p(256)(82),cout=>p(257)(83));
FA_ff_8125:FAff port map(x=>p(191)(83),y=>p(192)(83),Cin=>p(193)(83),clock=>clock,reset=>reset,s=>p(256)(83),cout=>p(257)(84));
FA_ff_8126:FAff port map(x=>p(191)(84),y=>p(192)(84),Cin=>p(193)(84),clock=>clock,reset=>reset,s=>p(256)(84),cout=>p(257)(85));
FA_ff_8127:FAff port map(x=>p(191)(85),y=>p(192)(85),Cin=>p(193)(85),clock=>clock,reset=>reset,s=>p(256)(85),cout=>p(257)(86));
FA_ff_8128:FAff port map(x=>p(191)(86),y=>p(192)(86),Cin=>p(193)(86),clock=>clock,reset=>reset,s=>p(256)(86),cout=>p(257)(87));
FA_ff_8129:FAff port map(x=>p(191)(87),y=>p(192)(87),Cin=>p(193)(87),clock=>clock,reset=>reset,s=>p(256)(87),cout=>p(257)(88));
FA_ff_8130:FAff port map(x=>p(191)(88),y=>p(192)(88),Cin=>p(193)(88),clock=>clock,reset=>reset,s=>p(256)(88),cout=>p(257)(89));
FA_ff_8131:FAff port map(x=>p(191)(89),y=>p(192)(89),Cin=>p(193)(89),clock=>clock,reset=>reset,s=>p(256)(89),cout=>p(257)(90));
FA_ff_8132:FAff port map(x=>p(191)(90),y=>p(192)(90),Cin=>p(193)(90),clock=>clock,reset=>reset,s=>p(256)(90),cout=>p(257)(91));
FA_ff_8133:FAff port map(x=>p(191)(91),y=>p(192)(91),Cin=>p(193)(91),clock=>clock,reset=>reset,s=>p(256)(91),cout=>p(257)(92));
FA_ff_8134:FAff port map(x=>p(191)(92),y=>p(192)(92),Cin=>p(193)(92),clock=>clock,reset=>reset,s=>p(256)(92),cout=>p(257)(93));
FA_ff_8135:FAff port map(x=>p(191)(93),y=>p(192)(93),Cin=>p(193)(93),clock=>clock,reset=>reset,s=>p(256)(93),cout=>p(257)(94));
FA_ff_8136:FAff port map(x=>p(191)(94),y=>p(192)(94),Cin=>p(193)(94),clock=>clock,reset=>reset,s=>p(256)(94),cout=>p(257)(95));
FA_ff_8137:FAff port map(x=>p(191)(95),y=>p(192)(95),Cin=>p(193)(95),clock=>clock,reset=>reset,s=>p(256)(95),cout=>p(257)(96));
FA_ff_8138:FAff port map(x=>p(191)(96),y=>p(192)(96),Cin=>p(193)(96),clock=>clock,reset=>reset,s=>p(256)(96),cout=>p(257)(97));
FA_ff_8139:FAff port map(x=>p(191)(97),y=>p(192)(97),Cin=>p(193)(97),clock=>clock,reset=>reset,s=>p(256)(97),cout=>p(257)(98));
FA_ff_8140:FAff port map(x=>p(191)(98),y=>p(192)(98),Cin=>p(193)(98),clock=>clock,reset=>reset,s=>p(256)(98),cout=>p(257)(99));
FA_ff_8141:FAff port map(x=>p(191)(99),y=>p(192)(99),Cin=>p(193)(99),clock=>clock,reset=>reset,s=>p(256)(99),cout=>p(257)(100));
FA_ff_8142:FAff port map(x=>p(191)(100),y=>p(192)(100),Cin=>p(193)(100),clock=>clock,reset=>reset,s=>p(256)(100),cout=>p(257)(101));
FA_ff_8143:FAff port map(x=>p(191)(101),y=>p(192)(101),Cin=>p(193)(101),clock=>clock,reset=>reset,s=>p(256)(101),cout=>p(257)(102));
FA_ff_8144:FAff port map(x=>p(191)(102),y=>p(192)(102),Cin=>p(193)(102),clock=>clock,reset=>reset,s=>p(256)(102),cout=>p(257)(103));
FA_ff_8145:FAff port map(x=>p(191)(103),y=>p(192)(103),Cin=>p(193)(103),clock=>clock,reset=>reset,s=>p(256)(103),cout=>p(257)(104));
FA_ff_8146:FAff port map(x=>p(191)(104),y=>p(192)(104),Cin=>p(193)(104),clock=>clock,reset=>reset,s=>p(256)(104),cout=>p(257)(105));
FA_ff_8147:FAff port map(x=>p(191)(105),y=>p(192)(105),Cin=>p(193)(105),clock=>clock,reset=>reset,s=>p(256)(105),cout=>p(257)(106));
FA_ff_8148:FAff port map(x=>p(191)(106),y=>p(192)(106),Cin=>p(193)(106),clock=>clock,reset=>reset,s=>p(256)(106),cout=>p(257)(107));
FA_ff_8149:FAff port map(x=>p(191)(107),y=>p(192)(107),Cin=>p(193)(107),clock=>clock,reset=>reset,s=>p(256)(107),cout=>p(257)(108));
FA_ff_8150:FAff port map(x=>p(191)(108),y=>p(192)(108),Cin=>p(193)(108),clock=>clock,reset=>reset,s=>p(256)(108),cout=>p(257)(109));
FA_ff_8151:FAff port map(x=>p(191)(109),y=>p(192)(109),Cin=>p(193)(109),clock=>clock,reset=>reset,s=>p(256)(109),cout=>p(257)(110));
FA_ff_8152:FAff port map(x=>p(191)(110),y=>p(192)(110),Cin=>p(193)(110),clock=>clock,reset=>reset,s=>p(256)(110),cout=>p(257)(111));
FA_ff_8153:FAff port map(x=>p(191)(111),y=>p(192)(111),Cin=>p(193)(111),clock=>clock,reset=>reset,s=>p(256)(111),cout=>p(257)(112));
FA_ff_8154:FAff port map(x=>p(191)(112),y=>p(192)(112),Cin=>p(193)(112),clock=>clock,reset=>reset,s=>p(256)(112),cout=>p(257)(113));
FA_ff_8155:FAff port map(x=>p(191)(113),y=>p(192)(113),Cin=>p(193)(113),clock=>clock,reset=>reset,s=>p(256)(113),cout=>p(257)(114));
FA_ff_8156:FAff port map(x=>p(191)(114),y=>p(192)(114),Cin=>p(193)(114),clock=>clock,reset=>reset,s=>p(256)(114),cout=>p(257)(115));
FA_ff_8157:FAff port map(x=>p(191)(115),y=>p(192)(115),Cin=>p(193)(115),clock=>clock,reset=>reset,s=>p(256)(115),cout=>p(257)(116));
FA_ff_8158:FAff port map(x=>p(191)(116),y=>p(192)(116),Cin=>p(193)(116),clock=>clock,reset=>reset,s=>p(256)(116),cout=>p(257)(117));
FA_ff_8159:FAff port map(x=>p(191)(117),y=>p(192)(117),Cin=>p(193)(117),clock=>clock,reset=>reset,s=>p(256)(117),cout=>p(257)(118));
FA_ff_8160:FAff port map(x=>p(191)(118),y=>p(192)(118),Cin=>p(193)(118),clock=>clock,reset=>reset,s=>p(256)(118),cout=>p(257)(119));
FA_ff_8161:FAff port map(x=>p(191)(119),y=>p(192)(119),Cin=>p(193)(119),clock=>clock,reset=>reset,s=>p(256)(119),cout=>p(257)(120));
FA_ff_8162:FAff port map(x=>p(191)(120),y=>p(192)(120),Cin=>p(193)(120),clock=>clock,reset=>reset,s=>p(256)(120),cout=>p(257)(121));
FA_ff_8163:FAff port map(x=>p(191)(121),y=>p(192)(121),Cin=>p(193)(121),clock=>clock,reset=>reset,s=>p(256)(121),cout=>p(257)(122));
FA_ff_8164:FAff port map(x=>p(191)(122),y=>p(192)(122),Cin=>p(193)(122),clock=>clock,reset=>reset,s=>p(256)(122),cout=>p(257)(123));
FA_ff_8165:FAff port map(x=>p(191)(123),y=>p(192)(123),Cin=>p(193)(123),clock=>clock,reset=>reset,s=>p(256)(123),cout=>p(257)(124));
FA_ff_8166:FAff port map(x=>p(191)(124),y=>p(192)(124),Cin=>p(193)(124),clock=>clock,reset=>reset,s=>p(256)(124),cout=>p(257)(125));
FA_ff_8167:FAff port map(x=>p(191)(125),y=>p(192)(125),Cin=>p(193)(125),clock=>clock,reset=>reset,s=>p(256)(125),cout=>p(257)(126));
FA_ff_8168:FAff port map(x=>p(191)(126),y=>p(192)(126),Cin=>p(193)(126),clock=>clock,reset=>reset,s=>p(256)(126),cout=>p(257)(127));
FA_ff_8169:FAff port map(x=>p(191)(127),y=>p(192)(127),Cin=>p(193)(127),clock=>clock,reset=>reset,s=>p(256)(127),cout=>p(257)(128));
HA_ff_21:HAff port map(x=>p(191)(128),y=>p(193)(128),clock=>clock,reset=>reset,s=>p(256)(128),c=>p(257)(129));
HA_ff_22:HAff port map(x=>p(194)(0),y=>p(196)(0),clock=>clock,reset=>reset,s=>p(258)(0),c=>p(259)(1));
FA_ff_8170:FAff port map(x=>p(194)(1),y=>p(195)(1),Cin=>p(196)(1),clock=>clock,reset=>reset,s=>p(258)(1),cout=>p(259)(2));
FA_ff_8171:FAff port map(x=>p(194)(2),y=>p(195)(2),Cin=>p(196)(2),clock=>clock,reset=>reset,s=>p(258)(2),cout=>p(259)(3));
FA_ff_8172:FAff port map(x=>p(194)(3),y=>p(195)(3),Cin=>p(196)(3),clock=>clock,reset=>reset,s=>p(258)(3),cout=>p(259)(4));
FA_ff_8173:FAff port map(x=>p(194)(4),y=>p(195)(4),Cin=>p(196)(4),clock=>clock,reset=>reset,s=>p(258)(4),cout=>p(259)(5));
FA_ff_8174:FAff port map(x=>p(194)(5),y=>p(195)(5),Cin=>p(196)(5),clock=>clock,reset=>reset,s=>p(258)(5),cout=>p(259)(6));
FA_ff_8175:FAff port map(x=>p(194)(6),y=>p(195)(6),Cin=>p(196)(6),clock=>clock,reset=>reset,s=>p(258)(6),cout=>p(259)(7));
FA_ff_8176:FAff port map(x=>p(194)(7),y=>p(195)(7),Cin=>p(196)(7),clock=>clock,reset=>reset,s=>p(258)(7),cout=>p(259)(8));
FA_ff_8177:FAff port map(x=>p(194)(8),y=>p(195)(8),Cin=>p(196)(8),clock=>clock,reset=>reset,s=>p(258)(8),cout=>p(259)(9));
FA_ff_8178:FAff port map(x=>p(194)(9),y=>p(195)(9),Cin=>p(196)(9),clock=>clock,reset=>reset,s=>p(258)(9),cout=>p(259)(10));
FA_ff_8179:FAff port map(x=>p(194)(10),y=>p(195)(10),Cin=>p(196)(10),clock=>clock,reset=>reset,s=>p(258)(10),cout=>p(259)(11));
FA_ff_8180:FAff port map(x=>p(194)(11),y=>p(195)(11),Cin=>p(196)(11),clock=>clock,reset=>reset,s=>p(258)(11),cout=>p(259)(12));
FA_ff_8181:FAff port map(x=>p(194)(12),y=>p(195)(12),Cin=>p(196)(12),clock=>clock,reset=>reset,s=>p(258)(12),cout=>p(259)(13));
FA_ff_8182:FAff port map(x=>p(194)(13),y=>p(195)(13),Cin=>p(196)(13),clock=>clock,reset=>reset,s=>p(258)(13),cout=>p(259)(14));
FA_ff_8183:FAff port map(x=>p(194)(14),y=>p(195)(14),Cin=>p(196)(14),clock=>clock,reset=>reset,s=>p(258)(14),cout=>p(259)(15));
FA_ff_8184:FAff port map(x=>p(194)(15),y=>p(195)(15),Cin=>p(196)(15),clock=>clock,reset=>reset,s=>p(258)(15),cout=>p(259)(16));
FA_ff_8185:FAff port map(x=>p(194)(16),y=>p(195)(16),Cin=>p(196)(16),clock=>clock,reset=>reset,s=>p(258)(16),cout=>p(259)(17));
FA_ff_8186:FAff port map(x=>p(194)(17),y=>p(195)(17),Cin=>p(196)(17),clock=>clock,reset=>reset,s=>p(258)(17),cout=>p(259)(18));
FA_ff_8187:FAff port map(x=>p(194)(18),y=>p(195)(18),Cin=>p(196)(18),clock=>clock,reset=>reset,s=>p(258)(18),cout=>p(259)(19));
FA_ff_8188:FAff port map(x=>p(194)(19),y=>p(195)(19),Cin=>p(196)(19),clock=>clock,reset=>reset,s=>p(258)(19),cout=>p(259)(20));
FA_ff_8189:FAff port map(x=>p(194)(20),y=>p(195)(20),Cin=>p(196)(20),clock=>clock,reset=>reset,s=>p(258)(20),cout=>p(259)(21));
FA_ff_8190:FAff port map(x=>p(194)(21),y=>p(195)(21),Cin=>p(196)(21),clock=>clock,reset=>reset,s=>p(258)(21),cout=>p(259)(22));
FA_ff_8191:FAff port map(x=>p(194)(22),y=>p(195)(22),Cin=>p(196)(22),clock=>clock,reset=>reset,s=>p(258)(22),cout=>p(259)(23));
FA_ff_8192:FAff port map(x=>p(194)(23),y=>p(195)(23),Cin=>p(196)(23),clock=>clock,reset=>reset,s=>p(258)(23),cout=>p(259)(24));
FA_ff_8193:FAff port map(x=>p(194)(24),y=>p(195)(24),Cin=>p(196)(24),clock=>clock,reset=>reset,s=>p(258)(24),cout=>p(259)(25));
FA_ff_8194:FAff port map(x=>p(194)(25),y=>p(195)(25),Cin=>p(196)(25),clock=>clock,reset=>reset,s=>p(258)(25),cout=>p(259)(26));
FA_ff_8195:FAff port map(x=>p(194)(26),y=>p(195)(26),Cin=>p(196)(26),clock=>clock,reset=>reset,s=>p(258)(26),cout=>p(259)(27));
FA_ff_8196:FAff port map(x=>p(194)(27),y=>p(195)(27),Cin=>p(196)(27),clock=>clock,reset=>reset,s=>p(258)(27),cout=>p(259)(28));
FA_ff_8197:FAff port map(x=>p(194)(28),y=>p(195)(28),Cin=>p(196)(28),clock=>clock,reset=>reset,s=>p(258)(28),cout=>p(259)(29));
FA_ff_8198:FAff port map(x=>p(194)(29),y=>p(195)(29),Cin=>p(196)(29),clock=>clock,reset=>reset,s=>p(258)(29),cout=>p(259)(30));
FA_ff_8199:FAff port map(x=>p(194)(30),y=>p(195)(30),Cin=>p(196)(30),clock=>clock,reset=>reset,s=>p(258)(30),cout=>p(259)(31));
FA_ff_8200:FAff port map(x=>p(194)(31),y=>p(195)(31),Cin=>p(196)(31),clock=>clock,reset=>reset,s=>p(258)(31),cout=>p(259)(32));
FA_ff_8201:FAff port map(x=>p(194)(32),y=>p(195)(32),Cin=>p(196)(32),clock=>clock,reset=>reset,s=>p(258)(32),cout=>p(259)(33));
FA_ff_8202:FAff port map(x=>p(194)(33),y=>p(195)(33),Cin=>p(196)(33),clock=>clock,reset=>reset,s=>p(258)(33),cout=>p(259)(34));
FA_ff_8203:FAff port map(x=>p(194)(34),y=>p(195)(34),Cin=>p(196)(34),clock=>clock,reset=>reset,s=>p(258)(34),cout=>p(259)(35));
FA_ff_8204:FAff port map(x=>p(194)(35),y=>p(195)(35),Cin=>p(196)(35),clock=>clock,reset=>reset,s=>p(258)(35),cout=>p(259)(36));
FA_ff_8205:FAff port map(x=>p(194)(36),y=>p(195)(36),Cin=>p(196)(36),clock=>clock,reset=>reset,s=>p(258)(36),cout=>p(259)(37));
FA_ff_8206:FAff port map(x=>p(194)(37),y=>p(195)(37),Cin=>p(196)(37),clock=>clock,reset=>reset,s=>p(258)(37),cout=>p(259)(38));
FA_ff_8207:FAff port map(x=>p(194)(38),y=>p(195)(38),Cin=>p(196)(38),clock=>clock,reset=>reset,s=>p(258)(38),cout=>p(259)(39));
FA_ff_8208:FAff port map(x=>p(194)(39),y=>p(195)(39),Cin=>p(196)(39),clock=>clock,reset=>reset,s=>p(258)(39),cout=>p(259)(40));
FA_ff_8209:FAff port map(x=>p(194)(40),y=>p(195)(40),Cin=>p(196)(40),clock=>clock,reset=>reset,s=>p(258)(40),cout=>p(259)(41));
FA_ff_8210:FAff port map(x=>p(194)(41),y=>p(195)(41),Cin=>p(196)(41),clock=>clock,reset=>reset,s=>p(258)(41),cout=>p(259)(42));
FA_ff_8211:FAff port map(x=>p(194)(42),y=>p(195)(42),Cin=>p(196)(42),clock=>clock,reset=>reset,s=>p(258)(42),cout=>p(259)(43));
FA_ff_8212:FAff port map(x=>p(194)(43),y=>p(195)(43),Cin=>p(196)(43),clock=>clock,reset=>reset,s=>p(258)(43),cout=>p(259)(44));
FA_ff_8213:FAff port map(x=>p(194)(44),y=>p(195)(44),Cin=>p(196)(44),clock=>clock,reset=>reset,s=>p(258)(44),cout=>p(259)(45));
FA_ff_8214:FAff port map(x=>p(194)(45),y=>p(195)(45),Cin=>p(196)(45),clock=>clock,reset=>reset,s=>p(258)(45),cout=>p(259)(46));
FA_ff_8215:FAff port map(x=>p(194)(46),y=>p(195)(46),Cin=>p(196)(46),clock=>clock,reset=>reset,s=>p(258)(46),cout=>p(259)(47));
FA_ff_8216:FAff port map(x=>p(194)(47),y=>p(195)(47),Cin=>p(196)(47),clock=>clock,reset=>reset,s=>p(258)(47),cout=>p(259)(48));
FA_ff_8217:FAff port map(x=>p(194)(48),y=>p(195)(48),Cin=>p(196)(48),clock=>clock,reset=>reset,s=>p(258)(48),cout=>p(259)(49));
FA_ff_8218:FAff port map(x=>p(194)(49),y=>p(195)(49),Cin=>p(196)(49),clock=>clock,reset=>reset,s=>p(258)(49),cout=>p(259)(50));
FA_ff_8219:FAff port map(x=>p(194)(50),y=>p(195)(50),Cin=>p(196)(50),clock=>clock,reset=>reset,s=>p(258)(50),cout=>p(259)(51));
FA_ff_8220:FAff port map(x=>p(194)(51),y=>p(195)(51),Cin=>p(196)(51),clock=>clock,reset=>reset,s=>p(258)(51),cout=>p(259)(52));
FA_ff_8221:FAff port map(x=>p(194)(52),y=>p(195)(52),Cin=>p(196)(52),clock=>clock,reset=>reset,s=>p(258)(52),cout=>p(259)(53));
FA_ff_8222:FAff port map(x=>p(194)(53),y=>p(195)(53),Cin=>p(196)(53),clock=>clock,reset=>reset,s=>p(258)(53),cout=>p(259)(54));
FA_ff_8223:FAff port map(x=>p(194)(54),y=>p(195)(54),Cin=>p(196)(54),clock=>clock,reset=>reset,s=>p(258)(54),cout=>p(259)(55));
FA_ff_8224:FAff port map(x=>p(194)(55),y=>p(195)(55),Cin=>p(196)(55),clock=>clock,reset=>reset,s=>p(258)(55),cout=>p(259)(56));
FA_ff_8225:FAff port map(x=>p(194)(56),y=>p(195)(56),Cin=>p(196)(56),clock=>clock,reset=>reset,s=>p(258)(56),cout=>p(259)(57));
FA_ff_8226:FAff port map(x=>p(194)(57),y=>p(195)(57),Cin=>p(196)(57),clock=>clock,reset=>reset,s=>p(258)(57),cout=>p(259)(58));
FA_ff_8227:FAff port map(x=>p(194)(58),y=>p(195)(58),Cin=>p(196)(58),clock=>clock,reset=>reset,s=>p(258)(58),cout=>p(259)(59));
FA_ff_8228:FAff port map(x=>p(194)(59),y=>p(195)(59),Cin=>p(196)(59),clock=>clock,reset=>reset,s=>p(258)(59),cout=>p(259)(60));
FA_ff_8229:FAff port map(x=>p(194)(60),y=>p(195)(60),Cin=>p(196)(60),clock=>clock,reset=>reset,s=>p(258)(60),cout=>p(259)(61));
FA_ff_8230:FAff port map(x=>p(194)(61),y=>p(195)(61),Cin=>p(196)(61),clock=>clock,reset=>reset,s=>p(258)(61),cout=>p(259)(62));
FA_ff_8231:FAff port map(x=>p(194)(62),y=>p(195)(62),Cin=>p(196)(62),clock=>clock,reset=>reset,s=>p(258)(62),cout=>p(259)(63));
FA_ff_8232:FAff port map(x=>p(194)(63),y=>p(195)(63),Cin=>p(196)(63),clock=>clock,reset=>reset,s=>p(258)(63),cout=>p(259)(64));
FA_ff_8233:FAff port map(x=>p(194)(64),y=>p(195)(64),Cin=>p(196)(64),clock=>clock,reset=>reset,s=>p(258)(64),cout=>p(259)(65));
FA_ff_8234:FAff port map(x=>p(194)(65),y=>p(195)(65),Cin=>p(196)(65),clock=>clock,reset=>reset,s=>p(258)(65),cout=>p(259)(66));
FA_ff_8235:FAff port map(x=>p(194)(66),y=>p(195)(66),Cin=>p(196)(66),clock=>clock,reset=>reset,s=>p(258)(66),cout=>p(259)(67));
FA_ff_8236:FAff port map(x=>p(194)(67),y=>p(195)(67),Cin=>p(196)(67),clock=>clock,reset=>reset,s=>p(258)(67),cout=>p(259)(68));
FA_ff_8237:FAff port map(x=>p(194)(68),y=>p(195)(68),Cin=>p(196)(68),clock=>clock,reset=>reset,s=>p(258)(68),cout=>p(259)(69));
FA_ff_8238:FAff port map(x=>p(194)(69),y=>p(195)(69),Cin=>p(196)(69),clock=>clock,reset=>reset,s=>p(258)(69),cout=>p(259)(70));
FA_ff_8239:FAff port map(x=>p(194)(70),y=>p(195)(70),Cin=>p(196)(70),clock=>clock,reset=>reset,s=>p(258)(70),cout=>p(259)(71));
FA_ff_8240:FAff port map(x=>p(194)(71),y=>p(195)(71),Cin=>p(196)(71),clock=>clock,reset=>reset,s=>p(258)(71),cout=>p(259)(72));
FA_ff_8241:FAff port map(x=>p(194)(72),y=>p(195)(72),Cin=>p(196)(72),clock=>clock,reset=>reset,s=>p(258)(72),cout=>p(259)(73));
FA_ff_8242:FAff port map(x=>p(194)(73),y=>p(195)(73),Cin=>p(196)(73),clock=>clock,reset=>reset,s=>p(258)(73),cout=>p(259)(74));
FA_ff_8243:FAff port map(x=>p(194)(74),y=>p(195)(74),Cin=>p(196)(74),clock=>clock,reset=>reset,s=>p(258)(74),cout=>p(259)(75));
FA_ff_8244:FAff port map(x=>p(194)(75),y=>p(195)(75),Cin=>p(196)(75),clock=>clock,reset=>reset,s=>p(258)(75),cout=>p(259)(76));
FA_ff_8245:FAff port map(x=>p(194)(76),y=>p(195)(76),Cin=>p(196)(76),clock=>clock,reset=>reset,s=>p(258)(76),cout=>p(259)(77));
FA_ff_8246:FAff port map(x=>p(194)(77),y=>p(195)(77),Cin=>p(196)(77),clock=>clock,reset=>reset,s=>p(258)(77),cout=>p(259)(78));
FA_ff_8247:FAff port map(x=>p(194)(78),y=>p(195)(78),Cin=>p(196)(78),clock=>clock,reset=>reset,s=>p(258)(78),cout=>p(259)(79));
FA_ff_8248:FAff port map(x=>p(194)(79),y=>p(195)(79),Cin=>p(196)(79),clock=>clock,reset=>reset,s=>p(258)(79),cout=>p(259)(80));
FA_ff_8249:FAff port map(x=>p(194)(80),y=>p(195)(80),Cin=>p(196)(80),clock=>clock,reset=>reset,s=>p(258)(80),cout=>p(259)(81));
FA_ff_8250:FAff port map(x=>p(194)(81),y=>p(195)(81),Cin=>p(196)(81),clock=>clock,reset=>reset,s=>p(258)(81),cout=>p(259)(82));
FA_ff_8251:FAff port map(x=>p(194)(82),y=>p(195)(82),Cin=>p(196)(82),clock=>clock,reset=>reset,s=>p(258)(82),cout=>p(259)(83));
FA_ff_8252:FAff port map(x=>p(194)(83),y=>p(195)(83),Cin=>p(196)(83),clock=>clock,reset=>reset,s=>p(258)(83),cout=>p(259)(84));
FA_ff_8253:FAff port map(x=>p(194)(84),y=>p(195)(84),Cin=>p(196)(84),clock=>clock,reset=>reset,s=>p(258)(84),cout=>p(259)(85));
FA_ff_8254:FAff port map(x=>p(194)(85),y=>p(195)(85),Cin=>p(196)(85),clock=>clock,reset=>reset,s=>p(258)(85),cout=>p(259)(86));
FA_ff_8255:FAff port map(x=>p(194)(86),y=>p(195)(86),Cin=>p(196)(86),clock=>clock,reset=>reset,s=>p(258)(86),cout=>p(259)(87));
FA_ff_8256:FAff port map(x=>p(194)(87),y=>p(195)(87),Cin=>p(196)(87),clock=>clock,reset=>reset,s=>p(258)(87),cout=>p(259)(88));
FA_ff_8257:FAff port map(x=>p(194)(88),y=>p(195)(88),Cin=>p(196)(88),clock=>clock,reset=>reset,s=>p(258)(88),cout=>p(259)(89));
FA_ff_8258:FAff port map(x=>p(194)(89),y=>p(195)(89),Cin=>p(196)(89),clock=>clock,reset=>reset,s=>p(258)(89),cout=>p(259)(90));
FA_ff_8259:FAff port map(x=>p(194)(90),y=>p(195)(90),Cin=>p(196)(90),clock=>clock,reset=>reset,s=>p(258)(90),cout=>p(259)(91));
FA_ff_8260:FAff port map(x=>p(194)(91),y=>p(195)(91),Cin=>p(196)(91),clock=>clock,reset=>reset,s=>p(258)(91),cout=>p(259)(92));
FA_ff_8261:FAff port map(x=>p(194)(92),y=>p(195)(92),Cin=>p(196)(92),clock=>clock,reset=>reset,s=>p(258)(92),cout=>p(259)(93));
FA_ff_8262:FAff port map(x=>p(194)(93),y=>p(195)(93),Cin=>p(196)(93),clock=>clock,reset=>reset,s=>p(258)(93),cout=>p(259)(94));
FA_ff_8263:FAff port map(x=>p(194)(94),y=>p(195)(94),Cin=>p(196)(94),clock=>clock,reset=>reset,s=>p(258)(94),cout=>p(259)(95));
FA_ff_8264:FAff port map(x=>p(194)(95),y=>p(195)(95),Cin=>p(196)(95),clock=>clock,reset=>reset,s=>p(258)(95),cout=>p(259)(96));
FA_ff_8265:FAff port map(x=>p(194)(96),y=>p(195)(96),Cin=>p(196)(96),clock=>clock,reset=>reset,s=>p(258)(96),cout=>p(259)(97));
FA_ff_8266:FAff port map(x=>p(194)(97),y=>p(195)(97),Cin=>p(196)(97),clock=>clock,reset=>reset,s=>p(258)(97),cout=>p(259)(98));
FA_ff_8267:FAff port map(x=>p(194)(98),y=>p(195)(98),Cin=>p(196)(98),clock=>clock,reset=>reset,s=>p(258)(98),cout=>p(259)(99));
FA_ff_8268:FAff port map(x=>p(194)(99),y=>p(195)(99),Cin=>p(196)(99),clock=>clock,reset=>reset,s=>p(258)(99),cout=>p(259)(100));
FA_ff_8269:FAff port map(x=>p(194)(100),y=>p(195)(100),Cin=>p(196)(100),clock=>clock,reset=>reset,s=>p(258)(100),cout=>p(259)(101));
FA_ff_8270:FAff port map(x=>p(194)(101),y=>p(195)(101),Cin=>p(196)(101),clock=>clock,reset=>reset,s=>p(258)(101),cout=>p(259)(102));
FA_ff_8271:FAff port map(x=>p(194)(102),y=>p(195)(102),Cin=>p(196)(102),clock=>clock,reset=>reset,s=>p(258)(102),cout=>p(259)(103));
FA_ff_8272:FAff port map(x=>p(194)(103),y=>p(195)(103),Cin=>p(196)(103),clock=>clock,reset=>reset,s=>p(258)(103),cout=>p(259)(104));
FA_ff_8273:FAff port map(x=>p(194)(104),y=>p(195)(104),Cin=>p(196)(104),clock=>clock,reset=>reset,s=>p(258)(104),cout=>p(259)(105));
FA_ff_8274:FAff port map(x=>p(194)(105),y=>p(195)(105),Cin=>p(196)(105),clock=>clock,reset=>reset,s=>p(258)(105),cout=>p(259)(106));
FA_ff_8275:FAff port map(x=>p(194)(106),y=>p(195)(106),Cin=>p(196)(106),clock=>clock,reset=>reset,s=>p(258)(106),cout=>p(259)(107));
FA_ff_8276:FAff port map(x=>p(194)(107),y=>p(195)(107),Cin=>p(196)(107),clock=>clock,reset=>reset,s=>p(258)(107),cout=>p(259)(108));
FA_ff_8277:FAff port map(x=>p(194)(108),y=>p(195)(108),Cin=>p(196)(108),clock=>clock,reset=>reset,s=>p(258)(108),cout=>p(259)(109));
FA_ff_8278:FAff port map(x=>p(194)(109),y=>p(195)(109),Cin=>p(196)(109),clock=>clock,reset=>reset,s=>p(258)(109),cout=>p(259)(110));
FA_ff_8279:FAff port map(x=>p(194)(110),y=>p(195)(110),Cin=>p(196)(110),clock=>clock,reset=>reset,s=>p(258)(110),cout=>p(259)(111));
FA_ff_8280:FAff port map(x=>p(194)(111),y=>p(195)(111),Cin=>p(196)(111),clock=>clock,reset=>reset,s=>p(258)(111),cout=>p(259)(112));
FA_ff_8281:FAff port map(x=>p(194)(112),y=>p(195)(112),Cin=>p(196)(112),clock=>clock,reset=>reset,s=>p(258)(112),cout=>p(259)(113));
FA_ff_8282:FAff port map(x=>p(194)(113),y=>p(195)(113),Cin=>p(196)(113),clock=>clock,reset=>reset,s=>p(258)(113),cout=>p(259)(114));
FA_ff_8283:FAff port map(x=>p(194)(114),y=>p(195)(114),Cin=>p(196)(114),clock=>clock,reset=>reset,s=>p(258)(114),cout=>p(259)(115));
FA_ff_8284:FAff port map(x=>p(194)(115),y=>p(195)(115),Cin=>p(196)(115),clock=>clock,reset=>reset,s=>p(258)(115),cout=>p(259)(116));
FA_ff_8285:FAff port map(x=>p(194)(116),y=>p(195)(116),Cin=>p(196)(116),clock=>clock,reset=>reset,s=>p(258)(116),cout=>p(259)(117));
FA_ff_8286:FAff port map(x=>p(194)(117),y=>p(195)(117),Cin=>p(196)(117),clock=>clock,reset=>reset,s=>p(258)(117),cout=>p(259)(118));
FA_ff_8287:FAff port map(x=>p(194)(118),y=>p(195)(118),Cin=>p(196)(118),clock=>clock,reset=>reset,s=>p(258)(118),cout=>p(259)(119));
FA_ff_8288:FAff port map(x=>p(194)(119),y=>p(195)(119),Cin=>p(196)(119),clock=>clock,reset=>reset,s=>p(258)(119),cout=>p(259)(120));
FA_ff_8289:FAff port map(x=>p(194)(120),y=>p(195)(120),Cin=>p(196)(120),clock=>clock,reset=>reset,s=>p(258)(120),cout=>p(259)(121));
FA_ff_8290:FAff port map(x=>p(194)(121),y=>p(195)(121),Cin=>p(196)(121),clock=>clock,reset=>reset,s=>p(258)(121),cout=>p(259)(122));
FA_ff_8291:FAff port map(x=>p(194)(122),y=>p(195)(122),Cin=>p(196)(122),clock=>clock,reset=>reset,s=>p(258)(122),cout=>p(259)(123));
FA_ff_8292:FAff port map(x=>p(194)(123),y=>p(195)(123),Cin=>p(196)(123),clock=>clock,reset=>reset,s=>p(258)(123),cout=>p(259)(124));
FA_ff_8293:FAff port map(x=>p(194)(124),y=>p(195)(124),Cin=>p(196)(124),clock=>clock,reset=>reset,s=>p(258)(124),cout=>p(259)(125));
FA_ff_8294:FAff port map(x=>p(194)(125),y=>p(195)(125),Cin=>p(196)(125),clock=>clock,reset=>reset,s=>p(258)(125),cout=>p(259)(126));
FA_ff_8295:FAff port map(x=>p(194)(126),y=>p(195)(126),Cin=>p(196)(126),clock=>clock,reset=>reset,s=>p(258)(126),cout=>p(259)(127));
FA_ff_8296:FAff port map(x=>p(194)(127),y=>p(195)(127),Cin=>p(196)(127),clock=>clock,reset=>reset,s=>p(258)(127),cout=>p(259)(128));
p(258)(128)<=p(195)(128);
p(260)(0)<=p(198)(0);
FA_ff_8297:FAff port map(x=>p(197)(1),y=>p(198)(1),Cin=>p(199)(1),clock=>clock,reset=>reset,s=>p(260)(1),cout=>p(261)(2));
FA_ff_8298:FAff port map(x=>p(197)(2),y=>p(198)(2),Cin=>p(199)(2),clock=>clock,reset=>reset,s=>p(260)(2),cout=>p(261)(3));
FA_ff_8299:FAff port map(x=>p(197)(3),y=>p(198)(3),Cin=>p(199)(3),clock=>clock,reset=>reset,s=>p(260)(3),cout=>p(261)(4));
FA_ff_8300:FAff port map(x=>p(197)(4),y=>p(198)(4),Cin=>p(199)(4),clock=>clock,reset=>reset,s=>p(260)(4),cout=>p(261)(5));
FA_ff_8301:FAff port map(x=>p(197)(5),y=>p(198)(5),Cin=>p(199)(5),clock=>clock,reset=>reset,s=>p(260)(5),cout=>p(261)(6));
FA_ff_8302:FAff port map(x=>p(197)(6),y=>p(198)(6),Cin=>p(199)(6),clock=>clock,reset=>reset,s=>p(260)(6),cout=>p(261)(7));
FA_ff_8303:FAff port map(x=>p(197)(7),y=>p(198)(7),Cin=>p(199)(7),clock=>clock,reset=>reset,s=>p(260)(7),cout=>p(261)(8));
FA_ff_8304:FAff port map(x=>p(197)(8),y=>p(198)(8),Cin=>p(199)(8),clock=>clock,reset=>reset,s=>p(260)(8),cout=>p(261)(9));
FA_ff_8305:FAff port map(x=>p(197)(9),y=>p(198)(9),Cin=>p(199)(9),clock=>clock,reset=>reset,s=>p(260)(9),cout=>p(261)(10));
FA_ff_8306:FAff port map(x=>p(197)(10),y=>p(198)(10),Cin=>p(199)(10),clock=>clock,reset=>reset,s=>p(260)(10),cout=>p(261)(11));
FA_ff_8307:FAff port map(x=>p(197)(11),y=>p(198)(11),Cin=>p(199)(11),clock=>clock,reset=>reset,s=>p(260)(11),cout=>p(261)(12));
FA_ff_8308:FAff port map(x=>p(197)(12),y=>p(198)(12),Cin=>p(199)(12),clock=>clock,reset=>reset,s=>p(260)(12),cout=>p(261)(13));
FA_ff_8309:FAff port map(x=>p(197)(13),y=>p(198)(13),Cin=>p(199)(13),clock=>clock,reset=>reset,s=>p(260)(13),cout=>p(261)(14));
FA_ff_8310:FAff port map(x=>p(197)(14),y=>p(198)(14),Cin=>p(199)(14),clock=>clock,reset=>reset,s=>p(260)(14),cout=>p(261)(15));
FA_ff_8311:FAff port map(x=>p(197)(15),y=>p(198)(15),Cin=>p(199)(15),clock=>clock,reset=>reset,s=>p(260)(15),cout=>p(261)(16));
FA_ff_8312:FAff port map(x=>p(197)(16),y=>p(198)(16),Cin=>p(199)(16),clock=>clock,reset=>reset,s=>p(260)(16),cout=>p(261)(17));
FA_ff_8313:FAff port map(x=>p(197)(17),y=>p(198)(17),Cin=>p(199)(17),clock=>clock,reset=>reset,s=>p(260)(17),cout=>p(261)(18));
FA_ff_8314:FAff port map(x=>p(197)(18),y=>p(198)(18),Cin=>p(199)(18),clock=>clock,reset=>reset,s=>p(260)(18),cout=>p(261)(19));
FA_ff_8315:FAff port map(x=>p(197)(19),y=>p(198)(19),Cin=>p(199)(19),clock=>clock,reset=>reset,s=>p(260)(19),cout=>p(261)(20));
FA_ff_8316:FAff port map(x=>p(197)(20),y=>p(198)(20),Cin=>p(199)(20),clock=>clock,reset=>reset,s=>p(260)(20),cout=>p(261)(21));
FA_ff_8317:FAff port map(x=>p(197)(21),y=>p(198)(21),Cin=>p(199)(21),clock=>clock,reset=>reset,s=>p(260)(21),cout=>p(261)(22));
FA_ff_8318:FAff port map(x=>p(197)(22),y=>p(198)(22),Cin=>p(199)(22),clock=>clock,reset=>reset,s=>p(260)(22),cout=>p(261)(23));
FA_ff_8319:FAff port map(x=>p(197)(23),y=>p(198)(23),Cin=>p(199)(23),clock=>clock,reset=>reset,s=>p(260)(23),cout=>p(261)(24));
FA_ff_8320:FAff port map(x=>p(197)(24),y=>p(198)(24),Cin=>p(199)(24),clock=>clock,reset=>reset,s=>p(260)(24),cout=>p(261)(25));
FA_ff_8321:FAff port map(x=>p(197)(25),y=>p(198)(25),Cin=>p(199)(25),clock=>clock,reset=>reset,s=>p(260)(25),cout=>p(261)(26));
FA_ff_8322:FAff port map(x=>p(197)(26),y=>p(198)(26),Cin=>p(199)(26),clock=>clock,reset=>reset,s=>p(260)(26),cout=>p(261)(27));
FA_ff_8323:FAff port map(x=>p(197)(27),y=>p(198)(27),Cin=>p(199)(27),clock=>clock,reset=>reset,s=>p(260)(27),cout=>p(261)(28));
FA_ff_8324:FAff port map(x=>p(197)(28),y=>p(198)(28),Cin=>p(199)(28),clock=>clock,reset=>reset,s=>p(260)(28),cout=>p(261)(29));
FA_ff_8325:FAff port map(x=>p(197)(29),y=>p(198)(29),Cin=>p(199)(29),clock=>clock,reset=>reset,s=>p(260)(29),cout=>p(261)(30));
FA_ff_8326:FAff port map(x=>p(197)(30),y=>p(198)(30),Cin=>p(199)(30),clock=>clock,reset=>reset,s=>p(260)(30),cout=>p(261)(31));
FA_ff_8327:FAff port map(x=>p(197)(31),y=>p(198)(31),Cin=>p(199)(31),clock=>clock,reset=>reset,s=>p(260)(31),cout=>p(261)(32));
FA_ff_8328:FAff port map(x=>p(197)(32),y=>p(198)(32),Cin=>p(199)(32),clock=>clock,reset=>reset,s=>p(260)(32),cout=>p(261)(33));
FA_ff_8329:FAff port map(x=>p(197)(33),y=>p(198)(33),Cin=>p(199)(33),clock=>clock,reset=>reset,s=>p(260)(33),cout=>p(261)(34));
FA_ff_8330:FAff port map(x=>p(197)(34),y=>p(198)(34),Cin=>p(199)(34),clock=>clock,reset=>reset,s=>p(260)(34),cout=>p(261)(35));
FA_ff_8331:FAff port map(x=>p(197)(35),y=>p(198)(35),Cin=>p(199)(35),clock=>clock,reset=>reset,s=>p(260)(35),cout=>p(261)(36));
FA_ff_8332:FAff port map(x=>p(197)(36),y=>p(198)(36),Cin=>p(199)(36),clock=>clock,reset=>reset,s=>p(260)(36),cout=>p(261)(37));
FA_ff_8333:FAff port map(x=>p(197)(37),y=>p(198)(37),Cin=>p(199)(37),clock=>clock,reset=>reset,s=>p(260)(37),cout=>p(261)(38));
FA_ff_8334:FAff port map(x=>p(197)(38),y=>p(198)(38),Cin=>p(199)(38),clock=>clock,reset=>reset,s=>p(260)(38),cout=>p(261)(39));
FA_ff_8335:FAff port map(x=>p(197)(39),y=>p(198)(39),Cin=>p(199)(39),clock=>clock,reset=>reset,s=>p(260)(39),cout=>p(261)(40));
FA_ff_8336:FAff port map(x=>p(197)(40),y=>p(198)(40),Cin=>p(199)(40),clock=>clock,reset=>reset,s=>p(260)(40),cout=>p(261)(41));
FA_ff_8337:FAff port map(x=>p(197)(41),y=>p(198)(41),Cin=>p(199)(41),clock=>clock,reset=>reset,s=>p(260)(41),cout=>p(261)(42));
FA_ff_8338:FAff port map(x=>p(197)(42),y=>p(198)(42),Cin=>p(199)(42),clock=>clock,reset=>reset,s=>p(260)(42),cout=>p(261)(43));
FA_ff_8339:FAff port map(x=>p(197)(43),y=>p(198)(43),Cin=>p(199)(43),clock=>clock,reset=>reset,s=>p(260)(43),cout=>p(261)(44));
FA_ff_8340:FAff port map(x=>p(197)(44),y=>p(198)(44),Cin=>p(199)(44),clock=>clock,reset=>reset,s=>p(260)(44),cout=>p(261)(45));
FA_ff_8341:FAff port map(x=>p(197)(45),y=>p(198)(45),Cin=>p(199)(45),clock=>clock,reset=>reset,s=>p(260)(45),cout=>p(261)(46));
FA_ff_8342:FAff port map(x=>p(197)(46),y=>p(198)(46),Cin=>p(199)(46),clock=>clock,reset=>reset,s=>p(260)(46),cout=>p(261)(47));
FA_ff_8343:FAff port map(x=>p(197)(47),y=>p(198)(47),Cin=>p(199)(47),clock=>clock,reset=>reset,s=>p(260)(47),cout=>p(261)(48));
FA_ff_8344:FAff port map(x=>p(197)(48),y=>p(198)(48),Cin=>p(199)(48),clock=>clock,reset=>reset,s=>p(260)(48),cout=>p(261)(49));
FA_ff_8345:FAff port map(x=>p(197)(49),y=>p(198)(49),Cin=>p(199)(49),clock=>clock,reset=>reset,s=>p(260)(49),cout=>p(261)(50));
FA_ff_8346:FAff port map(x=>p(197)(50),y=>p(198)(50),Cin=>p(199)(50),clock=>clock,reset=>reset,s=>p(260)(50),cout=>p(261)(51));
FA_ff_8347:FAff port map(x=>p(197)(51),y=>p(198)(51),Cin=>p(199)(51),clock=>clock,reset=>reset,s=>p(260)(51),cout=>p(261)(52));
FA_ff_8348:FAff port map(x=>p(197)(52),y=>p(198)(52),Cin=>p(199)(52),clock=>clock,reset=>reset,s=>p(260)(52),cout=>p(261)(53));
FA_ff_8349:FAff port map(x=>p(197)(53),y=>p(198)(53),Cin=>p(199)(53),clock=>clock,reset=>reset,s=>p(260)(53),cout=>p(261)(54));
FA_ff_8350:FAff port map(x=>p(197)(54),y=>p(198)(54),Cin=>p(199)(54),clock=>clock,reset=>reset,s=>p(260)(54),cout=>p(261)(55));
FA_ff_8351:FAff port map(x=>p(197)(55),y=>p(198)(55),Cin=>p(199)(55),clock=>clock,reset=>reset,s=>p(260)(55),cout=>p(261)(56));
FA_ff_8352:FAff port map(x=>p(197)(56),y=>p(198)(56),Cin=>p(199)(56),clock=>clock,reset=>reset,s=>p(260)(56),cout=>p(261)(57));
FA_ff_8353:FAff port map(x=>p(197)(57),y=>p(198)(57),Cin=>p(199)(57),clock=>clock,reset=>reset,s=>p(260)(57),cout=>p(261)(58));
FA_ff_8354:FAff port map(x=>p(197)(58),y=>p(198)(58),Cin=>p(199)(58),clock=>clock,reset=>reset,s=>p(260)(58),cout=>p(261)(59));
FA_ff_8355:FAff port map(x=>p(197)(59),y=>p(198)(59),Cin=>p(199)(59),clock=>clock,reset=>reset,s=>p(260)(59),cout=>p(261)(60));
FA_ff_8356:FAff port map(x=>p(197)(60),y=>p(198)(60),Cin=>p(199)(60),clock=>clock,reset=>reset,s=>p(260)(60),cout=>p(261)(61));
FA_ff_8357:FAff port map(x=>p(197)(61),y=>p(198)(61),Cin=>p(199)(61),clock=>clock,reset=>reset,s=>p(260)(61),cout=>p(261)(62));
FA_ff_8358:FAff port map(x=>p(197)(62),y=>p(198)(62),Cin=>p(199)(62),clock=>clock,reset=>reset,s=>p(260)(62),cout=>p(261)(63));
FA_ff_8359:FAff port map(x=>p(197)(63),y=>p(198)(63),Cin=>p(199)(63),clock=>clock,reset=>reset,s=>p(260)(63),cout=>p(261)(64));
FA_ff_8360:FAff port map(x=>p(197)(64),y=>p(198)(64),Cin=>p(199)(64),clock=>clock,reset=>reset,s=>p(260)(64),cout=>p(261)(65));
FA_ff_8361:FAff port map(x=>p(197)(65),y=>p(198)(65),Cin=>p(199)(65),clock=>clock,reset=>reset,s=>p(260)(65),cout=>p(261)(66));
FA_ff_8362:FAff port map(x=>p(197)(66),y=>p(198)(66),Cin=>p(199)(66),clock=>clock,reset=>reset,s=>p(260)(66),cout=>p(261)(67));
FA_ff_8363:FAff port map(x=>p(197)(67),y=>p(198)(67),Cin=>p(199)(67),clock=>clock,reset=>reset,s=>p(260)(67),cout=>p(261)(68));
FA_ff_8364:FAff port map(x=>p(197)(68),y=>p(198)(68),Cin=>p(199)(68),clock=>clock,reset=>reset,s=>p(260)(68),cout=>p(261)(69));
FA_ff_8365:FAff port map(x=>p(197)(69),y=>p(198)(69),Cin=>p(199)(69),clock=>clock,reset=>reset,s=>p(260)(69),cout=>p(261)(70));
FA_ff_8366:FAff port map(x=>p(197)(70),y=>p(198)(70),Cin=>p(199)(70),clock=>clock,reset=>reset,s=>p(260)(70),cout=>p(261)(71));
FA_ff_8367:FAff port map(x=>p(197)(71),y=>p(198)(71),Cin=>p(199)(71),clock=>clock,reset=>reset,s=>p(260)(71),cout=>p(261)(72));
FA_ff_8368:FAff port map(x=>p(197)(72),y=>p(198)(72),Cin=>p(199)(72),clock=>clock,reset=>reset,s=>p(260)(72),cout=>p(261)(73));
FA_ff_8369:FAff port map(x=>p(197)(73),y=>p(198)(73),Cin=>p(199)(73),clock=>clock,reset=>reset,s=>p(260)(73),cout=>p(261)(74));
FA_ff_8370:FAff port map(x=>p(197)(74),y=>p(198)(74),Cin=>p(199)(74),clock=>clock,reset=>reset,s=>p(260)(74),cout=>p(261)(75));
FA_ff_8371:FAff port map(x=>p(197)(75),y=>p(198)(75),Cin=>p(199)(75),clock=>clock,reset=>reset,s=>p(260)(75),cout=>p(261)(76));
FA_ff_8372:FAff port map(x=>p(197)(76),y=>p(198)(76),Cin=>p(199)(76),clock=>clock,reset=>reset,s=>p(260)(76),cout=>p(261)(77));
FA_ff_8373:FAff port map(x=>p(197)(77),y=>p(198)(77),Cin=>p(199)(77),clock=>clock,reset=>reset,s=>p(260)(77),cout=>p(261)(78));
FA_ff_8374:FAff port map(x=>p(197)(78),y=>p(198)(78),Cin=>p(199)(78),clock=>clock,reset=>reset,s=>p(260)(78),cout=>p(261)(79));
FA_ff_8375:FAff port map(x=>p(197)(79),y=>p(198)(79),Cin=>p(199)(79),clock=>clock,reset=>reset,s=>p(260)(79),cout=>p(261)(80));
FA_ff_8376:FAff port map(x=>p(197)(80),y=>p(198)(80),Cin=>p(199)(80),clock=>clock,reset=>reset,s=>p(260)(80),cout=>p(261)(81));
FA_ff_8377:FAff port map(x=>p(197)(81),y=>p(198)(81),Cin=>p(199)(81),clock=>clock,reset=>reset,s=>p(260)(81),cout=>p(261)(82));
FA_ff_8378:FAff port map(x=>p(197)(82),y=>p(198)(82),Cin=>p(199)(82),clock=>clock,reset=>reset,s=>p(260)(82),cout=>p(261)(83));
FA_ff_8379:FAff port map(x=>p(197)(83),y=>p(198)(83),Cin=>p(199)(83),clock=>clock,reset=>reset,s=>p(260)(83),cout=>p(261)(84));
FA_ff_8380:FAff port map(x=>p(197)(84),y=>p(198)(84),Cin=>p(199)(84),clock=>clock,reset=>reset,s=>p(260)(84),cout=>p(261)(85));
FA_ff_8381:FAff port map(x=>p(197)(85),y=>p(198)(85),Cin=>p(199)(85),clock=>clock,reset=>reset,s=>p(260)(85),cout=>p(261)(86));
FA_ff_8382:FAff port map(x=>p(197)(86),y=>p(198)(86),Cin=>p(199)(86),clock=>clock,reset=>reset,s=>p(260)(86),cout=>p(261)(87));
FA_ff_8383:FAff port map(x=>p(197)(87),y=>p(198)(87),Cin=>p(199)(87),clock=>clock,reset=>reset,s=>p(260)(87),cout=>p(261)(88));
FA_ff_8384:FAff port map(x=>p(197)(88),y=>p(198)(88),Cin=>p(199)(88),clock=>clock,reset=>reset,s=>p(260)(88),cout=>p(261)(89));
FA_ff_8385:FAff port map(x=>p(197)(89),y=>p(198)(89),Cin=>p(199)(89),clock=>clock,reset=>reset,s=>p(260)(89),cout=>p(261)(90));
FA_ff_8386:FAff port map(x=>p(197)(90),y=>p(198)(90),Cin=>p(199)(90),clock=>clock,reset=>reset,s=>p(260)(90),cout=>p(261)(91));
FA_ff_8387:FAff port map(x=>p(197)(91),y=>p(198)(91),Cin=>p(199)(91),clock=>clock,reset=>reset,s=>p(260)(91),cout=>p(261)(92));
FA_ff_8388:FAff port map(x=>p(197)(92),y=>p(198)(92),Cin=>p(199)(92),clock=>clock,reset=>reset,s=>p(260)(92),cout=>p(261)(93));
FA_ff_8389:FAff port map(x=>p(197)(93),y=>p(198)(93),Cin=>p(199)(93),clock=>clock,reset=>reset,s=>p(260)(93),cout=>p(261)(94));
FA_ff_8390:FAff port map(x=>p(197)(94),y=>p(198)(94),Cin=>p(199)(94),clock=>clock,reset=>reset,s=>p(260)(94),cout=>p(261)(95));
FA_ff_8391:FAff port map(x=>p(197)(95),y=>p(198)(95),Cin=>p(199)(95),clock=>clock,reset=>reset,s=>p(260)(95),cout=>p(261)(96));
FA_ff_8392:FAff port map(x=>p(197)(96),y=>p(198)(96),Cin=>p(199)(96),clock=>clock,reset=>reset,s=>p(260)(96),cout=>p(261)(97));
FA_ff_8393:FAff port map(x=>p(197)(97),y=>p(198)(97),Cin=>p(199)(97),clock=>clock,reset=>reset,s=>p(260)(97),cout=>p(261)(98));
FA_ff_8394:FAff port map(x=>p(197)(98),y=>p(198)(98),Cin=>p(199)(98),clock=>clock,reset=>reset,s=>p(260)(98),cout=>p(261)(99));
FA_ff_8395:FAff port map(x=>p(197)(99),y=>p(198)(99),Cin=>p(199)(99),clock=>clock,reset=>reset,s=>p(260)(99),cout=>p(261)(100));
FA_ff_8396:FAff port map(x=>p(197)(100),y=>p(198)(100),Cin=>p(199)(100),clock=>clock,reset=>reset,s=>p(260)(100),cout=>p(261)(101));
FA_ff_8397:FAff port map(x=>p(197)(101),y=>p(198)(101),Cin=>p(199)(101),clock=>clock,reset=>reset,s=>p(260)(101),cout=>p(261)(102));
FA_ff_8398:FAff port map(x=>p(197)(102),y=>p(198)(102),Cin=>p(199)(102),clock=>clock,reset=>reset,s=>p(260)(102),cout=>p(261)(103));
FA_ff_8399:FAff port map(x=>p(197)(103),y=>p(198)(103),Cin=>p(199)(103),clock=>clock,reset=>reset,s=>p(260)(103),cout=>p(261)(104));
FA_ff_8400:FAff port map(x=>p(197)(104),y=>p(198)(104),Cin=>p(199)(104),clock=>clock,reset=>reset,s=>p(260)(104),cout=>p(261)(105));
FA_ff_8401:FAff port map(x=>p(197)(105),y=>p(198)(105),Cin=>p(199)(105),clock=>clock,reset=>reset,s=>p(260)(105),cout=>p(261)(106));
FA_ff_8402:FAff port map(x=>p(197)(106),y=>p(198)(106),Cin=>p(199)(106),clock=>clock,reset=>reset,s=>p(260)(106),cout=>p(261)(107));
FA_ff_8403:FAff port map(x=>p(197)(107),y=>p(198)(107),Cin=>p(199)(107),clock=>clock,reset=>reset,s=>p(260)(107),cout=>p(261)(108));
FA_ff_8404:FAff port map(x=>p(197)(108),y=>p(198)(108),Cin=>p(199)(108),clock=>clock,reset=>reset,s=>p(260)(108),cout=>p(261)(109));
FA_ff_8405:FAff port map(x=>p(197)(109),y=>p(198)(109),Cin=>p(199)(109),clock=>clock,reset=>reset,s=>p(260)(109),cout=>p(261)(110));
FA_ff_8406:FAff port map(x=>p(197)(110),y=>p(198)(110),Cin=>p(199)(110),clock=>clock,reset=>reset,s=>p(260)(110),cout=>p(261)(111));
FA_ff_8407:FAff port map(x=>p(197)(111),y=>p(198)(111),Cin=>p(199)(111),clock=>clock,reset=>reset,s=>p(260)(111),cout=>p(261)(112));
FA_ff_8408:FAff port map(x=>p(197)(112),y=>p(198)(112),Cin=>p(199)(112),clock=>clock,reset=>reset,s=>p(260)(112),cout=>p(261)(113));
FA_ff_8409:FAff port map(x=>p(197)(113),y=>p(198)(113),Cin=>p(199)(113),clock=>clock,reset=>reset,s=>p(260)(113),cout=>p(261)(114));
FA_ff_8410:FAff port map(x=>p(197)(114),y=>p(198)(114),Cin=>p(199)(114),clock=>clock,reset=>reset,s=>p(260)(114),cout=>p(261)(115));
FA_ff_8411:FAff port map(x=>p(197)(115),y=>p(198)(115),Cin=>p(199)(115),clock=>clock,reset=>reset,s=>p(260)(115),cout=>p(261)(116));
FA_ff_8412:FAff port map(x=>p(197)(116),y=>p(198)(116),Cin=>p(199)(116),clock=>clock,reset=>reset,s=>p(260)(116),cout=>p(261)(117));
FA_ff_8413:FAff port map(x=>p(197)(117),y=>p(198)(117),Cin=>p(199)(117),clock=>clock,reset=>reset,s=>p(260)(117),cout=>p(261)(118));
FA_ff_8414:FAff port map(x=>p(197)(118),y=>p(198)(118),Cin=>p(199)(118),clock=>clock,reset=>reset,s=>p(260)(118),cout=>p(261)(119));
FA_ff_8415:FAff port map(x=>p(197)(119),y=>p(198)(119),Cin=>p(199)(119),clock=>clock,reset=>reset,s=>p(260)(119),cout=>p(261)(120));
FA_ff_8416:FAff port map(x=>p(197)(120),y=>p(198)(120),Cin=>p(199)(120),clock=>clock,reset=>reset,s=>p(260)(120),cout=>p(261)(121));
FA_ff_8417:FAff port map(x=>p(197)(121),y=>p(198)(121),Cin=>p(199)(121),clock=>clock,reset=>reset,s=>p(260)(121),cout=>p(261)(122));
FA_ff_8418:FAff port map(x=>p(197)(122),y=>p(198)(122),Cin=>p(199)(122),clock=>clock,reset=>reset,s=>p(260)(122),cout=>p(261)(123));
FA_ff_8419:FAff port map(x=>p(197)(123),y=>p(198)(123),Cin=>p(199)(123),clock=>clock,reset=>reset,s=>p(260)(123),cout=>p(261)(124));
FA_ff_8420:FAff port map(x=>p(197)(124),y=>p(198)(124),Cin=>p(199)(124),clock=>clock,reset=>reset,s=>p(260)(124),cout=>p(261)(125));
FA_ff_8421:FAff port map(x=>p(197)(125),y=>p(198)(125),Cin=>p(199)(125),clock=>clock,reset=>reset,s=>p(260)(125),cout=>p(261)(126));
FA_ff_8422:FAff port map(x=>p(197)(126),y=>p(198)(126),Cin=>p(199)(126),clock=>clock,reset=>reset,s=>p(260)(126),cout=>p(261)(127));
FA_ff_8423:FAff port map(x=>p(197)(127),y=>p(198)(127),Cin=>p(199)(127),clock=>clock,reset=>reset,s=>p(260)(127),cout=>p(261)(128));
HA_ff_23:HAff port map(x=>p(197)(128),y=>p(199)(128),clock=>clock,reset=>reset,s=>p(260)(128),c=>p(261)(129));
HA_ff_24:HAff port map(x=>p(200)(0),y=>p(202)(0),clock=>clock,reset=>reset,s=>p(262)(0),c=>p(263)(1));
FA_ff_8424:FAff port map(x=>p(200)(1),y=>p(201)(1),Cin=>p(202)(1),clock=>clock,reset=>reset,s=>p(262)(1),cout=>p(263)(2));
FA_ff_8425:FAff port map(x=>p(200)(2),y=>p(201)(2),Cin=>p(202)(2),clock=>clock,reset=>reset,s=>p(262)(2),cout=>p(263)(3));
FA_ff_8426:FAff port map(x=>p(200)(3),y=>p(201)(3),Cin=>p(202)(3),clock=>clock,reset=>reset,s=>p(262)(3),cout=>p(263)(4));
FA_ff_8427:FAff port map(x=>p(200)(4),y=>p(201)(4),Cin=>p(202)(4),clock=>clock,reset=>reset,s=>p(262)(4),cout=>p(263)(5));
FA_ff_8428:FAff port map(x=>p(200)(5),y=>p(201)(5),Cin=>p(202)(5),clock=>clock,reset=>reset,s=>p(262)(5),cout=>p(263)(6));
FA_ff_8429:FAff port map(x=>p(200)(6),y=>p(201)(6),Cin=>p(202)(6),clock=>clock,reset=>reset,s=>p(262)(6),cout=>p(263)(7));
FA_ff_8430:FAff port map(x=>p(200)(7),y=>p(201)(7),Cin=>p(202)(7),clock=>clock,reset=>reset,s=>p(262)(7),cout=>p(263)(8));
FA_ff_8431:FAff port map(x=>p(200)(8),y=>p(201)(8),Cin=>p(202)(8),clock=>clock,reset=>reset,s=>p(262)(8),cout=>p(263)(9));
FA_ff_8432:FAff port map(x=>p(200)(9),y=>p(201)(9),Cin=>p(202)(9),clock=>clock,reset=>reset,s=>p(262)(9),cout=>p(263)(10));
FA_ff_8433:FAff port map(x=>p(200)(10),y=>p(201)(10),Cin=>p(202)(10),clock=>clock,reset=>reset,s=>p(262)(10),cout=>p(263)(11));
FA_ff_8434:FAff port map(x=>p(200)(11),y=>p(201)(11),Cin=>p(202)(11),clock=>clock,reset=>reset,s=>p(262)(11),cout=>p(263)(12));
FA_ff_8435:FAff port map(x=>p(200)(12),y=>p(201)(12),Cin=>p(202)(12),clock=>clock,reset=>reset,s=>p(262)(12),cout=>p(263)(13));
FA_ff_8436:FAff port map(x=>p(200)(13),y=>p(201)(13),Cin=>p(202)(13),clock=>clock,reset=>reset,s=>p(262)(13),cout=>p(263)(14));
FA_ff_8437:FAff port map(x=>p(200)(14),y=>p(201)(14),Cin=>p(202)(14),clock=>clock,reset=>reset,s=>p(262)(14),cout=>p(263)(15));
FA_ff_8438:FAff port map(x=>p(200)(15),y=>p(201)(15),Cin=>p(202)(15),clock=>clock,reset=>reset,s=>p(262)(15),cout=>p(263)(16));
FA_ff_8439:FAff port map(x=>p(200)(16),y=>p(201)(16),Cin=>p(202)(16),clock=>clock,reset=>reset,s=>p(262)(16),cout=>p(263)(17));
FA_ff_8440:FAff port map(x=>p(200)(17),y=>p(201)(17),Cin=>p(202)(17),clock=>clock,reset=>reset,s=>p(262)(17),cout=>p(263)(18));
FA_ff_8441:FAff port map(x=>p(200)(18),y=>p(201)(18),Cin=>p(202)(18),clock=>clock,reset=>reset,s=>p(262)(18),cout=>p(263)(19));
FA_ff_8442:FAff port map(x=>p(200)(19),y=>p(201)(19),Cin=>p(202)(19),clock=>clock,reset=>reset,s=>p(262)(19),cout=>p(263)(20));
FA_ff_8443:FAff port map(x=>p(200)(20),y=>p(201)(20),Cin=>p(202)(20),clock=>clock,reset=>reset,s=>p(262)(20),cout=>p(263)(21));
FA_ff_8444:FAff port map(x=>p(200)(21),y=>p(201)(21),Cin=>p(202)(21),clock=>clock,reset=>reset,s=>p(262)(21),cout=>p(263)(22));
FA_ff_8445:FAff port map(x=>p(200)(22),y=>p(201)(22),Cin=>p(202)(22),clock=>clock,reset=>reset,s=>p(262)(22),cout=>p(263)(23));
FA_ff_8446:FAff port map(x=>p(200)(23),y=>p(201)(23),Cin=>p(202)(23),clock=>clock,reset=>reset,s=>p(262)(23),cout=>p(263)(24));
FA_ff_8447:FAff port map(x=>p(200)(24),y=>p(201)(24),Cin=>p(202)(24),clock=>clock,reset=>reset,s=>p(262)(24),cout=>p(263)(25));
FA_ff_8448:FAff port map(x=>p(200)(25),y=>p(201)(25),Cin=>p(202)(25),clock=>clock,reset=>reset,s=>p(262)(25),cout=>p(263)(26));
FA_ff_8449:FAff port map(x=>p(200)(26),y=>p(201)(26),Cin=>p(202)(26),clock=>clock,reset=>reset,s=>p(262)(26),cout=>p(263)(27));
FA_ff_8450:FAff port map(x=>p(200)(27),y=>p(201)(27),Cin=>p(202)(27),clock=>clock,reset=>reset,s=>p(262)(27),cout=>p(263)(28));
FA_ff_8451:FAff port map(x=>p(200)(28),y=>p(201)(28),Cin=>p(202)(28),clock=>clock,reset=>reset,s=>p(262)(28),cout=>p(263)(29));
FA_ff_8452:FAff port map(x=>p(200)(29),y=>p(201)(29),Cin=>p(202)(29),clock=>clock,reset=>reset,s=>p(262)(29),cout=>p(263)(30));
FA_ff_8453:FAff port map(x=>p(200)(30),y=>p(201)(30),Cin=>p(202)(30),clock=>clock,reset=>reset,s=>p(262)(30),cout=>p(263)(31));
FA_ff_8454:FAff port map(x=>p(200)(31),y=>p(201)(31),Cin=>p(202)(31),clock=>clock,reset=>reset,s=>p(262)(31),cout=>p(263)(32));
FA_ff_8455:FAff port map(x=>p(200)(32),y=>p(201)(32),Cin=>p(202)(32),clock=>clock,reset=>reset,s=>p(262)(32),cout=>p(263)(33));
FA_ff_8456:FAff port map(x=>p(200)(33),y=>p(201)(33),Cin=>p(202)(33),clock=>clock,reset=>reset,s=>p(262)(33),cout=>p(263)(34));
FA_ff_8457:FAff port map(x=>p(200)(34),y=>p(201)(34),Cin=>p(202)(34),clock=>clock,reset=>reset,s=>p(262)(34),cout=>p(263)(35));
FA_ff_8458:FAff port map(x=>p(200)(35),y=>p(201)(35),Cin=>p(202)(35),clock=>clock,reset=>reset,s=>p(262)(35),cout=>p(263)(36));
FA_ff_8459:FAff port map(x=>p(200)(36),y=>p(201)(36),Cin=>p(202)(36),clock=>clock,reset=>reset,s=>p(262)(36),cout=>p(263)(37));
FA_ff_8460:FAff port map(x=>p(200)(37),y=>p(201)(37),Cin=>p(202)(37),clock=>clock,reset=>reset,s=>p(262)(37),cout=>p(263)(38));
FA_ff_8461:FAff port map(x=>p(200)(38),y=>p(201)(38),Cin=>p(202)(38),clock=>clock,reset=>reset,s=>p(262)(38),cout=>p(263)(39));
FA_ff_8462:FAff port map(x=>p(200)(39),y=>p(201)(39),Cin=>p(202)(39),clock=>clock,reset=>reset,s=>p(262)(39),cout=>p(263)(40));
FA_ff_8463:FAff port map(x=>p(200)(40),y=>p(201)(40),Cin=>p(202)(40),clock=>clock,reset=>reset,s=>p(262)(40),cout=>p(263)(41));
FA_ff_8464:FAff port map(x=>p(200)(41),y=>p(201)(41),Cin=>p(202)(41),clock=>clock,reset=>reset,s=>p(262)(41),cout=>p(263)(42));
FA_ff_8465:FAff port map(x=>p(200)(42),y=>p(201)(42),Cin=>p(202)(42),clock=>clock,reset=>reset,s=>p(262)(42),cout=>p(263)(43));
FA_ff_8466:FAff port map(x=>p(200)(43),y=>p(201)(43),Cin=>p(202)(43),clock=>clock,reset=>reset,s=>p(262)(43),cout=>p(263)(44));
FA_ff_8467:FAff port map(x=>p(200)(44),y=>p(201)(44),Cin=>p(202)(44),clock=>clock,reset=>reset,s=>p(262)(44),cout=>p(263)(45));
FA_ff_8468:FAff port map(x=>p(200)(45),y=>p(201)(45),Cin=>p(202)(45),clock=>clock,reset=>reset,s=>p(262)(45),cout=>p(263)(46));
FA_ff_8469:FAff port map(x=>p(200)(46),y=>p(201)(46),Cin=>p(202)(46),clock=>clock,reset=>reset,s=>p(262)(46),cout=>p(263)(47));
FA_ff_8470:FAff port map(x=>p(200)(47),y=>p(201)(47),Cin=>p(202)(47),clock=>clock,reset=>reset,s=>p(262)(47),cout=>p(263)(48));
FA_ff_8471:FAff port map(x=>p(200)(48),y=>p(201)(48),Cin=>p(202)(48),clock=>clock,reset=>reset,s=>p(262)(48),cout=>p(263)(49));
FA_ff_8472:FAff port map(x=>p(200)(49),y=>p(201)(49),Cin=>p(202)(49),clock=>clock,reset=>reset,s=>p(262)(49),cout=>p(263)(50));
FA_ff_8473:FAff port map(x=>p(200)(50),y=>p(201)(50),Cin=>p(202)(50),clock=>clock,reset=>reset,s=>p(262)(50),cout=>p(263)(51));
FA_ff_8474:FAff port map(x=>p(200)(51),y=>p(201)(51),Cin=>p(202)(51),clock=>clock,reset=>reset,s=>p(262)(51),cout=>p(263)(52));
FA_ff_8475:FAff port map(x=>p(200)(52),y=>p(201)(52),Cin=>p(202)(52),clock=>clock,reset=>reset,s=>p(262)(52),cout=>p(263)(53));
FA_ff_8476:FAff port map(x=>p(200)(53),y=>p(201)(53),Cin=>p(202)(53),clock=>clock,reset=>reset,s=>p(262)(53),cout=>p(263)(54));
FA_ff_8477:FAff port map(x=>p(200)(54),y=>p(201)(54),Cin=>p(202)(54),clock=>clock,reset=>reset,s=>p(262)(54),cout=>p(263)(55));
FA_ff_8478:FAff port map(x=>p(200)(55),y=>p(201)(55),Cin=>p(202)(55),clock=>clock,reset=>reset,s=>p(262)(55),cout=>p(263)(56));
FA_ff_8479:FAff port map(x=>p(200)(56),y=>p(201)(56),Cin=>p(202)(56),clock=>clock,reset=>reset,s=>p(262)(56),cout=>p(263)(57));
FA_ff_8480:FAff port map(x=>p(200)(57),y=>p(201)(57),Cin=>p(202)(57),clock=>clock,reset=>reset,s=>p(262)(57),cout=>p(263)(58));
FA_ff_8481:FAff port map(x=>p(200)(58),y=>p(201)(58),Cin=>p(202)(58),clock=>clock,reset=>reset,s=>p(262)(58),cout=>p(263)(59));
FA_ff_8482:FAff port map(x=>p(200)(59),y=>p(201)(59),Cin=>p(202)(59),clock=>clock,reset=>reset,s=>p(262)(59),cout=>p(263)(60));
FA_ff_8483:FAff port map(x=>p(200)(60),y=>p(201)(60),Cin=>p(202)(60),clock=>clock,reset=>reset,s=>p(262)(60),cout=>p(263)(61));
FA_ff_8484:FAff port map(x=>p(200)(61),y=>p(201)(61),Cin=>p(202)(61),clock=>clock,reset=>reset,s=>p(262)(61),cout=>p(263)(62));
FA_ff_8485:FAff port map(x=>p(200)(62),y=>p(201)(62),Cin=>p(202)(62),clock=>clock,reset=>reset,s=>p(262)(62),cout=>p(263)(63));
FA_ff_8486:FAff port map(x=>p(200)(63),y=>p(201)(63),Cin=>p(202)(63),clock=>clock,reset=>reset,s=>p(262)(63),cout=>p(263)(64));
FA_ff_8487:FAff port map(x=>p(200)(64),y=>p(201)(64),Cin=>p(202)(64),clock=>clock,reset=>reset,s=>p(262)(64),cout=>p(263)(65));
FA_ff_8488:FAff port map(x=>p(200)(65),y=>p(201)(65),Cin=>p(202)(65),clock=>clock,reset=>reset,s=>p(262)(65),cout=>p(263)(66));
FA_ff_8489:FAff port map(x=>p(200)(66),y=>p(201)(66),Cin=>p(202)(66),clock=>clock,reset=>reset,s=>p(262)(66),cout=>p(263)(67));
FA_ff_8490:FAff port map(x=>p(200)(67),y=>p(201)(67),Cin=>p(202)(67),clock=>clock,reset=>reset,s=>p(262)(67),cout=>p(263)(68));
FA_ff_8491:FAff port map(x=>p(200)(68),y=>p(201)(68),Cin=>p(202)(68),clock=>clock,reset=>reset,s=>p(262)(68),cout=>p(263)(69));
FA_ff_8492:FAff port map(x=>p(200)(69),y=>p(201)(69),Cin=>p(202)(69),clock=>clock,reset=>reset,s=>p(262)(69),cout=>p(263)(70));
FA_ff_8493:FAff port map(x=>p(200)(70),y=>p(201)(70),Cin=>p(202)(70),clock=>clock,reset=>reset,s=>p(262)(70),cout=>p(263)(71));
FA_ff_8494:FAff port map(x=>p(200)(71),y=>p(201)(71),Cin=>p(202)(71),clock=>clock,reset=>reset,s=>p(262)(71),cout=>p(263)(72));
FA_ff_8495:FAff port map(x=>p(200)(72),y=>p(201)(72),Cin=>p(202)(72),clock=>clock,reset=>reset,s=>p(262)(72),cout=>p(263)(73));
FA_ff_8496:FAff port map(x=>p(200)(73),y=>p(201)(73),Cin=>p(202)(73),clock=>clock,reset=>reset,s=>p(262)(73),cout=>p(263)(74));
FA_ff_8497:FAff port map(x=>p(200)(74),y=>p(201)(74),Cin=>p(202)(74),clock=>clock,reset=>reset,s=>p(262)(74),cout=>p(263)(75));
FA_ff_8498:FAff port map(x=>p(200)(75),y=>p(201)(75),Cin=>p(202)(75),clock=>clock,reset=>reset,s=>p(262)(75),cout=>p(263)(76));
FA_ff_8499:FAff port map(x=>p(200)(76),y=>p(201)(76),Cin=>p(202)(76),clock=>clock,reset=>reset,s=>p(262)(76),cout=>p(263)(77));
FA_ff_8500:FAff port map(x=>p(200)(77),y=>p(201)(77),Cin=>p(202)(77),clock=>clock,reset=>reset,s=>p(262)(77),cout=>p(263)(78));
FA_ff_8501:FAff port map(x=>p(200)(78),y=>p(201)(78),Cin=>p(202)(78),clock=>clock,reset=>reset,s=>p(262)(78),cout=>p(263)(79));
FA_ff_8502:FAff port map(x=>p(200)(79),y=>p(201)(79),Cin=>p(202)(79),clock=>clock,reset=>reset,s=>p(262)(79),cout=>p(263)(80));
FA_ff_8503:FAff port map(x=>p(200)(80),y=>p(201)(80),Cin=>p(202)(80),clock=>clock,reset=>reset,s=>p(262)(80),cout=>p(263)(81));
FA_ff_8504:FAff port map(x=>p(200)(81),y=>p(201)(81),Cin=>p(202)(81),clock=>clock,reset=>reset,s=>p(262)(81),cout=>p(263)(82));
FA_ff_8505:FAff port map(x=>p(200)(82),y=>p(201)(82),Cin=>p(202)(82),clock=>clock,reset=>reset,s=>p(262)(82),cout=>p(263)(83));
FA_ff_8506:FAff port map(x=>p(200)(83),y=>p(201)(83),Cin=>p(202)(83),clock=>clock,reset=>reset,s=>p(262)(83),cout=>p(263)(84));
FA_ff_8507:FAff port map(x=>p(200)(84),y=>p(201)(84),Cin=>p(202)(84),clock=>clock,reset=>reset,s=>p(262)(84),cout=>p(263)(85));
FA_ff_8508:FAff port map(x=>p(200)(85),y=>p(201)(85),Cin=>p(202)(85),clock=>clock,reset=>reset,s=>p(262)(85),cout=>p(263)(86));
FA_ff_8509:FAff port map(x=>p(200)(86),y=>p(201)(86),Cin=>p(202)(86),clock=>clock,reset=>reset,s=>p(262)(86),cout=>p(263)(87));
FA_ff_8510:FAff port map(x=>p(200)(87),y=>p(201)(87),Cin=>p(202)(87),clock=>clock,reset=>reset,s=>p(262)(87),cout=>p(263)(88));
FA_ff_8511:FAff port map(x=>p(200)(88),y=>p(201)(88),Cin=>p(202)(88),clock=>clock,reset=>reset,s=>p(262)(88),cout=>p(263)(89));
FA_ff_8512:FAff port map(x=>p(200)(89),y=>p(201)(89),Cin=>p(202)(89),clock=>clock,reset=>reset,s=>p(262)(89),cout=>p(263)(90));
FA_ff_8513:FAff port map(x=>p(200)(90),y=>p(201)(90),Cin=>p(202)(90),clock=>clock,reset=>reset,s=>p(262)(90),cout=>p(263)(91));
FA_ff_8514:FAff port map(x=>p(200)(91),y=>p(201)(91),Cin=>p(202)(91),clock=>clock,reset=>reset,s=>p(262)(91),cout=>p(263)(92));
FA_ff_8515:FAff port map(x=>p(200)(92),y=>p(201)(92),Cin=>p(202)(92),clock=>clock,reset=>reset,s=>p(262)(92),cout=>p(263)(93));
FA_ff_8516:FAff port map(x=>p(200)(93),y=>p(201)(93),Cin=>p(202)(93),clock=>clock,reset=>reset,s=>p(262)(93),cout=>p(263)(94));
FA_ff_8517:FAff port map(x=>p(200)(94),y=>p(201)(94),Cin=>p(202)(94),clock=>clock,reset=>reset,s=>p(262)(94),cout=>p(263)(95));
FA_ff_8518:FAff port map(x=>p(200)(95),y=>p(201)(95),Cin=>p(202)(95),clock=>clock,reset=>reset,s=>p(262)(95),cout=>p(263)(96));
FA_ff_8519:FAff port map(x=>p(200)(96),y=>p(201)(96),Cin=>p(202)(96),clock=>clock,reset=>reset,s=>p(262)(96),cout=>p(263)(97));
FA_ff_8520:FAff port map(x=>p(200)(97),y=>p(201)(97),Cin=>p(202)(97),clock=>clock,reset=>reset,s=>p(262)(97),cout=>p(263)(98));
FA_ff_8521:FAff port map(x=>p(200)(98),y=>p(201)(98),Cin=>p(202)(98),clock=>clock,reset=>reset,s=>p(262)(98),cout=>p(263)(99));
FA_ff_8522:FAff port map(x=>p(200)(99),y=>p(201)(99),Cin=>p(202)(99),clock=>clock,reset=>reset,s=>p(262)(99),cout=>p(263)(100));
FA_ff_8523:FAff port map(x=>p(200)(100),y=>p(201)(100),Cin=>p(202)(100),clock=>clock,reset=>reset,s=>p(262)(100),cout=>p(263)(101));
FA_ff_8524:FAff port map(x=>p(200)(101),y=>p(201)(101),Cin=>p(202)(101),clock=>clock,reset=>reset,s=>p(262)(101),cout=>p(263)(102));
FA_ff_8525:FAff port map(x=>p(200)(102),y=>p(201)(102),Cin=>p(202)(102),clock=>clock,reset=>reset,s=>p(262)(102),cout=>p(263)(103));
FA_ff_8526:FAff port map(x=>p(200)(103),y=>p(201)(103),Cin=>p(202)(103),clock=>clock,reset=>reset,s=>p(262)(103),cout=>p(263)(104));
FA_ff_8527:FAff port map(x=>p(200)(104),y=>p(201)(104),Cin=>p(202)(104),clock=>clock,reset=>reset,s=>p(262)(104),cout=>p(263)(105));
FA_ff_8528:FAff port map(x=>p(200)(105),y=>p(201)(105),Cin=>p(202)(105),clock=>clock,reset=>reset,s=>p(262)(105),cout=>p(263)(106));
FA_ff_8529:FAff port map(x=>p(200)(106),y=>p(201)(106),Cin=>p(202)(106),clock=>clock,reset=>reset,s=>p(262)(106),cout=>p(263)(107));
FA_ff_8530:FAff port map(x=>p(200)(107),y=>p(201)(107),Cin=>p(202)(107),clock=>clock,reset=>reset,s=>p(262)(107),cout=>p(263)(108));
FA_ff_8531:FAff port map(x=>p(200)(108),y=>p(201)(108),Cin=>p(202)(108),clock=>clock,reset=>reset,s=>p(262)(108),cout=>p(263)(109));
FA_ff_8532:FAff port map(x=>p(200)(109),y=>p(201)(109),Cin=>p(202)(109),clock=>clock,reset=>reset,s=>p(262)(109),cout=>p(263)(110));
FA_ff_8533:FAff port map(x=>p(200)(110),y=>p(201)(110),Cin=>p(202)(110),clock=>clock,reset=>reset,s=>p(262)(110),cout=>p(263)(111));
FA_ff_8534:FAff port map(x=>p(200)(111),y=>p(201)(111),Cin=>p(202)(111),clock=>clock,reset=>reset,s=>p(262)(111),cout=>p(263)(112));
FA_ff_8535:FAff port map(x=>p(200)(112),y=>p(201)(112),Cin=>p(202)(112),clock=>clock,reset=>reset,s=>p(262)(112),cout=>p(263)(113));
FA_ff_8536:FAff port map(x=>p(200)(113),y=>p(201)(113),Cin=>p(202)(113),clock=>clock,reset=>reset,s=>p(262)(113),cout=>p(263)(114));
FA_ff_8537:FAff port map(x=>p(200)(114),y=>p(201)(114),Cin=>p(202)(114),clock=>clock,reset=>reset,s=>p(262)(114),cout=>p(263)(115));
FA_ff_8538:FAff port map(x=>p(200)(115),y=>p(201)(115),Cin=>p(202)(115),clock=>clock,reset=>reset,s=>p(262)(115),cout=>p(263)(116));
FA_ff_8539:FAff port map(x=>p(200)(116),y=>p(201)(116),Cin=>p(202)(116),clock=>clock,reset=>reset,s=>p(262)(116),cout=>p(263)(117));
FA_ff_8540:FAff port map(x=>p(200)(117),y=>p(201)(117),Cin=>p(202)(117),clock=>clock,reset=>reset,s=>p(262)(117),cout=>p(263)(118));
FA_ff_8541:FAff port map(x=>p(200)(118),y=>p(201)(118),Cin=>p(202)(118),clock=>clock,reset=>reset,s=>p(262)(118),cout=>p(263)(119));
FA_ff_8542:FAff port map(x=>p(200)(119),y=>p(201)(119),Cin=>p(202)(119),clock=>clock,reset=>reset,s=>p(262)(119),cout=>p(263)(120));
FA_ff_8543:FAff port map(x=>p(200)(120),y=>p(201)(120),Cin=>p(202)(120),clock=>clock,reset=>reset,s=>p(262)(120),cout=>p(263)(121));
FA_ff_8544:FAff port map(x=>p(200)(121),y=>p(201)(121),Cin=>p(202)(121),clock=>clock,reset=>reset,s=>p(262)(121),cout=>p(263)(122));
FA_ff_8545:FAff port map(x=>p(200)(122),y=>p(201)(122),Cin=>p(202)(122),clock=>clock,reset=>reset,s=>p(262)(122),cout=>p(263)(123));
FA_ff_8546:FAff port map(x=>p(200)(123),y=>p(201)(123),Cin=>p(202)(123),clock=>clock,reset=>reset,s=>p(262)(123),cout=>p(263)(124));
FA_ff_8547:FAff port map(x=>p(200)(124),y=>p(201)(124),Cin=>p(202)(124),clock=>clock,reset=>reset,s=>p(262)(124),cout=>p(263)(125));
FA_ff_8548:FAff port map(x=>p(200)(125),y=>p(201)(125),Cin=>p(202)(125),clock=>clock,reset=>reset,s=>p(262)(125),cout=>p(263)(126));
FA_ff_8549:FAff port map(x=>p(200)(126),y=>p(201)(126),Cin=>p(202)(126),clock=>clock,reset=>reset,s=>p(262)(126),cout=>p(263)(127));
FA_ff_8550:FAff port map(x=>p(200)(127),y=>p(201)(127),Cin=>p(202)(127),clock=>clock,reset=>reset,s=>p(262)(127),cout=>p(263)(128));
p(262)(128)<=p(201)(128);
p(264)(0)<=p(204)(0);
FA_ff_8551:FAff port map(x=>p(203)(1),y=>p(204)(1),Cin=>p(205)(1),clock=>clock,reset=>reset,s=>p(264)(1),cout=>p(265)(2));
FA_ff_8552:FAff port map(x=>p(203)(2),y=>p(204)(2),Cin=>p(205)(2),clock=>clock,reset=>reset,s=>p(264)(2),cout=>p(265)(3));
FA_ff_8553:FAff port map(x=>p(203)(3),y=>p(204)(3),Cin=>p(205)(3),clock=>clock,reset=>reset,s=>p(264)(3),cout=>p(265)(4));
FA_ff_8554:FAff port map(x=>p(203)(4),y=>p(204)(4),Cin=>p(205)(4),clock=>clock,reset=>reset,s=>p(264)(4),cout=>p(265)(5));
FA_ff_8555:FAff port map(x=>p(203)(5),y=>p(204)(5),Cin=>p(205)(5),clock=>clock,reset=>reset,s=>p(264)(5),cout=>p(265)(6));
FA_ff_8556:FAff port map(x=>p(203)(6),y=>p(204)(6),Cin=>p(205)(6),clock=>clock,reset=>reset,s=>p(264)(6),cout=>p(265)(7));
FA_ff_8557:FAff port map(x=>p(203)(7),y=>p(204)(7),Cin=>p(205)(7),clock=>clock,reset=>reset,s=>p(264)(7),cout=>p(265)(8));
FA_ff_8558:FAff port map(x=>p(203)(8),y=>p(204)(8),Cin=>p(205)(8),clock=>clock,reset=>reset,s=>p(264)(8),cout=>p(265)(9));
FA_ff_8559:FAff port map(x=>p(203)(9),y=>p(204)(9),Cin=>p(205)(9),clock=>clock,reset=>reset,s=>p(264)(9),cout=>p(265)(10));
FA_ff_8560:FAff port map(x=>p(203)(10),y=>p(204)(10),Cin=>p(205)(10),clock=>clock,reset=>reset,s=>p(264)(10),cout=>p(265)(11));
FA_ff_8561:FAff port map(x=>p(203)(11),y=>p(204)(11),Cin=>p(205)(11),clock=>clock,reset=>reset,s=>p(264)(11),cout=>p(265)(12));
FA_ff_8562:FAff port map(x=>p(203)(12),y=>p(204)(12),Cin=>p(205)(12),clock=>clock,reset=>reset,s=>p(264)(12),cout=>p(265)(13));
FA_ff_8563:FAff port map(x=>p(203)(13),y=>p(204)(13),Cin=>p(205)(13),clock=>clock,reset=>reset,s=>p(264)(13),cout=>p(265)(14));
FA_ff_8564:FAff port map(x=>p(203)(14),y=>p(204)(14),Cin=>p(205)(14),clock=>clock,reset=>reset,s=>p(264)(14),cout=>p(265)(15));
FA_ff_8565:FAff port map(x=>p(203)(15),y=>p(204)(15),Cin=>p(205)(15),clock=>clock,reset=>reset,s=>p(264)(15),cout=>p(265)(16));
FA_ff_8566:FAff port map(x=>p(203)(16),y=>p(204)(16),Cin=>p(205)(16),clock=>clock,reset=>reset,s=>p(264)(16),cout=>p(265)(17));
FA_ff_8567:FAff port map(x=>p(203)(17),y=>p(204)(17),Cin=>p(205)(17),clock=>clock,reset=>reset,s=>p(264)(17),cout=>p(265)(18));
FA_ff_8568:FAff port map(x=>p(203)(18),y=>p(204)(18),Cin=>p(205)(18),clock=>clock,reset=>reset,s=>p(264)(18),cout=>p(265)(19));
FA_ff_8569:FAff port map(x=>p(203)(19),y=>p(204)(19),Cin=>p(205)(19),clock=>clock,reset=>reset,s=>p(264)(19),cout=>p(265)(20));
FA_ff_8570:FAff port map(x=>p(203)(20),y=>p(204)(20),Cin=>p(205)(20),clock=>clock,reset=>reset,s=>p(264)(20),cout=>p(265)(21));
FA_ff_8571:FAff port map(x=>p(203)(21),y=>p(204)(21),Cin=>p(205)(21),clock=>clock,reset=>reset,s=>p(264)(21),cout=>p(265)(22));
FA_ff_8572:FAff port map(x=>p(203)(22),y=>p(204)(22),Cin=>p(205)(22),clock=>clock,reset=>reset,s=>p(264)(22),cout=>p(265)(23));
FA_ff_8573:FAff port map(x=>p(203)(23),y=>p(204)(23),Cin=>p(205)(23),clock=>clock,reset=>reset,s=>p(264)(23),cout=>p(265)(24));
FA_ff_8574:FAff port map(x=>p(203)(24),y=>p(204)(24),Cin=>p(205)(24),clock=>clock,reset=>reset,s=>p(264)(24),cout=>p(265)(25));
FA_ff_8575:FAff port map(x=>p(203)(25),y=>p(204)(25),Cin=>p(205)(25),clock=>clock,reset=>reset,s=>p(264)(25),cout=>p(265)(26));
FA_ff_8576:FAff port map(x=>p(203)(26),y=>p(204)(26),Cin=>p(205)(26),clock=>clock,reset=>reset,s=>p(264)(26),cout=>p(265)(27));
FA_ff_8577:FAff port map(x=>p(203)(27),y=>p(204)(27),Cin=>p(205)(27),clock=>clock,reset=>reset,s=>p(264)(27),cout=>p(265)(28));
FA_ff_8578:FAff port map(x=>p(203)(28),y=>p(204)(28),Cin=>p(205)(28),clock=>clock,reset=>reset,s=>p(264)(28),cout=>p(265)(29));
FA_ff_8579:FAff port map(x=>p(203)(29),y=>p(204)(29),Cin=>p(205)(29),clock=>clock,reset=>reset,s=>p(264)(29),cout=>p(265)(30));
FA_ff_8580:FAff port map(x=>p(203)(30),y=>p(204)(30),Cin=>p(205)(30),clock=>clock,reset=>reset,s=>p(264)(30),cout=>p(265)(31));
FA_ff_8581:FAff port map(x=>p(203)(31),y=>p(204)(31),Cin=>p(205)(31),clock=>clock,reset=>reset,s=>p(264)(31),cout=>p(265)(32));
FA_ff_8582:FAff port map(x=>p(203)(32),y=>p(204)(32),Cin=>p(205)(32),clock=>clock,reset=>reset,s=>p(264)(32),cout=>p(265)(33));
FA_ff_8583:FAff port map(x=>p(203)(33),y=>p(204)(33),Cin=>p(205)(33),clock=>clock,reset=>reset,s=>p(264)(33),cout=>p(265)(34));
FA_ff_8584:FAff port map(x=>p(203)(34),y=>p(204)(34),Cin=>p(205)(34),clock=>clock,reset=>reset,s=>p(264)(34),cout=>p(265)(35));
FA_ff_8585:FAff port map(x=>p(203)(35),y=>p(204)(35),Cin=>p(205)(35),clock=>clock,reset=>reset,s=>p(264)(35),cout=>p(265)(36));
FA_ff_8586:FAff port map(x=>p(203)(36),y=>p(204)(36),Cin=>p(205)(36),clock=>clock,reset=>reset,s=>p(264)(36),cout=>p(265)(37));
FA_ff_8587:FAff port map(x=>p(203)(37),y=>p(204)(37),Cin=>p(205)(37),clock=>clock,reset=>reset,s=>p(264)(37),cout=>p(265)(38));
FA_ff_8588:FAff port map(x=>p(203)(38),y=>p(204)(38),Cin=>p(205)(38),clock=>clock,reset=>reset,s=>p(264)(38),cout=>p(265)(39));
FA_ff_8589:FAff port map(x=>p(203)(39),y=>p(204)(39),Cin=>p(205)(39),clock=>clock,reset=>reset,s=>p(264)(39),cout=>p(265)(40));
FA_ff_8590:FAff port map(x=>p(203)(40),y=>p(204)(40),Cin=>p(205)(40),clock=>clock,reset=>reset,s=>p(264)(40),cout=>p(265)(41));
FA_ff_8591:FAff port map(x=>p(203)(41),y=>p(204)(41),Cin=>p(205)(41),clock=>clock,reset=>reset,s=>p(264)(41),cout=>p(265)(42));
FA_ff_8592:FAff port map(x=>p(203)(42),y=>p(204)(42),Cin=>p(205)(42),clock=>clock,reset=>reset,s=>p(264)(42),cout=>p(265)(43));
FA_ff_8593:FAff port map(x=>p(203)(43),y=>p(204)(43),Cin=>p(205)(43),clock=>clock,reset=>reset,s=>p(264)(43),cout=>p(265)(44));
FA_ff_8594:FAff port map(x=>p(203)(44),y=>p(204)(44),Cin=>p(205)(44),clock=>clock,reset=>reset,s=>p(264)(44),cout=>p(265)(45));
FA_ff_8595:FAff port map(x=>p(203)(45),y=>p(204)(45),Cin=>p(205)(45),clock=>clock,reset=>reset,s=>p(264)(45),cout=>p(265)(46));
FA_ff_8596:FAff port map(x=>p(203)(46),y=>p(204)(46),Cin=>p(205)(46),clock=>clock,reset=>reset,s=>p(264)(46),cout=>p(265)(47));
FA_ff_8597:FAff port map(x=>p(203)(47),y=>p(204)(47),Cin=>p(205)(47),clock=>clock,reset=>reset,s=>p(264)(47),cout=>p(265)(48));
FA_ff_8598:FAff port map(x=>p(203)(48),y=>p(204)(48),Cin=>p(205)(48),clock=>clock,reset=>reset,s=>p(264)(48),cout=>p(265)(49));
FA_ff_8599:FAff port map(x=>p(203)(49),y=>p(204)(49),Cin=>p(205)(49),clock=>clock,reset=>reset,s=>p(264)(49),cout=>p(265)(50));
FA_ff_8600:FAff port map(x=>p(203)(50),y=>p(204)(50),Cin=>p(205)(50),clock=>clock,reset=>reset,s=>p(264)(50),cout=>p(265)(51));
FA_ff_8601:FAff port map(x=>p(203)(51),y=>p(204)(51),Cin=>p(205)(51),clock=>clock,reset=>reset,s=>p(264)(51),cout=>p(265)(52));
FA_ff_8602:FAff port map(x=>p(203)(52),y=>p(204)(52),Cin=>p(205)(52),clock=>clock,reset=>reset,s=>p(264)(52),cout=>p(265)(53));
FA_ff_8603:FAff port map(x=>p(203)(53),y=>p(204)(53),Cin=>p(205)(53),clock=>clock,reset=>reset,s=>p(264)(53),cout=>p(265)(54));
FA_ff_8604:FAff port map(x=>p(203)(54),y=>p(204)(54),Cin=>p(205)(54),clock=>clock,reset=>reset,s=>p(264)(54),cout=>p(265)(55));
FA_ff_8605:FAff port map(x=>p(203)(55),y=>p(204)(55),Cin=>p(205)(55),clock=>clock,reset=>reset,s=>p(264)(55),cout=>p(265)(56));
FA_ff_8606:FAff port map(x=>p(203)(56),y=>p(204)(56),Cin=>p(205)(56),clock=>clock,reset=>reset,s=>p(264)(56),cout=>p(265)(57));
FA_ff_8607:FAff port map(x=>p(203)(57),y=>p(204)(57),Cin=>p(205)(57),clock=>clock,reset=>reset,s=>p(264)(57),cout=>p(265)(58));
FA_ff_8608:FAff port map(x=>p(203)(58),y=>p(204)(58),Cin=>p(205)(58),clock=>clock,reset=>reset,s=>p(264)(58),cout=>p(265)(59));
FA_ff_8609:FAff port map(x=>p(203)(59),y=>p(204)(59),Cin=>p(205)(59),clock=>clock,reset=>reset,s=>p(264)(59),cout=>p(265)(60));
FA_ff_8610:FAff port map(x=>p(203)(60),y=>p(204)(60),Cin=>p(205)(60),clock=>clock,reset=>reset,s=>p(264)(60),cout=>p(265)(61));
FA_ff_8611:FAff port map(x=>p(203)(61),y=>p(204)(61),Cin=>p(205)(61),clock=>clock,reset=>reset,s=>p(264)(61),cout=>p(265)(62));
FA_ff_8612:FAff port map(x=>p(203)(62),y=>p(204)(62),Cin=>p(205)(62),clock=>clock,reset=>reset,s=>p(264)(62),cout=>p(265)(63));
FA_ff_8613:FAff port map(x=>p(203)(63),y=>p(204)(63),Cin=>p(205)(63),clock=>clock,reset=>reset,s=>p(264)(63),cout=>p(265)(64));
FA_ff_8614:FAff port map(x=>p(203)(64),y=>p(204)(64),Cin=>p(205)(64),clock=>clock,reset=>reset,s=>p(264)(64),cout=>p(265)(65));
FA_ff_8615:FAff port map(x=>p(203)(65),y=>p(204)(65),Cin=>p(205)(65),clock=>clock,reset=>reset,s=>p(264)(65),cout=>p(265)(66));
FA_ff_8616:FAff port map(x=>p(203)(66),y=>p(204)(66),Cin=>p(205)(66),clock=>clock,reset=>reset,s=>p(264)(66),cout=>p(265)(67));
FA_ff_8617:FAff port map(x=>p(203)(67),y=>p(204)(67),Cin=>p(205)(67),clock=>clock,reset=>reset,s=>p(264)(67),cout=>p(265)(68));
FA_ff_8618:FAff port map(x=>p(203)(68),y=>p(204)(68),Cin=>p(205)(68),clock=>clock,reset=>reset,s=>p(264)(68),cout=>p(265)(69));
FA_ff_8619:FAff port map(x=>p(203)(69),y=>p(204)(69),Cin=>p(205)(69),clock=>clock,reset=>reset,s=>p(264)(69),cout=>p(265)(70));
FA_ff_8620:FAff port map(x=>p(203)(70),y=>p(204)(70),Cin=>p(205)(70),clock=>clock,reset=>reset,s=>p(264)(70),cout=>p(265)(71));
FA_ff_8621:FAff port map(x=>p(203)(71),y=>p(204)(71),Cin=>p(205)(71),clock=>clock,reset=>reset,s=>p(264)(71),cout=>p(265)(72));
FA_ff_8622:FAff port map(x=>p(203)(72),y=>p(204)(72),Cin=>p(205)(72),clock=>clock,reset=>reset,s=>p(264)(72),cout=>p(265)(73));
FA_ff_8623:FAff port map(x=>p(203)(73),y=>p(204)(73),Cin=>p(205)(73),clock=>clock,reset=>reset,s=>p(264)(73),cout=>p(265)(74));
FA_ff_8624:FAff port map(x=>p(203)(74),y=>p(204)(74),Cin=>p(205)(74),clock=>clock,reset=>reset,s=>p(264)(74),cout=>p(265)(75));
FA_ff_8625:FAff port map(x=>p(203)(75),y=>p(204)(75),Cin=>p(205)(75),clock=>clock,reset=>reset,s=>p(264)(75),cout=>p(265)(76));
FA_ff_8626:FAff port map(x=>p(203)(76),y=>p(204)(76),Cin=>p(205)(76),clock=>clock,reset=>reset,s=>p(264)(76),cout=>p(265)(77));
FA_ff_8627:FAff port map(x=>p(203)(77),y=>p(204)(77),Cin=>p(205)(77),clock=>clock,reset=>reset,s=>p(264)(77),cout=>p(265)(78));
FA_ff_8628:FAff port map(x=>p(203)(78),y=>p(204)(78),Cin=>p(205)(78),clock=>clock,reset=>reset,s=>p(264)(78),cout=>p(265)(79));
FA_ff_8629:FAff port map(x=>p(203)(79),y=>p(204)(79),Cin=>p(205)(79),clock=>clock,reset=>reset,s=>p(264)(79),cout=>p(265)(80));
FA_ff_8630:FAff port map(x=>p(203)(80),y=>p(204)(80),Cin=>p(205)(80),clock=>clock,reset=>reset,s=>p(264)(80),cout=>p(265)(81));
FA_ff_8631:FAff port map(x=>p(203)(81),y=>p(204)(81),Cin=>p(205)(81),clock=>clock,reset=>reset,s=>p(264)(81),cout=>p(265)(82));
FA_ff_8632:FAff port map(x=>p(203)(82),y=>p(204)(82),Cin=>p(205)(82),clock=>clock,reset=>reset,s=>p(264)(82),cout=>p(265)(83));
FA_ff_8633:FAff port map(x=>p(203)(83),y=>p(204)(83),Cin=>p(205)(83),clock=>clock,reset=>reset,s=>p(264)(83),cout=>p(265)(84));
FA_ff_8634:FAff port map(x=>p(203)(84),y=>p(204)(84),Cin=>p(205)(84),clock=>clock,reset=>reset,s=>p(264)(84),cout=>p(265)(85));
FA_ff_8635:FAff port map(x=>p(203)(85),y=>p(204)(85),Cin=>p(205)(85),clock=>clock,reset=>reset,s=>p(264)(85),cout=>p(265)(86));
FA_ff_8636:FAff port map(x=>p(203)(86),y=>p(204)(86),Cin=>p(205)(86),clock=>clock,reset=>reset,s=>p(264)(86),cout=>p(265)(87));
FA_ff_8637:FAff port map(x=>p(203)(87),y=>p(204)(87),Cin=>p(205)(87),clock=>clock,reset=>reset,s=>p(264)(87),cout=>p(265)(88));
FA_ff_8638:FAff port map(x=>p(203)(88),y=>p(204)(88),Cin=>p(205)(88),clock=>clock,reset=>reset,s=>p(264)(88),cout=>p(265)(89));
FA_ff_8639:FAff port map(x=>p(203)(89),y=>p(204)(89),Cin=>p(205)(89),clock=>clock,reset=>reset,s=>p(264)(89),cout=>p(265)(90));
FA_ff_8640:FAff port map(x=>p(203)(90),y=>p(204)(90),Cin=>p(205)(90),clock=>clock,reset=>reset,s=>p(264)(90),cout=>p(265)(91));
FA_ff_8641:FAff port map(x=>p(203)(91),y=>p(204)(91),Cin=>p(205)(91),clock=>clock,reset=>reset,s=>p(264)(91),cout=>p(265)(92));
FA_ff_8642:FAff port map(x=>p(203)(92),y=>p(204)(92),Cin=>p(205)(92),clock=>clock,reset=>reset,s=>p(264)(92),cout=>p(265)(93));
FA_ff_8643:FAff port map(x=>p(203)(93),y=>p(204)(93),Cin=>p(205)(93),clock=>clock,reset=>reset,s=>p(264)(93),cout=>p(265)(94));
FA_ff_8644:FAff port map(x=>p(203)(94),y=>p(204)(94),Cin=>p(205)(94),clock=>clock,reset=>reset,s=>p(264)(94),cout=>p(265)(95));
FA_ff_8645:FAff port map(x=>p(203)(95),y=>p(204)(95),Cin=>p(205)(95),clock=>clock,reset=>reset,s=>p(264)(95),cout=>p(265)(96));
FA_ff_8646:FAff port map(x=>p(203)(96),y=>p(204)(96),Cin=>p(205)(96),clock=>clock,reset=>reset,s=>p(264)(96),cout=>p(265)(97));
FA_ff_8647:FAff port map(x=>p(203)(97),y=>p(204)(97),Cin=>p(205)(97),clock=>clock,reset=>reset,s=>p(264)(97),cout=>p(265)(98));
FA_ff_8648:FAff port map(x=>p(203)(98),y=>p(204)(98),Cin=>p(205)(98),clock=>clock,reset=>reset,s=>p(264)(98),cout=>p(265)(99));
FA_ff_8649:FAff port map(x=>p(203)(99),y=>p(204)(99),Cin=>p(205)(99),clock=>clock,reset=>reset,s=>p(264)(99),cout=>p(265)(100));
FA_ff_8650:FAff port map(x=>p(203)(100),y=>p(204)(100),Cin=>p(205)(100),clock=>clock,reset=>reset,s=>p(264)(100),cout=>p(265)(101));
FA_ff_8651:FAff port map(x=>p(203)(101),y=>p(204)(101),Cin=>p(205)(101),clock=>clock,reset=>reset,s=>p(264)(101),cout=>p(265)(102));
FA_ff_8652:FAff port map(x=>p(203)(102),y=>p(204)(102),Cin=>p(205)(102),clock=>clock,reset=>reset,s=>p(264)(102),cout=>p(265)(103));
FA_ff_8653:FAff port map(x=>p(203)(103),y=>p(204)(103),Cin=>p(205)(103),clock=>clock,reset=>reset,s=>p(264)(103),cout=>p(265)(104));
FA_ff_8654:FAff port map(x=>p(203)(104),y=>p(204)(104),Cin=>p(205)(104),clock=>clock,reset=>reset,s=>p(264)(104),cout=>p(265)(105));
FA_ff_8655:FAff port map(x=>p(203)(105),y=>p(204)(105),Cin=>p(205)(105),clock=>clock,reset=>reset,s=>p(264)(105),cout=>p(265)(106));
FA_ff_8656:FAff port map(x=>p(203)(106),y=>p(204)(106),Cin=>p(205)(106),clock=>clock,reset=>reset,s=>p(264)(106),cout=>p(265)(107));
FA_ff_8657:FAff port map(x=>p(203)(107),y=>p(204)(107),Cin=>p(205)(107),clock=>clock,reset=>reset,s=>p(264)(107),cout=>p(265)(108));
FA_ff_8658:FAff port map(x=>p(203)(108),y=>p(204)(108),Cin=>p(205)(108),clock=>clock,reset=>reset,s=>p(264)(108),cout=>p(265)(109));
FA_ff_8659:FAff port map(x=>p(203)(109),y=>p(204)(109),Cin=>p(205)(109),clock=>clock,reset=>reset,s=>p(264)(109),cout=>p(265)(110));
FA_ff_8660:FAff port map(x=>p(203)(110),y=>p(204)(110),Cin=>p(205)(110),clock=>clock,reset=>reset,s=>p(264)(110),cout=>p(265)(111));
FA_ff_8661:FAff port map(x=>p(203)(111),y=>p(204)(111),Cin=>p(205)(111),clock=>clock,reset=>reset,s=>p(264)(111),cout=>p(265)(112));
FA_ff_8662:FAff port map(x=>p(203)(112),y=>p(204)(112),Cin=>p(205)(112),clock=>clock,reset=>reset,s=>p(264)(112),cout=>p(265)(113));
FA_ff_8663:FAff port map(x=>p(203)(113),y=>p(204)(113),Cin=>p(205)(113),clock=>clock,reset=>reset,s=>p(264)(113),cout=>p(265)(114));
FA_ff_8664:FAff port map(x=>p(203)(114),y=>p(204)(114),Cin=>p(205)(114),clock=>clock,reset=>reset,s=>p(264)(114),cout=>p(265)(115));
FA_ff_8665:FAff port map(x=>p(203)(115),y=>p(204)(115),Cin=>p(205)(115),clock=>clock,reset=>reset,s=>p(264)(115),cout=>p(265)(116));
FA_ff_8666:FAff port map(x=>p(203)(116),y=>p(204)(116),Cin=>p(205)(116),clock=>clock,reset=>reset,s=>p(264)(116),cout=>p(265)(117));
FA_ff_8667:FAff port map(x=>p(203)(117),y=>p(204)(117),Cin=>p(205)(117),clock=>clock,reset=>reset,s=>p(264)(117),cout=>p(265)(118));
FA_ff_8668:FAff port map(x=>p(203)(118),y=>p(204)(118),Cin=>p(205)(118),clock=>clock,reset=>reset,s=>p(264)(118),cout=>p(265)(119));
FA_ff_8669:FAff port map(x=>p(203)(119),y=>p(204)(119),Cin=>p(205)(119),clock=>clock,reset=>reset,s=>p(264)(119),cout=>p(265)(120));
FA_ff_8670:FAff port map(x=>p(203)(120),y=>p(204)(120),Cin=>p(205)(120),clock=>clock,reset=>reset,s=>p(264)(120),cout=>p(265)(121));
FA_ff_8671:FAff port map(x=>p(203)(121),y=>p(204)(121),Cin=>p(205)(121),clock=>clock,reset=>reset,s=>p(264)(121),cout=>p(265)(122));
FA_ff_8672:FAff port map(x=>p(203)(122),y=>p(204)(122),Cin=>p(205)(122),clock=>clock,reset=>reset,s=>p(264)(122),cout=>p(265)(123));
FA_ff_8673:FAff port map(x=>p(203)(123),y=>p(204)(123),Cin=>p(205)(123),clock=>clock,reset=>reset,s=>p(264)(123),cout=>p(265)(124));
FA_ff_8674:FAff port map(x=>p(203)(124),y=>p(204)(124),Cin=>p(205)(124),clock=>clock,reset=>reset,s=>p(264)(124),cout=>p(265)(125));
FA_ff_8675:FAff port map(x=>p(203)(125),y=>p(204)(125),Cin=>p(205)(125),clock=>clock,reset=>reset,s=>p(264)(125),cout=>p(265)(126));
FA_ff_8676:FAff port map(x=>p(203)(126),y=>p(204)(126),Cin=>p(205)(126),clock=>clock,reset=>reset,s=>p(264)(126),cout=>p(265)(127));
FA_ff_8677:FAff port map(x=>p(203)(127),y=>p(204)(127),Cin=>p(205)(127),clock=>clock,reset=>reset,s=>p(264)(127),cout=>p(265)(128));
HA_ff_25:HAff port map(x=>p(203)(128),y=>p(205)(128),clock=>clock,reset=>reset,s=>p(264)(128),c=>p(265)(129));
HA_ff_26:HAff port map(x=>p(206)(0),y=>p(208)(0),clock=>clock,reset=>reset,s=>p(266)(0),c=>p(267)(1));
FA_ff_8678:FAff port map(x=>p(206)(1),y=>p(207)(1),Cin=>p(208)(1),clock=>clock,reset=>reset,s=>p(266)(1),cout=>p(267)(2));
FA_ff_8679:FAff port map(x=>p(206)(2),y=>p(207)(2),Cin=>p(208)(2),clock=>clock,reset=>reset,s=>p(266)(2),cout=>p(267)(3));
FA_ff_8680:FAff port map(x=>p(206)(3),y=>p(207)(3),Cin=>p(208)(3),clock=>clock,reset=>reset,s=>p(266)(3),cout=>p(267)(4));
FA_ff_8681:FAff port map(x=>p(206)(4),y=>p(207)(4),Cin=>p(208)(4),clock=>clock,reset=>reset,s=>p(266)(4),cout=>p(267)(5));
FA_ff_8682:FAff port map(x=>p(206)(5),y=>p(207)(5),Cin=>p(208)(5),clock=>clock,reset=>reset,s=>p(266)(5),cout=>p(267)(6));
FA_ff_8683:FAff port map(x=>p(206)(6),y=>p(207)(6),Cin=>p(208)(6),clock=>clock,reset=>reset,s=>p(266)(6),cout=>p(267)(7));
FA_ff_8684:FAff port map(x=>p(206)(7),y=>p(207)(7),Cin=>p(208)(7),clock=>clock,reset=>reset,s=>p(266)(7),cout=>p(267)(8));
FA_ff_8685:FAff port map(x=>p(206)(8),y=>p(207)(8),Cin=>p(208)(8),clock=>clock,reset=>reset,s=>p(266)(8),cout=>p(267)(9));
FA_ff_8686:FAff port map(x=>p(206)(9),y=>p(207)(9),Cin=>p(208)(9),clock=>clock,reset=>reset,s=>p(266)(9),cout=>p(267)(10));
FA_ff_8687:FAff port map(x=>p(206)(10),y=>p(207)(10),Cin=>p(208)(10),clock=>clock,reset=>reset,s=>p(266)(10),cout=>p(267)(11));
FA_ff_8688:FAff port map(x=>p(206)(11),y=>p(207)(11),Cin=>p(208)(11),clock=>clock,reset=>reset,s=>p(266)(11),cout=>p(267)(12));
FA_ff_8689:FAff port map(x=>p(206)(12),y=>p(207)(12),Cin=>p(208)(12),clock=>clock,reset=>reset,s=>p(266)(12),cout=>p(267)(13));
FA_ff_8690:FAff port map(x=>p(206)(13),y=>p(207)(13),Cin=>p(208)(13),clock=>clock,reset=>reset,s=>p(266)(13),cout=>p(267)(14));
FA_ff_8691:FAff port map(x=>p(206)(14),y=>p(207)(14),Cin=>p(208)(14),clock=>clock,reset=>reset,s=>p(266)(14),cout=>p(267)(15));
FA_ff_8692:FAff port map(x=>p(206)(15),y=>p(207)(15),Cin=>p(208)(15),clock=>clock,reset=>reset,s=>p(266)(15),cout=>p(267)(16));
FA_ff_8693:FAff port map(x=>p(206)(16),y=>p(207)(16),Cin=>p(208)(16),clock=>clock,reset=>reset,s=>p(266)(16),cout=>p(267)(17));
FA_ff_8694:FAff port map(x=>p(206)(17),y=>p(207)(17),Cin=>p(208)(17),clock=>clock,reset=>reset,s=>p(266)(17),cout=>p(267)(18));
FA_ff_8695:FAff port map(x=>p(206)(18),y=>p(207)(18),Cin=>p(208)(18),clock=>clock,reset=>reset,s=>p(266)(18),cout=>p(267)(19));
FA_ff_8696:FAff port map(x=>p(206)(19),y=>p(207)(19),Cin=>p(208)(19),clock=>clock,reset=>reset,s=>p(266)(19),cout=>p(267)(20));
FA_ff_8697:FAff port map(x=>p(206)(20),y=>p(207)(20),Cin=>p(208)(20),clock=>clock,reset=>reset,s=>p(266)(20),cout=>p(267)(21));
FA_ff_8698:FAff port map(x=>p(206)(21),y=>p(207)(21),Cin=>p(208)(21),clock=>clock,reset=>reset,s=>p(266)(21),cout=>p(267)(22));
FA_ff_8699:FAff port map(x=>p(206)(22),y=>p(207)(22),Cin=>p(208)(22),clock=>clock,reset=>reset,s=>p(266)(22),cout=>p(267)(23));
FA_ff_8700:FAff port map(x=>p(206)(23),y=>p(207)(23),Cin=>p(208)(23),clock=>clock,reset=>reset,s=>p(266)(23),cout=>p(267)(24));
FA_ff_8701:FAff port map(x=>p(206)(24),y=>p(207)(24),Cin=>p(208)(24),clock=>clock,reset=>reset,s=>p(266)(24),cout=>p(267)(25));
FA_ff_8702:FAff port map(x=>p(206)(25),y=>p(207)(25),Cin=>p(208)(25),clock=>clock,reset=>reset,s=>p(266)(25),cout=>p(267)(26));
FA_ff_8703:FAff port map(x=>p(206)(26),y=>p(207)(26),Cin=>p(208)(26),clock=>clock,reset=>reset,s=>p(266)(26),cout=>p(267)(27));
FA_ff_8704:FAff port map(x=>p(206)(27),y=>p(207)(27),Cin=>p(208)(27),clock=>clock,reset=>reset,s=>p(266)(27),cout=>p(267)(28));
FA_ff_8705:FAff port map(x=>p(206)(28),y=>p(207)(28),Cin=>p(208)(28),clock=>clock,reset=>reset,s=>p(266)(28),cout=>p(267)(29));
FA_ff_8706:FAff port map(x=>p(206)(29),y=>p(207)(29),Cin=>p(208)(29),clock=>clock,reset=>reset,s=>p(266)(29),cout=>p(267)(30));
FA_ff_8707:FAff port map(x=>p(206)(30),y=>p(207)(30),Cin=>p(208)(30),clock=>clock,reset=>reset,s=>p(266)(30),cout=>p(267)(31));
FA_ff_8708:FAff port map(x=>p(206)(31),y=>p(207)(31),Cin=>p(208)(31),clock=>clock,reset=>reset,s=>p(266)(31),cout=>p(267)(32));
FA_ff_8709:FAff port map(x=>p(206)(32),y=>p(207)(32),Cin=>p(208)(32),clock=>clock,reset=>reset,s=>p(266)(32),cout=>p(267)(33));
FA_ff_8710:FAff port map(x=>p(206)(33),y=>p(207)(33),Cin=>p(208)(33),clock=>clock,reset=>reset,s=>p(266)(33),cout=>p(267)(34));
FA_ff_8711:FAff port map(x=>p(206)(34),y=>p(207)(34),Cin=>p(208)(34),clock=>clock,reset=>reset,s=>p(266)(34),cout=>p(267)(35));
FA_ff_8712:FAff port map(x=>p(206)(35),y=>p(207)(35),Cin=>p(208)(35),clock=>clock,reset=>reset,s=>p(266)(35),cout=>p(267)(36));
FA_ff_8713:FAff port map(x=>p(206)(36),y=>p(207)(36),Cin=>p(208)(36),clock=>clock,reset=>reset,s=>p(266)(36),cout=>p(267)(37));
FA_ff_8714:FAff port map(x=>p(206)(37),y=>p(207)(37),Cin=>p(208)(37),clock=>clock,reset=>reset,s=>p(266)(37),cout=>p(267)(38));
FA_ff_8715:FAff port map(x=>p(206)(38),y=>p(207)(38),Cin=>p(208)(38),clock=>clock,reset=>reset,s=>p(266)(38),cout=>p(267)(39));
FA_ff_8716:FAff port map(x=>p(206)(39),y=>p(207)(39),Cin=>p(208)(39),clock=>clock,reset=>reset,s=>p(266)(39),cout=>p(267)(40));
FA_ff_8717:FAff port map(x=>p(206)(40),y=>p(207)(40),Cin=>p(208)(40),clock=>clock,reset=>reset,s=>p(266)(40),cout=>p(267)(41));
FA_ff_8718:FAff port map(x=>p(206)(41),y=>p(207)(41),Cin=>p(208)(41),clock=>clock,reset=>reset,s=>p(266)(41),cout=>p(267)(42));
FA_ff_8719:FAff port map(x=>p(206)(42),y=>p(207)(42),Cin=>p(208)(42),clock=>clock,reset=>reset,s=>p(266)(42),cout=>p(267)(43));
FA_ff_8720:FAff port map(x=>p(206)(43),y=>p(207)(43),Cin=>p(208)(43),clock=>clock,reset=>reset,s=>p(266)(43),cout=>p(267)(44));
FA_ff_8721:FAff port map(x=>p(206)(44),y=>p(207)(44),Cin=>p(208)(44),clock=>clock,reset=>reset,s=>p(266)(44),cout=>p(267)(45));
FA_ff_8722:FAff port map(x=>p(206)(45),y=>p(207)(45),Cin=>p(208)(45),clock=>clock,reset=>reset,s=>p(266)(45),cout=>p(267)(46));
FA_ff_8723:FAff port map(x=>p(206)(46),y=>p(207)(46),Cin=>p(208)(46),clock=>clock,reset=>reset,s=>p(266)(46),cout=>p(267)(47));
FA_ff_8724:FAff port map(x=>p(206)(47),y=>p(207)(47),Cin=>p(208)(47),clock=>clock,reset=>reset,s=>p(266)(47),cout=>p(267)(48));
FA_ff_8725:FAff port map(x=>p(206)(48),y=>p(207)(48),Cin=>p(208)(48),clock=>clock,reset=>reset,s=>p(266)(48),cout=>p(267)(49));
FA_ff_8726:FAff port map(x=>p(206)(49),y=>p(207)(49),Cin=>p(208)(49),clock=>clock,reset=>reset,s=>p(266)(49),cout=>p(267)(50));
FA_ff_8727:FAff port map(x=>p(206)(50),y=>p(207)(50),Cin=>p(208)(50),clock=>clock,reset=>reset,s=>p(266)(50),cout=>p(267)(51));
FA_ff_8728:FAff port map(x=>p(206)(51),y=>p(207)(51),Cin=>p(208)(51),clock=>clock,reset=>reset,s=>p(266)(51),cout=>p(267)(52));
FA_ff_8729:FAff port map(x=>p(206)(52),y=>p(207)(52),Cin=>p(208)(52),clock=>clock,reset=>reset,s=>p(266)(52),cout=>p(267)(53));
FA_ff_8730:FAff port map(x=>p(206)(53),y=>p(207)(53),Cin=>p(208)(53),clock=>clock,reset=>reset,s=>p(266)(53),cout=>p(267)(54));
FA_ff_8731:FAff port map(x=>p(206)(54),y=>p(207)(54),Cin=>p(208)(54),clock=>clock,reset=>reset,s=>p(266)(54),cout=>p(267)(55));
FA_ff_8732:FAff port map(x=>p(206)(55),y=>p(207)(55),Cin=>p(208)(55),clock=>clock,reset=>reset,s=>p(266)(55),cout=>p(267)(56));
FA_ff_8733:FAff port map(x=>p(206)(56),y=>p(207)(56),Cin=>p(208)(56),clock=>clock,reset=>reset,s=>p(266)(56),cout=>p(267)(57));
FA_ff_8734:FAff port map(x=>p(206)(57),y=>p(207)(57),Cin=>p(208)(57),clock=>clock,reset=>reset,s=>p(266)(57),cout=>p(267)(58));
FA_ff_8735:FAff port map(x=>p(206)(58),y=>p(207)(58),Cin=>p(208)(58),clock=>clock,reset=>reset,s=>p(266)(58),cout=>p(267)(59));
FA_ff_8736:FAff port map(x=>p(206)(59),y=>p(207)(59),Cin=>p(208)(59),clock=>clock,reset=>reset,s=>p(266)(59),cout=>p(267)(60));
FA_ff_8737:FAff port map(x=>p(206)(60),y=>p(207)(60),Cin=>p(208)(60),clock=>clock,reset=>reset,s=>p(266)(60),cout=>p(267)(61));
FA_ff_8738:FAff port map(x=>p(206)(61),y=>p(207)(61),Cin=>p(208)(61),clock=>clock,reset=>reset,s=>p(266)(61),cout=>p(267)(62));
FA_ff_8739:FAff port map(x=>p(206)(62),y=>p(207)(62),Cin=>p(208)(62),clock=>clock,reset=>reset,s=>p(266)(62),cout=>p(267)(63));
FA_ff_8740:FAff port map(x=>p(206)(63),y=>p(207)(63),Cin=>p(208)(63),clock=>clock,reset=>reset,s=>p(266)(63),cout=>p(267)(64));
FA_ff_8741:FAff port map(x=>p(206)(64),y=>p(207)(64),Cin=>p(208)(64),clock=>clock,reset=>reset,s=>p(266)(64),cout=>p(267)(65));
FA_ff_8742:FAff port map(x=>p(206)(65),y=>p(207)(65),Cin=>p(208)(65),clock=>clock,reset=>reset,s=>p(266)(65),cout=>p(267)(66));
FA_ff_8743:FAff port map(x=>p(206)(66),y=>p(207)(66),Cin=>p(208)(66),clock=>clock,reset=>reset,s=>p(266)(66),cout=>p(267)(67));
FA_ff_8744:FAff port map(x=>p(206)(67),y=>p(207)(67),Cin=>p(208)(67),clock=>clock,reset=>reset,s=>p(266)(67),cout=>p(267)(68));
FA_ff_8745:FAff port map(x=>p(206)(68),y=>p(207)(68),Cin=>p(208)(68),clock=>clock,reset=>reset,s=>p(266)(68),cout=>p(267)(69));
FA_ff_8746:FAff port map(x=>p(206)(69),y=>p(207)(69),Cin=>p(208)(69),clock=>clock,reset=>reset,s=>p(266)(69),cout=>p(267)(70));
FA_ff_8747:FAff port map(x=>p(206)(70),y=>p(207)(70),Cin=>p(208)(70),clock=>clock,reset=>reset,s=>p(266)(70),cout=>p(267)(71));
FA_ff_8748:FAff port map(x=>p(206)(71),y=>p(207)(71),Cin=>p(208)(71),clock=>clock,reset=>reset,s=>p(266)(71),cout=>p(267)(72));
FA_ff_8749:FAff port map(x=>p(206)(72),y=>p(207)(72),Cin=>p(208)(72),clock=>clock,reset=>reset,s=>p(266)(72),cout=>p(267)(73));
FA_ff_8750:FAff port map(x=>p(206)(73),y=>p(207)(73),Cin=>p(208)(73),clock=>clock,reset=>reset,s=>p(266)(73),cout=>p(267)(74));
FA_ff_8751:FAff port map(x=>p(206)(74),y=>p(207)(74),Cin=>p(208)(74),clock=>clock,reset=>reset,s=>p(266)(74),cout=>p(267)(75));
FA_ff_8752:FAff port map(x=>p(206)(75),y=>p(207)(75),Cin=>p(208)(75),clock=>clock,reset=>reset,s=>p(266)(75),cout=>p(267)(76));
FA_ff_8753:FAff port map(x=>p(206)(76),y=>p(207)(76),Cin=>p(208)(76),clock=>clock,reset=>reset,s=>p(266)(76),cout=>p(267)(77));
FA_ff_8754:FAff port map(x=>p(206)(77),y=>p(207)(77),Cin=>p(208)(77),clock=>clock,reset=>reset,s=>p(266)(77),cout=>p(267)(78));
FA_ff_8755:FAff port map(x=>p(206)(78),y=>p(207)(78),Cin=>p(208)(78),clock=>clock,reset=>reset,s=>p(266)(78),cout=>p(267)(79));
FA_ff_8756:FAff port map(x=>p(206)(79),y=>p(207)(79),Cin=>p(208)(79),clock=>clock,reset=>reset,s=>p(266)(79),cout=>p(267)(80));
FA_ff_8757:FAff port map(x=>p(206)(80),y=>p(207)(80),Cin=>p(208)(80),clock=>clock,reset=>reset,s=>p(266)(80),cout=>p(267)(81));
FA_ff_8758:FAff port map(x=>p(206)(81),y=>p(207)(81),Cin=>p(208)(81),clock=>clock,reset=>reset,s=>p(266)(81),cout=>p(267)(82));
FA_ff_8759:FAff port map(x=>p(206)(82),y=>p(207)(82),Cin=>p(208)(82),clock=>clock,reset=>reset,s=>p(266)(82),cout=>p(267)(83));
FA_ff_8760:FAff port map(x=>p(206)(83),y=>p(207)(83),Cin=>p(208)(83),clock=>clock,reset=>reset,s=>p(266)(83),cout=>p(267)(84));
FA_ff_8761:FAff port map(x=>p(206)(84),y=>p(207)(84),Cin=>p(208)(84),clock=>clock,reset=>reset,s=>p(266)(84),cout=>p(267)(85));
FA_ff_8762:FAff port map(x=>p(206)(85),y=>p(207)(85),Cin=>p(208)(85),clock=>clock,reset=>reset,s=>p(266)(85),cout=>p(267)(86));
FA_ff_8763:FAff port map(x=>p(206)(86),y=>p(207)(86),Cin=>p(208)(86),clock=>clock,reset=>reset,s=>p(266)(86),cout=>p(267)(87));
FA_ff_8764:FAff port map(x=>p(206)(87),y=>p(207)(87),Cin=>p(208)(87),clock=>clock,reset=>reset,s=>p(266)(87),cout=>p(267)(88));
FA_ff_8765:FAff port map(x=>p(206)(88),y=>p(207)(88),Cin=>p(208)(88),clock=>clock,reset=>reset,s=>p(266)(88),cout=>p(267)(89));
FA_ff_8766:FAff port map(x=>p(206)(89),y=>p(207)(89),Cin=>p(208)(89),clock=>clock,reset=>reset,s=>p(266)(89),cout=>p(267)(90));
FA_ff_8767:FAff port map(x=>p(206)(90),y=>p(207)(90),Cin=>p(208)(90),clock=>clock,reset=>reset,s=>p(266)(90),cout=>p(267)(91));
FA_ff_8768:FAff port map(x=>p(206)(91),y=>p(207)(91),Cin=>p(208)(91),clock=>clock,reset=>reset,s=>p(266)(91),cout=>p(267)(92));
FA_ff_8769:FAff port map(x=>p(206)(92),y=>p(207)(92),Cin=>p(208)(92),clock=>clock,reset=>reset,s=>p(266)(92),cout=>p(267)(93));
FA_ff_8770:FAff port map(x=>p(206)(93),y=>p(207)(93),Cin=>p(208)(93),clock=>clock,reset=>reset,s=>p(266)(93),cout=>p(267)(94));
FA_ff_8771:FAff port map(x=>p(206)(94),y=>p(207)(94),Cin=>p(208)(94),clock=>clock,reset=>reset,s=>p(266)(94),cout=>p(267)(95));
FA_ff_8772:FAff port map(x=>p(206)(95),y=>p(207)(95),Cin=>p(208)(95),clock=>clock,reset=>reset,s=>p(266)(95),cout=>p(267)(96));
FA_ff_8773:FAff port map(x=>p(206)(96),y=>p(207)(96),Cin=>p(208)(96),clock=>clock,reset=>reset,s=>p(266)(96),cout=>p(267)(97));
FA_ff_8774:FAff port map(x=>p(206)(97),y=>p(207)(97),Cin=>p(208)(97),clock=>clock,reset=>reset,s=>p(266)(97),cout=>p(267)(98));
FA_ff_8775:FAff port map(x=>p(206)(98),y=>p(207)(98),Cin=>p(208)(98),clock=>clock,reset=>reset,s=>p(266)(98),cout=>p(267)(99));
FA_ff_8776:FAff port map(x=>p(206)(99),y=>p(207)(99),Cin=>p(208)(99),clock=>clock,reset=>reset,s=>p(266)(99),cout=>p(267)(100));
FA_ff_8777:FAff port map(x=>p(206)(100),y=>p(207)(100),Cin=>p(208)(100),clock=>clock,reset=>reset,s=>p(266)(100),cout=>p(267)(101));
FA_ff_8778:FAff port map(x=>p(206)(101),y=>p(207)(101),Cin=>p(208)(101),clock=>clock,reset=>reset,s=>p(266)(101),cout=>p(267)(102));
FA_ff_8779:FAff port map(x=>p(206)(102),y=>p(207)(102),Cin=>p(208)(102),clock=>clock,reset=>reset,s=>p(266)(102),cout=>p(267)(103));
FA_ff_8780:FAff port map(x=>p(206)(103),y=>p(207)(103),Cin=>p(208)(103),clock=>clock,reset=>reset,s=>p(266)(103),cout=>p(267)(104));
FA_ff_8781:FAff port map(x=>p(206)(104),y=>p(207)(104),Cin=>p(208)(104),clock=>clock,reset=>reset,s=>p(266)(104),cout=>p(267)(105));
FA_ff_8782:FAff port map(x=>p(206)(105),y=>p(207)(105),Cin=>p(208)(105),clock=>clock,reset=>reset,s=>p(266)(105),cout=>p(267)(106));
FA_ff_8783:FAff port map(x=>p(206)(106),y=>p(207)(106),Cin=>p(208)(106),clock=>clock,reset=>reset,s=>p(266)(106),cout=>p(267)(107));
FA_ff_8784:FAff port map(x=>p(206)(107),y=>p(207)(107),Cin=>p(208)(107),clock=>clock,reset=>reset,s=>p(266)(107),cout=>p(267)(108));
FA_ff_8785:FAff port map(x=>p(206)(108),y=>p(207)(108),Cin=>p(208)(108),clock=>clock,reset=>reset,s=>p(266)(108),cout=>p(267)(109));
FA_ff_8786:FAff port map(x=>p(206)(109),y=>p(207)(109),Cin=>p(208)(109),clock=>clock,reset=>reset,s=>p(266)(109),cout=>p(267)(110));
FA_ff_8787:FAff port map(x=>p(206)(110),y=>p(207)(110),Cin=>p(208)(110),clock=>clock,reset=>reset,s=>p(266)(110),cout=>p(267)(111));
FA_ff_8788:FAff port map(x=>p(206)(111),y=>p(207)(111),Cin=>p(208)(111),clock=>clock,reset=>reset,s=>p(266)(111),cout=>p(267)(112));
FA_ff_8789:FAff port map(x=>p(206)(112),y=>p(207)(112),Cin=>p(208)(112),clock=>clock,reset=>reset,s=>p(266)(112),cout=>p(267)(113));
FA_ff_8790:FAff port map(x=>p(206)(113),y=>p(207)(113),Cin=>p(208)(113),clock=>clock,reset=>reset,s=>p(266)(113),cout=>p(267)(114));
FA_ff_8791:FAff port map(x=>p(206)(114),y=>p(207)(114),Cin=>p(208)(114),clock=>clock,reset=>reset,s=>p(266)(114),cout=>p(267)(115));
FA_ff_8792:FAff port map(x=>p(206)(115),y=>p(207)(115),Cin=>p(208)(115),clock=>clock,reset=>reset,s=>p(266)(115),cout=>p(267)(116));
FA_ff_8793:FAff port map(x=>p(206)(116),y=>p(207)(116),Cin=>p(208)(116),clock=>clock,reset=>reset,s=>p(266)(116),cout=>p(267)(117));
FA_ff_8794:FAff port map(x=>p(206)(117),y=>p(207)(117),Cin=>p(208)(117),clock=>clock,reset=>reset,s=>p(266)(117),cout=>p(267)(118));
FA_ff_8795:FAff port map(x=>p(206)(118),y=>p(207)(118),Cin=>p(208)(118),clock=>clock,reset=>reset,s=>p(266)(118),cout=>p(267)(119));
FA_ff_8796:FAff port map(x=>p(206)(119),y=>p(207)(119),Cin=>p(208)(119),clock=>clock,reset=>reset,s=>p(266)(119),cout=>p(267)(120));
FA_ff_8797:FAff port map(x=>p(206)(120),y=>p(207)(120),Cin=>p(208)(120),clock=>clock,reset=>reset,s=>p(266)(120),cout=>p(267)(121));
FA_ff_8798:FAff port map(x=>p(206)(121),y=>p(207)(121),Cin=>p(208)(121),clock=>clock,reset=>reset,s=>p(266)(121),cout=>p(267)(122));
FA_ff_8799:FAff port map(x=>p(206)(122),y=>p(207)(122),Cin=>p(208)(122),clock=>clock,reset=>reset,s=>p(266)(122),cout=>p(267)(123));
FA_ff_8800:FAff port map(x=>p(206)(123),y=>p(207)(123),Cin=>p(208)(123),clock=>clock,reset=>reset,s=>p(266)(123),cout=>p(267)(124));
FA_ff_8801:FAff port map(x=>p(206)(124),y=>p(207)(124),Cin=>p(208)(124),clock=>clock,reset=>reset,s=>p(266)(124),cout=>p(267)(125));
FA_ff_8802:FAff port map(x=>p(206)(125),y=>p(207)(125),Cin=>p(208)(125),clock=>clock,reset=>reset,s=>p(266)(125),cout=>p(267)(126));
FA_ff_8803:FAff port map(x=>p(206)(126),y=>p(207)(126),Cin=>p(208)(126),clock=>clock,reset=>reset,s=>p(266)(126),cout=>p(267)(127));
FA_ff_8804:FAff port map(x=>p(206)(127),y=>p(207)(127),Cin=>p(208)(127),clock=>clock,reset=>reset,s=>p(266)(127),cout=>p(267)(128));
p(266)(128)<=p(207)(128);
p(268)(0)<=p(210)(0);
FA_ff_8805:FAff port map(x=>p(209)(1),y=>p(210)(1),Cin=>p(211)(1),clock=>clock,reset=>reset,s=>p(268)(1),cout=>p(269)(2));
FA_ff_8806:FAff port map(x=>p(209)(2),y=>p(210)(2),Cin=>p(211)(2),clock=>clock,reset=>reset,s=>p(268)(2),cout=>p(269)(3));
FA_ff_8807:FAff port map(x=>p(209)(3),y=>p(210)(3),Cin=>p(211)(3),clock=>clock,reset=>reset,s=>p(268)(3),cout=>p(269)(4));
FA_ff_8808:FAff port map(x=>p(209)(4),y=>p(210)(4),Cin=>p(211)(4),clock=>clock,reset=>reset,s=>p(268)(4),cout=>p(269)(5));
FA_ff_8809:FAff port map(x=>p(209)(5),y=>p(210)(5),Cin=>p(211)(5),clock=>clock,reset=>reset,s=>p(268)(5),cout=>p(269)(6));
FA_ff_8810:FAff port map(x=>p(209)(6),y=>p(210)(6),Cin=>p(211)(6),clock=>clock,reset=>reset,s=>p(268)(6),cout=>p(269)(7));
FA_ff_8811:FAff port map(x=>p(209)(7),y=>p(210)(7),Cin=>p(211)(7),clock=>clock,reset=>reset,s=>p(268)(7),cout=>p(269)(8));
FA_ff_8812:FAff port map(x=>p(209)(8),y=>p(210)(8),Cin=>p(211)(8),clock=>clock,reset=>reset,s=>p(268)(8),cout=>p(269)(9));
FA_ff_8813:FAff port map(x=>p(209)(9),y=>p(210)(9),Cin=>p(211)(9),clock=>clock,reset=>reset,s=>p(268)(9),cout=>p(269)(10));
FA_ff_8814:FAff port map(x=>p(209)(10),y=>p(210)(10),Cin=>p(211)(10),clock=>clock,reset=>reset,s=>p(268)(10),cout=>p(269)(11));
FA_ff_8815:FAff port map(x=>p(209)(11),y=>p(210)(11),Cin=>p(211)(11),clock=>clock,reset=>reset,s=>p(268)(11),cout=>p(269)(12));
FA_ff_8816:FAff port map(x=>p(209)(12),y=>p(210)(12),Cin=>p(211)(12),clock=>clock,reset=>reset,s=>p(268)(12),cout=>p(269)(13));
FA_ff_8817:FAff port map(x=>p(209)(13),y=>p(210)(13),Cin=>p(211)(13),clock=>clock,reset=>reset,s=>p(268)(13),cout=>p(269)(14));
FA_ff_8818:FAff port map(x=>p(209)(14),y=>p(210)(14),Cin=>p(211)(14),clock=>clock,reset=>reset,s=>p(268)(14),cout=>p(269)(15));
FA_ff_8819:FAff port map(x=>p(209)(15),y=>p(210)(15),Cin=>p(211)(15),clock=>clock,reset=>reset,s=>p(268)(15),cout=>p(269)(16));
FA_ff_8820:FAff port map(x=>p(209)(16),y=>p(210)(16),Cin=>p(211)(16),clock=>clock,reset=>reset,s=>p(268)(16),cout=>p(269)(17));
FA_ff_8821:FAff port map(x=>p(209)(17),y=>p(210)(17),Cin=>p(211)(17),clock=>clock,reset=>reset,s=>p(268)(17),cout=>p(269)(18));
FA_ff_8822:FAff port map(x=>p(209)(18),y=>p(210)(18),Cin=>p(211)(18),clock=>clock,reset=>reset,s=>p(268)(18),cout=>p(269)(19));
FA_ff_8823:FAff port map(x=>p(209)(19),y=>p(210)(19),Cin=>p(211)(19),clock=>clock,reset=>reset,s=>p(268)(19),cout=>p(269)(20));
FA_ff_8824:FAff port map(x=>p(209)(20),y=>p(210)(20),Cin=>p(211)(20),clock=>clock,reset=>reset,s=>p(268)(20),cout=>p(269)(21));
FA_ff_8825:FAff port map(x=>p(209)(21),y=>p(210)(21),Cin=>p(211)(21),clock=>clock,reset=>reset,s=>p(268)(21),cout=>p(269)(22));
FA_ff_8826:FAff port map(x=>p(209)(22),y=>p(210)(22),Cin=>p(211)(22),clock=>clock,reset=>reset,s=>p(268)(22),cout=>p(269)(23));
FA_ff_8827:FAff port map(x=>p(209)(23),y=>p(210)(23),Cin=>p(211)(23),clock=>clock,reset=>reset,s=>p(268)(23),cout=>p(269)(24));
FA_ff_8828:FAff port map(x=>p(209)(24),y=>p(210)(24),Cin=>p(211)(24),clock=>clock,reset=>reset,s=>p(268)(24),cout=>p(269)(25));
FA_ff_8829:FAff port map(x=>p(209)(25),y=>p(210)(25),Cin=>p(211)(25),clock=>clock,reset=>reset,s=>p(268)(25),cout=>p(269)(26));
FA_ff_8830:FAff port map(x=>p(209)(26),y=>p(210)(26),Cin=>p(211)(26),clock=>clock,reset=>reset,s=>p(268)(26),cout=>p(269)(27));
FA_ff_8831:FAff port map(x=>p(209)(27),y=>p(210)(27),Cin=>p(211)(27),clock=>clock,reset=>reset,s=>p(268)(27),cout=>p(269)(28));
FA_ff_8832:FAff port map(x=>p(209)(28),y=>p(210)(28),Cin=>p(211)(28),clock=>clock,reset=>reset,s=>p(268)(28),cout=>p(269)(29));
FA_ff_8833:FAff port map(x=>p(209)(29),y=>p(210)(29),Cin=>p(211)(29),clock=>clock,reset=>reset,s=>p(268)(29),cout=>p(269)(30));
FA_ff_8834:FAff port map(x=>p(209)(30),y=>p(210)(30),Cin=>p(211)(30),clock=>clock,reset=>reset,s=>p(268)(30),cout=>p(269)(31));
FA_ff_8835:FAff port map(x=>p(209)(31),y=>p(210)(31),Cin=>p(211)(31),clock=>clock,reset=>reset,s=>p(268)(31),cout=>p(269)(32));
FA_ff_8836:FAff port map(x=>p(209)(32),y=>p(210)(32),Cin=>p(211)(32),clock=>clock,reset=>reset,s=>p(268)(32),cout=>p(269)(33));
FA_ff_8837:FAff port map(x=>p(209)(33),y=>p(210)(33),Cin=>p(211)(33),clock=>clock,reset=>reset,s=>p(268)(33),cout=>p(269)(34));
FA_ff_8838:FAff port map(x=>p(209)(34),y=>p(210)(34),Cin=>p(211)(34),clock=>clock,reset=>reset,s=>p(268)(34),cout=>p(269)(35));
FA_ff_8839:FAff port map(x=>p(209)(35),y=>p(210)(35),Cin=>p(211)(35),clock=>clock,reset=>reset,s=>p(268)(35),cout=>p(269)(36));
FA_ff_8840:FAff port map(x=>p(209)(36),y=>p(210)(36),Cin=>p(211)(36),clock=>clock,reset=>reset,s=>p(268)(36),cout=>p(269)(37));
FA_ff_8841:FAff port map(x=>p(209)(37),y=>p(210)(37),Cin=>p(211)(37),clock=>clock,reset=>reset,s=>p(268)(37),cout=>p(269)(38));
FA_ff_8842:FAff port map(x=>p(209)(38),y=>p(210)(38),Cin=>p(211)(38),clock=>clock,reset=>reset,s=>p(268)(38),cout=>p(269)(39));
FA_ff_8843:FAff port map(x=>p(209)(39),y=>p(210)(39),Cin=>p(211)(39),clock=>clock,reset=>reset,s=>p(268)(39),cout=>p(269)(40));
FA_ff_8844:FAff port map(x=>p(209)(40),y=>p(210)(40),Cin=>p(211)(40),clock=>clock,reset=>reset,s=>p(268)(40),cout=>p(269)(41));
FA_ff_8845:FAff port map(x=>p(209)(41),y=>p(210)(41),Cin=>p(211)(41),clock=>clock,reset=>reset,s=>p(268)(41),cout=>p(269)(42));
FA_ff_8846:FAff port map(x=>p(209)(42),y=>p(210)(42),Cin=>p(211)(42),clock=>clock,reset=>reset,s=>p(268)(42),cout=>p(269)(43));
FA_ff_8847:FAff port map(x=>p(209)(43),y=>p(210)(43),Cin=>p(211)(43),clock=>clock,reset=>reset,s=>p(268)(43),cout=>p(269)(44));
FA_ff_8848:FAff port map(x=>p(209)(44),y=>p(210)(44),Cin=>p(211)(44),clock=>clock,reset=>reset,s=>p(268)(44),cout=>p(269)(45));
FA_ff_8849:FAff port map(x=>p(209)(45),y=>p(210)(45),Cin=>p(211)(45),clock=>clock,reset=>reset,s=>p(268)(45),cout=>p(269)(46));
FA_ff_8850:FAff port map(x=>p(209)(46),y=>p(210)(46),Cin=>p(211)(46),clock=>clock,reset=>reset,s=>p(268)(46),cout=>p(269)(47));
FA_ff_8851:FAff port map(x=>p(209)(47),y=>p(210)(47),Cin=>p(211)(47),clock=>clock,reset=>reset,s=>p(268)(47),cout=>p(269)(48));
FA_ff_8852:FAff port map(x=>p(209)(48),y=>p(210)(48),Cin=>p(211)(48),clock=>clock,reset=>reset,s=>p(268)(48),cout=>p(269)(49));
FA_ff_8853:FAff port map(x=>p(209)(49),y=>p(210)(49),Cin=>p(211)(49),clock=>clock,reset=>reset,s=>p(268)(49),cout=>p(269)(50));
FA_ff_8854:FAff port map(x=>p(209)(50),y=>p(210)(50),Cin=>p(211)(50),clock=>clock,reset=>reset,s=>p(268)(50),cout=>p(269)(51));
FA_ff_8855:FAff port map(x=>p(209)(51),y=>p(210)(51),Cin=>p(211)(51),clock=>clock,reset=>reset,s=>p(268)(51),cout=>p(269)(52));
FA_ff_8856:FAff port map(x=>p(209)(52),y=>p(210)(52),Cin=>p(211)(52),clock=>clock,reset=>reset,s=>p(268)(52),cout=>p(269)(53));
FA_ff_8857:FAff port map(x=>p(209)(53),y=>p(210)(53),Cin=>p(211)(53),clock=>clock,reset=>reset,s=>p(268)(53),cout=>p(269)(54));
FA_ff_8858:FAff port map(x=>p(209)(54),y=>p(210)(54),Cin=>p(211)(54),clock=>clock,reset=>reset,s=>p(268)(54),cout=>p(269)(55));
FA_ff_8859:FAff port map(x=>p(209)(55),y=>p(210)(55),Cin=>p(211)(55),clock=>clock,reset=>reset,s=>p(268)(55),cout=>p(269)(56));
FA_ff_8860:FAff port map(x=>p(209)(56),y=>p(210)(56),Cin=>p(211)(56),clock=>clock,reset=>reset,s=>p(268)(56),cout=>p(269)(57));
FA_ff_8861:FAff port map(x=>p(209)(57),y=>p(210)(57),Cin=>p(211)(57),clock=>clock,reset=>reset,s=>p(268)(57),cout=>p(269)(58));
FA_ff_8862:FAff port map(x=>p(209)(58),y=>p(210)(58),Cin=>p(211)(58),clock=>clock,reset=>reset,s=>p(268)(58),cout=>p(269)(59));
FA_ff_8863:FAff port map(x=>p(209)(59),y=>p(210)(59),Cin=>p(211)(59),clock=>clock,reset=>reset,s=>p(268)(59),cout=>p(269)(60));
FA_ff_8864:FAff port map(x=>p(209)(60),y=>p(210)(60),Cin=>p(211)(60),clock=>clock,reset=>reset,s=>p(268)(60),cout=>p(269)(61));
FA_ff_8865:FAff port map(x=>p(209)(61),y=>p(210)(61),Cin=>p(211)(61),clock=>clock,reset=>reset,s=>p(268)(61),cout=>p(269)(62));
FA_ff_8866:FAff port map(x=>p(209)(62),y=>p(210)(62),Cin=>p(211)(62),clock=>clock,reset=>reset,s=>p(268)(62),cout=>p(269)(63));
FA_ff_8867:FAff port map(x=>p(209)(63),y=>p(210)(63),Cin=>p(211)(63),clock=>clock,reset=>reset,s=>p(268)(63),cout=>p(269)(64));
FA_ff_8868:FAff port map(x=>p(209)(64),y=>p(210)(64),Cin=>p(211)(64),clock=>clock,reset=>reset,s=>p(268)(64),cout=>p(269)(65));
FA_ff_8869:FAff port map(x=>p(209)(65),y=>p(210)(65),Cin=>p(211)(65),clock=>clock,reset=>reset,s=>p(268)(65),cout=>p(269)(66));
FA_ff_8870:FAff port map(x=>p(209)(66),y=>p(210)(66),Cin=>p(211)(66),clock=>clock,reset=>reset,s=>p(268)(66),cout=>p(269)(67));
FA_ff_8871:FAff port map(x=>p(209)(67),y=>p(210)(67),Cin=>p(211)(67),clock=>clock,reset=>reset,s=>p(268)(67),cout=>p(269)(68));
FA_ff_8872:FAff port map(x=>p(209)(68),y=>p(210)(68),Cin=>p(211)(68),clock=>clock,reset=>reset,s=>p(268)(68),cout=>p(269)(69));
FA_ff_8873:FAff port map(x=>p(209)(69),y=>p(210)(69),Cin=>p(211)(69),clock=>clock,reset=>reset,s=>p(268)(69),cout=>p(269)(70));
FA_ff_8874:FAff port map(x=>p(209)(70),y=>p(210)(70),Cin=>p(211)(70),clock=>clock,reset=>reset,s=>p(268)(70),cout=>p(269)(71));
FA_ff_8875:FAff port map(x=>p(209)(71),y=>p(210)(71),Cin=>p(211)(71),clock=>clock,reset=>reset,s=>p(268)(71),cout=>p(269)(72));
FA_ff_8876:FAff port map(x=>p(209)(72),y=>p(210)(72),Cin=>p(211)(72),clock=>clock,reset=>reset,s=>p(268)(72),cout=>p(269)(73));
FA_ff_8877:FAff port map(x=>p(209)(73),y=>p(210)(73),Cin=>p(211)(73),clock=>clock,reset=>reset,s=>p(268)(73),cout=>p(269)(74));
FA_ff_8878:FAff port map(x=>p(209)(74),y=>p(210)(74),Cin=>p(211)(74),clock=>clock,reset=>reset,s=>p(268)(74),cout=>p(269)(75));
FA_ff_8879:FAff port map(x=>p(209)(75),y=>p(210)(75),Cin=>p(211)(75),clock=>clock,reset=>reset,s=>p(268)(75),cout=>p(269)(76));
FA_ff_8880:FAff port map(x=>p(209)(76),y=>p(210)(76),Cin=>p(211)(76),clock=>clock,reset=>reset,s=>p(268)(76),cout=>p(269)(77));
FA_ff_8881:FAff port map(x=>p(209)(77),y=>p(210)(77),Cin=>p(211)(77),clock=>clock,reset=>reset,s=>p(268)(77),cout=>p(269)(78));
FA_ff_8882:FAff port map(x=>p(209)(78),y=>p(210)(78),Cin=>p(211)(78),clock=>clock,reset=>reset,s=>p(268)(78),cout=>p(269)(79));
FA_ff_8883:FAff port map(x=>p(209)(79),y=>p(210)(79),Cin=>p(211)(79),clock=>clock,reset=>reset,s=>p(268)(79),cout=>p(269)(80));
FA_ff_8884:FAff port map(x=>p(209)(80),y=>p(210)(80),Cin=>p(211)(80),clock=>clock,reset=>reset,s=>p(268)(80),cout=>p(269)(81));
FA_ff_8885:FAff port map(x=>p(209)(81),y=>p(210)(81),Cin=>p(211)(81),clock=>clock,reset=>reset,s=>p(268)(81),cout=>p(269)(82));
FA_ff_8886:FAff port map(x=>p(209)(82),y=>p(210)(82),Cin=>p(211)(82),clock=>clock,reset=>reset,s=>p(268)(82),cout=>p(269)(83));
FA_ff_8887:FAff port map(x=>p(209)(83),y=>p(210)(83),Cin=>p(211)(83),clock=>clock,reset=>reset,s=>p(268)(83),cout=>p(269)(84));
FA_ff_8888:FAff port map(x=>p(209)(84),y=>p(210)(84),Cin=>p(211)(84),clock=>clock,reset=>reset,s=>p(268)(84),cout=>p(269)(85));
FA_ff_8889:FAff port map(x=>p(209)(85),y=>p(210)(85),Cin=>p(211)(85),clock=>clock,reset=>reset,s=>p(268)(85),cout=>p(269)(86));
FA_ff_8890:FAff port map(x=>p(209)(86),y=>p(210)(86),Cin=>p(211)(86),clock=>clock,reset=>reset,s=>p(268)(86),cout=>p(269)(87));
FA_ff_8891:FAff port map(x=>p(209)(87),y=>p(210)(87),Cin=>p(211)(87),clock=>clock,reset=>reset,s=>p(268)(87),cout=>p(269)(88));
FA_ff_8892:FAff port map(x=>p(209)(88),y=>p(210)(88),Cin=>p(211)(88),clock=>clock,reset=>reset,s=>p(268)(88),cout=>p(269)(89));
FA_ff_8893:FAff port map(x=>p(209)(89),y=>p(210)(89),Cin=>p(211)(89),clock=>clock,reset=>reset,s=>p(268)(89),cout=>p(269)(90));
FA_ff_8894:FAff port map(x=>p(209)(90),y=>p(210)(90),Cin=>p(211)(90),clock=>clock,reset=>reset,s=>p(268)(90),cout=>p(269)(91));
FA_ff_8895:FAff port map(x=>p(209)(91),y=>p(210)(91),Cin=>p(211)(91),clock=>clock,reset=>reset,s=>p(268)(91),cout=>p(269)(92));
FA_ff_8896:FAff port map(x=>p(209)(92),y=>p(210)(92),Cin=>p(211)(92),clock=>clock,reset=>reset,s=>p(268)(92),cout=>p(269)(93));
FA_ff_8897:FAff port map(x=>p(209)(93),y=>p(210)(93),Cin=>p(211)(93),clock=>clock,reset=>reset,s=>p(268)(93),cout=>p(269)(94));
FA_ff_8898:FAff port map(x=>p(209)(94),y=>p(210)(94),Cin=>p(211)(94),clock=>clock,reset=>reset,s=>p(268)(94),cout=>p(269)(95));
FA_ff_8899:FAff port map(x=>p(209)(95),y=>p(210)(95),Cin=>p(211)(95),clock=>clock,reset=>reset,s=>p(268)(95),cout=>p(269)(96));
FA_ff_8900:FAff port map(x=>p(209)(96),y=>p(210)(96),Cin=>p(211)(96),clock=>clock,reset=>reset,s=>p(268)(96),cout=>p(269)(97));
FA_ff_8901:FAff port map(x=>p(209)(97),y=>p(210)(97),Cin=>p(211)(97),clock=>clock,reset=>reset,s=>p(268)(97),cout=>p(269)(98));
FA_ff_8902:FAff port map(x=>p(209)(98),y=>p(210)(98),Cin=>p(211)(98),clock=>clock,reset=>reset,s=>p(268)(98),cout=>p(269)(99));
FA_ff_8903:FAff port map(x=>p(209)(99),y=>p(210)(99),Cin=>p(211)(99),clock=>clock,reset=>reset,s=>p(268)(99),cout=>p(269)(100));
FA_ff_8904:FAff port map(x=>p(209)(100),y=>p(210)(100),Cin=>p(211)(100),clock=>clock,reset=>reset,s=>p(268)(100),cout=>p(269)(101));
FA_ff_8905:FAff port map(x=>p(209)(101),y=>p(210)(101),Cin=>p(211)(101),clock=>clock,reset=>reset,s=>p(268)(101),cout=>p(269)(102));
FA_ff_8906:FAff port map(x=>p(209)(102),y=>p(210)(102),Cin=>p(211)(102),clock=>clock,reset=>reset,s=>p(268)(102),cout=>p(269)(103));
FA_ff_8907:FAff port map(x=>p(209)(103),y=>p(210)(103),Cin=>p(211)(103),clock=>clock,reset=>reset,s=>p(268)(103),cout=>p(269)(104));
FA_ff_8908:FAff port map(x=>p(209)(104),y=>p(210)(104),Cin=>p(211)(104),clock=>clock,reset=>reset,s=>p(268)(104),cout=>p(269)(105));
FA_ff_8909:FAff port map(x=>p(209)(105),y=>p(210)(105),Cin=>p(211)(105),clock=>clock,reset=>reset,s=>p(268)(105),cout=>p(269)(106));
FA_ff_8910:FAff port map(x=>p(209)(106),y=>p(210)(106),Cin=>p(211)(106),clock=>clock,reset=>reset,s=>p(268)(106),cout=>p(269)(107));
FA_ff_8911:FAff port map(x=>p(209)(107),y=>p(210)(107),Cin=>p(211)(107),clock=>clock,reset=>reset,s=>p(268)(107),cout=>p(269)(108));
FA_ff_8912:FAff port map(x=>p(209)(108),y=>p(210)(108),Cin=>p(211)(108),clock=>clock,reset=>reset,s=>p(268)(108),cout=>p(269)(109));
FA_ff_8913:FAff port map(x=>p(209)(109),y=>p(210)(109),Cin=>p(211)(109),clock=>clock,reset=>reset,s=>p(268)(109),cout=>p(269)(110));
FA_ff_8914:FAff port map(x=>p(209)(110),y=>p(210)(110),Cin=>p(211)(110),clock=>clock,reset=>reset,s=>p(268)(110),cout=>p(269)(111));
FA_ff_8915:FAff port map(x=>p(209)(111),y=>p(210)(111),Cin=>p(211)(111),clock=>clock,reset=>reset,s=>p(268)(111),cout=>p(269)(112));
FA_ff_8916:FAff port map(x=>p(209)(112),y=>p(210)(112),Cin=>p(211)(112),clock=>clock,reset=>reset,s=>p(268)(112),cout=>p(269)(113));
FA_ff_8917:FAff port map(x=>p(209)(113),y=>p(210)(113),Cin=>p(211)(113),clock=>clock,reset=>reset,s=>p(268)(113),cout=>p(269)(114));
FA_ff_8918:FAff port map(x=>p(209)(114),y=>p(210)(114),Cin=>p(211)(114),clock=>clock,reset=>reset,s=>p(268)(114),cout=>p(269)(115));
FA_ff_8919:FAff port map(x=>p(209)(115),y=>p(210)(115),Cin=>p(211)(115),clock=>clock,reset=>reset,s=>p(268)(115),cout=>p(269)(116));
FA_ff_8920:FAff port map(x=>p(209)(116),y=>p(210)(116),Cin=>p(211)(116),clock=>clock,reset=>reset,s=>p(268)(116),cout=>p(269)(117));
FA_ff_8921:FAff port map(x=>p(209)(117),y=>p(210)(117),Cin=>p(211)(117),clock=>clock,reset=>reset,s=>p(268)(117),cout=>p(269)(118));
FA_ff_8922:FAff port map(x=>p(209)(118),y=>p(210)(118),Cin=>p(211)(118),clock=>clock,reset=>reset,s=>p(268)(118),cout=>p(269)(119));
FA_ff_8923:FAff port map(x=>p(209)(119),y=>p(210)(119),Cin=>p(211)(119),clock=>clock,reset=>reset,s=>p(268)(119),cout=>p(269)(120));
FA_ff_8924:FAff port map(x=>p(209)(120),y=>p(210)(120),Cin=>p(211)(120),clock=>clock,reset=>reset,s=>p(268)(120),cout=>p(269)(121));
FA_ff_8925:FAff port map(x=>p(209)(121),y=>p(210)(121),Cin=>p(211)(121),clock=>clock,reset=>reset,s=>p(268)(121),cout=>p(269)(122));
FA_ff_8926:FAff port map(x=>p(209)(122),y=>p(210)(122),Cin=>p(211)(122),clock=>clock,reset=>reset,s=>p(268)(122),cout=>p(269)(123));
FA_ff_8927:FAff port map(x=>p(209)(123),y=>p(210)(123),Cin=>p(211)(123),clock=>clock,reset=>reset,s=>p(268)(123),cout=>p(269)(124));
FA_ff_8928:FAff port map(x=>p(209)(124),y=>p(210)(124),Cin=>p(211)(124),clock=>clock,reset=>reset,s=>p(268)(124),cout=>p(269)(125));
FA_ff_8929:FAff port map(x=>p(209)(125),y=>p(210)(125),Cin=>p(211)(125),clock=>clock,reset=>reset,s=>p(268)(125),cout=>p(269)(126));
FA_ff_8930:FAff port map(x=>p(209)(126),y=>p(210)(126),Cin=>p(211)(126),clock=>clock,reset=>reset,s=>p(268)(126),cout=>p(269)(127));
FA_ff_8931:FAff port map(x=>p(209)(127),y=>p(210)(127),Cin=>p(211)(127),clock=>clock,reset=>reset,s=>p(268)(127),cout=>p(269)(128));
HA_ff_27:HAff port map(x=>p(209)(128),y=>p(211)(128),clock=>clock,reset=>reset,s=>p(268)(128),c=>p(269)(129));
p(270)(0)<=p(212)(0);
p(270)(1)<=p(212)(1);
p(270)(2)<=p(212)(2);
p(270)(3)<=p(212)(3);
p(270)(4)<=p(212)(4);
p(270)(5)<=p(212)(5);
p(270)(6)<=p(212)(6);
p(270)(7)<=p(212)(7);
p(270)(8)<=p(212)(8);
p(270)(9)<=p(212)(9);
p(270)(10)<=p(212)(10);
p(270)(11)<=p(212)(11);
p(270)(12)<=p(212)(12);
p(270)(13)<=p(212)(13);
p(270)(14)<=p(212)(14);
p(270)(15)<=p(212)(15);
p(270)(16)<=p(212)(16);
p(270)(17)<=p(212)(17);
p(270)(18)<=p(212)(18);
p(270)(19)<=p(212)(19);
p(270)(20)<=p(212)(20);
p(270)(21)<=p(212)(21);
p(270)(22)<=p(212)(22);
p(270)(23)<=p(212)(23);
p(270)(24)<=p(212)(24);
p(270)(25)<=p(212)(25);
p(270)(26)<=p(212)(26);
p(270)(27)<=p(212)(27);
p(270)(28)<=p(212)(28);
p(270)(29)<=p(212)(29);
p(270)(30)<=p(212)(30);
p(270)(31)<=p(212)(31);
p(270)(32)<=p(212)(32);
p(270)(33)<=p(212)(33);
p(270)(34)<=p(212)(34);
p(270)(35)<=p(212)(35);
p(270)(36)<=p(212)(36);
p(270)(37)<=p(212)(37);
p(270)(38)<=p(212)(38);
p(270)(39)<=p(212)(39);
p(270)(40)<=p(212)(40);
p(270)(41)<=p(212)(41);
p(270)(42)<=p(212)(42);
p(270)(43)<=p(212)(43);
p(270)(44)<=p(212)(44);
p(270)(45)<=p(212)(45);
p(270)(46)<=p(212)(46);
p(270)(47)<=p(212)(47);
p(270)(48)<=p(212)(48);
p(270)(49)<=p(212)(49);
p(270)(50)<=p(212)(50);
p(270)(51)<=p(212)(51);
p(270)(52)<=p(212)(52);
p(270)(53)<=p(212)(53);
p(270)(54)<=p(212)(54);
p(270)(55)<=p(212)(55);
p(270)(56)<=p(212)(56);
p(270)(57)<=p(212)(57);
p(270)(58)<=p(212)(58);
p(270)(59)<=p(212)(59);
p(270)(60)<=p(212)(60);
p(270)(61)<=p(212)(61);
p(270)(62)<=p(212)(62);
p(270)(63)<=p(212)(63);
p(270)(64)<=p(212)(64);
p(270)(65)<=p(212)(65);
p(270)(66)<=p(212)(66);
p(270)(67)<=p(212)(67);
p(270)(68)<=p(212)(68);
p(270)(69)<=p(212)(69);
p(270)(70)<=p(212)(70);
p(270)(71)<=p(212)(71);
p(270)(72)<=p(212)(72);
p(270)(73)<=p(212)(73);
p(270)(74)<=p(212)(74);
p(270)(75)<=p(212)(75);
p(270)(76)<=p(212)(76);
p(270)(77)<=p(212)(77);
p(270)(78)<=p(212)(78);
p(270)(79)<=p(212)(79);
p(270)(80)<=p(212)(80);
p(270)(81)<=p(212)(81);
p(270)(82)<=p(212)(82);
p(270)(83)<=p(212)(83);
p(270)(84)<=p(212)(84);
p(270)(85)<=p(212)(85);
p(270)(86)<=p(212)(86);
p(270)(87)<=p(212)(87);
p(270)(88)<=p(212)(88);
p(270)(89)<=p(212)(89);
p(270)(90)<=p(212)(90);
p(270)(91)<=p(212)(91);
p(270)(92)<=p(212)(92);
p(270)(93)<=p(212)(93);
p(270)(94)<=p(212)(94);
p(270)(95)<=p(212)(95);
p(270)(96)<=p(212)(96);
p(270)(97)<=p(212)(97);
p(270)(98)<=p(212)(98);
p(270)(99)<=p(212)(99);
p(270)(100)<=p(212)(100);
p(270)(101)<=p(212)(101);
p(270)(102)<=p(212)(102);
p(270)(103)<=p(212)(103);
p(270)(104)<=p(212)(104);
p(270)(105)<=p(212)(105);
p(270)(106)<=p(212)(106);
p(270)(107)<=p(212)(107);
p(270)(108)<=p(212)(108);
p(270)(109)<=p(212)(109);
p(270)(110)<=p(212)(110);
p(270)(111)<=p(212)(111);
p(270)(112)<=p(212)(112);
p(270)(113)<=p(212)(113);
p(270)(114)<=p(212)(114);
p(270)(115)<=p(212)(115);
p(270)(116)<=p(212)(116);
p(270)(117)<=p(212)(117);
p(270)(118)<=p(212)(118);
p(270)(119)<=p(212)(119);
p(270)(120)<=p(212)(120);
p(270)(121)<=p(212)(121);
p(270)(122)<=p(212)(122);
p(270)(123)<=p(212)(123);
p(270)(124)<=p(212)(124);
p(270)(125)<=p(212)(125);
p(270)(126)<=p(212)(126);
p(270)(127)<=p(212)(127);
p(270)(128)<=p(212)(128);
p(270)(129)<=p(212)(129);
p(270)(130)<=p(212)(130);
p(270)(131)<=p(212)(131);
p(270)(132)<=p(212)(132);
p(270)(133)<=p(212)(133);
p(270)(134)<=p(212)(134);
p(271)(0)<=p(213)(0);
p(271)(1)<=p(213)(1);
p(271)(2)<=p(213)(2);
p(271)(3)<=p(213)(3);
p(271)(4)<=p(213)(4);
p(271)(5)<=p(213)(5);
p(271)(6)<=p(213)(6);
p(271)(7)<=p(213)(7);
p(271)(8)<=p(213)(8);
p(271)(9)<=p(213)(9);
p(271)(10)<=p(213)(10);
p(271)(11)<=p(213)(11);
p(271)(12)<=p(213)(12);
p(271)(13)<=p(213)(13);
p(271)(14)<=p(213)(14);
p(271)(15)<=p(213)(15);
p(271)(16)<=p(213)(16);
p(271)(17)<=p(213)(17);
p(271)(18)<=p(213)(18);
p(271)(19)<=p(213)(19);
p(271)(20)<=p(213)(20);
p(271)(21)<=p(213)(21);
p(271)(22)<=p(213)(22);
p(271)(23)<=p(213)(23);
p(271)(24)<=p(213)(24);
p(271)(25)<=p(213)(25);
p(271)(26)<=p(213)(26);
p(271)(27)<=p(213)(27);
p(271)(28)<=p(213)(28);
p(271)(29)<=p(213)(29);
p(271)(30)<=p(213)(30);
p(271)(31)<=p(213)(31);
p(271)(32)<=p(213)(32);
p(271)(33)<=p(213)(33);
p(271)(34)<=p(213)(34);
p(271)(35)<=p(213)(35);
p(271)(36)<=p(213)(36);
p(271)(37)<=p(213)(37);
p(271)(38)<=p(213)(38);
p(271)(39)<=p(213)(39);
p(271)(40)<=p(213)(40);
p(271)(41)<=p(213)(41);
p(271)(42)<=p(213)(42);
p(271)(43)<=p(213)(43);
p(271)(44)<=p(213)(44);
p(271)(45)<=p(213)(45);
p(271)(46)<=p(213)(46);
p(271)(47)<=p(213)(47);
p(271)(48)<=p(213)(48);
p(271)(49)<=p(213)(49);
p(271)(50)<=p(213)(50);
p(271)(51)<=p(213)(51);
p(271)(52)<=p(213)(52);
p(271)(53)<=p(213)(53);
p(271)(54)<=p(213)(54);
p(271)(55)<=p(213)(55);
p(271)(56)<=p(213)(56);
p(271)(57)<=p(213)(57);
p(271)(58)<=p(213)(58);
p(271)(59)<=p(213)(59);
p(271)(60)<=p(213)(60);
p(271)(61)<=p(213)(61);
p(271)(62)<=p(213)(62);
p(271)(63)<=p(213)(63);
p(271)(64)<=p(213)(64);
p(271)(65)<=p(213)(65);
p(271)(66)<=p(213)(66);
p(271)(67)<=p(213)(67);
p(271)(68)<=p(213)(68);
p(271)(69)<=p(213)(69);
p(271)(70)<=p(213)(70);
p(271)(71)<=p(213)(71);
p(271)(72)<=p(213)(72);
p(271)(73)<=p(213)(73);
p(271)(74)<=p(213)(74);
p(271)(75)<=p(213)(75);
p(271)(76)<=p(213)(76);
p(271)(77)<=p(213)(77);
p(271)(78)<=p(213)(78);
p(271)(79)<=p(213)(79);
p(271)(80)<=p(213)(80);
p(271)(81)<=p(213)(81);
p(271)(82)<=p(213)(82);
p(271)(83)<=p(213)(83);
p(271)(84)<=p(213)(84);
p(271)(85)<=p(213)(85);
p(271)(86)<=p(213)(86);
p(271)(87)<=p(213)(87);
p(271)(88)<=p(213)(88);
p(271)(89)<=p(213)(89);
p(271)(90)<=p(213)(90);
p(271)(91)<=p(213)(91);
p(271)(92)<=p(213)(92);
p(271)(93)<=p(213)(93);
p(271)(94)<=p(213)(94);
p(271)(95)<=p(213)(95);
p(271)(96)<=p(213)(96);
p(271)(97)<=p(213)(97);
p(271)(98)<=p(213)(98);
p(271)(99)<=p(213)(99);
p(271)(100)<=p(213)(100);
p(271)(101)<=p(213)(101);
p(271)(102)<=p(213)(102);
p(271)(103)<=p(213)(103);
p(271)(104)<=p(213)(104);
p(271)(105)<=p(213)(105);
p(271)(106)<=p(213)(106);
p(271)(107)<=p(213)(107);
p(271)(108)<=p(213)(108);
p(271)(109)<=p(213)(109);
p(271)(110)<=p(213)(110);
p(271)(111)<=p(213)(111);
p(271)(112)<=p(213)(112);
p(271)(113)<=p(213)(113);
p(271)(114)<=p(213)(114);
p(271)(115)<=p(213)(115);
p(271)(116)<=p(213)(116);
p(271)(117)<=p(213)(117);
p(271)(118)<=p(213)(118);
p(271)(119)<=p(213)(119);
p(271)(120)<=p(213)(120);
p(271)(121)<=p(213)(121);
p(271)(122)<=p(213)(122);
p(271)(123)<=p(213)(123);
p(271)(124)<=p(213)(124);
p(271)(125)<=p(213)(125);
p(271)(126)<=p(213)(126);
p(271)(127)<=p(213)(127);
p(271)(128)<=p(213)(128);
p(271)(129)<=p(213)(129);
p(271)(130)<=p(213)(130);
p(271)(131)<=p(213)(131);
p(271)(132)<=p(213)(132);
p(271)(133)<=p(213)(133);
p(271)(134)<=p(213)(134);
HA_ff_28:HAff port map(x=>p(214)(0),y=>p(216)(0),clock=>clock,reset=>reset,s=>p(272)(0),c=>p(273)(1));
FA_ff_8932:FAff port map(x=>p(214)(1),y=>p(215)(1),Cin=>p(216)(1),clock=>clock,reset=>reset,s=>p(272)(1),cout=>p(273)(2));
FA_ff_8933:FAff port map(x=>p(214)(2),y=>p(215)(2),Cin=>p(216)(2),clock=>clock,reset=>reset,s=>p(272)(2),cout=>p(273)(3));
FA_ff_8934:FAff port map(x=>p(214)(3),y=>p(215)(3),Cin=>p(216)(3),clock=>clock,reset=>reset,s=>p(272)(3),cout=>p(273)(4));
FA_ff_8935:FAff port map(x=>p(214)(4),y=>p(215)(4),Cin=>p(216)(4),clock=>clock,reset=>reset,s=>p(272)(4),cout=>p(273)(5));
FA_ff_8936:FAff port map(x=>p(214)(5),y=>p(215)(5),Cin=>p(216)(5),clock=>clock,reset=>reset,s=>p(272)(5),cout=>p(273)(6));
FA_ff_8937:FAff port map(x=>p(214)(6),y=>p(215)(6),Cin=>p(216)(6),clock=>clock,reset=>reset,s=>p(272)(6),cout=>p(273)(7));
FA_ff_8938:FAff port map(x=>p(214)(7),y=>p(215)(7),Cin=>p(216)(7),clock=>clock,reset=>reset,s=>p(272)(7),cout=>p(273)(8));
FA_ff_8939:FAff port map(x=>p(214)(8),y=>p(215)(8),Cin=>p(216)(8),clock=>clock,reset=>reset,s=>p(272)(8),cout=>p(273)(9));
FA_ff_8940:FAff port map(x=>p(214)(9),y=>p(215)(9),Cin=>p(216)(9),clock=>clock,reset=>reset,s=>p(272)(9),cout=>p(273)(10));
FA_ff_8941:FAff port map(x=>p(214)(10),y=>p(215)(10),Cin=>p(216)(10),clock=>clock,reset=>reset,s=>p(272)(10),cout=>p(273)(11));
FA_ff_8942:FAff port map(x=>p(214)(11),y=>p(215)(11),Cin=>p(216)(11),clock=>clock,reset=>reset,s=>p(272)(11),cout=>p(273)(12));
FA_ff_8943:FAff port map(x=>p(214)(12),y=>p(215)(12),Cin=>p(216)(12),clock=>clock,reset=>reset,s=>p(272)(12),cout=>p(273)(13));
FA_ff_8944:FAff port map(x=>p(214)(13),y=>p(215)(13),Cin=>p(216)(13),clock=>clock,reset=>reset,s=>p(272)(13),cout=>p(273)(14));
FA_ff_8945:FAff port map(x=>p(214)(14),y=>p(215)(14),Cin=>p(216)(14),clock=>clock,reset=>reset,s=>p(272)(14),cout=>p(273)(15));
FA_ff_8946:FAff port map(x=>p(214)(15),y=>p(215)(15),Cin=>p(216)(15),clock=>clock,reset=>reset,s=>p(272)(15),cout=>p(273)(16));
FA_ff_8947:FAff port map(x=>p(214)(16),y=>p(215)(16),Cin=>p(216)(16),clock=>clock,reset=>reset,s=>p(272)(16),cout=>p(273)(17));
FA_ff_8948:FAff port map(x=>p(214)(17),y=>p(215)(17),Cin=>p(216)(17),clock=>clock,reset=>reset,s=>p(272)(17),cout=>p(273)(18));
FA_ff_8949:FAff port map(x=>p(214)(18),y=>p(215)(18),Cin=>p(216)(18),clock=>clock,reset=>reset,s=>p(272)(18),cout=>p(273)(19));
FA_ff_8950:FAff port map(x=>p(214)(19),y=>p(215)(19),Cin=>p(216)(19),clock=>clock,reset=>reset,s=>p(272)(19),cout=>p(273)(20));
FA_ff_8951:FAff port map(x=>p(214)(20),y=>p(215)(20),Cin=>p(216)(20),clock=>clock,reset=>reset,s=>p(272)(20),cout=>p(273)(21));
FA_ff_8952:FAff port map(x=>p(214)(21),y=>p(215)(21),Cin=>p(216)(21),clock=>clock,reset=>reset,s=>p(272)(21),cout=>p(273)(22));
FA_ff_8953:FAff port map(x=>p(214)(22),y=>p(215)(22),Cin=>p(216)(22),clock=>clock,reset=>reset,s=>p(272)(22),cout=>p(273)(23));
FA_ff_8954:FAff port map(x=>p(214)(23),y=>p(215)(23),Cin=>p(216)(23),clock=>clock,reset=>reset,s=>p(272)(23),cout=>p(273)(24));
FA_ff_8955:FAff port map(x=>p(214)(24),y=>p(215)(24),Cin=>p(216)(24),clock=>clock,reset=>reset,s=>p(272)(24),cout=>p(273)(25));
FA_ff_8956:FAff port map(x=>p(214)(25),y=>p(215)(25),Cin=>p(216)(25),clock=>clock,reset=>reset,s=>p(272)(25),cout=>p(273)(26));
FA_ff_8957:FAff port map(x=>p(214)(26),y=>p(215)(26),Cin=>p(216)(26),clock=>clock,reset=>reset,s=>p(272)(26),cout=>p(273)(27));
FA_ff_8958:FAff port map(x=>p(214)(27),y=>p(215)(27),Cin=>p(216)(27),clock=>clock,reset=>reset,s=>p(272)(27),cout=>p(273)(28));
FA_ff_8959:FAff port map(x=>p(214)(28),y=>p(215)(28),Cin=>p(216)(28),clock=>clock,reset=>reset,s=>p(272)(28),cout=>p(273)(29));
FA_ff_8960:FAff port map(x=>p(214)(29),y=>p(215)(29),Cin=>p(216)(29),clock=>clock,reset=>reset,s=>p(272)(29),cout=>p(273)(30));
FA_ff_8961:FAff port map(x=>p(214)(30),y=>p(215)(30),Cin=>p(216)(30),clock=>clock,reset=>reset,s=>p(272)(30),cout=>p(273)(31));
FA_ff_8962:FAff port map(x=>p(214)(31),y=>p(215)(31),Cin=>p(216)(31),clock=>clock,reset=>reset,s=>p(272)(31),cout=>p(273)(32));
FA_ff_8963:FAff port map(x=>p(214)(32),y=>p(215)(32),Cin=>p(216)(32),clock=>clock,reset=>reset,s=>p(272)(32),cout=>p(273)(33));
FA_ff_8964:FAff port map(x=>p(214)(33),y=>p(215)(33),Cin=>p(216)(33),clock=>clock,reset=>reset,s=>p(272)(33),cout=>p(273)(34));
FA_ff_8965:FAff port map(x=>p(214)(34),y=>p(215)(34),Cin=>p(216)(34),clock=>clock,reset=>reset,s=>p(272)(34),cout=>p(273)(35));
FA_ff_8966:FAff port map(x=>p(214)(35),y=>p(215)(35),Cin=>p(216)(35),clock=>clock,reset=>reset,s=>p(272)(35),cout=>p(273)(36));
FA_ff_8967:FAff port map(x=>p(214)(36),y=>p(215)(36),Cin=>p(216)(36),clock=>clock,reset=>reset,s=>p(272)(36),cout=>p(273)(37));
FA_ff_8968:FAff port map(x=>p(214)(37),y=>p(215)(37),Cin=>p(216)(37),clock=>clock,reset=>reset,s=>p(272)(37),cout=>p(273)(38));
FA_ff_8969:FAff port map(x=>p(214)(38),y=>p(215)(38),Cin=>p(216)(38),clock=>clock,reset=>reset,s=>p(272)(38),cout=>p(273)(39));
FA_ff_8970:FAff port map(x=>p(214)(39),y=>p(215)(39),Cin=>p(216)(39),clock=>clock,reset=>reset,s=>p(272)(39),cout=>p(273)(40));
FA_ff_8971:FAff port map(x=>p(214)(40),y=>p(215)(40),Cin=>p(216)(40),clock=>clock,reset=>reset,s=>p(272)(40),cout=>p(273)(41));
FA_ff_8972:FAff port map(x=>p(214)(41),y=>p(215)(41),Cin=>p(216)(41),clock=>clock,reset=>reset,s=>p(272)(41),cout=>p(273)(42));
FA_ff_8973:FAff port map(x=>p(214)(42),y=>p(215)(42),Cin=>p(216)(42),clock=>clock,reset=>reset,s=>p(272)(42),cout=>p(273)(43));
FA_ff_8974:FAff port map(x=>p(214)(43),y=>p(215)(43),Cin=>p(216)(43),clock=>clock,reset=>reset,s=>p(272)(43),cout=>p(273)(44));
FA_ff_8975:FAff port map(x=>p(214)(44),y=>p(215)(44),Cin=>p(216)(44),clock=>clock,reset=>reset,s=>p(272)(44),cout=>p(273)(45));
FA_ff_8976:FAff port map(x=>p(214)(45),y=>p(215)(45),Cin=>p(216)(45),clock=>clock,reset=>reset,s=>p(272)(45),cout=>p(273)(46));
FA_ff_8977:FAff port map(x=>p(214)(46),y=>p(215)(46),Cin=>p(216)(46),clock=>clock,reset=>reset,s=>p(272)(46),cout=>p(273)(47));
FA_ff_8978:FAff port map(x=>p(214)(47),y=>p(215)(47),Cin=>p(216)(47),clock=>clock,reset=>reset,s=>p(272)(47),cout=>p(273)(48));
FA_ff_8979:FAff port map(x=>p(214)(48),y=>p(215)(48),Cin=>p(216)(48),clock=>clock,reset=>reset,s=>p(272)(48),cout=>p(273)(49));
FA_ff_8980:FAff port map(x=>p(214)(49),y=>p(215)(49),Cin=>p(216)(49),clock=>clock,reset=>reset,s=>p(272)(49),cout=>p(273)(50));
FA_ff_8981:FAff port map(x=>p(214)(50),y=>p(215)(50),Cin=>p(216)(50),clock=>clock,reset=>reset,s=>p(272)(50),cout=>p(273)(51));
FA_ff_8982:FAff port map(x=>p(214)(51),y=>p(215)(51),Cin=>p(216)(51),clock=>clock,reset=>reset,s=>p(272)(51),cout=>p(273)(52));
FA_ff_8983:FAff port map(x=>p(214)(52),y=>p(215)(52),Cin=>p(216)(52),clock=>clock,reset=>reset,s=>p(272)(52),cout=>p(273)(53));
FA_ff_8984:FAff port map(x=>p(214)(53),y=>p(215)(53),Cin=>p(216)(53),clock=>clock,reset=>reset,s=>p(272)(53),cout=>p(273)(54));
FA_ff_8985:FAff port map(x=>p(214)(54),y=>p(215)(54),Cin=>p(216)(54),clock=>clock,reset=>reset,s=>p(272)(54),cout=>p(273)(55));
FA_ff_8986:FAff port map(x=>p(214)(55),y=>p(215)(55),Cin=>p(216)(55),clock=>clock,reset=>reset,s=>p(272)(55),cout=>p(273)(56));
FA_ff_8987:FAff port map(x=>p(214)(56),y=>p(215)(56),Cin=>p(216)(56),clock=>clock,reset=>reset,s=>p(272)(56),cout=>p(273)(57));
FA_ff_8988:FAff port map(x=>p(214)(57),y=>p(215)(57),Cin=>p(216)(57),clock=>clock,reset=>reset,s=>p(272)(57),cout=>p(273)(58));
FA_ff_8989:FAff port map(x=>p(214)(58),y=>p(215)(58),Cin=>p(216)(58),clock=>clock,reset=>reset,s=>p(272)(58),cout=>p(273)(59));
FA_ff_8990:FAff port map(x=>p(214)(59),y=>p(215)(59),Cin=>p(216)(59),clock=>clock,reset=>reset,s=>p(272)(59),cout=>p(273)(60));
FA_ff_8991:FAff port map(x=>p(214)(60),y=>p(215)(60),Cin=>p(216)(60),clock=>clock,reset=>reset,s=>p(272)(60),cout=>p(273)(61));
FA_ff_8992:FAff port map(x=>p(214)(61),y=>p(215)(61),Cin=>p(216)(61),clock=>clock,reset=>reset,s=>p(272)(61),cout=>p(273)(62));
FA_ff_8993:FAff port map(x=>p(214)(62),y=>p(215)(62),Cin=>p(216)(62),clock=>clock,reset=>reset,s=>p(272)(62),cout=>p(273)(63));
FA_ff_8994:FAff port map(x=>p(214)(63),y=>p(215)(63),Cin=>p(216)(63),clock=>clock,reset=>reset,s=>p(272)(63),cout=>p(273)(64));
FA_ff_8995:FAff port map(x=>p(214)(64),y=>p(215)(64),Cin=>p(216)(64),clock=>clock,reset=>reset,s=>p(272)(64),cout=>p(273)(65));
FA_ff_8996:FAff port map(x=>p(214)(65),y=>p(215)(65),Cin=>p(216)(65),clock=>clock,reset=>reset,s=>p(272)(65),cout=>p(273)(66));
FA_ff_8997:FAff port map(x=>p(214)(66),y=>p(215)(66),Cin=>p(216)(66),clock=>clock,reset=>reset,s=>p(272)(66),cout=>p(273)(67));
FA_ff_8998:FAff port map(x=>p(214)(67),y=>p(215)(67),Cin=>p(216)(67),clock=>clock,reset=>reset,s=>p(272)(67),cout=>p(273)(68));
FA_ff_8999:FAff port map(x=>p(214)(68),y=>p(215)(68),Cin=>p(216)(68),clock=>clock,reset=>reset,s=>p(272)(68),cout=>p(273)(69));
FA_ff_9000:FAff port map(x=>p(214)(69),y=>p(215)(69),Cin=>p(216)(69),clock=>clock,reset=>reset,s=>p(272)(69),cout=>p(273)(70));
FA_ff_9001:FAff port map(x=>p(214)(70),y=>p(215)(70),Cin=>p(216)(70),clock=>clock,reset=>reset,s=>p(272)(70),cout=>p(273)(71));
FA_ff_9002:FAff port map(x=>p(214)(71),y=>p(215)(71),Cin=>p(216)(71),clock=>clock,reset=>reset,s=>p(272)(71),cout=>p(273)(72));
FA_ff_9003:FAff port map(x=>p(214)(72),y=>p(215)(72),Cin=>p(216)(72),clock=>clock,reset=>reset,s=>p(272)(72),cout=>p(273)(73));
FA_ff_9004:FAff port map(x=>p(214)(73),y=>p(215)(73),Cin=>p(216)(73),clock=>clock,reset=>reset,s=>p(272)(73),cout=>p(273)(74));
FA_ff_9005:FAff port map(x=>p(214)(74),y=>p(215)(74),Cin=>p(216)(74),clock=>clock,reset=>reset,s=>p(272)(74),cout=>p(273)(75));
FA_ff_9006:FAff port map(x=>p(214)(75),y=>p(215)(75),Cin=>p(216)(75),clock=>clock,reset=>reset,s=>p(272)(75),cout=>p(273)(76));
FA_ff_9007:FAff port map(x=>p(214)(76),y=>p(215)(76),Cin=>p(216)(76),clock=>clock,reset=>reset,s=>p(272)(76),cout=>p(273)(77));
FA_ff_9008:FAff port map(x=>p(214)(77),y=>p(215)(77),Cin=>p(216)(77),clock=>clock,reset=>reset,s=>p(272)(77),cout=>p(273)(78));
FA_ff_9009:FAff port map(x=>p(214)(78),y=>p(215)(78),Cin=>p(216)(78),clock=>clock,reset=>reset,s=>p(272)(78),cout=>p(273)(79));
FA_ff_9010:FAff port map(x=>p(214)(79),y=>p(215)(79),Cin=>p(216)(79),clock=>clock,reset=>reset,s=>p(272)(79),cout=>p(273)(80));
FA_ff_9011:FAff port map(x=>p(214)(80),y=>p(215)(80),Cin=>p(216)(80),clock=>clock,reset=>reset,s=>p(272)(80),cout=>p(273)(81));
FA_ff_9012:FAff port map(x=>p(214)(81),y=>p(215)(81),Cin=>p(216)(81),clock=>clock,reset=>reset,s=>p(272)(81),cout=>p(273)(82));
FA_ff_9013:FAff port map(x=>p(214)(82),y=>p(215)(82),Cin=>p(216)(82),clock=>clock,reset=>reset,s=>p(272)(82),cout=>p(273)(83));
FA_ff_9014:FAff port map(x=>p(214)(83),y=>p(215)(83),Cin=>p(216)(83),clock=>clock,reset=>reset,s=>p(272)(83),cout=>p(273)(84));
FA_ff_9015:FAff port map(x=>p(214)(84),y=>p(215)(84),Cin=>p(216)(84),clock=>clock,reset=>reset,s=>p(272)(84),cout=>p(273)(85));
FA_ff_9016:FAff port map(x=>p(214)(85),y=>p(215)(85),Cin=>p(216)(85),clock=>clock,reset=>reset,s=>p(272)(85),cout=>p(273)(86));
FA_ff_9017:FAff port map(x=>p(214)(86),y=>p(215)(86),Cin=>p(216)(86),clock=>clock,reset=>reset,s=>p(272)(86),cout=>p(273)(87));
FA_ff_9018:FAff port map(x=>p(214)(87),y=>p(215)(87),Cin=>p(216)(87),clock=>clock,reset=>reset,s=>p(272)(87),cout=>p(273)(88));
FA_ff_9019:FAff port map(x=>p(214)(88),y=>p(215)(88),Cin=>p(216)(88),clock=>clock,reset=>reset,s=>p(272)(88),cout=>p(273)(89));
FA_ff_9020:FAff port map(x=>p(214)(89),y=>p(215)(89),Cin=>p(216)(89),clock=>clock,reset=>reset,s=>p(272)(89),cout=>p(273)(90));
FA_ff_9021:FAff port map(x=>p(214)(90),y=>p(215)(90),Cin=>p(216)(90),clock=>clock,reset=>reset,s=>p(272)(90),cout=>p(273)(91));
FA_ff_9022:FAff port map(x=>p(214)(91),y=>p(215)(91),Cin=>p(216)(91),clock=>clock,reset=>reset,s=>p(272)(91),cout=>p(273)(92));
FA_ff_9023:FAff port map(x=>p(214)(92),y=>p(215)(92),Cin=>p(216)(92),clock=>clock,reset=>reset,s=>p(272)(92),cout=>p(273)(93));
FA_ff_9024:FAff port map(x=>p(214)(93),y=>p(215)(93),Cin=>p(216)(93),clock=>clock,reset=>reset,s=>p(272)(93),cout=>p(273)(94));
FA_ff_9025:FAff port map(x=>p(214)(94),y=>p(215)(94),Cin=>p(216)(94),clock=>clock,reset=>reset,s=>p(272)(94),cout=>p(273)(95));
FA_ff_9026:FAff port map(x=>p(214)(95),y=>p(215)(95),Cin=>p(216)(95),clock=>clock,reset=>reset,s=>p(272)(95),cout=>p(273)(96));
FA_ff_9027:FAff port map(x=>p(214)(96),y=>p(215)(96),Cin=>p(216)(96),clock=>clock,reset=>reset,s=>p(272)(96),cout=>p(273)(97));
FA_ff_9028:FAff port map(x=>p(214)(97),y=>p(215)(97),Cin=>p(216)(97),clock=>clock,reset=>reset,s=>p(272)(97),cout=>p(273)(98));
FA_ff_9029:FAff port map(x=>p(214)(98),y=>p(215)(98),Cin=>p(216)(98),clock=>clock,reset=>reset,s=>p(272)(98),cout=>p(273)(99));
FA_ff_9030:FAff port map(x=>p(214)(99),y=>p(215)(99),Cin=>p(216)(99),clock=>clock,reset=>reset,s=>p(272)(99),cout=>p(273)(100));
FA_ff_9031:FAff port map(x=>p(214)(100),y=>p(215)(100),Cin=>p(216)(100),clock=>clock,reset=>reset,s=>p(272)(100),cout=>p(273)(101));
FA_ff_9032:FAff port map(x=>p(214)(101),y=>p(215)(101),Cin=>p(216)(101),clock=>clock,reset=>reset,s=>p(272)(101),cout=>p(273)(102));
FA_ff_9033:FAff port map(x=>p(214)(102),y=>p(215)(102),Cin=>p(216)(102),clock=>clock,reset=>reset,s=>p(272)(102),cout=>p(273)(103));
FA_ff_9034:FAff port map(x=>p(214)(103),y=>p(215)(103),Cin=>p(216)(103),clock=>clock,reset=>reset,s=>p(272)(103),cout=>p(273)(104));
FA_ff_9035:FAff port map(x=>p(214)(104),y=>p(215)(104),Cin=>p(216)(104),clock=>clock,reset=>reset,s=>p(272)(104),cout=>p(273)(105));
FA_ff_9036:FAff port map(x=>p(214)(105),y=>p(215)(105),Cin=>p(216)(105),clock=>clock,reset=>reset,s=>p(272)(105),cout=>p(273)(106));
FA_ff_9037:FAff port map(x=>p(214)(106),y=>p(215)(106),Cin=>p(216)(106),clock=>clock,reset=>reset,s=>p(272)(106),cout=>p(273)(107));
FA_ff_9038:FAff port map(x=>p(214)(107),y=>p(215)(107),Cin=>p(216)(107),clock=>clock,reset=>reset,s=>p(272)(107),cout=>p(273)(108));
FA_ff_9039:FAff port map(x=>p(214)(108),y=>p(215)(108),Cin=>p(216)(108),clock=>clock,reset=>reset,s=>p(272)(108),cout=>p(273)(109));
FA_ff_9040:FAff port map(x=>p(214)(109),y=>p(215)(109),Cin=>p(216)(109),clock=>clock,reset=>reset,s=>p(272)(109),cout=>p(273)(110));
FA_ff_9041:FAff port map(x=>p(214)(110),y=>p(215)(110),Cin=>p(216)(110),clock=>clock,reset=>reset,s=>p(272)(110),cout=>p(273)(111));
FA_ff_9042:FAff port map(x=>p(214)(111),y=>p(215)(111),Cin=>p(216)(111),clock=>clock,reset=>reset,s=>p(272)(111),cout=>p(273)(112));
FA_ff_9043:FAff port map(x=>p(214)(112),y=>p(215)(112),Cin=>p(216)(112),clock=>clock,reset=>reset,s=>p(272)(112),cout=>p(273)(113));
FA_ff_9044:FAff port map(x=>p(214)(113),y=>p(215)(113),Cin=>p(216)(113),clock=>clock,reset=>reset,s=>p(272)(113),cout=>p(273)(114));
FA_ff_9045:FAff port map(x=>p(214)(114),y=>p(215)(114),Cin=>p(216)(114),clock=>clock,reset=>reset,s=>p(272)(114),cout=>p(273)(115));
FA_ff_9046:FAff port map(x=>p(214)(115),y=>p(215)(115),Cin=>p(216)(115),clock=>clock,reset=>reset,s=>p(272)(115),cout=>p(273)(116));
FA_ff_9047:FAff port map(x=>p(214)(116),y=>p(215)(116),Cin=>p(216)(116),clock=>clock,reset=>reset,s=>p(272)(116),cout=>p(273)(117));
FA_ff_9048:FAff port map(x=>p(214)(117),y=>p(215)(117),Cin=>p(216)(117),clock=>clock,reset=>reset,s=>p(272)(117),cout=>p(273)(118));
FA_ff_9049:FAff port map(x=>p(214)(118),y=>p(215)(118),Cin=>p(216)(118),clock=>clock,reset=>reset,s=>p(272)(118),cout=>p(273)(119));
FA_ff_9050:FAff port map(x=>p(214)(119),y=>p(215)(119),Cin=>p(216)(119),clock=>clock,reset=>reset,s=>p(272)(119),cout=>p(273)(120));
FA_ff_9051:FAff port map(x=>p(214)(120),y=>p(215)(120),Cin=>p(216)(120),clock=>clock,reset=>reset,s=>p(272)(120),cout=>p(273)(121));
FA_ff_9052:FAff port map(x=>p(214)(121),y=>p(215)(121),Cin=>p(216)(121),clock=>clock,reset=>reset,s=>p(272)(121),cout=>p(273)(122));
FA_ff_9053:FAff port map(x=>p(214)(122),y=>p(215)(122),Cin=>p(216)(122),clock=>clock,reset=>reset,s=>p(272)(122),cout=>p(273)(123));
FA_ff_9054:FAff port map(x=>p(214)(123),y=>p(215)(123),Cin=>p(216)(123),clock=>clock,reset=>reset,s=>p(272)(123),cout=>p(273)(124));
FA_ff_9055:FAff port map(x=>p(214)(124),y=>p(215)(124),Cin=>p(216)(124),clock=>clock,reset=>reset,s=>p(272)(124),cout=>p(273)(125));
FA_ff_9056:FAff port map(x=>p(214)(125),y=>p(215)(125),Cin=>p(216)(125),clock=>clock,reset=>reset,s=>p(272)(125),cout=>p(273)(126));
FA_ff_9057:FAff port map(x=>p(214)(126),y=>p(215)(126),Cin=>p(216)(126),clock=>clock,reset=>reset,s=>p(272)(126),cout=>p(273)(127));
FA_ff_9058:FAff port map(x=>p(214)(127),y=>p(215)(127),Cin=>p(216)(127),clock=>clock,reset=>reset,s=>p(272)(127),cout=>p(273)(128));
FA_ff_9059:FAff port map(x=>p(214)(128),y=>p(215)(128),Cin=>p(216)(128),clock=>clock,reset=>reset,s=>p(272)(128),cout=>p(273)(129));
p(274)(0)<=p(218)(0);
HA_ff_29:HAff port map(x=>p(218)(1),y=>p(219)(1),clock=>clock,reset=>reset,s=>p(274)(1),c=>p(275)(2));
FA_ff_9060:FAff port map(x=>p(217)(2),y=>p(218)(2),Cin=>p(219)(2),clock=>clock,reset=>reset,s=>p(274)(2),cout=>p(275)(3));
FA_ff_9061:FAff port map(x=>p(217)(3),y=>p(218)(3),Cin=>p(219)(3),clock=>clock,reset=>reset,s=>p(274)(3),cout=>p(275)(4));
FA_ff_9062:FAff port map(x=>p(217)(4),y=>p(218)(4),Cin=>p(219)(4),clock=>clock,reset=>reset,s=>p(274)(4),cout=>p(275)(5));
FA_ff_9063:FAff port map(x=>p(217)(5),y=>p(218)(5),Cin=>p(219)(5),clock=>clock,reset=>reset,s=>p(274)(5),cout=>p(275)(6));
FA_ff_9064:FAff port map(x=>p(217)(6),y=>p(218)(6),Cin=>p(219)(6),clock=>clock,reset=>reset,s=>p(274)(6),cout=>p(275)(7));
FA_ff_9065:FAff port map(x=>p(217)(7),y=>p(218)(7),Cin=>p(219)(7),clock=>clock,reset=>reset,s=>p(274)(7),cout=>p(275)(8));
FA_ff_9066:FAff port map(x=>p(217)(8),y=>p(218)(8),Cin=>p(219)(8),clock=>clock,reset=>reset,s=>p(274)(8),cout=>p(275)(9));
FA_ff_9067:FAff port map(x=>p(217)(9),y=>p(218)(9),Cin=>p(219)(9),clock=>clock,reset=>reset,s=>p(274)(9),cout=>p(275)(10));
FA_ff_9068:FAff port map(x=>p(217)(10),y=>p(218)(10),Cin=>p(219)(10),clock=>clock,reset=>reset,s=>p(274)(10),cout=>p(275)(11));
FA_ff_9069:FAff port map(x=>p(217)(11),y=>p(218)(11),Cin=>p(219)(11),clock=>clock,reset=>reset,s=>p(274)(11),cout=>p(275)(12));
FA_ff_9070:FAff port map(x=>p(217)(12),y=>p(218)(12),Cin=>p(219)(12),clock=>clock,reset=>reset,s=>p(274)(12),cout=>p(275)(13));
FA_ff_9071:FAff port map(x=>p(217)(13),y=>p(218)(13),Cin=>p(219)(13),clock=>clock,reset=>reset,s=>p(274)(13),cout=>p(275)(14));
FA_ff_9072:FAff port map(x=>p(217)(14),y=>p(218)(14),Cin=>p(219)(14),clock=>clock,reset=>reset,s=>p(274)(14),cout=>p(275)(15));
FA_ff_9073:FAff port map(x=>p(217)(15),y=>p(218)(15),Cin=>p(219)(15),clock=>clock,reset=>reset,s=>p(274)(15),cout=>p(275)(16));
FA_ff_9074:FAff port map(x=>p(217)(16),y=>p(218)(16),Cin=>p(219)(16),clock=>clock,reset=>reset,s=>p(274)(16),cout=>p(275)(17));
FA_ff_9075:FAff port map(x=>p(217)(17),y=>p(218)(17),Cin=>p(219)(17),clock=>clock,reset=>reset,s=>p(274)(17),cout=>p(275)(18));
FA_ff_9076:FAff port map(x=>p(217)(18),y=>p(218)(18),Cin=>p(219)(18),clock=>clock,reset=>reset,s=>p(274)(18),cout=>p(275)(19));
FA_ff_9077:FAff port map(x=>p(217)(19),y=>p(218)(19),Cin=>p(219)(19),clock=>clock,reset=>reset,s=>p(274)(19),cout=>p(275)(20));
FA_ff_9078:FAff port map(x=>p(217)(20),y=>p(218)(20),Cin=>p(219)(20),clock=>clock,reset=>reset,s=>p(274)(20),cout=>p(275)(21));
FA_ff_9079:FAff port map(x=>p(217)(21),y=>p(218)(21),Cin=>p(219)(21),clock=>clock,reset=>reset,s=>p(274)(21),cout=>p(275)(22));
FA_ff_9080:FAff port map(x=>p(217)(22),y=>p(218)(22),Cin=>p(219)(22),clock=>clock,reset=>reset,s=>p(274)(22),cout=>p(275)(23));
FA_ff_9081:FAff port map(x=>p(217)(23),y=>p(218)(23),Cin=>p(219)(23),clock=>clock,reset=>reset,s=>p(274)(23),cout=>p(275)(24));
FA_ff_9082:FAff port map(x=>p(217)(24),y=>p(218)(24),Cin=>p(219)(24),clock=>clock,reset=>reset,s=>p(274)(24),cout=>p(275)(25));
FA_ff_9083:FAff port map(x=>p(217)(25),y=>p(218)(25),Cin=>p(219)(25),clock=>clock,reset=>reset,s=>p(274)(25),cout=>p(275)(26));
FA_ff_9084:FAff port map(x=>p(217)(26),y=>p(218)(26),Cin=>p(219)(26),clock=>clock,reset=>reset,s=>p(274)(26),cout=>p(275)(27));
FA_ff_9085:FAff port map(x=>p(217)(27),y=>p(218)(27),Cin=>p(219)(27),clock=>clock,reset=>reset,s=>p(274)(27),cout=>p(275)(28));
FA_ff_9086:FAff port map(x=>p(217)(28),y=>p(218)(28),Cin=>p(219)(28),clock=>clock,reset=>reset,s=>p(274)(28),cout=>p(275)(29));
FA_ff_9087:FAff port map(x=>p(217)(29),y=>p(218)(29),Cin=>p(219)(29),clock=>clock,reset=>reset,s=>p(274)(29),cout=>p(275)(30));
FA_ff_9088:FAff port map(x=>p(217)(30),y=>p(218)(30),Cin=>p(219)(30),clock=>clock,reset=>reset,s=>p(274)(30),cout=>p(275)(31));
FA_ff_9089:FAff port map(x=>p(217)(31),y=>p(218)(31),Cin=>p(219)(31),clock=>clock,reset=>reset,s=>p(274)(31),cout=>p(275)(32));
FA_ff_9090:FAff port map(x=>p(217)(32),y=>p(218)(32),Cin=>p(219)(32),clock=>clock,reset=>reset,s=>p(274)(32),cout=>p(275)(33));
FA_ff_9091:FAff port map(x=>p(217)(33),y=>p(218)(33),Cin=>p(219)(33),clock=>clock,reset=>reset,s=>p(274)(33),cout=>p(275)(34));
FA_ff_9092:FAff port map(x=>p(217)(34),y=>p(218)(34),Cin=>p(219)(34),clock=>clock,reset=>reset,s=>p(274)(34),cout=>p(275)(35));
FA_ff_9093:FAff port map(x=>p(217)(35),y=>p(218)(35),Cin=>p(219)(35),clock=>clock,reset=>reset,s=>p(274)(35),cout=>p(275)(36));
FA_ff_9094:FAff port map(x=>p(217)(36),y=>p(218)(36),Cin=>p(219)(36),clock=>clock,reset=>reset,s=>p(274)(36),cout=>p(275)(37));
FA_ff_9095:FAff port map(x=>p(217)(37),y=>p(218)(37),Cin=>p(219)(37),clock=>clock,reset=>reset,s=>p(274)(37),cout=>p(275)(38));
FA_ff_9096:FAff port map(x=>p(217)(38),y=>p(218)(38),Cin=>p(219)(38),clock=>clock,reset=>reset,s=>p(274)(38),cout=>p(275)(39));
FA_ff_9097:FAff port map(x=>p(217)(39),y=>p(218)(39),Cin=>p(219)(39),clock=>clock,reset=>reset,s=>p(274)(39),cout=>p(275)(40));
FA_ff_9098:FAff port map(x=>p(217)(40),y=>p(218)(40),Cin=>p(219)(40),clock=>clock,reset=>reset,s=>p(274)(40),cout=>p(275)(41));
FA_ff_9099:FAff port map(x=>p(217)(41),y=>p(218)(41),Cin=>p(219)(41),clock=>clock,reset=>reset,s=>p(274)(41),cout=>p(275)(42));
FA_ff_9100:FAff port map(x=>p(217)(42),y=>p(218)(42),Cin=>p(219)(42),clock=>clock,reset=>reset,s=>p(274)(42),cout=>p(275)(43));
FA_ff_9101:FAff port map(x=>p(217)(43),y=>p(218)(43),Cin=>p(219)(43),clock=>clock,reset=>reset,s=>p(274)(43),cout=>p(275)(44));
FA_ff_9102:FAff port map(x=>p(217)(44),y=>p(218)(44),Cin=>p(219)(44),clock=>clock,reset=>reset,s=>p(274)(44),cout=>p(275)(45));
FA_ff_9103:FAff port map(x=>p(217)(45),y=>p(218)(45),Cin=>p(219)(45),clock=>clock,reset=>reset,s=>p(274)(45),cout=>p(275)(46));
FA_ff_9104:FAff port map(x=>p(217)(46),y=>p(218)(46),Cin=>p(219)(46),clock=>clock,reset=>reset,s=>p(274)(46),cout=>p(275)(47));
FA_ff_9105:FAff port map(x=>p(217)(47),y=>p(218)(47),Cin=>p(219)(47),clock=>clock,reset=>reset,s=>p(274)(47),cout=>p(275)(48));
FA_ff_9106:FAff port map(x=>p(217)(48),y=>p(218)(48),Cin=>p(219)(48),clock=>clock,reset=>reset,s=>p(274)(48),cout=>p(275)(49));
FA_ff_9107:FAff port map(x=>p(217)(49),y=>p(218)(49),Cin=>p(219)(49),clock=>clock,reset=>reset,s=>p(274)(49),cout=>p(275)(50));
FA_ff_9108:FAff port map(x=>p(217)(50),y=>p(218)(50),Cin=>p(219)(50),clock=>clock,reset=>reset,s=>p(274)(50),cout=>p(275)(51));
FA_ff_9109:FAff port map(x=>p(217)(51),y=>p(218)(51),Cin=>p(219)(51),clock=>clock,reset=>reset,s=>p(274)(51),cout=>p(275)(52));
FA_ff_9110:FAff port map(x=>p(217)(52),y=>p(218)(52),Cin=>p(219)(52),clock=>clock,reset=>reset,s=>p(274)(52),cout=>p(275)(53));
FA_ff_9111:FAff port map(x=>p(217)(53),y=>p(218)(53),Cin=>p(219)(53),clock=>clock,reset=>reset,s=>p(274)(53),cout=>p(275)(54));
FA_ff_9112:FAff port map(x=>p(217)(54),y=>p(218)(54),Cin=>p(219)(54),clock=>clock,reset=>reset,s=>p(274)(54),cout=>p(275)(55));
FA_ff_9113:FAff port map(x=>p(217)(55),y=>p(218)(55),Cin=>p(219)(55),clock=>clock,reset=>reset,s=>p(274)(55),cout=>p(275)(56));
FA_ff_9114:FAff port map(x=>p(217)(56),y=>p(218)(56),Cin=>p(219)(56),clock=>clock,reset=>reset,s=>p(274)(56),cout=>p(275)(57));
FA_ff_9115:FAff port map(x=>p(217)(57),y=>p(218)(57),Cin=>p(219)(57),clock=>clock,reset=>reset,s=>p(274)(57),cout=>p(275)(58));
FA_ff_9116:FAff port map(x=>p(217)(58),y=>p(218)(58),Cin=>p(219)(58),clock=>clock,reset=>reset,s=>p(274)(58),cout=>p(275)(59));
FA_ff_9117:FAff port map(x=>p(217)(59),y=>p(218)(59),Cin=>p(219)(59),clock=>clock,reset=>reset,s=>p(274)(59),cout=>p(275)(60));
FA_ff_9118:FAff port map(x=>p(217)(60),y=>p(218)(60),Cin=>p(219)(60),clock=>clock,reset=>reset,s=>p(274)(60),cout=>p(275)(61));
FA_ff_9119:FAff port map(x=>p(217)(61),y=>p(218)(61),Cin=>p(219)(61),clock=>clock,reset=>reset,s=>p(274)(61),cout=>p(275)(62));
FA_ff_9120:FAff port map(x=>p(217)(62),y=>p(218)(62),Cin=>p(219)(62),clock=>clock,reset=>reset,s=>p(274)(62),cout=>p(275)(63));
FA_ff_9121:FAff port map(x=>p(217)(63),y=>p(218)(63),Cin=>p(219)(63),clock=>clock,reset=>reset,s=>p(274)(63),cout=>p(275)(64));
FA_ff_9122:FAff port map(x=>p(217)(64),y=>p(218)(64),Cin=>p(219)(64),clock=>clock,reset=>reset,s=>p(274)(64),cout=>p(275)(65));
FA_ff_9123:FAff port map(x=>p(217)(65),y=>p(218)(65),Cin=>p(219)(65),clock=>clock,reset=>reset,s=>p(274)(65),cout=>p(275)(66));
FA_ff_9124:FAff port map(x=>p(217)(66),y=>p(218)(66),Cin=>p(219)(66),clock=>clock,reset=>reset,s=>p(274)(66),cout=>p(275)(67));
FA_ff_9125:FAff port map(x=>p(217)(67),y=>p(218)(67),Cin=>p(219)(67),clock=>clock,reset=>reset,s=>p(274)(67),cout=>p(275)(68));
FA_ff_9126:FAff port map(x=>p(217)(68),y=>p(218)(68),Cin=>p(219)(68),clock=>clock,reset=>reset,s=>p(274)(68),cout=>p(275)(69));
FA_ff_9127:FAff port map(x=>p(217)(69),y=>p(218)(69),Cin=>p(219)(69),clock=>clock,reset=>reset,s=>p(274)(69),cout=>p(275)(70));
FA_ff_9128:FAff port map(x=>p(217)(70),y=>p(218)(70),Cin=>p(219)(70),clock=>clock,reset=>reset,s=>p(274)(70),cout=>p(275)(71));
FA_ff_9129:FAff port map(x=>p(217)(71),y=>p(218)(71),Cin=>p(219)(71),clock=>clock,reset=>reset,s=>p(274)(71),cout=>p(275)(72));
FA_ff_9130:FAff port map(x=>p(217)(72),y=>p(218)(72),Cin=>p(219)(72),clock=>clock,reset=>reset,s=>p(274)(72),cout=>p(275)(73));
FA_ff_9131:FAff port map(x=>p(217)(73),y=>p(218)(73),Cin=>p(219)(73),clock=>clock,reset=>reset,s=>p(274)(73),cout=>p(275)(74));
FA_ff_9132:FAff port map(x=>p(217)(74),y=>p(218)(74),Cin=>p(219)(74),clock=>clock,reset=>reset,s=>p(274)(74),cout=>p(275)(75));
FA_ff_9133:FAff port map(x=>p(217)(75),y=>p(218)(75),Cin=>p(219)(75),clock=>clock,reset=>reset,s=>p(274)(75),cout=>p(275)(76));
FA_ff_9134:FAff port map(x=>p(217)(76),y=>p(218)(76),Cin=>p(219)(76),clock=>clock,reset=>reset,s=>p(274)(76),cout=>p(275)(77));
FA_ff_9135:FAff port map(x=>p(217)(77),y=>p(218)(77),Cin=>p(219)(77),clock=>clock,reset=>reset,s=>p(274)(77),cout=>p(275)(78));
FA_ff_9136:FAff port map(x=>p(217)(78),y=>p(218)(78),Cin=>p(219)(78),clock=>clock,reset=>reset,s=>p(274)(78),cout=>p(275)(79));
FA_ff_9137:FAff port map(x=>p(217)(79),y=>p(218)(79),Cin=>p(219)(79),clock=>clock,reset=>reset,s=>p(274)(79),cout=>p(275)(80));
FA_ff_9138:FAff port map(x=>p(217)(80),y=>p(218)(80),Cin=>p(219)(80),clock=>clock,reset=>reset,s=>p(274)(80),cout=>p(275)(81));
FA_ff_9139:FAff port map(x=>p(217)(81),y=>p(218)(81),Cin=>p(219)(81),clock=>clock,reset=>reset,s=>p(274)(81),cout=>p(275)(82));
FA_ff_9140:FAff port map(x=>p(217)(82),y=>p(218)(82),Cin=>p(219)(82),clock=>clock,reset=>reset,s=>p(274)(82),cout=>p(275)(83));
FA_ff_9141:FAff port map(x=>p(217)(83),y=>p(218)(83),Cin=>p(219)(83),clock=>clock,reset=>reset,s=>p(274)(83),cout=>p(275)(84));
FA_ff_9142:FAff port map(x=>p(217)(84),y=>p(218)(84),Cin=>p(219)(84),clock=>clock,reset=>reset,s=>p(274)(84),cout=>p(275)(85));
FA_ff_9143:FAff port map(x=>p(217)(85),y=>p(218)(85),Cin=>p(219)(85),clock=>clock,reset=>reset,s=>p(274)(85),cout=>p(275)(86));
FA_ff_9144:FAff port map(x=>p(217)(86),y=>p(218)(86),Cin=>p(219)(86),clock=>clock,reset=>reset,s=>p(274)(86),cout=>p(275)(87));
FA_ff_9145:FAff port map(x=>p(217)(87),y=>p(218)(87),Cin=>p(219)(87),clock=>clock,reset=>reset,s=>p(274)(87),cout=>p(275)(88));
FA_ff_9146:FAff port map(x=>p(217)(88),y=>p(218)(88),Cin=>p(219)(88),clock=>clock,reset=>reset,s=>p(274)(88),cout=>p(275)(89));
FA_ff_9147:FAff port map(x=>p(217)(89),y=>p(218)(89),Cin=>p(219)(89),clock=>clock,reset=>reset,s=>p(274)(89),cout=>p(275)(90));
FA_ff_9148:FAff port map(x=>p(217)(90),y=>p(218)(90),Cin=>p(219)(90),clock=>clock,reset=>reset,s=>p(274)(90),cout=>p(275)(91));
FA_ff_9149:FAff port map(x=>p(217)(91),y=>p(218)(91),Cin=>p(219)(91),clock=>clock,reset=>reset,s=>p(274)(91),cout=>p(275)(92));
FA_ff_9150:FAff port map(x=>p(217)(92),y=>p(218)(92),Cin=>p(219)(92),clock=>clock,reset=>reset,s=>p(274)(92),cout=>p(275)(93));
FA_ff_9151:FAff port map(x=>p(217)(93),y=>p(218)(93),Cin=>p(219)(93),clock=>clock,reset=>reset,s=>p(274)(93),cout=>p(275)(94));
FA_ff_9152:FAff port map(x=>p(217)(94),y=>p(218)(94),Cin=>p(219)(94),clock=>clock,reset=>reset,s=>p(274)(94),cout=>p(275)(95));
FA_ff_9153:FAff port map(x=>p(217)(95),y=>p(218)(95),Cin=>p(219)(95),clock=>clock,reset=>reset,s=>p(274)(95),cout=>p(275)(96));
FA_ff_9154:FAff port map(x=>p(217)(96),y=>p(218)(96),Cin=>p(219)(96),clock=>clock,reset=>reset,s=>p(274)(96),cout=>p(275)(97));
FA_ff_9155:FAff port map(x=>p(217)(97),y=>p(218)(97),Cin=>p(219)(97),clock=>clock,reset=>reset,s=>p(274)(97),cout=>p(275)(98));
FA_ff_9156:FAff port map(x=>p(217)(98),y=>p(218)(98),Cin=>p(219)(98),clock=>clock,reset=>reset,s=>p(274)(98),cout=>p(275)(99));
FA_ff_9157:FAff port map(x=>p(217)(99),y=>p(218)(99),Cin=>p(219)(99),clock=>clock,reset=>reset,s=>p(274)(99),cout=>p(275)(100));
FA_ff_9158:FAff port map(x=>p(217)(100),y=>p(218)(100),Cin=>p(219)(100),clock=>clock,reset=>reset,s=>p(274)(100),cout=>p(275)(101));
FA_ff_9159:FAff port map(x=>p(217)(101),y=>p(218)(101),Cin=>p(219)(101),clock=>clock,reset=>reset,s=>p(274)(101),cout=>p(275)(102));
FA_ff_9160:FAff port map(x=>p(217)(102),y=>p(218)(102),Cin=>p(219)(102),clock=>clock,reset=>reset,s=>p(274)(102),cout=>p(275)(103));
FA_ff_9161:FAff port map(x=>p(217)(103),y=>p(218)(103),Cin=>p(219)(103),clock=>clock,reset=>reset,s=>p(274)(103),cout=>p(275)(104));
FA_ff_9162:FAff port map(x=>p(217)(104),y=>p(218)(104),Cin=>p(219)(104),clock=>clock,reset=>reset,s=>p(274)(104),cout=>p(275)(105));
FA_ff_9163:FAff port map(x=>p(217)(105),y=>p(218)(105),Cin=>p(219)(105),clock=>clock,reset=>reset,s=>p(274)(105),cout=>p(275)(106));
FA_ff_9164:FAff port map(x=>p(217)(106),y=>p(218)(106),Cin=>p(219)(106),clock=>clock,reset=>reset,s=>p(274)(106),cout=>p(275)(107));
FA_ff_9165:FAff port map(x=>p(217)(107),y=>p(218)(107),Cin=>p(219)(107),clock=>clock,reset=>reset,s=>p(274)(107),cout=>p(275)(108));
FA_ff_9166:FAff port map(x=>p(217)(108),y=>p(218)(108),Cin=>p(219)(108),clock=>clock,reset=>reset,s=>p(274)(108),cout=>p(275)(109));
FA_ff_9167:FAff port map(x=>p(217)(109),y=>p(218)(109),Cin=>p(219)(109),clock=>clock,reset=>reset,s=>p(274)(109),cout=>p(275)(110));
FA_ff_9168:FAff port map(x=>p(217)(110),y=>p(218)(110),Cin=>p(219)(110),clock=>clock,reset=>reset,s=>p(274)(110),cout=>p(275)(111));
FA_ff_9169:FAff port map(x=>p(217)(111),y=>p(218)(111),Cin=>p(219)(111),clock=>clock,reset=>reset,s=>p(274)(111),cout=>p(275)(112));
FA_ff_9170:FAff port map(x=>p(217)(112),y=>p(218)(112),Cin=>p(219)(112),clock=>clock,reset=>reset,s=>p(274)(112),cout=>p(275)(113));
FA_ff_9171:FAff port map(x=>p(217)(113),y=>p(218)(113),Cin=>p(219)(113),clock=>clock,reset=>reset,s=>p(274)(113),cout=>p(275)(114));
FA_ff_9172:FAff port map(x=>p(217)(114),y=>p(218)(114),Cin=>p(219)(114),clock=>clock,reset=>reset,s=>p(274)(114),cout=>p(275)(115));
FA_ff_9173:FAff port map(x=>p(217)(115),y=>p(218)(115),Cin=>p(219)(115),clock=>clock,reset=>reset,s=>p(274)(115),cout=>p(275)(116));
FA_ff_9174:FAff port map(x=>p(217)(116),y=>p(218)(116),Cin=>p(219)(116),clock=>clock,reset=>reset,s=>p(274)(116),cout=>p(275)(117));
FA_ff_9175:FAff port map(x=>p(217)(117),y=>p(218)(117),Cin=>p(219)(117),clock=>clock,reset=>reset,s=>p(274)(117),cout=>p(275)(118));
FA_ff_9176:FAff port map(x=>p(217)(118),y=>p(218)(118),Cin=>p(219)(118),clock=>clock,reset=>reset,s=>p(274)(118),cout=>p(275)(119));
FA_ff_9177:FAff port map(x=>p(217)(119),y=>p(218)(119),Cin=>p(219)(119),clock=>clock,reset=>reset,s=>p(274)(119),cout=>p(275)(120));
FA_ff_9178:FAff port map(x=>p(217)(120),y=>p(218)(120),Cin=>p(219)(120),clock=>clock,reset=>reset,s=>p(274)(120),cout=>p(275)(121));
FA_ff_9179:FAff port map(x=>p(217)(121),y=>p(218)(121),Cin=>p(219)(121),clock=>clock,reset=>reset,s=>p(274)(121),cout=>p(275)(122));
FA_ff_9180:FAff port map(x=>p(217)(122),y=>p(218)(122),Cin=>p(219)(122),clock=>clock,reset=>reset,s=>p(274)(122),cout=>p(275)(123));
FA_ff_9181:FAff port map(x=>p(217)(123),y=>p(218)(123),Cin=>p(219)(123),clock=>clock,reset=>reset,s=>p(274)(123),cout=>p(275)(124));
FA_ff_9182:FAff port map(x=>p(217)(124),y=>p(218)(124),Cin=>p(219)(124),clock=>clock,reset=>reset,s=>p(274)(124),cout=>p(275)(125));
FA_ff_9183:FAff port map(x=>p(217)(125),y=>p(218)(125),Cin=>p(219)(125),clock=>clock,reset=>reset,s=>p(274)(125),cout=>p(275)(126));
FA_ff_9184:FAff port map(x=>p(217)(126),y=>p(218)(126),Cin=>p(219)(126),clock=>clock,reset=>reset,s=>p(274)(126),cout=>p(275)(127));
FA_ff_9185:FAff port map(x=>p(217)(127),y=>p(218)(127),Cin=>p(219)(127),clock=>clock,reset=>reset,s=>p(274)(127),cout=>p(275)(128));
FA_ff_9186:FAff port map(x=>p(217)(128),y=>p(218)(128),Cin=>p(219)(128),clock=>clock,reset=>reset,s=>p(274)(128),cout=>p(275)(129));
p(274)(129)<=p(217)(129);
HA_ff_30:HAff port map(x=>p(220)(0),y=>p(222)(0),clock=>clock,reset=>reset,s=>p(276)(0),c=>p(277)(1));
HA_ff_31:HAff port map(x=>p(220)(1),y=>p(222)(1),clock=>clock,reset=>reset,s=>p(276)(1),c=>p(277)(2));
FA_ff_9187:FAff port map(x=>p(220)(2),y=>p(221)(2),Cin=>p(222)(2),clock=>clock,reset=>reset,s=>p(276)(2),cout=>p(277)(3));
FA_ff_9188:FAff port map(x=>p(220)(3),y=>p(221)(3),Cin=>p(222)(3),clock=>clock,reset=>reset,s=>p(276)(3),cout=>p(277)(4));
FA_ff_9189:FAff port map(x=>p(220)(4),y=>p(221)(4),Cin=>p(222)(4),clock=>clock,reset=>reset,s=>p(276)(4),cout=>p(277)(5));
FA_ff_9190:FAff port map(x=>p(220)(5),y=>p(221)(5),Cin=>p(222)(5),clock=>clock,reset=>reset,s=>p(276)(5),cout=>p(277)(6));
FA_ff_9191:FAff port map(x=>p(220)(6),y=>p(221)(6),Cin=>p(222)(6),clock=>clock,reset=>reset,s=>p(276)(6),cout=>p(277)(7));
FA_ff_9192:FAff port map(x=>p(220)(7),y=>p(221)(7),Cin=>p(222)(7),clock=>clock,reset=>reset,s=>p(276)(7),cout=>p(277)(8));
FA_ff_9193:FAff port map(x=>p(220)(8),y=>p(221)(8),Cin=>p(222)(8),clock=>clock,reset=>reset,s=>p(276)(8),cout=>p(277)(9));
FA_ff_9194:FAff port map(x=>p(220)(9),y=>p(221)(9),Cin=>p(222)(9),clock=>clock,reset=>reset,s=>p(276)(9),cout=>p(277)(10));
FA_ff_9195:FAff port map(x=>p(220)(10),y=>p(221)(10),Cin=>p(222)(10),clock=>clock,reset=>reset,s=>p(276)(10),cout=>p(277)(11));
FA_ff_9196:FAff port map(x=>p(220)(11),y=>p(221)(11),Cin=>p(222)(11),clock=>clock,reset=>reset,s=>p(276)(11),cout=>p(277)(12));
FA_ff_9197:FAff port map(x=>p(220)(12),y=>p(221)(12),Cin=>p(222)(12),clock=>clock,reset=>reset,s=>p(276)(12),cout=>p(277)(13));
FA_ff_9198:FAff port map(x=>p(220)(13),y=>p(221)(13),Cin=>p(222)(13),clock=>clock,reset=>reset,s=>p(276)(13),cout=>p(277)(14));
FA_ff_9199:FAff port map(x=>p(220)(14),y=>p(221)(14),Cin=>p(222)(14),clock=>clock,reset=>reset,s=>p(276)(14),cout=>p(277)(15));
FA_ff_9200:FAff port map(x=>p(220)(15),y=>p(221)(15),Cin=>p(222)(15),clock=>clock,reset=>reset,s=>p(276)(15),cout=>p(277)(16));
FA_ff_9201:FAff port map(x=>p(220)(16),y=>p(221)(16),Cin=>p(222)(16),clock=>clock,reset=>reset,s=>p(276)(16),cout=>p(277)(17));
FA_ff_9202:FAff port map(x=>p(220)(17),y=>p(221)(17),Cin=>p(222)(17),clock=>clock,reset=>reset,s=>p(276)(17),cout=>p(277)(18));
FA_ff_9203:FAff port map(x=>p(220)(18),y=>p(221)(18),Cin=>p(222)(18),clock=>clock,reset=>reset,s=>p(276)(18),cout=>p(277)(19));
FA_ff_9204:FAff port map(x=>p(220)(19),y=>p(221)(19),Cin=>p(222)(19),clock=>clock,reset=>reset,s=>p(276)(19),cout=>p(277)(20));
FA_ff_9205:FAff port map(x=>p(220)(20),y=>p(221)(20),Cin=>p(222)(20),clock=>clock,reset=>reset,s=>p(276)(20),cout=>p(277)(21));
FA_ff_9206:FAff port map(x=>p(220)(21),y=>p(221)(21),Cin=>p(222)(21),clock=>clock,reset=>reset,s=>p(276)(21),cout=>p(277)(22));
FA_ff_9207:FAff port map(x=>p(220)(22),y=>p(221)(22),Cin=>p(222)(22),clock=>clock,reset=>reset,s=>p(276)(22),cout=>p(277)(23));
FA_ff_9208:FAff port map(x=>p(220)(23),y=>p(221)(23),Cin=>p(222)(23),clock=>clock,reset=>reset,s=>p(276)(23),cout=>p(277)(24));
FA_ff_9209:FAff port map(x=>p(220)(24),y=>p(221)(24),Cin=>p(222)(24),clock=>clock,reset=>reset,s=>p(276)(24),cout=>p(277)(25));
FA_ff_9210:FAff port map(x=>p(220)(25),y=>p(221)(25),Cin=>p(222)(25),clock=>clock,reset=>reset,s=>p(276)(25),cout=>p(277)(26));
FA_ff_9211:FAff port map(x=>p(220)(26),y=>p(221)(26),Cin=>p(222)(26),clock=>clock,reset=>reset,s=>p(276)(26),cout=>p(277)(27));
FA_ff_9212:FAff port map(x=>p(220)(27),y=>p(221)(27),Cin=>p(222)(27),clock=>clock,reset=>reset,s=>p(276)(27),cout=>p(277)(28));
FA_ff_9213:FAff port map(x=>p(220)(28),y=>p(221)(28),Cin=>p(222)(28),clock=>clock,reset=>reset,s=>p(276)(28),cout=>p(277)(29));
FA_ff_9214:FAff port map(x=>p(220)(29),y=>p(221)(29),Cin=>p(222)(29),clock=>clock,reset=>reset,s=>p(276)(29),cout=>p(277)(30));
FA_ff_9215:FAff port map(x=>p(220)(30),y=>p(221)(30),Cin=>p(222)(30),clock=>clock,reset=>reset,s=>p(276)(30),cout=>p(277)(31));
FA_ff_9216:FAff port map(x=>p(220)(31),y=>p(221)(31),Cin=>p(222)(31),clock=>clock,reset=>reset,s=>p(276)(31),cout=>p(277)(32));
FA_ff_9217:FAff port map(x=>p(220)(32),y=>p(221)(32),Cin=>p(222)(32),clock=>clock,reset=>reset,s=>p(276)(32),cout=>p(277)(33));
FA_ff_9218:FAff port map(x=>p(220)(33),y=>p(221)(33),Cin=>p(222)(33),clock=>clock,reset=>reset,s=>p(276)(33),cout=>p(277)(34));
FA_ff_9219:FAff port map(x=>p(220)(34),y=>p(221)(34),Cin=>p(222)(34),clock=>clock,reset=>reset,s=>p(276)(34),cout=>p(277)(35));
FA_ff_9220:FAff port map(x=>p(220)(35),y=>p(221)(35),Cin=>p(222)(35),clock=>clock,reset=>reset,s=>p(276)(35),cout=>p(277)(36));
FA_ff_9221:FAff port map(x=>p(220)(36),y=>p(221)(36),Cin=>p(222)(36),clock=>clock,reset=>reset,s=>p(276)(36),cout=>p(277)(37));
FA_ff_9222:FAff port map(x=>p(220)(37),y=>p(221)(37),Cin=>p(222)(37),clock=>clock,reset=>reset,s=>p(276)(37),cout=>p(277)(38));
FA_ff_9223:FAff port map(x=>p(220)(38),y=>p(221)(38),Cin=>p(222)(38),clock=>clock,reset=>reset,s=>p(276)(38),cout=>p(277)(39));
FA_ff_9224:FAff port map(x=>p(220)(39),y=>p(221)(39),Cin=>p(222)(39),clock=>clock,reset=>reset,s=>p(276)(39),cout=>p(277)(40));
FA_ff_9225:FAff port map(x=>p(220)(40),y=>p(221)(40),Cin=>p(222)(40),clock=>clock,reset=>reset,s=>p(276)(40),cout=>p(277)(41));
FA_ff_9226:FAff port map(x=>p(220)(41),y=>p(221)(41),Cin=>p(222)(41),clock=>clock,reset=>reset,s=>p(276)(41),cout=>p(277)(42));
FA_ff_9227:FAff port map(x=>p(220)(42),y=>p(221)(42),Cin=>p(222)(42),clock=>clock,reset=>reset,s=>p(276)(42),cout=>p(277)(43));
FA_ff_9228:FAff port map(x=>p(220)(43),y=>p(221)(43),Cin=>p(222)(43),clock=>clock,reset=>reset,s=>p(276)(43),cout=>p(277)(44));
FA_ff_9229:FAff port map(x=>p(220)(44),y=>p(221)(44),Cin=>p(222)(44),clock=>clock,reset=>reset,s=>p(276)(44),cout=>p(277)(45));
FA_ff_9230:FAff port map(x=>p(220)(45),y=>p(221)(45),Cin=>p(222)(45),clock=>clock,reset=>reset,s=>p(276)(45),cout=>p(277)(46));
FA_ff_9231:FAff port map(x=>p(220)(46),y=>p(221)(46),Cin=>p(222)(46),clock=>clock,reset=>reset,s=>p(276)(46),cout=>p(277)(47));
FA_ff_9232:FAff port map(x=>p(220)(47),y=>p(221)(47),Cin=>p(222)(47),clock=>clock,reset=>reset,s=>p(276)(47),cout=>p(277)(48));
FA_ff_9233:FAff port map(x=>p(220)(48),y=>p(221)(48),Cin=>p(222)(48),clock=>clock,reset=>reset,s=>p(276)(48),cout=>p(277)(49));
FA_ff_9234:FAff port map(x=>p(220)(49),y=>p(221)(49),Cin=>p(222)(49),clock=>clock,reset=>reset,s=>p(276)(49),cout=>p(277)(50));
FA_ff_9235:FAff port map(x=>p(220)(50),y=>p(221)(50),Cin=>p(222)(50),clock=>clock,reset=>reset,s=>p(276)(50),cout=>p(277)(51));
FA_ff_9236:FAff port map(x=>p(220)(51),y=>p(221)(51),Cin=>p(222)(51),clock=>clock,reset=>reset,s=>p(276)(51),cout=>p(277)(52));
FA_ff_9237:FAff port map(x=>p(220)(52),y=>p(221)(52),Cin=>p(222)(52),clock=>clock,reset=>reset,s=>p(276)(52),cout=>p(277)(53));
FA_ff_9238:FAff port map(x=>p(220)(53),y=>p(221)(53),Cin=>p(222)(53),clock=>clock,reset=>reset,s=>p(276)(53),cout=>p(277)(54));
FA_ff_9239:FAff port map(x=>p(220)(54),y=>p(221)(54),Cin=>p(222)(54),clock=>clock,reset=>reset,s=>p(276)(54),cout=>p(277)(55));
FA_ff_9240:FAff port map(x=>p(220)(55),y=>p(221)(55),Cin=>p(222)(55),clock=>clock,reset=>reset,s=>p(276)(55),cout=>p(277)(56));
FA_ff_9241:FAff port map(x=>p(220)(56),y=>p(221)(56),Cin=>p(222)(56),clock=>clock,reset=>reset,s=>p(276)(56),cout=>p(277)(57));
FA_ff_9242:FAff port map(x=>p(220)(57),y=>p(221)(57),Cin=>p(222)(57),clock=>clock,reset=>reset,s=>p(276)(57),cout=>p(277)(58));
FA_ff_9243:FAff port map(x=>p(220)(58),y=>p(221)(58),Cin=>p(222)(58),clock=>clock,reset=>reset,s=>p(276)(58),cout=>p(277)(59));
FA_ff_9244:FAff port map(x=>p(220)(59),y=>p(221)(59),Cin=>p(222)(59),clock=>clock,reset=>reset,s=>p(276)(59),cout=>p(277)(60));
FA_ff_9245:FAff port map(x=>p(220)(60),y=>p(221)(60),Cin=>p(222)(60),clock=>clock,reset=>reset,s=>p(276)(60),cout=>p(277)(61));
FA_ff_9246:FAff port map(x=>p(220)(61),y=>p(221)(61),Cin=>p(222)(61),clock=>clock,reset=>reset,s=>p(276)(61),cout=>p(277)(62));
FA_ff_9247:FAff port map(x=>p(220)(62),y=>p(221)(62),Cin=>p(222)(62),clock=>clock,reset=>reset,s=>p(276)(62),cout=>p(277)(63));
FA_ff_9248:FAff port map(x=>p(220)(63),y=>p(221)(63),Cin=>p(222)(63),clock=>clock,reset=>reset,s=>p(276)(63),cout=>p(277)(64));
FA_ff_9249:FAff port map(x=>p(220)(64),y=>p(221)(64),Cin=>p(222)(64),clock=>clock,reset=>reset,s=>p(276)(64),cout=>p(277)(65));
FA_ff_9250:FAff port map(x=>p(220)(65),y=>p(221)(65),Cin=>p(222)(65),clock=>clock,reset=>reset,s=>p(276)(65),cout=>p(277)(66));
FA_ff_9251:FAff port map(x=>p(220)(66),y=>p(221)(66),Cin=>p(222)(66),clock=>clock,reset=>reset,s=>p(276)(66),cout=>p(277)(67));
FA_ff_9252:FAff port map(x=>p(220)(67),y=>p(221)(67),Cin=>p(222)(67),clock=>clock,reset=>reset,s=>p(276)(67),cout=>p(277)(68));
FA_ff_9253:FAff port map(x=>p(220)(68),y=>p(221)(68),Cin=>p(222)(68),clock=>clock,reset=>reset,s=>p(276)(68),cout=>p(277)(69));
FA_ff_9254:FAff port map(x=>p(220)(69),y=>p(221)(69),Cin=>p(222)(69),clock=>clock,reset=>reset,s=>p(276)(69),cout=>p(277)(70));
FA_ff_9255:FAff port map(x=>p(220)(70),y=>p(221)(70),Cin=>p(222)(70),clock=>clock,reset=>reset,s=>p(276)(70),cout=>p(277)(71));
FA_ff_9256:FAff port map(x=>p(220)(71),y=>p(221)(71),Cin=>p(222)(71),clock=>clock,reset=>reset,s=>p(276)(71),cout=>p(277)(72));
FA_ff_9257:FAff port map(x=>p(220)(72),y=>p(221)(72),Cin=>p(222)(72),clock=>clock,reset=>reset,s=>p(276)(72),cout=>p(277)(73));
FA_ff_9258:FAff port map(x=>p(220)(73),y=>p(221)(73),Cin=>p(222)(73),clock=>clock,reset=>reset,s=>p(276)(73),cout=>p(277)(74));
FA_ff_9259:FAff port map(x=>p(220)(74),y=>p(221)(74),Cin=>p(222)(74),clock=>clock,reset=>reset,s=>p(276)(74),cout=>p(277)(75));
FA_ff_9260:FAff port map(x=>p(220)(75),y=>p(221)(75),Cin=>p(222)(75),clock=>clock,reset=>reset,s=>p(276)(75),cout=>p(277)(76));
FA_ff_9261:FAff port map(x=>p(220)(76),y=>p(221)(76),Cin=>p(222)(76),clock=>clock,reset=>reset,s=>p(276)(76),cout=>p(277)(77));
FA_ff_9262:FAff port map(x=>p(220)(77),y=>p(221)(77),Cin=>p(222)(77),clock=>clock,reset=>reset,s=>p(276)(77),cout=>p(277)(78));
FA_ff_9263:FAff port map(x=>p(220)(78),y=>p(221)(78),Cin=>p(222)(78),clock=>clock,reset=>reset,s=>p(276)(78),cout=>p(277)(79));
FA_ff_9264:FAff port map(x=>p(220)(79),y=>p(221)(79),Cin=>p(222)(79),clock=>clock,reset=>reset,s=>p(276)(79),cout=>p(277)(80));
FA_ff_9265:FAff port map(x=>p(220)(80),y=>p(221)(80),Cin=>p(222)(80),clock=>clock,reset=>reset,s=>p(276)(80),cout=>p(277)(81));
FA_ff_9266:FAff port map(x=>p(220)(81),y=>p(221)(81),Cin=>p(222)(81),clock=>clock,reset=>reset,s=>p(276)(81),cout=>p(277)(82));
FA_ff_9267:FAff port map(x=>p(220)(82),y=>p(221)(82),Cin=>p(222)(82),clock=>clock,reset=>reset,s=>p(276)(82),cout=>p(277)(83));
FA_ff_9268:FAff port map(x=>p(220)(83),y=>p(221)(83),Cin=>p(222)(83),clock=>clock,reset=>reset,s=>p(276)(83),cout=>p(277)(84));
FA_ff_9269:FAff port map(x=>p(220)(84),y=>p(221)(84),Cin=>p(222)(84),clock=>clock,reset=>reset,s=>p(276)(84),cout=>p(277)(85));
FA_ff_9270:FAff port map(x=>p(220)(85),y=>p(221)(85),Cin=>p(222)(85),clock=>clock,reset=>reset,s=>p(276)(85),cout=>p(277)(86));
FA_ff_9271:FAff port map(x=>p(220)(86),y=>p(221)(86),Cin=>p(222)(86),clock=>clock,reset=>reset,s=>p(276)(86),cout=>p(277)(87));
FA_ff_9272:FAff port map(x=>p(220)(87),y=>p(221)(87),Cin=>p(222)(87),clock=>clock,reset=>reset,s=>p(276)(87),cout=>p(277)(88));
FA_ff_9273:FAff port map(x=>p(220)(88),y=>p(221)(88),Cin=>p(222)(88),clock=>clock,reset=>reset,s=>p(276)(88),cout=>p(277)(89));
FA_ff_9274:FAff port map(x=>p(220)(89),y=>p(221)(89),Cin=>p(222)(89),clock=>clock,reset=>reset,s=>p(276)(89),cout=>p(277)(90));
FA_ff_9275:FAff port map(x=>p(220)(90),y=>p(221)(90),Cin=>p(222)(90),clock=>clock,reset=>reset,s=>p(276)(90),cout=>p(277)(91));
FA_ff_9276:FAff port map(x=>p(220)(91),y=>p(221)(91),Cin=>p(222)(91),clock=>clock,reset=>reset,s=>p(276)(91),cout=>p(277)(92));
FA_ff_9277:FAff port map(x=>p(220)(92),y=>p(221)(92),Cin=>p(222)(92),clock=>clock,reset=>reset,s=>p(276)(92),cout=>p(277)(93));
FA_ff_9278:FAff port map(x=>p(220)(93),y=>p(221)(93),Cin=>p(222)(93),clock=>clock,reset=>reset,s=>p(276)(93),cout=>p(277)(94));
FA_ff_9279:FAff port map(x=>p(220)(94),y=>p(221)(94),Cin=>p(222)(94),clock=>clock,reset=>reset,s=>p(276)(94),cout=>p(277)(95));
FA_ff_9280:FAff port map(x=>p(220)(95),y=>p(221)(95),Cin=>p(222)(95),clock=>clock,reset=>reset,s=>p(276)(95),cout=>p(277)(96));
FA_ff_9281:FAff port map(x=>p(220)(96),y=>p(221)(96),Cin=>p(222)(96),clock=>clock,reset=>reset,s=>p(276)(96),cout=>p(277)(97));
FA_ff_9282:FAff port map(x=>p(220)(97),y=>p(221)(97),Cin=>p(222)(97),clock=>clock,reset=>reset,s=>p(276)(97),cout=>p(277)(98));
FA_ff_9283:FAff port map(x=>p(220)(98),y=>p(221)(98),Cin=>p(222)(98),clock=>clock,reset=>reset,s=>p(276)(98),cout=>p(277)(99));
FA_ff_9284:FAff port map(x=>p(220)(99),y=>p(221)(99),Cin=>p(222)(99),clock=>clock,reset=>reset,s=>p(276)(99),cout=>p(277)(100));
FA_ff_9285:FAff port map(x=>p(220)(100),y=>p(221)(100),Cin=>p(222)(100),clock=>clock,reset=>reset,s=>p(276)(100),cout=>p(277)(101));
FA_ff_9286:FAff port map(x=>p(220)(101),y=>p(221)(101),Cin=>p(222)(101),clock=>clock,reset=>reset,s=>p(276)(101),cout=>p(277)(102));
FA_ff_9287:FAff port map(x=>p(220)(102),y=>p(221)(102),Cin=>p(222)(102),clock=>clock,reset=>reset,s=>p(276)(102),cout=>p(277)(103));
FA_ff_9288:FAff port map(x=>p(220)(103),y=>p(221)(103),Cin=>p(222)(103),clock=>clock,reset=>reset,s=>p(276)(103),cout=>p(277)(104));
FA_ff_9289:FAff port map(x=>p(220)(104),y=>p(221)(104),Cin=>p(222)(104),clock=>clock,reset=>reset,s=>p(276)(104),cout=>p(277)(105));
FA_ff_9290:FAff port map(x=>p(220)(105),y=>p(221)(105),Cin=>p(222)(105),clock=>clock,reset=>reset,s=>p(276)(105),cout=>p(277)(106));
FA_ff_9291:FAff port map(x=>p(220)(106),y=>p(221)(106),Cin=>p(222)(106),clock=>clock,reset=>reset,s=>p(276)(106),cout=>p(277)(107));
FA_ff_9292:FAff port map(x=>p(220)(107),y=>p(221)(107),Cin=>p(222)(107),clock=>clock,reset=>reset,s=>p(276)(107),cout=>p(277)(108));
FA_ff_9293:FAff port map(x=>p(220)(108),y=>p(221)(108),Cin=>p(222)(108),clock=>clock,reset=>reset,s=>p(276)(108),cout=>p(277)(109));
FA_ff_9294:FAff port map(x=>p(220)(109),y=>p(221)(109),Cin=>p(222)(109),clock=>clock,reset=>reset,s=>p(276)(109),cout=>p(277)(110));
FA_ff_9295:FAff port map(x=>p(220)(110),y=>p(221)(110),Cin=>p(222)(110),clock=>clock,reset=>reset,s=>p(276)(110),cout=>p(277)(111));
FA_ff_9296:FAff port map(x=>p(220)(111),y=>p(221)(111),Cin=>p(222)(111),clock=>clock,reset=>reset,s=>p(276)(111),cout=>p(277)(112));
FA_ff_9297:FAff port map(x=>p(220)(112),y=>p(221)(112),Cin=>p(222)(112),clock=>clock,reset=>reset,s=>p(276)(112),cout=>p(277)(113));
FA_ff_9298:FAff port map(x=>p(220)(113),y=>p(221)(113),Cin=>p(222)(113),clock=>clock,reset=>reset,s=>p(276)(113),cout=>p(277)(114));
FA_ff_9299:FAff port map(x=>p(220)(114),y=>p(221)(114),Cin=>p(222)(114),clock=>clock,reset=>reset,s=>p(276)(114),cout=>p(277)(115));
FA_ff_9300:FAff port map(x=>p(220)(115),y=>p(221)(115),Cin=>p(222)(115),clock=>clock,reset=>reset,s=>p(276)(115),cout=>p(277)(116));
FA_ff_9301:FAff port map(x=>p(220)(116),y=>p(221)(116),Cin=>p(222)(116),clock=>clock,reset=>reset,s=>p(276)(116),cout=>p(277)(117));
FA_ff_9302:FAff port map(x=>p(220)(117),y=>p(221)(117),Cin=>p(222)(117),clock=>clock,reset=>reset,s=>p(276)(117),cout=>p(277)(118));
FA_ff_9303:FAff port map(x=>p(220)(118),y=>p(221)(118),Cin=>p(222)(118),clock=>clock,reset=>reset,s=>p(276)(118),cout=>p(277)(119));
FA_ff_9304:FAff port map(x=>p(220)(119),y=>p(221)(119),Cin=>p(222)(119),clock=>clock,reset=>reset,s=>p(276)(119),cout=>p(277)(120));
FA_ff_9305:FAff port map(x=>p(220)(120),y=>p(221)(120),Cin=>p(222)(120),clock=>clock,reset=>reset,s=>p(276)(120),cout=>p(277)(121));
FA_ff_9306:FAff port map(x=>p(220)(121),y=>p(221)(121),Cin=>p(222)(121),clock=>clock,reset=>reset,s=>p(276)(121),cout=>p(277)(122));
FA_ff_9307:FAff port map(x=>p(220)(122),y=>p(221)(122),Cin=>p(222)(122),clock=>clock,reset=>reset,s=>p(276)(122),cout=>p(277)(123));
FA_ff_9308:FAff port map(x=>p(220)(123),y=>p(221)(123),Cin=>p(222)(123),clock=>clock,reset=>reset,s=>p(276)(123),cout=>p(277)(124));
FA_ff_9309:FAff port map(x=>p(220)(124),y=>p(221)(124),Cin=>p(222)(124),clock=>clock,reset=>reset,s=>p(276)(124),cout=>p(277)(125));
FA_ff_9310:FAff port map(x=>p(220)(125),y=>p(221)(125),Cin=>p(222)(125),clock=>clock,reset=>reset,s=>p(276)(125),cout=>p(277)(126));
FA_ff_9311:FAff port map(x=>p(220)(126),y=>p(221)(126),Cin=>p(222)(126),clock=>clock,reset=>reset,s=>p(276)(126),cout=>p(277)(127));
FA_ff_9312:FAff port map(x=>p(220)(127),y=>p(221)(127),Cin=>p(222)(127),clock=>clock,reset=>reset,s=>p(276)(127),cout=>p(277)(128));
FA_ff_9313:FAff port map(x=>p(220)(128),y=>p(221)(128),Cin=>p(222)(128),clock=>clock,reset=>reset,s=>p(276)(128),cout=>p(277)(129));
p(276)(129)<=p(221)(129);
p(278)(0)<=p(224)(0);
HA_ff_32:HAff port map(x=>p(223)(1),y=>p(224)(1),clock=>clock,reset=>reset,s=>p(278)(1),c=>p(279)(2));
FA_ff_9314:FAff port map(x=>p(223)(2),y=>p(224)(2),Cin=>p(225)(2),clock=>clock,reset=>reset,s=>p(278)(2),cout=>p(279)(3));
FA_ff_9315:FAff port map(x=>p(223)(3),y=>p(224)(3),Cin=>p(225)(3),clock=>clock,reset=>reset,s=>p(278)(3),cout=>p(279)(4));
FA_ff_9316:FAff port map(x=>p(223)(4),y=>p(224)(4),Cin=>p(225)(4),clock=>clock,reset=>reset,s=>p(278)(4),cout=>p(279)(5));
FA_ff_9317:FAff port map(x=>p(223)(5),y=>p(224)(5),Cin=>p(225)(5),clock=>clock,reset=>reset,s=>p(278)(5),cout=>p(279)(6));
FA_ff_9318:FAff port map(x=>p(223)(6),y=>p(224)(6),Cin=>p(225)(6),clock=>clock,reset=>reset,s=>p(278)(6),cout=>p(279)(7));
FA_ff_9319:FAff port map(x=>p(223)(7),y=>p(224)(7),Cin=>p(225)(7),clock=>clock,reset=>reset,s=>p(278)(7),cout=>p(279)(8));
FA_ff_9320:FAff port map(x=>p(223)(8),y=>p(224)(8),Cin=>p(225)(8),clock=>clock,reset=>reset,s=>p(278)(8),cout=>p(279)(9));
FA_ff_9321:FAff port map(x=>p(223)(9),y=>p(224)(9),Cin=>p(225)(9),clock=>clock,reset=>reset,s=>p(278)(9),cout=>p(279)(10));
FA_ff_9322:FAff port map(x=>p(223)(10),y=>p(224)(10),Cin=>p(225)(10),clock=>clock,reset=>reset,s=>p(278)(10),cout=>p(279)(11));
FA_ff_9323:FAff port map(x=>p(223)(11),y=>p(224)(11),Cin=>p(225)(11),clock=>clock,reset=>reset,s=>p(278)(11),cout=>p(279)(12));
FA_ff_9324:FAff port map(x=>p(223)(12),y=>p(224)(12),Cin=>p(225)(12),clock=>clock,reset=>reset,s=>p(278)(12),cout=>p(279)(13));
FA_ff_9325:FAff port map(x=>p(223)(13),y=>p(224)(13),Cin=>p(225)(13),clock=>clock,reset=>reset,s=>p(278)(13),cout=>p(279)(14));
FA_ff_9326:FAff port map(x=>p(223)(14),y=>p(224)(14),Cin=>p(225)(14),clock=>clock,reset=>reset,s=>p(278)(14),cout=>p(279)(15));
FA_ff_9327:FAff port map(x=>p(223)(15),y=>p(224)(15),Cin=>p(225)(15),clock=>clock,reset=>reset,s=>p(278)(15),cout=>p(279)(16));
FA_ff_9328:FAff port map(x=>p(223)(16),y=>p(224)(16),Cin=>p(225)(16),clock=>clock,reset=>reset,s=>p(278)(16),cout=>p(279)(17));
FA_ff_9329:FAff port map(x=>p(223)(17),y=>p(224)(17),Cin=>p(225)(17),clock=>clock,reset=>reset,s=>p(278)(17),cout=>p(279)(18));
FA_ff_9330:FAff port map(x=>p(223)(18),y=>p(224)(18),Cin=>p(225)(18),clock=>clock,reset=>reset,s=>p(278)(18),cout=>p(279)(19));
FA_ff_9331:FAff port map(x=>p(223)(19),y=>p(224)(19),Cin=>p(225)(19),clock=>clock,reset=>reset,s=>p(278)(19),cout=>p(279)(20));
FA_ff_9332:FAff port map(x=>p(223)(20),y=>p(224)(20),Cin=>p(225)(20),clock=>clock,reset=>reset,s=>p(278)(20),cout=>p(279)(21));
FA_ff_9333:FAff port map(x=>p(223)(21),y=>p(224)(21),Cin=>p(225)(21),clock=>clock,reset=>reset,s=>p(278)(21),cout=>p(279)(22));
FA_ff_9334:FAff port map(x=>p(223)(22),y=>p(224)(22),Cin=>p(225)(22),clock=>clock,reset=>reset,s=>p(278)(22),cout=>p(279)(23));
FA_ff_9335:FAff port map(x=>p(223)(23),y=>p(224)(23),Cin=>p(225)(23),clock=>clock,reset=>reset,s=>p(278)(23),cout=>p(279)(24));
FA_ff_9336:FAff port map(x=>p(223)(24),y=>p(224)(24),Cin=>p(225)(24),clock=>clock,reset=>reset,s=>p(278)(24),cout=>p(279)(25));
FA_ff_9337:FAff port map(x=>p(223)(25),y=>p(224)(25),Cin=>p(225)(25),clock=>clock,reset=>reset,s=>p(278)(25),cout=>p(279)(26));
FA_ff_9338:FAff port map(x=>p(223)(26),y=>p(224)(26),Cin=>p(225)(26),clock=>clock,reset=>reset,s=>p(278)(26),cout=>p(279)(27));
FA_ff_9339:FAff port map(x=>p(223)(27),y=>p(224)(27),Cin=>p(225)(27),clock=>clock,reset=>reset,s=>p(278)(27),cout=>p(279)(28));
FA_ff_9340:FAff port map(x=>p(223)(28),y=>p(224)(28),Cin=>p(225)(28),clock=>clock,reset=>reset,s=>p(278)(28),cout=>p(279)(29));
FA_ff_9341:FAff port map(x=>p(223)(29),y=>p(224)(29),Cin=>p(225)(29),clock=>clock,reset=>reset,s=>p(278)(29),cout=>p(279)(30));
FA_ff_9342:FAff port map(x=>p(223)(30),y=>p(224)(30),Cin=>p(225)(30),clock=>clock,reset=>reset,s=>p(278)(30),cout=>p(279)(31));
FA_ff_9343:FAff port map(x=>p(223)(31),y=>p(224)(31),Cin=>p(225)(31),clock=>clock,reset=>reset,s=>p(278)(31),cout=>p(279)(32));
FA_ff_9344:FAff port map(x=>p(223)(32),y=>p(224)(32),Cin=>p(225)(32),clock=>clock,reset=>reset,s=>p(278)(32),cout=>p(279)(33));
FA_ff_9345:FAff port map(x=>p(223)(33),y=>p(224)(33),Cin=>p(225)(33),clock=>clock,reset=>reset,s=>p(278)(33),cout=>p(279)(34));
FA_ff_9346:FAff port map(x=>p(223)(34),y=>p(224)(34),Cin=>p(225)(34),clock=>clock,reset=>reset,s=>p(278)(34),cout=>p(279)(35));
FA_ff_9347:FAff port map(x=>p(223)(35),y=>p(224)(35),Cin=>p(225)(35),clock=>clock,reset=>reset,s=>p(278)(35),cout=>p(279)(36));
FA_ff_9348:FAff port map(x=>p(223)(36),y=>p(224)(36),Cin=>p(225)(36),clock=>clock,reset=>reset,s=>p(278)(36),cout=>p(279)(37));
FA_ff_9349:FAff port map(x=>p(223)(37),y=>p(224)(37),Cin=>p(225)(37),clock=>clock,reset=>reset,s=>p(278)(37),cout=>p(279)(38));
FA_ff_9350:FAff port map(x=>p(223)(38),y=>p(224)(38),Cin=>p(225)(38),clock=>clock,reset=>reset,s=>p(278)(38),cout=>p(279)(39));
FA_ff_9351:FAff port map(x=>p(223)(39),y=>p(224)(39),Cin=>p(225)(39),clock=>clock,reset=>reset,s=>p(278)(39),cout=>p(279)(40));
FA_ff_9352:FAff port map(x=>p(223)(40),y=>p(224)(40),Cin=>p(225)(40),clock=>clock,reset=>reset,s=>p(278)(40),cout=>p(279)(41));
FA_ff_9353:FAff port map(x=>p(223)(41),y=>p(224)(41),Cin=>p(225)(41),clock=>clock,reset=>reset,s=>p(278)(41),cout=>p(279)(42));
FA_ff_9354:FAff port map(x=>p(223)(42),y=>p(224)(42),Cin=>p(225)(42),clock=>clock,reset=>reset,s=>p(278)(42),cout=>p(279)(43));
FA_ff_9355:FAff port map(x=>p(223)(43),y=>p(224)(43),Cin=>p(225)(43),clock=>clock,reset=>reset,s=>p(278)(43),cout=>p(279)(44));
FA_ff_9356:FAff port map(x=>p(223)(44),y=>p(224)(44),Cin=>p(225)(44),clock=>clock,reset=>reset,s=>p(278)(44),cout=>p(279)(45));
FA_ff_9357:FAff port map(x=>p(223)(45),y=>p(224)(45),Cin=>p(225)(45),clock=>clock,reset=>reset,s=>p(278)(45),cout=>p(279)(46));
FA_ff_9358:FAff port map(x=>p(223)(46),y=>p(224)(46),Cin=>p(225)(46),clock=>clock,reset=>reset,s=>p(278)(46),cout=>p(279)(47));
FA_ff_9359:FAff port map(x=>p(223)(47),y=>p(224)(47),Cin=>p(225)(47),clock=>clock,reset=>reset,s=>p(278)(47),cout=>p(279)(48));
FA_ff_9360:FAff port map(x=>p(223)(48),y=>p(224)(48),Cin=>p(225)(48),clock=>clock,reset=>reset,s=>p(278)(48),cout=>p(279)(49));
FA_ff_9361:FAff port map(x=>p(223)(49),y=>p(224)(49),Cin=>p(225)(49),clock=>clock,reset=>reset,s=>p(278)(49),cout=>p(279)(50));
FA_ff_9362:FAff port map(x=>p(223)(50),y=>p(224)(50),Cin=>p(225)(50),clock=>clock,reset=>reset,s=>p(278)(50),cout=>p(279)(51));
FA_ff_9363:FAff port map(x=>p(223)(51),y=>p(224)(51),Cin=>p(225)(51),clock=>clock,reset=>reset,s=>p(278)(51),cout=>p(279)(52));
FA_ff_9364:FAff port map(x=>p(223)(52),y=>p(224)(52),Cin=>p(225)(52),clock=>clock,reset=>reset,s=>p(278)(52),cout=>p(279)(53));
FA_ff_9365:FAff port map(x=>p(223)(53),y=>p(224)(53),Cin=>p(225)(53),clock=>clock,reset=>reset,s=>p(278)(53),cout=>p(279)(54));
FA_ff_9366:FAff port map(x=>p(223)(54),y=>p(224)(54),Cin=>p(225)(54),clock=>clock,reset=>reset,s=>p(278)(54),cout=>p(279)(55));
FA_ff_9367:FAff port map(x=>p(223)(55),y=>p(224)(55),Cin=>p(225)(55),clock=>clock,reset=>reset,s=>p(278)(55),cout=>p(279)(56));
FA_ff_9368:FAff port map(x=>p(223)(56),y=>p(224)(56),Cin=>p(225)(56),clock=>clock,reset=>reset,s=>p(278)(56),cout=>p(279)(57));
FA_ff_9369:FAff port map(x=>p(223)(57),y=>p(224)(57),Cin=>p(225)(57),clock=>clock,reset=>reset,s=>p(278)(57),cout=>p(279)(58));
FA_ff_9370:FAff port map(x=>p(223)(58),y=>p(224)(58),Cin=>p(225)(58),clock=>clock,reset=>reset,s=>p(278)(58),cout=>p(279)(59));
FA_ff_9371:FAff port map(x=>p(223)(59),y=>p(224)(59),Cin=>p(225)(59),clock=>clock,reset=>reset,s=>p(278)(59),cout=>p(279)(60));
FA_ff_9372:FAff port map(x=>p(223)(60),y=>p(224)(60),Cin=>p(225)(60),clock=>clock,reset=>reset,s=>p(278)(60),cout=>p(279)(61));
FA_ff_9373:FAff port map(x=>p(223)(61),y=>p(224)(61),Cin=>p(225)(61),clock=>clock,reset=>reset,s=>p(278)(61),cout=>p(279)(62));
FA_ff_9374:FAff port map(x=>p(223)(62),y=>p(224)(62),Cin=>p(225)(62),clock=>clock,reset=>reset,s=>p(278)(62),cout=>p(279)(63));
FA_ff_9375:FAff port map(x=>p(223)(63),y=>p(224)(63),Cin=>p(225)(63),clock=>clock,reset=>reset,s=>p(278)(63),cout=>p(279)(64));
FA_ff_9376:FAff port map(x=>p(223)(64),y=>p(224)(64),Cin=>p(225)(64),clock=>clock,reset=>reset,s=>p(278)(64),cout=>p(279)(65));
FA_ff_9377:FAff port map(x=>p(223)(65),y=>p(224)(65),Cin=>p(225)(65),clock=>clock,reset=>reset,s=>p(278)(65),cout=>p(279)(66));
FA_ff_9378:FAff port map(x=>p(223)(66),y=>p(224)(66),Cin=>p(225)(66),clock=>clock,reset=>reset,s=>p(278)(66),cout=>p(279)(67));
FA_ff_9379:FAff port map(x=>p(223)(67),y=>p(224)(67),Cin=>p(225)(67),clock=>clock,reset=>reset,s=>p(278)(67),cout=>p(279)(68));
FA_ff_9380:FAff port map(x=>p(223)(68),y=>p(224)(68),Cin=>p(225)(68),clock=>clock,reset=>reset,s=>p(278)(68),cout=>p(279)(69));
FA_ff_9381:FAff port map(x=>p(223)(69),y=>p(224)(69),Cin=>p(225)(69),clock=>clock,reset=>reset,s=>p(278)(69),cout=>p(279)(70));
FA_ff_9382:FAff port map(x=>p(223)(70),y=>p(224)(70),Cin=>p(225)(70),clock=>clock,reset=>reset,s=>p(278)(70),cout=>p(279)(71));
FA_ff_9383:FAff port map(x=>p(223)(71),y=>p(224)(71),Cin=>p(225)(71),clock=>clock,reset=>reset,s=>p(278)(71),cout=>p(279)(72));
FA_ff_9384:FAff port map(x=>p(223)(72),y=>p(224)(72),Cin=>p(225)(72),clock=>clock,reset=>reset,s=>p(278)(72),cout=>p(279)(73));
FA_ff_9385:FAff port map(x=>p(223)(73),y=>p(224)(73),Cin=>p(225)(73),clock=>clock,reset=>reset,s=>p(278)(73),cout=>p(279)(74));
FA_ff_9386:FAff port map(x=>p(223)(74),y=>p(224)(74),Cin=>p(225)(74),clock=>clock,reset=>reset,s=>p(278)(74),cout=>p(279)(75));
FA_ff_9387:FAff port map(x=>p(223)(75),y=>p(224)(75),Cin=>p(225)(75),clock=>clock,reset=>reset,s=>p(278)(75),cout=>p(279)(76));
FA_ff_9388:FAff port map(x=>p(223)(76),y=>p(224)(76),Cin=>p(225)(76),clock=>clock,reset=>reset,s=>p(278)(76),cout=>p(279)(77));
FA_ff_9389:FAff port map(x=>p(223)(77),y=>p(224)(77),Cin=>p(225)(77),clock=>clock,reset=>reset,s=>p(278)(77),cout=>p(279)(78));
FA_ff_9390:FAff port map(x=>p(223)(78),y=>p(224)(78),Cin=>p(225)(78),clock=>clock,reset=>reset,s=>p(278)(78),cout=>p(279)(79));
FA_ff_9391:FAff port map(x=>p(223)(79),y=>p(224)(79),Cin=>p(225)(79),clock=>clock,reset=>reset,s=>p(278)(79),cout=>p(279)(80));
FA_ff_9392:FAff port map(x=>p(223)(80),y=>p(224)(80),Cin=>p(225)(80),clock=>clock,reset=>reset,s=>p(278)(80),cout=>p(279)(81));
FA_ff_9393:FAff port map(x=>p(223)(81),y=>p(224)(81),Cin=>p(225)(81),clock=>clock,reset=>reset,s=>p(278)(81),cout=>p(279)(82));
FA_ff_9394:FAff port map(x=>p(223)(82),y=>p(224)(82),Cin=>p(225)(82),clock=>clock,reset=>reset,s=>p(278)(82),cout=>p(279)(83));
FA_ff_9395:FAff port map(x=>p(223)(83),y=>p(224)(83),Cin=>p(225)(83),clock=>clock,reset=>reset,s=>p(278)(83),cout=>p(279)(84));
FA_ff_9396:FAff port map(x=>p(223)(84),y=>p(224)(84),Cin=>p(225)(84),clock=>clock,reset=>reset,s=>p(278)(84),cout=>p(279)(85));
FA_ff_9397:FAff port map(x=>p(223)(85),y=>p(224)(85),Cin=>p(225)(85),clock=>clock,reset=>reset,s=>p(278)(85),cout=>p(279)(86));
FA_ff_9398:FAff port map(x=>p(223)(86),y=>p(224)(86),Cin=>p(225)(86),clock=>clock,reset=>reset,s=>p(278)(86),cout=>p(279)(87));
FA_ff_9399:FAff port map(x=>p(223)(87),y=>p(224)(87),Cin=>p(225)(87),clock=>clock,reset=>reset,s=>p(278)(87),cout=>p(279)(88));
FA_ff_9400:FAff port map(x=>p(223)(88),y=>p(224)(88),Cin=>p(225)(88),clock=>clock,reset=>reset,s=>p(278)(88),cout=>p(279)(89));
FA_ff_9401:FAff port map(x=>p(223)(89),y=>p(224)(89),Cin=>p(225)(89),clock=>clock,reset=>reset,s=>p(278)(89),cout=>p(279)(90));
FA_ff_9402:FAff port map(x=>p(223)(90),y=>p(224)(90),Cin=>p(225)(90),clock=>clock,reset=>reset,s=>p(278)(90),cout=>p(279)(91));
FA_ff_9403:FAff port map(x=>p(223)(91),y=>p(224)(91),Cin=>p(225)(91),clock=>clock,reset=>reset,s=>p(278)(91),cout=>p(279)(92));
FA_ff_9404:FAff port map(x=>p(223)(92),y=>p(224)(92),Cin=>p(225)(92),clock=>clock,reset=>reset,s=>p(278)(92),cout=>p(279)(93));
FA_ff_9405:FAff port map(x=>p(223)(93),y=>p(224)(93),Cin=>p(225)(93),clock=>clock,reset=>reset,s=>p(278)(93),cout=>p(279)(94));
FA_ff_9406:FAff port map(x=>p(223)(94),y=>p(224)(94),Cin=>p(225)(94),clock=>clock,reset=>reset,s=>p(278)(94),cout=>p(279)(95));
FA_ff_9407:FAff port map(x=>p(223)(95),y=>p(224)(95),Cin=>p(225)(95),clock=>clock,reset=>reset,s=>p(278)(95),cout=>p(279)(96));
FA_ff_9408:FAff port map(x=>p(223)(96),y=>p(224)(96),Cin=>p(225)(96),clock=>clock,reset=>reset,s=>p(278)(96),cout=>p(279)(97));
FA_ff_9409:FAff port map(x=>p(223)(97),y=>p(224)(97),Cin=>p(225)(97),clock=>clock,reset=>reset,s=>p(278)(97),cout=>p(279)(98));
FA_ff_9410:FAff port map(x=>p(223)(98),y=>p(224)(98),Cin=>p(225)(98),clock=>clock,reset=>reset,s=>p(278)(98),cout=>p(279)(99));
FA_ff_9411:FAff port map(x=>p(223)(99),y=>p(224)(99),Cin=>p(225)(99),clock=>clock,reset=>reset,s=>p(278)(99),cout=>p(279)(100));
FA_ff_9412:FAff port map(x=>p(223)(100),y=>p(224)(100),Cin=>p(225)(100),clock=>clock,reset=>reset,s=>p(278)(100),cout=>p(279)(101));
FA_ff_9413:FAff port map(x=>p(223)(101),y=>p(224)(101),Cin=>p(225)(101),clock=>clock,reset=>reset,s=>p(278)(101),cout=>p(279)(102));
FA_ff_9414:FAff port map(x=>p(223)(102),y=>p(224)(102),Cin=>p(225)(102),clock=>clock,reset=>reset,s=>p(278)(102),cout=>p(279)(103));
FA_ff_9415:FAff port map(x=>p(223)(103),y=>p(224)(103),Cin=>p(225)(103),clock=>clock,reset=>reset,s=>p(278)(103),cout=>p(279)(104));
FA_ff_9416:FAff port map(x=>p(223)(104),y=>p(224)(104),Cin=>p(225)(104),clock=>clock,reset=>reset,s=>p(278)(104),cout=>p(279)(105));
FA_ff_9417:FAff port map(x=>p(223)(105),y=>p(224)(105),Cin=>p(225)(105),clock=>clock,reset=>reset,s=>p(278)(105),cout=>p(279)(106));
FA_ff_9418:FAff port map(x=>p(223)(106),y=>p(224)(106),Cin=>p(225)(106),clock=>clock,reset=>reset,s=>p(278)(106),cout=>p(279)(107));
FA_ff_9419:FAff port map(x=>p(223)(107),y=>p(224)(107),Cin=>p(225)(107),clock=>clock,reset=>reset,s=>p(278)(107),cout=>p(279)(108));
FA_ff_9420:FAff port map(x=>p(223)(108),y=>p(224)(108),Cin=>p(225)(108),clock=>clock,reset=>reset,s=>p(278)(108),cout=>p(279)(109));
FA_ff_9421:FAff port map(x=>p(223)(109),y=>p(224)(109),Cin=>p(225)(109),clock=>clock,reset=>reset,s=>p(278)(109),cout=>p(279)(110));
FA_ff_9422:FAff port map(x=>p(223)(110),y=>p(224)(110),Cin=>p(225)(110),clock=>clock,reset=>reset,s=>p(278)(110),cout=>p(279)(111));
FA_ff_9423:FAff port map(x=>p(223)(111),y=>p(224)(111),Cin=>p(225)(111),clock=>clock,reset=>reset,s=>p(278)(111),cout=>p(279)(112));
FA_ff_9424:FAff port map(x=>p(223)(112),y=>p(224)(112),Cin=>p(225)(112),clock=>clock,reset=>reset,s=>p(278)(112),cout=>p(279)(113));
FA_ff_9425:FAff port map(x=>p(223)(113),y=>p(224)(113),Cin=>p(225)(113),clock=>clock,reset=>reset,s=>p(278)(113),cout=>p(279)(114));
FA_ff_9426:FAff port map(x=>p(223)(114),y=>p(224)(114),Cin=>p(225)(114),clock=>clock,reset=>reset,s=>p(278)(114),cout=>p(279)(115));
FA_ff_9427:FAff port map(x=>p(223)(115),y=>p(224)(115),Cin=>p(225)(115),clock=>clock,reset=>reset,s=>p(278)(115),cout=>p(279)(116));
FA_ff_9428:FAff port map(x=>p(223)(116),y=>p(224)(116),Cin=>p(225)(116),clock=>clock,reset=>reset,s=>p(278)(116),cout=>p(279)(117));
FA_ff_9429:FAff port map(x=>p(223)(117),y=>p(224)(117),Cin=>p(225)(117),clock=>clock,reset=>reset,s=>p(278)(117),cout=>p(279)(118));
FA_ff_9430:FAff port map(x=>p(223)(118),y=>p(224)(118),Cin=>p(225)(118),clock=>clock,reset=>reset,s=>p(278)(118),cout=>p(279)(119));
FA_ff_9431:FAff port map(x=>p(223)(119),y=>p(224)(119),Cin=>p(225)(119),clock=>clock,reset=>reset,s=>p(278)(119),cout=>p(279)(120));
FA_ff_9432:FAff port map(x=>p(223)(120),y=>p(224)(120),Cin=>p(225)(120),clock=>clock,reset=>reset,s=>p(278)(120),cout=>p(279)(121));
FA_ff_9433:FAff port map(x=>p(223)(121),y=>p(224)(121),Cin=>p(225)(121),clock=>clock,reset=>reset,s=>p(278)(121),cout=>p(279)(122));
FA_ff_9434:FAff port map(x=>p(223)(122),y=>p(224)(122),Cin=>p(225)(122),clock=>clock,reset=>reset,s=>p(278)(122),cout=>p(279)(123));
FA_ff_9435:FAff port map(x=>p(223)(123),y=>p(224)(123),Cin=>p(225)(123),clock=>clock,reset=>reset,s=>p(278)(123),cout=>p(279)(124));
FA_ff_9436:FAff port map(x=>p(223)(124),y=>p(224)(124),Cin=>p(225)(124),clock=>clock,reset=>reset,s=>p(278)(124),cout=>p(279)(125));
FA_ff_9437:FAff port map(x=>p(223)(125),y=>p(224)(125),Cin=>p(225)(125),clock=>clock,reset=>reset,s=>p(278)(125),cout=>p(279)(126));
FA_ff_9438:FAff port map(x=>p(223)(126),y=>p(224)(126),Cin=>p(225)(126),clock=>clock,reset=>reset,s=>p(278)(126),cout=>p(279)(127));
FA_ff_9439:FAff port map(x=>p(223)(127),y=>p(224)(127),Cin=>p(225)(127),clock=>clock,reset=>reset,s=>p(278)(127),cout=>p(279)(128));
FA_ff_9440:FAff port map(x=>p(223)(128),y=>p(224)(128),Cin=>p(225)(128),clock=>clock,reset=>reset,s=>p(278)(128),cout=>p(279)(129));
p(278)(129)<=p(225)(129);
HA_ff_33:HAff port map(x=>p(226)(0),y=>p(228)(0),clock=>clock,reset=>reset,s=>p(280)(0),c=>p(281)(1));
FA_ff_9441:FAff port map(x=>p(226)(1),y=>p(227)(1),Cin=>p(228)(1),clock=>clock,reset=>reset,s=>p(280)(1),cout=>p(281)(2));
FA_ff_9442:FAff port map(x=>p(226)(2),y=>p(227)(2),Cin=>p(228)(2),clock=>clock,reset=>reset,s=>p(280)(2),cout=>p(281)(3));
FA_ff_9443:FAff port map(x=>p(226)(3),y=>p(227)(3),Cin=>p(228)(3),clock=>clock,reset=>reset,s=>p(280)(3),cout=>p(281)(4));
FA_ff_9444:FAff port map(x=>p(226)(4),y=>p(227)(4),Cin=>p(228)(4),clock=>clock,reset=>reset,s=>p(280)(4),cout=>p(281)(5));
FA_ff_9445:FAff port map(x=>p(226)(5),y=>p(227)(5),Cin=>p(228)(5),clock=>clock,reset=>reset,s=>p(280)(5),cout=>p(281)(6));
FA_ff_9446:FAff port map(x=>p(226)(6),y=>p(227)(6),Cin=>p(228)(6),clock=>clock,reset=>reset,s=>p(280)(6),cout=>p(281)(7));
FA_ff_9447:FAff port map(x=>p(226)(7),y=>p(227)(7),Cin=>p(228)(7),clock=>clock,reset=>reset,s=>p(280)(7),cout=>p(281)(8));
FA_ff_9448:FAff port map(x=>p(226)(8),y=>p(227)(8),Cin=>p(228)(8),clock=>clock,reset=>reset,s=>p(280)(8),cout=>p(281)(9));
FA_ff_9449:FAff port map(x=>p(226)(9),y=>p(227)(9),Cin=>p(228)(9),clock=>clock,reset=>reset,s=>p(280)(9),cout=>p(281)(10));
FA_ff_9450:FAff port map(x=>p(226)(10),y=>p(227)(10),Cin=>p(228)(10),clock=>clock,reset=>reset,s=>p(280)(10),cout=>p(281)(11));
FA_ff_9451:FAff port map(x=>p(226)(11),y=>p(227)(11),Cin=>p(228)(11),clock=>clock,reset=>reset,s=>p(280)(11),cout=>p(281)(12));
FA_ff_9452:FAff port map(x=>p(226)(12),y=>p(227)(12),Cin=>p(228)(12),clock=>clock,reset=>reset,s=>p(280)(12),cout=>p(281)(13));
FA_ff_9453:FAff port map(x=>p(226)(13),y=>p(227)(13),Cin=>p(228)(13),clock=>clock,reset=>reset,s=>p(280)(13),cout=>p(281)(14));
FA_ff_9454:FAff port map(x=>p(226)(14),y=>p(227)(14),Cin=>p(228)(14),clock=>clock,reset=>reset,s=>p(280)(14),cout=>p(281)(15));
FA_ff_9455:FAff port map(x=>p(226)(15),y=>p(227)(15),Cin=>p(228)(15),clock=>clock,reset=>reset,s=>p(280)(15),cout=>p(281)(16));
FA_ff_9456:FAff port map(x=>p(226)(16),y=>p(227)(16),Cin=>p(228)(16),clock=>clock,reset=>reset,s=>p(280)(16),cout=>p(281)(17));
FA_ff_9457:FAff port map(x=>p(226)(17),y=>p(227)(17),Cin=>p(228)(17),clock=>clock,reset=>reset,s=>p(280)(17),cout=>p(281)(18));
FA_ff_9458:FAff port map(x=>p(226)(18),y=>p(227)(18),Cin=>p(228)(18),clock=>clock,reset=>reset,s=>p(280)(18),cout=>p(281)(19));
FA_ff_9459:FAff port map(x=>p(226)(19),y=>p(227)(19),Cin=>p(228)(19),clock=>clock,reset=>reset,s=>p(280)(19),cout=>p(281)(20));
FA_ff_9460:FAff port map(x=>p(226)(20),y=>p(227)(20),Cin=>p(228)(20),clock=>clock,reset=>reset,s=>p(280)(20),cout=>p(281)(21));
FA_ff_9461:FAff port map(x=>p(226)(21),y=>p(227)(21),Cin=>p(228)(21),clock=>clock,reset=>reset,s=>p(280)(21),cout=>p(281)(22));
FA_ff_9462:FAff port map(x=>p(226)(22),y=>p(227)(22),Cin=>p(228)(22),clock=>clock,reset=>reset,s=>p(280)(22),cout=>p(281)(23));
FA_ff_9463:FAff port map(x=>p(226)(23),y=>p(227)(23),Cin=>p(228)(23),clock=>clock,reset=>reset,s=>p(280)(23),cout=>p(281)(24));
FA_ff_9464:FAff port map(x=>p(226)(24),y=>p(227)(24),Cin=>p(228)(24),clock=>clock,reset=>reset,s=>p(280)(24),cout=>p(281)(25));
FA_ff_9465:FAff port map(x=>p(226)(25),y=>p(227)(25),Cin=>p(228)(25),clock=>clock,reset=>reset,s=>p(280)(25),cout=>p(281)(26));
FA_ff_9466:FAff port map(x=>p(226)(26),y=>p(227)(26),Cin=>p(228)(26),clock=>clock,reset=>reset,s=>p(280)(26),cout=>p(281)(27));
FA_ff_9467:FAff port map(x=>p(226)(27),y=>p(227)(27),Cin=>p(228)(27),clock=>clock,reset=>reset,s=>p(280)(27),cout=>p(281)(28));
FA_ff_9468:FAff port map(x=>p(226)(28),y=>p(227)(28),Cin=>p(228)(28),clock=>clock,reset=>reset,s=>p(280)(28),cout=>p(281)(29));
FA_ff_9469:FAff port map(x=>p(226)(29),y=>p(227)(29),Cin=>p(228)(29),clock=>clock,reset=>reset,s=>p(280)(29),cout=>p(281)(30));
FA_ff_9470:FAff port map(x=>p(226)(30),y=>p(227)(30),Cin=>p(228)(30),clock=>clock,reset=>reset,s=>p(280)(30),cout=>p(281)(31));
FA_ff_9471:FAff port map(x=>p(226)(31),y=>p(227)(31),Cin=>p(228)(31),clock=>clock,reset=>reset,s=>p(280)(31),cout=>p(281)(32));
FA_ff_9472:FAff port map(x=>p(226)(32),y=>p(227)(32),Cin=>p(228)(32),clock=>clock,reset=>reset,s=>p(280)(32),cout=>p(281)(33));
FA_ff_9473:FAff port map(x=>p(226)(33),y=>p(227)(33),Cin=>p(228)(33),clock=>clock,reset=>reset,s=>p(280)(33),cout=>p(281)(34));
FA_ff_9474:FAff port map(x=>p(226)(34),y=>p(227)(34),Cin=>p(228)(34),clock=>clock,reset=>reset,s=>p(280)(34),cout=>p(281)(35));
FA_ff_9475:FAff port map(x=>p(226)(35),y=>p(227)(35),Cin=>p(228)(35),clock=>clock,reset=>reset,s=>p(280)(35),cout=>p(281)(36));
FA_ff_9476:FAff port map(x=>p(226)(36),y=>p(227)(36),Cin=>p(228)(36),clock=>clock,reset=>reset,s=>p(280)(36),cout=>p(281)(37));
FA_ff_9477:FAff port map(x=>p(226)(37),y=>p(227)(37),Cin=>p(228)(37),clock=>clock,reset=>reset,s=>p(280)(37),cout=>p(281)(38));
FA_ff_9478:FAff port map(x=>p(226)(38),y=>p(227)(38),Cin=>p(228)(38),clock=>clock,reset=>reset,s=>p(280)(38),cout=>p(281)(39));
FA_ff_9479:FAff port map(x=>p(226)(39),y=>p(227)(39),Cin=>p(228)(39),clock=>clock,reset=>reset,s=>p(280)(39),cout=>p(281)(40));
FA_ff_9480:FAff port map(x=>p(226)(40),y=>p(227)(40),Cin=>p(228)(40),clock=>clock,reset=>reset,s=>p(280)(40),cout=>p(281)(41));
FA_ff_9481:FAff port map(x=>p(226)(41),y=>p(227)(41),Cin=>p(228)(41),clock=>clock,reset=>reset,s=>p(280)(41),cout=>p(281)(42));
FA_ff_9482:FAff port map(x=>p(226)(42),y=>p(227)(42),Cin=>p(228)(42),clock=>clock,reset=>reset,s=>p(280)(42),cout=>p(281)(43));
FA_ff_9483:FAff port map(x=>p(226)(43),y=>p(227)(43),Cin=>p(228)(43),clock=>clock,reset=>reset,s=>p(280)(43),cout=>p(281)(44));
FA_ff_9484:FAff port map(x=>p(226)(44),y=>p(227)(44),Cin=>p(228)(44),clock=>clock,reset=>reset,s=>p(280)(44),cout=>p(281)(45));
FA_ff_9485:FAff port map(x=>p(226)(45),y=>p(227)(45),Cin=>p(228)(45),clock=>clock,reset=>reset,s=>p(280)(45),cout=>p(281)(46));
FA_ff_9486:FAff port map(x=>p(226)(46),y=>p(227)(46),Cin=>p(228)(46),clock=>clock,reset=>reset,s=>p(280)(46),cout=>p(281)(47));
FA_ff_9487:FAff port map(x=>p(226)(47),y=>p(227)(47),Cin=>p(228)(47),clock=>clock,reset=>reset,s=>p(280)(47),cout=>p(281)(48));
FA_ff_9488:FAff port map(x=>p(226)(48),y=>p(227)(48),Cin=>p(228)(48),clock=>clock,reset=>reset,s=>p(280)(48),cout=>p(281)(49));
FA_ff_9489:FAff port map(x=>p(226)(49),y=>p(227)(49),Cin=>p(228)(49),clock=>clock,reset=>reset,s=>p(280)(49),cout=>p(281)(50));
FA_ff_9490:FAff port map(x=>p(226)(50),y=>p(227)(50),Cin=>p(228)(50),clock=>clock,reset=>reset,s=>p(280)(50),cout=>p(281)(51));
FA_ff_9491:FAff port map(x=>p(226)(51),y=>p(227)(51),Cin=>p(228)(51),clock=>clock,reset=>reset,s=>p(280)(51),cout=>p(281)(52));
FA_ff_9492:FAff port map(x=>p(226)(52),y=>p(227)(52),Cin=>p(228)(52),clock=>clock,reset=>reset,s=>p(280)(52),cout=>p(281)(53));
FA_ff_9493:FAff port map(x=>p(226)(53),y=>p(227)(53),Cin=>p(228)(53),clock=>clock,reset=>reset,s=>p(280)(53),cout=>p(281)(54));
FA_ff_9494:FAff port map(x=>p(226)(54),y=>p(227)(54),Cin=>p(228)(54),clock=>clock,reset=>reset,s=>p(280)(54),cout=>p(281)(55));
FA_ff_9495:FAff port map(x=>p(226)(55),y=>p(227)(55),Cin=>p(228)(55),clock=>clock,reset=>reset,s=>p(280)(55),cout=>p(281)(56));
FA_ff_9496:FAff port map(x=>p(226)(56),y=>p(227)(56),Cin=>p(228)(56),clock=>clock,reset=>reset,s=>p(280)(56),cout=>p(281)(57));
FA_ff_9497:FAff port map(x=>p(226)(57),y=>p(227)(57),Cin=>p(228)(57),clock=>clock,reset=>reset,s=>p(280)(57),cout=>p(281)(58));
FA_ff_9498:FAff port map(x=>p(226)(58),y=>p(227)(58),Cin=>p(228)(58),clock=>clock,reset=>reset,s=>p(280)(58),cout=>p(281)(59));
FA_ff_9499:FAff port map(x=>p(226)(59),y=>p(227)(59),Cin=>p(228)(59),clock=>clock,reset=>reset,s=>p(280)(59),cout=>p(281)(60));
FA_ff_9500:FAff port map(x=>p(226)(60),y=>p(227)(60),Cin=>p(228)(60),clock=>clock,reset=>reset,s=>p(280)(60),cout=>p(281)(61));
FA_ff_9501:FAff port map(x=>p(226)(61),y=>p(227)(61),Cin=>p(228)(61),clock=>clock,reset=>reset,s=>p(280)(61),cout=>p(281)(62));
FA_ff_9502:FAff port map(x=>p(226)(62),y=>p(227)(62),Cin=>p(228)(62),clock=>clock,reset=>reset,s=>p(280)(62),cout=>p(281)(63));
FA_ff_9503:FAff port map(x=>p(226)(63),y=>p(227)(63),Cin=>p(228)(63),clock=>clock,reset=>reset,s=>p(280)(63),cout=>p(281)(64));
FA_ff_9504:FAff port map(x=>p(226)(64),y=>p(227)(64),Cin=>p(228)(64),clock=>clock,reset=>reset,s=>p(280)(64),cout=>p(281)(65));
FA_ff_9505:FAff port map(x=>p(226)(65),y=>p(227)(65),Cin=>p(228)(65),clock=>clock,reset=>reset,s=>p(280)(65),cout=>p(281)(66));
FA_ff_9506:FAff port map(x=>p(226)(66),y=>p(227)(66),Cin=>p(228)(66),clock=>clock,reset=>reset,s=>p(280)(66),cout=>p(281)(67));
FA_ff_9507:FAff port map(x=>p(226)(67),y=>p(227)(67),Cin=>p(228)(67),clock=>clock,reset=>reset,s=>p(280)(67),cout=>p(281)(68));
FA_ff_9508:FAff port map(x=>p(226)(68),y=>p(227)(68),Cin=>p(228)(68),clock=>clock,reset=>reset,s=>p(280)(68),cout=>p(281)(69));
FA_ff_9509:FAff port map(x=>p(226)(69),y=>p(227)(69),Cin=>p(228)(69),clock=>clock,reset=>reset,s=>p(280)(69),cout=>p(281)(70));
FA_ff_9510:FAff port map(x=>p(226)(70),y=>p(227)(70),Cin=>p(228)(70),clock=>clock,reset=>reset,s=>p(280)(70),cout=>p(281)(71));
FA_ff_9511:FAff port map(x=>p(226)(71),y=>p(227)(71),Cin=>p(228)(71),clock=>clock,reset=>reset,s=>p(280)(71),cout=>p(281)(72));
FA_ff_9512:FAff port map(x=>p(226)(72),y=>p(227)(72),Cin=>p(228)(72),clock=>clock,reset=>reset,s=>p(280)(72),cout=>p(281)(73));
FA_ff_9513:FAff port map(x=>p(226)(73),y=>p(227)(73),Cin=>p(228)(73),clock=>clock,reset=>reset,s=>p(280)(73),cout=>p(281)(74));
FA_ff_9514:FAff port map(x=>p(226)(74),y=>p(227)(74),Cin=>p(228)(74),clock=>clock,reset=>reset,s=>p(280)(74),cout=>p(281)(75));
FA_ff_9515:FAff port map(x=>p(226)(75),y=>p(227)(75),Cin=>p(228)(75),clock=>clock,reset=>reset,s=>p(280)(75),cout=>p(281)(76));
FA_ff_9516:FAff port map(x=>p(226)(76),y=>p(227)(76),Cin=>p(228)(76),clock=>clock,reset=>reset,s=>p(280)(76),cout=>p(281)(77));
FA_ff_9517:FAff port map(x=>p(226)(77),y=>p(227)(77),Cin=>p(228)(77),clock=>clock,reset=>reset,s=>p(280)(77),cout=>p(281)(78));
FA_ff_9518:FAff port map(x=>p(226)(78),y=>p(227)(78),Cin=>p(228)(78),clock=>clock,reset=>reset,s=>p(280)(78),cout=>p(281)(79));
FA_ff_9519:FAff port map(x=>p(226)(79),y=>p(227)(79),Cin=>p(228)(79),clock=>clock,reset=>reset,s=>p(280)(79),cout=>p(281)(80));
FA_ff_9520:FAff port map(x=>p(226)(80),y=>p(227)(80),Cin=>p(228)(80),clock=>clock,reset=>reset,s=>p(280)(80),cout=>p(281)(81));
FA_ff_9521:FAff port map(x=>p(226)(81),y=>p(227)(81),Cin=>p(228)(81),clock=>clock,reset=>reset,s=>p(280)(81),cout=>p(281)(82));
FA_ff_9522:FAff port map(x=>p(226)(82),y=>p(227)(82),Cin=>p(228)(82),clock=>clock,reset=>reset,s=>p(280)(82),cout=>p(281)(83));
FA_ff_9523:FAff port map(x=>p(226)(83),y=>p(227)(83),Cin=>p(228)(83),clock=>clock,reset=>reset,s=>p(280)(83),cout=>p(281)(84));
FA_ff_9524:FAff port map(x=>p(226)(84),y=>p(227)(84),Cin=>p(228)(84),clock=>clock,reset=>reset,s=>p(280)(84),cout=>p(281)(85));
FA_ff_9525:FAff port map(x=>p(226)(85),y=>p(227)(85),Cin=>p(228)(85),clock=>clock,reset=>reset,s=>p(280)(85),cout=>p(281)(86));
FA_ff_9526:FAff port map(x=>p(226)(86),y=>p(227)(86),Cin=>p(228)(86),clock=>clock,reset=>reset,s=>p(280)(86),cout=>p(281)(87));
FA_ff_9527:FAff port map(x=>p(226)(87),y=>p(227)(87),Cin=>p(228)(87),clock=>clock,reset=>reset,s=>p(280)(87),cout=>p(281)(88));
FA_ff_9528:FAff port map(x=>p(226)(88),y=>p(227)(88),Cin=>p(228)(88),clock=>clock,reset=>reset,s=>p(280)(88),cout=>p(281)(89));
FA_ff_9529:FAff port map(x=>p(226)(89),y=>p(227)(89),Cin=>p(228)(89),clock=>clock,reset=>reset,s=>p(280)(89),cout=>p(281)(90));
FA_ff_9530:FAff port map(x=>p(226)(90),y=>p(227)(90),Cin=>p(228)(90),clock=>clock,reset=>reset,s=>p(280)(90),cout=>p(281)(91));
FA_ff_9531:FAff port map(x=>p(226)(91),y=>p(227)(91),Cin=>p(228)(91),clock=>clock,reset=>reset,s=>p(280)(91),cout=>p(281)(92));
FA_ff_9532:FAff port map(x=>p(226)(92),y=>p(227)(92),Cin=>p(228)(92),clock=>clock,reset=>reset,s=>p(280)(92),cout=>p(281)(93));
FA_ff_9533:FAff port map(x=>p(226)(93),y=>p(227)(93),Cin=>p(228)(93),clock=>clock,reset=>reset,s=>p(280)(93),cout=>p(281)(94));
FA_ff_9534:FAff port map(x=>p(226)(94),y=>p(227)(94),Cin=>p(228)(94),clock=>clock,reset=>reset,s=>p(280)(94),cout=>p(281)(95));
FA_ff_9535:FAff port map(x=>p(226)(95),y=>p(227)(95),Cin=>p(228)(95),clock=>clock,reset=>reset,s=>p(280)(95),cout=>p(281)(96));
FA_ff_9536:FAff port map(x=>p(226)(96),y=>p(227)(96),Cin=>p(228)(96),clock=>clock,reset=>reset,s=>p(280)(96),cout=>p(281)(97));
FA_ff_9537:FAff port map(x=>p(226)(97),y=>p(227)(97),Cin=>p(228)(97),clock=>clock,reset=>reset,s=>p(280)(97),cout=>p(281)(98));
FA_ff_9538:FAff port map(x=>p(226)(98),y=>p(227)(98),Cin=>p(228)(98),clock=>clock,reset=>reset,s=>p(280)(98),cout=>p(281)(99));
FA_ff_9539:FAff port map(x=>p(226)(99),y=>p(227)(99),Cin=>p(228)(99),clock=>clock,reset=>reset,s=>p(280)(99),cout=>p(281)(100));
FA_ff_9540:FAff port map(x=>p(226)(100),y=>p(227)(100),Cin=>p(228)(100),clock=>clock,reset=>reset,s=>p(280)(100),cout=>p(281)(101));
FA_ff_9541:FAff port map(x=>p(226)(101),y=>p(227)(101),Cin=>p(228)(101),clock=>clock,reset=>reset,s=>p(280)(101),cout=>p(281)(102));
FA_ff_9542:FAff port map(x=>p(226)(102),y=>p(227)(102),Cin=>p(228)(102),clock=>clock,reset=>reset,s=>p(280)(102),cout=>p(281)(103));
FA_ff_9543:FAff port map(x=>p(226)(103),y=>p(227)(103),Cin=>p(228)(103),clock=>clock,reset=>reset,s=>p(280)(103),cout=>p(281)(104));
FA_ff_9544:FAff port map(x=>p(226)(104),y=>p(227)(104),Cin=>p(228)(104),clock=>clock,reset=>reset,s=>p(280)(104),cout=>p(281)(105));
FA_ff_9545:FAff port map(x=>p(226)(105),y=>p(227)(105),Cin=>p(228)(105),clock=>clock,reset=>reset,s=>p(280)(105),cout=>p(281)(106));
FA_ff_9546:FAff port map(x=>p(226)(106),y=>p(227)(106),Cin=>p(228)(106),clock=>clock,reset=>reset,s=>p(280)(106),cout=>p(281)(107));
FA_ff_9547:FAff port map(x=>p(226)(107),y=>p(227)(107),Cin=>p(228)(107),clock=>clock,reset=>reset,s=>p(280)(107),cout=>p(281)(108));
FA_ff_9548:FAff port map(x=>p(226)(108),y=>p(227)(108),Cin=>p(228)(108),clock=>clock,reset=>reset,s=>p(280)(108),cout=>p(281)(109));
FA_ff_9549:FAff port map(x=>p(226)(109),y=>p(227)(109),Cin=>p(228)(109),clock=>clock,reset=>reset,s=>p(280)(109),cout=>p(281)(110));
FA_ff_9550:FAff port map(x=>p(226)(110),y=>p(227)(110),Cin=>p(228)(110),clock=>clock,reset=>reset,s=>p(280)(110),cout=>p(281)(111));
FA_ff_9551:FAff port map(x=>p(226)(111),y=>p(227)(111),Cin=>p(228)(111),clock=>clock,reset=>reset,s=>p(280)(111),cout=>p(281)(112));
FA_ff_9552:FAff port map(x=>p(226)(112),y=>p(227)(112),Cin=>p(228)(112),clock=>clock,reset=>reset,s=>p(280)(112),cout=>p(281)(113));
FA_ff_9553:FAff port map(x=>p(226)(113),y=>p(227)(113),Cin=>p(228)(113),clock=>clock,reset=>reset,s=>p(280)(113),cout=>p(281)(114));
FA_ff_9554:FAff port map(x=>p(226)(114),y=>p(227)(114),Cin=>p(228)(114),clock=>clock,reset=>reset,s=>p(280)(114),cout=>p(281)(115));
FA_ff_9555:FAff port map(x=>p(226)(115),y=>p(227)(115),Cin=>p(228)(115),clock=>clock,reset=>reset,s=>p(280)(115),cout=>p(281)(116));
FA_ff_9556:FAff port map(x=>p(226)(116),y=>p(227)(116),Cin=>p(228)(116),clock=>clock,reset=>reset,s=>p(280)(116),cout=>p(281)(117));
FA_ff_9557:FAff port map(x=>p(226)(117),y=>p(227)(117),Cin=>p(228)(117),clock=>clock,reset=>reset,s=>p(280)(117),cout=>p(281)(118));
FA_ff_9558:FAff port map(x=>p(226)(118),y=>p(227)(118),Cin=>p(228)(118),clock=>clock,reset=>reset,s=>p(280)(118),cout=>p(281)(119));
FA_ff_9559:FAff port map(x=>p(226)(119),y=>p(227)(119),Cin=>p(228)(119),clock=>clock,reset=>reset,s=>p(280)(119),cout=>p(281)(120));
FA_ff_9560:FAff port map(x=>p(226)(120),y=>p(227)(120),Cin=>p(228)(120),clock=>clock,reset=>reset,s=>p(280)(120),cout=>p(281)(121));
FA_ff_9561:FAff port map(x=>p(226)(121),y=>p(227)(121),Cin=>p(228)(121),clock=>clock,reset=>reset,s=>p(280)(121),cout=>p(281)(122));
FA_ff_9562:FAff port map(x=>p(226)(122),y=>p(227)(122),Cin=>p(228)(122),clock=>clock,reset=>reset,s=>p(280)(122),cout=>p(281)(123));
FA_ff_9563:FAff port map(x=>p(226)(123),y=>p(227)(123),Cin=>p(228)(123),clock=>clock,reset=>reset,s=>p(280)(123),cout=>p(281)(124));
FA_ff_9564:FAff port map(x=>p(226)(124),y=>p(227)(124),Cin=>p(228)(124),clock=>clock,reset=>reset,s=>p(280)(124),cout=>p(281)(125));
FA_ff_9565:FAff port map(x=>p(226)(125),y=>p(227)(125),Cin=>p(228)(125),clock=>clock,reset=>reset,s=>p(280)(125),cout=>p(281)(126));
FA_ff_9566:FAff port map(x=>p(226)(126),y=>p(227)(126),Cin=>p(228)(126),clock=>clock,reset=>reset,s=>p(280)(126),cout=>p(281)(127));
FA_ff_9567:FAff port map(x=>p(226)(127),y=>p(227)(127),Cin=>p(228)(127),clock=>clock,reset=>reset,s=>p(280)(127),cout=>p(281)(128));
FA_ff_9568:FAff port map(x=>p(226)(128),y=>p(227)(128),Cin=>p(228)(128),clock=>clock,reset=>reset,s=>p(280)(128),cout=>p(281)(129));
p(282)(0)<=p(230)(0);
HA_ff_34:HAff port map(x=>p(230)(1),y=>p(231)(1),clock=>clock,reset=>reset,s=>p(282)(1),c=>p(283)(2));
FA_ff_9569:FAff port map(x=>p(229)(2),y=>p(230)(2),Cin=>p(231)(2),clock=>clock,reset=>reset,s=>p(282)(2),cout=>p(283)(3));
FA_ff_9570:FAff port map(x=>p(229)(3),y=>p(230)(3),Cin=>p(231)(3),clock=>clock,reset=>reset,s=>p(282)(3),cout=>p(283)(4));
FA_ff_9571:FAff port map(x=>p(229)(4),y=>p(230)(4),Cin=>p(231)(4),clock=>clock,reset=>reset,s=>p(282)(4),cout=>p(283)(5));
FA_ff_9572:FAff port map(x=>p(229)(5),y=>p(230)(5),Cin=>p(231)(5),clock=>clock,reset=>reset,s=>p(282)(5),cout=>p(283)(6));
FA_ff_9573:FAff port map(x=>p(229)(6),y=>p(230)(6),Cin=>p(231)(6),clock=>clock,reset=>reset,s=>p(282)(6),cout=>p(283)(7));
FA_ff_9574:FAff port map(x=>p(229)(7),y=>p(230)(7),Cin=>p(231)(7),clock=>clock,reset=>reset,s=>p(282)(7),cout=>p(283)(8));
FA_ff_9575:FAff port map(x=>p(229)(8),y=>p(230)(8),Cin=>p(231)(8),clock=>clock,reset=>reset,s=>p(282)(8),cout=>p(283)(9));
FA_ff_9576:FAff port map(x=>p(229)(9),y=>p(230)(9),Cin=>p(231)(9),clock=>clock,reset=>reset,s=>p(282)(9),cout=>p(283)(10));
FA_ff_9577:FAff port map(x=>p(229)(10),y=>p(230)(10),Cin=>p(231)(10),clock=>clock,reset=>reset,s=>p(282)(10),cout=>p(283)(11));
FA_ff_9578:FAff port map(x=>p(229)(11),y=>p(230)(11),Cin=>p(231)(11),clock=>clock,reset=>reset,s=>p(282)(11),cout=>p(283)(12));
FA_ff_9579:FAff port map(x=>p(229)(12),y=>p(230)(12),Cin=>p(231)(12),clock=>clock,reset=>reset,s=>p(282)(12),cout=>p(283)(13));
FA_ff_9580:FAff port map(x=>p(229)(13),y=>p(230)(13),Cin=>p(231)(13),clock=>clock,reset=>reset,s=>p(282)(13),cout=>p(283)(14));
FA_ff_9581:FAff port map(x=>p(229)(14),y=>p(230)(14),Cin=>p(231)(14),clock=>clock,reset=>reset,s=>p(282)(14),cout=>p(283)(15));
FA_ff_9582:FAff port map(x=>p(229)(15),y=>p(230)(15),Cin=>p(231)(15),clock=>clock,reset=>reset,s=>p(282)(15),cout=>p(283)(16));
FA_ff_9583:FAff port map(x=>p(229)(16),y=>p(230)(16),Cin=>p(231)(16),clock=>clock,reset=>reset,s=>p(282)(16),cout=>p(283)(17));
FA_ff_9584:FAff port map(x=>p(229)(17),y=>p(230)(17),Cin=>p(231)(17),clock=>clock,reset=>reset,s=>p(282)(17),cout=>p(283)(18));
FA_ff_9585:FAff port map(x=>p(229)(18),y=>p(230)(18),Cin=>p(231)(18),clock=>clock,reset=>reset,s=>p(282)(18),cout=>p(283)(19));
FA_ff_9586:FAff port map(x=>p(229)(19),y=>p(230)(19),Cin=>p(231)(19),clock=>clock,reset=>reset,s=>p(282)(19),cout=>p(283)(20));
FA_ff_9587:FAff port map(x=>p(229)(20),y=>p(230)(20),Cin=>p(231)(20),clock=>clock,reset=>reset,s=>p(282)(20),cout=>p(283)(21));
FA_ff_9588:FAff port map(x=>p(229)(21),y=>p(230)(21),Cin=>p(231)(21),clock=>clock,reset=>reset,s=>p(282)(21),cout=>p(283)(22));
FA_ff_9589:FAff port map(x=>p(229)(22),y=>p(230)(22),Cin=>p(231)(22),clock=>clock,reset=>reset,s=>p(282)(22),cout=>p(283)(23));
FA_ff_9590:FAff port map(x=>p(229)(23),y=>p(230)(23),Cin=>p(231)(23),clock=>clock,reset=>reset,s=>p(282)(23),cout=>p(283)(24));
FA_ff_9591:FAff port map(x=>p(229)(24),y=>p(230)(24),Cin=>p(231)(24),clock=>clock,reset=>reset,s=>p(282)(24),cout=>p(283)(25));
FA_ff_9592:FAff port map(x=>p(229)(25),y=>p(230)(25),Cin=>p(231)(25),clock=>clock,reset=>reset,s=>p(282)(25),cout=>p(283)(26));
FA_ff_9593:FAff port map(x=>p(229)(26),y=>p(230)(26),Cin=>p(231)(26),clock=>clock,reset=>reset,s=>p(282)(26),cout=>p(283)(27));
FA_ff_9594:FAff port map(x=>p(229)(27),y=>p(230)(27),Cin=>p(231)(27),clock=>clock,reset=>reset,s=>p(282)(27),cout=>p(283)(28));
FA_ff_9595:FAff port map(x=>p(229)(28),y=>p(230)(28),Cin=>p(231)(28),clock=>clock,reset=>reset,s=>p(282)(28),cout=>p(283)(29));
FA_ff_9596:FAff port map(x=>p(229)(29),y=>p(230)(29),Cin=>p(231)(29),clock=>clock,reset=>reset,s=>p(282)(29),cout=>p(283)(30));
FA_ff_9597:FAff port map(x=>p(229)(30),y=>p(230)(30),Cin=>p(231)(30),clock=>clock,reset=>reset,s=>p(282)(30),cout=>p(283)(31));
FA_ff_9598:FAff port map(x=>p(229)(31),y=>p(230)(31),Cin=>p(231)(31),clock=>clock,reset=>reset,s=>p(282)(31),cout=>p(283)(32));
FA_ff_9599:FAff port map(x=>p(229)(32),y=>p(230)(32),Cin=>p(231)(32),clock=>clock,reset=>reset,s=>p(282)(32),cout=>p(283)(33));
FA_ff_9600:FAff port map(x=>p(229)(33),y=>p(230)(33),Cin=>p(231)(33),clock=>clock,reset=>reset,s=>p(282)(33),cout=>p(283)(34));
FA_ff_9601:FAff port map(x=>p(229)(34),y=>p(230)(34),Cin=>p(231)(34),clock=>clock,reset=>reset,s=>p(282)(34),cout=>p(283)(35));
FA_ff_9602:FAff port map(x=>p(229)(35),y=>p(230)(35),Cin=>p(231)(35),clock=>clock,reset=>reset,s=>p(282)(35),cout=>p(283)(36));
FA_ff_9603:FAff port map(x=>p(229)(36),y=>p(230)(36),Cin=>p(231)(36),clock=>clock,reset=>reset,s=>p(282)(36),cout=>p(283)(37));
FA_ff_9604:FAff port map(x=>p(229)(37),y=>p(230)(37),Cin=>p(231)(37),clock=>clock,reset=>reset,s=>p(282)(37),cout=>p(283)(38));
FA_ff_9605:FAff port map(x=>p(229)(38),y=>p(230)(38),Cin=>p(231)(38),clock=>clock,reset=>reset,s=>p(282)(38),cout=>p(283)(39));
FA_ff_9606:FAff port map(x=>p(229)(39),y=>p(230)(39),Cin=>p(231)(39),clock=>clock,reset=>reset,s=>p(282)(39),cout=>p(283)(40));
FA_ff_9607:FAff port map(x=>p(229)(40),y=>p(230)(40),Cin=>p(231)(40),clock=>clock,reset=>reset,s=>p(282)(40),cout=>p(283)(41));
FA_ff_9608:FAff port map(x=>p(229)(41),y=>p(230)(41),Cin=>p(231)(41),clock=>clock,reset=>reset,s=>p(282)(41),cout=>p(283)(42));
FA_ff_9609:FAff port map(x=>p(229)(42),y=>p(230)(42),Cin=>p(231)(42),clock=>clock,reset=>reset,s=>p(282)(42),cout=>p(283)(43));
FA_ff_9610:FAff port map(x=>p(229)(43),y=>p(230)(43),Cin=>p(231)(43),clock=>clock,reset=>reset,s=>p(282)(43),cout=>p(283)(44));
FA_ff_9611:FAff port map(x=>p(229)(44),y=>p(230)(44),Cin=>p(231)(44),clock=>clock,reset=>reset,s=>p(282)(44),cout=>p(283)(45));
FA_ff_9612:FAff port map(x=>p(229)(45),y=>p(230)(45),Cin=>p(231)(45),clock=>clock,reset=>reset,s=>p(282)(45),cout=>p(283)(46));
FA_ff_9613:FAff port map(x=>p(229)(46),y=>p(230)(46),Cin=>p(231)(46),clock=>clock,reset=>reset,s=>p(282)(46),cout=>p(283)(47));
FA_ff_9614:FAff port map(x=>p(229)(47),y=>p(230)(47),Cin=>p(231)(47),clock=>clock,reset=>reset,s=>p(282)(47),cout=>p(283)(48));
FA_ff_9615:FAff port map(x=>p(229)(48),y=>p(230)(48),Cin=>p(231)(48),clock=>clock,reset=>reset,s=>p(282)(48),cout=>p(283)(49));
FA_ff_9616:FAff port map(x=>p(229)(49),y=>p(230)(49),Cin=>p(231)(49),clock=>clock,reset=>reset,s=>p(282)(49),cout=>p(283)(50));
FA_ff_9617:FAff port map(x=>p(229)(50),y=>p(230)(50),Cin=>p(231)(50),clock=>clock,reset=>reset,s=>p(282)(50),cout=>p(283)(51));
FA_ff_9618:FAff port map(x=>p(229)(51),y=>p(230)(51),Cin=>p(231)(51),clock=>clock,reset=>reset,s=>p(282)(51),cout=>p(283)(52));
FA_ff_9619:FAff port map(x=>p(229)(52),y=>p(230)(52),Cin=>p(231)(52),clock=>clock,reset=>reset,s=>p(282)(52),cout=>p(283)(53));
FA_ff_9620:FAff port map(x=>p(229)(53),y=>p(230)(53),Cin=>p(231)(53),clock=>clock,reset=>reset,s=>p(282)(53),cout=>p(283)(54));
FA_ff_9621:FAff port map(x=>p(229)(54),y=>p(230)(54),Cin=>p(231)(54),clock=>clock,reset=>reset,s=>p(282)(54),cout=>p(283)(55));
FA_ff_9622:FAff port map(x=>p(229)(55),y=>p(230)(55),Cin=>p(231)(55),clock=>clock,reset=>reset,s=>p(282)(55),cout=>p(283)(56));
FA_ff_9623:FAff port map(x=>p(229)(56),y=>p(230)(56),Cin=>p(231)(56),clock=>clock,reset=>reset,s=>p(282)(56),cout=>p(283)(57));
FA_ff_9624:FAff port map(x=>p(229)(57),y=>p(230)(57),Cin=>p(231)(57),clock=>clock,reset=>reset,s=>p(282)(57),cout=>p(283)(58));
FA_ff_9625:FAff port map(x=>p(229)(58),y=>p(230)(58),Cin=>p(231)(58),clock=>clock,reset=>reset,s=>p(282)(58),cout=>p(283)(59));
FA_ff_9626:FAff port map(x=>p(229)(59),y=>p(230)(59),Cin=>p(231)(59),clock=>clock,reset=>reset,s=>p(282)(59),cout=>p(283)(60));
FA_ff_9627:FAff port map(x=>p(229)(60),y=>p(230)(60),Cin=>p(231)(60),clock=>clock,reset=>reset,s=>p(282)(60),cout=>p(283)(61));
FA_ff_9628:FAff port map(x=>p(229)(61),y=>p(230)(61),Cin=>p(231)(61),clock=>clock,reset=>reset,s=>p(282)(61),cout=>p(283)(62));
FA_ff_9629:FAff port map(x=>p(229)(62),y=>p(230)(62),Cin=>p(231)(62),clock=>clock,reset=>reset,s=>p(282)(62),cout=>p(283)(63));
FA_ff_9630:FAff port map(x=>p(229)(63),y=>p(230)(63),Cin=>p(231)(63),clock=>clock,reset=>reset,s=>p(282)(63),cout=>p(283)(64));
FA_ff_9631:FAff port map(x=>p(229)(64),y=>p(230)(64),Cin=>p(231)(64),clock=>clock,reset=>reset,s=>p(282)(64),cout=>p(283)(65));
FA_ff_9632:FAff port map(x=>p(229)(65),y=>p(230)(65),Cin=>p(231)(65),clock=>clock,reset=>reset,s=>p(282)(65),cout=>p(283)(66));
FA_ff_9633:FAff port map(x=>p(229)(66),y=>p(230)(66),Cin=>p(231)(66),clock=>clock,reset=>reset,s=>p(282)(66),cout=>p(283)(67));
FA_ff_9634:FAff port map(x=>p(229)(67),y=>p(230)(67),Cin=>p(231)(67),clock=>clock,reset=>reset,s=>p(282)(67),cout=>p(283)(68));
FA_ff_9635:FAff port map(x=>p(229)(68),y=>p(230)(68),Cin=>p(231)(68),clock=>clock,reset=>reset,s=>p(282)(68),cout=>p(283)(69));
FA_ff_9636:FAff port map(x=>p(229)(69),y=>p(230)(69),Cin=>p(231)(69),clock=>clock,reset=>reset,s=>p(282)(69),cout=>p(283)(70));
FA_ff_9637:FAff port map(x=>p(229)(70),y=>p(230)(70),Cin=>p(231)(70),clock=>clock,reset=>reset,s=>p(282)(70),cout=>p(283)(71));
FA_ff_9638:FAff port map(x=>p(229)(71),y=>p(230)(71),Cin=>p(231)(71),clock=>clock,reset=>reset,s=>p(282)(71),cout=>p(283)(72));
FA_ff_9639:FAff port map(x=>p(229)(72),y=>p(230)(72),Cin=>p(231)(72),clock=>clock,reset=>reset,s=>p(282)(72),cout=>p(283)(73));
FA_ff_9640:FAff port map(x=>p(229)(73),y=>p(230)(73),Cin=>p(231)(73),clock=>clock,reset=>reset,s=>p(282)(73),cout=>p(283)(74));
FA_ff_9641:FAff port map(x=>p(229)(74),y=>p(230)(74),Cin=>p(231)(74),clock=>clock,reset=>reset,s=>p(282)(74),cout=>p(283)(75));
FA_ff_9642:FAff port map(x=>p(229)(75),y=>p(230)(75),Cin=>p(231)(75),clock=>clock,reset=>reset,s=>p(282)(75),cout=>p(283)(76));
FA_ff_9643:FAff port map(x=>p(229)(76),y=>p(230)(76),Cin=>p(231)(76),clock=>clock,reset=>reset,s=>p(282)(76),cout=>p(283)(77));
FA_ff_9644:FAff port map(x=>p(229)(77),y=>p(230)(77),Cin=>p(231)(77),clock=>clock,reset=>reset,s=>p(282)(77),cout=>p(283)(78));
FA_ff_9645:FAff port map(x=>p(229)(78),y=>p(230)(78),Cin=>p(231)(78),clock=>clock,reset=>reset,s=>p(282)(78),cout=>p(283)(79));
FA_ff_9646:FAff port map(x=>p(229)(79),y=>p(230)(79),Cin=>p(231)(79),clock=>clock,reset=>reset,s=>p(282)(79),cout=>p(283)(80));
FA_ff_9647:FAff port map(x=>p(229)(80),y=>p(230)(80),Cin=>p(231)(80),clock=>clock,reset=>reset,s=>p(282)(80),cout=>p(283)(81));
FA_ff_9648:FAff port map(x=>p(229)(81),y=>p(230)(81),Cin=>p(231)(81),clock=>clock,reset=>reset,s=>p(282)(81),cout=>p(283)(82));
FA_ff_9649:FAff port map(x=>p(229)(82),y=>p(230)(82),Cin=>p(231)(82),clock=>clock,reset=>reset,s=>p(282)(82),cout=>p(283)(83));
FA_ff_9650:FAff port map(x=>p(229)(83),y=>p(230)(83),Cin=>p(231)(83),clock=>clock,reset=>reset,s=>p(282)(83),cout=>p(283)(84));
FA_ff_9651:FAff port map(x=>p(229)(84),y=>p(230)(84),Cin=>p(231)(84),clock=>clock,reset=>reset,s=>p(282)(84),cout=>p(283)(85));
FA_ff_9652:FAff port map(x=>p(229)(85),y=>p(230)(85),Cin=>p(231)(85),clock=>clock,reset=>reset,s=>p(282)(85),cout=>p(283)(86));
FA_ff_9653:FAff port map(x=>p(229)(86),y=>p(230)(86),Cin=>p(231)(86),clock=>clock,reset=>reset,s=>p(282)(86),cout=>p(283)(87));
FA_ff_9654:FAff port map(x=>p(229)(87),y=>p(230)(87),Cin=>p(231)(87),clock=>clock,reset=>reset,s=>p(282)(87),cout=>p(283)(88));
FA_ff_9655:FAff port map(x=>p(229)(88),y=>p(230)(88),Cin=>p(231)(88),clock=>clock,reset=>reset,s=>p(282)(88),cout=>p(283)(89));
FA_ff_9656:FAff port map(x=>p(229)(89),y=>p(230)(89),Cin=>p(231)(89),clock=>clock,reset=>reset,s=>p(282)(89),cout=>p(283)(90));
FA_ff_9657:FAff port map(x=>p(229)(90),y=>p(230)(90),Cin=>p(231)(90),clock=>clock,reset=>reset,s=>p(282)(90),cout=>p(283)(91));
FA_ff_9658:FAff port map(x=>p(229)(91),y=>p(230)(91),Cin=>p(231)(91),clock=>clock,reset=>reset,s=>p(282)(91),cout=>p(283)(92));
FA_ff_9659:FAff port map(x=>p(229)(92),y=>p(230)(92),Cin=>p(231)(92),clock=>clock,reset=>reset,s=>p(282)(92),cout=>p(283)(93));
FA_ff_9660:FAff port map(x=>p(229)(93),y=>p(230)(93),Cin=>p(231)(93),clock=>clock,reset=>reset,s=>p(282)(93),cout=>p(283)(94));
FA_ff_9661:FAff port map(x=>p(229)(94),y=>p(230)(94),Cin=>p(231)(94),clock=>clock,reset=>reset,s=>p(282)(94),cout=>p(283)(95));
FA_ff_9662:FAff port map(x=>p(229)(95),y=>p(230)(95),Cin=>p(231)(95),clock=>clock,reset=>reset,s=>p(282)(95),cout=>p(283)(96));
FA_ff_9663:FAff port map(x=>p(229)(96),y=>p(230)(96),Cin=>p(231)(96),clock=>clock,reset=>reset,s=>p(282)(96),cout=>p(283)(97));
FA_ff_9664:FAff port map(x=>p(229)(97),y=>p(230)(97),Cin=>p(231)(97),clock=>clock,reset=>reset,s=>p(282)(97),cout=>p(283)(98));
FA_ff_9665:FAff port map(x=>p(229)(98),y=>p(230)(98),Cin=>p(231)(98),clock=>clock,reset=>reset,s=>p(282)(98),cout=>p(283)(99));
FA_ff_9666:FAff port map(x=>p(229)(99),y=>p(230)(99),Cin=>p(231)(99),clock=>clock,reset=>reset,s=>p(282)(99),cout=>p(283)(100));
FA_ff_9667:FAff port map(x=>p(229)(100),y=>p(230)(100),Cin=>p(231)(100),clock=>clock,reset=>reset,s=>p(282)(100),cout=>p(283)(101));
FA_ff_9668:FAff port map(x=>p(229)(101),y=>p(230)(101),Cin=>p(231)(101),clock=>clock,reset=>reset,s=>p(282)(101),cout=>p(283)(102));
FA_ff_9669:FAff port map(x=>p(229)(102),y=>p(230)(102),Cin=>p(231)(102),clock=>clock,reset=>reset,s=>p(282)(102),cout=>p(283)(103));
FA_ff_9670:FAff port map(x=>p(229)(103),y=>p(230)(103),Cin=>p(231)(103),clock=>clock,reset=>reset,s=>p(282)(103),cout=>p(283)(104));
FA_ff_9671:FAff port map(x=>p(229)(104),y=>p(230)(104),Cin=>p(231)(104),clock=>clock,reset=>reset,s=>p(282)(104),cout=>p(283)(105));
FA_ff_9672:FAff port map(x=>p(229)(105),y=>p(230)(105),Cin=>p(231)(105),clock=>clock,reset=>reset,s=>p(282)(105),cout=>p(283)(106));
FA_ff_9673:FAff port map(x=>p(229)(106),y=>p(230)(106),Cin=>p(231)(106),clock=>clock,reset=>reset,s=>p(282)(106),cout=>p(283)(107));
FA_ff_9674:FAff port map(x=>p(229)(107),y=>p(230)(107),Cin=>p(231)(107),clock=>clock,reset=>reset,s=>p(282)(107),cout=>p(283)(108));
FA_ff_9675:FAff port map(x=>p(229)(108),y=>p(230)(108),Cin=>p(231)(108),clock=>clock,reset=>reset,s=>p(282)(108),cout=>p(283)(109));
FA_ff_9676:FAff port map(x=>p(229)(109),y=>p(230)(109),Cin=>p(231)(109),clock=>clock,reset=>reset,s=>p(282)(109),cout=>p(283)(110));
FA_ff_9677:FAff port map(x=>p(229)(110),y=>p(230)(110),Cin=>p(231)(110),clock=>clock,reset=>reset,s=>p(282)(110),cout=>p(283)(111));
FA_ff_9678:FAff port map(x=>p(229)(111),y=>p(230)(111),Cin=>p(231)(111),clock=>clock,reset=>reset,s=>p(282)(111),cout=>p(283)(112));
FA_ff_9679:FAff port map(x=>p(229)(112),y=>p(230)(112),Cin=>p(231)(112),clock=>clock,reset=>reset,s=>p(282)(112),cout=>p(283)(113));
FA_ff_9680:FAff port map(x=>p(229)(113),y=>p(230)(113),Cin=>p(231)(113),clock=>clock,reset=>reset,s=>p(282)(113),cout=>p(283)(114));
FA_ff_9681:FAff port map(x=>p(229)(114),y=>p(230)(114),Cin=>p(231)(114),clock=>clock,reset=>reset,s=>p(282)(114),cout=>p(283)(115));
FA_ff_9682:FAff port map(x=>p(229)(115),y=>p(230)(115),Cin=>p(231)(115),clock=>clock,reset=>reset,s=>p(282)(115),cout=>p(283)(116));
FA_ff_9683:FAff port map(x=>p(229)(116),y=>p(230)(116),Cin=>p(231)(116),clock=>clock,reset=>reset,s=>p(282)(116),cout=>p(283)(117));
FA_ff_9684:FAff port map(x=>p(229)(117),y=>p(230)(117),Cin=>p(231)(117),clock=>clock,reset=>reset,s=>p(282)(117),cout=>p(283)(118));
FA_ff_9685:FAff port map(x=>p(229)(118),y=>p(230)(118),Cin=>p(231)(118),clock=>clock,reset=>reset,s=>p(282)(118),cout=>p(283)(119));
FA_ff_9686:FAff port map(x=>p(229)(119),y=>p(230)(119),Cin=>p(231)(119),clock=>clock,reset=>reset,s=>p(282)(119),cout=>p(283)(120));
FA_ff_9687:FAff port map(x=>p(229)(120),y=>p(230)(120),Cin=>p(231)(120),clock=>clock,reset=>reset,s=>p(282)(120),cout=>p(283)(121));
FA_ff_9688:FAff port map(x=>p(229)(121),y=>p(230)(121),Cin=>p(231)(121),clock=>clock,reset=>reset,s=>p(282)(121),cout=>p(283)(122));
FA_ff_9689:FAff port map(x=>p(229)(122),y=>p(230)(122),Cin=>p(231)(122),clock=>clock,reset=>reset,s=>p(282)(122),cout=>p(283)(123));
FA_ff_9690:FAff port map(x=>p(229)(123),y=>p(230)(123),Cin=>p(231)(123),clock=>clock,reset=>reset,s=>p(282)(123),cout=>p(283)(124));
FA_ff_9691:FAff port map(x=>p(229)(124),y=>p(230)(124),Cin=>p(231)(124),clock=>clock,reset=>reset,s=>p(282)(124),cout=>p(283)(125));
FA_ff_9692:FAff port map(x=>p(229)(125),y=>p(230)(125),Cin=>p(231)(125),clock=>clock,reset=>reset,s=>p(282)(125),cout=>p(283)(126));
FA_ff_9693:FAff port map(x=>p(229)(126),y=>p(230)(126),Cin=>p(231)(126),clock=>clock,reset=>reset,s=>p(282)(126),cout=>p(283)(127));
FA_ff_9694:FAff port map(x=>p(229)(127),y=>p(230)(127),Cin=>p(231)(127),clock=>clock,reset=>reset,s=>p(282)(127),cout=>p(283)(128));
FA_ff_9695:FAff port map(x=>p(229)(128),y=>p(230)(128),Cin=>p(231)(128),clock=>clock,reset=>reset,s=>p(282)(128),cout=>p(283)(129));
p(282)(129)<=p(229)(129);
HA_ff_35:HAff port map(x=>p(232)(0),y=>p(234)(0),clock=>clock,reset=>reset,s=>p(284)(0),c=>p(285)(1));
HA_ff_36:HAff port map(x=>p(232)(1),y=>p(234)(1),clock=>clock,reset=>reset,s=>p(284)(1),c=>p(285)(2));
FA_ff_9696:FAff port map(x=>p(232)(2),y=>p(233)(2),Cin=>p(234)(2),clock=>clock,reset=>reset,s=>p(284)(2),cout=>p(285)(3));
FA_ff_9697:FAff port map(x=>p(232)(3),y=>p(233)(3),Cin=>p(234)(3),clock=>clock,reset=>reset,s=>p(284)(3),cout=>p(285)(4));
FA_ff_9698:FAff port map(x=>p(232)(4),y=>p(233)(4),Cin=>p(234)(4),clock=>clock,reset=>reset,s=>p(284)(4),cout=>p(285)(5));
FA_ff_9699:FAff port map(x=>p(232)(5),y=>p(233)(5),Cin=>p(234)(5),clock=>clock,reset=>reset,s=>p(284)(5),cout=>p(285)(6));
FA_ff_9700:FAff port map(x=>p(232)(6),y=>p(233)(6),Cin=>p(234)(6),clock=>clock,reset=>reset,s=>p(284)(6),cout=>p(285)(7));
FA_ff_9701:FAff port map(x=>p(232)(7),y=>p(233)(7),Cin=>p(234)(7),clock=>clock,reset=>reset,s=>p(284)(7),cout=>p(285)(8));
FA_ff_9702:FAff port map(x=>p(232)(8),y=>p(233)(8),Cin=>p(234)(8),clock=>clock,reset=>reset,s=>p(284)(8),cout=>p(285)(9));
FA_ff_9703:FAff port map(x=>p(232)(9),y=>p(233)(9),Cin=>p(234)(9),clock=>clock,reset=>reset,s=>p(284)(9),cout=>p(285)(10));
FA_ff_9704:FAff port map(x=>p(232)(10),y=>p(233)(10),Cin=>p(234)(10),clock=>clock,reset=>reset,s=>p(284)(10),cout=>p(285)(11));
FA_ff_9705:FAff port map(x=>p(232)(11),y=>p(233)(11),Cin=>p(234)(11),clock=>clock,reset=>reset,s=>p(284)(11),cout=>p(285)(12));
FA_ff_9706:FAff port map(x=>p(232)(12),y=>p(233)(12),Cin=>p(234)(12),clock=>clock,reset=>reset,s=>p(284)(12),cout=>p(285)(13));
FA_ff_9707:FAff port map(x=>p(232)(13),y=>p(233)(13),Cin=>p(234)(13),clock=>clock,reset=>reset,s=>p(284)(13),cout=>p(285)(14));
FA_ff_9708:FAff port map(x=>p(232)(14),y=>p(233)(14),Cin=>p(234)(14),clock=>clock,reset=>reset,s=>p(284)(14),cout=>p(285)(15));
FA_ff_9709:FAff port map(x=>p(232)(15),y=>p(233)(15),Cin=>p(234)(15),clock=>clock,reset=>reset,s=>p(284)(15),cout=>p(285)(16));
FA_ff_9710:FAff port map(x=>p(232)(16),y=>p(233)(16),Cin=>p(234)(16),clock=>clock,reset=>reset,s=>p(284)(16),cout=>p(285)(17));
FA_ff_9711:FAff port map(x=>p(232)(17),y=>p(233)(17),Cin=>p(234)(17),clock=>clock,reset=>reset,s=>p(284)(17),cout=>p(285)(18));
FA_ff_9712:FAff port map(x=>p(232)(18),y=>p(233)(18),Cin=>p(234)(18),clock=>clock,reset=>reset,s=>p(284)(18),cout=>p(285)(19));
FA_ff_9713:FAff port map(x=>p(232)(19),y=>p(233)(19),Cin=>p(234)(19),clock=>clock,reset=>reset,s=>p(284)(19),cout=>p(285)(20));
FA_ff_9714:FAff port map(x=>p(232)(20),y=>p(233)(20),Cin=>p(234)(20),clock=>clock,reset=>reset,s=>p(284)(20),cout=>p(285)(21));
FA_ff_9715:FAff port map(x=>p(232)(21),y=>p(233)(21),Cin=>p(234)(21),clock=>clock,reset=>reset,s=>p(284)(21),cout=>p(285)(22));
FA_ff_9716:FAff port map(x=>p(232)(22),y=>p(233)(22),Cin=>p(234)(22),clock=>clock,reset=>reset,s=>p(284)(22),cout=>p(285)(23));
FA_ff_9717:FAff port map(x=>p(232)(23),y=>p(233)(23),Cin=>p(234)(23),clock=>clock,reset=>reset,s=>p(284)(23),cout=>p(285)(24));
FA_ff_9718:FAff port map(x=>p(232)(24),y=>p(233)(24),Cin=>p(234)(24),clock=>clock,reset=>reset,s=>p(284)(24),cout=>p(285)(25));
FA_ff_9719:FAff port map(x=>p(232)(25),y=>p(233)(25),Cin=>p(234)(25),clock=>clock,reset=>reset,s=>p(284)(25),cout=>p(285)(26));
FA_ff_9720:FAff port map(x=>p(232)(26),y=>p(233)(26),Cin=>p(234)(26),clock=>clock,reset=>reset,s=>p(284)(26),cout=>p(285)(27));
FA_ff_9721:FAff port map(x=>p(232)(27),y=>p(233)(27),Cin=>p(234)(27),clock=>clock,reset=>reset,s=>p(284)(27),cout=>p(285)(28));
FA_ff_9722:FAff port map(x=>p(232)(28),y=>p(233)(28),Cin=>p(234)(28),clock=>clock,reset=>reset,s=>p(284)(28),cout=>p(285)(29));
FA_ff_9723:FAff port map(x=>p(232)(29),y=>p(233)(29),Cin=>p(234)(29),clock=>clock,reset=>reset,s=>p(284)(29),cout=>p(285)(30));
FA_ff_9724:FAff port map(x=>p(232)(30),y=>p(233)(30),Cin=>p(234)(30),clock=>clock,reset=>reset,s=>p(284)(30),cout=>p(285)(31));
FA_ff_9725:FAff port map(x=>p(232)(31),y=>p(233)(31),Cin=>p(234)(31),clock=>clock,reset=>reset,s=>p(284)(31),cout=>p(285)(32));
FA_ff_9726:FAff port map(x=>p(232)(32),y=>p(233)(32),Cin=>p(234)(32),clock=>clock,reset=>reset,s=>p(284)(32),cout=>p(285)(33));
FA_ff_9727:FAff port map(x=>p(232)(33),y=>p(233)(33),Cin=>p(234)(33),clock=>clock,reset=>reset,s=>p(284)(33),cout=>p(285)(34));
FA_ff_9728:FAff port map(x=>p(232)(34),y=>p(233)(34),Cin=>p(234)(34),clock=>clock,reset=>reset,s=>p(284)(34),cout=>p(285)(35));
FA_ff_9729:FAff port map(x=>p(232)(35),y=>p(233)(35),Cin=>p(234)(35),clock=>clock,reset=>reset,s=>p(284)(35),cout=>p(285)(36));
FA_ff_9730:FAff port map(x=>p(232)(36),y=>p(233)(36),Cin=>p(234)(36),clock=>clock,reset=>reset,s=>p(284)(36),cout=>p(285)(37));
FA_ff_9731:FAff port map(x=>p(232)(37),y=>p(233)(37),Cin=>p(234)(37),clock=>clock,reset=>reset,s=>p(284)(37),cout=>p(285)(38));
FA_ff_9732:FAff port map(x=>p(232)(38),y=>p(233)(38),Cin=>p(234)(38),clock=>clock,reset=>reset,s=>p(284)(38),cout=>p(285)(39));
FA_ff_9733:FAff port map(x=>p(232)(39),y=>p(233)(39),Cin=>p(234)(39),clock=>clock,reset=>reset,s=>p(284)(39),cout=>p(285)(40));
FA_ff_9734:FAff port map(x=>p(232)(40),y=>p(233)(40),Cin=>p(234)(40),clock=>clock,reset=>reset,s=>p(284)(40),cout=>p(285)(41));
FA_ff_9735:FAff port map(x=>p(232)(41),y=>p(233)(41),Cin=>p(234)(41),clock=>clock,reset=>reset,s=>p(284)(41),cout=>p(285)(42));
FA_ff_9736:FAff port map(x=>p(232)(42),y=>p(233)(42),Cin=>p(234)(42),clock=>clock,reset=>reset,s=>p(284)(42),cout=>p(285)(43));
FA_ff_9737:FAff port map(x=>p(232)(43),y=>p(233)(43),Cin=>p(234)(43),clock=>clock,reset=>reset,s=>p(284)(43),cout=>p(285)(44));
FA_ff_9738:FAff port map(x=>p(232)(44),y=>p(233)(44),Cin=>p(234)(44),clock=>clock,reset=>reset,s=>p(284)(44),cout=>p(285)(45));
FA_ff_9739:FAff port map(x=>p(232)(45),y=>p(233)(45),Cin=>p(234)(45),clock=>clock,reset=>reset,s=>p(284)(45),cout=>p(285)(46));
FA_ff_9740:FAff port map(x=>p(232)(46),y=>p(233)(46),Cin=>p(234)(46),clock=>clock,reset=>reset,s=>p(284)(46),cout=>p(285)(47));
FA_ff_9741:FAff port map(x=>p(232)(47),y=>p(233)(47),Cin=>p(234)(47),clock=>clock,reset=>reset,s=>p(284)(47),cout=>p(285)(48));
FA_ff_9742:FAff port map(x=>p(232)(48),y=>p(233)(48),Cin=>p(234)(48),clock=>clock,reset=>reset,s=>p(284)(48),cout=>p(285)(49));
FA_ff_9743:FAff port map(x=>p(232)(49),y=>p(233)(49),Cin=>p(234)(49),clock=>clock,reset=>reset,s=>p(284)(49),cout=>p(285)(50));
FA_ff_9744:FAff port map(x=>p(232)(50),y=>p(233)(50),Cin=>p(234)(50),clock=>clock,reset=>reset,s=>p(284)(50),cout=>p(285)(51));
FA_ff_9745:FAff port map(x=>p(232)(51),y=>p(233)(51),Cin=>p(234)(51),clock=>clock,reset=>reset,s=>p(284)(51),cout=>p(285)(52));
FA_ff_9746:FAff port map(x=>p(232)(52),y=>p(233)(52),Cin=>p(234)(52),clock=>clock,reset=>reset,s=>p(284)(52),cout=>p(285)(53));
FA_ff_9747:FAff port map(x=>p(232)(53),y=>p(233)(53),Cin=>p(234)(53),clock=>clock,reset=>reset,s=>p(284)(53),cout=>p(285)(54));
FA_ff_9748:FAff port map(x=>p(232)(54),y=>p(233)(54),Cin=>p(234)(54),clock=>clock,reset=>reset,s=>p(284)(54),cout=>p(285)(55));
FA_ff_9749:FAff port map(x=>p(232)(55),y=>p(233)(55),Cin=>p(234)(55),clock=>clock,reset=>reset,s=>p(284)(55),cout=>p(285)(56));
FA_ff_9750:FAff port map(x=>p(232)(56),y=>p(233)(56),Cin=>p(234)(56),clock=>clock,reset=>reset,s=>p(284)(56),cout=>p(285)(57));
FA_ff_9751:FAff port map(x=>p(232)(57),y=>p(233)(57),Cin=>p(234)(57),clock=>clock,reset=>reset,s=>p(284)(57),cout=>p(285)(58));
FA_ff_9752:FAff port map(x=>p(232)(58),y=>p(233)(58),Cin=>p(234)(58),clock=>clock,reset=>reset,s=>p(284)(58),cout=>p(285)(59));
FA_ff_9753:FAff port map(x=>p(232)(59),y=>p(233)(59),Cin=>p(234)(59),clock=>clock,reset=>reset,s=>p(284)(59),cout=>p(285)(60));
FA_ff_9754:FAff port map(x=>p(232)(60),y=>p(233)(60),Cin=>p(234)(60),clock=>clock,reset=>reset,s=>p(284)(60),cout=>p(285)(61));
FA_ff_9755:FAff port map(x=>p(232)(61),y=>p(233)(61),Cin=>p(234)(61),clock=>clock,reset=>reset,s=>p(284)(61),cout=>p(285)(62));
FA_ff_9756:FAff port map(x=>p(232)(62),y=>p(233)(62),Cin=>p(234)(62),clock=>clock,reset=>reset,s=>p(284)(62),cout=>p(285)(63));
FA_ff_9757:FAff port map(x=>p(232)(63),y=>p(233)(63),Cin=>p(234)(63),clock=>clock,reset=>reset,s=>p(284)(63),cout=>p(285)(64));
FA_ff_9758:FAff port map(x=>p(232)(64),y=>p(233)(64),Cin=>p(234)(64),clock=>clock,reset=>reset,s=>p(284)(64),cout=>p(285)(65));
FA_ff_9759:FAff port map(x=>p(232)(65),y=>p(233)(65),Cin=>p(234)(65),clock=>clock,reset=>reset,s=>p(284)(65),cout=>p(285)(66));
FA_ff_9760:FAff port map(x=>p(232)(66),y=>p(233)(66),Cin=>p(234)(66),clock=>clock,reset=>reset,s=>p(284)(66),cout=>p(285)(67));
FA_ff_9761:FAff port map(x=>p(232)(67),y=>p(233)(67),Cin=>p(234)(67),clock=>clock,reset=>reset,s=>p(284)(67),cout=>p(285)(68));
FA_ff_9762:FAff port map(x=>p(232)(68),y=>p(233)(68),Cin=>p(234)(68),clock=>clock,reset=>reset,s=>p(284)(68),cout=>p(285)(69));
FA_ff_9763:FAff port map(x=>p(232)(69),y=>p(233)(69),Cin=>p(234)(69),clock=>clock,reset=>reset,s=>p(284)(69),cout=>p(285)(70));
FA_ff_9764:FAff port map(x=>p(232)(70),y=>p(233)(70),Cin=>p(234)(70),clock=>clock,reset=>reset,s=>p(284)(70),cout=>p(285)(71));
FA_ff_9765:FAff port map(x=>p(232)(71),y=>p(233)(71),Cin=>p(234)(71),clock=>clock,reset=>reset,s=>p(284)(71),cout=>p(285)(72));
FA_ff_9766:FAff port map(x=>p(232)(72),y=>p(233)(72),Cin=>p(234)(72),clock=>clock,reset=>reset,s=>p(284)(72),cout=>p(285)(73));
FA_ff_9767:FAff port map(x=>p(232)(73),y=>p(233)(73),Cin=>p(234)(73),clock=>clock,reset=>reset,s=>p(284)(73),cout=>p(285)(74));
FA_ff_9768:FAff port map(x=>p(232)(74),y=>p(233)(74),Cin=>p(234)(74),clock=>clock,reset=>reset,s=>p(284)(74),cout=>p(285)(75));
FA_ff_9769:FAff port map(x=>p(232)(75),y=>p(233)(75),Cin=>p(234)(75),clock=>clock,reset=>reset,s=>p(284)(75),cout=>p(285)(76));
FA_ff_9770:FAff port map(x=>p(232)(76),y=>p(233)(76),Cin=>p(234)(76),clock=>clock,reset=>reset,s=>p(284)(76),cout=>p(285)(77));
FA_ff_9771:FAff port map(x=>p(232)(77),y=>p(233)(77),Cin=>p(234)(77),clock=>clock,reset=>reset,s=>p(284)(77),cout=>p(285)(78));
FA_ff_9772:FAff port map(x=>p(232)(78),y=>p(233)(78),Cin=>p(234)(78),clock=>clock,reset=>reset,s=>p(284)(78),cout=>p(285)(79));
FA_ff_9773:FAff port map(x=>p(232)(79),y=>p(233)(79),Cin=>p(234)(79),clock=>clock,reset=>reset,s=>p(284)(79),cout=>p(285)(80));
FA_ff_9774:FAff port map(x=>p(232)(80),y=>p(233)(80),Cin=>p(234)(80),clock=>clock,reset=>reset,s=>p(284)(80),cout=>p(285)(81));
FA_ff_9775:FAff port map(x=>p(232)(81),y=>p(233)(81),Cin=>p(234)(81),clock=>clock,reset=>reset,s=>p(284)(81),cout=>p(285)(82));
FA_ff_9776:FAff port map(x=>p(232)(82),y=>p(233)(82),Cin=>p(234)(82),clock=>clock,reset=>reset,s=>p(284)(82),cout=>p(285)(83));
FA_ff_9777:FAff port map(x=>p(232)(83),y=>p(233)(83),Cin=>p(234)(83),clock=>clock,reset=>reset,s=>p(284)(83),cout=>p(285)(84));
FA_ff_9778:FAff port map(x=>p(232)(84),y=>p(233)(84),Cin=>p(234)(84),clock=>clock,reset=>reset,s=>p(284)(84),cout=>p(285)(85));
FA_ff_9779:FAff port map(x=>p(232)(85),y=>p(233)(85),Cin=>p(234)(85),clock=>clock,reset=>reset,s=>p(284)(85),cout=>p(285)(86));
FA_ff_9780:FAff port map(x=>p(232)(86),y=>p(233)(86),Cin=>p(234)(86),clock=>clock,reset=>reset,s=>p(284)(86),cout=>p(285)(87));
FA_ff_9781:FAff port map(x=>p(232)(87),y=>p(233)(87),Cin=>p(234)(87),clock=>clock,reset=>reset,s=>p(284)(87),cout=>p(285)(88));
FA_ff_9782:FAff port map(x=>p(232)(88),y=>p(233)(88),Cin=>p(234)(88),clock=>clock,reset=>reset,s=>p(284)(88),cout=>p(285)(89));
FA_ff_9783:FAff port map(x=>p(232)(89),y=>p(233)(89),Cin=>p(234)(89),clock=>clock,reset=>reset,s=>p(284)(89),cout=>p(285)(90));
FA_ff_9784:FAff port map(x=>p(232)(90),y=>p(233)(90),Cin=>p(234)(90),clock=>clock,reset=>reset,s=>p(284)(90),cout=>p(285)(91));
FA_ff_9785:FAff port map(x=>p(232)(91),y=>p(233)(91),Cin=>p(234)(91),clock=>clock,reset=>reset,s=>p(284)(91),cout=>p(285)(92));
FA_ff_9786:FAff port map(x=>p(232)(92),y=>p(233)(92),Cin=>p(234)(92),clock=>clock,reset=>reset,s=>p(284)(92),cout=>p(285)(93));
FA_ff_9787:FAff port map(x=>p(232)(93),y=>p(233)(93),Cin=>p(234)(93),clock=>clock,reset=>reset,s=>p(284)(93),cout=>p(285)(94));
FA_ff_9788:FAff port map(x=>p(232)(94),y=>p(233)(94),Cin=>p(234)(94),clock=>clock,reset=>reset,s=>p(284)(94),cout=>p(285)(95));
FA_ff_9789:FAff port map(x=>p(232)(95),y=>p(233)(95),Cin=>p(234)(95),clock=>clock,reset=>reset,s=>p(284)(95),cout=>p(285)(96));
FA_ff_9790:FAff port map(x=>p(232)(96),y=>p(233)(96),Cin=>p(234)(96),clock=>clock,reset=>reset,s=>p(284)(96),cout=>p(285)(97));
FA_ff_9791:FAff port map(x=>p(232)(97),y=>p(233)(97),Cin=>p(234)(97),clock=>clock,reset=>reset,s=>p(284)(97),cout=>p(285)(98));
FA_ff_9792:FAff port map(x=>p(232)(98),y=>p(233)(98),Cin=>p(234)(98),clock=>clock,reset=>reset,s=>p(284)(98),cout=>p(285)(99));
FA_ff_9793:FAff port map(x=>p(232)(99),y=>p(233)(99),Cin=>p(234)(99),clock=>clock,reset=>reset,s=>p(284)(99),cout=>p(285)(100));
FA_ff_9794:FAff port map(x=>p(232)(100),y=>p(233)(100),Cin=>p(234)(100),clock=>clock,reset=>reset,s=>p(284)(100),cout=>p(285)(101));
FA_ff_9795:FAff port map(x=>p(232)(101),y=>p(233)(101),Cin=>p(234)(101),clock=>clock,reset=>reset,s=>p(284)(101),cout=>p(285)(102));
FA_ff_9796:FAff port map(x=>p(232)(102),y=>p(233)(102),Cin=>p(234)(102),clock=>clock,reset=>reset,s=>p(284)(102),cout=>p(285)(103));
FA_ff_9797:FAff port map(x=>p(232)(103),y=>p(233)(103),Cin=>p(234)(103),clock=>clock,reset=>reset,s=>p(284)(103),cout=>p(285)(104));
FA_ff_9798:FAff port map(x=>p(232)(104),y=>p(233)(104),Cin=>p(234)(104),clock=>clock,reset=>reset,s=>p(284)(104),cout=>p(285)(105));
FA_ff_9799:FAff port map(x=>p(232)(105),y=>p(233)(105),Cin=>p(234)(105),clock=>clock,reset=>reset,s=>p(284)(105),cout=>p(285)(106));
FA_ff_9800:FAff port map(x=>p(232)(106),y=>p(233)(106),Cin=>p(234)(106),clock=>clock,reset=>reset,s=>p(284)(106),cout=>p(285)(107));
FA_ff_9801:FAff port map(x=>p(232)(107),y=>p(233)(107),Cin=>p(234)(107),clock=>clock,reset=>reset,s=>p(284)(107),cout=>p(285)(108));
FA_ff_9802:FAff port map(x=>p(232)(108),y=>p(233)(108),Cin=>p(234)(108),clock=>clock,reset=>reset,s=>p(284)(108),cout=>p(285)(109));
FA_ff_9803:FAff port map(x=>p(232)(109),y=>p(233)(109),Cin=>p(234)(109),clock=>clock,reset=>reset,s=>p(284)(109),cout=>p(285)(110));
FA_ff_9804:FAff port map(x=>p(232)(110),y=>p(233)(110),Cin=>p(234)(110),clock=>clock,reset=>reset,s=>p(284)(110),cout=>p(285)(111));
FA_ff_9805:FAff port map(x=>p(232)(111),y=>p(233)(111),Cin=>p(234)(111),clock=>clock,reset=>reset,s=>p(284)(111),cout=>p(285)(112));
FA_ff_9806:FAff port map(x=>p(232)(112),y=>p(233)(112),Cin=>p(234)(112),clock=>clock,reset=>reset,s=>p(284)(112),cout=>p(285)(113));
FA_ff_9807:FAff port map(x=>p(232)(113),y=>p(233)(113),Cin=>p(234)(113),clock=>clock,reset=>reset,s=>p(284)(113),cout=>p(285)(114));
FA_ff_9808:FAff port map(x=>p(232)(114),y=>p(233)(114),Cin=>p(234)(114),clock=>clock,reset=>reset,s=>p(284)(114),cout=>p(285)(115));
FA_ff_9809:FAff port map(x=>p(232)(115),y=>p(233)(115),Cin=>p(234)(115),clock=>clock,reset=>reset,s=>p(284)(115),cout=>p(285)(116));
FA_ff_9810:FAff port map(x=>p(232)(116),y=>p(233)(116),Cin=>p(234)(116),clock=>clock,reset=>reset,s=>p(284)(116),cout=>p(285)(117));
FA_ff_9811:FAff port map(x=>p(232)(117),y=>p(233)(117),Cin=>p(234)(117),clock=>clock,reset=>reset,s=>p(284)(117),cout=>p(285)(118));
FA_ff_9812:FAff port map(x=>p(232)(118),y=>p(233)(118),Cin=>p(234)(118),clock=>clock,reset=>reset,s=>p(284)(118),cout=>p(285)(119));
FA_ff_9813:FAff port map(x=>p(232)(119),y=>p(233)(119),Cin=>p(234)(119),clock=>clock,reset=>reset,s=>p(284)(119),cout=>p(285)(120));
FA_ff_9814:FAff port map(x=>p(232)(120),y=>p(233)(120),Cin=>p(234)(120),clock=>clock,reset=>reset,s=>p(284)(120),cout=>p(285)(121));
FA_ff_9815:FAff port map(x=>p(232)(121),y=>p(233)(121),Cin=>p(234)(121),clock=>clock,reset=>reset,s=>p(284)(121),cout=>p(285)(122));
FA_ff_9816:FAff port map(x=>p(232)(122),y=>p(233)(122),Cin=>p(234)(122),clock=>clock,reset=>reset,s=>p(284)(122),cout=>p(285)(123));
FA_ff_9817:FAff port map(x=>p(232)(123),y=>p(233)(123),Cin=>p(234)(123),clock=>clock,reset=>reset,s=>p(284)(123),cout=>p(285)(124));
FA_ff_9818:FAff port map(x=>p(232)(124),y=>p(233)(124),Cin=>p(234)(124),clock=>clock,reset=>reset,s=>p(284)(124),cout=>p(285)(125));
FA_ff_9819:FAff port map(x=>p(232)(125),y=>p(233)(125),Cin=>p(234)(125),clock=>clock,reset=>reset,s=>p(284)(125),cout=>p(285)(126));
FA_ff_9820:FAff port map(x=>p(232)(126),y=>p(233)(126),Cin=>p(234)(126),clock=>clock,reset=>reset,s=>p(284)(126),cout=>p(285)(127));
FA_ff_9821:FAff port map(x=>p(232)(127),y=>p(233)(127),Cin=>p(234)(127),clock=>clock,reset=>reset,s=>p(284)(127),cout=>p(285)(128));
FA_ff_9822:FAff port map(x=>p(232)(128),y=>p(233)(128),Cin=>p(234)(128),clock=>clock,reset=>reset,s=>p(284)(128),cout=>p(285)(129));
p(284)(129)<=p(233)(129);
p(286)(0)<=p(236)(0);
HA_ff_37:HAff port map(x=>p(235)(1),y=>p(236)(1),clock=>clock,reset=>reset,s=>p(286)(1),c=>p(287)(2));
FA_ff_9823:FAff port map(x=>p(235)(2),y=>p(236)(2),Cin=>p(237)(2),clock=>clock,reset=>reset,s=>p(286)(2),cout=>p(287)(3));
FA_ff_9824:FAff port map(x=>p(235)(3),y=>p(236)(3),Cin=>p(237)(3),clock=>clock,reset=>reset,s=>p(286)(3),cout=>p(287)(4));
FA_ff_9825:FAff port map(x=>p(235)(4),y=>p(236)(4),Cin=>p(237)(4),clock=>clock,reset=>reset,s=>p(286)(4),cout=>p(287)(5));
FA_ff_9826:FAff port map(x=>p(235)(5),y=>p(236)(5),Cin=>p(237)(5),clock=>clock,reset=>reset,s=>p(286)(5),cout=>p(287)(6));
FA_ff_9827:FAff port map(x=>p(235)(6),y=>p(236)(6),Cin=>p(237)(6),clock=>clock,reset=>reset,s=>p(286)(6),cout=>p(287)(7));
FA_ff_9828:FAff port map(x=>p(235)(7),y=>p(236)(7),Cin=>p(237)(7),clock=>clock,reset=>reset,s=>p(286)(7),cout=>p(287)(8));
FA_ff_9829:FAff port map(x=>p(235)(8),y=>p(236)(8),Cin=>p(237)(8),clock=>clock,reset=>reset,s=>p(286)(8),cout=>p(287)(9));
FA_ff_9830:FAff port map(x=>p(235)(9),y=>p(236)(9),Cin=>p(237)(9),clock=>clock,reset=>reset,s=>p(286)(9),cout=>p(287)(10));
FA_ff_9831:FAff port map(x=>p(235)(10),y=>p(236)(10),Cin=>p(237)(10),clock=>clock,reset=>reset,s=>p(286)(10),cout=>p(287)(11));
FA_ff_9832:FAff port map(x=>p(235)(11),y=>p(236)(11),Cin=>p(237)(11),clock=>clock,reset=>reset,s=>p(286)(11),cout=>p(287)(12));
FA_ff_9833:FAff port map(x=>p(235)(12),y=>p(236)(12),Cin=>p(237)(12),clock=>clock,reset=>reset,s=>p(286)(12),cout=>p(287)(13));
FA_ff_9834:FAff port map(x=>p(235)(13),y=>p(236)(13),Cin=>p(237)(13),clock=>clock,reset=>reset,s=>p(286)(13),cout=>p(287)(14));
FA_ff_9835:FAff port map(x=>p(235)(14),y=>p(236)(14),Cin=>p(237)(14),clock=>clock,reset=>reset,s=>p(286)(14),cout=>p(287)(15));
FA_ff_9836:FAff port map(x=>p(235)(15),y=>p(236)(15),Cin=>p(237)(15),clock=>clock,reset=>reset,s=>p(286)(15),cout=>p(287)(16));
FA_ff_9837:FAff port map(x=>p(235)(16),y=>p(236)(16),Cin=>p(237)(16),clock=>clock,reset=>reset,s=>p(286)(16),cout=>p(287)(17));
FA_ff_9838:FAff port map(x=>p(235)(17),y=>p(236)(17),Cin=>p(237)(17),clock=>clock,reset=>reset,s=>p(286)(17),cout=>p(287)(18));
FA_ff_9839:FAff port map(x=>p(235)(18),y=>p(236)(18),Cin=>p(237)(18),clock=>clock,reset=>reset,s=>p(286)(18),cout=>p(287)(19));
FA_ff_9840:FAff port map(x=>p(235)(19),y=>p(236)(19),Cin=>p(237)(19),clock=>clock,reset=>reset,s=>p(286)(19),cout=>p(287)(20));
FA_ff_9841:FAff port map(x=>p(235)(20),y=>p(236)(20),Cin=>p(237)(20),clock=>clock,reset=>reset,s=>p(286)(20),cout=>p(287)(21));
FA_ff_9842:FAff port map(x=>p(235)(21),y=>p(236)(21),Cin=>p(237)(21),clock=>clock,reset=>reset,s=>p(286)(21),cout=>p(287)(22));
FA_ff_9843:FAff port map(x=>p(235)(22),y=>p(236)(22),Cin=>p(237)(22),clock=>clock,reset=>reset,s=>p(286)(22),cout=>p(287)(23));
FA_ff_9844:FAff port map(x=>p(235)(23),y=>p(236)(23),Cin=>p(237)(23),clock=>clock,reset=>reset,s=>p(286)(23),cout=>p(287)(24));
FA_ff_9845:FAff port map(x=>p(235)(24),y=>p(236)(24),Cin=>p(237)(24),clock=>clock,reset=>reset,s=>p(286)(24),cout=>p(287)(25));
FA_ff_9846:FAff port map(x=>p(235)(25),y=>p(236)(25),Cin=>p(237)(25),clock=>clock,reset=>reset,s=>p(286)(25),cout=>p(287)(26));
FA_ff_9847:FAff port map(x=>p(235)(26),y=>p(236)(26),Cin=>p(237)(26),clock=>clock,reset=>reset,s=>p(286)(26),cout=>p(287)(27));
FA_ff_9848:FAff port map(x=>p(235)(27),y=>p(236)(27),Cin=>p(237)(27),clock=>clock,reset=>reset,s=>p(286)(27),cout=>p(287)(28));
FA_ff_9849:FAff port map(x=>p(235)(28),y=>p(236)(28),Cin=>p(237)(28),clock=>clock,reset=>reset,s=>p(286)(28),cout=>p(287)(29));
FA_ff_9850:FAff port map(x=>p(235)(29),y=>p(236)(29),Cin=>p(237)(29),clock=>clock,reset=>reset,s=>p(286)(29),cout=>p(287)(30));
FA_ff_9851:FAff port map(x=>p(235)(30),y=>p(236)(30),Cin=>p(237)(30),clock=>clock,reset=>reset,s=>p(286)(30),cout=>p(287)(31));
FA_ff_9852:FAff port map(x=>p(235)(31),y=>p(236)(31),Cin=>p(237)(31),clock=>clock,reset=>reset,s=>p(286)(31),cout=>p(287)(32));
FA_ff_9853:FAff port map(x=>p(235)(32),y=>p(236)(32),Cin=>p(237)(32),clock=>clock,reset=>reset,s=>p(286)(32),cout=>p(287)(33));
FA_ff_9854:FAff port map(x=>p(235)(33),y=>p(236)(33),Cin=>p(237)(33),clock=>clock,reset=>reset,s=>p(286)(33),cout=>p(287)(34));
FA_ff_9855:FAff port map(x=>p(235)(34),y=>p(236)(34),Cin=>p(237)(34),clock=>clock,reset=>reset,s=>p(286)(34),cout=>p(287)(35));
FA_ff_9856:FAff port map(x=>p(235)(35),y=>p(236)(35),Cin=>p(237)(35),clock=>clock,reset=>reset,s=>p(286)(35),cout=>p(287)(36));
FA_ff_9857:FAff port map(x=>p(235)(36),y=>p(236)(36),Cin=>p(237)(36),clock=>clock,reset=>reset,s=>p(286)(36),cout=>p(287)(37));
FA_ff_9858:FAff port map(x=>p(235)(37),y=>p(236)(37),Cin=>p(237)(37),clock=>clock,reset=>reset,s=>p(286)(37),cout=>p(287)(38));
FA_ff_9859:FAff port map(x=>p(235)(38),y=>p(236)(38),Cin=>p(237)(38),clock=>clock,reset=>reset,s=>p(286)(38),cout=>p(287)(39));
FA_ff_9860:FAff port map(x=>p(235)(39),y=>p(236)(39),Cin=>p(237)(39),clock=>clock,reset=>reset,s=>p(286)(39),cout=>p(287)(40));
FA_ff_9861:FAff port map(x=>p(235)(40),y=>p(236)(40),Cin=>p(237)(40),clock=>clock,reset=>reset,s=>p(286)(40),cout=>p(287)(41));
FA_ff_9862:FAff port map(x=>p(235)(41),y=>p(236)(41),Cin=>p(237)(41),clock=>clock,reset=>reset,s=>p(286)(41),cout=>p(287)(42));
FA_ff_9863:FAff port map(x=>p(235)(42),y=>p(236)(42),Cin=>p(237)(42),clock=>clock,reset=>reset,s=>p(286)(42),cout=>p(287)(43));
FA_ff_9864:FAff port map(x=>p(235)(43),y=>p(236)(43),Cin=>p(237)(43),clock=>clock,reset=>reset,s=>p(286)(43),cout=>p(287)(44));
FA_ff_9865:FAff port map(x=>p(235)(44),y=>p(236)(44),Cin=>p(237)(44),clock=>clock,reset=>reset,s=>p(286)(44),cout=>p(287)(45));
FA_ff_9866:FAff port map(x=>p(235)(45),y=>p(236)(45),Cin=>p(237)(45),clock=>clock,reset=>reset,s=>p(286)(45),cout=>p(287)(46));
FA_ff_9867:FAff port map(x=>p(235)(46),y=>p(236)(46),Cin=>p(237)(46),clock=>clock,reset=>reset,s=>p(286)(46),cout=>p(287)(47));
FA_ff_9868:FAff port map(x=>p(235)(47),y=>p(236)(47),Cin=>p(237)(47),clock=>clock,reset=>reset,s=>p(286)(47),cout=>p(287)(48));
FA_ff_9869:FAff port map(x=>p(235)(48),y=>p(236)(48),Cin=>p(237)(48),clock=>clock,reset=>reset,s=>p(286)(48),cout=>p(287)(49));
FA_ff_9870:FAff port map(x=>p(235)(49),y=>p(236)(49),Cin=>p(237)(49),clock=>clock,reset=>reset,s=>p(286)(49),cout=>p(287)(50));
FA_ff_9871:FAff port map(x=>p(235)(50),y=>p(236)(50),Cin=>p(237)(50),clock=>clock,reset=>reset,s=>p(286)(50),cout=>p(287)(51));
FA_ff_9872:FAff port map(x=>p(235)(51),y=>p(236)(51),Cin=>p(237)(51),clock=>clock,reset=>reset,s=>p(286)(51),cout=>p(287)(52));
FA_ff_9873:FAff port map(x=>p(235)(52),y=>p(236)(52),Cin=>p(237)(52),clock=>clock,reset=>reset,s=>p(286)(52),cout=>p(287)(53));
FA_ff_9874:FAff port map(x=>p(235)(53),y=>p(236)(53),Cin=>p(237)(53),clock=>clock,reset=>reset,s=>p(286)(53),cout=>p(287)(54));
FA_ff_9875:FAff port map(x=>p(235)(54),y=>p(236)(54),Cin=>p(237)(54),clock=>clock,reset=>reset,s=>p(286)(54),cout=>p(287)(55));
FA_ff_9876:FAff port map(x=>p(235)(55),y=>p(236)(55),Cin=>p(237)(55),clock=>clock,reset=>reset,s=>p(286)(55),cout=>p(287)(56));
FA_ff_9877:FAff port map(x=>p(235)(56),y=>p(236)(56),Cin=>p(237)(56),clock=>clock,reset=>reset,s=>p(286)(56),cout=>p(287)(57));
FA_ff_9878:FAff port map(x=>p(235)(57),y=>p(236)(57),Cin=>p(237)(57),clock=>clock,reset=>reset,s=>p(286)(57),cout=>p(287)(58));
FA_ff_9879:FAff port map(x=>p(235)(58),y=>p(236)(58),Cin=>p(237)(58),clock=>clock,reset=>reset,s=>p(286)(58),cout=>p(287)(59));
FA_ff_9880:FAff port map(x=>p(235)(59),y=>p(236)(59),Cin=>p(237)(59),clock=>clock,reset=>reset,s=>p(286)(59),cout=>p(287)(60));
FA_ff_9881:FAff port map(x=>p(235)(60),y=>p(236)(60),Cin=>p(237)(60),clock=>clock,reset=>reset,s=>p(286)(60),cout=>p(287)(61));
FA_ff_9882:FAff port map(x=>p(235)(61),y=>p(236)(61),Cin=>p(237)(61),clock=>clock,reset=>reset,s=>p(286)(61),cout=>p(287)(62));
FA_ff_9883:FAff port map(x=>p(235)(62),y=>p(236)(62),Cin=>p(237)(62),clock=>clock,reset=>reset,s=>p(286)(62),cout=>p(287)(63));
FA_ff_9884:FAff port map(x=>p(235)(63),y=>p(236)(63),Cin=>p(237)(63),clock=>clock,reset=>reset,s=>p(286)(63),cout=>p(287)(64));
FA_ff_9885:FAff port map(x=>p(235)(64),y=>p(236)(64),Cin=>p(237)(64),clock=>clock,reset=>reset,s=>p(286)(64),cout=>p(287)(65));
FA_ff_9886:FAff port map(x=>p(235)(65),y=>p(236)(65),Cin=>p(237)(65),clock=>clock,reset=>reset,s=>p(286)(65),cout=>p(287)(66));
FA_ff_9887:FAff port map(x=>p(235)(66),y=>p(236)(66),Cin=>p(237)(66),clock=>clock,reset=>reset,s=>p(286)(66),cout=>p(287)(67));
FA_ff_9888:FAff port map(x=>p(235)(67),y=>p(236)(67),Cin=>p(237)(67),clock=>clock,reset=>reset,s=>p(286)(67),cout=>p(287)(68));
FA_ff_9889:FAff port map(x=>p(235)(68),y=>p(236)(68),Cin=>p(237)(68),clock=>clock,reset=>reset,s=>p(286)(68),cout=>p(287)(69));
FA_ff_9890:FAff port map(x=>p(235)(69),y=>p(236)(69),Cin=>p(237)(69),clock=>clock,reset=>reset,s=>p(286)(69),cout=>p(287)(70));
FA_ff_9891:FAff port map(x=>p(235)(70),y=>p(236)(70),Cin=>p(237)(70),clock=>clock,reset=>reset,s=>p(286)(70),cout=>p(287)(71));
FA_ff_9892:FAff port map(x=>p(235)(71),y=>p(236)(71),Cin=>p(237)(71),clock=>clock,reset=>reset,s=>p(286)(71),cout=>p(287)(72));
FA_ff_9893:FAff port map(x=>p(235)(72),y=>p(236)(72),Cin=>p(237)(72),clock=>clock,reset=>reset,s=>p(286)(72),cout=>p(287)(73));
FA_ff_9894:FAff port map(x=>p(235)(73),y=>p(236)(73),Cin=>p(237)(73),clock=>clock,reset=>reset,s=>p(286)(73),cout=>p(287)(74));
FA_ff_9895:FAff port map(x=>p(235)(74),y=>p(236)(74),Cin=>p(237)(74),clock=>clock,reset=>reset,s=>p(286)(74),cout=>p(287)(75));
FA_ff_9896:FAff port map(x=>p(235)(75),y=>p(236)(75),Cin=>p(237)(75),clock=>clock,reset=>reset,s=>p(286)(75),cout=>p(287)(76));
FA_ff_9897:FAff port map(x=>p(235)(76),y=>p(236)(76),Cin=>p(237)(76),clock=>clock,reset=>reset,s=>p(286)(76),cout=>p(287)(77));
FA_ff_9898:FAff port map(x=>p(235)(77),y=>p(236)(77),Cin=>p(237)(77),clock=>clock,reset=>reset,s=>p(286)(77),cout=>p(287)(78));
FA_ff_9899:FAff port map(x=>p(235)(78),y=>p(236)(78),Cin=>p(237)(78),clock=>clock,reset=>reset,s=>p(286)(78),cout=>p(287)(79));
FA_ff_9900:FAff port map(x=>p(235)(79),y=>p(236)(79),Cin=>p(237)(79),clock=>clock,reset=>reset,s=>p(286)(79),cout=>p(287)(80));
FA_ff_9901:FAff port map(x=>p(235)(80),y=>p(236)(80),Cin=>p(237)(80),clock=>clock,reset=>reset,s=>p(286)(80),cout=>p(287)(81));
FA_ff_9902:FAff port map(x=>p(235)(81),y=>p(236)(81),Cin=>p(237)(81),clock=>clock,reset=>reset,s=>p(286)(81),cout=>p(287)(82));
FA_ff_9903:FAff port map(x=>p(235)(82),y=>p(236)(82),Cin=>p(237)(82),clock=>clock,reset=>reset,s=>p(286)(82),cout=>p(287)(83));
FA_ff_9904:FAff port map(x=>p(235)(83),y=>p(236)(83),Cin=>p(237)(83),clock=>clock,reset=>reset,s=>p(286)(83),cout=>p(287)(84));
FA_ff_9905:FAff port map(x=>p(235)(84),y=>p(236)(84),Cin=>p(237)(84),clock=>clock,reset=>reset,s=>p(286)(84),cout=>p(287)(85));
FA_ff_9906:FAff port map(x=>p(235)(85),y=>p(236)(85),Cin=>p(237)(85),clock=>clock,reset=>reset,s=>p(286)(85),cout=>p(287)(86));
FA_ff_9907:FAff port map(x=>p(235)(86),y=>p(236)(86),Cin=>p(237)(86),clock=>clock,reset=>reset,s=>p(286)(86),cout=>p(287)(87));
FA_ff_9908:FAff port map(x=>p(235)(87),y=>p(236)(87),Cin=>p(237)(87),clock=>clock,reset=>reset,s=>p(286)(87),cout=>p(287)(88));
FA_ff_9909:FAff port map(x=>p(235)(88),y=>p(236)(88),Cin=>p(237)(88),clock=>clock,reset=>reset,s=>p(286)(88),cout=>p(287)(89));
FA_ff_9910:FAff port map(x=>p(235)(89),y=>p(236)(89),Cin=>p(237)(89),clock=>clock,reset=>reset,s=>p(286)(89),cout=>p(287)(90));
FA_ff_9911:FAff port map(x=>p(235)(90),y=>p(236)(90),Cin=>p(237)(90),clock=>clock,reset=>reset,s=>p(286)(90),cout=>p(287)(91));
FA_ff_9912:FAff port map(x=>p(235)(91),y=>p(236)(91),Cin=>p(237)(91),clock=>clock,reset=>reset,s=>p(286)(91),cout=>p(287)(92));
FA_ff_9913:FAff port map(x=>p(235)(92),y=>p(236)(92),Cin=>p(237)(92),clock=>clock,reset=>reset,s=>p(286)(92),cout=>p(287)(93));
FA_ff_9914:FAff port map(x=>p(235)(93),y=>p(236)(93),Cin=>p(237)(93),clock=>clock,reset=>reset,s=>p(286)(93),cout=>p(287)(94));
FA_ff_9915:FAff port map(x=>p(235)(94),y=>p(236)(94),Cin=>p(237)(94),clock=>clock,reset=>reset,s=>p(286)(94),cout=>p(287)(95));
FA_ff_9916:FAff port map(x=>p(235)(95),y=>p(236)(95),Cin=>p(237)(95),clock=>clock,reset=>reset,s=>p(286)(95),cout=>p(287)(96));
FA_ff_9917:FAff port map(x=>p(235)(96),y=>p(236)(96),Cin=>p(237)(96),clock=>clock,reset=>reset,s=>p(286)(96),cout=>p(287)(97));
FA_ff_9918:FAff port map(x=>p(235)(97),y=>p(236)(97),Cin=>p(237)(97),clock=>clock,reset=>reset,s=>p(286)(97),cout=>p(287)(98));
FA_ff_9919:FAff port map(x=>p(235)(98),y=>p(236)(98),Cin=>p(237)(98),clock=>clock,reset=>reset,s=>p(286)(98),cout=>p(287)(99));
FA_ff_9920:FAff port map(x=>p(235)(99),y=>p(236)(99),Cin=>p(237)(99),clock=>clock,reset=>reset,s=>p(286)(99),cout=>p(287)(100));
FA_ff_9921:FAff port map(x=>p(235)(100),y=>p(236)(100),Cin=>p(237)(100),clock=>clock,reset=>reset,s=>p(286)(100),cout=>p(287)(101));
FA_ff_9922:FAff port map(x=>p(235)(101),y=>p(236)(101),Cin=>p(237)(101),clock=>clock,reset=>reset,s=>p(286)(101),cout=>p(287)(102));
FA_ff_9923:FAff port map(x=>p(235)(102),y=>p(236)(102),Cin=>p(237)(102),clock=>clock,reset=>reset,s=>p(286)(102),cout=>p(287)(103));
FA_ff_9924:FAff port map(x=>p(235)(103),y=>p(236)(103),Cin=>p(237)(103),clock=>clock,reset=>reset,s=>p(286)(103),cout=>p(287)(104));
FA_ff_9925:FAff port map(x=>p(235)(104),y=>p(236)(104),Cin=>p(237)(104),clock=>clock,reset=>reset,s=>p(286)(104),cout=>p(287)(105));
FA_ff_9926:FAff port map(x=>p(235)(105),y=>p(236)(105),Cin=>p(237)(105),clock=>clock,reset=>reset,s=>p(286)(105),cout=>p(287)(106));
FA_ff_9927:FAff port map(x=>p(235)(106),y=>p(236)(106),Cin=>p(237)(106),clock=>clock,reset=>reset,s=>p(286)(106),cout=>p(287)(107));
FA_ff_9928:FAff port map(x=>p(235)(107),y=>p(236)(107),Cin=>p(237)(107),clock=>clock,reset=>reset,s=>p(286)(107),cout=>p(287)(108));
FA_ff_9929:FAff port map(x=>p(235)(108),y=>p(236)(108),Cin=>p(237)(108),clock=>clock,reset=>reset,s=>p(286)(108),cout=>p(287)(109));
FA_ff_9930:FAff port map(x=>p(235)(109),y=>p(236)(109),Cin=>p(237)(109),clock=>clock,reset=>reset,s=>p(286)(109),cout=>p(287)(110));
FA_ff_9931:FAff port map(x=>p(235)(110),y=>p(236)(110),Cin=>p(237)(110),clock=>clock,reset=>reset,s=>p(286)(110),cout=>p(287)(111));
FA_ff_9932:FAff port map(x=>p(235)(111),y=>p(236)(111),Cin=>p(237)(111),clock=>clock,reset=>reset,s=>p(286)(111),cout=>p(287)(112));
FA_ff_9933:FAff port map(x=>p(235)(112),y=>p(236)(112),Cin=>p(237)(112),clock=>clock,reset=>reset,s=>p(286)(112),cout=>p(287)(113));
FA_ff_9934:FAff port map(x=>p(235)(113),y=>p(236)(113),Cin=>p(237)(113),clock=>clock,reset=>reset,s=>p(286)(113),cout=>p(287)(114));
FA_ff_9935:FAff port map(x=>p(235)(114),y=>p(236)(114),Cin=>p(237)(114),clock=>clock,reset=>reset,s=>p(286)(114),cout=>p(287)(115));
FA_ff_9936:FAff port map(x=>p(235)(115),y=>p(236)(115),Cin=>p(237)(115),clock=>clock,reset=>reset,s=>p(286)(115),cout=>p(287)(116));
FA_ff_9937:FAff port map(x=>p(235)(116),y=>p(236)(116),Cin=>p(237)(116),clock=>clock,reset=>reset,s=>p(286)(116),cout=>p(287)(117));
FA_ff_9938:FAff port map(x=>p(235)(117),y=>p(236)(117),Cin=>p(237)(117),clock=>clock,reset=>reset,s=>p(286)(117),cout=>p(287)(118));
FA_ff_9939:FAff port map(x=>p(235)(118),y=>p(236)(118),Cin=>p(237)(118),clock=>clock,reset=>reset,s=>p(286)(118),cout=>p(287)(119));
FA_ff_9940:FAff port map(x=>p(235)(119),y=>p(236)(119),Cin=>p(237)(119),clock=>clock,reset=>reset,s=>p(286)(119),cout=>p(287)(120));
FA_ff_9941:FAff port map(x=>p(235)(120),y=>p(236)(120),Cin=>p(237)(120),clock=>clock,reset=>reset,s=>p(286)(120),cout=>p(287)(121));
FA_ff_9942:FAff port map(x=>p(235)(121),y=>p(236)(121),Cin=>p(237)(121),clock=>clock,reset=>reset,s=>p(286)(121),cout=>p(287)(122));
FA_ff_9943:FAff port map(x=>p(235)(122),y=>p(236)(122),Cin=>p(237)(122),clock=>clock,reset=>reset,s=>p(286)(122),cout=>p(287)(123));
FA_ff_9944:FAff port map(x=>p(235)(123),y=>p(236)(123),Cin=>p(237)(123),clock=>clock,reset=>reset,s=>p(286)(123),cout=>p(287)(124));
FA_ff_9945:FAff port map(x=>p(235)(124),y=>p(236)(124),Cin=>p(237)(124),clock=>clock,reset=>reset,s=>p(286)(124),cout=>p(287)(125));
FA_ff_9946:FAff port map(x=>p(235)(125),y=>p(236)(125),Cin=>p(237)(125),clock=>clock,reset=>reset,s=>p(286)(125),cout=>p(287)(126));
FA_ff_9947:FAff port map(x=>p(235)(126),y=>p(236)(126),Cin=>p(237)(126),clock=>clock,reset=>reset,s=>p(286)(126),cout=>p(287)(127));
FA_ff_9948:FAff port map(x=>p(235)(127),y=>p(236)(127),Cin=>p(237)(127),clock=>clock,reset=>reset,s=>p(286)(127),cout=>p(287)(128));
FA_ff_9949:FAff port map(x=>p(235)(128),y=>p(236)(128),Cin=>p(237)(128),clock=>clock,reset=>reset,s=>p(286)(128),cout=>p(287)(129));
p(286)(129)<=p(237)(129);
HA_ff_38:HAff port map(x=>p(238)(0),y=>p(240)(0),clock=>clock,reset=>reset,s=>p(288)(0),c=>p(289)(1));
FA_ff_9950:FAff port map(x=>p(238)(1),y=>p(239)(1),Cin=>p(240)(1),clock=>clock,reset=>reset,s=>p(288)(1),cout=>p(289)(2));
FA_ff_9951:FAff port map(x=>p(238)(2),y=>p(239)(2),Cin=>p(240)(2),clock=>clock,reset=>reset,s=>p(288)(2),cout=>p(289)(3));
FA_ff_9952:FAff port map(x=>p(238)(3),y=>p(239)(3),Cin=>p(240)(3),clock=>clock,reset=>reset,s=>p(288)(3),cout=>p(289)(4));
FA_ff_9953:FAff port map(x=>p(238)(4),y=>p(239)(4),Cin=>p(240)(4),clock=>clock,reset=>reset,s=>p(288)(4),cout=>p(289)(5));
FA_ff_9954:FAff port map(x=>p(238)(5),y=>p(239)(5),Cin=>p(240)(5),clock=>clock,reset=>reset,s=>p(288)(5),cout=>p(289)(6));
FA_ff_9955:FAff port map(x=>p(238)(6),y=>p(239)(6),Cin=>p(240)(6),clock=>clock,reset=>reset,s=>p(288)(6),cout=>p(289)(7));
FA_ff_9956:FAff port map(x=>p(238)(7),y=>p(239)(7),Cin=>p(240)(7),clock=>clock,reset=>reset,s=>p(288)(7),cout=>p(289)(8));
FA_ff_9957:FAff port map(x=>p(238)(8),y=>p(239)(8),Cin=>p(240)(8),clock=>clock,reset=>reset,s=>p(288)(8),cout=>p(289)(9));
FA_ff_9958:FAff port map(x=>p(238)(9),y=>p(239)(9),Cin=>p(240)(9),clock=>clock,reset=>reset,s=>p(288)(9),cout=>p(289)(10));
FA_ff_9959:FAff port map(x=>p(238)(10),y=>p(239)(10),Cin=>p(240)(10),clock=>clock,reset=>reset,s=>p(288)(10),cout=>p(289)(11));
FA_ff_9960:FAff port map(x=>p(238)(11),y=>p(239)(11),Cin=>p(240)(11),clock=>clock,reset=>reset,s=>p(288)(11),cout=>p(289)(12));
FA_ff_9961:FAff port map(x=>p(238)(12),y=>p(239)(12),Cin=>p(240)(12),clock=>clock,reset=>reset,s=>p(288)(12),cout=>p(289)(13));
FA_ff_9962:FAff port map(x=>p(238)(13),y=>p(239)(13),Cin=>p(240)(13),clock=>clock,reset=>reset,s=>p(288)(13),cout=>p(289)(14));
FA_ff_9963:FAff port map(x=>p(238)(14),y=>p(239)(14),Cin=>p(240)(14),clock=>clock,reset=>reset,s=>p(288)(14),cout=>p(289)(15));
FA_ff_9964:FAff port map(x=>p(238)(15),y=>p(239)(15),Cin=>p(240)(15),clock=>clock,reset=>reset,s=>p(288)(15),cout=>p(289)(16));
FA_ff_9965:FAff port map(x=>p(238)(16),y=>p(239)(16),Cin=>p(240)(16),clock=>clock,reset=>reset,s=>p(288)(16),cout=>p(289)(17));
FA_ff_9966:FAff port map(x=>p(238)(17),y=>p(239)(17),Cin=>p(240)(17),clock=>clock,reset=>reset,s=>p(288)(17),cout=>p(289)(18));
FA_ff_9967:FAff port map(x=>p(238)(18),y=>p(239)(18),Cin=>p(240)(18),clock=>clock,reset=>reset,s=>p(288)(18),cout=>p(289)(19));
FA_ff_9968:FAff port map(x=>p(238)(19),y=>p(239)(19),Cin=>p(240)(19),clock=>clock,reset=>reset,s=>p(288)(19),cout=>p(289)(20));
FA_ff_9969:FAff port map(x=>p(238)(20),y=>p(239)(20),Cin=>p(240)(20),clock=>clock,reset=>reset,s=>p(288)(20),cout=>p(289)(21));
FA_ff_9970:FAff port map(x=>p(238)(21),y=>p(239)(21),Cin=>p(240)(21),clock=>clock,reset=>reset,s=>p(288)(21),cout=>p(289)(22));
FA_ff_9971:FAff port map(x=>p(238)(22),y=>p(239)(22),Cin=>p(240)(22),clock=>clock,reset=>reset,s=>p(288)(22),cout=>p(289)(23));
FA_ff_9972:FAff port map(x=>p(238)(23),y=>p(239)(23),Cin=>p(240)(23),clock=>clock,reset=>reset,s=>p(288)(23),cout=>p(289)(24));
FA_ff_9973:FAff port map(x=>p(238)(24),y=>p(239)(24),Cin=>p(240)(24),clock=>clock,reset=>reset,s=>p(288)(24),cout=>p(289)(25));
FA_ff_9974:FAff port map(x=>p(238)(25),y=>p(239)(25),Cin=>p(240)(25),clock=>clock,reset=>reset,s=>p(288)(25),cout=>p(289)(26));
FA_ff_9975:FAff port map(x=>p(238)(26),y=>p(239)(26),Cin=>p(240)(26),clock=>clock,reset=>reset,s=>p(288)(26),cout=>p(289)(27));
FA_ff_9976:FAff port map(x=>p(238)(27),y=>p(239)(27),Cin=>p(240)(27),clock=>clock,reset=>reset,s=>p(288)(27),cout=>p(289)(28));
FA_ff_9977:FAff port map(x=>p(238)(28),y=>p(239)(28),Cin=>p(240)(28),clock=>clock,reset=>reset,s=>p(288)(28),cout=>p(289)(29));
FA_ff_9978:FAff port map(x=>p(238)(29),y=>p(239)(29),Cin=>p(240)(29),clock=>clock,reset=>reset,s=>p(288)(29),cout=>p(289)(30));
FA_ff_9979:FAff port map(x=>p(238)(30),y=>p(239)(30),Cin=>p(240)(30),clock=>clock,reset=>reset,s=>p(288)(30),cout=>p(289)(31));
FA_ff_9980:FAff port map(x=>p(238)(31),y=>p(239)(31),Cin=>p(240)(31),clock=>clock,reset=>reset,s=>p(288)(31),cout=>p(289)(32));
FA_ff_9981:FAff port map(x=>p(238)(32),y=>p(239)(32),Cin=>p(240)(32),clock=>clock,reset=>reset,s=>p(288)(32),cout=>p(289)(33));
FA_ff_9982:FAff port map(x=>p(238)(33),y=>p(239)(33),Cin=>p(240)(33),clock=>clock,reset=>reset,s=>p(288)(33),cout=>p(289)(34));
FA_ff_9983:FAff port map(x=>p(238)(34),y=>p(239)(34),Cin=>p(240)(34),clock=>clock,reset=>reset,s=>p(288)(34),cout=>p(289)(35));
FA_ff_9984:FAff port map(x=>p(238)(35),y=>p(239)(35),Cin=>p(240)(35),clock=>clock,reset=>reset,s=>p(288)(35),cout=>p(289)(36));
FA_ff_9985:FAff port map(x=>p(238)(36),y=>p(239)(36),Cin=>p(240)(36),clock=>clock,reset=>reset,s=>p(288)(36),cout=>p(289)(37));
FA_ff_9986:FAff port map(x=>p(238)(37),y=>p(239)(37),Cin=>p(240)(37),clock=>clock,reset=>reset,s=>p(288)(37),cout=>p(289)(38));
FA_ff_9987:FAff port map(x=>p(238)(38),y=>p(239)(38),Cin=>p(240)(38),clock=>clock,reset=>reset,s=>p(288)(38),cout=>p(289)(39));
FA_ff_9988:FAff port map(x=>p(238)(39),y=>p(239)(39),Cin=>p(240)(39),clock=>clock,reset=>reset,s=>p(288)(39),cout=>p(289)(40));
FA_ff_9989:FAff port map(x=>p(238)(40),y=>p(239)(40),Cin=>p(240)(40),clock=>clock,reset=>reset,s=>p(288)(40),cout=>p(289)(41));
FA_ff_9990:FAff port map(x=>p(238)(41),y=>p(239)(41),Cin=>p(240)(41),clock=>clock,reset=>reset,s=>p(288)(41),cout=>p(289)(42));
FA_ff_9991:FAff port map(x=>p(238)(42),y=>p(239)(42),Cin=>p(240)(42),clock=>clock,reset=>reset,s=>p(288)(42),cout=>p(289)(43));
FA_ff_9992:FAff port map(x=>p(238)(43),y=>p(239)(43),Cin=>p(240)(43),clock=>clock,reset=>reset,s=>p(288)(43),cout=>p(289)(44));
FA_ff_9993:FAff port map(x=>p(238)(44),y=>p(239)(44),Cin=>p(240)(44),clock=>clock,reset=>reset,s=>p(288)(44),cout=>p(289)(45));
FA_ff_9994:FAff port map(x=>p(238)(45),y=>p(239)(45),Cin=>p(240)(45),clock=>clock,reset=>reset,s=>p(288)(45),cout=>p(289)(46));
FA_ff_9995:FAff port map(x=>p(238)(46),y=>p(239)(46),Cin=>p(240)(46),clock=>clock,reset=>reset,s=>p(288)(46),cout=>p(289)(47));
FA_ff_9996:FAff port map(x=>p(238)(47),y=>p(239)(47),Cin=>p(240)(47),clock=>clock,reset=>reset,s=>p(288)(47),cout=>p(289)(48));
FA_ff_9997:FAff port map(x=>p(238)(48),y=>p(239)(48),Cin=>p(240)(48),clock=>clock,reset=>reset,s=>p(288)(48),cout=>p(289)(49));
FA_ff_9998:FAff port map(x=>p(238)(49),y=>p(239)(49),Cin=>p(240)(49),clock=>clock,reset=>reset,s=>p(288)(49),cout=>p(289)(50));
FA_ff_9999:FAff port map(x=>p(238)(50),y=>p(239)(50),Cin=>p(240)(50),clock=>clock,reset=>reset,s=>p(288)(50),cout=>p(289)(51));
FA_ff_10000:FAff port map(x=>p(238)(51),y=>p(239)(51),Cin=>p(240)(51),clock=>clock,reset=>reset,s=>p(288)(51),cout=>p(289)(52));
FA_ff_10001:FAff port map(x=>p(238)(52),y=>p(239)(52),Cin=>p(240)(52),clock=>clock,reset=>reset,s=>p(288)(52),cout=>p(289)(53));
FA_ff_10002:FAff port map(x=>p(238)(53),y=>p(239)(53),Cin=>p(240)(53),clock=>clock,reset=>reset,s=>p(288)(53),cout=>p(289)(54));
FA_ff_10003:FAff port map(x=>p(238)(54),y=>p(239)(54),Cin=>p(240)(54),clock=>clock,reset=>reset,s=>p(288)(54),cout=>p(289)(55));
FA_ff_10004:FAff port map(x=>p(238)(55),y=>p(239)(55),Cin=>p(240)(55),clock=>clock,reset=>reset,s=>p(288)(55),cout=>p(289)(56));
FA_ff_10005:FAff port map(x=>p(238)(56),y=>p(239)(56),Cin=>p(240)(56),clock=>clock,reset=>reset,s=>p(288)(56),cout=>p(289)(57));
FA_ff_10006:FAff port map(x=>p(238)(57),y=>p(239)(57),Cin=>p(240)(57),clock=>clock,reset=>reset,s=>p(288)(57),cout=>p(289)(58));
FA_ff_10007:FAff port map(x=>p(238)(58),y=>p(239)(58),Cin=>p(240)(58),clock=>clock,reset=>reset,s=>p(288)(58),cout=>p(289)(59));
FA_ff_10008:FAff port map(x=>p(238)(59),y=>p(239)(59),Cin=>p(240)(59),clock=>clock,reset=>reset,s=>p(288)(59),cout=>p(289)(60));
FA_ff_10009:FAff port map(x=>p(238)(60),y=>p(239)(60),Cin=>p(240)(60),clock=>clock,reset=>reset,s=>p(288)(60),cout=>p(289)(61));
FA_ff_10010:FAff port map(x=>p(238)(61),y=>p(239)(61),Cin=>p(240)(61),clock=>clock,reset=>reset,s=>p(288)(61),cout=>p(289)(62));
FA_ff_10011:FAff port map(x=>p(238)(62),y=>p(239)(62),Cin=>p(240)(62),clock=>clock,reset=>reset,s=>p(288)(62),cout=>p(289)(63));
FA_ff_10012:FAff port map(x=>p(238)(63),y=>p(239)(63),Cin=>p(240)(63),clock=>clock,reset=>reset,s=>p(288)(63),cout=>p(289)(64));
FA_ff_10013:FAff port map(x=>p(238)(64),y=>p(239)(64),Cin=>p(240)(64),clock=>clock,reset=>reset,s=>p(288)(64),cout=>p(289)(65));
FA_ff_10014:FAff port map(x=>p(238)(65),y=>p(239)(65),Cin=>p(240)(65),clock=>clock,reset=>reset,s=>p(288)(65),cout=>p(289)(66));
FA_ff_10015:FAff port map(x=>p(238)(66),y=>p(239)(66),Cin=>p(240)(66),clock=>clock,reset=>reset,s=>p(288)(66),cout=>p(289)(67));
FA_ff_10016:FAff port map(x=>p(238)(67),y=>p(239)(67),Cin=>p(240)(67),clock=>clock,reset=>reset,s=>p(288)(67),cout=>p(289)(68));
FA_ff_10017:FAff port map(x=>p(238)(68),y=>p(239)(68),Cin=>p(240)(68),clock=>clock,reset=>reset,s=>p(288)(68),cout=>p(289)(69));
FA_ff_10018:FAff port map(x=>p(238)(69),y=>p(239)(69),Cin=>p(240)(69),clock=>clock,reset=>reset,s=>p(288)(69),cout=>p(289)(70));
FA_ff_10019:FAff port map(x=>p(238)(70),y=>p(239)(70),Cin=>p(240)(70),clock=>clock,reset=>reset,s=>p(288)(70),cout=>p(289)(71));
FA_ff_10020:FAff port map(x=>p(238)(71),y=>p(239)(71),Cin=>p(240)(71),clock=>clock,reset=>reset,s=>p(288)(71),cout=>p(289)(72));
FA_ff_10021:FAff port map(x=>p(238)(72),y=>p(239)(72),Cin=>p(240)(72),clock=>clock,reset=>reset,s=>p(288)(72),cout=>p(289)(73));
FA_ff_10022:FAff port map(x=>p(238)(73),y=>p(239)(73),Cin=>p(240)(73),clock=>clock,reset=>reset,s=>p(288)(73),cout=>p(289)(74));
FA_ff_10023:FAff port map(x=>p(238)(74),y=>p(239)(74),Cin=>p(240)(74),clock=>clock,reset=>reset,s=>p(288)(74),cout=>p(289)(75));
FA_ff_10024:FAff port map(x=>p(238)(75),y=>p(239)(75),Cin=>p(240)(75),clock=>clock,reset=>reset,s=>p(288)(75),cout=>p(289)(76));
FA_ff_10025:FAff port map(x=>p(238)(76),y=>p(239)(76),Cin=>p(240)(76),clock=>clock,reset=>reset,s=>p(288)(76),cout=>p(289)(77));
FA_ff_10026:FAff port map(x=>p(238)(77),y=>p(239)(77),Cin=>p(240)(77),clock=>clock,reset=>reset,s=>p(288)(77),cout=>p(289)(78));
FA_ff_10027:FAff port map(x=>p(238)(78),y=>p(239)(78),Cin=>p(240)(78),clock=>clock,reset=>reset,s=>p(288)(78),cout=>p(289)(79));
FA_ff_10028:FAff port map(x=>p(238)(79),y=>p(239)(79),Cin=>p(240)(79),clock=>clock,reset=>reset,s=>p(288)(79),cout=>p(289)(80));
FA_ff_10029:FAff port map(x=>p(238)(80),y=>p(239)(80),Cin=>p(240)(80),clock=>clock,reset=>reset,s=>p(288)(80),cout=>p(289)(81));
FA_ff_10030:FAff port map(x=>p(238)(81),y=>p(239)(81),Cin=>p(240)(81),clock=>clock,reset=>reset,s=>p(288)(81),cout=>p(289)(82));
FA_ff_10031:FAff port map(x=>p(238)(82),y=>p(239)(82),Cin=>p(240)(82),clock=>clock,reset=>reset,s=>p(288)(82),cout=>p(289)(83));
FA_ff_10032:FAff port map(x=>p(238)(83),y=>p(239)(83),Cin=>p(240)(83),clock=>clock,reset=>reset,s=>p(288)(83),cout=>p(289)(84));
FA_ff_10033:FAff port map(x=>p(238)(84),y=>p(239)(84),Cin=>p(240)(84),clock=>clock,reset=>reset,s=>p(288)(84),cout=>p(289)(85));
FA_ff_10034:FAff port map(x=>p(238)(85),y=>p(239)(85),Cin=>p(240)(85),clock=>clock,reset=>reset,s=>p(288)(85),cout=>p(289)(86));
FA_ff_10035:FAff port map(x=>p(238)(86),y=>p(239)(86),Cin=>p(240)(86),clock=>clock,reset=>reset,s=>p(288)(86),cout=>p(289)(87));
FA_ff_10036:FAff port map(x=>p(238)(87),y=>p(239)(87),Cin=>p(240)(87),clock=>clock,reset=>reset,s=>p(288)(87),cout=>p(289)(88));
FA_ff_10037:FAff port map(x=>p(238)(88),y=>p(239)(88),Cin=>p(240)(88),clock=>clock,reset=>reset,s=>p(288)(88),cout=>p(289)(89));
FA_ff_10038:FAff port map(x=>p(238)(89),y=>p(239)(89),Cin=>p(240)(89),clock=>clock,reset=>reset,s=>p(288)(89),cout=>p(289)(90));
FA_ff_10039:FAff port map(x=>p(238)(90),y=>p(239)(90),Cin=>p(240)(90),clock=>clock,reset=>reset,s=>p(288)(90),cout=>p(289)(91));
FA_ff_10040:FAff port map(x=>p(238)(91),y=>p(239)(91),Cin=>p(240)(91),clock=>clock,reset=>reset,s=>p(288)(91),cout=>p(289)(92));
FA_ff_10041:FAff port map(x=>p(238)(92),y=>p(239)(92),Cin=>p(240)(92),clock=>clock,reset=>reset,s=>p(288)(92),cout=>p(289)(93));
FA_ff_10042:FAff port map(x=>p(238)(93),y=>p(239)(93),Cin=>p(240)(93),clock=>clock,reset=>reset,s=>p(288)(93),cout=>p(289)(94));
FA_ff_10043:FAff port map(x=>p(238)(94),y=>p(239)(94),Cin=>p(240)(94),clock=>clock,reset=>reset,s=>p(288)(94),cout=>p(289)(95));
FA_ff_10044:FAff port map(x=>p(238)(95),y=>p(239)(95),Cin=>p(240)(95),clock=>clock,reset=>reset,s=>p(288)(95),cout=>p(289)(96));
FA_ff_10045:FAff port map(x=>p(238)(96),y=>p(239)(96),Cin=>p(240)(96),clock=>clock,reset=>reset,s=>p(288)(96),cout=>p(289)(97));
FA_ff_10046:FAff port map(x=>p(238)(97),y=>p(239)(97),Cin=>p(240)(97),clock=>clock,reset=>reset,s=>p(288)(97),cout=>p(289)(98));
FA_ff_10047:FAff port map(x=>p(238)(98),y=>p(239)(98),Cin=>p(240)(98),clock=>clock,reset=>reset,s=>p(288)(98),cout=>p(289)(99));
FA_ff_10048:FAff port map(x=>p(238)(99),y=>p(239)(99),Cin=>p(240)(99),clock=>clock,reset=>reset,s=>p(288)(99),cout=>p(289)(100));
FA_ff_10049:FAff port map(x=>p(238)(100),y=>p(239)(100),Cin=>p(240)(100),clock=>clock,reset=>reset,s=>p(288)(100),cout=>p(289)(101));
FA_ff_10050:FAff port map(x=>p(238)(101),y=>p(239)(101),Cin=>p(240)(101),clock=>clock,reset=>reset,s=>p(288)(101),cout=>p(289)(102));
FA_ff_10051:FAff port map(x=>p(238)(102),y=>p(239)(102),Cin=>p(240)(102),clock=>clock,reset=>reset,s=>p(288)(102),cout=>p(289)(103));
FA_ff_10052:FAff port map(x=>p(238)(103),y=>p(239)(103),Cin=>p(240)(103),clock=>clock,reset=>reset,s=>p(288)(103),cout=>p(289)(104));
FA_ff_10053:FAff port map(x=>p(238)(104),y=>p(239)(104),Cin=>p(240)(104),clock=>clock,reset=>reset,s=>p(288)(104),cout=>p(289)(105));
FA_ff_10054:FAff port map(x=>p(238)(105),y=>p(239)(105),Cin=>p(240)(105),clock=>clock,reset=>reset,s=>p(288)(105),cout=>p(289)(106));
FA_ff_10055:FAff port map(x=>p(238)(106),y=>p(239)(106),Cin=>p(240)(106),clock=>clock,reset=>reset,s=>p(288)(106),cout=>p(289)(107));
FA_ff_10056:FAff port map(x=>p(238)(107),y=>p(239)(107),Cin=>p(240)(107),clock=>clock,reset=>reset,s=>p(288)(107),cout=>p(289)(108));
FA_ff_10057:FAff port map(x=>p(238)(108),y=>p(239)(108),Cin=>p(240)(108),clock=>clock,reset=>reset,s=>p(288)(108),cout=>p(289)(109));
FA_ff_10058:FAff port map(x=>p(238)(109),y=>p(239)(109),Cin=>p(240)(109),clock=>clock,reset=>reset,s=>p(288)(109),cout=>p(289)(110));
FA_ff_10059:FAff port map(x=>p(238)(110),y=>p(239)(110),Cin=>p(240)(110),clock=>clock,reset=>reset,s=>p(288)(110),cout=>p(289)(111));
FA_ff_10060:FAff port map(x=>p(238)(111),y=>p(239)(111),Cin=>p(240)(111),clock=>clock,reset=>reset,s=>p(288)(111),cout=>p(289)(112));
FA_ff_10061:FAff port map(x=>p(238)(112),y=>p(239)(112),Cin=>p(240)(112),clock=>clock,reset=>reset,s=>p(288)(112),cout=>p(289)(113));
FA_ff_10062:FAff port map(x=>p(238)(113),y=>p(239)(113),Cin=>p(240)(113),clock=>clock,reset=>reset,s=>p(288)(113),cout=>p(289)(114));
FA_ff_10063:FAff port map(x=>p(238)(114),y=>p(239)(114),Cin=>p(240)(114),clock=>clock,reset=>reset,s=>p(288)(114),cout=>p(289)(115));
FA_ff_10064:FAff port map(x=>p(238)(115),y=>p(239)(115),Cin=>p(240)(115),clock=>clock,reset=>reset,s=>p(288)(115),cout=>p(289)(116));
FA_ff_10065:FAff port map(x=>p(238)(116),y=>p(239)(116),Cin=>p(240)(116),clock=>clock,reset=>reset,s=>p(288)(116),cout=>p(289)(117));
FA_ff_10066:FAff port map(x=>p(238)(117),y=>p(239)(117),Cin=>p(240)(117),clock=>clock,reset=>reset,s=>p(288)(117),cout=>p(289)(118));
FA_ff_10067:FAff port map(x=>p(238)(118),y=>p(239)(118),Cin=>p(240)(118),clock=>clock,reset=>reset,s=>p(288)(118),cout=>p(289)(119));
FA_ff_10068:FAff port map(x=>p(238)(119),y=>p(239)(119),Cin=>p(240)(119),clock=>clock,reset=>reset,s=>p(288)(119),cout=>p(289)(120));
FA_ff_10069:FAff port map(x=>p(238)(120),y=>p(239)(120),Cin=>p(240)(120),clock=>clock,reset=>reset,s=>p(288)(120),cout=>p(289)(121));
FA_ff_10070:FAff port map(x=>p(238)(121),y=>p(239)(121),Cin=>p(240)(121),clock=>clock,reset=>reset,s=>p(288)(121),cout=>p(289)(122));
FA_ff_10071:FAff port map(x=>p(238)(122),y=>p(239)(122),Cin=>p(240)(122),clock=>clock,reset=>reset,s=>p(288)(122),cout=>p(289)(123));
FA_ff_10072:FAff port map(x=>p(238)(123),y=>p(239)(123),Cin=>p(240)(123),clock=>clock,reset=>reset,s=>p(288)(123),cout=>p(289)(124));
FA_ff_10073:FAff port map(x=>p(238)(124),y=>p(239)(124),Cin=>p(240)(124),clock=>clock,reset=>reset,s=>p(288)(124),cout=>p(289)(125));
FA_ff_10074:FAff port map(x=>p(238)(125),y=>p(239)(125),Cin=>p(240)(125),clock=>clock,reset=>reset,s=>p(288)(125),cout=>p(289)(126));
FA_ff_10075:FAff port map(x=>p(238)(126),y=>p(239)(126),Cin=>p(240)(126),clock=>clock,reset=>reset,s=>p(288)(126),cout=>p(289)(127));
FA_ff_10076:FAff port map(x=>p(238)(127),y=>p(239)(127),Cin=>p(240)(127),clock=>clock,reset=>reset,s=>p(288)(127),cout=>p(289)(128));
FA_ff_10077:FAff port map(x=>p(238)(128),y=>p(239)(128),Cin=>p(240)(128),clock=>clock,reset=>reset,s=>p(288)(128),cout=>p(289)(129));
p(290)(0)<=p(242)(0);
HA_ff_39:HAff port map(x=>p(242)(1),y=>p(243)(1),clock=>clock,reset=>reset,s=>p(290)(1),c=>p(291)(2));
FA_ff_10078:FAff port map(x=>p(241)(2),y=>p(242)(2),Cin=>p(243)(2),clock=>clock,reset=>reset,s=>p(290)(2),cout=>p(291)(3));
FA_ff_10079:FAff port map(x=>p(241)(3),y=>p(242)(3),Cin=>p(243)(3),clock=>clock,reset=>reset,s=>p(290)(3),cout=>p(291)(4));
FA_ff_10080:FAff port map(x=>p(241)(4),y=>p(242)(4),Cin=>p(243)(4),clock=>clock,reset=>reset,s=>p(290)(4),cout=>p(291)(5));
FA_ff_10081:FAff port map(x=>p(241)(5),y=>p(242)(5),Cin=>p(243)(5),clock=>clock,reset=>reset,s=>p(290)(5),cout=>p(291)(6));
FA_ff_10082:FAff port map(x=>p(241)(6),y=>p(242)(6),Cin=>p(243)(6),clock=>clock,reset=>reset,s=>p(290)(6),cout=>p(291)(7));
FA_ff_10083:FAff port map(x=>p(241)(7),y=>p(242)(7),Cin=>p(243)(7),clock=>clock,reset=>reset,s=>p(290)(7),cout=>p(291)(8));
FA_ff_10084:FAff port map(x=>p(241)(8),y=>p(242)(8),Cin=>p(243)(8),clock=>clock,reset=>reset,s=>p(290)(8),cout=>p(291)(9));
FA_ff_10085:FAff port map(x=>p(241)(9),y=>p(242)(9),Cin=>p(243)(9),clock=>clock,reset=>reset,s=>p(290)(9),cout=>p(291)(10));
FA_ff_10086:FAff port map(x=>p(241)(10),y=>p(242)(10),Cin=>p(243)(10),clock=>clock,reset=>reset,s=>p(290)(10),cout=>p(291)(11));
FA_ff_10087:FAff port map(x=>p(241)(11),y=>p(242)(11),Cin=>p(243)(11),clock=>clock,reset=>reset,s=>p(290)(11),cout=>p(291)(12));
FA_ff_10088:FAff port map(x=>p(241)(12),y=>p(242)(12),Cin=>p(243)(12),clock=>clock,reset=>reset,s=>p(290)(12),cout=>p(291)(13));
FA_ff_10089:FAff port map(x=>p(241)(13),y=>p(242)(13),Cin=>p(243)(13),clock=>clock,reset=>reset,s=>p(290)(13),cout=>p(291)(14));
FA_ff_10090:FAff port map(x=>p(241)(14),y=>p(242)(14),Cin=>p(243)(14),clock=>clock,reset=>reset,s=>p(290)(14),cout=>p(291)(15));
FA_ff_10091:FAff port map(x=>p(241)(15),y=>p(242)(15),Cin=>p(243)(15),clock=>clock,reset=>reset,s=>p(290)(15),cout=>p(291)(16));
FA_ff_10092:FAff port map(x=>p(241)(16),y=>p(242)(16),Cin=>p(243)(16),clock=>clock,reset=>reset,s=>p(290)(16),cout=>p(291)(17));
FA_ff_10093:FAff port map(x=>p(241)(17),y=>p(242)(17),Cin=>p(243)(17),clock=>clock,reset=>reset,s=>p(290)(17),cout=>p(291)(18));
FA_ff_10094:FAff port map(x=>p(241)(18),y=>p(242)(18),Cin=>p(243)(18),clock=>clock,reset=>reset,s=>p(290)(18),cout=>p(291)(19));
FA_ff_10095:FAff port map(x=>p(241)(19),y=>p(242)(19),Cin=>p(243)(19),clock=>clock,reset=>reset,s=>p(290)(19),cout=>p(291)(20));
FA_ff_10096:FAff port map(x=>p(241)(20),y=>p(242)(20),Cin=>p(243)(20),clock=>clock,reset=>reset,s=>p(290)(20),cout=>p(291)(21));
FA_ff_10097:FAff port map(x=>p(241)(21),y=>p(242)(21),Cin=>p(243)(21),clock=>clock,reset=>reset,s=>p(290)(21),cout=>p(291)(22));
FA_ff_10098:FAff port map(x=>p(241)(22),y=>p(242)(22),Cin=>p(243)(22),clock=>clock,reset=>reset,s=>p(290)(22),cout=>p(291)(23));
FA_ff_10099:FAff port map(x=>p(241)(23),y=>p(242)(23),Cin=>p(243)(23),clock=>clock,reset=>reset,s=>p(290)(23),cout=>p(291)(24));
FA_ff_10100:FAff port map(x=>p(241)(24),y=>p(242)(24),Cin=>p(243)(24),clock=>clock,reset=>reset,s=>p(290)(24),cout=>p(291)(25));
FA_ff_10101:FAff port map(x=>p(241)(25),y=>p(242)(25),Cin=>p(243)(25),clock=>clock,reset=>reset,s=>p(290)(25),cout=>p(291)(26));
FA_ff_10102:FAff port map(x=>p(241)(26),y=>p(242)(26),Cin=>p(243)(26),clock=>clock,reset=>reset,s=>p(290)(26),cout=>p(291)(27));
FA_ff_10103:FAff port map(x=>p(241)(27),y=>p(242)(27),Cin=>p(243)(27),clock=>clock,reset=>reset,s=>p(290)(27),cout=>p(291)(28));
FA_ff_10104:FAff port map(x=>p(241)(28),y=>p(242)(28),Cin=>p(243)(28),clock=>clock,reset=>reset,s=>p(290)(28),cout=>p(291)(29));
FA_ff_10105:FAff port map(x=>p(241)(29),y=>p(242)(29),Cin=>p(243)(29),clock=>clock,reset=>reset,s=>p(290)(29),cout=>p(291)(30));
FA_ff_10106:FAff port map(x=>p(241)(30),y=>p(242)(30),Cin=>p(243)(30),clock=>clock,reset=>reset,s=>p(290)(30),cout=>p(291)(31));
FA_ff_10107:FAff port map(x=>p(241)(31),y=>p(242)(31),Cin=>p(243)(31),clock=>clock,reset=>reset,s=>p(290)(31),cout=>p(291)(32));
FA_ff_10108:FAff port map(x=>p(241)(32),y=>p(242)(32),Cin=>p(243)(32),clock=>clock,reset=>reset,s=>p(290)(32),cout=>p(291)(33));
FA_ff_10109:FAff port map(x=>p(241)(33),y=>p(242)(33),Cin=>p(243)(33),clock=>clock,reset=>reset,s=>p(290)(33),cout=>p(291)(34));
FA_ff_10110:FAff port map(x=>p(241)(34),y=>p(242)(34),Cin=>p(243)(34),clock=>clock,reset=>reset,s=>p(290)(34),cout=>p(291)(35));
FA_ff_10111:FAff port map(x=>p(241)(35),y=>p(242)(35),Cin=>p(243)(35),clock=>clock,reset=>reset,s=>p(290)(35),cout=>p(291)(36));
FA_ff_10112:FAff port map(x=>p(241)(36),y=>p(242)(36),Cin=>p(243)(36),clock=>clock,reset=>reset,s=>p(290)(36),cout=>p(291)(37));
FA_ff_10113:FAff port map(x=>p(241)(37),y=>p(242)(37),Cin=>p(243)(37),clock=>clock,reset=>reset,s=>p(290)(37),cout=>p(291)(38));
FA_ff_10114:FAff port map(x=>p(241)(38),y=>p(242)(38),Cin=>p(243)(38),clock=>clock,reset=>reset,s=>p(290)(38),cout=>p(291)(39));
FA_ff_10115:FAff port map(x=>p(241)(39),y=>p(242)(39),Cin=>p(243)(39),clock=>clock,reset=>reset,s=>p(290)(39),cout=>p(291)(40));
FA_ff_10116:FAff port map(x=>p(241)(40),y=>p(242)(40),Cin=>p(243)(40),clock=>clock,reset=>reset,s=>p(290)(40),cout=>p(291)(41));
FA_ff_10117:FAff port map(x=>p(241)(41),y=>p(242)(41),Cin=>p(243)(41),clock=>clock,reset=>reset,s=>p(290)(41),cout=>p(291)(42));
FA_ff_10118:FAff port map(x=>p(241)(42),y=>p(242)(42),Cin=>p(243)(42),clock=>clock,reset=>reset,s=>p(290)(42),cout=>p(291)(43));
FA_ff_10119:FAff port map(x=>p(241)(43),y=>p(242)(43),Cin=>p(243)(43),clock=>clock,reset=>reset,s=>p(290)(43),cout=>p(291)(44));
FA_ff_10120:FAff port map(x=>p(241)(44),y=>p(242)(44),Cin=>p(243)(44),clock=>clock,reset=>reset,s=>p(290)(44),cout=>p(291)(45));
FA_ff_10121:FAff port map(x=>p(241)(45),y=>p(242)(45),Cin=>p(243)(45),clock=>clock,reset=>reset,s=>p(290)(45),cout=>p(291)(46));
FA_ff_10122:FAff port map(x=>p(241)(46),y=>p(242)(46),Cin=>p(243)(46),clock=>clock,reset=>reset,s=>p(290)(46),cout=>p(291)(47));
FA_ff_10123:FAff port map(x=>p(241)(47),y=>p(242)(47),Cin=>p(243)(47),clock=>clock,reset=>reset,s=>p(290)(47),cout=>p(291)(48));
FA_ff_10124:FAff port map(x=>p(241)(48),y=>p(242)(48),Cin=>p(243)(48),clock=>clock,reset=>reset,s=>p(290)(48),cout=>p(291)(49));
FA_ff_10125:FAff port map(x=>p(241)(49),y=>p(242)(49),Cin=>p(243)(49),clock=>clock,reset=>reset,s=>p(290)(49),cout=>p(291)(50));
FA_ff_10126:FAff port map(x=>p(241)(50),y=>p(242)(50),Cin=>p(243)(50),clock=>clock,reset=>reset,s=>p(290)(50),cout=>p(291)(51));
FA_ff_10127:FAff port map(x=>p(241)(51),y=>p(242)(51),Cin=>p(243)(51),clock=>clock,reset=>reset,s=>p(290)(51),cout=>p(291)(52));
FA_ff_10128:FAff port map(x=>p(241)(52),y=>p(242)(52),Cin=>p(243)(52),clock=>clock,reset=>reset,s=>p(290)(52),cout=>p(291)(53));
FA_ff_10129:FAff port map(x=>p(241)(53),y=>p(242)(53),Cin=>p(243)(53),clock=>clock,reset=>reset,s=>p(290)(53),cout=>p(291)(54));
FA_ff_10130:FAff port map(x=>p(241)(54),y=>p(242)(54),Cin=>p(243)(54),clock=>clock,reset=>reset,s=>p(290)(54),cout=>p(291)(55));
FA_ff_10131:FAff port map(x=>p(241)(55),y=>p(242)(55),Cin=>p(243)(55),clock=>clock,reset=>reset,s=>p(290)(55),cout=>p(291)(56));
FA_ff_10132:FAff port map(x=>p(241)(56),y=>p(242)(56),Cin=>p(243)(56),clock=>clock,reset=>reset,s=>p(290)(56),cout=>p(291)(57));
FA_ff_10133:FAff port map(x=>p(241)(57),y=>p(242)(57),Cin=>p(243)(57),clock=>clock,reset=>reset,s=>p(290)(57),cout=>p(291)(58));
FA_ff_10134:FAff port map(x=>p(241)(58),y=>p(242)(58),Cin=>p(243)(58),clock=>clock,reset=>reset,s=>p(290)(58),cout=>p(291)(59));
FA_ff_10135:FAff port map(x=>p(241)(59),y=>p(242)(59),Cin=>p(243)(59),clock=>clock,reset=>reset,s=>p(290)(59),cout=>p(291)(60));
FA_ff_10136:FAff port map(x=>p(241)(60),y=>p(242)(60),Cin=>p(243)(60),clock=>clock,reset=>reset,s=>p(290)(60),cout=>p(291)(61));
FA_ff_10137:FAff port map(x=>p(241)(61),y=>p(242)(61),Cin=>p(243)(61),clock=>clock,reset=>reset,s=>p(290)(61),cout=>p(291)(62));
FA_ff_10138:FAff port map(x=>p(241)(62),y=>p(242)(62),Cin=>p(243)(62),clock=>clock,reset=>reset,s=>p(290)(62),cout=>p(291)(63));
FA_ff_10139:FAff port map(x=>p(241)(63),y=>p(242)(63),Cin=>p(243)(63),clock=>clock,reset=>reset,s=>p(290)(63),cout=>p(291)(64));
FA_ff_10140:FAff port map(x=>p(241)(64),y=>p(242)(64),Cin=>p(243)(64),clock=>clock,reset=>reset,s=>p(290)(64),cout=>p(291)(65));
FA_ff_10141:FAff port map(x=>p(241)(65),y=>p(242)(65),Cin=>p(243)(65),clock=>clock,reset=>reset,s=>p(290)(65),cout=>p(291)(66));
FA_ff_10142:FAff port map(x=>p(241)(66),y=>p(242)(66),Cin=>p(243)(66),clock=>clock,reset=>reset,s=>p(290)(66),cout=>p(291)(67));
FA_ff_10143:FAff port map(x=>p(241)(67),y=>p(242)(67),Cin=>p(243)(67),clock=>clock,reset=>reset,s=>p(290)(67),cout=>p(291)(68));
FA_ff_10144:FAff port map(x=>p(241)(68),y=>p(242)(68),Cin=>p(243)(68),clock=>clock,reset=>reset,s=>p(290)(68),cout=>p(291)(69));
FA_ff_10145:FAff port map(x=>p(241)(69),y=>p(242)(69),Cin=>p(243)(69),clock=>clock,reset=>reset,s=>p(290)(69),cout=>p(291)(70));
FA_ff_10146:FAff port map(x=>p(241)(70),y=>p(242)(70),Cin=>p(243)(70),clock=>clock,reset=>reset,s=>p(290)(70),cout=>p(291)(71));
FA_ff_10147:FAff port map(x=>p(241)(71),y=>p(242)(71),Cin=>p(243)(71),clock=>clock,reset=>reset,s=>p(290)(71),cout=>p(291)(72));
FA_ff_10148:FAff port map(x=>p(241)(72),y=>p(242)(72),Cin=>p(243)(72),clock=>clock,reset=>reset,s=>p(290)(72),cout=>p(291)(73));
FA_ff_10149:FAff port map(x=>p(241)(73),y=>p(242)(73),Cin=>p(243)(73),clock=>clock,reset=>reset,s=>p(290)(73),cout=>p(291)(74));
FA_ff_10150:FAff port map(x=>p(241)(74),y=>p(242)(74),Cin=>p(243)(74),clock=>clock,reset=>reset,s=>p(290)(74),cout=>p(291)(75));
FA_ff_10151:FAff port map(x=>p(241)(75),y=>p(242)(75),Cin=>p(243)(75),clock=>clock,reset=>reset,s=>p(290)(75),cout=>p(291)(76));
FA_ff_10152:FAff port map(x=>p(241)(76),y=>p(242)(76),Cin=>p(243)(76),clock=>clock,reset=>reset,s=>p(290)(76),cout=>p(291)(77));
FA_ff_10153:FAff port map(x=>p(241)(77),y=>p(242)(77),Cin=>p(243)(77),clock=>clock,reset=>reset,s=>p(290)(77),cout=>p(291)(78));
FA_ff_10154:FAff port map(x=>p(241)(78),y=>p(242)(78),Cin=>p(243)(78),clock=>clock,reset=>reset,s=>p(290)(78),cout=>p(291)(79));
FA_ff_10155:FAff port map(x=>p(241)(79),y=>p(242)(79),Cin=>p(243)(79),clock=>clock,reset=>reset,s=>p(290)(79),cout=>p(291)(80));
FA_ff_10156:FAff port map(x=>p(241)(80),y=>p(242)(80),Cin=>p(243)(80),clock=>clock,reset=>reset,s=>p(290)(80),cout=>p(291)(81));
FA_ff_10157:FAff port map(x=>p(241)(81),y=>p(242)(81),Cin=>p(243)(81),clock=>clock,reset=>reset,s=>p(290)(81),cout=>p(291)(82));
FA_ff_10158:FAff port map(x=>p(241)(82),y=>p(242)(82),Cin=>p(243)(82),clock=>clock,reset=>reset,s=>p(290)(82),cout=>p(291)(83));
FA_ff_10159:FAff port map(x=>p(241)(83),y=>p(242)(83),Cin=>p(243)(83),clock=>clock,reset=>reset,s=>p(290)(83),cout=>p(291)(84));
FA_ff_10160:FAff port map(x=>p(241)(84),y=>p(242)(84),Cin=>p(243)(84),clock=>clock,reset=>reset,s=>p(290)(84),cout=>p(291)(85));
FA_ff_10161:FAff port map(x=>p(241)(85),y=>p(242)(85),Cin=>p(243)(85),clock=>clock,reset=>reset,s=>p(290)(85),cout=>p(291)(86));
FA_ff_10162:FAff port map(x=>p(241)(86),y=>p(242)(86),Cin=>p(243)(86),clock=>clock,reset=>reset,s=>p(290)(86),cout=>p(291)(87));
FA_ff_10163:FAff port map(x=>p(241)(87),y=>p(242)(87),Cin=>p(243)(87),clock=>clock,reset=>reset,s=>p(290)(87),cout=>p(291)(88));
FA_ff_10164:FAff port map(x=>p(241)(88),y=>p(242)(88),Cin=>p(243)(88),clock=>clock,reset=>reset,s=>p(290)(88),cout=>p(291)(89));
FA_ff_10165:FAff port map(x=>p(241)(89),y=>p(242)(89),Cin=>p(243)(89),clock=>clock,reset=>reset,s=>p(290)(89),cout=>p(291)(90));
FA_ff_10166:FAff port map(x=>p(241)(90),y=>p(242)(90),Cin=>p(243)(90),clock=>clock,reset=>reset,s=>p(290)(90),cout=>p(291)(91));
FA_ff_10167:FAff port map(x=>p(241)(91),y=>p(242)(91),Cin=>p(243)(91),clock=>clock,reset=>reset,s=>p(290)(91),cout=>p(291)(92));
FA_ff_10168:FAff port map(x=>p(241)(92),y=>p(242)(92),Cin=>p(243)(92),clock=>clock,reset=>reset,s=>p(290)(92),cout=>p(291)(93));
FA_ff_10169:FAff port map(x=>p(241)(93),y=>p(242)(93),Cin=>p(243)(93),clock=>clock,reset=>reset,s=>p(290)(93),cout=>p(291)(94));
FA_ff_10170:FAff port map(x=>p(241)(94),y=>p(242)(94),Cin=>p(243)(94),clock=>clock,reset=>reset,s=>p(290)(94),cout=>p(291)(95));
FA_ff_10171:FAff port map(x=>p(241)(95),y=>p(242)(95),Cin=>p(243)(95),clock=>clock,reset=>reset,s=>p(290)(95),cout=>p(291)(96));
FA_ff_10172:FAff port map(x=>p(241)(96),y=>p(242)(96),Cin=>p(243)(96),clock=>clock,reset=>reset,s=>p(290)(96),cout=>p(291)(97));
FA_ff_10173:FAff port map(x=>p(241)(97),y=>p(242)(97),Cin=>p(243)(97),clock=>clock,reset=>reset,s=>p(290)(97),cout=>p(291)(98));
FA_ff_10174:FAff port map(x=>p(241)(98),y=>p(242)(98),Cin=>p(243)(98),clock=>clock,reset=>reset,s=>p(290)(98),cout=>p(291)(99));
FA_ff_10175:FAff port map(x=>p(241)(99),y=>p(242)(99),Cin=>p(243)(99),clock=>clock,reset=>reset,s=>p(290)(99),cout=>p(291)(100));
FA_ff_10176:FAff port map(x=>p(241)(100),y=>p(242)(100),Cin=>p(243)(100),clock=>clock,reset=>reset,s=>p(290)(100),cout=>p(291)(101));
FA_ff_10177:FAff port map(x=>p(241)(101),y=>p(242)(101),Cin=>p(243)(101),clock=>clock,reset=>reset,s=>p(290)(101),cout=>p(291)(102));
FA_ff_10178:FAff port map(x=>p(241)(102),y=>p(242)(102),Cin=>p(243)(102),clock=>clock,reset=>reset,s=>p(290)(102),cout=>p(291)(103));
FA_ff_10179:FAff port map(x=>p(241)(103),y=>p(242)(103),Cin=>p(243)(103),clock=>clock,reset=>reset,s=>p(290)(103),cout=>p(291)(104));
FA_ff_10180:FAff port map(x=>p(241)(104),y=>p(242)(104),Cin=>p(243)(104),clock=>clock,reset=>reset,s=>p(290)(104),cout=>p(291)(105));
FA_ff_10181:FAff port map(x=>p(241)(105),y=>p(242)(105),Cin=>p(243)(105),clock=>clock,reset=>reset,s=>p(290)(105),cout=>p(291)(106));
FA_ff_10182:FAff port map(x=>p(241)(106),y=>p(242)(106),Cin=>p(243)(106),clock=>clock,reset=>reset,s=>p(290)(106),cout=>p(291)(107));
FA_ff_10183:FAff port map(x=>p(241)(107),y=>p(242)(107),Cin=>p(243)(107),clock=>clock,reset=>reset,s=>p(290)(107),cout=>p(291)(108));
FA_ff_10184:FAff port map(x=>p(241)(108),y=>p(242)(108),Cin=>p(243)(108),clock=>clock,reset=>reset,s=>p(290)(108),cout=>p(291)(109));
FA_ff_10185:FAff port map(x=>p(241)(109),y=>p(242)(109),Cin=>p(243)(109),clock=>clock,reset=>reset,s=>p(290)(109),cout=>p(291)(110));
FA_ff_10186:FAff port map(x=>p(241)(110),y=>p(242)(110),Cin=>p(243)(110),clock=>clock,reset=>reset,s=>p(290)(110),cout=>p(291)(111));
FA_ff_10187:FAff port map(x=>p(241)(111),y=>p(242)(111),Cin=>p(243)(111),clock=>clock,reset=>reset,s=>p(290)(111),cout=>p(291)(112));
FA_ff_10188:FAff port map(x=>p(241)(112),y=>p(242)(112),Cin=>p(243)(112),clock=>clock,reset=>reset,s=>p(290)(112),cout=>p(291)(113));
FA_ff_10189:FAff port map(x=>p(241)(113),y=>p(242)(113),Cin=>p(243)(113),clock=>clock,reset=>reset,s=>p(290)(113),cout=>p(291)(114));
FA_ff_10190:FAff port map(x=>p(241)(114),y=>p(242)(114),Cin=>p(243)(114),clock=>clock,reset=>reset,s=>p(290)(114),cout=>p(291)(115));
FA_ff_10191:FAff port map(x=>p(241)(115),y=>p(242)(115),Cin=>p(243)(115),clock=>clock,reset=>reset,s=>p(290)(115),cout=>p(291)(116));
FA_ff_10192:FAff port map(x=>p(241)(116),y=>p(242)(116),Cin=>p(243)(116),clock=>clock,reset=>reset,s=>p(290)(116),cout=>p(291)(117));
FA_ff_10193:FAff port map(x=>p(241)(117),y=>p(242)(117),Cin=>p(243)(117),clock=>clock,reset=>reset,s=>p(290)(117),cout=>p(291)(118));
FA_ff_10194:FAff port map(x=>p(241)(118),y=>p(242)(118),Cin=>p(243)(118),clock=>clock,reset=>reset,s=>p(290)(118),cout=>p(291)(119));
FA_ff_10195:FAff port map(x=>p(241)(119),y=>p(242)(119),Cin=>p(243)(119),clock=>clock,reset=>reset,s=>p(290)(119),cout=>p(291)(120));
FA_ff_10196:FAff port map(x=>p(241)(120),y=>p(242)(120),Cin=>p(243)(120),clock=>clock,reset=>reset,s=>p(290)(120),cout=>p(291)(121));
FA_ff_10197:FAff port map(x=>p(241)(121),y=>p(242)(121),Cin=>p(243)(121),clock=>clock,reset=>reset,s=>p(290)(121),cout=>p(291)(122));
FA_ff_10198:FAff port map(x=>p(241)(122),y=>p(242)(122),Cin=>p(243)(122),clock=>clock,reset=>reset,s=>p(290)(122),cout=>p(291)(123));
FA_ff_10199:FAff port map(x=>p(241)(123),y=>p(242)(123),Cin=>p(243)(123),clock=>clock,reset=>reset,s=>p(290)(123),cout=>p(291)(124));
FA_ff_10200:FAff port map(x=>p(241)(124),y=>p(242)(124),Cin=>p(243)(124),clock=>clock,reset=>reset,s=>p(290)(124),cout=>p(291)(125));
FA_ff_10201:FAff port map(x=>p(241)(125),y=>p(242)(125),Cin=>p(243)(125),clock=>clock,reset=>reset,s=>p(290)(125),cout=>p(291)(126));
FA_ff_10202:FAff port map(x=>p(241)(126),y=>p(242)(126),Cin=>p(243)(126),clock=>clock,reset=>reset,s=>p(290)(126),cout=>p(291)(127));
FA_ff_10203:FAff port map(x=>p(241)(127),y=>p(242)(127),Cin=>p(243)(127),clock=>clock,reset=>reset,s=>p(290)(127),cout=>p(291)(128));
FA_ff_10204:FAff port map(x=>p(241)(128),y=>p(242)(128),Cin=>p(243)(128),clock=>clock,reset=>reset,s=>p(290)(128),cout=>p(291)(129));
p(290)(129)<=p(241)(129);
HA_ff_40:HAff port map(x=>p(244)(0),y=>p(246)(0),clock=>clock,reset=>reset,s=>p(292)(0),c=>p(293)(1));
HA_ff_41:HAff port map(x=>p(244)(1),y=>p(246)(1),clock=>clock,reset=>reset,s=>p(292)(1),c=>p(293)(2));
FA_ff_10205:FAff port map(x=>p(244)(2),y=>p(245)(2),Cin=>p(246)(2),clock=>clock,reset=>reset,s=>p(292)(2),cout=>p(293)(3));
FA_ff_10206:FAff port map(x=>p(244)(3),y=>p(245)(3),Cin=>p(246)(3),clock=>clock,reset=>reset,s=>p(292)(3),cout=>p(293)(4));
FA_ff_10207:FAff port map(x=>p(244)(4),y=>p(245)(4),Cin=>p(246)(4),clock=>clock,reset=>reset,s=>p(292)(4),cout=>p(293)(5));
FA_ff_10208:FAff port map(x=>p(244)(5),y=>p(245)(5),Cin=>p(246)(5),clock=>clock,reset=>reset,s=>p(292)(5),cout=>p(293)(6));
FA_ff_10209:FAff port map(x=>p(244)(6),y=>p(245)(6),Cin=>p(246)(6),clock=>clock,reset=>reset,s=>p(292)(6),cout=>p(293)(7));
FA_ff_10210:FAff port map(x=>p(244)(7),y=>p(245)(7),Cin=>p(246)(7),clock=>clock,reset=>reset,s=>p(292)(7),cout=>p(293)(8));
FA_ff_10211:FAff port map(x=>p(244)(8),y=>p(245)(8),Cin=>p(246)(8),clock=>clock,reset=>reset,s=>p(292)(8),cout=>p(293)(9));
FA_ff_10212:FAff port map(x=>p(244)(9),y=>p(245)(9),Cin=>p(246)(9),clock=>clock,reset=>reset,s=>p(292)(9),cout=>p(293)(10));
FA_ff_10213:FAff port map(x=>p(244)(10),y=>p(245)(10),Cin=>p(246)(10),clock=>clock,reset=>reset,s=>p(292)(10),cout=>p(293)(11));
FA_ff_10214:FAff port map(x=>p(244)(11),y=>p(245)(11),Cin=>p(246)(11),clock=>clock,reset=>reset,s=>p(292)(11),cout=>p(293)(12));
FA_ff_10215:FAff port map(x=>p(244)(12),y=>p(245)(12),Cin=>p(246)(12),clock=>clock,reset=>reset,s=>p(292)(12),cout=>p(293)(13));
FA_ff_10216:FAff port map(x=>p(244)(13),y=>p(245)(13),Cin=>p(246)(13),clock=>clock,reset=>reset,s=>p(292)(13),cout=>p(293)(14));
FA_ff_10217:FAff port map(x=>p(244)(14),y=>p(245)(14),Cin=>p(246)(14),clock=>clock,reset=>reset,s=>p(292)(14),cout=>p(293)(15));
FA_ff_10218:FAff port map(x=>p(244)(15),y=>p(245)(15),Cin=>p(246)(15),clock=>clock,reset=>reset,s=>p(292)(15),cout=>p(293)(16));
FA_ff_10219:FAff port map(x=>p(244)(16),y=>p(245)(16),Cin=>p(246)(16),clock=>clock,reset=>reset,s=>p(292)(16),cout=>p(293)(17));
FA_ff_10220:FAff port map(x=>p(244)(17),y=>p(245)(17),Cin=>p(246)(17),clock=>clock,reset=>reset,s=>p(292)(17),cout=>p(293)(18));
FA_ff_10221:FAff port map(x=>p(244)(18),y=>p(245)(18),Cin=>p(246)(18),clock=>clock,reset=>reset,s=>p(292)(18),cout=>p(293)(19));
FA_ff_10222:FAff port map(x=>p(244)(19),y=>p(245)(19),Cin=>p(246)(19),clock=>clock,reset=>reset,s=>p(292)(19),cout=>p(293)(20));
FA_ff_10223:FAff port map(x=>p(244)(20),y=>p(245)(20),Cin=>p(246)(20),clock=>clock,reset=>reset,s=>p(292)(20),cout=>p(293)(21));
FA_ff_10224:FAff port map(x=>p(244)(21),y=>p(245)(21),Cin=>p(246)(21),clock=>clock,reset=>reset,s=>p(292)(21),cout=>p(293)(22));
FA_ff_10225:FAff port map(x=>p(244)(22),y=>p(245)(22),Cin=>p(246)(22),clock=>clock,reset=>reset,s=>p(292)(22),cout=>p(293)(23));
FA_ff_10226:FAff port map(x=>p(244)(23),y=>p(245)(23),Cin=>p(246)(23),clock=>clock,reset=>reset,s=>p(292)(23),cout=>p(293)(24));
FA_ff_10227:FAff port map(x=>p(244)(24),y=>p(245)(24),Cin=>p(246)(24),clock=>clock,reset=>reset,s=>p(292)(24),cout=>p(293)(25));
FA_ff_10228:FAff port map(x=>p(244)(25),y=>p(245)(25),Cin=>p(246)(25),clock=>clock,reset=>reset,s=>p(292)(25),cout=>p(293)(26));
FA_ff_10229:FAff port map(x=>p(244)(26),y=>p(245)(26),Cin=>p(246)(26),clock=>clock,reset=>reset,s=>p(292)(26),cout=>p(293)(27));
FA_ff_10230:FAff port map(x=>p(244)(27),y=>p(245)(27),Cin=>p(246)(27),clock=>clock,reset=>reset,s=>p(292)(27),cout=>p(293)(28));
FA_ff_10231:FAff port map(x=>p(244)(28),y=>p(245)(28),Cin=>p(246)(28),clock=>clock,reset=>reset,s=>p(292)(28),cout=>p(293)(29));
FA_ff_10232:FAff port map(x=>p(244)(29),y=>p(245)(29),Cin=>p(246)(29),clock=>clock,reset=>reset,s=>p(292)(29),cout=>p(293)(30));
FA_ff_10233:FAff port map(x=>p(244)(30),y=>p(245)(30),Cin=>p(246)(30),clock=>clock,reset=>reset,s=>p(292)(30),cout=>p(293)(31));
FA_ff_10234:FAff port map(x=>p(244)(31),y=>p(245)(31),Cin=>p(246)(31),clock=>clock,reset=>reset,s=>p(292)(31),cout=>p(293)(32));
FA_ff_10235:FAff port map(x=>p(244)(32),y=>p(245)(32),Cin=>p(246)(32),clock=>clock,reset=>reset,s=>p(292)(32),cout=>p(293)(33));
FA_ff_10236:FAff port map(x=>p(244)(33),y=>p(245)(33),Cin=>p(246)(33),clock=>clock,reset=>reset,s=>p(292)(33),cout=>p(293)(34));
FA_ff_10237:FAff port map(x=>p(244)(34),y=>p(245)(34),Cin=>p(246)(34),clock=>clock,reset=>reset,s=>p(292)(34),cout=>p(293)(35));
FA_ff_10238:FAff port map(x=>p(244)(35),y=>p(245)(35),Cin=>p(246)(35),clock=>clock,reset=>reset,s=>p(292)(35),cout=>p(293)(36));
FA_ff_10239:FAff port map(x=>p(244)(36),y=>p(245)(36),Cin=>p(246)(36),clock=>clock,reset=>reset,s=>p(292)(36),cout=>p(293)(37));
FA_ff_10240:FAff port map(x=>p(244)(37),y=>p(245)(37),Cin=>p(246)(37),clock=>clock,reset=>reset,s=>p(292)(37),cout=>p(293)(38));
FA_ff_10241:FAff port map(x=>p(244)(38),y=>p(245)(38),Cin=>p(246)(38),clock=>clock,reset=>reset,s=>p(292)(38),cout=>p(293)(39));
FA_ff_10242:FAff port map(x=>p(244)(39),y=>p(245)(39),Cin=>p(246)(39),clock=>clock,reset=>reset,s=>p(292)(39),cout=>p(293)(40));
FA_ff_10243:FAff port map(x=>p(244)(40),y=>p(245)(40),Cin=>p(246)(40),clock=>clock,reset=>reset,s=>p(292)(40),cout=>p(293)(41));
FA_ff_10244:FAff port map(x=>p(244)(41),y=>p(245)(41),Cin=>p(246)(41),clock=>clock,reset=>reset,s=>p(292)(41),cout=>p(293)(42));
FA_ff_10245:FAff port map(x=>p(244)(42),y=>p(245)(42),Cin=>p(246)(42),clock=>clock,reset=>reset,s=>p(292)(42),cout=>p(293)(43));
FA_ff_10246:FAff port map(x=>p(244)(43),y=>p(245)(43),Cin=>p(246)(43),clock=>clock,reset=>reset,s=>p(292)(43),cout=>p(293)(44));
FA_ff_10247:FAff port map(x=>p(244)(44),y=>p(245)(44),Cin=>p(246)(44),clock=>clock,reset=>reset,s=>p(292)(44),cout=>p(293)(45));
FA_ff_10248:FAff port map(x=>p(244)(45),y=>p(245)(45),Cin=>p(246)(45),clock=>clock,reset=>reset,s=>p(292)(45),cout=>p(293)(46));
FA_ff_10249:FAff port map(x=>p(244)(46),y=>p(245)(46),Cin=>p(246)(46),clock=>clock,reset=>reset,s=>p(292)(46),cout=>p(293)(47));
FA_ff_10250:FAff port map(x=>p(244)(47),y=>p(245)(47),Cin=>p(246)(47),clock=>clock,reset=>reset,s=>p(292)(47),cout=>p(293)(48));
FA_ff_10251:FAff port map(x=>p(244)(48),y=>p(245)(48),Cin=>p(246)(48),clock=>clock,reset=>reset,s=>p(292)(48),cout=>p(293)(49));
FA_ff_10252:FAff port map(x=>p(244)(49),y=>p(245)(49),Cin=>p(246)(49),clock=>clock,reset=>reset,s=>p(292)(49),cout=>p(293)(50));
FA_ff_10253:FAff port map(x=>p(244)(50),y=>p(245)(50),Cin=>p(246)(50),clock=>clock,reset=>reset,s=>p(292)(50),cout=>p(293)(51));
FA_ff_10254:FAff port map(x=>p(244)(51),y=>p(245)(51),Cin=>p(246)(51),clock=>clock,reset=>reset,s=>p(292)(51),cout=>p(293)(52));
FA_ff_10255:FAff port map(x=>p(244)(52),y=>p(245)(52),Cin=>p(246)(52),clock=>clock,reset=>reset,s=>p(292)(52),cout=>p(293)(53));
FA_ff_10256:FAff port map(x=>p(244)(53),y=>p(245)(53),Cin=>p(246)(53),clock=>clock,reset=>reset,s=>p(292)(53),cout=>p(293)(54));
FA_ff_10257:FAff port map(x=>p(244)(54),y=>p(245)(54),Cin=>p(246)(54),clock=>clock,reset=>reset,s=>p(292)(54),cout=>p(293)(55));
FA_ff_10258:FAff port map(x=>p(244)(55),y=>p(245)(55),Cin=>p(246)(55),clock=>clock,reset=>reset,s=>p(292)(55),cout=>p(293)(56));
FA_ff_10259:FAff port map(x=>p(244)(56),y=>p(245)(56),Cin=>p(246)(56),clock=>clock,reset=>reset,s=>p(292)(56),cout=>p(293)(57));
FA_ff_10260:FAff port map(x=>p(244)(57),y=>p(245)(57),Cin=>p(246)(57),clock=>clock,reset=>reset,s=>p(292)(57),cout=>p(293)(58));
FA_ff_10261:FAff port map(x=>p(244)(58),y=>p(245)(58),Cin=>p(246)(58),clock=>clock,reset=>reset,s=>p(292)(58),cout=>p(293)(59));
FA_ff_10262:FAff port map(x=>p(244)(59),y=>p(245)(59),Cin=>p(246)(59),clock=>clock,reset=>reset,s=>p(292)(59),cout=>p(293)(60));
FA_ff_10263:FAff port map(x=>p(244)(60),y=>p(245)(60),Cin=>p(246)(60),clock=>clock,reset=>reset,s=>p(292)(60),cout=>p(293)(61));
FA_ff_10264:FAff port map(x=>p(244)(61),y=>p(245)(61),Cin=>p(246)(61),clock=>clock,reset=>reset,s=>p(292)(61),cout=>p(293)(62));
FA_ff_10265:FAff port map(x=>p(244)(62),y=>p(245)(62),Cin=>p(246)(62),clock=>clock,reset=>reset,s=>p(292)(62),cout=>p(293)(63));
FA_ff_10266:FAff port map(x=>p(244)(63),y=>p(245)(63),Cin=>p(246)(63),clock=>clock,reset=>reset,s=>p(292)(63),cout=>p(293)(64));
FA_ff_10267:FAff port map(x=>p(244)(64),y=>p(245)(64),Cin=>p(246)(64),clock=>clock,reset=>reset,s=>p(292)(64),cout=>p(293)(65));
FA_ff_10268:FAff port map(x=>p(244)(65),y=>p(245)(65),Cin=>p(246)(65),clock=>clock,reset=>reset,s=>p(292)(65),cout=>p(293)(66));
FA_ff_10269:FAff port map(x=>p(244)(66),y=>p(245)(66),Cin=>p(246)(66),clock=>clock,reset=>reset,s=>p(292)(66),cout=>p(293)(67));
FA_ff_10270:FAff port map(x=>p(244)(67),y=>p(245)(67),Cin=>p(246)(67),clock=>clock,reset=>reset,s=>p(292)(67),cout=>p(293)(68));
FA_ff_10271:FAff port map(x=>p(244)(68),y=>p(245)(68),Cin=>p(246)(68),clock=>clock,reset=>reset,s=>p(292)(68),cout=>p(293)(69));
FA_ff_10272:FAff port map(x=>p(244)(69),y=>p(245)(69),Cin=>p(246)(69),clock=>clock,reset=>reset,s=>p(292)(69),cout=>p(293)(70));
FA_ff_10273:FAff port map(x=>p(244)(70),y=>p(245)(70),Cin=>p(246)(70),clock=>clock,reset=>reset,s=>p(292)(70),cout=>p(293)(71));
FA_ff_10274:FAff port map(x=>p(244)(71),y=>p(245)(71),Cin=>p(246)(71),clock=>clock,reset=>reset,s=>p(292)(71),cout=>p(293)(72));
FA_ff_10275:FAff port map(x=>p(244)(72),y=>p(245)(72),Cin=>p(246)(72),clock=>clock,reset=>reset,s=>p(292)(72),cout=>p(293)(73));
FA_ff_10276:FAff port map(x=>p(244)(73),y=>p(245)(73),Cin=>p(246)(73),clock=>clock,reset=>reset,s=>p(292)(73),cout=>p(293)(74));
FA_ff_10277:FAff port map(x=>p(244)(74),y=>p(245)(74),Cin=>p(246)(74),clock=>clock,reset=>reset,s=>p(292)(74),cout=>p(293)(75));
FA_ff_10278:FAff port map(x=>p(244)(75),y=>p(245)(75),Cin=>p(246)(75),clock=>clock,reset=>reset,s=>p(292)(75),cout=>p(293)(76));
FA_ff_10279:FAff port map(x=>p(244)(76),y=>p(245)(76),Cin=>p(246)(76),clock=>clock,reset=>reset,s=>p(292)(76),cout=>p(293)(77));
FA_ff_10280:FAff port map(x=>p(244)(77),y=>p(245)(77),Cin=>p(246)(77),clock=>clock,reset=>reset,s=>p(292)(77),cout=>p(293)(78));
FA_ff_10281:FAff port map(x=>p(244)(78),y=>p(245)(78),Cin=>p(246)(78),clock=>clock,reset=>reset,s=>p(292)(78),cout=>p(293)(79));
FA_ff_10282:FAff port map(x=>p(244)(79),y=>p(245)(79),Cin=>p(246)(79),clock=>clock,reset=>reset,s=>p(292)(79),cout=>p(293)(80));
FA_ff_10283:FAff port map(x=>p(244)(80),y=>p(245)(80),Cin=>p(246)(80),clock=>clock,reset=>reset,s=>p(292)(80),cout=>p(293)(81));
FA_ff_10284:FAff port map(x=>p(244)(81),y=>p(245)(81),Cin=>p(246)(81),clock=>clock,reset=>reset,s=>p(292)(81),cout=>p(293)(82));
FA_ff_10285:FAff port map(x=>p(244)(82),y=>p(245)(82),Cin=>p(246)(82),clock=>clock,reset=>reset,s=>p(292)(82),cout=>p(293)(83));
FA_ff_10286:FAff port map(x=>p(244)(83),y=>p(245)(83),Cin=>p(246)(83),clock=>clock,reset=>reset,s=>p(292)(83),cout=>p(293)(84));
FA_ff_10287:FAff port map(x=>p(244)(84),y=>p(245)(84),Cin=>p(246)(84),clock=>clock,reset=>reset,s=>p(292)(84),cout=>p(293)(85));
FA_ff_10288:FAff port map(x=>p(244)(85),y=>p(245)(85),Cin=>p(246)(85),clock=>clock,reset=>reset,s=>p(292)(85),cout=>p(293)(86));
FA_ff_10289:FAff port map(x=>p(244)(86),y=>p(245)(86),Cin=>p(246)(86),clock=>clock,reset=>reset,s=>p(292)(86),cout=>p(293)(87));
FA_ff_10290:FAff port map(x=>p(244)(87),y=>p(245)(87),Cin=>p(246)(87),clock=>clock,reset=>reset,s=>p(292)(87),cout=>p(293)(88));
FA_ff_10291:FAff port map(x=>p(244)(88),y=>p(245)(88),Cin=>p(246)(88),clock=>clock,reset=>reset,s=>p(292)(88),cout=>p(293)(89));
FA_ff_10292:FAff port map(x=>p(244)(89),y=>p(245)(89),Cin=>p(246)(89),clock=>clock,reset=>reset,s=>p(292)(89),cout=>p(293)(90));
FA_ff_10293:FAff port map(x=>p(244)(90),y=>p(245)(90),Cin=>p(246)(90),clock=>clock,reset=>reset,s=>p(292)(90),cout=>p(293)(91));
FA_ff_10294:FAff port map(x=>p(244)(91),y=>p(245)(91),Cin=>p(246)(91),clock=>clock,reset=>reset,s=>p(292)(91),cout=>p(293)(92));
FA_ff_10295:FAff port map(x=>p(244)(92),y=>p(245)(92),Cin=>p(246)(92),clock=>clock,reset=>reset,s=>p(292)(92),cout=>p(293)(93));
FA_ff_10296:FAff port map(x=>p(244)(93),y=>p(245)(93),Cin=>p(246)(93),clock=>clock,reset=>reset,s=>p(292)(93),cout=>p(293)(94));
FA_ff_10297:FAff port map(x=>p(244)(94),y=>p(245)(94),Cin=>p(246)(94),clock=>clock,reset=>reset,s=>p(292)(94),cout=>p(293)(95));
FA_ff_10298:FAff port map(x=>p(244)(95),y=>p(245)(95),Cin=>p(246)(95),clock=>clock,reset=>reset,s=>p(292)(95),cout=>p(293)(96));
FA_ff_10299:FAff port map(x=>p(244)(96),y=>p(245)(96),Cin=>p(246)(96),clock=>clock,reset=>reset,s=>p(292)(96),cout=>p(293)(97));
FA_ff_10300:FAff port map(x=>p(244)(97),y=>p(245)(97),Cin=>p(246)(97),clock=>clock,reset=>reset,s=>p(292)(97),cout=>p(293)(98));
FA_ff_10301:FAff port map(x=>p(244)(98),y=>p(245)(98),Cin=>p(246)(98),clock=>clock,reset=>reset,s=>p(292)(98),cout=>p(293)(99));
FA_ff_10302:FAff port map(x=>p(244)(99),y=>p(245)(99),Cin=>p(246)(99),clock=>clock,reset=>reset,s=>p(292)(99),cout=>p(293)(100));
FA_ff_10303:FAff port map(x=>p(244)(100),y=>p(245)(100),Cin=>p(246)(100),clock=>clock,reset=>reset,s=>p(292)(100),cout=>p(293)(101));
FA_ff_10304:FAff port map(x=>p(244)(101),y=>p(245)(101),Cin=>p(246)(101),clock=>clock,reset=>reset,s=>p(292)(101),cout=>p(293)(102));
FA_ff_10305:FAff port map(x=>p(244)(102),y=>p(245)(102),Cin=>p(246)(102),clock=>clock,reset=>reset,s=>p(292)(102),cout=>p(293)(103));
FA_ff_10306:FAff port map(x=>p(244)(103),y=>p(245)(103),Cin=>p(246)(103),clock=>clock,reset=>reset,s=>p(292)(103),cout=>p(293)(104));
FA_ff_10307:FAff port map(x=>p(244)(104),y=>p(245)(104),Cin=>p(246)(104),clock=>clock,reset=>reset,s=>p(292)(104),cout=>p(293)(105));
FA_ff_10308:FAff port map(x=>p(244)(105),y=>p(245)(105),Cin=>p(246)(105),clock=>clock,reset=>reset,s=>p(292)(105),cout=>p(293)(106));
FA_ff_10309:FAff port map(x=>p(244)(106),y=>p(245)(106),Cin=>p(246)(106),clock=>clock,reset=>reset,s=>p(292)(106),cout=>p(293)(107));
FA_ff_10310:FAff port map(x=>p(244)(107),y=>p(245)(107),Cin=>p(246)(107),clock=>clock,reset=>reset,s=>p(292)(107),cout=>p(293)(108));
FA_ff_10311:FAff port map(x=>p(244)(108),y=>p(245)(108),Cin=>p(246)(108),clock=>clock,reset=>reset,s=>p(292)(108),cout=>p(293)(109));
FA_ff_10312:FAff port map(x=>p(244)(109),y=>p(245)(109),Cin=>p(246)(109),clock=>clock,reset=>reset,s=>p(292)(109),cout=>p(293)(110));
FA_ff_10313:FAff port map(x=>p(244)(110),y=>p(245)(110),Cin=>p(246)(110),clock=>clock,reset=>reset,s=>p(292)(110),cout=>p(293)(111));
FA_ff_10314:FAff port map(x=>p(244)(111),y=>p(245)(111),Cin=>p(246)(111),clock=>clock,reset=>reset,s=>p(292)(111),cout=>p(293)(112));
FA_ff_10315:FAff port map(x=>p(244)(112),y=>p(245)(112),Cin=>p(246)(112),clock=>clock,reset=>reset,s=>p(292)(112),cout=>p(293)(113));
FA_ff_10316:FAff port map(x=>p(244)(113),y=>p(245)(113),Cin=>p(246)(113),clock=>clock,reset=>reset,s=>p(292)(113),cout=>p(293)(114));
FA_ff_10317:FAff port map(x=>p(244)(114),y=>p(245)(114),Cin=>p(246)(114),clock=>clock,reset=>reset,s=>p(292)(114),cout=>p(293)(115));
FA_ff_10318:FAff port map(x=>p(244)(115),y=>p(245)(115),Cin=>p(246)(115),clock=>clock,reset=>reset,s=>p(292)(115),cout=>p(293)(116));
FA_ff_10319:FAff port map(x=>p(244)(116),y=>p(245)(116),Cin=>p(246)(116),clock=>clock,reset=>reset,s=>p(292)(116),cout=>p(293)(117));
FA_ff_10320:FAff port map(x=>p(244)(117),y=>p(245)(117),Cin=>p(246)(117),clock=>clock,reset=>reset,s=>p(292)(117),cout=>p(293)(118));
FA_ff_10321:FAff port map(x=>p(244)(118),y=>p(245)(118),Cin=>p(246)(118),clock=>clock,reset=>reset,s=>p(292)(118),cout=>p(293)(119));
FA_ff_10322:FAff port map(x=>p(244)(119),y=>p(245)(119),Cin=>p(246)(119),clock=>clock,reset=>reset,s=>p(292)(119),cout=>p(293)(120));
FA_ff_10323:FAff port map(x=>p(244)(120),y=>p(245)(120),Cin=>p(246)(120),clock=>clock,reset=>reset,s=>p(292)(120),cout=>p(293)(121));
FA_ff_10324:FAff port map(x=>p(244)(121),y=>p(245)(121),Cin=>p(246)(121),clock=>clock,reset=>reset,s=>p(292)(121),cout=>p(293)(122));
FA_ff_10325:FAff port map(x=>p(244)(122),y=>p(245)(122),Cin=>p(246)(122),clock=>clock,reset=>reset,s=>p(292)(122),cout=>p(293)(123));
FA_ff_10326:FAff port map(x=>p(244)(123),y=>p(245)(123),Cin=>p(246)(123),clock=>clock,reset=>reset,s=>p(292)(123),cout=>p(293)(124));
FA_ff_10327:FAff port map(x=>p(244)(124),y=>p(245)(124),Cin=>p(246)(124),clock=>clock,reset=>reset,s=>p(292)(124),cout=>p(293)(125));
FA_ff_10328:FAff port map(x=>p(244)(125),y=>p(245)(125),Cin=>p(246)(125),clock=>clock,reset=>reset,s=>p(292)(125),cout=>p(293)(126));
FA_ff_10329:FAff port map(x=>p(244)(126),y=>p(245)(126),Cin=>p(246)(126),clock=>clock,reset=>reset,s=>p(292)(126),cout=>p(293)(127));
FA_ff_10330:FAff port map(x=>p(244)(127),y=>p(245)(127),Cin=>p(246)(127),clock=>clock,reset=>reset,s=>p(292)(127),cout=>p(293)(128));
FA_ff_10331:FAff port map(x=>p(244)(128),y=>p(245)(128),Cin=>p(246)(128),clock=>clock,reset=>reset,s=>p(292)(128),cout=>p(293)(129));
p(292)(129)<=p(245)(129);
p(294)(0)<=p(248)(0);
HA_ff_42:HAff port map(x=>p(247)(1),y=>p(248)(1),clock=>clock,reset=>reset,s=>p(294)(1),c=>p(295)(2));
FA_ff_10332:FAff port map(x=>p(247)(2),y=>p(248)(2),Cin=>p(249)(2),clock=>clock,reset=>reset,s=>p(294)(2),cout=>p(295)(3));
FA_ff_10333:FAff port map(x=>p(247)(3),y=>p(248)(3),Cin=>p(249)(3),clock=>clock,reset=>reset,s=>p(294)(3),cout=>p(295)(4));
FA_ff_10334:FAff port map(x=>p(247)(4),y=>p(248)(4),Cin=>p(249)(4),clock=>clock,reset=>reset,s=>p(294)(4),cout=>p(295)(5));
FA_ff_10335:FAff port map(x=>p(247)(5),y=>p(248)(5),Cin=>p(249)(5),clock=>clock,reset=>reset,s=>p(294)(5),cout=>p(295)(6));
FA_ff_10336:FAff port map(x=>p(247)(6),y=>p(248)(6),Cin=>p(249)(6),clock=>clock,reset=>reset,s=>p(294)(6),cout=>p(295)(7));
FA_ff_10337:FAff port map(x=>p(247)(7),y=>p(248)(7),Cin=>p(249)(7),clock=>clock,reset=>reset,s=>p(294)(7),cout=>p(295)(8));
FA_ff_10338:FAff port map(x=>p(247)(8),y=>p(248)(8),Cin=>p(249)(8),clock=>clock,reset=>reset,s=>p(294)(8),cout=>p(295)(9));
FA_ff_10339:FAff port map(x=>p(247)(9),y=>p(248)(9),Cin=>p(249)(9),clock=>clock,reset=>reset,s=>p(294)(9),cout=>p(295)(10));
FA_ff_10340:FAff port map(x=>p(247)(10),y=>p(248)(10),Cin=>p(249)(10),clock=>clock,reset=>reset,s=>p(294)(10),cout=>p(295)(11));
FA_ff_10341:FAff port map(x=>p(247)(11),y=>p(248)(11),Cin=>p(249)(11),clock=>clock,reset=>reset,s=>p(294)(11),cout=>p(295)(12));
FA_ff_10342:FAff port map(x=>p(247)(12),y=>p(248)(12),Cin=>p(249)(12),clock=>clock,reset=>reset,s=>p(294)(12),cout=>p(295)(13));
FA_ff_10343:FAff port map(x=>p(247)(13),y=>p(248)(13),Cin=>p(249)(13),clock=>clock,reset=>reset,s=>p(294)(13),cout=>p(295)(14));
FA_ff_10344:FAff port map(x=>p(247)(14),y=>p(248)(14),Cin=>p(249)(14),clock=>clock,reset=>reset,s=>p(294)(14),cout=>p(295)(15));
FA_ff_10345:FAff port map(x=>p(247)(15),y=>p(248)(15),Cin=>p(249)(15),clock=>clock,reset=>reset,s=>p(294)(15),cout=>p(295)(16));
FA_ff_10346:FAff port map(x=>p(247)(16),y=>p(248)(16),Cin=>p(249)(16),clock=>clock,reset=>reset,s=>p(294)(16),cout=>p(295)(17));
FA_ff_10347:FAff port map(x=>p(247)(17),y=>p(248)(17),Cin=>p(249)(17),clock=>clock,reset=>reset,s=>p(294)(17),cout=>p(295)(18));
FA_ff_10348:FAff port map(x=>p(247)(18),y=>p(248)(18),Cin=>p(249)(18),clock=>clock,reset=>reset,s=>p(294)(18),cout=>p(295)(19));
FA_ff_10349:FAff port map(x=>p(247)(19),y=>p(248)(19),Cin=>p(249)(19),clock=>clock,reset=>reset,s=>p(294)(19),cout=>p(295)(20));
FA_ff_10350:FAff port map(x=>p(247)(20),y=>p(248)(20),Cin=>p(249)(20),clock=>clock,reset=>reset,s=>p(294)(20),cout=>p(295)(21));
FA_ff_10351:FAff port map(x=>p(247)(21),y=>p(248)(21),Cin=>p(249)(21),clock=>clock,reset=>reset,s=>p(294)(21),cout=>p(295)(22));
FA_ff_10352:FAff port map(x=>p(247)(22),y=>p(248)(22),Cin=>p(249)(22),clock=>clock,reset=>reset,s=>p(294)(22),cout=>p(295)(23));
FA_ff_10353:FAff port map(x=>p(247)(23),y=>p(248)(23),Cin=>p(249)(23),clock=>clock,reset=>reset,s=>p(294)(23),cout=>p(295)(24));
FA_ff_10354:FAff port map(x=>p(247)(24),y=>p(248)(24),Cin=>p(249)(24),clock=>clock,reset=>reset,s=>p(294)(24),cout=>p(295)(25));
FA_ff_10355:FAff port map(x=>p(247)(25),y=>p(248)(25),Cin=>p(249)(25),clock=>clock,reset=>reset,s=>p(294)(25),cout=>p(295)(26));
FA_ff_10356:FAff port map(x=>p(247)(26),y=>p(248)(26),Cin=>p(249)(26),clock=>clock,reset=>reset,s=>p(294)(26),cout=>p(295)(27));
FA_ff_10357:FAff port map(x=>p(247)(27),y=>p(248)(27),Cin=>p(249)(27),clock=>clock,reset=>reset,s=>p(294)(27),cout=>p(295)(28));
FA_ff_10358:FAff port map(x=>p(247)(28),y=>p(248)(28),Cin=>p(249)(28),clock=>clock,reset=>reset,s=>p(294)(28),cout=>p(295)(29));
FA_ff_10359:FAff port map(x=>p(247)(29),y=>p(248)(29),Cin=>p(249)(29),clock=>clock,reset=>reset,s=>p(294)(29),cout=>p(295)(30));
FA_ff_10360:FAff port map(x=>p(247)(30),y=>p(248)(30),Cin=>p(249)(30),clock=>clock,reset=>reset,s=>p(294)(30),cout=>p(295)(31));
FA_ff_10361:FAff port map(x=>p(247)(31),y=>p(248)(31),Cin=>p(249)(31),clock=>clock,reset=>reset,s=>p(294)(31),cout=>p(295)(32));
FA_ff_10362:FAff port map(x=>p(247)(32),y=>p(248)(32),Cin=>p(249)(32),clock=>clock,reset=>reset,s=>p(294)(32),cout=>p(295)(33));
FA_ff_10363:FAff port map(x=>p(247)(33),y=>p(248)(33),Cin=>p(249)(33),clock=>clock,reset=>reset,s=>p(294)(33),cout=>p(295)(34));
FA_ff_10364:FAff port map(x=>p(247)(34),y=>p(248)(34),Cin=>p(249)(34),clock=>clock,reset=>reset,s=>p(294)(34),cout=>p(295)(35));
FA_ff_10365:FAff port map(x=>p(247)(35),y=>p(248)(35),Cin=>p(249)(35),clock=>clock,reset=>reset,s=>p(294)(35),cout=>p(295)(36));
FA_ff_10366:FAff port map(x=>p(247)(36),y=>p(248)(36),Cin=>p(249)(36),clock=>clock,reset=>reset,s=>p(294)(36),cout=>p(295)(37));
FA_ff_10367:FAff port map(x=>p(247)(37),y=>p(248)(37),Cin=>p(249)(37),clock=>clock,reset=>reset,s=>p(294)(37),cout=>p(295)(38));
FA_ff_10368:FAff port map(x=>p(247)(38),y=>p(248)(38),Cin=>p(249)(38),clock=>clock,reset=>reset,s=>p(294)(38),cout=>p(295)(39));
FA_ff_10369:FAff port map(x=>p(247)(39),y=>p(248)(39),Cin=>p(249)(39),clock=>clock,reset=>reset,s=>p(294)(39),cout=>p(295)(40));
FA_ff_10370:FAff port map(x=>p(247)(40),y=>p(248)(40),Cin=>p(249)(40),clock=>clock,reset=>reset,s=>p(294)(40),cout=>p(295)(41));
FA_ff_10371:FAff port map(x=>p(247)(41),y=>p(248)(41),Cin=>p(249)(41),clock=>clock,reset=>reset,s=>p(294)(41),cout=>p(295)(42));
FA_ff_10372:FAff port map(x=>p(247)(42),y=>p(248)(42),Cin=>p(249)(42),clock=>clock,reset=>reset,s=>p(294)(42),cout=>p(295)(43));
FA_ff_10373:FAff port map(x=>p(247)(43),y=>p(248)(43),Cin=>p(249)(43),clock=>clock,reset=>reset,s=>p(294)(43),cout=>p(295)(44));
FA_ff_10374:FAff port map(x=>p(247)(44),y=>p(248)(44),Cin=>p(249)(44),clock=>clock,reset=>reset,s=>p(294)(44),cout=>p(295)(45));
FA_ff_10375:FAff port map(x=>p(247)(45),y=>p(248)(45),Cin=>p(249)(45),clock=>clock,reset=>reset,s=>p(294)(45),cout=>p(295)(46));
FA_ff_10376:FAff port map(x=>p(247)(46),y=>p(248)(46),Cin=>p(249)(46),clock=>clock,reset=>reset,s=>p(294)(46),cout=>p(295)(47));
FA_ff_10377:FAff port map(x=>p(247)(47),y=>p(248)(47),Cin=>p(249)(47),clock=>clock,reset=>reset,s=>p(294)(47),cout=>p(295)(48));
FA_ff_10378:FAff port map(x=>p(247)(48),y=>p(248)(48),Cin=>p(249)(48),clock=>clock,reset=>reset,s=>p(294)(48),cout=>p(295)(49));
FA_ff_10379:FAff port map(x=>p(247)(49),y=>p(248)(49),Cin=>p(249)(49),clock=>clock,reset=>reset,s=>p(294)(49),cout=>p(295)(50));
FA_ff_10380:FAff port map(x=>p(247)(50),y=>p(248)(50),Cin=>p(249)(50),clock=>clock,reset=>reset,s=>p(294)(50),cout=>p(295)(51));
FA_ff_10381:FAff port map(x=>p(247)(51),y=>p(248)(51),Cin=>p(249)(51),clock=>clock,reset=>reset,s=>p(294)(51),cout=>p(295)(52));
FA_ff_10382:FAff port map(x=>p(247)(52),y=>p(248)(52),Cin=>p(249)(52),clock=>clock,reset=>reset,s=>p(294)(52),cout=>p(295)(53));
FA_ff_10383:FAff port map(x=>p(247)(53),y=>p(248)(53),Cin=>p(249)(53),clock=>clock,reset=>reset,s=>p(294)(53),cout=>p(295)(54));
FA_ff_10384:FAff port map(x=>p(247)(54),y=>p(248)(54),Cin=>p(249)(54),clock=>clock,reset=>reset,s=>p(294)(54),cout=>p(295)(55));
FA_ff_10385:FAff port map(x=>p(247)(55),y=>p(248)(55),Cin=>p(249)(55),clock=>clock,reset=>reset,s=>p(294)(55),cout=>p(295)(56));
FA_ff_10386:FAff port map(x=>p(247)(56),y=>p(248)(56),Cin=>p(249)(56),clock=>clock,reset=>reset,s=>p(294)(56),cout=>p(295)(57));
FA_ff_10387:FAff port map(x=>p(247)(57),y=>p(248)(57),Cin=>p(249)(57),clock=>clock,reset=>reset,s=>p(294)(57),cout=>p(295)(58));
FA_ff_10388:FAff port map(x=>p(247)(58),y=>p(248)(58),Cin=>p(249)(58),clock=>clock,reset=>reset,s=>p(294)(58),cout=>p(295)(59));
FA_ff_10389:FAff port map(x=>p(247)(59),y=>p(248)(59),Cin=>p(249)(59),clock=>clock,reset=>reset,s=>p(294)(59),cout=>p(295)(60));
FA_ff_10390:FAff port map(x=>p(247)(60),y=>p(248)(60),Cin=>p(249)(60),clock=>clock,reset=>reset,s=>p(294)(60),cout=>p(295)(61));
FA_ff_10391:FAff port map(x=>p(247)(61),y=>p(248)(61),Cin=>p(249)(61),clock=>clock,reset=>reset,s=>p(294)(61),cout=>p(295)(62));
FA_ff_10392:FAff port map(x=>p(247)(62),y=>p(248)(62),Cin=>p(249)(62),clock=>clock,reset=>reset,s=>p(294)(62),cout=>p(295)(63));
FA_ff_10393:FAff port map(x=>p(247)(63),y=>p(248)(63),Cin=>p(249)(63),clock=>clock,reset=>reset,s=>p(294)(63),cout=>p(295)(64));
FA_ff_10394:FAff port map(x=>p(247)(64),y=>p(248)(64),Cin=>p(249)(64),clock=>clock,reset=>reset,s=>p(294)(64),cout=>p(295)(65));
FA_ff_10395:FAff port map(x=>p(247)(65),y=>p(248)(65),Cin=>p(249)(65),clock=>clock,reset=>reset,s=>p(294)(65),cout=>p(295)(66));
FA_ff_10396:FAff port map(x=>p(247)(66),y=>p(248)(66),Cin=>p(249)(66),clock=>clock,reset=>reset,s=>p(294)(66),cout=>p(295)(67));
FA_ff_10397:FAff port map(x=>p(247)(67),y=>p(248)(67),Cin=>p(249)(67),clock=>clock,reset=>reset,s=>p(294)(67),cout=>p(295)(68));
FA_ff_10398:FAff port map(x=>p(247)(68),y=>p(248)(68),Cin=>p(249)(68),clock=>clock,reset=>reset,s=>p(294)(68),cout=>p(295)(69));
FA_ff_10399:FAff port map(x=>p(247)(69),y=>p(248)(69),Cin=>p(249)(69),clock=>clock,reset=>reset,s=>p(294)(69),cout=>p(295)(70));
FA_ff_10400:FAff port map(x=>p(247)(70),y=>p(248)(70),Cin=>p(249)(70),clock=>clock,reset=>reset,s=>p(294)(70),cout=>p(295)(71));
FA_ff_10401:FAff port map(x=>p(247)(71),y=>p(248)(71),Cin=>p(249)(71),clock=>clock,reset=>reset,s=>p(294)(71),cout=>p(295)(72));
FA_ff_10402:FAff port map(x=>p(247)(72),y=>p(248)(72),Cin=>p(249)(72),clock=>clock,reset=>reset,s=>p(294)(72),cout=>p(295)(73));
FA_ff_10403:FAff port map(x=>p(247)(73),y=>p(248)(73),Cin=>p(249)(73),clock=>clock,reset=>reset,s=>p(294)(73),cout=>p(295)(74));
FA_ff_10404:FAff port map(x=>p(247)(74),y=>p(248)(74),Cin=>p(249)(74),clock=>clock,reset=>reset,s=>p(294)(74),cout=>p(295)(75));
FA_ff_10405:FAff port map(x=>p(247)(75),y=>p(248)(75),Cin=>p(249)(75),clock=>clock,reset=>reset,s=>p(294)(75),cout=>p(295)(76));
FA_ff_10406:FAff port map(x=>p(247)(76),y=>p(248)(76),Cin=>p(249)(76),clock=>clock,reset=>reset,s=>p(294)(76),cout=>p(295)(77));
FA_ff_10407:FAff port map(x=>p(247)(77),y=>p(248)(77),Cin=>p(249)(77),clock=>clock,reset=>reset,s=>p(294)(77),cout=>p(295)(78));
FA_ff_10408:FAff port map(x=>p(247)(78),y=>p(248)(78),Cin=>p(249)(78),clock=>clock,reset=>reset,s=>p(294)(78),cout=>p(295)(79));
FA_ff_10409:FAff port map(x=>p(247)(79),y=>p(248)(79),Cin=>p(249)(79),clock=>clock,reset=>reset,s=>p(294)(79),cout=>p(295)(80));
FA_ff_10410:FAff port map(x=>p(247)(80),y=>p(248)(80),Cin=>p(249)(80),clock=>clock,reset=>reset,s=>p(294)(80),cout=>p(295)(81));
FA_ff_10411:FAff port map(x=>p(247)(81),y=>p(248)(81),Cin=>p(249)(81),clock=>clock,reset=>reset,s=>p(294)(81),cout=>p(295)(82));
FA_ff_10412:FAff port map(x=>p(247)(82),y=>p(248)(82),Cin=>p(249)(82),clock=>clock,reset=>reset,s=>p(294)(82),cout=>p(295)(83));
FA_ff_10413:FAff port map(x=>p(247)(83),y=>p(248)(83),Cin=>p(249)(83),clock=>clock,reset=>reset,s=>p(294)(83),cout=>p(295)(84));
FA_ff_10414:FAff port map(x=>p(247)(84),y=>p(248)(84),Cin=>p(249)(84),clock=>clock,reset=>reset,s=>p(294)(84),cout=>p(295)(85));
FA_ff_10415:FAff port map(x=>p(247)(85),y=>p(248)(85),Cin=>p(249)(85),clock=>clock,reset=>reset,s=>p(294)(85),cout=>p(295)(86));
FA_ff_10416:FAff port map(x=>p(247)(86),y=>p(248)(86),Cin=>p(249)(86),clock=>clock,reset=>reset,s=>p(294)(86),cout=>p(295)(87));
FA_ff_10417:FAff port map(x=>p(247)(87),y=>p(248)(87),Cin=>p(249)(87),clock=>clock,reset=>reset,s=>p(294)(87),cout=>p(295)(88));
FA_ff_10418:FAff port map(x=>p(247)(88),y=>p(248)(88),Cin=>p(249)(88),clock=>clock,reset=>reset,s=>p(294)(88),cout=>p(295)(89));
FA_ff_10419:FAff port map(x=>p(247)(89),y=>p(248)(89),Cin=>p(249)(89),clock=>clock,reset=>reset,s=>p(294)(89),cout=>p(295)(90));
FA_ff_10420:FAff port map(x=>p(247)(90),y=>p(248)(90),Cin=>p(249)(90),clock=>clock,reset=>reset,s=>p(294)(90),cout=>p(295)(91));
FA_ff_10421:FAff port map(x=>p(247)(91),y=>p(248)(91),Cin=>p(249)(91),clock=>clock,reset=>reset,s=>p(294)(91),cout=>p(295)(92));
FA_ff_10422:FAff port map(x=>p(247)(92),y=>p(248)(92),Cin=>p(249)(92),clock=>clock,reset=>reset,s=>p(294)(92),cout=>p(295)(93));
FA_ff_10423:FAff port map(x=>p(247)(93),y=>p(248)(93),Cin=>p(249)(93),clock=>clock,reset=>reset,s=>p(294)(93),cout=>p(295)(94));
FA_ff_10424:FAff port map(x=>p(247)(94),y=>p(248)(94),Cin=>p(249)(94),clock=>clock,reset=>reset,s=>p(294)(94),cout=>p(295)(95));
FA_ff_10425:FAff port map(x=>p(247)(95),y=>p(248)(95),Cin=>p(249)(95),clock=>clock,reset=>reset,s=>p(294)(95),cout=>p(295)(96));
FA_ff_10426:FAff port map(x=>p(247)(96),y=>p(248)(96),Cin=>p(249)(96),clock=>clock,reset=>reset,s=>p(294)(96),cout=>p(295)(97));
FA_ff_10427:FAff port map(x=>p(247)(97),y=>p(248)(97),Cin=>p(249)(97),clock=>clock,reset=>reset,s=>p(294)(97),cout=>p(295)(98));
FA_ff_10428:FAff port map(x=>p(247)(98),y=>p(248)(98),Cin=>p(249)(98),clock=>clock,reset=>reset,s=>p(294)(98),cout=>p(295)(99));
FA_ff_10429:FAff port map(x=>p(247)(99),y=>p(248)(99),Cin=>p(249)(99),clock=>clock,reset=>reset,s=>p(294)(99),cout=>p(295)(100));
FA_ff_10430:FAff port map(x=>p(247)(100),y=>p(248)(100),Cin=>p(249)(100),clock=>clock,reset=>reset,s=>p(294)(100),cout=>p(295)(101));
FA_ff_10431:FAff port map(x=>p(247)(101),y=>p(248)(101),Cin=>p(249)(101),clock=>clock,reset=>reset,s=>p(294)(101),cout=>p(295)(102));
FA_ff_10432:FAff port map(x=>p(247)(102),y=>p(248)(102),Cin=>p(249)(102),clock=>clock,reset=>reset,s=>p(294)(102),cout=>p(295)(103));
FA_ff_10433:FAff port map(x=>p(247)(103),y=>p(248)(103),Cin=>p(249)(103),clock=>clock,reset=>reset,s=>p(294)(103),cout=>p(295)(104));
FA_ff_10434:FAff port map(x=>p(247)(104),y=>p(248)(104),Cin=>p(249)(104),clock=>clock,reset=>reset,s=>p(294)(104),cout=>p(295)(105));
FA_ff_10435:FAff port map(x=>p(247)(105),y=>p(248)(105),Cin=>p(249)(105),clock=>clock,reset=>reset,s=>p(294)(105),cout=>p(295)(106));
FA_ff_10436:FAff port map(x=>p(247)(106),y=>p(248)(106),Cin=>p(249)(106),clock=>clock,reset=>reset,s=>p(294)(106),cout=>p(295)(107));
FA_ff_10437:FAff port map(x=>p(247)(107),y=>p(248)(107),Cin=>p(249)(107),clock=>clock,reset=>reset,s=>p(294)(107),cout=>p(295)(108));
FA_ff_10438:FAff port map(x=>p(247)(108),y=>p(248)(108),Cin=>p(249)(108),clock=>clock,reset=>reset,s=>p(294)(108),cout=>p(295)(109));
FA_ff_10439:FAff port map(x=>p(247)(109),y=>p(248)(109),Cin=>p(249)(109),clock=>clock,reset=>reset,s=>p(294)(109),cout=>p(295)(110));
FA_ff_10440:FAff port map(x=>p(247)(110),y=>p(248)(110),Cin=>p(249)(110),clock=>clock,reset=>reset,s=>p(294)(110),cout=>p(295)(111));
FA_ff_10441:FAff port map(x=>p(247)(111),y=>p(248)(111),Cin=>p(249)(111),clock=>clock,reset=>reset,s=>p(294)(111),cout=>p(295)(112));
FA_ff_10442:FAff port map(x=>p(247)(112),y=>p(248)(112),Cin=>p(249)(112),clock=>clock,reset=>reset,s=>p(294)(112),cout=>p(295)(113));
FA_ff_10443:FAff port map(x=>p(247)(113),y=>p(248)(113),Cin=>p(249)(113),clock=>clock,reset=>reset,s=>p(294)(113),cout=>p(295)(114));
FA_ff_10444:FAff port map(x=>p(247)(114),y=>p(248)(114),Cin=>p(249)(114),clock=>clock,reset=>reset,s=>p(294)(114),cout=>p(295)(115));
FA_ff_10445:FAff port map(x=>p(247)(115),y=>p(248)(115),Cin=>p(249)(115),clock=>clock,reset=>reset,s=>p(294)(115),cout=>p(295)(116));
FA_ff_10446:FAff port map(x=>p(247)(116),y=>p(248)(116),Cin=>p(249)(116),clock=>clock,reset=>reset,s=>p(294)(116),cout=>p(295)(117));
FA_ff_10447:FAff port map(x=>p(247)(117),y=>p(248)(117),Cin=>p(249)(117),clock=>clock,reset=>reset,s=>p(294)(117),cout=>p(295)(118));
FA_ff_10448:FAff port map(x=>p(247)(118),y=>p(248)(118),Cin=>p(249)(118),clock=>clock,reset=>reset,s=>p(294)(118),cout=>p(295)(119));
FA_ff_10449:FAff port map(x=>p(247)(119),y=>p(248)(119),Cin=>p(249)(119),clock=>clock,reset=>reset,s=>p(294)(119),cout=>p(295)(120));
FA_ff_10450:FAff port map(x=>p(247)(120),y=>p(248)(120),Cin=>p(249)(120),clock=>clock,reset=>reset,s=>p(294)(120),cout=>p(295)(121));
FA_ff_10451:FAff port map(x=>p(247)(121),y=>p(248)(121),Cin=>p(249)(121),clock=>clock,reset=>reset,s=>p(294)(121),cout=>p(295)(122));
FA_ff_10452:FAff port map(x=>p(247)(122),y=>p(248)(122),Cin=>p(249)(122),clock=>clock,reset=>reset,s=>p(294)(122),cout=>p(295)(123));
FA_ff_10453:FAff port map(x=>p(247)(123),y=>p(248)(123),Cin=>p(249)(123),clock=>clock,reset=>reset,s=>p(294)(123),cout=>p(295)(124));
FA_ff_10454:FAff port map(x=>p(247)(124),y=>p(248)(124),Cin=>p(249)(124),clock=>clock,reset=>reset,s=>p(294)(124),cout=>p(295)(125));
FA_ff_10455:FAff port map(x=>p(247)(125),y=>p(248)(125),Cin=>p(249)(125),clock=>clock,reset=>reset,s=>p(294)(125),cout=>p(295)(126));
FA_ff_10456:FAff port map(x=>p(247)(126),y=>p(248)(126),Cin=>p(249)(126),clock=>clock,reset=>reset,s=>p(294)(126),cout=>p(295)(127));
FA_ff_10457:FAff port map(x=>p(247)(127),y=>p(248)(127),Cin=>p(249)(127),clock=>clock,reset=>reset,s=>p(294)(127),cout=>p(295)(128));
FA_ff_10458:FAff port map(x=>p(247)(128),y=>p(248)(128),Cin=>p(249)(128),clock=>clock,reset=>reset,s=>p(294)(128),cout=>p(295)(129));
p(294)(129)<=p(249)(129);
HA_ff_43:HAff port map(x=>p(250)(0),y=>p(252)(0),clock=>clock,reset=>reset,s=>p(296)(0),c=>p(297)(1));
FA_ff_10459:FAff port map(x=>p(250)(1),y=>p(251)(1),Cin=>p(252)(1),clock=>clock,reset=>reset,s=>p(296)(1),cout=>p(297)(2));
FA_ff_10460:FAff port map(x=>p(250)(2),y=>p(251)(2),Cin=>p(252)(2),clock=>clock,reset=>reset,s=>p(296)(2),cout=>p(297)(3));
FA_ff_10461:FAff port map(x=>p(250)(3),y=>p(251)(3),Cin=>p(252)(3),clock=>clock,reset=>reset,s=>p(296)(3),cout=>p(297)(4));
FA_ff_10462:FAff port map(x=>p(250)(4),y=>p(251)(4),Cin=>p(252)(4),clock=>clock,reset=>reset,s=>p(296)(4),cout=>p(297)(5));
FA_ff_10463:FAff port map(x=>p(250)(5),y=>p(251)(5),Cin=>p(252)(5),clock=>clock,reset=>reset,s=>p(296)(5),cout=>p(297)(6));
FA_ff_10464:FAff port map(x=>p(250)(6),y=>p(251)(6),Cin=>p(252)(6),clock=>clock,reset=>reset,s=>p(296)(6),cout=>p(297)(7));
FA_ff_10465:FAff port map(x=>p(250)(7),y=>p(251)(7),Cin=>p(252)(7),clock=>clock,reset=>reset,s=>p(296)(7),cout=>p(297)(8));
FA_ff_10466:FAff port map(x=>p(250)(8),y=>p(251)(8),Cin=>p(252)(8),clock=>clock,reset=>reset,s=>p(296)(8),cout=>p(297)(9));
FA_ff_10467:FAff port map(x=>p(250)(9),y=>p(251)(9),Cin=>p(252)(9),clock=>clock,reset=>reset,s=>p(296)(9),cout=>p(297)(10));
FA_ff_10468:FAff port map(x=>p(250)(10),y=>p(251)(10),Cin=>p(252)(10),clock=>clock,reset=>reset,s=>p(296)(10),cout=>p(297)(11));
FA_ff_10469:FAff port map(x=>p(250)(11),y=>p(251)(11),Cin=>p(252)(11),clock=>clock,reset=>reset,s=>p(296)(11),cout=>p(297)(12));
FA_ff_10470:FAff port map(x=>p(250)(12),y=>p(251)(12),Cin=>p(252)(12),clock=>clock,reset=>reset,s=>p(296)(12),cout=>p(297)(13));
FA_ff_10471:FAff port map(x=>p(250)(13),y=>p(251)(13),Cin=>p(252)(13),clock=>clock,reset=>reset,s=>p(296)(13),cout=>p(297)(14));
FA_ff_10472:FAff port map(x=>p(250)(14),y=>p(251)(14),Cin=>p(252)(14),clock=>clock,reset=>reset,s=>p(296)(14),cout=>p(297)(15));
FA_ff_10473:FAff port map(x=>p(250)(15),y=>p(251)(15),Cin=>p(252)(15),clock=>clock,reset=>reset,s=>p(296)(15),cout=>p(297)(16));
FA_ff_10474:FAff port map(x=>p(250)(16),y=>p(251)(16),Cin=>p(252)(16),clock=>clock,reset=>reset,s=>p(296)(16),cout=>p(297)(17));
FA_ff_10475:FAff port map(x=>p(250)(17),y=>p(251)(17),Cin=>p(252)(17),clock=>clock,reset=>reset,s=>p(296)(17),cout=>p(297)(18));
FA_ff_10476:FAff port map(x=>p(250)(18),y=>p(251)(18),Cin=>p(252)(18),clock=>clock,reset=>reset,s=>p(296)(18),cout=>p(297)(19));
FA_ff_10477:FAff port map(x=>p(250)(19),y=>p(251)(19),Cin=>p(252)(19),clock=>clock,reset=>reset,s=>p(296)(19),cout=>p(297)(20));
FA_ff_10478:FAff port map(x=>p(250)(20),y=>p(251)(20),Cin=>p(252)(20),clock=>clock,reset=>reset,s=>p(296)(20),cout=>p(297)(21));
FA_ff_10479:FAff port map(x=>p(250)(21),y=>p(251)(21),Cin=>p(252)(21),clock=>clock,reset=>reset,s=>p(296)(21),cout=>p(297)(22));
FA_ff_10480:FAff port map(x=>p(250)(22),y=>p(251)(22),Cin=>p(252)(22),clock=>clock,reset=>reset,s=>p(296)(22),cout=>p(297)(23));
FA_ff_10481:FAff port map(x=>p(250)(23),y=>p(251)(23),Cin=>p(252)(23),clock=>clock,reset=>reset,s=>p(296)(23),cout=>p(297)(24));
FA_ff_10482:FAff port map(x=>p(250)(24),y=>p(251)(24),Cin=>p(252)(24),clock=>clock,reset=>reset,s=>p(296)(24),cout=>p(297)(25));
FA_ff_10483:FAff port map(x=>p(250)(25),y=>p(251)(25),Cin=>p(252)(25),clock=>clock,reset=>reset,s=>p(296)(25),cout=>p(297)(26));
FA_ff_10484:FAff port map(x=>p(250)(26),y=>p(251)(26),Cin=>p(252)(26),clock=>clock,reset=>reset,s=>p(296)(26),cout=>p(297)(27));
FA_ff_10485:FAff port map(x=>p(250)(27),y=>p(251)(27),Cin=>p(252)(27),clock=>clock,reset=>reset,s=>p(296)(27),cout=>p(297)(28));
FA_ff_10486:FAff port map(x=>p(250)(28),y=>p(251)(28),Cin=>p(252)(28),clock=>clock,reset=>reset,s=>p(296)(28),cout=>p(297)(29));
FA_ff_10487:FAff port map(x=>p(250)(29),y=>p(251)(29),Cin=>p(252)(29),clock=>clock,reset=>reset,s=>p(296)(29),cout=>p(297)(30));
FA_ff_10488:FAff port map(x=>p(250)(30),y=>p(251)(30),Cin=>p(252)(30),clock=>clock,reset=>reset,s=>p(296)(30),cout=>p(297)(31));
FA_ff_10489:FAff port map(x=>p(250)(31),y=>p(251)(31),Cin=>p(252)(31),clock=>clock,reset=>reset,s=>p(296)(31),cout=>p(297)(32));
FA_ff_10490:FAff port map(x=>p(250)(32),y=>p(251)(32),Cin=>p(252)(32),clock=>clock,reset=>reset,s=>p(296)(32),cout=>p(297)(33));
FA_ff_10491:FAff port map(x=>p(250)(33),y=>p(251)(33),Cin=>p(252)(33),clock=>clock,reset=>reset,s=>p(296)(33),cout=>p(297)(34));
FA_ff_10492:FAff port map(x=>p(250)(34),y=>p(251)(34),Cin=>p(252)(34),clock=>clock,reset=>reset,s=>p(296)(34),cout=>p(297)(35));
FA_ff_10493:FAff port map(x=>p(250)(35),y=>p(251)(35),Cin=>p(252)(35),clock=>clock,reset=>reset,s=>p(296)(35),cout=>p(297)(36));
FA_ff_10494:FAff port map(x=>p(250)(36),y=>p(251)(36),Cin=>p(252)(36),clock=>clock,reset=>reset,s=>p(296)(36),cout=>p(297)(37));
FA_ff_10495:FAff port map(x=>p(250)(37),y=>p(251)(37),Cin=>p(252)(37),clock=>clock,reset=>reset,s=>p(296)(37),cout=>p(297)(38));
FA_ff_10496:FAff port map(x=>p(250)(38),y=>p(251)(38),Cin=>p(252)(38),clock=>clock,reset=>reset,s=>p(296)(38),cout=>p(297)(39));
FA_ff_10497:FAff port map(x=>p(250)(39),y=>p(251)(39),Cin=>p(252)(39),clock=>clock,reset=>reset,s=>p(296)(39),cout=>p(297)(40));
FA_ff_10498:FAff port map(x=>p(250)(40),y=>p(251)(40),Cin=>p(252)(40),clock=>clock,reset=>reset,s=>p(296)(40),cout=>p(297)(41));
FA_ff_10499:FAff port map(x=>p(250)(41),y=>p(251)(41),Cin=>p(252)(41),clock=>clock,reset=>reset,s=>p(296)(41),cout=>p(297)(42));
FA_ff_10500:FAff port map(x=>p(250)(42),y=>p(251)(42),Cin=>p(252)(42),clock=>clock,reset=>reset,s=>p(296)(42),cout=>p(297)(43));
FA_ff_10501:FAff port map(x=>p(250)(43),y=>p(251)(43),Cin=>p(252)(43),clock=>clock,reset=>reset,s=>p(296)(43),cout=>p(297)(44));
FA_ff_10502:FAff port map(x=>p(250)(44),y=>p(251)(44),Cin=>p(252)(44),clock=>clock,reset=>reset,s=>p(296)(44),cout=>p(297)(45));
FA_ff_10503:FAff port map(x=>p(250)(45),y=>p(251)(45),Cin=>p(252)(45),clock=>clock,reset=>reset,s=>p(296)(45),cout=>p(297)(46));
FA_ff_10504:FAff port map(x=>p(250)(46),y=>p(251)(46),Cin=>p(252)(46),clock=>clock,reset=>reset,s=>p(296)(46),cout=>p(297)(47));
FA_ff_10505:FAff port map(x=>p(250)(47),y=>p(251)(47),Cin=>p(252)(47),clock=>clock,reset=>reset,s=>p(296)(47),cout=>p(297)(48));
FA_ff_10506:FAff port map(x=>p(250)(48),y=>p(251)(48),Cin=>p(252)(48),clock=>clock,reset=>reset,s=>p(296)(48),cout=>p(297)(49));
FA_ff_10507:FAff port map(x=>p(250)(49),y=>p(251)(49),Cin=>p(252)(49),clock=>clock,reset=>reset,s=>p(296)(49),cout=>p(297)(50));
FA_ff_10508:FAff port map(x=>p(250)(50),y=>p(251)(50),Cin=>p(252)(50),clock=>clock,reset=>reset,s=>p(296)(50),cout=>p(297)(51));
FA_ff_10509:FAff port map(x=>p(250)(51),y=>p(251)(51),Cin=>p(252)(51),clock=>clock,reset=>reset,s=>p(296)(51),cout=>p(297)(52));
FA_ff_10510:FAff port map(x=>p(250)(52),y=>p(251)(52),Cin=>p(252)(52),clock=>clock,reset=>reset,s=>p(296)(52),cout=>p(297)(53));
FA_ff_10511:FAff port map(x=>p(250)(53),y=>p(251)(53),Cin=>p(252)(53),clock=>clock,reset=>reset,s=>p(296)(53),cout=>p(297)(54));
FA_ff_10512:FAff port map(x=>p(250)(54),y=>p(251)(54),Cin=>p(252)(54),clock=>clock,reset=>reset,s=>p(296)(54),cout=>p(297)(55));
FA_ff_10513:FAff port map(x=>p(250)(55),y=>p(251)(55),Cin=>p(252)(55),clock=>clock,reset=>reset,s=>p(296)(55),cout=>p(297)(56));
FA_ff_10514:FAff port map(x=>p(250)(56),y=>p(251)(56),Cin=>p(252)(56),clock=>clock,reset=>reset,s=>p(296)(56),cout=>p(297)(57));
FA_ff_10515:FAff port map(x=>p(250)(57),y=>p(251)(57),Cin=>p(252)(57),clock=>clock,reset=>reset,s=>p(296)(57),cout=>p(297)(58));
FA_ff_10516:FAff port map(x=>p(250)(58),y=>p(251)(58),Cin=>p(252)(58),clock=>clock,reset=>reset,s=>p(296)(58),cout=>p(297)(59));
FA_ff_10517:FAff port map(x=>p(250)(59),y=>p(251)(59),Cin=>p(252)(59),clock=>clock,reset=>reset,s=>p(296)(59),cout=>p(297)(60));
FA_ff_10518:FAff port map(x=>p(250)(60),y=>p(251)(60),Cin=>p(252)(60),clock=>clock,reset=>reset,s=>p(296)(60),cout=>p(297)(61));
FA_ff_10519:FAff port map(x=>p(250)(61),y=>p(251)(61),Cin=>p(252)(61),clock=>clock,reset=>reset,s=>p(296)(61),cout=>p(297)(62));
FA_ff_10520:FAff port map(x=>p(250)(62),y=>p(251)(62),Cin=>p(252)(62),clock=>clock,reset=>reset,s=>p(296)(62),cout=>p(297)(63));
FA_ff_10521:FAff port map(x=>p(250)(63),y=>p(251)(63),Cin=>p(252)(63),clock=>clock,reset=>reset,s=>p(296)(63),cout=>p(297)(64));
FA_ff_10522:FAff port map(x=>p(250)(64),y=>p(251)(64),Cin=>p(252)(64),clock=>clock,reset=>reset,s=>p(296)(64),cout=>p(297)(65));
FA_ff_10523:FAff port map(x=>p(250)(65),y=>p(251)(65),Cin=>p(252)(65),clock=>clock,reset=>reset,s=>p(296)(65),cout=>p(297)(66));
FA_ff_10524:FAff port map(x=>p(250)(66),y=>p(251)(66),Cin=>p(252)(66),clock=>clock,reset=>reset,s=>p(296)(66),cout=>p(297)(67));
FA_ff_10525:FAff port map(x=>p(250)(67),y=>p(251)(67),Cin=>p(252)(67),clock=>clock,reset=>reset,s=>p(296)(67),cout=>p(297)(68));
FA_ff_10526:FAff port map(x=>p(250)(68),y=>p(251)(68),Cin=>p(252)(68),clock=>clock,reset=>reset,s=>p(296)(68),cout=>p(297)(69));
FA_ff_10527:FAff port map(x=>p(250)(69),y=>p(251)(69),Cin=>p(252)(69),clock=>clock,reset=>reset,s=>p(296)(69),cout=>p(297)(70));
FA_ff_10528:FAff port map(x=>p(250)(70),y=>p(251)(70),Cin=>p(252)(70),clock=>clock,reset=>reset,s=>p(296)(70),cout=>p(297)(71));
FA_ff_10529:FAff port map(x=>p(250)(71),y=>p(251)(71),Cin=>p(252)(71),clock=>clock,reset=>reset,s=>p(296)(71),cout=>p(297)(72));
FA_ff_10530:FAff port map(x=>p(250)(72),y=>p(251)(72),Cin=>p(252)(72),clock=>clock,reset=>reset,s=>p(296)(72),cout=>p(297)(73));
FA_ff_10531:FAff port map(x=>p(250)(73),y=>p(251)(73),Cin=>p(252)(73),clock=>clock,reset=>reset,s=>p(296)(73),cout=>p(297)(74));
FA_ff_10532:FAff port map(x=>p(250)(74),y=>p(251)(74),Cin=>p(252)(74),clock=>clock,reset=>reset,s=>p(296)(74),cout=>p(297)(75));
FA_ff_10533:FAff port map(x=>p(250)(75),y=>p(251)(75),Cin=>p(252)(75),clock=>clock,reset=>reset,s=>p(296)(75),cout=>p(297)(76));
FA_ff_10534:FAff port map(x=>p(250)(76),y=>p(251)(76),Cin=>p(252)(76),clock=>clock,reset=>reset,s=>p(296)(76),cout=>p(297)(77));
FA_ff_10535:FAff port map(x=>p(250)(77),y=>p(251)(77),Cin=>p(252)(77),clock=>clock,reset=>reset,s=>p(296)(77),cout=>p(297)(78));
FA_ff_10536:FAff port map(x=>p(250)(78),y=>p(251)(78),Cin=>p(252)(78),clock=>clock,reset=>reset,s=>p(296)(78),cout=>p(297)(79));
FA_ff_10537:FAff port map(x=>p(250)(79),y=>p(251)(79),Cin=>p(252)(79),clock=>clock,reset=>reset,s=>p(296)(79),cout=>p(297)(80));
FA_ff_10538:FAff port map(x=>p(250)(80),y=>p(251)(80),Cin=>p(252)(80),clock=>clock,reset=>reset,s=>p(296)(80),cout=>p(297)(81));
FA_ff_10539:FAff port map(x=>p(250)(81),y=>p(251)(81),Cin=>p(252)(81),clock=>clock,reset=>reset,s=>p(296)(81),cout=>p(297)(82));
FA_ff_10540:FAff port map(x=>p(250)(82),y=>p(251)(82),Cin=>p(252)(82),clock=>clock,reset=>reset,s=>p(296)(82),cout=>p(297)(83));
FA_ff_10541:FAff port map(x=>p(250)(83),y=>p(251)(83),Cin=>p(252)(83),clock=>clock,reset=>reset,s=>p(296)(83),cout=>p(297)(84));
FA_ff_10542:FAff port map(x=>p(250)(84),y=>p(251)(84),Cin=>p(252)(84),clock=>clock,reset=>reset,s=>p(296)(84),cout=>p(297)(85));
FA_ff_10543:FAff port map(x=>p(250)(85),y=>p(251)(85),Cin=>p(252)(85),clock=>clock,reset=>reset,s=>p(296)(85),cout=>p(297)(86));
FA_ff_10544:FAff port map(x=>p(250)(86),y=>p(251)(86),Cin=>p(252)(86),clock=>clock,reset=>reset,s=>p(296)(86),cout=>p(297)(87));
FA_ff_10545:FAff port map(x=>p(250)(87),y=>p(251)(87),Cin=>p(252)(87),clock=>clock,reset=>reset,s=>p(296)(87),cout=>p(297)(88));
FA_ff_10546:FAff port map(x=>p(250)(88),y=>p(251)(88),Cin=>p(252)(88),clock=>clock,reset=>reset,s=>p(296)(88),cout=>p(297)(89));
FA_ff_10547:FAff port map(x=>p(250)(89),y=>p(251)(89),Cin=>p(252)(89),clock=>clock,reset=>reset,s=>p(296)(89),cout=>p(297)(90));
FA_ff_10548:FAff port map(x=>p(250)(90),y=>p(251)(90),Cin=>p(252)(90),clock=>clock,reset=>reset,s=>p(296)(90),cout=>p(297)(91));
FA_ff_10549:FAff port map(x=>p(250)(91),y=>p(251)(91),Cin=>p(252)(91),clock=>clock,reset=>reset,s=>p(296)(91),cout=>p(297)(92));
FA_ff_10550:FAff port map(x=>p(250)(92),y=>p(251)(92),Cin=>p(252)(92),clock=>clock,reset=>reset,s=>p(296)(92),cout=>p(297)(93));
FA_ff_10551:FAff port map(x=>p(250)(93),y=>p(251)(93),Cin=>p(252)(93),clock=>clock,reset=>reset,s=>p(296)(93),cout=>p(297)(94));
FA_ff_10552:FAff port map(x=>p(250)(94),y=>p(251)(94),Cin=>p(252)(94),clock=>clock,reset=>reset,s=>p(296)(94),cout=>p(297)(95));
FA_ff_10553:FAff port map(x=>p(250)(95),y=>p(251)(95),Cin=>p(252)(95),clock=>clock,reset=>reset,s=>p(296)(95),cout=>p(297)(96));
FA_ff_10554:FAff port map(x=>p(250)(96),y=>p(251)(96),Cin=>p(252)(96),clock=>clock,reset=>reset,s=>p(296)(96),cout=>p(297)(97));
FA_ff_10555:FAff port map(x=>p(250)(97),y=>p(251)(97),Cin=>p(252)(97),clock=>clock,reset=>reset,s=>p(296)(97),cout=>p(297)(98));
FA_ff_10556:FAff port map(x=>p(250)(98),y=>p(251)(98),Cin=>p(252)(98),clock=>clock,reset=>reset,s=>p(296)(98),cout=>p(297)(99));
FA_ff_10557:FAff port map(x=>p(250)(99),y=>p(251)(99),Cin=>p(252)(99),clock=>clock,reset=>reset,s=>p(296)(99),cout=>p(297)(100));
FA_ff_10558:FAff port map(x=>p(250)(100),y=>p(251)(100),Cin=>p(252)(100),clock=>clock,reset=>reset,s=>p(296)(100),cout=>p(297)(101));
FA_ff_10559:FAff port map(x=>p(250)(101),y=>p(251)(101),Cin=>p(252)(101),clock=>clock,reset=>reset,s=>p(296)(101),cout=>p(297)(102));
FA_ff_10560:FAff port map(x=>p(250)(102),y=>p(251)(102),Cin=>p(252)(102),clock=>clock,reset=>reset,s=>p(296)(102),cout=>p(297)(103));
FA_ff_10561:FAff port map(x=>p(250)(103),y=>p(251)(103),Cin=>p(252)(103),clock=>clock,reset=>reset,s=>p(296)(103),cout=>p(297)(104));
FA_ff_10562:FAff port map(x=>p(250)(104),y=>p(251)(104),Cin=>p(252)(104),clock=>clock,reset=>reset,s=>p(296)(104),cout=>p(297)(105));
FA_ff_10563:FAff port map(x=>p(250)(105),y=>p(251)(105),Cin=>p(252)(105),clock=>clock,reset=>reset,s=>p(296)(105),cout=>p(297)(106));
FA_ff_10564:FAff port map(x=>p(250)(106),y=>p(251)(106),Cin=>p(252)(106),clock=>clock,reset=>reset,s=>p(296)(106),cout=>p(297)(107));
FA_ff_10565:FAff port map(x=>p(250)(107),y=>p(251)(107),Cin=>p(252)(107),clock=>clock,reset=>reset,s=>p(296)(107),cout=>p(297)(108));
FA_ff_10566:FAff port map(x=>p(250)(108),y=>p(251)(108),Cin=>p(252)(108),clock=>clock,reset=>reset,s=>p(296)(108),cout=>p(297)(109));
FA_ff_10567:FAff port map(x=>p(250)(109),y=>p(251)(109),Cin=>p(252)(109),clock=>clock,reset=>reset,s=>p(296)(109),cout=>p(297)(110));
FA_ff_10568:FAff port map(x=>p(250)(110),y=>p(251)(110),Cin=>p(252)(110),clock=>clock,reset=>reset,s=>p(296)(110),cout=>p(297)(111));
FA_ff_10569:FAff port map(x=>p(250)(111),y=>p(251)(111),Cin=>p(252)(111),clock=>clock,reset=>reset,s=>p(296)(111),cout=>p(297)(112));
FA_ff_10570:FAff port map(x=>p(250)(112),y=>p(251)(112),Cin=>p(252)(112),clock=>clock,reset=>reset,s=>p(296)(112),cout=>p(297)(113));
FA_ff_10571:FAff port map(x=>p(250)(113),y=>p(251)(113),Cin=>p(252)(113),clock=>clock,reset=>reset,s=>p(296)(113),cout=>p(297)(114));
FA_ff_10572:FAff port map(x=>p(250)(114),y=>p(251)(114),Cin=>p(252)(114),clock=>clock,reset=>reset,s=>p(296)(114),cout=>p(297)(115));
FA_ff_10573:FAff port map(x=>p(250)(115),y=>p(251)(115),Cin=>p(252)(115),clock=>clock,reset=>reset,s=>p(296)(115),cout=>p(297)(116));
FA_ff_10574:FAff port map(x=>p(250)(116),y=>p(251)(116),Cin=>p(252)(116),clock=>clock,reset=>reset,s=>p(296)(116),cout=>p(297)(117));
FA_ff_10575:FAff port map(x=>p(250)(117),y=>p(251)(117),Cin=>p(252)(117),clock=>clock,reset=>reset,s=>p(296)(117),cout=>p(297)(118));
FA_ff_10576:FAff port map(x=>p(250)(118),y=>p(251)(118),Cin=>p(252)(118),clock=>clock,reset=>reset,s=>p(296)(118),cout=>p(297)(119));
FA_ff_10577:FAff port map(x=>p(250)(119),y=>p(251)(119),Cin=>p(252)(119),clock=>clock,reset=>reset,s=>p(296)(119),cout=>p(297)(120));
FA_ff_10578:FAff port map(x=>p(250)(120),y=>p(251)(120),Cin=>p(252)(120),clock=>clock,reset=>reset,s=>p(296)(120),cout=>p(297)(121));
FA_ff_10579:FAff port map(x=>p(250)(121),y=>p(251)(121),Cin=>p(252)(121),clock=>clock,reset=>reset,s=>p(296)(121),cout=>p(297)(122));
FA_ff_10580:FAff port map(x=>p(250)(122),y=>p(251)(122),Cin=>p(252)(122),clock=>clock,reset=>reset,s=>p(296)(122),cout=>p(297)(123));
FA_ff_10581:FAff port map(x=>p(250)(123),y=>p(251)(123),Cin=>p(252)(123),clock=>clock,reset=>reset,s=>p(296)(123),cout=>p(297)(124));
FA_ff_10582:FAff port map(x=>p(250)(124),y=>p(251)(124),Cin=>p(252)(124),clock=>clock,reset=>reset,s=>p(296)(124),cout=>p(297)(125));
FA_ff_10583:FAff port map(x=>p(250)(125),y=>p(251)(125),Cin=>p(252)(125),clock=>clock,reset=>reset,s=>p(296)(125),cout=>p(297)(126));
FA_ff_10584:FAff port map(x=>p(250)(126),y=>p(251)(126),Cin=>p(252)(126),clock=>clock,reset=>reset,s=>p(296)(126),cout=>p(297)(127));
FA_ff_10585:FAff port map(x=>p(250)(127),y=>p(251)(127),Cin=>p(252)(127),clock=>clock,reset=>reset,s=>p(296)(127),cout=>p(297)(128));
FA_ff_10586:FAff port map(x=>p(250)(128),y=>p(251)(128),Cin=>p(252)(128),clock=>clock,reset=>reset,s=>p(296)(128),cout=>p(297)(129));
p(298)(0)<=p(254)(0);
HA_ff_44:HAff port map(x=>p(254)(1),y=>p(255)(1),clock=>clock,reset=>reset,s=>p(298)(1),c=>p(299)(2));
FA_ff_10587:FAff port map(x=>p(253)(2),y=>p(254)(2),Cin=>p(255)(2),clock=>clock,reset=>reset,s=>p(298)(2),cout=>p(299)(3));
FA_ff_10588:FAff port map(x=>p(253)(3),y=>p(254)(3),Cin=>p(255)(3),clock=>clock,reset=>reset,s=>p(298)(3),cout=>p(299)(4));
FA_ff_10589:FAff port map(x=>p(253)(4),y=>p(254)(4),Cin=>p(255)(4),clock=>clock,reset=>reset,s=>p(298)(4),cout=>p(299)(5));
FA_ff_10590:FAff port map(x=>p(253)(5),y=>p(254)(5),Cin=>p(255)(5),clock=>clock,reset=>reset,s=>p(298)(5),cout=>p(299)(6));
FA_ff_10591:FAff port map(x=>p(253)(6),y=>p(254)(6),Cin=>p(255)(6),clock=>clock,reset=>reset,s=>p(298)(6),cout=>p(299)(7));
FA_ff_10592:FAff port map(x=>p(253)(7),y=>p(254)(7),Cin=>p(255)(7),clock=>clock,reset=>reset,s=>p(298)(7),cout=>p(299)(8));
FA_ff_10593:FAff port map(x=>p(253)(8),y=>p(254)(8),Cin=>p(255)(8),clock=>clock,reset=>reset,s=>p(298)(8),cout=>p(299)(9));
FA_ff_10594:FAff port map(x=>p(253)(9),y=>p(254)(9),Cin=>p(255)(9),clock=>clock,reset=>reset,s=>p(298)(9),cout=>p(299)(10));
FA_ff_10595:FAff port map(x=>p(253)(10),y=>p(254)(10),Cin=>p(255)(10),clock=>clock,reset=>reset,s=>p(298)(10),cout=>p(299)(11));
FA_ff_10596:FAff port map(x=>p(253)(11),y=>p(254)(11),Cin=>p(255)(11),clock=>clock,reset=>reset,s=>p(298)(11),cout=>p(299)(12));
FA_ff_10597:FAff port map(x=>p(253)(12),y=>p(254)(12),Cin=>p(255)(12),clock=>clock,reset=>reset,s=>p(298)(12),cout=>p(299)(13));
FA_ff_10598:FAff port map(x=>p(253)(13),y=>p(254)(13),Cin=>p(255)(13),clock=>clock,reset=>reset,s=>p(298)(13),cout=>p(299)(14));
FA_ff_10599:FAff port map(x=>p(253)(14),y=>p(254)(14),Cin=>p(255)(14),clock=>clock,reset=>reset,s=>p(298)(14),cout=>p(299)(15));
FA_ff_10600:FAff port map(x=>p(253)(15),y=>p(254)(15),Cin=>p(255)(15),clock=>clock,reset=>reset,s=>p(298)(15),cout=>p(299)(16));
FA_ff_10601:FAff port map(x=>p(253)(16),y=>p(254)(16),Cin=>p(255)(16),clock=>clock,reset=>reset,s=>p(298)(16),cout=>p(299)(17));
FA_ff_10602:FAff port map(x=>p(253)(17),y=>p(254)(17),Cin=>p(255)(17),clock=>clock,reset=>reset,s=>p(298)(17),cout=>p(299)(18));
FA_ff_10603:FAff port map(x=>p(253)(18),y=>p(254)(18),Cin=>p(255)(18),clock=>clock,reset=>reset,s=>p(298)(18),cout=>p(299)(19));
FA_ff_10604:FAff port map(x=>p(253)(19),y=>p(254)(19),Cin=>p(255)(19),clock=>clock,reset=>reset,s=>p(298)(19),cout=>p(299)(20));
FA_ff_10605:FAff port map(x=>p(253)(20),y=>p(254)(20),Cin=>p(255)(20),clock=>clock,reset=>reset,s=>p(298)(20),cout=>p(299)(21));
FA_ff_10606:FAff port map(x=>p(253)(21),y=>p(254)(21),Cin=>p(255)(21),clock=>clock,reset=>reset,s=>p(298)(21),cout=>p(299)(22));
FA_ff_10607:FAff port map(x=>p(253)(22),y=>p(254)(22),Cin=>p(255)(22),clock=>clock,reset=>reset,s=>p(298)(22),cout=>p(299)(23));
FA_ff_10608:FAff port map(x=>p(253)(23),y=>p(254)(23),Cin=>p(255)(23),clock=>clock,reset=>reset,s=>p(298)(23),cout=>p(299)(24));
FA_ff_10609:FAff port map(x=>p(253)(24),y=>p(254)(24),Cin=>p(255)(24),clock=>clock,reset=>reset,s=>p(298)(24),cout=>p(299)(25));
FA_ff_10610:FAff port map(x=>p(253)(25),y=>p(254)(25),Cin=>p(255)(25),clock=>clock,reset=>reset,s=>p(298)(25),cout=>p(299)(26));
FA_ff_10611:FAff port map(x=>p(253)(26),y=>p(254)(26),Cin=>p(255)(26),clock=>clock,reset=>reset,s=>p(298)(26),cout=>p(299)(27));
FA_ff_10612:FAff port map(x=>p(253)(27),y=>p(254)(27),Cin=>p(255)(27),clock=>clock,reset=>reset,s=>p(298)(27),cout=>p(299)(28));
FA_ff_10613:FAff port map(x=>p(253)(28),y=>p(254)(28),Cin=>p(255)(28),clock=>clock,reset=>reset,s=>p(298)(28),cout=>p(299)(29));
FA_ff_10614:FAff port map(x=>p(253)(29),y=>p(254)(29),Cin=>p(255)(29),clock=>clock,reset=>reset,s=>p(298)(29),cout=>p(299)(30));
FA_ff_10615:FAff port map(x=>p(253)(30),y=>p(254)(30),Cin=>p(255)(30),clock=>clock,reset=>reset,s=>p(298)(30),cout=>p(299)(31));
FA_ff_10616:FAff port map(x=>p(253)(31),y=>p(254)(31),Cin=>p(255)(31),clock=>clock,reset=>reset,s=>p(298)(31),cout=>p(299)(32));
FA_ff_10617:FAff port map(x=>p(253)(32),y=>p(254)(32),Cin=>p(255)(32),clock=>clock,reset=>reset,s=>p(298)(32),cout=>p(299)(33));
FA_ff_10618:FAff port map(x=>p(253)(33),y=>p(254)(33),Cin=>p(255)(33),clock=>clock,reset=>reset,s=>p(298)(33),cout=>p(299)(34));
FA_ff_10619:FAff port map(x=>p(253)(34),y=>p(254)(34),Cin=>p(255)(34),clock=>clock,reset=>reset,s=>p(298)(34),cout=>p(299)(35));
FA_ff_10620:FAff port map(x=>p(253)(35),y=>p(254)(35),Cin=>p(255)(35),clock=>clock,reset=>reset,s=>p(298)(35),cout=>p(299)(36));
FA_ff_10621:FAff port map(x=>p(253)(36),y=>p(254)(36),Cin=>p(255)(36),clock=>clock,reset=>reset,s=>p(298)(36),cout=>p(299)(37));
FA_ff_10622:FAff port map(x=>p(253)(37),y=>p(254)(37),Cin=>p(255)(37),clock=>clock,reset=>reset,s=>p(298)(37),cout=>p(299)(38));
FA_ff_10623:FAff port map(x=>p(253)(38),y=>p(254)(38),Cin=>p(255)(38),clock=>clock,reset=>reset,s=>p(298)(38),cout=>p(299)(39));
FA_ff_10624:FAff port map(x=>p(253)(39),y=>p(254)(39),Cin=>p(255)(39),clock=>clock,reset=>reset,s=>p(298)(39),cout=>p(299)(40));
FA_ff_10625:FAff port map(x=>p(253)(40),y=>p(254)(40),Cin=>p(255)(40),clock=>clock,reset=>reset,s=>p(298)(40),cout=>p(299)(41));
FA_ff_10626:FAff port map(x=>p(253)(41),y=>p(254)(41),Cin=>p(255)(41),clock=>clock,reset=>reset,s=>p(298)(41),cout=>p(299)(42));
FA_ff_10627:FAff port map(x=>p(253)(42),y=>p(254)(42),Cin=>p(255)(42),clock=>clock,reset=>reset,s=>p(298)(42),cout=>p(299)(43));
FA_ff_10628:FAff port map(x=>p(253)(43),y=>p(254)(43),Cin=>p(255)(43),clock=>clock,reset=>reset,s=>p(298)(43),cout=>p(299)(44));
FA_ff_10629:FAff port map(x=>p(253)(44),y=>p(254)(44),Cin=>p(255)(44),clock=>clock,reset=>reset,s=>p(298)(44),cout=>p(299)(45));
FA_ff_10630:FAff port map(x=>p(253)(45),y=>p(254)(45),Cin=>p(255)(45),clock=>clock,reset=>reset,s=>p(298)(45),cout=>p(299)(46));
FA_ff_10631:FAff port map(x=>p(253)(46),y=>p(254)(46),Cin=>p(255)(46),clock=>clock,reset=>reset,s=>p(298)(46),cout=>p(299)(47));
FA_ff_10632:FAff port map(x=>p(253)(47),y=>p(254)(47),Cin=>p(255)(47),clock=>clock,reset=>reset,s=>p(298)(47),cout=>p(299)(48));
FA_ff_10633:FAff port map(x=>p(253)(48),y=>p(254)(48),Cin=>p(255)(48),clock=>clock,reset=>reset,s=>p(298)(48),cout=>p(299)(49));
FA_ff_10634:FAff port map(x=>p(253)(49),y=>p(254)(49),Cin=>p(255)(49),clock=>clock,reset=>reset,s=>p(298)(49),cout=>p(299)(50));
FA_ff_10635:FAff port map(x=>p(253)(50),y=>p(254)(50),Cin=>p(255)(50),clock=>clock,reset=>reset,s=>p(298)(50),cout=>p(299)(51));
FA_ff_10636:FAff port map(x=>p(253)(51),y=>p(254)(51),Cin=>p(255)(51),clock=>clock,reset=>reset,s=>p(298)(51),cout=>p(299)(52));
FA_ff_10637:FAff port map(x=>p(253)(52),y=>p(254)(52),Cin=>p(255)(52),clock=>clock,reset=>reset,s=>p(298)(52),cout=>p(299)(53));
FA_ff_10638:FAff port map(x=>p(253)(53),y=>p(254)(53),Cin=>p(255)(53),clock=>clock,reset=>reset,s=>p(298)(53),cout=>p(299)(54));
FA_ff_10639:FAff port map(x=>p(253)(54),y=>p(254)(54),Cin=>p(255)(54),clock=>clock,reset=>reset,s=>p(298)(54),cout=>p(299)(55));
FA_ff_10640:FAff port map(x=>p(253)(55),y=>p(254)(55),Cin=>p(255)(55),clock=>clock,reset=>reset,s=>p(298)(55),cout=>p(299)(56));
FA_ff_10641:FAff port map(x=>p(253)(56),y=>p(254)(56),Cin=>p(255)(56),clock=>clock,reset=>reset,s=>p(298)(56),cout=>p(299)(57));
FA_ff_10642:FAff port map(x=>p(253)(57),y=>p(254)(57),Cin=>p(255)(57),clock=>clock,reset=>reset,s=>p(298)(57),cout=>p(299)(58));
FA_ff_10643:FAff port map(x=>p(253)(58),y=>p(254)(58),Cin=>p(255)(58),clock=>clock,reset=>reset,s=>p(298)(58),cout=>p(299)(59));
FA_ff_10644:FAff port map(x=>p(253)(59),y=>p(254)(59),Cin=>p(255)(59),clock=>clock,reset=>reset,s=>p(298)(59),cout=>p(299)(60));
FA_ff_10645:FAff port map(x=>p(253)(60),y=>p(254)(60),Cin=>p(255)(60),clock=>clock,reset=>reset,s=>p(298)(60),cout=>p(299)(61));
FA_ff_10646:FAff port map(x=>p(253)(61),y=>p(254)(61),Cin=>p(255)(61),clock=>clock,reset=>reset,s=>p(298)(61),cout=>p(299)(62));
FA_ff_10647:FAff port map(x=>p(253)(62),y=>p(254)(62),Cin=>p(255)(62),clock=>clock,reset=>reset,s=>p(298)(62),cout=>p(299)(63));
FA_ff_10648:FAff port map(x=>p(253)(63),y=>p(254)(63),Cin=>p(255)(63),clock=>clock,reset=>reset,s=>p(298)(63),cout=>p(299)(64));
FA_ff_10649:FAff port map(x=>p(253)(64),y=>p(254)(64),Cin=>p(255)(64),clock=>clock,reset=>reset,s=>p(298)(64),cout=>p(299)(65));
FA_ff_10650:FAff port map(x=>p(253)(65),y=>p(254)(65),Cin=>p(255)(65),clock=>clock,reset=>reset,s=>p(298)(65),cout=>p(299)(66));
FA_ff_10651:FAff port map(x=>p(253)(66),y=>p(254)(66),Cin=>p(255)(66),clock=>clock,reset=>reset,s=>p(298)(66),cout=>p(299)(67));
FA_ff_10652:FAff port map(x=>p(253)(67),y=>p(254)(67),Cin=>p(255)(67),clock=>clock,reset=>reset,s=>p(298)(67),cout=>p(299)(68));
FA_ff_10653:FAff port map(x=>p(253)(68),y=>p(254)(68),Cin=>p(255)(68),clock=>clock,reset=>reset,s=>p(298)(68),cout=>p(299)(69));
FA_ff_10654:FAff port map(x=>p(253)(69),y=>p(254)(69),Cin=>p(255)(69),clock=>clock,reset=>reset,s=>p(298)(69),cout=>p(299)(70));
FA_ff_10655:FAff port map(x=>p(253)(70),y=>p(254)(70),Cin=>p(255)(70),clock=>clock,reset=>reset,s=>p(298)(70),cout=>p(299)(71));
FA_ff_10656:FAff port map(x=>p(253)(71),y=>p(254)(71),Cin=>p(255)(71),clock=>clock,reset=>reset,s=>p(298)(71),cout=>p(299)(72));
FA_ff_10657:FAff port map(x=>p(253)(72),y=>p(254)(72),Cin=>p(255)(72),clock=>clock,reset=>reset,s=>p(298)(72),cout=>p(299)(73));
FA_ff_10658:FAff port map(x=>p(253)(73),y=>p(254)(73),Cin=>p(255)(73),clock=>clock,reset=>reset,s=>p(298)(73),cout=>p(299)(74));
FA_ff_10659:FAff port map(x=>p(253)(74),y=>p(254)(74),Cin=>p(255)(74),clock=>clock,reset=>reset,s=>p(298)(74),cout=>p(299)(75));
FA_ff_10660:FAff port map(x=>p(253)(75),y=>p(254)(75),Cin=>p(255)(75),clock=>clock,reset=>reset,s=>p(298)(75),cout=>p(299)(76));
FA_ff_10661:FAff port map(x=>p(253)(76),y=>p(254)(76),Cin=>p(255)(76),clock=>clock,reset=>reset,s=>p(298)(76),cout=>p(299)(77));
FA_ff_10662:FAff port map(x=>p(253)(77),y=>p(254)(77),Cin=>p(255)(77),clock=>clock,reset=>reset,s=>p(298)(77),cout=>p(299)(78));
FA_ff_10663:FAff port map(x=>p(253)(78),y=>p(254)(78),Cin=>p(255)(78),clock=>clock,reset=>reset,s=>p(298)(78),cout=>p(299)(79));
FA_ff_10664:FAff port map(x=>p(253)(79),y=>p(254)(79),Cin=>p(255)(79),clock=>clock,reset=>reset,s=>p(298)(79),cout=>p(299)(80));
FA_ff_10665:FAff port map(x=>p(253)(80),y=>p(254)(80),Cin=>p(255)(80),clock=>clock,reset=>reset,s=>p(298)(80),cout=>p(299)(81));
FA_ff_10666:FAff port map(x=>p(253)(81),y=>p(254)(81),Cin=>p(255)(81),clock=>clock,reset=>reset,s=>p(298)(81),cout=>p(299)(82));
FA_ff_10667:FAff port map(x=>p(253)(82),y=>p(254)(82),Cin=>p(255)(82),clock=>clock,reset=>reset,s=>p(298)(82),cout=>p(299)(83));
FA_ff_10668:FAff port map(x=>p(253)(83),y=>p(254)(83),Cin=>p(255)(83),clock=>clock,reset=>reset,s=>p(298)(83),cout=>p(299)(84));
FA_ff_10669:FAff port map(x=>p(253)(84),y=>p(254)(84),Cin=>p(255)(84),clock=>clock,reset=>reset,s=>p(298)(84),cout=>p(299)(85));
FA_ff_10670:FAff port map(x=>p(253)(85),y=>p(254)(85),Cin=>p(255)(85),clock=>clock,reset=>reset,s=>p(298)(85),cout=>p(299)(86));
FA_ff_10671:FAff port map(x=>p(253)(86),y=>p(254)(86),Cin=>p(255)(86),clock=>clock,reset=>reset,s=>p(298)(86),cout=>p(299)(87));
FA_ff_10672:FAff port map(x=>p(253)(87),y=>p(254)(87),Cin=>p(255)(87),clock=>clock,reset=>reset,s=>p(298)(87),cout=>p(299)(88));
FA_ff_10673:FAff port map(x=>p(253)(88),y=>p(254)(88),Cin=>p(255)(88),clock=>clock,reset=>reset,s=>p(298)(88),cout=>p(299)(89));
FA_ff_10674:FAff port map(x=>p(253)(89),y=>p(254)(89),Cin=>p(255)(89),clock=>clock,reset=>reset,s=>p(298)(89),cout=>p(299)(90));
FA_ff_10675:FAff port map(x=>p(253)(90),y=>p(254)(90),Cin=>p(255)(90),clock=>clock,reset=>reset,s=>p(298)(90),cout=>p(299)(91));
FA_ff_10676:FAff port map(x=>p(253)(91),y=>p(254)(91),Cin=>p(255)(91),clock=>clock,reset=>reset,s=>p(298)(91),cout=>p(299)(92));
FA_ff_10677:FAff port map(x=>p(253)(92),y=>p(254)(92),Cin=>p(255)(92),clock=>clock,reset=>reset,s=>p(298)(92),cout=>p(299)(93));
FA_ff_10678:FAff port map(x=>p(253)(93),y=>p(254)(93),Cin=>p(255)(93),clock=>clock,reset=>reset,s=>p(298)(93),cout=>p(299)(94));
FA_ff_10679:FAff port map(x=>p(253)(94),y=>p(254)(94),Cin=>p(255)(94),clock=>clock,reset=>reset,s=>p(298)(94),cout=>p(299)(95));
FA_ff_10680:FAff port map(x=>p(253)(95),y=>p(254)(95),Cin=>p(255)(95),clock=>clock,reset=>reset,s=>p(298)(95),cout=>p(299)(96));
FA_ff_10681:FAff port map(x=>p(253)(96),y=>p(254)(96),Cin=>p(255)(96),clock=>clock,reset=>reset,s=>p(298)(96),cout=>p(299)(97));
FA_ff_10682:FAff port map(x=>p(253)(97),y=>p(254)(97),Cin=>p(255)(97),clock=>clock,reset=>reset,s=>p(298)(97),cout=>p(299)(98));
FA_ff_10683:FAff port map(x=>p(253)(98),y=>p(254)(98),Cin=>p(255)(98),clock=>clock,reset=>reset,s=>p(298)(98),cout=>p(299)(99));
FA_ff_10684:FAff port map(x=>p(253)(99),y=>p(254)(99),Cin=>p(255)(99),clock=>clock,reset=>reset,s=>p(298)(99),cout=>p(299)(100));
FA_ff_10685:FAff port map(x=>p(253)(100),y=>p(254)(100),Cin=>p(255)(100),clock=>clock,reset=>reset,s=>p(298)(100),cout=>p(299)(101));
FA_ff_10686:FAff port map(x=>p(253)(101),y=>p(254)(101),Cin=>p(255)(101),clock=>clock,reset=>reset,s=>p(298)(101),cout=>p(299)(102));
FA_ff_10687:FAff port map(x=>p(253)(102),y=>p(254)(102),Cin=>p(255)(102),clock=>clock,reset=>reset,s=>p(298)(102),cout=>p(299)(103));
FA_ff_10688:FAff port map(x=>p(253)(103),y=>p(254)(103),Cin=>p(255)(103),clock=>clock,reset=>reset,s=>p(298)(103),cout=>p(299)(104));
FA_ff_10689:FAff port map(x=>p(253)(104),y=>p(254)(104),Cin=>p(255)(104),clock=>clock,reset=>reset,s=>p(298)(104),cout=>p(299)(105));
FA_ff_10690:FAff port map(x=>p(253)(105),y=>p(254)(105),Cin=>p(255)(105),clock=>clock,reset=>reset,s=>p(298)(105),cout=>p(299)(106));
FA_ff_10691:FAff port map(x=>p(253)(106),y=>p(254)(106),Cin=>p(255)(106),clock=>clock,reset=>reset,s=>p(298)(106),cout=>p(299)(107));
FA_ff_10692:FAff port map(x=>p(253)(107),y=>p(254)(107),Cin=>p(255)(107),clock=>clock,reset=>reset,s=>p(298)(107),cout=>p(299)(108));
FA_ff_10693:FAff port map(x=>p(253)(108),y=>p(254)(108),Cin=>p(255)(108),clock=>clock,reset=>reset,s=>p(298)(108),cout=>p(299)(109));
FA_ff_10694:FAff port map(x=>p(253)(109),y=>p(254)(109),Cin=>p(255)(109),clock=>clock,reset=>reset,s=>p(298)(109),cout=>p(299)(110));
FA_ff_10695:FAff port map(x=>p(253)(110),y=>p(254)(110),Cin=>p(255)(110),clock=>clock,reset=>reset,s=>p(298)(110),cout=>p(299)(111));
FA_ff_10696:FAff port map(x=>p(253)(111),y=>p(254)(111),Cin=>p(255)(111),clock=>clock,reset=>reset,s=>p(298)(111),cout=>p(299)(112));
FA_ff_10697:FAff port map(x=>p(253)(112),y=>p(254)(112),Cin=>p(255)(112),clock=>clock,reset=>reset,s=>p(298)(112),cout=>p(299)(113));
FA_ff_10698:FAff port map(x=>p(253)(113),y=>p(254)(113),Cin=>p(255)(113),clock=>clock,reset=>reset,s=>p(298)(113),cout=>p(299)(114));
FA_ff_10699:FAff port map(x=>p(253)(114),y=>p(254)(114),Cin=>p(255)(114),clock=>clock,reset=>reset,s=>p(298)(114),cout=>p(299)(115));
FA_ff_10700:FAff port map(x=>p(253)(115),y=>p(254)(115),Cin=>p(255)(115),clock=>clock,reset=>reset,s=>p(298)(115),cout=>p(299)(116));
FA_ff_10701:FAff port map(x=>p(253)(116),y=>p(254)(116),Cin=>p(255)(116),clock=>clock,reset=>reset,s=>p(298)(116),cout=>p(299)(117));
FA_ff_10702:FAff port map(x=>p(253)(117),y=>p(254)(117),Cin=>p(255)(117),clock=>clock,reset=>reset,s=>p(298)(117),cout=>p(299)(118));
FA_ff_10703:FAff port map(x=>p(253)(118),y=>p(254)(118),Cin=>p(255)(118),clock=>clock,reset=>reset,s=>p(298)(118),cout=>p(299)(119));
FA_ff_10704:FAff port map(x=>p(253)(119),y=>p(254)(119),Cin=>p(255)(119),clock=>clock,reset=>reset,s=>p(298)(119),cout=>p(299)(120));
FA_ff_10705:FAff port map(x=>p(253)(120),y=>p(254)(120),Cin=>p(255)(120),clock=>clock,reset=>reset,s=>p(298)(120),cout=>p(299)(121));
FA_ff_10706:FAff port map(x=>p(253)(121),y=>p(254)(121),Cin=>p(255)(121),clock=>clock,reset=>reset,s=>p(298)(121),cout=>p(299)(122));
FA_ff_10707:FAff port map(x=>p(253)(122),y=>p(254)(122),Cin=>p(255)(122),clock=>clock,reset=>reset,s=>p(298)(122),cout=>p(299)(123));
FA_ff_10708:FAff port map(x=>p(253)(123),y=>p(254)(123),Cin=>p(255)(123),clock=>clock,reset=>reset,s=>p(298)(123),cout=>p(299)(124));
FA_ff_10709:FAff port map(x=>p(253)(124),y=>p(254)(124),Cin=>p(255)(124),clock=>clock,reset=>reset,s=>p(298)(124),cout=>p(299)(125));
FA_ff_10710:FAff port map(x=>p(253)(125),y=>p(254)(125),Cin=>p(255)(125),clock=>clock,reset=>reset,s=>p(298)(125),cout=>p(299)(126));
FA_ff_10711:FAff port map(x=>p(253)(126),y=>p(254)(126),Cin=>p(255)(126),clock=>clock,reset=>reset,s=>p(298)(126),cout=>p(299)(127));
FA_ff_10712:FAff port map(x=>p(253)(127),y=>p(254)(127),Cin=>p(255)(127),clock=>clock,reset=>reset,s=>p(298)(127),cout=>p(299)(128));
FA_ff_10713:FAff port map(x=>p(253)(128),y=>p(254)(128),Cin=>p(255)(128),clock=>clock,reset=>reset,s=>p(298)(128),cout=>p(299)(129));
p(298)(129)<=p(253)(129);
HA_ff_45:HAff port map(x=>p(256)(0),y=>p(258)(0),clock=>clock,reset=>reset,s=>p(300)(0),c=>p(301)(1));
HA_ff_46:HAff port map(x=>p(256)(1),y=>p(258)(1),clock=>clock,reset=>reset,s=>p(300)(1),c=>p(301)(2));
FA_ff_10714:FAff port map(x=>p(256)(2),y=>p(257)(2),Cin=>p(258)(2),clock=>clock,reset=>reset,s=>p(300)(2),cout=>p(301)(3));
FA_ff_10715:FAff port map(x=>p(256)(3),y=>p(257)(3),Cin=>p(258)(3),clock=>clock,reset=>reset,s=>p(300)(3),cout=>p(301)(4));
FA_ff_10716:FAff port map(x=>p(256)(4),y=>p(257)(4),Cin=>p(258)(4),clock=>clock,reset=>reset,s=>p(300)(4),cout=>p(301)(5));
FA_ff_10717:FAff port map(x=>p(256)(5),y=>p(257)(5),Cin=>p(258)(5),clock=>clock,reset=>reset,s=>p(300)(5),cout=>p(301)(6));
FA_ff_10718:FAff port map(x=>p(256)(6),y=>p(257)(6),Cin=>p(258)(6),clock=>clock,reset=>reset,s=>p(300)(6),cout=>p(301)(7));
FA_ff_10719:FAff port map(x=>p(256)(7),y=>p(257)(7),Cin=>p(258)(7),clock=>clock,reset=>reset,s=>p(300)(7),cout=>p(301)(8));
FA_ff_10720:FAff port map(x=>p(256)(8),y=>p(257)(8),Cin=>p(258)(8),clock=>clock,reset=>reset,s=>p(300)(8),cout=>p(301)(9));
FA_ff_10721:FAff port map(x=>p(256)(9),y=>p(257)(9),Cin=>p(258)(9),clock=>clock,reset=>reset,s=>p(300)(9),cout=>p(301)(10));
FA_ff_10722:FAff port map(x=>p(256)(10),y=>p(257)(10),Cin=>p(258)(10),clock=>clock,reset=>reset,s=>p(300)(10),cout=>p(301)(11));
FA_ff_10723:FAff port map(x=>p(256)(11),y=>p(257)(11),Cin=>p(258)(11),clock=>clock,reset=>reset,s=>p(300)(11),cout=>p(301)(12));
FA_ff_10724:FAff port map(x=>p(256)(12),y=>p(257)(12),Cin=>p(258)(12),clock=>clock,reset=>reset,s=>p(300)(12),cout=>p(301)(13));
FA_ff_10725:FAff port map(x=>p(256)(13),y=>p(257)(13),Cin=>p(258)(13),clock=>clock,reset=>reset,s=>p(300)(13),cout=>p(301)(14));
FA_ff_10726:FAff port map(x=>p(256)(14),y=>p(257)(14),Cin=>p(258)(14),clock=>clock,reset=>reset,s=>p(300)(14),cout=>p(301)(15));
FA_ff_10727:FAff port map(x=>p(256)(15),y=>p(257)(15),Cin=>p(258)(15),clock=>clock,reset=>reset,s=>p(300)(15),cout=>p(301)(16));
FA_ff_10728:FAff port map(x=>p(256)(16),y=>p(257)(16),Cin=>p(258)(16),clock=>clock,reset=>reset,s=>p(300)(16),cout=>p(301)(17));
FA_ff_10729:FAff port map(x=>p(256)(17),y=>p(257)(17),Cin=>p(258)(17),clock=>clock,reset=>reset,s=>p(300)(17),cout=>p(301)(18));
FA_ff_10730:FAff port map(x=>p(256)(18),y=>p(257)(18),Cin=>p(258)(18),clock=>clock,reset=>reset,s=>p(300)(18),cout=>p(301)(19));
FA_ff_10731:FAff port map(x=>p(256)(19),y=>p(257)(19),Cin=>p(258)(19),clock=>clock,reset=>reset,s=>p(300)(19),cout=>p(301)(20));
FA_ff_10732:FAff port map(x=>p(256)(20),y=>p(257)(20),Cin=>p(258)(20),clock=>clock,reset=>reset,s=>p(300)(20),cout=>p(301)(21));
FA_ff_10733:FAff port map(x=>p(256)(21),y=>p(257)(21),Cin=>p(258)(21),clock=>clock,reset=>reset,s=>p(300)(21),cout=>p(301)(22));
FA_ff_10734:FAff port map(x=>p(256)(22),y=>p(257)(22),Cin=>p(258)(22),clock=>clock,reset=>reset,s=>p(300)(22),cout=>p(301)(23));
FA_ff_10735:FAff port map(x=>p(256)(23),y=>p(257)(23),Cin=>p(258)(23),clock=>clock,reset=>reset,s=>p(300)(23),cout=>p(301)(24));
FA_ff_10736:FAff port map(x=>p(256)(24),y=>p(257)(24),Cin=>p(258)(24),clock=>clock,reset=>reset,s=>p(300)(24),cout=>p(301)(25));
FA_ff_10737:FAff port map(x=>p(256)(25),y=>p(257)(25),Cin=>p(258)(25),clock=>clock,reset=>reset,s=>p(300)(25),cout=>p(301)(26));
FA_ff_10738:FAff port map(x=>p(256)(26),y=>p(257)(26),Cin=>p(258)(26),clock=>clock,reset=>reset,s=>p(300)(26),cout=>p(301)(27));
FA_ff_10739:FAff port map(x=>p(256)(27),y=>p(257)(27),Cin=>p(258)(27),clock=>clock,reset=>reset,s=>p(300)(27),cout=>p(301)(28));
FA_ff_10740:FAff port map(x=>p(256)(28),y=>p(257)(28),Cin=>p(258)(28),clock=>clock,reset=>reset,s=>p(300)(28),cout=>p(301)(29));
FA_ff_10741:FAff port map(x=>p(256)(29),y=>p(257)(29),Cin=>p(258)(29),clock=>clock,reset=>reset,s=>p(300)(29),cout=>p(301)(30));
FA_ff_10742:FAff port map(x=>p(256)(30),y=>p(257)(30),Cin=>p(258)(30),clock=>clock,reset=>reset,s=>p(300)(30),cout=>p(301)(31));
FA_ff_10743:FAff port map(x=>p(256)(31),y=>p(257)(31),Cin=>p(258)(31),clock=>clock,reset=>reset,s=>p(300)(31),cout=>p(301)(32));
FA_ff_10744:FAff port map(x=>p(256)(32),y=>p(257)(32),Cin=>p(258)(32),clock=>clock,reset=>reset,s=>p(300)(32),cout=>p(301)(33));
FA_ff_10745:FAff port map(x=>p(256)(33),y=>p(257)(33),Cin=>p(258)(33),clock=>clock,reset=>reset,s=>p(300)(33),cout=>p(301)(34));
FA_ff_10746:FAff port map(x=>p(256)(34),y=>p(257)(34),Cin=>p(258)(34),clock=>clock,reset=>reset,s=>p(300)(34),cout=>p(301)(35));
FA_ff_10747:FAff port map(x=>p(256)(35),y=>p(257)(35),Cin=>p(258)(35),clock=>clock,reset=>reset,s=>p(300)(35),cout=>p(301)(36));
FA_ff_10748:FAff port map(x=>p(256)(36),y=>p(257)(36),Cin=>p(258)(36),clock=>clock,reset=>reset,s=>p(300)(36),cout=>p(301)(37));
FA_ff_10749:FAff port map(x=>p(256)(37),y=>p(257)(37),Cin=>p(258)(37),clock=>clock,reset=>reset,s=>p(300)(37),cout=>p(301)(38));
FA_ff_10750:FAff port map(x=>p(256)(38),y=>p(257)(38),Cin=>p(258)(38),clock=>clock,reset=>reset,s=>p(300)(38),cout=>p(301)(39));
FA_ff_10751:FAff port map(x=>p(256)(39),y=>p(257)(39),Cin=>p(258)(39),clock=>clock,reset=>reset,s=>p(300)(39),cout=>p(301)(40));
FA_ff_10752:FAff port map(x=>p(256)(40),y=>p(257)(40),Cin=>p(258)(40),clock=>clock,reset=>reset,s=>p(300)(40),cout=>p(301)(41));
FA_ff_10753:FAff port map(x=>p(256)(41),y=>p(257)(41),Cin=>p(258)(41),clock=>clock,reset=>reset,s=>p(300)(41),cout=>p(301)(42));
FA_ff_10754:FAff port map(x=>p(256)(42),y=>p(257)(42),Cin=>p(258)(42),clock=>clock,reset=>reset,s=>p(300)(42),cout=>p(301)(43));
FA_ff_10755:FAff port map(x=>p(256)(43),y=>p(257)(43),Cin=>p(258)(43),clock=>clock,reset=>reset,s=>p(300)(43),cout=>p(301)(44));
FA_ff_10756:FAff port map(x=>p(256)(44),y=>p(257)(44),Cin=>p(258)(44),clock=>clock,reset=>reset,s=>p(300)(44),cout=>p(301)(45));
FA_ff_10757:FAff port map(x=>p(256)(45),y=>p(257)(45),Cin=>p(258)(45),clock=>clock,reset=>reset,s=>p(300)(45),cout=>p(301)(46));
FA_ff_10758:FAff port map(x=>p(256)(46),y=>p(257)(46),Cin=>p(258)(46),clock=>clock,reset=>reset,s=>p(300)(46),cout=>p(301)(47));
FA_ff_10759:FAff port map(x=>p(256)(47),y=>p(257)(47),Cin=>p(258)(47),clock=>clock,reset=>reset,s=>p(300)(47),cout=>p(301)(48));
FA_ff_10760:FAff port map(x=>p(256)(48),y=>p(257)(48),Cin=>p(258)(48),clock=>clock,reset=>reset,s=>p(300)(48),cout=>p(301)(49));
FA_ff_10761:FAff port map(x=>p(256)(49),y=>p(257)(49),Cin=>p(258)(49),clock=>clock,reset=>reset,s=>p(300)(49),cout=>p(301)(50));
FA_ff_10762:FAff port map(x=>p(256)(50),y=>p(257)(50),Cin=>p(258)(50),clock=>clock,reset=>reset,s=>p(300)(50),cout=>p(301)(51));
FA_ff_10763:FAff port map(x=>p(256)(51),y=>p(257)(51),Cin=>p(258)(51),clock=>clock,reset=>reset,s=>p(300)(51),cout=>p(301)(52));
FA_ff_10764:FAff port map(x=>p(256)(52),y=>p(257)(52),Cin=>p(258)(52),clock=>clock,reset=>reset,s=>p(300)(52),cout=>p(301)(53));
FA_ff_10765:FAff port map(x=>p(256)(53),y=>p(257)(53),Cin=>p(258)(53),clock=>clock,reset=>reset,s=>p(300)(53),cout=>p(301)(54));
FA_ff_10766:FAff port map(x=>p(256)(54),y=>p(257)(54),Cin=>p(258)(54),clock=>clock,reset=>reset,s=>p(300)(54),cout=>p(301)(55));
FA_ff_10767:FAff port map(x=>p(256)(55),y=>p(257)(55),Cin=>p(258)(55),clock=>clock,reset=>reset,s=>p(300)(55),cout=>p(301)(56));
FA_ff_10768:FAff port map(x=>p(256)(56),y=>p(257)(56),Cin=>p(258)(56),clock=>clock,reset=>reset,s=>p(300)(56),cout=>p(301)(57));
FA_ff_10769:FAff port map(x=>p(256)(57),y=>p(257)(57),Cin=>p(258)(57),clock=>clock,reset=>reset,s=>p(300)(57),cout=>p(301)(58));
FA_ff_10770:FAff port map(x=>p(256)(58),y=>p(257)(58),Cin=>p(258)(58),clock=>clock,reset=>reset,s=>p(300)(58),cout=>p(301)(59));
FA_ff_10771:FAff port map(x=>p(256)(59),y=>p(257)(59),Cin=>p(258)(59),clock=>clock,reset=>reset,s=>p(300)(59),cout=>p(301)(60));
FA_ff_10772:FAff port map(x=>p(256)(60),y=>p(257)(60),Cin=>p(258)(60),clock=>clock,reset=>reset,s=>p(300)(60),cout=>p(301)(61));
FA_ff_10773:FAff port map(x=>p(256)(61),y=>p(257)(61),Cin=>p(258)(61),clock=>clock,reset=>reset,s=>p(300)(61),cout=>p(301)(62));
FA_ff_10774:FAff port map(x=>p(256)(62),y=>p(257)(62),Cin=>p(258)(62),clock=>clock,reset=>reset,s=>p(300)(62),cout=>p(301)(63));
FA_ff_10775:FAff port map(x=>p(256)(63),y=>p(257)(63),Cin=>p(258)(63),clock=>clock,reset=>reset,s=>p(300)(63),cout=>p(301)(64));
FA_ff_10776:FAff port map(x=>p(256)(64),y=>p(257)(64),Cin=>p(258)(64),clock=>clock,reset=>reset,s=>p(300)(64),cout=>p(301)(65));
FA_ff_10777:FAff port map(x=>p(256)(65),y=>p(257)(65),Cin=>p(258)(65),clock=>clock,reset=>reset,s=>p(300)(65),cout=>p(301)(66));
FA_ff_10778:FAff port map(x=>p(256)(66),y=>p(257)(66),Cin=>p(258)(66),clock=>clock,reset=>reset,s=>p(300)(66),cout=>p(301)(67));
FA_ff_10779:FAff port map(x=>p(256)(67),y=>p(257)(67),Cin=>p(258)(67),clock=>clock,reset=>reset,s=>p(300)(67),cout=>p(301)(68));
FA_ff_10780:FAff port map(x=>p(256)(68),y=>p(257)(68),Cin=>p(258)(68),clock=>clock,reset=>reset,s=>p(300)(68),cout=>p(301)(69));
FA_ff_10781:FAff port map(x=>p(256)(69),y=>p(257)(69),Cin=>p(258)(69),clock=>clock,reset=>reset,s=>p(300)(69),cout=>p(301)(70));
FA_ff_10782:FAff port map(x=>p(256)(70),y=>p(257)(70),Cin=>p(258)(70),clock=>clock,reset=>reset,s=>p(300)(70),cout=>p(301)(71));
FA_ff_10783:FAff port map(x=>p(256)(71),y=>p(257)(71),Cin=>p(258)(71),clock=>clock,reset=>reset,s=>p(300)(71),cout=>p(301)(72));
FA_ff_10784:FAff port map(x=>p(256)(72),y=>p(257)(72),Cin=>p(258)(72),clock=>clock,reset=>reset,s=>p(300)(72),cout=>p(301)(73));
FA_ff_10785:FAff port map(x=>p(256)(73),y=>p(257)(73),Cin=>p(258)(73),clock=>clock,reset=>reset,s=>p(300)(73),cout=>p(301)(74));
FA_ff_10786:FAff port map(x=>p(256)(74),y=>p(257)(74),Cin=>p(258)(74),clock=>clock,reset=>reset,s=>p(300)(74),cout=>p(301)(75));
FA_ff_10787:FAff port map(x=>p(256)(75),y=>p(257)(75),Cin=>p(258)(75),clock=>clock,reset=>reset,s=>p(300)(75),cout=>p(301)(76));
FA_ff_10788:FAff port map(x=>p(256)(76),y=>p(257)(76),Cin=>p(258)(76),clock=>clock,reset=>reset,s=>p(300)(76),cout=>p(301)(77));
FA_ff_10789:FAff port map(x=>p(256)(77),y=>p(257)(77),Cin=>p(258)(77),clock=>clock,reset=>reset,s=>p(300)(77),cout=>p(301)(78));
FA_ff_10790:FAff port map(x=>p(256)(78),y=>p(257)(78),Cin=>p(258)(78),clock=>clock,reset=>reset,s=>p(300)(78),cout=>p(301)(79));
FA_ff_10791:FAff port map(x=>p(256)(79),y=>p(257)(79),Cin=>p(258)(79),clock=>clock,reset=>reset,s=>p(300)(79),cout=>p(301)(80));
FA_ff_10792:FAff port map(x=>p(256)(80),y=>p(257)(80),Cin=>p(258)(80),clock=>clock,reset=>reset,s=>p(300)(80),cout=>p(301)(81));
FA_ff_10793:FAff port map(x=>p(256)(81),y=>p(257)(81),Cin=>p(258)(81),clock=>clock,reset=>reset,s=>p(300)(81),cout=>p(301)(82));
FA_ff_10794:FAff port map(x=>p(256)(82),y=>p(257)(82),Cin=>p(258)(82),clock=>clock,reset=>reset,s=>p(300)(82),cout=>p(301)(83));
FA_ff_10795:FAff port map(x=>p(256)(83),y=>p(257)(83),Cin=>p(258)(83),clock=>clock,reset=>reset,s=>p(300)(83),cout=>p(301)(84));
FA_ff_10796:FAff port map(x=>p(256)(84),y=>p(257)(84),Cin=>p(258)(84),clock=>clock,reset=>reset,s=>p(300)(84),cout=>p(301)(85));
FA_ff_10797:FAff port map(x=>p(256)(85),y=>p(257)(85),Cin=>p(258)(85),clock=>clock,reset=>reset,s=>p(300)(85),cout=>p(301)(86));
FA_ff_10798:FAff port map(x=>p(256)(86),y=>p(257)(86),Cin=>p(258)(86),clock=>clock,reset=>reset,s=>p(300)(86),cout=>p(301)(87));
FA_ff_10799:FAff port map(x=>p(256)(87),y=>p(257)(87),Cin=>p(258)(87),clock=>clock,reset=>reset,s=>p(300)(87),cout=>p(301)(88));
FA_ff_10800:FAff port map(x=>p(256)(88),y=>p(257)(88),Cin=>p(258)(88),clock=>clock,reset=>reset,s=>p(300)(88),cout=>p(301)(89));
FA_ff_10801:FAff port map(x=>p(256)(89),y=>p(257)(89),Cin=>p(258)(89),clock=>clock,reset=>reset,s=>p(300)(89),cout=>p(301)(90));
FA_ff_10802:FAff port map(x=>p(256)(90),y=>p(257)(90),Cin=>p(258)(90),clock=>clock,reset=>reset,s=>p(300)(90),cout=>p(301)(91));
FA_ff_10803:FAff port map(x=>p(256)(91),y=>p(257)(91),Cin=>p(258)(91),clock=>clock,reset=>reset,s=>p(300)(91),cout=>p(301)(92));
FA_ff_10804:FAff port map(x=>p(256)(92),y=>p(257)(92),Cin=>p(258)(92),clock=>clock,reset=>reset,s=>p(300)(92),cout=>p(301)(93));
FA_ff_10805:FAff port map(x=>p(256)(93),y=>p(257)(93),Cin=>p(258)(93),clock=>clock,reset=>reset,s=>p(300)(93),cout=>p(301)(94));
FA_ff_10806:FAff port map(x=>p(256)(94),y=>p(257)(94),Cin=>p(258)(94),clock=>clock,reset=>reset,s=>p(300)(94),cout=>p(301)(95));
FA_ff_10807:FAff port map(x=>p(256)(95),y=>p(257)(95),Cin=>p(258)(95),clock=>clock,reset=>reset,s=>p(300)(95),cout=>p(301)(96));
FA_ff_10808:FAff port map(x=>p(256)(96),y=>p(257)(96),Cin=>p(258)(96),clock=>clock,reset=>reset,s=>p(300)(96),cout=>p(301)(97));
FA_ff_10809:FAff port map(x=>p(256)(97),y=>p(257)(97),Cin=>p(258)(97),clock=>clock,reset=>reset,s=>p(300)(97),cout=>p(301)(98));
FA_ff_10810:FAff port map(x=>p(256)(98),y=>p(257)(98),Cin=>p(258)(98),clock=>clock,reset=>reset,s=>p(300)(98),cout=>p(301)(99));
FA_ff_10811:FAff port map(x=>p(256)(99),y=>p(257)(99),Cin=>p(258)(99),clock=>clock,reset=>reset,s=>p(300)(99),cout=>p(301)(100));
FA_ff_10812:FAff port map(x=>p(256)(100),y=>p(257)(100),Cin=>p(258)(100),clock=>clock,reset=>reset,s=>p(300)(100),cout=>p(301)(101));
FA_ff_10813:FAff port map(x=>p(256)(101),y=>p(257)(101),Cin=>p(258)(101),clock=>clock,reset=>reset,s=>p(300)(101),cout=>p(301)(102));
FA_ff_10814:FAff port map(x=>p(256)(102),y=>p(257)(102),Cin=>p(258)(102),clock=>clock,reset=>reset,s=>p(300)(102),cout=>p(301)(103));
FA_ff_10815:FAff port map(x=>p(256)(103),y=>p(257)(103),Cin=>p(258)(103),clock=>clock,reset=>reset,s=>p(300)(103),cout=>p(301)(104));
FA_ff_10816:FAff port map(x=>p(256)(104),y=>p(257)(104),Cin=>p(258)(104),clock=>clock,reset=>reset,s=>p(300)(104),cout=>p(301)(105));
FA_ff_10817:FAff port map(x=>p(256)(105),y=>p(257)(105),Cin=>p(258)(105),clock=>clock,reset=>reset,s=>p(300)(105),cout=>p(301)(106));
FA_ff_10818:FAff port map(x=>p(256)(106),y=>p(257)(106),Cin=>p(258)(106),clock=>clock,reset=>reset,s=>p(300)(106),cout=>p(301)(107));
FA_ff_10819:FAff port map(x=>p(256)(107),y=>p(257)(107),Cin=>p(258)(107),clock=>clock,reset=>reset,s=>p(300)(107),cout=>p(301)(108));
FA_ff_10820:FAff port map(x=>p(256)(108),y=>p(257)(108),Cin=>p(258)(108),clock=>clock,reset=>reset,s=>p(300)(108),cout=>p(301)(109));
FA_ff_10821:FAff port map(x=>p(256)(109),y=>p(257)(109),Cin=>p(258)(109),clock=>clock,reset=>reset,s=>p(300)(109),cout=>p(301)(110));
FA_ff_10822:FAff port map(x=>p(256)(110),y=>p(257)(110),Cin=>p(258)(110),clock=>clock,reset=>reset,s=>p(300)(110),cout=>p(301)(111));
FA_ff_10823:FAff port map(x=>p(256)(111),y=>p(257)(111),Cin=>p(258)(111),clock=>clock,reset=>reset,s=>p(300)(111),cout=>p(301)(112));
FA_ff_10824:FAff port map(x=>p(256)(112),y=>p(257)(112),Cin=>p(258)(112),clock=>clock,reset=>reset,s=>p(300)(112),cout=>p(301)(113));
FA_ff_10825:FAff port map(x=>p(256)(113),y=>p(257)(113),Cin=>p(258)(113),clock=>clock,reset=>reset,s=>p(300)(113),cout=>p(301)(114));
FA_ff_10826:FAff port map(x=>p(256)(114),y=>p(257)(114),Cin=>p(258)(114),clock=>clock,reset=>reset,s=>p(300)(114),cout=>p(301)(115));
FA_ff_10827:FAff port map(x=>p(256)(115),y=>p(257)(115),Cin=>p(258)(115),clock=>clock,reset=>reset,s=>p(300)(115),cout=>p(301)(116));
FA_ff_10828:FAff port map(x=>p(256)(116),y=>p(257)(116),Cin=>p(258)(116),clock=>clock,reset=>reset,s=>p(300)(116),cout=>p(301)(117));
FA_ff_10829:FAff port map(x=>p(256)(117),y=>p(257)(117),Cin=>p(258)(117),clock=>clock,reset=>reset,s=>p(300)(117),cout=>p(301)(118));
FA_ff_10830:FAff port map(x=>p(256)(118),y=>p(257)(118),Cin=>p(258)(118),clock=>clock,reset=>reset,s=>p(300)(118),cout=>p(301)(119));
FA_ff_10831:FAff port map(x=>p(256)(119),y=>p(257)(119),Cin=>p(258)(119),clock=>clock,reset=>reset,s=>p(300)(119),cout=>p(301)(120));
FA_ff_10832:FAff port map(x=>p(256)(120),y=>p(257)(120),Cin=>p(258)(120),clock=>clock,reset=>reset,s=>p(300)(120),cout=>p(301)(121));
FA_ff_10833:FAff port map(x=>p(256)(121),y=>p(257)(121),Cin=>p(258)(121),clock=>clock,reset=>reset,s=>p(300)(121),cout=>p(301)(122));
FA_ff_10834:FAff port map(x=>p(256)(122),y=>p(257)(122),Cin=>p(258)(122),clock=>clock,reset=>reset,s=>p(300)(122),cout=>p(301)(123));
FA_ff_10835:FAff port map(x=>p(256)(123),y=>p(257)(123),Cin=>p(258)(123),clock=>clock,reset=>reset,s=>p(300)(123),cout=>p(301)(124));
FA_ff_10836:FAff port map(x=>p(256)(124),y=>p(257)(124),Cin=>p(258)(124),clock=>clock,reset=>reset,s=>p(300)(124),cout=>p(301)(125));
FA_ff_10837:FAff port map(x=>p(256)(125),y=>p(257)(125),Cin=>p(258)(125),clock=>clock,reset=>reset,s=>p(300)(125),cout=>p(301)(126));
FA_ff_10838:FAff port map(x=>p(256)(126),y=>p(257)(126),Cin=>p(258)(126),clock=>clock,reset=>reset,s=>p(300)(126),cout=>p(301)(127));
FA_ff_10839:FAff port map(x=>p(256)(127),y=>p(257)(127),Cin=>p(258)(127),clock=>clock,reset=>reset,s=>p(300)(127),cout=>p(301)(128));
FA_ff_10840:FAff port map(x=>p(256)(128),y=>p(257)(128),Cin=>p(258)(128),clock=>clock,reset=>reset,s=>p(300)(128),cout=>p(301)(129));
p(300)(129)<=p(257)(129);
p(302)(0)<=p(260)(0);
HA_ff_47:HAff port map(x=>p(259)(1),y=>p(260)(1),clock=>clock,reset=>reset,s=>p(302)(1),c=>p(303)(2));
FA_ff_10841:FAff port map(x=>p(259)(2),y=>p(260)(2),Cin=>p(261)(2),clock=>clock,reset=>reset,s=>p(302)(2),cout=>p(303)(3));
FA_ff_10842:FAff port map(x=>p(259)(3),y=>p(260)(3),Cin=>p(261)(3),clock=>clock,reset=>reset,s=>p(302)(3),cout=>p(303)(4));
FA_ff_10843:FAff port map(x=>p(259)(4),y=>p(260)(4),Cin=>p(261)(4),clock=>clock,reset=>reset,s=>p(302)(4),cout=>p(303)(5));
FA_ff_10844:FAff port map(x=>p(259)(5),y=>p(260)(5),Cin=>p(261)(5),clock=>clock,reset=>reset,s=>p(302)(5),cout=>p(303)(6));
FA_ff_10845:FAff port map(x=>p(259)(6),y=>p(260)(6),Cin=>p(261)(6),clock=>clock,reset=>reset,s=>p(302)(6),cout=>p(303)(7));
FA_ff_10846:FAff port map(x=>p(259)(7),y=>p(260)(7),Cin=>p(261)(7),clock=>clock,reset=>reset,s=>p(302)(7),cout=>p(303)(8));
FA_ff_10847:FAff port map(x=>p(259)(8),y=>p(260)(8),Cin=>p(261)(8),clock=>clock,reset=>reset,s=>p(302)(8),cout=>p(303)(9));
FA_ff_10848:FAff port map(x=>p(259)(9),y=>p(260)(9),Cin=>p(261)(9),clock=>clock,reset=>reset,s=>p(302)(9),cout=>p(303)(10));
FA_ff_10849:FAff port map(x=>p(259)(10),y=>p(260)(10),Cin=>p(261)(10),clock=>clock,reset=>reset,s=>p(302)(10),cout=>p(303)(11));
FA_ff_10850:FAff port map(x=>p(259)(11),y=>p(260)(11),Cin=>p(261)(11),clock=>clock,reset=>reset,s=>p(302)(11),cout=>p(303)(12));
FA_ff_10851:FAff port map(x=>p(259)(12),y=>p(260)(12),Cin=>p(261)(12),clock=>clock,reset=>reset,s=>p(302)(12),cout=>p(303)(13));
FA_ff_10852:FAff port map(x=>p(259)(13),y=>p(260)(13),Cin=>p(261)(13),clock=>clock,reset=>reset,s=>p(302)(13),cout=>p(303)(14));
FA_ff_10853:FAff port map(x=>p(259)(14),y=>p(260)(14),Cin=>p(261)(14),clock=>clock,reset=>reset,s=>p(302)(14),cout=>p(303)(15));
FA_ff_10854:FAff port map(x=>p(259)(15),y=>p(260)(15),Cin=>p(261)(15),clock=>clock,reset=>reset,s=>p(302)(15),cout=>p(303)(16));
FA_ff_10855:FAff port map(x=>p(259)(16),y=>p(260)(16),Cin=>p(261)(16),clock=>clock,reset=>reset,s=>p(302)(16),cout=>p(303)(17));
FA_ff_10856:FAff port map(x=>p(259)(17),y=>p(260)(17),Cin=>p(261)(17),clock=>clock,reset=>reset,s=>p(302)(17),cout=>p(303)(18));
FA_ff_10857:FAff port map(x=>p(259)(18),y=>p(260)(18),Cin=>p(261)(18),clock=>clock,reset=>reset,s=>p(302)(18),cout=>p(303)(19));
FA_ff_10858:FAff port map(x=>p(259)(19),y=>p(260)(19),Cin=>p(261)(19),clock=>clock,reset=>reset,s=>p(302)(19),cout=>p(303)(20));
FA_ff_10859:FAff port map(x=>p(259)(20),y=>p(260)(20),Cin=>p(261)(20),clock=>clock,reset=>reset,s=>p(302)(20),cout=>p(303)(21));
FA_ff_10860:FAff port map(x=>p(259)(21),y=>p(260)(21),Cin=>p(261)(21),clock=>clock,reset=>reset,s=>p(302)(21),cout=>p(303)(22));
FA_ff_10861:FAff port map(x=>p(259)(22),y=>p(260)(22),Cin=>p(261)(22),clock=>clock,reset=>reset,s=>p(302)(22),cout=>p(303)(23));
FA_ff_10862:FAff port map(x=>p(259)(23),y=>p(260)(23),Cin=>p(261)(23),clock=>clock,reset=>reset,s=>p(302)(23),cout=>p(303)(24));
FA_ff_10863:FAff port map(x=>p(259)(24),y=>p(260)(24),Cin=>p(261)(24),clock=>clock,reset=>reset,s=>p(302)(24),cout=>p(303)(25));
FA_ff_10864:FAff port map(x=>p(259)(25),y=>p(260)(25),Cin=>p(261)(25),clock=>clock,reset=>reset,s=>p(302)(25),cout=>p(303)(26));
FA_ff_10865:FAff port map(x=>p(259)(26),y=>p(260)(26),Cin=>p(261)(26),clock=>clock,reset=>reset,s=>p(302)(26),cout=>p(303)(27));
FA_ff_10866:FAff port map(x=>p(259)(27),y=>p(260)(27),Cin=>p(261)(27),clock=>clock,reset=>reset,s=>p(302)(27),cout=>p(303)(28));
FA_ff_10867:FAff port map(x=>p(259)(28),y=>p(260)(28),Cin=>p(261)(28),clock=>clock,reset=>reset,s=>p(302)(28),cout=>p(303)(29));
FA_ff_10868:FAff port map(x=>p(259)(29),y=>p(260)(29),Cin=>p(261)(29),clock=>clock,reset=>reset,s=>p(302)(29),cout=>p(303)(30));
FA_ff_10869:FAff port map(x=>p(259)(30),y=>p(260)(30),Cin=>p(261)(30),clock=>clock,reset=>reset,s=>p(302)(30),cout=>p(303)(31));
FA_ff_10870:FAff port map(x=>p(259)(31),y=>p(260)(31),Cin=>p(261)(31),clock=>clock,reset=>reset,s=>p(302)(31),cout=>p(303)(32));
FA_ff_10871:FAff port map(x=>p(259)(32),y=>p(260)(32),Cin=>p(261)(32),clock=>clock,reset=>reset,s=>p(302)(32),cout=>p(303)(33));
FA_ff_10872:FAff port map(x=>p(259)(33),y=>p(260)(33),Cin=>p(261)(33),clock=>clock,reset=>reset,s=>p(302)(33),cout=>p(303)(34));
FA_ff_10873:FAff port map(x=>p(259)(34),y=>p(260)(34),Cin=>p(261)(34),clock=>clock,reset=>reset,s=>p(302)(34),cout=>p(303)(35));
FA_ff_10874:FAff port map(x=>p(259)(35),y=>p(260)(35),Cin=>p(261)(35),clock=>clock,reset=>reset,s=>p(302)(35),cout=>p(303)(36));
FA_ff_10875:FAff port map(x=>p(259)(36),y=>p(260)(36),Cin=>p(261)(36),clock=>clock,reset=>reset,s=>p(302)(36),cout=>p(303)(37));
FA_ff_10876:FAff port map(x=>p(259)(37),y=>p(260)(37),Cin=>p(261)(37),clock=>clock,reset=>reset,s=>p(302)(37),cout=>p(303)(38));
FA_ff_10877:FAff port map(x=>p(259)(38),y=>p(260)(38),Cin=>p(261)(38),clock=>clock,reset=>reset,s=>p(302)(38),cout=>p(303)(39));
FA_ff_10878:FAff port map(x=>p(259)(39),y=>p(260)(39),Cin=>p(261)(39),clock=>clock,reset=>reset,s=>p(302)(39),cout=>p(303)(40));
FA_ff_10879:FAff port map(x=>p(259)(40),y=>p(260)(40),Cin=>p(261)(40),clock=>clock,reset=>reset,s=>p(302)(40),cout=>p(303)(41));
FA_ff_10880:FAff port map(x=>p(259)(41),y=>p(260)(41),Cin=>p(261)(41),clock=>clock,reset=>reset,s=>p(302)(41),cout=>p(303)(42));
FA_ff_10881:FAff port map(x=>p(259)(42),y=>p(260)(42),Cin=>p(261)(42),clock=>clock,reset=>reset,s=>p(302)(42),cout=>p(303)(43));
FA_ff_10882:FAff port map(x=>p(259)(43),y=>p(260)(43),Cin=>p(261)(43),clock=>clock,reset=>reset,s=>p(302)(43),cout=>p(303)(44));
FA_ff_10883:FAff port map(x=>p(259)(44),y=>p(260)(44),Cin=>p(261)(44),clock=>clock,reset=>reset,s=>p(302)(44),cout=>p(303)(45));
FA_ff_10884:FAff port map(x=>p(259)(45),y=>p(260)(45),Cin=>p(261)(45),clock=>clock,reset=>reset,s=>p(302)(45),cout=>p(303)(46));
FA_ff_10885:FAff port map(x=>p(259)(46),y=>p(260)(46),Cin=>p(261)(46),clock=>clock,reset=>reset,s=>p(302)(46),cout=>p(303)(47));
FA_ff_10886:FAff port map(x=>p(259)(47),y=>p(260)(47),Cin=>p(261)(47),clock=>clock,reset=>reset,s=>p(302)(47),cout=>p(303)(48));
FA_ff_10887:FAff port map(x=>p(259)(48),y=>p(260)(48),Cin=>p(261)(48),clock=>clock,reset=>reset,s=>p(302)(48),cout=>p(303)(49));
FA_ff_10888:FAff port map(x=>p(259)(49),y=>p(260)(49),Cin=>p(261)(49),clock=>clock,reset=>reset,s=>p(302)(49),cout=>p(303)(50));
FA_ff_10889:FAff port map(x=>p(259)(50),y=>p(260)(50),Cin=>p(261)(50),clock=>clock,reset=>reset,s=>p(302)(50),cout=>p(303)(51));
FA_ff_10890:FAff port map(x=>p(259)(51),y=>p(260)(51),Cin=>p(261)(51),clock=>clock,reset=>reset,s=>p(302)(51),cout=>p(303)(52));
FA_ff_10891:FAff port map(x=>p(259)(52),y=>p(260)(52),Cin=>p(261)(52),clock=>clock,reset=>reset,s=>p(302)(52),cout=>p(303)(53));
FA_ff_10892:FAff port map(x=>p(259)(53),y=>p(260)(53),Cin=>p(261)(53),clock=>clock,reset=>reset,s=>p(302)(53),cout=>p(303)(54));
FA_ff_10893:FAff port map(x=>p(259)(54),y=>p(260)(54),Cin=>p(261)(54),clock=>clock,reset=>reset,s=>p(302)(54),cout=>p(303)(55));
FA_ff_10894:FAff port map(x=>p(259)(55),y=>p(260)(55),Cin=>p(261)(55),clock=>clock,reset=>reset,s=>p(302)(55),cout=>p(303)(56));
FA_ff_10895:FAff port map(x=>p(259)(56),y=>p(260)(56),Cin=>p(261)(56),clock=>clock,reset=>reset,s=>p(302)(56),cout=>p(303)(57));
FA_ff_10896:FAff port map(x=>p(259)(57),y=>p(260)(57),Cin=>p(261)(57),clock=>clock,reset=>reset,s=>p(302)(57),cout=>p(303)(58));
FA_ff_10897:FAff port map(x=>p(259)(58),y=>p(260)(58),Cin=>p(261)(58),clock=>clock,reset=>reset,s=>p(302)(58),cout=>p(303)(59));
FA_ff_10898:FAff port map(x=>p(259)(59),y=>p(260)(59),Cin=>p(261)(59),clock=>clock,reset=>reset,s=>p(302)(59),cout=>p(303)(60));
FA_ff_10899:FAff port map(x=>p(259)(60),y=>p(260)(60),Cin=>p(261)(60),clock=>clock,reset=>reset,s=>p(302)(60),cout=>p(303)(61));
FA_ff_10900:FAff port map(x=>p(259)(61),y=>p(260)(61),Cin=>p(261)(61),clock=>clock,reset=>reset,s=>p(302)(61),cout=>p(303)(62));
FA_ff_10901:FAff port map(x=>p(259)(62),y=>p(260)(62),Cin=>p(261)(62),clock=>clock,reset=>reset,s=>p(302)(62),cout=>p(303)(63));
FA_ff_10902:FAff port map(x=>p(259)(63),y=>p(260)(63),Cin=>p(261)(63),clock=>clock,reset=>reset,s=>p(302)(63),cout=>p(303)(64));
FA_ff_10903:FAff port map(x=>p(259)(64),y=>p(260)(64),Cin=>p(261)(64),clock=>clock,reset=>reset,s=>p(302)(64),cout=>p(303)(65));
FA_ff_10904:FAff port map(x=>p(259)(65),y=>p(260)(65),Cin=>p(261)(65),clock=>clock,reset=>reset,s=>p(302)(65),cout=>p(303)(66));
FA_ff_10905:FAff port map(x=>p(259)(66),y=>p(260)(66),Cin=>p(261)(66),clock=>clock,reset=>reset,s=>p(302)(66),cout=>p(303)(67));
FA_ff_10906:FAff port map(x=>p(259)(67),y=>p(260)(67),Cin=>p(261)(67),clock=>clock,reset=>reset,s=>p(302)(67),cout=>p(303)(68));
FA_ff_10907:FAff port map(x=>p(259)(68),y=>p(260)(68),Cin=>p(261)(68),clock=>clock,reset=>reset,s=>p(302)(68),cout=>p(303)(69));
FA_ff_10908:FAff port map(x=>p(259)(69),y=>p(260)(69),Cin=>p(261)(69),clock=>clock,reset=>reset,s=>p(302)(69),cout=>p(303)(70));
FA_ff_10909:FAff port map(x=>p(259)(70),y=>p(260)(70),Cin=>p(261)(70),clock=>clock,reset=>reset,s=>p(302)(70),cout=>p(303)(71));
FA_ff_10910:FAff port map(x=>p(259)(71),y=>p(260)(71),Cin=>p(261)(71),clock=>clock,reset=>reset,s=>p(302)(71),cout=>p(303)(72));
FA_ff_10911:FAff port map(x=>p(259)(72),y=>p(260)(72),Cin=>p(261)(72),clock=>clock,reset=>reset,s=>p(302)(72),cout=>p(303)(73));
FA_ff_10912:FAff port map(x=>p(259)(73),y=>p(260)(73),Cin=>p(261)(73),clock=>clock,reset=>reset,s=>p(302)(73),cout=>p(303)(74));
FA_ff_10913:FAff port map(x=>p(259)(74),y=>p(260)(74),Cin=>p(261)(74),clock=>clock,reset=>reset,s=>p(302)(74),cout=>p(303)(75));
FA_ff_10914:FAff port map(x=>p(259)(75),y=>p(260)(75),Cin=>p(261)(75),clock=>clock,reset=>reset,s=>p(302)(75),cout=>p(303)(76));
FA_ff_10915:FAff port map(x=>p(259)(76),y=>p(260)(76),Cin=>p(261)(76),clock=>clock,reset=>reset,s=>p(302)(76),cout=>p(303)(77));
FA_ff_10916:FAff port map(x=>p(259)(77),y=>p(260)(77),Cin=>p(261)(77),clock=>clock,reset=>reset,s=>p(302)(77),cout=>p(303)(78));
FA_ff_10917:FAff port map(x=>p(259)(78),y=>p(260)(78),Cin=>p(261)(78),clock=>clock,reset=>reset,s=>p(302)(78),cout=>p(303)(79));
FA_ff_10918:FAff port map(x=>p(259)(79),y=>p(260)(79),Cin=>p(261)(79),clock=>clock,reset=>reset,s=>p(302)(79),cout=>p(303)(80));
FA_ff_10919:FAff port map(x=>p(259)(80),y=>p(260)(80),Cin=>p(261)(80),clock=>clock,reset=>reset,s=>p(302)(80),cout=>p(303)(81));
FA_ff_10920:FAff port map(x=>p(259)(81),y=>p(260)(81),Cin=>p(261)(81),clock=>clock,reset=>reset,s=>p(302)(81),cout=>p(303)(82));
FA_ff_10921:FAff port map(x=>p(259)(82),y=>p(260)(82),Cin=>p(261)(82),clock=>clock,reset=>reset,s=>p(302)(82),cout=>p(303)(83));
FA_ff_10922:FAff port map(x=>p(259)(83),y=>p(260)(83),Cin=>p(261)(83),clock=>clock,reset=>reset,s=>p(302)(83),cout=>p(303)(84));
FA_ff_10923:FAff port map(x=>p(259)(84),y=>p(260)(84),Cin=>p(261)(84),clock=>clock,reset=>reset,s=>p(302)(84),cout=>p(303)(85));
FA_ff_10924:FAff port map(x=>p(259)(85),y=>p(260)(85),Cin=>p(261)(85),clock=>clock,reset=>reset,s=>p(302)(85),cout=>p(303)(86));
FA_ff_10925:FAff port map(x=>p(259)(86),y=>p(260)(86),Cin=>p(261)(86),clock=>clock,reset=>reset,s=>p(302)(86),cout=>p(303)(87));
FA_ff_10926:FAff port map(x=>p(259)(87),y=>p(260)(87),Cin=>p(261)(87),clock=>clock,reset=>reset,s=>p(302)(87),cout=>p(303)(88));
FA_ff_10927:FAff port map(x=>p(259)(88),y=>p(260)(88),Cin=>p(261)(88),clock=>clock,reset=>reset,s=>p(302)(88),cout=>p(303)(89));
FA_ff_10928:FAff port map(x=>p(259)(89),y=>p(260)(89),Cin=>p(261)(89),clock=>clock,reset=>reset,s=>p(302)(89),cout=>p(303)(90));
FA_ff_10929:FAff port map(x=>p(259)(90),y=>p(260)(90),Cin=>p(261)(90),clock=>clock,reset=>reset,s=>p(302)(90),cout=>p(303)(91));
FA_ff_10930:FAff port map(x=>p(259)(91),y=>p(260)(91),Cin=>p(261)(91),clock=>clock,reset=>reset,s=>p(302)(91),cout=>p(303)(92));
FA_ff_10931:FAff port map(x=>p(259)(92),y=>p(260)(92),Cin=>p(261)(92),clock=>clock,reset=>reset,s=>p(302)(92),cout=>p(303)(93));
FA_ff_10932:FAff port map(x=>p(259)(93),y=>p(260)(93),Cin=>p(261)(93),clock=>clock,reset=>reset,s=>p(302)(93),cout=>p(303)(94));
FA_ff_10933:FAff port map(x=>p(259)(94),y=>p(260)(94),Cin=>p(261)(94),clock=>clock,reset=>reset,s=>p(302)(94),cout=>p(303)(95));
FA_ff_10934:FAff port map(x=>p(259)(95),y=>p(260)(95),Cin=>p(261)(95),clock=>clock,reset=>reset,s=>p(302)(95),cout=>p(303)(96));
FA_ff_10935:FAff port map(x=>p(259)(96),y=>p(260)(96),Cin=>p(261)(96),clock=>clock,reset=>reset,s=>p(302)(96),cout=>p(303)(97));
FA_ff_10936:FAff port map(x=>p(259)(97),y=>p(260)(97),Cin=>p(261)(97),clock=>clock,reset=>reset,s=>p(302)(97),cout=>p(303)(98));
FA_ff_10937:FAff port map(x=>p(259)(98),y=>p(260)(98),Cin=>p(261)(98),clock=>clock,reset=>reset,s=>p(302)(98),cout=>p(303)(99));
FA_ff_10938:FAff port map(x=>p(259)(99),y=>p(260)(99),Cin=>p(261)(99),clock=>clock,reset=>reset,s=>p(302)(99),cout=>p(303)(100));
FA_ff_10939:FAff port map(x=>p(259)(100),y=>p(260)(100),Cin=>p(261)(100),clock=>clock,reset=>reset,s=>p(302)(100),cout=>p(303)(101));
FA_ff_10940:FAff port map(x=>p(259)(101),y=>p(260)(101),Cin=>p(261)(101),clock=>clock,reset=>reset,s=>p(302)(101),cout=>p(303)(102));
FA_ff_10941:FAff port map(x=>p(259)(102),y=>p(260)(102),Cin=>p(261)(102),clock=>clock,reset=>reset,s=>p(302)(102),cout=>p(303)(103));
FA_ff_10942:FAff port map(x=>p(259)(103),y=>p(260)(103),Cin=>p(261)(103),clock=>clock,reset=>reset,s=>p(302)(103),cout=>p(303)(104));
FA_ff_10943:FAff port map(x=>p(259)(104),y=>p(260)(104),Cin=>p(261)(104),clock=>clock,reset=>reset,s=>p(302)(104),cout=>p(303)(105));
FA_ff_10944:FAff port map(x=>p(259)(105),y=>p(260)(105),Cin=>p(261)(105),clock=>clock,reset=>reset,s=>p(302)(105),cout=>p(303)(106));
FA_ff_10945:FAff port map(x=>p(259)(106),y=>p(260)(106),Cin=>p(261)(106),clock=>clock,reset=>reset,s=>p(302)(106),cout=>p(303)(107));
FA_ff_10946:FAff port map(x=>p(259)(107),y=>p(260)(107),Cin=>p(261)(107),clock=>clock,reset=>reset,s=>p(302)(107),cout=>p(303)(108));
FA_ff_10947:FAff port map(x=>p(259)(108),y=>p(260)(108),Cin=>p(261)(108),clock=>clock,reset=>reset,s=>p(302)(108),cout=>p(303)(109));
FA_ff_10948:FAff port map(x=>p(259)(109),y=>p(260)(109),Cin=>p(261)(109),clock=>clock,reset=>reset,s=>p(302)(109),cout=>p(303)(110));
FA_ff_10949:FAff port map(x=>p(259)(110),y=>p(260)(110),Cin=>p(261)(110),clock=>clock,reset=>reset,s=>p(302)(110),cout=>p(303)(111));
FA_ff_10950:FAff port map(x=>p(259)(111),y=>p(260)(111),Cin=>p(261)(111),clock=>clock,reset=>reset,s=>p(302)(111),cout=>p(303)(112));
FA_ff_10951:FAff port map(x=>p(259)(112),y=>p(260)(112),Cin=>p(261)(112),clock=>clock,reset=>reset,s=>p(302)(112),cout=>p(303)(113));
FA_ff_10952:FAff port map(x=>p(259)(113),y=>p(260)(113),Cin=>p(261)(113),clock=>clock,reset=>reset,s=>p(302)(113),cout=>p(303)(114));
FA_ff_10953:FAff port map(x=>p(259)(114),y=>p(260)(114),Cin=>p(261)(114),clock=>clock,reset=>reset,s=>p(302)(114),cout=>p(303)(115));
FA_ff_10954:FAff port map(x=>p(259)(115),y=>p(260)(115),Cin=>p(261)(115),clock=>clock,reset=>reset,s=>p(302)(115),cout=>p(303)(116));
FA_ff_10955:FAff port map(x=>p(259)(116),y=>p(260)(116),Cin=>p(261)(116),clock=>clock,reset=>reset,s=>p(302)(116),cout=>p(303)(117));
FA_ff_10956:FAff port map(x=>p(259)(117),y=>p(260)(117),Cin=>p(261)(117),clock=>clock,reset=>reset,s=>p(302)(117),cout=>p(303)(118));
FA_ff_10957:FAff port map(x=>p(259)(118),y=>p(260)(118),Cin=>p(261)(118),clock=>clock,reset=>reset,s=>p(302)(118),cout=>p(303)(119));
FA_ff_10958:FAff port map(x=>p(259)(119),y=>p(260)(119),Cin=>p(261)(119),clock=>clock,reset=>reset,s=>p(302)(119),cout=>p(303)(120));
FA_ff_10959:FAff port map(x=>p(259)(120),y=>p(260)(120),Cin=>p(261)(120),clock=>clock,reset=>reset,s=>p(302)(120),cout=>p(303)(121));
FA_ff_10960:FAff port map(x=>p(259)(121),y=>p(260)(121),Cin=>p(261)(121),clock=>clock,reset=>reset,s=>p(302)(121),cout=>p(303)(122));
FA_ff_10961:FAff port map(x=>p(259)(122),y=>p(260)(122),Cin=>p(261)(122),clock=>clock,reset=>reset,s=>p(302)(122),cout=>p(303)(123));
FA_ff_10962:FAff port map(x=>p(259)(123),y=>p(260)(123),Cin=>p(261)(123),clock=>clock,reset=>reset,s=>p(302)(123),cout=>p(303)(124));
FA_ff_10963:FAff port map(x=>p(259)(124),y=>p(260)(124),Cin=>p(261)(124),clock=>clock,reset=>reset,s=>p(302)(124),cout=>p(303)(125));
FA_ff_10964:FAff port map(x=>p(259)(125),y=>p(260)(125),Cin=>p(261)(125),clock=>clock,reset=>reset,s=>p(302)(125),cout=>p(303)(126));
FA_ff_10965:FAff port map(x=>p(259)(126),y=>p(260)(126),Cin=>p(261)(126),clock=>clock,reset=>reset,s=>p(302)(126),cout=>p(303)(127));
FA_ff_10966:FAff port map(x=>p(259)(127),y=>p(260)(127),Cin=>p(261)(127),clock=>clock,reset=>reset,s=>p(302)(127),cout=>p(303)(128));
FA_ff_10967:FAff port map(x=>p(259)(128),y=>p(260)(128),Cin=>p(261)(128),clock=>clock,reset=>reset,s=>p(302)(128),cout=>p(303)(129));
p(302)(129)<=p(261)(129);
HA_ff_48:HAff port map(x=>p(262)(0),y=>p(264)(0),clock=>clock,reset=>reset,s=>p(304)(0),c=>p(305)(1));
FA_ff_10968:FAff port map(x=>p(262)(1),y=>p(263)(1),Cin=>p(264)(1),clock=>clock,reset=>reset,s=>p(304)(1),cout=>p(305)(2));
FA_ff_10969:FAff port map(x=>p(262)(2),y=>p(263)(2),Cin=>p(264)(2),clock=>clock,reset=>reset,s=>p(304)(2),cout=>p(305)(3));
FA_ff_10970:FAff port map(x=>p(262)(3),y=>p(263)(3),Cin=>p(264)(3),clock=>clock,reset=>reset,s=>p(304)(3),cout=>p(305)(4));
FA_ff_10971:FAff port map(x=>p(262)(4),y=>p(263)(4),Cin=>p(264)(4),clock=>clock,reset=>reset,s=>p(304)(4),cout=>p(305)(5));
FA_ff_10972:FAff port map(x=>p(262)(5),y=>p(263)(5),Cin=>p(264)(5),clock=>clock,reset=>reset,s=>p(304)(5),cout=>p(305)(6));
FA_ff_10973:FAff port map(x=>p(262)(6),y=>p(263)(6),Cin=>p(264)(6),clock=>clock,reset=>reset,s=>p(304)(6),cout=>p(305)(7));
FA_ff_10974:FAff port map(x=>p(262)(7),y=>p(263)(7),Cin=>p(264)(7),clock=>clock,reset=>reset,s=>p(304)(7),cout=>p(305)(8));
FA_ff_10975:FAff port map(x=>p(262)(8),y=>p(263)(8),Cin=>p(264)(8),clock=>clock,reset=>reset,s=>p(304)(8),cout=>p(305)(9));
FA_ff_10976:FAff port map(x=>p(262)(9),y=>p(263)(9),Cin=>p(264)(9),clock=>clock,reset=>reset,s=>p(304)(9),cout=>p(305)(10));
FA_ff_10977:FAff port map(x=>p(262)(10),y=>p(263)(10),Cin=>p(264)(10),clock=>clock,reset=>reset,s=>p(304)(10),cout=>p(305)(11));
FA_ff_10978:FAff port map(x=>p(262)(11),y=>p(263)(11),Cin=>p(264)(11),clock=>clock,reset=>reset,s=>p(304)(11),cout=>p(305)(12));
FA_ff_10979:FAff port map(x=>p(262)(12),y=>p(263)(12),Cin=>p(264)(12),clock=>clock,reset=>reset,s=>p(304)(12),cout=>p(305)(13));
FA_ff_10980:FAff port map(x=>p(262)(13),y=>p(263)(13),Cin=>p(264)(13),clock=>clock,reset=>reset,s=>p(304)(13),cout=>p(305)(14));
FA_ff_10981:FAff port map(x=>p(262)(14),y=>p(263)(14),Cin=>p(264)(14),clock=>clock,reset=>reset,s=>p(304)(14),cout=>p(305)(15));
FA_ff_10982:FAff port map(x=>p(262)(15),y=>p(263)(15),Cin=>p(264)(15),clock=>clock,reset=>reset,s=>p(304)(15),cout=>p(305)(16));
FA_ff_10983:FAff port map(x=>p(262)(16),y=>p(263)(16),Cin=>p(264)(16),clock=>clock,reset=>reset,s=>p(304)(16),cout=>p(305)(17));
FA_ff_10984:FAff port map(x=>p(262)(17),y=>p(263)(17),Cin=>p(264)(17),clock=>clock,reset=>reset,s=>p(304)(17),cout=>p(305)(18));
FA_ff_10985:FAff port map(x=>p(262)(18),y=>p(263)(18),Cin=>p(264)(18),clock=>clock,reset=>reset,s=>p(304)(18),cout=>p(305)(19));
FA_ff_10986:FAff port map(x=>p(262)(19),y=>p(263)(19),Cin=>p(264)(19),clock=>clock,reset=>reset,s=>p(304)(19),cout=>p(305)(20));
FA_ff_10987:FAff port map(x=>p(262)(20),y=>p(263)(20),Cin=>p(264)(20),clock=>clock,reset=>reset,s=>p(304)(20),cout=>p(305)(21));
FA_ff_10988:FAff port map(x=>p(262)(21),y=>p(263)(21),Cin=>p(264)(21),clock=>clock,reset=>reset,s=>p(304)(21),cout=>p(305)(22));
FA_ff_10989:FAff port map(x=>p(262)(22),y=>p(263)(22),Cin=>p(264)(22),clock=>clock,reset=>reset,s=>p(304)(22),cout=>p(305)(23));
FA_ff_10990:FAff port map(x=>p(262)(23),y=>p(263)(23),Cin=>p(264)(23),clock=>clock,reset=>reset,s=>p(304)(23),cout=>p(305)(24));
FA_ff_10991:FAff port map(x=>p(262)(24),y=>p(263)(24),Cin=>p(264)(24),clock=>clock,reset=>reset,s=>p(304)(24),cout=>p(305)(25));
FA_ff_10992:FAff port map(x=>p(262)(25),y=>p(263)(25),Cin=>p(264)(25),clock=>clock,reset=>reset,s=>p(304)(25),cout=>p(305)(26));
FA_ff_10993:FAff port map(x=>p(262)(26),y=>p(263)(26),Cin=>p(264)(26),clock=>clock,reset=>reset,s=>p(304)(26),cout=>p(305)(27));
FA_ff_10994:FAff port map(x=>p(262)(27),y=>p(263)(27),Cin=>p(264)(27),clock=>clock,reset=>reset,s=>p(304)(27),cout=>p(305)(28));
FA_ff_10995:FAff port map(x=>p(262)(28),y=>p(263)(28),Cin=>p(264)(28),clock=>clock,reset=>reset,s=>p(304)(28),cout=>p(305)(29));
FA_ff_10996:FAff port map(x=>p(262)(29),y=>p(263)(29),Cin=>p(264)(29),clock=>clock,reset=>reset,s=>p(304)(29),cout=>p(305)(30));
FA_ff_10997:FAff port map(x=>p(262)(30),y=>p(263)(30),Cin=>p(264)(30),clock=>clock,reset=>reset,s=>p(304)(30),cout=>p(305)(31));
FA_ff_10998:FAff port map(x=>p(262)(31),y=>p(263)(31),Cin=>p(264)(31),clock=>clock,reset=>reset,s=>p(304)(31),cout=>p(305)(32));
FA_ff_10999:FAff port map(x=>p(262)(32),y=>p(263)(32),Cin=>p(264)(32),clock=>clock,reset=>reset,s=>p(304)(32),cout=>p(305)(33));
FA_ff_11000:FAff port map(x=>p(262)(33),y=>p(263)(33),Cin=>p(264)(33),clock=>clock,reset=>reset,s=>p(304)(33),cout=>p(305)(34));
FA_ff_11001:FAff port map(x=>p(262)(34),y=>p(263)(34),Cin=>p(264)(34),clock=>clock,reset=>reset,s=>p(304)(34),cout=>p(305)(35));
FA_ff_11002:FAff port map(x=>p(262)(35),y=>p(263)(35),Cin=>p(264)(35),clock=>clock,reset=>reset,s=>p(304)(35),cout=>p(305)(36));
FA_ff_11003:FAff port map(x=>p(262)(36),y=>p(263)(36),Cin=>p(264)(36),clock=>clock,reset=>reset,s=>p(304)(36),cout=>p(305)(37));
FA_ff_11004:FAff port map(x=>p(262)(37),y=>p(263)(37),Cin=>p(264)(37),clock=>clock,reset=>reset,s=>p(304)(37),cout=>p(305)(38));
FA_ff_11005:FAff port map(x=>p(262)(38),y=>p(263)(38),Cin=>p(264)(38),clock=>clock,reset=>reset,s=>p(304)(38),cout=>p(305)(39));
FA_ff_11006:FAff port map(x=>p(262)(39),y=>p(263)(39),Cin=>p(264)(39),clock=>clock,reset=>reset,s=>p(304)(39),cout=>p(305)(40));
FA_ff_11007:FAff port map(x=>p(262)(40),y=>p(263)(40),Cin=>p(264)(40),clock=>clock,reset=>reset,s=>p(304)(40),cout=>p(305)(41));
FA_ff_11008:FAff port map(x=>p(262)(41),y=>p(263)(41),Cin=>p(264)(41),clock=>clock,reset=>reset,s=>p(304)(41),cout=>p(305)(42));
FA_ff_11009:FAff port map(x=>p(262)(42),y=>p(263)(42),Cin=>p(264)(42),clock=>clock,reset=>reset,s=>p(304)(42),cout=>p(305)(43));
FA_ff_11010:FAff port map(x=>p(262)(43),y=>p(263)(43),Cin=>p(264)(43),clock=>clock,reset=>reset,s=>p(304)(43),cout=>p(305)(44));
FA_ff_11011:FAff port map(x=>p(262)(44),y=>p(263)(44),Cin=>p(264)(44),clock=>clock,reset=>reset,s=>p(304)(44),cout=>p(305)(45));
FA_ff_11012:FAff port map(x=>p(262)(45),y=>p(263)(45),Cin=>p(264)(45),clock=>clock,reset=>reset,s=>p(304)(45),cout=>p(305)(46));
FA_ff_11013:FAff port map(x=>p(262)(46),y=>p(263)(46),Cin=>p(264)(46),clock=>clock,reset=>reset,s=>p(304)(46),cout=>p(305)(47));
FA_ff_11014:FAff port map(x=>p(262)(47),y=>p(263)(47),Cin=>p(264)(47),clock=>clock,reset=>reset,s=>p(304)(47),cout=>p(305)(48));
FA_ff_11015:FAff port map(x=>p(262)(48),y=>p(263)(48),Cin=>p(264)(48),clock=>clock,reset=>reset,s=>p(304)(48),cout=>p(305)(49));
FA_ff_11016:FAff port map(x=>p(262)(49),y=>p(263)(49),Cin=>p(264)(49),clock=>clock,reset=>reset,s=>p(304)(49),cout=>p(305)(50));
FA_ff_11017:FAff port map(x=>p(262)(50),y=>p(263)(50),Cin=>p(264)(50),clock=>clock,reset=>reset,s=>p(304)(50),cout=>p(305)(51));
FA_ff_11018:FAff port map(x=>p(262)(51),y=>p(263)(51),Cin=>p(264)(51),clock=>clock,reset=>reset,s=>p(304)(51),cout=>p(305)(52));
FA_ff_11019:FAff port map(x=>p(262)(52),y=>p(263)(52),Cin=>p(264)(52),clock=>clock,reset=>reset,s=>p(304)(52),cout=>p(305)(53));
FA_ff_11020:FAff port map(x=>p(262)(53),y=>p(263)(53),Cin=>p(264)(53),clock=>clock,reset=>reset,s=>p(304)(53),cout=>p(305)(54));
FA_ff_11021:FAff port map(x=>p(262)(54),y=>p(263)(54),Cin=>p(264)(54),clock=>clock,reset=>reset,s=>p(304)(54),cout=>p(305)(55));
FA_ff_11022:FAff port map(x=>p(262)(55),y=>p(263)(55),Cin=>p(264)(55),clock=>clock,reset=>reset,s=>p(304)(55),cout=>p(305)(56));
FA_ff_11023:FAff port map(x=>p(262)(56),y=>p(263)(56),Cin=>p(264)(56),clock=>clock,reset=>reset,s=>p(304)(56),cout=>p(305)(57));
FA_ff_11024:FAff port map(x=>p(262)(57),y=>p(263)(57),Cin=>p(264)(57),clock=>clock,reset=>reset,s=>p(304)(57),cout=>p(305)(58));
FA_ff_11025:FAff port map(x=>p(262)(58),y=>p(263)(58),Cin=>p(264)(58),clock=>clock,reset=>reset,s=>p(304)(58),cout=>p(305)(59));
FA_ff_11026:FAff port map(x=>p(262)(59),y=>p(263)(59),Cin=>p(264)(59),clock=>clock,reset=>reset,s=>p(304)(59),cout=>p(305)(60));
FA_ff_11027:FAff port map(x=>p(262)(60),y=>p(263)(60),Cin=>p(264)(60),clock=>clock,reset=>reset,s=>p(304)(60),cout=>p(305)(61));
FA_ff_11028:FAff port map(x=>p(262)(61),y=>p(263)(61),Cin=>p(264)(61),clock=>clock,reset=>reset,s=>p(304)(61),cout=>p(305)(62));
FA_ff_11029:FAff port map(x=>p(262)(62),y=>p(263)(62),Cin=>p(264)(62),clock=>clock,reset=>reset,s=>p(304)(62),cout=>p(305)(63));
FA_ff_11030:FAff port map(x=>p(262)(63),y=>p(263)(63),Cin=>p(264)(63),clock=>clock,reset=>reset,s=>p(304)(63),cout=>p(305)(64));
FA_ff_11031:FAff port map(x=>p(262)(64),y=>p(263)(64),Cin=>p(264)(64),clock=>clock,reset=>reset,s=>p(304)(64),cout=>p(305)(65));
FA_ff_11032:FAff port map(x=>p(262)(65),y=>p(263)(65),Cin=>p(264)(65),clock=>clock,reset=>reset,s=>p(304)(65),cout=>p(305)(66));
FA_ff_11033:FAff port map(x=>p(262)(66),y=>p(263)(66),Cin=>p(264)(66),clock=>clock,reset=>reset,s=>p(304)(66),cout=>p(305)(67));
FA_ff_11034:FAff port map(x=>p(262)(67),y=>p(263)(67),Cin=>p(264)(67),clock=>clock,reset=>reset,s=>p(304)(67),cout=>p(305)(68));
FA_ff_11035:FAff port map(x=>p(262)(68),y=>p(263)(68),Cin=>p(264)(68),clock=>clock,reset=>reset,s=>p(304)(68),cout=>p(305)(69));
FA_ff_11036:FAff port map(x=>p(262)(69),y=>p(263)(69),Cin=>p(264)(69),clock=>clock,reset=>reset,s=>p(304)(69),cout=>p(305)(70));
FA_ff_11037:FAff port map(x=>p(262)(70),y=>p(263)(70),Cin=>p(264)(70),clock=>clock,reset=>reset,s=>p(304)(70),cout=>p(305)(71));
FA_ff_11038:FAff port map(x=>p(262)(71),y=>p(263)(71),Cin=>p(264)(71),clock=>clock,reset=>reset,s=>p(304)(71),cout=>p(305)(72));
FA_ff_11039:FAff port map(x=>p(262)(72),y=>p(263)(72),Cin=>p(264)(72),clock=>clock,reset=>reset,s=>p(304)(72),cout=>p(305)(73));
FA_ff_11040:FAff port map(x=>p(262)(73),y=>p(263)(73),Cin=>p(264)(73),clock=>clock,reset=>reset,s=>p(304)(73),cout=>p(305)(74));
FA_ff_11041:FAff port map(x=>p(262)(74),y=>p(263)(74),Cin=>p(264)(74),clock=>clock,reset=>reset,s=>p(304)(74),cout=>p(305)(75));
FA_ff_11042:FAff port map(x=>p(262)(75),y=>p(263)(75),Cin=>p(264)(75),clock=>clock,reset=>reset,s=>p(304)(75),cout=>p(305)(76));
FA_ff_11043:FAff port map(x=>p(262)(76),y=>p(263)(76),Cin=>p(264)(76),clock=>clock,reset=>reset,s=>p(304)(76),cout=>p(305)(77));
FA_ff_11044:FAff port map(x=>p(262)(77),y=>p(263)(77),Cin=>p(264)(77),clock=>clock,reset=>reset,s=>p(304)(77),cout=>p(305)(78));
FA_ff_11045:FAff port map(x=>p(262)(78),y=>p(263)(78),Cin=>p(264)(78),clock=>clock,reset=>reset,s=>p(304)(78),cout=>p(305)(79));
FA_ff_11046:FAff port map(x=>p(262)(79),y=>p(263)(79),Cin=>p(264)(79),clock=>clock,reset=>reset,s=>p(304)(79),cout=>p(305)(80));
FA_ff_11047:FAff port map(x=>p(262)(80),y=>p(263)(80),Cin=>p(264)(80),clock=>clock,reset=>reset,s=>p(304)(80),cout=>p(305)(81));
FA_ff_11048:FAff port map(x=>p(262)(81),y=>p(263)(81),Cin=>p(264)(81),clock=>clock,reset=>reset,s=>p(304)(81),cout=>p(305)(82));
FA_ff_11049:FAff port map(x=>p(262)(82),y=>p(263)(82),Cin=>p(264)(82),clock=>clock,reset=>reset,s=>p(304)(82),cout=>p(305)(83));
FA_ff_11050:FAff port map(x=>p(262)(83),y=>p(263)(83),Cin=>p(264)(83),clock=>clock,reset=>reset,s=>p(304)(83),cout=>p(305)(84));
FA_ff_11051:FAff port map(x=>p(262)(84),y=>p(263)(84),Cin=>p(264)(84),clock=>clock,reset=>reset,s=>p(304)(84),cout=>p(305)(85));
FA_ff_11052:FAff port map(x=>p(262)(85),y=>p(263)(85),Cin=>p(264)(85),clock=>clock,reset=>reset,s=>p(304)(85),cout=>p(305)(86));
FA_ff_11053:FAff port map(x=>p(262)(86),y=>p(263)(86),Cin=>p(264)(86),clock=>clock,reset=>reset,s=>p(304)(86),cout=>p(305)(87));
FA_ff_11054:FAff port map(x=>p(262)(87),y=>p(263)(87),Cin=>p(264)(87),clock=>clock,reset=>reset,s=>p(304)(87),cout=>p(305)(88));
FA_ff_11055:FAff port map(x=>p(262)(88),y=>p(263)(88),Cin=>p(264)(88),clock=>clock,reset=>reset,s=>p(304)(88),cout=>p(305)(89));
FA_ff_11056:FAff port map(x=>p(262)(89),y=>p(263)(89),Cin=>p(264)(89),clock=>clock,reset=>reset,s=>p(304)(89),cout=>p(305)(90));
FA_ff_11057:FAff port map(x=>p(262)(90),y=>p(263)(90),Cin=>p(264)(90),clock=>clock,reset=>reset,s=>p(304)(90),cout=>p(305)(91));
FA_ff_11058:FAff port map(x=>p(262)(91),y=>p(263)(91),Cin=>p(264)(91),clock=>clock,reset=>reset,s=>p(304)(91),cout=>p(305)(92));
FA_ff_11059:FAff port map(x=>p(262)(92),y=>p(263)(92),Cin=>p(264)(92),clock=>clock,reset=>reset,s=>p(304)(92),cout=>p(305)(93));
FA_ff_11060:FAff port map(x=>p(262)(93),y=>p(263)(93),Cin=>p(264)(93),clock=>clock,reset=>reset,s=>p(304)(93),cout=>p(305)(94));
FA_ff_11061:FAff port map(x=>p(262)(94),y=>p(263)(94),Cin=>p(264)(94),clock=>clock,reset=>reset,s=>p(304)(94),cout=>p(305)(95));
FA_ff_11062:FAff port map(x=>p(262)(95),y=>p(263)(95),Cin=>p(264)(95),clock=>clock,reset=>reset,s=>p(304)(95),cout=>p(305)(96));
FA_ff_11063:FAff port map(x=>p(262)(96),y=>p(263)(96),Cin=>p(264)(96),clock=>clock,reset=>reset,s=>p(304)(96),cout=>p(305)(97));
FA_ff_11064:FAff port map(x=>p(262)(97),y=>p(263)(97),Cin=>p(264)(97),clock=>clock,reset=>reset,s=>p(304)(97),cout=>p(305)(98));
FA_ff_11065:FAff port map(x=>p(262)(98),y=>p(263)(98),Cin=>p(264)(98),clock=>clock,reset=>reset,s=>p(304)(98),cout=>p(305)(99));
FA_ff_11066:FAff port map(x=>p(262)(99),y=>p(263)(99),Cin=>p(264)(99),clock=>clock,reset=>reset,s=>p(304)(99),cout=>p(305)(100));
FA_ff_11067:FAff port map(x=>p(262)(100),y=>p(263)(100),Cin=>p(264)(100),clock=>clock,reset=>reset,s=>p(304)(100),cout=>p(305)(101));
FA_ff_11068:FAff port map(x=>p(262)(101),y=>p(263)(101),Cin=>p(264)(101),clock=>clock,reset=>reset,s=>p(304)(101),cout=>p(305)(102));
FA_ff_11069:FAff port map(x=>p(262)(102),y=>p(263)(102),Cin=>p(264)(102),clock=>clock,reset=>reset,s=>p(304)(102),cout=>p(305)(103));
FA_ff_11070:FAff port map(x=>p(262)(103),y=>p(263)(103),Cin=>p(264)(103),clock=>clock,reset=>reset,s=>p(304)(103),cout=>p(305)(104));
FA_ff_11071:FAff port map(x=>p(262)(104),y=>p(263)(104),Cin=>p(264)(104),clock=>clock,reset=>reset,s=>p(304)(104),cout=>p(305)(105));
FA_ff_11072:FAff port map(x=>p(262)(105),y=>p(263)(105),Cin=>p(264)(105),clock=>clock,reset=>reset,s=>p(304)(105),cout=>p(305)(106));
FA_ff_11073:FAff port map(x=>p(262)(106),y=>p(263)(106),Cin=>p(264)(106),clock=>clock,reset=>reset,s=>p(304)(106),cout=>p(305)(107));
FA_ff_11074:FAff port map(x=>p(262)(107),y=>p(263)(107),Cin=>p(264)(107),clock=>clock,reset=>reset,s=>p(304)(107),cout=>p(305)(108));
FA_ff_11075:FAff port map(x=>p(262)(108),y=>p(263)(108),Cin=>p(264)(108),clock=>clock,reset=>reset,s=>p(304)(108),cout=>p(305)(109));
FA_ff_11076:FAff port map(x=>p(262)(109),y=>p(263)(109),Cin=>p(264)(109),clock=>clock,reset=>reset,s=>p(304)(109),cout=>p(305)(110));
FA_ff_11077:FAff port map(x=>p(262)(110),y=>p(263)(110),Cin=>p(264)(110),clock=>clock,reset=>reset,s=>p(304)(110),cout=>p(305)(111));
FA_ff_11078:FAff port map(x=>p(262)(111),y=>p(263)(111),Cin=>p(264)(111),clock=>clock,reset=>reset,s=>p(304)(111),cout=>p(305)(112));
FA_ff_11079:FAff port map(x=>p(262)(112),y=>p(263)(112),Cin=>p(264)(112),clock=>clock,reset=>reset,s=>p(304)(112),cout=>p(305)(113));
FA_ff_11080:FAff port map(x=>p(262)(113),y=>p(263)(113),Cin=>p(264)(113),clock=>clock,reset=>reset,s=>p(304)(113),cout=>p(305)(114));
FA_ff_11081:FAff port map(x=>p(262)(114),y=>p(263)(114),Cin=>p(264)(114),clock=>clock,reset=>reset,s=>p(304)(114),cout=>p(305)(115));
FA_ff_11082:FAff port map(x=>p(262)(115),y=>p(263)(115),Cin=>p(264)(115),clock=>clock,reset=>reset,s=>p(304)(115),cout=>p(305)(116));
FA_ff_11083:FAff port map(x=>p(262)(116),y=>p(263)(116),Cin=>p(264)(116),clock=>clock,reset=>reset,s=>p(304)(116),cout=>p(305)(117));
FA_ff_11084:FAff port map(x=>p(262)(117),y=>p(263)(117),Cin=>p(264)(117),clock=>clock,reset=>reset,s=>p(304)(117),cout=>p(305)(118));
FA_ff_11085:FAff port map(x=>p(262)(118),y=>p(263)(118),Cin=>p(264)(118),clock=>clock,reset=>reset,s=>p(304)(118),cout=>p(305)(119));
FA_ff_11086:FAff port map(x=>p(262)(119),y=>p(263)(119),Cin=>p(264)(119),clock=>clock,reset=>reset,s=>p(304)(119),cout=>p(305)(120));
FA_ff_11087:FAff port map(x=>p(262)(120),y=>p(263)(120),Cin=>p(264)(120),clock=>clock,reset=>reset,s=>p(304)(120),cout=>p(305)(121));
FA_ff_11088:FAff port map(x=>p(262)(121),y=>p(263)(121),Cin=>p(264)(121),clock=>clock,reset=>reset,s=>p(304)(121),cout=>p(305)(122));
FA_ff_11089:FAff port map(x=>p(262)(122),y=>p(263)(122),Cin=>p(264)(122),clock=>clock,reset=>reset,s=>p(304)(122),cout=>p(305)(123));
FA_ff_11090:FAff port map(x=>p(262)(123),y=>p(263)(123),Cin=>p(264)(123),clock=>clock,reset=>reset,s=>p(304)(123),cout=>p(305)(124));
FA_ff_11091:FAff port map(x=>p(262)(124),y=>p(263)(124),Cin=>p(264)(124),clock=>clock,reset=>reset,s=>p(304)(124),cout=>p(305)(125));
FA_ff_11092:FAff port map(x=>p(262)(125),y=>p(263)(125),Cin=>p(264)(125),clock=>clock,reset=>reset,s=>p(304)(125),cout=>p(305)(126));
FA_ff_11093:FAff port map(x=>p(262)(126),y=>p(263)(126),Cin=>p(264)(126),clock=>clock,reset=>reset,s=>p(304)(126),cout=>p(305)(127));
FA_ff_11094:FAff port map(x=>p(262)(127),y=>p(263)(127),Cin=>p(264)(127),clock=>clock,reset=>reset,s=>p(304)(127),cout=>p(305)(128));
FA_ff_11095:FAff port map(x=>p(262)(128),y=>p(263)(128),Cin=>p(264)(128),clock=>clock,reset=>reset,s=>p(304)(128),cout=>p(305)(129));
p(306)(0)<=p(266)(0);
HA_ff_49:HAff port map(x=>p(266)(1),y=>p(267)(1),clock=>clock,reset=>reset,s=>p(306)(1),c=>p(307)(2));
FA_ff_11096:FAff port map(x=>p(265)(2),y=>p(266)(2),Cin=>p(267)(2),clock=>clock,reset=>reset,s=>p(306)(2),cout=>p(307)(3));
FA_ff_11097:FAff port map(x=>p(265)(3),y=>p(266)(3),Cin=>p(267)(3),clock=>clock,reset=>reset,s=>p(306)(3),cout=>p(307)(4));
FA_ff_11098:FAff port map(x=>p(265)(4),y=>p(266)(4),Cin=>p(267)(4),clock=>clock,reset=>reset,s=>p(306)(4),cout=>p(307)(5));
FA_ff_11099:FAff port map(x=>p(265)(5),y=>p(266)(5),Cin=>p(267)(5),clock=>clock,reset=>reset,s=>p(306)(5),cout=>p(307)(6));
FA_ff_11100:FAff port map(x=>p(265)(6),y=>p(266)(6),Cin=>p(267)(6),clock=>clock,reset=>reset,s=>p(306)(6),cout=>p(307)(7));
FA_ff_11101:FAff port map(x=>p(265)(7),y=>p(266)(7),Cin=>p(267)(7),clock=>clock,reset=>reset,s=>p(306)(7),cout=>p(307)(8));
FA_ff_11102:FAff port map(x=>p(265)(8),y=>p(266)(8),Cin=>p(267)(8),clock=>clock,reset=>reset,s=>p(306)(8),cout=>p(307)(9));
FA_ff_11103:FAff port map(x=>p(265)(9),y=>p(266)(9),Cin=>p(267)(9),clock=>clock,reset=>reset,s=>p(306)(9),cout=>p(307)(10));
FA_ff_11104:FAff port map(x=>p(265)(10),y=>p(266)(10),Cin=>p(267)(10),clock=>clock,reset=>reset,s=>p(306)(10),cout=>p(307)(11));
FA_ff_11105:FAff port map(x=>p(265)(11),y=>p(266)(11),Cin=>p(267)(11),clock=>clock,reset=>reset,s=>p(306)(11),cout=>p(307)(12));
FA_ff_11106:FAff port map(x=>p(265)(12),y=>p(266)(12),Cin=>p(267)(12),clock=>clock,reset=>reset,s=>p(306)(12),cout=>p(307)(13));
FA_ff_11107:FAff port map(x=>p(265)(13),y=>p(266)(13),Cin=>p(267)(13),clock=>clock,reset=>reset,s=>p(306)(13),cout=>p(307)(14));
FA_ff_11108:FAff port map(x=>p(265)(14),y=>p(266)(14),Cin=>p(267)(14),clock=>clock,reset=>reset,s=>p(306)(14),cout=>p(307)(15));
FA_ff_11109:FAff port map(x=>p(265)(15),y=>p(266)(15),Cin=>p(267)(15),clock=>clock,reset=>reset,s=>p(306)(15),cout=>p(307)(16));
FA_ff_11110:FAff port map(x=>p(265)(16),y=>p(266)(16),Cin=>p(267)(16),clock=>clock,reset=>reset,s=>p(306)(16),cout=>p(307)(17));
FA_ff_11111:FAff port map(x=>p(265)(17),y=>p(266)(17),Cin=>p(267)(17),clock=>clock,reset=>reset,s=>p(306)(17),cout=>p(307)(18));
FA_ff_11112:FAff port map(x=>p(265)(18),y=>p(266)(18),Cin=>p(267)(18),clock=>clock,reset=>reset,s=>p(306)(18),cout=>p(307)(19));
FA_ff_11113:FAff port map(x=>p(265)(19),y=>p(266)(19),Cin=>p(267)(19),clock=>clock,reset=>reset,s=>p(306)(19),cout=>p(307)(20));
FA_ff_11114:FAff port map(x=>p(265)(20),y=>p(266)(20),Cin=>p(267)(20),clock=>clock,reset=>reset,s=>p(306)(20),cout=>p(307)(21));
FA_ff_11115:FAff port map(x=>p(265)(21),y=>p(266)(21),Cin=>p(267)(21),clock=>clock,reset=>reset,s=>p(306)(21),cout=>p(307)(22));
FA_ff_11116:FAff port map(x=>p(265)(22),y=>p(266)(22),Cin=>p(267)(22),clock=>clock,reset=>reset,s=>p(306)(22),cout=>p(307)(23));
FA_ff_11117:FAff port map(x=>p(265)(23),y=>p(266)(23),Cin=>p(267)(23),clock=>clock,reset=>reset,s=>p(306)(23),cout=>p(307)(24));
FA_ff_11118:FAff port map(x=>p(265)(24),y=>p(266)(24),Cin=>p(267)(24),clock=>clock,reset=>reset,s=>p(306)(24),cout=>p(307)(25));
FA_ff_11119:FAff port map(x=>p(265)(25),y=>p(266)(25),Cin=>p(267)(25),clock=>clock,reset=>reset,s=>p(306)(25),cout=>p(307)(26));
FA_ff_11120:FAff port map(x=>p(265)(26),y=>p(266)(26),Cin=>p(267)(26),clock=>clock,reset=>reset,s=>p(306)(26),cout=>p(307)(27));
FA_ff_11121:FAff port map(x=>p(265)(27),y=>p(266)(27),Cin=>p(267)(27),clock=>clock,reset=>reset,s=>p(306)(27),cout=>p(307)(28));
FA_ff_11122:FAff port map(x=>p(265)(28),y=>p(266)(28),Cin=>p(267)(28),clock=>clock,reset=>reset,s=>p(306)(28),cout=>p(307)(29));
FA_ff_11123:FAff port map(x=>p(265)(29),y=>p(266)(29),Cin=>p(267)(29),clock=>clock,reset=>reset,s=>p(306)(29),cout=>p(307)(30));
FA_ff_11124:FAff port map(x=>p(265)(30),y=>p(266)(30),Cin=>p(267)(30),clock=>clock,reset=>reset,s=>p(306)(30),cout=>p(307)(31));
FA_ff_11125:FAff port map(x=>p(265)(31),y=>p(266)(31),Cin=>p(267)(31),clock=>clock,reset=>reset,s=>p(306)(31),cout=>p(307)(32));
FA_ff_11126:FAff port map(x=>p(265)(32),y=>p(266)(32),Cin=>p(267)(32),clock=>clock,reset=>reset,s=>p(306)(32),cout=>p(307)(33));
FA_ff_11127:FAff port map(x=>p(265)(33),y=>p(266)(33),Cin=>p(267)(33),clock=>clock,reset=>reset,s=>p(306)(33),cout=>p(307)(34));
FA_ff_11128:FAff port map(x=>p(265)(34),y=>p(266)(34),Cin=>p(267)(34),clock=>clock,reset=>reset,s=>p(306)(34),cout=>p(307)(35));
FA_ff_11129:FAff port map(x=>p(265)(35),y=>p(266)(35),Cin=>p(267)(35),clock=>clock,reset=>reset,s=>p(306)(35),cout=>p(307)(36));
FA_ff_11130:FAff port map(x=>p(265)(36),y=>p(266)(36),Cin=>p(267)(36),clock=>clock,reset=>reset,s=>p(306)(36),cout=>p(307)(37));
FA_ff_11131:FAff port map(x=>p(265)(37),y=>p(266)(37),Cin=>p(267)(37),clock=>clock,reset=>reset,s=>p(306)(37),cout=>p(307)(38));
FA_ff_11132:FAff port map(x=>p(265)(38),y=>p(266)(38),Cin=>p(267)(38),clock=>clock,reset=>reset,s=>p(306)(38),cout=>p(307)(39));
FA_ff_11133:FAff port map(x=>p(265)(39),y=>p(266)(39),Cin=>p(267)(39),clock=>clock,reset=>reset,s=>p(306)(39),cout=>p(307)(40));
FA_ff_11134:FAff port map(x=>p(265)(40),y=>p(266)(40),Cin=>p(267)(40),clock=>clock,reset=>reset,s=>p(306)(40),cout=>p(307)(41));
FA_ff_11135:FAff port map(x=>p(265)(41),y=>p(266)(41),Cin=>p(267)(41),clock=>clock,reset=>reset,s=>p(306)(41),cout=>p(307)(42));
FA_ff_11136:FAff port map(x=>p(265)(42),y=>p(266)(42),Cin=>p(267)(42),clock=>clock,reset=>reset,s=>p(306)(42),cout=>p(307)(43));
FA_ff_11137:FAff port map(x=>p(265)(43),y=>p(266)(43),Cin=>p(267)(43),clock=>clock,reset=>reset,s=>p(306)(43),cout=>p(307)(44));
FA_ff_11138:FAff port map(x=>p(265)(44),y=>p(266)(44),Cin=>p(267)(44),clock=>clock,reset=>reset,s=>p(306)(44),cout=>p(307)(45));
FA_ff_11139:FAff port map(x=>p(265)(45),y=>p(266)(45),Cin=>p(267)(45),clock=>clock,reset=>reset,s=>p(306)(45),cout=>p(307)(46));
FA_ff_11140:FAff port map(x=>p(265)(46),y=>p(266)(46),Cin=>p(267)(46),clock=>clock,reset=>reset,s=>p(306)(46),cout=>p(307)(47));
FA_ff_11141:FAff port map(x=>p(265)(47),y=>p(266)(47),Cin=>p(267)(47),clock=>clock,reset=>reset,s=>p(306)(47),cout=>p(307)(48));
FA_ff_11142:FAff port map(x=>p(265)(48),y=>p(266)(48),Cin=>p(267)(48),clock=>clock,reset=>reset,s=>p(306)(48),cout=>p(307)(49));
FA_ff_11143:FAff port map(x=>p(265)(49),y=>p(266)(49),Cin=>p(267)(49),clock=>clock,reset=>reset,s=>p(306)(49),cout=>p(307)(50));
FA_ff_11144:FAff port map(x=>p(265)(50),y=>p(266)(50),Cin=>p(267)(50),clock=>clock,reset=>reset,s=>p(306)(50),cout=>p(307)(51));
FA_ff_11145:FAff port map(x=>p(265)(51),y=>p(266)(51),Cin=>p(267)(51),clock=>clock,reset=>reset,s=>p(306)(51),cout=>p(307)(52));
FA_ff_11146:FAff port map(x=>p(265)(52),y=>p(266)(52),Cin=>p(267)(52),clock=>clock,reset=>reset,s=>p(306)(52),cout=>p(307)(53));
FA_ff_11147:FAff port map(x=>p(265)(53),y=>p(266)(53),Cin=>p(267)(53),clock=>clock,reset=>reset,s=>p(306)(53),cout=>p(307)(54));
FA_ff_11148:FAff port map(x=>p(265)(54),y=>p(266)(54),Cin=>p(267)(54),clock=>clock,reset=>reset,s=>p(306)(54),cout=>p(307)(55));
FA_ff_11149:FAff port map(x=>p(265)(55),y=>p(266)(55),Cin=>p(267)(55),clock=>clock,reset=>reset,s=>p(306)(55),cout=>p(307)(56));
FA_ff_11150:FAff port map(x=>p(265)(56),y=>p(266)(56),Cin=>p(267)(56),clock=>clock,reset=>reset,s=>p(306)(56),cout=>p(307)(57));
FA_ff_11151:FAff port map(x=>p(265)(57),y=>p(266)(57),Cin=>p(267)(57),clock=>clock,reset=>reset,s=>p(306)(57),cout=>p(307)(58));
FA_ff_11152:FAff port map(x=>p(265)(58),y=>p(266)(58),Cin=>p(267)(58),clock=>clock,reset=>reset,s=>p(306)(58),cout=>p(307)(59));
FA_ff_11153:FAff port map(x=>p(265)(59),y=>p(266)(59),Cin=>p(267)(59),clock=>clock,reset=>reset,s=>p(306)(59),cout=>p(307)(60));
FA_ff_11154:FAff port map(x=>p(265)(60),y=>p(266)(60),Cin=>p(267)(60),clock=>clock,reset=>reset,s=>p(306)(60),cout=>p(307)(61));
FA_ff_11155:FAff port map(x=>p(265)(61),y=>p(266)(61),Cin=>p(267)(61),clock=>clock,reset=>reset,s=>p(306)(61),cout=>p(307)(62));
FA_ff_11156:FAff port map(x=>p(265)(62),y=>p(266)(62),Cin=>p(267)(62),clock=>clock,reset=>reset,s=>p(306)(62),cout=>p(307)(63));
FA_ff_11157:FAff port map(x=>p(265)(63),y=>p(266)(63),Cin=>p(267)(63),clock=>clock,reset=>reset,s=>p(306)(63),cout=>p(307)(64));
FA_ff_11158:FAff port map(x=>p(265)(64),y=>p(266)(64),Cin=>p(267)(64),clock=>clock,reset=>reset,s=>p(306)(64),cout=>p(307)(65));
FA_ff_11159:FAff port map(x=>p(265)(65),y=>p(266)(65),Cin=>p(267)(65),clock=>clock,reset=>reset,s=>p(306)(65),cout=>p(307)(66));
FA_ff_11160:FAff port map(x=>p(265)(66),y=>p(266)(66),Cin=>p(267)(66),clock=>clock,reset=>reset,s=>p(306)(66),cout=>p(307)(67));
FA_ff_11161:FAff port map(x=>p(265)(67),y=>p(266)(67),Cin=>p(267)(67),clock=>clock,reset=>reset,s=>p(306)(67),cout=>p(307)(68));
FA_ff_11162:FAff port map(x=>p(265)(68),y=>p(266)(68),Cin=>p(267)(68),clock=>clock,reset=>reset,s=>p(306)(68),cout=>p(307)(69));
FA_ff_11163:FAff port map(x=>p(265)(69),y=>p(266)(69),Cin=>p(267)(69),clock=>clock,reset=>reset,s=>p(306)(69),cout=>p(307)(70));
FA_ff_11164:FAff port map(x=>p(265)(70),y=>p(266)(70),Cin=>p(267)(70),clock=>clock,reset=>reset,s=>p(306)(70),cout=>p(307)(71));
FA_ff_11165:FAff port map(x=>p(265)(71),y=>p(266)(71),Cin=>p(267)(71),clock=>clock,reset=>reset,s=>p(306)(71),cout=>p(307)(72));
FA_ff_11166:FAff port map(x=>p(265)(72),y=>p(266)(72),Cin=>p(267)(72),clock=>clock,reset=>reset,s=>p(306)(72),cout=>p(307)(73));
FA_ff_11167:FAff port map(x=>p(265)(73),y=>p(266)(73),Cin=>p(267)(73),clock=>clock,reset=>reset,s=>p(306)(73),cout=>p(307)(74));
FA_ff_11168:FAff port map(x=>p(265)(74),y=>p(266)(74),Cin=>p(267)(74),clock=>clock,reset=>reset,s=>p(306)(74),cout=>p(307)(75));
FA_ff_11169:FAff port map(x=>p(265)(75),y=>p(266)(75),Cin=>p(267)(75),clock=>clock,reset=>reset,s=>p(306)(75),cout=>p(307)(76));
FA_ff_11170:FAff port map(x=>p(265)(76),y=>p(266)(76),Cin=>p(267)(76),clock=>clock,reset=>reset,s=>p(306)(76),cout=>p(307)(77));
FA_ff_11171:FAff port map(x=>p(265)(77),y=>p(266)(77),Cin=>p(267)(77),clock=>clock,reset=>reset,s=>p(306)(77),cout=>p(307)(78));
FA_ff_11172:FAff port map(x=>p(265)(78),y=>p(266)(78),Cin=>p(267)(78),clock=>clock,reset=>reset,s=>p(306)(78),cout=>p(307)(79));
FA_ff_11173:FAff port map(x=>p(265)(79),y=>p(266)(79),Cin=>p(267)(79),clock=>clock,reset=>reset,s=>p(306)(79),cout=>p(307)(80));
FA_ff_11174:FAff port map(x=>p(265)(80),y=>p(266)(80),Cin=>p(267)(80),clock=>clock,reset=>reset,s=>p(306)(80),cout=>p(307)(81));
FA_ff_11175:FAff port map(x=>p(265)(81),y=>p(266)(81),Cin=>p(267)(81),clock=>clock,reset=>reset,s=>p(306)(81),cout=>p(307)(82));
FA_ff_11176:FAff port map(x=>p(265)(82),y=>p(266)(82),Cin=>p(267)(82),clock=>clock,reset=>reset,s=>p(306)(82),cout=>p(307)(83));
FA_ff_11177:FAff port map(x=>p(265)(83),y=>p(266)(83),Cin=>p(267)(83),clock=>clock,reset=>reset,s=>p(306)(83),cout=>p(307)(84));
FA_ff_11178:FAff port map(x=>p(265)(84),y=>p(266)(84),Cin=>p(267)(84),clock=>clock,reset=>reset,s=>p(306)(84),cout=>p(307)(85));
FA_ff_11179:FAff port map(x=>p(265)(85),y=>p(266)(85),Cin=>p(267)(85),clock=>clock,reset=>reset,s=>p(306)(85),cout=>p(307)(86));
FA_ff_11180:FAff port map(x=>p(265)(86),y=>p(266)(86),Cin=>p(267)(86),clock=>clock,reset=>reset,s=>p(306)(86),cout=>p(307)(87));
FA_ff_11181:FAff port map(x=>p(265)(87),y=>p(266)(87),Cin=>p(267)(87),clock=>clock,reset=>reset,s=>p(306)(87),cout=>p(307)(88));
FA_ff_11182:FAff port map(x=>p(265)(88),y=>p(266)(88),Cin=>p(267)(88),clock=>clock,reset=>reset,s=>p(306)(88),cout=>p(307)(89));
FA_ff_11183:FAff port map(x=>p(265)(89),y=>p(266)(89),Cin=>p(267)(89),clock=>clock,reset=>reset,s=>p(306)(89),cout=>p(307)(90));
FA_ff_11184:FAff port map(x=>p(265)(90),y=>p(266)(90),Cin=>p(267)(90),clock=>clock,reset=>reset,s=>p(306)(90),cout=>p(307)(91));
FA_ff_11185:FAff port map(x=>p(265)(91),y=>p(266)(91),Cin=>p(267)(91),clock=>clock,reset=>reset,s=>p(306)(91),cout=>p(307)(92));
FA_ff_11186:FAff port map(x=>p(265)(92),y=>p(266)(92),Cin=>p(267)(92),clock=>clock,reset=>reset,s=>p(306)(92),cout=>p(307)(93));
FA_ff_11187:FAff port map(x=>p(265)(93),y=>p(266)(93),Cin=>p(267)(93),clock=>clock,reset=>reset,s=>p(306)(93),cout=>p(307)(94));
FA_ff_11188:FAff port map(x=>p(265)(94),y=>p(266)(94),Cin=>p(267)(94),clock=>clock,reset=>reset,s=>p(306)(94),cout=>p(307)(95));
FA_ff_11189:FAff port map(x=>p(265)(95),y=>p(266)(95),Cin=>p(267)(95),clock=>clock,reset=>reset,s=>p(306)(95),cout=>p(307)(96));
FA_ff_11190:FAff port map(x=>p(265)(96),y=>p(266)(96),Cin=>p(267)(96),clock=>clock,reset=>reset,s=>p(306)(96),cout=>p(307)(97));
FA_ff_11191:FAff port map(x=>p(265)(97),y=>p(266)(97),Cin=>p(267)(97),clock=>clock,reset=>reset,s=>p(306)(97),cout=>p(307)(98));
FA_ff_11192:FAff port map(x=>p(265)(98),y=>p(266)(98),Cin=>p(267)(98),clock=>clock,reset=>reset,s=>p(306)(98),cout=>p(307)(99));
FA_ff_11193:FAff port map(x=>p(265)(99),y=>p(266)(99),Cin=>p(267)(99),clock=>clock,reset=>reset,s=>p(306)(99),cout=>p(307)(100));
FA_ff_11194:FAff port map(x=>p(265)(100),y=>p(266)(100),Cin=>p(267)(100),clock=>clock,reset=>reset,s=>p(306)(100),cout=>p(307)(101));
FA_ff_11195:FAff port map(x=>p(265)(101),y=>p(266)(101),Cin=>p(267)(101),clock=>clock,reset=>reset,s=>p(306)(101),cout=>p(307)(102));
FA_ff_11196:FAff port map(x=>p(265)(102),y=>p(266)(102),Cin=>p(267)(102),clock=>clock,reset=>reset,s=>p(306)(102),cout=>p(307)(103));
FA_ff_11197:FAff port map(x=>p(265)(103),y=>p(266)(103),Cin=>p(267)(103),clock=>clock,reset=>reset,s=>p(306)(103),cout=>p(307)(104));
FA_ff_11198:FAff port map(x=>p(265)(104),y=>p(266)(104),Cin=>p(267)(104),clock=>clock,reset=>reset,s=>p(306)(104),cout=>p(307)(105));
FA_ff_11199:FAff port map(x=>p(265)(105),y=>p(266)(105),Cin=>p(267)(105),clock=>clock,reset=>reset,s=>p(306)(105),cout=>p(307)(106));
FA_ff_11200:FAff port map(x=>p(265)(106),y=>p(266)(106),Cin=>p(267)(106),clock=>clock,reset=>reset,s=>p(306)(106),cout=>p(307)(107));
FA_ff_11201:FAff port map(x=>p(265)(107),y=>p(266)(107),Cin=>p(267)(107),clock=>clock,reset=>reset,s=>p(306)(107),cout=>p(307)(108));
FA_ff_11202:FAff port map(x=>p(265)(108),y=>p(266)(108),Cin=>p(267)(108),clock=>clock,reset=>reset,s=>p(306)(108),cout=>p(307)(109));
FA_ff_11203:FAff port map(x=>p(265)(109),y=>p(266)(109),Cin=>p(267)(109),clock=>clock,reset=>reset,s=>p(306)(109),cout=>p(307)(110));
FA_ff_11204:FAff port map(x=>p(265)(110),y=>p(266)(110),Cin=>p(267)(110),clock=>clock,reset=>reset,s=>p(306)(110),cout=>p(307)(111));
FA_ff_11205:FAff port map(x=>p(265)(111),y=>p(266)(111),Cin=>p(267)(111),clock=>clock,reset=>reset,s=>p(306)(111),cout=>p(307)(112));
FA_ff_11206:FAff port map(x=>p(265)(112),y=>p(266)(112),Cin=>p(267)(112),clock=>clock,reset=>reset,s=>p(306)(112),cout=>p(307)(113));
FA_ff_11207:FAff port map(x=>p(265)(113),y=>p(266)(113),Cin=>p(267)(113),clock=>clock,reset=>reset,s=>p(306)(113),cout=>p(307)(114));
FA_ff_11208:FAff port map(x=>p(265)(114),y=>p(266)(114),Cin=>p(267)(114),clock=>clock,reset=>reset,s=>p(306)(114),cout=>p(307)(115));
FA_ff_11209:FAff port map(x=>p(265)(115),y=>p(266)(115),Cin=>p(267)(115),clock=>clock,reset=>reset,s=>p(306)(115),cout=>p(307)(116));
FA_ff_11210:FAff port map(x=>p(265)(116),y=>p(266)(116),Cin=>p(267)(116),clock=>clock,reset=>reset,s=>p(306)(116),cout=>p(307)(117));
FA_ff_11211:FAff port map(x=>p(265)(117),y=>p(266)(117),Cin=>p(267)(117),clock=>clock,reset=>reset,s=>p(306)(117),cout=>p(307)(118));
FA_ff_11212:FAff port map(x=>p(265)(118),y=>p(266)(118),Cin=>p(267)(118),clock=>clock,reset=>reset,s=>p(306)(118),cout=>p(307)(119));
FA_ff_11213:FAff port map(x=>p(265)(119),y=>p(266)(119),Cin=>p(267)(119),clock=>clock,reset=>reset,s=>p(306)(119),cout=>p(307)(120));
FA_ff_11214:FAff port map(x=>p(265)(120),y=>p(266)(120),Cin=>p(267)(120),clock=>clock,reset=>reset,s=>p(306)(120),cout=>p(307)(121));
FA_ff_11215:FAff port map(x=>p(265)(121),y=>p(266)(121),Cin=>p(267)(121),clock=>clock,reset=>reset,s=>p(306)(121),cout=>p(307)(122));
FA_ff_11216:FAff port map(x=>p(265)(122),y=>p(266)(122),Cin=>p(267)(122),clock=>clock,reset=>reset,s=>p(306)(122),cout=>p(307)(123));
FA_ff_11217:FAff port map(x=>p(265)(123),y=>p(266)(123),Cin=>p(267)(123),clock=>clock,reset=>reset,s=>p(306)(123),cout=>p(307)(124));
FA_ff_11218:FAff port map(x=>p(265)(124),y=>p(266)(124),Cin=>p(267)(124),clock=>clock,reset=>reset,s=>p(306)(124),cout=>p(307)(125));
FA_ff_11219:FAff port map(x=>p(265)(125),y=>p(266)(125),Cin=>p(267)(125),clock=>clock,reset=>reset,s=>p(306)(125),cout=>p(307)(126));
FA_ff_11220:FAff port map(x=>p(265)(126),y=>p(266)(126),Cin=>p(267)(126),clock=>clock,reset=>reset,s=>p(306)(126),cout=>p(307)(127));
FA_ff_11221:FAff port map(x=>p(265)(127),y=>p(266)(127),Cin=>p(267)(127),clock=>clock,reset=>reset,s=>p(306)(127),cout=>p(307)(128));
FA_ff_11222:FAff port map(x=>p(265)(128),y=>p(266)(128),Cin=>p(267)(128),clock=>clock,reset=>reset,s=>p(306)(128),cout=>p(307)(129));
p(306)(129)<=p(265)(129);
HA_ff_50:HAff port map(x=>p(268)(0),y=>p(270)(0),clock=>clock,reset=>reset,s=>p(308)(0),c=>p(309)(1));
HA_ff_51:HAff port map(x=>p(268)(1),y=>p(270)(1),clock=>clock,reset=>reset,s=>p(308)(1),c=>p(309)(2));
FA_ff_11223:FAff port map(x=>p(268)(2),y=>p(269)(2),Cin=>p(270)(2),clock=>clock,reset=>reset,s=>p(308)(2),cout=>p(309)(3));
FA_ff_11224:FAff port map(x=>p(268)(3),y=>p(269)(3),Cin=>p(270)(3),clock=>clock,reset=>reset,s=>p(308)(3),cout=>p(309)(4));
FA_ff_11225:FAff port map(x=>p(268)(4),y=>p(269)(4),Cin=>p(270)(4),clock=>clock,reset=>reset,s=>p(308)(4),cout=>p(309)(5));
FA_ff_11226:FAff port map(x=>p(268)(5),y=>p(269)(5),Cin=>p(270)(5),clock=>clock,reset=>reset,s=>p(308)(5),cout=>p(309)(6));
FA_ff_11227:FAff port map(x=>p(268)(6),y=>p(269)(6),Cin=>p(270)(6),clock=>clock,reset=>reset,s=>p(308)(6),cout=>p(309)(7));
FA_ff_11228:FAff port map(x=>p(268)(7),y=>p(269)(7),Cin=>p(270)(7),clock=>clock,reset=>reset,s=>p(308)(7),cout=>p(309)(8));
FA_ff_11229:FAff port map(x=>p(268)(8),y=>p(269)(8),Cin=>p(270)(8),clock=>clock,reset=>reset,s=>p(308)(8),cout=>p(309)(9));
FA_ff_11230:FAff port map(x=>p(268)(9),y=>p(269)(9),Cin=>p(270)(9),clock=>clock,reset=>reset,s=>p(308)(9),cout=>p(309)(10));
FA_ff_11231:FAff port map(x=>p(268)(10),y=>p(269)(10),Cin=>p(270)(10),clock=>clock,reset=>reset,s=>p(308)(10),cout=>p(309)(11));
FA_ff_11232:FAff port map(x=>p(268)(11),y=>p(269)(11),Cin=>p(270)(11),clock=>clock,reset=>reset,s=>p(308)(11),cout=>p(309)(12));
FA_ff_11233:FAff port map(x=>p(268)(12),y=>p(269)(12),Cin=>p(270)(12),clock=>clock,reset=>reset,s=>p(308)(12),cout=>p(309)(13));
FA_ff_11234:FAff port map(x=>p(268)(13),y=>p(269)(13),Cin=>p(270)(13),clock=>clock,reset=>reset,s=>p(308)(13),cout=>p(309)(14));
FA_ff_11235:FAff port map(x=>p(268)(14),y=>p(269)(14),Cin=>p(270)(14),clock=>clock,reset=>reset,s=>p(308)(14),cout=>p(309)(15));
FA_ff_11236:FAff port map(x=>p(268)(15),y=>p(269)(15),Cin=>p(270)(15),clock=>clock,reset=>reset,s=>p(308)(15),cout=>p(309)(16));
FA_ff_11237:FAff port map(x=>p(268)(16),y=>p(269)(16),Cin=>p(270)(16),clock=>clock,reset=>reset,s=>p(308)(16),cout=>p(309)(17));
FA_ff_11238:FAff port map(x=>p(268)(17),y=>p(269)(17),Cin=>p(270)(17),clock=>clock,reset=>reset,s=>p(308)(17),cout=>p(309)(18));
FA_ff_11239:FAff port map(x=>p(268)(18),y=>p(269)(18),Cin=>p(270)(18),clock=>clock,reset=>reset,s=>p(308)(18),cout=>p(309)(19));
FA_ff_11240:FAff port map(x=>p(268)(19),y=>p(269)(19),Cin=>p(270)(19),clock=>clock,reset=>reset,s=>p(308)(19),cout=>p(309)(20));
FA_ff_11241:FAff port map(x=>p(268)(20),y=>p(269)(20),Cin=>p(270)(20),clock=>clock,reset=>reset,s=>p(308)(20),cout=>p(309)(21));
FA_ff_11242:FAff port map(x=>p(268)(21),y=>p(269)(21),Cin=>p(270)(21),clock=>clock,reset=>reset,s=>p(308)(21),cout=>p(309)(22));
FA_ff_11243:FAff port map(x=>p(268)(22),y=>p(269)(22),Cin=>p(270)(22),clock=>clock,reset=>reset,s=>p(308)(22),cout=>p(309)(23));
FA_ff_11244:FAff port map(x=>p(268)(23),y=>p(269)(23),Cin=>p(270)(23),clock=>clock,reset=>reset,s=>p(308)(23),cout=>p(309)(24));
FA_ff_11245:FAff port map(x=>p(268)(24),y=>p(269)(24),Cin=>p(270)(24),clock=>clock,reset=>reset,s=>p(308)(24),cout=>p(309)(25));
FA_ff_11246:FAff port map(x=>p(268)(25),y=>p(269)(25),Cin=>p(270)(25),clock=>clock,reset=>reset,s=>p(308)(25),cout=>p(309)(26));
FA_ff_11247:FAff port map(x=>p(268)(26),y=>p(269)(26),Cin=>p(270)(26),clock=>clock,reset=>reset,s=>p(308)(26),cout=>p(309)(27));
FA_ff_11248:FAff port map(x=>p(268)(27),y=>p(269)(27),Cin=>p(270)(27),clock=>clock,reset=>reset,s=>p(308)(27),cout=>p(309)(28));
FA_ff_11249:FAff port map(x=>p(268)(28),y=>p(269)(28),Cin=>p(270)(28),clock=>clock,reset=>reset,s=>p(308)(28),cout=>p(309)(29));
FA_ff_11250:FAff port map(x=>p(268)(29),y=>p(269)(29),Cin=>p(270)(29),clock=>clock,reset=>reset,s=>p(308)(29),cout=>p(309)(30));
FA_ff_11251:FAff port map(x=>p(268)(30),y=>p(269)(30),Cin=>p(270)(30),clock=>clock,reset=>reset,s=>p(308)(30),cout=>p(309)(31));
FA_ff_11252:FAff port map(x=>p(268)(31),y=>p(269)(31),Cin=>p(270)(31),clock=>clock,reset=>reset,s=>p(308)(31),cout=>p(309)(32));
FA_ff_11253:FAff port map(x=>p(268)(32),y=>p(269)(32),Cin=>p(270)(32),clock=>clock,reset=>reset,s=>p(308)(32),cout=>p(309)(33));
FA_ff_11254:FAff port map(x=>p(268)(33),y=>p(269)(33),Cin=>p(270)(33),clock=>clock,reset=>reset,s=>p(308)(33),cout=>p(309)(34));
FA_ff_11255:FAff port map(x=>p(268)(34),y=>p(269)(34),Cin=>p(270)(34),clock=>clock,reset=>reset,s=>p(308)(34),cout=>p(309)(35));
FA_ff_11256:FAff port map(x=>p(268)(35),y=>p(269)(35),Cin=>p(270)(35),clock=>clock,reset=>reset,s=>p(308)(35),cout=>p(309)(36));
FA_ff_11257:FAff port map(x=>p(268)(36),y=>p(269)(36),Cin=>p(270)(36),clock=>clock,reset=>reset,s=>p(308)(36),cout=>p(309)(37));
FA_ff_11258:FAff port map(x=>p(268)(37),y=>p(269)(37),Cin=>p(270)(37),clock=>clock,reset=>reset,s=>p(308)(37),cout=>p(309)(38));
FA_ff_11259:FAff port map(x=>p(268)(38),y=>p(269)(38),Cin=>p(270)(38),clock=>clock,reset=>reset,s=>p(308)(38),cout=>p(309)(39));
FA_ff_11260:FAff port map(x=>p(268)(39),y=>p(269)(39),Cin=>p(270)(39),clock=>clock,reset=>reset,s=>p(308)(39),cout=>p(309)(40));
FA_ff_11261:FAff port map(x=>p(268)(40),y=>p(269)(40),Cin=>p(270)(40),clock=>clock,reset=>reset,s=>p(308)(40),cout=>p(309)(41));
FA_ff_11262:FAff port map(x=>p(268)(41),y=>p(269)(41),Cin=>p(270)(41),clock=>clock,reset=>reset,s=>p(308)(41),cout=>p(309)(42));
FA_ff_11263:FAff port map(x=>p(268)(42),y=>p(269)(42),Cin=>p(270)(42),clock=>clock,reset=>reset,s=>p(308)(42),cout=>p(309)(43));
FA_ff_11264:FAff port map(x=>p(268)(43),y=>p(269)(43),Cin=>p(270)(43),clock=>clock,reset=>reset,s=>p(308)(43),cout=>p(309)(44));
FA_ff_11265:FAff port map(x=>p(268)(44),y=>p(269)(44),Cin=>p(270)(44),clock=>clock,reset=>reset,s=>p(308)(44),cout=>p(309)(45));
FA_ff_11266:FAff port map(x=>p(268)(45),y=>p(269)(45),Cin=>p(270)(45),clock=>clock,reset=>reset,s=>p(308)(45),cout=>p(309)(46));
FA_ff_11267:FAff port map(x=>p(268)(46),y=>p(269)(46),Cin=>p(270)(46),clock=>clock,reset=>reset,s=>p(308)(46),cout=>p(309)(47));
FA_ff_11268:FAff port map(x=>p(268)(47),y=>p(269)(47),Cin=>p(270)(47),clock=>clock,reset=>reset,s=>p(308)(47),cout=>p(309)(48));
FA_ff_11269:FAff port map(x=>p(268)(48),y=>p(269)(48),Cin=>p(270)(48),clock=>clock,reset=>reset,s=>p(308)(48),cout=>p(309)(49));
FA_ff_11270:FAff port map(x=>p(268)(49),y=>p(269)(49),Cin=>p(270)(49),clock=>clock,reset=>reset,s=>p(308)(49),cout=>p(309)(50));
FA_ff_11271:FAff port map(x=>p(268)(50),y=>p(269)(50),Cin=>p(270)(50),clock=>clock,reset=>reset,s=>p(308)(50),cout=>p(309)(51));
FA_ff_11272:FAff port map(x=>p(268)(51),y=>p(269)(51),Cin=>p(270)(51),clock=>clock,reset=>reset,s=>p(308)(51),cout=>p(309)(52));
FA_ff_11273:FAff port map(x=>p(268)(52),y=>p(269)(52),Cin=>p(270)(52),clock=>clock,reset=>reset,s=>p(308)(52),cout=>p(309)(53));
FA_ff_11274:FAff port map(x=>p(268)(53),y=>p(269)(53),Cin=>p(270)(53),clock=>clock,reset=>reset,s=>p(308)(53),cout=>p(309)(54));
FA_ff_11275:FAff port map(x=>p(268)(54),y=>p(269)(54),Cin=>p(270)(54),clock=>clock,reset=>reset,s=>p(308)(54),cout=>p(309)(55));
FA_ff_11276:FAff port map(x=>p(268)(55),y=>p(269)(55),Cin=>p(270)(55),clock=>clock,reset=>reset,s=>p(308)(55),cout=>p(309)(56));
FA_ff_11277:FAff port map(x=>p(268)(56),y=>p(269)(56),Cin=>p(270)(56),clock=>clock,reset=>reset,s=>p(308)(56),cout=>p(309)(57));
FA_ff_11278:FAff port map(x=>p(268)(57),y=>p(269)(57),Cin=>p(270)(57),clock=>clock,reset=>reset,s=>p(308)(57),cout=>p(309)(58));
FA_ff_11279:FAff port map(x=>p(268)(58),y=>p(269)(58),Cin=>p(270)(58),clock=>clock,reset=>reset,s=>p(308)(58),cout=>p(309)(59));
FA_ff_11280:FAff port map(x=>p(268)(59),y=>p(269)(59),Cin=>p(270)(59),clock=>clock,reset=>reset,s=>p(308)(59),cout=>p(309)(60));
FA_ff_11281:FAff port map(x=>p(268)(60),y=>p(269)(60),Cin=>p(270)(60),clock=>clock,reset=>reset,s=>p(308)(60),cout=>p(309)(61));
FA_ff_11282:FAff port map(x=>p(268)(61),y=>p(269)(61),Cin=>p(270)(61),clock=>clock,reset=>reset,s=>p(308)(61),cout=>p(309)(62));
FA_ff_11283:FAff port map(x=>p(268)(62),y=>p(269)(62),Cin=>p(270)(62),clock=>clock,reset=>reset,s=>p(308)(62),cout=>p(309)(63));
FA_ff_11284:FAff port map(x=>p(268)(63),y=>p(269)(63),Cin=>p(270)(63),clock=>clock,reset=>reset,s=>p(308)(63),cout=>p(309)(64));
FA_ff_11285:FAff port map(x=>p(268)(64),y=>p(269)(64),Cin=>p(270)(64),clock=>clock,reset=>reset,s=>p(308)(64),cout=>p(309)(65));
FA_ff_11286:FAff port map(x=>p(268)(65),y=>p(269)(65),Cin=>p(270)(65),clock=>clock,reset=>reset,s=>p(308)(65),cout=>p(309)(66));
FA_ff_11287:FAff port map(x=>p(268)(66),y=>p(269)(66),Cin=>p(270)(66),clock=>clock,reset=>reset,s=>p(308)(66),cout=>p(309)(67));
FA_ff_11288:FAff port map(x=>p(268)(67),y=>p(269)(67),Cin=>p(270)(67),clock=>clock,reset=>reset,s=>p(308)(67),cout=>p(309)(68));
FA_ff_11289:FAff port map(x=>p(268)(68),y=>p(269)(68),Cin=>p(270)(68),clock=>clock,reset=>reset,s=>p(308)(68),cout=>p(309)(69));
FA_ff_11290:FAff port map(x=>p(268)(69),y=>p(269)(69),Cin=>p(270)(69),clock=>clock,reset=>reset,s=>p(308)(69),cout=>p(309)(70));
FA_ff_11291:FAff port map(x=>p(268)(70),y=>p(269)(70),Cin=>p(270)(70),clock=>clock,reset=>reset,s=>p(308)(70),cout=>p(309)(71));
FA_ff_11292:FAff port map(x=>p(268)(71),y=>p(269)(71),Cin=>p(270)(71),clock=>clock,reset=>reset,s=>p(308)(71),cout=>p(309)(72));
FA_ff_11293:FAff port map(x=>p(268)(72),y=>p(269)(72),Cin=>p(270)(72),clock=>clock,reset=>reset,s=>p(308)(72),cout=>p(309)(73));
FA_ff_11294:FAff port map(x=>p(268)(73),y=>p(269)(73),Cin=>p(270)(73),clock=>clock,reset=>reset,s=>p(308)(73),cout=>p(309)(74));
FA_ff_11295:FAff port map(x=>p(268)(74),y=>p(269)(74),Cin=>p(270)(74),clock=>clock,reset=>reset,s=>p(308)(74),cout=>p(309)(75));
FA_ff_11296:FAff port map(x=>p(268)(75),y=>p(269)(75),Cin=>p(270)(75),clock=>clock,reset=>reset,s=>p(308)(75),cout=>p(309)(76));
FA_ff_11297:FAff port map(x=>p(268)(76),y=>p(269)(76),Cin=>p(270)(76),clock=>clock,reset=>reset,s=>p(308)(76),cout=>p(309)(77));
FA_ff_11298:FAff port map(x=>p(268)(77),y=>p(269)(77),Cin=>p(270)(77),clock=>clock,reset=>reset,s=>p(308)(77),cout=>p(309)(78));
FA_ff_11299:FAff port map(x=>p(268)(78),y=>p(269)(78),Cin=>p(270)(78),clock=>clock,reset=>reset,s=>p(308)(78),cout=>p(309)(79));
FA_ff_11300:FAff port map(x=>p(268)(79),y=>p(269)(79),Cin=>p(270)(79),clock=>clock,reset=>reset,s=>p(308)(79),cout=>p(309)(80));
FA_ff_11301:FAff port map(x=>p(268)(80),y=>p(269)(80),Cin=>p(270)(80),clock=>clock,reset=>reset,s=>p(308)(80),cout=>p(309)(81));
FA_ff_11302:FAff port map(x=>p(268)(81),y=>p(269)(81),Cin=>p(270)(81),clock=>clock,reset=>reset,s=>p(308)(81),cout=>p(309)(82));
FA_ff_11303:FAff port map(x=>p(268)(82),y=>p(269)(82),Cin=>p(270)(82),clock=>clock,reset=>reset,s=>p(308)(82),cout=>p(309)(83));
FA_ff_11304:FAff port map(x=>p(268)(83),y=>p(269)(83),Cin=>p(270)(83),clock=>clock,reset=>reset,s=>p(308)(83),cout=>p(309)(84));
FA_ff_11305:FAff port map(x=>p(268)(84),y=>p(269)(84),Cin=>p(270)(84),clock=>clock,reset=>reset,s=>p(308)(84),cout=>p(309)(85));
FA_ff_11306:FAff port map(x=>p(268)(85),y=>p(269)(85),Cin=>p(270)(85),clock=>clock,reset=>reset,s=>p(308)(85),cout=>p(309)(86));
FA_ff_11307:FAff port map(x=>p(268)(86),y=>p(269)(86),Cin=>p(270)(86),clock=>clock,reset=>reset,s=>p(308)(86),cout=>p(309)(87));
FA_ff_11308:FAff port map(x=>p(268)(87),y=>p(269)(87),Cin=>p(270)(87),clock=>clock,reset=>reset,s=>p(308)(87),cout=>p(309)(88));
FA_ff_11309:FAff port map(x=>p(268)(88),y=>p(269)(88),Cin=>p(270)(88),clock=>clock,reset=>reset,s=>p(308)(88),cout=>p(309)(89));
FA_ff_11310:FAff port map(x=>p(268)(89),y=>p(269)(89),Cin=>p(270)(89),clock=>clock,reset=>reset,s=>p(308)(89),cout=>p(309)(90));
FA_ff_11311:FAff port map(x=>p(268)(90),y=>p(269)(90),Cin=>p(270)(90),clock=>clock,reset=>reset,s=>p(308)(90),cout=>p(309)(91));
FA_ff_11312:FAff port map(x=>p(268)(91),y=>p(269)(91),Cin=>p(270)(91),clock=>clock,reset=>reset,s=>p(308)(91),cout=>p(309)(92));
FA_ff_11313:FAff port map(x=>p(268)(92),y=>p(269)(92),Cin=>p(270)(92),clock=>clock,reset=>reset,s=>p(308)(92),cout=>p(309)(93));
FA_ff_11314:FAff port map(x=>p(268)(93),y=>p(269)(93),Cin=>p(270)(93),clock=>clock,reset=>reset,s=>p(308)(93),cout=>p(309)(94));
FA_ff_11315:FAff port map(x=>p(268)(94),y=>p(269)(94),Cin=>p(270)(94),clock=>clock,reset=>reset,s=>p(308)(94),cout=>p(309)(95));
FA_ff_11316:FAff port map(x=>p(268)(95),y=>p(269)(95),Cin=>p(270)(95),clock=>clock,reset=>reset,s=>p(308)(95),cout=>p(309)(96));
FA_ff_11317:FAff port map(x=>p(268)(96),y=>p(269)(96),Cin=>p(270)(96),clock=>clock,reset=>reset,s=>p(308)(96),cout=>p(309)(97));
FA_ff_11318:FAff port map(x=>p(268)(97),y=>p(269)(97),Cin=>p(270)(97),clock=>clock,reset=>reset,s=>p(308)(97),cout=>p(309)(98));
FA_ff_11319:FAff port map(x=>p(268)(98),y=>p(269)(98),Cin=>p(270)(98),clock=>clock,reset=>reset,s=>p(308)(98),cout=>p(309)(99));
FA_ff_11320:FAff port map(x=>p(268)(99),y=>p(269)(99),Cin=>p(270)(99),clock=>clock,reset=>reset,s=>p(308)(99),cout=>p(309)(100));
FA_ff_11321:FAff port map(x=>p(268)(100),y=>p(269)(100),Cin=>p(270)(100),clock=>clock,reset=>reset,s=>p(308)(100),cout=>p(309)(101));
FA_ff_11322:FAff port map(x=>p(268)(101),y=>p(269)(101),Cin=>p(270)(101),clock=>clock,reset=>reset,s=>p(308)(101),cout=>p(309)(102));
FA_ff_11323:FAff port map(x=>p(268)(102),y=>p(269)(102),Cin=>p(270)(102),clock=>clock,reset=>reset,s=>p(308)(102),cout=>p(309)(103));
FA_ff_11324:FAff port map(x=>p(268)(103),y=>p(269)(103),Cin=>p(270)(103),clock=>clock,reset=>reset,s=>p(308)(103),cout=>p(309)(104));
FA_ff_11325:FAff port map(x=>p(268)(104),y=>p(269)(104),Cin=>p(270)(104),clock=>clock,reset=>reset,s=>p(308)(104),cout=>p(309)(105));
FA_ff_11326:FAff port map(x=>p(268)(105),y=>p(269)(105),Cin=>p(270)(105),clock=>clock,reset=>reset,s=>p(308)(105),cout=>p(309)(106));
FA_ff_11327:FAff port map(x=>p(268)(106),y=>p(269)(106),Cin=>p(270)(106),clock=>clock,reset=>reset,s=>p(308)(106),cout=>p(309)(107));
FA_ff_11328:FAff port map(x=>p(268)(107),y=>p(269)(107),Cin=>p(270)(107),clock=>clock,reset=>reset,s=>p(308)(107),cout=>p(309)(108));
FA_ff_11329:FAff port map(x=>p(268)(108),y=>p(269)(108),Cin=>p(270)(108),clock=>clock,reset=>reset,s=>p(308)(108),cout=>p(309)(109));
FA_ff_11330:FAff port map(x=>p(268)(109),y=>p(269)(109),Cin=>p(270)(109),clock=>clock,reset=>reset,s=>p(308)(109),cout=>p(309)(110));
FA_ff_11331:FAff port map(x=>p(268)(110),y=>p(269)(110),Cin=>p(270)(110),clock=>clock,reset=>reset,s=>p(308)(110),cout=>p(309)(111));
FA_ff_11332:FAff port map(x=>p(268)(111),y=>p(269)(111),Cin=>p(270)(111),clock=>clock,reset=>reset,s=>p(308)(111),cout=>p(309)(112));
FA_ff_11333:FAff port map(x=>p(268)(112),y=>p(269)(112),Cin=>p(270)(112),clock=>clock,reset=>reset,s=>p(308)(112),cout=>p(309)(113));
FA_ff_11334:FAff port map(x=>p(268)(113),y=>p(269)(113),Cin=>p(270)(113),clock=>clock,reset=>reset,s=>p(308)(113),cout=>p(309)(114));
FA_ff_11335:FAff port map(x=>p(268)(114),y=>p(269)(114),Cin=>p(270)(114),clock=>clock,reset=>reset,s=>p(308)(114),cout=>p(309)(115));
FA_ff_11336:FAff port map(x=>p(268)(115),y=>p(269)(115),Cin=>p(270)(115),clock=>clock,reset=>reset,s=>p(308)(115),cout=>p(309)(116));
FA_ff_11337:FAff port map(x=>p(268)(116),y=>p(269)(116),Cin=>p(270)(116),clock=>clock,reset=>reset,s=>p(308)(116),cout=>p(309)(117));
FA_ff_11338:FAff port map(x=>p(268)(117),y=>p(269)(117),Cin=>p(270)(117),clock=>clock,reset=>reset,s=>p(308)(117),cout=>p(309)(118));
FA_ff_11339:FAff port map(x=>p(268)(118),y=>p(269)(118),Cin=>p(270)(118),clock=>clock,reset=>reset,s=>p(308)(118),cout=>p(309)(119));
FA_ff_11340:FAff port map(x=>p(268)(119),y=>p(269)(119),Cin=>p(270)(119),clock=>clock,reset=>reset,s=>p(308)(119),cout=>p(309)(120));
FA_ff_11341:FAff port map(x=>p(268)(120),y=>p(269)(120),Cin=>p(270)(120),clock=>clock,reset=>reset,s=>p(308)(120),cout=>p(309)(121));
FA_ff_11342:FAff port map(x=>p(268)(121),y=>p(269)(121),Cin=>p(270)(121),clock=>clock,reset=>reset,s=>p(308)(121),cout=>p(309)(122));
FA_ff_11343:FAff port map(x=>p(268)(122),y=>p(269)(122),Cin=>p(270)(122),clock=>clock,reset=>reset,s=>p(308)(122),cout=>p(309)(123));
FA_ff_11344:FAff port map(x=>p(268)(123),y=>p(269)(123),Cin=>p(270)(123),clock=>clock,reset=>reset,s=>p(308)(123),cout=>p(309)(124));
FA_ff_11345:FAff port map(x=>p(268)(124),y=>p(269)(124),Cin=>p(270)(124),clock=>clock,reset=>reset,s=>p(308)(124),cout=>p(309)(125));
FA_ff_11346:FAff port map(x=>p(268)(125),y=>p(269)(125),Cin=>p(270)(125),clock=>clock,reset=>reset,s=>p(308)(125),cout=>p(309)(126));
FA_ff_11347:FAff port map(x=>p(268)(126),y=>p(269)(126),Cin=>p(270)(126),clock=>clock,reset=>reset,s=>p(308)(126),cout=>p(309)(127));
FA_ff_11348:FAff port map(x=>p(268)(127),y=>p(269)(127),Cin=>p(270)(127),clock=>clock,reset=>reset,s=>p(308)(127),cout=>p(309)(128));
HA_ff_52:HAff port map(x=>p(268)(128),y=>p(269)(128),clock=>clock,reset=>reset,s=>p(308)(128),c=>p(309)(129));
p(308)(129)<=p(269)(129);
p(310)(0)<=p(271)(0);
p(310)(1)<=p(271)(1);
p(310)(2)<=p(271)(2);
p(310)(3)<=p(271)(3);
p(310)(4)<=p(271)(4);
p(310)(5)<=p(271)(5);
p(310)(6)<=p(271)(6);
p(310)(7)<=p(271)(7);
p(310)(8)<=p(271)(8);
p(310)(9)<=p(271)(9);
p(310)(10)<=p(271)(10);
p(310)(11)<=p(271)(11);
p(310)(12)<=p(271)(12);
p(310)(13)<=p(271)(13);
p(310)(14)<=p(271)(14);
p(310)(15)<=p(271)(15);
p(310)(16)<=p(271)(16);
p(310)(17)<=p(271)(17);
p(310)(18)<=p(271)(18);
p(310)(19)<=p(271)(19);
p(310)(20)<=p(271)(20);
p(310)(21)<=p(271)(21);
p(310)(22)<=p(271)(22);
p(310)(23)<=p(271)(23);
p(310)(24)<=p(271)(24);
p(310)(25)<=p(271)(25);
p(310)(26)<=p(271)(26);
p(310)(27)<=p(271)(27);
p(310)(28)<=p(271)(28);
p(310)(29)<=p(271)(29);
p(310)(30)<=p(271)(30);
p(310)(31)<=p(271)(31);
p(310)(32)<=p(271)(32);
p(310)(33)<=p(271)(33);
p(310)(34)<=p(271)(34);
p(310)(35)<=p(271)(35);
p(310)(36)<=p(271)(36);
p(310)(37)<=p(271)(37);
p(310)(38)<=p(271)(38);
p(310)(39)<=p(271)(39);
p(310)(40)<=p(271)(40);
p(310)(41)<=p(271)(41);
p(310)(42)<=p(271)(42);
p(310)(43)<=p(271)(43);
p(310)(44)<=p(271)(44);
p(310)(45)<=p(271)(45);
p(310)(46)<=p(271)(46);
p(310)(47)<=p(271)(47);
p(310)(48)<=p(271)(48);
p(310)(49)<=p(271)(49);
p(310)(50)<=p(271)(50);
p(310)(51)<=p(271)(51);
p(310)(52)<=p(271)(52);
p(310)(53)<=p(271)(53);
p(310)(54)<=p(271)(54);
p(310)(55)<=p(271)(55);
p(310)(56)<=p(271)(56);
p(310)(57)<=p(271)(57);
p(310)(58)<=p(271)(58);
p(310)(59)<=p(271)(59);
p(310)(60)<=p(271)(60);
p(310)(61)<=p(271)(61);
p(310)(62)<=p(271)(62);
p(310)(63)<=p(271)(63);
p(310)(64)<=p(271)(64);
p(310)(65)<=p(271)(65);
p(310)(66)<=p(271)(66);
p(310)(67)<=p(271)(67);
p(310)(68)<=p(271)(68);
p(310)(69)<=p(271)(69);
p(310)(70)<=p(271)(70);
p(310)(71)<=p(271)(71);
p(310)(72)<=p(271)(72);
p(310)(73)<=p(271)(73);
p(310)(74)<=p(271)(74);
p(310)(75)<=p(271)(75);
p(310)(76)<=p(271)(76);
p(310)(77)<=p(271)(77);
p(310)(78)<=p(271)(78);
p(310)(79)<=p(271)(79);
p(310)(80)<=p(271)(80);
p(310)(81)<=p(271)(81);
p(310)(82)<=p(271)(82);
p(310)(83)<=p(271)(83);
p(310)(84)<=p(271)(84);
p(310)(85)<=p(271)(85);
p(310)(86)<=p(271)(86);
p(310)(87)<=p(271)(87);
p(310)(88)<=p(271)(88);
p(310)(89)<=p(271)(89);
p(310)(90)<=p(271)(90);
p(310)(91)<=p(271)(91);
p(310)(92)<=p(271)(92);
p(310)(93)<=p(271)(93);
p(310)(94)<=p(271)(94);
p(310)(95)<=p(271)(95);
p(310)(96)<=p(271)(96);
p(310)(97)<=p(271)(97);
p(310)(98)<=p(271)(98);
p(310)(99)<=p(271)(99);
p(310)(100)<=p(271)(100);
p(310)(101)<=p(271)(101);
p(310)(102)<=p(271)(102);
p(310)(103)<=p(271)(103);
p(310)(104)<=p(271)(104);
p(310)(105)<=p(271)(105);
p(310)(106)<=p(271)(106);
p(310)(107)<=p(271)(107);
p(310)(108)<=p(271)(108);
p(310)(109)<=p(271)(109);
p(310)(110)<=p(271)(110);
p(310)(111)<=p(271)(111);
p(310)(112)<=p(271)(112);
p(310)(113)<=p(271)(113);
p(310)(114)<=p(271)(114);
p(310)(115)<=p(271)(115);
p(310)(116)<=p(271)(116);
p(310)(117)<=p(271)(117);
p(310)(118)<=p(271)(118);
p(310)(119)<=p(271)(119);
p(310)(120)<=p(271)(120);
p(310)(121)<=p(271)(121);
p(310)(122)<=p(271)(122);
p(310)(123)<=p(271)(123);
p(310)(124)<=p(271)(124);
p(310)(125)<=p(271)(125);
p(310)(126)<=p(271)(126);
p(310)(127)<=p(271)(127);
p(310)(128)<=p(271)(128);
p(310)(129)<=p(271)(129);
p(310)(130)<=p(271)(130);
p(310)(131)<=p(271)(131);
p(310)(132)<=p(271)(132);
p(310)(133)<=p(271)(133);
p(310)(134)<=p(271)(134);
HA_ff_53:HAff port map(x=>p(272)(0),y=>p(274)(0),clock=>clock,reset=>reset,s=>p(311)(0),c=>p(312)(1));
FA_ff_11349:FAff port map(x=>p(272)(1),y=>p(273)(1),Cin=>p(274)(1),clock=>clock,reset=>reset,s=>p(311)(1),cout=>p(312)(2));
FA_ff_11350:FAff port map(x=>p(272)(2),y=>p(273)(2),Cin=>p(274)(2),clock=>clock,reset=>reset,s=>p(311)(2),cout=>p(312)(3));
FA_ff_11351:FAff port map(x=>p(272)(3),y=>p(273)(3),Cin=>p(274)(3),clock=>clock,reset=>reset,s=>p(311)(3),cout=>p(312)(4));
FA_ff_11352:FAff port map(x=>p(272)(4),y=>p(273)(4),Cin=>p(274)(4),clock=>clock,reset=>reset,s=>p(311)(4),cout=>p(312)(5));
FA_ff_11353:FAff port map(x=>p(272)(5),y=>p(273)(5),Cin=>p(274)(5),clock=>clock,reset=>reset,s=>p(311)(5),cout=>p(312)(6));
FA_ff_11354:FAff port map(x=>p(272)(6),y=>p(273)(6),Cin=>p(274)(6),clock=>clock,reset=>reset,s=>p(311)(6),cout=>p(312)(7));
FA_ff_11355:FAff port map(x=>p(272)(7),y=>p(273)(7),Cin=>p(274)(7),clock=>clock,reset=>reset,s=>p(311)(7),cout=>p(312)(8));
FA_ff_11356:FAff port map(x=>p(272)(8),y=>p(273)(8),Cin=>p(274)(8),clock=>clock,reset=>reset,s=>p(311)(8),cout=>p(312)(9));
FA_ff_11357:FAff port map(x=>p(272)(9),y=>p(273)(9),Cin=>p(274)(9),clock=>clock,reset=>reset,s=>p(311)(9),cout=>p(312)(10));
FA_ff_11358:FAff port map(x=>p(272)(10),y=>p(273)(10),Cin=>p(274)(10),clock=>clock,reset=>reset,s=>p(311)(10),cout=>p(312)(11));
FA_ff_11359:FAff port map(x=>p(272)(11),y=>p(273)(11),Cin=>p(274)(11),clock=>clock,reset=>reset,s=>p(311)(11),cout=>p(312)(12));
FA_ff_11360:FAff port map(x=>p(272)(12),y=>p(273)(12),Cin=>p(274)(12),clock=>clock,reset=>reset,s=>p(311)(12),cout=>p(312)(13));
FA_ff_11361:FAff port map(x=>p(272)(13),y=>p(273)(13),Cin=>p(274)(13),clock=>clock,reset=>reset,s=>p(311)(13),cout=>p(312)(14));
FA_ff_11362:FAff port map(x=>p(272)(14),y=>p(273)(14),Cin=>p(274)(14),clock=>clock,reset=>reset,s=>p(311)(14),cout=>p(312)(15));
FA_ff_11363:FAff port map(x=>p(272)(15),y=>p(273)(15),Cin=>p(274)(15),clock=>clock,reset=>reset,s=>p(311)(15),cout=>p(312)(16));
FA_ff_11364:FAff port map(x=>p(272)(16),y=>p(273)(16),Cin=>p(274)(16),clock=>clock,reset=>reset,s=>p(311)(16),cout=>p(312)(17));
FA_ff_11365:FAff port map(x=>p(272)(17),y=>p(273)(17),Cin=>p(274)(17),clock=>clock,reset=>reset,s=>p(311)(17),cout=>p(312)(18));
FA_ff_11366:FAff port map(x=>p(272)(18),y=>p(273)(18),Cin=>p(274)(18),clock=>clock,reset=>reset,s=>p(311)(18),cout=>p(312)(19));
FA_ff_11367:FAff port map(x=>p(272)(19),y=>p(273)(19),Cin=>p(274)(19),clock=>clock,reset=>reset,s=>p(311)(19),cout=>p(312)(20));
FA_ff_11368:FAff port map(x=>p(272)(20),y=>p(273)(20),Cin=>p(274)(20),clock=>clock,reset=>reset,s=>p(311)(20),cout=>p(312)(21));
FA_ff_11369:FAff port map(x=>p(272)(21),y=>p(273)(21),Cin=>p(274)(21),clock=>clock,reset=>reset,s=>p(311)(21),cout=>p(312)(22));
FA_ff_11370:FAff port map(x=>p(272)(22),y=>p(273)(22),Cin=>p(274)(22),clock=>clock,reset=>reset,s=>p(311)(22),cout=>p(312)(23));
FA_ff_11371:FAff port map(x=>p(272)(23),y=>p(273)(23),Cin=>p(274)(23),clock=>clock,reset=>reset,s=>p(311)(23),cout=>p(312)(24));
FA_ff_11372:FAff port map(x=>p(272)(24),y=>p(273)(24),Cin=>p(274)(24),clock=>clock,reset=>reset,s=>p(311)(24),cout=>p(312)(25));
FA_ff_11373:FAff port map(x=>p(272)(25),y=>p(273)(25),Cin=>p(274)(25),clock=>clock,reset=>reset,s=>p(311)(25),cout=>p(312)(26));
FA_ff_11374:FAff port map(x=>p(272)(26),y=>p(273)(26),Cin=>p(274)(26),clock=>clock,reset=>reset,s=>p(311)(26),cout=>p(312)(27));
FA_ff_11375:FAff port map(x=>p(272)(27),y=>p(273)(27),Cin=>p(274)(27),clock=>clock,reset=>reset,s=>p(311)(27),cout=>p(312)(28));
FA_ff_11376:FAff port map(x=>p(272)(28),y=>p(273)(28),Cin=>p(274)(28),clock=>clock,reset=>reset,s=>p(311)(28),cout=>p(312)(29));
FA_ff_11377:FAff port map(x=>p(272)(29),y=>p(273)(29),Cin=>p(274)(29),clock=>clock,reset=>reset,s=>p(311)(29),cout=>p(312)(30));
FA_ff_11378:FAff port map(x=>p(272)(30),y=>p(273)(30),Cin=>p(274)(30),clock=>clock,reset=>reset,s=>p(311)(30),cout=>p(312)(31));
FA_ff_11379:FAff port map(x=>p(272)(31),y=>p(273)(31),Cin=>p(274)(31),clock=>clock,reset=>reset,s=>p(311)(31),cout=>p(312)(32));
FA_ff_11380:FAff port map(x=>p(272)(32),y=>p(273)(32),Cin=>p(274)(32),clock=>clock,reset=>reset,s=>p(311)(32),cout=>p(312)(33));
FA_ff_11381:FAff port map(x=>p(272)(33),y=>p(273)(33),Cin=>p(274)(33),clock=>clock,reset=>reset,s=>p(311)(33),cout=>p(312)(34));
FA_ff_11382:FAff port map(x=>p(272)(34),y=>p(273)(34),Cin=>p(274)(34),clock=>clock,reset=>reset,s=>p(311)(34),cout=>p(312)(35));
FA_ff_11383:FAff port map(x=>p(272)(35),y=>p(273)(35),Cin=>p(274)(35),clock=>clock,reset=>reset,s=>p(311)(35),cout=>p(312)(36));
FA_ff_11384:FAff port map(x=>p(272)(36),y=>p(273)(36),Cin=>p(274)(36),clock=>clock,reset=>reset,s=>p(311)(36),cout=>p(312)(37));
FA_ff_11385:FAff port map(x=>p(272)(37),y=>p(273)(37),Cin=>p(274)(37),clock=>clock,reset=>reset,s=>p(311)(37),cout=>p(312)(38));
FA_ff_11386:FAff port map(x=>p(272)(38),y=>p(273)(38),Cin=>p(274)(38),clock=>clock,reset=>reset,s=>p(311)(38),cout=>p(312)(39));
FA_ff_11387:FAff port map(x=>p(272)(39),y=>p(273)(39),Cin=>p(274)(39),clock=>clock,reset=>reset,s=>p(311)(39),cout=>p(312)(40));
FA_ff_11388:FAff port map(x=>p(272)(40),y=>p(273)(40),Cin=>p(274)(40),clock=>clock,reset=>reset,s=>p(311)(40),cout=>p(312)(41));
FA_ff_11389:FAff port map(x=>p(272)(41),y=>p(273)(41),Cin=>p(274)(41),clock=>clock,reset=>reset,s=>p(311)(41),cout=>p(312)(42));
FA_ff_11390:FAff port map(x=>p(272)(42),y=>p(273)(42),Cin=>p(274)(42),clock=>clock,reset=>reset,s=>p(311)(42),cout=>p(312)(43));
FA_ff_11391:FAff port map(x=>p(272)(43),y=>p(273)(43),Cin=>p(274)(43),clock=>clock,reset=>reset,s=>p(311)(43),cout=>p(312)(44));
FA_ff_11392:FAff port map(x=>p(272)(44),y=>p(273)(44),Cin=>p(274)(44),clock=>clock,reset=>reset,s=>p(311)(44),cout=>p(312)(45));
FA_ff_11393:FAff port map(x=>p(272)(45),y=>p(273)(45),Cin=>p(274)(45),clock=>clock,reset=>reset,s=>p(311)(45),cout=>p(312)(46));
FA_ff_11394:FAff port map(x=>p(272)(46),y=>p(273)(46),Cin=>p(274)(46),clock=>clock,reset=>reset,s=>p(311)(46),cout=>p(312)(47));
FA_ff_11395:FAff port map(x=>p(272)(47),y=>p(273)(47),Cin=>p(274)(47),clock=>clock,reset=>reset,s=>p(311)(47),cout=>p(312)(48));
FA_ff_11396:FAff port map(x=>p(272)(48),y=>p(273)(48),Cin=>p(274)(48),clock=>clock,reset=>reset,s=>p(311)(48),cout=>p(312)(49));
FA_ff_11397:FAff port map(x=>p(272)(49),y=>p(273)(49),Cin=>p(274)(49),clock=>clock,reset=>reset,s=>p(311)(49),cout=>p(312)(50));
FA_ff_11398:FAff port map(x=>p(272)(50),y=>p(273)(50),Cin=>p(274)(50),clock=>clock,reset=>reset,s=>p(311)(50),cout=>p(312)(51));
FA_ff_11399:FAff port map(x=>p(272)(51),y=>p(273)(51),Cin=>p(274)(51),clock=>clock,reset=>reset,s=>p(311)(51),cout=>p(312)(52));
FA_ff_11400:FAff port map(x=>p(272)(52),y=>p(273)(52),Cin=>p(274)(52),clock=>clock,reset=>reset,s=>p(311)(52),cout=>p(312)(53));
FA_ff_11401:FAff port map(x=>p(272)(53),y=>p(273)(53),Cin=>p(274)(53),clock=>clock,reset=>reset,s=>p(311)(53),cout=>p(312)(54));
FA_ff_11402:FAff port map(x=>p(272)(54),y=>p(273)(54),Cin=>p(274)(54),clock=>clock,reset=>reset,s=>p(311)(54),cout=>p(312)(55));
FA_ff_11403:FAff port map(x=>p(272)(55),y=>p(273)(55),Cin=>p(274)(55),clock=>clock,reset=>reset,s=>p(311)(55),cout=>p(312)(56));
FA_ff_11404:FAff port map(x=>p(272)(56),y=>p(273)(56),Cin=>p(274)(56),clock=>clock,reset=>reset,s=>p(311)(56),cout=>p(312)(57));
FA_ff_11405:FAff port map(x=>p(272)(57),y=>p(273)(57),Cin=>p(274)(57),clock=>clock,reset=>reset,s=>p(311)(57),cout=>p(312)(58));
FA_ff_11406:FAff port map(x=>p(272)(58),y=>p(273)(58),Cin=>p(274)(58),clock=>clock,reset=>reset,s=>p(311)(58),cout=>p(312)(59));
FA_ff_11407:FAff port map(x=>p(272)(59),y=>p(273)(59),Cin=>p(274)(59),clock=>clock,reset=>reset,s=>p(311)(59),cout=>p(312)(60));
FA_ff_11408:FAff port map(x=>p(272)(60),y=>p(273)(60),Cin=>p(274)(60),clock=>clock,reset=>reset,s=>p(311)(60),cout=>p(312)(61));
FA_ff_11409:FAff port map(x=>p(272)(61),y=>p(273)(61),Cin=>p(274)(61),clock=>clock,reset=>reset,s=>p(311)(61),cout=>p(312)(62));
FA_ff_11410:FAff port map(x=>p(272)(62),y=>p(273)(62),Cin=>p(274)(62),clock=>clock,reset=>reset,s=>p(311)(62),cout=>p(312)(63));
FA_ff_11411:FAff port map(x=>p(272)(63),y=>p(273)(63),Cin=>p(274)(63),clock=>clock,reset=>reset,s=>p(311)(63),cout=>p(312)(64));
FA_ff_11412:FAff port map(x=>p(272)(64),y=>p(273)(64),Cin=>p(274)(64),clock=>clock,reset=>reset,s=>p(311)(64),cout=>p(312)(65));
FA_ff_11413:FAff port map(x=>p(272)(65),y=>p(273)(65),Cin=>p(274)(65),clock=>clock,reset=>reset,s=>p(311)(65),cout=>p(312)(66));
FA_ff_11414:FAff port map(x=>p(272)(66),y=>p(273)(66),Cin=>p(274)(66),clock=>clock,reset=>reset,s=>p(311)(66),cout=>p(312)(67));
FA_ff_11415:FAff port map(x=>p(272)(67),y=>p(273)(67),Cin=>p(274)(67),clock=>clock,reset=>reset,s=>p(311)(67),cout=>p(312)(68));
FA_ff_11416:FAff port map(x=>p(272)(68),y=>p(273)(68),Cin=>p(274)(68),clock=>clock,reset=>reset,s=>p(311)(68),cout=>p(312)(69));
FA_ff_11417:FAff port map(x=>p(272)(69),y=>p(273)(69),Cin=>p(274)(69),clock=>clock,reset=>reset,s=>p(311)(69),cout=>p(312)(70));
FA_ff_11418:FAff port map(x=>p(272)(70),y=>p(273)(70),Cin=>p(274)(70),clock=>clock,reset=>reset,s=>p(311)(70),cout=>p(312)(71));
FA_ff_11419:FAff port map(x=>p(272)(71),y=>p(273)(71),Cin=>p(274)(71),clock=>clock,reset=>reset,s=>p(311)(71),cout=>p(312)(72));
FA_ff_11420:FAff port map(x=>p(272)(72),y=>p(273)(72),Cin=>p(274)(72),clock=>clock,reset=>reset,s=>p(311)(72),cout=>p(312)(73));
FA_ff_11421:FAff port map(x=>p(272)(73),y=>p(273)(73),Cin=>p(274)(73),clock=>clock,reset=>reset,s=>p(311)(73),cout=>p(312)(74));
FA_ff_11422:FAff port map(x=>p(272)(74),y=>p(273)(74),Cin=>p(274)(74),clock=>clock,reset=>reset,s=>p(311)(74),cout=>p(312)(75));
FA_ff_11423:FAff port map(x=>p(272)(75),y=>p(273)(75),Cin=>p(274)(75),clock=>clock,reset=>reset,s=>p(311)(75),cout=>p(312)(76));
FA_ff_11424:FAff port map(x=>p(272)(76),y=>p(273)(76),Cin=>p(274)(76),clock=>clock,reset=>reset,s=>p(311)(76),cout=>p(312)(77));
FA_ff_11425:FAff port map(x=>p(272)(77),y=>p(273)(77),Cin=>p(274)(77),clock=>clock,reset=>reset,s=>p(311)(77),cout=>p(312)(78));
FA_ff_11426:FAff port map(x=>p(272)(78),y=>p(273)(78),Cin=>p(274)(78),clock=>clock,reset=>reset,s=>p(311)(78),cout=>p(312)(79));
FA_ff_11427:FAff port map(x=>p(272)(79),y=>p(273)(79),Cin=>p(274)(79),clock=>clock,reset=>reset,s=>p(311)(79),cout=>p(312)(80));
FA_ff_11428:FAff port map(x=>p(272)(80),y=>p(273)(80),Cin=>p(274)(80),clock=>clock,reset=>reset,s=>p(311)(80),cout=>p(312)(81));
FA_ff_11429:FAff port map(x=>p(272)(81),y=>p(273)(81),Cin=>p(274)(81),clock=>clock,reset=>reset,s=>p(311)(81),cout=>p(312)(82));
FA_ff_11430:FAff port map(x=>p(272)(82),y=>p(273)(82),Cin=>p(274)(82),clock=>clock,reset=>reset,s=>p(311)(82),cout=>p(312)(83));
FA_ff_11431:FAff port map(x=>p(272)(83),y=>p(273)(83),Cin=>p(274)(83),clock=>clock,reset=>reset,s=>p(311)(83),cout=>p(312)(84));
FA_ff_11432:FAff port map(x=>p(272)(84),y=>p(273)(84),Cin=>p(274)(84),clock=>clock,reset=>reset,s=>p(311)(84),cout=>p(312)(85));
FA_ff_11433:FAff port map(x=>p(272)(85),y=>p(273)(85),Cin=>p(274)(85),clock=>clock,reset=>reset,s=>p(311)(85),cout=>p(312)(86));
FA_ff_11434:FAff port map(x=>p(272)(86),y=>p(273)(86),Cin=>p(274)(86),clock=>clock,reset=>reset,s=>p(311)(86),cout=>p(312)(87));
FA_ff_11435:FAff port map(x=>p(272)(87),y=>p(273)(87),Cin=>p(274)(87),clock=>clock,reset=>reset,s=>p(311)(87),cout=>p(312)(88));
FA_ff_11436:FAff port map(x=>p(272)(88),y=>p(273)(88),Cin=>p(274)(88),clock=>clock,reset=>reset,s=>p(311)(88),cout=>p(312)(89));
FA_ff_11437:FAff port map(x=>p(272)(89),y=>p(273)(89),Cin=>p(274)(89),clock=>clock,reset=>reset,s=>p(311)(89),cout=>p(312)(90));
FA_ff_11438:FAff port map(x=>p(272)(90),y=>p(273)(90),Cin=>p(274)(90),clock=>clock,reset=>reset,s=>p(311)(90),cout=>p(312)(91));
FA_ff_11439:FAff port map(x=>p(272)(91),y=>p(273)(91),Cin=>p(274)(91),clock=>clock,reset=>reset,s=>p(311)(91),cout=>p(312)(92));
FA_ff_11440:FAff port map(x=>p(272)(92),y=>p(273)(92),Cin=>p(274)(92),clock=>clock,reset=>reset,s=>p(311)(92),cout=>p(312)(93));
FA_ff_11441:FAff port map(x=>p(272)(93),y=>p(273)(93),Cin=>p(274)(93),clock=>clock,reset=>reset,s=>p(311)(93),cout=>p(312)(94));
FA_ff_11442:FAff port map(x=>p(272)(94),y=>p(273)(94),Cin=>p(274)(94),clock=>clock,reset=>reset,s=>p(311)(94),cout=>p(312)(95));
FA_ff_11443:FAff port map(x=>p(272)(95),y=>p(273)(95),Cin=>p(274)(95),clock=>clock,reset=>reset,s=>p(311)(95),cout=>p(312)(96));
FA_ff_11444:FAff port map(x=>p(272)(96),y=>p(273)(96),Cin=>p(274)(96),clock=>clock,reset=>reset,s=>p(311)(96),cout=>p(312)(97));
FA_ff_11445:FAff port map(x=>p(272)(97),y=>p(273)(97),Cin=>p(274)(97),clock=>clock,reset=>reset,s=>p(311)(97),cout=>p(312)(98));
FA_ff_11446:FAff port map(x=>p(272)(98),y=>p(273)(98),Cin=>p(274)(98),clock=>clock,reset=>reset,s=>p(311)(98),cout=>p(312)(99));
FA_ff_11447:FAff port map(x=>p(272)(99),y=>p(273)(99),Cin=>p(274)(99),clock=>clock,reset=>reset,s=>p(311)(99),cout=>p(312)(100));
FA_ff_11448:FAff port map(x=>p(272)(100),y=>p(273)(100),Cin=>p(274)(100),clock=>clock,reset=>reset,s=>p(311)(100),cout=>p(312)(101));
FA_ff_11449:FAff port map(x=>p(272)(101),y=>p(273)(101),Cin=>p(274)(101),clock=>clock,reset=>reset,s=>p(311)(101),cout=>p(312)(102));
FA_ff_11450:FAff port map(x=>p(272)(102),y=>p(273)(102),Cin=>p(274)(102),clock=>clock,reset=>reset,s=>p(311)(102),cout=>p(312)(103));
FA_ff_11451:FAff port map(x=>p(272)(103),y=>p(273)(103),Cin=>p(274)(103),clock=>clock,reset=>reset,s=>p(311)(103),cout=>p(312)(104));
FA_ff_11452:FAff port map(x=>p(272)(104),y=>p(273)(104),Cin=>p(274)(104),clock=>clock,reset=>reset,s=>p(311)(104),cout=>p(312)(105));
FA_ff_11453:FAff port map(x=>p(272)(105),y=>p(273)(105),Cin=>p(274)(105),clock=>clock,reset=>reset,s=>p(311)(105),cout=>p(312)(106));
FA_ff_11454:FAff port map(x=>p(272)(106),y=>p(273)(106),Cin=>p(274)(106),clock=>clock,reset=>reset,s=>p(311)(106),cout=>p(312)(107));
FA_ff_11455:FAff port map(x=>p(272)(107),y=>p(273)(107),Cin=>p(274)(107),clock=>clock,reset=>reset,s=>p(311)(107),cout=>p(312)(108));
FA_ff_11456:FAff port map(x=>p(272)(108),y=>p(273)(108),Cin=>p(274)(108),clock=>clock,reset=>reset,s=>p(311)(108),cout=>p(312)(109));
FA_ff_11457:FAff port map(x=>p(272)(109),y=>p(273)(109),Cin=>p(274)(109),clock=>clock,reset=>reset,s=>p(311)(109),cout=>p(312)(110));
FA_ff_11458:FAff port map(x=>p(272)(110),y=>p(273)(110),Cin=>p(274)(110),clock=>clock,reset=>reset,s=>p(311)(110),cout=>p(312)(111));
FA_ff_11459:FAff port map(x=>p(272)(111),y=>p(273)(111),Cin=>p(274)(111),clock=>clock,reset=>reset,s=>p(311)(111),cout=>p(312)(112));
FA_ff_11460:FAff port map(x=>p(272)(112),y=>p(273)(112),Cin=>p(274)(112),clock=>clock,reset=>reset,s=>p(311)(112),cout=>p(312)(113));
FA_ff_11461:FAff port map(x=>p(272)(113),y=>p(273)(113),Cin=>p(274)(113),clock=>clock,reset=>reset,s=>p(311)(113),cout=>p(312)(114));
FA_ff_11462:FAff port map(x=>p(272)(114),y=>p(273)(114),Cin=>p(274)(114),clock=>clock,reset=>reset,s=>p(311)(114),cout=>p(312)(115));
FA_ff_11463:FAff port map(x=>p(272)(115),y=>p(273)(115),Cin=>p(274)(115),clock=>clock,reset=>reset,s=>p(311)(115),cout=>p(312)(116));
FA_ff_11464:FAff port map(x=>p(272)(116),y=>p(273)(116),Cin=>p(274)(116),clock=>clock,reset=>reset,s=>p(311)(116),cout=>p(312)(117));
FA_ff_11465:FAff port map(x=>p(272)(117),y=>p(273)(117),Cin=>p(274)(117),clock=>clock,reset=>reset,s=>p(311)(117),cout=>p(312)(118));
FA_ff_11466:FAff port map(x=>p(272)(118),y=>p(273)(118),Cin=>p(274)(118),clock=>clock,reset=>reset,s=>p(311)(118),cout=>p(312)(119));
FA_ff_11467:FAff port map(x=>p(272)(119),y=>p(273)(119),Cin=>p(274)(119),clock=>clock,reset=>reset,s=>p(311)(119),cout=>p(312)(120));
FA_ff_11468:FAff port map(x=>p(272)(120),y=>p(273)(120),Cin=>p(274)(120),clock=>clock,reset=>reset,s=>p(311)(120),cout=>p(312)(121));
FA_ff_11469:FAff port map(x=>p(272)(121),y=>p(273)(121),Cin=>p(274)(121),clock=>clock,reset=>reset,s=>p(311)(121),cout=>p(312)(122));
FA_ff_11470:FAff port map(x=>p(272)(122),y=>p(273)(122),Cin=>p(274)(122),clock=>clock,reset=>reset,s=>p(311)(122),cout=>p(312)(123));
FA_ff_11471:FAff port map(x=>p(272)(123),y=>p(273)(123),Cin=>p(274)(123),clock=>clock,reset=>reset,s=>p(311)(123),cout=>p(312)(124));
FA_ff_11472:FAff port map(x=>p(272)(124),y=>p(273)(124),Cin=>p(274)(124),clock=>clock,reset=>reset,s=>p(311)(124),cout=>p(312)(125));
FA_ff_11473:FAff port map(x=>p(272)(125),y=>p(273)(125),Cin=>p(274)(125),clock=>clock,reset=>reset,s=>p(311)(125),cout=>p(312)(126));
FA_ff_11474:FAff port map(x=>p(272)(126),y=>p(273)(126),Cin=>p(274)(126),clock=>clock,reset=>reset,s=>p(311)(126),cout=>p(312)(127));
FA_ff_11475:FAff port map(x=>p(272)(127),y=>p(273)(127),Cin=>p(274)(127),clock=>clock,reset=>reset,s=>p(311)(127),cout=>p(312)(128));
FA_ff_11476:FAff port map(x=>p(272)(128),y=>p(273)(128),Cin=>p(274)(128),clock=>clock,reset=>reset,s=>p(311)(128),cout=>p(312)(129));
HA_ff_54:HAff port map(x=>p(273)(129),y=>p(274)(129),clock=>clock,reset=>reset,s=>p(311)(129),c=>p(312)(130));
p(313)(0)<=p(276)(0);
HA_ff_55:HAff port map(x=>p(276)(1),y=>p(277)(1),clock=>clock,reset=>reset,s=>p(313)(1),c=>p(314)(2));
FA_ff_11477:FAff port map(x=>p(275)(2),y=>p(276)(2),Cin=>p(277)(2),clock=>clock,reset=>reset,s=>p(313)(2),cout=>p(314)(3));
FA_ff_11478:FAff port map(x=>p(275)(3),y=>p(276)(3),Cin=>p(277)(3),clock=>clock,reset=>reset,s=>p(313)(3),cout=>p(314)(4));
FA_ff_11479:FAff port map(x=>p(275)(4),y=>p(276)(4),Cin=>p(277)(4),clock=>clock,reset=>reset,s=>p(313)(4),cout=>p(314)(5));
FA_ff_11480:FAff port map(x=>p(275)(5),y=>p(276)(5),Cin=>p(277)(5),clock=>clock,reset=>reset,s=>p(313)(5),cout=>p(314)(6));
FA_ff_11481:FAff port map(x=>p(275)(6),y=>p(276)(6),Cin=>p(277)(6),clock=>clock,reset=>reset,s=>p(313)(6),cout=>p(314)(7));
FA_ff_11482:FAff port map(x=>p(275)(7),y=>p(276)(7),Cin=>p(277)(7),clock=>clock,reset=>reset,s=>p(313)(7),cout=>p(314)(8));
FA_ff_11483:FAff port map(x=>p(275)(8),y=>p(276)(8),Cin=>p(277)(8),clock=>clock,reset=>reset,s=>p(313)(8),cout=>p(314)(9));
FA_ff_11484:FAff port map(x=>p(275)(9),y=>p(276)(9),Cin=>p(277)(9),clock=>clock,reset=>reset,s=>p(313)(9),cout=>p(314)(10));
FA_ff_11485:FAff port map(x=>p(275)(10),y=>p(276)(10),Cin=>p(277)(10),clock=>clock,reset=>reset,s=>p(313)(10),cout=>p(314)(11));
FA_ff_11486:FAff port map(x=>p(275)(11),y=>p(276)(11),Cin=>p(277)(11),clock=>clock,reset=>reset,s=>p(313)(11),cout=>p(314)(12));
FA_ff_11487:FAff port map(x=>p(275)(12),y=>p(276)(12),Cin=>p(277)(12),clock=>clock,reset=>reset,s=>p(313)(12),cout=>p(314)(13));
FA_ff_11488:FAff port map(x=>p(275)(13),y=>p(276)(13),Cin=>p(277)(13),clock=>clock,reset=>reset,s=>p(313)(13),cout=>p(314)(14));
FA_ff_11489:FAff port map(x=>p(275)(14),y=>p(276)(14),Cin=>p(277)(14),clock=>clock,reset=>reset,s=>p(313)(14),cout=>p(314)(15));
FA_ff_11490:FAff port map(x=>p(275)(15),y=>p(276)(15),Cin=>p(277)(15),clock=>clock,reset=>reset,s=>p(313)(15),cout=>p(314)(16));
FA_ff_11491:FAff port map(x=>p(275)(16),y=>p(276)(16),Cin=>p(277)(16),clock=>clock,reset=>reset,s=>p(313)(16),cout=>p(314)(17));
FA_ff_11492:FAff port map(x=>p(275)(17),y=>p(276)(17),Cin=>p(277)(17),clock=>clock,reset=>reset,s=>p(313)(17),cout=>p(314)(18));
FA_ff_11493:FAff port map(x=>p(275)(18),y=>p(276)(18),Cin=>p(277)(18),clock=>clock,reset=>reset,s=>p(313)(18),cout=>p(314)(19));
FA_ff_11494:FAff port map(x=>p(275)(19),y=>p(276)(19),Cin=>p(277)(19),clock=>clock,reset=>reset,s=>p(313)(19),cout=>p(314)(20));
FA_ff_11495:FAff port map(x=>p(275)(20),y=>p(276)(20),Cin=>p(277)(20),clock=>clock,reset=>reset,s=>p(313)(20),cout=>p(314)(21));
FA_ff_11496:FAff port map(x=>p(275)(21),y=>p(276)(21),Cin=>p(277)(21),clock=>clock,reset=>reset,s=>p(313)(21),cout=>p(314)(22));
FA_ff_11497:FAff port map(x=>p(275)(22),y=>p(276)(22),Cin=>p(277)(22),clock=>clock,reset=>reset,s=>p(313)(22),cout=>p(314)(23));
FA_ff_11498:FAff port map(x=>p(275)(23),y=>p(276)(23),Cin=>p(277)(23),clock=>clock,reset=>reset,s=>p(313)(23),cout=>p(314)(24));
FA_ff_11499:FAff port map(x=>p(275)(24),y=>p(276)(24),Cin=>p(277)(24),clock=>clock,reset=>reset,s=>p(313)(24),cout=>p(314)(25));
FA_ff_11500:FAff port map(x=>p(275)(25),y=>p(276)(25),Cin=>p(277)(25),clock=>clock,reset=>reset,s=>p(313)(25),cout=>p(314)(26));
FA_ff_11501:FAff port map(x=>p(275)(26),y=>p(276)(26),Cin=>p(277)(26),clock=>clock,reset=>reset,s=>p(313)(26),cout=>p(314)(27));
FA_ff_11502:FAff port map(x=>p(275)(27),y=>p(276)(27),Cin=>p(277)(27),clock=>clock,reset=>reset,s=>p(313)(27),cout=>p(314)(28));
FA_ff_11503:FAff port map(x=>p(275)(28),y=>p(276)(28),Cin=>p(277)(28),clock=>clock,reset=>reset,s=>p(313)(28),cout=>p(314)(29));
FA_ff_11504:FAff port map(x=>p(275)(29),y=>p(276)(29),Cin=>p(277)(29),clock=>clock,reset=>reset,s=>p(313)(29),cout=>p(314)(30));
FA_ff_11505:FAff port map(x=>p(275)(30),y=>p(276)(30),Cin=>p(277)(30),clock=>clock,reset=>reset,s=>p(313)(30),cout=>p(314)(31));
FA_ff_11506:FAff port map(x=>p(275)(31),y=>p(276)(31),Cin=>p(277)(31),clock=>clock,reset=>reset,s=>p(313)(31),cout=>p(314)(32));
FA_ff_11507:FAff port map(x=>p(275)(32),y=>p(276)(32),Cin=>p(277)(32),clock=>clock,reset=>reset,s=>p(313)(32),cout=>p(314)(33));
FA_ff_11508:FAff port map(x=>p(275)(33),y=>p(276)(33),Cin=>p(277)(33),clock=>clock,reset=>reset,s=>p(313)(33),cout=>p(314)(34));
FA_ff_11509:FAff port map(x=>p(275)(34),y=>p(276)(34),Cin=>p(277)(34),clock=>clock,reset=>reset,s=>p(313)(34),cout=>p(314)(35));
FA_ff_11510:FAff port map(x=>p(275)(35),y=>p(276)(35),Cin=>p(277)(35),clock=>clock,reset=>reset,s=>p(313)(35),cout=>p(314)(36));
FA_ff_11511:FAff port map(x=>p(275)(36),y=>p(276)(36),Cin=>p(277)(36),clock=>clock,reset=>reset,s=>p(313)(36),cout=>p(314)(37));
FA_ff_11512:FAff port map(x=>p(275)(37),y=>p(276)(37),Cin=>p(277)(37),clock=>clock,reset=>reset,s=>p(313)(37),cout=>p(314)(38));
FA_ff_11513:FAff port map(x=>p(275)(38),y=>p(276)(38),Cin=>p(277)(38),clock=>clock,reset=>reset,s=>p(313)(38),cout=>p(314)(39));
FA_ff_11514:FAff port map(x=>p(275)(39),y=>p(276)(39),Cin=>p(277)(39),clock=>clock,reset=>reset,s=>p(313)(39),cout=>p(314)(40));
FA_ff_11515:FAff port map(x=>p(275)(40),y=>p(276)(40),Cin=>p(277)(40),clock=>clock,reset=>reset,s=>p(313)(40),cout=>p(314)(41));
FA_ff_11516:FAff port map(x=>p(275)(41),y=>p(276)(41),Cin=>p(277)(41),clock=>clock,reset=>reset,s=>p(313)(41),cout=>p(314)(42));
FA_ff_11517:FAff port map(x=>p(275)(42),y=>p(276)(42),Cin=>p(277)(42),clock=>clock,reset=>reset,s=>p(313)(42),cout=>p(314)(43));
FA_ff_11518:FAff port map(x=>p(275)(43),y=>p(276)(43),Cin=>p(277)(43),clock=>clock,reset=>reset,s=>p(313)(43),cout=>p(314)(44));
FA_ff_11519:FAff port map(x=>p(275)(44),y=>p(276)(44),Cin=>p(277)(44),clock=>clock,reset=>reset,s=>p(313)(44),cout=>p(314)(45));
FA_ff_11520:FAff port map(x=>p(275)(45),y=>p(276)(45),Cin=>p(277)(45),clock=>clock,reset=>reset,s=>p(313)(45),cout=>p(314)(46));
FA_ff_11521:FAff port map(x=>p(275)(46),y=>p(276)(46),Cin=>p(277)(46),clock=>clock,reset=>reset,s=>p(313)(46),cout=>p(314)(47));
FA_ff_11522:FAff port map(x=>p(275)(47),y=>p(276)(47),Cin=>p(277)(47),clock=>clock,reset=>reset,s=>p(313)(47),cout=>p(314)(48));
FA_ff_11523:FAff port map(x=>p(275)(48),y=>p(276)(48),Cin=>p(277)(48),clock=>clock,reset=>reset,s=>p(313)(48),cout=>p(314)(49));
FA_ff_11524:FAff port map(x=>p(275)(49),y=>p(276)(49),Cin=>p(277)(49),clock=>clock,reset=>reset,s=>p(313)(49),cout=>p(314)(50));
FA_ff_11525:FAff port map(x=>p(275)(50),y=>p(276)(50),Cin=>p(277)(50),clock=>clock,reset=>reset,s=>p(313)(50),cout=>p(314)(51));
FA_ff_11526:FAff port map(x=>p(275)(51),y=>p(276)(51),Cin=>p(277)(51),clock=>clock,reset=>reset,s=>p(313)(51),cout=>p(314)(52));
FA_ff_11527:FAff port map(x=>p(275)(52),y=>p(276)(52),Cin=>p(277)(52),clock=>clock,reset=>reset,s=>p(313)(52),cout=>p(314)(53));
FA_ff_11528:FAff port map(x=>p(275)(53),y=>p(276)(53),Cin=>p(277)(53),clock=>clock,reset=>reset,s=>p(313)(53),cout=>p(314)(54));
FA_ff_11529:FAff port map(x=>p(275)(54),y=>p(276)(54),Cin=>p(277)(54),clock=>clock,reset=>reset,s=>p(313)(54),cout=>p(314)(55));
FA_ff_11530:FAff port map(x=>p(275)(55),y=>p(276)(55),Cin=>p(277)(55),clock=>clock,reset=>reset,s=>p(313)(55),cout=>p(314)(56));
FA_ff_11531:FAff port map(x=>p(275)(56),y=>p(276)(56),Cin=>p(277)(56),clock=>clock,reset=>reset,s=>p(313)(56),cout=>p(314)(57));
FA_ff_11532:FAff port map(x=>p(275)(57),y=>p(276)(57),Cin=>p(277)(57),clock=>clock,reset=>reset,s=>p(313)(57),cout=>p(314)(58));
FA_ff_11533:FAff port map(x=>p(275)(58),y=>p(276)(58),Cin=>p(277)(58),clock=>clock,reset=>reset,s=>p(313)(58),cout=>p(314)(59));
FA_ff_11534:FAff port map(x=>p(275)(59),y=>p(276)(59),Cin=>p(277)(59),clock=>clock,reset=>reset,s=>p(313)(59),cout=>p(314)(60));
FA_ff_11535:FAff port map(x=>p(275)(60),y=>p(276)(60),Cin=>p(277)(60),clock=>clock,reset=>reset,s=>p(313)(60),cout=>p(314)(61));
FA_ff_11536:FAff port map(x=>p(275)(61),y=>p(276)(61),Cin=>p(277)(61),clock=>clock,reset=>reset,s=>p(313)(61),cout=>p(314)(62));
FA_ff_11537:FAff port map(x=>p(275)(62),y=>p(276)(62),Cin=>p(277)(62),clock=>clock,reset=>reset,s=>p(313)(62),cout=>p(314)(63));
FA_ff_11538:FAff port map(x=>p(275)(63),y=>p(276)(63),Cin=>p(277)(63),clock=>clock,reset=>reset,s=>p(313)(63),cout=>p(314)(64));
FA_ff_11539:FAff port map(x=>p(275)(64),y=>p(276)(64),Cin=>p(277)(64),clock=>clock,reset=>reset,s=>p(313)(64),cout=>p(314)(65));
FA_ff_11540:FAff port map(x=>p(275)(65),y=>p(276)(65),Cin=>p(277)(65),clock=>clock,reset=>reset,s=>p(313)(65),cout=>p(314)(66));
FA_ff_11541:FAff port map(x=>p(275)(66),y=>p(276)(66),Cin=>p(277)(66),clock=>clock,reset=>reset,s=>p(313)(66),cout=>p(314)(67));
FA_ff_11542:FAff port map(x=>p(275)(67),y=>p(276)(67),Cin=>p(277)(67),clock=>clock,reset=>reset,s=>p(313)(67),cout=>p(314)(68));
FA_ff_11543:FAff port map(x=>p(275)(68),y=>p(276)(68),Cin=>p(277)(68),clock=>clock,reset=>reset,s=>p(313)(68),cout=>p(314)(69));
FA_ff_11544:FAff port map(x=>p(275)(69),y=>p(276)(69),Cin=>p(277)(69),clock=>clock,reset=>reset,s=>p(313)(69),cout=>p(314)(70));
FA_ff_11545:FAff port map(x=>p(275)(70),y=>p(276)(70),Cin=>p(277)(70),clock=>clock,reset=>reset,s=>p(313)(70),cout=>p(314)(71));
FA_ff_11546:FAff port map(x=>p(275)(71),y=>p(276)(71),Cin=>p(277)(71),clock=>clock,reset=>reset,s=>p(313)(71),cout=>p(314)(72));
FA_ff_11547:FAff port map(x=>p(275)(72),y=>p(276)(72),Cin=>p(277)(72),clock=>clock,reset=>reset,s=>p(313)(72),cout=>p(314)(73));
FA_ff_11548:FAff port map(x=>p(275)(73),y=>p(276)(73),Cin=>p(277)(73),clock=>clock,reset=>reset,s=>p(313)(73),cout=>p(314)(74));
FA_ff_11549:FAff port map(x=>p(275)(74),y=>p(276)(74),Cin=>p(277)(74),clock=>clock,reset=>reset,s=>p(313)(74),cout=>p(314)(75));
FA_ff_11550:FAff port map(x=>p(275)(75),y=>p(276)(75),Cin=>p(277)(75),clock=>clock,reset=>reset,s=>p(313)(75),cout=>p(314)(76));
FA_ff_11551:FAff port map(x=>p(275)(76),y=>p(276)(76),Cin=>p(277)(76),clock=>clock,reset=>reset,s=>p(313)(76),cout=>p(314)(77));
FA_ff_11552:FAff port map(x=>p(275)(77),y=>p(276)(77),Cin=>p(277)(77),clock=>clock,reset=>reset,s=>p(313)(77),cout=>p(314)(78));
FA_ff_11553:FAff port map(x=>p(275)(78),y=>p(276)(78),Cin=>p(277)(78),clock=>clock,reset=>reset,s=>p(313)(78),cout=>p(314)(79));
FA_ff_11554:FAff port map(x=>p(275)(79),y=>p(276)(79),Cin=>p(277)(79),clock=>clock,reset=>reset,s=>p(313)(79),cout=>p(314)(80));
FA_ff_11555:FAff port map(x=>p(275)(80),y=>p(276)(80),Cin=>p(277)(80),clock=>clock,reset=>reset,s=>p(313)(80),cout=>p(314)(81));
FA_ff_11556:FAff port map(x=>p(275)(81),y=>p(276)(81),Cin=>p(277)(81),clock=>clock,reset=>reset,s=>p(313)(81),cout=>p(314)(82));
FA_ff_11557:FAff port map(x=>p(275)(82),y=>p(276)(82),Cin=>p(277)(82),clock=>clock,reset=>reset,s=>p(313)(82),cout=>p(314)(83));
FA_ff_11558:FAff port map(x=>p(275)(83),y=>p(276)(83),Cin=>p(277)(83),clock=>clock,reset=>reset,s=>p(313)(83),cout=>p(314)(84));
FA_ff_11559:FAff port map(x=>p(275)(84),y=>p(276)(84),Cin=>p(277)(84),clock=>clock,reset=>reset,s=>p(313)(84),cout=>p(314)(85));
FA_ff_11560:FAff port map(x=>p(275)(85),y=>p(276)(85),Cin=>p(277)(85),clock=>clock,reset=>reset,s=>p(313)(85),cout=>p(314)(86));
FA_ff_11561:FAff port map(x=>p(275)(86),y=>p(276)(86),Cin=>p(277)(86),clock=>clock,reset=>reset,s=>p(313)(86),cout=>p(314)(87));
FA_ff_11562:FAff port map(x=>p(275)(87),y=>p(276)(87),Cin=>p(277)(87),clock=>clock,reset=>reset,s=>p(313)(87),cout=>p(314)(88));
FA_ff_11563:FAff port map(x=>p(275)(88),y=>p(276)(88),Cin=>p(277)(88),clock=>clock,reset=>reset,s=>p(313)(88),cout=>p(314)(89));
FA_ff_11564:FAff port map(x=>p(275)(89),y=>p(276)(89),Cin=>p(277)(89),clock=>clock,reset=>reset,s=>p(313)(89),cout=>p(314)(90));
FA_ff_11565:FAff port map(x=>p(275)(90),y=>p(276)(90),Cin=>p(277)(90),clock=>clock,reset=>reset,s=>p(313)(90),cout=>p(314)(91));
FA_ff_11566:FAff port map(x=>p(275)(91),y=>p(276)(91),Cin=>p(277)(91),clock=>clock,reset=>reset,s=>p(313)(91),cout=>p(314)(92));
FA_ff_11567:FAff port map(x=>p(275)(92),y=>p(276)(92),Cin=>p(277)(92),clock=>clock,reset=>reset,s=>p(313)(92),cout=>p(314)(93));
FA_ff_11568:FAff port map(x=>p(275)(93),y=>p(276)(93),Cin=>p(277)(93),clock=>clock,reset=>reset,s=>p(313)(93),cout=>p(314)(94));
FA_ff_11569:FAff port map(x=>p(275)(94),y=>p(276)(94),Cin=>p(277)(94),clock=>clock,reset=>reset,s=>p(313)(94),cout=>p(314)(95));
FA_ff_11570:FAff port map(x=>p(275)(95),y=>p(276)(95),Cin=>p(277)(95),clock=>clock,reset=>reset,s=>p(313)(95),cout=>p(314)(96));
FA_ff_11571:FAff port map(x=>p(275)(96),y=>p(276)(96),Cin=>p(277)(96),clock=>clock,reset=>reset,s=>p(313)(96),cout=>p(314)(97));
FA_ff_11572:FAff port map(x=>p(275)(97),y=>p(276)(97),Cin=>p(277)(97),clock=>clock,reset=>reset,s=>p(313)(97),cout=>p(314)(98));
FA_ff_11573:FAff port map(x=>p(275)(98),y=>p(276)(98),Cin=>p(277)(98),clock=>clock,reset=>reset,s=>p(313)(98),cout=>p(314)(99));
FA_ff_11574:FAff port map(x=>p(275)(99),y=>p(276)(99),Cin=>p(277)(99),clock=>clock,reset=>reset,s=>p(313)(99),cout=>p(314)(100));
FA_ff_11575:FAff port map(x=>p(275)(100),y=>p(276)(100),Cin=>p(277)(100),clock=>clock,reset=>reset,s=>p(313)(100),cout=>p(314)(101));
FA_ff_11576:FAff port map(x=>p(275)(101),y=>p(276)(101),Cin=>p(277)(101),clock=>clock,reset=>reset,s=>p(313)(101),cout=>p(314)(102));
FA_ff_11577:FAff port map(x=>p(275)(102),y=>p(276)(102),Cin=>p(277)(102),clock=>clock,reset=>reset,s=>p(313)(102),cout=>p(314)(103));
FA_ff_11578:FAff port map(x=>p(275)(103),y=>p(276)(103),Cin=>p(277)(103),clock=>clock,reset=>reset,s=>p(313)(103),cout=>p(314)(104));
FA_ff_11579:FAff port map(x=>p(275)(104),y=>p(276)(104),Cin=>p(277)(104),clock=>clock,reset=>reset,s=>p(313)(104),cout=>p(314)(105));
FA_ff_11580:FAff port map(x=>p(275)(105),y=>p(276)(105),Cin=>p(277)(105),clock=>clock,reset=>reset,s=>p(313)(105),cout=>p(314)(106));
FA_ff_11581:FAff port map(x=>p(275)(106),y=>p(276)(106),Cin=>p(277)(106),clock=>clock,reset=>reset,s=>p(313)(106),cout=>p(314)(107));
FA_ff_11582:FAff port map(x=>p(275)(107),y=>p(276)(107),Cin=>p(277)(107),clock=>clock,reset=>reset,s=>p(313)(107),cout=>p(314)(108));
FA_ff_11583:FAff port map(x=>p(275)(108),y=>p(276)(108),Cin=>p(277)(108),clock=>clock,reset=>reset,s=>p(313)(108),cout=>p(314)(109));
FA_ff_11584:FAff port map(x=>p(275)(109),y=>p(276)(109),Cin=>p(277)(109),clock=>clock,reset=>reset,s=>p(313)(109),cout=>p(314)(110));
FA_ff_11585:FAff port map(x=>p(275)(110),y=>p(276)(110),Cin=>p(277)(110),clock=>clock,reset=>reset,s=>p(313)(110),cout=>p(314)(111));
FA_ff_11586:FAff port map(x=>p(275)(111),y=>p(276)(111),Cin=>p(277)(111),clock=>clock,reset=>reset,s=>p(313)(111),cout=>p(314)(112));
FA_ff_11587:FAff port map(x=>p(275)(112),y=>p(276)(112),Cin=>p(277)(112),clock=>clock,reset=>reset,s=>p(313)(112),cout=>p(314)(113));
FA_ff_11588:FAff port map(x=>p(275)(113),y=>p(276)(113),Cin=>p(277)(113),clock=>clock,reset=>reset,s=>p(313)(113),cout=>p(314)(114));
FA_ff_11589:FAff port map(x=>p(275)(114),y=>p(276)(114),Cin=>p(277)(114),clock=>clock,reset=>reset,s=>p(313)(114),cout=>p(314)(115));
FA_ff_11590:FAff port map(x=>p(275)(115),y=>p(276)(115),Cin=>p(277)(115),clock=>clock,reset=>reset,s=>p(313)(115),cout=>p(314)(116));
FA_ff_11591:FAff port map(x=>p(275)(116),y=>p(276)(116),Cin=>p(277)(116),clock=>clock,reset=>reset,s=>p(313)(116),cout=>p(314)(117));
FA_ff_11592:FAff port map(x=>p(275)(117),y=>p(276)(117),Cin=>p(277)(117),clock=>clock,reset=>reset,s=>p(313)(117),cout=>p(314)(118));
FA_ff_11593:FAff port map(x=>p(275)(118),y=>p(276)(118),Cin=>p(277)(118),clock=>clock,reset=>reset,s=>p(313)(118),cout=>p(314)(119));
FA_ff_11594:FAff port map(x=>p(275)(119),y=>p(276)(119),Cin=>p(277)(119),clock=>clock,reset=>reset,s=>p(313)(119),cout=>p(314)(120));
FA_ff_11595:FAff port map(x=>p(275)(120),y=>p(276)(120),Cin=>p(277)(120),clock=>clock,reset=>reset,s=>p(313)(120),cout=>p(314)(121));
FA_ff_11596:FAff port map(x=>p(275)(121),y=>p(276)(121),Cin=>p(277)(121),clock=>clock,reset=>reset,s=>p(313)(121),cout=>p(314)(122));
FA_ff_11597:FAff port map(x=>p(275)(122),y=>p(276)(122),Cin=>p(277)(122),clock=>clock,reset=>reset,s=>p(313)(122),cout=>p(314)(123));
FA_ff_11598:FAff port map(x=>p(275)(123),y=>p(276)(123),Cin=>p(277)(123),clock=>clock,reset=>reset,s=>p(313)(123),cout=>p(314)(124));
FA_ff_11599:FAff port map(x=>p(275)(124),y=>p(276)(124),Cin=>p(277)(124),clock=>clock,reset=>reset,s=>p(313)(124),cout=>p(314)(125));
FA_ff_11600:FAff port map(x=>p(275)(125),y=>p(276)(125),Cin=>p(277)(125),clock=>clock,reset=>reset,s=>p(313)(125),cout=>p(314)(126));
FA_ff_11601:FAff port map(x=>p(275)(126),y=>p(276)(126),Cin=>p(277)(126),clock=>clock,reset=>reset,s=>p(313)(126),cout=>p(314)(127));
FA_ff_11602:FAff port map(x=>p(275)(127),y=>p(276)(127),Cin=>p(277)(127),clock=>clock,reset=>reset,s=>p(313)(127),cout=>p(314)(128));
FA_ff_11603:FAff port map(x=>p(275)(128),y=>p(276)(128),Cin=>p(277)(128),clock=>clock,reset=>reset,s=>p(313)(128),cout=>p(314)(129));
FA_ff_11604:FAff port map(x=>p(275)(129),y=>p(276)(129),Cin=>p(277)(129),clock=>clock,reset=>reset,s=>p(313)(129),cout=>p(314)(130));
HA_ff_56:HAff port map(x=>p(278)(0),y=>p(280)(0),clock=>clock,reset=>reset,s=>p(315)(0),c=>p(316)(1));
HA_ff_57:HAff port map(x=>p(278)(1),y=>p(280)(1),clock=>clock,reset=>reset,s=>p(315)(1),c=>p(316)(2));
FA_ff_11605:FAff port map(x=>p(278)(2),y=>p(279)(2),Cin=>p(280)(2),clock=>clock,reset=>reset,s=>p(315)(2),cout=>p(316)(3));
FA_ff_11606:FAff port map(x=>p(278)(3),y=>p(279)(3),Cin=>p(280)(3),clock=>clock,reset=>reset,s=>p(315)(3),cout=>p(316)(4));
FA_ff_11607:FAff port map(x=>p(278)(4),y=>p(279)(4),Cin=>p(280)(4),clock=>clock,reset=>reset,s=>p(315)(4),cout=>p(316)(5));
FA_ff_11608:FAff port map(x=>p(278)(5),y=>p(279)(5),Cin=>p(280)(5),clock=>clock,reset=>reset,s=>p(315)(5),cout=>p(316)(6));
FA_ff_11609:FAff port map(x=>p(278)(6),y=>p(279)(6),Cin=>p(280)(6),clock=>clock,reset=>reset,s=>p(315)(6),cout=>p(316)(7));
FA_ff_11610:FAff port map(x=>p(278)(7),y=>p(279)(7),Cin=>p(280)(7),clock=>clock,reset=>reset,s=>p(315)(7),cout=>p(316)(8));
FA_ff_11611:FAff port map(x=>p(278)(8),y=>p(279)(8),Cin=>p(280)(8),clock=>clock,reset=>reset,s=>p(315)(8),cout=>p(316)(9));
FA_ff_11612:FAff port map(x=>p(278)(9),y=>p(279)(9),Cin=>p(280)(9),clock=>clock,reset=>reset,s=>p(315)(9),cout=>p(316)(10));
FA_ff_11613:FAff port map(x=>p(278)(10),y=>p(279)(10),Cin=>p(280)(10),clock=>clock,reset=>reset,s=>p(315)(10),cout=>p(316)(11));
FA_ff_11614:FAff port map(x=>p(278)(11),y=>p(279)(11),Cin=>p(280)(11),clock=>clock,reset=>reset,s=>p(315)(11),cout=>p(316)(12));
FA_ff_11615:FAff port map(x=>p(278)(12),y=>p(279)(12),Cin=>p(280)(12),clock=>clock,reset=>reset,s=>p(315)(12),cout=>p(316)(13));
FA_ff_11616:FAff port map(x=>p(278)(13),y=>p(279)(13),Cin=>p(280)(13),clock=>clock,reset=>reset,s=>p(315)(13),cout=>p(316)(14));
FA_ff_11617:FAff port map(x=>p(278)(14),y=>p(279)(14),Cin=>p(280)(14),clock=>clock,reset=>reset,s=>p(315)(14),cout=>p(316)(15));
FA_ff_11618:FAff port map(x=>p(278)(15),y=>p(279)(15),Cin=>p(280)(15),clock=>clock,reset=>reset,s=>p(315)(15),cout=>p(316)(16));
FA_ff_11619:FAff port map(x=>p(278)(16),y=>p(279)(16),Cin=>p(280)(16),clock=>clock,reset=>reset,s=>p(315)(16),cout=>p(316)(17));
FA_ff_11620:FAff port map(x=>p(278)(17),y=>p(279)(17),Cin=>p(280)(17),clock=>clock,reset=>reset,s=>p(315)(17),cout=>p(316)(18));
FA_ff_11621:FAff port map(x=>p(278)(18),y=>p(279)(18),Cin=>p(280)(18),clock=>clock,reset=>reset,s=>p(315)(18),cout=>p(316)(19));
FA_ff_11622:FAff port map(x=>p(278)(19),y=>p(279)(19),Cin=>p(280)(19),clock=>clock,reset=>reset,s=>p(315)(19),cout=>p(316)(20));
FA_ff_11623:FAff port map(x=>p(278)(20),y=>p(279)(20),Cin=>p(280)(20),clock=>clock,reset=>reset,s=>p(315)(20),cout=>p(316)(21));
FA_ff_11624:FAff port map(x=>p(278)(21),y=>p(279)(21),Cin=>p(280)(21),clock=>clock,reset=>reset,s=>p(315)(21),cout=>p(316)(22));
FA_ff_11625:FAff port map(x=>p(278)(22),y=>p(279)(22),Cin=>p(280)(22),clock=>clock,reset=>reset,s=>p(315)(22),cout=>p(316)(23));
FA_ff_11626:FAff port map(x=>p(278)(23),y=>p(279)(23),Cin=>p(280)(23),clock=>clock,reset=>reset,s=>p(315)(23),cout=>p(316)(24));
FA_ff_11627:FAff port map(x=>p(278)(24),y=>p(279)(24),Cin=>p(280)(24),clock=>clock,reset=>reset,s=>p(315)(24),cout=>p(316)(25));
FA_ff_11628:FAff port map(x=>p(278)(25),y=>p(279)(25),Cin=>p(280)(25),clock=>clock,reset=>reset,s=>p(315)(25),cout=>p(316)(26));
FA_ff_11629:FAff port map(x=>p(278)(26),y=>p(279)(26),Cin=>p(280)(26),clock=>clock,reset=>reset,s=>p(315)(26),cout=>p(316)(27));
FA_ff_11630:FAff port map(x=>p(278)(27),y=>p(279)(27),Cin=>p(280)(27),clock=>clock,reset=>reset,s=>p(315)(27),cout=>p(316)(28));
FA_ff_11631:FAff port map(x=>p(278)(28),y=>p(279)(28),Cin=>p(280)(28),clock=>clock,reset=>reset,s=>p(315)(28),cout=>p(316)(29));
FA_ff_11632:FAff port map(x=>p(278)(29),y=>p(279)(29),Cin=>p(280)(29),clock=>clock,reset=>reset,s=>p(315)(29),cout=>p(316)(30));
FA_ff_11633:FAff port map(x=>p(278)(30),y=>p(279)(30),Cin=>p(280)(30),clock=>clock,reset=>reset,s=>p(315)(30),cout=>p(316)(31));
FA_ff_11634:FAff port map(x=>p(278)(31),y=>p(279)(31),Cin=>p(280)(31),clock=>clock,reset=>reset,s=>p(315)(31),cout=>p(316)(32));
FA_ff_11635:FAff port map(x=>p(278)(32),y=>p(279)(32),Cin=>p(280)(32),clock=>clock,reset=>reset,s=>p(315)(32),cout=>p(316)(33));
FA_ff_11636:FAff port map(x=>p(278)(33),y=>p(279)(33),Cin=>p(280)(33),clock=>clock,reset=>reset,s=>p(315)(33),cout=>p(316)(34));
FA_ff_11637:FAff port map(x=>p(278)(34),y=>p(279)(34),Cin=>p(280)(34),clock=>clock,reset=>reset,s=>p(315)(34),cout=>p(316)(35));
FA_ff_11638:FAff port map(x=>p(278)(35),y=>p(279)(35),Cin=>p(280)(35),clock=>clock,reset=>reset,s=>p(315)(35),cout=>p(316)(36));
FA_ff_11639:FAff port map(x=>p(278)(36),y=>p(279)(36),Cin=>p(280)(36),clock=>clock,reset=>reset,s=>p(315)(36),cout=>p(316)(37));
FA_ff_11640:FAff port map(x=>p(278)(37),y=>p(279)(37),Cin=>p(280)(37),clock=>clock,reset=>reset,s=>p(315)(37),cout=>p(316)(38));
FA_ff_11641:FAff port map(x=>p(278)(38),y=>p(279)(38),Cin=>p(280)(38),clock=>clock,reset=>reset,s=>p(315)(38),cout=>p(316)(39));
FA_ff_11642:FAff port map(x=>p(278)(39),y=>p(279)(39),Cin=>p(280)(39),clock=>clock,reset=>reset,s=>p(315)(39),cout=>p(316)(40));
FA_ff_11643:FAff port map(x=>p(278)(40),y=>p(279)(40),Cin=>p(280)(40),clock=>clock,reset=>reset,s=>p(315)(40),cout=>p(316)(41));
FA_ff_11644:FAff port map(x=>p(278)(41),y=>p(279)(41),Cin=>p(280)(41),clock=>clock,reset=>reset,s=>p(315)(41),cout=>p(316)(42));
FA_ff_11645:FAff port map(x=>p(278)(42),y=>p(279)(42),Cin=>p(280)(42),clock=>clock,reset=>reset,s=>p(315)(42),cout=>p(316)(43));
FA_ff_11646:FAff port map(x=>p(278)(43),y=>p(279)(43),Cin=>p(280)(43),clock=>clock,reset=>reset,s=>p(315)(43),cout=>p(316)(44));
FA_ff_11647:FAff port map(x=>p(278)(44),y=>p(279)(44),Cin=>p(280)(44),clock=>clock,reset=>reset,s=>p(315)(44),cout=>p(316)(45));
FA_ff_11648:FAff port map(x=>p(278)(45),y=>p(279)(45),Cin=>p(280)(45),clock=>clock,reset=>reset,s=>p(315)(45),cout=>p(316)(46));
FA_ff_11649:FAff port map(x=>p(278)(46),y=>p(279)(46),Cin=>p(280)(46),clock=>clock,reset=>reset,s=>p(315)(46),cout=>p(316)(47));
FA_ff_11650:FAff port map(x=>p(278)(47),y=>p(279)(47),Cin=>p(280)(47),clock=>clock,reset=>reset,s=>p(315)(47),cout=>p(316)(48));
FA_ff_11651:FAff port map(x=>p(278)(48),y=>p(279)(48),Cin=>p(280)(48),clock=>clock,reset=>reset,s=>p(315)(48),cout=>p(316)(49));
FA_ff_11652:FAff port map(x=>p(278)(49),y=>p(279)(49),Cin=>p(280)(49),clock=>clock,reset=>reset,s=>p(315)(49),cout=>p(316)(50));
FA_ff_11653:FAff port map(x=>p(278)(50),y=>p(279)(50),Cin=>p(280)(50),clock=>clock,reset=>reset,s=>p(315)(50),cout=>p(316)(51));
FA_ff_11654:FAff port map(x=>p(278)(51),y=>p(279)(51),Cin=>p(280)(51),clock=>clock,reset=>reset,s=>p(315)(51),cout=>p(316)(52));
FA_ff_11655:FAff port map(x=>p(278)(52),y=>p(279)(52),Cin=>p(280)(52),clock=>clock,reset=>reset,s=>p(315)(52),cout=>p(316)(53));
FA_ff_11656:FAff port map(x=>p(278)(53),y=>p(279)(53),Cin=>p(280)(53),clock=>clock,reset=>reset,s=>p(315)(53),cout=>p(316)(54));
FA_ff_11657:FAff port map(x=>p(278)(54),y=>p(279)(54),Cin=>p(280)(54),clock=>clock,reset=>reset,s=>p(315)(54),cout=>p(316)(55));
FA_ff_11658:FAff port map(x=>p(278)(55),y=>p(279)(55),Cin=>p(280)(55),clock=>clock,reset=>reset,s=>p(315)(55),cout=>p(316)(56));
FA_ff_11659:FAff port map(x=>p(278)(56),y=>p(279)(56),Cin=>p(280)(56),clock=>clock,reset=>reset,s=>p(315)(56),cout=>p(316)(57));
FA_ff_11660:FAff port map(x=>p(278)(57),y=>p(279)(57),Cin=>p(280)(57),clock=>clock,reset=>reset,s=>p(315)(57),cout=>p(316)(58));
FA_ff_11661:FAff port map(x=>p(278)(58),y=>p(279)(58),Cin=>p(280)(58),clock=>clock,reset=>reset,s=>p(315)(58),cout=>p(316)(59));
FA_ff_11662:FAff port map(x=>p(278)(59),y=>p(279)(59),Cin=>p(280)(59),clock=>clock,reset=>reset,s=>p(315)(59),cout=>p(316)(60));
FA_ff_11663:FAff port map(x=>p(278)(60),y=>p(279)(60),Cin=>p(280)(60),clock=>clock,reset=>reset,s=>p(315)(60),cout=>p(316)(61));
FA_ff_11664:FAff port map(x=>p(278)(61),y=>p(279)(61),Cin=>p(280)(61),clock=>clock,reset=>reset,s=>p(315)(61),cout=>p(316)(62));
FA_ff_11665:FAff port map(x=>p(278)(62),y=>p(279)(62),Cin=>p(280)(62),clock=>clock,reset=>reset,s=>p(315)(62),cout=>p(316)(63));
FA_ff_11666:FAff port map(x=>p(278)(63),y=>p(279)(63),Cin=>p(280)(63),clock=>clock,reset=>reset,s=>p(315)(63),cout=>p(316)(64));
FA_ff_11667:FAff port map(x=>p(278)(64),y=>p(279)(64),Cin=>p(280)(64),clock=>clock,reset=>reset,s=>p(315)(64),cout=>p(316)(65));
FA_ff_11668:FAff port map(x=>p(278)(65),y=>p(279)(65),Cin=>p(280)(65),clock=>clock,reset=>reset,s=>p(315)(65),cout=>p(316)(66));
FA_ff_11669:FAff port map(x=>p(278)(66),y=>p(279)(66),Cin=>p(280)(66),clock=>clock,reset=>reset,s=>p(315)(66),cout=>p(316)(67));
FA_ff_11670:FAff port map(x=>p(278)(67),y=>p(279)(67),Cin=>p(280)(67),clock=>clock,reset=>reset,s=>p(315)(67),cout=>p(316)(68));
FA_ff_11671:FAff port map(x=>p(278)(68),y=>p(279)(68),Cin=>p(280)(68),clock=>clock,reset=>reset,s=>p(315)(68),cout=>p(316)(69));
FA_ff_11672:FAff port map(x=>p(278)(69),y=>p(279)(69),Cin=>p(280)(69),clock=>clock,reset=>reset,s=>p(315)(69),cout=>p(316)(70));
FA_ff_11673:FAff port map(x=>p(278)(70),y=>p(279)(70),Cin=>p(280)(70),clock=>clock,reset=>reset,s=>p(315)(70),cout=>p(316)(71));
FA_ff_11674:FAff port map(x=>p(278)(71),y=>p(279)(71),Cin=>p(280)(71),clock=>clock,reset=>reset,s=>p(315)(71),cout=>p(316)(72));
FA_ff_11675:FAff port map(x=>p(278)(72),y=>p(279)(72),Cin=>p(280)(72),clock=>clock,reset=>reset,s=>p(315)(72),cout=>p(316)(73));
FA_ff_11676:FAff port map(x=>p(278)(73),y=>p(279)(73),Cin=>p(280)(73),clock=>clock,reset=>reset,s=>p(315)(73),cout=>p(316)(74));
FA_ff_11677:FAff port map(x=>p(278)(74),y=>p(279)(74),Cin=>p(280)(74),clock=>clock,reset=>reset,s=>p(315)(74),cout=>p(316)(75));
FA_ff_11678:FAff port map(x=>p(278)(75),y=>p(279)(75),Cin=>p(280)(75),clock=>clock,reset=>reset,s=>p(315)(75),cout=>p(316)(76));
FA_ff_11679:FAff port map(x=>p(278)(76),y=>p(279)(76),Cin=>p(280)(76),clock=>clock,reset=>reset,s=>p(315)(76),cout=>p(316)(77));
FA_ff_11680:FAff port map(x=>p(278)(77),y=>p(279)(77),Cin=>p(280)(77),clock=>clock,reset=>reset,s=>p(315)(77),cout=>p(316)(78));
FA_ff_11681:FAff port map(x=>p(278)(78),y=>p(279)(78),Cin=>p(280)(78),clock=>clock,reset=>reset,s=>p(315)(78),cout=>p(316)(79));
FA_ff_11682:FAff port map(x=>p(278)(79),y=>p(279)(79),Cin=>p(280)(79),clock=>clock,reset=>reset,s=>p(315)(79),cout=>p(316)(80));
FA_ff_11683:FAff port map(x=>p(278)(80),y=>p(279)(80),Cin=>p(280)(80),clock=>clock,reset=>reset,s=>p(315)(80),cout=>p(316)(81));
FA_ff_11684:FAff port map(x=>p(278)(81),y=>p(279)(81),Cin=>p(280)(81),clock=>clock,reset=>reset,s=>p(315)(81),cout=>p(316)(82));
FA_ff_11685:FAff port map(x=>p(278)(82),y=>p(279)(82),Cin=>p(280)(82),clock=>clock,reset=>reset,s=>p(315)(82),cout=>p(316)(83));
FA_ff_11686:FAff port map(x=>p(278)(83),y=>p(279)(83),Cin=>p(280)(83),clock=>clock,reset=>reset,s=>p(315)(83),cout=>p(316)(84));
FA_ff_11687:FAff port map(x=>p(278)(84),y=>p(279)(84),Cin=>p(280)(84),clock=>clock,reset=>reset,s=>p(315)(84),cout=>p(316)(85));
FA_ff_11688:FAff port map(x=>p(278)(85),y=>p(279)(85),Cin=>p(280)(85),clock=>clock,reset=>reset,s=>p(315)(85),cout=>p(316)(86));
FA_ff_11689:FAff port map(x=>p(278)(86),y=>p(279)(86),Cin=>p(280)(86),clock=>clock,reset=>reset,s=>p(315)(86),cout=>p(316)(87));
FA_ff_11690:FAff port map(x=>p(278)(87),y=>p(279)(87),Cin=>p(280)(87),clock=>clock,reset=>reset,s=>p(315)(87),cout=>p(316)(88));
FA_ff_11691:FAff port map(x=>p(278)(88),y=>p(279)(88),Cin=>p(280)(88),clock=>clock,reset=>reset,s=>p(315)(88),cout=>p(316)(89));
FA_ff_11692:FAff port map(x=>p(278)(89),y=>p(279)(89),Cin=>p(280)(89),clock=>clock,reset=>reset,s=>p(315)(89),cout=>p(316)(90));
FA_ff_11693:FAff port map(x=>p(278)(90),y=>p(279)(90),Cin=>p(280)(90),clock=>clock,reset=>reset,s=>p(315)(90),cout=>p(316)(91));
FA_ff_11694:FAff port map(x=>p(278)(91),y=>p(279)(91),Cin=>p(280)(91),clock=>clock,reset=>reset,s=>p(315)(91),cout=>p(316)(92));
FA_ff_11695:FAff port map(x=>p(278)(92),y=>p(279)(92),Cin=>p(280)(92),clock=>clock,reset=>reset,s=>p(315)(92),cout=>p(316)(93));
FA_ff_11696:FAff port map(x=>p(278)(93),y=>p(279)(93),Cin=>p(280)(93),clock=>clock,reset=>reset,s=>p(315)(93),cout=>p(316)(94));
FA_ff_11697:FAff port map(x=>p(278)(94),y=>p(279)(94),Cin=>p(280)(94),clock=>clock,reset=>reset,s=>p(315)(94),cout=>p(316)(95));
FA_ff_11698:FAff port map(x=>p(278)(95),y=>p(279)(95),Cin=>p(280)(95),clock=>clock,reset=>reset,s=>p(315)(95),cout=>p(316)(96));
FA_ff_11699:FAff port map(x=>p(278)(96),y=>p(279)(96),Cin=>p(280)(96),clock=>clock,reset=>reset,s=>p(315)(96),cout=>p(316)(97));
FA_ff_11700:FAff port map(x=>p(278)(97),y=>p(279)(97),Cin=>p(280)(97),clock=>clock,reset=>reset,s=>p(315)(97),cout=>p(316)(98));
FA_ff_11701:FAff port map(x=>p(278)(98),y=>p(279)(98),Cin=>p(280)(98),clock=>clock,reset=>reset,s=>p(315)(98),cout=>p(316)(99));
FA_ff_11702:FAff port map(x=>p(278)(99),y=>p(279)(99),Cin=>p(280)(99),clock=>clock,reset=>reset,s=>p(315)(99),cout=>p(316)(100));
FA_ff_11703:FAff port map(x=>p(278)(100),y=>p(279)(100),Cin=>p(280)(100),clock=>clock,reset=>reset,s=>p(315)(100),cout=>p(316)(101));
FA_ff_11704:FAff port map(x=>p(278)(101),y=>p(279)(101),Cin=>p(280)(101),clock=>clock,reset=>reset,s=>p(315)(101),cout=>p(316)(102));
FA_ff_11705:FAff port map(x=>p(278)(102),y=>p(279)(102),Cin=>p(280)(102),clock=>clock,reset=>reset,s=>p(315)(102),cout=>p(316)(103));
FA_ff_11706:FAff port map(x=>p(278)(103),y=>p(279)(103),Cin=>p(280)(103),clock=>clock,reset=>reset,s=>p(315)(103),cout=>p(316)(104));
FA_ff_11707:FAff port map(x=>p(278)(104),y=>p(279)(104),Cin=>p(280)(104),clock=>clock,reset=>reset,s=>p(315)(104),cout=>p(316)(105));
FA_ff_11708:FAff port map(x=>p(278)(105),y=>p(279)(105),Cin=>p(280)(105),clock=>clock,reset=>reset,s=>p(315)(105),cout=>p(316)(106));
FA_ff_11709:FAff port map(x=>p(278)(106),y=>p(279)(106),Cin=>p(280)(106),clock=>clock,reset=>reset,s=>p(315)(106),cout=>p(316)(107));
FA_ff_11710:FAff port map(x=>p(278)(107),y=>p(279)(107),Cin=>p(280)(107),clock=>clock,reset=>reset,s=>p(315)(107),cout=>p(316)(108));
FA_ff_11711:FAff port map(x=>p(278)(108),y=>p(279)(108),Cin=>p(280)(108),clock=>clock,reset=>reset,s=>p(315)(108),cout=>p(316)(109));
FA_ff_11712:FAff port map(x=>p(278)(109),y=>p(279)(109),Cin=>p(280)(109),clock=>clock,reset=>reset,s=>p(315)(109),cout=>p(316)(110));
FA_ff_11713:FAff port map(x=>p(278)(110),y=>p(279)(110),Cin=>p(280)(110),clock=>clock,reset=>reset,s=>p(315)(110),cout=>p(316)(111));
FA_ff_11714:FAff port map(x=>p(278)(111),y=>p(279)(111),Cin=>p(280)(111),clock=>clock,reset=>reset,s=>p(315)(111),cout=>p(316)(112));
FA_ff_11715:FAff port map(x=>p(278)(112),y=>p(279)(112),Cin=>p(280)(112),clock=>clock,reset=>reset,s=>p(315)(112),cout=>p(316)(113));
FA_ff_11716:FAff port map(x=>p(278)(113),y=>p(279)(113),Cin=>p(280)(113),clock=>clock,reset=>reset,s=>p(315)(113),cout=>p(316)(114));
FA_ff_11717:FAff port map(x=>p(278)(114),y=>p(279)(114),Cin=>p(280)(114),clock=>clock,reset=>reset,s=>p(315)(114),cout=>p(316)(115));
FA_ff_11718:FAff port map(x=>p(278)(115),y=>p(279)(115),Cin=>p(280)(115),clock=>clock,reset=>reset,s=>p(315)(115),cout=>p(316)(116));
FA_ff_11719:FAff port map(x=>p(278)(116),y=>p(279)(116),Cin=>p(280)(116),clock=>clock,reset=>reset,s=>p(315)(116),cout=>p(316)(117));
FA_ff_11720:FAff port map(x=>p(278)(117),y=>p(279)(117),Cin=>p(280)(117),clock=>clock,reset=>reset,s=>p(315)(117),cout=>p(316)(118));
FA_ff_11721:FAff port map(x=>p(278)(118),y=>p(279)(118),Cin=>p(280)(118),clock=>clock,reset=>reset,s=>p(315)(118),cout=>p(316)(119));
FA_ff_11722:FAff port map(x=>p(278)(119),y=>p(279)(119),Cin=>p(280)(119),clock=>clock,reset=>reset,s=>p(315)(119),cout=>p(316)(120));
FA_ff_11723:FAff port map(x=>p(278)(120),y=>p(279)(120),Cin=>p(280)(120),clock=>clock,reset=>reset,s=>p(315)(120),cout=>p(316)(121));
FA_ff_11724:FAff port map(x=>p(278)(121),y=>p(279)(121),Cin=>p(280)(121),clock=>clock,reset=>reset,s=>p(315)(121),cout=>p(316)(122));
FA_ff_11725:FAff port map(x=>p(278)(122),y=>p(279)(122),Cin=>p(280)(122),clock=>clock,reset=>reset,s=>p(315)(122),cout=>p(316)(123));
FA_ff_11726:FAff port map(x=>p(278)(123),y=>p(279)(123),Cin=>p(280)(123),clock=>clock,reset=>reset,s=>p(315)(123),cout=>p(316)(124));
FA_ff_11727:FAff port map(x=>p(278)(124),y=>p(279)(124),Cin=>p(280)(124),clock=>clock,reset=>reset,s=>p(315)(124),cout=>p(316)(125));
FA_ff_11728:FAff port map(x=>p(278)(125),y=>p(279)(125),Cin=>p(280)(125),clock=>clock,reset=>reset,s=>p(315)(125),cout=>p(316)(126));
FA_ff_11729:FAff port map(x=>p(278)(126),y=>p(279)(126),Cin=>p(280)(126),clock=>clock,reset=>reset,s=>p(315)(126),cout=>p(316)(127));
FA_ff_11730:FAff port map(x=>p(278)(127),y=>p(279)(127),Cin=>p(280)(127),clock=>clock,reset=>reset,s=>p(315)(127),cout=>p(316)(128));
FA_ff_11731:FAff port map(x=>p(278)(128),y=>p(279)(128),Cin=>p(280)(128),clock=>clock,reset=>reset,s=>p(315)(128),cout=>p(316)(129));
HA_ff_58:HAff port map(x=>p(278)(129),y=>p(279)(129),clock=>clock,reset=>reset,s=>p(315)(129),c=>p(316)(130));
p(317)(0)<=p(282)(0);
HA_ff_59:HAff port map(x=>p(281)(1),y=>p(282)(1),clock=>clock,reset=>reset,s=>p(317)(1),c=>p(318)(2));
FA_ff_11732:FAff port map(x=>p(281)(2),y=>p(282)(2),Cin=>p(283)(2),clock=>clock,reset=>reset,s=>p(317)(2),cout=>p(318)(3));
FA_ff_11733:FAff port map(x=>p(281)(3),y=>p(282)(3),Cin=>p(283)(3),clock=>clock,reset=>reset,s=>p(317)(3),cout=>p(318)(4));
FA_ff_11734:FAff port map(x=>p(281)(4),y=>p(282)(4),Cin=>p(283)(4),clock=>clock,reset=>reset,s=>p(317)(4),cout=>p(318)(5));
FA_ff_11735:FAff port map(x=>p(281)(5),y=>p(282)(5),Cin=>p(283)(5),clock=>clock,reset=>reset,s=>p(317)(5),cout=>p(318)(6));
FA_ff_11736:FAff port map(x=>p(281)(6),y=>p(282)(6),Cin=>p(283)(6),clock=>clock,reset=>reset,s=>p(317)(6),cout=>p(318)(7));
FA_ff_11737:FAff port map(x=>p(281)(7),y=>p(282)(7),Cin=>p(283)(7),clock=>clock,reset=>reset,s=>p(317)(7),cout=>p(318)(8));
FA_ff_11738:FAff port map(x=>p(281)(8),y=>p(282)(8),Cin=>p(283)(8),clock=>clock,reset=>reset,s=>p(317)(8),cout=>p(318)(9));
FA_ff_11739:FAff port map(x=>p(281)(9),y=>p(282)(9),Cin=>p(283)(9),clock=>clock,reset=>reset,s=>p(317)(9),cout=>p(318)(10));
FA_ff_11740:FAff port map(x=>p(281)(10),y=>p(282)(10),Cin=>p(283)(10),clock=>clock,reset=>reset,s=>p(317)(10),cout=>p(318)(11));
FA_ff_11741:FAff port map(x=>p(281)(11),y=>p(282)(11),Cin=>p(283)(11),clock=>clock,reset=>reset,s=>p(317)(11),cout=>p(318)(12));
FA_ff_11742:FAff port map(x=>p(281)(12),y=>p(282)(12),Cin=>p(283)(12),clock=>clock,reset=>reset,s=>p(317)(12),cout=>p(318)(13));
FA_ff_11743:FAff port map(x=>p(281)(13),y=>p(282)(13),Cin=>p(283)(13),clock=>clock,reset=>reset,s=>p(317)(13),cout=>p(318)(14));
FA_ff_11744:FAff port map(x=>p(281)(14),y=>p(282)(14),Cin=>p(283)(14),clock=>clock,reset=>reset,s=>p(317)(14),cout=>p(318)(15));
FA_ff_11745:FAff port map(x=>p(281)(15),y=>p(282)(15),Cin=>p(283)(15),clock=>clock,reset=>reset,s=>p(317)(15),cout=>p(318)(16));
FA_ff_11746:FAff port map(x=>p(281)(16),y=>p(282)(16),Cin=>p(283)(16),clock=>clock,reset=>reset,s=>p(317)(16),cout=>p(318)(17));
FA_ff_11747:FAff port map(x=>p(281)(17),y=>p(282)(17),Cin=>p(283)(17),clock=>clock,reset=>reset,s=>p(317)(17),cout=>p(318)(18));
FA_ff_11748:FAff port map(x=>p(281)(18),y=>p(282)(18),Cin=>p(283)(18),clock=>clock,reset=>reset,s=>p(317)(18),cout=>p(318)(19));
FA_ff_11749:FAff port map(x=>p(281)(19),y=>p(282)(19),Cin=>p(283)(19),clock=>clock,reset=>reset,s=>p(317)(19),cout=>p(318)(20));
FA_ff_11750:FAff port map(x=>p(281)(20),y=>p(282)(20),Cin=>p(283)(20),clock=>clock,reset=>reset,s=>p(317)(20),cout=>p(318)(21));
FA_ff_11751:FAff port map(x=>p(281)(21),y=>p(282)(21),Cin=>p(283)(21),clock=>clock,reset=>reset,s=>p(317)(21),cout=>p(318)(22));
FA_ff_11752:FAff port map(x=>p(281)(22),y=>p(282)(22),Cin=>p(283)(22),clock=>clock,reset=>reset,s=>p(317)(22),cout=>p(318)(23));
FA_ff_11753:FAff port map(x=>p(281)(23),y=>p(282)(23),Cin=>p(283)(23),clock=>clock,reset=>reset,s=>p(317)(23),cout=>p(318)(24));
FA_ff_11754:FAff port map(x=>p(281)(24),y=>p(282)(24),Cin=>p(283)(24),clock=>clock,reset=>reset,s=>p(317)(24),cout=>p(318)(25));
FA_ff_11755:FAff port map(x=>p(281)(25),y=>p(282)(25),Cin=>p(283)(25),clock=>clock,reset=>reset,s=>p(317)(25),cout=>p(318)(26));
FA_ff_11756:FAff port map(x=>p(281)(26),y=>p(282)(26),Cin=>p(283)(26),clock=>clock,reset=>reset,s=>p(317)(26),cout=>p(318)(27));
FA_ff_11757:FAff port map(x=>p(281)(27),y=>p(282)(27),Cin=>p(283)(27),clock=>clock,reset=>reset,s=>p(317)(27),cout=>p(318)(28));
FA_ff_11758:FAff port map(x=>p(281)(28),y=>p(282)(28),Cin=>p(283)(28),clock=>clock,reset=>reset,s=>p(317)(28),cout=>p(318)(29));
FA_ff_11759:FAff port map(x=>p(281)(29),y=>p(282)(29),Cin=>p(283)(29),clock=>clock,reset=>reset,s=>p(317)(29),cout=>p(318)(30));
FA_ff_11760:FAff port map(x=>p(281)(30),y=>p(282)(30),Cin=>p(283)(30),clock=>clock,reset=>reset,s=>p(317)(30),cout=>p(318)(31));
FA_ff_11761:FAff port map(x=>p(281)(31),y=>p(282)(31),Cin=>p(283)(31),clock=>clock,reset=>reset,s=>p(317)(31),cout=>p(318)(32));
FA_ff_11762:FAff port map(x=>p(281)(32),y=>p(282)(32),Cin=>p(283)(32),clock=>clock,reset=>reset,s=>p(317)(32),cout=>p(318)(33));
FA_ff_11763:FAff port map(x=>p(281)(33),y=>p(282)(33),Cin=>p(283)(33),clock=>clock,reset=>reset,s=>p(317)(33),cout=>p(318)(34));
FA_ff_11764:FAff port map(x=>p(281)(34),y=>p(282)(34),Cin=>p(283)(34),clock=>clock,reset=>reset,s=>p(317)(34),cout=>p(318)(35));
FA_ff_11765:FAff port map(x=>p(281)(35),y=>p(282)(35),Cin=>p(283)(35),clock=>clock,reset=>reset,s=>p(317)(35),cout=>p(318)(36));
FA_ff_11766:FAff port map(x=>p(281)(36),y=>p(282)(36),Cin=>p(283)(36),clock=>clock,reset=>reset,s=>p(317)(36),cout=>p(318)(37));
FA_ff_11767:FAff port map(x=>p(281)(37),y=>p(282)(37),Cin=>p(283)(37),clock=>clock,reset=>reset,s=>p(317)(37),cout=>p(318)(38));
FA_ff_11768:FAff port map(x=>p(281)(38),y=>p(282)(38),Cin=>p(283)(38),clock=>clock,reset=>reset,s=>p(317)(38),cout=>p(318)(39));
FA_ff_11769:FAff port map(x=>p(281)(39),y=>p(282)(39),Cin=>p(283)(39),clock=>clock,reset=>reset,s=>p(317)(39),cout=>p(318)(40));
FA_ff_11770:FAff port map(x=>p(281)(40),y=>p(282)(40),Cin=>p(283)(40),clock=>clock,reset=>reset,s=>p(317)(40),cout=>p(318)(41));
FA_ff_11771:FAff port map(x=>p(281)(41),y=>p(282)(41),Cin=>p(283)(41),clock=>clock,reset=>reset,s=>p(317)(41),cout=>p(318)(42));
FA_ff_11772:FAff port map(x=>p(281)(42),y=>p(282)(42),Cin=>p(283)(42),clock=>clock,reset=>reset,s=>p(317)(42),cout=>p(318)(43));
FA_ff_11773:FAff port map(x=>p(281)(43),y=>p(282)(43),Cin=>p(283)(43),clock=>clock,reset=>reset,s=>p(317)(43),cout=>p(318)(44));
FA_ff_11774:FAff port map(x=>p(281)(44),y=>p(282)(44),Cin=>p(283)(44),clock=>clock,reset=>reset,s=>p(317)(44),cout=>p(318)(45));
FA_ff_11775:FAff port map(x=>p(281)(45),y=>p(282)(45),Cin=>p(283)(45),clock=>clock,reset=>reset,s=>p(317)(45),cout=>p(318)(46));
FA_ff_11776:FAff port map(x=>p(281)(46),y=>p(282)(46),Cin=>p(283)(46),clock=>clock,reset=>reset,s=>p(317)(46),cout=>p(318)(47));
FA_ff_11777:FAff port map(x=>p(281)(47),y=>p(282)(47),Cin=>p(283)(47),clock=>clock,reset=>reset,s=>p(317)(47),cout=>p(318)(48));
FA_ff_11778:FAff port map(x=>p(281)(48),y=>p(282)(48),Cin=>p(283)(48),clock=>clock,reset=>reset,s=>p(317)(48),cout=>p(318)(49));
FA_ff_11779:FAff port map(x=>p(281)(49),y=>p(282)(49),Cin=>p(283)(49),clock=>clock,reset=>reset,s=>p(317)(49),cout=>p(318)(50));
FA_ff_11780:FAff port map(x=>p(281)(50),y=>p(282)(50),Cin=>p(283)(50),clock=>clock,reset=>reset,s=>p(317)(50),cout=>p(318)(51));
FA_ff_11781:FAff port map(x=>p(281)(51),y=>p(282)(51),Cin=>p(283)(51),clock=>clock,reset=>reset,s=>p(317)(51),cout=>p(318)(52));
FA_ff_11782:FAff port map(x=>p(281)(52),y=>p(282)(52),Cin=>p(283)(52),clock=>clock,reset=>reset,s=>p(317)(52),cout=>p(318)(53));
FA_ff_11783:FAff port map(x=>p(281)(53),y=>p(282)(53),Cin=>p(283)(53),clock=>clock,reset=>reset,s=>p(317)(53),cout=>p(318)(54));
FA_ff_11784:FAff port map(x=>p(281)(54),y=>p(282)(54),Cin=>p(283)(54),clock=>clock,reset=>reset,s=>p(317)(54),cout=>p(318)(55));
FA_ff_11785:FAff port map(x=>p(281)(55),y=>p(282)(55),Cin=>p(283)(55),clock=>clock,reset=>reset,s=>p(317)(55),cout=>p(318)(56));
FA_ff_11786:FAff port map(x=>p(281)(56),y=>p(282)(56),Cin=>p(283)(56),clock=>clock,reset=>reset,s=>p(317)(56),cout=>p(318)(57));
FA_ff_11787:FAff port map(x=>p(281)(57),y=>p(282)(57),Cin=>p(283)(57),clock=>clock,reset=>reset,s=>p(317)(57),cout=>p(318)(58));
FA_ff_11788:FAff port map(x=>p(281)(58),y=>p(282)(58),Cin=>p(283)(58),clock=>clock,reset=>reset,s=>p(317)(58),cout=>p(318)(59));
FA_ff_11789:FAff port map(x=>p(281)(59),y=>p(282)(59),Cin=>p(283)(59),clock=>clock,reset=>reset,s=>p(317)(59),cout=>p(318)(60));
FA_ff_11790:FAff port map(x=>p(281)(60),y=>p(282)(60),Cin=>p(283)(60),clock=>clock,reset=>reset,s=>p(317)(60),cout=>p(318)(61));
FA_ff_11791:FAff port map(x=>p(281)(61),y=>p(282)(61),Cin=>p(283)(61),clock=>clock,reset=>reset,s=>p(317)(61),cout=>p(318)(62));
FA_ff_11792:FAff port map(x=>p(281)(62),y=>p(282)(62),Cin=>p(283)(62),clock=>clock,reset=>reset,s=>p(317)(62),cout=>p(318)(63));
FA_ff_11793:FAff port map(x=>p(281)(63),y=>p(282)(63),Cin=>p(283)(63),clock=>clock,reset=>reset,s=>p(317)(63),cout=>p(318)(64));
FA_ff_11794:FAff port map(x=>p(281)(64),y=>p(282)(64),Cin=>p(283)(64),clock=>clock,reset=>reset,s=>p(317)(64),cout=>p(318)(65));
FA_ff_11795:FAff port map(x=>p(281)(65),y=>p(282)(65),Cin=>p(283)(65),clock=>clock,reset=>reset,s=>p(317)(65),cout=>p(318)(66));
FA_ff_11796:FAff port map(x=>p(281)(66),y=>p(282)(66),Cin=>p(283)(66),clock=>clock,reset=>reset,s=>p(317)(66),cout=>p(318)(67));
FA_ff_11797:FAff port map(x=>p(281)(67),y=>p(282)(67),Cin=>p(283)(67),clock=>clock,reset=>reset,s=>p(317)(67),cout=>p(318)(68));
FA_ff_11798:FAff port map(x=>p(281)(68),y=>p(282)(68),Cin=>p(283)(68),clock=>clock,reset=>reset,s=>p(317)(68),cout=>p(318)(69));
FA_ff_11799:FAff port map(x=>p(281)(69),y=>p(282)(69),Cin=>p(283)(69),clock=>clock,reset=>reset,s=>p(317)(69),cout=>p(318)(70));
FA_ff_11800:FAff port map(x=>p(281)(70),y=>p(282)(70),Cin=>p(283)(70),clock=>clock,reset=>reset,s=>p(317)(70),cout=>p(318)(71));
FA_ff_11801:FAff port map(x=>p(281)(71),y=>p(282)(71),Cin=>p(283)(71),clock=>clock,reset=>reset,s=>p(317)(71),cout=>p(318)(72));
FA_ff_11802:FAff port map(x=>p(281)(72),y=>p(282)(72),Cin=>p(283)(72),clock=>clock,reset=>reset,s=>p(317)(72),cout=>p(318)(73));
FA_ff_11803:FAff port map(x=>p(281)(73),y=>p(282)(73),Cin=>p(283)(73),clock=>clock,reset=>reset,s=>p(317)(73),cout=>p(318)(74));
FA_ff_11804:FAff port map(x=>p(281)(74),y=>p(282)(74),Cin=>p(283)(74),clock=>clock,reset=>reset,s=>p(317)(74),cout=>p(318)(75));
FA_ff_11805:FAff port map(x=>p(281)(75),y=>p(282)(75),Cin=>p(283)(75),clock=>clock,reset=>reset,s=>p(317)(75),cout=>p(318)(76));
FA_ff_11806:FAff port map(x=>p(281)(76),y=>p(282)(76),Cin=>p(283)(76),clock=>clock,reset=>reset,s=>p(317)(76),cout=>p(318)(77));
FA_ff_11807:FAff port map(x=>p(281)(77),y=>p(282)(77),Cin=>p(283)(77),clock=>clock,reset=>reset,s=>p(317)(77),cout=>p(318)(78));
FA_ff_11808:FAff port map(x=>p(281)(78),y=>p(282)(78),Cin=>p(283)(78),clock=>clock,reset=>reset,s=>p(317)(78),cout=>p(318)(79));
FA_ff_11809:FAff port map(x=>p(281)(79),y=>p(282)(79),Cin=>p(283)(79),clock=>clock,reset=>reset,s=>p(317)(79),cout=>p(318)(80));
FA_ff_11810:FAff port map(x=>p(281)(80),y=>p(282)(80),Cin=>p(283)(80),clock=>clock,reset=>reset,s=>p(317)(80),cout=>p(318)(81));
FA_ff_11811:FAff port map(x=>p(281)(81),y=>p(282)(81),Cin=>p(283)(81),clock=>clock,reset=>reset,s=>p(317)(81),cout=>p(318)(82));
FA_ff_11812:FAff port map(x=>p(281)(82),y=>p(282)(82),Cin=>p(283)(82),clock=>clock,reset=>reset,s=>p(317)(82),cout=>p(318)(83));
FA_ff_11813:FAff port map(x=>p(281)(83),y=>p(282)(83),Cin=>p(283)(83),clock=>clock,reset=>reset,s=>p(317)(83),cout=>p(318)(84));
FA_ff_11814:FAff port map(x=>p(281)(84),y=>p(282)(84),Cin=>p(283)(84),clock=>clock,reset=>reset,s=>p(317)(84),cout=>p(318)(85));
FA_ff_11815:FAff port map(x=>p(281)(85),y=>p(282)(85),Cin=>p(283)(85),clock=>clock,reset=>reset,s=>p(317)(85),cout=>p(318)(86));
FA_ff_11816:FAff port map(x=>p(281)(86),y=>p(282)(86),Cin=>p(283)(86),clock=>clock,reset=>reset,s=>p(317)(86),cout=>p(318)(87));
FA_ff_11817:FAff port map(x=>p(281)(87),y=>p(282)(87),Cin=>p(283)(87),clock=>clock,reset=>reset,s=>p(317)(87),cout=>p(318)(88));
FA_ff_11818:FAff port map(x=>p(281)(88),y=>p(282)(88),Cin=>p(283)(88),clock=>clock,reset=>reset,s=>p(317)(88),cout=>p(318)(89));
FA_ff_11819:FAff port map(x=>p(281)(89),y=>p(282)(89),Cin=>p(283)(89),clock=>clock,reset=>reset,s=>p(317)(89),cout=>p(318)(90));
FA_ff_11820:FAff port map(x=>p(281)(90),y=>p(282)(90),Cin=>p(283)(90),clock=>clock,reset=>reset,s=>p(317)(90),cout=>p(318)(91));
FA_ff_11821:FAff port map(x=>p(281)(91),y=>p(282)(91),Cin=>p(283)(91),clock=>clock,reset=>reset,s=>p(317)(91),cout=>p(318)(92));
FA_ff_11822:FAff port map(x=>p(281)(92),y=>p(282)(92),Cin=>p(283)(92),clock=>clock,reset=>reset,s=>p(317)(92),cout=>p(318)(93));
FA_ff_11823:FAff port map(x=>p(281)(93),y=>p(282)(93),Cin=>p(283)(93),clock=>clock,reset=>reset,s=>p(317)(93),cout=>p(318)(94));
FA_ff_11824:FAff port map(x=>p(281)(94),y=>p(282)(94),Cin=>p(283)(94),clock=>clock,reset=>reset,s=>p(317)(94),cout=>p(318)(95));
FA_ff_11825:FAff port map(x=>p(281)(95),y=>p(282)(95),Cin=>p(283)(95),clock=>clock,reset=>reset,s=>p(317)(95),cout=>p(318)(96));
FA_ff_11826:FAff port map(x=>p(281)(96),y=>p(282)(96),Cin=>p(283)(96),clock=>clock,reset=>reset,s=>p(317)(96),cout=>p(318)(97));
FA_ff_11827:FAff port map(x=>p(281)(97),y=>p(282)(97),Cin=>p(283)(97),clock=>clock,reset=>reset,s=>p(317)(97),cout=>p(318)(98));
FA_ff_11828:FAff port map(x=>p(281)(98),y=>p(282)(98),Cin=>p(283)(98),clock=>clock,reset=>reset,s=>p(317)(98),cout=>p(318)(99));
FA_ff_11829:FAff port map(x=>p(281)(99),y=>p(282)(99),Cin=>p(283)(99),clock=>clock,reset=>reset,s=>p(317)(99),cout=>p(318)(100));
FA_ff_11830:FAff port map(x=>p(281)(100),y=>p(282)(100),Cin=>p(283)(100),clock=>clock,reset=>reset,s=>p(317)(100),cout=>p(318)(101));
FA_ff_11831:FAff port map(x=>p(281)(101),y=>p(282)(101),Cin=>p(283)(101),clock=>clock,reset=>reset,s=>p(317)(101),cout=>p(318)(102));
FA_ff_11832:FAff port map(x=>p(281)(102),y=>p(282)(102),Cin=>p(283)(102),clock=>clock,reset=>reset,s=>p(317)(102),cout=>p(318)(103));
FA_ff_11833:FAff port map(x=>p(281)(103),y=>p(282)(103),Cin=>p(283)(103),clock=>clock,reset=>reset,s=>p(317)(103),cout=>p(318)(104));
FA_ff_11834:FAff port map(x=>p(281)(104),y=>p(282)(104),Cin=>p(283)(104),clock=>clock,reset=>reset,s=>p(317)(104),cout=>p(318)(105));
FA_ff_11835:FAff port map(x=>p(281)(105),y=>p(282)(105),Cin=>p(283)(105),clock=>clock,reset=>reset,s=>p(317)(105),cout=>p(318)(106));
FA_ff_11836:FAff port map(x=>p(281)(106),y=>p(282)(106),Cin=>p(283)(106),clock=>clock,reset=>reset,s=>p(317)(106),cout=>p(318)(107));
FA_ff_11837:FAff port map(x=>p(281)(107),y=>p(282)(107),Cin=>p(283)(107),clock=>clock,reset=>reset,s=>p(317)(107),cout=>p(318)(108));
FA_ff_11838:FAff port map(x=>p(281)(108),y=>p(282)(108),Cin=>p(283)(108),clock=>clock,reset=>reset,s=>p(317)(108),cout=>p(318)(109));
FA_ff_11839:FAff port map(x=>p(281)(109),y=>p(282)(109),Cin=>p(283)(109),clock=>clock,reset=>reset,s=>p(317)(109),cout=>p(318)(110));
FA_ff_11840:FAff port map(x=>p(281)(110),y=>p(282)(110),Cin=>p(283)(110),clock=>clock,reset=>reset,s=>p(317)(110),cout=>p(318)(111));
FA_ff_11841:FAff port map(x=>p(281)(111),y=>p(282)(111),Cin=>p(283)(111),clock=>clock,reset=>reset,s=>p(317)(111),cout=>p(318)(112));
FA_ff_11842:FAff port map(x=>p(281)(112),y=>p(282)(112),Cin=>p(283)(112),clock=>clock,reset=>reset,s=>p(317)(112),cout=>p(318)(113));
FA_ff_11843:FAff port map(x=>p(281)(113),y=>p(282)(113),Cin=>p(283)(113),clock=>clock,reset=>reset,s=>p(317)(113),cout=>p(318)(114));
FA_ff_11844:FAff port map(x=>p(281)(114),y=>p(282)(114),Cin=>p(283)(114),clock=>clock,reset=>reset,s=>p(317)(114),cout=>p(318)(115));
FA_ff_11845:FAff port map(x=>p(281)(115),y=>p(282)(115),Cin=>p(283)(115),clock=>clock,reset=>reset,s=>p(317)(115),cout=>p(318)(116));
FA_ff_11846:FAff port map(x=>p(281)(116),y=>p(282)(116),Cin=>p(283)(116),clock=>clock,reset=>reset,s=>p(317)(116),cout=>p(318)(117));
FA_ff_11847:FAff port map(x=>p(281)(117),y=>p(282)(117),Cin=>p(283)(117),clock=>clock,reset=>reset,s=>p(317)(117),cout=>p(318)(118));
FA_ff_11848:FAff port map(x=>p(281)(118),y=>p(282)(118),Cin=>p(283)(118),clock=>clock,reset=>reset,s=>p(317)(118),cout=>p(318)(119));
FA_ff_11849:FAff port map(x=>p(281)(119),y=>p(282)(119),Cin=>p(283)(119),clock=>clock,reset=>reset,s=>p(317)(119),cout=>p(318)(120));
FA_ff_11850:FAff port map(x=>p(281)(120),y=>p(282)(120),Cin=>p(283)(120),clock=>clock,reset=>reset,s=>p(317)(120),cout=>p(318)(121));
FA_ff_11851:FAff port map(x=>p(281)(121),y=>p(282)(121),Cin=>p(283)(121),clock=>clock,reset=>reset,s=>p(317)(121),cout=>p(318)(122));
FA_ff_11852:FAff port map(x=>p(281)(122),y=>p(282)(122),Cin=>p(283)(122),clock=>clock,reset=>reset,s=>p(317)(122),cout=>p(318)(123));
FA_ff_11853:FAff port map(x=>p(281)(123),y=>p(282)(123),Cin=>p(283)(123),clock=>clock,reset=>reset,s=>p(317)(123),cout=>p(318)(124));
FA_ff_11854:FAff port map(x=>p(281)(124),y=>p(282)(124),Cin=>p(283)(124),clock=>clock,reset=>reset,s=>p(317)(124),cout=>p(318)(125));
FA_ff_11855:FAff port map(x=>p(281)(125),y=>p(282)(125),Cin=>p(283)(125),clock=>clock,reset=>reset,s=>p(317)(125),cout=>p(318)(126));
FA_ff_11856:FAff port map(x=>p(281)(126),y=>p(282)(126),Cin=>p(283)(126),clock=>clock,reset=>reset,s=>p(317)(126),cout=>p(318)(127));
FA_ff_11857:FAff port map(x=>p(281)(127),y=>p(282)(127),Cin=>p(283)(127),clock=>clock,reset=>reset,s=>p(317)(127),cout=>p(318)(128));
FA_ff_11858:FAff port map(x=>p(281)(128),y=>p(282)(128),Cin=>p(283)(128),clock=>clock,reset=>reset,s=>p(317)(128),cout=>p(318)(129));
FA_ff_11859:FAff port map(x=>p(281)(129),y=>p(282)(129),Cin=>p(283)(129),clock=>clock,reset=>reset,s=>p(317)(129),cout=>p(318)(130));
HA_ff_60:HAff port map(x=>p(284)(0),y=>p(286)(0),clock=>clock,reset=>reset,s=>p(319)(0),c=>p(320)(1));
FA_ff_11860:FAff port map(x=>p(284)(1),y=>p(285)(1),Cin=>p(286)(1),clock=>clock,reset=>reset,s=>p(319)(1),cout=>p(320)(2));
FA_ff_11861:FAff port map(x=>p(284)(2),y=>p(285)(2),Cin=>p(286)(2),clock=>clock,reset=>reset,s=>p(319)(2),cout=>p(320)(3));
FA_ff_11862:FAff port map(x=>p(284)(3),y=>p(285)(3),Cin=>p(286)(3),clock=>clock,reset=>reset,s=>p(319)(3),cout=>p(320)(4));
FA_ff_11863:FAff port map(x=>p(284)(4),y=>p(285)(4),Cin=>p(286)(4),clock=>clock,reset=>reset,s=>p(319)(4),cout=>p(320)(5));
FA_ff_11864:FAff port map(x=>p(284)(5),y=>p(285)(5),Cin=>p(286)(5),clock=>clock,reset=>reset,s=>p(319)(5),cout=>p(320)(6));
FA_ff_11865:FAff port map(x=>p(284)(6),y=>p(285)(6),Cin=>p(286)(6),clock=>clock,reset=>reset,s=>p(319)(6),cout=>p(320)(7));
FA_ff_11866:FAff port map(x=>p(284)(7),y=>p(285)(7),Cin=>p(286)(7),clock=>clock,reset=>reset,s=>p(319)(7),cout=>p(320)(8));
FA_ff_11867:FAff port map(x=>p(284)(8),y=>p(285)(8),Cin=>p(286)(8),clock=>clock,reset=>reset,s=>p(319)(8),cout=>p(320)(9));
FA_ff_11868:FAff port map(x=>p(284)(9),y=>p(285)(9),Cin=>p(286)(9),clock=>clock,reset=>reset,s=>p(319)(9),cout=>p(320)(10));
FA_ff_11869:FAff port map(x=>p(284)(10),y=>p(285)(10),Cin=>p(286)(10),clock=>clock,reset=>reset,s=>p(319)(10),cout=>p(320)(11));
FA_ff_11870:FAff port map(x=>p(284)(11),y=>p(285)(11),Cin=>p(286)(11),clock=>clock,reset=>reset,s=>p(319)(11),cout=>p(320)(12));
FA_ff_11871:FAff port map(x=>p(284)(12),y=>p(285)(12),Cin=>p(286)(12),clock=>clock,reset=>reset,s=>p(319)(12),cout=>p(320)(13));
FA_ff_11872:FAff port map(x=>p(284)(13),y=>p(285)(13),Cin=>p(286)(13),clock=>clock,reset=>reset,s=>p(319)(13),cout=>p(320)(14));
FA_ff_11873:FAff port map(x=>p(284)(14),y=>p(285)(14),Cin=>p(286)(14),clock=>clock,reset=>reset,s=>p(319)(14),cout=>p(320)(15));
FA_ff_11874:FAff port map(x=>p(284)(15),y=>p(285)(15),Cin=>p(286)(15),clock=>clock,reset=>reset,s=>p(319)(15),cout=>p(320)(16));
FA_ff_11875:FAff port map(x=>p(284)(16),y=>p(285)(16),Cin=>p(286)(16),clock=>clock,reset=>reset,s=>p(319)(16),cout=>p(320)(17));
FA_ff_11876:FAff port map(x=>p(284)(17),y=>p(285)(17),Cin=>p(286)(17),clock=>clock,reset=>reset,s=>p(319)(17),cout=>p(320)(18));
FA_ff_11877:FAff port map(x=>p(284)(18),y=>p(285)(18),Cin=>p(286)(18),clock=>clock,reset=>reset,s=>p(319)(18),cout=>p(320)(19));
FA_ff_11878:FAff port map(x=>p(284)(19),y=>p(285)(19),Cin=>p(286)(19),clock=>clock,reset=>reset,s=>p(319)(19),cout=>p(320)(20));
FA_ff_11879:FAff port map(x=>p(284)(20),y=>p(285)(20),Cin=>p(286)(20),clock=>clock,reset=>reset,s=>p(319)(20),cout=>p(320)(21));
FA_ff_11880:FAff port map(x=>p(284)(21),y=>p(285)(21),Cin=>p(286)(21),clock=>clock,reset=>reset,s=>p(319)(21),cout=>p(320)(22));
FA_ff_11881:FAff port map(x=>p(284)(22),y=>p(285)(22),Cin=>p(286)(22),clock=>clock,reset=>reset,s=>p(319)(22),cout=>p(320)(23));
FA_ff_11882:FAff port map(x=>p(284)(23),y=>p(285)(23),Cin=>p(286)(23),clock=>clock,reset=>reset,s=>p(319)(23),cout=>p(320)(24));
FA_ff_11883:FAff port map(x=>p(284)(24),y=>p(285)(24),Cin=>p(286)(24),clock=>clock,reset=>reset,s=>p(319)(24),cout=>p(320)(25));
FA_ff_11884:FAff port map(x=>p(284)(25),y=>p(285)(25),Cin=>p(286)(25),clock=>clock,reset=>reset,s=>p(319)(25),cout=>p(320)(26));
FA_ff_11885:FAff port map(x=>p(284)(26),y=>p(285)(26),Cin=>p(286)(26),clock=>clock,reset=>reset,s=>p(319)(26),cout=>p(320)(27));
FA_ff_11886:FAff port map(x=>p(284)(27),y=>p(285)(27),Cin=>p(286)(27),clock=>clock,reset=>reset,s=>p(319)(27),cout=>p(320)(28));
FA_ff_11887:FAff port map(x=>p(284)(28),y=>p(285)(28),Cin=>p(286)(28),clock=>clock,reset=>reset,s=>p(319)(28),cout=>p(320)(29));
FA_ff_11888:FAff port map(x=>p(284)(29),y=>p(285)(29),Cin=>p(286)(29),clock=>clock,reset=>reset,s=>p(319)(29),cout=>p(320)(30));
FA_ff_11889:FAff port map(x=>p(284)(30),y=>p(285)(30),Cin=>p(286)(30),clock=>clock,reset=>reset,s=>p(319)(30),cout=>p(320)(31));
FA_ff_11890:FAff port map(x=>p(284)(31),y=>p(285)(31),Cin=>p(286)(31),clock=>clock,reset=>reset,s=>p(319)(31),cout=>p(320)(32));
FA_ff_11891:FAff port map(x=>p(284)(32),y=>p(285)(32),Cin=>p(286)(32),clock=>clock,reset=>reset,s=>p(319)(32),cout=>p(320)(33));
FA_ff_11892:FAff port map(x=>p(284)(33),y=>p(285)(33),Cin=>p(286)(33),clock=>clock,reset=>reset,s=>p(319)(33),cout=>p(320)(34));
FA_ff_11893:FAff port map(x=>p(284)(34),y=>p(285)(34),Cin=>p(286)(34),clock=>clock,reset=>reset,s=>p(319)(34),cout=>p(320)(35));
FA_ff_11894:FAff port map(x=>p(284)(35),y=>p(285)(35),Cin=>p(286)(35),clock=>clock,reset=>reset,s=>p(319)(35),cout=>p(320)(36));
FA_ff_11895:FAff port map(x=>p(284)(36),y=>p(285)(36),Cin=>p(286)(36),clock=>clock,reset=>reset,s=>p(319)(36),cout=>p(320)(37));
FA_ff_11896:FAff port map(x=>p(284)(37),y=>p(285)(37),Cin=>p(286)(37),clock=>clock,reset=>reset,s=>p(319)(37),cout=>p(320)(38));
FA_ff_11897:FAff port map(x=>p(284)(38),y=>p(285)(38),Cin=>p(286)(38),clock=>clock,reset=>reset,s=>p(319)(38),cout=>p(320)(39));
FA_ff_11898:FAff port map(x=>p(284)(39),y=>p(285)(39),Cin=>p(286)(39),clock=>clock,reset=>reset,s=>p(319)(39),cout=>p(320)(40));
FA_ff_11899:FAff port map(x=>p(284)(40),y=>p(285)(40),Cin=>p(286)(40),clock=>clock,reset=>reset,s=>p(319)(40),cout=>p(320)(41));
FA_ff_11900:FAff port map(x=>p(284)(41),y=>p(285)(41),Cin=>p(286)(41),clock=>clock,reset=>reset,s=>p(319)(41),cout=>p(320)(42));
FA_ff_11901:FAff port map(x=>p(284)(42),y=>p(285)(42),Cin=>p(286)(42),clock=>clock,reset=>reset,s=>p(319)(42),cout=>p(320)(43));
FA_ff_11902:FAff port map(x=>p(284)(43),y=>p(285)(43),Cin=>p(286)(43),clock=>clock,reset=>reset,s=>p(319)(43),cout=>p(320)(44));
FA_ff_11903:FAff port map(x=>p(284)(44),y=>p(285)(44),Cin=>p(286)(44),clock=>clock,reset=>reset,s=>p(319)(44),cout=>p(320)(45));
FA_ff_11904:FAff port map(x=>p(284)(45),y=>p(285)(45),Cin=>p(286)(45),clock=>clock,reset=>reset,s=>p(319)(45),cout=>p(320)(46));
FA_ff_11905:FAff port map(x=>p(284)(46),y=>p(285)(46),Cin=>p(286)(46),clock=>clock,reset=>reset,s=>p(319)(46),cout=>p(320)(47));
FA_ff_11906:FAff port map(x=>p(284)(47),y=>p(285)(47),Cin=>p(286)(47),clock=>clock,reset=>reset,s=>p(319)(47),cout=>p(320)(48));
FA_ff_11907:FAff port map(x=>p(284)(48),y=>p(285)(48),Cin=>p(286)(48),clock=>clock,reset=>reset,s=>p(319)(48),cout=>p(320)(49));
FA_ff_11908:FAff port map(x=>p(284)(49),y=>p(285)(49),Cin=>p(286)(49),clock=>clock,reset=>reset,s=>p(319)(49),cout=>p(320)(50));
FA_ff_11909:FAff port map(x=>p(284)(50),y=>p(285)(50),Cin=>p(286)(50),clock=>clock,reset=>reset,s=>p(319)(50),cout=>p(320)(51));
FA_ff_11910:FAff port map(x=>p(284)(51),y=>p(285)(51),Cin=>p(286)(51),clock=>clock,reset=>reset,s=>p(319)(51),cout=>p(320)(52));
FA_ff_11911:FAff port map(x=>p(284)(52),y=>p(285)(52),Cin=>p(286)(52),clock=>clock,reset=>reset,s=>p(319)(52),cout=>p(320)(53));
FA_ff_11912:FAff port map(x=>p(284)(53),y=>p(285)(53),Cin=>p(286)(53),clock=>clock,reset=>reset,s=>p(319)(53),cout=>p(320)(54));
FA_ff_11913:FAff port map(x=>p(284)(54),y=>p(285)(54),Cin=>p(286)(54),clock=>clock,reset=>reset,s=>p(319)(54),cout=>p(320)(55));
FA_ff_11914:FAff port map(x=>p(284)(55),y=>p(285)(55),Cin=>p(286)(55),clock=>clock,reset=>reset,s=>p(319)(55),cout=>p(320)(56));
FA_ff_11915:FAff port map(x=>p(284)(56),y=>p(285)(56),Cin=>p(286)(56),clock=>clock,reset=>reset,s=>p(319)(56),cout=>p(320)(57));
FA_ff_11916:FAff port map(x=>p(284)(57),y=>p(285)(57),Cin=>p(286)(57),clock=>clock,reset=>reset,s=>p(319)(57),cout=>p(320)(58));
FA_ff_11917:FAff port map(x=>p(284)(58),y=>p(285)(58),Cin=>p(286)(58),clock=>clock,reset=>reset,s=>p(319)(58),cout=>p(320)(59));
FA_ff_11918:FAff port map(x=>p(284)(59),y=>p(285)(59),Cin=>p(286)(59),clock=>clock,reset=>reset,s=>p(319)(59),cout=>p(320)(60));
FA_ff_11919:FAff port map(x=>p(284)(60),y=>p(285)(60),Cin=>p(286)(60),clock=>clock,reset=>reset,s=>p(319)(60),cout=>p(320)(61));
FA_ff_11920:FAff port map(x=>p(284)(61),y=>p(285)(61),Cin=>p(286)(61),clock=>clock,reset=>reset,s=>p(319)(61),cout=>p(320)(62));
FA_ff_11921:FAff port map(x=>p(284)(62),y=>p(285)(62),Cin=>p(286)(62),clock=>clock,reset=>reset,s=>p(319)(62),cout=>p(320)(63));
FA_ff_11922:FAff port map(x=>p(284)(63),y=>p(285)(63),Cin=>p(286)(63),clock=>clock,reset=>reset,s=>p(319)(63),cout=>p(320)(64));
FA_ff_11923:FAff port map(x=>p(284)(64),y=>p(285)(64),Cin=>p(286)(64),clock=>clock,reset=>reset,s=>p(319)(64),cout=>p(320)(65));
FA_ff_11924:FAff port map(x=>p(284)(65),y=>p(285)(65),Cin=>p(286)(65),clock=>clock,reset=>reset,s=>p(319)(65),cout=>p(320)(66));
FA_ff_11925:FAff port map(x=>p(284)(66),y=>p(285)(66),Cin=>p(286)(66),clock=>clock,reset=>reset,s=>p(319)(66),cout=>p(320)(67));
FA_ff_11926:FAff port map(x=>p(284)(67),y=>p(285)(67),Cin=>p(286)(67),clock=>clock,reset=>reset,s=>p(319)(67),cout=>p(320)(68));
FA_ff_11927:FAff port map(x=>p(284)(68),y=>p(285)(68),Cin=>p(286)(68),clock=>clock,reset=>reset,s=>p(319)(68),cout=>p(320)(69));
FA_ff_11928:FAff port map(x=>p(284)(69),y=>p(285)(69),Cin=>p(286)(69),clock=>clock,reset=>reset,s=>p(319)(69),cout=>p(320)(70));
FA_ff_11929:FAff port map(x=>p(284)(70),y=>p(285)(70),Cin=>p(286)(70),clock=>clock,reset=>reset,s=>p(319)(70),cout=>p(320)(71));
FA_ff_11930:FAff port map(x=>p(284)(71),y=>p(285)(71),Cin=>p(286)(71),clock=>clock,reset=>reset,s=>p(319)(71),cout=>p(320)(72));
FA_ff_11931:FAff port map(x=>p(284)(72),y=>p(285)(72),Cin=>p(286)(72),clock=>clock,reset=>reset,s=>p(319)(72),cout=>p(320)(73));
FA_ff_11932:FAff port map(x=>p(284)(73),y=>p(285)(73),Cin=>p(286)(73),clock=>clock,reset=>reset,s=>p(319)(73),cout=>p(320)(74));
FA_ff_11933:FAff port map(x=>p(284)(74),y=>p(285)(74),Cin=>p(286)(74),clock=>clock,reset=>reset,s=>p(319)(74),cout=>p(320)(75));
FA_ff_11934:FAff port map(x=>p(284)(75),y=>p(285)(75),Cin=>p(286)(75),clock=>clock,reset=>reset,s=>p(319)(75),cout=>p(320)(76));
FA_ff_11935:FAff port map(x=>p(284)(76),y=>p(285)(76),Cin=>p(286)(76),clock=>clock,reset=>reset,s=>p(319)(76),cout=>p(320)(77));
FA_ff_11936:FAff port map(x=>p(284)(77),y=>p(285)(77),Cin=>p(286)(77),clock=>clock,reset=>reset,s=>p(319)(77),cout=>p(320)(78));
FA_ff_11937:FAff port map(x=>p(284)(78),y=>p(285)(78),Cin=>p(286)(78),clock=>clock,reset=>reset,s=>p(319)(78),cout=>p(320)(79));
FA_ff_11938:FAff port map(x=>p(284)(79),y=>p(285)(79),Cin=>p(286)(79),clock=>clock,reset=>reset,s=>p(319)(79),cout=>p(320)(80));
FA_ff_11939:FAff port map(x=>p(284)(80),y=>p(285)(80),Cin=>p(286)(80),clock=>clock,reset=>reset,s=>p(319)(80),cout=>p(320)(81));
FA_ff_11940:FAff port map(x=>p(284)(81),y=>p(285)(81),Cin=>p(286)(81),clock=>clock,reset=>reset,s=>p(319)(81),cout=>p(320)(82));
FA_ff_11941:FAff port map(x=>p(284)(82),y=>p(285)(82),Cin=>p(286)(82),clock=>clock,reset=>reset,s=>p(319)(82),cout=>p(320)(83));
FA_ff_11942:FAff port map(x=>p(284)(83),y=>p(285)(83),Cin=>p(286)(83),clock=>clock,reset=>reset,s=>p(319)(83),cout=>p(320)(84));
FA_ff_11943:FAff port map(x=>p(284)(84),y=>p(285)(84),Cin=>p(286)(84),clock=>clock,reset=>reset,s=>p(319)(84),cout=>p(320)(85));
FA_ff_11944:FAff port map(x=>p(284)(85),y=>p(285)(85),Cin=>p(286)(85),clock=>clock,reset=>reset,s=>p(319)(85),cout=>p(320)(86));
FA_ff_11945:FAff port map(x=>p(284)(86),y=>p(285)(86),Cin=>p(286)(86),clock=>clock,reset=>reset,s=>p(319)(86),cout=>p(320)(87));
FA_ff_11946:FAff port map(x=>p(284)(87),y=>p(285)(87),Cin=>p(286)(87),clock=>clock,reset=>reset,s=>p(319)(87),cout=>p(320)(88));
FA_ff_11947:FAff port map(x=>p(284)(88),y=>p(285)(88),Cin=>p(286)(88),clock=>clock,reset=>reset,s=>p(319)(88),cout=>p(320)(89));
FA_ff_11948:FAff port map(x=>p(284)(89),y=>p(285)(89),Cin=>p(286)(89),clock=>clock,reset=>reset,s=>p(319)(89),cout=>p(320)(90));
FA_ff_11949:FAff port map(x=>p(284)(90),y=>p(285)(90),Cin=>p(286)(90),clock=>clock,reset=>reset,s=>p(319)(90),cout=>p(320)(91));
FA_ff_11950:FAff port map(x=>p(284)(91),y=>p(285)(91),Cin=>p(286)(91),clock=>clock,reset=>reset,s=>p(319)(91),cout=>p(320)(92));
FA_ff_11951:FAff port map(x=>p(284)(92),y=>p(285)(92),Cin=>p(286)(92),clock=>clock,reset=>reset,s=>p(319)(92),cout=>p(320)(93));
FA_ff_11952:FAff port map(x=>p(284)(93),y=>p(285)(93),Cin=>p(286)(93),clock=>clock,reset=>reset,s=>p(319)(93),cout=>p(320)(94));
FA_ff_11953:FAff port map(x=>p(284)(94),y=>p(285)(94),Cin=>p(286)(94),clock=>clock,reset=>reset,s=>p(319)(94),cout=>p(320)(95));
FA_ff_11954:FAff port map(x=>p(284)(95),y=>p(285)(95),Cin=>p(286)(95),clock=>clock,reset=>reset,s=>p(319)(95),cout=>p(320)(96));
FA_ff_11955:FAff port map(x=>p(284)(96),y=>p(285)(96),Cin=>p(286)(96),clock=>clock,reset=>reset,s=>p(319)(96),cout=>p(320)(97));
FA_ff_11956:FAff port map(x=>p(284)(97),y=>p(285)(97),Cin=>p(286)(97),clock=>clock,reset=>reset,s=>p(319)(97),cout=>p(320)(98));
FA_ff_11957:FAff port map(x=>p(284)(98),y=>p(285)(98),Cin=>p(286)(98),clock=>clock,reset=>reset,s=>p(319)(98),cout=>p(320)(99));
FA_ff_11958:FAff port map(x=>p(284)(99),y=>p(285)(99),Cin=>p(286)(99),clock=>clock,reset=>reset,s=>p(319)(99),cout=>p(320)(100));
FA_ff_11959:FAff port map(x=>p(284)(100),y=>p(285)(100),Cin=>p(286)(100),clock=>clock,reset=>reset,s=>p(319)(100),cout=>p(320)(101));
FA_ff_11960:FAff port map(x=>p(284)(101),y=>p(285)(101),Cin=>p(286)(101),clock=>clock,reset=>reset,s=>p(319)(101),cout=>p(320)(102));
FA_ff_11961:FAff port map(x=>p(284)(102),y=>p(285)(102),Cin=>p(286)(102),clock=>clock,reset=>reset,s=>p(319)(102),cout=>p(320)(103));
FA_ff_11962:FAff port map(x=>p(284)(103),y=>p(285)(103),Cin=>p(286)(103),clock=>clock,reset=>reset,s=>p(319)(103),cout=>p(320)(104));
FA_ff_11963:FAff port map(x=>p(284)(104),y=>p(285)(104),Cin=>p(286)(104),clock=>clock,reset=>reset,s=>p(319)(104),cout=>p(320)(105));
FA_ff_11964:FAff port map(x=>p(284)(105),y=>p(285)(105),Cin=>p(286)(105),clock=>clock,reset=>reset,s=>p(319)(105),cout=>p(320)(106));
FA_ff_11965:FAff port map(x=>p(284)(106),y=>p(285)(106),Cin=>p(286)(106),clock=>clock,reset=>reset,s=>p(319)(106),cout=>p(320)(107));
FA_ff_11966:FAff port map(x=>p(284)(107),y=>p(285)(107),Cin=>p(286)(107),clock=>clock,reset=>reset,s=>p(319)(107),cout=>p(320)(108));
FA_ff_11967:FAff port map(x=>p(284)(108),y=>p(285)(108),Cin=>p(286)(108),clock=>clock,reset=>reset,s=>p(319)(108),cout=>p(320)(109));
FA_ff_11968:FAff port map(x=>p(284)(109),y=>p(285)(109),Cin=>p(286)(109),clock=>clock,reset=>reset,s=>p(319)(109),cout=>p(320)(110));
FA_ff_11969:FAff port map(x=>p(284)(110),y=>p(285)(110),Cin=>p(286)(110),clock=>clock,reset=>reset,s=>p(319)(110),cout=>p(320)(111));
FA_ff_11970:FAff port map(x=>p(284)(111),y=>p(285)(111),Cin=>p(286)(111),clock=>clock,reset=>reset,s=>p(319)(111),cout=>p(320)(112));
FA_ff_11971:FAff port map(x=>p(284)(112),y=>p(285)(112),Cin=>p(286)(112),clock=>clock,reset=>reset,s=>p(319)(112),cout=>p(320)(113));
FA_ff_11972:FAff port map(x=>p(284)(113),y=>p(285)(113),Cin=>p(286)(113),clock=>clock,reset=>reset,s=>p(319)(113),cout=>p(320)(114));
FA_ff_11973:FAff port map(x=>p(284)(114),y=>p(285)(114),Cin=>p(286)(114),clock=>clock,reset=>reset,s=>p(319)(114),cout=>p(320)(115));
FA_ff_11974:FAff port map(x=>p(284)(115),y=>p(285)(115),Cin=>p(286)(115),clock=>clock,reset=>reset,s=>p(319)(115),cout=>p(320)(116));
FA_ff_11975:FAff port map(x=>p(284)(116),y=>p(285)(116),Cin=>p(286)(116),clock=>clock,reset=>reset,s=>p(319)(116),cout=>p(320)(117));
FA_ff_11976:FAff port map(x=>p(284)(117),y=>p(285)(117),Cin=>p(286)(117),clock=>clock,reset=>reset,s=>p(319)(117),cout=>p(320)(118));
FA_ff_11977:FAff port map(x=>p(284)(118),y=>p(285)(118),Cin=>p(286)(118),clock=>clock,reset=>reset,s=>p(319)(118),cout=>p(320)(119));
FA_ff_11978:FAff port map(x=>p(284)(119),y=>p(285)(119),Cin=>p(286)(119),clock=>clock,reset=>reset,s=>p(319)(119),cout=>p(320)(120));
FA_ff_11979:FAff port map(x=>p(284)(120),y=>p(285)(120),Cin=>p(286)(120),clock=>clock,reset=>reset,s=>p(319)(120),cout=>p(320)(121));
FA_ff_11980:FAff port map(x=>p(284)(121),y=>p(285)(121),Cin=>p(286)(121),clock=>clock,reset=>reset,s=>p(319)(121),cout=>p(320)(122));
FA_ff_11981:FAff port map(x=>p(284)(122),y=>p(285)(122),Cin=>p(286)(122),clock=>clock,reset=>reset,s=>p(319)(122),cout=>p(320)(123));
FA_ff_11982:FAff port map(x=>p(284)(123),y=>p(285)(123),Cin=>p(286)(123),clock=>clock,reset=>reset,s=>p(319)(123),cout=>p(320)(124));
FA_ff_11983:FAff port map(x=>p(284)(124),y=>p(285)(124),Cin=>p(286)(124),clock=>clock,reset=>reset,s=>p(319)(124),cout=>p(320)(125));
FA_ff_11984:FAff port map(x=>p(284)(125),y=>p(285)(125),Cin=>p(286)(125),clock=>clock,reset=>reset,s=>p(319)(125),cout=>p(320)(126));
FA_ff_11985:FAff port map(x=>p(284)(126),y=>p(285)(126),Cin=>p(286)(126),clock=>clock,reset=>reset,s=>p(319)(126),cout=>p(320)(127));
FA_ff_11986:FAff port map(x=>p(284)(127),y=>p(285)(127),Cin=>p(286)(127),clock=>clock,reset=>reset,s=>p(319)(127),cout=>p(320)(128));
FA_ff_11987:FAff port map(x=>p(284)(128),y=>p(285)(128),Cin=>p(286)(128),clock=>clock,reset=>reset,s=>p(319)(128),cout=>p(320)(129));
FA_ff_11988:FAff port map(x=>p(284)(129),y=>p(285)(129),Cin=>p(286)(129),clock=>clock,reset=>reset,s=>p(319)(129),cout=>p(320)(130));
p(321)(0)<=p(288)(0);
HA_ff_61:HAff port map(x=>p(288)(1),y=>p(289)(1),clock=>clock,reset=>reset,s=>p(321)(1),c=>p(322)(2));
FA_ff_11989:FAff port map(x=>p(287)(2),y=>p(288)(2),Cin=>p(289)(2),clock=>clock,reset=>reset,s=>p(321)(2),cout=>p(322)(3));
FA_ff_11990:FAff port map(x=>p(287)(3),y=>p(288)(3),Cin=>p(289)(3),clock=>clock,reset=>reset,s=>p(321)(3),cout=>p(322)(4));
FA_ff_11991:FAff port map(x=>p(287)(4),y=>p(288)(4),Cin=>p(289)(4),clock=>clock,reset=>reset,s=>p(321)(4),cout=>p(322)(5));
FA_ff_11992:FAff port map(x=>p(287)(5),y=>p(288)(5),Cin=>p(289)(5),clock=>clock,reset=>reset,s=>p(321)(5),cout=>p(322)(6));
FA_ff_11993:FAff port map(x=>p(287)(6),y=>p(288)(6),Cin=>p(289)(6),clock=>clock,reset=>reset,s=>p(321)(6),cout=>p(322)(7));
FA_ff_11994:FAff port map(x=>p(287)(7),y=>p(288)(7),Cin=>p(289)(7),clock=>clock,reset=>reset,s=>p(321)(7),cout=>p(322)(8));
FA_ff_11995:FAff port map(x=>p(287)(8),y=>p(288)(8),Cin=>p(289)(8),clock=>clock,reset=>reset,s=>p(321)(8),cout=>p(322)(9));
FA_ff_11996:FAff port map(x=>p(287)(9),y=>p(288)(9),Cin=>p(289)(9),clock=>clock,reset=>reset,s=>p(321)(9),cout=>p(322)(10));
FA_ff_11997:FAff port map(x=>p(287)(10),y=>p(288)(10),Cin=>p(289)(10),clock=>clock,reset=>reset,s=>p(321)(10),cout=>p(322)(11));
FA_ff_11998:FAff port map(x=>p(287)(11),y=>p(288)(11),Cin=>p(289)(11),clock=>clock,reset=>reset,s=>p(321)(11),cout=>p(322)(12));
FA_ff_11999:FAff port map(x=>p(287)(12),y=>p(288)(12),Cin=>p(289)(12),clock=>clock,reset=>reset,s=>p(321)(12),cout=>p(322)(13));
FA_ff_12000:FAff port map(x=>p(287)(13),y=>p(288)(13),Cin=>p(289)(13),clock=>clock,reset=>reset,s=>p(321)(13),cout=>p(322)(14));
FA_ff_12001:FAff port map(x=>p(287)(14),y=>p(288)(14),Cin=>p(289)(14),clock=>clock,reset=>reset,s=>p(321)(14),cout=>p(322)(15));
FA_ff_12002:FAff port map(x=>p(287)(15),y=>p(288)(15),Cin=>p(289)(15),clock=>clock,reset=>reset,s=>p(321)(15),cout=>p(322)(16));
FA_ff_12003:FAff port map(x=>p(287)(16),y=>p(288)(16),Cin=>p(289)(16),clock=>clock,reset=>reset,s=>p(321)(16),cout=>p(322)(17));
FA_ff_12004:FAff port map(x=>p(287)(17),y=>p(288)(17),Cin=>p(289)(17),clock=>clock,reset=>reset,s=>p(321)(17),cout=>p(322)(18));
FA_ff_12005:FAff port map(x=>p(287)(18),y=>p(288)(18),Cin=>p(289)(18),clock=>clock,reset=>reset,s=>p(321)(18),cout=>p(322)(19));
FA_ff_12006:FAff port map(x=>p(287)(19),y=>p(288)(19),Cin=>p(289)(19),clock=>clock,reset=>reset,s=>p(321)(19),cout=>p(322)(20));
FA_ff_12007:FAff port map(x=>p(287)(20),y=>p(288)(20),Cin=>p(289)(20),clock=>clock,reset=>reset,s=>p(321)(20),cout=>p(322)(21));
FA_ff_12008:FAff port map(x=>p(287)(21),y=>p(288)(21),Cin=>p(289)(21),clock=>clock,reset=>reset,s=>p(321)(21),cout=>p(322)(22));
FA_ff_12009:FAff port map(x=>p(287)(22),y=>p(288)(22),Cin=>p(289)(22),clock=>clock,reset=>reset,s=>p(321)(22),cout=>p(322)(23));
FA_ff_12010:FAff port map(x=>p(287)(23),y=>p(288)(23),Cin=>p(289)(23),clock=>clock,reset=>reset,s=>p(321)(23),cout=>p(322)(24));
FA_ff_12011:FAff port map(x=>p(287)(24),y=>p(288)(24),Cin=>p(289)(24),clock=>clock,reset=>reset,s=>p(321)(24),cout=>p(322)(25));
FA_ff_12012:FAff port map(x=>p(287)(25),y=>p(288)(25),Cin=>p(289)(25),clock=>clock,reset=>reset,s=>p(321)(25),cout=>p(322)(26));
FA_ff_12013:FAff port map(x=>p(287)(26),y=>p(288)(26),Cin=>p(289)(26),clock=>clock,reset=>reset,s=>p(321)(26),cout=>p(322)(27));
FA_ff_12014:FAff port map(x=>p(287)(27),y=>p(288)(27),Cin=>p(289)(27),clock=>clock,reset=>reset,s=>p(321)(27),cout=>p(322)(28));
FA_ff_12015:FAff port map(x=>p(287)(28),y=>p(288)(28),Cin=>p(289)(28),clock=>clock,reset=>reset,s=>p(321)(28),cout=>p(322)(29));
FA_ff_12016:FAff port map(x=>p(287)(29),y=>p(288)(29),Cin=>p(289)(29),clock=>clock,reset=>reset,s=>p(321)(29),cout=>p(322)(30));
FA_ff_12017:FAff port map(x=>p(287)(30),y=>p(288)(30),Cin=>p(289)(30),clock=>clock,reset=>reset,s=>p(321)(30),cout=>p(322)(31));
FA_ff_12018:FAff port map(x=>p(287)(31),y=>p(288)(31),Cin=>p(289)(31),clock=>clock,reset=>reset,s=>p(321)(31),cout=>p(322)(32));
FA_ff_12019:FAff port map(x=>p(287)(32),y=>p(288)(32),Cin=>p(289)(32),clock=>clock,reset=>reset,s=>p(321)(32),cout=>p(322)(33));
FA_ff_12020:FAff port map(x=>p(287)(33),y=>p(288)(33),Cin=>p(289)(33),clock=>clock,reset=>reset,s=>p(321)(33),cout=>p(322)(34));
FA_ff_12021:FAff port map(x=>p(287)(34),y=>p(288)(34),Cin=>p(289)(34),clock=>clock,reset=>reset,s=>p(321)(34),cout=>p(322)(35));
FA_ff_12022:FAff port map(x=>p(287)(35),y=>p(288)(35),Cin=>p(289)(35),clock=>clock,reset=>reset,s=>p(321)(35),cout=>p(322)(36));
FA_ff_12023:FAff port map(x=>p(287)(36),y=>p(288)(36),Cin=>p(289)(36),clock=>clock,reset=>reset,s=>p(321)(36),cout=>p(322)(37));
FA_ff_12024:FAff port map(x=>p(287)(37),y=>p(288)(37),Cin=>p(289)(37),clock=>clock,reset=>reset,s=>p(321)(37),cout=>p(322)(38));
FA_ff_12025:FAff port map(x=>p(287)(38),y=>p(288)(38),Cin=>p(289)(38),clock=>clock,reset=>reset,s=>p(321)(38),cout=>p(322)(39));
FA_ff_12026:FAff port map(x=>p(287)(39),y=>p(288)(39),Cin=>p(289)(39),clock=>clock,reset=>reset,s=>p(321)(39),cout=>p(322)(40));
FA_ff_12027:FAff port map(x=>p(287)(40),y=>p(288)(40),Cin=>p(289)(40),clock=>clock,reset=>reset,s=>p(321)(40),cout=>p(322)(41));
FA_ff_12028:FAff port map(x=>p(287)(41),y=>p(288)(41),Cin=>p(289)(41),clock=>clock,reset=>reset,s=>p(321)(41),cout=>p(322)(42));
FA_ff_12029:FAff port map(x=>p(287)(42),y=>p(288)(42),Cin=>p(289)(42),clock=>clock,reset=>reset,s=>p(321)(42),cout=>p(322)(43));
FA_ff_12030:FAff port map(x=>p(287)(43),y=>p(288)(43),Cin=>p(289)(43),clock=>clock,reset=>reset,s=>p(321)(43),cout=>p(322)(44));
FA_ff_12031:FAff port map(x=>p(287)(44),y=>p(288)(44),Cin=>p(289)(44),clock=>clock,reset=>reset,s=>p(321)(44),cout=>p(322)(45));
FA_ff_12032:FAff port map(x=>p(287)(45),y=>p(288)(45),Cin=>p(289)(45),clock=>clock,reset=>reset,s=>p(321)(45),cout=>p(322)(46));
FA_ff_12033:FAff port map(x=>p(287)(46),y=>p(288)(46),Cin=>p(289)(46),clock=>clock,reset=>reset,s=>p(321)(46),cout=>p(322)(47));
FA_ff_12034:FAff port map(x=>p(287)(47),y=>p(288)(47),Cin=>p(289)(47),clock=>clock,reset=>reset,s=>p(321)(47),cout=>p(322)(48));
FA_ff_12035:FAff port map(x=>p(287)(48),y=>p(288)(48),Cin=>p(289)(48),clock=>clock,reset=>reset,s=>p(321)(48),cout=>p(322)(49));
FA_ff_12036:FAff port map(x=>p(287)(49),y=>p(288)(49),Cin=>p(289)(49),clock=>clock,reset=>reset,s=>p(321)(49),cout=>p(322)(50));
FA_ff_12037:FAff port map(x=>p(287)(50),y=>p(288)(50),Cin=>p(289)(50),clock=>clock,reset=>reset,s=>p(321)(50),cout=>p(322)(51));
FA_ff_12038:FAff port map(x=>p(287)(51),y=>p(288)(51),Cin=>p(289)(51),clock=>clock,reset=>reset,s=>p(321)(51),cout=>p(322)(52));
FA_ff_12039:FAff port map(x=>p(287)(52),y=>p(288)(52),Cin=>p(289)(52),clock=>clock,reset=>reset,s=>p(321)(52),cout=>p(322)(53));
FA_ff_12040:FAff port map(x=>p(287)(53),y=>p(288)(53),Cin=>p(289)(53),clock=>clock,reset=>reset,s=>p(321)(53),cout=>p(322)(54));
FA_ff_12041:FAff port map(x=>p(287)(54),y=>p(288)(54),Cin=>p(289)(54),clock=>clock,reset=>reset,s=>p(321)(54),cout=>p(322)(55));
FA_ff_12042:FAff port map(x=>p(287)(55),y=>p(288)(55),Cin=>p(289)(55),clock=>clock,reset=>reset,s=>p(321)(55),cout=>p(322)(56));
FA_ff_12043:FAff port map(x=>p(287)(56),y=>p(288)(56),Cin=>p(289)(56),clock=>clock,reset=>reset,s=>p(321)(56),cout=>p(322)(57));
FA_ff_12044:FAff port map(x=>p(287)(57),y=>p(288)(57),Cin=>p(289)(57),clock=>clock,reset=>reset,s=>p(321)(57),cout=>p(322)(58));
FA_ff_12045:FAff port map(x=>p(287)(58),y=>p(288)(58),Cin=>p(289)(58),clock=>clock,reset=>reset,s=>p(321)(58),cout=>p(322)(59));
FA_ff_12046:FAff port map(x=>p(287)(59),y=>p(288)(59),Cin=>p(289)(59),clock=>clock,reset=>reset,s=>p(321)(59),cout=>p(322)(60));
FA_ff_12047:FAff port map(x=>p(287)(60),y=>p(288)(60),Cin=>p(289)(60),clock=>clock,reset=>reset,s=>p(321)(60),cout=>p(322)(61));
FA_ff_12048:FAff port map(x=>p(287)(61),y=>p(288)(61),Cin=>p(289)(61),clock=>clock,reset=>reset,s=>p(321)(61),cout=>p(322)(62));
FA_ff_12049:FAff port map(x=>p(287)(62),y=>p(288)(62),Cin=>p(289)(62),clock=>clock,reset=>reset,s=>p(321)(62),cout=>p(322)(63));
FA_ff_12050:FAff port map(x=>p(287)(63),y=>p(288)(63),Cin=>p(289)(63),clock=>clock,reset=>reset,s=>p(321)(63),cout=>p(322)(64));
FA_ff_12051:FAff port map(x=>p(287)(64),y=>p(288)(64),Cin=>p(289)(64),clock=>clock,reset=>reset,s=>p(321)(64),cout=>p(322)(65));
FA_ff_12052:FAff port map(x=>p(287)(65),y=>p(288)(65),Cin=>p(289)(65),clock=>clock,reset=>reset,s=>p(321)(65),cout=>p(322)(66));
FA_ff_12053:FAff port map(x=>p(287)(66),y=>p(288)(66),Cin=>p(289)(66),clock=>clock,reset=>reset,s=>p(321)(66),cout=>p(322)(67));
FA_ff_12054:FAff port map(x=>p(287)(67),y=>p(288)(67),Cin=>p(289)(67),clock=>clock,reset=>reset,s=>p(321)(67),cout=>p(322)(68));
FA_ff_12055:FAff port map(x=>p(287)(68),y=>p(288)(68),Cin=>p(289)(68),clock=>clock,reset=>reset,s=>p(321)(68),cout=>p(322)(69));
FA_ff_12056:FAff port map(x=>p(287)(69),y=>p(288)(69),Cin=>p(289)(69),clock=>clock,reset=>reset,s=>p(321)(69),cout=>p(322)(70));
FA_ff_12057:FAff port map(x=>p(287)(70),y=>p(288)(70),Cin=>p(289)(70),clock=>clock,reset=>reset,s=>p(321)(70),cout=>p(322)(71));
FA_ff_12058:FAff port map(x=>p(287)(71),y=>p(288)(71),Cin=>p(289)(71),clock=>clock,reset=>reset,s=>p(321)(71),cout=>p(322)(72));
FA_ff_12059:FAff port map(x=>p(287)(72),y=>p(288)(72),Cin=>p(289)(72),clock=>clock,reset=>reset,s=>p(321)(72),cout=>p(322)(73));
FA_ff_12060:FAff port map(x=>p(287)(73),y=>p(288)(73),Cin=>p(289)(73),clock=>clock,reset=>reset,s=>p(321)(73),cout=>p(322)(74));
FA_ff_12061:FAff port map(x=>p(287)(74),y=>p(288)(74),Cin=>p(289)(74),clock=>clock,reset=>reset,s=>p(321)(74),cout=>p(322)(75));
FA_ff_12062:FAff port map(x=>p(287)(75),y=>p(288)(75),Cin=>p(289)(75),clock=>clock,reset=>reset,s=>p(321)(75),cout=>p(322)(76));
FA_ff_12063:FAff port map(x=>p(287)(76),y=>p(288)(76),Cin=>p(289)(76),clock=>clock,reset=>reset,s=>p(321)(76),cout=>p(322)(77));
FA_ff_12064:FAff port map(x=>p(287)(77),y=>p(288)(77),Cin=>p(289)(77),clock=>clock,reset=>reset,s=>p(321)(77),cout=>p(322)(78));
FA_ff_12065:FAff port map(x=>p(287)(78),y=>p(288)(78),Cin=>p(289)(78),clock=>clock,reset=>reset,s=>p(321)(78),cout=>p(322)(79));
FA_ff_12066:FAff port map(x=>p(287)(79),y=>p(288)(79),Cin=>p(289)(79),clock=>clock,reset=>reset,s=>p(321)(79),cout=>p(322)(80));
FA_ff_12067:FAff port map(x=>p(287)(80),y=>p(288)(80),Cin=>p(289)(80),clock=>clock,reset=>reset,s=>p(321)(80),cout=>p(322)(81));
FA_ff_12068:FAff port map(x=>p(287)(81),y=>p(288)(81),Cin=>p(289)(81),clock=>clock,reset=>reset,s=>p(321)(81),cout=>p(322)(82));
FA_ff_12069:FAff port map(x=>p(287)(82),y=>p(288)(82),Cin=>p(289)(82),clock=>clock,reset=>reset,s=>p(321)(82),cout=>p(322)(83));
FA_ff_12070:FAff port map(x=>p(287)(83),y=>p(288)(83),Cin=>p(289)(83),clock=>clock,reset=>reset,s=>p(321)(83),cout=>p(322)(84));
FA_ff_12071:FAff port map(x=>p(287)(84),y=>p(288)(84),Cin=>p(289)(84),clock=>clock,reset=>reset,s=>p(321)(84),cout=>p(322)(85));
FA_ff_12072:FAff port map(x=>p(287)(85),y=>p(288)(85),Cin=>p(289)(85),clock=>clock,reset=>reset,s=>p(321)(85),cout=>p(322)(86));
FA_ff_12073:FAff port map(x=>p(287)(86),y=>p(288)(86),Cin=>p(289)(86),clock=>clock,reset=>reset,s=>p(321)(86),cout=>p(322)(87));
FA_ff_12074:FAff port map(x=>p(287)(87),y=>p(288)(87),Cin=>p(289)(87),clock=>clock,reset=>reset,s=>p(321)(87),cout=>p(322)(88));
FA_ff_12075:FAff port map(x=>p(287)(88),y=>p(288)(88),Cin=>p(289)(88),clock=>clock,reset=>reset,s=>p(321)(88),cout=>p(322)(89));
FA_ff_12076:FAff port map(x=>p(287)(89),y=>p(288)(89),Cin=>p(289)(89),clock=>clock,reset=>reset,s=>p(321)(89),cout=>p(322)(90));
FA_ff_12077:FAff port map(x=>p(287)(90),y=>p(288)(90),Cin=>p(289)(90),clock=>clock,reset=>reset,s=>p(321)(90),cout=>p(322)(91));
FA_ff_12078:FAff port map(x=>p(287)(91),y=>p(288)(91),Cin=>p(289)(91),clock=>clock,reset=>reset,s=>p(321)(91),cout=>p(322)(92));
FA_ff_12079:FAff port map(x=>p(287)(92),y=>p(288)(92),Cin=>p(289)(92),clock=>clock,reset=>reset,s=>p(321)(92),cout=>p(322)(93));
FA_ff_12080:FAff port map(x=>p(287)(93),y=>p(288)(93),Cin=>p(289)(93),clock=>clock,reset=>reset,s=>p(321)(93),cout=>p(322)(94));
FA_ff_12081:FAff port map(x=>p(287)(94),y=>p(288)(94),Cin=>p(289)(94),clock=>clock,reset=>reset,s=>p(321)(94),cout=>p(322)(95));
FA_ff_12082:FAff port map(x=>p(287)(95),y=>p(288)(95),Cin=>p(289)(95),clock=>clock,reset=>reset,s=>p(321)(95),cout=>p(322)(96));
FA_ff_12083:FAff port map(x=>p(287)(96),y=>p(288)(96),Cin=>p(289)(96),clock=>clock,reset=>reset,s=>p(321)(96),cout=>p(322)(97));
FA_ff_12084:FAff port map(x=>p(287)(97),y=>p(288)(97),Cin=>p(289)(97),clock=>clock,reset=>reset,s=>p(321)(97),cout=>p(322)(98));
FA_ff_12085:FAff port map(x=>p(287)(98),y=>p(288)(98),Cin=>p(289)(98),clock=>clock,reset=>reset,s=>p(321)(98),cout=>p(322)(99));
FA_ff_12086:FAff port map(x=>p(287)(99),y=>p(288)(99),Cin=>p(289)(99),clock=>clock,reset=>reset,s=>p(321)(99),cout=>p(322)(100));
FA_ff_12087:FAff port map(x=>p(287)(100),y=>p(288)(100),Cin=>p(289)(100),clock=>clock,reset=>reset,s=>p(321)(100),cout=>p(322)(101));
FA_ff_12088:FAff port map(x=>p(287)(101),y=>p(288)(101),Cin=>p(289)(101),clock=>clock,reset=>reset,s=>p(321)(101),cout=>p(322)(102));
FA_ff_12089:FAff port map(x=>p(287)(102),y=>p(288)(102),Cin=>p(289)(102),clock=>clock,reset=>reset,s=>p(321)(102),cout=>p(322)(103));
FA_ff_12090:FAff port map(x=>p(287)(103),y=>p(288)(103),Cin=>p(289)(103),clock=>clock,reset=>reset,s=>p(321)(103),cout=>p(322)(104));
FA_ff_12091:FAff port map(x=>p(287)(104),y=>p(288)(104),Cin=>p(289)(104),clock=>clock,reset=>reset,s=>p(321)(104),cout=>p(322)(105));
FA_ff_12092:FAff port map(x=>p(287)(105),y=>p(288)(105),Cin=>p(289)(105),clock=>clock,reset=>reset,s=>p(321)(105),cout=>p(322)(106));
FA_ff_12093:FAff port map(x=>p(287)(106),y=>p(288)(106),Cin=>p(289)(106),clock=>clock,reset=>reset,s=>p(321)(106),cout=>p(322)(107));
FA_ff_12094:FAff port map(x=>p(287)(107),y=>p(288)(107),Cin=>p(289)(107),clock=>clock,reset=>reset,s=>p(321)(107),cout=>p(322)(108));
FA_ff_12095:FAff port map(x=>p(287)(108),y=>p(288)(108),Cin=>p(289)(108),clock=>clock,reset=>reset,s=>p(321)(108),cout=>p(322)(109));
FA_ff_12096:FAff port map(x=>p(287)(109),y=>p(288)(109),Cin=>p(289)(109),clock=>clock,reset=>reset,s=>p(321)(109),cout=>p(322)(110));
FA_ff_12097:FAff port map(x=>p(287)(110),y=>p(288)(110),Cin=>p(289)(110),clock=>clock,reset=>reset,s=>p(321)(110),cout=>p(322)(111));
FA_ff_12098:FAff port map(x=>p(287)(111),y=>p(288)(111),Cin=>p(289)(111),clock=>clock,reset=>reset,s=>p(321)(111),cout=>p(322)(112));
FA_ff_12099:FAff port map(x=>p(287)(112),y=>p(288)(112),Cin=>p(289)(112),clock=>clock,reset=>reset,s=>p(321)(112),cout=>p(322)(113));
FA_ff_12100:FAff port map(x=>p(287)(113),y=>p(288)(113),Cin=>p(289)(113),clock=>clock,reset=>reset,s=>p(321)(113),cout=>p(322)(114));
FA_ff_12101:FAff port map(x=>p(287)(114),y=>p(288)(114),Cin=>p(289)(114),clock=>clock,reset=>reset,s=>p(321)(114),cout=>p(322)(115));
FA_ff_12102:FAff port map(x=>p(287)(115),y=>p(288)(115),Cin=>p(289)(115),clock=>clock,reset=>reset,s=>p(321)(115),cout=>p(322)(116));
FA_ff_12103:FAff port map(x=>p(287)(116),y=>p(288)(116),Cin=>p(289)(116),clock=>clock,reset=>reset,s=>p(321)(116),cout=>p(322)(117));
FA_ff_12104:FAff port map(x=>p(287)(117),y=>p(288)(117),Cin=>p(289)(117),clock=>clock,reset=>reset,s=>p(321)(117),cout=>p(322)(118));
FA_ff_12105:FAff port map(x=>p(287)(118),y=>p(288)(118),Cin=>p(289)(118),clock=>clock,reset=>reset,s=>p(321)(118),cout=>p(322)(119));
FA_ff_12106:FAff port map(x=>p(287)(119),y=>p(288)(119),Cin=>p(289)(119),clock=>clock,reset=>reset,s=>p(321)(119),cout=>p(322)(120));
FA_ff_12107:FAff port map(x=>p(287)(120),y=>p(288)(120),Cin=>p(289)(120),clock=>clock,reset=>reset,s=>p(321)(120),cout=>p(322)(121));
FA_ff_12108:FAff port map(x=>p(287)(121),y=>p(288)(121),Cin=>p(289)(121),clock=>clock,reset=>reset,s=>p(321)(121),cout=>p(322)(122));
FA_ff_12109:FAff port map(x=>p(287)(122),y=>p(288)(122),Cin=>p(289)(122),clock=>clock,reset=>reset,s=>p(321)(122),cout=>p(322)(123));
FA_ff_12110:FAff port map(x=>p(287)(123),y=>p(288)(123),Cin=>p(289)(123),clock=>clock,reset=>reset,s=>p(321)(123),cout=>p(322)(124));
FA_ff_12111:FAff port map(x=>p(287)(124),y=>p(288)(124),Cin=>p(289)(124),clock=>clock,reset=>reset,s=>p(321)(124),cout=>p(322)(125));
FA_ff_12112:FAff port map(x=>p(287)(125),y=>p(288)(125),Cin=>p(289)(125),clock=>clock,reset=>reset,s=>p(321)(125),cout=>p(322)(126));
FA_ff_12113:FAff port map(x=>p(287)(126),y=>p(288)(126),Cin=>p(289)(126),clock=>clock,reset=>reset,s=>p(321)(126),cout=>p(322)(127));
FA_ff_12114:FAff port map(x=>p(287)(127),y=>p(288)(127),Cin=>p(289)(127),clock=>clock,reset=>reset,s=>p(321)(127),cout=>p(322)(128));
FA_ff_12115:FAff port map(x=>p(287)(128),y=>p(288)(128),Cin=>p(289)(128),clock=>clock,reset=>reset,s=>p(321)(128),cout=>p(322)(129));
HA_ff_62:HAff port map(x=>p(287)(129),y=>p(289)(129),clock=>clock,reset=>reset,s=>p(321)(129),c=>p(322)(130));
HA_ff_63:HAff port map(x=>p(290)(0),y=>p(292)(0),clock=>clock,reset=>reset,s=>p(323)(0),c=>p(324)(1));
HA_ff_64:HAff port map(x=>p(290)(1),y=>p(292)(1),clock=>clock,reset=>reset,s=>p(323)(1),c=>p(324)(2));
FA_ff_12116:FAff port map(x=>p(290)(2),y=>p(291)(2),Cin=>p(292)(2),clock=>clock,reset=>reset,s=>p(323)(2),cout=>p(324)(3));
FA_ff_12117:FAff port map(x=>p(290)(3),y=>p(291)(3),Cin=>p(292)(3),clock=>clock,reset=>reset,s=>p(323)(3),cout=>p(324)(4));
FA_ff_12118:FAff port map(x=>p(290)(4),y=>p(291)(4),Cin=>p(292)(4),clock=>clock,reset=>reset,s=>p(323)(4),cout=>p(324)(5));
FA_ff_12119:FAff port map(x=>p(290)(5),y=>p(291)(5),Cin=>p(292)(5),clock=>clock,reset=>reset,s=>p(323)(5),cout=>p(324)(6));
FA_ff_12120:FAff port map(x=>p(290)(6),y=>p(291)(6),Cin=>p(292)(6),clock=>clock,reset=>reset,s=>p(323)(6),cout=>p(324)(7));
FA_ff_12121:FAff port map(x=>p(290)(7),y=>p(291)(7),Cin=>p(292)(7),clock=>clock,reset=>reset,s=>p(323)(7),cout=>p(324)(8));
FA_ff_12122:FAff port map(x=>p(290)(8),y=>p(291)(8),Cin=>p(292)(8),clock=>clock,reset=>reset,s=>p(323)(8),cout=>p(324)(9));
FA_ff_12123:FAff port map(x=>p(290)(9),y=>p(291)(9),Cin=>p(292)(9),clock=>clock,reset=>reset,s=>p(323)(9),cout=>p(324)(10));
FA_ff_12124:FAff port map(x=>p(290)(10),y=>p(291)(10),Cin=>p(292)(10),clock=>clock,reset=>reset,s=>p(323)(10),cout=>p(324)(11));
FA_ff_12125:FAff port map(x=>p(290)(11),y=>p(291)(11),Cin=>p(292)(11),clock=>clock,reset=>reset,s=>p(323)(11),cout=>p(324)(12));
FA_ff_12126:FAff port map(x=>p(290)(12),y=>p(291)(12),Cin=>p(292)(12),clock=>clock,reset=>reset,s=>p(323)(12),cout=>p(324)(13));
FA_ff_12127:FAff port map(x=>p(290)(13),y=>p(291)(13),Cin=>p(292)(13),clock=>clock,reset=>reset,s=>p(323)(13),cout=>p(324)(14));
FA_ff_12128:FAff port map(x=>p(290)(14),y=>p(291)(14),Cin=>p(292)(14),clock=>clock,reset=>reset,s=>p(323)(14),cout=>p(324)(15));
FA_ff_12129:FAff port map(x=>p(290)(15),y=>p(291)(15),Cin=>p(292)(15),clock=>clock,reset=>reset,s=>p(323)(15),cout=>p(324)(16));
FA_ff_12130:FAff port map(x=>p(290)(16),y=>p(291)(16),Cin=>p(292)(16),clock=>clock,reset=>reset,s=>p(323)(16),cout=>p(324)(17));
FA_ff_12131:FAff port map(x=>p(290)(17),y=>p(291)(17),Cin=>p(292)(17),clock=>clock,reset=>reset,s=>p(323)(17),cout=>p(324)(18));
FA_ff_12132:FAff port map(x=>p(290)(18),y=>p(291)(18),Cin=>p(292)(18),clock=>clock,reset=>reset,s=>p(323)(18),cout=>p(324)(19));
FA_ff_12133:FAff port map(x=>p(290)(19),y=>p(291)(19),Cin=>p(292)(19),clock=>clock,reset=>reset,s=>p(323)(19),cout=>p(324)(20));
FA_ff_12134:FAff port map(x=>p(290)(20),y=>p(291)(20),Cin=>p(292)(20),clock=>clock,reset=>reset,s=>p(323)(20),cout=>p(324)(21));
FA_ff_12135:FAff port map(x=>p(290)(21),y=>p(291)(21),Cin=>p(292)(21),clock=>clock,reset=>reset,s=>p(323)(21),cout=>p(324)(22));
FA_ff_12136:FAff port map(x=>p(290)(22),y=>p(291)(22),Cin=>p(292)(22),clock=>clock,reset=>reset,s=>p(323)(22),cout=>p(324)(23));
FA_ff_12137:FAff port map(x=>p(290)(23),y=>p(291)(23),Cin=>p(292)(23),clock=>clock,reset=>reset,s=>p(323)(23),cout=>p(324)(24));
FA_ff_12138:FAff port map(x=>p(290)(24),y=>p(291)(24),Cin=>p(292)(24),clock=>clock,reset=>reset,s=>p(323)(24),cout=>p(324)(25));
FA_ff_12139:FAff port map(x=>p(290)(25),y=>p(291)(25),Cin=>p(292)(25),clock=>clock,reset=>reset,s=>p(323)(25),cout=>p(324)(26));
FA_ff_12140:FAff port map(x=>p(290)(26),y=>p(291)(26),Cin=>p(292)(26),clock=>clock,reset=>reset,s=>p(323)(26),cout=>p(324)(27));
FA_ff_12141:FAff port map(x=>p(290)(27),y=>p(291)(27),Cin=>p(292)(27),clock=>clock,reset=>reset,s=>p(323)(27),cout=>p(324)(28));
FA_ff_12142:FAff port map(x=>p(290)(28),y=>p(291)(28),Cin=>p(292)(28),clock=>clock,reset=>reset,s=>p(323)(28),cout=>p(324)(29));
FA_ff_12143:FAff port map(x=>p(290)(29),y=>p(291)(29),Cin=>p(292)(29),clock=>clock,reset=>reset,s=>p(323)(29),cout=>p(324)(30));
FA_ff_12144:FAff port map(x=>p(290)(30),y=>p(291)(30),Cin=>p(292)(30),clock=>clock,reset=>reset,s=>p(323)(30),cout=>p(324)(31));
FA_ff_12145:FAff port map(x=>p(290)(31),y=>p(291)(31),Cin=>p(292)(31),clock=>clock,reset=>reset,s=>p(323)(31),cout=>p(324)(32));
FA_ff_12146:FAff port map(x=>p(290)(32),y=>p(291)(32),Cin=>p(292)(32),clock=>clock,reset=>reset,s=>p(323)(32),cout=>p(324)(33));
FA_ff_12147:FAff port map(x=>p(290)(33),y=>p(291)(33),Cin=>p(292)(33),clock=>clock,reset=>reset,s=>p(323)(33),cout=>p(324)(34));
FA_ff_12148:FAff port map(x=>p(290)(34),y=>p(291)(34),Cin=>p(292)(34),clock=>clock,reset=>reset,s=>p(323)(34),cout=>p(324)(35));
FA_ff_12149:FAff port map(x=>p(290)(35),y=>p(291)(35),Cin=>p(292)(35),clock=>clock,reset=>reset,s=>p(323)(35),cout=>p(324)(36));
FA_ff_12150:FAff port map(x=>p(290)(36),y=>p(291)(36),Cin=>p(292)(36),clock=>clock,reset=>reset,s=>p(323)(36),cout=>p(324)(37));
FA_ff_12151:FAff port map(x=>p(290)(37),y=>p(291)(37),Cin=>p(292)(37),clock=>clock,reset=>reset,s=>p(323)(37),cout=>p(324)(38));
FA_ff_12152:FAff port map(x=>p(290)(38),y=>p(291)(38),Cin=>p(292)(38),clock=>clock,reset=>reset,s=>p(323)(38),cout=>p(324)(39));
FA_ff_12153:FAff port map(x=>p(290)(39),y=>p(291)(39),Cin=>p(292)(39),clock=>clock,reset=>reset,s=>p(323)(39),cout=>p(324)(40));
FA_ff_12154:FAff port map(x=>p(290)(40),y=>p(291)(40),Cin=>p(292)(40),clock=>clock,reset=>reset,s=>p(323)(40),cout=>p(324)(41));
FA_ff_12155:FAff port map(x=>p(290)(41),y=>p(291)(41),Cin=>p(292)(41),clock=>clock,reset=>reset,s=>p(323)(41),cout=>p(324)(42));
FA_ff_12156:FAff port map(x=>p(290)(42),y=>p(291)(42),Cin=>p(292)(42),clock=>clock,reset=>reset,s=>p(323)(42),cout=>p(324)(43));
FA_ff_12157:FAff port map(x=>p(290)(43),y=>p(291)(43),Cin=>p(292)(43),clock=>clock,reset=>reset,s=>p(323)(43),cout=>p(324)(44));
FA_ff_12158:FAff port map(x=>p(290)(44),y=>p(291)(44),Cin=>p(292)(44),clock=>clock,reset=>reset,s=>p(323)(44),cout=>p(324)(45));
FA_ff_12159:FAff port map(x=>p(290)(45),y=>p(291)(45),Cin=>p(292)(45),clock=>clock,reset=>reset,s=>p(323)(45),cout=>p(324)(46));
FA_ff_12160:FAff port map(x=>p(290)(46),y=>p(291)(46),Cin=>p(292)(46),clock=>clock,reset=>reset,s=>p(323)(46),cout=>p(324)(47));
FA_ff_12161:FAff port map(x=>p(290)(47),y=>p(291)(47),Cin=>p(292)(47),clock=>clock,reset=>reset,s=>p(323)(47),cout=>p(324)(48));
FA_ff_12162:FAff port map(x=>p(290)(48),y=>p(291)(48),Cin=>p(292)(48),clock=>clock,reset=>reset,s=>p(323)(48),cout=>p(324)(49));
FA_ff_12163:FAff port map(x=>p(290)(49),y=>p(291)(49),Cin=>p(292)(49),clock=>clock,reset=>reset,s=>p(323)(49),cout=>p(324)(50));
FA_ff_12164:FAff port map(x=>p(290)(50),y=>p(291)(50),Cin=>p(292)(50),clock=>clock,reset=>reset,s=>p(323)(50),cout=>p(324)(51));
FA_ff_12165:FAff port map(x=>p(290)(51),y=>p(291)(51),Cin=>p(292)(51),clock=>clock,reset=>reset,s=>p(323)(51),cout=>p(324)(52));
FA_ff_12166:FAff port map(x=>p(290)(52),y=>p(291)(52),Cin=>p(292)(52),clock=>clock,reset=>reset,s=>p(323)(52),cout=>p(324)(53));
FA_ff_12167:FAff port map(x=>p(290)(53),y=>p(291)(53),Cin=>p(292)(53),clock=>clock,reset=>reset,s=>p(323)(53),cout=>p(324)(54));
FA_ff_12168:FAff port map(x=>p(290)(54),y=>p(291)(54),Cin=>p(292)(54),clock=>clock,reset=>reset,s=>p(323)(54),cout=>p(324)(55));
FA_ff_12169:FAff port map(x=>p(290)(55),y=>p(291)(55),Cin=>p(292)(55),clock=>clock,reset=>reset,s=>p(323)(55),cout=>p(324)(56));
FA_ff_12170:FAff port map(x=>p(290)(56),y=>p(291)(56),Cin=>p(292)(56),clock=>clock,reset=>reset,s=>p(323)(56),cout=>p(324)(57));
FA_ff_12171:FAff port map(x=>p(290)(57),y=>p(291)(57),Cin=>p(292)(57),clock=>clock,reset=>reset,s=>p(323)(57),cout=>p(324)(58));
FA_ff_12172:FAff port map(x=>p(290)(58),y=>p(291)(58),Cin=>p(292)(58),clock=>clock,reset=>reset,s=>p(323)(58),cout=>p(324)(59));
FA_ff_12173:FAff port map(x=>p(290)(59),y=>p(291)(59),Cin=>p(292)(59),clock=>clock,reset=>reset,s=>p(323)(59),cout=>p(324)(60));
FA_ff_12174:FAff port map(x=>p(290)(60),y=>p(291)(60),Cin=>p(292)(60),clock=>clock,reset=>reset,s=>p(323)(60),cout=>p(324)(61));
FA_ff_12175:FAff port map(x=>p(290)(61),y=>p(291)(61),Cin=>p(292)(61),clock=>clock,reset=>reset,s=>p(323)(61),cout=>p(324)(62));
FA_ff_12176:FAff port map(x=>p(290)(62),y=>p(291)(62),Cin=>p(292)(62),clock=>clock,reset=>reset,s=>p(323)(62),cout=>p(324)(63));
FA_ff_12177:FAff port map(x=>p(290)(63),y=>p(291)(63),Cin=>p(292)(63),clock=>clock,reset=>reset,s=>p(323)(63),cout=>p(324)(64));
FA_ff_12178:FAff port map(x=>p(290)(64),y=>p(291)(64),Cin=>p(292)(64),clock=>clock,reset=>reset,s=>p(323)(64),cout=>p(324)(65));
FA_ff_12179:FAff port map(x=>p(290)(65),y=>p(291)(65),Cin=>p(292)(65),clock=>clock,reset=>reset,s=>p(323)(65),cout=>p(324)(66));
FA_ff_12180:FAff port map(x=>p(290)(66),y=>p(291)(66),Cin=>p(292)(66),clock=>clock,reset=>reset,s=>p(323)(66),cout=>p(324)(67));
FA_ff_12181:FAff port map(x=>p(290)(67),y=>p(291)(67),Cin=>p(292)(67),clock=>clock,reset=>reset,s=>p(323)(67),cout=>p(324)(68));
FA_ff_12182:FAff port map(x=>p(290)(68),y=>p(291)(68),Cin=>p(292)(68),clock=>clock,reset=>reset,s=>p(323)(68),cout=>p(324)(69));
FA_ff_12183:FAff port map(x=>p(290)(69),y=>p(291)(69),Cin=>p(292)(69),clock=>clock,reset=>reset,s=>p(323)(69),cout=>p(324)(70));
FA_ff_12184:FAff port map(x=>p(290)(70),y=>p(291)(70),Cin=>p(292)(70),clock=>clock,reset=>reset,s=>p(323)(70),cout=>p(324)(71));
FA_ff_12185:FAff port map(x=>p(290)(71),y=>p(291)(71),Cin=>p(292)(71),clock=>clock,reset=>reset,s=>p(323)(71),cout=>p(324)(72));
FA_ff_12186:FAff port map(x=>p(290)(72),y=>p(291)(72),Cin=>p(292)(72),clock=>clock,reset=>reset,s=>p(323)(72),cout=>p(324)(73));
FA_ff_12187:FAff port map(x=>p(290)(73),y=>p(291)(73),Cin=>p(292)(73),clock=>clock,reset=>reset,s=>p(323)(73),cout=>p(324)(74));
FA_ff_12188:FAff port map(x=>p(290)(74),y=>p(291)(74),Cin=>p(292)(74),clock=>clock,reset=>reset,s=>p(323)(74),cout=>p(324)(75));
FA_ff_12189:FAff port map(x=>p(290)(75),y=>p(291)(75),Cin=>p(292)(75),clock=>clock,reset=>reset,s=>p(323)(75),cout=>p(324)(76));
FA_ff_12190:FAff port map(x=>p(290)(76),y=>p(291)(76),Cin=>p(292)(76),clock=>clock,reset=>reset,s=>p(323)(76),cout=>p(324)(77));
FA_ff_12191:FAff port map(x=>p(290)(77),y=>p(291)(77),Cin=>p(292)(77),clock=>clock,reset=>reset,s=>p(323)(77),cout=>p(324)(78));
FA_ff_12192:FAff port map(x=>p(290)(78),y=>p(291)(78),Cin=>p(292)(78),clock=>clock,reset=>reset,s=>p(323)(78),cout=>p(324)(79));
FA_ff_12193:FAff port map(x=>p(290)(79),y=>p(291)(79),Cin=>p(292)(79),clock=>clock,reset=>reset,s=>p(323)(79),cout=>p(324)(80));
FA_ff_12194:FAff port map(x=>p(290)(80),y=>p(291)(80),Cin=>p(292)(80),clock=>clock,reset=>reset,s=>p(323)(80),cout=>p(324)(81));
FA_ff_12195:FAff port map(x=>p(290)(81),y=>p(291)(81),Cin=>p(292)(81),clock=>clock,reset=>reset,s=>p(323)(81),cout=>p(324)(82));
FA_ff_12196:FAff port map(x=>p(290)(82),y=>p(291)(82),Cin=>p(292)(82),clock=>clock,reset=>reset,s=>p(323)(82),cout=>p(324)(83));
FA_ff_12197:FAff port map(x=>p(290)(83),y=>p(291)(83),Cin=>p(292)(83),clock=>clock,reset=>reset,s=>p(323)(83),cout=>p(324)(84));
FA_ff_12198:FAff port map(x=>p(290)(84),y=>p(291)(84),Cin=>p(292)(84),clock=>clock,reset=>reset,s=>p(323)(84),cout=>p(324)(85));
FA_ff_12199:FAff port map(x=>p(290)(85),y=>p(291)(85),Cin=>p(292)(85),clock=>clock,reset=>reset,s=>p(323)(85),cout=>p(324)(86));
FA_ff_12200:FAff port map(x=>p(290)(86),y=>p(291)(86),Cin=>p(292)(86),clock=>clock,reset=>reset,s=>p(323)(86),cout=>p(324)(87));
FA_ff_12201:FAff port map(x=>p(290)(87),y=>p(291)(87),Cin=>p(292)(87),clock=>clock,reset=>reset,s=>p(323)(87),cout=>p(324)(88));
FA_ff_12202:FAff port map(x=>p(290)(88),y=>p(291)(88),Cin=>p(292)(88),clock=>clock,reset=>reset,s=>p(323)(88),cout=>p(324)(89));
FA_ff_12203:FAff port map(x=>p(290)(89),y=>p(291)(89),Cin=>p(292)(89),clock=>clock,reset=>reset,s=>p(323)(89),cout=>p(324)(90));
FA_ff_12204:FAff port map(x=>p(290)(90),y=>p(291)(90),Cin=>p(292)(90),clock=>clock,reset=>reset,s=>p(323)(90),cout=>p(324)(91));
FA_ff_12205:FAff port map(x=>p(290)(91),y=>p(291)(91),Cin=>p(292)(91),clock=>clock,reset=>reset,s=>p(323)(91),cout=>p(324)(92));
FA_ff_12206:FAff port map(x=>p(290)(92),y=>p(291)(92),Cin=>p(292)(92),clock=>clock,reset=>reset,s=>p(323)(92),cout=>p(324)(93));
FA_ff_12207:FAff port map(x=>p(290)(93),y=>p(291)(93),Cin=>p(292)(93),clock=>clock,reset=>reset,s=>p(323)(93),cout=>p(324)(94));
FA_ff_12208:FAff port map(x=>p(290)(94),y=>p(291)(94),Cin=>p(292)(94),clock=>clock,reset=>reset,s=>p(323)(94),cout=>p(324)(95));
FA_ff_12209:FAff port map(x=>p(290)(95),y=>p(291)(95),Cin=>p(292)(95),clock=>clock,reset=>reset,s=>p(323)(95),cout=>p(324)(96));
FA_ff_12210:FAff port map(x=>p(290)(96),y=>p(291)(96),Cin=>p(292)(96),clock=>clock,reset=>reset,s=>p(323)(96),cout=>p(324)(97));
FA_ff_12211:FAff port map(x=>p(290)(97),y=>p(291)(97),Cin=>p(292)(97),clock=>clock,reset=>reset,s=>p(323)(97),cout=>p(324)(98));
FA_ff_12212:FAff port map(x=>p(290)(98),y=>p(291)(98),Cin=>p(292)(98),clock=>clock,reset=>reset,s=>p(323)(98),cout=>p(324)(99));
FA_ff_12213:FAff port map(x=>p(290)(99),y=>p(291)(99),Cin=>p(292)(99),clock=>clock,reset=>reset,s=>p(323)(99),cout=>p(324)(100));
FA_ff_12214:FAff port map(x=>p(290)(100),y=>p(291)(100),Cin=>p(292)(100),clock=>clock,reset=>reset,s=>p(323)(100),cout=>p(324)(101));
FA_ff_12215:FAff port map(x=>p(290)(101),y=>p(291)(101),Cin=>p(292)(101),clock=>clock,reset=>reset,s=>p(323)(101),cout=>p(324)(102));
FA_ff_12216:FAff port map(x=>p(290)(102),y=>p(291)(102),Cin=>p(292)(102),clock=>clock,reset=>reset,s=>p(323)(102),cout=>p(324)(103));
FA_ff_12217:FAff port map(x=>p(290)(103),y=>p(291)(103),Cin=>p(292)(103),clock=>clock,reset=>reset,s=>p(323)(103),cout=>p(324)(104));
FA_ff_12218:FAff port map(x=>p(290)(104),y=>p(291)(104),Cin=>p(292)(104),clock=>clock,reset=>reset,s=>p(323)(104),cout=>p(324)(105));
FA_ff_12219:FAff port map(x=>p(290)(105),y=>p(291)(105),Cin=>p(292)(105),clock=>clock,reset=>reset,s=>p(323)(105),cout=>p(324)(106));
FA_ff_12220:FAff port map(x=>p(290)(106),y=>p(291)(106),Cin=>p(292)(106),clock=>clock,reset=>reset,s=>p(323)(106),cout=>p(324)(107));
FA_ff_12221:FAff port map(x=>p(290)(107),y=>p(291)(107),Cin=>p(292)(107),clock=>clock,reset=>reset,s=>p(323)(107),cout=>p(324)(108));
FA_ff_12222:FAff port map(x=>p(290)(108),y=>p(291)(108),Cin=>p(292)(108),clock=>clock,reset=>reset,s=>p(323)(108),cout=>p(324)(109));
FA_ff_12223:FAff port map(x=>p(290)(109),y=>p(291)(109),Cin=>p(292)(109),clock=>clock,reset=>reset,s=>p(323)(109),cout=>p(324)(110));
FA_ff_12224:FAff port map(x=>p(290)(110),y=>p(291)(110),Cin=>p(292)(110),clock=>clock,reset=>reset,s=>p(323)(110),cout=>p(324)(111));
FA_ff_12225:FAff port map(x=>p(290)(111),y=>p(291)(111),Cin=>p(292)(111),clock=>clock,reset=>reset,s=>p(323)(111),cout=>p(324)(112));
FA_ff_12226:FAff port map(x=>p(290)(112),y=>p(291)(112),Cin=>p(292)(112),clock=>clock,reset=>reset,s=>p(323)(112),cout=>p(324)(113));
FA_ff_12227:FAff port map(x=>p(290)(113),y=>p(291)(113),Cin=>p(292)(113),clock=>clock,reset=>reset,s=>p(323)(113),cout=>p(324)(114));
FA_ff_12228:FAff port map(x=>p(290)(114),y=>p(291)(114),Cin=>p(292)(114),clock=>clock,reset=>reset,s=>p(323)(114),cout=>p(324)(115));
FA_ff_12229:FAff port map(x=>p(290)(115),y=>p(291)(115),Cin=>p(292)(115),clock=>clock,reset=>reset,s=>p(323)(115),cout=>p(324)(116));
FA_ff_12230:FAff port map(x=>p(290)(116),y=>p(291)(116),Cin=>p(292)(116),clock=>clock,reset=>reset,s=>p(323)(116),cout=>p(324)(117));
FA_ff_12231:FAff port map(x=>p(290)(117),y=>p(291)(117),Cin=>p(292)(117),clock=>clock,reset=>reset,s=>p(323)(117),cout=>p(324)(118));
FA_ff_12232:FAff port map(x=>p(290)(118),y=>p(291)(118),Cin=>p(292)(118),clock=>clock,reset=>reset,s=>p(323)(118),cout=>p(324)(119));
FA_ff_12233:FAff port map(x=>p(290)(119),y=>p(291)(119),Cin=>p(292)(119),clock=>clock,reset=>reset,s=>p(323)(119),cout=>p(324)(120));
FA_ff_12234:FAff port map(x=>p(290)(120),y=>p(291)(120),Cin=>p(292)(120),clock=>clock,reset=>reset,s=>p(323)(120),cout=>p(324)(121));
FA_ff_12235:FAff port map(x=>p(290)(121),y=>p(291)(121),Cin=>p(292)(121),clock=>clock,reset=>reset,s=>p(323)(121),cout=>p(324)(122));
FA_ff_12236:FAff port map(x=>p(290)(122),y=>p(291)(122),Cin=>p(292)(122),clock=>clock,reset=>reset,s=>p(323)(122),cout=>p(324)(123));
FA_ff_12237:FAff port map(x=>p(290)(123),y=>p(291)(123),Cin=>p(292)(123),clock=>clock,reset=>reset,s=>p(323)(123),cout=>p(324)(124));
FA_ff_12238:FAff port map(x=>p(290)(124),y=>p(291)(124),Cin=>p(292)(124),clock=>clock,reset=>reset,s=>p(323)(124),cout=>p(324)(125));
FA_ff_12239:FAff port map(x=>p(290)(125),y=>p(291)(125),Cin=>p(292)(125),clock=>clock,reset=>reset,s=>p(323)(125),cout=>p(324)(126));
FA_ff_12240:FAff port map(x=>p(290)(126),y=>p(291)(126),Cin=>p(292)(126),clock=>clock,reset=>reset,s=>p(323)(126),cout=>p(324)(127));
FA_ff_12241:FAff port map(x=>p(290)(127),y=>p(291)(127),Cin=>p(292)(127),clock=>clock,reset=>reset,s=>p(323)(127),cout=>p(324)(128));
FA_ff_12242:FAff port map(x=>p(290)(128),y=>p(291)(128),Cin=>p(292)(128),clock=>clock,reset=>reset,s=>p(323)(128),cout=>p(324)(129));
FA_ff_12243:FAff port map(x=>p(290)(129),y=>p(291)(129),Cin=>p(292)(129),clock=>clock,reset=>reset,s=>p(323)(129),cout=>p(324)(130));
p(325)(0)<=p(294)(0);
HA_ff_65:HAff port map(x=>p(293)(1),y=>p(294)(1),clock=>clock,reset=>reset,s=>p(325)(1),c=>p(326)(2));
FA_ff_12244:FAff port map(x=>p(293)(2),y=>p(294)(2),Cin=>p(295)(2),clock=>clock,reset=>reset,s=>p(325)(2),cout=>p(326)(3));
FA_ff_12245:FAff port map(x=>p(293)(3),y=>p(294)(3),Cin=>p(295)(3),clock=>clock,reset=>reset,s=>p(325)(3),cout=>p(326)(4));
FA_ff_12246:FAff port map(x=>p(293)(4),y=>p(294)(4),Cin=>p(295)(4),clock=>clock,reset=>reset,s=>p(325)(4),cout=>p(326)(5));
FA_ff_12247:FAff port map(x=>p(293)(5),y=>p(294)(5),Cin=>p(295)(5),clock=>clock,reset=>reset,s=>p(325)(5),cout=>p(326)(6));
FA_ff_12248:FAff port map(x=>p(293)(6),y=>p(294)(6),Cin=>p(295)(6),clock=>clock,reset=>reset,s=>p(325)(6),cout=>p(326)(7));
FA_ff_12249:FAff port map(x=>p(293)(7),y=>p(294)(7),Cin=>p(295)(7),clock=>clock,reset=>reset,s=>p(325)(7),cout=>p(326)(8));
FA_ff_12250:FAff port map(x=>p(293)(8),y=>p(294)(8),Cin=>p(295)(8),clock=>clock,reset=>reset,s=>p(325)(8),cout=>p(326)(9));
FA_ff_12251:FAff port map(x=>p(293)(9),y=>p(294)(9),Cin=>p(295)(9),clock=>clock,reset=>reset,s=>p(325)(9),cout=>p(326)(10));
FA_ff_12252:FAff port map(x=>p(293)(10),y=>p(294)(10),Cin=>p(295)(10),clock=>clock,reset=>reset,s=>p(325)(10),cout=>p(326)(11));
FA_ff_12253:FAff port map(x=>p(293)(11),y=>p(294)(11),Cin=>p(295)(11),clock=>clock,reset=>reset,s=>p(325)(11),cout=>p(326)(12));
FA_ff_12254:FAff port map(x=>p(293)(12),y=>p(294)(12),Cin=>p(295)(12),clock=>clock,reset=>reset,s=>p(325)(12),cout=>p(326)(13));
FA_ff_12255:FAff port map(x=>p(293)(13),y=>p(294)(13),Cin=>p(295)(13),clock=>clock,reset=>reset,s=>p(325)(13),cout=>p(326)(14));
FA_ff_12256:FAff port map(x=>p(293)(14),y=>p(294)(14),Cin=>p(295)(14),clock=>clock,reset=>reset,s=>p(325)(14),cout=>p(326)(15));
FA_ff_12257:FAff port map(x=>p(293)(15),y=>p(294)(15),Cin=>p(295)(15),clock=>clock,reset=>reset,s=>p(325)(15),cout=>p(326)(16));
FA_ff_12258:FAff port map(x=>p(293)(16),y=>p(294)(16),Cin=>p(295)(16),clock=>clock,reset=>reset,s=>p(325)(16),cout=>p(326)(17));
FA_ff_12259:FAff port map(x=>p(293)(17),y=>p(294)(17),Cin=>p(295)(17),clock=>clock,reset=>reset,s=>p(325)(17),cout=>p(326)(18));
FA_ff_12260:FAff port map(x=>p(293)(18),y=>p(294)(18),Cin=>p(295)(18),clock=>clock,reset=>reset,s=>p(325)(18),cout=>p(326)(19));
FA_ff_12261:FAff port map(x=>p(293)(19),y=>p(294)(19),Cin=>p(295)(19),clock=>clock,reset=>reset,s=>p(325)(19),cout=>p(326)(20));
FA_ff_12262:FAff port map(x=>p(293)(20),y=>p(294)(20),Cin=>p(295)(20),clock=>clock,reset=>reset,s=>p(325)(20),cout=>p(326)(21));
FA_ff_12263:FAff port map(x=>p(293)(21),y=>p(294)(21),Cin=>p(295)(21),clock=>clock,reset=>reset,s=>p(325)(21),cout=>p(326)(22));
FA_ff_12264:FAff port map(x=>p(293)(22),y=>p(294)(22),Cin=>p(295)(22),clock=>clock,reset=>reset,s=>p(325)(22),cout=>p(326)(23));
FA_ff_12265:FAff port map(x=>p(293)(23),y=>p(294)(23),Cin=>p(295)(23),clock=>clock,reset=>reset,s=>p(325)(23),cout=>p(326)(24));
FA_ff_12266:FAff port map(x=>p(293)(24),y=>p(294)(24),Cin=>p(295)(24),clock=>clock,reset=>reset,s=>p(325)(24),cout=>p(326)(25));
FA_ff_12267:FAff port map(x=>p(293)(25),y=>p(294)(25),Cin=>p(295)(25),clock=>clock,reset=>reset,s=>p(325)(25),cout=>p(326)(26));
FA_ff_12268:FAff port map(x=>p(293)(26),y=>p(294)(26),Cin=>p(295)(26),clock=>clock,reset=>reset,s=>p(325)(26),cout=>p(326)(27));
FA_ff_12269:FAff port map(x=>p(293)(27),y=>p(294)(27),Cin=>p(295)(27),clock=>clock,reset=>reset,s=>p(325)(27),cout=>p(326)(28));
FA_ff_12270:FAff port map(x=>p(293)(28),y=>p(294)(28),Cin=>p(295)(28),clock=>clock,reset=>reset,s=>p(325)(28),cout=>p(326)(29));
FA_ff_12271:FAff port map(x=>p(293)(29),y=>p(294)(29),Cin=>p(295)(29),clock=>clock,reset=>reset,s=>p(325)(29),cout=>p(326)(30));
FA_ff_12272:FAff port map(x=>p(293)(30),y=>p(294)(30),Cin=>p(295)(30),clock=>clock,reset=>reset,s=>p(325)(30),cout=>p(326)(31));
FA_ff_12273:FAff port map(x=>p(293)(31),y=>p(294)(31),Cin=>p(295)(31),clock=>clock,reset=>reset,s=>p(325)(31),cout=>p(326)(32));
FA_ff_12274:FAff port map(x=>p(293)(32),y=>p(294)(32),Cin=>p(295)(32),clock=>clock,reset=>reset,s=>p(325)(32),cout=>p(326)(33));
FA_ff_12275:FAff port map(x=>p(293)(33),y=>p(294)(33),Cin=>p(295)(33),clock=>clock,reset=>reset,s=>p(325)(33),cout=>p(326)(34));
FA_ff_12276:FAff port map(x=>p(293)(34),y=>p(294)(34),Cin=>p(295)(34),clock=>clock,reset=>reset,s=>p(325)(34),cout=>p(326)(35));
FA_ff_12277:FAff port map(x=>p(293)(35),y=>p(294)(35),Cin=>p(295)(35),clock=>clock,reset=>reset,s=>p(325)(35),cout=>p(326)(36));
FA_ff_12278:FAff port map(x=>p(293)(36),y=>p(294)(36),Cin=>p(295)(36),clock=>clock,reset=>reset,s=>p(325)(36),cout=>p(326)(37));
FA_ff_12279:FAff port map(x=>p(293)(37),y=>p(294)(37),Cin=>p(295)(37),clock=>clock,reset=>reset,s=>p(325)(37),cout=>p(326)(38));
FA_ff_12280:FAff port map(x=>p(293)(38),y=>p(294)(38),Cin=>p(295)(38),clock=>clock,reset=>reset,s=>p(325)(38),cout=>p(326)(39));
FA_ff_12281:FAff port map(x=>p(293)(39),y=>p(294)(39),Cin=>p(295)(39),clock=>clock,reset=>reset,s=>p(325)(39),cout=>p(326)(40));
FA_ff_12282:FAff port map(x=>p(293)(40),y=>p(294)(40),Cin=>p(295)(40),clock=>clock,reset=>reset,s=>p(325)(40),cout=>p(326)(41));
FA_ff_12283:FAff port map(x=>p(293)(41),y=>p(294)(41),Cin=>p(295)(41),clock=>clock,reset=>reset,s=>p(325)(41),cout=>p(326)(42));
FA_ff_12284:FAff port map(x=>p(293)(42),y=>p(294)(42),Cin=>p(295)(42),clock=>clock,reset=>reset,s=>p(325)(42),cout=>p(326)(43));
FA_ff_12285:FAff port map(x=>p(293)(43),y=>p(294)(43),Cin=>p(295)(43),clock=>clock,reset=>reset,s=>p(325)(43),cout=>p(326)(44));
FA_ff_12286:FAff port map(x=>p(293)(44),y=>p(294)(44),Cin=>p(295)(44),clock=>clock,reset=>reset,s=>p(325)(44),cout=>p(326)(45));
FA_ff_12287:FAff port map(x=>p(293)(45),y=>p(294)(45),Cin=>p(295)(45),clock=>clock,reset=>reset,s=>p(325)(45),cout=>p(326)(46));
FA_ff_12288:FAff port map(x=>p(293)(46),y=>p(294)(46),Cin=>p(295)(46),clock=>clock,reset=>reset,s=>p(325)(46),cout=>p(326)(47));
FA_ff_12289:FAff port map(x=>p(293)(47),y=>p(294)(47),Cin=>p(295)(47),clock=>clock,reset=>reset,s=>p(325)(47),cout=>p(326)(48));
FA_ff_12290:FAff port map(x=>p(293)(48),y=>p(294)(48),Cin=>p(295)(48),clock=>clock,reset=>reset,s=>p(325)(48),cout=>p(326)(49));
FA_ff_12291:FAff port map(x=>p(293)(49),y=>p(294)(49),Cin=>p(295)(49),clock=>clock,reset=>reset,s=>p(325)(49),cout=>p(326)(50));
FA_ff_12292:FAff port map(x=>p(293)(50),y=>p(294)(50),Cin=>p(295)(50),clock=>clock,reset=>reset,s=>p(325)(50),cout=>p(326)(51));
FA_ff_12293:FAff port map(x=>p(293)(51),y=>p(294)(51),Cin=>p(295)(51),clock=>clock,reset=>reset,s=>p(325)(51),cout=>p(326)(52));
FA_ff_12294:FAff port map(x=>p(293)(52),y=>p(294)(52),Cin=>p(295)(52),clock=>clock,reset=>reset,s=>p(325)(52),cout=>p(326)(53));
FA_ff_12295:FAff port map(x=>p(293)(53),y=>p(294)(53),Cin=>p(295)(53),clock=>clock,reset=>reset,s=>p(325)(53),cout=>p(326)(54));
FA_ff_12296:FAff port map(x=>p(293)(54),y=>p(294)(54),Cin=>p(295)(54),clock=>clock,reset=>reset,s=>p(325)(54),cout=>p(326)(55));
FA_ff_12297:FAff port map(x=>p(293)(55),y=>p(294)(55),Cin=>p(295)(55),clock=>clock,reset=>reset,s=>p(325)(55),cout=>p(326)(56));
FA_ff_12298:FAff port map(x=>p(293)(56),y=>p(294)(56),Cin=>p(295)(56),clock=>clock,reset=>reset,s=>p(325)(56),cout=>p(326)(57));
FA_ff_12299:FAff port map(x=>p(293)(57),y=>p(294)(57),Cin=>p(295)(57),clock=>clock,reset=>reset,s=>p(325)(57),cout=>p(326)(58));
FA_ff_12300:FAff port map(x=>p(293)(58),y=>p(294)(58),Cin=>p(295)(58),clock=>clock,reset=>reset,s=>p(325)(58),cout=>p(326)(59));
FA_ff_12301:FAff port map(x=>p(293)(59),y=>p(294)(59),Cin=>p(295)(59),clock=>clock,reset=>reset,s=>p(325)(59),cout=>p(326)(60));
FA_ff_12302:FAff port map(x=>p(293)(60),y=>p(294)(60),Cin=>p(295)(60),clock=>clock,reset=>reset,s=>p(325)(60),cout=>p(326)(61));
FA_ff_12303:FAff port map(x=>p(293)(61),y=>p(294)(61),Cin=>p(295)(61),clock=>clock,reset=>reset,s=>p(325)(61),cout=>p(326)(62));
FA_ff_12304:FAff port map(x=>p(293)(62),y=>p(294)(62),Cin=>p(295)(62),clock=>clock,reset=>reset,s=>p(325)(62),cout=>p(326)(63));
FA_ff_12305:FAff port map(x=>p(293)(63),y=>p(294)(63),Cin=>p(295)(63),clock=>clock,reset=>reset,s=>p(325)(63),cout=>p(326)(64));
FA_ff_12306:FAff port map(x=>p(293)(64),y=>p(294)(64),Cin=>p(295)(64),clock=>clock,reset=>reset,s=>p(325)(64),cout=>p(326)(65));
FA_ff_12307:FAff port map(x=>p(293)(65),y=>p(294)(65),Cin=>p(295)(65),clock=>clock,reset=>reset,s=>p(325)(65),cout=>p(326)(66));
FA_ff_12308:FAff port map(x=>p(293)(66),y=>p(294)(66),Cin=>p(295)(66),clock=>clock,reset=>reset,s=>p(325)(66),cout=>p(326)(67));
FA_ff_12309:FAff port map(x=>p(293)(67),y=>p(294)(67),Cin=>p(295)(67),clock=>clock,reset=>reset,s=>p(325)(67),cout=>p(326)(68));
FA_ff_12310:FAff port map(x=>p(293)(68),y=>p(294)(68),Cin=>p(295)(68),clock=>clock,reset=>reset,s=>p(325)(68),cout=>p(326)(69));
FA_ff_12311:FAff port map(x=>p(293)(69),y=>p(294)(69),Cin=>p(295)(69),clock=>clock,reset=>reset,s=>p(325)(69),cout=>p(326)(70));
FA_ff_12312:FAff port map(x=>p(293)(70),y=>p(294)(70),Cin=>p(295)(70),clock=>clock,reset=>reset,s=>p(325)(70),cout=>p(326)(71));
FA_ff_12313:FAff port map(x=>p(293)(71),y=>p(294)(71),Cin=>p(295)(71),clock=>clock,reset=>reset,s=>p(325)(71),cout=>p(326)(72));
FA_ff_12314:FAff port map(x=>p(293)(72),y=>p(294)(72),Cin=>p(295)(72),clock=>clock,reset=>reset,s=>p(325)(72),cout=>p(326)(73));
FA_ff_12315:FAff port map(x=>p(293)(73),y=>p(294)(73),Cin=>p(295)(73),clock=>clock,reset=>reset,s=>p(325)(73),cout=>p(326)(74));
FA_ff_12316:FAff port map(x=>p(293)(74),y=>p(294)(74),Cin=>p(295)(74),clock=>clock,reset=>reset,s=>p(325)(74),cout=>p(326)(75));
FA_ff_12317:FAff port map(x=>p(293)(75),y=>p(294)(75),Cin=>p(295)(75),clock=>clock,reset=>reset,s=>p(325)(75),cout=>p(326)(76));
FA_ff_12318:FAff port map(x=>p(293)(76),y=>p(294)(76),Cin=>p(295)(76),clock=>clock,reset=>reset,s=>p(325)(76),cout=>p(326)(77));
FA_ff_12319:FAff port map(x=>p(293)(77),y=>p(294)(77),Cin=>p(295)(77),clock=>clock,reset=>reset,s=>p(325)(77),cout=>p(326)(78));
FA_ff_12320:FAff port map(x=>p(293)(78),y=>p(294)(78),Cin=>p(295)(78),clock=>clock,reset=>reset,s=>p(325)(78),cout=>p(326)(79));
FA_ff_12321:FAff port map(x=>p(293)(79),y=>p(294)(79),Cin=>p(295)(79),clock=>clock,reset=>reset,s=>p(325)(79),cout=>p(326)(80));
FA_ff_12322:FAff port map(x=>p(293)(80),y=>p(294)(80),Cin=>p(295)(80),clock=>clock,reset=>reset,s=>p(325)(80),cout=>p(326)(81));
FA_ff_12323:FAff port map(x=>p(293)(81),y=>p(294)(81),Cin=>p(295)(81),clock=>clock,reset=>reset,s=>p(325)(81),cout=>p(326)(82));
FA_ff_12324:FAff port map(x=>p(293)(82),y=>p(294)(82),Cin=>p(295)(82),clock=>clock,reset=>reset,s=>p(325)(82),cout=>p(326)(83));
FA_ff_12325:FAff port map(x=>p(293)(83),y=>p(294)(83),Cin=>p(295)(83),clock=>clock,reset=>reset,s=>p(325)(83),cout=>p(326)(84));
FA_ff_12326:FAff port map(x=>p(293)(84),y=>p(294)(84),Cin=>p(295)(84),clock=>clock,reset=>reset,s=>p(325)(84),cout=>p(326)(85));
FA_ff_12327:FAff port map(x=>p(293)(85),y=>p(294)(85),Cin=>p(295)(85),clock=>clock,reset=>reset,s=>p(325)(85),cout=>p(326)(86));
FA_ff_12328:FAff port map(x=>p(293)(86),y=>p(294)(86),Cin=>p(295)(86),clock=>clock,reset=>reset,s=>p(325)(86),cout=>p(326)(87));
FA_ff_12329:FAff port map(x=>p(293)(87),y=>p(294)(87),Cin=>p(295)(87),clock=>clock,reset=>reset,s=>p(325)(87),cout=>p(326)(88));
FA_ff_12330:FAff port map(x=>p(293)(88),y=>p(294)(88),Cin=>p(295)(88),clock=>clock,reset=>reset,s=>p(325)(88),cout=>p(326)(89));
FA_ff_12331:FAff port map(x=>p(293)(89),y=>p(294)(89),Cin=>p(295)(89),clock=>clock,reset=>reset,s=>p(325)(89),cout=>p(326)(90));
FA_ff_12332:FAff port map(x=>p(293)(90),y=>p(294)(90),Cin=>p(295)(90),clock=>clock,reset=>reset,s=>p(325)(90),cout=>p(326)(91));
FA_ff_12333:FAff port map(x=>p(293)(91),y=>p(294)(91),Cin=>p(295)(91),clock=>clock,reset=>reset,s=>p(325)(91),cout=>p(326)(92));
FA_ff_12334:FAff port map(x=>p(293)(92),y=>p(294)(92),Cin=>p(295)(92),clock=>clock,reset=>reset,s=>p(325)(92),cout=>p(326)(93));
FA_ff_12335:FAff port map(x=>p(293)(93),y=>p(294)(93),Cin=>p(295)(93),clock=>clock,reset=>reset,s=>p(325)(93),cout=>p(326)(94));
FA_ff_12336:FAff port map(x=>p(293)(94),y=>p(294)(94),Cin=>p(295)(94),clock=>clock,reset=>reset,s=>p(325)(94),cout=>p(326)(95));
FA_ff_12337:FAff port map(x=>p(293)(95),y=>p(294)(95),Cin=>p(295)(95),clock=>clock,reset=>reset,s=>p(325)(95),cout=>p(326)(96));
FA_ff_12338:FAff port map(x=>p(293)(96),y=>p(294)(96),Cin=>p(295)(96),clock=>clock,reset=>reset,s=>p(325)(96),cout=>p(326)(97));
FA_ff_12339:FAff port map(x=>p(293)(97),y=>p(294)(97),Cin=>p(295)(97),clock=>clock,reset=>reset,s=>p(325)(97),cout=>p(326)(98));
FA_ff_12340:FAff port map(x=>p(293)(98),y=>p(294)(98),Cin=>p(295)(98),clock=>clock,reset=>reset,s=>p(325)(98),cout=>p(326)(99));
FA_ff_12341:FAff port map(x=>p(293)(99),y=>p(294)(99),Cin=>p(295)(99),clock=>clock,reset=>reset,s=>p(325)(99),cout=>p(326)(100));
FA_ff_12342:FAff port map(x=>p(293)(100),y=>p(294)(100),Cin=>p(295)(100),clock=>clock,reset=>reset,s=>p(325)(100),cout=>p(326)(101));
FA_ff_12343:FAff port map(x=>p(293)(101),y=>p(294)(101),Cin=>p(295)(101),clock=>clock,reset=>reset,s=>p(325)(101),cout=>p(326)(102));
FA_ff_12344:FAff port map(x=>p(293)(102),y=>p(294)(102),Cin=>p(295)(102),clock=>clock,reset=>reset,s=>p(325)(102),cout=>p(326)(103));
FA_ff_12345:FAff port map(x=>p(293)(103),y=>p(294)(103),Cin=>p(295)(103),clock=>clock,reset=>reset,s=>p(325)(103),cout=>p(326)(104));
FA_ff_12346:FAff port map(x=>p(293)(104),y=>p(294)(104),Cin=>p(295)(104),clock=>clock,reset=>reset,s=>p(325)(104),cout=>p(326)(105));
FA_ff_12347:FAff port map(x=>p(293)(105),y=>p(294)(105),Cin=>p(295)(105),clock=>clock,reset=>reset,s=>p(325)(105),cout=>p(326)(106));
FA_ff_12348:FAff port map(x=>p(293)(106),y=>p(294)(106),Cin=>p(295)(106),clock=>clock,reset=>reset,s=>p(325)(106),cout=>p(326)(107));
FA_ff_12349:FAff port map(x=>p(293)(107),y=>p(294)(107),Cin=>p(295)(107),clock=>clock,reset=>reset,s=>p(325)(107),cout=>p(326)(108));
FA_ff_12350:FAff port map(x=>p(293)(108),y=>p(294)(108),Cin=>p(295)(108),clock=>clock,reset=>reset,s=>p(325)(108),cout=>p(326)(109));
FA_ff_12351:FAff port map(x=>p(293)(109),y=>p(294)(109),Cin=>p(295)(109),clock=>clock,reset=>reset,s=>p(325)(109),cout=>p(326)(110));
FA_ff_12352:FAff port map(x=>p(293)(110),y=>p(294)(110),Cin=>p(295)(110),clock=>clock,reset=>reset,s=>p(325)(110),cout=>p(326)(111));
FA_ff_12353:FAff port map(x=>p(293)(111),y=>p(294)(111),Cin=>p(295)(111),clock=>clock,reset=>reset,s=>p(325)(111),cout=>p(326)(112));
FA_ff_12354:FAff port map(x=>p(293)(112),y=>p(294)(112),Cin=>p(295)(112),clock=>clock,reset=>reset,s=>p(325)(112),cout=>p(326)(113));
FA_ff_12355:FAff port map(x=>p(293)(113),y=>p(294)(113),Cin=>p(295)(113),clock=>clock,reset=>reset,s=>p(325)(113),cout=>p(326)(114));
FA_ff_12356:FAff port map(x=>p(293)(114),y=>p(294)(114),Cin=>p(295)(114),clock=>clock,reset=>reset,s=>p(325)(114),cout=>p(326)(115));
FA_ff_12357:FAff port map(x=>p(293)(115),y=>p(294)(115),Cin=>p(295)(115),clock=>clock,reset=>reset,s=>p(325)(115),cout=>p(326)(116));
FA_ff_12358:FAff port map(x=>p(293)(116),y=>p(294)(116),Cin=>p(295)(116),clock=>clock,reset=>reset,s=>p(325)(116),cout=>p(326)(117));
FA_ff_12359:FAff port map(x=>p(293)(117),y=>p(294)(117),Cin=>p(295)(117),clock=>clock,reset=>reset,s=>p(325)(117),cout=>p(326)(118));
FA_ff_12360:FAff port map(x=>p(293)(118),y=>p(294)(118),Cin=>p(295)(118),clock=>clock,reset=>reset,s=>p(325)(118),cout=>p(326)(119));
FA_ff_12361:FAff port map(x=>p(293)(119),y=>p(294)(119),Cin=>p(295)(119),clock=>clock,reset=>reset,s=>p(325)(119),cout=>p(326)(120));
FA_ff_12362:FAff port map(x=>p(293)(120),y=>p(294)(120),Cin=>p(295)(120),clock=>clock,reset=>reset,s=>p(325)(120),cout=>p(326)(121));
FA_ff_12363:FAff port map(x=>p(293)(121),y=>p(294)(121),Cin=>p(295)(121),clock=>clock,reset=>reset,s=>p(325)(121),cout=>p(326)(122));
FA_ff_12364:FAff port map(x=>p(293)(122),y=>p(294)(122),Cin=>p(295)(122),clock=>clock,reset=>reset,s=>p(325)(122),cout=>p(326)(123));
FA_ff_12365:FAff port map(x=>p(293)(123),y=>p(294)(123),Cin=>p(295)(123),clock=>clock,reset=>reset,s=>p(325)(123),cout=>p(326)(124));
FA_ff_12366:FAff port map(x=>p(293)(124),y=>p(294)(124),Cin=>p(295)(124),clock=>clock,reset=>reset,s=>p(325)(124),cout=>p(326)(125));
FA_ff_12367:FAff port map(x=>p(293)(125),y=>p(294)(125),Cin=>p(295)(125),clock=>clock,reset=>reset,s=>p(325)(125),cout=>p(326)(126));
FA_ff_12368:FAff port map(x=>p(293)(126),y=>p(294)(126),Cin=>p(295)(126),clock=>clock,reset=>reset,s=>p(325)(126),cout=>p(326)(127));
FA_ff_12369:FAff port map(x=>p(293)(127),y=>p(294)(127),Cin=>p(295)(127),clock=>clock,reset=>reset,s=>p(325)(127),cout=>p(326)(128));
FA_ff_12370:FAff port map(x=>p(293)(128),y=>p(294)(128),Cin=>p(295)(128),clock=>clock,reset=>reset,s=>p(325)(128),cout=>p(326)(129));
FA_ff_12371:FAff port map(x=>p(293)(129),y=>p(294)(129),Cin=>p(295)(129),clock=>clock,reset=>reset,s=>p(325)(129),cout=>p(326)(130));
HA_ff_66:HAff port map(x=>p(296)(0),y=>p(298)(0),clock=>clock,reset=>reset,s=>p(327)(0),c=>p(328)(1));
FA_ff_12372:FAff port map(x=>p(296)(1),y=>p(297)(1),Cin=>p(298)(1),clock=>clock,reset=>reset,s=>p(327)(1),cout=>p(328)(2));
FA_ff_12373:FAff port map(x=>p(296)(2),y=>p(297)(2),Cin=>p(298)(2),clock=>clock,reset=>reset,s=>p(327)(2),cout=>p(328)(3));
FA_ff_12374:FAff port map(x=>p(296)(3),y=>p(297)(3),Cin=>p(298)(3),clock=>clock,reset=>reset,s=>p(327)(3),cout=>p(328)(4));
FA_ff_12375:FAff port map(x=>p(296)(4),y=>p(297)(4),Cin=>p(298)(4),clock=>clock,reset=>reset,s=>p(327)(4),cout=>p(328)(5));
FA_ff_12376:FAff port map(x=>p(296)(5),y=>p(297)(5),Cin=>p(298)(5),clock=>clock,reset=>reset,s=>p(327)(5),cout=>p(328)(6));
FA_ff_12377:FAff port map(x=>p(296)(6),y=>p(297)(6),Cin=>p(298)(6),clock=>clock,reset=>reset,s=>p(327)(6),cout=>p(328)(7));
FA_ff_12378:FAff port map(x=>p(296)(7),y=>p(297)(7),Cin=>p(298)(7),clock=>clock,reset=>reset,s=>p(327)(7),cout=>p(328)(8));
FA_ff_12379:FAff port map(x=>p(296)(8),y=>p(297)(8),Cin=>p(298)(8),clock=>clock,reset=>reset,s=>p(327)(8),cout=>p(328)(9));
FA_ff_12380:FAff port map(x=>p(296)(9),y=>p(297)(9),Cin=>p(298)(9),clock=>clock,reset=>reset,s=>p(327)(9),cout=>p(328)(10));
FA_ff_12381:FAff port map(x=>p(296)(10),y=>p(297)(10),Cin=>p(298)(10),clock=>clock,reset=>reset,s=>p(327)(10),cout=>p(328)(11));
FA_ff_12382:FAff port map(x=>p(296)(11),y=>p(297)(11),Cin=>p(298)(11),clock=>clock,reset=>reset,s=>p(327)(11),cout=>p(328)(12));
FA_ff_12383:FAff port map(x=>p(296)(12),y=>p(297)(12),Cin=>p(298)(12),clock=>clock,reset=>reset,s=>p(327)(12),cout=>p(328)(13));
FA_ff_12384:FAff port map(x=>p(296)(13),y=>p(297)(13),Cin=>p(298)(13),clock=>clock,reset=>reset,s=>p(327)(13),cout=>p(328)(14));
FA_ff_12385:FAff port map(x=>p(296)(14),y=>p(297)(14),Cin=>p(298)(14),clock=>clock,reset=>reset,s=>p(327)(14),cout=>p(328)(15));
FA_ff_12386:FAff port map(x=>p(296)(15),y=>p(297)(15),Cin=>p(298)(15),clock=>clock,reset=>reset,s=>p(327)(15),cout=>p(328)(16));
FA_ff_12387:FAff port map(x=>p(296)(16),y=>p(297)(16),Cin=>p(298)(16),clock=>clock,reset=>reset,s=>p(327)(16),cout=>p(328)(17));
FA_ff_12388:FAff port map(x=>p(296)(17),y=>p(297)(17),Cin=>p(298)(17),clock=>clock,reset=>reset,s=>p(327)(17),cout=>p(328)(18));
FA_ff_12389:FAff port map(x=>p(296)(18),y=>p(297)(18),Cin=>p(298)(18),clock=>clock,reset=>reset,s=>p(327)(18),cout=>p(328)(19));
FA_ff_12390:FAff port map(x=>p(296)(19),y=>p(297)(19),Cin=>p(298)(19),clock=>clock,reset=>reset,s=>p(327)(19),cout=>p(328)(20));
FA_ff_12391:FAff port map(x=>p(296)(20),y=>p(297)(20),Cin=>p(298)(20),clock=>clock,reset=>reset,s=>p(327)(20),cout=>p(328)(21));
FA_ff_12392:FAff port map(x=>p(296)(21),y=>p(297)(21),Cin=>p(298)(21),clock=>clock,reset=>reset,s=>p(327)(21),cout=>p(328)(22));
FA_ff_12393:FAff port map(x=>p(296)(22),y=>p(297)(22),Cin=>p(298)(22),clock=>clock,reset=>reset,s=>p(327)(22),cout=>p(328)(23));
FA_ff_12394:FAff port map(x=>p(296)(23),y=>p(297)(23),Cin=>p(298)(23),clock=>clock,reset=>reset,s=>p(327)(23),cout=>p(328)(24));
FA_ff_12395:FAff port map(x=>p(296)(24),y=>p(297)(24),Cin=>p(298)(24),clock=>clock,reset=>reset,s=>p(327)(24),cout=>p(328)(25));
FA_ff_12396:FAff port map(x=>p(296)(25),y=>p(297)(25),Cin=>p(298)(25),clock=>clock,reset=>reset,s=>p(327)(25),cout=>p(328)(26));
FA_ff_12397:FAff port map(x=>p(296)(26),y=>p(297)(26),Cin=>p(298)(26),clock=>clock,reset=>reset,s=>p(327)(26),cout=>p(328)(27));
FA_ff_12398:FAff port map(x=>p(296)(27),y=>p(297)(27),Cin=>p(298)(27),clock=>clock,reset=>reset,s=>p(327)(27),cout=>p(328)(28));
FA_ff_12399:FAff port map(x=>p(296)(28),y=>p(297)(28),Cin=>p(298)(28),clock=>clock,reset=>reset,s=>p(327)(28),cout=>p(328)(29));
FA_ff_12400:FAff port map(x=>p(296)(29),y=>p(297)(29),Cin=>p(298)(29),clock=>clock,reset=>reset,s=>p(327)(29),cout=>p(328)(30));
FA_ff_12401:FAff port map(x=>p(296)(30),y=>p(297)(30),Cin=>p(298)(30),clock=>clock,reset=>reset,s=>p(327)(30),cout=>p(328)(31));
FA_ff_12402:FAff port map(x=>p(296)(31),y=>p(297)(31),Cin=>p(298)(31),clock=>clock,reset=>reset,s=>p(327)(31),cout=>p(328)(32));
FA_ff_12403:FAff port map(x=>p(296)(32),y=>p(297)(32),Cin=>p(298)(32),clock=>clock,reset=>reset,s=>p(327)(32),cout=>p(328)(33));
FA_ff_12404:FAff port map(x=>p(296)(33),y=>p(297)(33),Cin=>p(298)(33),clock=>clock,reset=>reset,s=>p(327)(33),cout=>p(328)(34));
FA_ff_12405:FAff port map(x=>p(296)(34),y=>p(297)(34),Cin=>p(298)(34),clock=>clock,reset=>reset,s=>p(327)(34),cout=>p(328)(35));
FA_ff_12406:FAff port map(x=>p(296)(35),y=>p(297)(35),Cin=>p(298)(35),clock=>clock,reset=>reset,s=>p(327)(35),cout=>p(328)(36));
FA_ff_12407:FAff port map(x=>p(296)(36),y=>p(297)(36),Cin=>p(298)(36),clock=>clock,reset=>reset,s=>p(327)(36),cout=>p(328)(37));
FA_ff_12408:FAff port map(x=>p(296)(37),y=>p(297)(37),Cin=>p(298)(37),clock=>clock,reset=>reset,s=>p(327)(37),cout=>p(328)(38));
FA_ff_12409:FAff port map(x=>p(296)(38),y=>p(297)(38),Cin=>p(298)(38),clock=>clock,reset=>reset,s=>p(327)(38),cout=>p(328)(39));
FA_ff_12410:FAff port map(x=>p(296)(39),y=>p(297)(39),Cin=>p(298)(39),clock=>clock,reset=>reset,s=>p(327)(39),cout=>p(328)(40));
FA_ff_12411:FAff port map(x=>p(296)(40),y=>p(297)(40),Cin=>p(298)(40),clock=>clock,reset=>reset,s=>p(327)(40),cout=>p(328)(41));
FA_ff_12412:FAff port map(x=>p(296)(41),y=>p(297)(41),Cin=>p(298)(41),clock=>clock,reset=>reset,s=>p(327)(41),cout=>p(328)(42));
FA_ff_12413:FAff port map(x=>p(296)(42),y=>p(297)(42),Cin=>p(298)(42),clock=>clock,reset=>reset,s=>p(327)(42),cout=>p(328)(43));
FA_ff_12414:FAff port map(x=>p(296)(43),y=>p(297)(43),Cin=>p(298)(43),clock=>clock,reset=>reset,s=>p(327)(43),cout=>p(328)(44));
FA_ff_12415:FAff port map(x=>p(296)(44),y=>p(297)(44),Cin=>p(298)(44),clock=>clock,reset=>reset,s=>p(327)(44),cout=>p(328)(45));
FA_ff_12416:FAff port map(x=>p(296)(45),y=>p(297)(45),Cin=>p(298)(45),clock=>clock,reset=>reset,s=>p(327)(45),cout=>p(328)(46));
FA_ff_12417:FAff port map(x=>p(296)(46),y=>p(297)(46),Cin=>p(298)(46),clock=>clock,reset=>reset,s=>p(327)(46),cout=>p(328)(47));
FA_ff_12418:FAff port map(x=>p(296)(47),y=>p(297)(47),Cin=>p(298)(47),clock=>clock,reset=>reset,s=>p(327)(47),cout=>p(328)(48));
FA_ff_12419:FAff port map(x=>p(296)(48),y=>p(297)(48),Cin=>p(298)(48),clock=>clock,reset=>reset,s=>p(327)(48),cout=>p(328)(49));
FA_ff_12420:FAff port map(x=>p(296)(49),y=>p(297)(49),Cin=>p(298)(49),clock=>clock,reset=>reset,s=>p(327)(49),cout=>p(328)(50));
FA_ff_12421:FAff port map(x=>p(296)(50),y=>p(297)(50),Cin=>p(298)(50),clock=>clock,reset=>reset,s=>p(327)(50),cout=>p(328)(51));
FA_ff_12422:FAff port map(x=>p(296)(51),y=>p(297)(51),Cin=>p(298)(51),clock=>clock,reset=>reset,s=>p(327)(51),cout=>p(328)(52));
FA_ff_12423:FAff port map(x=>p(296)(52),y=>p(297)(52),Cin=>p(298)(52),clock=>clock,reset=>reset,s=>p(327)(52),cout=>p(328)(53));
FA_ff_12424:FAff port map(x=>p(296)(53),y=>p(297)(53),Cin=>p(298)(53),clock=>clock,reset=>reset,s=>p(327)(53),cout=>p(328)(54));
FA_ff_12425:FAff port map(x=>p(296)(54),y=>p(297)(54),Cin=>p(298)(54),clock=>clock,reset=>reset,s=>p(327)(54),cout=>p(328)(55));
FA_ff_12426:FAff port map(x=>p(296)(55),y=>p(297)(55),Cin=>p(298)(55),clock=>clock,reset=>reset,s=>p(327)(55),cout=>p(328)(56));
FA_ff_12427:FAff port map(x=>p(296)(56),y=>p(297)(56),Cin=>p(298)(56),clock=>clock,reset=>reset,s=>p(327)(56),cout=>p(328)(57));
FA_ff_12428:FAff port map(x=>p(296)(57),y=>p(297)(57),Cin=>p(298)(57),clock=>clock,reset=>reset,s=>p(327)(57),cout=>p(328)(58));
FA_ff_12429:FAff port map(x=>p(296)(58),y=>p(297)(58),Cin=>p(298)(58),clock=>clock,reset=>reset,s=>p(327)(58),cout=>p(328)(59));
FA_ff_12430:FAff port map(x=>p(296)(59),y=>p(297)(59),Cin=>p(298)(59),clock=>clock,reset=>reset,s=>p(327)(59),cout=>p(328)(60));
FA_ff_12431:FAff port map(x=>p(296)(60),y=>p(297)(60),Cin=>p(298)(60),clock=>clock,reset=>reset,s=>p(327)(60),cout=>p(328)(61));
FA_ff_12432:FAff port map(x=>p(296)(61),y=>p(297)(61),Cin=>p(298)(61),clock=>clock,reset=>reset,s=>p(327)(61),cout=>p(328)(62));
FA_ff_12433:FAff port map(x=>p(296)(62),y=>p(297)(62),Cin=>p(298)(62),clock=>clock,reset=>reset,s=>p(327)(62),cout=>p(328)(63));
FA_ff_12434:FAff port map(x=>p(296)(63),y=>p(297)(63),Cin=>p(298)(63),clock=>clock,reset=>reset,s=>p(327)(63),cout=>p(328)(64));
FA_ff_12435:FAff port map(x=>p(296)(64),y=>p(297)(64),Cin=>p(298)(64),clock=>clock,reset=>reset,s=>p(327)(64),cout=>p(328)(65));
FA_ff_12436:FAff port map(x=>p(296)(65),y=>p(297)(65),Cin=>p(298)(65),clock=>clock,reset=>reset,s=>p(327)(65),cout=>p(328)(66));
FA_ff_12437:FAff port map(x=>p(296)(66),y=>p(297)(66),Cin=>p(298)(66),clock=>clock,reset=>reset,s=>p(327)(66),cout=>p(328)(67));
FA_ff_12438:FAff port map(x=>p(296)(67),y=>p(297)(67),Cin=>p(298)(67),clock=>clock,reset=>reset,s=>p(327)(67),cout=>p(328)(68));
FA_ff_12439:FAff port map(x=>p(296)(68),y=>p(297)(68),Cin=>p(298)(68),clock=>clock,reset=>reset,s=>p(327)(68),cout=>p(328)(69));
FA_ff_12440:FAff port map(x=>p(296)(69),y=>p(297)(69),Cin=>p(298)(69),clock=>clock,reset=>reset,s=>p(327)(69),cout=>p(328)(70));
FA_ff_12441:FAff port map(x=>p(296)(70),y=>p(297)(70),Cin=>p(298)(70),clock=>clock,reset=>reset,s=>p(327)(70),cout=>p(328)(71));
FA_ff_12442:FAff port map(x=>p(296)(71),y=>p(297)(71),Cin=>p(298)(71),clock=>clock,reset=>reset,s=>p(327)(71),cout=>p(328)(72));
FA_ff_12443:FAff port map(x=>p(296)(72),y=>p(297)(72),Cin=>p(298)(72),clock=>clock,reset=>reset,s=>p(327)(72),cout=>p(328)(73));
FA_ff_12444:FAff port map(x=>p(296)(73),y=>p(297)(73),Cin=>p(298)(73),clock=>clock,reset=>reset,s=>p(327)(73),cout=>p(328)(74));
FA_ff_12445:FAff port map(x=>p(296)(74),y=>p(297)(74),Cin=>p(298)(74),clock=>clock,reset=>reset,s=>p(327)(74),cout=>p(328)(75));
FA_ff_12446:FAff port map(x=>p(296)(75),y=>p(297)(75),Cin=>p(298)(75),clock=>clock,reset=>reset,s=>p(327)(75),cout=>p(328)(76));
FA_ff_12447:FAff port map(x=>p(296)(76),y=>p(297)(76),Cin=>p(298)(76),clock=>clock,reset=>reset,s=>p(327)(76),cout=>p(328)(77));
FA_ff_12448:FAff port map(x=>p(296)(77),y=>p(297)(77),Cin=>p(298)(77),clock=>clock,reset=>reset,s=>p(327)(77),cout=>p(328)(78));
FA_ff_12449:FAff port map(x=>p(296)(78),y=>p(297)(78),Cin=>p(298)(78),clock=>clock,reset=>reset,s=>p(327)(78),cout=>p(328)(79));
FA_ff_12450:FAff port map(x=>p(296)(79),y=>p(297)(79),Cin=>p(298)(79),clock=>clock,reset=>reset,s=>p(327)(79),cout=>p(328)(80));
FA_ff_12451:FAff port map(x=>p(296)(80),y=>p(297)(80),Cin=>p(298)(80),clock=>clock,reset=>reset,s=>p(327)(80),cout=>p(328)(81));
FA_ff_12452:FAff port map(x=>p(296)(81),y=>p(297)(81),Cin=>p(298)(81),clock=>clock,reset=>reset,s=>p(327)(81),cout=>p(328)(82));
FA_ff_12453:FAff port map(x=>p(296)(82),y=>p(297)(82),Cin=>p(298)(82),clock=>clock,reset=>reset,s=>p(327)(82),cout=>p(328)(83));
FA_ff_12454:FAff port map(x=>p(296)(83),y=>p(297)(83),Cin=>p(298)(83),clock=>clock,reset=>reset,s=>p(327)(83),cout=>p(328)(84));
FA_ff_12455:FAff port map(x=>p(296)(84),y=>p(297)(84),Cin=>p(298)(84),clock=>clock,reset=>reset,s=>p(327)(84),cout=>p(328)(85));
FA_ff_12456:FAff port map(x=>p(296)(85),y=>p(297)(85),Cin=>p(298)(85),clock=>clock,reset=>reset,s=>p(327)(85),cout=>p(328)(86));
FA_ff_12457:FAff port map(x=>p(296)(86),y=>p(297)(86),Cin=>p(298)(86),clock=>clock,reset=>reset,s=>p(327)(86),cout=>p(328)(87));
FA_ff_12458:FAff port map(x=>p(296)(87),y=>p(297)(87),Cin=>p(298)(87),clock=>clock,reset=>reset,s=>p(327)(87),cout=>p(328)(88));
FA_ff_12459:FAff port map(x=>p(296)(88),y=>p(297)(88),Cin=>p(298)(88),clock=>clock,reset=>reset,s=>p(327)(88),cout=>p(328)(89));
FA_ff_12460:FAff port map(x=>p(296)(89),y=>p(297)(89),Cin=>p(298)(89),clock=>clock,reset=>reset,s=>p(327)(89),cout=>p(328)(90));
FA_ff_12461:FAff port map(x=>p(296)(90),y=>p(297)(90),Cin=>p(298)(90),clock=>clock,reset=>reset,s=>p(327)(90),cout=>p(328)(91));
FA_ff_12462:FAff port map(x=>p(296)(91),y=>p(297)(91),Cin=>p(298)(91),clock=>clock,reset=>reset,s=>p(327)(91),cout=>p(328)(92));
FA_ff_12463:FAff port map(x=>p(296)(92),y=>p(297)(92),Cin=>p(298)(92),clock=>clock,reset=>reset,s=>p(327)(92),cout=>p(328)(93));
FA_ff_12464:FAff port map(x=>p(296)(93),y=>p(297)(93),Cin=>p(298)(93),clock=>clock,reset=>reset,s=>p(327)(93),cout=>p(328)(94));
FA_ff_12465:FAff port map(x=>p(296)(94),y=>p(297)(94),Cin=>p(298)(94),clock=>clock,reset=>reset,s=>p(327)(94),cout=>p(328)(95));
FA_ff_12466:FAff port map(x=>p(296)(95),y=>p(297)(95),Cin=>p(298)(95),clock=>clock,reset=>reset,s=>p(327)(95),cout=>p(328)(96));
FA_ff_12467:FAff port map(x=>p(296)(96),y=>p(297)(96),Cin=>p(298)(96),clock=>clock,reset=>reset,s=>p(327)(96),cout=>p(328)(97));
FA_ff_12468:FAff port map(x=>p(296)(97),y=>p(297)(97),Cin=>p(298)(97),clock=>clock,reset=>reset,s=>p(327)(97),cout=>p(328)(98));
FA_ff_12469:FAff port map(x=>p(296)(98),y=>p(297)(98),Cin=>p(298)(98),clock=>clock,reset=>reset,s=>p(327)(98),cout=>p(328)(99));
FA_ff_12470:FAff port map(x=>p(296)(99),y=>p(297)(99),Cin=>p(298)(99),clock=>clock,reset=>reset,s=>p(327)(99),cout=>p(328)(100));
FA_ff_12471:FAff port map(x=>p(296)(100),y=>p(297)(100),Cin=>p(298)(100),clock=>clock,reset=>reset,s=>p(327)(100),cout=>p(328)(101));
FA_ff_12472:FAff port map(x=>p(296)(101),y=>p(297)(101),Cin=>p(298)(101),clock=>clock,reset=>reset,s=>p(327)(101),cout=>p(328)(102));
FA_ff_12473:FAff port map(x=>p(296)(102),y=>p(297)(102),Cin=>p(298)(102),clock=>clock,reset=>reset,s=>p(327)(102),cout=>p(328)(103));
FA_ff_12474:FAff port map(x=>p(296)(103),y=>p(297)(103),Cin=>p(298)(103),clock=>clock,reset=>reset,s=>p(327)(103),cout=>p(328)(104));
FA_ff_12475:FAff port map(x=>p(296)(104),y=>p(297)(104),Cin=>p(298)(104),clock=>clock,reset=>reset,s=>p(327)(104),cout=>p(328)(105));
FA_ff_12476:FAff port map(x=>p(296)(105),y=>p(297)(105),Cin=>p(298)(105),clock=>clock,reset=>reset,s=>p(327)(105),cout=>p(328)(106));
FA_ff_12477:FAff port map(x=>p(296)(106),y=>p(297)(106),Cin=>p(298)(106),clock=>clock,reset=>reset,s=>p(327)(106),cout=>p(328)(107));
FA_ff_12478:FAff port map(x=>p(296)(107),y=>p(297)(107),Cin=>p(298)(107),clock=>clock,reset=>reset,s=>p(327)(107),cout=>p(328)(108));
FA_ff_12479:FAff port map(x=>p(296)(108),y=>p(297)(108),Cin=>p(298)(108),clock=>clock,reset=>reset,s=>p(327)(108),cout=>p(328)(109));
FA_ff_12480:FAff port map(x=>p(296)(109),y=>p(297)(109),Cin=>p(298)(109),clock=>clock,reset=>reset,s=>p(327)(109),cout=>p(328)(110));
FA_ff_12481:FAff port map(x=>p(296)(110),y=>p(297)(110),Cin=>p(298)(110),clock=>clock,reset=>reset,s=>p(327)(110),cout=>p(328)(111));
FA_ff_12482:FAff port map(x=>p(296)(111),y=>p(297)(111),Cin=>p(298)(111),clock=>clock,reset=>reset,s=>p(327)(111),cout=>p(328)(112));
FA_ff_12483:FAff port map(x=>p(296)(112),y=>p(297)(112),Cin=>p(298)(112),clock=>clock,reset=>reset,s=>p(327)(112),cout=>p(328)(113));
FA_ff_12484:FAff port map(x=>p(296)(113),y=>p(297)(113),Cin=>p(298)(113),clock=>clock,reset=>reset,s=>p(327)(113),cout=>p(328)(114));
FA_ff_12485:FAff port map(x=>p(296)(114),y=>p(297)(114),Cin=>p(298)(114),clock=>clock,reset=>reset,s=>p(327)(114),cout=>p(328)(115));
FA_ff_12486:FAff port map(x=>p(296)(115),y=>p(297)(115),Cin=>p(298)(115),clock=>clock,reset=>reset,s=>p(327)(115),cout=>p(328)(116));
FA_ff_12487:FAff port map(x=>p(296)(116),y=>p(297)(116),Cin=>p(298)(116),clock=>clock,reset=>reset,s=>p(327)(116),cout=>p(328)(117));
FA_ff_12488:FAff port map(x=>p(296)(117),y=>p(297)(117),Cin=>p(298)(117),clock=>clock,reset=>reset,s=>p(327)(117),cout=>p(328)(118));
FA_ff_12489:FAff port map(x=>p(296)(118),y=>p(297)(118),Cin=>p(298)(118),clock=>clock,reset=>reset,s=>p(327)(118),cout=>p(328)(119));
FA_ff_12490:FAff port map(x=>p(296)(119),y=>p(297)(119),Cin=>p(298)(119),clock=>clock,reset=>reset,s=>p(327)(119),cout=>p(328)(120));
FA_ff_12491:FAff port map(x=>p(296)(120),y=>p(297)(120),Cin=>p(298)(120),clock=>clock,reset=>reset,s=>p(327)(120),cout=>p(328)(121));
FA_ff_12492:FAff port map(x=>p(296)(121),y=>p(297)(121),Cin=>p(298)(121),clock=>clock,reset=>reset,s=>p(327)(121),cout=>p(328)(122));
FA_ff_12493:FAff port map(x=>p(296)(122),y=>p(297)(122),Cin=>p(298)(122),clock=>clock,reset=>reset,s=>p(327)(122),cout=>p(328)(123));
FA_ff_12494:FAff port map(x=>p(296)(123),y=>p(297)(123),Cin=>p(298)(123),clock=>clock,reset=>reset,s=>p(327)(123),cout=>p(328)(124));
FA_ff_12495:FAff port map(x=>p(296)(124),y=>p(297)(124),Cin=>p(298)(124),clock=>clock,reset=>reset,s=>p(327)(124),cout=>p(328)(125));
FA_ff_12496:FAff port map(x=>p(296)(125),y=>p(297)(125),Cin=>p(298)(125),clock=>clock,reset=>reset,s=>p(327)(125),cout=>p(328)(126));
FA_ff_12497:FAff port map(x=>p(296)(126),y=>p(297)(126),Cin=>p(298)(126),clock=>clock,reset=>reset,s=>p(327)(126),cout=>p(328)(127));
FA_ff_12498:FAff port map(x=>p(296)(127),y=>p(297)(127),Cin=>p(298)(127),clock=>clock,reset=>reset,s=>p(327)(127),cout=>p(328)(128));
FA_ff_12499:FAff port map(x=>p(296)(128),y=>p(297)(128),Cin=>p(298)(128),clock=>clock,reset=>reset,s=>p(327)(128),cout=>p(328)(129));
HA_ff_67:HAff port map(x=>p(297)(129),y=>p(298)(129),clock=>clock,reset=>reset,s=>p(327)(129),c=>p(328)(130));
p(329)(0)<=p(300)(0);
HA_ff_68:HAff port map(x=>p(300)(1),y=>p(301)(1),clock=>clock,reset=>reset,s=>p(329)(1),c=>p(330)(2));
FA_ff_12500:FAff port map(x=>p(299)(2),y=>p(300)(2),Cin=>p(301)(2),clock=>clock,reset=>reset,s=>p(329)(2),cout=>p(330)(3));
FA_ff_12501:FAff port map(x=>p(299)(3),y=>p(300)(3),Cin=>p(301)(3),clock=>clock,reset=>reset,s=>p(329)(3),cout=>p(330)(4));
FA_ff_12502:FAff port map(x=>p(299)(4),y=>p(300)(4),Cin=>p(301)(4),clock=>clock,reset=>reset,s=>p(329)(4),cout=>p(330)(5));
FA_ff_12503:FAff port map(x=>p(299)(5),y=>p(300)(5),Cin=>p(301)(5),clock=>clock,reset=>reset,s=>p(329)(5),cout=>p(330)(6));
FA_ff_12504:FAff port map(x=>p(299)(6),y=>p(300)(6),Cin=>p(301)(6),clock=>clock,reset=>reset,s=>p(329)(6),cout=>p(330)(7));
FA_ff_12505:FAff port map(x=>p(299)(7),y=>p(300)(7),Cin=>p(301)(7),clock=>clock,reset=>reset,s=>p(329)(7),cout=>p(330)(8));
FA_ff_12506:FAff port map(x=>p(299)(8),y=>p(300)(8),Cin=>p(301)(8),clock=>clock,reset=>reset,s=>p(329)(8),cout=>p(330)(9));
FA_ff_12507:FAff port map(x=>p(299)(9),y=>p(300)(9),Cin=>p(301)(9),clock=>clock,reset=>reset,s=>p(329)(9),cout=>p(330)(10));
FA_ff_12508:FAff port map(x=>p(299)(10),y=>p(300)(10),Cin=>p(301)(10),clock=>clock,reset=>reset,s=>p(329)(10),cout=>p(330)(11));
FA_ff_12509:FAff port map(x=>p(299)(11),y=>p(300)(11),Cin=>p(301)(11),clock=>clock,reset=>reset,s=>p(329)(11),cout=>p(330)(12));
FA_ff_12510:FAff port map(x=>p(299)(12),y=>p(300)(12),Cin=>p(301)(12),clock=>clock,reset=>reset,s=>p(329)(12),cout=>p(330)(13));
FA_ff_12511:FAff port map(x=>p(299)(13),y=>p(300)(13),Cin=>p(301)(13),clock=>clock,reset=>reset,s=>p(329)(13),cout=>p(330)(14));
FA_ff_12512:FAff port map(x=>p(299)(14),y=>p(300)(14),Cin=>p(301)(14),clock=>clock,reset=>reset,s=>p(329)(14),cout=>p(330)(15));
FA_ff_12513:FAff port map(x=>p(299)(15),y=>p(300)(15),Cin=>p(301)(15),clock=>clock,reset=>reset,s=>p(329)(15),cout=>p(330)(16));
FA_ff_12514:FAff port map(x=>p(299)(16),y=>p(300)(16),Cin=>p(301)(16),clock=>clock,reset=>reset,s=>p(329)(16),cout=>p(330)(17));
FA_ff_12515:FAff port map(x=>p(299)(17),y=>p(300)(17),Cin=>p(301)(17),clock=>clock,reset=>reset,s=>p(329)(17),cout=>p(330)(18));
FA_ff_12516:FAff port map(x=>p(299)(18),y=>p(300)(18),Cin=>p(301)(18),clock=>clock,reset=>reset,s=>p(329)(18),cout=>p(330)(19));
FA_ff_12517:FAff port map(x=>p(299)(19),y=>p(300)(19),Cin=>p(301)(19),clock=>clock,reset=>reset,s=>p(329)(19),cout=>p(330)(20));
FA_ff_12518:FAff port map(x=>p(299)(20),y=>p(300)(20),Cin=>p(301)(20),clock=>clock,reset=>reset,s=>p(329)(20),cout=>p(330)(21));
FA_ff_12519:FAff port map(x=>p(299)(21),y=>p(300)(21),Cin=>p(301)(21),clock=>clock,reset=>reset,s=>p(329)(21),cout=>p(330)(22));
FA_ff_12520:FAff port map(x=>p(299)(22),y=>p(300)(22),Cin=>p(301)(22),clock=>clock,reset=>reset,s=>p(329)(22),cout=>p(330)(23));
FA_ff_12521:FAff port map(x=>p(299)(23),y=>p(300)(23),Cin=>p(301)(23),clock=>clock,reset=>reset,s=>p(329)(23),cout=>p(330)(24));
FA_ff_12522:FAff port map(x=>p(299)(24),y=>p(300)(24),Cin=>p(301)(24),clock=>clock,reset=>reset,s=>p(329)(24),cout=>p(330)(25));
FA_ff_12523:FAff port map(x=>p(299)(25),y=>p(300)(25),Cin=>p(301)(25),clock=>clock,reset=>reset,s=>p(329)(25),cout=>p(330)(26));
FA_ff_12524:FAff port map(x=>p(299)(26),y=>p(300)(26),Cin=>p(301)(26),clock=>clock,reset=>reset,s=>p(329)(26),cout=>p(330)(27));
FA_ff_12525:FAff port map(x=>p(299)(27),y=>p(300)(27),Cin=>p(301)(27),clock=>clock,reset=>reset,s=>p(329)(27),cout=>p(330)(28));
FA_ff_12526:FAff port map(x=>p(299)(28),y=>p(300)(28),Cin=>p(301)(28),clock=>clock,reset=>reset,s=>p(329)(28),cout=>p(330)(29));
FA_ff_12527:FAff port map(x=>p(299)(29),y=>p(300)(29),Cin=>p(301)(29),clock=>clock,reset=>reset,s=>p(329)(29),cout=>p(330)(30));
FA_ff_12528:FAff port map(x=>p(299)(30),y=>p(300)(30),Cin=>p(301)(30),clock=>clock,reset=>reset,s=>p(329)(30),cout=>p(330)(31));
FA_ff_12529:FAff port map(x=>p(299)(31),y=>p(300)(31),Cin=>p(301)(31),clock=>clock,reset=>reset,s=>p(329)(31),cout=>p(330)(32));
FA_ff_12530:FAff port map(x=>p(299)(32),y=>p(300)(32),Cin=>p(301)(32),clock=>clock,reset=>reset,s=>p(329)(32),cout=>p(330)(33));
FA_ff_12531:FAff port map(x=>p(299)(33),y=>p(300)(33),Cin=>p(301)(33),clock=>clock,reset=>reset,s=>p(329)(33),cout=>p(330)(34));
FA_ff_12532:FAff port map(x=>p(299)(34),y=>p(300)(34),Cin=>p(301)(34),clock=>clock,reset=>reset,s=>p(329)(34),cout=>p(330)(35));
FA_ff_12533:FAff port map(x=>p(299)(35),y=>p(300)(35),Cin=>p(301)(35),clock=>clock,reset=>reset,s=>p(329)(35),cout=>p(330)(36));
FA_ff_12534:FAff port map(x=>p(299)(36),y=>p(300)(36),Cin=>p(301)(36),clock=>clock,reset=>reset,s=>p(329)(36),cout=>p(330)(37));
FA_ff_12535:FAff port map(x=>p(299)(37),y=>p(300)(37),Cin=>p(301)(37),clock=>clock,reset=>reset,s=>p(329)(37),cout=>p(330)(38));
FA_ff_12536:FAff port map(x=>p(299)(38),y=>p(300)(38),Cin=>p(301)(38),clock=>clock,reset=>reset,s=>p(329)(38),cout=>p(330)(39));
FA_ff_12537:FAff port map(x=>p(299)(39),y=>p(300)(39),Cin=>p(301)(39),clock=>clock,reset=>reset,s=>p(329)(39),cout=>p(330)(40));
FA_ff_12538:FAff port map(x=>p(299)(40),y=>p(300)(40),Cin=>p(301)(40),clock=>clock,reset=>reset,s=>p(329)(40),cout=>p(330)(41));
FA_ff_12539:FAff port map(x=>p(299)(41),y=>p(300)(41),Cin=>p(301)(41),clock=>clock,reset=>reset,s=>p(329)(41),cout=>p(330)(42));
FA_ff_12540:FAff port map(x=>p(299)(42),y=>p(300)(42),Cin=>p(301)(42),clock=>clock,reset=>reset,s=>p(329)(42),cout=>p(330)(43));
FA_ff_12541:FAff port map(x=>p(299)(43),y=>p(300)(43),Cin=>p(301)(43),clock=>clock,reset=>reset,s=>p(329)(43),cout=>p(330)(44));
FA_ff_12542:FAff port map(x=>p(299)(44),y=>p(300)(44),Cin=>p(301)(44),clock=>clock,reset=>reset,s=>p(329)(44),cout=>p(330)(45));
FA_ff_12543:FAff port map(x=>p(299)(45),y=>p(300)(45),Cin=>p(301)(45),clock=>clock,reset=>reset,s=>p(329)(45),cout=>p(330)(46));
FA_ff_12544:FAff port map(x=>p(299)(46),y=>p(300)(46),Cin=>p(301)(46),clock=>clock,reset=>reset,s=>p(329)(46),cout=>p(330)(47));
FA_ff_12545:FAff port map(x=>p(299)(47),y=>p(300)(47),Cin=>p(301)(47),clock=>clock,reset=>reset,s=>p(329)(47),cout=>p(330)(48));
FA_ff_12546:FAff port map(x=>p(299)(48),y=>p(300)(48),Cin=>p(301)(48),clock=>clock,reset=>reset,s=>p(329)(48),cout=>p(330)(49));
FA_ff_12547:FAff port map(x=>p(299)(49),y=>p(300)(49),Cin=>p(301)(49),clock=>clock,reset=>reset,s=>p(329)(49),cout=>p(330)(50));
FA_ff_12548:FAff port map(x=>p(299)(50),y=>p(300)(50),Cin=>p(301)(50),clock=>clock,reset=>reset,s=>p(329)(50),cout=>p(330)(51));
FA_ff_12549:FAff port map(x=>p(299)(51),y=>p(300)(51),Cin=>p(301)(51),clock=>clock,reset=>reset,s=>p(329)(51),cout=>p(330)(52));
FA_ff_12550:FAff port map(x=>p(299)(52),y=>p(300)(52),Cin=>p(301)(52),clock=>clock,reset=>reset,s=>p(329)(52),cout=>p(330)(53));
FA_ff_12551:FAff port map(x=>p(299)(53),y=>p(300)(53),Cin=>p(301)(53),clock=>clock,reset=>reset,s=>p(329)(53),cout=>p(330)(54));
FA_ff_12552:FAff port map(x=>p(299)(54),y=>p(300)(54),Cin=>p(301)(54),clock=>clock,reset=>reset,s=>p(329)(54),cout=>p(330)(55));
FA_ff_12553:FAff port map(x=>p(299)(55),y=>p(300)(55),Cin=>p(301)(55),clock=>clock,reset=>reset,s=>p(329)(55),cout=>p(330)(56));
FA_ff_12554:FAff port map(x=>p(299)(56),y=>p(300)(56),Cin=>p(301)(56),clock=>clock,reset=>reset,s=>p(329)(56),cout=>p(330)(57));
FA_ff_12555:FAff port map(x=>p(299)(57),y=>p(300)(57),Cin=>p(301)(57),clock=>clock,reset=>reset,s=>p(329)(57),cout=>p(330)(58));
FA_ff_12556:FAff port map(x=>p(299)(58),y=>p(300)(58),Cin=>p(301)(58),clock=>clock,reset=>reset,s=>p(329)(58),cout=>p(330)(59));
FA_ff_12557:FAff port map(x=>p(299)(59),y=>p(300)(59),Cin=>p(301)(59),clock=>clock,reset=>reset,s=>p(329)(59),cout=>p(330)(60));
FA_ff_12558:FAff port map(x=>p(299)(60),y=>p(300)(60),Cin=>p(301)(60),clock=>clock,reset=>reset,s=>p(329)(60),cout=>p(330)(61));
FA_ff_12559:FAff port map(x=>p(299)(61),y=>p(300)(61),Cin=>p(301)(61),clock=>clock,reset=>reset,s=>p(329)(61),cout=>p(330)(62));
FA_ff_12560:FAff port map(x=>p(299)(62),y=>p(300)(62),Cin=>p(301)(62),clock=>clock,reset=>reset,s=>p(329)(62),cout=>p(330)(63));
FA_ff_12561:FAff port map(x=>p(299)(63),y=>p(300)(63),Cin=>p(301)(63),clock=>clock,reset=>reset,s=>p(329)(63),cout=>p(330)(64));
FA_ff_12562:FAff port map(x=>p(299)(64),y=>p(300)(64),Cin=>p(301)(64),clock=>clock,reset=>reset,s=>p(329)(64),cout=>p(330)(65));
FA_ff_12563:FAff port map(x=>p(299)(65),y=>p(300)(65),Cin=>p(301)(65),clock=>clock,reset=>reset,s=>p(329)(65),cout=>p(330)(66));
FA_ff_12564:FAff port map(x=>p(299)(66),y=>p(300)(66),Cin=>p(301)(66),clock=>clock,reset=>reset,s=>p(329)(66),cout=>p(330)(67));
FA_ff_12565:FAff port map(x=>p(299)(67),y=>p(300)(67),Cin=>p(301)(67),clock=>clock,reset=>reset,s=>p(329)(67),cout=>p(330)(68));
FA_ff_12566:FAff port map(x=>p(299)(68),y=>p(300)(68),Cin=>p(301)(68),clock=>clock,reset=>reset,s=>p(329)(68),cout=>p(330)(69));
FA_ff_12567:FAff port map(x=>p(299)(69),y=>p(300)(69),Cin=>p(301)(69),clock=>clock,reset=>reset,s=>p(329)(69),cout=>p(330)(70));
FA_ff_12568:FAff port map(x=>p(299)(70),y=>p(300)(70),Cin=>p(301)(70),clock=>clock,reset=>reset,s=>p(329)(70),cout=>p(330)(71));
FA_ff_12569:FAff port map(x=>p(299)(71),y=>p(300)(71),Cin=>p(301)(71),clock=>clock,reset=>reset,s=>p(329)(71),cout=>p(330)(72));
FA_ff_12570:FAff port map(x=>p(299)(72),y=>p(300)(72),Cin=>p(301)(72),clock=>clock,reset=>reset,s=>p(329)(72),cout=>p(330)(73));
FA_ff_12571:FAff port map(x=>p(299)(73),y=>p(300)(73),Cin=>p(301)(73),clock=>clock,reset=>reset,s=>p(329)(73),cout=>p(330)(74));
FA_ff_12572:FAff port map(x=>p(299)(74),y=>p(300)(74),Cin=>p(301)(74),clock=>clock,reset=>reset,s=>p(329)(74),cout=>p(330)(75));
FA_ff_12573:FAff port map(x=>p(299)(75),y=>p(300)(75),Cin=>p(301)(75),clock=>clock,reset=>reset,s=>p(329)(75),cout=>p(330)(76));
FA_ff_12574:FAff port map(x=>p(299)(76),y=>p(300)(76),Cin=>p(301)(76),clock=>clock,reset=>reset,s=>p(329)(76),cout=>p(330)(77));
FA_ff_12575:FAff port map(x=>p(299)(77),y=>p(300)(77),Cin=>p(301)(77),clock=>clock,reset=>reset,s=>p(329)(77),cout=>p(330)(78));
FA_ff_12576:FAff port map(x=>p(299)(78),y=>p(300)(78),Cin=>p(301)(78),clock=>clock,reset=>reset,s=>p(329)(78),cout=>p(330)(79));
FA_ff_12577:FAff port map(x=>p(299)(79),y=>p(300)(79),Cin=>p(301)(79),clock=>clock,reset=>reset,s=>p(329)(79),cout=>p(330)(80));
FA_ff_12578:FAff port map(x=>p(299)(80),y=>p(300)(80),Cin=>p(301)(80),clock=>clock,reset=>reset,s=>p(329)(80),cout=>p(330)(81));
FA_ff_12579:FAff port map(x=>p(299)(81),y=>p(300)(81),Cin=>p(301)(81),clock=>clock,reset=>reset,s=>p(329)(81),cout=>p(330)(82));
FA_ff_12580:FAff port map(x=>p(299)(82),y=>p(300)(82),Cin=>p(301)(82),clock=>clock,reset=>reset,s=>p(329)(82),cout=>p(330)(83));
FA_ff_12581:FAff port map(x=>p(299)(83),y=>p(300)(83),Cin=>p(301)(83),clock=>clock,reset=>reset,s=>p(329)(83),cout=>p(330)(84));
FA_ff_12582:FAff port map(x=>p(299)(84),y=>p(300)(84),Cin=>p(301)(84),clock=>clock,reset=>reset,s=>p(329)(84),cout=>p(330)(85));
FA_ff_12583:FAff port map(x=>p(299)(85),y=>p(300)(85),Cin=>p(301)(85),clock=>clock,reset=>reset,s=>p(329)(85),cout=>p(330)(86));
FA_ff_12584:FAff port map(x=>p(299)(86),y=>p(300)(86),Cin=>p(301)(86),clock=>clock,reset=>reset,s=>p(329)(86),cout=>p(330)(87));
FA_ff_12585:FAff port map(x=>p(299)(87),y=>p(300)(87),Cin=>p(301)(87),clock=>clock,reset=>reset,s=>p(329)(87),cout=>p(330)(88));
FA_ff_12586:FAff port map(x=>p(299)(88),y=>p(300)(88),Cin=>p(301)(88),clock=>clock,reset=>reset,s=>p(329)(88),cout=>p(330)(89));
FA_ff_12587:FAff port map(x=>p(299)(89),y=>p(300)(89),Cin=>p(301)(89),clock=>clock,reset=>reset,s=>p(329)(89),cout=>p(330)(90));
FA_ff_12588:FAff port map(x=>p(299)(90),y=>p(300)(90),Cin=>p(301)(90),clock=>clock,reset=>reset,s=>p(329)(90),cout=>p(330)(91));
FA_ff_12589:FAff port map(x=>p(299)(91),y=>p(300)(91),Cin=>p(301)(91),clock=>clock,reset=>reset,s=>p(329)(91),cout=>p(330)(92));
FA_ff_12590:FAff port map(x=>p(299)(92),y=>p(300)(92),Cin=>p(301)(92),clock=>clock,reset=>reset,s=>p(329)(92),cout=>p(330)(93));
FA_ff_12591:FAff port map(x=>p(299)(93),y=>p(300)(93),Cin=>p(301)(93),clock=>clock,reset=>reset,s=>p(329)(93),cout=>p(330)(94));
FA_ff_12592:FAff port map(x=>p(299)(94),y=>p(300)(94),Cin=>p(301)(94),clock=>clock,reset=>reset,s=>p(329)(94),cout=>p(330)(95));
FA_ff_12593:FAff port map(x=>p(299)(95),y=>p(300)(95),Cin=>p(301)(95),clock=>clock,reset=>reset,s=>p(329)(95),cout=>p(330)(96));
FA_ff_12594:FAff port map(x=>p(299)(96),y=>p(300)(96),Cin=>p(301)(96),clock=>clock,reset=>reset,s=>p(329)(96),cout=>p(330)(97));
FA_ff_12595:FAff port map(x=>p(299)(97),y=>p(300)(97),Cin=>p(301)(97),clock=>clock,reset=>reset,s=>p(329)(97),cout=>p(330)(98));
FA_ff_12596:FAff port map(x=>p(299)(98),y=>p(300)(98),Cin=>p(301)(98),clock=>clock,reset=>reset,s=>p(329)(98),cout=>p(330)(99));
FA_ff_12597:FAff port map(x=>p(299)(99),y=>p(300)(99),Cin=>p(301)(99),clock=>clock,reset=>reset,s=>p(329)(99),cout=>p(330)(100));
FA_ff_12598:FAff port map(x=>p(299)(100),y=>p(300)(100),Cin=>p(301)(100),clock=>clock,reset=>reset,s=>p(329)(100),cout=>p(330)(101));
FA_ff_12599:FAff port map(x=>p(299)(101),y=>p(300)(101),Cin=>p(301)(101),clock=>clock,reset=>reset,s=>p(329)(101),cout=>p(330)(102));
FA_ff_12600:FAff port map(x=>p(299)(102),y=>p(300)(102),Cin=>p(301)(102),clock=>clock,reset=>reset,s=>p(329)(102),cout=>p(330)(103));
FA_ff_12601:FAff port map(x=>p(299)(103),y=>p(300)(103),Cin=>p(301)(103),clock=>clock,reset=>reset,s=>p(329)(103),cout=>p(330)(104));
FA_ff_12602:FAff port map(x=>p(299)(104),y=>p(300)(104),Cin=>p(301)(104),clock=>clock,reset=>reset,s=>p(329)(104),cout=>p(330)(105));
FA_ff_12603:FAff port map(x=>p(299)(105),y=>p(300)(105),Cin=>p(301)(105),clock=>clock,reset=>reset,s=>p(329)(105),cout=>p(330)(106));
FA_ff_12604:FAff port map(x=>p(299)(106),y=>p(300)(106),Cin=>p(301)(106),clock=>clock,reset=>reset,s=>p(329)(106),cout=>p(330)(107));
FA_ff_12605:FAff port map(x=>p(299)(107),y=>p(300)(107),Cin=>p(301)(107),clock=>clock,reset=>reset,s=>p(329)(107),cout=>p(330)(108));
FA_ff_12606:FAff port map(x=>p(299)(108),y=>p(300)(108),Cin=>p(301)(108),clock=>clock,reset=>reset,s=>p(329)(108),cout=>p(330)(109));
FA_ff_12607:FAff port map(x=>p(299)(109),y=>p(300)(109),Cin=>p(301)(109),clock=>clock,reset=>reset,s=>p(329)(109),cout=>p(330)(110));
FA_ff_12608:FAff port map(x=>p(299)(110),y=>p(300)(110),Cin=>p(301)(110),clock=>clock,reset=>reset,s=>p(329)(110),cout=>p(330)(111));
FA_ff_12609:FAff port map(x=>p(299)(111),y=>p(300)(111),Cin=>p(301)(111),clock=>clock,reset=>reset,s=>p(329)(111),cout=>p(330)(112));
FA_ff_12610:FAff port map(x=>p(299)(112),y=>p(300)(112),Cin=>p(301)(112),clock=>clock,reset=>reset,s=>p(329)(112),cout=>p(330)(113));
FA_ff_12611:FAff port map(x=>p(299)(113),y=>p(300)(113),Cin=>p(301)(113),clock=>clock,reset=>reset,s=>p(329)(113),cout=>p(330)(114));
FA_ff_12612:FAff port map(x=>p(299)(114),y=>p(300)(114),Cin=>p(301)(114),clock=>clock,reset=>reset,s=>p(329)(114),cout=>p(330)(115));
FA_ff_12613:FAff port map(x=>p(299)(115),y=>p(300)(115),Cin=>p(301)(115),clock=>clock,reset=>reset,s=>p(329)(115),cout=>p(330)(116));
FA_ff_12614:FAff port map(x=>p(299)(116),y=>p(300)(116),Cin=>p(301)(116),clock=>clock,reset=>reset,s=>p(329)(116),cout=>p(330)(117));
FA_ff_12615:FAff port map(x=>p(299)(117),y=>p(300)(117),Cin=>p(301)(117),clock=>clock,reset=>reset,s=>p(329)(117),cout=>p(330)(118));
FA_ff_12616:FAff port map(x=>p(299)(118),y=>p(300)(118),Cin=>p(301)(118),clock=>clock,reset=>reset,s=>p(329)(118),cout=>p(330)(119));
FA_ff_12617:FAff port map(x=>p(299)(119),y=>p(300)(119),Cin=>p(301)(119),clock=>clock,reset=>reset,s=>p(329)(119),cout=>p(330)(120));
FA_ff_12618:FAff port map(x=>p(299)(120),y=>p(300)(120),Cin=>p(301)(120),clock=>clock,reset=>reset,s=>p(329)(120),cout=>p(330)(121));
FA_ff_12619:FAff port map(x=>p(299)(121),y=>p(300)(121),Cin=>p(301)(121),clock=>clock,reset=>reset,s=>p(329)(121),cout=>p(330)(122));
FA_ff_12620:FAff port map(x=>p(299)(122),y=>p(300)(122),Cin=>p(301)(122),clock=>clock,reset=>reset,s=>p(329)(122),cout=>p(330)(123));
FA_ff_12621:FAff port map(x=>p(299)(123),y=>p(300)(123),Cin=>p(301)(123),clock=>clock,reset=>reset,s=>p(329)(123),cout=>p(330)(124));
FA_ff_12622:FAff port map(x=>p(299)(124),y=>p(300)(124),Cin=>p(301)(124),clock=>clock,reset=>reset,s=>p(329)(124),cout=>p(330)(125));
FA_ff_12623:FAff port map(x=>p(299)(125),y=>p(300)(125),Cin=>p(301)(125),clock=>clock,reset=>reset,s=>p(329)(125),cout=>p(330)(126));
FA_ff_12624:FAff port map(x=>p(299)(126),y=>p(300)(126),Cin=>p(301)(126),clock=>clock,reset=>reset,s=>p(329)(126),cout=>p(330)(127));
FA_ff_12625:FAff port map(x=>p(299)(127),y=>p(300)(127),Cin=>p(301)(127),clock=>clock,reset=>reset,s=>p(329)(127),cout=>p(330)(128));
FA_ff_12626:FAff port map(x=>p(299)(128),y=>p(300)(128),Cin=>p(301)(128),clock=>clock,reset=>reset,s=>p(329)(128),cout=>p(330)(129));
FA_ff_12627:FAff port map(x=>p(299)(129),y=>p(300)(129),Cin=>p(301)(129),clock=>clock,reset=>reset,s=>p(329)(129),cout=>p(330)(130));
HA_ff_69:HAff port map(x=>p(302)(0),y=>p(304)(0),clock=>clock,reset=>reset,s=>p(331)(0),c=>p(332)(1));
HA_ff_70:HAff port map(x=>p(302)(1),y=>p(304)(1),clock=>clock,reset=>reset,s=>p(331)(1),c=>p(332)(2));
FA_ff_12628:FAff port map(x=>p(302)(2),y=>p(303)(2),Cin=>p(304)(2),clock=>clock,reset=>reset,s=>p(331)(2),cout=>p(332)(3));
FA_ff_12629:FAff port map(x=>p(302)(3),y=>p(303)(3),Cin=>p(304)(3),clock=>clock,reset=>reset,s=>p(331)(3),cout=>p(332)(4));
FA_ff_12630:FAff port map(x=>p(302)(4),y=>p(303)(4),Cin=>p(304)(4),clock=>clock,reset=>reset,s=>p(331)(4),cout=>p(332)(5));
FA_ff_12631:FAff port map(x=>p(302)(5),y=>p(303)(5),Cin=>p(304)(5),clock=>clock,reset=>reset,s=>p(331)(5),cout=>p(332)(6));
FA_ff_12632:FAff port map(x=>p(302)(6),y=>p(303)(6),Cin=>p(304)(6),clock=>clock,reset=>reset,s=>p(331)(6),cout=>p(332)(7));
FA_ff_12633:FAff port map(x=>p(302)(7),y=>p(303)(7),Cin=>p(304)(7),clock=>clock,reset=>reset,s=>p(331)(7),cout=>p(332)(8));
FA_ff_12634:FAff port map(x=>p(302)(8),y=>p(303)(8),Cin=>p(304)(8),clock=>clock,reset=>reset,s=>p(331)(8),cout=>p(332)(9));
FA_ff_12635:FAff port map(x=>p(302)(9),y=>p(303)(9),Cin=>p(304)(9),clock=>clock,reset=>reset,s=>p(331)(9),cout=>p(332)(10));
FA_ff_12636:FAff port map(x=>p(302)(10),y=>p(303)(10),Cin=>p(304)(10),clock=>clock,reset=>reset,s=>p(331)(10),cout=>p(332)(11));
FA_ff_12637:FAff port map(x=>p(302)(11),y=>p(303)(11),Cin=>p(304)(11),clock=>clock,reset=>reset,s=>p(331)(11),cout=>p(332)(12));
FA_ff_12638:FAff port map(x=>p(302)(12),y=>p(303)(12),Cin=>p(304)(12),clock=>clock,reset=>reset,s=>p(331)(12),cout=>p(332)(13));
FA_ff_12639:FAff port map(x=>p(302)(13),y=>p(303)(13),Cin=>p(304)(13),clock=>clock,reset=>reset,s=>p(331)(13),cout=>p(332)(14));
FA_ff_12640:FAff port map(x=>p(302)(14),y=>p(303)(14),Cin=>p(304)(14),clock=>clock,reset=>reset,s=>p(331)(14),cout=>p(332)(15));
FA_ff_12641:FAff port map(x=>p(302)(15),y=>p(303)(15),Cin=>p(304)(15),clock=>clock,reset=>reset,s=>p(331)(15),cout=>p(332)(16));
FA_ff_12642:FAff port map(x=>p(302)(16),y=>p(303)(16),Cin=>p(304)(16),clock=>clock,reset=>reset,s=>p(331)(16),cout=>p(332)(17));
FA_ff_12643:FAff port map(x=>p(302)(17),y=>p(303)(17),Cin=>p(304)(17),clock=>clock,reset=>reset,s=>p(331)(17),cout=>p(332)(18));
FA_ff_12644:FAff port map(x=>p(302)(18),y=>p(303)(18),Cin=>p(304)(18),clock=>clock,reset=>reset,s=>p(331)(18),cout=>p(332)(19));
FA_ff_12645:FAff port map(x=>p(302)(19),y=>p(303)(19),Cin=>p(304)(19),clock=>clock,reset=>reset,s=>p(331)(19),cout=>p(332)(20));
FA_ff_12646:FAff port map(x=>p(302)(20),y=>p(303)(20),Cin=>p(304)(20),clock=>clock,reset=>reset,s=>p(331)(20),cout=>p(332)(21));
FA_ff_12647:FAff port map(x=>p(302)(21),y=>p(303)(21),Cin=>p(304)(21),clock=>clock,reset=>reset,s=>p(331)(21),cout=>p(332)(22));
FA_ff_12648:FAff port map(x=>p(302)(22),y=>p(303)(22),Cin=>p(304)(22),clock=>clock,reset=>reset,s=>p(331)(22),cout=>p(332)(23));
FA_ff_12649:FAff port map(x=>p(302)(23),y=>p(303)(23),Cin=>p(304)(23),clock=>clock,reset=>reset,s=>p(331)(23),cout=>p(332)(24));
FA_ff_12650:FAff port map(x=>p(302)(24),y=>p(303)(24),Cin=>p(304)(24),clock=>clock,reset=>reset,s=>p(331)(24),cout=>p(332)(25));
FA_ff_12651:FAff port map(x=>p(302)(25),y=>p(303)(25),Cin=>p(304)(25),clock=>clock,reset=>reset,s=>p(331)(25),cout=>p(332)(26));
FA_ff_12652:FAff port map(x=>p(302)(26),y=>p(303)(26),Cin=>p(304)(26),clock=>clock,reset=>reset,s=>p(331)(26),cout=>p(332)(27));
FA_ff_12653:FAff port map(x=>p(302)(27),y=>p(303)(27),Cin=>p(304)(27),clock=>clock,reset=>reset,s=>p(331)(27),cout=>p(332)(28));
FA_ff_12654:FAff port map(x=>p(302)(28),y=>p(303)(28),Cin=>p(304)(28),clock=>clock,reset=>reset,s=>p(331)(28),cout=>p(332)(29));
FA_ff_12655:FAff port map(x=>p(302)(29),y=>p(303)(29),Cin=>p(304)(29),clock=>clock,reset=>reset,s=>p(331)(29),cout=>p(332)(30));
FA_ff_12656:FAff port map(x=>p(302)(30),y=>p(303)(30),Cin=>p(304)(30),clock=>clock,reset=>reset,s=>p(331)(30),cout=>p(332)(31));
FA_ff_12657:FAff port map(x=>p(302)(31),y=>p(303)(31),Cin=>p(304)(31),clock=>clock,reset=>reset,s=>p(331)(31),cout=>p(332)(32));
FA_ff_12658:FAff port map(x=>p(302)(32),y=>p(303)(32),Cin=>p(304)(32),clock=>clock,reset=>reset,s=>p(331)(32),cout=>p(332)(33));
FA_ff_12659:FAff port map(x=>p(302)(33),y=>p(303)(33),Cin=>p(304)(33),clock=>clock,reset=>reset,s=>p(331)(33),cout=>p(332)(34));
FA_ff_12660:FAff port map(x=>p(302)(34),y=>p(303)(34),Cin=>p(304)(34),clock=>clock,reset=>reset,s=>p(331)(34),cout=>p(332)(35));
FA_ff_12661:FAff port map(x=>p(302)(35),y=>p(303)(35),Cin=>p(304)(35),clock=>clock,reset=>reset,s=>p(331)(35),cout=>p(332)(36));
FA_ff_12662:FAff port map(x=>p(302)(36),y=>p(303)(36),Cin=>p(304)(36),clock=>clock,reset=>reset,s=>p(331)(36),cout=>p(332)(37));
FA_ff_12663:FAff port map(x=>p(302)(37),y=>p(303)(37),Cin=>p(304)(37),clock=>clock,reset=>reset,s=>p(331)(37),cout=>p(332)(38));
FA_ff_12664:FAff port map(x=>p(302)(38),y=>p(303)(38),Cin=>p(304)(38),clock=>clock,reset=>reset,s=>p(331)(38),cout=>p(332)(39));
FA_ff_12665:FAff port map(x=>p(302)(39),y=>p(303)(39),Cin=>p(304)(39),clock=>clock,reset=>reset,s=>p(331)(39),cout=>p(332)(40));
FA_ff_12666:FAff port map(x=>p(302)(40),y=>p(303)(40),Cin=>p(304)(40),clock=>clock,reset=>reset,s=>p(331)(40),cout=>p(332)(41));
FA_ff_12667:FAff port map(x=>p(302)(41),y=>p(303)(41),Cin=>p(304)(41),clock=>clock,reset=>reset,s=>p(331)(41),cout=>p(332)(42));
FA_ff_12668:FAff port map(x=>p(302)(42),y=>p(303)(42),Cin=>p(304)(42),clock=>clock,reset=>reset,s=>p(331)(42),cout=>p(332)(43));
FA_ff_12669:FAff port map(x=>p(302)(43),y=>p(303)(43),Cin=>p(304)(43),clock=>clock,reset=>reset,s=>p(331)(43),cout=>p(332)(44));
FA_ff_12670:FAff port map(x=>p(302)(44),y=>p(303)(44),Cin=>p(304)(44),clock=>clock,reset=>reset,s=>p(331)(44),cout=>p(332)(45));
FA_ff_12671:FAff port map(x=>p(302)(45),y=>p(303)(45),Cin=>p(304)(45),clock=>clock,reset=>reset,s=>p(331)(45),cout=>p(332)(46));
FA_ff_12672:FAff port map(x=>p(302)(46),y=>p(303)(46),Cin=>p(304)(46),clock=>clock,reset=>reset,s=>p(331)(46),cout=>p(332)(47));
FA_ff_12673:FAff port map(x=>p(302)(47),y=>p(303)(47),Cin=>p(304)(47),clock=>clock,reset=>reset,s=>p(331)(47),cout=>p(332)(48));
FA_ff_12674:FAff port map(x=>p(302)(48),y=>p(303)(48),Cin=>p(304)(48),clock=>clock,reset=>reset,s=>p(331)(48),cout=>p(332)(49));
FA_ff_12675:FAff port map(x=>p(302)(49),y=>p(303)(49),Cin=>p(304)(49),clock=>clock,reset=>reset,s=>p(331)(49),cout=>p(332)(50));
FA_ff_12676:FAff port map(x=>p(302)(50),y=>p(303)(50),Cin=>p(304)(50),clock=>clock,reset=>reset,s=>p(331)(50),cout=>p(332)(51));
FA_ff_12677:FAff port map(x=>p(302)(51),y=>p(303)(51),Cin=>p(304)(51),clock=>clock,reset=>reset,s=>p(331)(51),cout=>p(332)(52));
FA_ff_12678:FAff port map(x=>p(302)(52),y=>p(303)(52),Cin=>p(304)(52),clock=>clock,reset=>reset,s=>p(331)(52),cout=>p(332)(53));
FA_ff_12679:FAff port map(x=>p(302)(53),y=>p(303)(53),Cin=>p(304)(53),clock=>clock,reset=>reset,s=>p(331)(53),cout=>p(332)(54));
FA_ff_12680:FAff port map(x=>p(302)(54),y=>p(303)(54),Cin=>p(304)(54),clock=>clock,reset=>reset,s=>p(331)(54),cout=>p(332)(55));
FA_ff_12681:FAff port map(x=>p(302)(55),y=>p(303)(55),Cin=>p(304)(55),clock=>clock,reset=>reset,s=>p(331)(55),cout=>p(332)(56));
FA_ff_12682:FAff port map(x=>p(302)(56),y=>p(303)(56),Cin=>p(304)(56),clock=>clock,reset=>reset,s=>p(331)(56),cout=>p(332)(57));
FA_ff_12683:FAff port map(x=>p(302)(57),y=>p(303)(57),Cin=>p(304)(57),clock=>clock,reset=>reset,s=>p(331)(57),cout=>p(332)(58));
FA_ff_12684:FAff port map(x=>p(302)(58),y=>p(303)(58),Cin=>p(304)(58),clock=>clock,reset=>reset,s=>p(331)(58),cout=>p(332)(59));
FA_ff_12685:FAff port map(x=>p(302)(59),y=>p(303)(59),Cin=>p(304)(59),clock=>clock,reset=>reset,s=>p(331)(59),cout=>p(332)(60));
FA_ff_12686:FAff port map(x=>p(302)(60),y=>p(303)(60),Cin=>p(304)(60),clock=>clock,reset=>reset,s=>p(331)(60),cout=>p(332)(61));
FA_ff_12687:FAff port map(x=>p(302)(61),y=>p(303)(61),Cin=>p(304)(61),clock=>clock,reset=>reset,s=>p(331)(61),cout=>p(332)(62));
FA_ff_12688:FAff port map(x=>p(302)(62),y=>p(303)(62),Cin=>p(304)(62),clock=>clock,reset=>reset,s=>p(331)(62),cout=>p(332)(63));
FA_ff_12689:FAff port map(x=>p(302)(63),y=>p(303)(63),Cin=>p(304)(63),clock=>clock,reset=>reset,s=>p(331)(63),cout=>p(332)(64));
FA_ff_12690:FAff port map(x=>p(302)(64),y=>p(303)(64),Cin=>p(304)(64),clock=>clock,reset=>reset,s=>p(331)(64),cout=>p(332)(65));
FA_ff_12691:FAff port map(x=>p(302)(65),y=>p(303)(65),Cin=>p(304)(65),clock=>clock,reset=>reset,s=>p(331)(65),cout=>p(332)(66));
FA_ff_12692:FAff port map(x=>p(302)(66),y=>p(303)(66),Cin=>p(304)(66),clock=>clock,reset=>reset,s=>p(331)(66),cout=>p(332)(67));
FA_ff_12693:FAff port map(x=>p(302)(67),y=>p(303)(67),Cin=>p(304)(67),clock=>clock,reset=>reset,s=>p(331)(67),cout=>p(332)(68));
FA_ff_12694:FAff port map(x=>p(302)(68),y=>p(303)(68),Cin=>p(304)(68),clock=>clock,reset=>reset,s=>p(331)(68),cout=>p(332)(69));
FA_ff_12695:FAff port map(x=>p(302)(69),y=>p(303)(69),Cin=>p(304)(69),clock=>clock,reset=>reset,s=>p(331)(69),cout=>p(332)(70));
FA_ff_12696:FAff port map(x=>p(302)(70),y=>p(303)(70),Cin=>p(304)(70),clock=>clock,reset=>reset,s=>p(331)(70),cout=>p(332)(71));
FA_ff_12697:FAff port map(x=>p(302)(71),y=>p(303)(71),Cin=>p(304)(71),clock=>clock,reset=>reset,s=>p(331)(71),cout=>p(332)(72));
FA_ff_12698:FAff port map(x=>p(302)(72),y=>p(303)(72),Cin=>p(304)(72),clock=>clock,reset=>reset,s=>p(331)(72),cout=>p(332)(73));
FA_ff_12699:FAff port map(x=>p(302)(73),y=>p(303)(73),Cin=>p(304)(73),clock=>clock,reset=>reset,s=>p(331)(73),cout=>p(332)(74));
FA_ff_12700:FAff port map(x=>p(302)(74),y=>p(303)(74),Cin=>p(304)(74),clock=>clock,reset=>reset,s=>p(331)(74),cout=>p(332)(75));
FA_ff_12701:FAff port map(x=>p(302)(75),y=>p(303)(75),Cin=>p(304)(75),clock=>clock,reset=>reset,s=>p(331)(75),cout=>p(332)(76));
FA_ff_12702:FAff port map(x=>p(302)(76),y=>p(303)(76),Cin=>p(304)(76),clock=>clock,reset=>reset,s=>p(331)(76),cout=>p(332)(77));
FA_ff_12703:FAff port map(x=>p(302)(77),y=>p(303)(77),Cin=>p(304)(77),clock=>clock,reset=>reset,s=>p(331)(77),cout=>p(332)(78));
FA_ff_12704:FAff port map(x=>p(302)(78),y=>p(303)(78),Cin=>p(304)(78),clock=>clock,reset=>reset,s=>p(331)(78),cout=>p(332)(79));
FA_ff_12705:FAff port map(x=>p(302)(79),y=>p(303)(79),Cin=>p(304)(79),clock=>clock,reset=>reset,s=>p(331)(79),cout=>p(332)(80));
FA_ff_12706:FAff port map(x=>p(302)(80),y=>p(303)(80),Cin=>p(304)(80),clock=>clock,reset=>reset,s=>p(331)(80),cout=>p(332)(81));
FA_ff_12707:FAff port map(x=>p(302)(81),y=>p(303)(81),Cin=>p(304)(81),clock=>clock,reset=>reset,s=>p(331)(81),cout=>p(332)(82));
FA_ff_12708:FAff port map(x=>p(302)(82),y=>p(303)(82),Cin=>p(304)(82),clock=>clock,reset=>reset,s=>p(331)(82),cout=>p(332)(83));
FA_ff_12709:FAff port map(x=>p(302)(83),y=>p(303)(83),Cin=>p(304)(83),clock=>clock,reset=>reset,s=>p(331)(83),cout=>p(332)(84));
FA_ff_12710:FAff port map(x=>p(302)(84),y=>p(303)(84),Cin=>p(304)(84),clock=>clock,reset=>reset,s=>p(331)(84),cout=>p(332)(85));
FA_ff_12711:FAff port map(x=>p(302)(85),y=>p(303)(85),Cin=>p(304)(85),clock=>clock,reset=>reset,s=>p(331)(85),cout=>p(332)(86));
FA_ff_12712:FAff port map(x=>p(302)(86),y=>p(303)(86),Cin=>p(304)(86),clock=>clock,reset=>reset,s=>p(331)(86),cout=>p(332)(87));
FA_ff_12713:FAff port map(x=>p(302)(87),y=>p(303)(87),Cin=>p(304)(87),clock=>clock,reset=>reset,s=>p(331)(87),cout=>p(332)(88));
FA_ff_12714:FAff port map(x=>p(302)(88),y=>p(303)(88),Cin=>p(304)(88),clock=>clock,reset=>reset,s=>p(331)(88),cout=>p(332)(89));
FA_ff_12715:FAff port map(x=>p(302)(89),y=>p(303)(89),Cin=>p(304)(89),clock=>clock,reset=>reset,s=>p(331)(89),cout=>p(332)(90));
FA_ff_12716:FAff port map(x=>p(302)(90),y=>p(303)(90),Cin=>p(304)(90),clock=>clock,reset=>reset,s=>p(331)(90),cout=>p(332)(91));
FA_ff_12717:FAff port map(x=>p(302)(91),y=>p(303)(91),Cin=>p(304)(91),clock=>clock,reset=>reset,s=>p(331)(91),cout=>p(332)(92));
FA_ff_12718:FAff port map(x=>p(302)(92),y=>p(303)(92),Cin=>p(304)(92),clock=>clock,reset=>reset,s=>p(331)(92),cout=>p(332)(93));
FA_ff_12719:FAff port map(x=>p(302)(93),y=>p(303)(93),Cin=>p(304)(93),clock=>clock,reset=>reset,s=>p(331)(93),cout=>p(332)(94));
FA_ff_12720:FAff port map(x=>p(302)(94),y=>p(303)(94),Cin=>p(304)(94),clock=>clock,reset=>reset,s=>p(331)(94),cout=>p(332)(95));
FA_ff_12721:FAff port map(x=>p(302)(95),y=>p(303)(95),Cin=>p(304)(95),clock=>clock,reset=>reset,s=>p(331)(95),cout=>p(332)(96));
FA_ff_12722:FAff port map(x=>p(302)(96),y=>p(303)(96),Cin=>p(304)(96),clock=>clock,reset=>reset,s=>p(331)(96),cout=>p(332)(97));
FA_ff_12723:FAff port map(x=>p(302)(97),y=>p(303)(97),Cin=>p(304)(97),clock=>clock,reset=>reset,s=>p(331)(97),cout=>p(332)(98));
FA_ff_12724:FAff port map(x=>p(302)(98),y=>p(303)(98),Cin=>p(304)(98),clock=>clock,reset=>reset,s=>p(331)(98),cout=>p(332)(99));
FA_ff_12725:FAff port map(x=>p(302)(99),y=>p(303)(99),Cin=>p(304)(99),clock=>clock,reset=>reset,s=>p(331)(99),cout=>p(332)(100));
FA_ff_12726:FAff port map(x=>p(302)(100),y=>p(303)(100),Cin=>p(304)(100),clock=>clock,reset=>reset,s=>p(331)(100),cout=>p(332)(101));
FA_ff_12727:FAff port map(x=>p(302)(101),y=>p(303)(101),Cin=>p(304)(101),clock=>clock,reset=>reset,s=>p(331)(101),cout=>p(332)(102));
FA_ff_12728:FAff port map(x=>p(302)(102),y=>p(303)(102),Cin=>p(304)(102),clock=>clock,reset=>reset,s=>p(331)(102),cout=>p(332)(103));
FA_ff_12729:FAff port map(x=>p(302)(103),y=>p(303)(103),Cin=>p(304)(103),clock=>clock,reset=>reset,s=>p(331)(103),cout=>p(332)(104));
FA_ff_12730:FAff port map(x=>p(302)(104),y=>p(303)(104),Cin=>p(304)(104),clock=>clock,reset=>reset,s=>p(331)(104),cout=>p(332)(105));
FA_ff_12731:FAff port map(x=>p(302)(105),y=>p(303)(105),Cin=>p(304)(105),clock=>clock,reset=>reset,s=>p(331)(105),cout=>p(332)(106));
FA_ff_12732:FAff port map(x=>p(302)(106),y=>p(303)(106),Cin=>p(304)(106),clock=>clock,reset=>reset,s=>p(331)(106),cout=>p(332)(107));
FA_ff_12733:FAff port map(x=>p(302)(107),y=>p(303)(107),Cin=>p(304)(107),clock=>clock,reset=>reset,s=>p(331)(107),cout=>p(332)(108));
FA_ff_12734:FAff port map(x=>p(302)(108),y=>p(303)(108),Cin=>p(304)(108),clock=>clock,reset=>reset,s=>p(331)(108),cout=>p(332)(109));
FA_ff_12735:FAff port map(x=>p(302)(109),y=>p(303)(109),Cin=>p(304)(109),clock=>clock,reset=>reset,s=>p(331)(109),cout=>p(332)(110));
FA_ff_12736:FAff port map(x=>p(302)(110),y=>p(303)(110),Cin=>p(304)(110),clock=>clock,reset=>reset,s=>p(331)(110),cout=>p(332)(111));
FA_ff_12737:FAff port map(x=>p(302)(111),y=>p(303)(111),Cin=>p(304)(111),clock=>clock,reset=>reset,s=>p(331)(111),cout=>p(332)(112));
FA_ff_12738:FAff port map(x=>p(302)(112),y=>p(303)(112),Cin=>p(304)(112),clock=>clock,reset=>reset,s=>p(331)(112),cout=>p(332)(113));
FA_ff_12739:FAff port map(x=>p(302)(113),y=>p(303)(113),Cin=>p(304)(113),clock=>clock,reset=>reset,s=>p(331)(113),cout=>p(332)(114));
FA_ff_12740:FAff port map(x=>p(302)(114),y=>p(303)(114),Cin=>p(304)(114),clock=>clock,reset=>reset,s=>p(331)(114),cout=>p(332)(115));
FA_ff_12741:FAff port map(x=>p(302)(115),y=>p(303)(115),Cin=>p(304)(115),clock=>clock,reset=>reset,s=>p(331)(115),cout=>p(332)(116));
FA_ff_12742:FAff port map(x=>p(302)(116),y=>p(303)(116),Cin=>p(304)(116),clock=>clock,reset=>reset,s=>p(331)(116),cout=>p(332)(117));
FA_ff_12743:FAff port map(x=>p(302)(117),y=>p(303)(117),Cin=>p(304)(117),clock=>clock,reset=>reset,s=>p(331)(117),cout=>p(332)(118));
FA_ff_12744:FAff port map(x=>p(302)(118),y=>p(303)(118),Cin=>p(304)(118),clock=>clock,reset=>reset,s=>p(331)(118),cout=>p(332)(119));
FA_ff_12745:FAff port map(x=>p(302)(119),y=>p(303)(119),Cin=>p(304)(119),clock=>clock,reset=>reset,s=>p(331)(119),cout=>p(332)(120));
FA_ff_12746:FAff port map(x=>p(302)(120),y=>p(303)(120),Cin=>p(304)(120),clock=>clock,reset=>reset,s=>p(331)(120),cout=>p(332)(121));
FA_ff_12747:FAff port map(x=>p(302)(121),y=>p(303)(121),Cin=>p(304)(121),clock=>clock,reset=>reset,s=>p(331)(121),cout=>p(332)(122));
FA_ff_12748:FAff port map(x=>p(302)(122),y=>p(303)(122),Cin=>p(304)(122),clock=>clock,reset=>reset,s=>p(331)(122),cout=>p(332)(123));
FA_ff_12749:FAff port map(x=>p(302)(123),y=>p(303)(123),Cin=>p(304)(123),clock=>clock,reset=>reset,s=>p(331)(123),cout=>p(332)(124));
FA_ff_12750:FAff port map(x=>p(302)(124),y=>p(303)(124),Cin=>p(304)(124),clock=>clock,reset=>reset,s=>p(331)(124),cout=>p(332)(125));
FA_ff_12751:FAff port map(x=>p(302)(125),y=>p(303)(125),Cin=>p(304)(125),clock=>clock,reset=>reset,s=>p(331)(125),cout=>p(332)(126));
FA_ff_12752:FAff port map(x=>p(302)(126),y=>p(303)(126),Cin=>p(304)(126),clock=>clock,reset=>reset,s=>p(331)(126),cout=>p(332)(127));
FA_ff_12753:FAff port map(x=>p(302)(127),y=>p(303)(127),Cin=>p(304)(127),clock=>clock,reset=>reset,s=>p(331)(127),cout=>p(332)(128));
FA_ff_12754:FAff port map(x=>p(302)(128),y=>p(303)(128),Cin=>p(304)(128),clock=>clock,reset=>reset,s=>p(331)(128),cout=>p(332)(129));
HA_ff_71:HAff port map(x=>p(302)(129),y=>p(303)(129),clock=>clock,reset=>reset,s=>p(331)(129),c=>p(332)(130));
p(333)(0)<=p(306)(0);
HA_ff_72:HAff port map(x=>p(305)(1),y=>p(306)(1),clock=>clock,reset=>reset,s=>p(333)(1),c=>p(334)(2));
FA_ff_12755:FAff port map(x=>p(305)(2),y=>p(306)(2),Cin=>p(307)(2),clock=>clock,reset=>reset,s=>p(333)(2),cout=>p(334)(3));
FA_ff_12756:FAff port map(x=>p(305)(3),y=>p(306)(3),Cin=>p(307)(3),clock=>clock,reset=>reset,s=>p(333)(3),cout=>p(334)(4));
FA_ff_12757:FAff port map(x=>p(305)(4),y=>p(306)(4),Cin=>p(307)(4),clock=>clock,reset=>reset,s=>p(333)(4),cout=>p(334)(5));
FA_ff_12758:FAff port map(x=>p(305)(5),y=>p(306)(5),Cin=>p(307)(5),clock=>clock,reset=>reset,s=>p(333)(5),cout=>p(334)(6));
FA_ff_12759:FAff port map(x=>p(305)(6),y=>p(306)(6),Cin=>p(307)(6),clock=>clock,reset=>reset,s=>p(333)(6),cout=>p(334)(7));
FA_ff_12760:FAff port map(x=>p(305)(7),y=>p(306)(7),Cin=>p(307)(7),clock=>clock,reset=>reset,s=>p(333)(7),cout=>p(334)(8));
FA_ff_12761:FAff port map(x=>p(305)(8),y=>p(306)(8),Cin=>p(307)(8),clock=>clock,reset=>reset,s=>p(333)(8),cout=>p(334)(9));
FA_ff_12762:FAff port map(x=>p(305)(9),y=>p(306)(9),Cin=>p(307)(9),clock=>clock,reset=>reset,s=>p(333)(9),cout=>p(334)(10));
FA_ff_12763:FAff port map(x=>p(305)(10),y=>p(306)(10),Cin=>p(307)(10),clock=>clock,reset=>reset,s=>p(333)(10),cout=>p(334)(11));
FA_ff_12764:FAff port map(x=>p(305)(11),y=>p(306)(11),Cin=>p(307)(11),clock=>clock,reset=>reset,s=>p(333)(11),cout=>p(334)(12));
FA_ff_12765:FAff port map(x=>p(305)(12),y=>p(306)(12),Cin=>p(307)(12),clock=>clock,reset=>reset,s=>p(333)(12),cout=>p(334)(13));
FA_ff_12766:FAff port map(x=>p(305)(13),y=>p(306)(13),Cin=>p(307)(13),clock=>clock,reset=>reset,s=>p(333)(13),cout=>p(334)(14));
FA_ff_12767:FAff port map(x=>p(305)(14),y=>p(306)(14),Cin=>p(307)(14),clock=>clock,reset=>reset,s=>p(333)(14),cout=>p(334)(15));
FA_ff_12768:FAff port map(x=>p(305)(15),y=>p(306)(15),Cin=>p(307)(15),clock=>clock,reset=>reset,s=>p(333)(15),cout=>p(334)(16));
FA_ff_12769:FAff port map(x=>p(305)(16),y=>p(306)(16),Cin=>p(307)(16),clock=>clock,reset=>reset,s=>p(333)(16),cout=>p(334)(17));
FA_ff_12770:FAff port map(x=>p(305)(17),y=>p(306)(17),Cin=>p(307)(17),clock=>clock,reset=>reset,s=>p(333)(17),cout=>p(334)(18));
FA_ff_12771:FAff port map(x=>p(305)(18),y=>p(306)(18),Cin=>p(307)(18),clock=>clock,reset=>reset,s=>p(333)(18),cout=>p(334)(19));
FA_ff_12772:FAff port map(x=>p(305)(19),y=>p(306)(19),Cin=>p(307)(19),clock=>clock,reset=>reset,s=>p(333)(19),cout=>p(334)(20));
FA_ff_12773:FAff port map(x=>p(305)(20),y=>p(306)(20),Cin=>p(307)(20),clock=>clock,reset=>reset,s=>p(333)(20),cout=>p(334)(21));
FA_ff_12774:FAff port map(x=>p(305)(21),y=>p(306)(21),Cin=>p(307)(21),clock=>clock,reset=>reset,s=>p(333)(21),cout=>p(334)(22));
FA_ff_12775:FAff port map(x=>p(305)(22),y=>p(306)(22),Cin=>p(307)(22),clock=>clock,reset=>reset,s=>p(333)(22),cout=>p(334)(23));
FA_ff_12776:FAff port map(x=>p(305)(23),y=>p(306)(23),Cin=>p(307)(23),clock=>clock,reset=>reset,s=>p(333)(23),cout=>p(334)(24));
FA_ff_12777:FAff port map(x=>p(305)(24),y=>p(306)(24),Cin=>p(307)(24),clock=>clock,reset=>reset,s=>p(333)(24),cout=>p(334)(25));
FA_ff_12778:FAff port map(x=>p(305)(25),y=>p(306)(25),Cin=>p(307)(25),clock=>clock,reset=>reset,s=>p(333)(25),cout=>p(334)(26));
FA_ff_12779:FAff port map(x=>p(305)(26),y=>p(306)(26),Cin=>p(307)(26),clock=>clock,reset=>reset,s=>p(333)(26),cout=>p(334)(27));
FA_ff_12780:FAff port map(x=>p(305)(27),y=>p(306)(27),Cin=>p(307)(27),clock=>clock,reset=>reset,s=>p(333)(27),cout=>p(334)(28));
FA_ff_12781:FAff port map(x=>p(305)(28),y=>p(306)(28),Cin=>p(307)(28),clock=>clock,reset=>reset,s=>p(333)(28),cout=>p(334)(29));
FA_ff_12782:FAff port map(x=>p(305)(29),y=>p(306)(29),Cin=>p(307)(29),clock=>clock,reset=>reset,s=>p(333)(29),cout=>p(334)(30));
FA_ff_12783:FAff port map(x=>p(305)(30),y=>p(306)(30),Cin=>p(307)(30),clock=>clock,reset=>reset,s=>p(333)(30),cout=>p(334)(31));
FA_ff_12784:FAff port map(x=>p(305)(31),y=>p(306)(31),Cin=>p(307)(31),clock=>clock,reset=>reset,s=>p(333)(31),cout=>p(334)(32));
FA_ff_12785:FAff port map(x=>p(305)(32),y=>p(306)(32),Cin=>p(307)(32),clock=>clock,reset=>reset,s=>p(333)(32),cout=>p(334)(33));
FA_ff_12786:FAff port map(x=>p(305)(33),y=>p(306)(33),Cin=>p(307)(33),clock=>clock,reset=>reset,s=>p(333)(33),cout=>p(334)(34));
FA_ff_12787:FAff port map(x=>p(305)(34),y=>p(306)(34),Cin=>p(307)(34),clock=>clock,reset=>reset,s=>p(333)(34),cout=>p(334)(35));
FA_ff_12788:FAff port map(x=>p(305)(35),y=>p(306)(35),Cin=>p(307)(35),clock=>clock,reset=>reset,s=>p(333)(35),cout=>p(334)(36));
FA_ff_12789:FAff port map(x=>p(305)(36),y=>p(306)(36),Cin=>p(307)(36),clock=>clock,reset=>reset,s=>p(333)(36),cout=>p(334)(37));
FA_ff_12790:FAff port map(x=>p(305)(37),y=>p(306)(37),Cin=>p(307)(37),clock=>clock,reset=>reset,s=>p(333)(37),cout=>p(334)(38));
FA_ff_12791:FAff port map(x=>p(305)(38),y=>p(306)(38),Cin=>p(307)(38),clock=>clock,reset=>reset,s=>p(333)(38),cout=>p(334)(39));
FA_ff_12792:FAff port map(x=>p(305)(39),y=>p(306)(39),Cin=>p(307)(39),clock=>clock,reset=>reset,s=>p(333)(39),cout=>p(334)(40));
FA_ff_12793:FAff port map(x=>p(305)(40),y=>p(306)(40),Cin=>p(307)(40),clock=>clock,reset=>reset,s=>p(333)(40),cout=>p(334)(41));
FA_ff_12794:FAff port map(x=>p(305)(41),y=>p(306)(41),Cin=>p(307)(41),clock=>clock,reset=>reset,s=>p(333)(41),cout=>p(334)(42));
FA_ff_12795:FAff port map(x=>p(305)(42),y=>p(306)(42),Cin=>p(307)(42),clock=>clock,reset=>reset,s=>p(333)(42),cout=>p(334)(43));
FA_ff_12796:FAff port map(x=>p(305)(43),y=>p(306)(43),Cin=>p(307)(43),clock=>clock,reset=>reset,s=>p(333)(43),cout=>p(334)(44));
FA_ff_12797:FAff port map(x=>p(305)(44),y=>p(306)(44),Cin=>p(307)(44),clock=>clock,reset=>reset,s=>p(333)(44),cout=>p(334)(45));
FA_ff_12798:FAff port map(x=>p(305)(45),y=>p(306)(45),Cin=>p(307)(45),clock=>clock,reset=>reset,s=>p(333)(45),cout=>p(334)(46));
FA_ff_12799:FAff port map(x=>p(305)(46),y=>p(306)(46),Cin=>p(307)(46),clock=>clock,reset=>reset,s=>p(333)(46),cout=>p(334)(47));
FA_ff_12800:FAff port map(x=>p(305)(47),y=>p(306)(47),Cin=>p(307)(47),clock=>clock,reset=>reset,s=>p(333)(47),cout=>p(334)(48));
FA_ff_12801:FAff port map(x=>p(305)(48),y=>p(306)(48),Cin=>p(307)(48),clock=>clock,reset=>reset,s=>p(333)(48),cout=>p(334)(49));
FA_ff_12802:FAff port map(x=>p(305)(49),y=>p(306)(49),Cin=>p(307)(49),clock=>clock,reset=>reset,s=>p(333)(49),cout=>p(334)(50));
FA_ff_12803:FAff port map(x=>p(305)(50),y=>p(306)(50),Cin=>p(307)(50),clock=>clock,reset=>reset,s=>p(333)(50),cout=>p(334)(51));
FA_ff_12804:FAff port map(x=>p(305)(51),y=>p(306)(51),Cin=>p(307)(51),clock=>clock,reset=>reset,s=>p(333)(51),cout=>p(334)(52));
FA_ff_12805:FAff port map(x=>p(305)(52),y=>p(306)(52),Cin=>p(307)(52),clock=>clock,reset=>reset,s=>p(333)(52),cout=>p(334)(53));
FA_ff_12806:FAff port map(x=>p(305)(53),y=>p(306)(53),Cin=>p(307)(53),clock=>clock,reset=>reset,s=>p(333)(53),cout=>p(334)(54));
FA_ff_12807:FAff port map(x=>p(305)(54),y=>p(306)(54),Cin=>p(307)(54),clock=>clock,reset=>reset,s=>p(333)(54),cout=>p(334)(55));
FA_ff_12808:FAff port map(x=>p(305)(55),y=>p(306)(55),Cin=>p(307)(55),clock=>clock,reset=>reset,s=>p(333)(55),cout=>p(334)(56));
FA_ff_12809:FAff port map(x=>p(305)(56),y=>p(306)(56),Cin=>p(307)(56),clock=>clock,reset=>reset,s=>p(333)(56),cout=>p(334)(57));
FA_ff_12810:FAff port map(x=>p(305)(57),y=>p(306)(57),Cin=>p(307)(57),clock=>clock,reset=>reset,s=>p(333)(57),cout=>p(334)(58));
FA_ff_12811:FAff port map(x=>p(305)(58),y=>p(306)(58),Cin=>p(307)(58),clock=>clock,reset=>reset,s=>p(333)(58),cout=>p(334)(59));
FA_ff_12812:FAff port map(x=>p(305)(59),y=>p(306)(59),Cin=>p(307)(59),clock=>clock,reset=>reset,s=>p(333)(59),cout=>p(334)(60));
FA_ff_12813:FAff port map(x=>p(305)(60),y=>p(306)(60),Cin=>p(307)(60),clock=>clock,reset=>reset,s=>p(333)(60),cout=>p(334)(61));
FA_ff_12814:FAff port map(x=>p(305)(61),y=>p(306)(61),Cin=>p(307)(61),clock=>clock,reset=>reset,s=>p(333)(61),cout=>p(334)(62));
FA_ff_12815:FAff port map(x=>p(305)(62),y=>p(306)(62),Cin=>p(307)(62),clock=>clock,reset=>reset,s=>p(333)(62),cout=>p(334)(63));
FA_ff_12816:FAff port map(x=>p(305)(63),y=>p(306)(63),Cin=>p(307)(63),clock=>clock,reset=>reset,s=>p(333)(63),cout=>p(334)(64));
FA_ff_12817:FAff port map(x=>p(305)(64),y=>p(306)(64),Cin=>p(307)(64),clock=>clock,reset=>reset,s=>p(333)(64),cout=>p(334)(65));
FA_ff_12818:FAff port map(x=>p(305)(65),y=>p(306)(65),Cin=>p(307)(65),clock=>clock,reset=>reset,s=>p(333)(65),cout=>p(334)(66));
FA_ff_12819:FAff port map(x=>p(305)(66),y=>p(306)(66),Cin=>p(307)(66),clock=>clock,reset=>reset,s=>p(333)(66),cout=>p(334)(67));
FA_ff_12820:FAff port map(x=>p(305)(67),y=>p(306)(67),Cin=>p(307)(67),clock=>clock,reset=>reset,s=>p(333)(67),cout=>p(334)(68));
FA_ff_12821:FAff port map(x=>p(305)(68),y=>p(306)(68),Cin=>p(307)(68),clock=>clock,reset=>reset,s=>p(333)(68),cout=>p(334)(69));
FA_ff_12822:FAff port map(x=>p(305)(69),y=>p(306)(69),Cin=>p(307)(69),clock=>clock,reset=>reset,s=>p(333)(69),cout=>p(334)(70));
FA_ff_12823:FAff port map(x=>p(305)(70),y=>p(306)(70),Cin=>p(307)(70),clock=>clock,reset=>reset,s=>p(333)(70),cout=>p(334)(71));
FA_ff_12824:FAff port map(x=>p(305)(71),y=>p(306)(71),Cin=>p(307)(71),clock=>clock,reset=>reset,s=>p(333)(71),cout=>p(334)(72));
FA_ff_12825:FAff port map(x=>p(305)(72),y=>p(306)(72),Cin=>p(307)(72),clock=>clock,reset=>reset,s=>p(333)(72),cout=>p(334)(73));
FA_ff_12826:FAff port map(x=>p(305)(73),y=>p(306)(73),Cin=>p(307)(73),clock=>clock,reset=>reset,s=>p(333)(73),cout=>p(334)(74));
FA_ff_12827:FAff port map(x=>p(305)(74),y=>p(306)(74),Cin=>p(307)(74),clock=>clock,reset=>reset,s=>p(333)(74),cout=>p(334)(75));
FA_ff_12828:FAff port map(x=>p(305)(75),y=>p(306)(75),Cin=>p(307)(75),clock=>clock,reset=>reset,s=>p(333)(75),cout=>p(334)(76));
FA_ff_12829:FAff port map(x=>p(305)(76),y=>p(306)(76),Cin=>p(307)(76),clock=>clock,reset=>reset,s=>p(333)(76),cout=>p(334)(77));
FA_ff_12830:FAff port map(x=>p(305)(77),y=>p(306)(77),Cin=>p(307)(77),clock=>clock,reset=>reset,s=>p(333)(77),cout=>p(334)(78));
FA_ff_12831:FAff port map(x=>p(305)(78),y=>p(306)(78),Cin=>p(307)(78),clock=>clock,reset=>reset,s=>p(333)(78),cout=>p(334)(79));
FA_ff_12832:FAff port map(x=>p(305)(79),y=>p(306)(79),Cin=>p(307)(79),clock=>clock,reset=>reset,s=>p(333)(79),cout=>p(334)(80));
FA_ff_12833:FAff port map(x=>p(305)(80),y=>p(306)(80),Cin=>p(307)(80),clock=>clock,reset=>reset,s=>p(333)(80),cout=>p(334)(81));
FA_ff_12834:FAff port map(x=>p(305)(81),y=>p(306)(81),Cin=>p(307)(81),clock=>clock,reset=>reset,s=>p(333)(81),cout=>p(334)(82));
FA_ff_12835:FAff port map(x=>p(305)(82),y=>p(306)(82),Cin=>p(307)(82),clock=>clock,reset=>reset,s=>p(333)(82),cout=>p(334)(83));
FA_ff_12836:FAff port map(x=>p(305)(83),y=>p(306)(83),Cin=>p(307)(83),clock=>clock,reset=>reset,s=>p(333)(83),cout=>p(334)(84));
FA_ff_12837:FAff port map(x=>p(305)(84),y=>p(306)(84),Cin=>p(307)(84),clock=>clock,reset=>reset,s=>p(333)(84),cout=>p(334)(85));
FA_ff_12838:FAff port map(x=>p(305)(85),y=>p(306)(85),Cin=>p(307)(85),clock=>clock,reset=>reset,s=>p(333)(85),cout=>p(334)(86));
FA_ff_12839:FAff port map(x=>p(305)(86),y=>p(306)(86),Cin=>p(307)(86),clock=>clock,reset=>reset,s=>p(333)(86),cout=>p(334)(87));
FA_ff_12840:FAff port map(x=>p(305)(87),y=>p(306)(87),Cin=>p(307)(87),clock=>clock,reset=>reset,s=>p(333)(87),cout=>p(334)(88));
FA_ff_12841:FAff port map(x=>p(305)(88),y=>p(306)(88),Cin=>p(307)(88),clock=>clock,reset=>reset,s=>p(333)(88),cout=>p(334)(89));
FA_ff_12842:FAff port map(x=>p(305)(89),y=>p(306)(89),Cin=>p(307)(89),clock=>clock,reset=>reset,s=>p(333)(89),cout=>p(334)(90));
FA_ff_12843:FAff port map(x=>p(305)(90),y=>p(306)(90),Cin=>p(307)(90),clock=>clock,reset=>reset,s=>p(333)(90),cout=>p(334)(91));
FA_ff_12844:FAff port map(x=>p(305)(91),y=>p(306)(91),Cin=>p(307)(91),clock=>clock,reset=>reset,s=>p(333)(91),cout=>p(334)(92));
FA_ff_12845:FAff port map(x=>p(305)(92),y=>p(306)(92),Cin=>p(307)(92),clock=>clock,reset=>reset,s=>p(333)(92),cout=>p(334)(93));
FA_ff_12846:FAff port map(x=>p(305)(93),y=>p(306)(93),Cin=>p(307)(93),clock=>clock,reset=>reset,s=>p(333)(93),cout=>p(334)(94));
FA_ff_12847:FAff port map(x=>p(305)(94),y=>p(306)(94),Cin=>p(307)(94),clock=>clock,reset=>reset,s=>p(333)(94),cout=>p(334)(95));
FA_ff_12848:FAff port map(x=>p(305)(95),y=>p(306)(95),Cin=>p(307)(95),clock=>clock,reset=>reset,s=>p(333)(95),cout=>p(334)(96));
FA_ff_12849:FAff port map(x=>p(305)(96),y=>p(306)(96),Cin=>p(307)(96),clock=>clock,reset=>reset,s=>p(333)(96),cout=>p(334)(97));
FA_ff_12850:FAff port map(x=>p(305)(97),y=>p(306)(97),Cin=>p(307)(97),clock=>clock,reset=>reset,s=>p(333)(97),cout=>p(334)(98));
FA_ff_12851:FAff port map(x=>p(305)(98),y=>p(306)(98),Cin=>p(307)(98),clock=>clock,reset=>reset,s=>p(333)(98),cout=>p(334)(99));
FA_ff_12852:FAff port map(x=>p(305)(99),y=>p(306)(99),Cin=>p(307)(99),clock=>clock,reset=>reset,s=>p(333)(99),cout=>p(334)(100));
FA_ff_12853:FAff port map(x=>p(305)(100),y=>p(306)(100),Cin=>p(307)(100),clock=>clock,reset=>reset,s=>p(333)(100),cout=>p(334)(101));
FA_ff_12854:FAff port map(x=>p(305)(101),y=>p(306)(101),Cin=>p(307)(101),clock=>clock,reset=>reset,s=>p(333)(101),cout=>p(334)(102));
FA_ff_12855:FAff port map(x=>p(305)(102),y=>p(306)(102),Cin=>p(307)(102),clock=>clock,reset=>reset,s=>p(333)(102),cout=>p(334)(103));
FA_ff_12856:FAff port map(x=>p(305)(103),y=>p(306)(103),Cin=>p(307)(103),clock=>clock,reset=>reset,s=>p(333)(103),cout=>p(334)(104));
FA_ff_12857:FAff port map(x=>p(305)(104),y=>p(306)(104),Cin=>p(307)(104),clock=>clock,reset=>reset,s=>p(333)(104),cout=>p(334)(105));
FA_ff_12858:FAff port map(x=>p(305)(105),y=>p(306)(105),Cin=>p(307)(105),clock=>clock,reset=>reset,s=>p(333)(105),cout=>p(334)(106));
FA_ff_12859:FAff port map(x=>p(305)(106),y=>p(306)(106),Cin=>p(307)(106),clock=>clock,reset=>reset,s=>p(333)(106),cout=>p(334)(107));
FA_ff_12860:FAff port map(x=>p(305)(107),y=>p(306)(107),Cin=>p(307)(107),clock=>clock,reset=>reset,s=>p(333)(107),cout=>p(334)(108));
FA_ff_12861:FAff port map(x=>p(305)(108),y=>p(306)(108),Cin=>p(307)(108),clock=>clock,reset=>reset,s=>p(333)(108),cout=>p(334)(109));
FA_ff_12862:FAff port map(x=>p(305)(109),y=>p(306)(109),Cin=>p(307)(109),clock=>clock,reset=>reset,s=>p(333)(109),cout=>p(334)(110));
FA_ff_12863:FAff port map(x=>p(305)(110),y=>p(306)(110),Cin=>p(307)(110),clock=>clock,reset=>reset,s=>p(333)(110),cout=>p(334)(111));
FA_ff_12864:FAff port map(x=>p(305)(111),y=>p(306)(111),Cin=>p(307)(111),clock=>clock,reset=>reset,s=>p(333)(111),cout=>p(334)(112));
FA_ff_12865:FAff port map(x=>p(305)(112),y=>p(306)(112),Cin=>p(307)(112),clock=>clock,reset=>reset,s=>p(333)(112),cout=>p(334)(113));
FA_ff_12866:FAff port map(x=>p(305)(113),y=>p(306)(113),Cin=>p(307)(113),clock=>clock,reset=>reset,s=>p(333)(113),cout=>p(334)(114));
FA_ff_12867:FAff port map(x=>p(305)(114),y=>p(306)(114),Cin=>p(307)(114),clock=>clock,reset=>reset,s=>p(333)(114),cout=>p(334)(115));
FA_ff_12868:FAff port map(x=>p(305)(115),y=>p(306)(115),Cin=>p(307)(115),clock=>clock,reset=>reset,s=>p(333)(115),cout=>p(334)(116));
FA_ff_12869:FAff port map(x=>p(305)(116),y=>p(306)(116),Cin=>p(307)(116),clock=>clock,reset=>reset,s=>p(333)(116),cout=>p(334)(117));
FA_ff_12870:FAff port map(x=>p(305)(117),y=>p(306)(117),Cin=>p(307)(117),clock=>clock,reset=>reset,s=>p(333)(117),cout=>p(334)(118));
FA_ff_12871:FAff port map(x=>p(305)(118),y=>p(306)(118),Cin=>p(307)(118),clock=>clock,reset=>reset,s=>p(333)(118),cout=>p(334)(119));
FA_ff_12872:FAff port map(x=>p(305)(119),y=>p(306)(119),Cin=>p(307)(119),clock=>clock,reset=>reset,s=>p(333)(119),cout=>p(334)(120));
FA_ff_12873:FAff port map(x=>p(305)(120),y=>p(306)(120),Cin=>p(307)(120),clock=>clock,reset=>reset,s=>p(333)(120),cout=>p(334)(121));
FA_ff_12874:FAff port map(x=>p(305)(121),y=>p(306)(121),Cin=>p(307)(121),clock=>clock,reset=>reset,s=>p(333)(121),cout=>p(334)(122));
FA_ff_12875:FAff port map(x=>p(305)(122),y=>p(306)(122),Cin=>p(307)(122),clock=>clock,reset=>reset,s=>p(333)(122),cout=>p(334)(123));
FA_ff_12876:FAff port map(x=>p(305)(123),y=>p(306)(123),Cin=>p(307)(123),clock=>clock,reset=>reset,s=>p(333)(123),cout=>p(334)(124));
FA_ff_12877:FAff port map(x=>p(305)(124),y=>p(306)(124),Cin=>p(307)(124),clock=>clock,reset=>reset,s=>p(333)(124),cout=>p(334)(125));
FA_ff_12878:FAff port map(x=>p(305)(125),y=>p(306)(125),Cin=>p(307)(125),clock=>clock,reset=>reset,s=>p(333)(125),cout=>p(334)(126));
FA_ff_12879:FAff port map(x=>p(305)(126),y=>p(306)(126),Cin=>p(307)(126),clock=>clock,reset=>reset,s=>p(333)(126),cout=>p(334)(127));
FA_ff_12880:FAff port map(x=>p(305)(127),y=>p(306)(127),Cin=>p(307)(127),clock=>clock,reset=>reset,s=>p(333)(127),cout=>p(334)(128));
FA_ff_12881:FAff port map(x=>p(305)(128),y=>p(306)(128),Cin=>p(307)(128),clock=>clock,reset=>reset,s=>p(333)(128),cout=>p(334)(129));
FA_ff_12882:FAff port map(x=>p(305)(129),y=>p(306)(129),Cin=>p(307)(129),clock=>clock,reset=>reset,s=>p(333)(129),cout=>p(334)(130));
HA_ff_73:HAff port map(x=>p(308)(0),y=>p(310)(0),clock=>clock,reset=>reset,s=>p(335)(0),c=>p(336)(1));
FA_ff_12883:FAff port map(x=>p(308)(1),y=>p(309)(1),Cin=>p(310)(1),clock=>clock,reset=>reset,s=>p(335)(1),cout=>p(336)(2));
FA_ff_12884:FAff port map(x=>p(308)(2),y=>p(309)(2),Cin=>p(310)(2),clock=>clock,reset=>reset,s=>p(335)(2),cout=>p(336)(3));
FA_ff_12885:FAff port map(x=>p(308)(3),y=>p(309)(3),Cin=>p(310)(3),clock=>clock,reset=>reset,s=>p(335)(3),cout=>p(336)(4));
FA_ff_12886:FAff port map(x=>p(308)(4),y=>p(309)(4),Cin=>p(310)(4),clock=>clock,reset=>reset,s=>p(335)(4),cout=>p(336)(5));
FA_ff_12887:FAff port map(x=>p(308)(5),y=>p(309)(5),Cin=>p(310)(5),clock=>clock,reset=>reset,s=>p(335)(5),cout=>p(336)(6));
FA_ff_12888:FAff port map(x=>p(308)(6),y=>p(309)(6),Cin=>p(310)(6),clock=>clock,reset=>reset,s=>p(335)(6),cout=>p(336)(7));
FA_ff_12889:FAff port map(x=>p(308)(7),y=>p(309)(7),Cin=>p(310)(7),clock=>clock,reset=>reset,s=>p(335)(7),cout=>p(336)(8));
FA_ff_12890:FAff port map(x=>p(308)(8),y=>p(309)(8),Cin=>p(310)(8),clock=>clock,reset=>reset,s=>p(335)(8),cout=>p(336)(9));
FA_ff_12891:FAff port map(x=>p(308)(9),y=>p(309)(9),Cin=>p(310)(9),clock=>clock,reset=>reset,s=>p(335)(9),cout=>p(336)(10));
FA_ff_12892:FAff port map(x=>p(308)(10),y=>p(309)(10),Cin=>p(310)(10),clock=>clock,reset=>reset,s=>p(335)(10),cout=>p(336)(11));
FA_ff_12893:FAff port map(x=>p(308)(11),y=>p(309)(11),Cin=>p(310)(11),clock=>clock,reset=>reset,s=>p(335)(11),cout=>p(336)(12));
FA_ff_12894:FAff port map(x=>p(308)(12),y=>p(309)(12),Cin=>p(310)(12),clock=>clock,reset=>reset,s=>p(335)(12),cout=>p(336)(13));
FA_ff_12895:FAff port map(x=>p(308)(13),y=>p(309)(13),Cin=>p(310)(13),clock=>clock,reset=>reset,s=>p(335)(13),cout=>p(336)(14));
FA_ff_12896:FAff port map(x=>p(308)(14),y=>p(309)(14),Cin=>p(310)(14),clock=>clock,reset=>reset,s=>p(335)(14),cout=>p(336)(15));
FA_ff_12897:FAff port map(x=>p(308)(15),y=>p(309)(15),Cin=>p(310)(15),clock=>clock,reset=>reset,s=>p(335)(15),cout=>p(336)(16));
FA_ff_12898:FAff port map(x=>p(308)(16),y=>p(309)(16),Cin=>p(310)(16),clock=>clock,reset=>reset,s=>p(335)(16),cout=>p(336)(17));
FA_ff_12899:FAff port map(x=>p(308)(17),y=>p(309)(17),Cin=>p(310)(17),clock=>clock,reset=>reset,s=>p(335)(17),cout=>p(336)(18));
FA_ff_12900:FAff port map(x=>p(308)(18),y=>p(309)(18),Cin=>p(310)(18),clock=>clock,reset=>reset,s=>p(335)(18),cout=>p(336)(19));
FA_ff_12901:FAff port map(x=>p(308)(19),y=>p(309)(19),Cin=>p(310)(19),clock=>clock,reset=>reset,s=>p(335)(19),cout=>p(336)(20));
FA_ff_12902:FAff port map(x=>p(308)(20),y=>p(309)(20),Cin=>p(310)(20),clock=>clock,reset=>reset,s=>p(335)(20),cout=>p(336)(21));
FA_ff_12903:FAff port map(x=>p(308)(21),y=>p(309)(21),Cin=>p(310)(21),clock=>clock,reset=>reset,s=>p(335)(21),cout=>p(336)(22));
FA_ff_12904:FAff port map(x=>p(308)(22),y=>p(309)(22),Cin=>p(310)(22),clock=>clock,reset=>reset,s=>p(335)(22),cout=>p(336)(23));
FA_ff_12905:FAff port map(x=>p(308)(23),y=>p(309)(23),Cin=>p(310)(23),clock=>clock,reset=>reset,s=>p(335)(23),cout=>p(336)(24));
FA_ff_12906:FAff port map(x=>p(308)(24),y=>p(309)(24),Cin=>p(310)(24),clock=>clock,reset=>reset,s=>p(335)(24),cout=>p(336)(25));
FA_ff_12907:FAff port map(x=>p(308)(25),y=>p(309)(25),Cin=>p(310)(25),clock=>clock,reset=>reset,s=>p(335)(25),cout=>p(336)(26));
FA_ff_12908:FAff port map(x=>p(308)(26),y=>p(309)(26),Cin=>p(310)(26),clock=>clock,reset=>reset,s=>p(335)(26),cout=>p(336)(27));
FA_ff_12909:FAff port map(x=>p(308)(27),y=>p(309)(27),Cin=>p(310)(27),clock=>clock,reset=>reset,s=>p(335)(27),cout=>p(336)(28));
FA_ff_12910:FAff port map(x=>p(308)(28),y=>p(309)(28),Cin=>p(310)(28),clock=>clock,reset=>reset,s=>p(335)(28),cout=>p(336)(29));
FA_ff_12911:FAff port map(x=>p(308)(29),y=>p(309)(29),Cin=>p(310)(29),clock=>clock,reset=>reset,s=>p(335)(29),cout=>p(336)(30));
FA_ff_12912:FAff port map(x=>p(308)(30),y=>p(309)(30),Cin=>p(310)(30),clock=>clock,reset=>reset,s=>p(335)(30),cout=>p(336)(31));
FA_ff_12913:FAff port map(x=>p(308)(31),y=>p(309)(31),Cin=>p(310)(31),clock=>clock,reset=>reset,s=>p(335)(31),cout=>p(336)(32));
FA_ff_12914:FAff port map(x=>p(308)(32),y=>p(309)(32),Cin=>p(310)(32),clock=>clock,reset=>reset,s=>p(335)(32),cout=>p(336)(33));
FA_ff_12915:FAff port map(x=>p(308)(33),y=>p(309)(33),Cin=>p(310)(33),clock=>clock,reset=>reset,s=>p(335)(33),cout=>p(336)(34));
FA_ff_12916:FAff port map(x=>p(308)(34),y=>p(309)(34),Cin=>p(310)(34),clock=>clock,reset=>reset,s=>p(335)(34),cout=>p(336)(35));
FA_ff_12917:FAff port map(x=>p(308)(35),y=>p(309)(35),Cin=>p(310)(35),clock=>clock,reset=>reset,s=>p(335)(35),cout=>p(336)(36));
FA_ff_12918:FAff port map(x=>p(308)(36),y=>p(309)(36),Cin=>p(310)(36),clock=>clock,reset=>reset,s=>p(335)(36),cout=>p(336)(37));
FA_ff_12919:FAff port map(x=>p(308)(37),y=>p(309)(37),Cin=>p(310)(37),clock=>clock,reset=>reset,s=>p(335)(37),cout=>p(336)(38));
FA_ff_12920:FAff port map(x=>p(308)(38),y=>p(309)(38),Cin=>p(310)(38),clock=>clock,reset=>reset,s=>p(335)(38),cout=>p(336)(39));
FA_ff_12921:FAff port map(x=>p(308)(39),y=>p(309)(39),Cin=>p(310)(39),clock=>clock,reset=>reset,s=>p(335)(39),cout=>p(336)(40));
FA_ff_12922:FAff port map(x=>p(308)(40),y=>p(309)(40),Cin=>p(310)(40),clock=>clock,reset=>reset,s=>p(335)(40),cout=>p(336)(41));
FA_ff_12923:FAff port map(x=>p(308)(41),y=>p(309)(41),Cin=>p(310)(41),clock=>clock,reset=>reset,s=>p(335)(41),cout=>p(336)(42));
FA_ff_12924:FAff port map(x=>p(308)(42),y=>p(309)(42),Cin=>p(310)(42),clock=>clock,reset=>reset,s=>p(335)(42),cout=>p(336)(43));
FA_ff_12925:FAff port map(x=>p(308)(43),y=>p(309)(43),Cin=>p(310)(43),clock=>clock,reset=>reset,s=>p(335)(43),cout=>p(336)(44));
FA_ff_12926:FAff port map(x=>p(308)(44),y=>p(309)(44),Cin=>p(310)(44),clock=>clock,reset=>reset,s=>p(335)(44),cout=>p(336)(45));
FA_ff_12927:FAff port map(x=>p(308)(45),y=>p(309)(45),Cin=>p(310)(45),clock=>clock,reset=>reset,s=>p(335)(45),cout=>p(336)(46));
FA_ff_12928:FAff port map(x=>p(308)(46),y=>p(309)(46),Cin=>p(310)(46),clock=>clock,reset=>reset,s=>p(335)(46),cout=>p(336)(47));
FA_ff_12929:FAff port map(x=>p(308)(47),y=>p(309)(47),Cin=>p(310)(47),clock=>clock,reset=>reset,s=>p(335)(47),cout=>p(336)(48));
FA_ff_12930:FAff port map(x=>p(308)(48),y=>p(309)(48),Cin=>p(310)(48),clock=>clock,reset=>reset,s=>p(335)(48),cout=>p(336)(49));
FA_ff_12931:FAff port map(x=>p(308)(49),y=>p(309)(49),Cin=>p(310)(49),clock=>clock,reset=>reset,s=>p(335)(49),cout=>p(336)(50));
FA_ff_12932:FAff port map(x=>p(308)(50),y=>p(309)(50),Cin=>p(310)(50),clock=>clock,reset=>reset,s=>p(335)(50),cout=>p(336)(51));
FA_ff_12933:FAff port map(x=>p(308)(51),y=>p(309)(51),Cin=>p(310)(51),clock=>clock,reset=>reset,s=>p(335)(51),cout=>p(336)(52));
FA_ff_12934:FAff port map(x=>p(308)(52),y=>p(309)(52),Cin=>p(310)(52),clock=>clock,reset=>reset,s=>p(335)(52),cout=>p(336)(53));
FA_ff_12935:FAff port map(x=>p(308)(53),y=>p(309)(53),Cin=>p(310)(53),clock=>clock,reset=>reset,s=>p(335)(53),cout=>p(336)(54));
FA_ff_12936:FAff port map(x=>p(308)(54),y=>p(309)(54),Cin=>p(310)(54),clock=>clock,reset=>reset,s=>p(335)(54),cout=>p(336)(55));
FA_ff_12937:FAff port map(x=>p(308)(55),y=>p(309)(55),Cin=>p(310)(55),clock=>clock,reset=>reset,s=>p(335)(55),cout=>p(336)(56));
FA_ff_12938:FAff port map(x=>p(308)(56),y=>p(309)(56),Cin=>p(310)(56),clock=>clock,reset=>reset,s=>p(335)(56),cout=>p(336)(57));
FA_ff_12939:FAff port map(x=>p(308)(57),y=>p(309)(57),Cin=>p(310)(57),clock=>clock,reset=>reset,s=>p(335)(57),cout=>p(336)(58));
FA_ff_12940:FAff port map(x=>p(308)(58),y=>p(309)(58),Cin=>p(310)(58),clock=>clock,reset=>reset,s=>p(335)(58),cout=>p(336)(59));
FA_ff_12941:FAff port map(x=>p(308)(59),y=>p(309)(59),Cin=>p(310)(59),clock=>clock,reset=>reset,s=>p(335)(59),cout=>p(336)(60));
FA_ff_12942:FAff port map(x=>p(308)(60),y=>p(309)(60),Cin=>p(310)(60),clock=>clock,reset=>reset,s=>p(335)(60),cout=>p(336)(61));
FA_ff_12943:FAff port map(x=>p(308)(61),y=>p(309)(61),Cin=>p(310)(61),clock=>clock,reset=>reset,s=>p(335)(61),cout=>p(336)(62));
FA_ff_12944:FAff port map(x=>p(308)(62),y=>p(309)(62),Cin=>p(310)(62),clock=>clock,reset=>reset,s=>p(335)(62),cout=>p(336)(63));
FA_ff_12945:FAff port map(x=>p(308)(63),y=>p(309)(63),Cin=>p(310)(63),clock=>clock,reset=>reset,s=>p(335)(63),cout=>p(336)(64));
FA_ff_12946:FAff port map(x=>p(308)(64),y=>p(309)(64),Cin=>p(310)(64),clock=>clock,reset=>reset,s=>p(335)(64),cout=>p(336)(65));
FA_ff_12947:FAff port map(x=>p(308)(65),y=>p(309)(65),Cin=>p(310)(65),clock=>clock,reset=>reset,s=>p(335)(65),cout=>p(336)(66));
FA_ff_12948:FAff port map(x=>p(308)(66),y=>p(309)(66),Cin=>p(310)(66),clock=>clock,reset=>reset,s=>p(335)(66),cout=>p(336)(67));
FA_ff_12949:FAff port map(x=>p(308)(67),y=>p(309)(67),Cin=>p(310)(67),clock=>clock,reset=>reset,s=>p(335)(67),cout=>p(336)(68));
FA_ff_12950:FAff port map(x=>p(308)(68),y=>p(309)(68),Cin=>p(310)(68),clock=>clock,reset=>reset,s=>p(335)(68),cout=>p(336)(69));
FA_ff_12951:FAff port map(x=>p(308)(69),y=>p(309)(69),Cin=>p(310)(69),clock=>clock,reset=>reset,s=>p(335)(69),cout=>p(336)(70));
FA_ff_12952:FAff port map(x=>p(308)(70),y=>p(309)(70),Cin=>p(310)(70),clock=>clock,reset=>reset,s=>p(335)(70),cout=>p(336)(71));
FA_ff_12953:FAff port map(x=>p(308)(71),y=>p(309)(71),Cin=>p(310)(71),clock=>clock,reset=>reset,s=>p(335)(71),cout=>p(336)(72));
FA_ff_12954:FAff port map(x=>p(308)(72),y=>p(309)(72),Cin=>p(310)(72),clock=>clock,reset=>reset,s=>p(335)(72),cout=>p(336)(73));
FA_ff_12955:FAff port map(x=>p(308)(73),y=>p(309)(73),Cin=>p(310)(73),clock=>clock,reset=>reset,s=>p(335)(73),cout=>p(336)(74));
FA_ff_12956:FAff port map(x=>p(308)(74),y=>p(309)(74),Cin=>p(310)(74),clock=>clock,reset=>reset,s=>p(335)(74),cout=>p(336)(75));
FA_ff_12957:FAff port map(x=>p(308)(75),y=>p(309)(75),Cin=>p(310)(75),clock=>clock,reset=>reset,s=>p(335)(75),cout=>p(336)(76));
FA_ff_12958:FAff port map(x=>p(308)(76),y=>p(309)(76),Cin=>p(310)(76),clock=>clock,reset=>reset,s=>p(335)(76),cout=>p(336)(77));
FA_ff_12959:FAff port map(x=>p(308)(77),y=>p(309)(77),Cin=>p(310)(77),clock=>clock,reset=>reset,s=>p(335)(77),cout=>p(336)(78));
FA_ff_12960:FAff port map(x=>p(308)(78),y=>p(309)(78),Cin=>p(310)(78),clock=>clock,reset=>reset,s=>p(335)(78),cout=>p(336)(79));
FA_ff_12961:FAff port map(x=>p(308)(79),y=>p(309)(79),Cin=>p(310)(79),clock=>clock,reset=>reset,s=>p(335)(79),cout=>p(336)(80));
FA_ff_12962:FAff port map(x=>p(308)(80),y=>p(309)(80),Cin=>p(310)(80),clock=>clock,reset=>reset,s=>p(335)(80),cout=>p(336)(81));
FA_ff_12963:FAff port map(x=>p(308)(81),y=>p(309)(81),Cin=>p(310)(81),clock=>clock,reset=>reset,s=>p(335)(81),cout=>p(336)(82));
FA_ff_12964:FAff port map(x=>p(308)(82),y=>p(309)(82),Cin=>p(310)(82),clock=>clock,reset=>reset,s=>p(335)(82),cout=>p(336)(83));
FA_ff_12965:FAff port map(x=>p(308)(83),y=>p(309)(83),Cin=>p(310)(83),clock=>clock,reset=>reset,s=>p(335)(83),cout=>p(336)(84));
FA_ff_12966:FAff port map(x=>p(308)(84),y=>p(309)(84),Cin=>p(310)(84),clock=>clock,reset=>reset,s=>p(335)(84),cout=>p(336)(85));
FA_ff_12967:FAff port map(x=>p(308)(85),y=>p(309)(85),Cin=>p(310)(85),clock=>clock,reset=>reset,s=>p(335)(85),cout=>p(336)(86));
FA_ff_12968:FAff port map(x=>p(308)(86),y=>p(309)(86),Cin=>p(310)(86),clock=>clock,reset=>reset,s=>p(335)(86),cout=>p(336)(87));
FA_ff_12969:FAff port map(x=>p(308)(87),y=>p(309)(87),Cin=>p(310)(87),clock=>clock,reset=>reset,s=>p(335)(87),cout=>p(336)(88));
FA_ff_12970:FAff port map(x=>p(308)(88),y=>p(309)(88),Cin=>p(310)(88),clock=>clock,reset=>reset,s=>p(335)(88),cout=>p(336)(89));
FA_ff_12971:FAff port map(x=>p(308)(89),y=>p(309)(89),Cin=>p(310)(89),clock=>clock,reset=>reset,s=>p(335)(89),cout=>p(336)(90));
FA_ff_12972:FAff port map(x=>p(308)(90),y=>p(309)(90),Cin=>p(310)(90),clock=>clock,reset=>reset,s=>p(335)(90),cout=>p(336)(91));
FA_ff_12973:FAff port map(x=>p(308)(91),y=>p(309)(91),Cin=>p(310)(91),clock=>clock,reset=>reset,s=>p(335)(91),cout=>p(336)(92));
FA_ff_12974:FAff port map(x=>p(308)(92),y=>p(309)(92),Cin=>p(310)(92),clock=>clock,reset=>reset,s=>p(335)(92),cout=>p(336)(93));
FA_ff_12975:FAff port map(x=>p(308)(93),y=>p(309)(93),Cin=>p(310)(93),clock=>clock,reset=>reset,s=>p(335)(93),cout=>p(336)(94));
FA_ff_12976:FAff port map(x=>p(308)(94),y=>p(309)(94),Cin=>p(310)(94),clock=>clock,reset=>reset,s=>p(335)(94),cout=>p(336)(95));
FA_ff_12977:FAff port map(x=>p(308)(95),y=>p(309)(95),Cin=>p(310)(95),clock=>clock,reset=>reset,s=>p(335)(95),cout=>p(336)(96));
FA_ff_12978:FAff port map(x=>p(308)(96),y=>p(309)(96),Cin=>p(310)(96),clock=>clock,reset=>reset,s=>p(335)(96),cout=>p(336)(97));
FA_ff_12979:FAff port map(x=>p(308)(97),y=>p(309)(97),Cin=>p(310)(97),clock=>clock,reset=>reset,s=>p(335)(97),cout=>p(336)(98));
FA_ff_12980:FAff port map(x=>p(308)(98),y=>p(309)(98),Cin=>p(310)(98),clock=>clock,reset=>reset,s=>p(335)(98),cout=>p(336)(99));
FA_ff_12981:FAff port map(x=>p(308)(99),y=>p(309)(99),Cin=>p(310)(99),clock=>clock,reset=>reset,s=>p(335)(99),cout=>p(336)(100));
FA_ff_12982:FAff port map(x=>p(308)(100),y=>p(309)(100),Cin=>p(310)(100),clock=>clock,reset=>reset,s=>p(335)(100),cout=>p(336)(101));
FA_ff_12983:FAff port map(x=>p(308)(101),y=>p(309)(101),Cin=>p(310)(101),clock=>clock,reset=>reset,s=>p(335)(101),cout=>p(336)(102));
FA_ff_12984:FAff port map(x=>p(308)(102),y=>p(309)(102),Cin=>p(310)(102),clock=>clock,reset=>reset,s=>p(335)(102),cout=>p(336)(103));
FA_ff_12985:FAff port map(x=>p(308)(103),y=>p(309)(103),Cin=>p(310)(103),clock=>clock,reset=>reset,s=>p(335)(103),cout=>p(336)(104));
FA_ff_12986:FAff port map(x=>p(308)(104),y=>p(309)(104),Cin=>p(310)(104),clock=>clock,reset=>reset,s=>p(335)(104),cout=>p(336)(105));
FA_ff_12987:FAff port map(x=>p(308)(105),y=>p(309)(105),Cin=>p(310)(105),clock=>clock,reset=>reset,s=>p(335)(105),cout=>p(336)(106));
FA_ff_12988:FAff port map(x=>p(308)(106),y=>p(309)(106),Cin=>p(310)(106),clock=>clock,reset=>reset,s=>p(335)(106),cout=>p(336)(107));
FA_ff_12989:FAff port map(x=>p(308)(107),y=>p(309)(107),Cin=>p(310)(107),clock=>clock,reset=>reset,s=>p(335)(107),cout=>p(336)(108));
FA_ff_12990:FAff port map(x=>p(308)(108),y=>p(309)(108),Cin=>p(310)(108),clock=>clock,reset=>reset,s=>p(335)(108),cout=>p(336)(109));
FA_ff_12991:FAff port map(x=>p(308)(109),y=>p(309)(109),Cin=>p(310)(109),clock=>clock,reset=>reset,s=>p(335)(109),cout=>p(336)(110));
FA_ff_12992:FAff port map(x=>p(308)(110),y=>p(309)(110),Cin=>p(310)(110),clock=>clock,reset=>reset,s=>p(335)(110),cout=>p(336)(111));
FA_ff_12993:FAff port map(x=>p(308)(111),y=>p(309)(111),Cin=>p(310)(111),clock=>clock,reset=>reset,s=>p(335)(111),cout=>p(336)(112));
FA_ff_12994:FAff port map(x=>p(308)(112),y=>p(309)(112),Cin=>p(310)(112),clock=>clock,reset=>reset,s=>p(335)(112),cout=>p(336)(113));
FA_ff_12995:FAff port map(x=>p(308)(113),y=>p(309)(113),Cin=>p(310)(113),clock=>clock,reset=>reset,s=>p(335)(113),cout=>p(336)(114));
FA_ff_12996:FAff port map(x=>p(308)(114),y=>p(309)(114),Cin=>p(310)(114),clock=>clock,reset=>reset,s=>p(335)(114),cout=>p(336)(115));
FA_ff_12997:FAff port map(x=>p(308)(115),y=>p(309)(115),Cin=>p(310)(115),clock=>clock,reset=>reset,s=>p(335)(115),cout=>p(336)(116));
FA_ff_12998:FAff port map(x=>p(308)(116),y=>p(309)(116),Cin=>p(310)(116),clock=>clock,reset=>reset,s=>p(335)(116),cout=>p(336)(117));
FA_ff_12999:FAff port map(x=>p(308)(117),y=>p(309)(117),Cin=>p(310)(117),clock=>clock,reset=>reset,s=>p(335)(117),cout=>p(336)(118));
FA_ff_13000:FAff port map(x=>p(308)(118),y=>p(309)(118),Cin=>p(310)(118),clock=>clock,reset=>reset,s=>p(335)(118),cout=>p(336)(119));
FA_ff_13001:FAff port map(x=>p(308)(119),y=>p(309)(119),Cin=>p(310)(119),clock=>clock,reset=>reset,s=>p(335)(119),cout=>p(336)(120));
FA_ff_13002:FAff port map(x=>p(308)(120),y=>p(309)(120),Cin=>p(310)(120),clock=>clock,reset=>reset,s=>p(335)(120),cout=>p(336)(121));
FA_ff_13003:FAff port map(x=>p(308)(121),y=>p(309)(121),Cin=>p(310)(121),clock=>clock,reset=>reset,s=>p(335)(121),cout=>p(336)(122));
FA_ff_13004:FAff port map(x=>p(308)(122),y=>p(309)(122),Cin=>p(310)(122),clock=>clock,reset=>reset,s=>p(335)(122),cout=>p(336)(123));
FA_ff_13005:FAff port map(x=>p(308)(123),y=>p(309)(123),Cin=>p(310)(123),clock=>clock,reset=>reset,s=>p(335)(123),cout=>p(336)(124));
FA_ff_13006:FAff port map(x=>p(308)(124),y=>p(309)(124),Cin=>p(310)(124),clock=>clock,reset=>reset,s=>p(335)(124),cout=>p(336)(125));
FA_ff_13007:FAff port map(x=>p(308)(125),y=>p(309)(125),Cin=>p(310)(125),clock=>clock,reset=>reset,s=>p(335)(125),cout=>p(336)(126));
FA_ff_13008:FAff port map(x=>p(308)(126),y=>p(309)(126),Cin=>p(310)(126),clock=>clock,reset=>reset,s=>p(335)(126),cout=>p(336)(127));
FA_ff_13009:FAff port map(x=>p(308)(127),y=>p(309)(127),Cin=>p(310)(127),clock=>clock,reset=>reset,s=>p(335)(127),cout=>p(336)(128));
HA_ff_74:HAff port map(x=>p(308)(128),y=>p(309)(128),clock=>clock,reset=>reset,s=>p(335)(128),c=>p(336)(129));
HA_ff_75:HAff port map(x=>p(308)(129),y=>p(309)(129),clock=>clock,reset=>reset,s=>p(335)(129),c=>p(336)(130));
HA_ff_76:HAff port map(x=>p(311)(0),y=>p(313)(0),clock=>clock,reset=>reset,s=>p(337)(0),c=>p(338)(1));
FA_ff_13010:FAff port map(x=>p(311)(1),y=>p(312)(1),Cin=>p(313)(1),clock=>clock,reset=>reset,s=>p(337)(1),cout=>p(338)(2));
FA_ff_13011:FAff port map(x=>p(311)(2),y=>p(312)(2),Cin=>p(313)(2),clock=>clock,reset=>reset,s=>p(337)(2),cout=>p(338)(3));
FA_ff_13012:FAff port map(x=>p(311)(3),y=>p(312)(3),Cin=>p(313)(3),clock=>clock,reset=>reset,s=>p(337)(3),cout=>p(338)(4));
FA_ff_13013:FAff port map(x=>p(311)(4),y=>p(312)(4),Cin=>p(313)(4),clock=>clock,reset=>reset,s=>p(337)(4),cout=>p(338)(5));
FA_ff_13014:FAff port map(x=>p(311)(5),y=>p(312)(5),Cin=>p(313)(5),clock=>clock,reset=>reset,s=>p(337)(5),cout=>p(338)(6));
FA_ff_13015:FAff port map(x=>p(311)(6),y=>p(312)(6),Cin=>p(313)(6),clock=>clock,reset=>reset,s=>p(337)(6),cout=>p(338)(7));
FA_ff_13016:FAff port map(x=>p(311)(7),y=>p(312)(7),Cin=>p(313)(7),clock=>clock,reset=>reset,s=>p(337)(7),cout=>p(338)(8));
FA_ff_13017:FAff port map(x=>p(311)(8),y=>p(312)(8),Cin=>p(313)(8),clock=>clock,reset=>reset,s=>p(337)(8),cout=>p(338)(9));
FA_ff_13018:FAff port map(x=>p(311)(9),y=>p(312)(9),Cin=>p(313)(9),clock=>clock,reset=>reset,s=>p(337)(9),cout=>p(338)(10));
FA_ff_13019:FAff port map(x=>p(311)(10),y=>p(312)(10),Cin=>p(313)(10),clock=>clock,reset=>reset,s=>p(337)(10),cout=>p(338)(11));
FA_ff_13020:FAff port map(x=>p(311)(11),y=>p(312)(11),Cin=>p(313)(11),clock=>clock,reset=>reset,s=>p(337)(11),cout=>p(338)(12));
FA_ff_13021:FAff port map(x=>p(311)(12),y=>p(312)(12),Cin=>p(313)(12),clock=>clock,reset=>reset,s=>p(337)(12),cout=>p(338)(13));
FA_ff_13022:FAff port map(x=>p(311)(13),y=>p(312)(13),Cin=>p(313)(13),clock=>clock,reset=>reset,s=>p(337)(13),cout=>p(338)(14));
FA_ff_13023:FAff port map(x=>p(311)(14),y=>p(312)(14),Cin=>p(313)(14),clock=>clock,reset=>reset,s=>p(337)(14),cout=>p(338)(15));
FA_ff_13024:FAff port map(x=>p(311)(15),y=>p(312)(15),Cin=>p(313)(15),clock=>clock,reset=>reset,s=>p(337)(15),cout=>p(338)(16));
FA_ff_13025:FAff port map(x=>p(311)(16),y=>p(312)(16),Cin=>p(313)(16),clock=>clock,reset=>reset,s=>p(337)(16),cout=>p(338)(17));
FA_ff_13026:FAff port map(x=>p(311)(17),y=>p(312)(17),Cin=>p(313)(17),clock=>clock,reset=>reset,s=>p(337)(17),cout=>p(338)(18));
FA_ff_13027:FAff port map(x=>p(311)(18),y=>p(312)(18),Cin=>p(313)(18),clock=>clock,reset=>reset,s=>p(337)(18),cout=>p(338)(19));
FA_ff_13028:FAff port map(x=>p(311)(19),y=>p(312)(19),Cin=>p(313)(19),clock=>clock,reset=>reset,s=>p(337)(19),cout=>p(338)(20));
FA_ff_13029:FAff port map(x=>p(311)(20),y=>p(312)(20),Cin=>p(313)(20),clock=>clock,reset=>reset,s=>p(337)(20),cout=>p(338)(21));
FA_ff_13030:FAff port map(x=>p(311)(21),y=>p(312)(21),Cin=>p(313)(21),clock=>clock,reset=>reset,s=>p(337)(21),cout=>p(338)(22));
FA_ff_13031:FAff port map(x=>p(311)(22),y=>p(312)(22),Cin=>p(313)(22),clock=>clock,reset=>reset,s=>p(337)(22),cout=>p(338)(23));
FA_ff_13032:FAff port map(x=>p(311)(23),y=>p(312)(23),Cin=>p(313)(23),clock=>clock,reset=>reset,s=>p(337)(23),cout=>p(338)(24));
FA_ff_13033:FAff port map(x=>p(311)(24),y=>p(312)(24),Cin=>p(313)(24),clock=>clock,reset=>reset,s=>p(337)(24),cout=>p(338)(25));
FA_ff_13034:FAff port map(x=>p(311)(25),y=>p(312)(25),Cin=>p(313)(25),clock=>clock,reset=>reset,s=>p(337)(25),cout=>p(338)(26));
FA_ff_13035:FAff port map(x=>p(311)(26),y=>p(312)(26),Cin=>p(313)(26),clock=>clock,reset=>reset,s=>p(337)(26),cout=>p(338)(27));
FA_ff_13036:FAff port map(x=>p(311)(27),y=>p(312)(27),Cin=>p(313)(27),clock=>clock,reset=>reset,s=>p(337)(27),cout=>p(338)(28));
FA_ff_13037:FAff port map(x=>p(311)(28),y=>p(312)(28),Cin=>p(313)(28),clock=>clock,reset=>reset,s=>p(337)(28),cout=>p(338)(29));
FA_ff_13038:FAff port map(x=>p(311)(29),y=>p(312)(29),Cin=>p(313)(29),clock=>clock,reset=>reset,s=>p(337)(29),cout=>p(338)(30));
FA_ff_13039:FAff port map(x=>p(311)(30),y=>p(312)(30),Cin=>p(313)(30),clock=>clock,reset=>reset,s=>p(337)(30),cout=>p(338)(31));
FA_ff_13040:FAff port map(x=>p(311)(31),y=>p(312)(31),Cin=>p(313)(31),clock=>clock,reset=>reset,s=>p(337)(31),cout=>p(338)(32));
FA_ff_13041:FAff port map(x=>p(311)(32),y=>p(312)(32),Cin=>p(313)(32),clock=>clock,reset=>reset,s=>p(337)(32),cout=>p(338)(33));
FA_ff_13042:FAff port map(x=>p(311)(33),y=>p(312)(33),Cin=>p(313)(33),clock=>clock,reset=>reset,s=>p(337)(33),cout=>p(338)(34));
FA_ff_13043:FAff port map(x=>p(311)(34),y=>p(312)(34),Cin=>p(313)(34),clock=>clock,reset=>reset,s=>p(337)(34),cout=>p(338)(35));
FA_ff_13044:FAff port map(x=>p(311)(35),y=>p(312)(35),Cin=>p(313)(35),clock=>clock,reset=>reset,s=>p(337)(35),cout=>p(338)(36));
FA_ff_13045:FAff port map(x=>p(311)(36),y=>p(312)(36),Cin=>p(313)(36),clock=>clock,reset=>reset,s=>p(337)(36),cout=>p(338)(37));
FA_ff_13046:FAff port map(x=>p(311)(37),y=>p(312)(37),Cin=>p(313)(37),clock=>clock,reset=>reset,s=>p(337)(37),cout=>p(338)(38));
FA_ff_13047:FAff port map(x=>p(311)(38),y=>p(312)(38),Cin=>p(313)(38),clock=>clock,reset=>reset,s=>p(337)(38),cout=>p(338)(39));
FA_ff_13048:FAff port map(x=>p(311)(39),y=>p(312)(39),Cin=>p(313)(39),clock=>clock,reset=>reset,s=>p(337)(39),cout=>p(338)(40));
FA_ff_13049:FAff port map(x=>p(311)(40),y=>p(312)(40),Cin=>p(313)(40),clock=>clock,reset=>reset,s=>p(337)(40),cout=>p(338)(41));
FA_ff_13050:FAff port map(x=>p(311)(41),y=>p(312)(41),Cin=>p(313)(41),clock=>clock,reset=>reset,s=>p(337)(41),cout=>p(338)(42));
FA_ff_13051:FAff port map(x=>p(311)(42),y=>p(312)(42),Cin=>p(313)(42),clock=>clock,reset=>reset,s=>p(337)(42),cout=>p(338)(43));
FA_ff_13052:FAff port map(x=>p(311)(43),y=>p(312)(43),Cin=>p(313)(43),clock=>clock,reset=>reset,s=>p(337)(43),cout=>p(338)(44));
FA_ff_13053:FAff port map(x=>p(311)(44),y=>p(312)(44),Cin=>p(313)(44),clock=>clock,reset=>reset,s=>p(337)(44),cout=>p(338)(45));
FA_ff_13054:FAff port map(x=>p(311)(45),y=>p(312)(45),Cin=>p(313)(45),clock=>clock,reset=>reset,s=>p(337)(45),cout=>p(338)(46));
FA_ff_13055:FAff port map(x=>p(311)(46),y=>p(312)(46),Cin=>p(313)(46),clock=>clock,reset=>reset,s=>p(337)(46),cout=>p(338)(47));
FA_ff_13056:FAff port map(x=>p(311)(47),y=>p(312)(47),Cin=>p(313)(47),clock=>clock,reset=>reset,s=>p(337)(47),cout=>p(338)(48));
FA_ff_13057:FAff port map(x=>p(311)(48),y=>p(312)(48),Cin=>p(313)(48),clock=>clock,reset=>reset,s=>p(337)(48),cout=>p(338)(49));
FA_ff_13058:FAff port map(x=>p(311)(49),y=>p(312)(49),Cin=>p(313)(49),clock=>clock,reset=>reset,s=>p(337)(49),cout=>p(338)(50));
FA_ff_13059:FAff port map(x=>p(311)(50),y=>p(312)(50),Cin=>p(313)(50),clock=>clock,reset=>reset,s=>p(337)(50),cout=>p(338)(51));
FA_ff_13060:FAff port map(x=>p(311)(51),y=>p(312)(51),Cin=>p(313)(51),clock=>clock,reset=>reset,s=>p(337)(51),cout=>p(338)(52));
FA_ff_13061:FAff port map(x=>p(311)(52),y=>p(312)(52),Cin=>p(313)(52),clock=>clock,reset=>reset,s=>p(337)(52),cout=>p(338)(53));
FA_ff_13062:FAff port map(x=>p(311)(53),y=>p(312)(53),Cin=>p(313)(53),clock=>clock,reset=>reset,s=>p(337)(53),cout=>p(338)(54));
FA_ff_13063:FAff port map(x=>p(311)(54),y=>p(312)(54),Cin=>p(313)(54),clock=>clock,reset=>reset,s=>p(337)(54),cout=>p(338)(55));
FA_ff_13064:FAff port map(x=>p(311)(55),y=>p(312)(55),Cin=>p(313)(55),clock=>clock,reset=>reset,s=>p(337)(55),cout=>p(338)(56));
FA_ff_13065:FAff port map(x=>p(311)(56),y=>p(312)(56),Cin=>p(313)(56),clock=>clock,reset=>reset,s=>p(337)(56),cout=>p(338)(57));
FA_ff_13066:FAff port map(x=>p(311)(57),y=>p(312)(57),Cin=>p(313)(57),clock=>clock,reset=>reset,s=>p(337)(57),cout=>p(338)(58));
FA_ff_13067:FAff port map(x=>p(311)(58),y=>p(312)(58),Cin=>p(313)(58),clock=>clock,reset=>reset,s=>p(337)(58),cout=>p(338)(59));
FA_ff_13068:FAff port map(x=>p(311)(59),y=>p(312)(59),Cin=>p(313)(59),clock=>clock,reset=>reset,s=>p(337)(59),cout=>p(338)(60));
FA_ff_13069:FAff port map(x=>p(311)(60),y=>p(312)(60),Cin=>p(313)(60),clock=>clock,reset=>reset,s=>p(337)(60),cout=>p(338)(61));
FA_ff_13070:FAff port map(x=>p(311)(61),y=>p(312)(61),Cin=>p(313)(61),clock=>clock,reset=>reset,s=>p(337)(61),cout=>p(338)(62));
FA_ff_13071:FAff port map(x=>p(311)(62),y=>p(312)(62),Cin=>p(313)(62),clock=>clock,reset=>reset,s=>p(337)(62),cout=>p(338)(63));
FA_ff_13072:FAff port map(x=>p(311)(63),y=>p(312)(63),Cin=>p(313)(63),clock=>clock,reset=>reset,s=>p(337)(63),cout=>p(338)(64));
FA_ff_13073:FAff port map(x=>p(311)(64),y=>p(312)(64),Cin=>p(313)(64),clock=>clock,reset=>reset,s=>p(337)(64),cout=>p(338)(65));
FA_ff_13074:FAff port map(x=>p(311)(65),y=>p(312)(65),Cin=>p(313)(65),clock=>clock,reset=>reset,s=>p(337)(65),cout=>p(338)(66));
FA_ff_13075:FAff port map(x=>p(311)(66),y=>p(312)(66),Cin=>p(313)(66),clock=>clock,reset=>reset,s=>p(337)(66),cout=>p(338)(67));
FA_ff_13076:FAff port map(x=>p(311)(67),y=>p(312)(67),Cin=>p(313)(67),clock=>clock,reset=>reset,s=>p(337)(67),cout=>p(338)(68));
FA_ff_13077:FAff port map(x=>p(311)(68),y=>p(312)(68),Cin=>p(313)(68),clock=>clock,reset=>reset,s=>p(337)(68),cout=>p(338)(69));
FA_ff_13078:FAff port map(x=>p(311)(69),y=>p(312)(69),Cin=>p(313)(69),clock=>clock,reset=>reset,s=>p(337)(69),cout=>p(338)(70));
FA_ff_13079:FAff port map(x=>p(311)(70),y=>p(312)(70),Cin=>p(313)(70),clock=>clock,reset=>reset,s=>p(337)(70),cout=>p(338)(71));
FA_ff_13080:FAff port map(x=>p(311)(71),y=>p(312)(71),Cin=>p(313)(71),clock=>clock,reset=>reset,s=>p(337)(71),cout=>p(338)(72));
FA_ff_13081:FAff port map(x=>p(311)(72),y=>p(312)(72),Cin=>p(313)(72),clock=>clock,reset=>reset,s=>p(337)(72),cout=>p(338)(73));
FA_ff_13082:FAff port map(x=>p(311)(73),y=>p(312)(73),Cin=>p(313)(73),clock=>clock,reset=>reset,s=>p(337)(73),cout=>p(338)(74));
FA_ff_13083:FAff port map(x=>p(311)(74),y=>p(312)(74),Cin=>p(313)(74),clock=>clock,reset=>reset,s=>p(337)(74),cout=>p(338)(75));
FA_ff_13084:FAff port map(x=>p(311)(75),y=>p(312)(75),Cin=>p(313)(75),clock=>clock,reset=>reset,s=>p(337)(75),cout=>p(338)(76));
FA_ff_13085:FAff port map(x=>p(311)(76),y=>p(312)(76),Cin=>p(313)(76),clock=>clock,reset=>reset,s=>p(337)(76),cout=>p(338)(77));
FA_ff_13086:FAff port map(x=>p(311)(77),y=>p(312)(77),Cin=>p(313)(77),clock=>clock,reset=>reset,s=>p(337)(77),cout=>p(338)(78));
FA_ff_13087:FAff port map(x=>p(311)(78),y=>p(312)(78),Cin=>p(313)(78),clock=>clock,reset=>reset,s=>p(337)(78),cout=>p(338)(79));
FA_ff_13088:FAff port map(x=>p(311)(79),y=>p(312)(79),Cin=>p(313)(79),clock=>clock,reset=>reset,s=>p(337)(79),cout=>p(338)(80));
FA_ff_13089:FAff port map(x=>p(311)(80),y=>p(312)(80),Cin=>p(313)(80),clock=>clock,reset=>reset,s=>p(337)(80),cout=>p(338)(81));
FA_ff_13090:FAff port map(x=>p(311)(81),y=>p(312)(81),Cin=>p(313)(81),clock=>clock,reset=>reset,s=>p(337)(81),cout=>p(338)(82));
FA_ff_13091:FAff port map(x=>p(311)(82),y=>p(312)(82),Cin=>p(313)(82),clock=>clock,reset=>reset,s=>p(337)(82),cout=>p(338)(83));
FA_ff_13092:FAff port map(x=>p(311)(83),y=>p(312)(83),Cin=>p(313)(83),clock=>clock,reset=>reset,s=>p(337)(83),cout=>p(338)(84));
FA_ff_13093:FAff port map(x=>p(311)(84),y=>p(312)(84),Cin=>p(313)(84),clock=>clock,reset=>reset,s=>p(337)(84),cout=>p(338)(85));
FA_ff_13094:FAff port map(x=>p(311)(85),y=>p(312)(85),Cin=>p(313)(85),clock=>clock,reset=>reset,s=>p(337)(85),cout=>p(338)(86));
FA_ff_13095:FAff port map(x=>p(311)(86),y=>p(312)(86),Cin=>p(313)(86),clock=>clock,reset=>reset,s=>p(337)(86),cout=>p(338)(87));
FA_ff_13096:FAff port map(x=>p(311)(87),y=>p(312)(87),Cin=>p(313)(87),clock=>clock,reset=>reset,s=>p(337)(87),cout=>p(338)(88));
FA_ff_13097:FAff port map(x=>p(311)(88),y=>p(312)(88),Cin=>p(313)(88),clock=>clock,reset=>reset,s=>p(337)(88),cout=>p(338)(89));
FA_ff_13098:FAff port map(x=>p(311)(89),y=>p(312)(89),Cin=>p(313)(89),clock=>clock,reset=>reset,s=>p(337)(89),cout=>p(338)(90));
FA_ff_13099:FAff port map(x=>p(311)(90),y=>p(312)(90),Cin=>p(313)(90),clock=>clock,reset=>reset,s=>p(337)(90),cout=>p(338)(91));
FA_ff_13100:FAff port map(x=>p(311)(91),y=>p(312)(91),Cin=>p(313)(91),clock=>clock,reset=>reset,s=>p(337)(91),cout=>p(338)(92));
FA_ff_13101:FAff port map(x=>p(311)(92),y=>p(312)(92),Cin=>p(313)(92),clock=>clock,reset=>reset,s=>p(337)(92),cout=>p(338)(93));
FA_ff_13102:FAff port map(x=>p(311)(93),y=>p(312)(93),Cin=>p(313)(93),clock=>clock,reset=>reset,s=>p(337)(93),cout=>p(338)(94));
FA_ff_13103:FAff port map(x=>p(311)(94),y=>p(312)(94),Cin=>p(313)(94),clock=>clock,reset=>reset,s=>p(337)(94),cout=>p(338)(95));
FA_ff_13104:FAff port map(x=>p(311)(95),y=>p(312)(95),Cin=>p(313)(95),clock=>clock,reset=>reset,s=>p(337)(95),cout=>p(338)(96));
FA_ff_13105:FAff port map(x=>p(311)(96),y=>p(312)(96),Cin=>p(313)(96),clock=>clock,reset=>reset,s=>p(337)(96),cout=>p(338)(97));
FA_ff_13106:FAff port map(x=>p(311)(97),y=>p(312)(97),Cin=>p(313)(97),clock=>clock,reset=>reset,s=>p(337)(97),cout=>p(338)(98));
FA_ff_13107:FAff port map(x=>p(311)(98),y=>p(312)(98),Cin=>p(313)(98),clock=>clock,reset=>reset,s=>p(337)(98),cout=>p(338)(99));
FA_ff_13108:FAff port map(x=>p(311)(99),y=>p(312)(99),Cin=>p(313)(99),clock=>clock,reset=>reset,s=>p(337)(99),cout=>p(338)(100));
FA_ff_13109:FAff port map(x=>p(311)(100),y=>p(312)(100),Cin=>p(313)(100),clock=>clock,reset=>reset,s=>p(337)(100),cout=>p(338)(101));
FA_ff_13110:FAff port map(x=>p(311)(101),y=>p(312)(101),Cin=>p(313)(101),clock=>clock,reset=>reset,s=>p(337)(101),cout=>p(338)(102));
FA_ff_13111:FAff port map(x=>p(311)(102),y=>p(312)(102),Cin=>p(313)(102),clock=>clock,reset=>reset,s=>p(337)(102),cout=>p(338)(103));
FA_ff_13112:FAff port map(x=>p(311)(103),y=>p(312)(103),Cin=>p(313)(103),clock=>clock,reset=>reset,s=>p(337)(103),cout=>p(338)(104));
FA_ff_13113:FAff port map(x=>p(311)(104),y=>p(312)(104),Cin=>p(313)(104),clock=>clock,reset=>reset,s=>p(337)(104),cout=>p(338)(105));
FA_ff_13114:FAff port map(x=>p(311)(105),y=>p(312)(105),Cin=>p(313)(105),clock=>clock,reset=>reset,s=>p(337)(105),cout=>p(338)(106));
FA_ff_13115:FAff port map(x=>p(311)(106),y=>p(312)(106),Cin=>p(313)(106),clock=>clock,reset=>reset,s=>p(337)(106),cout=>p(338)(107));
FA_ff_13116:FAff port map(x=>p(311)(107),y=>p(312)(107),Cin=>p(313)(107),clock=>clock,reset=>reset,s=>p(337)(107),cout=>p(338)(108));
FA_ff_13117:FAff port map(x=>p(311)(108),y=>p(312)(108),Cin=>p(313)(108),clock=>clock,reset=>reset,s=>p(337)(108),cout=>p(338)(109));
FA_ff_13118:FAff port map(x=>p(311)(109),y=>p(312)(109),Cin=>p(313)(109),clock=>clock,reset=>reset,s=>p(337)(109),cout=>p(338)(110));
FA_ff_13119:FAff port map(x=>p(311)(110),y=>p(312)(110),Cin=>p(313)(110),clock=>clock,reset=>reset,s=>p(337)(110),cout=>p(338)(111));
FA_ff_13120:FAff port map(x=>p(311)(111),y=>p(312)(111),Cin=>p(313)(111),clock=>clock,reset=>reset,s=>p(337)(111),cout=>p(338)(112));
FA_ff_13121:FAff port map(x=>p(311)(112),y=>p(312)(112),Cin=>p(313)(112),clock=>clock,reset=>reset,s=>p(337)(112),cout=>p(338)(113));
FA_ff_13122:FAff port map(x=>p(311)(113),y=>p(312)(113),Cin=>p(313)(113),clock=>clock,reset=>reset,s=>p(337)(113),cout=>p(338)(114));
FA_ff_13123:FAff port map(x=>p(311)(114),y=>p(312)(114),Cin=>p(313)(114),clock=>clock,reset=>reset,s=>p(337)(114),cout=>p(338)(115));
FA_ff_13124:FAff port map(x=>p(311)(115),y=>p(312)(115),Cin=>p(313)(115),clock=>clock,reset=>reset,s=>p(337)(115),cout=>p(338)(116));
FA_ff_13125:FAff port map(x=>p(311)(116),y=>p(312)(116),Cin=>p(313)(116),clock=>clock,reset=>reset,s=>p(337)(116),cout=>p(338)(117));
FA_ff_13126:FAff port map(x=>p(311)(117),y=>p(312)(117),Cin=>p(313)(117),clock=>clock,reset=>reset,s=>p(337)(117),cout=>p(338)(118));
FA_ff_13127:FAff port map(x=>p(311)(118),y=>p(312)(118),Cin=>p(313)(118),clock=>clock,reset=>reset,s=>p(337)(118),cout=>p(338)(119));
FA_ff_13128:FAff port map(x=>p(311)(119),y=>p(312)(119),Cin=>p(313)(119),clock=>clock,reset=>reset,s=>p(337)(119),cout=>p(338)(120));
FA_ff_13129:FAff port map(x=>p(311)(120),y=>p(312)(120),Cin=>p(313)(120),clock=>clock,reset=>reset,s=>p(337)(120),cout=>p(338)(121));
FA_ff_13130:FAff port map(x=>p(311)(121),y=>p(312)(121),Cin=>p(313)(121),clock=>clock,reset=>reset,s=>p(337)(121),cout=>p(338)(122));
FA_ff_13131:FAff port map(x=>p(311)(122),y=>p(312)(122),Cin=>p(313)(122),clock=>clock,reset=>reset,s=>p(337)(122),cout=>p(338)(123));
FA_ff_13132:FAff port map(x=>p(311)(123),y=>p(312)(123),Cin=>p(313)(123),clock=>clock,reset=>reset,s=>p(337)(123),cout=>p(338)(124));
FA_ff_13133:FAff port map(x=>p(311)(124),y=>p(312)(124),Cin=>p(313)(124),clock=>clock,reset=>reset,s=>p(337)(124),cout=>p(338)(125));
FA_ff_13134:FAff port map(x=>p(311)(125),y=>p(312)(125),Cin=>p(313)(125),clock=>clock,reset=>reset,s=>p(337)(125),cout=>p(338)(126));
FA_ff_13135:FAff port map(x=>p(311)(126),y=>p(312)(126),Cin=>p(313)(126),clock=>clock,reset=>reset,s=>p(337)(126),cout=>p(338)(127));
FA_ff_13136:FAff port map(x=>p(311)(127),y=>p(312)(127),Cin=>p(313)(127),clock=>clock,reset=>reset,s=>p(337)(127),cout=>p(338)(128));
FA_ff_13137:FAff port map(x=>p(311)(128),y=>p(312)(128),Cin=>p(313)(128),clock=>clock,reset=>reset,s=>p(337)(128),cout=>p(338)(129));
FA_ff_13138:FAff port map(x=>p(311)(129),y=>p(312)(129),Cin=>p(313)(129),clock=>clock,reset=>reset,s=>p(337)(129),cout=>p(338)(130));
p(337)(130)<=p(312)(130);
p(339)(0)<=p(315)(0);
HA_ff_77:HAff port map(x=>p(315)(1),y=>p(316)(1),clock=>clock,reset=>reset,s=>p(339)(1),c=>p(340)(2));
FA_ff_13139:FAff port map(x=>p(314)(2),y=>p(315)(2),Cin=>p(316)(2),clock=>clock,reset=>reset,s=>p(339)(2),cout=>p(340)(3));
FA_ff_13140:FAff port map(x=>p(314)(3),y=>p(315)(3),Cin=>p(316)(3),clock=>clock,reset=>reset,s=>p(339)(3),cout=>p(340)(4));
FA_ff_13141:FAff port map(x=>p(314)(4),y=>p(315)(4),Cin=>p(316)(4),clock=>clock,reset=>reset,s=>p(339)(4),cout=>p(340)(5));
FA_ff_13142:FAff port map(x=>p(314)(5),y=>p(315)(5),Cin=>p(316)(5),clock=>clock,reset=>reset,s=>p(339)(5),cout=>p(340)(6));
FA_ff_13143:FAff port map(x=>p(314)(6),y=>p(315)(6),Cin=>p(316)(6),clock=>clock,reset=>reset,s=>p(339)(6),cout=>p(340)(7));
FA_ff_13144:FAff port map(x=>p(314)(7),y=>p(315)(7),Cin=>p(316)(7),clock=>clock,reset=>reset,s=>p(339)(7),cout=>p(340)(8));
FA_ff_13145:FAff port map(x=>p(314)(8),y=>p(315)(8),Cin=>p(316)(8),clock=>clock,reset=>reset,s=>p(339)(8),cout=>p(340)(9));
FA_ff_13146:FAff port map(x=>p(314)(9),y=>p(315)(9),Cin=>p(316)(9),clock=>clock,reset=>reset,s=>p(339)(9),cout=>p(340)(10));
FA_ff_13147:FAff port map(x=>p(314)(10),y=>p(315)(10),Cin=>p(316)(10),clock=>clock,reset=>reset,s=>p(339)(10),cout=>p(340)(11));
FA_ff_13148:FAff port map(x=>p(314)(11),y=>p(315)(11),Cin=>p(316)(11),clock=>clock,reset=>reset,s=>p(339)(11),cout=>p(340)(12));
FA_ff_13149:FAff port map(x=>p(314)(12),y=>p(315)(12),Cin=>p(316)(12),clock=>clock,reset=>reset,s=>p(339)(12),cout=>p(340)(13));
FA_ff_13150:FAff port map(x=>p(314)(13),y=>p(315)(13),Cin=>p(316)(13),clock=>clock,reset=>reset,s=>p(339)(13),cout=>p(340)(14));
FA_ff_13151:FAff port map(x=>p(314)(14),y=>p(315)(14),Cin=>p(316)(14),clock=>clock,reset=>reset,s=>p(339)(14),cout=>p(340)(15));
FA_ff_13152:FAff port map(x=>p(314)(15),y=>p(315)(15),Cin=>p(316)(15),clock=>clock,reset=>reset,s=>p(339)(15),cout=>p(340)(16));
FA_ff_13153:FAff port map(x=>p(314)(16),y=>p(315)(16),Cin=>p(316)(16),clock=>clock,reset=>reset,s=>p(339)(16),cout=>p(340)(17));
FA_ff_13154:FAff port map(x=>p(314)(17),y=>p(315)(17),Cin=>p(316)(17),clock=>clock,reset=>reset,s=>p(339)(17),cout=>p(340)(18));
FA_ff_13155:FAff port map(x=>p(314)(18),y=>p(315)(18),Cin=>p(316)(18),clock=>clock,reset=>reset,s=>p(339)(18),cout=>p(340)(19));
FA_ff_13156:FAff port map(x=>p(314)(19),y=>p(315)(19),Cin=>p(316)(19),clock=>clock,reset=>reset,s=>p(339)(19),cout=>p(340)(20));
FA_ff_13157:FAff port map(x=>p(314)(20),y=>p(315)(20),Cin=>p(316)(20),clock=>clock,reset=>reset,s=>p(339)(20),cout=>p(340)(21));
FA_ff_13158:FAff port map(x=>p(314)(21),y=>p(315)(21),Cin=>p(316)(21),clock=>clock,reset=>reset,s=>p(339)(21),cout=>p(340)(22));
FA_ff_13159:FAff port map(x=>p(314)(22),y=>p(315)(22),Cin=>p(316)(22),clock=>clock,reset=>reset,s=>p(339)(22),cout=>p(340)(23));
FA_ff_13160:FAff port map(x=>p(314)(23),y=>p(315)(23),Cin=>p(316)(23),clock=>clock,reset=>reset,s=>p(339)(23),cout=>p(340)(24));
FA_ff_13161:FAff port map(x=>p(314)(24),y=>p(315)(24),Cin=>p(316)(24),clock=>clock,reset=>reset,s=>p(339)(24),cout=>p(340)(25));
FA_ff_13162:FAff port map(x=>p(314)(25),y=>p(315)(25),Cin=>p(316)(25),clock=>clock,reset=>reset,s=>p(339)(25),cout=>p(340)(26));
FA_ff_13163:FAff port map(x=>p(314)(26),y=>p(315)(26),Cin=>p(316)(26),clock=>clock,reset=>reset,s=>p(339)(26),cout=>p(340)(27));
FA_ff_13164:FAff port map(x=>p(314)(27),y=>p(315)(27),Cin=>p(316)(27),clock=>clock,reset=>reset,s=>p(339)(27),cout=>p(340)(28));
FA_ff_13165:FAff port map(x=>p(314)(28),y=>p(315)(28),Cin=>p(316)(28),clock=>clock,reset=>reset,s=>p(339)(28),cout=>p(340)(29));
FA_ff_13166:FAff port map(x=>p(314)(29),y=>p(315)(29),Cin=>p(316)(29),clock=>clock,reset=>reset,s=>p(339)(29),cout=>p(340)(30));
FA_ff_13167:FAff port map(x=>p(314)(30),y=>p(315)(30),Cin=>p(316)(30),clock=>clock,reset=>reset,s=>p(339)(30),cout=>p(340)(31));
FA_ff_13168:FAff port map(x=>p(314)(31),y=>p(315)(31),Cin=>p(316)(31),clock=>clock,reset=>reset,s=>p(339)(31),cout=>p(340)(32));
FA_ff_13169:FAff port map(x=>p(314)(32),y=>p(315)(32),Cin=>p(316)(32),clock=>clock,reset=>reset,s=>p(339)(32),cout=>p(340)(33));
FA_ff_13170:FAff port map(x=>p(314)(33),y=>p(315)(33),Cin=>p(316)(33),clock=>clock,reset=>reset,s=>p(339)(33),cout=>p(340)(34));
FA_ff_13171:FAff port map(x=>p(314)(34),y=>p(315)(34),Cin=>p(316)(34),clock=>clock,reset=>reset,s=>p(339)(34),cout=>p(340)(35));
FA_ff_13172:FAff port map(x=>p(314)(35),y=>p(315)(35),Cin=>p(316)(35),clock=>clock,reset=>reset,s=>p(339)(35),cout=>p(340)(36));
FA_ff_13173:FAff port map(x=>p(314)(36),y=>p(315)(36),Cin=>p(316)(36),clock=>clock,reset=>reset,s=>p(339)(36),cout=>p(340)(37));
FA_ff_13174:FAff port map(x=>p(314)(37),y=>p(315)(37),Cin=>p(316)(37),clock=>clock,reset=>reset,s=>p(339)(37),cout=>p(340)(38));
FA_ff_13175:FAff port map(x=>p(314)(38),y=>p(315)(38),Cin=>p(316)(38),clock=>clock,reset=>reset,s=>p(339)(38),cout=>p(340)(39));
FA_ff_13176:FAff port map(x=>p(314)(39),y=>p(315)(39),Cin=>p(316)(39),clock=>clock,reset=>reset,s=>p(339)(39),cout=>p(340)(40));
FA_ff_13177:FAff port map(x=>p(314)(40),y=>p(315)(40),Cin=>p(316)(40),clock=>clock,reset=>reset,s=>p(339)(40),cout=>p(340)(41));
FA_ff_13178:FAff port map(x=>p(314)(41),y=>p(315)(41),Cin=>p(316)(41),clock=>clock,reset=>reset,s=>p(339)(41),cout=>p(340)(42));
FA_ff_13179:FAff port map(x=>p(314)(42),y=>p(315)(42),Cin=>p(316)(42),clock=>clock,reset=>reset,s=>p(339)(42),cout=>p(340)(43));
FA_ff_13180:FAff port map(x=>p(314)(43),y=>p(315)(43),Cin=>p(316)(43),clock=>clock,reset=>reset,s=>p(339)(43),cout=>p(340)(44));
FA_ff_13181:FAff port map(x=>p(314)(44),y=>p(315)(44),Cin=>p(316)(44),clock=>clock,reset=>reset,s=>p(339)(44),cout=>p(340)(45));
FA_ff_13182:FAff port map(x=>p(314)(45),y=>p(315)(45),Cin=>p(316)(45),clock=>clock,reset=>reset,s=>p(339)(45),cout=>p(340)(46));
FA_ff_13183:FAff port map(x=>p(314)(46),y=>p(315)(46),Cin=>p(316)(46),clock=>clock,reset=>reset,s=>p(339)(46),cout=>p(340)(47));
FA_ff_13184:FAff port map(x=>p(314)(47),y=>p(315)(47),Cin=>p(316)(47),clock=>clock,reset=>reset,s=>p(339)(47),cout=>p(340)(48));
FA_ff_13185:FAff port map(x=>p(314)(48),y=>p(315)(48),Cin=>p(316)(48),clock=>clock,reset=>reset,s=>p(339)(48),cout=>p(340)(49));
FA_ff_13186:FAff port map(x=>p(314)(49),y=>p(315)(49),Cin=>p(316)(49),clock=>clock,reset=>reset,s=>p(339)(49),cout=>p(340)(50));
FA_ff_13187:FAff port map(x=>p(314)(50),y=>p(315)(50),Cin=>p(316)(50),clock=>clock,reset=>reset,s=>p(339)(50),cout=>p(340)(51));
FA_ff_13188:FAff port map(x=>p(314)(51),y=>p(315)(51),Cin=>p(316)(51),clock=>clock,reset=>reset,s=>p(339)(51),cout=>p(340)(52));
FA_ff_13189:FAff port map(x=>p(314)(52),y=>p(315)(52),Cin=>p(316)(52),clock=>clock,reset=>reset,s=>p(339)(52),cout=>p(340)(53));
FA_ff_13190:FAff port map(x=>p(314)(53),y=>p(315)(53),Cin=>p(316)(53),clock=>clock,reset=>reset,s=>p(339)(53),cout=>p(340)(54));
FA_ff_13191:FAff port map(x=>p(314)(54),y=>p(315)(54),Cin=>p(316)(54),clock=>clock,reset=>reset,s=>p(339)(54),cout=>p(340)(55));
FA_ff_13192:FAff port map(x=>p(314)(55),y=>p(315)(55),Cin=>p(316)(55),clock=>clock,reset=>reset,s=>p(339)(55),cout=>p(340)(56));
FA_ff_13193:FAff port map(x=>p(314)(56),y=>p(315)(56),Cin=>p(316)(56),clock=>clock,reset=>reset,s=>p(339)(56),cout=>p(340)(57));
FA_ff_13194:FAff port map(x=>p(314)(57),y=>p(315)(57),Cin=>p(316)(57),clock=>clock,reset=>reset,s=>p(339)(57),cout=>p(340)(58));
FA_ff_13195:FAff port map(x=>p(314)(58),y=>p(315)(58),Cin=>p(316)(58),clock=>clock,reset=>reset,s=>p(339)(58),cout=>p(340)(59));
FA_ff_13196:FAff port map(x=>p(314)(59),y=>p(315)(59),Cin=>p(316)(59),clock=>clock,reset=>reset,s=>p(339)(59),cout=>p(340)(60));
FA_ff_13197:FAff port map(x=>p(314)(60),y=>p(315)(60),Cin=>p(316)(60),clock=>clock,reset=>reset,s=>p(339)(60),cout=>p(340)(61));
FA_ff_13198:FAff port map(x=>p(314)(61),y=>p(315)(61),Cin=>p(316)(61),clock=>clock,reset=>reset,s=>p(339)(61),cout=>p(340)(62));
FA_ff_13199:FAff port map(x=>p(314)(62),y=>p(315)(62),Cin=>p(316)(62),clock=>clock,reset=>reset,s=>p(339)(62),cout=>p(340)(63));
FA_ff_13200:FAff port map(x=>p(314)(63),y=>p(315)(63),Cin=>p(316)(63),clock=>clock,reset=>reset,s=>p(339)(63),cout=>p(340)(64));
FA_ff_13201:FAff port map(x=>p(314)(64),y=>p(315)(64),Cin=>p(316)(64),clock=>clock,reset=>reset,s=>p(339)(64),cout=>p(340)(65));
FA_ff_13202:FAff port map(x=>p(314)(65),y=>p(315)(65),Cin=>p(316)(65),clock=>clock,reset=>reset,s=>p(339)(65),cout=>p(340)(66));
FA_ff_13203:FAff port map(x=>p(314)(66),y=>p(315)(66),Cin=>p(316)(66),clock=>clock,reset=>reset,s=>p(339)(66),cout=>p(340)(67));
FA_ff_13204:FAff port map(x=>p(314)(67),y=>p(315)(67),Cin=>p(316)(67),clock=>clock,reset=>reset,s=>p(339)(67),cout=>p(340)(68));
FA_ff_13205:FAff port map(x=>p(314)(68),y=>p(315)(68),Cin=>p(316)(68),clock=>clock,reset=>reset,s=>p(339)(68),cout=>p(340)(69));
FA_ff_13206:FAff port map(x=>p(314)(69),y=>p(315)(69),Cin=>p(316)(69),clock=>clock,reset=>reset,s=>p(339)(69),cout=>p(340)(70));
FA_ff_13207:FAff port map(x=>p(314)(70),y=>p(315)(70),Cin=>p(316)(70),clock=>clock,reset=>reset,s=>p(339)(70),cout=>p(340)(71));
FA_ff_13208:FAff port map(x=>p(314)(71),y=>p(315)(71),Cin=>p(316)(71),clock=>clock,reset=>reset,s=>p(339)(71),cout=>p(340)(72));
FA_ff_13209:FAff port map(x=>p(314)(72),y=>p(315)(72),Cin=>p(316)(72),clock=>clock,reset=>reset,s=>p(339)(72),cout=>p(340)(73));
FA_ff_13210:FAff port map(x=>p(314)(73),y=>p(315)(73),Cin=>p(316)(73),clock=>clock,reset=>reset,s=>p(339)(73),cout=>p(340)(74));
FA_ff_13211:FAff port map(x=>p(314)(74),y=>p(315)(74),Cin=>p(316)(74),clock=>clock,reset=>reset,s=>p(339)(74),cout=>p(340)(75));
FA_ff_13212:FAff port map(x=>p(314)(75),y=>p(315)(75),Cin=>p(316)(75),clock=>clock,reset=>reset,s=>p(339)(75),cout=>p(340)(76));
FA_ff_13213:FAff port map(x=>p(314)(76),y=>p(315)(76),Cin=>p(316)(76),clock=>clock,reset=>reset,s=>p(339)(76),cout=>p(340)(77));
FA_ff_13214:FAff port map(x=>p(314)(77),y=>p(315)(77),Cin=>p(316)(77),clock=>clock,reset=>reset,s=>p(339)(77),cout=>p(340)(78));
FA_ff_13215:FAff port map(x=>p(314)(78),y=>p(315)(78),Cin=>p(316)(78),clock=>clock,reset=>reset,s=>p(339)(78),cout=>p(340)(79));
FA_ff_13216:FAff port map(x=>p(314)(79),y=>p(315)(79),Cin=>p(316)(79),clock=>clock,reset=>reset,s=>p(339)(79),cout=>p(340)(80));
FA_ff_13217:FAff port map(x=>p(314)(80),y=>p(315)(80),Cin=>p(316)(80),clock=>clock,reset=>reset,s=>p(339)(80),cout=>p(340)(81));
FA_ff_13218:FAff port map(x=>p(314)(81),y=>p(315)(81),Cin=>p(316)(81),clock=>clock,reset=>reset,s=>p(339)(81),cout=>p(340)(82));
FA_ff_13219:FAff port map(x=>p(314)(82),y=>p(315)(82),Cin=>p(316)(82),clock=>clock,reset=>reset,s=>p(339)(82),cout=>p(340)(83));
FA_ff_13220:FAff port map(x=>p(314)(83),y=>p(315)(83),Cin=>p(316)(83),clock=>clock,reset=>reset,s=>p(339)(83),cout=>p(340)(84));
FA_ff_13221:FAff port map(x=>p(314)(84),y=>p(315)(84),Cin=>p(316)(84),clock=>clock,reset=>reset,s=>p(339)(84),cout=>p(340)(85));
FA_ff_13222:FAff port map(x=>p(314)(85),y=>p(315)(85),Cin=>p(316)(85),clock=>clock,reset=>reset,s=>p(339)(85),cout=>p(340)(86));
FA_ff_13223:FAff port map(x=>p(314)(86),y=>p(315)(86),Cin=>p(316)(86),clock=>clock,reset=>reset,s=>p(339)(86),cout=>p(340)(87));
FA_ff_13224:FAff port map(x=>p(314)(87),y=>p(315)(87),Cin=>p(316)(87),clock=>clock,reset=>reset,s=>p(339)(87),cout=>p(340)(88));
FA_ff_13225:FAff port map(x=>p(314)(88),y=>p(315)(88),Cin=>p(316)(88),clock=>clock,reset=>reset,s=>p(339)(88),cout=>p(340)(89));
FA_ff_13226:FAff port map(x=>p(314)(89),y=>p(315)(89),Cin=>p(316)(89),clock=>clock,reset=>reset,s=>p(339)(89),cout=>p(340)(90));
FA_ff_13227:FAff port map(x=>p(314)(90),y=>p(315)(90),Cin=>p(316)(90),clock=>clock,reset=>reset,s=>p(339)(90),cout=>p(340)(91));
FA_ff_13228:FAff port map(x=>p(314)(91),y=>p(315)(91),Cin=>p(316)(91),clock=>clock,reset=>reset,s=>p(339)(91),cout=>p(340)(92));
FA_ff_13229:FAff port map(x=>p(314)(92),y=>p(315)(92),Cin=>p(316)(92),clock=>clock,reset=>reset,s=>p(339)(92),cout=>p(340)(93));
FA_ff_13230:FAff port map(x=>p(314)(93),y=>p(315)(93),Cin=>p(316)(93),clock=>clock,reset=>reset,s=>p(339)(93),cout=>p(340)(94));
FA_ff_13231:FAff port map(x=>p(314)(94),y=>p(315)(94),Cin=>p(316)(94),clock=>clock,reset=>reset,s=>p(339)(94),cout=>p(340)(95));
FA_ff_13232:FAff port map(x=>p(314)(95),y=>p(315)(95),Cin=>p(316)(95),clock=>clock,reset=>reset,s=>p(339)(95),cout=>p(340)(96));
FA_ff_13233:FAff port map(x=>p(314)(96),y=>p(315)(96),Cin=>p(316)(96),clock=>clock,reset=>reset,s=>p(339)(96),cout=>p(340)(97));
FA_ff_13234:FAff port map(x=>p(314)(97),y=>p(315)(97),Cin=>p(316)(97),clock=>clock,reset=>reset,s=>p(339)(97),cout=>p(340)(98));
FA_ff_13235:FAff port map(x=>p(314)(98),y=>p(315)(98),Cin=>p(316)(98),clock=>clock,reset=>reset,s=>p(339)(98),cout=>p(340)(99));
FA_ff_13236:FAff port map(x=>p(314)(99),y=>p(315)(99),Cin=>p(316)(99),clock=>clock,reset=>reset,s=>p(339)(99),cout=>p(340)(100));
FA_ff_13237:FAff port map(x=>p(314)(100),y=>p(315)(100),Cin=>p(316)(100),clock=>clock,reset=>reset,s=>p(339)(100),cout=>p(340)(101));
FA_ff_13238:FAff port map(x=>p(314)(101),y=>p(315)(101),Cin=>p(316)(101),clock=>clock,reset=>reset,s=>p(339)(101),cout=>p(340)(102));
FA_ff_13239:FAff port map(x=>p(314)(102),y=>p(315)(102),Cin=>p(316)(102),clock=>clock,reset=>reset,s=>p(339)(102),cout=>p(340)(103));
FA_ff_13240:FAff port map(x=>p(314)(103),y=>p(315)(103),Cin=>p(316)(103),clock=>clock,reset=>reset,s=>p(339)(103),cout=>p(340)(104));
FA_ff_13241:FAff port map(x=>p(314)(104),y=>p(315)(104),Cin=>p(316)(104),clock=>clock,reset=>reset,s=>p(339)(104),cout=>p(340)(105));
FA_ff_13242:FAff port map(x=>p(314)(105),y=>p(315)(105),Cin=>p(316)(105),clock=>clock,reset=>reset,s=>p(339)(105),cout=>p(340)(106));
FA_ff_13243:FAff port map(x=>p(314)(106),y=>p(315)(106),Cin=>p(316)(106),clock=>clock,reset=>reset,s=>p(339)(106),cout=>p(340)(107));
FA_ff_13244:FAff port map(x=>p(314)(107),y=>p(315)(107),Cin=>p(316)(107),clock=>clock,reset=>reset,s=>p(339)(107),cout=>p(340)(108));
FA_ff_13245:FAff port map(x=>p(314)(108),y=>p(315)(108),Cin=>p(316)(108),clock=>clock,reset=>reset,s=>p(339)(108),cout=>p(340)(109));
FA_ff_13246:FAff port map(x=>p(314)(109),y=>p(315)(109),Cin=>p(316)(109),clock=>clock,reset=>reset,s=>p(339)(109),cout=>p(340)(110));
FA_ff_13247:FAff port map(x=>p(314)(110),y=>p(315)(110),Cin=>p(316)(110),clock=>clock,reset=>reset,s=>p(339)(110),cout=>p(340)(111));
FA_ff_13248:FAff port map(x=>p(314)(111),y=>p(315)(111),Cin=>p(316)(111),clock=>clock,reset=>reset,s=>p(339)(111),cout=>p(340)(112));
FA_ff_13249:FAff port map(x=>p(314)(112),y=>p(315)(112),Cin=>p(316)(112),clock=>clock,reset=>reset,s=>p(339)(112),cout=>p(340)(113));
FA_ff_13250:FAff port map(x=>p(314)(113),y=>p(315)(113),Cin=>p(316)(113),clock=>clock,reset=>reset,s=>p(339)(113),cout=>p(340)(114));
FA_ff_13251:FAff port map(x=>p(314)(114),y=>p(315)(114),Cin=>p(316)(114),clock=>clock,reset=>reset,s=>p(339)(114),cout=>p(340)(115));
FA_ff_13252:FAff port map(x=>p(314)(115),y=>p(315)(115),Cin=>p(316)(115),clock=>clock,reset=>reset,s=>p(339)(115),cout=>p(340)(116));
FA_ff_13253:FAff port map(x=>p(314)(116),y=>p(315)(116),Cin=>p(316)(116),clock=>clock,reset=>reset,s=>p(339)(116),cout=>p(340)(117));
FA_ff_13254:FAff port map(x=>p(314)(117),y=>p(315)(117),Cin=>p(316)(117),clock=>clock,reset=>reset,s=>p(339)(117),cout=>p(340)(118));
FA_ff_13255:FAff port map(x=>p(314)(118),y=>p(315)(118),Cin=>p(316)(118),clock=>clock,reset=>reset,s=>p(339)(118),cout=>p(340)(119));
FA_ff_13256:FAff port map(x=>p(314)(119),y=>p(315)(119),Cin=>p(316)(119),clock=>clock,reset=>reset,s=>p(339)(119),cout=>p(340)(120));
FA_ff_13257:FAff port map(x=>p(314)(120),y=>p(315)(120),Cin=>p(316)(120),clock=>clock,reset=>reset,s=>p(339)(120),cout=>p(340)(121));
FA_ff_13258:FAff port map(x=>p(314)(121),y=>p(315)(121),Cin=>p(316)(121),clock=>clock,reset=>reset,s=>p(339)(121),cout=>p(340)(122));
FA_ff_13259:FAff port map(x=>p(314)(122),y=>p(315)(122),Cin=>p(316)(122),clock=>clock,reset=>reset,s=>p(339)(122),cout=>p(340)(123));
FA_ff_13260:FAff port map(x=>p(314)(123),y=>p(315)(123),Cin=>p(316)(123),clock=>clock,reset=>reset,s=>p(339)(123),cout=>p(340)(124));
FA_ff_13261:FAff port map(x=>p(314)(124),y=>p(315)(124),Cin=>p(316)(124),clock=>clock,reset=>reset,s=>p(339)(124),cout=>p(340)(125));
FA_ff_13262:FAff port map(x=>p(314)(125),y=>p(315)(125),Cin=>p(316)(125),clock=>clock,reset=>reset,s=>p(339)(125),cout=>p(340)(126));
FA_ff_13263:FAff port map(x=>p(314)(126),y=>p(315)(126),Cin=>p(316)(126),clock=>clock,reset=>reset,s=>p(339)(126),cout=>p(340)(127));
FA_ff_13264:FAff port map(x=>p(314)(127),y=>p(315)(127),Cin=>p(316)(127),clock=>clock,reset=>reset,s=>p(339)(127),cout=>p(340)(128));
FA_ff_13265:FAff port map(x=>p(314)(128),y=>p(315)(128),Cin=>p(316)(128),clock=>clock,reset=>reset,s=>p(339)(128),cout=>p(340)(129));
FA_ff_13266:FAff port map(x=>p(314)(129),y=>p(315)(129),Cin=>p(316)(129),clock=>clock,reset=>reset,s=>p(339)(129),cout=>p(340)(130));
HA_ff_78:HAff port map(x=>p(314)(130),y=>p(316)(130),clock=>clock,reset=>reset,s=>p(339)(130),c=>p(340)(131));
HA_ff_79:HAff port map(x=>p(317)(0),y=>p(319)(0),clock=>clock,reset=>reset,s=>p(341)(0),c=>p(342)(1));
HA_ff_80:HAff port map(x=>p(317)(1),y=>p(319)(1),clock=>clock,reset=>reset,s=>p(341)(1),c=>p(342)(2));
FA_ff_13267:FAff port map(x=>p(317)(2),y=>p(318)(2),Cin=>p(319)(2),clock=>clock,reset=>reset,s=>p(341)(2),cout=>p(342)(3));
FA_ff_13268:FAff port map(x=>p(317)(3),y=>p(318)(3),Cin=>p(319)(3),clock=>clock,reset=>reset,s=>p(341)(3),cout=>p(342)(4));
FA_ff_13269:FAff port map(x=>p(317)(4),y=>p(318)(4),Cin=>p(319)(4),clock=>clock,reset=>reset,s=>p(341)(4),cout=>p(342)(5));
FA_ff_13270:FAff port map(x=>p(317)(5),y=>p(318)(5),Cin=>p(319)(5),clock=>clock,reset=>reset,s=>p(341)(5),cout=>p(342)(6));
FA_ff_13271:FAff port map(x=>p(317)(6),y=>p(318)(6),Cin=>p(319)(6),clock=>clock,reset=>reset,s=>p(341)(6),cout=>p(342)(7));
FA_ff_13272:FAff port map(x=>p(317)(7),y=>p(318)(7),Cin=>p(319)(7),clock=>clock,reset=>reset,s=>p(341)(7),cout=>p(342)(8));
FA_ff_13273:FAff port map(x=>p(317)(8),y=>p(318)(8),Cin=>p(319)(8),clock=>clock,reset=>reset,s=>p(341)(8),cout=>p(342)(9));
FA_ff_13274:FAff port map(x=>p(317)(9),y=>p(318)(9),Cin=>p(319)(9),clock=>clock,reset=>reset,s=>p(341)(9),cout=>p(342)(10));
FA_ff_13275:FAff port map(x=>p(317)(10),y=>p(318)(10),Cin=>p(319)(10),clock=>clock,reset=>reset,s=>p(341)(10),cout=>p(342)(11));
FA_ff_13276:FAff port map(x=>p(317)(11),y=>p(318)(11),Cin=>p(319)(11),clock=>clock,reset=>reset,s=>p(341)(11),cout=>p(342)(12));
FA_ff_13277:FAff port map(x=>p(317)(12),y=>p(318)(12),Cin=>p(319)(12),clock=>clock,reset=>reset,s=>p(341)(12),cout=>p(342)(13));
FA_ff_13278:FAff port map(x=>p(317)(13),y=>p(318)(13),Cin=>p(319)(13),clock=>clock,reset=>reset,s=>p(341)(13),cout=>p(342)(14));
FA_ff_13279:FAff port map(x=>p(317)(14),y=>p(318)(14),Cin=>p(319)(14),clock=>clock,reset=>reset,s=>p(341)(14),cout=>p(342)(15));
FA_ff_13280:FAff port map(x=>p(317)(15),y=>p(318)(15),Cin=>p(319)(15),clock=>clock,reset=>reset,s=>p(341)(15),cout=>p(342)(16));
FA_ff_13281:FAff port map(x=>p(317)(16),y=>p(318)(16),Cin=>p(319)(16),clock=>clock,reset=>reset,s=>p(341)(16),cout=>p(342)(17));
FA_ff_13282:FAff port map(x=>p(317)(17),y=>p(318)(17),Cin=>p(319)(17),clock=>clock,reset=>reset,s=>p(341)(17),cout=>p(342)(18));
FA_ff_13283:FAff port map(x=>p(317)(18),y=>p(318)(18),Cin=>p(319)(18),clock=>clock,reset=>reset,s=>p(341)(18),cout=>p(342)(19));
FA_ff_13284:FAff port map(x=>p(317)(19),y=>p(318)(19),Cin=>p(319)(19),clock=>clock,reset=>reset,s=>p(341)(19),cout=>p(342)(20));
FA_ff_13285:FAff port map(x=>p(317)(20),y=>p(318)(20),Cin=>p(319)(20),clock=>clock,reset=>reset,s=>p(341)(20),cout=>p(342)(21));
FA_ff_13286:FAff port map(x=>p(317)(21),y=>p(318)(21),Cin=>p(319)(21),clock=>clock,reset=>reset,s=>p(341)(21),cout=>p(342)(22));
FA_ff_13287:FAff port map(x=>p(317)(22),y=>p(318)(22),Cin=>p(319)(22),clock=>clock,reset=>reset,s=>p(341)(22),cout=>p(342)(23));
FA_ff_13288:FAff port map(x=>p(317)(23),y=>p(318)(23),Cin=>p(319)(23),clock=>clock,reset=>reset,s=>p(341)(23),cout=>p(342)(24));
FA_ff_13289:FAff port map(x=>p(317)(24),y=>p(318)(24),Cin=>p(319)(24),clock=>clock,reset=>reset,s=>p(341)(24),cout=>p(342)(25));
FA_ff_13290:FAff port map(x=>p(317)(25),y=>p(318)(25),Cin=>p(319)(25),clock=>clock,reset=>reset,s=>p(341)(25),cout=>p(342)(26));
FA_ff_13291:FAff port map(x=>p(317)(26),y=>p(318)(26),Cin=>p(319)(26),clock=>clock,reset=>reset,s=>p(341)(26),cout=>p(342)(27));
FA_ff_13292:FAff port map(x=>p(317)(27),y=>p(318)(27),Cin=>p(319)(27),clock=>clock,reset=>reset,s=>p(341)(27),cout=>p(342)(28));
FA_ff_13293:FAff port map(x=>p(317)(28),y=>p(318)(28),Cin=>p(319)(28),clock=>clock,reset=>reset,s=>p(341)(28),cout=>p(342)(29));
FA_ff_13294:FAff port map(x=>p(317)(29),y=>p(318)(29),Cin=>p(319)(29),clock=>clock,reset=>reset,s=>p(341)(29),cout=>p(342)(30));
FA_ff_13295:FAff port map(x=>p(317)(30),y=>p(318)(30),Cin=>p(319)(30),clock=>clock,reset=>reset,s=>p(341)(30),cout=>p(342)(31));
FA_ff_13296:FAff port map(x=>p(317)(31),y=>p(318)(31),Cin=>p(319)(31),clock=>clock,reset=>reset,s=>p(341)(31),cout=>p(342)(32));
FA_ff_13297:FAff port map(x=>p(317)(32),y=>p(318)(32),Cin=>p(319)(32),clock=>clock,reset=>reset,s=>p(341)(32),cout=>p(342)(33));
FA_ff_13298:FAff port map(x=>p(317)(33),y=>p(318)(33),Cin=>p(319)(33),clock=>clock,reset=>reset,s=>p(341)(33),cout=>p(342)(34));
FA_ff_13299:FAff port map(x=>p(317)(34),y=>p(318)(34),Cin=>p(319)(34),clock=>clock,reset=>reset,s=>p(341)(34),cout=>p(342)(35));
FA_ff_13300:FAff port map(x=>p(317)(35),y=>p(318)(35),Cin=>p(319)(35),clock=>clock,reset=>reset,s=>p(341)(35),cout=>p(342)(36));
FA_ff_13301:FAff port map(x=>p(317)(36),y=>p(318)(36),Cin=>p(319)(36),clock=>clock,reset=>reset,s=>p(341)(36),cout=>p(342)(37));
FA_ff_13302:FAff port map(x=>p(317)(37),y=>p(318)(37),Cin=>p(319)(37),clock=>clock,reset=>reset,s=>p(341)(37),cout=>p(342)(38));
FA_ff_13303:FAff port map(x=>p(317)(38),y=>p(318)(38),Cin=>p(319)(38),clock=>clock,reset=>reset,s=>p(341)(38),cout=>p(342)(39));
FA_ff_13304:FAff port map(x=>p(317)(39),y=>p(318)(39),Cin=>p(319)(39),clock=>clock,reset=>reset,s=>p(341)(39),cout=>p(342)(40));
FA_ff_13305:FAff port map(x=>p(317)(40),y=>p(318)(40),Cin=>p(319)(40),clock=>clock,reset=>reset,s=>p(341)(40),cout=>p(342)(41));
FA_ff_13306:FAff port map(x=>p(317)(41),y=>p(318)(41),Cin=>p(319)(41),clock=>clock,reset=>reset,s=>p(341)(41),cout=>p(342)(42));
FA_ff_13307:FAff port map(x=>p(317)(42),y=>p(318)(42),Cin=>p(319)(42),clock=>clock,reset=>reset,s=>p(341)(42),cout=>p(342)(43));
FA_ff_13308:FAff port map(x=>p(317)(43),y=>p(318)(43),Cin=>p(319)(43),clock=>clock,reset=>reset,s=>p(341)(43),cout=>p(342)(44));
FA_ff_13309:FAff port map(x=>p(317)(44),y=>p(318)(44),Cin=>p(319)(44),clock=>clock,reset=>reset,s=>p(341)(44),cout=>p(342)(45));
FA_ff_13310:FAff port map(x=>p(317)(45),y=>p(318)(45),Cin=>p(319)(45),clock=>clock,reset=>reset,s=>p(341)(45),cout=>p(342)(46));
FA_ff_13311:FAff port map(x=>p(317)(46),y=>p(318)(46),Cin=>p(319)(46),clock=>clock,reset=>reset,s=>p(341)(46),cout=>p(342)(47));
FA_ff_13312:FAff port map(x=>p(317)(47),y=>p(318)(47),Cin=>p(319)(47),clock=>clock,reset=>reset,s=>p(341)(47),cout=>p(342)(48));
FA_ff_13313:FAff port map(x=>p(317)(48),y=>p(318)(48),Cin=>p(319)(48),clock=>clock,reset=>reset,s=>p(341)(48),cout=>p(342)(49));
FA_ff_13314:FAff port map(x=>p(317)(49),y=>p(318)(49),Cin=>p(319)(49),clock=>clock,reset=>reset,s=>p(341)(49),cout=>p(342)(50));
FA_ff_13315:FAff port map(x=>p(317)(50),y=>p(318)(50),Cin=>p(319)(50),clock=>clock,reset=>reset,s=>p(341)(50),cout=>p(342)(51));
FA_ff_13316:FAff port map(x=>p(317)(51),y=>p(318)(51),Cin=>p(319)(51),clock=>clock,reset=>reset,s=>p(341)(51),cout=>p(342)(52));
FA_ff_13317:FAff port map(x=>p(317)(52),y=>p(318)(52),Cin=>p(319)(52),clock=>clock,reset=>reset,s=>p(341)(52),cout=>p(342)(53));
FA_ff_13318:FAff port map(x=>p(317)(53),y=>p(318)(53),Cin=>p(319)(53),clock=>clock,reset=>reset,s=>p(341)(53),cout=>p(342)(54));
FA_ff_13319:FAff port map(x=>p(317)(54),y=>p(318)(54),Cin=>p(319)(54),clock=>clock,reset=>reset,s=>p(341)(54),cout=>p(342)(55));
FA_ff_13320:FAff port map(x=>p(317)(55),y=>p(318)(55),Cin=>p(319)(55),clock=>clock,reset=>reset,s=>p(341)(55),cout=>p(342)(56));
FA_ff_13321:FAff port map(x=>p(317)(56),y=>p(318)(56),Cin=>p(319)(56),clock=>clock,reset=>reset,s=>p(341)(56),cout=>p(342)(57));
FA_ff_13322:FAff port map(x=>p(317)(57),y=>p(318)(57),Cin=>p(319)(57),clock=>clock,reset=>reset,s=>p(341)(57),cout=>p(342)(58));
FA_ff_13323:FAff port map(x=>p(317)(58),y=>p(318)(58),Cin=>p(319)(58),clock=>clock,reset=>reset,s=>p(341)(58),cout=>p(342)(59));
FA_ff_13324:FAff port map(x=>p(317)(59),y=>p(318)(59),Cin=>p(319)(59),clock=>clock,reset=>reset,s=>p(341)(59),cout=>p(342)(60));
FA_ff_13325:FAff port map(x=>p(317)(60),y=>p(318)(60),Cin=>p(319)(60),clock=>clock,reset=>reset,s=>p(341)(60),cout=>p(342)(61));
FA_ff_13326:FAff port map(x=>p(317)(61),y=>p(318)(61),Cin=>p(319)(61),clock=>clock,reset=>reset,s=>p(341)(61),cout=>p(342)(62));
FA_ff_13327:FAff port map(x=>p(317)(62),y=>p(318)(62),Cin=>p(319)(62),clock=>clock,reset=>reset,s=>p(341)(62),cout=>p(342)(63));
FA_ff_13328:FAff port map(x=>p(317)(63),y=>p(318)(63),Cin=>p(319)(63),clock=>clock,reset=>reset,s=>p(341)(63),cout=>p(342)(64));
FA_ff_13329:FAff port map(x=>p(317)(64),y=>p(318)(64),Cin=>p(319)(64),clock=>clock,reset=>reset,s=>p(341)(64),cout=>p(342)(65));
FA_ff_13330:FAff port map(x=>p(317)(65),y=>p(318)(65),Cin=>p(319)(65),clock=>clock,reset=>reset,s=>p(341)(65),cout=>p(342)(66));
FA_ff_13331:FAff port map(x=>p(317)(66),y=>p(318)(66),Cin=>p(319)(66),clock=>clock,reset=>reset,s=>p(341)(66),cout=>p(342)(67));
FA_ff_13332:FAff port map(x=>p(317)(67),y=>p(318)(67),Cin=>p(319)(67),clock=>clock,reset=>reset,s=>p(341)(67),cout=>p(342)(68));
FA_ff_13333:FAff port map(x=>p(317)(68),y=>p(318)(68),Cin=>p(319)(68),clock=>clock,reset=>reset,s=>p(341)(68),cout=>p(342)(69));
FA_ff_13334:FAff port map(x=>p(317)(69),y=>p(318)(69),Cin=>p(319)(69),clock=>clock,reset=>reset,s=>p(341)(69),cout=>p(342)(70));
FA_ff_13335:FAff port map(x=>p(317)(70),y=>p(318)(70),Cin=>p(319)(70),clock=>clock,reset=>reset,s=>p(341)(70),cout=>p(342)(71));
FA_ff_13336:FAff port map(x=>p(317)(71),y=>p(318)(71),Cin=>p(319)(71),clock=>clock,reset=>reset,s=>p(341)(71),cout=>p(342)(72));
FA_ff_13337:FAff port map(x=>p(317)(72),y=>p(318)(72),Cin=>p(319)(72),clock=>clock,reset=>reset,s=>p(341)(72),cout=>p(342)(73));
FA_ff_13338:FAff port map(x=>p(317)(73),y=>p(318)(73),Cin=>p(319)(73),clock=>clock,reset=>reset,s=>p(341)(73),cout=>p(342)(74));
FA_ff_13339:FAff port map(x=>p(317)(74),y=>p(318)(74),Cin=>p(319)(74),clock=>clock,reset=>reset,s=>p(341)(74),cout=>p(342)(75));
FA_ff_13340:FAff port map(x=>p(317)(75),y=>p(318)(75),Cin=>p(319)(75),clock=>clock,reset=>reset,s=>p(341)(75),cout=>p(342)(76));
FA_ff_13341:FAff port map(x=>p(317)(76),y=>p(318)(76),Cin=>p(319)(76),clock=>clock,reset=>reset,s=>p(341)(76),cout=>p(342)(77));
FA_ff_13342:FAff port map(x=>p(317)(77),y=>p(318)(77),Cin=>p(319)(77),clock=>clock,reset=>reset,s=>p(341)(77),cout=>p(342)(78));
FA_ff_13343:FAff port map(x=>p(317)(78),y=>p(318)(78),Cin=>p(319)(78),clock=>clock,reset=>reset,s=>p(341)(78),cout=>p(342)(79));
FA_ff_13344:FAff port map(x=>p(317)(79),y=>p(318)(79),Cin=>p(319)(79),clock=>clock,reset=>reset,s=>p(341)(79),cout=>p(342)(80));
FA_ff_13345:FAff port map(x=>p(317)(80),y=>p(318)(80),Cin=>p(319)(80),clock=>clock,reset=>reset,s=>p(341)(80),cout=>p(342)(81));
FA_ff_13346:FAff port map(x=>p(317)(81),y=>p(318)(81),Cin=>p(319)(81),clock=>clock,reset=>reset,s=>p(341)(81),cout=>p(342)(82));
FA_ff_13347:FAff port map(x=>p(317)(82),y=>p(318)(82),Cin=>p(319)(82),clock=>clock,reset=>reset,s=>p(341)(82),cout=>p(342)(83));
FA_ff_13348:FAff port map(x=>p(317)(83),y=>p(318)(83),Cin=>p(319)(83),clock=>clock,reset=>reset,s=>p(341)(83),cout=>p(342)(84));
FA_ff_13349:FAff port map(x=>p(317)(84),y=>p(318)(84),Cin=>p(319)(84),clock=>clock,reset=>reset,s=>p(341)(84),cout=>p(342)(85));
FA_ff_13350:FAff port map(x=>p(317)(85),y=>p(318)(85),Cin=>p(319)(85),clock=>clock,reset=>reset,s=>p(341)(85),cout=>p(342)(86));
FA_ff_13351:FAff port map(x=>p(317)(86),y=>p(318)(86),Cin=>p(319)(86),clock=>clock,reset=>reset,s=>p(341)(86),cout=>p(342)(87));
FA_ff_13352:FAff port map(x=>p(317)(87),y=>p(318)(87),Cin=>p(319)(87),clock=>clock,reset=>reset,s=>p(341)(87),cout=>p(342)(88));
FA_ff_13353:FAff port map(x=>p(317)(88),y=>p(318)(88),Cin=>p(319)(88),clock=>clock,reset=>reset,s=>p(341)(88),cout=>p(342)(89));
FA_ff_13354:FAff port map(x=>p(317)(89),y=>p(318)(89),Cin=>p(319)(89),clock=>clock,reset=>reset,s=>p(341)(89),cout=>p(342)(90));
FA_ff_13355:FAff port map(x=>p(317)(90),y=>p(318)(90),Cin=>p(319)(90),clock=>clock,reset=>reset,s=>p(341)(90),cout=>p(342)(91));
FA_ff_13356:FAff port map(x=>p(317)(91),y=>p(318)(91),Cin=>p(319)(91),clock=>clock,reset=>reset,s=>p(341)(91),cout=>p(342)(92));
FA_ff_13357:FAff port map(x=>p(317)(92),y=>p(318)(92),Cin=>p(319)(92),clock=>clock,reset=>reset,s=>p(341)(92),cout=>p(342)(93));
FA_ff_13358:FAff port map(x=>p(317)(93),y=>p(318)(93),Cin=>p(319)(93),clock=>clock,reset=>reset,s=>p(341)(93),cout=>p(342)(94));
FA_ff_13359:FAff port map(x=>p(317)(94),y=>p(318)(94),Cin=>p(319)(94),clock=>clock,reset=>reset,s=>p(341)(94),cout=>p(342)(95));
FA_ff_13360:FAff port map(x=>p(317)(95),y=>p(318)(95),Cin=>p(319)(95),clock=>clock,reset=>reset,s=>p(341)(95),cout=>p(342)(96));
FA_ff_13361:FAff port map(x=>p(317)(96),y=>p(318)(96),Cin=>p(319)(96),clock=>clock,reset=>reset,s=>p(341)(96),cout=>p(342)(97));
FA_ff_13362:FAff port map(x=>p(317)(97),y=>p(318)(97),Cin=>p(319)(97),clock=>clock,reset=>reset,s=>p(341)(97),cout=>p(342)(98));
FA_ff_13363:FAff port map(x=>p(317)(98),y=>p(318)(98),Cin=>p(319)(98),clock=>clock,reset=>reset,s=>p(341)(98),cout=>p(342)(99));
FA_ff_13364:FAff port map(x=>p(317)(99),y=>p(318)(99),Cin=>p(319)(99),clock=>clock,reset=>reset,s=>p(341)(99),cout=>p(342)(100));
FA_ff_13365:FAff port map(x=>p(317)(100),y=>p(318)(100),Cin=>p(319)(100),clock=>clock,reset=>reset,s=>p(341)(100),cout=>p(342)(101));
FA_ff_13366:FAff port map(x=>p(317)(101),y=>p(318)(101),Cin=>p(319)(101),clock=>clock,reset=>reset,s=>p(341)(101),cout=>p(342)(102));
FA_ff_13367:FAff port map(x=>p(317)(102),y=>p(318)(102),Cin=>p(319)(102),clock=>clock,reset=>reset,s=>p(341)(102),cout=>p(342)(103));
FA_ff_13368:FAff port map(x=>p(317)(103),y=>p(318)(103),Cin=>p(319)(103),clock=>clock,reset=>reset,s=>p(341)(103),cout=>p(342)(104));
FA_ff_13369:FAff port map(x=>p(317)(104),y=>p(318)(104),Cin=>p(319)(104),clock=>clock,reset=>reset,s=>p(341)(104),cout=>p(342)(105));
FA_ff_13370:FAff port map(x=>p(317)(105),y=>p(318)(105),Cin=>p(319)(105),clock=>clock,reset=>reset,s=>p(341)(105),cout=>p(342)(106));
FA_ff_13371:FAff port map(x=>p(317)(106),y=>p(318)(106),Cin=>p(319)(106),clock=>clock,reset=>reset,s=>p(341)(106),cout=>p(342)(107));
FA_ff_13372:FAff port map(x=>p(317)(107),y=>p(318)(107),Cin=>p(319)(107),clock=>clock,reset=>reset,s=>p(341)(107),cout=>p(342)(108));
FA_ff_13373:FAff port map(x=>p(317)(108),y=>p(318)(108),Cin=>p(319)(108),clock=>clock,reset=>reset,s=>p(341)(108),cout=>p(342)(109));
FA_ff_13374:FAff port map(x=>p(317)(109),y=>p(318)(109),Cin=>p(319)(109),clock=>clock,reset=>reset,s=>p(341)(109),cout=>p(342)(110));
FA_ff_13375:FAff port map(x=>p(317)(110),y=>p(318)(110),Cin=>p(319)(110),clock=>clock,reset=>reset,s=>p(341)(110),cout=>p(342)(111));
FA_ff_13376:FAff port map(x=>p(317)(111),y=>p(318)(111),Cin=>p(319)(111),clock=>clock,reset=>reset,s=>p(341)(111),cout=>p(342)(112));
FA_ff_13377:FAff port map(x=>p(317)(112),y=>p(318)(112),Cin=>p(319)(112),clock=>clock,reset=>reset,s=>p(341)(112),cout=>p(342)(113));
FA_ff_13378:FAff port map(x=>p(317)(113),y=>p(318)(113),Cin=>p(319)(113),clock=>clock,reset=>reset,s=>p(341)(113),cout=>p(342)(114));
FA_ff_13379:FAff port map(x=>p(317)(114),y=>p(318)(114),Cin=>p(319)(114),clock=>clock,reset=>reset,s=>p(341)(114),cout=>p(342)(115));
FA_ff_13380:FAff port map(x=>p(317)(115),y=>p(318)(115),Cin=>p(319)(115),clock=>clock,reset=>reset,s=>p(341)(115),cout=>p(342)(116));
FA_ff_13381:FAff port map(x=>p(317)(116),y=>p(318)(116),Cin=>p(319)(116),clock=>clock,reset=>reset,s=>p(341)(116),cout=>p(342)(117));
FA_ff_13382:FAff port map(x=>p(317)(117),y=>p(318)(117),Cin=>p(319)(117),clock=>clock,reset=>reset,s=>p(341)(117),cout=>p(342)(118));
FA_ff_13383:FAff port map(x=>p(317)(118),y=>p(318)(118),Cin=>p(319)(118),clock=>clock,reset=>reset,s=>p(341)(118),cout=>p(342)(119));
FA_ff_13384:FAff port map(x=>p(317)(119),y=>p(318)(119),Cin=>p(319)(119),clock=>clock,reset=>reset,s=>p(341)(119),cout=>p(342)(120));
FA_ff_13385:FAff port map(x=>p(317)(120),y=>p(318)(120),Cin=>p(319)(120),clock=>clock,reset=>reset,s=>p(341)(120),cout=>p(342)(121));
FA_ff_13386:FAff port map(x=>p(317)(121),y=>p(318)(121),Cin=>p(319)(121),clock=>clock,reset=>reset,s=>p(341)(121),cout=>p(342)(122));
FA_ff_13387:FAff port map(x=>p(317)(122),y=>p(318)(122),Cin=>p(319)(122),clock=>clock,reset=>reset,s=>p(341)(122),cout=>p(342)(123));
FA_ff_13388:FAff port map(x=>p(317)(123),y=>p(318)(123),Cin=>p(319)(123),clock=>clock,reset=>reset,s=>p(341)(123),cout=>p(342)(124));
FA_ff_13389:FAff port map(x=>p(317)(124),y=>p(318)(124),Cin=>p(319)(124),clock=>clock,reset=>reset,s=>p(341)(124),cout=>p(342)(125));
FA_ff_13390:FAff port map(x=>p(317)(125),y=>p(318)(125),Cin=>p(319)(125),clock=>clock,reset=>reset,s=>p(341)(125),cout=>p(342)(126));
FA_ff_13391:FAff port map(x=>p(317)(126),y=>p(318)(126),Cin=>p(319)(126),clock=>clock,reset=>reset,s=>p(341)(126),cout=>p(342)(127));
FA_ff_13392:FAff port map(x=>p(317)(127),y=>p(318)(127),Cin=>p(319)(127),clock=>clock,reset=>reset,s=>p(341)(127),cout=>p(342)(128));
FA_ff_13393:FAff port map(x=>p(317)(128),y=>p(318)(128),Cin=>p(319)(128),clock=>clock,reset=>reset,s=>p(341)(128),cout=>p(342)(129));
FA_ff_13394:FAff port map(x=>p(317)(129),y=>p(318)(129),Cin=>p(319)(129),clock=>clock,reset=>reset,s=>p(341)(129),cout=>p(342)(130));
p(341)(130)<=p(318)(130);
p(343)(0)<=p(321)(0);
HA_ff_81:HAff port map(x=>p(320)(1),y=>p(321)(1),clock=>clock,reset=>reset,s=>p(343)(1),c=>p(344)(2));
FA_ff_13395:FAff port map(x=>p(320)(2),y=>p(321)(2),Cin=>p(322)(2),clock=>clock,reset=>reset,s=>p(343)(2),cout=>p(344)(3));
FA_ff_13396:FAff port map(x=>p(320)(3),y=>p(321)(3),Cin=>p(322)(3),clock=>clock,reset=>reset,s=>p(343)(3),cout=>p(344)(4));
FA_ff_13397:FAff port map(x=>p(320)(4),y=>p(321)(4),Cin=>p(322)(4),clock=>clock,reset=>reset,s=>p(343)(4),cout=>p(344)(5));
FA_ff_13398:FAff port map(x=>p(320)(5),y=>p(321)(5),Cin=>p(322)(5),clock=>clock,reset=>reset,s=>p(343)(5),cout=>p(344)(6));
FA_ff_13399:FAff port map(x=>p(320)(6),y=>p(321)(6),Cin=>p(322)(6),clock=>clock,reset=>reset,s=>p(343)(6),cout=>p(344)(7));
FA_ff_13400:FAff port map(x=>p(320)(7),y=>p(321)(7),Cin=>p(322)(7),clock=>clock,reset=>reset,s=>p(343)(7),cout=>p(344)(8));
FA_ff_13401:FAff port map(x=>p(320)(8),y=>p(321)(8),Cin=>p(322)(8),clock=>clock,reset=>reset,s=>p(343)(8),cout=>p(344)(9));
FA_ff_13402:FAff port map(x=>p(320)(9),y=>p(321)(9),Cin=>p(322)(9),clock=>clock,reset=>reset,s=>p(343)(9),cout=>p(344)(10));
FA_ff_13403:FAff port map(x=>p(320)(10),y=>p(321)(10),Cin=>p(322)(10),clock=>clock,reset=>reset,s=>p(343)(10),cout=>p(344)(11));
FA_ff_13404:FAff port map(x=>p(320)(11),y=>p(321)(11),Cin=>p(322)(11),clock=>clock,reset=>reset,s=>p(343)(11),cout=>p(344)(12));
FA_ff_13405:FAff port map(x=>p(320)(12),y=>p(321)(12),Cin=>p(322)(12),clock=>clock,reset=>reset,s=>p(343)(12),cout=>p(344)(13));
FA_ff_13406:FAff port map(x=>p(320)(13),y=>p(321)(13),Cin=>p(322)(13),clock=>clock,reset=>reset,s=>p(343)(13),cout=>p(344)(14));
FA_ff_13407:FAff port map(x=>p(320)(14),y=>p(321)(14),Cin=>p(322)(14),clock=>clock,reset=>reset,s=>p(343)(14),cout=>p(344)(15));
FA_ff_13408:FAff port map(x=>p(320)(15),y=>p(321)(15),Cin=>p(322)(15),clock=>clock,reset=>reset,s=>p(343)(15),cout=>p(344)(16));
FA_ff_13409:FAff port map(x=>p(320)(16),y=>p(321)(16),Cin=>p(322)(16),clock=>clock,reset=>reset,s=>p(343)(16),cout=>p(344)(17));
FA_ff_13410:FAff port map(x=>p(320)(17),y=>p(321)(17),Cin=>p(322)(17),clock=>clock,reset=>reset,s=>p(343)(17),cout=>p(344)(18));
FA_ff_13411:FAff port map(x=>p(320)(18),y=>p(321)(18),Cin=>p(322)(18),clock=>clock,reset=>reset,s=>p(343)(18),cout=>p(344)(19));
FA_ff_13412:FAff port map(x=>p(320)(19),y=>p(321)(19),Cin=>p(322)(19),clock=>clock,reset=>reset,s=>p(343)(19),cout=>p(344)(20));
FA_ff_13413:FAff port map(x=>p(320)(20),y=>p(321)(20),Cin=>p(322)(20),clock=>clock,reset=>reset,s=>p(343)(20),cout=>p(344)(21));
FA_ff_13414:FAff port map(x=>p(320)(21),y=>p(321)(21),Cin=>p(322)(21),clock=>clock,reset=>reset,s=>p(343)(21),cout=>p(344)(22));
FA_ff_13415:FAff port map(x=>p(320)(22),y=>p(321)(22),Cin=>p(322)(22),clock=>clock,reset=>reset,s=>p(343)(22),cout=>p(344)(23));
FA_ff_13416:FAff port map(x=>p(320)(23),y=>p(321)(23),Cin=>p(322)(23),clock=>clock,reset=>reset,s=>p(343)(23),cout=>p(344)(24));
FA_ff_13417:FAff port map(x=>p(320)(24),y=>p(321)(24),Cin=>p(322)(24),clock=>clock,reset=>reset,s=>p(343)(24),cout=>p(344)(25));
FA_ff_13418:FAff port map(x=>p(320)(25),y=>p(321)(25),Cin=>p(322)(25),clock=>clock,reset=>reset,s=>p(343)(25),cout=>p(344)(26));
FA_ff_13419:FAff port map(x=>p(320)(26),y=>p(321)(26),Cin=>p(322)(26),clock=>clock,reset=>reset,s=>p(343)(26),cout=>p(344)(27));
FA_ff_13420:FAff port map(x=>p(320)(27),y=>p(321)(27),Cin=>p(322)(27),clock=>clock,reset=>reset,s=>p(343)(27),cout=>p(344)(28));
FA_ff_13421:FAff port map(x=>p(320)(28),y=>p(321)(28),Cin=>p(322)(28),clock=>clock,reset=>reset,s=>p(343)(28),cout=>p(344)(29));
FA_ff_13422:FAff port map(x=>p(320)(29),y=>p(321)(29),Cin=>p(322)(29),clock=>clock,reset=>reset,s=>p(343)(29),cout=>p(344)(30));
FA_ff_13423:FAff port map(x=>p(320)(30),y=>p(321)(30),Cin=>p(322)(30),clock=>clock,reset=>reset,s=>p(343)(30),cout=>p(344)(31));
FA_ff_13424:FAff port map(x=>p(320)(31),y=>p(321)(31),Cin=>p(322)(31),clock=>clock,reset=>reset,s=>p(343)(31),cout=>p(344)(32));
FA_ff_13425:FAff port map(x=>p(320)(32),y=>p(321)(32),Cin=>p(322)(32),clock=>clock,reset=>reset,s=>p(343)(32),cout=>p(344)(33));
FA_ff_13426:FAff port map(x=>p(320)(33),y=>p(321)(33),Cin=>p(322)(33),clock=>clock,reset=>reset,s=>p(343)(33),cout=>p(344)(34));
FA_ff_13427:FAff port map(x=>p(320)(34),y=>p(321)(34),Cin=>p(322)(34),clock=>clock,reset=>reset,s=>p(343)(34),cout=>p(344)(35));
FA_ff_13428:FAff port map(x=>p(320)(35),y=>p(321)(35),Cin=>p(322)(35),clock=>clock,reset=>reset,s=>p(343)(35),cout=>p(344)(36));
FA_ff_13429:FAff port map(x=>p(320)(36),y=>p(321)(36),Cin=>p(322)(36),clock=>clock,reset=>reset,s=>p(343)(36),cout=>p(344)(37));
FA_ff_13430:FAff port map(x=>p(320)(37),y=>p(321)(37),Cin=>p(322)(37),clock=>clock,reset=>reset,s=>p(343)(37),cout=>p(344)(38));
FA_ff_13431:FAff port map(x=>p(320)(38),y=>p(321)(38),Cin=>p(322)(38),clock=>clock,reset=>reset,s=>p(343)(38),cout=>p(344)(39));
FA_ff_13432:FAff port map(x=>p(320)(39),y=>p(321)(39),Cin=>p(322)(39),clock=>clock,reset=>reset,s=>p(343)(39),cout=>p(344)(40));
FA_ff_13433:FAff port map(x=>p(320)(40),y=>p(321)(40),Cin=>p(322)(40),clock=>clock,reset=>reset,s=>p(343)(40),cout=>p(344)(41));
FA_ff_13434:FAff port map(x=>p(320)(41),y=>p(321)(41),Cin=>p(322)(41),clock=>clock,reset=>reset,s=>p(343)(41),cout=>p(344)(42));
FA_ff_13435:FAff port map(x=>p(320)(42),y=>p(321)(42),Cin=>p(322)(42),clock=>clock,reset=>reset,s=>p(343)(42),cout=>p(344)(43));
FA_ff_13436:FAff port map(x=>p(320)(43),y=>p(321)(43),Cin=>p(322)(43),clock=>clock,reset=>reset,s=>p(343)(43),cout=>p(344)(44));
FA_ff_13437:FAff port map(x=>p(320)(44),y=>p(321)(44),Cin=>p(322)(44),clock=>clock,reset=>reset,s=>p(343)(44),cout=>p(344)(45));
FA_ff_13438:FAff port map(x=>p(320)(45),y=>p(321)(45),Cin=>p(322)(45),clock=>clock,reset=>reset,s=>p(343)(45),cout=>p(344)(46));
FA_ff_13439:FAff port map(x=>p(320)(46),y=>p(321)(46),Cin=>p(322)(46),clock=>clock,reset=>reset,s=>p(343)(46),cout=>p(344)(47));
FA_ff_13440:FAff port map(x=>p(320)(47),y=>p(321)(47),Cin=>p(322)(47),clock=>clock,reset=>reset,s=>p(343)(47),cout=>p(344)(48));
FA_ff_13441:FAff port map(x=>p(320)(48),y=>p(321)(48),Cin=>p(322)(48),clock=>clock,reset=>reset,s=>p(343)(48),cout=>p(344)(49));
FA_ff_13442:FAff port map(x=>p(320)(49),y=>p(321)(49),Cin=>p(322)(49),clock=>clock,reset=>reset,s=>p(343)(49),cout=>p(344)(50));
FA_ff_13443:FAff port map(x=>p(320)(50),y=>p(321)(50),Cin=>p(322)(50),clock=>clock,reset=>reset,s=>p(343)(50),cout=>p(344)(51));
FA_ff_13444:FAff port map(x=>p(320)(51),y=>p(321)(51),Cin=>p(322)(51),clock=>clock,reset=>reset,s=>p(343)(51),cout=>p(344)(52));
FA_ff_13445:FAff port map(x=>p(320)(52),y=>p(321)(52),Cin=>p(322)(52),clock=>clock,reset=>reset,s=>p(343)(52),cout=>p(344)(53));
FA_ff_13446:FAff port map(x=>p(320)(53),y=>p(321)(53),Cin=>p(322)(53),clock=>clock,reset=>reset,s=>p(343)(53),cout=>p(344)(54));
FA_ff_13447:FAff port map(x=>p(320)(54),y=>p(321)(54),Cin=>p(322)(54),clock=>clock,reset=>reset,s=>p(343)(54),cout=>p(344)(55));
FA_ff_13448:FAff port map(x=>p(320)(55),y=>p(321)(55),Cin=>p(322)(55),clock=>clock,reset=>reset,s=>p(343)(55),cout=>p(344)(56));
FA_ff_13449:FAff port map(x=>p(320)(56),y=>p(321)(56),Cin=>p(322)(56),clock=>clock,reset=>reset,s=>p(343)(56),cout=>p(344)(57));
FA_ff_13450:FAff port map(x=>p(320)(57),y=>p(321)(57),Cin=>p(322)(57),clock=>clock,reset=>reset,s=>p(343)(57),cout=>p(344)(58));
FA_ff_13451:FAff port map(x=>p(320)(58),y=>p(321)(58),Cin=>p(322)(58),clock=>clock,reset=>reset,s=>p(343)(58),cout=>p(344)(59));
FA_ff_13452:FAff port map(x=>p(320)(59),y=>p(321)(59),Cin=>p(322)(59),clock=>clock,reset=>reset,s=>p(343)(59),cout=>p(344)(60));
FA_ff_13453:FAff port map(x=>p(320)(60),y=>p(321)(60),Cin=>p(322)(60),clock=>clock,reset=>reset,s=>p(343)(60),cout=>p(344)(61));
FA_ff_13454:FAff port map(x=>p(320)(61),y=>p(321)(61),Cin=>p(322)(61),clock=>clock,reset=>reset,s=>p(343)(61),cout=>p(344)(62));
FA_ff_13455:FAff port map(x=>p(320)(62),y=>p(321)(62),Cin=>p(322)(62),clock=>clock,reset=>reset,s=>p(343)(62),cout=>p(344)(63));
FA_ff_13456:FAff port map(x=>p(320)(63),y=>p(321)(63),Cin=>p(322)(63),clock=>clock,reset=>reset,s=>p(343)(63),cout=>p(344)(64));
FA_ff_13457:FAff port map(x=>p(320)(64),y=>p(321)(64),Cin=>p(322)(64),clock=>clock,reset=>reset,s=>p(343)(64),cout=>p(344)(65));
FA_ff_13458:FAff port map(x=>p(320)(65),y=>p(321)(65),Cin=>p(322)(65),clock=>clock,reset=>reset,s=>p(343)(65),cout=>p(344)(66));
FA_ff_13459:FAff port map(x=>p(320)(66),y=>p(321)(66),Cin=>p(322)(66),clock=>clock,reset=>reset,s=>p(343)(66),cout=>p(344)(67));
FA_ff_13460:FAff port map(x=>p(320)(67),y=>p(321)(67),Cin=>p(322)(67),clock=>clock,reset=>reset,s=>p(343)(67),cout=>p(344)(68));
FA_ff_13461:FAff port map(x=>p(320)(68),y=>p(321)(68),Cin=>p(322)(68),clock=>clock,reset=>reset,s=>p(343)(68),cout=>p(344)(69));
FA_ff_13462:FAff port map(x=>p(320)(69),y=>p(321)(69),Cin=>p(322)(69),clock=>clock,reset=>reset,s=>p(343)(69),cout=>p(344)(70));
FA_ff_13463:FAff port map(x=>p(320)(70),y=>p(321)(70),Cin=>p(322)(70),clock=>clock,reset=>reset,s=>p(343)(70),cout=>p(344)(71));
FA_ff_13464:FAff port map(x=>p(320)(71),y=>p(321)(71),Cin=>p(322)(71),clock=>clock,reset=>reset,s=>p(343)(71),cout=>p(344)(72));
FA_ff_13465:FAff port map(x=>p(320)(72),y=>p(321)(72),Cin=>p(322)(72),clock=>clock,reset=>reset,s=>p(343)(72),cout=>p(344)(73));
FA_ff_13466:FAff port map(x=>p(320)(73),y=>p(321)(73),Cin=>p(322)(73),clock=>clock,reset=>reset,s=>p(343)(73),cout=>p(344)(74));
FA_ff_13467:FAff port map(x=>p(320)(74),y=>p(321)(74),Cin=>p(322)(74),clock=>clock,reset=>reset,s=>p(343)(74),cout=>p(344)(75));
FA_ff_13468:FAff port map(x=>p(320)(75),y=>p(321)(75),Cin=>p(322)(75),clock=>clock,reset=>reset,s=>p(343)(75),cout=>p(344)(76));
FA_ff_13469:FAff port map(x=>p(320)(76),y=>p(321)(76),Cin=>p(322)(76),clock=>clock,reset=>reset,s=>p(343)(76),cout=>p(344)(77));
FA_ff_13470:FAff port map(x=>p(320)(77),y=>p(321)(77),Cin=>p(322)(77),clock=>clock,reset=>reset,s=>p(343)(77),cout=>p(344)(78));
FA_ff_13471:FAff port map(x=>p(320)(78),y=>p(321)(78),Cin=>p(322)(78),clock=>clock,reset=>reset,s=>p(343)(78),cout=>p(344)(79));
FA_ff_13472:FAff port map(x=>p(320)(79),y=>p(321)(79),Cin=>p(322)(79),clock=>clock,reset=>reset,s=>p(343)(79),cout=>p(344)(80));
FA_ff_13473:FAff port map(x=>p(320)(80),y=>p(321)(80),Cin=>p(322)(80),clock=>clock,reset=>reset,s=>p(343)(80),cout=>p(344)(81));
FA_ff_13474:FAff port map(x=>p(320)(81),y=>p(321)(81),Cin=>p(322)(81),clock=>clock,reset=>reset,s=>p(343)(81),cout=>p(344)(82));
FA_ff_13475:FAff port map(x=>p(320)(82),y=>p(321)(82),Cin=>p(322)(82),clock=>clock,reset=>reset,s=>p(343)(82),cout=>p(344)(83));
FA_ff_13476:FAff port map(x=>p(320)(83),y=>p(321)(83),Cin=>p(322)(83),clock=>clock,reset=>reset,s=>p(343)(83),cout=>p(344)(84));
FA_ff_13477:FAff port map(x=>p(320)(84),y=>p(321)(84),Cin=>p(322)(84),clock=>clock,reset=>reset,s=>p(343)(84),cout=>p(344)(85));
FA_ff_13478:FAff port map(x=>p(320)(85),y=>p(321)(85),Cin=>p(322)(85),clock=>clock,reset=>reset,s=>p(343)(85),cout=>p(344)(86));
FA_ff_13479:FAff port map(x=>p(320)(86),y=>p(321)(86),Cin=>p(322)(86),clock=>clock,reset=>reset,s=>p(343)(86),cout=>p(344)(87));
FA_ff_13480:FAff port map(x=>p(320)(87),y=>p(321)(87),Cin=>p(322)(87),clock=>clock,reset=>reset,s=>p(343)(87),cout=>p(344)(88));
FA_ff_13481:FAff port map(x=>p(320)(88),y=>p(321)(88),Cin=>p(322)(88),clock=>clock,reset=>reset,s=>p(343)(88),cout=>p(344)(89));
FA_ff_13482:FAff port map(x=>p(320)(89),y=>p(321)(89),Cin=>p(322)(89),clock=>clock,reset=>reset,s=>p(343)(89),cout=>p(344)(90));
FA_ff_13483:FAff port map(x=>p(320)(90),y=>p(321)(90),Cin=>p(322)(90),clock=>clock,reset=>reset,s=>p(343)(90),cout=>p(344)(91));
FA_ff_13484:FAff port map(x=>p(320)(91),y=>p(321)(91),Cin=>p(322)(91),clock=>clock,reset=>reset,s=>p(343)(91),cout=>p(344)(92));
FA_ff_13485:FAff port map(x=>p(320)(92),y=>p(321)(92),Cin=>p(322)(92),clock=>clock,reset=>reset,s=>p(343)(92),cout=>p(344)(93));
FA_ff_13486:FAff port map(x=>p(320)(93),y=>p(321)(93),Cin=>p(322)(93),clock=>clock,reset=>reset,s=>p(343)(93),cout=>p(344)(94));
FA_ff_13487:FAff port map(x=>p(320)(94),y=>p(321)(94),Cin=>p(322)(94),clock=>clock,reset=>reset,s=>p(343)(94),cout=>p(344)(95));
FA_ff_13488:FAff port map(x=>p(320)(95),y=>p(321)(95),Cin=>p(322)(95),clock=>clock,reset=>reset,s=>p(343)(95),cout=>p(344)(96));
FA_ff_13489:FAff port map(x=>p(320)(96),y=>p(321)(96),Cin=>p(322)(96),clock=>clock,reset=>reset,s=>p(343)(96),cout=>p(344)(97));
FA_ff_13490:FAff port map(x=>p(320)(97),y=>p(321)(97),Cin=>p(322)(97),clock=>clock,reset=>reset,s=>p(343)(97),cout=>p(344)(98));
FA_ff_13491:FAff port map(x=>p(320)(98),y=>p(321)(98),Cin=>p(322)(98),clock=>clock,reset=>reset,s=>p(343)(98),cout=>p(344)(99));
FA_ff_13492:FAff port map(x=>p(320)(99),y=>p(321)(99),Cin=>p(322)(99),clock=>clock,reset=>reset,s=>p(343)(99),cout=>p(344)(100));
FA_ff_13493:FAff port map(x=>p(320)(100),y=>p(321)(100),Cin=>p(322)(100),clock=>clock,reset=>reset,s=>p(343)(100),cout=>p(344)(101));
FA_ff_13494:FAff port map(x=>p(320)(101),y=>p(321)(101),Cin=>p(322)(101),clock=>clock,reset=>reset,s=>p(343)(101),cout=>p(344)(102));
FA_ff_13495:FAff port map(x=>p(320)(102),y=>p(321)(102),Cin=>p(322)(102),clock=>clock,reset=>reset,s=>p(343)(102),cout=>p(344)(103));
FA_ff_13496:FAff port map(x=>p(320)(103),y=>p(321)(103),Cin=>p(322)(103),clock=>clock,reset=>reset,s=>p(343)(103),cout=>p(344)(104));
FA_ff_13497:FAff port map(x=>p(320)(104),y=>p(321)(104),Cin=>p(322)(104),clock=>clock,reset=>reset,s=>p(343)(104),cout=>p(344)(105));
FA_ff_13498:FAff port map(x=>p(320)(105),y=>p(321)(105),Cin=>p(322)(105),clock=>clock,reset=>reset,s=>p(343)(105),cout=>p(344)(106));
FA_ff_13499:FAff port map(x=>p(320)(106),y=>p(321)(106),Cin=>p(322)(106),clock=>clock,reset=>reset,s=>p(343)(106),cout=>p(344)(107));
FA_ff_13500:FAff port map(x=>p(320)(107),y=>p(321)(107),Cin=>p(322)(107),clock=>clock,reset=>reset,s=>p(343)(107),cout=>p(344)(108));
FA_ff_13501:FAff port map(x=>p(320)(108),y=>p(321)(108),Cin=>p(322)(108),clock=>clock,reset=>reset,s=>p(343)(108),cout=>p(344)(109));
FA_ff_13502:FAff port map(x=>p(320)(109),y=>p(321)(109),Cin=>p(322)(109),clock=>clock,reset=>reset,s=>p(343)(109),cout=>p(344)(110));
FA_ff_13503:FAff port map(x=>p(320)(110),y=>p(321)(110),Cin=>p(322)(110),clock=>clock,reset=>reset,s=>p(343)(110),cout=>p(344)(111));
FA_ff_13504:FAff port map(x=>p(320)(111),y=>p(321)(111),Cin=>p(322)(111),clock=>clock,reset=>reset,s=>p(343)(111),cout=>p(344)(112));
FA_ff_13505:FAff port map(x=>p(320)(112),y=>p(321)(112),Cin=>p(322)(112),clock=>clock,reset=>reset,s=>p(343)(112),cout=>p(344)(113));
FA_ff_13506:FAff port map(x=>p(320)(113),y=>p(321)(113),Cin=>p(322)(113),clock=>clock,reset=>reset,s=>p(343)(113),cout=>p(344)(114));
FA_ff_13507:FAff port map(x=>p(320)(114),y=>p(321)(114),Cin=>p(322)(114),clock=>clock,reset=>reset,s=>p(343)(114),cout=>p(344)(115));
FA_ff_13508:FAff port map(x=>p(320)(115),y=>p(321)(115),Cin=>p(322)(115),clock=>clock,reset=>reset,s=>p(343)(115),cout=>p(344)(116));
FA_ff_13509:FAff port map(x=>p(320)(116),y=>p(321)(116),Cin=>p(322)(116),clock=>clock,reset=>reset,s=>p(343)(116),cout=>p(344)(117));
FA_ff_13510:FAff port map(x=>p(320)(117),y=>p(321)(117),Cin=>p(322)(117),clock=>clock,reset=>reset,s=>p(343)(117),cout=>p(344)(118));
FA_ff_13511:FAff port map(x=>p(320)(118),y=>p(321)(118),Cin=>p(322)(118),clock=>clock,reset=>reset,s=>p(343)(118),cout=>p(344)(119));
FA_ff_13512:FAff port map(x=>p(320)(119),y=>p(321)(119),Cin=>p(322)(119),clock=>clock,reset=>reset,s=>p(343)(119),cout=>p(344)(120));
FA_ff_13513:FAff port map(x=>p(320)(120),y=>p(321)(120),Cin=>p(322)(120),clock=>clock,reset=>reset,s=>p(343)(120),cout=>p(344)(121));
FA_ff_13514:FAff port map(x=>p(320)(121),y=>p(321)(121),Cin=>p(322)(121),clock=>clock,reset=>reset,s=>p(343)(121),cout=>p(344)(122));
FA_ff_13515:FAff port map(x=>p(320)(122),y=>p(321)(122),Cin=>p(322)(122),clock=>clock,reset=>reset,s=>p(343)(122),cout=>p(344)(123));
FA_ff_13516:FAff port map(x=>p(320)(123),y=>p(321)(123),Cin=>p(322)(123),clock=>clock,reset=>reset,s=>p(343)(123),cout=>p(344)(124));
FA_ff_13517:FAff port map(x=>p(320)(124),y=>p(321)(124),Cin=>p(322)(124),clock=>clock,reset=>reset,s=>p(343)(124),cout=>p(344)(125));
FA_ff_13518:FAff port map(x=>p(320)(125),y=>p(321)(125),Cin=>p(322)(125),clock=>clock,reset=>reset,s=>p(343)(125),cout=>p(344)(126));
FA_ff_13519:FAff port map(x=>p(320)(126),y=>p(321)(126),Cin=>p(322)(126),clock=>clock,reset=>reset,s=>p(343)(126),cout=>p(344)(127));
FA_ff_13520:FAff port map(x=>p(320)(127),y=>p(321)(127),Cin=>p(322)(127),clock=>clock,reset=>reset,s=>p(343)(127),cout=>p(344)(128));
FA_ff_13521:FAff port map(x=>p(320)(128),y=>p(321)(128),Cin=>p(322)(128),clock=>clock,reset=>reset,s=>p(343)(128),cout=>p(344)(129));
FA_ff_13522:FAff port map(x=>p(320)(129),y=>p(321)(129),Cin=>p(322)(129),clock=>clock,reset=>reset,s=>p(343)(129),cout=>p(344)(130));
HA_ff_82:HAff port map(x=>p(320)(130),y=>p(322)(130),clock=>clock,reset=>reset,s=>p(343)(130),c=>p(344)(131));
HA_ff_83:HAff port map(x=>p(323)(0),y=>p(325)(0),clock=>clock,reset=>reset,s=>p(345)(0),c=>p(346)(1));
FA_ff_13523:FAff port map(x=>p(323)(1),y=>p(324)(1),Cin=>p(325)(1),clock=>clock,reset=>reset,s=>p(345)(1),cout=>p(346)(2));
FA_ff_13524:FAff port map(x=>p(323)(2),y=>p(324)(2),Cin=>p(325)(2),clock=>clock,reset=>reset,s=>p(345)(2),cout=>p(346)(3));
FA_ff_13525:FAff port map(x=>p(323)(3),y=>p(324)(3),Cin=>p(325)(3),clock=>clock,reset=>reset,s=>p(345)(3),cout=>p(346)(4));
FA_ff_13526:FAff port map(x=>p(323)(4),y=>p(324)(4),Cin=>p(325)(4),clock=>clock,reset=>reset,s=>p(345)(4),cout=>p(346)(5));
FA_ff_13527:FAff port map(x=>p(323)(5),y=>p(324)(5),Cin=>p(325)(5),clock=>clock,reset=>reset,s=>p(345)(5),cout=>p(346)(6));
FA_ff_13528:FAff port map(x=>p(323)(6),y=>p(324)(6),Cin=>p(325)(6),clock=>clock,reset=>reset,s=>p(345)(6),cout=>p(346)(7));
FA_ff_13529:FAff port map(x=>p(323)(7),y=>p(324)(7),Cin=>p(325)(7),clock=>clock,reset=>reset,s=>p(345)(7),cout=>p(346)(8));
FA_ff_13530:FAff port map(x=>p(323)(8),y=>p(324)(8),Cin=>p(325)(8),clock=>clock,reset=>reset,s=>p(345)(8),cout=>p(346)(9));
FA_ff_13531:FAff port map(x=>p(323)(9),y=>p(324)(9),Cin=>p(325)(9),clock=>clock,reset=>reset,s=>p(345)(9),cout=>p(346)(10));
FA_ff_13532:FAff port map(x=>p(323)(10),y=>p(324)(10),Cin=>p(325)(10),clock=>clock,reset=>reset,s=>p(345)(10),cout=>p(346)(11));
FA_ff_13533:FAff port map(x=>p(323)(11),y=>p(324)(11),Cin=>p(325)(11),clock=>clock,reset=>reset,s=>p(345)(11),cout=>p(346)(12));
FA_ff_13534:FAff port map(x=>p(323)(12),y=>p(324)(12),Cin=>p(325)(12),clock=>clock,reset=>reset,s=>p(345)(12),cout=>p(346)(13));
FA_ff_13535:FAff port map(x=>p(323)(13),y=>p(324)(13),Cin=>p(325)(13),clock=>clock,reset=>reset,s=>p(345)(13),cout=>p(346)(14));
FA_ff_13536:FAff port map(x=>p(323)(14),y=>p(324)(14),Cin=>p(325)(14),clock=>clock,reset=>reset,s=>p(345)(14),cout=>p(346)(15));
FA_ff_13537:FAff port map(x=>p(323)(15),y=>p(324)(15),Cin=>p(325)(15),clock=>clock,reset=>reset,s=>p(345)(15),cout=>p(346)(16));
FA_ff_13538:FAff port map(x=>p(323)(16),y=>p(324)(16),Cin=>p(325)(16),clock=>clock,reset=>reset,s=>p(345)(16),cout=>p(346)(17));
FA_ff_13539:FAff port map(x=>p(323)(17),y=>p(324)(17),Cin=>p(325)(17),clock=>clock,reset=>reset,s=>p(345)(17),cout=>p(346)(18));
FA_ff_13540:FAff port map(x=>p(323)(18),y=>p(324)(18),Cin=>p(325)(18),clock=>clock,reset=>reset,s=>p(345)(18),cout=>p(346)(19));
FA_ff_13541:FAff port map(x=>p(323)(19),y=>p(324)(19),Cin=>p(325)(19),clock=>clock,reset=>reset,s=>p(345)(19),cout=>p(346)(20));
FA_ff_13542:FAff port map(x=>p(323)(20),y=>p(324)(20),Cin=>p(325)(20),clock=>clock,reset=>reset,s=>p(345)(20),cout=>p(346)(21));
FA_ff_13543:FAff port map(x=>p(323)(21),y=>p(324)(21),Cin=>p(325)(21),clock=>clock,reset=>reset,s=>p(345)(21),cout=>p(346)(22));
FA_ff_13544:FAff port map(x=>p(323)(22),y=>p(324)(22),Cin=>p(325)(22),clock=>clock,reset=>reset,s=>p(345)(22),cout=>p(346)(23));
FA_ff_13545:FAff port map(x=>p(323)(23),y=>p(324)(23),Cin=>p(325)(23),clock=>clock,reset=>reset,s=>p(345)(23),cout=>p(346)(24));
FA_ff_13546:FAff port map(x=>p(323)(24),y=>p(324)(24),Cin=>p(325)(24),clock=>clock,reset=>reset,s=>p(345)(24),cout=>p(346)(25));
FA_ff_13547:FAff port map(x=>p(323)(25),y=>p(324)(25),Cin=>p(325)(25),clock=>clock,reset=>reset,s=>p(345)(25),cout=>p(346)(26));
FA_ff_13548:FAff port map(x=>p(323)(26),y=>p(324)(26),Cin=>p(325)(26),clock=>clock,reset=>reset,s=>p(345)(26),cout=>p(346)(27));
FA_ff_13549:FAff port map(x=>p(323)(27),y=>p(324)(27),Cin=>p(325)(27),clock=>clock,reset=>reset,s=>p(345)(27),cout=>p(346)(28));
FA_ff_13550:FAff port map(x=>p(323)(28),y=>p(324)(28),Cin=>p(325)(28),clock=>clock,reset=>reset,s=>p(345)(28),cout=>p(346)(29));
FA_ff_13551:FAff port map(x=>p(323)(29),y=>p(324)(29),Cin=>p(325)(29),clock=>clock,reset=>reset,s=>p(345)(29),cout=>p(346)(30));
FA_ff_13552:FAff port map(x=>p(323)(30),y=>p(324)(30),Cin=>p(325)(30),clock=>clock,reset=>reset,s=>p(345)(30),cout=>p(346)(31));
FA_ff_13553:FAff port map(x=>p(323)(31),y=>p(324)(31),Cin=>p(325)(31),clock=>clock,reset=>reset,s=>p(345)(31),cout=>p(346)(32));
FA_ff_13554:FAff port map(x=>p(323)(32),y=>p(324)(32),Cin=>p(325)(32),clock=>clock,reset=>reset,s=>p(345)(32),cout=>p(346)(33));
FA_ff_13555:FAff port map(x=>p(323)(33),y=>p(324)(33),Cin=>p(325)(33),clock=>clock,reset=>reset,s=>p(345)(33),cout=>p(346)(34));
FA_ff_13556:FAff port map(x=>p(323)(34),y=>p(324)(34),Cin=>p(325)(34),clock=>clock,reset=>reset,s=>p(345)(34),cout=>p(346)(35));
FA_ff_13557:FAff port map(x=>p(323)(35),y=>p(324)(35),Cin=>p(325)(35),clock=>clock,reset=>reset,s=>p(345)(35),cout=>p(346)(36));
FA_ff_13558:FAff port map(x=>p(323)(36),y=>p(324)(36),Cin=>p(325)(36),clock=>clock,reset=>reset,s=>p(345)(36),cout=>p(346)(37));
FA_ff_13559:FAff port map(x=>p(323)(37),y=>p(324)(37),Cin=>p(325)(37),clock=>clock,reset=>reset,s=>p(345)(37),cout=>p(346)(38));
FA_ff_13560:FAff port map(x=>p(323)(38),y=>p(324)(38),Cin=>p(325)(38),clock=>clock,reset=>reset,s=>p(345)(38),cout=>p(346)(39));
FA_ff_13561:FAff port map(x=>p(323)(39),y=>p(324)(39),Cin=>p(325)(39),clock=>clock,reset=>reset,s=>p(345)(39),cout=>p(346)(40));
FA_ff_13562:FAff port map(x=>p(323)(40),y=>p(324)(40),Cin=>p(325)(40),clock=>clock,reset=>reset,s=>p(345)(40),cout=>p(346)(41));
FA_ff_13563:FAff port map(x=>p(323)(41),y=>p(324)(41),Cin=>p(325)(41),clock=>clock,reset=>reset,s=>p(345)(41),cout=>p(346)(42));
FA_ff_13564:FAff port map(x=>p(323)(42),y=>p(324)(42),Cin=>p(325)(42),clock=>clock,reset=>reset,s=>p(345)(42),cout=>p(346)(43));
FA_ff_13565:FAff port map(x=>p(323)(43),y=>p(324)(43),Cin=>p(325)(43),clock=>clock,reset=>reset,s=>p(345)(43),cout=>p(346)(44));
FA_ff_13566:FAff port map(x=>p(323)(44),y=>p(324)(44),Cin=>p(325)(44),clock=>clock,reset=>reset,s=>p(345)(44),cout=>p(346)(45));
FA_ff_13567:FAff port map(x=>p(323)(45),y=>p(324)(45),Cin=>p(325)(45),clock=>clock,reset=>reset,s=>p(345)(45),cout=>p(346)(46));
FA_ff_13568:FAff port map(x=>p(323)(46),y=>p(324)(46),Cin=>p(325)(46),clock=>clock,reset=>reset,s=>p(345)(46),cout=>p(346)(47));
FA_ff_13569:FAff port map(x=>p(323)(47),y=>p(324)(47),Cin=>p(325)(47),clock=>clock,reset=>reset,s=>p(345)(47),cout=>p(346)(48));
FA_ff_13570:FAff port map(x=>p(323)(48),y=>p(324)(48),Cin=>p(325)(48),clock=>clock,reset=>reset,s=>p(345)(48),cout=>p(346)(49));
FA_ff_13571:FAff port map(x=>p(323)(49),y=>p(324)(49),Cin=>p(325)(49),clock=>clock,reset=>reset,s=>p(345)(49),cout=>p(346)(50));
FA_ff_13572:FAff port map(x=>p(323)(50),y=>p(324)(50),Cin=>p(325)(50),clock=>clock,reset=>reset,s=>p(345)(50),cout=>p(346)(51));
FA_ff_13573:FAff port map(x=>p(323)(51),y=>p(324)(51),Cin=>p(325)(51),clock=>clock,reset=>reset,s=>p(345)(51),cout=>p(346)(52));
FA_ff_13574:FAff port map(x=>p(323)(52),y=>p(324)(52),Cin=>p(325)(52),clock=>clock,reset=>reset,s=>p(345)(52),cout=>p(346)(53));
FA_ff_13575:FAff port map(x=>p(323)(53),y=>p(324)(53),Cin=>p(325)(53),clock=>clock,reset=>reset,s=>p(345)(53),cout=>p(346)(54));
FA_ff_13576:FAff port map(x=>p(323)(54),y=>p(324)(54),Cin=>p(325)(54),clock=>clock,reset=>reset,s=>p(345)(54),cout=>p(346)(55));
FA_ff_13577:FAff port map(x=>p(323)(55),y=>p(324)(55),Cin=>p(325)(55),clock=>clock,reset=>reset,s=>p(345)(55),cout=>p(346)(56));
FA_ff_13578:FAff port map(x=>p(323)(56),y=>p(324)(56),Cin=>p(325)(56),clock=>clock,reset=>reset,s=>p(345)(56),cout=>p(346)(57));
FA_ff_13579:FAff port map(x=>p(323)(57),y=>p(324)(57),Cin=>p(325)(57),clock=>clock,reset=>reset,s=>p(345)(57),cout=>p(346)(58));
FA_ff_13580:FAff port map(x=>p(323)(58),y=>p(324)(58),Cin=>p(325)(58),clock=>clock,reset=>reset,s=>p(345)(58),cout=>p(346)(59));
FA_ff_13581:FAff port map(x=>p(323)(59),y=>p(324)(59),Cin=>p(325)(59),clock=>clock,reset=>reset,s=>p(345)(59),cout=>p(346)(60));
FA_ff_13582:FAff port map(x=>p(323)(60),y=>p(324)(60),Cin=>p(325)(60),clock=>clock,reset=>reset,s=>p(345)(60),cout=>p(346)(61));
FA_ff_13583:FAff port map(x=>p(323)(61),y=>p(324)(61),Cin=>p(325)(61),clock=>clock,reset=>reset,s=>p(345)(61),cout=>p(346)(62));
FA_ff_13584:FAff port map(x=>p(323)(62),y=>p(324)(62),Cin=>p(325)(62),clock=>clock,reset=>reset,s=>p(345)(62),cout=>p(346)(63));
FA_ff_13585:FAff port map(x=>p(323)(63),y=>p(324)(63),Cin=>p(325)(63),clock=>clock,reset=>reset,s=>p(345)(63),cout=>p(346)(64));
FA_ff_13586:FAff port map(x=>p(323)(64),y=>p(324)(64),Cin=>p(325)(64),clock=>clock,reset=>reset,s=>p(345)(64),cout=>p(346)(65));
FA_ff_13587:FAff port map(x=>p(323)(65),y=>p(324)(65),Cin=>p(325)(65),clock=>clock,reset=>reset,s=>p(345)(65),cout=>p(346)(66));
FA_ff_13588:FAff port map(x=>p(323)(66),y=>p(324)(66),Cin=>p(325)(66),clock=>clock,reset=>reset,s=>p(345)(66),cout=>p(346)(67));
FA_ff_13589:FAff port map(x=>p(323)(67),y=>p(324)(67),Cin=>p(325)(67),clock=>clock,reset=>reset,s=>p(345)(67),cout=>p(346)(68));
FA_ff_13590:FAff port map(x=>p(323)(68),y=>p(324)(68),Cin=>p(325)(68),clock=>clock,reset=>reset,s=>p(345)(68),cout=>p(346)(69));
FA_ff_13591:FAff port map(x=>p(323)(69),y=>p(324)(69),Cin=>p(325)(69),clock=>clock,reset=>reset,s=>p(345)(69),cout=>p(346)(70));
FA_ff_13592:FAff port map(x=>p(323)(70),y=>p(324)(70),Cin=>p(325)(70),clock=>clock,reset=>reset,s=>p(345)(70),cout=>p(346)(71));
FA_ff_13593:FAff port map(x=>p(323)(71),y=>p(324)(71),Cin=>p(325)(71),clock=>clock,reset=>reset,s=>p(345)(71),cout=>p(346)(72));
FA_ff_13594:FAff port map(x=>p(323)(72),y=>p(324)(72),Cin=>p(325)(72),clock=>clock,reset=>reset,s=>p(345)(72),cout=>p(346)(73));
FA_ff_13595:FAff port map(x=>p(323)(73),y=>p(324)(73),Cin=>p(325)(73),clock=>clock,reset=>reset,s=>p(345)(73),cout=>p(346)(74));
FA_ff_13596:FAff port map(x=>p(323)(74),y=>p(324)(74),Cin=>p(325)(74),clock=>clock,reset=>reset,s=>p(345)(74),cout=>p(346)(75));
FA_ff_13597:FAff port map(x=>p(323)(75),y=>p(324)(75),Cin=>p(325)(75),clock=>clock,reset=>reset,s=>p(345)(75),cout=>p(346)(76));
FA_ff_13598:FAff port map(x=>p(323)(76),y=>p(324)(76),Cin=>p(325)(76),clock=>clock,reset=>reset,s=>p(345)(76),cout=>p(346)(77));
FA_ff_13599:FAff port map(x=>p(323)(77),y=>p(324)(77),Cin=>p(325)(77),clock=>clock,reset=>reset,s=>p(345)(77),cout=>p(346)(78));
FA_ff_13600:FAff port map(x=>p(323)(78),y=>p(324)(78),Cin=>p(325)(78),clock=>clock,reset=>reset,s=>p(345)(78),cout=>p(346)(79));
FA_ff_13601:FAff port map(x=>p(323)(79),y=>p(324)(79),Cin=>p(325)(79),clock=>clock,reset=>reset,s=>p(345)(79),cout=>p(346)(80));
FA_ff_13602:FAff port map(x=>p(323)(80),y=>p(324)(80),Cin=>p(325)(80),clock=>clock,reset=>reset,s=>p(345)(80),cout=>p(346)(81));
FA_ff_13603:FAff port map(x=>p(323)(81),y=>p(324)(81),Cin=>p(325)(81),clock=>clock,reset=>reset,s=>p(345)(81),cout=>p(346)(82));
FA_ff_13604:FAff port map(x=>p(323)(82),y=>p(324)(82),Cin=>p(325)(82),clock=>clock,reset=>reset,s=>p(345)(82),cout=>p(346)(83));
FA_ff_13605:FAff port map(x=>p(323)(83),y=>p(324)(83),Cin=>p(325)(83),clock=>clock,reset=>reset,s=>p(345)(83),cout=>p(346)(84));
FA_ff_13606:FAff port map(x=>p(323)(84),y=>p(324)(84),Cin=>p(325)(84),clock=>clock,reset=>reset,s=>p(345)(84),cout=>p(346)(85));
FA_ff_13607:FAff port map(x=>p(323)(85),y=>p(324)(85),Cin=>p(325)(85),clock=>clock,reset=>reset,s=>p(345)(85),cout=>p(346)(86));
FA_ff_13608:FAff port map(x=>p(323)(86),y=>p(324)(86),Cin=>p(325)(86),clock=>clock,reset=>reset,s=>p(345)(86),cout=>p(346)(87));
FA_ff_13609:FAff port map(x=>p(323)(87),y=>p(324)(87),Cin=>p(325)(87),clock=>clock,reset=>reset,s=>p(345)(87),cout=>p(346)(88));
FA_ff_13610:FAff port map(x=>p(323)(88),y=>p(324)(88),Cin=>p(325)(88),clock=>clock,reset=>reset,s=>p(345)(88),cout=>p(346)(89));
FA_ff_13611:FAff port map(x=>p(323)(89),y=>p(324)(89),Cin=>p(325)(89),clock=>clock,reset=>reset,s=>p(345)(89),cout=>p(346)(90));
FA_ff_13612:FAff port map(x=>p(323)(90),y=>p(324)(90),Cin=>p(325)(90),clock=>clock,reset=>reset,s=>p(345)(90),cout=>p(346)(91));
FA_ff_13613:FAff port map(x=>p(323)(91),y=>p(324)(91),Cin=>p(325)(91),clock=>clock,reset=>reset,s=>p(345)(91),cout=>p(346)(92));
FA_ff_13614:FAff port map(x=>p(323)(92),y=>p(324)(92),Cin=>p(325)(92),clock=>clock,reset=>reset,s=>p(345)(92),cout=>p(346)(93));
FA_ff_13615:FAff port map(x=>p(323)(93),y=>p(324)(93),Cin=>p(325)(93),clock=>clock,reset=>reset,s=>p(345)(93),cout=>p(346)(94));
FA_ff_13616:FAff port map(x=>p(323)(94),y=>p(324)(94),Cin=>p(325)(94),clock=>clock,reset=>reset,s=>p(345)(94),cout=>p(346)(95));
FA_ff_13617:FAff port map(x=>p(323)(95),y=>p(324)(95),Cin=>p(325)(95),clock=>clock,reset=>reset,s=>p(345)(95),cout=>p(346)(96));
FA_ff_13618:FAff port map(x=>p(323)(96),y=>p(324)(96),Cin=>p(325)(96),clock=>clock,reset=>reset,s=>p(345)(96),cout=>p(346)(97));
FA_ff_13619:FAff port map(x=>p(323)(97),y=>p(324)(97),Cin=>p(325)(97),clock=>clock,reset=>reset,s=>p(345)(97),cout=>p(346)(98));
FA_ff_13620:FAff port map(x=>p(323)(98),y=>p(324)(98),Cin=>p(325)(98),clock=>clock,reset=>reset,s=>p(345)(98),cout=>p(346)(99));
FA_ff_13621:FAff port map(x=>p(323)(99),y=>p(324)(99),Cin=>p(325)(99),clock=>clock,reset=>reset,s=>p(345)(99),cout=>p(346)(100));
FA_ff_13622:FAff port map(x=>p(323)(100),y=>p(324)(100),Cin=>p(325)(100),clock=>clock,reset=>reset,s=>p(345)(100),cout=>p(346)(101));
FA_ff_13623:FAff port map(x=>p(323)(101),y=>p(324)(101),Cin=>p(325)(101),clock=>clock,reset=>reset,s=>p(345)(101),cout=>p(346)(102));
FA_ff_13624:FAff port map(x=>p(323)(102),y=>p(324)(102),Cin=>p(325)(102),clock=>clock,reset=>reset,s=>p(345)(102),cout=>p(346)(103));
FA_ff_13625:FAff port map(x=>p(323)(103),y=>p(324)(103),Cin=>p(325)(103),clock=>clock,reset=>reset,s=>p(345)(103),cout=>p(346)(104));
FA_ff_13626:FAff port map(x=>p(323)(104),y=>p(324)(104),Cin=>p(325)(104),clock=>clock,reset=>reset,s=>p(345)(104),cout=>p(346)(105));
FA_ff_13627:FAff port map(x=>p(323)(105),y=>p(324)(105),Cin=>p(325)(105),clock=>clock,reset=>reset,s=>p(345)(105),cout=>p(346)(106));
FA_ff_13628:FAff port map(x=>p(323)(106),y=>p(324)(106),Cin=>p(325)(106),clock=>clock,reset=>reset,s=>p(345)(106),cout=>p(346)(107));
FA_ff_13629:FAff port map(x=>p(323)(107),y=>p(324)(107),Cin=>p(325)(107),clock=>clock,reset=>reset,s=>p(345)(107),cout=>p(346)(108));
FA_ff_13630:FAff port map(x=>p(323)(108),y=>p(324)(108),Cin=>p(325)(108),clock=>clock,reset=>reset,s=>p(345)(108),cout=>p(346)(109));
FA_ff_13631:FAff port map(x=>p(323)(109),y=>p(324)(109),Cin=>p(325)(109),clock=>clock,reset=>reset,s=>p(345)(109),cout=>p(346)(110));
FA_ff_13632:FAff port map(x=>p(323)(110),y=>p(324)(110),Cin=>p(325)(110),clock=>clock,reset=>reset,s=>p(345)(110),cout=>p(346)(111));
FA_ff_13633:FAff port map(x=>p(323)(111),y=>p(324)(111),Cin=>p(325)(111),clock=>clock,reset=>reset,s=>p(345)(111),cout=>p(346)(112));
FA_ff_13634:FAff port map(x=>p(323)(112),y=>p(324)(112),Cin=>p(325)(112),clock=>clock,reset=>reset,s=>p(345)(112),cout=>p(346)(113));
FA_ff_13635:FAff port map(x=>p(323)(113),y=>p(324)(113),Cin=>p(325)(113),clock=>clock,reset=>reset,s=>p(345)(113),cout=>p(346)(114));
FA_ff_13636:FAff port map(x=>p(323)(114),y=>p(324)(114),Cin=>p(325)(114),clock=>clock,reset=>reset,s=>p(345)(114),cout=>p(346)(115));
FA_ff_13637:FAff port map(x=>p(323)(115),y=>p(324)(115),Cin=>p(325)(115),clock=>clock,reset=>reset,s=>p(345)(115),cout=>p(346)(116));
FA_ff_13638:FAff port map(x=>p(323)(116),y=>p(324)(116),Cin=>p(325)(116),clock=>clock,reset=>reset,s=>p(345)(116),cout=>p(346)(117));
FA_ff_13639:FAff port map(x=>p(323)(117),y=>p(324)(117),Cin=>p(325)(117),clock=>clock,reset=>reset,s=>p(345)(117),cout=>p(346)(118));
FA_ff_13640:FAff port map(x=>p(323)(118),y=>p(324)(118),Cin=>p(325)(118),clock=>clock,reset=>reset,s=>p(345)(118),cout=>p(346)(119));
FA_ff_13641:FAff port map(x=>p(323)(119),y=>p(324)(119),Cin=>p(325)(119),clock=>clock,reset=>reset,s=>p(345)(119),cout=>p(346)(120));
FA_ff_13642:FAff port map(x=>p(323)(120),y=>p(324)(120),Cin=>p(325)(120),clock=>clock,reset=>reset,s=>p(345)(120),cout=>p(346)(121));
FA_ff_13643:FAff port map(x=>p(323)(121),y=>p(324)(121),Cin=>p(325)(121),clock=>clock,reset=>reset,s=>p(345)(121),cout=>p(346)(122));
FA_ff_13644:FAff port map(x=>p(323)(122),y=>p(324)(122),Cin=>p(325)(122),clock=>clock,reset=>reset,s=>p(345)(122),cout=>p(346)(123));
FA_ff_13645:FAff port map(x=>p(323)(123),y=>p(324)(123),Cin=>p(325)(123),clock=>clock,reset=>reset,s=>p(345)(123),cout=>p(346)(124));
FA_ff_13646:FAff port map(x=>p(323)(124),y=>p(324)(124),Cin=>p(325)(124),clock=>clock,reset=>reset,s=>p(345)(124),cout=>p(346)(125));
FA_ff_13647:FAff port map(x=>p(323)(125),y=>p(324)(125),Cin=>p(325)(125),clock=>clock,reset=>reset,s=>p(345)(125),cout=>p(346)(126));
FA_ff_13648:FAff port map(x=>p(323)(126),y=>p(324)(126),Cin=>p(325)(126),clock=>clock,reset=>reset,s=>p(345)(126),cout=>p(346)(127));
FA_ff_13649:FAff port map(x=>p(323)(127),y=>p(324)(127),Cin=>p(325)(127),clock=>clock,reset=>reset,s=>p(345)(127),cout=>p(346)(128));
FA_ff_13650:FAff port map(x=>p(323)(128),y=>p(324)(128),Cin=>p(325)(128),clock=>clock,reset=>reset,s=>p(345)(128),cout=>p(346)(129));
FA_ff_13651:FAff port map(x=>p(323)(129),y=>p(324)(129),Cin=>p(325)(129),clock=>clock,reset=>reset,s=>p(345)(129),cout=>p(346)(130));
p(345)(130)<=p(324)(130);
p(347)(0)<=p(327)(0);
HA_ff_84:HAff port map(x=>p(327)(1),y=>p(328)(1),clock=>clock,reset=>reset,s=>p(347)(1),c=>p(348)(2));
FA_ff_13652:FAff port map(x=>p(326)(2),y=>p(327)(2),Cin=>p(328)(2),clock=>clock,reset=>reset,s=>p(347)(2),cout=>p(348)(3));
FA_ff_13653:FAff port map(x=>p(326)(3),y=>p(327)(3),Cin=>p(328)(3),clock=>clock,reset=>reset,s=>p(347)(3),cout=>p(348)(4));
FA_ff_13654:FAff port map(x=>p(326)(4),y=>p(327)(4),Cin=>p(328)(4),clock=>clock,reset=>reset,s=>p(347)(4),cout=>p(348)(5));
FA_ff_13655:FAff port map(x=>p(326)(5),y=>p(327)(5),Cin=>p(328)(5),clock=>clock,reset=>reset,s=>p(347)(5),cout=>p(348)(6));
FA_ff_13656:FAff port map(x=>p(326)(6),y=>p(327)(6),Cin=>p(328)(6),clock=>clock,reset=>reset,s=>p(347)(6),cout=>p(348)(7));
FA_ff_13657:FAff port map(x=>p(326)(7),y=>p(327)(7),Cin=>p(328)(7),clock=>clock,reset=>reset,s=>p(347)(7),cout=>p(348)(8));
FA_ff_13658:FAff port map(x=>p(326)(8),y=>p(327)(8),Cin=>p(328)(8),clock=>clock,reset=>reset,s=>p(347)(8),cout=>p(348)(9));
FA_ff_13659:FAff port map(x=>p(326)(9),y=>p(327)(9),Cin=>p(328)(9),clock=>clock,reset=>reset,s=>p(347)(9),cout=>p(348)(10));
FA_ff_13660:FAff port map(x=>p(326)(10),y=>p(327)(10),Cin=>p(328)(10),clock=>clock,reset=>reset,s=>p(347)(10),cout=>p(348)(11));
FA_ff_13661:FAff port map(x=>p(326)(11),y=>p(327)(11),Cin=>p(328)(11),clock=>clock,reset=>reset,s=>p(347)(11),cout=>p(348)(12));
FA_ff_13662:FAff port map(x=>p(326)(12),y=>p(327)(12),Cin=>p(328)(12),clock=>clock,reset=>reset,s=>p(347)(12),cout=>p(348)(13));
FA_ff_13663:FAff port map(x=>p(326)(13),y=>p(327)(13),Cin=>p(328)(13),clock=>clock,reset=>reset,s=>p(347)(13),cout=>p(348)(14));
FA_ff_13664:FAff port map(x=>p(326)(14),y=>p(327)(14),Cin=>p(328)(14),clock=>clock,reset=>reset,s=>p(347)(14),cout=>p(348)(15));
FA_ff_13665:FAff port map(x=>p(326)(15),y=>p(327)(15),Cin=>p(328)(15),clock=>clock,reset=>reset,s=>p(347)(15),cout=>p(348)(16));
FA_ff_13666:FAff port map(x=>p(326)(16),y=>p(327)(16),Cin=>p(328)(16),clock=>clock,reset=>reset,s=>p(347)(16),cout=>p(348)(17));
FA_ff_13667:FAff port map(x=>p(326)(17),y=>p(327)(17),Cin=>p(328)(17),clock=>clock,reset=>reset,s=>p(347)(17),cout=>p(348)(18));
FA_ff_13668:FAff port map(x=>p(326)(18),y=>p(327)(18),Cin=>p(328)(18),clock=>clock,reset=>reset,s=>p(347)(18),cout=>p(348)(19));
FA_ff_13669:FAff port map(x=>p(326)(19),y=>p(327)(19),Cin=>p(328)(19),clock=>clock,reset=>reset,s=>p(347)(19),cout=>p(348)(20));
FA_ff_13670:FAff port map(x=>p(326)(20),y=>p(327)(20),Cin=>p(328)(20),clock=>clock,reset=>reset,s=>p(347)(20),cout=>p(348)(21));
FA_ff_13671:FAff port map(x=>p(326)(21),y=>p(327)(21),Cin=>p(328)(21),clock=>clock,reset=>reset,s=>p(347)(21),cout=>p(348)(22));
FA_ff_13672:FAff port map(x=>p(326)(22),y=>p(327)(22),Cin=>p(328)(22),clock=>clock,reset=>reset,s=>p(347)(22),cout=>p(348)(23));
FA_ff_13673:FAff port map(x=>p(326)(23),y=>p(327)(23),Cin=>p(328)(23),clock=>clock,reset=>reset,s=>p(347)(23),cout=>p(348)(24));
FA_ff_13674:FAff port map(x=>p(326)(24),y=>p(327)(24),Cin=>p(328)(24),clock=>clock,reset=>reset,s=>p(347)(24),cout=>p(348)(25));
FA_ff_13675:FAff port map(x=>p(326)(25),y=>p(327)(25),Cin=>p(328)(25),clock=>clock,reset=>reset,s=>p(347)(25),cout=>p(348)(26));
FA_ff_13676:FAff port map(x=>p(326)(26),y=>p(327)(26),Cin=>p(328)(26),clock=>clock,reset=>reset,s=>p(347)(26),cout=>p(348)(27));
FA_ff_13677:FAff port map(x=>p(326)(27),y=>p(327)(27),Cin=>p(328)(27),clock=>clock,reset=>reset,s=>p(347)(27),cout=>p(348)(28));
FA_ff_13678:FAff port map(x=>p(326)(28),y=>p(327)(28),Cin=>p(328)(28),clock=>clock,reset=>reset,s=>p(347)(28),cout=>p(348)(29));
FA_ff_13679:FAff port map(x=>p(326)(29),y=>p(327)(29),Cin=>p(328)(29),clock=>clock,reset=>reset,s=>p(347)(29),cout=>p(348)(30));
FA_ff_13680:FAff port map(x=>p(326)(30),y=>p(327)(30),Cin=>p(328)(30),clock=>clock,reset=>reset,s=>p(347)(30),cout=>p(348)(31));
FA_ff_13681:FAff port map(x=>p(326)(31),y=>p(327)(31),Cin=>p(328)(31),clock=>clock,reset=>reset,s=>p(347)(31),cout=>p(348)(32));
FA_ff_13682:FAff port map(x=>p(326)(32),y=>p(327)(32),Cin=>p(328)(32),clock=>clock,reset=>reset,s=>p(347)(32),cout=>p(348)(33));
FA_ff_13683:FAff port map(x=>p(326)(33),y=>p(327)(33),Cin=>p(328)(33),clock=>clock,reset=>reset,s=>p(347)(33),cout=>p(348)(34));
FA_ff_13684:FAff port map(x=>p(326)(34),y=>p(327)(34),Cin=>p(328)(34),clock=>clock,reset=>reset,s=>p(347)(34),cout=>p(348)(35));
FA_ff_13685:FAff port map(x=>p(326)(35),y=>p(327)(35),Cin=>p(328)(35),clock=>clock,reset=>reset,s=>p(347)(35),cout=>p(348)(36));
FA_ff_13686:FAff port map(x=>p(326)(36),y=>p(327)(36),Cin=>p(328)(36),clock=>clock,reset=>reset,s=>p(347)(36),cout=>p(348)(37));
FA_ff_13687:FAff port map(x=>p(326)(37),y=>p(327)(37),Cin=>p(328)(37),clock=>clock,reset=>reset,s=>p(347)(37),cout=>p(348)(38));
FA_ff_13688:FAff port map(x=>p(326)(38),y=>p(327)(38),Cin=>p(328)(38),clock=>clock,reset=>reset,s=>p(347)(38),cout=>p(348)(39));
FA_ff_13689:FAff port map(x=>p(326)(39),y=>p(327)(39),Cin=>p(328)(39),clock=>clock,reset=>reset,s=>p(347)(39),cout=>p(348)(40));
FA_ff_13690:FAff port map(x=>p(326)(40),y=>p(327)(40),Cin=>p(328)(40),clock=>clock,reset=>reset,s=>p(347)(40),cout=>p(348)(41));
FA_ff_13691:FAff port map(x=>p(326)(41),y=>p(327)(41),Cin=>p(328)(41),clock=>clock,reset=>reset,s=>p(347)(41),cout=>p(348)(42));
FA_ff_13692:FAff port map(x=>p(326)(42),y=>p(327)(42),Cin=>p(328)(42),clock=>clock,reset=>reset,s=>p(347)(42),cout=>p(348)(43));
FA_ff_13693:FAff port map(x=>p(326)(43),y=>p(327)(43),Cin=>p(328)(43),clock=>clock,reset=>reset,s=>p(347)(43),cout=>p(348)(44));
FA_ff_13694:FAff port map(x=>p(326)(44),y=>p(327)(44),Cin=>p(328)(44),clock=>clock,reset=>reset,s=>p(347)(44),cout=>p(348)(45));
FA_ff_13695:FAff port map(x=>p(326)(45),y=>p(327)(45),Cin=>p(328)(45),clock=>clock,reset=>reset,s=>p(347)(45),cout=>p(348)(46));
FA_ff_13696:FAff port map(x=>p(326)(46),y=>p(327)(46),Cin=>p(328)(46),clock=>clock,reset=>reset,s=>p(347)(46),cout=>p(348)(47));
FA_ff_13697:FAff port map(x=>p(326)(47),y=>p(327)(47),Cin=>p(328)(47),clock=>clock,reset=>reset,s=>p(347)(47),cout=>p(348)(48));
FA_ff_13698:FAff port map(x=>p(326)(48),y=>p(327)(48),Cin=>p(328)(48),clock=>clock,reset=>reset,s=>p(347)(48),cout=>p(348)(49));
FA_ff_13699:FAff port map(x=>p(326)(49),y=>p(327)(49),Cin=>p(328)(49),clock=>clock,reset=>reset,s=>p(347)(49),cout=>p(348)(50));
FA_ff_13700:FAff port map(x=>p(326)(50),y=>p(327)(50),Cin=>p(328)(50),clock=>clock,reset=>reset,s=>p(347)(50),cout=>p(348)(51));
FA_ff_13701:FAff port map(x=>p(326)(51),y=>p(327)(51),Cin=>p(328)(51),clock=>clock,reset=>reset,s=>p(347)(51),cout=>p(348)(52));
FA_ff_13702:FAff port map(x=>p(326)(52),y=>p(327)(52),Cin=>p(328)(52),clock=>clock,reset=>reset,s=>p(347)(52),cout=>p(348)(53));
FA_ff_13703:FAff port map(x=>p(326)(53),y=>p(327)(53),Cin=>p(328)(53),clock=>clock,reset=>reset,s=>p(347)(53),cout=>p(348)(54));
FA_ff_13704:FAff port map(x=>p(326)(54),y=>p(327)(54),Cin=>p(328)(54),clock=>clock,reset=>reset,s=>p(347)(54),cout=>p(348)(55));
FA_ff_13705:FAff port map(x=>p(326)(55),y=>p(327)(55),Cin=>p(328)(55),clock=>clock,reset=>reset,s=>p(347)(55),cout=>p(348)(56));
FA_ff_13706:FAff port map(x=>p(326)(56),y=>p(327)(56),Cin=>p(328)(56),clock=>clock,reset=>reset,s=>p(347)(56),cout=>p(348)(57));
FA_ff_13707:FAff port map(x=>p(326)(57),y=>p(327)(57),Cin=>p(328)(57),clock=>clock,reset=>reset,s=>p(347)(57),cout=>p(348)(58));
FA_ff_13708:FAff port map(x=>p(326)(58),y=>p(327)(58),Cin=>p(328)(58),clock=>clock,reset=>reset,s=>p(347)(58),cout=>p(348)(59));
FA_ff_13709:FAff port map(x=>p(326)(59),y=>p(327)(59),Cin=>p(328)(59),clock=>clock,reset=>reset,s=>p(347)(59),cout=>p(348)(60));
FA_ff_13710:FAff port map(x=>p(326)(60),y=>p(327)(60),Cin=>p(328)(60),clock=>clock,reset=>reset,s=>p(347)(60),cout=>p(348)(61));
FA_ff_13711:FAff port map(x=>p(326)(61),y=>p(327)(61),Cin=>p(328)(61),clock=>clock,reset=>reset,s=>p(347)(61),cout=>p(348)(62));
FA_ff_13712:FAff port map(x=>p(326)(62),y=>p(327)(62),Cin=>p(328)(62),clock=>clock,reset=>reset,s=>p(347)(62),cout=>p(348)(63));
FA_ff_13713:FAff port map(x=>p(326)(63),y=>p(327)(63),Cin=>p(328)(63),clock=>clock,reset=>reset,s=>p(347)(63),cout=>p(348)(64));
FA_ff_13714:FAff port map(x=>p(326)(64),y=>p(327)(64),Cin=>p(328)(64),clock=>clock,reset=>reset,s=>p(347)(64),cout=>p(348)(65));
FA_ff_13715:FAff port map(x=>p(326)(65),y=>p(327)(65),Cin=>p(328)(65),clock=>clock,reset=>reset,s=>p(347)(65),cout=>p(348)(66));
FA_ff_13716:FAff port map(x=>p(326)(66),y=>p(327)(66),Cin=>p(328)(66),clock=>clock,reset=>reset,s=>p(347)(66),cout=>p(348)(67));
FA_ff_13717:FAff port map(x=>p(326)(67),y=>p(327)(67),Cin=>p(328)(67),clock=>clock,reset=>reset,s=>p(347)(67),cout=>p(348)(68));
FA_ff_13718:FAff port map(x=>p(326)(68),y=>p(327)(68),Cin=>p(328)(68),clock=>clock,reset=>reset,s=>p(347)(68),cout=>p(348)(69));
FA_ff_13719:FAff port map(x=>p(326)(69),y=>p(327)(69),Cin=>p(328)(69),clock=>clock,reset=>reset,s=>p(347)(69),cout=>p(348)(70));
FA_ff_13720:FAff port map(x=>p(326)(70),y=>p(327)(70),Cin=>p(328)(70),clock=>clock,reset=>reset,s=>p(347)(70),cout=>p(348)(71));
FA_ff_13721:FAff port map(x=>p(326)(71),y=>p(327)(71),Cin=>p(328)(71),clock=>clock,reset=>reset,s=>p(347)(71),cout=>p(348)(72));
FA_ff_13722:FAff port map(x=>p(326)(72),y=>p(327)(72),Cin=>p(328)(72),clock=>clock,reset=>reset,s=>p(347)(72),cout=>p(348)(73));
FA_ff_13723:FAff port map(x=>p(326)(73),y=>p(327)(73),Cin=>p(328)(73),clock=>clock,reset=>reset,s=>p(347)(73),cout=>p(348)(74));
FA_ff_13724:FAff port map(x=>p(326)(74),y=>p(327)(74),Cin=>p(328)(74),clock=>clock,reset=>reset,s=>p(347)(74),cout=>p(348)(75));
FA_ff_13725:FAff port map(x=>p(326)(75),y=>p(327)(75),Cin=>p(328)(75),clock=>clock,reset=>reset,s=>p(347)(75),cout=>p(348)(76));
FA_ff_13726:FAff port map(x=>p(326)(76),y=>p(327)(76),Cin=>p(328)(76),clock=>clock,reset=>reset,s=>p(347)(76),cout=>p(348)(77));
FA_ff_13727:FAff port map(x=>p(326)(77),y=>p(327)(77),Cin=>p(328)(77),clock=>clock,reset=>reset,s=>p(347)(77),cout=>p(348)(78));
FA_ff_13728:FAff port map(x=>p(326)(78),y=>p(327)(78),Cin=>p(328)(78),clock=>clock,reset=>reset,s=>p(347)(78),cout=>p(348)(79));
FA_ff_13729:FAff port map(x=>p(326)(79),y=>p(327)(79),Cin=>p(328)(79),clock=>clock,reset=>reset,s=>p(347)(79),cout=>p(348)(80));
FA_ff_13730:FAff port map(x=>p(326)(80),y=>p(327)(80),Cin=>p(328)(80),clock=>clock,reset=>reset,s=>p(347)(80),cout=>p(348)(81));
FA_ff_13731:FAff port map(x=>p(326)(81),y=>p(327)(81),Cin=>p(328)(81),clock=>clock,reset=>reset,s=>p(347)(81),cout=>p(348)(82));
FA_ff_13732:FAff port map(x=>p(326)(82),y=>p(327)(82),Cin=>p(328)(82),clock=>clock,reset=>reset,s=>p(347)(82),cout=>p(348)(83));
FA_ff_13733:FAff port map(x=>p(326)(83),y=>p(327)(83),Cin=>p(328)(83),clock=>clock,reset=>reset,s=>p(347)(83),cout=>p(348)(84));
FA_ff_13734:FAff port map(x=>p(326)(84),y=>p(327)(84),Cin=>p(328)(84),clock=>clock,reset=>reset,s=>p(347)(84),cout=>p(348)(85));
FA_ff_13735:FAff port map(x=>p(326)(85),y=>p(327)(85),Cin=>p(328)(85),clock=>clock,reset=>reset,s=>p(347)(85),cout=>p(348)(86));
FA_ff_13736:FAff port map(x=>p(326)(86),y=>p(327)(86),Cin=>p(328)(86),clock=>clock,reset=>reset,s=>p(347)(86),cout=>p(348)(87));
FA_ff_13737:FAff port map(x=>p(326)(87),y=>p(327)(87),Cin=>p(328)(87),clock=>clock,reset=>reset,s=>p(347)(87),cout=>p(348)(88));
FA_ff_13738:FAff port map(x=>p(326)(88),y=>p(327)(88),Cin=>p(328)(88),clock=>clock,reset=>reset,s=>p(347)(88),cout=>p(348)(89));
FA_ff_13739:FAff port map(x=>p(326)(89),y=>p(327)(89),Cin=>p(328)(89),clock=>clock,reset=>reset,s=>p(347)(89),cout=>p(348)(90));
FA_ff_13740:FAff port map(x=>p(326)(90),y=>p(327)(90),Cin=>p(328)(90),clock=>clock,reset=>reset,s=>p(347)(90),cout=>p(348)(91));
FA_ff_13741:FAff port map(x=>p(326)(91),y=>p(327)(91),Cin=>p(328)(91),clock=>clock,reset=>reset,s=>p(347)(91),cout=>p(348)(92));
FA_ff_13742:FAff port map(x=>p(326)(92),y=>p(327)(92),Cin=>p(328)(92),clock=>clock,reset=>reset,s=>p(347)(92),cout=>p(348)(93));
FA_ff_13743:FAff port map(x=>p(326)(93),y=>p(327)(93),Cin=>p(328)(93),clock=>clock,reset=>reset,s=>p(347)(93),cout=>p(348)(94));
FA_ff_13744:FAff port map(x=>p(326)(94),y=>p(327)(94),Cin=>p(328)(94),clock=>clock,reset=>reset,s=>p(347)(94),cout=>p(348)(95));
FA_ff_13745:FAff port map(x=>p(326)(95),y=>p(327)(95),Cin=>p(328)(95),clock=>clock,reset=>reset,s=>p(347)(95),cout=>p(348)(96));
FA_ff_13746:FAff port map(x=>p(326)(96),y=>p(327)(96),Cin=>p(328)(96),clock=>clock,reset=>reset,s=>p(347)(96),cout=>p(348)(97));
FA_ff_13747:FAff port map(x=>p(326)(97),y=>p(327)(97),Cin=>p(328)(97),clock=>clock,reset=>reset,s=>p(347)(97),cout=>p(348)(98));
FA_ff_13748:FAff port map(x=>p(326)(98),y=>p(327)(98),Cin=>p(328)(98),clock=>clock,reset=>reset,s=>p(347)(98),cout=>p(348)(99));
FA_ff_13749:FAff port map(x=>p(326)(99),y=>p(327)(99),Cin=>p(328)(99),clock=>clock,reset=>reset,s=>p(347)(99),cout=>p(348)(100));
FA_ff_13750:FAff port map(x=>p(326)(100),y=>p(327)(100),Cin=>p(328)(100),clock=>clock,reset=>reset,s=>p(347)(100),cout=>p(348)(101));
FA_ff_13751:FAff port map(x=>p(326)(101),y=>p(327)(101),Cin=>p(328)(101),clock=>clock,reset=>reset,s=>p(347)(101),cout=>p(348)(102));
FA_ff_13752:FAff port map(x=>p(326)(102),y=>p(327)(102),Cin=>p(328)(102),clock=>clock,reset=>reset,s=>p(347)(102),cout=>p(348)(103));
FA_ff_13753:FAff port map(x=>p(326)(103),y=>p(327)(103),Cin=>p(328)(103),clock=>clock,reset=>reset,s=>p(347)(103),cout=>p(348)(104));
FA_ff_13754:FAff port map(x=>p(326)(104),y=>p(327)(104),Cin=>p(328)(104),clock=>clock,reset=>reset,s=>p(347)(104),cout=>p(348)(105));
FA_ff_13755:FAff port map(x=>p(326)(105),y=>p(327)(105),Cin=>p(328)(105),clock=>clock,reset=>reset,s=>p(347)(105),cout=>p(348)(106));
FA_ff_13756:FAff port map(x=>p(326)(106),y=>p(327)(106),Cin=>p(328)(106),clock=>clock,reset=>reset,s=>p(347)(106),cout=>p(348)(107));
FA_ff_13757:FAff port map(x=>p(326)(107),y=>p(327)(107),Cin=>p(328)(107),clock=>clock,reset=>reset,s=>p(347)(107),cout=>p(348)(108));
FA_ff_13758:FAff port map(x=>p(326)(108),y=>p(327)(108),Cin=>p(328)(108),clock=>clock,reset=>reset,s=>p(347)(108),cout=>p(348)(109));
FA_ff_13759:FAff port map(x=>p(326)(109),y=>p(327)(109),Cin=>p(328)(109),clock=>clock,reset=>reset,s=>p(347)(109),cout=>p(348)(110));
FA_ff_13760:FAff port map(x=>p(326)(110),y=>p(327)(110),Cin=>p(328)(110),clock=>clock,reset=>reset,s=>p(347)(110),cout=>p(348)(111));
FA_ff_13761:FAff port map(x=>p(326)(111),y=>p(327)(111),Cin=>p(328)(111),clock=>clock,reset=>reset,s=>p(347)(111),cout=>p(348)(112));
FA_ff_13762:FAff port map(x=>p(326)(112),y=>p(327)(112),Cin=>p(328)(112),clock=>clock,reset=>reset,s=>p(347)(112),cout=>p(348)(113));
FA_ff_13763:FAff port map(x=>p(326)(113),y=>p(327)(113),Cin=>p(328)(113),clock=>clock,reset=>reset,s=>p(347)(113),cout=>p(348)(114));
FA_ff_13764:FAff port map(x=>p(326)(114),y=>p(327)(114),Cin=>p(328)(114),clock=>clock,reset=>reset,s=>p(347)(114),cout=>p(348)(115));
FA_ff_13765:FAff port map(x=>p(326)(115),y=>p(327)(115),Cin=>p(328)(115),clock=>clock,reset=>reset,s=>p(347)(115),cout=>p(348)(116));
FA_ff_13766:FAff port map(x=>p(326)(116),y=>p(327)(116),Cin=>p(328)(116),clock=>clock,reset=>reset,s=>p(347)(116),cout=>p(348)(117));
FA_ff_13767:FAff port map(x=>p(326)(117),y=>p(327)(117),Cin=>p(328)(117),clock=>clock,reset=>reset,s=>p(347)(117),cout=>p(348)(118));
FA_ff_13768:FAff port map(x=>p(326)(118),y=>p(327)(118),Cin=>p(328)(118),clock=>clock,reset=>reset,s=>p(347)(118),cout=>p(348)(119));
FA_ff_13769:FAff port map(x=>p(326)(119),y=>p(327)(119),Cin=>p(328)(119),clock=>clock,reset=>reset,s=>p(347)(119),cout=>p(348)(120));
FA_ff_13770:FAff port map(x=>p(326)(120),y=>p(327)(120),Cin=>p(328)(120),clock=>clock,reset=>reset,s=>p(347)(120),cout=>p(348)(121));
FA_ff_13771:FAff port map(x=>p(326)(121),y=>p(327)(121),Cin=>p(328)(121),clock=>clock,reset=>reset,s=>p(347)(121),cout=>p(348)(122));
FA_ff_13772:FAff port map(x=>p(326)(122),y=>p(327)(122),Cin=>p(328)(122),clock=>clock,reset=>reset,s=>p(347)(122),cout=>p(348)(123));
FA_ff_13773:FAff port map(x=>p(326)(123),y=>p(327)(123),Cin=>p(328)(123),clock=>clock,reset=>reset,s=>p(347)(123),cout=>p(348)(124));
FA_ff_13774:FAff port map(x=>p(326)(124),y=>p(327)(124),Cin=>p(328)(124),clock=>clock,reset=>reset,s=>p(347)(124),cout=>p(348)(125));
FA_ff_13775:FAff port map(x=>p(326)(125),y=>p(327)(125),Cin=>p(328)(125),clock=>clock,reset=>reset,s=>p(347)(125),cout=>p(348)(126));
FA_ff_13776:FAff port map(x=>p(326)(126),y=>p(327)(126),Cin=>p(328)(126),clock=>clock,reset=>reset,s=>p(347)(126),cout=>p(348)(127));
FA_ff_13777:FAff port map(x=>p(326)(127),y=>p(327)(127),Cin=>p(328)(127),clock=>clock,reset=>reset,s=>p(347)(127),cout=>p(348)(128));
FA_ff_13778:FAff port map(x=>p(326)(128),y=>p(327)(128),Cin=>p(328)(128),clock=>clock,reset=>reset,s=>p(347)(128),cout=>p(348)(129));
FA_ff_13779:FAff port map(x=>p(326)(129),y=>p(327)(129),Cin=>p(328)(129),clock=>clock,reset=>reset,s=>p(347)(129),cout=>p(348)(130));
HA_ff_85:HAff port map(x=>p(326)(130),y=>p(328)(130),clock=>clock,reset=>reset,s=>p(347)(130),c=>p(348)(131));
HA_ff_86:HAff port map(x=>p(329)(0),y=>p(331)(0),clock=>clock,reset=>reset,s=>p(349)(0),c=>p(350)(1));
HA_ff_87:HAff port map(x=>p(329)(1),y=>p(331)(1),clock=>clock,reset=>reset,s=>p(349)(1),c=>p(350)(2));
FA_ff_13780:FAff port map(x=>p(329)(2),y=>p(330)(2),Cin=>p(331)(2),clock=>clock,reset=>reset,s=>p(349)(2),cout=>p(350)(3));
FA_ff_13781:FAff port map(x=>p(329)(3),y=>p(330)(3),Cin=>p(331)(3),clock=>clock,reset=>reset,s=>p(349)(3),cout=>p(350)(4));
FA_ff_13782:FAff port map(x=>p(329)(4),y=>p(330)(4),Cin=>p(331)(4),clock=>clock,reset=>reset,s=>p(349)(4),cout=>p(350)(5));
FA_ff_13783:FAff port map(x=>p(329)(5),y=>p(330)(5),Cin=>p(331)(5),clock=>clock,reset=>reset,s=>p(349)(5),cout=>p(350)(6));
FA_ff_13784:FAff port map(x=>p(329)(6),y=>p(330)(6),Cin=>p(331)(6),clock=>clock,reset=>reset,s=>p(349)(6),cout=>p(350)(7));
FA_ff_13785:FAff port map(x=>p(329)(7),y=>p(330)(7),Cin=>p(331)(7),clock=>clock,reset=>reset,s=>p(349)(7),cout=>p(350)(8));
FA_ff_13786:FAff port map(x=>p(329)(8),y=>p(330)(8),Cin=>p(331)(8),clock=>clock,reset=>reset,s=>p(349)(8),cout=>p(350)(9));
FA_ff_13787:FAff port map(x=>p(329)(9),y=>p(330)(9),Cin=>p(331)(9),clock=>clock,reset=>reset,s=>p(349)(9),cout=>p(350)(10));
FA_ff_13788:FAff port map(x=>p(329)(10),y=>p(330)(10),Cin=>p(331)(10),clock=>clock,reset=>reset,s=>p(349)(10),cout=>p(350)(11));
FA_ff_13789:FAff port map(x=>p(329)(11),y=>p(330)(11),Cin=>p(331)(11),clock=>clock,reset=>reset,s=>p(349)(11),cout=>p(350)(12));
FA_ff_13790:FAff port map(x=>p(329)(12),y=>p(330)(12),Cin=>p(331)(12),clock=>clock,reset=>reset,s=>p(349)(12),cout=>p(350)(13));
FA_ff_13791:FAff port map(x=>p(329)(13),y=>p(330)(13),Cin=>p(331)(13),clock=>clock,reset=>reset,s=>p(349)(13),cout=>p(350)(14));
FA_ff_13792:FAff port map(x=>p(329)(14),y=>p(330)(14),Cin=>p(331)(14),clock=>clock,reset=>reset,s=>p(349)(14),cout=>p(350)(15));
FA_ff_13793:FAff port map(x=>p(329)(15),y=>p(330)(15),Cin=>p(331)(15),clock=>clock,reset=>reset,s=>p(349)(15),cout=>p(350)(16));
FA_ff_13794:FAff port map(x=>p(329)(16),y=>p(330)(16),Cin=>p(331)(16),clock=>clock,reset=>reset,s=>p(349)(16),cout=>p(350)(17));
FA_ff_13795:FAff port map(x=>p(329)(17),y=>p(330)(17),Cin=>p(331)(17),clock=>clock,reset=>reset,s=>p(349)(17),cout=>p(350)(18));
FA_ff_13796:FAff port map(x=>p(329)(18),y=>p(330)(18),Cin=>p(331)(18),clock=>clock,reset=>reset,s=>p(349)(18),cout=>p(350)(19));
FA_ff_13797:FAff port map(x=>p(329)(19),y=>p(330)(19),Cin=>p(331)(19),clock=>clock,reset=>reset,s=>p(349)(19),cout=>p(350)(20));
FA_ff_13798:FAff port map(x=>p(329)(20),y=>p(330)(20),Cin=>p(331)(20),clock=>clock,reset=>reset,s=>p(349)(20),cout=>p(350)(21));
FA_ff_13799:FAff port map(x=>p(329)(21),y=>p(330)(21),Cin=>p(331)(21),clock=>clock,reset=>reset,s=>p(349)(21),cout=>p(350)(22));
FA_ff_13800:FAff port map(x=>p(329)(22),y=>p(330)(22),Cin=>p(331)(22),clock=>clock,reset=>reset,s=>p(349)(22),cout=>p(350)(23));
FA_ff_13801:FAff port map(x=>p(329)(23),y=>p(330)(23),Cin=>p(331)(23),clock=>clock,reset=>reset,s=>p(349)(23),cout=>p(350)(24));
FA_ff_13802:FAff port map(x=>p(329)(24),y=>p(330)(24),Cin=>p(331)(24),clock=>clock,reset=>reset,s=>p(349)(24),cout=>p(350)(25));
FA_ff_13803:FAff port map(x=>p(329)(25),y=>p(330)(25),Cin=>p(331)(25),clock=>clock,reset=>reset,s=>p(349)(25),cout=>p(350)(26));
FA_ff_13804:FAff port map(x=>p(329)(26),y=>p(330)(26),Cin=>p(331)(26),clock=>clock,reset=>reset,s=>p(349)(26),cout=>p(350)(27));
FA_ff_13805:FAff port map(x=>p(329)(27),y=>p(330)(27),Cin=>p(331)(27),clock=>clock,reset=>reset,s=>p(349)(27),cout=>p(350)(28));
FA_ff_13806:FAff port map(x=>p(329)(28),y=>p(330)(28),Cin=>p(331)(28),clock=>clock,reset=>reset,s=>p(349)(28),cout=>p(350)(29));
FA_ff_13807:FAff port map(x=>p(329)(29),y=>p(330)(29),Cin=>p(331)(29),clock=>clock,reset=>reset,s=>p(349)(29),cout=>p(350)(30));
FA_ff_13808:FAff port map(x=>p(329)(30),y=>p(330)(30),Cin=>p(331)(30),clock=>clock,reset=>reset,s=>p(349)(30),cout=>p(350)(31));
FA_ff_13809:FAff port map(x=>p(329)(31),y=>p(330)(31),Cin=>p(331)(31),clock=>clock,reset=>reset,s=>p(349)(31),cout=>p(350)(32));
FA_ff_13810:FAff port map(x=>p(329)(32),y=>p(330)(32),Cin=>p(331)(32),clock=>clock,reset=>reset,s=>p(349)(32),cout=>p(350)(33));
FA_ff_13811:FAff port map(x=>p(329)(33),y=>p(330)(33),Cin=>p(331)(33),clock=>clock,reset=>reset,s=>p(349)(33),cout=>p(350)(34));
FA_ff_13812:FAff port map(x=>p(329)(34),y=>p(330)(34),Cin=>p(331)(34),clock=>clock,reset=>reset,s=>p(349)(34),cout=>p(350)(35));
FA_ff_13813:FAff port map(x=>p(329)(35),y=>p(330)(35),Cin=>p(331)(35),clock=>clock,reset=>reset,s=>p(349)(35),cout=>p(350)(36));
FA_ff_13814:FAff port map(x=>p(329)(36),y=>p(330)(36),Cin=>p(331)(36),clock=>clock,reset=>reset,s=>p(349)(36),cout=>p(350)(37));
FA_ff_13815:FAff port map(x=>p(329)(37),y=>p(330)(37),Cin=>p(331)(37),clock=>clock,reset=>reset,s=>p(349)(37),cout=>p(350)(38));
FA_ff_13816:FAff port map(x=>p(329)(38),y=>p(330)(38),Cin=>p(331)(38),clock=>clock,reset=>reset,s=>p(349)(38),cout=>p(350)(39));
FA_ff_13817:FAff port map(x=>p(329)(39),y=>p(330)(39),Cin=>p(331)(39),clock=>clock,reset=>reset,s=>p(349)(39),cout=>p(350)(40));
FA_ff_13818:FAff port map(x=>p(329)(40),y=>p(330)(40),Cin=>p(331)(40),clock=>clock,reset=>reset,s=>p(349)(40),cout=>p(350)(41));
FA_ff_13819:FAff port map(x=>p(329)(41),y=>p(330)(41),Cin=>p(331)(41),clock=>clock,reset=>reset,s=>p(349)(41),cout=>p(350)(42));
FA_ff_13820:FAff port map(x=>p(329)(42),y=>p(330)(42),Cin=>p(331)(42),clock=>clock,reset=>reset,s=>p(349)(42),cout=>p(350)(43));
FA_ff_13821:FAff port map(x=>p(329)(43),y=>p(330)(43),Cin=>p(331)(43),clock=>clock,reset=>reset,s=>p(349)(43),cout=>p(350)(44));
FA_ff_13822:FAff port map(x=>p(329)(44),y=>p(330)(44),Cin=>p(331)(44),clock=>clock,reset=>reset,s=>p(349)(44),cout=>p(350)(45));
FA_ff_13823:FAff port map(x=>p(329)(45),y=>p(330)(45),Cin=>p(331)(45),clock=>clock,reset=>reset,s=>p(349)(45),cout=>p(350)(46));
FA_ff_13824:FAff port map(x=>p(329)(46),y=>p(330)(46),Cin=>p(331)(46),clock=>clock,reset=>reset,s=>p(349)(46),cout=>p(350)(47));
FA_ff_13825:FAff port map(x=>p(329)(47),y=>p(330)(47),Cin=>p(331)(47),clock=>clock,reset=>reset,s=>p(349)(47),cout=>p(350)(48));
FA_ff_13826:FAff port map(x=>p(329)(48),y=>p(330)(48),Cin=>p(331)(48),clock=>clock,reset=>reset,s=>p(349)(48),cout=>p(350)(49));
FA_ff_13827:FAff port map(x=>p(329)(49),y=>p(330)(49),Cin=>p(331)(49),clock=>clock,reset=>reset,s=>p(349)(49),cout=>p(350)(50));
FA_ff_13828:FAff port map(x=>p(329)(50),y=>p(330)(50),Cin=>p(331)(50),clock=>clock,reset=>reset,s=>p(349)(50),cout=>p(350)(51));
FA_ff_13829:FAff port map(x=>p(329)(51),y=>p(330)(51),Cin=>p(331)(51),clock=>clock,reset=>reset,s=>p(349)(51),cout=>p(350)(52));
FA_ff_13830:FAff port map(x=>p(329)(52),y=>p(330)(52),Cin=>p(331)(52),clock=>clock,reset=>reset,s=>p(349)(52),cout=>p(350)(53));
FA_ff_13831:FAff port map(x=>p(329)(53),y=>p(330)(53),Cin=>p(331)(53),clock=>clock,reset=>reset,s=>p(349)(53),cout=>p(350)(54));
FA_ff_13832:FAff port map(x=>p(329)(54),y=>p(330)(54),Cin=>p(331)(54),clock=>clock,reset=>reset,s=>p(349)(54),cout=>p(350)(55));
FA_ff_13833:FAff port map(x=>p(329)(55),y=>p(330)(55),Cin=>p(331)(55),clock=>clock,reset=>reset,s=>p(349)(55),cout=>p(350)(56));
FA_ff_13834:FAff port map(x=>p(329)(56),y=>p(330)(56),Cin=>p(331)(56),clock=>clock,reset=>reset,s=>p(349)(56),cout=>p(350)(57));
FA_ff_13835:FAff port map(x=>p(329)(57),y=>p(330)(57),Cin=>p(331)(57),clock=>clock,reset=>reset,s=>p(349)(57),cout=>p(350)(58));
FA_ff_13836:FAff port map(x=>p(329)(58),y=>p(330)(58),Cin=>p(331)(58),clock=>clock,reset=>reset,s=>p(349)(58),cout=>p(350)(59));
FA_ff_13837:FAff port map(x=>p(329)(59),y=>p(330)(59),Cin=>p(331)(59),clock=>clock,reset=>reset,s=>p(349)(59),cout=>p(350)(60));
FA_ff_13838:FAff port map(x=>p(329)(60),y=>p(330)(60),Cin=>p(331)(60),clock=>clock,reset=>reset,s=>p(349)(60),cout=>p(350)(61));
FA_ff_13839:FAff port map(x=>p(329)(61),y=>p(330)(61),Cin=>p(331)(61),clock=>clock,reset=>reset,s=>p(349)(61),cout=>p(350)(62));
FA_ff_13840:FAff port map(x=>p(329)(62),y=>p(330)(62),Cin=>p(331)(62),clock=>clock,reset=>reset,s=>p(349)(62),cout=>p(350)(63));
FA_ff_13841:FAff port map(x=>p(329)(63),y=>p(330)(63),Cin=>p(331)(63),clock=>clock,reset=>reset,s=>p(349)(63),cout=>p(350)(64));
FA_ff_13842:FAff port map(x=>p(329)(64),y=>p(330)(64),Cin=>p(331)(64),clock=>clock,reset=>reset,s=>p(349)(64),cout=>p(350)(65));
FA_ff_13843:FAff port map(x=>p(329)(65),y=>p(330)(65),Cin=>p(331)(65),clock=>clock,reset=>reset,s=>p(349)(65),cout=>p(350)(66));
FA_ff_13844:FAff port map(x=>p(329)(66),y=>p(330)(66),Cin=>p(331)(66),clock=>clock,reset=>reset,s=>p(349)(66),cout=>p(350)(67));
FA_ff_13845:FAff port map(x=>p(329)(67),y=>p(330)(67),Cin=>p(331)(67),clock=>clock,reset=>reset,s=>p(349)(67),cout=>p(350)(68));
FA_ff_13846:FAff port map(x=>p(329)(68),y=>p(330)(68),Cin=>p(331)(68),clock=>clock,reset=>reset,s=>p(349)(68),cout=>p(350)(69));
FA_ff_13847:FAff port map(x=>p(329)(69),y=>p(330)(69),Cin=>p(331)(69),clock=>clock,reset=>reset,s=>p(349)(69),cout=>p(350)(70));
FA_ff_13848:FAff port map(x=>p(329)(70),y=>p(330)(70),Cin=>p(331)(70),clock=>clock,reset=>reset,s=>p(349)(70),cout=>p(350)(71));
FA_ff_13849:FAff port map(x=>p(329)(71),y=>p(330)(71),Cin=>p(331)(71),clock=>clock,reset=>reset,s=>p(349)(71),cout=>p(350)(72));
FA_ff_13850:FAff port map(x=>p(329)(72),y=>p(330)(72),Cin=>p(331)(72),clock=>clock,reset=>reset,s=>p(349)(72),cout=>p(350)(73));
FA_ff_13851:FAff port map(x=>p(329)(73),y=>p(330)(73),Cin=>p(331)(73),clock=>clock,reset=>reset,s=>p(349)(73),cout=>p(350)(74));
FA_ff_13852:FAff port map(x=>p(329)(74),y=>p(330)(74),Cin=>p(331)(74),clock=>clock,reset=>reset,s=>p(349)(74),cout=>p(350)(75));
FA_ff_13853:FAff port map(x=>p(329)(75),y=>p(330)(75),Cin=>p(331)(75),clock=>clock,reset=>reset,s=>p(349)(75),cout=>p(350)(76));
FA_ff_13854:FAff port map(x=>p(329)(76),y=>p(330)(76),Cin=>p(331)(76),clock=>clock,reset=>reset,s=>p(349)(76),cout=>p(350)(77));
FA_ff_13855:FAff port map(x=>p(329)(77),y=>p(330)(77),Cin=>p(331)(77),clock=>clock,reset=>reset,s=>p(349)(77),cout=>p(350)(78));
FA_ff_13856:FAff port map(x=>p(329)(78),y=>p(330)(78),Cin=>p(331)(78),clock=>clock,reset=>reset,s=>p(349)(78),cout=>p(350)(79));
FA_ff_13857:FAff port map(x=>p(329)(79),y=>p(330)(79),Cin=>p(331)(79),clock=>clock,reset=>reset,s=>p(349)(79),cout=>p(350)(80));
FA_ff_13858:FAff port map(x=>p(329)(80),y=>p(330)(80),Cin=>p(331)(80),clock=>clock,reset=>reset,s=>p(349)(80),cout=>p(350)(81));
FA_ff_13859:FAff port map(x=>p(329)(81),y=>p(330)(81),Cin=>p(331)(81),clock=>clock,reset=>reset,s=>p(349)(81),cout=>p(350)(82));
FA_ff_13860:FAff port map(x=>p(329)(82),y=>p(330)(82),Cin=>p(331)(82),clock=>clock,reset=>reset,s=>p(349)(82),cout=>p(350)(83));
FA_ff_13861:FAff port map(x=>p(329)(83),y=>p(330)(83),Cin=>p(331)(83),clock=>clock,reset=>reset,s=>p(349)(83),cout=>p(350)(84));
FA_ff_13862:FAff port map(x=>p(329)(84),y=>p(330)(84),Cin=>p(331)(84),clock=>clock,reset=>reset,s=>p(349)(84),cout=>p(350)(85));
FA_ff_13863:FAff port map(x=>p(329)(85),y=>p(330)(85),Cin=>p(331)(85),clock=>clock,reset=>reset,s=>p(349)(85),cout=>p(350)(86));
FA_ff_13864:FAff port map(x=>p(329)(86),y=>p(330)(86),Cin=>p(331)(86),clock=>clock,reset=>reset,s=>p(349)(86),cout=>p(350)(87));
FA_ff_13865:FAff port map(x=>p(329)(87),y=>p(330)(87),Cin=>p(331)(87),clock=>clock,reset=>reset,s=>p(349)(87),cout=>p(350)(88));
FA_ff_13866:FAff port map(x=>p(329)(88),y=>p(330)(88),Cin=>p(331)(88),clock=>clock,reset=>reset,s=>p(349)(88),cout=>p(350)(89));
FA_ff_13867:FAff port map(x=>p(329)(89),y=>p(330)(89),Cin=>p(331)(89),clock=>clock,reset=>reset,s=>p(349)(89),cout=>p(350)(90));
FA_ff_13868:FAff port map(x=>p(329)(90),y=>p(330)(90),Cin=>p(331)(90),clock=>clock,reset=>reset,s=>p(349)(90),cout=>p(350)(91));
FA_ff_13869:FAff port map(x=>p(329)(91),y=>p(330)(91),Cin=>p(331)(91),clock=>clock,reset=>reset,s=>p(349)(91),cout=>p(350)(92));
FA_ff_13870:FAff port map(x=>p(329)(92),y=>p(330)(92),Cin=>p(331)(92),clock=>clock,reset=>reset,s=>p(349)(92),cout=>p(350)(93));
FA_ff_13871:FAff port map(x=>p(329)(93),y=>p(330)(93),Cin=>p(331)(93),clock=>clock,reset=>reset,s=>p(349)(93),cout=>p(350)(94));
FA_ff_13872:FAff port map(x=>p(329)(94),y=>p(330)(94),Cin=>p(331)(94),clock=>clock,reset=>reset,s=>p(349)(94),cout=>p(350)(95));
FA_ff_13873:FAff port map(x=>p(329)(95),y=>p(330)(95),Cin=>p(331)(95),clock=>clock,reset=>reset,s=>p(349)(95),cout=>p(350)(96));
FA_ff_13874:FAff port map(x=>p(329)(96),y=>p(330)(96),Cin=>p(331)(96),clock=>clock,reset=>reset,s=>p(349)(96),cout=>p(350)(97));
FA_ff_13875:FAff port map(x=>p(329)(97),y=>p(330)(97),Cin=>p(331)(97),clock=>clock,reset=>reset,s=>p(349)(97),cout=>p(350)(98));
FA_ff_13876:FAff port map(x=>p(329)(98),y=>p(330)(98),Cin=>p(331)(98),clock=>clock,reset=>reset,s=>p(349)(98),cout=>p(350)(99));
FA_ff_13877:FAff port map(x=>p(329)(99),y=>p(330)(99),Cin=>p(331)(99),clock=>clock,reset=>reset,s=>p(349)(99),cout=>p(350)(100));
FA_ff_13878:FAff port map(x=>p(329)(100),y=>p(330)(100),Cin=>p(331)(100),clock=>clock,reset=>reset,s=>p(349)(100),cout=>p(350)(101));
FA_ff_13879:FAff port map(x=>p(329)(101),y=>p(330)(101),Cin=>p(331)(101),clock=>clock,reset=>reset,s=>p(349)(101),cout=>p(350)(102));
FA_ff_13880:FAff port map(x=>p(329)(102),y=>p(330)(102),Cin=>p(331)(102),clock=>clock,reset=>reset,s=>p(349)(102),cout=>p(350)(103));
FA_ff_13881:FAff port map(x=>p(329)(103),y=>p(330)(103),Cin=>p(331)(103),clock=>clock,reset=>reset,s=>p(349)(103),cout=>p(350)(104));
FA_ff_13882:FAff port map(x=>p(329)(104),y=>p(330)(104),Cin=>p(331)(104),clock=>clock,reset=>reset,s=>p(349)(104),cout=>p(350)(105));
FA_ff_13883:FAff port map(x=>p(329)(105),y=>p(330)(105),Cin=>p(331)(105),clock=>clock,reset=>reset,s=>p(349)(105),cout=>p(350)(106));
FA_ff_13884:FAff port map(x=>p(329)(106),y=>p(330)(106),Cin=>p(331)(106),clock=>clock,reset=>reset,s=>p(349)(106),cout=>p(350)(107));
FA_ff_13885:FAff port map(x=>p(329)(107),y=>p(330)(107),Cin=>p(331)(107),clock=>clock,reset=>reset,s=>p(349)(107),cout=>p(350)(108));
FA_ff_13886:FAff port map(x=>p(329)(108),y=>p(330)(108),Cin=>p(331)(108),clock=>clock,reset=>reset,s=>p(349)(108),cout=>p(350)(109));
FA_ff_13887:FAff port map(x=>p(329)(109),y=>p(330)(109),Cin=>p(331)(109),clock=>clock,reset=>reset,s=>p(349)(109),cout=>p(350)(110));
FA_ff_13888:FAff port map(x=>p(329)(110),y=>p(330)(110),Cin=>p(331)(110),clock=>clock,reset=>reset,s=>p(349)(110),cout=>p(350)(111));
FA_ff_13889:FAff port map(x=>p(329)(111),y=>p(330)(111),Cin=>p(331)(111),clock=>clock,reset=>reset,s=>p(349)(111),cout=>p(350)(112));
FA_ff_13890:FAff port map(x=>p(329)(112),y=>p(330)(112),Cin=>p(331)(112),clock=>clock,reset=>reset,s=>p(349)(112),cout=>p(350)(113));
FA_ff_13891:FAff port map(x=>p(329)(113),y=>p(330)(113),Cin=>p(331)(113),clock=>clock,reset=>reset,s=>p(349)(113),cout=>p(350)(114));
FA_ff_13892:FAff port map(x=>p(329)(114),y=>p(330)(114),Cin=>p(331)(114),clock=>clock,reset=>reset,s=>p(349)(114),cout=>p(350)(115));
FA_ff_13893:FAff port map(x=>p(329)(115),y=>p(330)(115),Cin=>p(331)(115),clock=>clock,reset=>reset,s=>p(349)(115),cout=>p(350)(116));
FA_ff_13894:FAff port map(x=>p(329)(116),y=>p(330)(116),Cin=>p(331)(116),clock=>clock,reset=>reset,s=>p(349)(116),cout=>p(350)(117));
FA_ff_13895:FAff port map(x=>p(329)(117),y=>p(330)(117),Cin=>p(331)(117),clock=>clock,reset=>reset,s=>p(349)(117),cout=>p(350)(118));
FA_ff_13896:FAff port map(x=>p(329)(118),y=>p(330)(118),Cin=>p(331)(118),clock=>clock,reset=>reset,s=>p(349)(118),cout=>p(350)(119));
FA_ff_13897:FAff port map(x=>p(329)(119),y=>p(330)(119),Cin=>p(331)(119),clock=>clock,reset=>reset,s=>p(349)(119),cout=>p(350)(120));
FA_ff_13898:FAff port map(x=>p(329)(120),y=>p(330)(120),Cin=>p(331)(120),clock=>clock,reset=>reset,s=>p(349)(120),cout=>p(350)(121));
FA_ff_13899:FAff port map(x=>p(329)(121),y=>p(330)(121),Cin=>p(331)(121),clock=>clock,reset=>reset,s=>p(349)(121),cout=>p(350)(122));
FA_ff_13900:FAff port map(x=>p(329)(122),y=>p(330)(122),Cin=>p(331)(122),clock=>clock,reset=>reset,s=>p(349)(122),cout=>p(350)(123));
FA_ff_13901:FAff port map(x=>p(329)(123),y=>p(330)(123),Cin=>p(331)(123),clock=>clock,reset=>reset,s=>p(349)(123),cout=>p(350)(124));
FA_ff_13902:FAff port map(x=>p(329)(124),y=>p(330)(124),Cin=>p(331)(124),clock=>clock,reset=>reset,s=>p(349)(124),cout=>p(350)(125));
FA_ff_13903:FAff port map(x=>p(329)(125),y=>p(330)(125),Cin=>p(331)(125),clock=>clock,reset=>reset,s=>p(349)(125),cout=>p(350)(126));
FA_ff_13904:FAff port map(x=>p(329)(126),y=>p(330)(126),Cin=>p(331)(126),clock=>clock,reset=>reset,s=>p(349)(126),cout=>p(350)(127));
FA_ff_13905:FAff port map(x=>p(329)(127),y=>p(330)(127),Cin=>p(331)(127),clock=>clock,reset=>reset,s=>p(349)(127),cout=>p(350)(128));
FA_ff_13906:FAff port map(x=>p(329)(128),y=>p(330)(128),Cin=>p(331)(128),clock=>clock,reset=>reset,s=>p(349)(128),cout=>p(350)(129));
FA_ff_13907:FAff port map(x=>p(329)(129),y=>p(330)(129),Cin=>p(331)(129),clock=>clock,reset=>reset,s=>p(349)(129),cout=>p(350)(130));
p(349)(130)<=p(330)(130);
p(351)(0)<=p(333)(0);
HA_ff_88:HAff port map(x=>p(332)(1),y=>p(333)(1),clock=>clock,reset=>reset,s=>p(351)(1),c=>p(352)(2));
FA_ff_13908:FAff port map(x=>p(332)(2),y=>p(333)(2),Cin=>p(334)(2),clock=>clock,reset=>reset,s=>p(351)(2),cout=>p(352)(3));
FA_ff_13909:FAff port map(x=>p(332)(3),y=>p(333)(3),Cin=>p(334)(3),clock=>clock,reset=>reset,s=>p(351)(3),cout=>p(352)(4));
FA_ff_13910:FAff port map(x=>p(332)(4),y=>p(333)(4),Cin=>p(334)(4),clock=>clock,reset=>reset,s=>p(351)(4),cout=>p(352)(5));
FA_ff_13911:FAff port map(x=>p(332)(5),y=>p(333)(5),Cin=>p(334)(5),clock=>clock,reset=>reset,s=>p(351)(5),cout=>p(352)(6));
FA_ff_13912:FAff port map(x=>p(332)(6),y=>p(333)(6),Cin=>p(334)(6),clock=>clock,reset=>reset,s=>p(351)(6),cout=>p(352)(7));
FA_ff_13913:FAff port map(x=>p(332)(7),y=>p(333)(7),Cin=>p(334)(7),clock=>clock,reset=>reset,s=>p(351)(7),cout=>p(352)(8));
FA_ff_13914:FAff port map(x=>p(332)(8),y=>p(333)(8),Cin=>p(334)(8),clock=>clock,reset=>reset,s=>p(351)(8),cout=>p(352)(9));
FA_ff_13915:FAff port map(x=>p(332)(9),y=>p(333)(9),Cin=>p(334)(9),clock=>clock,reset=>reset,s=>p(351)(9),cout=>p(352)(10));
FA_ff_13916:FAff port map(x=>p(332)(10),y=>p(333)(10),Cin=>p(334)(10),clock=>clock,reset=>reset,s=>p(351)(10),cout=>p(352)(11));
FA_ff_13917:FAff port map(x=>p(332)(11),y=>p(333)(11),Cin=>p(334)(11),clock=>clock,reset=>reset,s=>p(351)(11),cout=>p(352)(12));
FA_ff_13918:FAff port map(x=>p(332)(12),y=>p(333)(12),Cin=>p(334)(12),clock=>clock,reset=>reset,s=>p(351)(12),cout=>p(352)(13));
FA_ff_13919:FAff port map(x=>p(332)(13),y=>p(333)(13),Cin=>p(334)(13),clock=>clock,reset=>reset,s=>p(351)(13),cout=>p(352)(14));
FA_ff_13920:FAff port map(x=>p(332)(14),y=>p(333)(14),Cin=>p(334)(14),clock=>clock,reset=>reset,s=>p(351)(14),cout=>p(352)(15));
FA_ff_13921:FAff port map(x=>p(332)(15),y=>p(333)(15),Cin=>p(334)(15),clock=>clock,reset=>reset,s=>p(351)(15),cout=>p(352)(16));
FA_ff_13922:FAff port map(x=>p(332)(16),y=>p(333)(16),Cin=>p(334)(16),clock=>clock,reset=>reset,s=>p(351)(16),cout=>p(352)(17));
FA_ff_13923:FAff port map(x=>p(332)(17),y=>p(333)(17),Cin=>p(334)(17),clock=>clock,reset=>reset,s=>p(351)(17),cout=>p(352)(18));
FA_ff_13924:FAff port map(x=>p(332)(18),y=>p(333)(18),Cin=>p(334)(18),clock=>clock,reset=>reset,s=>p(351)(18),cout=>p(352)(19));
FA_ff_13925:FAff port map(x=>p(332)(19),y=>p(333)(19),Cin=>p(334)(19),clock=>clock,reset=>reset,s=>p(351)(19),cout=>p(352)(20));
FA_ff_13926:FAff port map(x=>p(332)(20),y=>p(333)(20),Cin=>p(334)(20),clock=>clock,reset=>reset,s=>p(351)(20),cout=>p(352)(21));
FA_ff_13927:FAff port map(x=>p(332)(21),y=>p(333)(21),Cin=>p(334)(21),clock=>clock,reset=>reset,s=>p(351)(21),cout=>p(352)(22));
FA_ff_13928:FAff port map(x=>p(332)(22),y=>p(333)(22),Cin=>p(334)(22),clock=>clock,reset=>reset,s=>p(351)(22),cout=>p(352)(23));
FA_ff_13929:FAff port map(x=>p(332)(23),y=>p(333)(23),Cin=>p(334)(23),clock=>clock,reset=>reset,s=>p(351)(23),cout=>p(352)(24));
FA_ff_13930:FAff port map(x=>p(332)(24),y=>p(333)(24),Cin=>p(334)(24),clock=>clock,reset=>reset,s=>p(351)(24),cout=>p(352)(25));
FA_ff_13931:FAff port map(x=>p(332)(25),y=>p(333)(25),Cin=>p(334)(25),clock=>clock,reset=>reset,s=>p(351)(25),cout=>p(352)(26));
FA_ff_13932:FAff port map(x=>p(332)(26),y=>p(333)(26),Cin=>p(334)(26),clock=>clock,reset=>reset,s=>p(351)(26),cout=>p(352)(27));
FA_ff_13933:FAff port map(x=>p(332)(27),y=>p(333)(27),Cin=>p(334)(27),clock=>clock,reset=>reset,s=>p(351)(27),cout=>p(352)(28));
FA_ff_13934:FAff port map(x=>p(332)(28),y=>p(333)(28),Cin=>p(334)(28),clock=>clock,reset=>reset,s=>p(351)(28),cout=>p(352)(29));
FA_ff_13935:FAff port map(x=>p(332)(29),y=>p(333)(29),Cin=>p(334)(29),clock=>clock,reset=>reset,s=>p(351)(29),cout=>p(352)(30));
FA_ff_13936:FAff port map(x=>p(332)(30),y=>p(333)(30),Cin=>p(334)(30),clock=>clock,reset=>reset,s=>p(351)(30),cout=>p(352)(31));
FA_ff_13937:FAff port map(x=>p(332)(31),y=>p(333)(31),Cin=>p(334)(31),clock=>clock,reset=>reset,s=>p(351)(31),cout=>p(352)(32));
FA_ff_13938:FAff port map(x=>p(332)(32),y=>p(333)(32),Cin=>p(334)(32),clock=>clock,reset=>reset,s=>p(351)(32),cout=>p(352)(33));
FA_ff_13939:FAff port map(x=>p(332)(33),y=>p(333)(33),Cin=>p(334)(33),clock=>clock,reset=>reset,s=>p(351)(33),cout=>p(352)(34));
FA_ff_13940:FAff port map(x=>p(332)(34),y=>p(333)(34),Cin=>p(334)(34),clock=>clock,reset=>reset,s=>p(351)(34),cout=>p(352)(35));
FA_ff_13941:FAff port map(x=>p(332)(35),y=>p(333)(35),Cin=>p(334)(35),clock=>clock,reset=>reset,s=>p(351)(35),cout=>p(352)(36));
FA_ff_13942:FAff port map(x=>p(332)(36),y=>p(333)(36),Cin=>p(334)(36),clock=>clock,reset=>reset,s=>p(351)(36),cout=>p(352)(37));
FA_ff_13943:FAff port map(x=>p(332)(37),y=>p(333)(37),Cin=>p(334)(37),clock=>clock,reset=>reset,s=>p(351)(37),cout=>p(352)(38));
FA_ff_13944:FAff port map(x=>p(332)(38),y=>p(333)(38),Cin=>p(334)(38),clock=>clock,reset=>reset,s=>p(351)(38),cout=>p(352)(39));
FA_ff_13945:FAff port map(x=>p(332)(39),y=>p(333)(39),Cin=>p(334)(39),clock=>clock,reset=>reset,s=>p(351)(39),cout=>p(352)(40));
FA_ff_13946:FAff port map(x=>p(332)(40),y=>p(333)(40),Cin=>p(334)(40),clock=>clock,reset=>reset,s=>p(351)(40),cout=>p(352)(41));
FA_ff_13947:FAff port map(x=>p(332)(41),y=>p(333)(41),Cin=>p(334)(41),clock=>clock,reset=>reset,s=>p(351)(41),cout=>p(352)(42));
FA_ff_13948:FAff port map(x=>p(332)(42),y=>p(333)(42),Cin=>p(334)(42),clock=>clock,reset=>reset,s=>p(351)(42),cout=>p(352)(43));
FA_ff_13949:FAff port map(x=>p(332)(43),y=>p(333)(43),Cin=>p(334)(43),clock=>clock,reset=>reset,s=>p(351)(43),cout=>p(352)(44));
FA_ff_13950:FAff port map(x=>p(332)(44),y=>p(333)(44),Cin=>p(334)(44),clock=>clock,reset=>reset,s=>p(351)(44),cout=>p(352)(45));
FA_ff_13951:FAff port map(x=>p(332)(45),y=>p(333)(45),Cin=>p(334)(45),clock=>clock,reset=>reset,s=>p(351)(45),cout=>p(352)(46));
FA_ff_13952:FAff port map(x=>p(332)(46),y=>p(333)(46),Cin=>p(334)(46),clock=>clock,reset=>reset,s=>p(351)(46),cout=>p(352)(47));
FA_ff_13953:FAff port map(x=>p(332)(47),y=>p(333)(47),Cin=>p(334)(47),clock=>clock,reset=>reset,s=>p(351)(47),cout=>p(352)(48));
FA_ff_13954:FAff port map(x=>p(332)(48),y=>p(333)(48),Cin=>p(334)(48),clock=>clock,reset=>reset,s=>p(351)(48),cout=>p(352)(49));
FA_ff_13955:FAff port map(x=>p(332)(49),y=>p(333)(49),Cin=>p(334)(49),clock=>clock,reset=>reset,s=>p(351)(49),cout=>p(352)(50));
FA_ff_13956:FAff port map(x=>p(332)(50),y=>p(333)(50),Cin=>p(334)(50),clock=>clock,reset=>reset,s=>p(351)(50),cout=>p(352)(51));
FA_ff_13957:FAff port map(x=>p(332)(51),y=>p(333)(51),Cin=>p(334)(51),clock=>clock,reset=>reset,s=>p(351)(51),cout=>p(352)(52));
FA_ff_13958:FAff port map(x=>p(332)(52),y=>p(333)(52),Cin=>p(334)(52),clock=>clock,reset=>reset,s=>p(351)(52),cout=>p(352)(53));
FA_ff_13959:FAff port map(x=>p(332)(53),y=>p(333)(53),Cin=>p(334)(53),clock=>clock,reset=>reset,s=>p(351)(53),cout=>p(352)(54));
FA_ff_13960:FAff port map(x=>p(332)(54),y=>p(333)(54),Cin=>p(334)(54),clock=>clock,reset=>reset,s=>p(351)(54),cout=>p(352)(55));
FA_ff_13961:FAff port map(x=>p(332)(55),y=>p(333)(55),Cin=>p(334)(55),clock=>clock,reset=>reset,s=>p(351)(55),cout=>p(352)(56));
FA_ff_13962:FAff port map(x=>p(332)(56),y=>p(333)(56),Cin=>p(334)(56),clock=>clock,reset=>reset,s=>p(351)(56),cout=>p(352)(57));
FA_ff_13963:FAff port map(x=>p(332)(57),y=>p(333)(57),Cin=>p(334)(57),clock=>clock,reset=>reset,s=>p(351)(57),cout=>p(352)(58));
FA_ff_13964:FAff port map(x=>p(332)(58),y=>p(333)(58),Cin=>p(334)(58),clock=>clock,reset=>reset,s=>p(351)(58),cout=>p(352)(59));
FA_ff_13965:FAff port map(x=>p(332)(59),y=>p(333)(59),Cin=>p(334)(59),clock=>clock,reset=>reset,s=>p(351)(59),cout=>p(352)(60));
FA_ff_13966:FAff port map(x=>p(332)(60),y=>p(333)(60),Cin=>p(334)(60),clock=>clock,reset=>reset,s=>p(351)(60),cout=>p(352)(61));
FA_ff_13967:FAff port map(x=>p(332)(61),y=>p(333)(61),Cin=>p(334)(61),clock=>clock,reset=>reset,s=>p(351)(61),cout=>p(352)(62));
FA_ff_13968:FAff port map(x=>p(332)(62),y=>p(333)(62),Cin=>p(334)(62),clock=>clock,reset=>reset,s=>p(351)(62),cout=>p(352)(63));
FA_ff_13969:FAff port map(x=>p(332)(63),y=>p(333)(63),Cin=>p(334)(63),clock=>clock,reset=>reset,s=>p(351)(63),cout=>p(352)(64));
FA_ff_13970:FAff port map(x=>p(332)(64),y=>p(333)(64),Cin=>p(334)(64),clock=>clock,reset=>reset,s=>p(351)(64),cout=>p(352)(65));
FA_ff_13971:FAff port map(x=>p(332)(65),y=>p(333)(65),Cin=>p(334)(65),clock=>clock,reset=>reset,s=>p(351)(65),cout=>p(352)(66));
FA_ff_13972:FAff port map(x=>p(332)(66),y=>p(333)(66),Cin=>p(334)(66),clock=>clock,reset=>reset,s=>p(351)(66),cout=>p(352)(67));
FA_ff_13973:FAff port map(x=>p(332)(67),y=>p(333)(67),Cin=>p(334)(67),clock=>clock,reset=>reset,s=>p(351)(67),cout=>p(352)(68));
FA_ff_13974:FAff port map(x=>p(332)(68),y=>p(333)(68),Cin=>p(334)(68),clock=>clock,reset=>reset,s=>p(351)(68),cout=>p(352)(69));
FA_ff_13975:FAff port map(x=>p(332)(69),y=>p(333)(69),Cin=>p(334)(69),clock=>clock,reset=>reset,s=>p(351)(69),cout=>p(352)(70));
FA_ff_13976:FAff port map(x=>p(332)(70),y=>p(333)(70),Cin=>p(334)(70),clock=>clock,reset=>reset,s=>p(351)(70),cout=>p(352)(71));
FA_ff_13977:FAff port map(x=>p(332)(71),y=>p(333)(71),Cin=>p(334)(71),clock=>clock,reset=>reset,s=>p(351)(71),cout=>p(352)(72));
FA_ff_13978:FAff port map(x=>p(332)(72),y=>p(333)(72),Cin=>p(334)(72),clock=>clock,reset=>reset,s=>p(351)(72),cout=>p(352)(73));
FA_ff_13979:FAff port map(x=>p(332)(73),y=>p(333)(73),Cin=>p(334)(73),clock=>clock,reset=>reset,s=>p(351)(73),cout=>p(352)(74));
FA_ff_13980:FAff port map(x=>p(332)(74),y=>p(333)(74),Cin=>p(334)(74),clock=>clock,reset=>reset,s=>p(351)(74),cout=>p(352)(75));
FA_ff_13981:FAff port map(x=>p(332)(75),y=>p(333)(75),Cin=>p(334)(75),clock=>clock,reset=>reset,s=>p(351)(75),cout=>p(352)(76));
FA_ff_13982:FAff port map(x=>p(332)(76),y=>p(333)(76),Cin=>p(334)(76),clock=>clock,reset=>reset,s=>p(351)(76),cout=>p(352)(77));
FA_ff_13983:FAff port map(x=>p(332)(77),y=>p(333)(77),Cin=>p(334)(77),clock=>clock,reset=>reset,s=>p(351)(77),cout=>p(352)(78));
FA_ff_13984:FAff port map(x=>p(332)(78),y=>p(333)(78),Cin=>p(334)(78),clock=>clock,reset=>reset,s=>p(351)(78),cout=>p(352)(79));
FA_ff_13985:FAff port map(x=>p(332)(79),y=>p(333)(79),Cin=>p(334)(79),clock=>clock,reset=>reset,s=>p(351)(79),cout=>p(352)(80));
FA_ff_13986:FAff port map(x=>p(332)(80),y=>p(333)(80),Cin=>p(334)(80),clock=>clock,reset=>reset,s=>p(351)(80),cout=>p(352)(81));
FA_ff_13987:FAff port map(x=>p(332)(81),y=>p(333)(81),Cin=>p(334)(81),clock=>clock,reset=>reset,s=>p(351)(81),cout=>p(352)(82));
FA_ff_13988:FAff port map(x=>p(332)(82),y=>p(333)(82),Cin=>p(334)(82),clock=>clock,reset=>reset,s=>p(351)(82),cout=>p(352)(83));
FA_ff_13989:FAff port map(x=>p(332)(83),y=>p(333)(83),Cin=>p(334)(83),clock=>clock,reset=>reset,s=>p(351)(83),cout=>p(352)(84));
FA_ff_13990:FAff port map(x=>p(332)(84),y=>p(333)(84),Cin=>p(334)(84),clock=>clock,reset=>reset,s=>p(351)(84),cout=>p(352)(85));
FA_ff_13991:FAff port map(x=>p(332)(85),y=>p(333)(85),Cin=>p(334)(85),clock=>clock,reset=>reset,s=>p(351)(85),cout=>p(352)(86));
FA_ff_13992:FAff port map(x=>p(332)(86),y=>p(333)(86),Cin=>p(334)(86),clock=>clock,reset=>reset,s=>p(351)(86),cout=>p(352)(87));
FA_ff_13993:FAff port map(x=>p(332)(87),y=>p(333)(87),Cin=>p(334)(87),clock=>clock,reset=>reset,s=>p(351)(87),cout=>p(352)(88));
FA_ff_13994:FAff port map(x=>p(332)(88),y=>p(333)(88),Cin=>p(334)(88),clock=>clock,reset=>reset,s=>p(351)(88),cout=>p(352)(89));
FA_ff_13995:FAff port map(x=>p(332)(89),y=>p(333)(89),Cin=>p(334)(89),clock=>clock,reset=>reset,s=>p(351)(89),cout=>p(352)(90));
FA_ff_13996:FAff port map(x=>p(332)(90),y=>p(333)(90),Cin=>p(334)(90),clock=>clock,reset=>reset,s=>p(351)(90),cout=>p(352)(91));
FA_ff_13997:FAff port map(x=>p(332)(91),y=>p(333)(91),Cin=>p(334)(91),clock=>clock,reset=>reset,s=>p(351)(91),cout=>p(352)(92));
FA_ff_13998:FAff port map(x=>p(332)(92),y=>p(333)(92),Cin=>p(334)(92),clock=>clock,reset=>reset,s=>p(351)(92),cout=>p(352)(93));
FA_ff_13999:FAff port map(x=>p(332)(93),y=>p(333)(93),Cin=>p(334)(93),clock=>clock,reset=>reset,s=>p(351)(93),cout=>p(352)(94));
FA_ff_14000:FAff port map(x=>p(332)(94),y=>p(333)(94),Cin=>p(334)(94),clock=>clock,reset=>reset,s=>p(351)(94),cout=>p(352)(95));
FA_ff_14001:FAff port map(x=>p(332)(95),y=>p(333)(95),Cin=>p(334)(95),clock=>clock,reset=>reset,s=>p(351)(95),cout=>p(352)(96));
FA_ff_14002:FAff port map(x=>p(332)(96),y=>p(333)(96),Cin=>p(334)(96),clock=>clock,reset=>reset,s=>p(351)(96),cout=>p(352)(97));
FA_ff_14003:FAff port map(x=>p(332)(97),y=>p(333)(97),Cin=>p(334)(97),clock=>clock,reset=>reset,s=>p(351)(97),cout=>p(352)(98));
FA_ff_14004:FAff port map(x=>p(332)(98),y=>p(333)(98),Cin=>p(334)(98),clock=>clock,reset=>reset,s=>p(351)(98),cout=>p(352)(99));
FA_ff_14005:FAff port map(x=>p(332)(99),y=>p(333)(99),Cin=>p(334)(99),clock=>clock,reset=>reset,s=>p(351)(99),cout=>p(352)(100));
FA_ff_14006:FAff port map(x=>p(332)(100),y=>p(333)(100),Cin=>p(334)(100),clock=>clock,reset=>reset,s=>p(351)(100),cout=>p(352)(101));
FA_ff_14007:FAff port map(x=>p(332)(101),y=>p(333)(101),Cin=>p(334)(101),clock=>clock,reset=>reset,s=>p(351)(101),cout=>p(352)(102));
FA_ff_14008:FAff port map(x=>p(332)(102),y=>p(333)(102),Cin=>p(334)(102),clock=>clock,reset=>reset,s=>p(351)(102),cout=>p(352)(103));
FA_ff_14009:FAff port map(x=>p(332)(103),y=>p(333)(103),Cin=>p(334)(103),clock=>clock,reset=>reset,s=>p(351)(103),cout=>p(352)(104));
FA_ff_14010:FAff port map(x=>p(332)(104),y=>p(333)(104),Cin=>p(334)(104),clock=>clock,reset=>reset,s=>p(351)(104),cout=>p(352)(105));
FA_ff_14011:FAff port map(x=>p(332)(105),y=>p(333)(105),Cin=>p(334)(105),clock=>clock,reset=>reset,s=>p(351)(105),cout=>p(352)(106));
FA_ff_14012:FAff port map(x=>p(332)(106),y=>p(333)(106),Cin=>p(334)(106),clock=>clock,reset=>reset,s=>p(351)(106),cout=>p(352)(107));
FA_ff_14013:FAff port map(x=>p(332)(107),y=>p(333)(107),Cin=>p(334)(107),clock=>clock,reset=>reset,s=>p(351)(107),cout=>p(352)(108));
FA_ff_14014:FAff port map(x=>p(332)(108),y=>p(333)(108),Cin=>p(334)(108),clock=>clock,reset=>reset,s=>p(351)(108),cout=>p(352)(109));
FA_ff_14015:FAff port map(x=>p(332)(109),y=>p(333)(109),Cin=>p(334)(109),clock=>clock,reset=>reset,s=>p(351)(109),cout=>p(352)(110));
FA_ff_14016:FAff port map(x=>p(332)(110),y=>p(333)(110),Cin=>p(334)(110),clock=>clock,reset=>reset,s=>p(351)(110),cout=>p(352)(111));
FA_ff_14017:FAff port map(x=>p(332)(111),y=>p(333)(111),Cin=>p(334)(111),clock=>clock,reset=>reset,s=>p(351)(111),cout=>p(352)(112));
FA_ff_14018:FAff port map(x=>p(332)(112),y=>p(333)(112),Cin=>p(334)(112),clock=>clock,reset=>reset,s=>p(351)(112),cout=>p(352)(113));
FA_ff_14019:FAff port map(x=>p(332)(113),y=>p(333)(113),Cin=>p(334)(113),clock=>clock,reset=>reset,s=>p(351)(113),cout=>p(352)(114));
FA_ff_14020:FAff port map(x=>p(332)(114),y=>p(333)(114),Cin=>p(334)(114),clock=>clock,reset=>reset,s=>p(351)(114),cout=>p(352)(115));
FA_ff_14021:FAff port map(x=>p(332)(115),y=>p(333)(115),Cin=>p(334)(115),clock=>clock,reset=>reset,s=>p(351)(115),cout=>p(352)(116));
FA_ff_14022:FAff port map(x=>p(332)(116),y=>p(333)(116),Cin=>p(334)(116),clock=>clock,reset=>reset,s=>p(351)(116),cout=>p(352)(117));
FA_ff_14023:FAff port map(x=>p(332)(117),y=>p(333)(117),Cin=>p(334)(117),clock=>clock,reset=>reset,s=>p(351)(117),cout=>p(352)(118));
FA_ff_14024:FAff port map(x=>p(332)(118),y=>p(333)(118),Cin=>p(334)(118),clock=>clock,reset=>reset,s=>p(351)(118),cout=>p(352)(119));
FA_ff_14025:FAff port map(x=>p(332)(119),y=>p(333)(119),Cin=>p(334)(119),clock=>clock,reset=>reset,s=>p(351)(119),cout=>p(352)(120));
FA_ff_14026:FAff port map(x=>p(332)(120),y=>p(333)(120),Cin=>p(334)(120),clock=>clock,reset=>reset,s=>p(351)(120),cout=>p(352)(121));
FA_ff_14027:FAff port map(x=>p(332)(121),y=>p(333)(121),Cin=>p(334)(121),clock=>clock,reset=>reset,s=>p(351)(121),cout=>p(352)(122));
FA_ff_14028:FAff port map(x=>p(332)(122),y=>p(333)(122),Cin=>p(334)(122),clock=>clock,reset=>reset,s=>p(351)(122),cout=>p(352)(123));
FA_ff_14029:FAff port map(x=>p(332)(123),y=>p(333)(123),Cin=>p(334)(123),clock=>clock,reset=>reset,s=>p(351)(123),cout=>p(352)(124));
FA_ff_14030:FAff port map(x=>p(332)(124),y=>p(333)(124),Cin=>p(334)(124),clock=>clock,reset=>reset,s=>p(351)(124),cout=>p(352)(125));
FA_ff_14031:FAff port map(x=>p(332)(125),y=>p(333)(125),Cin=>p(334)(125),clock=>clock,reset=>reset,s=>p(351)(125),cout=>p(352)(126));
FA_ff_14032:FAff port map(x=>p(332)(126),y=>p(333)(126),Cin=>p(334)(126),clock=>clock,reset=>reset,s=>p(351)(126),cout=>p(352)(127));
FA_ff_14033:FAff port map(x=>p(332)(127),y=>p(333)(127),Cin=>p(334)(127),clock=>clock,reset=>reset,s=>p(351)(127),cout=>p(352)(128));
FA_ff_14034:FAff port map(x=>p(332)(128),y=>p(333)(128),Cin=>p(334)(128),clock=>clock,reset=>reset,s=>p(351)(128),cout=>p(352)(129));
FA_ff_14035:FAff port map(x=>p(332)(129),y=>p(333)(129),Cin=>p(334)(129),clock=>clock,reset=>reset,s=>p(351)(129),cout=>p(352)(130));
HA_ff_89:HAff port map(x=>p(332)(130),y=>p(334)(130),clock=>clock,reset=>reset,s=>p(351)(130),c=>p(352)(131));
p(353)(0)<=p(335)(0);
p(353)(1)<=p(335)(1);
p(353)(2)<=p(335)(2);
p(353)(3)<=p(335)(3);
p(353)(4)<=p(335)(4);
p(353)(5)<=p(335)(5);
p(353)(6)<=p(335)(6);
p(353)(7)<=p(335)(7);
p(353)(8)<=p(335)(8);
p(353)(9)<=p(335)(9);
p(353)(10)<=p(335)(10);
p(353)(11)<=p(335)(11);
p(353)(12)<=p(335)(12);
p(353)(13)<=p(335)(13);
p(353)(14)<=p(335)(14);
p(353)(15)<=p(335)(15);
p(353)(16)<=p(335)(16);
p(353)(17)<=p(335)(17);
p(353)(18)<=p(335)(18);
p(353)(19)<=p(335)(19);
p(353)(20)<=p(335)(20);
p(353)(21)<=p(335)(21);
p(353)(22)<=p(335)(22);
p(353)(23)<=p(335)(23);
p(353)(24)<=p(335)(24);
p(353)(25)<=p(335)(25);
p(353)(26)<=p(335)(26);
p(353)(27)<=p(335)(27);
p(353)(28)<=p(335)(28);
p(353)(29)<=p(335)(29);
p(353)(30)<=p(335)(30);
p(353)(31)<=p(335)(31);
p(353)(32)<=p(335)(32);
p(353)(33)<=p(335)(33);
p(353)(34)<=p(335)(34);
p(353)(35)<=p(335)(35);
p(353)(36)<=p(335)(36);
p(353)(37)<=p(335)(37);
p(353)(38)<=p(335)(38);
p(353)(39)<=p(335)(39);
p(353)(40)<=p(335)(40);
p(353)(41)<=p(335)(41);
p(353)(42)<=p(335)(42);
p(353)(43)<=p(335)(43);
p(353)(44)<=p(335)(44);
p(353)(45)<=p(335)(45);
p(353)(46)<=p(335)(46);
p(353)(47)<=p(335)(47);
p(353)(48)<=p(335)(48);
p(353)(49)<=p(335)(49);
p(353)(50)<=p(335)(50);
p(353)(51)<=p(335)(51);
p(353)(52)<=p(335)(52);
p(353)(53)<=p(335)(53);
p(353)(54)<=p(335)(54);
p(353)(55)<=p(335)(55);
p(353)(56)<=p(335)(56);
p(353)(57)<=p(335)(57);
p(353)(58)<=p(335)(58);
p(353)(59)<=p(335)(59);
p(353)(60)<=p(335)(60);
p(353)(61)<=p(335)(61);
p(353)(62)<=p(335)(62);
p(353)(63)<=p(335)(63);
p(353)(64)<=p(335)(64);
p(353)(65)<=p(335)(65);
p(353)(66)<=p(335)(66);
p(353)(67)<=p(335)(67);
p(353)(68)<=p(335)(68);
p(353)(69)<=p(335)(69);
p(353)(70)<=p(335)(70);
p(353)(71)<=p(335)(71);
p(353)(72)<=p(335)(72);
p(353)(73)<=p(335)(73);
p(353)(74)<=p(335)(74);
p(353)(75)<=p(335)(75);
p(353)(76)<=p(335)(76);
p(353)(77)<=p(335)(77);
p(353)(78)<=p(335)(78);
p(353)(79)<=p(335)(79);
p(353)(80)<=p(335)(80);
p(353)(81)<=p(335)(81);
p(353)(82)<=p(335)(82);
p(353)(83)<=p(335)(83);
p(353)(84)<=p(335)(84);
p(353)(85)<=p(335)(85);
p(353)(86)<=p(335)(86);
p(353)(87)<=p(335)(87);
p(353)(88)<=p(335)(88);
p(353)(89)<=p(335)(89);
p(353)(90)<=p(335)(90);
p(353)(91)<=p(335)(91);
p(353)(92)<=p(335)(92);
p(353)(93)<=p(335)(93);
p(353)(94)<=p(335)(94);
p(353)(95)<=p(335)(95);
p(353)(96)<=p(335)(96);
p(353)(97)<=p(335)(97);
p(353)(98)<=p(335)(98);
p(353)(99)<=p(335)(99);
p(353)(100)<=p(335)(100);
p(353)(101)<=p(335)(101);
p(353)(102)<=p(335)(102);
p(353)(103)<=p(335)(103);
p(353)(104)<=p(335)(104);
p(353)(105)<=p(335)(105);
p(353)(106)<=p(335)(106);
p(353)(107)<=p(335)(107);
p(353)(108)<=p(335)(108);
p(353)(109)<=p(335)(109);
p(353)(110)<=p(335)(110);
p(353)(111)<=p(335)(111);
p(353)(112)<=p(335)(112);
p(353)(113)<=p(335)(113);
p(353)(114)<=p(335)(114);
p(353)(115)<=p(335)(115);
p(353)(116)<=p(335)(116);
p(353)(117)<=p(335)(117);
p(353)(118)<=p(335)(118);
p(353)(119)<=p(335)(119);
p(353)(120)<=p(335)(120);
p(353)(121)<=p(335)(121);
p(353)(122)<=p(335)(122);
p(353)(123)<=p(335)(123);
p(353)(124)<=p(335)(124);
p(353)(125)<=p(335)(125);
p(353)(126)<=p(335)(126);
p(353)(127)<=p(335)(127);
p(353)(128)<=p(335)(128);
p(353)(129)<=p(335)(129);
p(353)(130)<=p(335)(130);
p(353)(131)<=p(335)(131);
p(353)(132)<=p(335)(132);
p(353)(133)<=p(335)(133);
p(353)(134)<=p(335)(134);
p(354)(0)<=p(336)(0);
p(354)(1)<=p(336)(1);
p(354)(2)<=p(336)(2);
p(354)(3)<=p(336)(3);
p(354)(4)<=p(336)(4);
p(354)(5)<=p(336)(5);
p(354)(6)<=p(336)(6);
p(354)(7)<=p(336)(7);
p(354)(8)<=p(336)(8);
p(354)(9)<=p(336)(9);
p(354)(10)<=p(336)(10);
p(354)(11)<=p(336)(11);
p(354)(12)<=p(336)(12);
p(354)(13)<=p(336)(13);
p(354)(14)<=p(336)(14);
p(354)(15)<=p(336)(15);
p(354)(16)<=p(336)(16);
p(354)(17)<=p(336)(17);
p(354)(18)<=p(336)(18);
p(354)(19)<=p(336)(19);
p(354)(20)<=p(336)(20);
p(354)(21)<=p(336)(21);
p(354)(22)<=p(336)(22);
p(354)(23)<=p(336)(23);
p(354)(24)<=p(336)(24);
p(354)(25)<=p(336)(25);
p(354)(26)<=p(336)(26);
p(354)(27)<=p(336)(27);
p(354)(28)<=p(336)(28);
p(354)(29)<=p(336)(29);
p(354)(30)<=p(336)(30);
p(354)(31)<=p(336)(31);
p(354)(32)<=p(336)(32);
p(354)(33)<=p(336)(33);
p(354)(34)<=p(336)(34);
p(354)(35)<=p(336)(35);
p(354)(36)<=p(336)(36);
p(354)(37)<=p(336)(37);
p(354)(38)<=p(336)(38);
p(354)(39)<=p(336)(39);
p(354)(40)<=p(336)(40);
p(354)(41)<=p(336)(41);
p(354)(42)<=p(336)(42);
p(354)(43)<=p(336)(43);
p(354)(44)<=p(336)(44);
p(354)(45)<=p(336)(45);
p(354)(46)<=p(336)(46);
p(354)(47)<=p(336)(47);
p(354)(48)<=p(336)(48);
p(354)(49)<=p(336)(49);
p(354)(50)<=p(336)(50);
p(354)(51)<=p(336)(51);
p(354)(52)<=p(336)(52);
p(354)(53)<=p(336)(53);
p(354)(54)<=p(336)(54);
p(354)(55)<=p(336)(55);
p(354)(56)<=p(336)(56);
p(354)(57)<=p(336)(57);
p(354)(58)<=p(336)(58);
p(354)(59)<=p(336)(59);
p(354)(60)<=p(336)(60);
p(354)(61)<=p(336)(61);
p(354)(62)<=p(336)(62);
p(354)(63)<=p(336)(63);
p(354)(64)<=p(336)(64);
p(354)(65)<=p(336)(65);
p(354)(66)<=p(336)(66);
p(354)(67)<=p(336)(67);
p(354)(68)<=p(336)(68);
p(354)(69)<=p(336)(69);
p(354)(70)<=p(336)(70);
p(354)(71)<=p(336)(71);
p(354)(72)<=p(336)(72);
p(354)(73)<=p(336)(73);
p(354)(74)<=p(336)(74);
p(354)(75)<=p(336)(75);
p(354)(76)<=p(336)(76);
p(354)(77)<=p(336)(77);
p(354)(78)<=p(336)(78);
p(354)(79)<=p(336)(79);
p(354)(80)<=p(336)(80);
p(354)(81)<=p(336)(81);
p(354)(82)<=p(336)(82);
p(354)(83)<=p(336)(83);
p(354)(84)<=p(336)(84);
p(354)(85)<=p(336)(85);
p(354)(86)<=p(336)(86);
p(354)(87)<=p(336)(87);
p(354)(88)<=p(336)(88);
p(354)(89)<=p(336)(89);
p(354)(90)<=p(336)(90);
p(354)(91)<=p(336)(91);
p(354)(92)<=p(336)(92);
p(354)(93)<=p(336)(93);
p(354)(94)<=p(336)(94);
p(354)(95)<=p(336)(95);
p(354)(96)<=p(336)(96);
p(354)(97)<=p(336)(97);
p(354)(98)<=p(336)(98);
p(354)(99)<=p(336)(99);
p(354)(100)<=p(336)(100);
p(354)(101)<=p(336)(101);
p(354)(102)<=p(336)(102);
p(354)(103)<=p(336)(103);
p(354)(104)<=p(336)(104);
p(354)(105)<=p(336)(105);
p(354)(106)<=p(336)(106);
p(354)(107)<=p(336)(107);
p(354)(108)<=p(336)(108);
p(354)(109)<=p(336)(109);
p(354)(110)<=p(336)(110);
p(354)(111)<=p(336)(111);
p(354)(112)<=p(336)(112);
p(354)(113)<=p(336)(113);
p(354)(114)<=p(336)(114);
p(354)(115)<=p(336)(115);
p(354)(116)<=p(336)(116);
p(354)(117)<=p(336)(117);
p(354)(118)<=p(336)(118);
p(354)(119)<=p(336)(119);
p(354)(120)<=p(336)(120);
p(354)(121)<=p(336)(121);
p(354)(122)<=p(336)(122);
p(354)(123)<=p(336)(123);
p(354)(124)<=p(336)(124);
p(354)(125)<=p(336)(125);
p(354)(126)<=p(336)(126);
p(354)(127)<=p(336)(127);
p(354)(128)<=p(336)(128);
p(354)(129)<=p(336)(129);
p(354)(130)<=p(336)(130);
p(354)(131)<=p(336)(131);
p(354)(132)<=p(336)(132);
p(354)(133)<=p(336)(133);
p(354)(134)<=p(336)(134);
HA_ff_90:HAff port map(x=>p(337)(0),y=>p(339)(0),clock=>clock,reset=>reset,s=>p(355)(0),c=>p(356)(1));
FA_ff_14036:FAff port map(x=>p(337)(1),y=>p(338)(1),Cin=>p(339)(1),clock=>clock,reset=>reset,s=>p(355)(1),cout=>p(356)(2));
FA_ff_14037:FAff port map(x=>p(337)(2),y=>p(338)(2),Cin=>p(339)(2),clock=>clock,reset=>reset,s=>p(355)(2),cout=>p(356)(3));
FA_ff_14038:FAff port map(x=>p(337)(3),y=>p(338)(3),Cin=>p(339)(3),clock=>clock,reset=>reset,s=>p(355)(3),cout=>p(356)(4));
FA_ff_14039:FAff port map(x=>p(337)(4),y=>p(338)(4),Cin=>p(339)(4),clock=>clock,reset=>reset,s=>p(355)(4),cout=>p(356)(5));
FA_ff_14040:FAff port map(x=>p(337)(5),y=>p(338)(5),Cin=>p(339)(5),clock=>clock,reset=>reset,s=>p(355)(5),cout=>p(356)(6));
FA_ff_14041:FAff port map(x=>p(337)(6),y=>p(338)(6),Cin=>p(339)(6),clock=>clock,reset=>reset,s=>p(355)(6),cout=>p(356)(7));
FA_ff_14042:FAff port map(x=>p(337)(7),y=>p(338)(7),Cin=>p(339)(7),clock=>clock,reset=>reset,s=>p(355)(7),cout=>p(356)(8));
FA_ff_14043:FAff port map(x=>p(337)(8),y=>p(338)(8),Cin=>p(339)(8),clock=>clock,reset=>reset,s=>p(355)(8),cout=>p(356)(9));
FA_ff_14044:FAff port map(x=>p(337)(9),y=>p(338)(9),Cin=>p(339)(9),clock=>clock,reset=>reset,s=>p(355)(9),cout=>p(356)(10));
FA_ff_14045:FAff port map(x=>p(337)(10),y=>p(338)(10),Cin=>p(339)(10),clock=>clock,reset=>reset,s=>p(355)(10),cout=>p(356)(11));
FA_ff_14046:FAff port map(x=>p(337)(11),y=>p(338)(11),Cin=>p(339)(11),clock=>clock,reset=>reset,s=>p(355)(11),cout=>p(356)(12));
FA_ff_14047:FAff port map(x=>p(337)(12),y=>p(338)(12),Cin=>p(339)(12),clock=>clock,reset=>reset,s=>p(355)(12),cout=>p(356)(13));
FA_ff_14048:FAff port map(x=>p(337)(13),y=>p(338)(13),Cin=>p(339)(13),clock=>clock,reset=>reset,s=>p(355)(13),cout=>p(356)(14));
FA_ff_14049:FAff port map(x=>p(337)(14),y=>p(338)(14),Cin=>p(339)(14),clock=>clock,reset=>reset,s=>p(355)(14),cout=>p(356)(15));
FA_ff_14050:FAff port map(x=>p(337)(15),y=>p(338)(15),Cin=>p(339)(15),clock=>clock,reset=>reset,s=>p(355)(15),cout=>p(356)(16));
FA_ff_14051:FAff port map(x=>p(337)(16),y=>p(338)(16),Cin=>p(339)(16),clock=>clock,reset=>reset,s=>p(355)(16),cout=>p(356)(17));
FA_ff_14052:FAff port map(x=>p(337)(17),y=>p(338)(17),Cin=>p(339)(17),clock=>clock,reset=>reset,s=>p(355)(17),cout=>p(356)(18));
FA_ff_14053:FAff port map(x=>p(337)(18),y=>p(338)(18),Cin=>p(339)(18),clock=>clock,reset=>reset,s=>p(355)(18),cout=>p(356)(19));
FA_ff_14054:FAff port map(x=>p(337)(19),y=>p(338)(19),Cin=>p(339)(19),clock=>clock,reset=>reset,s=>p(355)(19),cout=>p(356)(20));
FA_ff_14055:FAff port map(x=>p(337)(20),y=>p(338)(20),Cin=>p(339)(20),clock=>clock,reset=>reset,s=>p(355)(20),cout=>p(356)(21));
FA_ff_14056:FAff port map(x=>p(337)(21),y=>p(338)(21),Cin=>p(339)(21),clock=>clock,reset=>reset,s=>p(355)(21),cout=>p(356)(22));
FA_ff_14057:FAff port map(x=>p(337)(22),y=>p(338)(22),Cin=>p(339)(22),clock=>clock,reset=>reset,s=>p(355)(22),cout=>p(356)(23));
FA_ff_14058:FAff port map(x=>p(337)(23),y=>p(338)(23),Cin=>p(339)(23),clock=>clock,reset=>reset,s=>p(355)(23),cout=>p(356)(24));
FA_ff_14059:FAff port map(x=>p(337)(24),y=>p(338)(24),Cin=>p(339)(24),clock=>clock,reset=>reset,s=>p(355)(24),cout=>p(356)(25));
FA_ff_14060:FAff port map(x=>p(337)(25),y=>p(338)(25),Cin=>p(339)(25),clock=>clock,reset=>reset,s=>p(355)(25),cout=>p(356)(26));
FA_ff_14061:FAff port map(x=>p(337)(26),y=>p(338)(26),Cin=>p(339)(26),clock=>clock,reset=>reset,s=>p(355)(26),cout=>p(356)(27));
FA_ff_14062:FAff port map(x=>p(337)(27),y=>p(338)(27),Cin=>p(339)(27),clock=>clock,reset=>reset,s=>p(355)(27),cout=>p(356)(28));
FA_ff_14063:FAff port map(x=>p(337)(28),y=>p(338)(28),Cin=>p(339)(28),clock=>clock,reset=>reset,s=>p(355)(28),cout=>p(356)(29));
FA_ff_14064:FAff port map(x=>p(337)(29),y=>p(338)(29),Cin=>p(339)(29),clock=>clock,reset=>reset,s=>p(355)(29),cout=>p(356)(30));
FA_ff_14065:FAff port map(x=>p(337)(30),y=>p(338)(30),Cin=>p(339)(30),clock=>clock,reset=>reset,s=>p(355)(30),cout=>p(356)(31));
FA_ff_14066:FAff port map(x=>p(337)(31),y=>p(338)(31),Cin=>p(339)(31),clock=>clock,reset=>reset,s=>p(355)(31),cout=>p(356)(32));
FA_ff_14067:FAff port map(x=>p(337)(32),y=>p(338)(32),Cin=>p(339)(32),clock=>clock,reset=>reset,s=>p(355)(32),cout=>p(356)(33));
FA_ff_14068:FAff port map(x=>p(337)(33),y=>p(338)(33),Cin=>p(339)(33),clock=>clock,reset=>reset,s=>p(355)(33),cout=>p(356)(34));
FA_ff_14069:FAff port map(x=>p(337)(34),y=>p(338)(34),Cin=>p(339)(34),clock=>clock,reset=>reset,s=>p(355)(34),cout=>p(356)(35));
FA_ff_14070:FAff port map(x=>p(337)(35),y=>p(338)(35),Cin=>p(339)(35),clock=>clock,reset=>reset,s=>p(355)(35),cout=>p(356)(36));
FA_ff_14071:FAff port map(x=>p(337)(36),y=>p(338)(36),Cin=>p(339)(36),clock=>clock,reset=>reset,s=>p(355)(36),cout=>p(356)(37));
FA_ff_14072:FAff port map(x=>p(337)(37),y=>p(338)(37),Cin=>p(339)(37),clock=>clock,reset=>reset,s=>p(355)(37),cout=>p(356)(38));
FA_ff_14073:FAff port map(x=>p(337)(38),y=>p(338)(38),Cin=>p(339)(38),clock=>clock,reset=>reset,s=>p(355)(38),cout=>p(356)(39));
FA_ff_14074:FAff port map(x=>p(337)(39),y=>p(338)(39),Cin=>p(339)(39),clock=>clock,reset=>reset,s=>p(355)(39),cout=>p(356)(40));
FA_ff_14075:FAff port map(x=>p(337)(40),y=>p(338)(40),Cin=>p(339)(40),clock=>clock,reset=>reset,s=>p(355)(40),cout=>p(356)(41));
FA_ff_14076:FAff port map(x=>p(337)(41),y=>p(338)(41),Cin=>p(339)(41),clock=>clock,reset=>reset,s=>p(355)(41),cout=>p(356)(42));
FA_ff_14077:FAff port map(x=>p(337)(42),y=>p(338)(42),Cin=>p(339)(42),clock=>clock,reset=>reset,s=>p(355)(42),cout=>p(356)(43));
FA_ff_14078:FAff port map(x=>p(337)(43),y=>p(338)(43),Cin=>p(339)(43),clock=>clock,reset=>reset,s=>p(355)(43),cout=>p(356)(44));
FA_ff_14079:FAff port map(x=>p(337)(44),y=>p(338)(44),Cin=>p(339)(44),clock=>clock,reset=>reset,s=>p(355)(44),cout=>p(356)(45));
FA_ff_14080:FAff port map(x=>p(337)(45),y=>p(338)(45),Cin=>p(339)(45),clock=>clock,reset=>reset,s=>p(355)(45),cout=>p(356)(46));
FA_ff_14081:FAff port map(x=>p(337)(46),y=>p(338)(46),Cin=>p(339)(46),clock=>clock,reset=>reset,s=>p(355)(46),cout=>p(356)(47));
FA_ff_14082:FAff port map(x=>p(337)(47),y=>p(338)(47),Cin=>p(339)(47),clock=>clock,reset=>reset,s=>p(355)(47),cout=>p(356)(48));
FA_ff_14083:FAff port map(x=>p(337)(48),y=>p(338)(48),Cin=>p(339)(48),clock=>clock,reset=>reset,s=>p(355)(48),cout=>p(356)(49));
FA_ff_14084:FAff port map(x=>p(337)(49),y=>p(338)(49),Cin=>p(339)(49),clock=>clock,reset=>reset,s=>p(355)(49),cout=>p(356)(50));
FA_ff_14085:FAff port map(x=>p(337)(50),y=>p(338)(50),Cin=>p(339)(50),clock=>clock,reset=>reset,s=>p(355)(50),cout=>p(356)(51));
FA_ff_14086:FAff port map(x=>p(337)(51),y=>p(338)(51),Cin=>p(339)(51),clock=>clock,reset=>reset,s=>p(355)(51),cout=>p(356)(52));
FA_ff_14087:FAff port map(x=>p(337)(52),y=>p(338)(52),Cin=>p(339)(52),clock=>clock,reset=>reset,s=>p(355)(52),cout=>p(356)(53));
FA_ff_14088:FAff port map(x=>p(337)(53),y=>p(338)(53),Cin=>p(339)(53),clock=>clock,reset=>reset,s=>p(355)(53),cout=>p(356)(54));
FA_ff_14089:FAff port map(x=>p(337)(54),y=>p(338)(54),Cin=>p(339)(54),clock=>clock,reset=>reset,s=>p(355)(54),cout=>p(356)(55));
FA_ff_14090:FAff port map(x=>p(337)(55),y=>p(338)(55),Cin=>p(339)(55),clock=>clock,reset=>reset,s=>p(355)(55),cout=>p(356)(56));
FA_ff_14091:FAff port map(x=>p(337)(56),y=>p(338)(56),Cin=>p(339)(56),clock=>clock,reset=>reset,s=>p(355)(56),cout=>p(356)(57));
FA_ff_14092:FAff port map(x=>p(337)(57),y=>p(338)(57),Cin=>p(339)(57),clock=>clock,reset=>reset,s=>p(355)(57),cout=>p(356)(58));
FA_ff_14093:FAff port map(x=>p(337)(58),y=>p(338)(58),Cin=>p(339)(58),clock=>clock,reset=>reset,s=>p(355)(58),cout=>p(356)(59));
FA_ff_14094:FAff port map(x=>p(337)(59),y=>p(338)(59),Cin=>p(339)(59),clock=>clock,reset=>reset,s=>p(355)(59),cout=>p(356)(60));
FA_ff_14095:FAff port map(x=>p(337)(60),y=>p(338)(60),Cin=>p(339)(60),clock=>clock,reset=>reset,s=>p(355)(60),cout=>p(356)(61));
FA_ff_14096:FAff port map(x=>p(337)(61),y=>p(338)(61),Cin=>p(339)(61),clock=>clock,reset=>reset,s=>p(355)(61),cout=>p(356)(62));
FA_ff_14097:FAff port map(x=>p(337)(62),y=>p(338)(62),Cin=>p(339)(62),clock=>clock,reset=>reset,s=>p(355)(62),cout=>p(356)(63));
FA_ff_14098:FAff port map(x=>p(337)(63),y=>p(338)(63),Cin=>p(339)(63),clock=>clock,reset=>reset,s=>p(355)(63),cout=>p(356)(64));
FA_ff_14099:FAff port map(x=>p(337)(64),y=>p(338)(64),Cin=>p(339)(64),clock=>clock,reset=>reset,s=>p(355)(64),cout=>p(356)(65));
FA_ff_14100:FAff port map(x=>p(337)(65),y=>p(338)(65),Cin=>p(339)(65),clock=>clock,reset=>reset,s=>p(355)(65),cout=>p(356)(66));
FA_ff_14101:FAff port map(x=>p(337)(66),y=>p(338)(66),Cin=>p(339)(66),clock=>clock,reset=>reset,s=>p(355)(66),cout=>p(356)(67));
FA_ff_14102:FAff port map(x=>p(337)(67),y=>p(338)(67),Cin=>p(339)(67),clock=>clock,reset=>reset,s=>p(355)(67),cout=>p(356)(68));
FA_ff_14103:FAff port map(x=>p(337)(68),y=>p(338)(68),Cin=>p(339)(68),clock=>clock,reset=>reset,s=>p(355)(68),cout=>p(356)(69));
FA_ff_14104:FAff port map(x=>p(337)(69),y=>p(338)(69),Cin=>p(339)(69),clock=>clock,reset=>reset,s=>p(355)(69),cout=>p(356)(70));
FA_ff_14105:FAff port map(x=>p(337)(70),y=>p(338)(70),Cin=>p(339)(70),clock=>clock,reset=>reset,s=>p(355)(70),cout=>p(356)(71));
FA_ff_14106:FAff port map(x=>p(337)(71),y=>p(338)(71),Cin=>p(339)(71),clock=>clock,reset=>reset,s=>p(355)(71),cout=>p(356)(72));
FA_ff_14107:FAff port map(x=>p(337)(72),y=>p(338)(72),Cin=>p(339)(72),clock=>clock,reset=>reset,s=>p(355)(72),cout=>p(356)(73));
FA_ff_14108:FAff port map(x=>p(337)(73),y=>p(338)(73),Cin=>p(339)(73),clock=>clock,reset=>reset,s=>p(355)(73),cout=>p(356)(74));
FA_ff_14109:FAff port map(x=>p(337)(74),y=>p(338)(74),Cin=>p(339)(74),clock=>clock,reset=>reset,s=>p(355)(74),cout=>p(356)(75));
FA_ff_14110:FAff port map(x=>p(337)(75),y=>p(338)(75),Cin=>p(339)(75),clock=>clock,reset=>reset,s=>p(355)(75),cout=>p(356)(76));
FA_ff_14111:FAff port map(x=>p(337)(76),y=>p(338)(76),Cin=>p(339)(76),clock=>clock,reset=>reset,s=>p(355)(76),cout=>p(356)(77));
FA_ff_14112:FAff port map(x=>p(337)(77),y=>p(338)(77),Cin=>p(339)(77),clock=>clock,reset=>reset,s=>p(355)(77),cout=>p(356)(78));
FA_ff_14113:FAff port map(x=>p(337)(78),y=>p(338)(78),Cin=>p(339)(78),clock=>clock,reset=>reset,s=>p(355)(78),cout=>p(356)(79));
FA_ff_14114:FAff port map(x=>p(337)(79),y=>p(338)(79),Cin=>p(339)(79),clock=>clock,reset=>reset,s=>p(355)(79),cout=>p(356)(80));
FA_ff_14115:FAff port map(x=>p(337)(80),y=>p(338)(80),Cin=>p(339)(80),clock=>clock,reset=>reset,s=>p(355)(80),cout=>p(356)(81));
FA_ff_14116:FAff port map(x=>p(337)(81),y=>p(338)(81),Cin=>p(339)(81),clock=>clock,reset=>reset,s=>p(355)(81),cout=>p(356)(82));
FA_ff_14117:FAff port map(x=>p(337)(82),y=>p(338)(82),Cin=>p(339)(82),clock=>clock,reset=>reset,s=>p(355)(82),cout=>p(356)(83));
FA_ff_14118:FAff port map(x=>p(337)(83),y=>p(338)(83),Cin=>p(339)(83),clock=>clock,reset=>reset,s=>p(355)(83),cout=>p(356)(84));
FA_ff_14119:FAff port map(x=>p(337)(84),y=>p(338)(84),Cin=>p(339)(84),clock=>clock,reset=>reset,s=>p(355)(84),cout=>p(356)(85));
FA_ff_14120:FAff port map(x=>p(337)(85),y=>p(338)(85),Cin=>p(339)(85),clock=>clock,reset=>reset,s=>p(355)(85),cout=>p(356)(86));
FA_ff_14121:FAff port map(x=>p(337)(86),y=>p(338)(86),Cin=>p(339)(86),clock=>clock,reset=>reset,s=>p(355)(86),cout=>p(356)(87));
FA_ff_14122:FAff port map(x=>p(337)(87),y=>p(338)(87),Cin=>p(339)(87),clock=>clock,reset=>reset,s=>p(355)(87),cout=>p(356)(88));
FA_ff_14123:FAff port map(x=>p(337)(88),y=>p(338)(88),Cin=>p(339)(88),clock=>clock,reset=>reset,s=>p(355)(88),cout=>p(356)(89));
FA_ff_14124:FAff port map(x=>p(337)(89),y=>p(338)(89),Cin=>p(339)(89),clock=>clock,reset=>reset,s=>p(355)(89),cout=>p(356)(90));
FA_ff_14125:FAff port map(x=>p(337)(90),y=>p(338)(90),Cin=>p(339)(90),clock=>clock,reset=>reset,s=>p(355)(90),cout=>p(356)(91));
FA_ff_14126:FAff port map(x=>p(337)(91),y=>p(338)(91),Cin=>p(339)(91),clock=>clock,reset=>reset,s=>p(355)(91),cout=>p(356)(92));
FA_ff_14127:FAff port map(x=>p(337)(92),y=>p(338)(92),Cin=>p(339)(92),clock=>clock,reset=>reset,s=>p(355)(92),cout=>p(356)(93));
FA_ff_14128:FAff port map(x=>p(337)(93),y=>p(338)(93),Cin=>p(339)(93),clock=>clock,reset=>reset,s=>p(355)(93),cout=>p(356)(94));
FA_ff_14129:FAff port map(x=>p(337)(94),y=>p(338)(94),Cin=>p(339)(94),clock=>clock,reset=>reset,s=>p(355)(94),cout=>p(356)(95));
FA_ff_14130:FAff port map(x=>p(337)(95),y=>p(338)(95),Cin=>p(339)(95),clock=>clock,reset=>reset,s=>p(355)(95),cout=>p(356)(96));
FA_ff_14131:FAff port map(x=>p(337)(96),y=>p(338)(96),Cin=>p(339)(96),clock=>clock,reset=>reset,s=>p(355)(96),cout=>p(356)(97));
FA_ff_14132:FAff port map(x=>p(337)(97),y=>p(338)(97),Cin=>p(339)(97),clock=>clock,reset=>reset,s=>p(355)(97),cout=>p(356)(98));
FA_ff_14133:FAff port map(x=>p(337)(98),y=>p(338)(98),Cin=>p(339)(98),clock=>clock,reset=>reset,s=>p(355)(98),cout=>p(356)(99));
FA_ff_14134:FAff port map(x=>p(337)(99),y=>p(338)(99),Cin=>p(339)(99),clock=>clock,reset=>reset,s=>p(355)(99),cout=>p(356)(100));
FA_ff_14135:FAff port map(x=>p(337)(100),y=>p(338)(100),Cin=>p(339)(100),clock=>clock,reset=>reset,s=>p(355)(100),cout=>p(356)(101));
FA_ff_14136:FAff port map(x=>p(337)(101),y=>p(338)(101),Cin=>p(339)(101),clock=>clock,reset=>reset,s=>p(355)(101),cout=>p(356)(102));
FA_ff_14137:FAff port map(x=>p(337)(102),y=>p(338)(102),Cin=>p(339)(102),clock=>clock,reset=>reset,s=>p(355)(102),cout=>p(356)(103));
FA_ff_14138:FAff port map(x=>p(337)(103),y=>p(338)(103),Cin=>p(339)(103),clock=>clock,reset=>reset,s=>p(355)(103),cout=>p(356)(104));
FA_ff_14139:FAff port map(x=>p(337)(104),y=>p(338)(104),Cin=>p(339)(104),clock=>clock,reset=>reset,s=>p(355)(104),cout=>p(356)(105));
FA_ff_14140:FAff port map(x=>p(337)(105),y=>p(338)(105),Cin=>p(339)(105),clock=>clock,reset=>reset,s=>p(355)(105),cout=>p(356)(106));
FA_ff_14141:FAff port map(x=>p(337)(106),y=>p(338)(106),Cin=>p(339)(106),clock=>clock,reset=>reset,s=>p(355)(106),cout=>p(356)(107));
FA_ff_14142:FAff port map(x=>p(337)(107),y=>p(338)(107),Cin=>p(339)(107),clock=>clock,reset=>reset,s=>p(355)(107),cout=>p(356)(108));
FA_ff_14143:FAff port map(x=>p(337)(108),y=>p(338)(108),Cin=>p(339)(108),clock=>clock,reset=>reset,s=>p(355)(108),cout=>p(356)(109));
FA_ff_14144:FAff port map(x=>p(337)(109),y=>p(338)(109),Cin=>p(339)(109),clock=>clock,reset=>reset,s=>p(355)(109),cout=>p(356)(110));
FA_ff_14145:FAff port map(x=>p(337)(110),y=>p(338)(110),Cin=>p(339)(110),clock=>clock,reset=>reset,s=>p(355)(110),cout=>p(356)(111));
FA_ff_14146:FAff port map(x=>p(337)(111),y=>p(338)(111),Cin=>p(339)(111),clock=>clock,reset=>reset,s=>p(355)(111),cout=>p(356)(112));
FA_ff_14147:FAff port map(x=>p(337)(112),y=>p(338)(112),Cin=>p(339)(112),clock=>clock,reset=>reset,s=>p(355)(112),cout=>p(356)(113));
FA_ff_14148:FAff port map(x=>p(337)(113),y=>p(338)(113),Cin=>p(339)(113),clock=>clock,reset=>reset,s=>p(355)(113),cout=>p(356)(114));
FA_ff_14149:FAff port map(x=>p(337)(114),y=>p(338)(114),Cin=>p(339)(114),clock=>clock,reset=>reset,s=>p(355)(114),cout=>p(356)(115));
FA_ff_14150:FAff port map(x=>p(337)(115),y=>p(338)(115),Cin=>p(339)(115),clock=>clock,reset=>reset,s=>p(355)(115),cout=>p(356)(116));
FA_ff_14151:FAff port map(x=>p(337)(116),y=>p(338)(116),Cin=>p(339)(116),clock=>clock,reset=>reset,s=>p(355)(116),cout=>p(356)(117));
FA_ff_14152:FAff port map(x=>p(337)(117),y=>p(338)(117),Cin=>p(339)(117),clock=>clock,reset=>reset,s=>p(355)(117),cout=>p(356)(118));
FA_ff_14153:FAff port map(x=>p(337)(118),y=>p(338)(118),Cin=>p(339)(118),clock=>clock,reset=>reset,s=>p(355)(118),cout=>p(356)(119));
FA_ff_14154:FAff port map(x=>p(337)(119),y=>p(338)(119),Cin=>p(339)(119),clock=>clock,reset=>reset,s=>p(355)(119),cout=>p(356)(120));
FA_ff_14155:FAff port map(x=>p(337)(120),y=>p(338)(120),Cin=>p(339)(120),clock=>clock,reset=>reset,s=>p(355)(120),cout=>p(356)(121));
FA_ff_14156:FAff port map(x=>p(337)(121),y=>p(338)(121),Cin=>p(339)(121),clock=>clock,reset=>reset,s=>p(355)(121),cout=>p(356)(122));
FA_ff_14157:FAff port map(x=>p(337)(122),y=>p(338)(122),Cin=>p(339)(122),clock=>clock,reset=>reset,s=>p(355)(122),cout=>p(356)(123));
FA_ff_14158:FAff port map(x=>p(337)(123),y=>p(338)(123),Cin=>p(339)(123),clock=>clock,reset=>reset,s=>p(355)(123),cout=>p(356)(124));
FA_ff_14159:FAff port map(x=>p(337)(124),y=>p(338)(124),Cin=>p(339)(124),clock=>clock,reset=>reset,s=>p(355)(124),cout=>p(356)(125));
FA_ff_14160:FAff port map(x=>p(337)(125),y=>p(338)(125),Cin=>p(339)(125),clock=>clock,reset=>reset,s=>p(355)(125),cout=>p(356)(126));
FA_ff_14161:FAff port map(x=>p(337)(126),y=>p(338)(126),Cin=>p(339)(126),clock=>clock,reset=>reset,s=>p(355)(126),cout=>p(356)(127));
FA_ff_14162:FAff port map(x=>p(337)(127),y=>p(338)(127),Cin=>p(339)(127),clock=>clock,reset=>reset,s=>p(355)(127),cout=>p(356)(128));
FA_ff_14163:FAff port map(x=>p(337)(128),y=>p(338)(128),Cin=>p(339)(128),clock=>clock,reset=>reset,s=>p(355)(128),cout=>p(356)(129));
FA_ff_14164:FAff port map(x=>p(337)(129),y=>p(338)(129),Cin=>p(339)(129),clock=>clock,reset=>reset,s=>p(355)(129),cout=>p(356)(130));
FA_ff_14165:FAff port map(x=>p(337)(130),y=>p(338)(130),Cin=>p(339)(130),clock=>clock,reset=>reset,s=>p(355)(130),cout=>p(356)(131));
p(357)(0)<=p(341)(0);
HA_ff_91:HAff port map(x=>p(341)(1),y=>p(342)(1),clock=>clock,reset=>reset,s=>p(357)(1),c=>p(358)(2));
FA_ff_14166:FAff port map(x=>p(340)(2),y=>p(341)(2),Cin=>p(342)(2),clock=>clock,reset=>reset,s=>p(357)(2),cout=>p(358)(3));
FA_ff_14167:FAff port map(x=>p(340)(3),y=>p(341)(3),Cin=>p(342)(3),clock=>clock,reset=>reset,s=>p(357)(3),cout=>p(358)(4));
FA_ff_14168:FAff port map(x=>p(340)(4),y=>p(341)(4),Cin=>p(342)(4),clock=>clock,reset=>reset,s=>p(357)(4),cout=>p(358)(5));
FA_ff_14169:FAff port map(x=>p(340)(5),y=>p(341)(5),Cin=>p(342)(5),clock=>clock,reset=>reset,s=>p(357)(5),cout=>p(358)(6));
FA_ff_14170:FAff port map(x=>p(340)(6),y=>p(341)(6),Cin=>p(342)(6),clock=>clock,reset=>reset,s=>p(357)(6),cout=>p(358)(7));
FA_ff_14171:FAff port map(x=>p(340)(7),y=>p(341)(7),Cin=>p(342)(7),clock=>clock,reset=>reset,s=>p(357)(7),cout=>p(358)(8));
FA_ff_14172:FAff port map(x=>p(340)(8),y=>p(341)(8),Cin=>p(342)(8),clock=>clock,reset=>reset,s=>p(357)(8),cout=>p(358)(9));
FA_ff_14173:FAff port map(x=>p(340)(9),y=>p(341)(9),Cin=>p(342)(9),clock=>clock,reset=>reset,s=>p(357)(9),cout=>p(358)(10));
FA_ff_14174:FAff port map(x=>p(340)(10),y=>p(341)(10),Cin=>p(342)(10),clock=>clock,reset=>reset,s=>p(357)(10),cout=>p(358)(11));
FA_ff_14175:FAff port map(x=>p(340)(11),y=>p(341)(11),Cin=>p(342)(11),clock=>clock,reset=>reset,s=>p(357)(11),cout=>p(358)(12));
FA_ff_14176:FAff port map(x=>p(340)(12),y=>p(341)(12),Cin=>p(342)(12),clock=>clock,reset=>reset,s=>p(357)(12),cout=>p(358)(13));
FA_ff_14177:FAff port map(x=>p(340)(13),y=>p(341)(13),Cin=>p(342)(13),clock=>clock,reset=>reset,s=>p(357)(13),cout=>p(358)(14));
FA_ff_14178:FAff port map(x=>p(340)(14),y=>p(341)(14),Cin=>p(342)(14),clock=>clock,reset=>reset,s=>p(357)(14),cout=>p(358)(15));
FA_ff_14179:FAff port map(x=>p(340)(15),y=>p(341)(15),Cin=>p(342)(15),clock=>clock,reset=>reset,s=>p(357)(15),cout=>p(358)(16));
FA_ff_14180:FAff port map(x=>p(340)(16),y=>p(341)(16),Cin=>p(342)(16),clock=>clock,reset=>reset,s=>p(357)(16),cout=>p(358)(17));
FA_ff_14181:FAff port map(x=>p(340)(17),y=>p(341)(17),Cin=>p(342)(17),clock=>clock,reset=>reset,s=>p(357)(17),cout=>p(358)(18));
FA_ff_14182:FAff port map(x=>p(340)(18),y=>p(341)(18),Cin=>p(342)(18),clock=>clock,reset=>reset,s=>p(357)(18),cout=>p(358)(19));
FA_ff_14183:FAff port map(x=>p(340)(19),y=>p(341)(19),Cin=>p(342)(19),clock=>clock,reset=>reset,s=>p(357)(19),cout=>p(358)(20));
FA_ff_14184:FAff port map(x=>p(340)(20),y=>p(341)(20),Cin=>p(342)(20),clock=>clock,reset=>reset,s=>p(357)(20),cout=>p(358)(21));
FA_ff_14185:FAff port map(x=>p(340)(21),y=>p(341)(21),Cin=>p(342)(21),clock=>clock,reset=>reset,s=>p(357)(21),cout=>p(358)(22));
FA_ff_14186:FAff port map(x=>p(340)(22),y=>p(341)(22),Cin=>p(342)(22),clock=>clock,reset=>reset,s=>p(357)(22),cout=>p(358)(23));
FA_ff_14187:FAff port map(x=>p(340)(23),y=>p(341)(23),Cin=>p(342)(23),clock=>clock,reset=>reset,s=>p(357)(23),cout=>p(358)(24));
FA_ff_14188:FAff port map(x=>p(340)(24),y=>p(341)(24),Cin=>p(342)(24),clock=>clock,reset=>reset,s=>p(357)(24),cout=>p(358)(25));
FA_ff_14189:FAff port map(x=>p(340)(25),y=>p(341)(25),Cin=>p(342)(25),clock=>clock,reset=>reset,s=>p(357)(25),cout=>p(358)(26));
FA_ff_14190:FAff port map(x=>p(340)(26),y=>p(341)(26),Cin=>p(342)(26),clock=>clock,reset=>reset,s=>p(357)(26),cout=>p(358)(27));
FA_ff_14191:FAff port map(x=>p(340)(27),y=>p(341)(27),Cin=>p(342)(27),clock=>clock,reset=>reset,s=>p(357)(27),cout=>p(358)(28));
FA_ff_14192:FAff port map(x=>p(340)(28),y=>p(341)(28),Cin=>p(342)(28),clock=>clock,reset=>reset,s=>p(357)(28),cout=>p(358)(29));
FA_ff_14193:FAff port map(x=>p(340)(29),y=>p(341)(29),Cin=>p(342)(29),clock=>clock,reset=>reset,s=>p(357)(29),cout=>p(358)(30));
FA_ff_14194:FAff port map(x=>p(340)(30),y=>p(341)(30),Cin=>p(342)(30),clock=>clock,reset=>reset,s=>p(357)(30),cout=>p(358)(31));
FA_ff_14195:FAff port map(x=>p(340)(31),y=>p(341)(31),Cin=>p(342)(31),clock=>clock,reset=>reset,s=>p(357)(31),cout=>p(358)(32));
FA_ff_14196:FAff port map(x=>p(340)(32),y=>p(341)(32),Cin=>p(342)(32),clock=>clock,reset=>reset,s=>p(357)(32),cout=>p(358)(33));
FA_ff_14197:FAff port map(x=>p(340)(33),y=>p(341)(33),Cin=>p(342)(33),clock=>clock,reset=>reset,s=>p(357)(33),cout=>p(358)(34));
FA_ff_14198:FAff port map(x=>p(340)(34),y=>p(341)(34),Cin=>p(342)(34),clock=>clock,reset=>reset,s=>p(357)(34),cout=>p(358)(35));
FA_ff_14199:FAff port map(x=>p(340)(35),y=>p(341)(35),Cin=>p(342)(35),clock=>clock,reset=>reset,s=>p(357)(35),cout=>p(358)(36));
FA_ff_14200:FAff port map(x=>p(340)(36),y=>p(341)(36),Cin=>p(342)(36),clock=>clock,reset=>reset,s=>p(357)(36),cout=>p(358)(37));
FA_ff_14201:FAff port map(x=>p(340)(37),y=>p(341)(37),Cin=>p(342)(37),clock=>clock,reset=>reset,s=>p(357)(37),cout=>p(358)(38));
FA_ff_14202:FAff port map(x=>p(340)(38),y=>p(341)(38),Cin=>p(342)(38),clock=>clock,reset=>reset,s=>p(357)(38),cout=>p(358)(39));
FA_ff_14203:FAff port map(x=>p(340)(39),y=>p(341)(39),Cin=>p(342)(39),clock=>clock,reset=>reset,s=>p(357)(39),cout=>p(358)(40));
FA_ff_14204:FAff port map(x=>p(340)(40),y=>p(341)(40),Cin=>p(342)(40),clock=>clock,reset=>reset,s=>p(357)(40),cout=>p(358)(41));
FA_ff_14205:FAff port map(x=>p(340)(41),y=>p(341)(41),Cin=>p(342)(41),clock=>clock,reset=>reset,s=>p(357)(41),cout=>p(358)(42));
FA_ff_14206:FAff port map(x=>p(340)(42),y=>p(341)(42),Cin=>p(342)(42),clock=>clock,reset=>reset,s=>p(357)(42),cout=>p(358)(43));
FA_ff_14207:FAff port map(x=>p(340)(43),y=>p(341)(43),Cin=>p(342)(43),clock=>clock,reset=>reset,s=>p(357)(43),cout=>p(358)(44));
FA_ff_14208:FAff port map(x=>p(340)(44),y=>p(341)(44),Cin=>p(342)(44),clock=>clock,reset=>reset,s=>p(357)(44),cout=>p(358)(45));
FA_ff_14209:FAff port map(x=>p(340)(45),y=>p(341)(45),Cin=>p(342)(45),clock=>clock,reset=>reset,s=>p(357)(45),cout=>p(358)(46));
FA_ff_14210:FAff port map(x=>p(340)(46),y=>p(341)(46),Cin=>p(342)(46),clock=>clock,reset=>reset,s=>p(357)(46),cout=>p(358)(47));
FA_ff_14211:FAff port map(x=>p(340)(47),y=>p(341)(47),Cin=>p(342)(47),clock=>clock,reset=>reset,s=>p(357)(47),cout=>p(358)(48));
FA_ff_14212:FAff port map(x=>p(340)(48),y=>p(341)(48),Cin=>p(342)(48),clock=>clock,reset=>reset,s=>p(357)(48),cout=>p(358)(49));
FA_ff_14213:FAff port map(x=>p(340)(49),y=>p(341)(49),Cin=>p(342)(49),clock=>clock,reset=>reset,s=>p(357)(49),cout=>p(358)(50));
FA_ff_14214:FAff port map(x=>p(340)(50),y=>p(341)(50),Cin=>p(342)(50),clock=>clock,reset=>reset,s=>p(357)(50),cout=>p(358)(51));
FA_ff_14215:FAff port map(x=>p(340)(51),y=>p(341)(51),Cin=>p(342)(51),clock=>clock,reset=>reset,s=>p(357)(51),cout=>p(358)(52));
FA_ff_14216:FAff port map(x=>p(340)(52),y=>p(341)(52),Cin=>p(342)(52),clock=>clock,reset=>reset,s=>p(357)(52),cout=>p(358)(53));
FA_ff_14217:FAff port map(x=>p(340)(53),y=>p(341)(53),Cin=>p(342)(53),clock=>clock,reset=>reset,s=>p(357)(53),cout=>p(358)(54));
FA_ff_14218:FAff port map(x=>p(340)(54),y=>p(341)(54),Cin=>p(342)(54),clock=>clock,reset=>reset,s=>p(357)(54),cout=>p(358)(55));
FA_ff_14219:FAff port map(x=>p(340)(55),y=>p(341)(55),Cin=>p(342)(55),clock=>clock,reset=>reset,s=>p(357)(55),cout=>p(358)(56));
FA_ff_14220:FAff port map(x=>p(340)(56),y=>p(341)(56),Cin=>p(342)(56),clock=>clock,reset=>reset,s=>p(357)(56),cout=>p(358)(57));
FA_ff_14221:FAff port map(x=>p(340)(57),y=>p(341)(57),Cin=>p(342)(57),clock=>clock,reset=>reset,s=>p(357)(57),cout=>p(358)(58));
FA_ff_14222:FAff port map(x=>p(340)(58),y=>p(341)(58),Cin=>p(342)(58),clock=>clock,reset=>reset,s=>p(357)(58),cout=>p(358)(59));
FA_ff_14223:FAff port map(x=>p(340)(59),y=>p(341)(59),Cin=>p(342)(59),clock=>clock,reset=>reset,s=>p(357)(59),cout=>p(358)(60));
FA_ff_14224:FAff port map(x=>p(340)(60),y=>p(341)(60),Cin=>p(342)(60),clock=>clock,reset=>reset,s=>p(357)(60),cout=>p(358)(61));
FA_ff_14225:FAff port map(x=>p(340)(61),y=>p(341)(61),Cin=>p(342)(61),clock=>clock,reset=>reset,s=>p(357)(61),cout=>p(358)(62));
FA_ff_14226:FAff port map(x=>p(340)(62),y=>p(341)(62),Cin=>p(342)(62),clock=>clock,reset=>reset,s=>p(357)(62),cout=>p(358)(63));
FA_ff_14227:FAff port map(x=>p(340)(63),y=>p(341)(63),Cin=>p(342)(63),clock=>clock,reset=>reset,s=>p(357)(63),cout=>p(358)(64));
FA_ff_14228:FAff port map(x=>p(340)(64),y=>p(341)(64),Cin=>p(342)(64),clock=>clock,reset=>reset,s=>p(357)(64),cout=>p(358)(65));
FA_ff_14229:FAff port map(x=>p(340)(65),y=>p(341)(65),Cin=>p(342)(65),clock=>clock,reset=>reset,s=>p(357)(65),cout=>p(358)(66));
FA_ff_14230:FAff port map(x=>p(340)(66),y=>p(341)(66),Cin=>p(342)(66),clock=>clock,reset=>reset,s=>p(357)(66),cout=>p(358)(67));
FA_ff_14231:FAff port map(x=>p(340)(67),y=>p(341)(67),Cin=>p(342)(67),clock=>clock,reset=>reset,s=>p(357)(67),cout=>p(358)(68));
FA_ff_14232:FAff port map(x=>p(340)(68),y=>p(341)(68),Cin=>p(342)(68),clock=>clock,reset=>reset,s=>p(357)(68),cout=>p(358)(69));
FA_ff_14233:FAff port map(x=>p(340)(69),y=>p(341)(69),Cin=>p(342)(69),clock=>clock,reset=>reset,s=>p(357)(69),cout=>p(358)(70));
FA_ff_14234:FAff port map(x=>p(340)(70),y=>p(341)(70),Cin=>p(342)(70),clock=>clock,reset=>reset,s=>p(357)(70),cout=>p(358)(71));
FA_ff_14235:FAff port map(x=>p(340)(71),y=>p(341)(71),Cin=>p(342)(71),clock=>clock,reset=>reset,s=>p(357)(71),cout=>p(358)(72));
FA_ff_14236:FAff port map(x=>p(340)(72),y=>p(341)(72),Cin=>p(342)(72),clock=>clock,reset=>reset,s=>p(357)(72),cout=>p(358)(73));
FA_ff_14237:FAff port map(x=>p(340)(73),y=>p(341)(73),Cin=>p(342)(73),clock=>clock,reset=>reset,s=>p(357)(73),cout=>p(358)(74));
FA_ff_14238:FAff port map(x=>p(340)(74),y=>p(341)(74),Cin=>p(342)(74),clock=>clock,reset=>reset,s=>p(357)(74),cout=>p(358)(75));
FA_ff_14239:FAff port map(x=>p(340)(75),y=>p(341)(75),Cin=>p(342)(75),clock=>clock,reset=>reset,s=>p(357)(75),cout=>p(358)(76));
FA_ff_14240:FAff port map(x=>p(340)(76),y=>p(341)(76),Cin=>p(342)(76),clock=>clock,reset=>reset,s=>p(357)(76),cout=>p(358)(77));
FA_ff_14241:FAff port map(x=>p(340)(77),y=>p(341)(77),Cin=>p(342)(77),clock=>clock,reset=>reset,s=>p(357)(77),cout=>p(358)(78));
FA_ff_14242:FAff port map(x=>p(340)(78),y=>p(341)(78),Cin=>p(342)(78),clock=>clock,reset=>reset,s=>p(357)(78),cout=>p(358)(79));
FA_ff_14243:FAff port map(x=>p(340)(79),y=>p(341)(79),Cin=>p(342)(79),clock=>clock,reset=>reset,s=>p(357)(79),cout=>p(358)(80));
FA_ff_14244:FAff port map(x=>p(340)(80),y=>p(341)(80),Cin=>p(342)(80),clock=>clock,reset=>reset,s=>p(357)(80),cout=>p(358)(81));
FA_ff_14245:FAff port map(x=>p(340)(81),y=>p(341)(81),Cin=>p(342)(81),clock=>clock,reset=>reset,s=>p(357)(81),cout=>p(358)(82));
FA_ff_14246:FAff port map(x=>p(340)(82),y=>p(341)(82),Cin=>p(342)(82),clock=>clock,reset=>reset,s=>p(357)(82),cout=>p(358)(83));
FA_ff_14247:FAff port map(x=>p(340)(83),y=>p(341)(83),Cin=>p(342)(83),clock=>clock,reset=>reset,s=>p(357)(83),cout=>p(358)(84));
FA_ff_14248:FAff port map(x=>p(340)(84),y=>p(341)(84),Cin=>p(342)(84),clock=>clock,reset=>reset,s=>p(357)(84),cout=>p(358)(85));
FA_ff_14249:FAff port map(x=>p(340)(85),y=>p(341)(85),Cin=>p(342)(85),clock=>clock,reset=>reset,s=>p(357)(85),cout=>p(358)(86));
FA_ff_14250:FAff port map(x=>p(340)(86),y=>p(341)(86),Cin=>p(342)(86),clock=>clock,reset=>reset,s=>p(357)(86),cout=>p(358)(87));
FA_ff_14251:FAff port map(x=>p(340)(87),y=>p(341)(87),Cin=>p(342)(87),clock=>clock,reset=>reset,s=>p(357)(87),cout=>p(358)(88));
FA_ff_14252:FAff port map(x=>p(340)(88),y=>p(341)(88),Cin=>p(342)(88),clock=>clock,reset=>reset,s=>p(357)(88),cout=>p(358)(89));
FA_ff_14253:FAff port map(x=>p(340)(89),y=>p(341)(89),Cin=>p(342)(89),clock=>clock,reset=>reset,s=>p(357)(89),cout=>p(358)(90));
FA_ff_14254:FAff port map(x=>p(340)(90),y=>p(341)(90),Cin=>p(342)(90),clock=>clock,reset=>reset,s=>p(357)(90),cout=>p(358)(91));
FA_ff_14255:FAff port map(x=>p(340)(91),y=>p(341)(91),Cin=>p(342)(91),clock=>clock,reset=>reset,s=>p(357)(91),cout=>p(358)(92));
FA_ff_14256:FAff port map(x=>p(340)(92),y=>p(341)(92),Cin=>p(342)(92),clock=>clock,reset=>reset,s=>p(357)(92),cout=>p(358)(93));
FA_ff_14257:FAff port map(x=>p(340)(93),y=>p(341)(93),Cin=>p(342)(93),clock=>clock,reset=>reset,s=>p(357)(93),cout=>p(358)(94));
FA_ff_14258:FAff port map(x=>p(340)(94),y=>p(341)(94),Cin=>p(342)(94),clock=>clock,reset=>reset,s=>p(357)(94),cout=>p(358)(95));
FA_ff_14259:FAff port map(x=>p(340)(95),y=>p(341)(95),Cin=>p(342)(95),clock=>clock,reset=>reset,s=>p(357)(95),cout=>p(358)(96));
FA_ff_14260:FAff port map(x=>p(340)(96),y=>p(341)(96),Cin=>p(342)(96),clock=>clock,reset=>reset,s=>p(357)(96),cout=>p(358)(97));
FA_ff_14261:FAff port map(x=>p(340)(97),y=>p(341)(97),Cin=>p(342)(97),clock=>clock,reset=>reset,s=>p(357)(97),cout=>p(358)(98));
FA_ff_14262:FAff port map(x=>p(340)(98),y=>p(341)(98),Cin=>p(342)(98),clock=>clock,reset=>reset,s=>p(357)(98),cout=>p(358)(99));
FA_ff_14263:FAff port map(x=>p(340)(99),y=>p(341)(99),Cin=>p(342)(99),clock=>clock,reset=>reset,s=>p(357)(99),cout=>p(358)(100));
FA_ff_14264:FAff port map(x=>p(340)(100),y=>p(341)(100),Cin=>p(342)(100),clock=>clock,reset=>reset,s=>p(357)(100),cout=>p(358)(101));
FA_ff_14265:FAff port map(x=>p(340)(101),y=>p(341)(101),Cin=>p(342)(101),clock=>clock,reset=>reset,s=>p(357)(101),cout=>p(358)(102));
FA_ff_14266:FAff port map(x=>p(340)(102),y=>p(341)(102),Cin=>p(342)(102),clock=>clock,reset=>reset,s=>p(357)(102),cout=>p(358)(103));
FA_ff_14267:FAff port map(x=>p(340)(103),y=>p(341)(103),Cin=>p(342)(103),clock=>clock,reset=>reset,s=>p(357)(103),cout=>p(358)(104));
FA_ff_14268:FAff port map(x=>p(340)(104),y=>p(341)(104),Cin=>p(342)(104),clock=>clock,reset=>reset,s=>p(357)(104),cout=>p(358)(105));
FA_ff_14269:FAff port map(x=>p(340)(105),y=>p(341)(105),Cin=>p(342)(105),clock=>clock,reset=>reset,s=>p(357)(105),cout=>p(358)(106));
FA_ff_14270:FAff port map(x=>p(340)(106),y=>p(341)(106),Cin=>p(342)(106),clock=>clock,reset=>reset,s=>p(357)(106),cout=>p(358)(107));
FA_ff_14271:FAff port map(x=>p(340)(107),y=>p(341)(107),Cin=>p(342)(107),clock=>clock,reset=>reset,s=>p(357)(107),cout=>p(358)(108));
FA_ff_14272:FAff port map(x=>p(340)(108),y=>p(341)(108),Cin=>p(342)(108),clock=>clock,reset=>reset,s=>p(357)(108),cout=>p(358)(109));
FA_ff_14273:FAff port map(x=>p(340)(109),y=>p(341)(109),Cin=>p(342)(109),clock=>clock,reset=>reset,s=>p(357)(109),cout=>p(358)(110));
FA_ff_14274:FAff port map(x=>p(340)(110),y=>p(341)(110),Cin=>p(342)(110),clock=>clock,reset=>reset,s=>p(357)(110),cout=>p(358)(111));
FA_ff_14275:FAff port map(x=>p(340)(111),y=>p(341)(111),Cin=>p(342)(111),clock=>clock,reset=>reset,s=>p(357)(111),cout=>p(358)(112));
FA_ff_14276:FAff port map(x=>p(340)(112),y=>p(341)(112),Cin=>p(342)(112),clock=>clock,reset=>reset,s=>p(357)(112),cout=>p(358)(113));
FA_ff_14277:FAff port map(x=>p(340)(113),y=>p(341)(113),Cin=>p(342)(113),clock=>clock,reset=>reset,s=>p(357)(113),cout=>p(358)(114));
FA_ff_14278:FAff port map(x=>p(340)(114),y=>p(341)(114),Cin=>p(342)(114),clock=>clock,reset=>reset,s=>p(357)(114),cout=>p(358)(115));
FA_ff_14279:FAff port map(x=>p(340)(115),y=>p(341)(115),Cin=>p(342)(115),clock=>clock,reset=>reset,s=>p(357)(115),cout=>p(358)(116));
FA_ff_14280:FAff port map(x=>p(340)(116),y=>p(341)(116),Cin=>p(342)(116),clock=>clock,reset=>reset,s=>p(357)(116),cout=>p(358)(117));
FA_ff_14281:FAff port map(x=>p(340)(117),y=>p(341)(117),Cin=>p(342)(117),clock=>clock,reset=>reset,s=>p(357)(117),cout=>p(358)(118));
FA_ff_14282:FAff port map(x=>p(340)(118),y=>p(341)(118),Cin=>p(342)(118),clock=>clock,reset=>reset,s=>p(357)(118),cout=>p(358)(119));
FA_ff_14283:FAff port map(x=>p(340)(119),y=>p(341)(119),Cin=>p(342)(119),clock=>clock,reset=>reset,s=>p(357)(119),cout=>p(358)(120));
FA_ff_14284:FAff port map(x=>p(340)(120),y=>p(341)(120),Cin=>p(342)(120),clock=>clock,reset=>reset,s=>p(357)(120),cout=>p(358)(121));
FA_ff_14285:FAff port map(x=>p(340)(121),y=>p(341)(121),Cin=>p(342)(121),clock=>clock,reset=>reset,s=>p(357)(121),cout=>p(358)(122));
FA_ff_14286:FAff port map(x=>p(340)(122),y=>p(341)(122),Cin=>p(342)(122),clock=>clock,reset=>reset,s=>p(357)(122),cout=>p(358)(123));
FA_ff_14287:FAff port map(x=>p(340)(123),y=>p(341)(123),Cin=>p(342)(123),clock=>clock,reset=>reset,s=>p(357)(123),cout=>p(358)(124));
FA_ff_14288:FAff port map(x=>p(340)(124),y=>p(341)(124),Cin=>p(342)(124),clock=>clock,reset=>reset,s=>p(357)(124),cout=>p(358)(125));
FA_ff_14289:FAff port map(x=>p(340)(125),y=>p(341)(125),Cin=>p(342)(125),clock=>clock,reset=>reset,s=>p(357)(125),cout=>p(358)(126));
FA_ff_14290:FAff port map(x=>p(340)(126),y=>p(341)(126),Cin=>p(342)(126),clock=>clock,reset=>reset,s=>p(357)(126),cout=>p(358)(127));
FA_ff_14291:FAff port map(x=>p(340)(127),y=>p(341)(127),Cin=>p(342)(127),clock=>clock,reset=>reset,s=>p(357)(127),cout=>p(358)(128));
FA_ff_14292:FAff port map(x=>p(340)(128),y=>p(341)(128),Cin=>p(342)(128),clock=>clock,reset=>reset,s=>p(357)(128),cout=>p(358)(129));
FA_ff_14293:FAff port map(x=>p(340)(129),y=>p(341)(129),Cin=>p(342)(129),clock=>clock,reset=>reset,s=>p(357)(129),cout=>p(358)(130));
FA_ff_14294:FAff port map(x=>p(340)(130),y=>p(341)(130),Cin=>p(342)(130),clock=>clock,reset=>reset,s=>p(357)(130),cout=>p(358)(131));
p(357)(131)<=p(340)(131);
HA_ff_92:HAff port map(x=>p(343)(0),y=>p(345)(0),clock=>clock,reset=>reset,s=>p(359)(0),c=>p(360)(1));
HA_ff_93:HAff port map(x=>p(343)(1),y=>p(345)(1),clock=>clock,reset=>reset,s=>p(359)(1),c=>p(360)(2));
FA_ff_14295:FAff port map(x=>p(343)(2),y=>p(344)(2),Cin=>p(345)(2),clock=>clock,reset=>reset,s=>p(359)(2),cout=>p(360)(3));
FA_ff_14296:FAff port map(x=>p(343)(3),y=>p(344)(3),Cin=>p(345)(3),clock=>clock,reset=>reset,s=>p(359)(3),cout=>p(360)(4));
FA_ff_14297:FAff port map(x=>p(343)(4),y=>p(344)(4),Cin=>p(345)(4),clock=>clock,reset=>reset,s=>p(359)(4),cout=>p(360)(5));
FA_ff_14298:FAff port map(x=>p(343)(5),y=>p(344)(5),Cin=>p(345)(5),clock=>clock,reset=>reset,s=>p(359)(5),cout=>p(360)(6));
FA_ff_14299:FAff port map(x=>p(343)(6),y=>p(344)(6),Cin=>p(345)(6),clock=>clock,reset=>reset,s=>p(359)(6),cout=>p(360)(7));
FA_ff_14300:FAff port map(x=>p(343)(7),y=>p(344)(7),Cin=>p(345)(7),clock=>clock,reset=>reset,s=>p(359)(7),cout=>p(360)(8));
FA_ff_14301:FAff port map(x=>p(343)(8),y=>p(344)(8),Cin=>p(345)(8),clock=>clock,reset=>reset,s=>p(359)(8),cout=>p(360)(9));
FA_ff_14302:FAff port map(x=>p(343)(9),y=>p(344)(9),Cin=>p(345)(9),clock=>clock,reset=>reset,s=>p(359)(9),cout=>p(360)(10));
FA_ff_14303:FAff port map(x=>p(343)(10),y=>p(344)(10),Cin=>p(345)(10),clock=>clock,reset=>reset,s=>p(359)(10),cout=>p(360)(11));
FA_ff_14304:FAff port map(x=>p(343)(11),y=>p(344)(11),Cin=>p(345)(11),clock=>clock,reset=>reset,s=>p(359)(11),cout=>p(360)(12));
FA_ff_14305:FAff port map(x=>p(343)(12),y=>p(344)(12),Cin=>p(345)(12),clock=>clock,reset=>reset,s=>p(359)(12),cout=>p(360)(13));
FA_ff_14306:FAff port map(x=>p(343)(13),y=>p(344)(13),Cin=>p(345)(13),clock=>clock,reset=>reset,s=>p(359)(13),cout=>p(360)(14));
FA_ff_14307:FAff port map(x=>p(343)(14),y=>p(344)(14),Cin=>p(345)(14),clock=>clock,reset=>reset,s=>p(359)(14),cout=>p(360)(15));
FA_ff_14308:FAff port map(x=>p(343)(15),y=>p(344)(15),Cin=>p(345)(15),clock=>clock,reset=>reset,s=>p(359)(15),cout=>p(360)(16));
FA_ff_14309:FAff port map(x=>p(343)(16),y=>p(344)(16),Cin=>p(345)(16),clock=>clock,reset=>reset,s=>p(359)(16),cout=>p(360)(17));
FA_ff_14310:FAff port map(x=>p(343)(17),y=>p(344)(17),Cin=>p(345)(17),clock=>clock,reset=>reset,s=>p(359)(17),cout=>p(360)(18));
FA_ff_14311:FAff port map(x=>p(343)(18),y=>p(344)(18),Cin=>p(345)(18),clock=>clock,reset=>reset,s=>p(359)(18),cout=>p(360)(19));
FA_ff_14312:FAff port map(x=>p(343)(19),y=>p(344)(19),Cin=>p(345)(19),clock=>clock,reset=>reset,s=>p(359)(19),cout=>p(360)(20));
FA_ff_14313:FAff port map(x=>p(343)(20),y=>p(344)(20),Cin=>p(345)(20),clock=>clock,reset=>reset,s=>p(359)(20),cout=>p(360)(21));
FA_ff_14314:FAff port map(x=>p(343)(21),y=>p(344)(21),Cin=>p(345)(21),clock=>clock,reset=>reset,s=>p(359)(21),cout=>p(360)(22));
FA_ff_14315:FAff port map(x=>p(343)(22),y=>p(344)(22),Cin=>p(345)(22),clock=>clock,reset=>reset,s=>p(359)(22),cout=>p(360)(23));
FA_ff_14316:FAff port map(x=>p(343)(23),y=>p(344)(23),Cin=>p(345)(23),clock=>clock,reset=>reset,s=>p(359)(23),cout=>p(360)(24));
FA_ff_14317:FAff port map(x=>p(343)(24),y=>p(344)(24),Cin=>p(345)(24),clock=>clock,reset=>reset,s=>p(359)(24),cout=>p(360)(25));
FA_ff_14318:FAff port map(x=>p(343)(25),y=>p(344)(25),Cin=>p(345)(25),clock=>clock,reset=>reset,s=>p(359)(25),cout=>p(360)(26));
FA_ff_14319:FAff port map(x=>p(343)(26),y=>p(344)(26),Cin=>p(345)(26),clock=>clock,reset=>reset,s=>p(359)(26),cout=>p(360)(27));
FA_ff_14320:FAff port map(x=>p(343)(27),y=>p(344)(27),Cin=>p(345)(27),clock=>clock,reset=>reset,s=>p(359)(27),cout=>p(360)(28));
FA_ff_14321:FAff port map(x=>p(343)(28),y=>p(344)(28),Cin=>p(345)(28),clock=>clock,reset=>reset,s=>p(359)(28),cout=>p(360)(29));
FA_ff_14322:FAff port map(x=>p(343)(29),y=>p(344)(29),Cin=>p(345)(29),clock=>clock,reset=>reset,s=>p(359)(29),cout=>p(360)(30));
FA_ff_14323:FAff port map(x=>p(343)(30),y=>p(344)(30),Cin=>p(345)(30),clock=>clock,reset=>reset,s=>p(359)(30),cout=>p(360)(31));
FA_ff_14324:FAff port map(x=>p(343)(31),y=>p(344)(31),Cin=>p(345)(31),clock=>clock,reset=>reset,s=>p(359)(31),cout=>p(360)(32));
FA_ff_14325:FAff port map(x=>p(343)(32),y=>p(344)(32),Cin=>p(345)(32),clock=>clock,reset=>reset,s=>p(359)(32),cout=>p(360)(33));
FA_ff_14326:FAff port map(x=>p(343)(33),y=>p(344)(33),Cin=>p(345)(33),clock=>clock,reset=>reset,s=>p(359)(33),cout=>p(360)(34));
FA_ff_14327:FAff port map(x=>p(343)(34),y=>p(344)(34),Cin=>p(345)(34),clock=>clock,reset=>reset,s=>p(359)(34),cout=>p(360)(35));
FA_ff_14328:FAff port map(x=>p(343)(35),y=>p(344)(35),Cin=>p(345)(35),clock=>clock,reset=>reset,s=>p(359)(35),cout=>p(360)(36));
FA_ff_14329:FAff port map(x=>p(343)(36),y=>p(344)(36),Cin=>p(345)(36),clock=>clock,reset=>reset,s=>p(359)(36),cout=>p(360)(37));
FA_ff_14330:FAff port map(x=>p(343)(37),y=>p(344)(37),Cin=>p(345)(37),clock=>clock,reset=>reset,s=>p(359)(37),cout=>p(360)(38));
FA_ff_14331:FAff port map(x=>p(343)(38),y=>p(344)(38),Cin=>p(345)(38),clock=>clock,reset=>reset,s=>p(359)(38),cout=>p(360)(39));
FA_ff_14332:FAff port map(x=>p(343)(39),y=>p(344)(39),Cin=>p(345)(39),clock=>clock,reset=>reset,s=>p(359)(39),cout=>p(360)(40));
FA_ff_14333:FAff port map(x=>p(343)(40),y=>p(344)(40),Cin=>p(345)(40),clock=>clock,reset=>reset,s=>p(359)(40),cout=>p(360)(41));
FA_ff_14334:FAff port map(x=>p(343)(41),y=>p(344)(41),Cin=>p(345)(41),clock=>clock,reset=>reset,s=>p(359)(41),cout=>p(360)(42));
FA_ff_14335:FAff port map(x=>p(343)(42),y=>p(344)(42),Cin=>p(345)(42),clock=>clock,reset=>reset,s=>p(359)(42),cout=>p(360)(43));
FA_ff_14336:FAff port map(x=>p(343)(43),y=>p(344)(43),Cin=>p(345)(43),clock=>clock,reset=>reset,s=>p(359)(43),cout=>p(360)(44));
FA_ff_14337:FAff port map(x=>p(343)(44),y=>p(344)(44),Cin=>p(345)(44),clock=>clock,reset=>reset,s=>p(359)(44),cout=>p(360)(45));
FA_ff_14338:FAff port map(x=>p(343)(45),y=>p(344)(45),Cin=>p(345)(45),clock=>clock,reset=>reset,s=>p(359)(45),cout=>p(360)(46));
FA_ff_14339:FAff port map(x=>p(343)(46),y=>p(344)(46),Cin=>p(345)(46),clock=>clock,reset=>reset,s=>p(359)(46),cout=>p(360)(47));
FA_ff_14340:FAff port map(x=>p(343)(47),y=>p(344)(47),Cin=>p(345)(47),clock=>clock,reset=>reset,s=>p(359)(47),cout=>p(360)(48));
FA_ff_14341:FAff port map(x=>p(343)(48),y=>p(344)(48),Cin=>p(345)(48),clock=>clock,reset=>reset,s=>p(359)(48),cout=>p(360)(49));
FA_ff_14342:FAff port map(x=>p(343)(49),y=>p(344)(49),Cin=>p(345)(49),clock=>clock,reset=>reset,s=>p(359)(49),cout=>p(360)(50));
FA_ff_14343:FAff port map(x=>p(343)(50),y=>p(344)(50),Cin=>p(345)(50),clock=>clock,reset=>reset,s=>p(359)(50),cout=>p(360)(51));
FA_ff_14344:FAff port map(x=>p(343)(51),y=>p(344)(51),Cin=>p(345)(51),clock=>clock,reset=>reset,s=>p(359)(51),cout=>p(360)(52));
FA_ff_14345:FAff port map(x=>p(343)(52),y=>p(344)(52),Cin=>p(345)(52),clock=>clock,reset=>reset,s=>p(359)(52),cout=>p(360)(53));
FA_ff_14346:FAff port map(x=>p(343)(53),y=>p(344)(53),Cin=>p(345)(53),clock=>clock,reset=>reset,s=>p(359)(53),cout=>p(360)(54));
FA_ff_14347:FAff port map(x=>p(343)(54),y=>p(344)(54),Cin=>p(345)(54),clock=>clock,reset=>reset,s=>p(359)(54),cout=>p(360)(55));
FA_ff_14348:FAff port map(x=>p(343)(55),y=>p(344)(55),Cin=>p(345)(55),clock=>clock,reset=>reset,s=>p(359)(55),cout=>p(360)(56));
FA_ff_14349:FAff port map(x=>p(343)(56),y=>p(344)(56),Cin=>p(345)(56),clock=>clock,reset=>reset,s=>p(359)(56),cout=>p(360)(57));
FA_ff_14350:FAff port map(x=>p(343)(57),y=>p(344)(57),Cin=>p(345)(57),clock=>clock,reset=>reset,s=>p(359)(57),cout=>p(360)(58));
FA_ff_14351:FAff port map(x=>p(343)(58),y=>p(344)(58),Cin=>p(345)(58),clock=>clock,reset=>reset,s=>p(359)(58),cout=>p(360)(59));
FA_ff_14352:FAff port map(x=>p(343)(59),y=>p(344)(59),Cin=>p(345)(59),clock=>clock,reset=>reset,s=>p(359)(59),cout=>p(360)(60));
FA_ff_14353:FAff port map(x=>p(343)(60),y=>p(344)(60),Cin=>p(345)(60),clock=>clock,reset=>reset,s=>p(359)(60),cout=>p(360)(61));
FA_ff_14354:FAff port map(x=>p(343)(61),y=>p(344)(61),Cin=>p(345)(61),clock=>clock,reset=>reset,s=>p(359)(61),cout=>p(360)(62));
FA_ff_14355:FAff port map(x=>p(343)(62),y=>p(344)(62),Cin=>p(345)(62),clock=>clock,reset=>reset,s=>p(359)(62),cout=>p(360)(63));
FA_ff_14356:FAff port map(x=>p(343)(63),y=>p(344)(63),Cin=>p(345)(63),clock=>clock,reset=>reset,s=>p(359)(63),cout=>p(360)(64));
FA_ff_14357:FAff port map(x=>p(343)(64),y=>p(344)(64),Cin=>p(345)(64),clock=>clock,reset=>reset,s=>p(359)(64),cout=>p(360)(65));
FA_ff_14358:FAff port map(x=>p(343)(65),y=>p(344)(65),Cin=>p(345)(65),clock=>clock,reset=>reset,s=>p(359)(65),cout=>p(360)(66));
FA_ff_14359:FAff port map(x=>p(343)(66),y=>p(344)(66),Cin=>p(345)(66),clock=>clock,reset=>reset,s=>p(359)(66),cout=>p(360)(67));
FA_ff_14360:FAff port map(x=>p(343)(67),y=>p(344)(67),Cin=>p(345)(67),clock=>clock,reset=>reset,s=>p(359)(67),cout=>p(360)(68));
FA_ff_14361:FAff port map(x=>p(343)(68),y=>p(344)(68),Cin=>p(345)(68),clock=>clock,reset=>reset,s=>p(359)(68),cout=>p(360)(69));
FA_ff_14362:FAff port map(x=>p(343)(69),y=>p(344)(69),Cin=>p(345)(69),clock=>clock,reset=>reset,s=>p(359)(69),cout=>p(360)(70));
FA_ff_14363:FAff port map(x=>p(343)(70),y=>p(344)(70),Cin=>p(345)(70),clock=>clock,reset=>reset,s=>p(359)(70),cout=>p(360)(71));
FA_ff_14364:FAff port map(x=>p(343)(71),y=>p(344)(71),Cin=>p(345)(71),clock=>clock,reset=>reset,s=>p(359)(71),cout=>p(360)(72));
FA_ff_14365:FAff port map(x=>p(343)(72),y=>p(344)(72),Cin=>p(345)(72),clock=>clock,reset=>reset,s=>p(359)(72),cout=>p(360)(73));
FA_ff_14366:FAff port map(x=>p(343)(73),y=>p(344)(73),Cin=>p(345)(73),clock=>clock,reset=>reset,s=>p(359)(73),cout=>p(360)(74));
FA_ff_14367:FAff port map(x=>p(343)(74),y=>p(344)(74),Cin=>p(345)(74),clock=>clock,reset=>reset,s=>p(359)(74),cout=>p(360)(75));
FA_ff_14368:FAff port map(x=>p(343)(75),y=>p(344)(75),Cin=>p(345)(75),clock=>clock,reset=>reset,s=>p(359)(75),cout=>p(360)(76));
FA_ff_14369:FAff port map(x=>p(343)(76),y=>p(344)(76),Cin=>p(345)(76),clock=>clock,reset=>reset,s=>p(359)(76),cout=>p(360)(77));
FA_ff_14370:FAff port map(x=>p(343)(77),y=>p(344)(77),Cin=>p(345)(77),clock=>clock,reset=>reset,s=>p(359)(77),cout=>p(360)(78));
FA_ff_14371:FAff port map(x=>p(343)(78),y=>p(344)(78),Cin=>p(345)(78),clock=>clock,reset=>reset,s=>p(359)(78),cout=>p(360)(79));
FA_ff_14372:FAff port map(x=>p(343)(79),y=>p(344)(79),Cin=>p(345)(79),clock=>clock,reset=>reset,s=>p(359)(79),cout=>p(360)(80));
FA_ff_14373:FAff port map(x=>p(343)(80),y=>p(344)(80),Cin=>p(345)(80),clock=>clock,reset=>reset,s=>p(359)(80),cout=>p(360)(81));
FA_ff_14374:FAff port map(x=>p(343)(81),y=>p(344)(81),Cin=>p(345)(81),clock=>clock,reset=>reset,s=>p(359)(81),cout=>p(360)(82));
FA_ff_14375:FAff port map(x=>p(343)(82),y=>p(344)(82),Cin=>p(345)(82),clock=>clock,reset=>reset,s=>p(359)(82),cout=>p(360)(83));
FA_ff_14376:FAff port map(x=>p(343)(83),y=>p(344)(83),Cin=>p(345)(83),clock=>clock,reset=>reset,s=>p(359)(83),cout=>p(360)(84));
FA_ff_14377:FAff port map(x=>p(343)(84),y=>p(344)(84),Cin=>p(345)(84),clock=>clock,reset=>reset,s=>p(359)(84),cout=>p(360)(85));
FA_ff_14378:FAff port map(x=>p(343)(85),y=>p(344)(85),Cin=>p(345)(85),clock=>clock,reset=>reset,s=>p(359)(85),cout=>p(360)(86));
FA_ff_14379:FAff port map(x=>p(343)(86),y=>p(344)(86),Cin=>p(345)(86),clock=>clock,reset=>reset,s=>p(359)(86),cout=>p(360)(87));
FA_ff_14380:FAff port map(x=>p(343)(87),y=>p(344)(87),Cin=>p(345)(87),clock=>clock,reset=>reset,s=>p(359)(87),cout=>p(360)(88));
FA_ff_14381:FAff port map(x=>p(343)(88),y=>p(344)(88),Cin=>p(345)(88),clock=>clock,reset=>reset,s=>p(359)(88),cout=>p(360)(89));
FA_ff_14382:FAff port map(x=>p(343)(89),y=>p(344)(89),Cin=>p(345)(89),clock=>clock,reset=>reset,s=>p(359)(89),cout=>p(360)(90));
FA_ff_14383:FAff port map(x=>p(343)(90),y=>p(344)(90),Cin=>p(345)(90),clock=>clock,reset=>reset,s=>p(359)(90),cout=>p(360)(91));
FA_ff_14384:FAff port map(x=>p(343)(91),y=>p(344)(91),Cin=>p(345)(91),clock=>clock,reset=>reset,s=>p(359)(91),cout=>p(360)(92));
FA_ff_14385:FAff port map(x=>p(343)(92),y=>p(344)(92),Cin=>p(345)(92),clock=>clock,reset=>reset,s=>p(359)(92),cout=>p(360)(93));
FA_ff_14386:FAff port map(x=>p(343)(93),y=>p(344)(93),Cin=>p(345)(93),clock=>clock,reset=>reset,s=>p(359)(93),cout=>p(360)(94));
FA_ff_14387:FAff port map(x=>p(343)(94),y=>p(344)(94),Cin=>p(345)(94),clock=>clock,reset=>reset,s=>p(359)(94),cout=>p(360)(95));
FA_ff_14388:FAff port map(x=>p(343)(95),y=>p(344)(95),Cin=>p(345)(95),clock=>clock,reset=>reset,s=>p(359)(95),cout=>p(360)(96));
FA_ff_14389:FAff port map(x=>p(343)(96),y=>p(344)(96),Cin=>p(345)(96),clock=>clock,reset=>reset,s=>p(359)(96),cout=>p(360)(97));
FA_ff_14390:FAff port map(x=>p(343)(97),y=>p(344)(97),Cin=>p(345)(97),clock=>clock,reset=>reset,s=>p(359)(97),cout=>p(360)(98));
FA_ff_14391:FAff port map(x=>p(343)(98),y=>p(344)(98),Cin=>p(345)(98),clock=>clock,reset=>reset,s=>p(359)(98),cout=>p(360)(99));
FA_ff_14392:FAff port map(x=>p(343)(99),y=>p(344)(99),Cin=>p(345)(99),clock=>clock,reset=>reset,s=>p(359)(99),cout=>p(360)(100));
FA_ff_14393:FAff port map(x=>p(343)(100),y=>p(344)(100),Cin=>p(345)(100),clock=>clock,reset=>reset,s=>p(359)(100),cout=>p(360)(101));
FA_ff_14394:FAff port map(x=>p(343)(101),y=>p(344)(101),Cin=>p(345)(101),clock=>clock,reset=>reset,s=>p(359)(101),cout=>p(360)(102));
FA_ff_14395:FAff port map(x=>p(343)(102),y=>p(344)(102),Cin=>p(345)(102),clock=>clock,reset=>reset,s=>p(359)(102),cout=>p(360)(103));
FA_ff_14396:FAff port map(x=>p(343)(103),y=>p(344)(103),Cin=>p(345)(103),clock=>clock,reset=>reset,s=>p(359)(103),cout=>p(360)(104));
FA_ff_14397:FAff port map(x=>p(343)(104),y=>p(344)(104),Cin=>p(345)(104),clock=>clock,reset=>reset,s=>p(359)(104),cout=>p(360)(105));
FA_ff_14398:FAff port map(x=>p(343)(105),y=>p(344)(105),Cin=>p(345)(105),clock=>clock,reset=>reset,s=>p(359)(105),cout=>p(360)(106));
FA_ff_14399:FAff port map(x=>p(343)(106),y=>p(344)(106),Cin=>p(345)(106),clock=>clock,reset=>reset,s=>p(359)(106),cout=>p(360)(107));
FA_ff_14400:FAff port map(x=>p(343)(107),y=>p(344)(107),Cin=>p(345)(107),clock=>clock,reset=>reset,s=>p(359)(107),cout=>p(360)(108));
FA_ff_14401:FAff port map(x=>p(343)(108),y=>p(344)(108),Cin=>p(345)(108),clock=>clock,reset=>reset,s=>p(359)(108),cout=>p(360)(109));
FA_ff_14402:FAff port map(x=>p(343)(109),y=>p(344)(109),Cin=>p(345)(109),clock=>clock,reset=>reset,s=>p(359)(109),cout=>p(360)(110));
FA_ff_14403:FAff port map(x=>p(343)(110),y=>p(344)(110),Cin=>p(345)(110),clock=>clock,reset=>reset,s=>p(359)(110),cout=>p(360)(111));
FA_ff_14404:FAff port map(x=>p(343)(111),y=>p(344)(111),Cin=>p(345)(111),clock=>clock,reset=>reset,s=>p(359)(111),cout=>p(360)(112));
FA_ff_14405:FAff port map(x=>p(343)(112),y=>p(344)(112),Cin=>p(345)(112),clock=>clock,reset=>reset,s=>p(359)(112),cout=>p(360)(113));
FA_ff_14406:FAff port map(x=>p(343)(113),y=>p(344)(113),Cin=>p(345)(113),clock=>clock,reset=>reset,s=>p(359)(113),cout=>p(360)(114));
FA_ff_14407:FAff port map(x=>p(343)(114),y=>p(344)(114),Cin=>p(345)(114),clock=>clock,reset=>reset,s=>p(359)(114),cout=>p(360)(115));
FA_ff_14408:FAff port map(x=>p(343)(115),y=>p(344)(115),Cin=>p(345)(115),clock=>clock,reset=>reset,s=>p(359)(115),cout=>p(360)(116));
FA_ff_14409:FAff port map(x=>p(343)(116),y=>p(344)(116),Cin=>p(345)(116),clock=>clock,reset=>reset,s=>p(359)(116),cout=>p(360)(117));
FA_ff_14410:FAff port map(x=>p(343)(117),y=>p(344)(117),Cin=>p(345)(117),clock=>clock,reset=>reset,s=>p(359)(117),cout=>p(360)(118));
FA_ff_14411:FAff port map(x=>p(343)(118),y=>p(344)(118),Cin=>p(345)(118),clock=>clock,reset=>reset,s=>p(359)(118),cout=>p(360)(119));
FA_ff_14412:FAff port map(x=>p(343)(119),y=>p(344)(119),Cin=>p(345)(119),clock=>clock,reset=>reset,s=>p(359)(119),cout=>p(360)(120));
FA_ff_14413:FAff port map(x=>p(343)(120),y=>p(344)(120),Cin=>p(345)(120),clock=>clock,reset=>reset,s=>p(359)(120),cout=>p(360)(121));
FA_ff_14414:FAff port map(x=>p(343)(121),y=>p(344)(121),Cin=>p(345)(121),clock=>clock,reset=>reset,s=>p(359)(121),cout=>p(360)(122));
FA_ff_14415:FAff port map(x=>p(343)(122),y=>p(344)(122),Cin=>p(345)(122),clock=>clock,reset=>reset,s=>p(359)(122),cout=>p(360)(123));
FA_ff_14416:FAff port map(x=>p(343)(123),y=>p(344)(123),Cin=>p(345)(123),clock=>clock,reset=>reset,s=>p(359)(123),cout=>p(360)(124));
FA_ff_14417:FAff port map(x=>p(343)(124),y=>p(344)(124),Cin=>p(345)(124),clock=>clock,reset=>reset,s=>p(359)(124),cout=>p(360)(125));
FA_ff_14418:FAff port map(x=>p(343)(125),y=>p(344)(125),Cin=>p(345)(125),clock=>clock,reset=>reset,s=>p(359)(125),cout=>p(360)(126));
FA_ff_14419:FAff port map(x=>p(343)(126),y=>p(344)(126),Cin=>p(345)(126),clock=>clock,reset=>reset,s=>p(359)(126),cout=>p(360)(127));
FA_ff_14420:FAff port map(x=>p(343)(127),y=>p(344)(127),Cin=>p(345)(127),clock=>clock,reset=>reset,s=>p(359)(127),cout=>p(360)(128));
FA_ff_14421:FAff port map(x=>p(343)(128),y=>p(344)(128),Cin=>p(345)(128),clock=>clock,reset=>reset,s=>p(359)(128),cout=>p(360)(129));
FA_ff_14422:FAff port map(x=>p(343)(129),y=>p(344)(129),Cin=>p(345)(129),clock=>clock,reset=>reset,s=>p(359)(129),cout=>p(360)(130));
FA_ff_14423:FAff port map(x=>p(343)(130),y=>p(344)(130),Cin=>p(345)(130),clock=>clock,reset=>reset,s=>p(359)(130),cout=>p(360)(131));
p(359)(131)<=p(344)(131);
p(361)(0)<=p(347)(0);
HA_ff_94:HAff port map(x=>p(346)(1),y=>p(347)(1),clock=>clock,reset=>reset,s=>p(361)(1),c=>p(362)(2));
FA_ff_14424:FAff port map(x=>p(346)(2),y=>p(347)(2),Cin=>p(348)(2),clock=>clock,reset=>reset,s=>p(361)(2),cout=>p(362)(3));
FA_ff_14425:FAff port map(x=>p(346)(3),y=>p(347)(3),Cin=>p(348)(3),clock=>clock,reset=>reset,s=>p(361)(3),cout=>p(362)(4));
FA_ff_14426:FAff port map(x=>p(346)(4),y=>p(347)(4),Cin=>p(348)(4),clock=>clock,reset=>reset,s=>p(361)(4),cout=>p(362)(5));
FA_ff_14427:FAff port map(x=>p(346)(5),y=>p(347)(5),Cin=>p(348)(5),clock=>clock,reset=>reset,s=>p(361)(5),cout=>p(362)(6));
FA_ff_14428:FAff port map(x=>p(346)(6),y=>p(347)(6),Cin=>p(348)(6),clock=>clock,reset=>reset,s=>p(361)(6),cout=>p(362)(7));
FA_ff_14429:FAff port map(x=>p(346)(7),y=>p(347)(7),Cin=>p(348)(7),clock=>clock,reset=>reset,s=>p(361)(7),cout=>p(362)(8));
FA_ff_14430:FAff port map(x=>p(346)(8),y=>p(347)(8),Cin=>p(348)(8),clock=>clock,reset=>reset,s=>p(361)(8),cout=>p(362)(9));
FA_ff_14431:FAff port map(x=>p(346)(9),y=>p(347)(9),Cin=>p(348)(9),clock=>clock,reset=>reset,s=>p(361)(9),cout=>p(362)(10));
FA_ff_14432:FAff port map(x=>p(346)(10),y=>p(347)(10),Cin=>p(348)(10),clock=>clock,reset=>reset,s=>p(361)(10),cout=>p(362)(11));
FA_ff_14433:FAff port map(x=>p(346)(11),y=>p(347)(11),Cin=>p(348)(11),clock=>clock,reset=>reset,s=>p(361)(11),cout=>p(362)(12));
FA_ff_14434:FAff port map(x=>p(346)(12),y=>p(347)(12),Cin=>p(348)(12),clock=>clock,reset=>reset,s=>p(361)(12),cout=>p(362)(13));
FA_ff_14435:FAff port map(x=>p(346)(13),y=>p(347)(13),Cin=>p(348)(13),clock=>clock,reset=>reset,s=>p(361)(13),cout=>p(362)(14));
FA_ff_14436:FAff port map(x=>p(346)(14),y=>p(347)(14),Cin=>p(348)(14),clock=>clock,reset=>reset,s=>p(361)(14),cout=>p(362)(15));
FA_ff_14437:FAff port map(x=>p(346)(15),y=>p(347)(15),Cin=>p(348)(15),clock=>clock,reset=>reset,s=>p(361)(15),cout=>p(362)(16));
FA_ff_14438:FAff port map(x=>p(346)(16),y=>p(347)(16),Cin=>p(348)(16),clock=>clock,reset=>reset,s=>p(361)(16),cout=>p(362)(17));
FA_ff_14439:FAff port map(x=>p(346)(17),y=>p(347)(17),Cin=>p(348)(17),clock=>clock,reset=>reset,s=>p(361)(17),cout=>p(362)(18));
FA_ff_14440:FAff port map(x=>p(346)(18),y=>p(347)(18),Cin=>p(348)(18),clock=>clock,reset=>reset,s=>p(361)(18),cout=>p(362)(19));
FA_ff_14441:FAff port map(x=>p(346)(19),y=>p(347)(19),Cin=>p(348)(19),clock=>clock,reset=>reset,s=>p(361)(19),cout=>p(362)(20));
FA_ff_14442:FAff port map(x=>p(346)(20),y=>p(347)(20),Cin=>p(348)(20),clock=>clock,reset=>reset,s=>p(361)(20),cout=>p(362)(21));
FA_ff_14443:FAff port map(x=>p(346)(21),y=>p(347)(21),Cin=>p(348)(21),clock=>clock,reset=>reset,s=>p(361)(21),cout=>p(362)(22));
FA_ff_14444:FAff port map(x=>p(346)(22),y=>p(347)(22),Cin=>p(348)(22),clock=>clock,reset=>reset,s=>p(361)(22),cout=>p(362)(23));
FA_ff_14445:FAff port map(x=>p(346)(23),y=>p(347)(23),Cin=>p(348)(23),clock=>clock,reset=>reset,s=>p(361)(23),cout=>p(362)(24));
FA_ff_14446:FAff port map(x=>p(346)(24),y=>p(347)(24),Cin=>p(348)(24),clock=>clock,reset=>reset,s=>p(361)(24),cout=>p(362)(25));
FA_ff_14447:FAff port map(x=>p(346)(25),y=>p(347)(25),Cin=>p(348)(25),clock=>clock,reset=>reset,s=>p(361)(25),cout=>p(362)(26));
FA_ff_14448:FAff port map(x=>p(346)(26),y=>p(347)(26),Cin=>p(348)(26),clock=>clock,reset=>reset,s=>p(361)(26),cout=>p(362)(27));
FA_ff_14449:FAff port map(x=>p(346)(27),y=>p(347)(27),Cin=>p(348)(27),clock=>clock,reset=>reset,s=>p(361)(27),cout=>p(362)(28));
FA_ff_14450:FAff port map(x=>p(346)(28),y=>p(347)(28),Cin=>p(348)(28),clock=>clock,reset=>reset,s=>p(361)(28),cout=>p(362)(29));
FA_ff_14451:FAff port map(x=>p(346)(29),y=>p(347)(29),Cin=>p(348)(29),clock=>clock,reset=>reset,s=>p(361)(29),cout=>p(362)(30));
FA_ff_14452:FAff port map(x=>p(346)(30),y=>p(347)(30),Cin=>p(348)(30),clock=>clock,reset=>reset,s=>p(361)(30),cout=>p(362)(31));
FA_ff_14453:FAff port map(x=>p(346)(31),y=>p(347)(31),Cin=>p(348)(31),clock=>clock,reset=>reset,s=>p(361)(31),cout=>p(362)(32));
FA_ff_14454:FAff port map(x=>p(346)(32),y=>p(347)(32),Cin=>p(348)(32),clock=>clock,reset=>reset,s=>p(361)(32),cout=>p(362)(33));
FA_ff_14455:FAff port map(x=>p(346)(33),y=>p(347)(33),Cin=>p(348)(33),clock=>clock,reset=>reset,s=>p(361)(33),cout=>p(362)(34));
FA_ff_14456:FAff port map(x=>p(346)(34),y=>p(347)(34),Cin=>p(348)(34),clock=>clock,reset=>reset,s=>p(361)(34),cout=>p(362)(35));
FA_ff_14457:FAff port map(x=>p(346)(35),y=>p(347)(35),Cin=>p(348)(35),clock=>clock,reset=>reset,s=>p(361)(35),cout=>p(362)(36));
FA_ff_14458:FAff port map(x=>p(346)(36),y=>p(347)(36),Cin=>p(348)(36),clock=>clock,reset=>reset,s=>p(361)(36),cout=>p(362)(37));
FA_ff_14459:FAff port map(x=>p(346)(37),y=>p(347)(37),Cin=>p(348)(37),clock=>clock,reset=>reset,s=>p(361)(37),cout=>p(362)(38));
FA_ff_14460:FAff port map(x=>p(346)(38),y=>p(347)(38),Cin=>p(348)(38),clock=>clock,reset=>reset,s=>p(361)(38),cout=>p(362)(39));
FA_ff_14461:FAff port map(x=>p(346)(39),y=>p(347)(39),Cin=>p(348)(39),clock=>clock,reset=>reset,s=>p(361)(39),cout=>p(362)(40));
FA_ff_14462:FAff port map(x=>p(346)(40),y=>p(347)(40),Cin=>p(348)(40),clock=>clock,reset=>reset,s=>p(361)(40),cout=>p(362)(41));
FA_ff_14463:FAff port map(x=>p(346)(41),y=>p(347)(41),Cin=>p(348)(41),clock=>clock,reset=>reset,s=>p(361)(41),cout=>p(362)(42));
FA_ff_14464:FAff port map(x=>p(346)(42),y=>p(347)(42),Cin=>p(348)(42),clock=>clock,reset=>reset,s=>p(361)(42),cout=>p(362)(43));
FA_ff_14465:FAff port map(x=>p(346)(43),y=>p(347)(43),Cin=>p(348)(43),clock=>clock,reset=>reset,s=>p(361)(43),cout=>p(362)(44));
FA_ff_14466:FAff port map(x=>p(346)(44),y=>p(347)(44),Cin=>p(348)(44),clock=>clock,reset=>reset,s=>p(361)(44),cout=>p(362)(45));
FA_ff_14467:FAff port map(x=>p(346)(45),y=>p(347)(45),Cin=>p(348)(45),clock=>clock,reset=>reset,s=>p(361)(45),cout=>p(362)(46));
FA_ff_14468:FAff port map(x=>p(346)(46),y=>p(347)(46),Cin=>p(348)(46),clock=>clock,reset=>reset,s=>p(361)(46),cout=>p(362)(47));
FA_ff_14469:FAff port map(x=>p(346)(47),y=>p(347)(47),Cin=>p(348)(47),clock=>clock,reset=>reset,s=>p(361)(47),cout=>p(362)(48));
FA_ff_14470:FAff port map(x=>p(346)(48),y=>p(347)(48),Cin=>p(348)(48),clock=>clock,reset=>reset,s=>p(361)(48),cout=>p(362)(49));
FA_ff_14471:FAff port map(x=>p(346)(49),y=>p(347)(49),Cin=>p(348)(49),clock=>clock,reset=>reset,s=>p(361)(49),cout=>p(362)(50));
FA_ff_14472:FAff port map(x=>p(346)(50),y=>p(347)(50),Cin=>p(348)(50),clock=>clock,reset=>reset,s=>p(361)(50),cout=>p(362)(51));
FA_ff_14473:FAff port map(x=>p(346)(51),y=>p(347)(51),Cin=>p(348)(51),clock=>clock,reset=>reset,s=>p(361)(51),cout=>p(362)(52));
FA_ff_14474:FAff port map(x=>p(346)(52),y=>p(347)(52),Cin=>p(348)(52),clock=>clock,reset=>reset,s=>p(361)(52),cout=>p(362)(53));
FA_ff_14475:FAff port map(x=>p(346)(53),y=>p(347)(53),Cin=>p(348)(53),clock=>clock,reset=>reset,s=>p(361)(53),cout=>p(362)(54));
FA_ff_14476:FAff port map(x=>p(346)(54),y=>p(347)(54),Cin=>p(348)(54),clock=>clock,reset=>reset,s=>p(361)(54),cout=>p(362)(55));
FA_ff_14477:FAff port map(x=>p(346)(55),y=>p(347)(55),Cin=>p(348)(55),clock=>clock,reset=>reset,s=>p(361)(55),cout=>p(362)(56));
FA_ff_14478:FAff port map(x=>p(346)(56),y=>p(347)(56),Cin=>p(348)(56),clock=>clock,reset=>reset,s=>p(361)(56),cout=>p(362)(57));
FA_ff_14479:FAff port map(x=>p(346)(57),y=>p(347)(57),Cin=>p(348)(57),clock=>clock,reset=>reset,s=>p(361)(57),cout=>p(362)(58));
FA_ff_14480:FAff port map(x=>p(346)(58),y=>p(347)(58),Cin=>p(348)(58),clock=>clock,reset=>reset,s=>p(361)(58),cout=>p(362)(59));
FA_ff_14481:FAff port map(x=>p(346)(59),y=>p(347)(59),Cin=>p(348)(59),clock=>clock,reset=>reset,s=>p(361)(59),cout=>p(362)(60));
FA_ff_14482:FAff port map(x=>p(346)(60),y=>p(347)(60),Cin=>p(348)(60),clock=>clock,reset=>reset,s=>p(361)(60),cout=>p(362)(61));
FA_ff_14483:FAff port map(x=>p(346)(61),y=>p(347)(61),Cin=>p(348)(61),clock=>clock,reset=>reset,s=>p(361)(61),cout=>p(362)(62));
FA_ff_14484:FAff port map(x=>p(346)(62),y=>p(347)(62),Cin=>p(348)(62),clock=>clock,reset=>reset,s=>p(361)(62),cout=>p(362)(63));
FA_ff_14485:FAff port map(x=>p(346)(63),y=>p(347)(63),Cin=>p(348)(63),clock=>clock,reset=>reset,s=>p(361)(63),cout=>p(362)(64));
FA_ff_14486:FAff port map(x=>p(346)(64),y=>p(347)(64),Cin=>p(348)(64),clock=>clock,reset=>reset,s=>p(361)(64),cout=>p(362)(65));
FA_ff_14487:FAff port map(x=>p(346)(65),y=>p(347)(65),Cin=>p(348)(65),clock=>clock,reset=>reset,s=>p(361)(65),cout=>p(362)(66));
FA_ff_14488:FAff port map(x=>p(346)(66),y=>p(347)(66),Cin=>p(348)(66),clock=>clock,reset=>reset,s=>p(361)(66),cout=>p(362)(67));
FA_ff_14489:FAff port map(x=>p(346)(67),y=>p(347)(67),Cin=>p(348)(67),clock=>clock,reset=>reset,s=>p(361)(67),cout=>p(362)(68));
FA_ff_14490:FAff port map(x=>p(346)(68),y=>p(347)(68),Cin=>p(348)(68),clock=>clock,reset=>reset,s=>p(361)(68),cout=>p(362)(69));
FA_ff_14491:FAff port map(x=>p(346)(69),y=>p(347)(69),Cin=>p(348)(69),clock=>clock,reset=>reset,s=>p(361)(69),cout=>p(362)(70));
FA_ff_14492:FAff port map(x=>p(346)(70),y=>p(347)(70),Cin=>p(348)(70),clock=>clock,reset=>reset,s=>p(361)(70),cout=>p(362)(71));
FA_ff_14493:FAff port map(x=>p(346)(71),y=>p(347)(71),Cin=>p(348)(71),clock=>clock,reset=>reset,s=>p(361)(71),cout=>p(362)(72));
FA_ff_14494:FAff port map(x=>p(346)(72),y=>p(347)(72),Cin=>p(348)(72),clock=>clock,reset=>reset,s=>p(361)(72),cout=>p(362)(73));
FA_ff_14495:FAff port map(x=>p(346)(73),y=>p(347)(73),Cin=>p(348)(73),clock=>clock,reset=>reset,s=>p(361)(73),cout=>p(362)(74));
FA_ff_14496:FAff port map(x=>p(346)(74),y=>p(347)(74),Cin=>p(348)(74),clock=>clock,reset=>reset,s=>p(361)(74),cout=>p(362)(75));
FA_ff_14497:FAff port map(x=>p(346)(75),y=>p(347)(75),Cin=>p(348)(75),clock=>clock,reset=>reset,s=>p(361)(75),cout=>p(362)(76));
FA_ff_14498:FAff port map(x=>p(346)(76),y=>p(347)(76),Cin=>p(348)(76),clock=>clock,reset=>reset,s=>p(361)(76),cout=>p(362)(77));
FA_ff_14499:FAff port map(x=>p(346)(77),y=>p(347)(77),Cin=>p(348)(77),clock=>clock,reset=>reset,s=>p(361)(77),cout=>p(362)(78));
FA_ff_14500:FAff port map(x=>p(346)(78),y=>p(347)(78),Cin=>p(348)(78),clock=>clock,reset=>reset,s=>p(361)(78),cout=>p(362)(79));
FA_ff_14501:FAff port map(x=>p(346)(79),y=>p(347)(79),Cin=>p(348)(79),clock=>clock,reset=>reset,s=>p(361)(79),cout=>p(362)(80));
FA_ff_14502:FAff port map(x=>p(346)(80),y=>p(347)(80),Cin=>p(348)(80),clock=>clock,reset=>reset,s=>p(361)(80),cout=>p(362)(81));
FA_ff_14503:FAff port map(x=>p(346)(81),y=>p(347)(81),Cin=>p(348)(81),clock=>clock,reset=>reset,s=>p(361)(81),cout=>p(362)(82));
FA_ff_14504:FAff port map(x=>p(346)(82),y=>p(347)(82),Cin=>p(348)(82),clock=>clock,reset=>reset,s=>p(361)(82),cout=>p(362)(83));
FA_ff_14505:FAff port map(x=>p(346)(83),y=>p(347)(83),Cin=>p(348)(83),clock=>clock,reset=>reset,s=>p(361)(83),cout=>p(362)(84));
FA_ff_14506:FAff port map(x=>p(346)(84),y=>p(347)(84),Cin=>p(348)(84),clock=>clock,reset=>reset,s=>p(361)(84),cout=>p(362)(85));
FA_ff_14507:FAff port map(x=>p(346)(85),y=>p(347)(85),Cin=>p(348)(85),clock=>clock,reset=>reset,s=>p(361)(85),cout=>p(362)(86));
FA_ff_14508:FAff port map(x=>p(346)(86),y=>p(347)(86),Cin=>p(348)(86),clock=>clock,reset=>reset,s=>p(361)(86),cout=>p(362)(87));
FA_ff_14509:FAff port map(x=>p(346)(87),y=>p(347)(87),Cin=>p(348)(87),clock=>clock,reset=>reset,s=>p(361)(87),cout=>p(362)(88));
FA_ff_14510:FAff port map(x=>p(346)(88),y=>p(347)(88),Cin=>p(348)(88),clock=>clock,reset=>reset,s=>p(361)(88),cout=>p(362)(89));
FA_ff_14511:FAff port map(x=>p(346)(89),y=>p(347)(89),Cin=>p(348)(89),clock=>clock,reset=>reset,s=>p(361)(89),cout=>p(362)(90));
FA_ff_14512:FAff port map(x=>p(346)(90),y=>p(347)(90),Cin=>p(348)(90),clock=>clock,reset=>reset,s=>p(361)(90),cout=>p(362)(91));
FA_ff_14513:FAff port map(x=>p(346)(91),y=>p(347)(91),Cin=>p(348)(91),clock=>clock,reset=>reset,s=>p(361)(91),cout=>p(362)(92));
FA_ff_14514:FAff port map(x=>p(346)(92),y=>p(347)(92),Cin=>p(348)(92),clock=>clock,reset=>reset,s=>p(361)(92),cout=>p(362)(93));
FA_ff_14515:FAff port map(x=>p(346)(93),y=>p(347)(93),Cin=>p(348)(93),clock=>clock,reset=>reset,s=>p(361)(93),cout=>p(362)(94));
FA_ff_14516:FAff port map(x=>p(346)(94),y=>p(347)(94),Cin=>p(348)(94),clock=>clock,reset=>reset,s=>p(361)(94),cout=>p(362)(95));
FA_ff_14517:FAff port map(x=>p(346)(95),y=>p(347)(95),Cin=>p(348)(95),clock=>clock,reset=>reset,s=>p(361)(95),cout=>p(362)(96));
FA_ff_14518:FAff port map(x=>p(346)(96),y=>p(347)(96),Cin=>p(348)(96),clock=>clock,reset=>reset,s=>p(361)(96),cout=>p(362)(97));
FA_ff_14519:FAff port map(x=>p(346)(97),y=>p(347)(97),Cin=>p(348)(97),clock=>clock,reset=>reset,s=>p(361)(97),cout=>p(362)(98));
FA_ff_14520:FAff port map(x=>p(346)(98),y=>p(347)(98),Cin=>p(348)(98),clock=>clock,reset=>reset,s=>p(361)(98),cout=>p(362)(99));
FA_ff_14521:FAff port map(x=>p(346)(99),y=>p(347)(99),Cin=>p(348)(99),clock=>clock,reset=>reset,s=>p(361)(99),cout=>p(362)(100));
FA_ff_14522:FAff port map(x=>p(346)(100),y=>p(347)(100),Cin=>p(348)(100),clock=>clock,reset=>reset,s=>p(361)(100),cout=>p(362)(101));
FA_ff_14523:FAff port map(x=>p(346)(101),y=>p(347)(101),Cin=>p(348)(101),clock=>clock,reset=>reset,s=>p(361)(101),cout=>p(362)(102));
FA_ff_14524:FAff port map(x=>p(346)(102),y=>p(347)(102),Cin=>p(348)(102),clock=>clock,reset=>reset,s=>p(361)(102),cout=>p(362)(103));
FA_ff_14525:FAff port map(x=>p(346)(103),y=>p(347)(103),Cin=>p(348)(103),clock=>clock,reset=>reset,s=>p(361)(103),cout=>p(362)(104));
FA_ff_14526:FAff port map(x=>p(346)(104),y=>p(347)(104),Cin=>p(348)(104),clock=>clock,reset=>reset,s=>p(361)(104),cout=>p(362)(105));
FA_ff_14527:FAff port map(x=>p(346)(105),y=>p(347)(105),Cin=>p(348)(105),clock=>clock,reset=>reset,s=>p(361)(105),cout=>p(362)(106));
FA_ff_14528:FAff port map(x=>p(346)(106),y=>p(347)(106),Cin=>p(348)(106),clock=>clock,reset=>reset,s=>p(361)(106),cout=>p(362)(107));
FA_ff_14529:FAff port map(x=>p(346)(107),y=>p(347)(107),Cin=>p(348)(107),clock=>clock,reset=>reset,s=>p(361)(107),cout=>p(362)(108));
FA_ff_14530:FAff port map(x=>p(346)(108),y=>p(347)(108),Cin=>p(348)(108),clock=>clock,reset=>reset,s=>p(361)(108),cout=>p(362)(109));
FA_ff_14531:FAff port map(x=>p(346)(109),y=>p(347)(109),Cin=>p(348)(109),clock=>clock,reset=>reset,s=>p(361)(109),cout=>p(362)(110));
FA_ff_14532:FAff port map(x=>p(346)(110),y=>p(347)(110),Cin=>p(348)(110),clock=>clock,reset=>reset,s=>p(361)(110),cout=>p(362)(111));
FA_ff_14533:FAff port map(x=>p(346)(111),y=>p(347)(111),Cin=>p(348)(111),clock=>clock,reset=>reset,s=>p(361)(111),cout=>p(362)(112));
FA_ff_14534:FAff port map(x=>p(346)(112),y=>p(347)(112),Cin=>p(348)(112),clock=>clock,reset=>reset,s=>p(361)(112),cout=>p(362)(113));
FA_ff_14535:FAff port map(x=>p(346)(113),y=>p(347)(113),Cin=>p(348)(113),clock=>clock,reset=>reset,s=>p(361)(113),cout=>p(362)(114));
FA_ff_14536:FAff port map(x=>p(346)(114),y=>p(347)(114),Cin=>p(348)(114),clock=>clock,reset=>reset,s=>p(361)(114),cout=>p(362)(115));
FA_ff_14537:FAff port map(x=>p(346)(115),y=>p(347)(115),Cin=>p(348)(115),clock=>clock,reset=>reset,s=>p(361)(115),cout=>p(362)(116));
FA_ff_14538:FAff port map(x=>p(346)(116),y=>p(347)(116),Cin=>p(348)(116),clock=>clock,reset=>reset,s=>p(361)(116),cout=>p(362)(117));
FA_ff_14539:FAff port map(x=>p(346)(117),y=>p(347)(117),Cin=>p(348)(117),clock=>clock,reset=>reset,s=>p(361)(117),cout=>p(362)(118));
FA_ff_14540:FAff port map(x=>p(346)(118),y=>p(347)(118),Cin=>p(348)(118),clock=>clock,reset=>reset,s=>p(361)(118),cout=>p(362)(119));
FA_ff_14541:FAff port map(x=>p(346)(119),y=>p(347)(119),Cin=>p(348)(119),clock=>clock,reset=>reset,s=>p(361)(119),cout=>p(362)(120));
FA_ff_14542:FAff port map(x=>p(346)(120),y=>p(347)(120),Cin=>p(348)(120),clock=>clock,reset=>reset,s=>p(361)(120),cout=>p(362)(121));
FA_ff_14543:FAff port map(x=>p(346)(121),y=>p(347)(121),Cin=>p(348)(121),clock=>clock,reset=>reset,s=>p(361)(121),cout=>p(362)(122));
FA_ff_14544:FAff port map(x=>p(346)(122),y=>p(347)(122),Cin=>p(348)(122),clock=>clock,reset=>reset,s=>p(361)(122),cout=>p(362)(123));
FA_ff_14545:FAff port map(x=>p(346)(123),y=>p(347)(123),Cin=>p(348)(123),clock=>clock,reset=>reset,s=>p(361)(123),cout=>p(362)(124));
FA_ff_14546:FAff port map(x=>p(346)(124),y=>p(347)(124),Cin=>p(348)(124),clock=>clock,reset=>reset,s=>p(361)(124),cout=>p(362)(125));
FA_ff_14547:FAff port map(x=>p(346)(125),y=>p(347)(125),Cin=>p(348)(125),clock=>clock,reset=>reset,s=>p(361)(125),cout=>p(362)(126));
FA_ff_14548:FAff port map(x=>p(346)(126),y=>p(347)(126),Cin=>p(348)(126),clock=>clock,reset=>reset,s=>p(361)(126),cout=>p(362)(127));
FA_ff_14549:FAff port map(x=>p(346)(127),y=>p(347)(127),Cin=>p(348)(127),clock=>clock,reset=>reset,s=>p(361)(127),cout=>p(362)(128));
FA_ff_14550:FAff port map(x=>p(346)(128),y=>p(347)(128),Cin=>p(348)(128),clock=>clock,reset=>reset,s=>p(361)(128),cout=>p(362)(129));
FA_ff_14551:FAff port map(x=>p(346)(129),y=>p(347)(129),Cin=>p(348)(129),clock=>clock,reset=>reset,s=>p(361)(129),cout=>p(362)(130));
FA_ff_14552:FAff port map(x=>p(346)(130),y=>p(347)(130),Cin=>p(348)(130),clock=>clock,reset=>reset,s=>p(361)(130),cout=>p(362)(131));
p(361)(131)<=p(348)(131);
HA_ff_95:HAff port map(x=>p(349)(0),y=>p(351)(0),clock=>clock,reset=>reset,s=>p(363)(0),c=>p(364)(1));
FA_ff_14553:FAff port map(x=>p(349)(1),y=>p(350)(1),Cin=>p(351)(1),clock=>clock,reset=>reset,s=>p(363)(1),cout=>p(364)(2));
FA_ff_14554:FAff port map(x=>p(349)(2),y=>p(350)(2),Cin=>p(351)(2),clock=>clock,reset=>reset,s=>p(363)(2),cout=>p(364)(3));
FA_ff_14555:FAff port map(x=>p(349)(3),y=>p(350)(3),Cin=>p(351)(3),clock=>clock,reset=>reset,s=>p(363)(3),cout=>p(364)(4));
FA_ff_14556:FAff port map(x=>p(349)(4),y=>p(350)(4),Cin=>p(351)(4),clock=>clock,reset=>reset,s=>p(363)(4),cout=>p(364)(5));
FA_ff_14557:FAff port map(x=>p(349)(5),y=>p(350)(5),Cin=>p(351)(5),clock=>clock,reset=>reset,s=>p(363)(5),cout=>p(364)(6));
FA_ff_14558:FAff port map(x=>p(349)(6),y=>p(350)(6),Cin=>p(351)(6),clock=>clock,reset=>reset,s=>p(363)(6),cout=>p(364)(7));
FA_ff_14559:FAff port map(x=>p(349)(7),y=>p(350)(7),Cin=>p(351)(7),clock=>clock,reset=>reset,s=>p(363)(7),cout=>p(364)(8));
FA_ff_14560:FAff port map(x=>p(349)(8),y=>p(350)(8),Cin=>p(351)(8),clock=>clock,reset=>reset,s=>p(363)(8),cout=>p(364)(9));
FA_ff_14561:FAff port map(x=>p(349)(9),y=>p(350)(9),Cin=>p(351)(9),clock=>clock,reset=>reset,s=>p(363)(9),cout=>p(364)(10));
FA_ff_14562:FAff port map(x=>p(349)(10),y=>p(350)(10),Cin=>p(351)(10),clock=>clock,reset=>reset,s=>p(363)(10),cout=>p(364)(11));
FA_ff_14563:FAff port map(x=>p(349)(11),y=>p(350)(11),Cin=>p(351)(11),clock=>clock,reset=>reset,s=>p(363)(11),cout=>p(364)(12));
FA_ff_14564:FAff port map(x=>p(349)(12),y=>p(350)(12),Cin=>p(351)(12),clock=>clock,reset=>reset,s=>p(363)(12),cout=>p(364)(13));
FA_ff_14565:FAff port map(x=>p(349)(13),y=>p(350)(13),Cin=>p(351)(13),clock=>clock,reset=>reset,s=>p(363)(13),cout=>p(364)(14));
FA_ff_14566:FAff port map(x=>p(349)(14),y=>p(350)(14),Cin=>p(351)(14),clock=>clock,reset=>reset,s=>p(363)(14),cout=>p(364)(15));
FA_ff_14567:FAff port map(x=>p(349)(15),y=>p(350)(15),Cin=>p(351)(15),clock=>clock,reset=>reset,s=>p(363)(15),cout=>p(364)(16));
FA_ff_14568:FAff port map(x=>p(349)(16),y=>p(350)(16),Cin=>p(351)(16),clock=>clock,reset=>reset,s=>p(363)(16),cout=>p(364)(17));
FA_ff_14569:FAff port map(x=>p(349)(17),y=>p(350)(17),Cin=>p(351)(17),clock=>clock,reset=>reset,s=>p(363)(17),cout=>p(364)(18));
FA_ff_14570:FAff port map(x=>p(349)(18),y=>p(350)(18),Cin=>p(351)(18),clock=>clock,reset=>reset,s=>p(363)(18),cout=>p(364)(19));
FA_ff_14571:FAff port map(x=>p(349)(19),y=>p(350)(19),Cin=>p(351)(19),clock=>clock,reset=>reset,s=>p(363)(19),cout=>p(364)(20));
FA_ff_14572:FAff port map(x=>p(349)(20),y=>p(350)(20),Cin=>p(351)(20),clock=>clock,reset=>reset,s=>p(363)(20),cout=>p(364)(21));
FA_ff_14573:FAff port map(x=>p(349)(21),y=>p(350)(21),Cin=>p(351)(21),clock=>clock,reset=>reset,s=>p(363)(21),cout=>p(364)(22));
FA_ff_14574:FAff port map(x=>p(349)(22),y=>p(350)(22),Cin=>p(351)(22),clock=>clock,reset=>reset,s=>p(363)(22),cout=>p(364)(23));
FA_ff_14575:FAff port map(x=>p(349)(23),y=>p(350)(23),Cin=>p(351)(23),clock=>clock,reset=>reset,s=>p(363)(23),cout=>p(364)(24));
FA_ff_14576:FAff port map(x=>p(349)(24),y=>p(350)(24),Cin=>p(351)(24),clock=>clock,reset=>reset,s=>p(363)(24),cout=>p(364)(25));
FA_ff_14577:FAff port map(x=>p(349)(25),y=>p(350)(25),Cin=>p(351)(25),clock=>clock,reset=>reset,s=>p(363)(25),cout=>p(364)(26));
FA_ff_14578:FAff port map(x=>p(349)(26),y=>p(350)(26),Cin=>p(351)(26),clock=>clock,reset=>reset,s=>p(363)(26),cout=>p(364)(27));
FA_ff_14579:FAff port map(x=>p(349)(27),y=>p(350)(27),Cin=>p(351)(27),clock=>clock,reset=>reset,s=>p(363)(27),cout=>p(364)(28));
FA_ff_14580:FAff port map(x=>p(349)(28),y=>p(350)(28),Cin=>p(351)(28),clock=>clock,reset=>reset,s=>p(363)(28),cout=>p(364)(29));
FA_ff_14581:FAff port map(x=>p(349)(29),y=>p(350)(29),Cin=>p(351)(29),clock=>clock,reset=>reset,s=>p(363)(29),cout=>p(364)(30));
FA_ff_14582:FAff port map(x=>p(349)(30),y=>p(350)(30),Cin=>p(351)(30),clock=>clock,reset=>reset,s=>p(363)(30),cout=>p(364)(31));
FA_ff_14583:FAff port map(x=>p(349)(31),y=>p(350)(31),Cin=>p(351)(31),clock=>clock,reset=>reset,s=>p(363)(31),cout=>p(364)(32));
FA_ff_14584:FAff port map(x=>p(349)(32),y=>p(350)(32),Cin=>p(351)(32),clock=>clock,reset=>reset,s=>p(363)(32),cout=>p(364)(33));
FA_ff_14585:FAff port map(x=>p(349)(33),y=>p(350)(33),Cin=>p(351)(33),clock=>clock,reset=>reset,s=>p(363)(33),cout=>p(364)(34));
FA_ff_14586:FAff port map(x=>p(349)(34),y=>p(350)(34),Cin=>p(351)(34),clock=>clock,reset=>reset,s=>p(363)(34),cout=>p(364)(35));
FA_ff_14587:FAff port map(x=>p(349)(35),y=>p(350)(35),Cin=>p(351)(35),clock=>clock,reset=>reset,s=>p(363)(35),cout=>p(364)(36));
FA_ff_14588:FAff port map(x=>p(349)(36),y=>p(350)(36),Cin=>p(351)(36),clock=>clock,reset=>reset,s=>p(363)(36),cout=>p(364)(37));
FA_ff_14589:FAff port map(x=>p(349)(37),y=>p(350)(37),Cin=>p(351)(37),clock=>clock,reset=>reset,s=>p(363)(37),cout=>p(364)(38));
FA_ff_14590:FAff port map(x=>p(349)(38),y=>p(350)(38),Cin=>p(351)(38),clock=>clock,reset=>reset,s=>p(363)(38),cout=>p(364)(39));
FA_ff_14591:FAff port map(x=>p(349)(39),y=>p(350)(39),Cin=>p(351)(39),clock=>clock,reset=>reset,s=>p(363)(39),cout=>p(364)(40));
FA_ff_14592:FAff port map(x=>p(349)(40),y=>p(350)(40),Cin=>p(351)(40),clock=>clock,reset=>reset,s=>p(363)(40),cout=>p(364)(41));
FA_ff_14593:FAff port map(x=>p(349)(41),y=>p(350)(41),Cin=>p(351)(41),clock=>clock,reset=>reset,s=>p(363)(41),cout=>p(364)(42));
FA_ff_14594:FAff port map(x=>p(349)(42),y=>p(350)(42),Cin=>p(351)(42),clock=>clock,reset=>reset,s=>p(363)(42),cout=>p(364)(43));
FA_ff_14595:FAff port map(x=>p(349)(43),y=>p(350)(43),Cin=>p(351)(43),clock=>clock,reset=>reset,s=>p(363)(43),cout=>p(364)(44));
FA_ff_14596:FAff port map(x=>p(349)(44),y=>p(350)(44),Cin=>p(351)(44),clock=>clock,reset=>reset,s=>p(363)(44),cout=>p(364)(45));
FA_ff_14597:FAff port map(x=>p(349)(45),y=>p(350)(45),Cin=>p(351)(45),clock=>clock,reset=>reset,s=>p(363)(45),cout=>p(364)(46));
FA_ff_14598:FAff port map(x=>p(349)(46),y=>p(350)(46),Cin=>p(351)(46),clock=>clock,reset=>reset,s=>p(363)(46),cout=>p(364)(47));
FA_ff_14599:FAff port map(x=>p(349)(47),y=>p(350)(47),Cin=>p(351)(47),clock=>clock,reset=>reset,s=>p(363)(47),cout=>p(364)(48));
FA_ff_14600:FAff port map(x=>p(349)(48),y=>p(350)(48),Cin=>p(351)(48),clock=>clock,reset=>reset,s=>p(363)(48),cout=>p(364)(49));
FA_ff_14601:FAff port map(x=>p(349)(49),y=>p(350)(49),Cin=>p(351)(49),clock=>clock,reset=>reset,s=>p(363)(49),cout=>p(364)(50));
FA_ff_14602:FAff port map(x=>p(349)(50),y=>p(350)(50),Cin=>p(351)(50),clock=>clock,reset=>reset,s=>p(363)(50),cout=>p(364)(51));
FA_ff_14603:FAff port map(x=>p(349)(51),y=>p(350)(51),Cin=>p(351)(51),clock=>clock,reset=>reset,s=>p(363)(51),cout=>p(364)(52));
FA_ff_14604:FAff port map(x=>p(349)(52),y=>p(350)(52),Cin=>p(351)(52),clock=>clock,reset=>reset,s=>p(363)(52),cout=>p(364)(53));
FA_ff_14605:FAff port map(x=>p(349)(53),y=>p(350)(53),Cin=>p(351)(53),clock=>clock,reset=>reset,s=>p(363)(53),cout=>p(364)(54));
FA_ff_14606:FAff port map(x=>p(349)(54),y=>p(350)(54),Cin=>p(351)(54),clock=>clock,reset=>reset,s=>p(363)(54),cout=>p(364)(55));
FA_ff_14607:FAff port map(x=>p(349)(55),y=>p(350)(55),Cin=>p(351)(55),clock=>clock,reset=>reset,s=>p(363)(55),cout=>p(364)(56));
FA_ff_14608:FAff port map(x=>p(349)(56),y=>p(350)(56),Cin=>p(351)(56),clock=>clock,reset=>reset,s=>p(363)(56),cout=>p(364)(57));
FA_ff_14609:FAff port map(x=>p(349)(57),y=>p(350)(57),Cin=>p(351)(57),clock=>clock,reset=>reset,s=>p(363)(57),cout=>p(364)(58));
FA_ff_14610:FAff port map(x=>p(349)(58),y=>p(350)(58),Cin=>p(351)(58),clock=>clock,reset=>reset,s=>p(363)(58),cout=>p(364)(59));
FA_ff_14611:FAff port map(x=>p(349)(59),y=>p(350)(59),Cin=>p(351)(59),clock=>clock,reset=>reset,s=>p(363)(59),cout=>p(364)(60));
FA_ff_14612:FAff port map(x=>p(349)(60),y=>p(350)(60),Cin=>p(351)(60),clock=>clock,reset=>reset,s=>p(363)(60),cout=>p(364)(61));
FA_ff_14613:FAff port map(x=>p(349)(61),y=>p(350)(61),Cin=>p(351)(61),clock=>clock,reset=>reset,s=>p(363)(61),cout=>p(364)(62));
FA_ff_14614:FAff port map(x=>p(349)(62),y=>p(350)(62),Cin=>p(351)(62),clock=>clock,reset=>reset,s=>p(363)(62),cout=>p(364)(63));
FA_ff_14615:FAff port map(x=>p(349)(63),y=>p(350)(63),Cin=>p(351)(63),clock=>clock,reset=>reset,s=>p(363)(63),cout=>p(364)(64));
FA_ff_14616:FAff port map(x=>p(349)(64),y=>p(350)(64),Cin=>p(351)(64),clock=>clock,reset=>reset,s=>p(363)(64),cout=>p(364)(65));
FA_ff_14617:FAff port map(x=>p(349)(65),y=>p(350)(65),Cin=>p(351)(65),clock=>clock,reset=>reset,s=>p(363)(65),cout=>p(364)(66));
FA_ff_14618:FAff port map(x=>p(349)(66),y=>p(350)(66),Cin=>p(351)(66),clock=>clock,reset=>reset,s=>p(363)(66),cout=>p(364)(67));
FA_ff_14619:FAff port map(x=>p(349)(67),y=>p(350)(67),Cin=>p(351)(67),clock=>clock,reset=>reset,s=>p(363)(67),cout=>p(364)(68));
FA_ff_14620:FAff port map(x=>p(349)(68),y=>p(350)(68),Cin=>p(351)(68),clock=>clock,reset=>reset,s=>p(363)(68),cout=>p(364)(69));
FA_ff_14621:FAff port map(x=>p(349)(69),y=>p(350)(69),Cin=>p(351)(69),clock=>clock,reset=>reset,s=>p(363)(69),cout=>p(364)(70));
FA_ff_14622:FAff port map(x=>p(349)(70),y=>p(350)(70),Cin=>p(351)(70),clock=>clock,reset=>reset,s=>p(363)(70),cout=>p(364)(71));
FA_ff_14623:FAff port map(x=>p(349)(71),y=>p(350)(71),Cin=>p(351)(71),clock=>clock,reset=>reset,s=>p(363)(71),cout=>p(364)(72));
FA_ff_14624:FAff port map(x=>p(349)(72),y=>p(350)(72),Cin=>p(351)(72),clock=>clock,reset=>reset,s=>p(363)(72),cout=>p(364)(73));
FA_ff_14625:FAff port map(x=>p(349)(73),y=>p(350)(73),Cin=>p(351)(73),clock=>clock,reset=>reset,s=>p(363)(73),cout=>p(364)(74));
FA_ff_14626:FAff port map(x=>p(349)(74),y=>p(350)(74),Cin=>p(351)(74),clock=>clock,reset=>reset,s=>p(363)(74),cout=>p(364)(75));
FA_ff_14627:FAff port map(x=>p(349)(75),y=>p(350)(75),Cin=>p(351)(75),clock=>clock,reset=>reset,s=>p(363)(75),cout=>p(364)(76));
FA_ff_14628:FAff port map(x=>p(349)(76),y=>p(350)(76),Cin=>p(351)(76),clock=>clock,reset=>reset,s=>p(363)(76),cout=>p(364)(77));
FA_ff_14629:FAff port map(x=>p(349)(77),y=>p(350)(77),Cin=>p(351)(77),clock=>clock,reset=>reset,s=>p(363)(77),cout=>p(364)(78));
FA_ff_14630:FAff port map(x=>p(349)(78),y=>p(350)(78),Cin=>p(351)(78),clock=>clock,reset=>reset,s=>p(363)(78),cout=>p(364)(79));
FA_ff_14631:FAff port map(x=>p(349)(79),y=>p(350)(79),Cin=>p(351)(79),clock=>clock,reset=>reset,s=>p(363)(79),cout=>p(364)(80));
FA_ff_14632:FAff port map(x=>p(349)(80),y=>p(350)(80),Cin=>p(351)(80),clock=>clock,reset=>reset,s=>p(363)(80),cout=>p(364)(81));
FA_ff_14633:FAff port map(x=>p(349)(81),y=>p(350)(81),Cin=>p(351)(81),clock=>clock,reset=>reset,s=>p(363)(81),cout=>p(364)(82));
FA_ff_14634:FAff port map(x=>p(349)(82),y=>p(350)(82),Cin=>p(351)(82),clock=>clock,reset=>reset,s=>p(363)(82),cout=>p(364)(83));
FA_ff_14635:FAff port map(x=>p(349)(83),y=>p(350)(83),Cin=>p(351)(83),clock=>clock,reset=>reset,s=>p(363)(83),cout=>p(364)(84));
FA_ff_14636:FAff port map(x=>p(349)(84),y=>p(350)(84),Cin=>p(351)(84),clock=>clock,reset=>reset,s=>p(363)(84),cout=>p(364)(85));
FA_ff_14637:FAff port map(x=>p(349)(85),y=>p(350)(85),Cin=>p(351)(85),clock=>clock,reset=>reset,s=>p(363)(85),cout=>p(364)(86));
FA_ff_14638:FAff port map(x=>p(349)(86),y=>p(350)(86),Cin=>p(351)(86),clock=>clock,reset=>reset,s=>p(363)(86),cout=>p(364)(87));
FA_ff_14639:FAff port map(x=>p(349)(87),y=>p(350)(87),Cin=>p(351)(87),clock=>clock,reset=>reset,s=>p(363)(87),cout=>p(364)(88));
FA_ff_14640:FAff port map(x=>p(349)(88),y=>p(350)(88),Cin=>p(351)(88),clock=>clock,reset=>reset,s=>p(363)(88),cout=>p(364)(89));
FA_ff_14641:FAff port map(x=>p(349)(89),y=>p(350)(89),Cin=>p(351)(89),clock=>clock,reset=>reset,s=>p(363)(89),cout=>p(364)(90));
FA_ff_14642:FAff port map(x=>p(349)(90),y=>p(350)(90),Cin=>p(351)(90),clock=>clock,reset=>reset,s=>p(363)(90),cout=>p(364)(91));
FA_ff_14643:FAff port map(x=>p(349)(91),y=>p(350)(91),Cin=>p(351)(91),clock=>clock,reset=>reset,s=>p(363)(91),cout=>p(364)(92));
FA_ff_14644:FAff port map(x=>p(349)(92),y=>p(350)(92),Cin=>p(351)(92),clock=>clock,reset=>reset,s=>p(363)(92),cout=>p(364)(93));
FA_ff_14645:FAff port map(x=>p(349)(93),y=>p(350)(93),Cin=>p(351)(93),clock=>clock,reset=>reset,s=>p(363)(93),cout=>p(364)(94));
FA_ff_14646:FAff port map(x=>p(349)(94),y=>p(350)(94),Cin=>p(351)(94),clock=>clock,reset=>reset,s=>p(363)(94),cout=>p(364)(95));
FA_ff_14647:FAff port map(x=>p(349)(95),y=>p(350)(95),Cin=>p(351)(95),clock=>clock,reset=>reset,s=>p(363)(95),cout=>p(364)(96));
FA_ff_14648:FAff port map(x=>p(349)(96),y=>p(350)(96),Cin=>p(351)(96),clock=>clock,reset=>reset,s=>p(363)(96),cout=>p(364)(97));
FA_ff_14649:FAff port map(x=>p(349)(97),y=>p(350)(97),Cin=>p(351)(97),clock=>clock,reset=>reset,s=>p(363)(97),cout=>p(364)(98));
FA_ff_14650:FAff port map(x=>p(349)(98),y=>p(350)(98),Cin=>p(351)(98),clock=>clock,reset=>reset,s=>p(363)(98),cout=>p(364)(99));
FA_ff_14651:FAff port map(x=>p(349)(99),y=>p(350)(99),Cin=>p(351)(99),clock=>clock,reset=>reset,s=>p(363)(99),cout=>p(364)(100));
FA_ff_14652:FAff port map(x=>p(349)(100),y=>p(350)(100),Cin=>p(351)(100),clock=>clock,reset=>reset,s=>p(363)(100),cout=>p(364)(101));
FA_ff_14653:FAff port map(x=>p(349)(101),y=>p(350)(101),Cin=>p(351)(101),clock=>clock,reset=>reset,s=>p(363)(101),cout=>p(364)(102));
FA_ff_14654:FAff port map(x=>p(349)(102),y=>p(350)(102),Cin=>p(351)(102),clock=>clock,reset=>reset,s=>p(363)(102),cout=>p(364)(103));
FA_ff_14655:FAff port map(x=>p(349)(103),y=>p(350)(103),Cin=>p(351)(103),clock=>clock,reset=>reset,s=>p(363)(103),cout=>p(364)(104));
FA_ff_14656:FAff port map(x=>p(349)(104),y=>p(350)(104),Cin=>p(351)(104),clock=>clock,reset=>reset,s=>p(363)(104),cout=>p(364)(105));
FA_ff_14657:FAff port map(x=>p(349)(105),y=>p(350)(105),Cin=>p(351)(105),clock=>clock,reset=>reset,s=>p(363)(105),cout=>p(364)(106));
FA_ff_14658:FAff port map(x=>p(349)(106),y=>p(350)(106),Cin=>p(351)(106),clock=>clock,reset=>reset,s=>p(363)(106),cout=>p(364)(107));
FA_ff_14659:FAff port map(x=>p(349)(107),y=>p(350)(107),Cin=>p(351)(107),clock=>clock,reset=>reset,s=>p(363)(107),cout=>p(364)(108));
FA_ff_14660:FAff port map(x=>p(349)(108),y=>p(350)(108),Cin=>p(351)(108),clock=>clock,reset=>reset,s=>p(363)(108),cout=>p(364)(109));
FA_ff_14661:FAff port map(x=>p(349)(109),y=>p(350)(109),Cin=>p(351)(109),clock=>clock,reset=>reset,s=>p(363)(109),cout=>p(364)(110));
FA_ff_14662:FAff port map(x=>p(349)(110),y=>p(350)(110),Cin=>p(351)(110),clock=>clock,reset=>reset,s=>p(363)(110),cout=>p(364)(111));
FA_ff_14663:FAff port map(x=>p(349)(111),y=>p(350)(111),Cin=>p(351)(111),clock=>clock,reset=>reset,s=>p(363)(111),cout=>p(364)(112));
FA_ff_14664:FAff port map(x=>p(349)(112),y=>p(350)(112),Cin=>p(351)(112),clock=>clock,reset=>reset,s=>p(363)(112),cout=>p(364)(113));
FA_ff_14665:FAff port map(x=>p(349)(113),y=>p(350)(113),Cin=>p(351)(113),clock=>clock,reset=>reset,s=>p(363)(113),cout=>p(364)(114));
FA_ff_14666:FAff port map(x=>p(349)(114),y=>p(350)(114),Cin=>p(351)(114),clock=>clock,reset=>reset,s=>p(363)(114),cout=>p(364)(115));
FA_ff_14667:FAff port map(x=>p(349)(115),y=>p(350)(115),Cin=>p(351)(115),clock=>clock,reset=>reset,s=>p(363)(115),cout=>p(364)(116));
FA_ff_14668:FAff port map(x=>p(349)(116),y=>p(350)(116),Cin=>p(351)(116),clock=>clock,reset=>reset,s=>p(363)(116),cout=>p(364)(117));
FA_ff_14669:FAff port map(x=>p(349)(117),y=>p(350)(117),Cin=>p(351)(117),clock=>clock,reset=>reset,s=>p(363)(117),cout=>p(364)(118));
FA_ff_14670:FAff port map(x=>p(349)(118),y=>p(350)(118),Cin=>p(351)(118),clock=>clock,reset=>reset,s=>p(363)(118),cout=>p(364)(119));
FA_ff_14671:FAff port map(x=>p(349)(119),y=>p(350)(119),Cin=>p(351)(119),clock=>clock,reset=>reset,s=>p(363)(119),cout=>p(364)(120));
FA_ff_14672:FAff port map(x=>p(349)(120),y=>p(350)(120),Cin=>p(351)(120),clock=>clock,reset=>reset,s=>p(363)(120),cout=>p(364)(121));
FA_ff_14673:FAff port map(x=>p(349)(121),y=>p(350)(121),Cin=>p(351)(121),clock=>clock,reset=>reset,s=>p(363)(121),cout=>p(364)(122));
FA_ff_14674:FAff port map(x=>p(349)(122),y=>p(350)(122),Cin=>p(351)(122),clock=>clock,reset=>reset,s=>p(363)(122),cout=>p(364)(123));
FA_ff_14675:FAff port map(x=>p(349)(123),y=>p(350)(123),Cin=>p(351)(123),clock=>clock,reset=>reset,s=>p(363)(123),cout=>p(364)(124));
FA_ff_14676:FAff port map(x=>p(349)(124),y=>p(350)(124),Cin=>p(351)(124),clock=>clock,reset=>reset,s=>p(363)(124),cout=>p(364)(125));
FA_ff_14677:FAff port map(x=>p(349)(125),y=>p(350)(125),Cin=>p(351)(125),clock=>clock,reset=>reset,s=>p(363)(125),cout=>p(364)(126));
FA_ff_14678:FAff port map(x=>p(349)(126),y=>p(350)(126),Cin=>p(351)(126),clock=>clock,reset=>reset,s=>p(363)(126),cout=>p(364)(127));
FA_ff_14679:FAff port map(x=>p(349)(127),y=>p(350)(127),Cin=>p(351)(127),clock=>clock,reset=>reset,s=>p(363)(127),cout=>p(364)(128));
FA_ff_14680:FAff port map(x=>p(349)(128),y=>p(350)(128),Cin=>p(351)(128),clock=>clock,reset=>reset,s=>p(363)(128),cout=>p(364)(129));
FA_ff_14681:FAff port map(x=>p(349)(129),y=>p(350)(129),Cin=>p(351)(129),clock=>clock,reset=>reset,s=>p(363)(129),cout=>p(364)(130));
FA_ff_14682:FAff port map(x=>p(349)(130),y=>p(350)(130),Cin=>p(351)(130),clock=>clock,reset=>reset,s=>p(363)(130),cout=>p(364)(131));
p(365)(0)<=p(353)(0);
HA_ff_96:HAff port map(x=>p(353)(1),y=>p(354)(1),clock=>clock,reset=>reset,s=>p(365)(1),c=>p(366)(2));
FA_ff_14683:FAff port map(x=>p(352)(2),y=>p(353)(2),Cin=>p(354)(2),clock=>clock,reset=>reset,s=>p(365)(2),cout=>p(366)(3));
FA_ff_14684:FAff port map(x=>p(352)(3),y=>p(353)(3),Cin=>p(354)(3),clock=>clock,reset=>reset,s=>p(365)(3),cout=>p(366)(4));
FA_ff_14685:FAff port map(x=>p(352)(4),y=>p(353)(4),Cin=>p(354)(4),clock=>clock,reset=>reset,s=>p(365)(4),cout=>p(366)(5));
FA_ff_14686:FAff port map(x=>p(352)(5),y=>p(353)(5),Cin=>p(354)(5),clock=>clock,reset=>reset,s=>p(365)(5),cout=>p(366)(6));
FA_ff_14687:FAff port map(x=>p(352)(6),y=>p(353)(6),Cin=>p(354)(6),clock=>clock,reset=>reset,s=>p(365)(6),cout=>p(366)(7));
FA_ff_14688:FAff port map(x=>p(352)(7),y=>p(353)(7),Cin=>p(354)(7),clock=>clock,reset=>reset,s=>p(365)(7),cout=>p(366)(8));
FA_ff_14689:FAff port map(x=>p(352)(8),y=>p(353)(8),Cin=>p(354)(8),clock=>clock,reset=>reset,s=>p(365)(8),cout=>p(366)(9));
FA_ff_14690:FAff port map(x=>p(352)(9),y=>p(353)(9),Cin=>p(354)(9),clock=>clock,reset=>reset,s=>p(365)(9),cout=>p(366)(10));
FA_ff_14691:FAff port map(x=>p(352)(10),y=>p(353)(10),Cin=>p(354)(10),clock=>clock,reset=>reset,s=>p(365)(10),cout=>p(366)(11));
FA_ff_14692:FAff port map(x=>p(352)(11),y=>p(353)(11),Cin=>p(354)(11),clock=>clock,reset=>reset,s=>p(365)(11),cout=>p(366)(12));
FA_ff_14693:FAff port map(x=>p(352)(12),y=>p(353)(12),Cin=>p(354)(12),clock=>clock,reset=>reset,s=>p(365)(12),cout=>p(366)(13));
FA_ff_14694:FAff port map(x=>p(352)(13),y=>p(353)(13),Cin=>p(354)(13),clock=>clock,reset=>reset,s=>p(365)(13),cout=>p(366)(14));
FA_ff_14695:FAff port map(x=>p(352)(14),y=>p(353)(14),Cin=>p(354)(14),clock=>clock,reset=>reset,s=>p(365)(14),cout=>p(366)(15));
FA_ff_14696:FAff port map(x=>p(352)(15),y=>p(353)(15),Cin=>p(354)(15),clock=>clock,reset=>reset,s=>p(365)(15),cout=>p(366)(16));
FA_ff_14697:FAff port map(x=>p(352)(16),y=>p(353)(16),Cin=>p(354)(16),clock=>clock,reset=>reset,s=>p(365)(16),cout=>p(366)(17));
FA_ff_14698:FAff port map(x=>p(352)(17),y=>p(353)(17),Cin=>p(354)(17),clock=>clock,reset=>reset,s=>p(365)(17),cout=>p(366)(18));
FA_ff_14699:FAff port map(x=>p(352)(18),y=>p(353)(18),Cin=>p(354)(18),clock=>clock,reset=>reset,s=>p(365)(18),cout=>p(366)(19));
FA_ff_14700:FAff port map(x=>p(352)(19),y=>p(353)(19),Cin=>p(354)(19),clock=>clock,reset=>reset,s=>p(365)(19),cout=>p(366)(20));
FA_ff_14701:FAff port map(x=>p(352)(20),y=>p(353)(20),Cin=>p(354)(20),clock=>clock,reset=>reset,s=>p(365)(20),cout=>p(366)(21));
FA_ff_14702:FAff port map(x=>p(352)(21),y=>p(353)(21),Cin=>p(354)(21),clock=>clock,reset=>reset,s=>p(365)(21),cout=>p(366)(22));
FA_ff_14703:FAff port map(x=>p(352)(22),y=>p(353)(22),Cin=>p(354)(22),clock=>clock,reset=>reset,s=>p(365)(22),cout=>p(366)(23));
FA_ff_14704:FAff port map(x=>p(352)(23),y=>p(353)(23),Cin=>p(354)(23),clock=>clock,reset=>reset,s=>p(365)(23),cout=>p(366)(24));
FA_ff_14705:FAff port map(x=>p(352)(24),y=>p(353)(24),Cin=>p(354)(24),clock=>clock,reset=>reset,s=>p(365)(24),cout=>p(366)(25));
FA_ff_14706:FAff port map(x=>p(352)(25),y=>p(353)(25),Cin=>p(354)(25),clock=>clock,reset=>reset,s=>p(365)(25),cout=>p(366)(26));
FA_ff_14707:FAff port map(x=>p(352)(26),y=>p(353)(26),Cin=>p(354)(26),clock=>clock,reset=>reset,s=>p(365)(26),cout=>p(366)(27));
FA_ff_14708:FAff port map(x=>p(352)(27),y=>p(353)(27),Cin=>p(354)(27),clock=>clock,reset=>reset,s=>p(365)(27),cout=>p(366)(28));
FA_ff_14709:FAff port map(x=>p(352)(28),y=>p(353)(28),Cin=>p(354)(28),clock=>clock,reset=>reset,s=>p(365)(28),cout=>p(366)(29));
FA_ff_14710:FAff port map(x=>p(352)(29),y=>p(353)(29),Cin=>p(354)(29),clock=>clock,reset=>reset,s=>p(365)(29),cout=>p(366)(30));
FA_ff_14711:FAff port map(x=>p(352)(30),y=>p(353)(30),Cin=>p(354)(30),clock=>clock,reset=>reset,s=>p(365)(30),cout=>p(366)(31));
FA_ff_14712:FAff port map(x=>p(352)(31),y=>p(353)(31),Cin=>p(354)(31),clock=>clock,reset=>reset,s=>p(365)(31),cout=>p(366)(32));
FA_ff_14713:FAff port map(x=>p(352)(32),y=>p(353)(32),Cin=>p(354)(32),clock=>clock,reset=>reset,s=>p(365)(32),cout=>p(366)(33));
FA_ff_14714:FAff port map(x=>p(352)(33),y=>p(353)(33),Cin=>p(354)(33),clock=>clock,reset=>reset,s=>p(365)(33),cout=>p(366)(34));
FA_ff_14715:FAff port map(x=>p(352)(34),y=>p(353)(34),Cin=>p(354)(34),clock=>clock,reset=>reset,s=>p(365)(34),cout=>p(366)(35));
FA_ff_14716:FAff port map(x=>p(352)(35),y=>p(353)(35),Cin=>p(354)(35),clock=>clock,reset=>reset,s=>p(365)(35),cout=>p(366)(36));
FA_ff_14717:FAff port map(x=>p(352)(36),y=>p(353)(36),Cin=>p(354)(36),clock=>clock,reset=>reset,s=>p(365)(36),cout=>p(366)(37));
FA_ff_14718:FAff port map(x=>p(352)(37),y=>p(353)(37),Cin=>p(354)(37),clock=>clock,reset=>reset,s=>p(365)(37),cout=>p(366)(38));
FA_ff_14719:FAff port map(x=>p(352)(38),y=>p(353)(38),Cin=>p(354)(38),clock=>clock,reset=>reset,s=>p(365)(38),cout=>p(366)(39));
FA_ff_14720:FAff port map(x=>p(352)(39),y=>p(353)(39),Cin=>p(354)(39),clock=>clock,reset=>reset,s=>p(365)(39),cout=>p(366)(40));
FA_ff_14721:FAff port map(x=>p(352)(40),y=>p(353)(40),Cin=>p(354)(40),clock=>clock,reset=>reset,s=>p(365)(40),cout=>p(366)(41));
FA_ff_14722:FAff port map(x=>p(352)(41),y=>p(353)(41),Cin=>p(354)(41),clock=>clock,reset=>reset,s=>p(365)(41),cout=>p(366)(42));
FA_ff_14723:FAff port map(x=>p(352)(42),y=>p(353)(42),Cin=>p(354)(42),clock=>clock,reset=>reset,s=>p(365)(42),cout=>p(366)(43));
FA_ff_14724:FAff port map(x=>p(352)(43),y=>p(353)(43),Cin=>p(354)(43),clock=>clock,reset=>reset,s=>p(365)(43),cout=>p(366)(44));
FA_ff_14725:FAff port map(x=>p(352)(44),y=>p(353)(44),Cin=>p(354)(44),clock=>clock,reset=>reset,s=>p(365)(44),cout=>p(366)(45));
FA_ff_14726:FAff port map(x=>p(352)(45),y=>p(353)(45),Cin=>p(354)(45),clock=>clock,reset=>reset,s=>p(365)(45),cout=>p(366)(46));
FA_ff_14727:FAff port map(x=>p(352)(46),y=>p(353)(46),Cin=>p(354)(46),clock=>clock,reset=>reset,s=>p(365)(46),cout=>p(366)(47));
FA_ff_14728:FAff port map(x=>p(352)(47),y=>p(353)(47),Cin=>p(354)(47),clock=>clock,reset=>reset,s=>p(365)(47),cout=>p(366)(48));
FA_ff_14729:FAff port map(x=>p(352)(48),y=>p(353)(48),Cin=>p(354)(48),clock=>clock,reset=>reset,s=>p(365)(48),cout=>p(366)(49));
FA_ff_14730:FAff port map(x=>p(352)(49),y=>p(353)(49),Cin=>p(354)(49),clock=>clock,reset=>reset,s=>p(365)(49),cout=>p(366)(50));
FA_ff_14731:FAff port map(x=>p(352)(50),y=>p(353)(50),Cin=>p(354)(50),clock=>clock,reset=>reset,s=>p(365)(50),cout=>p(366)(51));
FA_ff_14732:FAff port map(x=>p(352)(51),y=>p(353)(51),Cin=>p(354)(51),clock=>clock,reset=>reset,s=>p(365)(51),cout=>p(366)(52));
FA_ff_14733:FAff port map(x=>p(352)(52),y=>p(353)(52),Cin=>p(354)(52),clock=>clock,reset=>reset,s=>p(365)(52),cout=>p(366)(53));
FA_ff_14734:FAff port map(x=>p(352)(53),y=>p(353)(53),Cin=>p(354)(53),clock=>clock,reset=>reset,s=>p(365)(53),cout=>p(366)(54));
FA_ff_14735:FAff port map(x=>p(352)(54),y=>p(353)(54),Cin=>p(354)(54),clock=>clock,reset=>reset,s=>p(365)(54),cout=>p(366)(55));
FA_ff_14736:FAff port map(x=>p(352)(55),y=>p(353)(55),Cin=>p(354)(55),clock=>clock,reset=>reset,s=>p(365)(55),cout=>p(366)(56));
FA_ff_14737:FAff port map(x=>p(352)(56),y=>p(353)(56),Cin=>p(354)(56),clock=>clock,reset=>reset,s=>p(365)(56),cout=>p(366)(57));
FA_ff_14738:FAff port map(x=>p(352)(57),y=>p(353)(57),Cin=>p(354)(57),clock=>clock,reset=>reset,s=>p(365)(57),cout=>p(366)(58));
FA_ff_14739:FAff port map(x=>p(352)(58),y=>p(353)(58),Cin=>p(354)(58),clock=>clock,reset=>reset,s=>p(365)(58),cout=>p(366)(59));
FA_ff_14740:FAff port map(x=>p(352)(59),y=>p(353)(59),Cin=>p(354)(59),clock=>clock,reset=>reset,s=>p(365)(59),cout=>p(366)(60));
FA_ff_14741:FAff port map(x=>p(352)(60),y=>p(353)(60),Cin=>p(354)(60),clock=>clock,reset=>reset,s=>p(365)(60),cout=>p(366)(61));
FA_ff_14742:FAff port map(x=>p(352)(61),y=>p(353)(61),Cin=>p(354)(61),clock=>clock,reset=>reset,s=>p(365)(61),cout=>p(366)(62));
FA_ff_14743:FAff port map(x=>p(352)(62),y=>p(353)(62),Cin=>p(354)(62),clock=>clock,reset=>reset,s=>p(365)(62),cout=>p(366)(63));
FA_ff_14744:FAff port map(x=>p(352)(63),y=>p(353)(63),Cin=>p(354)(63),clock=>clock,reset=>reset,s=>p(365)(63),cout=>p(366)(64));
FA_ff_14745:FAff port map(x=>p(352)(64),y=>p(353)(64),Cin=>p(354)(64),clock=>clock,reset=>reset,s=>p(365)(64),cout=>p(366)(65));
FA_ff_14746:FAff port map(x=>p(352)(65),y=>p(353)(65),Cin=>p(354)(65),clock=>clock,reset=>reset,s=>p(365)(65),cout=>p(366)(66));
FA_ff_14747:FAff port map(x=>p(352)(66),y=>p(353)(66),Cin=>p(354)(66),clock=>clock,reset=>reset,s=>p(365)(66),cout=>p(366)(67));
FA_ff_14748:FAff port map(x=>p(352)(67),y=>p(353)(67),Cin=>p(354)(67),clock=>clock,reset=>reset,s=>p(365)(67),cout=>p(366)(68));
FA_ff_14749:FAff port map(x=>p(352)(68),y=>p(353)(68),Cin=>p(354)(68),clock=>clock,reset=>reset,s=>p(365)(68),cout=>p(366)(69));
FA_ff_14750:FAff port map(x=>p(352)(69),y=>p(353)(69),Cin=>p(354)(69),clock=>clock,reset=>reset,s=>p(365)(69),cout=>p(366)(70));
FA_ff_14751:FAff port map(x=>p(352)(70),y=>p(353)(70),Cin=>p(354)(70),clock=>clock,reset=>reset,s=>p(365)(70),cout=>p(366)(71));
FA_ff_14752:FAff port map(x=>p(352)(71),y=>p(353)(71),Cin=>p(354)(71),clock=>clock,reset=>reset,s=>p(365)(71),cout=>p(366)(72));
FA_ff_14753:FAff port map(x=>p(352)(72),y=>p(353)(72),Cin=>p(354)(72),clock=>clock,reset=>reset,s=>p(365)(72),cout=>p(366)(73));
FA_ff_14754:FAff port map(x=>p(352)(73),y=>p(353)(73),Cin=>p(354)(73),clock=>clock,reset=>reset,s=>p(365)(73),cout=>p(366)(74));
FA_ff_14755:FAff port map(x=>p(352)(74),y=>p(353)(74),Cin=>p(354)(74),clock=>clock,reset=>reset,s=>p(365)(74),cout=>p(366)(75));
FA_ff_14756:FAff port map(x=>p(352)(75),y=>p(353)(75),Cin=>p(354)(75),clock=>clock,reset=>reset,s=>p(365)(75),cout=>p(366)(76));
FA_ff_14757:FAff port map(x=>p(352)(76),y=>p(353)(76),Cin=>p(354)(76),clock=>clock,reset=>reset,s=>p(365)(76),cout=>p(366)(77));
FA_ff_14758:FAff port map(x=>p(352)(77),y=>p(353)(77),Cin=>p(354)(77),clock=>clock,reset=>reset,s=>p(365)(77),cout=>p(366)(78));
FA_ff_14759:FAff port map(x=>p(352)(78),y=>p(353)(78),Cin=>p(354)(78),clock=>clock,reset=>reset,s=>p(365)(78),cout=>p(366)(79));
FA_ff_14760:FAff port map(x=>p(352)(79),y=>p(353)(79),Cin=>p(354)(79),clock=>clock,reset=>reset,s=>p(365)(79),cout=>p(366)(80));
FA_ff_14761:FAff port map(x=>p(352)(80),y=>p(353)(80),Cin=>p(354)(80),clock=>clock,reset=>reset,s=>p(365)(80),cout=>p(366)(81));
FA_ff_14762:FAff port map(x=>p(352)(81),y=>p(353)(81),Cin=>p(354)(81),clock=>clock,reset=>reset,s=>p(365)(81),cout=>p(366)(82));
FA_ff_14763:FAff port map(x=>p(352)(82),y=>p(353)(82),Cin=>p(354)(82),clock=>clock,reset=>reset,s=>p(365)(82),cout=>p(366)(83));
FA_ff_14764:FAff port map(x=>p(352)(83),y=>p(353)(83),Cin=>p(354)(83),clock=>clock,reset=>reset,s=>p(365)(83),cout=>p(366)(84));
FA_ff_14765:FAff port map(x=>p(352)(84),y=>p(353)(84),Cin=>p(354)(84),clock=>clock,reset=>reset,s=>p(365)(84),cout=>p(366)(85));
FA_ff_14766:FAff port map(x=>p(352)(85),y=>p(353)(85),Cin=>p(354)(85),clock=>clock,reset=>reset,s=>p(365)(85),cout=>p(366)(86));
FA_ff_14767:FAff port map(x=>p(352)(86),y=>p(353)(86),Cin=>p(354)(86),clock=>clock,reset=>reset,s=>p(365)(86),cout=>p(366)(87));
FA_ff_14768:FAff port map(x=>p(352)(87),y=>p(353)(87),Cin=>p(354)(87),clock=>clock,reset=>reset,s=>p(365)(87),cout=>p(366)(88));
FA_ff_14769:FAff port map(x=>p(352)(88),y=>p(353)(88),Cin=>p(354)(88),clock=>clock,reset=>reset,s=>p(365)(88),cout=>p(366)(89));
FA_ff_14770:FAff port map(x=>p(352)(89),y=>p(353)(89),Cin=>p(354)(89),clock=>clock,reset=>reset,s=>p(365)(89),cout=>p(366)(90));
FA_ff_14771:FAff port map(x=>p(352)(90),y=>p(353)(90),Cin=>p(354)(90),clock=>clock,reset=>reset,s=>p(365)(90),cout=>p(366)(91));
FA_ff_14772:FAff port map(x=>p(352)(91),y=>p(353)(91),Cin=>p(354)(91),clock=>clock,reset=>reset,s=>p(365)(91),cout=>p(366)(92));
FA_ff_14773:FAff port map(x=>p(352)(92),y=>p(353)(92),Cin=>p(354)(92),clock=>clock,reset=>reset,s=>p(365)(92),cout=>p(366)(93));
FA_ff_14774:FAff port map(x=>p(352)(93),y=>p(353)(93),Cin=>p(354)(93),clock=>clock,reset=>reset,s=>p(365)(93),cout=>p(366)(94));
FA_ff_14775:FAff port map(x=>p(352)(94),y=>p(353)(94),Cin=>p(354)(94),clock=>clock,reset=>reset,s=>p(365)(94),cout=>p(366)(95));
FA_ff_14776:FAff port map(x=>p(352)(95),y=>p(353)(95),Cin=>p(354)(95),clock=>clock,reset=>reset,s=>p(365)(95),cout=>p(366)(96));
FA_ff_14777:FAff port map(x=>p(352)(96),y=>p(353)(96),Cin=>p(354)(96),clock=>clock,reset=>reset,s=>p(365)(96),cout=>p(366)(97));
FA_ff_14778:FAff port map(x=>p(352)(97),y=>p(353)(97),Cin=>p(354)(97),clock=>clock,reset=>reset,s=>p(365)(97),cout=>p(366)(98));
FA_ff_14779:FAff port map(x=>p(352)(98),y=>p(353)(98),Cin=>p(354)(98),clock=>clock,reset=>reset,s=>p(365)(98),cout=>p(366)(99));
FA_ff_14780:FAff port map(x=>p(352)(99),y=>p(353)(99),Cin=>p(354)(99),clock=>clock,reset=>reset,s=>p(365)(99),cout=>p(366)(100));
FA_ff_14781:FAff port map(x=>p(352)(100),y=>p(353)(100),Cin=>p(354)(100),clock=>clock,reset=>reset,s=>p(365)(100),cout=>p(366)(101));
FA_ff_14782:FAff port map(x=>p(352)(101),y=>p(353)(101),Cin=>p(354)(101),clock=>clock,reset=>reset,s=>p(365)(101),cout=>p(366)(102));
FA_ff_14783:FAff port map(x=>p(352)(102),y=>p(353)(102),Cin=>p(354)(102),clock=>clock,reset=>reset,s=>p(365)(102),cout=>p(366)(103));
FA_ff_14784:FAff port map(x=>p(352)(103),y=>p(353)(103),Cin=>p(354)(103),clock=>clock,reset=>reset,s=>p(365)(103),cout=>p(366)(104));
FA_ff_14785:FAff port map(x=>p(352)(104),y=>p(353)(104),Cin=>p(354)(104),clock=>clock,reset=>reset,s=>p(365)(104),cout=>p(366)(105));
FA_ff_14786:FAff port map(x=>p(352)(105),y=>p(353)(105),Cin=>p(354)(105),clock=>clock,reset=>reset,s=>p(365)(105),cout=>p(366)(106));
FA_ff_14787:FAff port map(x=>p(352)(106),y=>p(353)(106),Cin=>p(354)(106),clock=>clock,reset=>reset,s=>p(365)(106),cout=>p(366)(107));
FA_ff_14788:FAff port map(x=>p(352)(107),y=>p(353)(107),Cin=>p(354)(107),clock=>clock,reset=>reset,s=>p(365)(107),cout=>p(366)(108));
FA_ff_14789:FAff port map(x=>p(352)(108),y=>p(353)(108),Cin=>p(354)(108),clock=>clock,reset=>reset,s=>p(365)(108),cout=>p(366)(109));
FA_ff_14790:FAff port map(x=>p(352)(109),y=>p(353)(109),Cin=>p(354)(109),clock=>clock,reset=>reset,s=>p(365)(109),cout=>p(366)(110));
FA_ff_14791:FAff port map(x=>p(352)(110),y=>p(353)(110),Cin=>p(354)(110),clock=>clock,reset=>reset,s=>p(365)(110),cout=>p(366)(111));
FA_ff_14792:FAff port map(x=>p(352)(111),y=>p(353)(111),Cin=>p(354)(111),clock=>clock,reset=>reset,s=>p(365)(111),cout=>p(366)(112));
FA_ff_14793:FAff port map(x=>p(352)(112),y=>p(353)(112),Cin=>p(354)(112),clock=>clock,reset=>reset,s=>p(365)(112),cout=>p(366)(113));
FA_ff_14794:FAff port map(x=>p(352)(113),y=>p(353)(113),Cin=>p(354)(113),clock=>clock,reset=>reset,s=>p(365)(113),cout=>p(366)(114));
FA_ff_14795:FAff port map(x=>p(352)(114),y=>p(353)(114),Cin=>p(354)(114),clock=>clock,reset=>reset,s=>p(365)(114),cout=>p(366)(115));
FA_ff_14796:FAff port map(x=>p(352)(115),y=>p(353)(115),Cin=>p(354)(115),clock=>clock,reset=>reset,s=>p(365)(115),cout=>p(366)(116));
FA_ff_14797:FAff port map(x=>p(352)(116),y=>p(353)(116),Cin=>p(354)(116),clock=>clock,reset=>reset,s=>p(365)(116),cout=>p(366)(117));
FA_ff_14798:FAff port map(x=>p(352)(117),y=>p(353)(117),Cin=>p(354)(117),clock=>clock,reset=>reset,s=>p(365)(117),cout=>p(366)(118));
FA_ff_14799:FAff port map(x=>p(352)(118),y=>p(353)(118),Cin=>p(354)(118),clock=>clock,reset=>reset,s=>p(365)(118),cout=>p(366)(119));
FA_ff_14800:FAff port map(x=>p(352)(119),y=>p(353)(119),Cin=>p(354)(119),clock=>clock,reset=>reset,s=>p(365)(119),cout=>p(366)(120));
FA_ff_14801:FAff port map(x=>p(352)(120),y=>p(353)(120),Cin=>p(354)(120),clock=>clock,reset=>reset,s=>p(365)(120),cout=>p(366)(121));
FA_ff_14802:FAff port map(x=>p(352)(121),y=>p(353)(121),Cin=>p(354)(121),clock=>clock,reset=>reset,s=>p(365)(121),cout=>p(366)(122));
FA_ff_14803:FAff port map(x=>p(352)(122),y=>p(353)(122),Cin=>p(354)(122),clock=>clock,reset=>reset,s=>p(365)(122),cout=>p(366)(123));
FA_ff_14804:FAff port map(x=>p(352)(123),y=>p(353)(123),Cin=>p(354)(123),clock=>clock,reset=>reset,s=>p(365)(123),cout=>p(366)(124));
FA_ff_14805:FAff port map(x=>p(352)(124),y=>p(353)(124),Cin=>p(354)(124),clock=>clock,reset=>reset,s=>p(365)(124),cout=>p(366)(125));
FA_ff_14806:FAff port map(x=>p(352)(125),y=>p(353)(125),Cin=>p(354)(125),clock=>clock,reset=>reset,s=>p(365)(125),cout=>p(366)(126));
FA_ff_14807:FAff port map(x=>p(352)(126),y=>p(353)(126),Cin=>p(354)(126),clock=>clock,reset=>reset,s=>p(365)(126),cout=>p(366)(127));
FA_ff_14808:FAff port map(x=>p(352)(127),y=>p(353)(127),Cin=>p(354)(127),clock=>clock,reset=>reset,s=>p(365)(127),cout=>p(366)(128));
FA_ff_14809:FAff port map(x=>p(352)(128),y=>p(353)(128),Cin=>p(354)(128),clock=>clock,reset=>reset,s=>p(365)(128),cout=>p(366)(129));
FA_ff_14810:FAff port map(x=>p(352)(129),y=>p(353)(129),Cin=>p(354)(129),clock=>clock,reset=>reset,s=>p(365)(129),cout=>p(366)(130));
HA_ff_97:HAff port map(x=>p(352)(130),y=>p(354)(130),clock=>clock,reset=>reset,s=>p(365)(130),c=>p(366)(131));
p(365)(131)<=p(352)(131);
HA_ff_98:HAff port map(x=>p(355)(0),y=>p(357)(0),clock=>clock,reset=>reset,s=>p(367)(0),c=>p(368)(1));
FA_ff_14811:FAff port map(x=>p(355)(1),y=>p(356)(1),Cin=>p(357)(1),clock=>clock,reset=>reset,s=>p(367)(1),cout=>p(368)(2));
FA_ff_14812:FAff port map(x=>p(355)(2),y=>p(356)(2),Cin=>p(357)(2),clock=>clock,reset=>reset,s=>p(367)(2),cout=>p(368)(3));
FA_ff_14813:FAff port map(x=>p(355)(3),y=>p(356)(3),Cin=>p(357)(3),clock=>clock,reset=>reset,s=>p(367)(3),cout=>p(368)(4));
FA_ff_14814:FAff port map(x=>p(355)(4),y=>p(356)(4),Cin=>p(357)(4),clock=>clock,reset=>reset,s=>p(367)(4),cout=>p(368)(5));
FA_ff_14815:FAff port map(x=>p(355)(5),y=>p(356)(5),Cin=>p(357)(5),clock=>clock,reset=>reset,s=>p(367)(5),cout=>p(368)(6));
FA_ff_14816:FAff port map(x=>p(355)(6),y=>p(356)(6),Cin=>p(357)(6),clock=>clock,reset=>reset,s=>p(367)(6),cout=>p(368)(7));
FA_ff_14817:FAff port map(x=>p(355)(7),y=>p(356)(7),Cin=>p(357)(7),clock=>clock,reset=>reset,s=>p(367)(7),cout=>p(368)(8));
FA_ff_14818:FAff port map(x=>p(355)(8),y=>p(356)(8),Cin=>p(357)(8),clock=>clock,reset=>reset,s=>p(367)(8),cout=>p(368)(9));
FA_ff_14819:FAff port map(x=>p(355)(9),y=>p(356)(9),Cin=>p(357)(9),clock=>clock,reset=>reset,s=>p(367)(9),cout=>p(368)(10));
FA_ff_14820:FAff port map(x=>p(355)(10),y=>p(356)(10),Cin=>p(357)(10),clock=>clock,reset=>reset,s=>p(367)(10),cout=>p(368)(11));
FA_ff_14821:FAff port map(x=>p(355)(11),y=>p(356)(11),Cin=>p(357)(11),clock=>clock,reset=>reset,s=>p(367)(11),cout=>p(368)(12));
FA_ff_14822:FAff port map(x=>p(355)(12),y=>p(356)(12),Cin=>p(357)(12),clock=>clock,reset=>reset,s=>p(367)(12),cout=>p(368)(13));
FA_ff_14823:FAff port map(x=>p(355)(13),y=>p(356)(13),Cin=>p(357)(13),clock=>clock,reset=>reset,s=>p(367)(13),cout=>p(368)(14));
FA_ff_14824:FAff port map(x=>p(355)(14),y=>p(356)(14),Cin=>p(357)(14),clock=>clock,reset=>reset,s=>p(367)(14),cout=>p(368)(15));
FA_ff_14825:FAff port map(x=>p(355)(15),y=>p(356)(15),Cin=>p(357)(15),clock=>clock,reset=>reset,s=>p(367)(15),cout=>p(368)(16));
FA_ff_14826:FAff port map(x=>p(355)(16),y=>p(356)(16),Cin=>p(357)(16),clock=>clock,reset=>reset,s=>p(367)(16),cout=>p(368)(17));
FA_ff_14827:FAff port map(x=>p(355)(17),y=>p(356)(17),Cin=>p(357)(17),clock=>clock,reset=>reset,s=>p(367)(17),cout=>p(368)(18));
FA_ff_14828:FAff port map(x=>p(355)(18),y=>p(356)(18),Cin=>p(357)(18),clock=>clock,reset=>reset,s=>p(367)(18),cout=>p(368)(19));
FA_ff_14829:FAff port map(x=>p(355)(19),y=>p(356)(19),Cin=>p(357)(19),clock=>clock,reset=>reset,s=>p(367)(19),cout=>p(368)(20));
FA_ff_14830:FAff port map(x=>p(355)(20),y=>p(356)(20),Cin=>p(357)(20),clock=>clock,reset=>reset,s=>p(367)(20),cout=>p(368)(21));
FA_ff_14831:FAff port map(x=>p(355)(21),y=>p(356)(21),Cin=>p(357)(21),clock=>clock,reset=>reset,s=>p(367)(21),cout=>p(368)(22));
FA_ff_14832:FAff port map(x=>p(355)(22),y=>p(356)(22),Cin=>p(357)(22),clock=>clock,reset=>reset,s=>p(367)(22),cout=>p(368)(23));
FA_ff_14833:FAff port map(x=>p(355)(23),y=>p(356)(23),Cin=>p(357)(23),clock=>clock,reset=>reset,s=>p(367)(23),cout=>p(368)(24));
FA_ff_14834:FAff port map(x=>p(355)(24),y=>p(356)(24),Cin=>p(357)(24),clock=>clock,reset=>reset,s=>p(367)(24),cout=>p(368)(25));
FA_ff_14835:FAff port map(x=>p(355)(25),y=>p(356)(25),Cin=>p(357)(25),clock=>clock,reset=>reset,s=>p(367)(25),cout=>p(368)(26));
FA_ff_14836:FAff port map(x=>p(355)(26),y=>p(356)(26),Cin=>p(357)(26),clock=>clock,reset=>reset,s=>p(367)(26),cout=>p(368)(27));
FA_ff_14837:FAff port map(x=>p(355)(27),y=>p(356)(27),Cin=>p(357)(27),clock=>clock,reset=>reset,s=>p(367)(27),cout=>p(368)(28));
FA_ff_14838:FAff port map(x=>p(355)(28),y=>p(356)(28),Cin=>p(357)(28),clock=>clock,reset=>reset,s=>p(367)(28),cout=>p(368)(29));
FA_ff_14839:FAff port map(x=>p(355)(29),y=>p(356)(29),Cin=>p(357)(29),clock=>clock,reset=>reset,s=>p(367)(29),cout=>p(368)(30));
FA_ff_14840:FAff port map(x=>p(355)(30),y=>p(356)(30),Cin=>p(357)(30),clock=>clock,reset=>reset,s=>p(367)(30),cout=>p(368)(31));
FA_ff_14841:FAff port map(x=>p(355)(31),y=>p(356)(31),Cin=>p(357)(31),clock=>clock,reset=>reset,s=>p(367)(31),cout=>p(368)(32));
FA_ff_14842:FAff port map(x=>p(355)(32),y=>p(356)(32),Cin=>p(357)(32),clock=>clock,reset=>reset,s=>p(367)(32),cout=>p(368)(33));
FA_ff_14843:FAff port map(x=>p(355)(33),y=>p(356)(33),Cin=>p(357)(33),clock=>clock,reset=>reset,s=>p(367)(33),cout=>p(368)(34));
FA_ff_14844:FAff port map(x=>p(355)(34),y=>p(356)(34),Cin=>p(357)(34),clock=>clock,reset=>reset,s=>p(367)(34),cout=>p(368)(35));
FA_ff_14845:FAff port map(x=>p(355)(35),y=>p(356)(35),Cin=>p(357)(35),clock=>clock,reset=>reset,s=>p(367)(35),cout=>p(368)(36));
FA_ff_14846:FAff port map(x=>p(355)(36),y=>p(356)(36),Cin=>p(357)(36),clock=>clock,reset=>reset,s=>p(367)(36),cout=>p(368)(37));
FA_ff_14847:FAff port map(x=>p(355)(37),y=>p(356)(37),Cin=>p(357)(37),clock=>clock,reset=>reset,s=>p(367)(37),cout=>p(368)(38));
FA_ff_14848:FAff port map(x=>p(355)(38),y=>p(356)(38),Cin=>p(357)(38),clock=>clock,reset=>reset,s=>p(367)(38),cout=>p(368)(39));
FA_ff_14849:FAff port map(x=>p(355)(39),y=>p(356)(39),Cin=>p(357)(39),clock=>clock,reset=>reset,s=>p(367)(39),cout=>p(368)(40));
FA_ff_14850:FAff port map(x=>p(355)(40),y=>p(356)(40),Cin=>p(357)(40),clock=>clock,reset=>reset,s=>p(367)(40),cout=>p(368)(41));
FA_ff_14851:FAff port map(x=>p(355)(41),y=>p(356)(41),Cin=>p(357)(41),clock=>clock,reset=>reset,s=>p(367)(41),cout=>p(368)(42));
FA_ff_14852:FAff port map(x=>p(355)(42),y=>p(356)(42),Cin=>p(357)(42),clock=>clock,reset=>reset,s=>p(367)(42),cout=>p(368)(43));
FA_ff_14853:FAff port map(x=>p(355)(43),y=>p(356)(43),Cin=>p(357)(43),clock=>clock,reset=>reset,s=>p(367)(43),cout=>p(368)(44));
FA_ff_14854:FAff port map(x=>p(355)(44),y=>p(356)(44),Cin=>p(357)(44),clock=>clock,reset=>reset,s=>p(367)(44),cout=>p(368)(45));
FA_ff_14855:FAff port map(x=>p(355)(45),y=>p(356)(45),Cin=>p(357)(45),clock=>clock,reset=>reset,s=>p(367)(45),cout=>p(368)(46));
FA_ff_14856:FAff port map(x=>p(355)(46),y=>p(356)(46),Cin=>p(357)(46),clock=>clock,reset=>reset,s=>p(367)(46),cout=>p(368)(47));
FA_ff_14857:FAff port map(x=>p(355)(47),y=>p(356)(47),Cin=>p(357)(47),clock=>clock,reset=>reset,s=>p(367)(47),cout=>p(368)(48));
FA_ff_14858:FAff port map(x=>p(355)(48),y=>p(356)(48),Cin=>p(357)(48),clock=>clock,reset=>reset,s=>p(367)(48),cout=>p(368)(49));
FA_ff_14859:FAff port map(x=>p(355)(49),y=>p(356)(49),Cin=>p(357)(49),clock=>clock,reset=>reset,s=>p(367)(49),cout=>p(368)(50));
FA_ff_14860:FAff port map(x=>p(355)(50),y=>p(356)(50),Cin=>p(357)(50),clock=>clock,reset=>reset,s=>p(367)(50),cout=>p(368)(51));
FA_ff_14861:FAff port map(x=>p(355)(51),y=>p(356)(51),Cin=>p(357)(51),clock=>clock,reset=>reset,s=>p(367)(51),cout=>p(368)(52));
FA_ff_14862:FAff port map(x=>p(355)(52),y=>p(356)(52),Cin=>p(357)(52),clock=>clock,reset=>reset,s=>p(367)(52),cout=>p(368)(53));
FA_ff_14863:FAff port map(x=>p(355)(53),y=>p(356)(53),Cin=>p(357)(53),clock=>clock,reset=>reset,s=>p(367)(53),cout=>p(368)(54));
FA_ff_14864:FAff port map(x=>p(355)(54),y=>p(356)(54),Cin=>p(357)(54),clock=>clock,reset=>reset,s=>p(367)(54),cout=>p(368)(55));
FA_ff_14865:FAff port map(x=>p(355)(55),y=>p(356)(55),Cin=>p(357)(55),clock=>clock,reset=>reset,s=>p(367)(55),cout=>p(368)(56));
FA_ff_14866:FAff port map(x=>p(355)(56),y=>p(356)(56),Cin=>p(357)(56),clock=>clock,reset=>reset,s=>p(367)(56),cout=>p(368)(57));
FA_ff_14867:FAff port map(x=>p(355)(57),y=>p(356)(57),Cin=>p(357)(57),clock=>clock,reset=>reset,s=>p(367)(57),cout=>p(368)(58));
FA_ff_14868:FAff port map(x=>p(355)(58),y=>p(356)(58),Cin=>p(357)(58),clock=>clock,reset=>reset,s=>p(367)(58),cout=>p(368)(59));
FA_ff_14869:FAff port map(x=>p(355)(59),y=>p(356)(59),Cin=>p(357)(59),clock=>clock,reset=>reset,s=>p(367)(59),cout=>p(368)(60));
FA_ff_14870:FAff port map(x=>p(355)(60),y=>p(356)(60),Cin=>p(357)(60),clock=>clock,reset=>reset,s=>p(367)(60),cout=>p(368)(61));
FA_ff_14871:FAff port map(x=>p(355)(61),y=>p(356)(61),Cin=>p(357)(61),clock=>clock,reset=>reset,s=>p(367)(61),cout=>p(368)(62));
FA_ff_14872:FAff port map(x=>p(355)(62),y=>p(356)(62),Cin=>p(357)(62),clock=>clock,reset=>reset,s=>p(367)(62),cout=>p(368)(63));
FA_ff_14873:FAff port map(x=>p(355)(63),y=>p(356)(63),Cin=>p(357)(63),clock=>clock,reset=>reset,s=>p(367)(63),cout=>p(368)(64));
FA_ff_14874:FAff port map(x=>p(355)(64),y=>p(356)(64),Cin=>p(357)(64),clock=>clock,reset=>reset,s=>p(367)(64),cout=>p(368)(65));
FA_ff_14875:FAff port map(x=>p(355)(65),y=>p(356)(65),Cin=>p(357)(65),clock=>clock,reset=>reset,s=>p(367)(65),cout=>p(368)(66));
FA_ff_14876:FAff port map(x=>p(355)(66),y=>p(356)(66),Cin=>p(357)(66),clock=>clock,reset=>reset,s=>p(367)(66),cout=>p(368)(67));
FA_ff_14877:FAff port map(x=>p(355)(67),y=>p(356)(67),Cin=>p(357)(67),clock=>clock,reset=>reset,s=>p(367)(67),cout=>p(368)(68));
FA_ff_14878:FAff port map(x=>p(355)(68),y=>p(356)(68),Cin=>p(357)(68),clock=>clock,reset=>reset,s=>p(367)(68),cout=>p(368)(69));
FA_ff_14879:FAff port map(x=>p(355)(69),y=>p(356)(69),Cin=>p(357)(69),clock=>clock,reset=>reset,s=>p(367)(69),cout=>p(368)(70));
FA_ff_14880:FAff port map(x=>p(355)(70),y=>p(356)(70),Cin=>p(357)(70),clock=>clock,reset=>reset,s=>p(367)(70),cout=>p(368)(71));
FA_ff_14881:FAff port map(x=>p(355)(71),y=>p(356)(71),Cin=>p(357)(71),clock=>clock,reset=>reset,s=>p(367)(71),cout=>p(368)(72));
FA_ff_14882:FAff port map(x=>p(355)(72),y=>p(356)(72),Cin=>p(357)(72),clock=>clock,reset=>reset,s=>p(367)(72),cout=>p(368)(73));
FA_ff_14883:FAff port map(x=>p(355)(73),y=>p(356)(73),Cin=>p(357)(73),clock=>clock,reset=>reset,s=>p(367)(73),cout=>p(368)(74));
FA_ff_14884:FAff port map(x=>p(355)(74),y=>p(356)(74),Cin=>p(357)(74),clock=>clock,reset=>reset,s=>p(367)(74),cout=>p(368)(75));
FA_ff_14885:FAff port map(x=>p(355)(75),y=>p(356)(75),Cin=>p(357)(75),clock=>clock,reset=>reset,s=>p(367)(75),cout=>p(368)(76));
FA_ff_14886:FAff port map(x=>p(355)(76),y=>p(356)(76),Cin=>p(357)(76),clock=>clock,reset=>reset,s=>p(367)(76),cout=>p(368)(77));
FA_ff_14887:FAff port map(x=>p(355)(77),y=>p(356)(77),Cin=>p(357)(77),clock=>clock,reset=>reset,s=>p(367)(77),cout=>p(368)(78));
FA_ff_14888:FAff port map(x=>p(355)(78),y=>p(356)(78),Cin=>p(357)(78),clock=>clock,reset=>reset,s=>p(367)(78),cout=>p(368)(79));
FA_ff_14889:FAff port map(x=>p(355)(79),y=>p(356)(79),Cin=>p(357)(79),clock=>clock,reset=>reset,s=>p(367)(79),cout=>p(368)(80));
FA_ff_14890:FAff port map(x=>p(355)(80),y=>p(356)(80),Cin=>p(357)(80),clock=>clock,reset=>reset,s=>p(367)(80),cout=>p(368)(81));
FA_ff_14891:FAff port map(x=>p(355)(81),y=>p(356)(81),Cin=>p(357)(81),clock=>clock,reset=>reset,s=>p(367)(81),cout=>p(368)(82));
FA_ff_14892:FAff port map(x=>p(355)(82),y=>p(356)(82),Cin=>p(357)(82),clock=>clock,reset=>reset,s=>p(367)(82),cout=>p(368)(83));
FA_ff_14893:FAff port map(x=>p(355)(83),y=>p(356)(83),Cin=>p(357)(83),clock=>clock,reset=>reset,s=>p(367)(83),cout=>p(368)(84));
FA_ff_14894:FAff port map(x=>p(355)(84),y=>p(356)(84),Cin=>p(357)(84),clock=>clock,reset=>reset,s=>p(367)(84),cout=>p(368)(85));
FA_ff_14895:FAff port map(x=>p(355)(85),y=>p(356)(85),Cin=>p(357)(85),clock=>clock,reset=>reset,s=>p(367)(85),cout=>p(368)(86));
FA_ff_14896:FAff port map(x=>p(355)(86),y=>p(356)(86),Cin=>p(357)(86),clock=>clock,reset=>reset,s=>p(367)(86),cout=>p(368)(87));
FA_ff_14897:FAff port map(x=>p(355)(87),y=>p(356)(87),Cin=>p(357)(87),clock=>clock,reset=>reset,s=>p(367)(87),cout=>p(368)(88));
FA_ff_14898:FAff port map(x=>p(355)(88),y=>p(356)(88),Cin=>p(357)(88),clock=>clock,reset=>reset,s=>p(367)(88),cout=>p(368)(89));
FA_ff_14899:FAff port map(x=>p(355)(89),y=>p(356)(89),Cin=>p(357)(89),clock=>clock,reset=>reset,s=>p(367)(89),cout=>p(368)(90));
FA_ff_14900:FAff port map(x=>p(355)(90),y=>p(356)(90),Cin=>p(357)(90),clock=>clock,reset=>reset,s=>p(367)(90),cout=>p(368)(91));
FA_ff_14901:FAff port map(x=>p(355)(91),y=>p(356)(91),Cin=>p(357)(91),clock=>clock,reset=>reset,s=>p(367)(91),cout=>p(368)(92));
FA_ff_14902:FAff port map(x=>p(355)(92),y=>p(356)(92),Cin=>p(357)(92),clock=>clock,reset=>reset,s=>p(367)(92),cout=>p(368)(93));
FA_ff_14903:FAff port map(x=>p(355)(93),y=>p(356)(93),Cin=>p(357)(93),clock=>clock,reset=>reset,s=>p(367)(93),cout=>p(368)(94));
FA_ff_14904:FAff port map(x=>p(355)(94),y=>p(356)(94),Cin=>p(357)(94),clock=>clock,reset=>reset,s=>p(367)(94),cout=>p(368)(95));
FA_ff_14905:FAff port map(x=>p(355)(95),y=>p(356)(95),Cin=>p(357)(95),clock=>clock,reset=>reset,s=>p(367)(95),cout=>p(368)(96));
FA_ff_14906:FAff port map(x=>p(355)(96),y=>p(356)(96),Cin=>p(357)(96),clock=>clock,reset=>reset,s=>p(367)(96),cout=>p(368)(97));
FA_ff_14907:FAff port map(x=>p(355)(97),y=>p(356)(97),Cin=>p(357)(97),clock=>clock,reset=>reset,s=>p(367)(97),cout=>p(368)(98));
FA_ff_14908:FAff port map(x=>p(355)(98),y=>p(356)(98),Cin=>p(357)(98),clock=>clock,reset=>reset,s=>p(367)(98),cout=>p(368)(99));
FA_ff_14909:FAff port map(x=>p(355)(99),y=>p(356)(99),Cin=>p(357)(99),clock=>clock,reset=>reset,s=>p(367)(99),cout=>p(368)(100));
FA_ff_14910:FAff port map(x=>p(355)(100),y=>p(356)(100),Cin=>p(357)(100),clock=>clock,reset=>reset,s=>p(367)(100),cout=>p(368)(101));
FA_ff_14911:FAff port map(x=>p(355)(101),y=>p(356)(101),Cin=>p(357)(101),clock=>clock,reset=>reset,s=>p(367)(101),cout=>p(368)(102));
FA_ff_14912:FAff port map(x=>p(355)(102),y=>p(356)(102),Cin=>p(357)(102),clock=>clock,reset=>reset,s=>p(367)(102),cout=>p(368)(103));
FA_ff_14913:FAff port map(x=>p(355)(103),y=>p(356)(103),Cin=>p(357)(103),clock=>clock,reset=>reset,s=>p(367)(103),cout=>p(368)(104));
FA_ff_14914:FAff port map(x=>p(355)(104),y=>p(356)(104),Cin=>p(357)(104),clock=>clock,reset=>reset,s=>p(367)(104),cout=>p(368)(105));
FA_ff_14915:FAff port map(x=>p(355)(105),y=>p(356)(105),Cin=>p(357)(105),clock=>clock,reset=>reset,s=>p(367)(105),cout=>p(368)(106));
FA_ff_14916:FAff port map(x=>p(355)(106),y=>p(356)(106),Cin=>p(357)(106),clock=>clock,reset=>reset,s=>p(367)(106),cout=>p(368)(107));
FA_ff_14917:FAff port map(x=>p(355)(107),y=>p(356)(107),Cin=>p(357)(107),clock=>clock,reset=>reset,s=>p(367)(107),cout=>p(368)(108));
FA_ff_14918:FAff port map(x=>p(355)(108),y=>p(356)(108),Cin=>p(357)(108),clock=>clock,reset=>reset,s=>p(367)(108),cout=>p(368)(109));
FA_ff_14919:FAff port map(x=>p(355)(109),y=>p(356)(109),Cin=>p(357)(109),clock=>clock,reset=>reset,s=>p(367)(109),cout=>p(368)(110));
FA_ff_14920:FAff port map(x=>p(355)(110),y=>p(356)(110),Cin=>p(357)(110),clock=>clock,reset=>reset,s=>p(367)(110),cout=>p(368)(111));
FA_ff_14921:FAff port map(x=>p(355)(111),y=>p(356)(111),Cin=>p(357)(111),clock=>clock,reset=>reset,s=>p(367)(111),cout=>p(368)(112));
FA_ff_14922:FAff port map(x=>p(355)(112),y=>p(356)(112),Cin=>p(357)(112),clock=>clock,reset=>reset,s=>p(367)(112),cout=>p(368)(113));
FA_ff_14923:FAff port map(x=>p(355)(113),y=>p(356)(113),Cin=>p(357)(113),clock=>clock,reset=>reset,s=>p(367)(113),cout=>p(368)(114));
FA_ff_14924:FAff port map(x=>p(355)(114),y=>p(356)(114),Cin=>p(357)(114),clock=>clock,reset=>reset,s=>p(367)(114),cout=>p(368)(115));
FA_ff_14925:FAff port map(x=>p(355)(115),y=>p(356)(115),Cin=>p(357)(115),clock=>clock,reset=>reset,s=>p(367)(115),cout=>p(368)(116));
FA_ff_14926:FAff port map(x=>p(355)(116),y=>p(356)(116),Cin=>p(357)(116),clock=>clock,reset=>reset,s=>p(367)(116),cout=>p(368)(117));
FA_ff_14927:FAff port map(x=>p(355)(117),y=>p(356)(117),Cin=>p(357)(117),clock=>clock,reset=>reset,s=>p(367)(117),cout=>p(368)(118));
FA_ff_14928:FAff port map(x=>p(355)(118),y=>p(356)(118),Cin=>p(357)(118),clock=>clock,reset=>reset,s=>p(367)(118),cout=>p(368)(119));
FA_ff_14929:FAff port map(x=>p(355)(119),y=>p(356)(119),Cin=>p(357)(119),clock=>clock,reset=>reset,s=>p(367)(119),cout=>p(368)(120));
FA_ff_14930:FAff port map(x=>p(355)(120),y=>p(356)(120),Cin=>p(357)(120),clock=>clock,reset=>reset,s=>p(367)(120),cout=>p(368)(121));
FA_ff_14931:FAff port map(x=>p(355)(121),y=>p(356)(121),Cin=>p(357)(121),clock=>clock,reset=>reset,s=>p(367)(121),cout=>p(368)(122));
FA_ff_14932:FAff port map(x=>p(355)(122),y=>p(356)(122),Cin=>p(357)(122),clock=>clock,reset=>reset,s=>p(367)(122),cout=>p(368)(123));
FA_ff_14933:FAff port map(x=>p(355)(123),y=>p(356)(123),Cin=>p(357)(123),clock=>clock,reset=>reset,s=>p(367)(123),cout=>p(368)(124));
FA_ff_14934:FAff port map(x=>p(355)(124),y=>p(356)(124),Cin=>p(357)(124),clock=>clock,reset=>reset,s=>p(367)(124),cout=>p(368)(125));
FA_ff_14935:FAff port map(x=>p(355)(125),y=>p(356)(125),Cin=>p(357)(125),clock=>clock,reset=>reset,s=>p(367)(125),cout=>p(368)(126));
FA_ff_14936:FAff port map(x=>p(355)(126),y=>p(356)(126),Cin=>p(357)(126),clock=>clock,reset=>reset,s=>p(367)(126),cout=>p(368)(127));
FA_ff_14937:FAff port map(x=>p(355)(127),y=>p(356)(127),Cin=>p(357)(127),clock=>clock,reset=>reset,s=>p(367)(127),cout=>p(368)(128));
FA_ff_14938:FAff port map(x=>p(355)(128),y=>p(356)(128),Cin=>p(357)(128),clock=>clock,reset=>reset,s=>p(367)(128),cout=>p(368)(129));
FA_ff_14939:FAff port map(x=>p(355)(129),y=>p(356)(129),Cin=>p(357)(129),clock=>clock,reset=>reset,s=>p(367)(129),cout=>p(368)(130));
FA_ff_14940:FAff port map(x=>p(355)(130),y=>p(356)(130),Cin=>p(357)(130),clock=>clock,reset=>reset,s=>p(367)(130),cout=>p(368)(131));
HA_ff_99:HAff port map(x=>p(356)(131),y=>p(357)(131),clock=>clock,reset=>reset,s=>p(367)(131),c=>p(368)(132));
p(369)(0)<=p(359)(0);
HA_ff_100:HAff port map(x=>p(359)(1),y=>p(360)(1),clock=>clock,reset=>reset,s=>p(369)(1),c=>p(370)(2));
FA_ff_14941:FAff port map(x=>p(358)(2),y=>p(359)(2),Cin=>p(360)(2),clock=>clock,reset=>reset,s=>p(369)(2),cout=>p(370)(3));
FA_ff_14942:FAff port map(x=>p(358)(3),y=>p(359)(3),Cin=>p(360)(3),clock=>clock,reset=>reset,s=>p(369)(3),cout=>p(370)(4));
FA_ff_14943:FAff port map(x=>p(358)(4),y=>p(359)(4),Cin=>p(360)(4),clock=>clock,reset=>reset,s=>p(369)(4),cout=>p(370)(5));
FA_ff_14944:FAff port map(x=>p(358)(5),y=>p(359)(5),Cin=>p(360)(5),clock=>clock,reset=>reset,s=>p(369)(5),cout=>p(370)(6));
FA_ff_14945:FAff port map(x=>p(358)(6),y=>p(359)(6),Cin=>p(360)(6),clock=>clock,reset=>reset,s=>p(369)(6),cout=>p(370)(7));
FA_ff_14946:FAff port map(x=>p(358)(7),y=>p(359)(7),Cin=>p(360)(7),clock=>clock,reset=>reset,s=>p(369)(7),cout=>p(370)(8));
FA_ff_14947:FAff port map(x=>p(358)(8),y=>p(359)(8),Cin=>p(360)(8),clock=>clock,reset=>reset,s=>p(369)(8),cout=>p(370)(9));
FA_ff_14948:FAff port map(x=>p(358)(9),y=>p(359)(9),Cin=>p(360)(9),clock=>clock,reset=>reset,s=>p(369)(9),cout=>p(370)(10));
FA_ff_14949:FAff port map(x=>p(358)(10),y=>p(359)(10),Cin=>p(360)(10),clock=>clock,reset=>reset,s=>p(369)(10),cout=>p(370)(11));
FA_ff_14950:FAff port map(x=>p(358)(11),y=>p(359)(11),Cin=>p(360)(11),clock=>clock,reset=>reset,s=>p(369)(11),cout=>p(370)(12));
FA_ff_14951:FAff port map(x=>p(358)(12),y=>p(359)(12),Cin=>p(360)(12),clock=>clock,reset=>reset,s=>p(369)(12),cout=>p(370)(13));
FA_ff_14952:FAff port map(x=>p(358)(13),y=>p(359)(13),Cin=>p(360)(13),clock=>clock,reset=>reset,s=>p(369)(13),cout=>p(370)(14));
FA_ff_14953:FAff port map(x=>p(358)(14),y=>p(359)(14),Cin=>p(360)(14),clock=>clock,reset=>reset,s=>p(369)(14),cout=>p(370)(15));
FA_ff_14954:FAff port map(x=>p(358)(15),y=>p(359)(15),Cin=>p(360)(15),clock=>clock,reset=>reset,s=>p(369)(15),cout=>p(370)(16));
FA_ff_14955:FAff port map(x=>p(358)(16),y=>p(359)(16),Cin=>p(360)(16),clock=>clock,reset=>reset,s=>p(369)(16),cout=>p(370)(17));
FA_ff_14956:FAff port map(x=>p(358)(17),y=>p(359)(17),Cin=>p(360)(17),clock=>clock,reset=>reset,s=>p(369)(17),cout=>p(370)(18));
FA_ff_14957:FAff port map(x=>p(358)(18),y=>p(359)(18),Cin=>p(360)(18),clock=>clock,reset=>reset,s=>p(369)(18),cout=>p(370)(19));
FA_ff_14958:FAff port map(x=>p(358)(19),y=>p(359)(19),Cin=>p(360)(19),clock=>clock,reset=>reset,s=>p(369)(19),cout=>p(370)(20));
FA_ff_14959:FAff port map(x=>p(358)(20),y=>p(359)(20),Cin=>p(360)(20),clock=>clock,reset=>reset,s=>p(369)(20),cout=>p(370)(21));
FA_ff_14960:FAff port map(x=>p(358)(21),y=>p(359)(21),Cin=>p(360)(21),clock=>clock,reset=>reset,s=>p(369)(21),cout=>p(370)(22));
FA_ff_14961:FAff port map(x=>p(358)(22),y=>p(359)(22),Cin=>p(360)(22),clock=>clock,reset=>reset,s=>p(369)(22),cout=>p(370)(23));
FA_ff_14962:FAff port map(x=>p(358)(23),y=>p(359)(23),Cin=>p(360)(23),clock=>clock,reset=>reset,s=>p(369)(23),cout=>p(370)(24));
FA_ff_14963:FAff port map(x=>p(358)(24),y=>p(359)(24),Cin=>p(360)(24),clock=>clock,reset=>reset,s=>p(369)(24),cout=>p(370)(25));
FA_ff_14964:FAff port map(x=>p(358)(25),y=>p(359)(25),Cin=>p(360)(25),clock=>clock,reset=>reset,s=>p(369)(25),cout=>p(370)(26));
FA_ff_14965:FAff port map(x=>p(358)(26),y=>p(359)(26),Cin=>p(360)(26),clock=>clock,reset=>reset,s=>p(369)(26),cout=>p(370)(27));
FA_ff_14966:FAff port map(x=>p(358)(27),y=>p(359)(27),Cin=>p(360)(27),clock=>clock,reset=>reset,s=>p(369)(27),cout=>p(370)(28));
FA_ff_14967:FAff port map(x=>p(358)(28),y=>p(359)(28),Cin=>p(360)(28),clock=>clock,reset=>reset,s=>p(369)(28),cout=>p(370)(29));
FA_ff_14968:FAff port map(x=>p(358)(29),y=>p(359)(29),Cin=>p(360)(29),clock=>clock,reset=>reset,s=>p(369)(29),cout=>p(370)(30));
FA_ff_14969:FAff port map(x=>p(358)(30),y=>p(359)(30),Cin=>p(360)(30),clock=>clock,reset=>reset,s=>p(369)(30),cout=>p(370)(31));
FA_ff_14970:FAff port map(x=>p(358)(31),y=>p(359)(31),Cin=>p(360)(31),clock=>clock,reset=>reset,s=>p(369)(31),cout=>p(370)(32));
FA_ff_14971:FAff port map(x=>p(358)(32),y=>p(359)(32),Cin=>p(360)(32),clock=>clock,reset=>reset,s=>p(369)(32),cout=>p(370)(33));
FA_ff_14972:FAff port map(x=>p(358)(33),y=>p(359)(33),Cin=>p(360)(33),clock=>clock,reset=>reset,s=>p(369)(33),cout=>p(370)(34));
FA_ff_14973:FAff port map(x=>p(358)(34),y=>p(359)(34),Cin=>p(360)(34),clock=>clock,reset=>reset,s=>p(369)(34),cout=>p(370)(35));
FA_ff_14974:FAff port map(x=>p(358)(35),y=>p(359)(35),Cin=>p(360)(35),clock=>clock,reset=>reset,s=>p(369)(35),cout=>p(370)(36));
FA_ff_14975:FAff port map(x=>p(358)(36),y=>p(359)(36),Cin=>p(360)(36),clock=>clock,reset=>reset,s=>p(369)(36),cout=>p(370)(37));
FA_ff_14976:FAff port map(x=>p(358)(37),y=>p(359)(37),Cin=>p(360)(37),clock=>clock,reset=>reset,s=>p(369)(37),cout=>p(370)(38));
FA_ff_14977:FAff port map(x=>p(358)(38),y=>p(359)(38),Cin=>p(360)(38),clock=>clock,reset=>reset,s=>p(369)(38),cout=>p(370)(39));
FA_ff_14978:FAff port map(x=>p(358)(39),y=>p(359)(39),Cin=>p(360)(39),clock=>clock,reset=>reset,s=>p(369)(39),cout=>p(370)(40));
FA_ff_14979:FAff port map(x=>p(358)(40),y=>p(359)(40),Cin=>p(360)(40),clock=>clock,reset=>reset,s=>p(369)(40),cout=>p(370)(41));
FA_ff_14980:FAff port map(x=>p(358)(41),y=>p(359)(41),Cin=>p(360)(41),clock=>clock,reset=>reset,s=>p(369)(41),cout=>p(370)(42));
FA_ff_14981:FAff port map(x=>p(358)(42),y=>p(359)(42),Cin=>p(360)(42),clock=>clock,reset=>reset,s=>p(369)(42),cout=>p(370)(43));
FA_ff_14982:FAff port map(x=>p(358)(43),y=>p(359)(43),Cin=>p(360)(43),clock=>clock,reset=>reset,s=>p(369)(43),cout=>p(370)(44));
FA_ff_14983:FAff port map(x=>p(358)(44),y=>p(359)(44),Cin=>p(360)(44),clock=>clock,reset=>reset,s=>p(369)(44),cout=>p(370)(45));
FA_ff_14984:FAff port map(x=>p(358)(45),y=>p(359)(45),Cin=>p(360)(45),clock=>clock,reset=>reset,s=>p(369)(45),cout=>p(370)(46));
FA_ff_14985:FAff port map(x=>p(358)(46),y=>p(359)(46),Cin=>p(360)(46),clock=>clock,reset=>reset,s=>p(369)(46),cout=>p(370)(47));
FA_ff_14986:FAff port map(x=>p(358)(47),y=>p(359)(47),Cin=>p(360)(47),clock=>clock,reset=>reset,s=>p(369)(47),cout=>p(370)(48));
FA_ff_14987:FAff port map(x=>p(358)(48),y=>p(359)(48),Cin=>p(360)(48),clock=>clock,reset=>reset,s=>p(369)(48),cout=>p(370)(49));
FA_ff_14988:FAff port map(x=>p(358)(49),y=>p(359)(49),Cin=>p(360)(49),clock=>clock,reset=>reset,s=>p(369)(49),cout=>p(370)(50));
FA_ff_14989:FAff port map(x=>p(358)(50),y=>p(359)(50),Cin=>p(360)(50),clock=>clock,reset=>reset,s=>p(369)(50),cout=>p(370)(51));
FA_ff_14990:FAff port map(x=>p(358)(51),y=>p(359)(51),Cin=>p(360)(51),clock=>clock,reset=>reset,s=>p(369)(51),cout=>p(370)(52));
FA_ff_14991:FAff port map(x=>p(358)(52),y=>p(359)(52),Cin=>p(360)(52),clock=>clock,reset=>reset,s=>p(369)(52),cout=>p(370)(53));
FA_ff_14992:FAff port map(x=>p(358)(53),y=>p(359)(53),Cin=>p(360)(53),clock=>clock,reset=>reset,s=>p(369)(53),cout=>p(370)(54));
FA_ff_14993:FAff port map(x=>p(358)(54),y=>p(359)(54),Cin=>p(360)(54),clock=>clock,reset=>reset,s=>p(369)(54),cout=>p(370)(55));
FA_ff_14994:FAff port map(x=>p(358)(55),y=>p(359)(55),Cin=>p(360)(55),clock=>clock,reset=>reset,s=>p(369)(55),cout=>p(370)(56));
FA_ff_14995:FAff port map(x=>p(358)(56),y=>p(359)(56),Cin=>p(360)(56),clock=>clock,reset=>reset,s=>p(369)(56),cout=>p(370)(57));
FA_ff_14996:FAff port map(x=>p(358)(57),y=>p(359)(57),Cin=>p(360)(57),clock=>clock,reset=>reset,s=>p(369)(57),cout=>p(370)(58));
FA_ff_14997:FAff port map(x=>p(358)(58),y=>p(359)(58),Cin=>p(360)(58),clock=>clock,reset=>reset,s=>p(369)(58),cout=>p(370)(59));
FA_ff_14998:FAff port map(x=>p(358)(59),y=>p(359)(59),Cin=>p(360)(59),clock=>clock,reset=>reset,s=>p(369)(59),cout=>p(370)(60));
FA_ff_14999:FAff port map(x=>p(358)(60),y=>p(359)(60),Cin=>p(360)(60),clock=>clock,reset=>reset,s=>p(369)(60),cout=>p(370)(61));
FA_ff_15000:FAff port map(x=>p(358)(61),y=>p(359)(61),Cin=>p(360)(61),clock=>clock,reset=>reset,s=>p(369)(61),cout=>p(370)(62));
FA_ff_15001:FAff port map(x=>p(358)(62),y=>p(359)(62),Cin=>p(360)(62),clock=>clock,reset=>reset,s=>p(369)(62),cout=>p(370)(63));
FA_ff_15002:FAff port map(x=>p(358)(63),y=>p(359)(63),Cin=>p(360)(63),clock=>clock,reset=>reset,s=>p(369)(63),cout=>p(370)(64));
FA_ff_15003:FAff port map(x=>p(358)(64),y=>p(359)(64),Cin=>p(360)(64),clock=>clock,reset=>reset,s=>p(369)(64),cout=>p(370)(65));
FA_ff_15004:FAff port map(x=>p(358)(65),y=>p(359)(65),Cin=>p(360)(65),clock=>clock,reset=>reset,s=>p(369)(65),cout=>p(370)(66));
FA_ff_15005:FAff port map(x=>p(358)(66),y=>p(359)(66),Cin=>p(360)(66),clock=>clock,reset=>reset,s=>p(369)(66),cout=>p(370)(67));
FA_ff_15006:FAff port map(x=>p(358)(67),y=>p(359)(67),Cin=>p(360)(67),clock=>clock,reset=>reset,s=>p(369)(67),cout=>p(370)(68));
FA_ff_15007:FAff port map(x=>p(358)(68),y=>p(359)(68),Cin=>p(360)(68),clock=>clock,reset=>reset,s=>p(369)(68),cout=>p(370)(69));
FA_ff_15008:FAff port map(x=>p(358)(69),y=>p(359)(69),Cin=>p(360)(69),clock=>clock,reset=>reset,s=>p(369)(69),cout=>p(370)(70));
FA_ff_15009:FAff port map(x=>p(358)(70),y=>p(359)(70),Cin=>p(360)(70),clock=>clock,reset=>reset,s=>p(369)(70),cout=>p(370)(71));
FA_ff_15010:FAff port map(x=>p(358)(71),y=>p(359)(71),Cin=>p(360)(71),clock=>clock,reset=>reset,s=>p(369)(71),cout=>p(370)(72));
FA_ff_15011:FAff port map(x=>p(358)(72),y=>p(359)(72),Cin=>p(360)(72),clock=>clock,reset=>reset,s=>p(369)(72),cout=>p(370)(73));
FA_ff_15012:FAff port map(x=>p(358)(73),y=>p(359)(73),Cin=>p(360)(73),clock=>clock,reset=>reset,s=>p(369)(73),cout=>p(370)(74));
FA_ff_15013:FAff port map(x=>p(358)(74),y=>p(359)(74),Cin=>p(360)(74),clock=>clock,reset=>reset,s=>p(369)(74),cout=>p(370)(75));
FA_ff_15014:FAff port map(x=>p(358)(75),y=>p(359)(75),Cin=>p(360)(75),clock=>clock,reset=>reset,s=>p(369)(75),cout=>p(370)(76));
FA_ff_15015:FAff port map(x=>p(358)(76),y=>p(359)(76),Cin=>p(360)(76),clock=>clock,reset=>reset,s=>p(369)(76),cout=>p(370)(77));
FA_ff_15016:FAff port map(x=>p(358)(77),y=>p(359)(77),Cin=>p(360)(77),clock=>clock,reset=>reset,s=>p(369)(77),cout=>p(370)(78));
FA_ff_15017:FAff port map(x=>p(358)(78),y=>p(359)(78),Cin=>p(360)(78),clock=>clock,reset=>reset,s=>p(369)(78),cout=>p(370)(79));
FA_ff_15018:FAff port map(x=>p(358)(79),y=>p(359)(79),Cin=>p(360)(79),clock=>clock,reset=>reset,s=>p(369)(79),cout=>p(370)(80));
FA_ff_15019:FAff port map(x=>p(358)(80),y=>p(359)(80),Cin=>p(360)(80),clock=>clock,reset=>reset,s=>p(369)(80),cout=>p(370)(81));
FA_ff_15020:FAff port map(x=>p(358)(81),y=>p(359)(81),Cin=>p(360)(81),clock=>clock,reset=>reset,s=>p(369)(81),cout=>p(370)(82));
FA_ff_15021:FAff port map(x=>p(358)(82),y=>p(359)(82),Cin=>p(360)(82),clock=>clock,reset=>reset,s=>p(369)(82),cout=>p(370)(83));
FA_ff_15022:FAff port map(x=>p(358)(83),y=>p(359)(83),Cin=>p(360)(83),clock=>clock,reset=>reset,s=>p(369)(83),cout=>p(370)(84));
FA_ff_15023:FAff port map(x=>p(358)(84),y=>p(359)(84),Cin=>p(360)(84),clock=>clock,reset=>reset,s=>p(369)(84),cout=>p(370)(85));
FA_ff_15024:FAff port map(x=>p(358)(85),y=>p(359)(85),Cin=>p(360)(85),clock=>clock,reset=>reset,s=>p(369)(85),cout=>p(370)(86));
FA_ff_15025:FAff port map(x=>p(358)(86),y=>p(359)(86),Cin=>p(360)(86),clock=>clock,reset=>reset,s=>p(369)(86),cout=>p(370)(87));
FA_ff_15026:FAff port map(x=>p(358)(87),y=>p(359)(87),Cin=>p(360)(87),clock=>clock,reset=>reset,s=>p(369)(87),cout=>p(370)(88));
FA_ff_15027:FAff port map(x=>p(358)(88),y=>p(359)(88),Cin=>p(360)(88),clock=>clock,reset=>reset,s=>p(369)(88),cout=>p(370)(89));
FA_ff_15028:FAff port map(x=>p(358)(89),y=>p(359)(89),Cin=>p(360)(89),clock=>clock,reset=>reset,s=>p(369)(89),cout=>p(370)(90));
FA_ff_15029:FAff port map(x=>p(358)(90),y=>p(359)(90),Cin=>p(360)(90),clock=>clock,reset=>reset,s=>p(369)(90),cout=>p(370)(91));
FA_ff_15030:FAff port map(x=>p(358)(91),y=>p(359)(91),Cin=>p(360)(91),clock=>clock,reset=>reset,s=>p(369)(91),cout=>p(370)(92));
FA_ff_15031:FAff port map(x=>p(358)(92),y=>p(359)(92),Cin=>p(360)(92),clock=>clock,reset=>reset,s=>p(369)(92),cout=>p(370)(93));
FA_ff_15032:FAff port map(x=>p(358)(93),y=>p(359)(93),Cin=>p(360)(93),clock=>clock,reset=>reset,s=>p(369)(93),cout=>p(370)(94));
FA_ff_15033:FAff port map(x=>p(358)(94),y=>p(359)(94),Cin=>p(360)(94),clock=>clock,reset=>reset,s=>p(369)(94),cout=>p(370)(95));
FA_ff_15034:FAff port map(x=>p(358)(95),y=>p(359)(95),Cin=>p(360)(95),clock=>clock,reset=>reset,s=>p(369)(95),cout=>p(370)(96));
FA_ff_15035:FAff port map(x=>p(358)(96),y=>p(359)(96),Cin=>p(360)(96),clock=>clock,reset=>reset,s=>p(369)(96),cout=>p(370)(97));
FA_ff_15036:FAff port map(x=>p(358)(97),y=>p(359)(97),Cin=>p(360)(97),clock=>clock,reset=>reset,s=>p(369)(97),cout=>p(370)(98));
FA_ff_15037:FAff port map(x=>p(358)(98),y=>p(359)(98),Cin=>p(360)(98),clock=>clock,reset=>reset,s=>p(369)(98),cout=>p(370)(99));
FA_ff_15038:FAff port map(x=>p(358)(99),y=>p(359)(99),Cin=>p(360)(99),clock=>clock,reset=>reset,s=>p(369)(99),cout=>p(370)(100));
FA_ff_15039:FAff port map(x=>p(358)(100),y=>p(359)(100),Cin=>p(360)(100),clock=>clock,reset=>reset,s=>p(369)(100),cout=>p(370)(101));
FA_ff_15040:FAff port map(x=>p(358)(101),y=>p(359)(101),Cin=>p(360)(101),clock=>clock,reset=>reset,s=>p(369)(101),cout=>p(370)(102));
FA_ff_15041:FAff port map(x=>p(358)(102),y=>p(359)(102),Cin=>p(360)(102),clock=>clock,reset=>reset,s=>p(369)(102),cout=>p(370)(103));
FA_ff_15042:FAff port map(x=>p(358)(103),y=>p(359)(103),Cin=>p(360)(103),clock=>clock,reset=>reset,s=>p(369)(103),cout=>p(370)(104));
FA_ff_15043:FAff port map(x=>p(358)(104),y=>p(359)(104),Cin=>p(360)(104),clock=>clock,reset=>reset,s=>p(369)(104),cout=>p(370)(105));
FA_ff_15044:FAff port map(x=>p(358)(105),y=>p(359)(105),Cin=>p(360)(105),clock=>clock,reset=>reset,s=>p(369)(105),cout=>p(370)(106));
FA_ff_15045:FAff port map(x=>p(358)(106),y=>p(359)(106),Cin=>p(360)(106),clock=>clock,reset=>reset,s=>p(369)(106),cout=>p(370)(107));
FA_ff_15046:FAff port map(x=>p(358)(107),y=>p(359)(107),Cin=>p(360)(107),clock=>clock,reset=>reset,s=>p(369)(107),cout=>p(370)(108));
FA_ff_15047:FAff port map(x=>p(358)(108),y=>p(359)(108),Cin=>p(360)(108),clock=>clock,reset=>reset,s=>p(369)(108),cout=>p(370)(109));
FA_ff_15048:FAff port map(x=>p(358)(109),y=>p(359)(109),Cin=>p(360)(109),clock=>clock,reset=>reset,s=>p(369)(109),cout=>p(370)(110));
FA_ff_15049:FAff port map(x=>p(358)(110),y=>p(359)(110),Cin=>p(360)(110),clock=>clock,reset=>reset,s=>p(369)(110),cout=>p(370)(111));
FA_ff_15050:FAff port map(x=>p(358)(111),y=>p(359)(111),Cin=>p(360)(111),clock=>clock,reset=>reset,s=>p(369)(111),cout=>p(370)(112));
FA_ff_15051:FAff port map(x=>p(358)(112),y=>p(359)(112),Cin=>p(360)(112),clock=>clock,reset=>reset,s=>p(369)(112),cout=>p(370)(113));
FA_ff_15052:FAff port map(x=>p(358)(113),y=>p(359)(113),Cin=>p(360)(113),clock=>clock,reset=>reset,s=>p(369)(113),cout=>p(370)(114));
FA_ff_15053:FAff port map(x=>p(358)(114),y=>p(359)(114),Cin=>p(360)(114),clock=>clock,reset=>reset,s=>p(369)(114),cout=>p(370)(115));
FA_ff_15054:FAff port map(x=>p(358)(115),y=>p(359)(115),Cin=>p(360)(115),clock=>clock,reset=>reset,s=>p(369)(115),cout=>p(370)(116));
FA_ff_15055:FAff port map(x=>p(358)(116),y=>p(359)(116),Cin=>p(360)(116),clock=>clock,reset=>reset,s=>p(369)(116),cout=>p(370)(117));
FA_ff_15056:FAff port map(x=>p(358)(117),y=>p(359)(117),Cin=>p(360)(117),clock=>clock,reset=>reset,s=>p(369)(117),cout=>p(370)(118));
FA_ff_15057:FAff port map(x=>p(358)(118),y=>p(359)(118),Cin=>p(360)(118),clock=>clock,reset=>reset,s=>p(369)(118),cout=>p(370)(119));
FA_ff_15058:FAff port map(x=>p(358)(119),y=>p(359)(119),Cin=>p(360)(119),clock=>clock,reset=>reset,s=>p(369)(119),cout=>p(370)(120));
FA_ff_15059:FAff port map(x=>p(358)(120),y=>p(359)(120),Cin=>p(360)(120),clock=>clock,reset=>reset,s=>p(369)(120),cout=>p(370)(121));
FA_ff_15060:FAff port map(x=>p(358)(121),y=>p(359)(121),Cin=>p(360)(121),clock=>clock,reset=>reset,s=>p(369)(121),cout=>p(370)(122));
FA_ff_15061:FAff port map(x=>p(358)(122),y=>p(359)(122),Cin=>p(360)(122),clock=>clock,reset=>reset,s=>p(369)(122),cout=>p(370)(123));
FA_ff_15062:FAff port map(x=>p(358)(123),y=>p(359)(123),Cin=>p(360)(123),clock=>clock,reset=>reset,s=>p(369)(123),cout=>p(370)(124));
FA_ff_15063:FAff port map(x=>p(358)(124),y=>p(359)(124),Cin=>p(360)(124),clock=>clock,reset=>reset,s=>p(369)(124),cout=>p(370)(125));
FA_ff_15064:FAff port map(x=>p(358)(125),y=>p(359)(125),Cin=>p(360)(125),clock=>clock,reset=>reset,s=>p(369)(125),cout=>p(370)(126));
FA_ff_15065:FAff port map(x=>p(358)(126),y=>p(359)(126),Cin=>p(360)(126),clock=>clock,reset=>reset,s=>p(369)(126),cout=>p(370)(127));
FA_ff_15066:FAff port map(x=>p(358)(127),y=>p(359)(127),Cin=>p(360)(127),clock=>clock,reset=>reset,s=>p(369)(127),cout=>p(370)(128));
FA_ff_15067:FAff port map(x=>p(358)(128),y=>p(359)(128),Cin=>p(360)(128),clock=>clock,reset=>reset,s=>p(369)(128),cout=>p(370)(129));
FA_ff_15068:FAff port map(x=>p(358)(129),y=>p(359)(129),Cin=>p(360)(129),clock=>clock,reset=>reset,s=>p(369)(129),cout=>p(370)(130));
FA_ff_15069:FAff port map(x=>p(358)(130),y=>p(359)(130),Cin=>p(360)(130),clock=>clock,reset=>reset,s=>p(369)(130),cout=>p(370)(131));
FA_ff_15070:FAff port map(x=>p(358)(131),y=>p(359)(131),Cin=>p(360)(131),clock=>clock,reset=>reset,s=>p(369)(131),cout=>p(370)(132));
HA_ff_101:HAff port map(x=>p(361)(0),y=>p(363)(0),clock=>clock,reset=>reset,s=>p(371)(0),c=>p(372)(1));
HA_ff_102:HAff port map(x=>p(361)(1),y=>p(363)(1),clock=>clock,reset=>reset,s=>p(371)(1),c=>p(372)(2));
FA_ff_15071:FAff port map(x=>p(361)(2),y=>p(362)(2),Cin=>p(363)(2),clock=>clock,reset=>reset,s=>p(371)(2),cout=>p(372)(3));
FA_ff_15072:FAff port map(x=>p(361)(3),y=>p(362)(3),Cin=>p(363)(3),clock=>clock,reset=>reset,s=>p(371)(3),cout=>p(372)(4));
FA_ff_15073:FAff port map(x=>p(361)(4),y=>p(362)(4),Cin=>p(363)(4),clock=>clock,reset=>reset,s=>p(371)(4),cout=>p(372)(5));
FA_ff_15074:FAff port map(x=>p(361)(5),y=>p(362)(5),Cin=>p(363)(5),clock=>clock,reset=>reset,s=>p(371)(5),cout=>p(372)(6));
FA_ff_15075:FAff port map(x=>p(361)(6),y=>p(362)(6),Cin=>p(363)(6),clock=>clock,reset=>reset,s=>p(371)(6),cout=>p(372)(7));
FA_ff_15076:FAff port map(x=>p(361)(7),y=>p(362)(7),Cin=>p(363)(7),clock=>clock,reset=>reset,s=>p(371)(7),cout=>p(372)(8));
FA_ff_15077:FAff port map(x=>p(361)(8),y=>p(362)(8),Cin=>p(363)(8),clock=>clock,reset=>reset,s=>p(371)(8),cout=>p(372)(9));
FA_ff_15078:FAff port map(x=>p(361)(9),y=>p(362)(9),Cin=>p(363)(9),clock=>clock,reset=>reset,s=>p(371)(9),cout=>p(372)(10));
FA_ff_15079:FAff port map(x=>p(361)(10),y=>p(362)(10),Cin=>p(363)(10),clock=>clock,reset=>reset,s=>p(371)(10),cout=>p(372)(11));
FA_ff_15080:FAff port map(x=>p(361)(11),y=>p(362)(11),Cin=>p(363)(11),clock=>clock,reset=>reset,s=>p(371)(11),cout=>p(372)(12));
FA_ff_15081:FAff port map(x=>p(361)(12),y=>p(362)(12),Cin=>p(363)(12),clock=>clock,reset=>reset,s=>p(371)(12),cout=>p(372)(13));
FA_ff_15082:FAff port map(x=>p(361)(13),y=>p(362)(13),Cin=>p(363)(13),clock=>clock,reset=>reset,s=>p(371)(13),cout=>p(372)(14));
FA_ff_15083:FAff port map(x=>p(361)(14),y=>p(362)(14),Cin=>p(363)(14),clock=>clock,reset=>reset,s=>p(371)(14),cout=>p(372)(15));
FA_ff_15084:FAff port map(x=>p(361)(15),y=>p(362)(15),Cin=>p(363)(15),clock=>clock,reset=>reset,s=>p(371)(15),cout=>p(372)(16));
FA_ff_15085:FAff port map(x=>p(361)(16),y=>p(362)(16),Cin=>p(363)(16),clock=>clock,reset=>reset,s=>p(371)(16),cout=>p(372)(17));
FA_ff_15086:FAff port map(x=>p(361)(17),y=>p(362)(17),Cin=>p(363)(17),clock=>clock,reset=>reset,s=>p(371)(17),cout=>p(372)(18));
FA_ff_15087:FAff port map(x=>p(361)(18),y=>p(362)(18),Cin=>p(363)(18),clock=>clock,reset=>reset,s=>p(371)(18),cout=>p(372)(19));
FA_ff_15088:FAff port map(x=>p(361)(19),y=>p(362)(19),Cin=>p(363)(19),clock=>clock,reset=>reset,s=>p(371)(19),cout=>p(372)(20));
FA_ff_15089:FAff port map(x=>p(361)(20),y=>p(362)(20),Cin=>p(363)(20),clock=>clock,reset=>reset,s=>p(371)(20),cout=>p(372)(21));
FA_ff_15090:FAff port map(x=>p(361)(21),y=>p(362)(21),Cin=>p(363)(21),clock=>clock,reset=>reset,s=>p(371)(21),cout=>p(372)(22));
FA_ff_15091:FAff port map(x=>p(361)(22),y=>p(362)(22),Cin=>p(363)(22),clock=>clock,reset=>reset,s=>p(371)(22),cout=>p(372)(23));
FA_ff_15092:FAff port map(x=>p(361)(23),y=>p(362)(23),Cin=>p(363)(23),clock=>clock,reset=>reset,s=>p(371)(23),cout=>p(372)(24));
FA_ff_15093:FAff port map(x=>p(361)(24),y=>p(362)(24),Cin=>p(363)(24),clock=>clock,reset=>reset,s=>p(371)(24),cout=>p(372)(25));
FA_ff_15094:FAff port map(x=>p(361)(25),y=>p(362)(25),Cin=>p(363)(25),clock=>clock,reset=>reset,s=>p(371)(25),cout=>p(372)(26));
FA_ff_15095:FAff port map(x=>p(361)(26),y=>p(362)(26),Cin=>p(363)(26),clock=>clock,reset=>reset,s=>p(371)(26),cout=>p(372)(27));
FA_ff_15096:FAff port map(x=>p(361)(27),y=>p(362)(27),Cin=>p(363)(27),clock=>clock,reset=>reset,s=>p(371)(27),cout=>p(372)(28));
FA_ff_15097:FAff port map(x=>p(361)(28),y=>p(362)(28),Cin=>p(363)(28),clock=>clock,reset=>reset,s=>p(371)(28),cout=>p(372)(29));
FA_ff_15098:FAff port map(x=>p(361)(29),y=>p(362)(29),Cin=>p(363)(29),clock=>clock,reset=>reset,s=>p(371)(29),cout=>p(372)(30));
FA_ff_15099:FAff port map(x=>p(361)(30),y=>p(362)(30),Cin=>p(363)(30),clock=>clock,reset=>reset,s=>p(371)(30),cout=>p(372)(31));
FA_ff_15100:FAff port map(x=>p(361)(31),y=>p(362)(31),Cin=>p(363)(31),clock=>clock,reset=>reset,s=>p(371)(31),cout=>p(372)(32));
FA_ff_15101:FAff port map(x=>p(361)(32),y=>p(362)(32),Cin=>p(363)(32),clock=>clock,reset=>reset,s=>p(371)(32),cout=>p(372)(33));
FA_ff_15102:FAff port map(x=>p(361)(33),y=>p(362)(33),Cin=>p(363)(33),clock=>clock,reset=>reset,s=>p(371)(33),cout=>p(372)(34));
FA_ff_15103:FAff port map(x=>p(361)(34),y=>p(362)(34),Cin=>p(363)(34),clock=>clock,reset=>reset,s=>p(371)(34),cout=>p(372)(35));
FA_ff_15104:FAff port map(x=>p(361)(35),y=>p(362)(35),Cin=>p(363)(35),clock=>clock,reset=>reset,s=>p(371)(35),cout=>p(372)(36));
FA_ff_15105:FAff port map(x=>p(361)(36),y=>p(362)(36),Cin=>p(363)(36),clock=>clock,reset=>reset,s=>p(371)(36),cout=>p(372)(37));
FA_ff_15106:FAff port map(x=>p(361)(37),y=>p(362)(37),Cin=>p(363)(37),clock=>clock,reset=>reset,s=>p(371)(37),cout=>p(372)(38));
FA_ff_15107:FAff port map(x=>p(361)(38),y=>p(362)(38),Cin=>p(363)(38),clock=>clock,reset=>reset,s=>p(371)(38),cout=>p(372)(39));
FA_ff_15108:FAff port map(x=>p(361)(39),y=>p(362)(39),Cin=>p(363)(39),clock=>clock,reset=>reset,s=>p(371)(39),cout=>p(372)(40));
FA_ff_15109:FAff port map(x=>p(361)(40),y=>p(362)(40),Cin=>p(363)(40),clock=>clock,reset=>reset,s=>p(371)(40),cout=>p(372)(41));
FA_ff_15110:FAff port map(x=>p(361)(41),y=>p(362)(41),Cin=>p(363)(41),clock=>clock,reset=>reset,s=>p(371)(41),cout=>p(372)(42));
FA_ff_15111:FAff port map(x=>p(361)(42),y=>p(362)(42),Cin=>p(363)(42),clock=>clock,reset=>reset,s=>p(371)(42),cout=>p(372)(43));
FA_ff_15112:FAff port map(x=>p(361)(43),y=>p(362)(43),Cin=>p(363)(43),clock=>clock,reset=>reset,s=>p(371)(43),cout=>p(372)(44));
FA_ff_15113:FAff port map(x=>p(361)(44),y=>p(362)(44),Cin=>p(363)(44),clock=>clock,reset=>reset,s=>p(371)(44),cout=>p(372)(45));
FA_ff_15114:FAff port map(x=>p(361)(45),y=>p(362)(45),Cin=>p(363)(45),clock=>clock,reset=>reset,s=>p(371)(45),cout=>p(372)(46));
FA_ff_15115:FAff port map(x=>p(361)(46),y=>p(362)(46),Cin=>p(363)(46),clock=>clock,reset=>reset,s=>p(371)(46),cout=>p(372)(47));
FA_ff_15116:FAff port map(x=>p(361)(47),y=>p(362)(47),Cin=>p(363)(47),clock=>clock,reset=>reset,s=>p(371)(47),cout=>p(372)(48));
FA_ff_15117:FAff port map(x=>p(361)(48),y=>p(362)(48),Cin=>p(363)(48),clock=>clock,reset=>reset,s=>p(371)(48),cout=>p(372)(49));
FA_ff_15118:FAff port map(x=>p(361)(49),y=>p(362)(49),Cin=>p(363)(49),clock=>clock,reset=>reset,s=>p(371)(49),cout=>p(372)(50));
FA_ff_15119:FAff port map(x=>p(361)(50),y=>p(362)(50),Cin=>p(363)(50),clock=>clock,reset=>reset,s=>p(371)(50),cout=>p(372)(51));
FA_ff_15120:FAff port map(x=>p(361)(51),y=>p(362)(51),Cin=>p(363)(51),clock=>clock,reset=>reset,s=>p(371)(51),cout=>p(372)(52));
FA_ff_15121:FAff port map(x=>p(361)(52),y=>p(362)(52),Cin=>p(363)(52),clock=>clock,reset=>reset,s=>p(371)(52),cout=>p(372)(53));
FA_ff_15122:FAff port map(x=>p(361)(53),y=>p(362)(53),Cin=>p(363)(53),clock=>clock,reset=>reset,s=>p(371)(53),cout=>p(372)(54));
FA_ff_15123:FAff port map(x=>p(361)(54),y=>p(362)(54),Cin=>p(363)(54),clock=>clock,reset=>reset,s=>p(371)(54),cout=>p(372)(55));
FA_ff_15124:FAff port map(x=>p(361)(55),y=>p(362)(55),Cin=>p(363)(55),clock=>clock,reset=>reset,s=>p(371)(55),cout=>p(372)(56));
FA_ff_15125:FAff port map(x=>p(361)(56),y=>p(362)(56),Cin=>p(363)(56),clock=>clock,reset=>reset,s=>p(371)(56),cout=>p(372)(57));
FA_ff_15126:FAff port map(x=>p(361)(57),y=>p(362)(57),Cin=>p(363)(57),clock=>clock,reset=>reset,s=>p(371)(57),cout=>p(372)(58));
FA_ff_15127:FAff port map(x=>p(361)(58),y=>p(362)(58),Cin=>p(363)(58),clock=>clock,reset=>reset,s=>p(371)(58),cout=>p(372)(59));
FA_ff_15128:FAff port map(x=>p(361)(59),y=>p(362)(59),Cin=>p(363)(59),clock=>clock,reset=>reset,s=>p(371)(59),cout=>p(372)(60));
FA_ff_15129:FAff port map(x=>p(361)(60),y=>p(362)(60),Cin=>p(363)(60),clock=>clock,reset=>reset,s=>p(371)(60),cout=>p(372)(61));
FA_ff_15130:FAff port map(x=>p(361)(61),y=>p(362)(61),Cin=>p(363)(61),clock=>clock,reset=>reset,s=>p(371)(61),cout=>p(372)(62));
FA_ff_15131:FAff port map(x=>p(361)(62),y=>p(362)(62),Cin=>p(363)(62),clock=>clock,reset=>reset,s=>p(371)(62),cout=>p(372)(63));
FA_ff_15132:FAff port map(x=>p(361)(63),y=>p(362)(63),Cin=>p(363)(63),clock=>clock,reset=>reset,s=>p(371)(63),cout=>p(372)(64));
FA_ff_15133:FAff port map(x=>p(361)(64),y=>p(362)(64),Cin=>p(363)(64),clock=>clock,reset=>reset,s=>p(371)(64),cout=>p(372)(65));
FA_ff_15134:FAff port map(x=>p(361)(65),y=>p(362)(65),Cin=>p(363)(65),clock=>clock,reset=>reset,s=>p(371)(65),cout=>p(372)(66));
FA_ff_15135:FAff port map(x=>p(361)(66),y=>p(362)(66),Cin=>p(363)(66),clock=>clock,reset=>reset,s=>p(371)(66),cout=>p(372)(67));
FA_ff_15136:FAff port map(x=>p(361)(67),y=>p(362)(67),Cin=>p(363)(67),clock=>clock,reset=>reset,s=>p(371)(67),cout=>p(372)(68));
FA_ff_15137:FAff port map(x=>p(361)(68),y=>p(362)(68),Cin=>p(363)(68),clock=>clock,reset=>reset,s=>p(371)(68),cout=>p(372)(69));
FA_ff_15138:FAff port map(x=>p(361)(69),y=>p(362)(69),Cin=>p(363)(69),clock=>clock,reset=>reset,s=>p(371)(69),cout=>p(372)(70));
FA_ff_15139:FAff port map(x=>p(361)(70),y=>p(362)(70),Cin=>p(363)(70),clock=>clock,reset=>reset,s=>p(371)(70),cout=>p(372)(71));
FA_ff_15140:FAff port map(x=>p(361)(71),y=>p(362)(71),Cin=>p(363)(71),clock=>clock,reset=>reset,s=>p(371)(71),cout=>p(372)(72));
FA_ff_15141:FAff port map(x=>p(361)(72),y=>p(362)(72),Cin=>p(363)(72),clock=>clock,reset=>reset,s=>p(371)(72),cout=>p(372)(73));
FA_ff_15142:FAff port map(x=>p(361)(73),y=>p(362)(73),Cin=>p(363)(73),clock=>clock,reset=>reset,s=>p(371)(73),cout=>p(372)(74));
FA_ff_15143:FAff port map(x=>p(361)(74),y=>p(362)(74),Cin=>p(363)(74),clock=>clock,reset=>reset,s=>p(371)(74),cout=>p(372)(75));
FA_ff_15144:FAff port map(x=>p(361)(75),y=>p(362)(75),Cin=>p(363)(75),clock=>clock,reset=>reset,s=>p(371)(75),cout=>p(372)(76));
FA_ff_15145:FAff port map(x=>p(361)(76),y=>p(362)(76),Cin=>p(363)(76),clock=>clock,reset=>reset,s=>p(371)(76),cout=>p(372)(77));
FA_ff_15146:FAff port map(x=>p(361)(77),y=>p(362)(77),Cin=>p(363)(77),clock=>clock,reset=>reset,s=>p(371)(77),cout=>p(372)(78));
FA_ff_15147:FAff port map(x=>p(361)(78),y=>p(362)(78),Cin=>p(363)(78),clock=>clock,reset=>reset,s=>p(371)(78),cout=>p(372)(79));
FA_ff_15148:FAff port map(x=>p(361)(79),y=>p(362)(79),Cin=>p(363)(79),clock=>clock,reset=>reset,s=>p(371)(79),cout=>p(372)(80));
FA_ff_15149:FAff port map(x=>p(361)(80),y=>p(362)(80),Cin=>p(363)(80),clock=>clock,reset=>reset,s=>p(371)(80),cout=>p(372)(81));
FA_ff_15150:FAff port map(x=>p(361)(81),y=>p(362)(81),Cin=>p(363)(81),clock=>clock,reset=>reset,s=>p(371)(81),cout=>p(372)(82));
FA_ff_15151:FAff port map(x=>p(361)(82),y=>p(362)(82),Cin=>p(363)(82),clock=>clock,reset=>reset,s=>p(371)(82),cout=>p(372)(83));
FA_ff_15152:FAff port map(x=>p(361)(83),y=>p(362)(83),Cin=>p(363)(83),clock=>clock,reset=>reset,s=>p(371)(83),cout=>p(372)(84));
FA_ff_15153:FAff port map(x=>p(361)(84),y=>p(362)(84),Cin=>p(363)(84),clock=>clock,reset=>reset,s=>p(371)(84),cout=>p(372)(85));
FA_ff_15154:FAff port map(x=>p(361)(85),y=>p(362)(85),Cin=>p(363)(85),clock=>clock,reset=>reset,s=>p(371)(85),cout=>p(372)(86));
FA_ff_15155:FAff port map(x=>p(361)(86),y=>p(362)(86),Cin=>p(363)(86),clock=>clock,reset=>reset,s=>p(371)(86),cout=>p(372)(87));
FA_ff_15156:FAff port map(x=>p(361)(87),y=>p(362)(87),Cin=>p(363)(87),clock=>clock,reset=>reset,s=>p(371)(87),cout=>p(372)(88));
FA_ff_15157:FAff port map(x=>p(361)(88),y=>p(362)(88),Cin=>p(363)(88),clock=>clock,reset=>reset,s=>p(371)(88),cout=>p(372)(89));
FA_ff_15158:FAff port map(x=>p(361)(89),y=>p(362)(89),Cin=>p(363)(89),clock=>clock,reset=>reset,s=>p(371)(89),cout=>p(372)(90));
FA_ff_15159:FAff port map(x=>p(361)(90),y=>p(362)(90),Cin=>p(363)(90),clock=>clock,reset=>reset,s=>p(371)(90),cout=>p(372)(91));
FA_ff_15160:FAff port map(x=>p(361)(91),y=>p(362)(91),Cin=>p(363)(91),clock=>clock,reset=>reset,s=>p(371)(91),cout=>p(372)(92));
FA_ff_15161:FAff port map(x=>p(361)(92),y=>p(362)(92),Cin=>p(363)(92),clock=>clock,reset=>reset,s=>p(371)(92),cout=>p(372)(93));
FA_ff_15162:FAff port map(x=>p(361)(93),y=>p(362)(93),Cin=>p(363)(93),clock=>clock,reset=>reset,s=>p(371)(93),cout=>p(372)(94));
FA_ff_15163:FAff port map(x=>p(361)(94),y=>p(362)(94),Cin=>p(363)(94),clock=>clock,reset=>reset,s=>p(371)(94),cout=>p(372)(95));
FA_ff_15164:FAff port map(x=>p(361)(95),y=>p(362)(95),Cin=>p(363)(95),clock=>clock,reset=>reset,s=>p(371)(95),cout=>p(372)(96));
FA_ff_15165:FAff port map(x=>p(361)(96),y=>p(362)(96),Cin=>p(363)(96),clock=>clock,reset=>reset,s=>p(371)(96),cout=>p(372)(97));
FA_ff_15166:FAff port map(x=>p(361)(97),y=>p(362)(97),Cin=>p(363)(97),clock=>clock,reset=>reset,s=>p(371)(97),cout=>p(372)(98));
FA_ff_15167:FAff port map(x=>p(361)(98),y=>p(362)(98),Cin=>p(363)(98),clock=>clock,reset=>reset,s=>p(371)(98),cout=>p(372)(99));
FA_ff_15168:FAff port map(x=>p(361)(99),y=>p(362)(99),Cin=>p(363)(99),clock=>clock,reset=>reset,s=>p(371)(99),cout=>p(372)(100));
FA_ff_15169:FAff port map(x=>p(361)(100),y=>p(362)(100),Cin=>p(363)(100),clock=>clock,reset=>reset,s=>p(371)(100),cout=>p(372)(101));
FA_ff_15170:FAff port map(x=>p(361)(101),y=>p(362)(101),Cin=>p(363)(101),clock=>clock,reset=>reset,s=>p(371)(101),cout=>p(372)(102));
FA_ff_15171:FAff port map(x=>p(361)(102),y=>p(362)(102),Cin=>p(363)(102),clock=>clock,reset=>reset,s=>p(371)(102),cout=>p(372)(103));
FA_ff_15172:FAff port map(x=>p(361)(103),y=>p(362)(103),Cin=>p(363)(103),clock=>clock,reset=>reset,s=>p(371)(103),cout=>p(372)(104));
FA_ff_15173:FAff port map(x=>p(361)(104),y=>p(362)(104),Cin=>p(363)(104),clock=>clock,reset=>reset,s=>p(371)(104),cout=>p(372)(105));
FA_ff_15174:FAff port map(x=>p(361)(105),y=>p(362)(105),Cin=>p(363)(105),clock=>clock,reset=>reset,s=>p(371)(105),cout=>p(372)(106));
FA_ff_15175:FAff port map(x=>p(361)(106),y=>p(362)(106),Cin=>p(363)(106),clock=>clock,reset=>reset,s=>p(371)(106),cout=>p(372)(107));
FA_ff_15176:FAff port map(x=>p(361)(107),y=>p(362)(107),Cin=>p(363)(107),clock=>clock,reset=>reset,s=>p(371)(107),cout=>p(372)(108));
FA_ff_15177:FAff port map(x=>p(361)(108),y=>p(362)(108),Cin=>p(363)(108),clock=>clock,reset=>reset,s=>p(371)(108),cout=>p(372)(109));
FA_ff_15178:FAff port map(x=>p(361)(109),y=>p(362)(109),Cin=>p(363)(109),clock=>clock,reset=>reset,s=>p(371)(109),cout=>p(372)(110));
FA_ff_15179:FAff port map(x=>p(361)(110),y=>p(362)(110),Cin=>p(363)(110),clock=>clock,reset=>reset,s=>p(371)(110),cout=>p(372)(111));
FA_ff_15180:FAff port map(x=>p(361)(111),y=>p(362)(111),Cin=>p(363)(111),clock=>clock,reset=>reset,s=>p(371)(111),cout=>p(372)(112));
FA_ff_15181:FAff port map(x=>p(361)(112),y=>p(362)(112),Cin=>p(363)(112),clock=>clock,reset=>reset,s=>p(371)(112),cout=>p(372)(113));
FA_ff_15182:FAff port map(x=>p(361)(113),y=>p(362)(113),Cin=>p(363)(113),clock=>clock,reset=>reset,s=>p(371)(113),cout=>p(372)(114));
FA_ff_15183:FAff port map(x=>p(361)(114),y=>p(362)(114),Cin=>p(363)(114),clock=>clock,reset=>reset,s=>p(371)(114),cout=>p(372)(115));
FA_ff_15184:FAff port map(x=>p(361)(115),y=>p(362)(115),Cin=>p(363)(115),clock=>clock,reset=>reset,s=>p(371)(115),cout=>p(372)(116));
FA_ff_15185:FAff port map(x=>p(361)(116),y=>p(362)(116),Cin=>p(363)(116),clock=>clock,reset=>reset,s=>p(371)(116),cout=>p(372)(117));
FA_ff_15186:FAff port map(x=>p(361)(117),y=>p(362)(117),Cin=>p(363)(117),clock=>clock,reset=>reset,s=>p(371)(117),cout=>p(372)(118));
FA_ff_15187:FAff port map(x=>p(361)(118),y=>p(362)(118),Cin=>p(363)(118),clock=>clock,reset=>reset,s=>p(371)(118),cout=>p(372)(119));
FA_ff_15188:FAff port map(x=>p(361)(119),y=>p(362)(119),Cin=>p(363)(119),clock=>clock,reset=>reset,s=>p(371)(119),cout=>p(372)(120));
FA_ff_15189:FAff port map(x=>p(361)(120),y=>p(362)(120),Cin=>p(363)(120),clock=>clock,reset=>reset,s=>p(371)(120),cout=>p(372)(121));
FA_ff_15190:FAff port map(x=>p(361)(121),y=>p(362)(121),Cin=>p(363)(121),clock=>clock,reset=>reset,s=>p(371)(121),cout=>p(372)(122));
FA_ff_15191:FAff port map(x=>p(361)(122),y=>p(362)(122),Cin=>p(363)(122),clock=>clock,reset=>reset,s=>p(371)(122),cout=>p(372)(123));
FA_ff_15192:FAff port map(x=>p(361)(123),y=>p(362)(123),Cin=>p(363)(123),clock=>clock,reset=>reset,s=>p(371)(123),cout=>p(372)(124));
FA_ff_15193:FAff port map(x=>p(361)(124),y=>p(362)(124),Cin=>p(363)(124),clock=>clock,reset=>reset,s=>p(371)(124),cout=>p(372)(125));
FA_ff_15194:FAff port map(x=>p(361)(125),y=>p(362)(125),Cin=>p(363)(125),clock=>clock,reset=>reset,s=>p(371)(125),cout=>p(372)(126));
FA_ff_15195:FAff port map(x=>p(361)(126),y=>p(362)(126),Cin=>p(363)(126),clock=>clock,reset=>reset,s=>p(371)(126),cout=>p(372)(127));
FA_ff_15196:FAff port map(x=>p(361)(127),y=>p(362)(127),Cin=>p(363)(127),clock=>clock,reset=>reset,s=>p(371)(127),cout=>p(372)(128));
FA_ff_15197:FAff port map(x=>p(361)(128),y=>p(362)(128),Cin=>p(363)(128),clock=>clock,reset=>reset,s=>p(371)(128),cout=>p(372)(129));
FA_ff_15198:FAff port map(x=>p(361)(129),y=>p(362)(129),Cin=>p(363)(129),clock=>clock,reset=>reset,s=>p(371)(129),cout=>p(372)(130));
FA_ff_15199:FAff port map(x=>p(361)(130),y=>p(362)(130),Cin=>p(363)(130),clock=>clock,reset=>reset,s=>p(371)(130),cout=>p(372)(131));
HA_ff_103:HAff port map(x=>p(361)(131),y=>p(362)(131),clock=>clock,reset=>reset,s=>p(371)(131),c=>p(372)(132));
p(373)(0)<=p(365)(0);
HA_ff_104:HAff port map(x=>p(364)(1),y=>p(365)(1),clock=>clock,reset=>reset,s=>p(373)(1),c=>p(374)(2));
FA_ff_15200:FAff port map(x=>p(364)(2),y=>p(365)(2),Cin=>p(366)(2),clock=>clock,reset=>reset,s=>p(373)(2),cout=>p(374)(3));
FA_ff_15201:FAff port map(x=>p(364)(3),y=>p(365)(3),Cin=>p(366)(3),clock=>clock,reset=>reset,s=>p(373)(3),cout=>p(374)(4));
FA_ff_15202:FAff port map(x=>p(364)(4),y=>p(365)(4),Cin=>p(366)(4),clock=>clock,reset=>reset,s=>p(373)(4),cout=>p(374)(5));
FA_ff_15203:FAff port map(x=>p(364)(5),y=>p(365)(5),Cin=>p(366)(5),clock=>clock,reset=>reset,s=>p(373)(5),cout=>p(374)(6));
FA_ff_15204:FAff port map(x=>p(364)(6),y=>p(365)(6),Cin=>p(366)(6),clock=>clock,reset=>reset,s=>p(373)(6),cout=>p(374)(7));
FA_ff_15205:FAff port map(x=>p(364)(7),y=>p(365)(7),Cin=>p(366)(7),clock=>clock,reset=>reset,s=>p(373)(7),cout=>p(374)(8));
FA_ff_15206:FAff port map(x=>p(364)(8),y=>p(365)(8),Cin=>p(366)(8),clock=>clock,reset=>reset,s=>p(373)(8),cout=>p(374)(9));
FA_ff_15207:FAff port map(x=>p(364)(9),y=>p(365)(9),Cin=>p(366)(9),clock=>clock,reset=>reset,s=>p(373)(9),cout=>p(374)(10));
FA_ff_15208:FAff port map(x=>p(364)(10),y=>p(365)(10),Cin=>p(366)(10),clock=>clock,reset=>reset,s=>p(373)(10),cout=>p(374)(11));
FA_ff_15209:FAff port map(x=>p(364)(11),y=>p(365)(11),Cin=>p(366)(11),clock=>clock,reset=>reset,s=>p(373)(11),cout=>p(374)(12));
FA_ff_15210:FAff port map(x=>p(364)(12),y=>p(365)(12),Cin=>p(366)(12),clock=>clock,reset=>reset,s=>p(373)(12),cout=>p(374)(13));
FA_ff_15211:FAff port map(x=>p(364)(13),y=>p(365)(13),Cin=>p(366)(13),clock=>clock,reset=>reset,s=>p(373)(13),cout=>p(374)(14));
FA_ff_15212:FAff port map(x=>p(364)(14),y=>p(365)(14),Cin=>p(366)(14),clock=>clock,reset=>reset,s=>p(373)(14),cout=>p(374)(15));
FA_ff_15213:FAff port map(x=>p(364)(15),y=>p(365)(15),Cin=>p(366)(15),clock=>clock,reset=>reset,s=>p(373)(15),cout=>p(374)(16));
FA_ff_15214:FAff port map(x=>p(364)(16),y=>p(365)(16),Cin=>p(366)(16),clock=>clock,reset=>reset,s=>p(373)(16),cout=>p(374)(17));
FA_ff_15215:FAff port map(x=>p(364)(17),y=>p(365)(17),Cin=>p(366)(17),clock=>clock,reset=>reset,s=>p(373)(17),cout=>p(374)(18));
FA_ff_15216:FAff port map(x=>p(364)(18),y=>p(365)(18),Cin=>p(366)(18),clock=>clock,reset=>reset,s=>p(373)(18),cout=>p(374)(19));
FA_ff_15217:FAff port map(x=>p(364)(19),y=>p(365)(19),Cin=>p(366)(19),clock=>clock,reset=>reset,s=>p(373)(19),cout=>p(374)(20));
FA_ff_15218:FAff port map(x=>p(364)(20),y=>p(365)(20),Cin=>p(366)(20),clock=>clock,reset=>reset,s=>p(373)(20),cout=>p(374)(21));
FA_ff_15219:FAff port map(x=>p(364)(21),y=>p(365)(21),Cin=>p(366)(21),clock=>clock,reset=>reset,s=>p(373)(21),cout=>p(374)(22));
FA_ff_15220:FAff port map(x=>p(364)(22),y=>p(365)(22),Cin=>p(366)(22),clock=>clock,reset=>reset,s=>p(373)(22),cout=>p(374)(23));
FA_ff_15221:FAff port map(x=>p(364)(23),y=>p(365)(23),Cin=>p(366)(23),clock=>clock,reset=>reset,s=>p(373)(23),cout=>p(374)(24));
FA_ff_15222:FAff port map(x=>p(364)(24),y=>p(365)(24),Cin=>p(366)(24),clock=>clock,reset=>reset,s=>p(373)(24),cout=>p(374)(25));
FA_ff_15223:FAff port map(x=>p(364)(25),y=>p(365)(25),Cin=>p(366)(25),clock=>clock,reset=>reset,s=>p(373)(25),cout=>p(374)(26));
FA_ff_15224:FAff port map(x=>p(364)(26),y=>p(365)(26),Cin=>p(366)(26),clock=>clock,reset=>reset,s=>p(373)(26),cout=>p(374)(27));
FA_ff_15225:FAff port map(x=>p(364)(27),y=>p(365)(27),Cin=>p(366)(27),clock=>clock,reset=>reset,s=>p(373)(27),cout=>p(374)(28));
FA_ff_15226:FAff port map(x=>p(364)(28),y=>p(365)(28),Cin=>p(366)(28),clock=>clock,reset=>reset,s=>p(373)(28),cout=>p(374)(29));
FA_ff_15227:FAff port map(x=>p(364)(29),y=>p(365)(29),Cin=>p(366)(29),clock=>clock,reset=>reset,s=>p(373)(29),cout=>p(374)(30));
FA_ff_15228:FAff port map(x=>p(364)(30),y=>p(365)(30),Cin=>p(366)(30),clock=>clock,reset=>reset,s=>p(373)(30),cout=>p(374)(31));
FA_ff_15229:FAff port map(x=>p(364)(31),y=>p(365)(31),Cin=>p(366)(31),clock=>clock,reset=>reset,s=>p(373)(31),cout=>p(374)(32));
FA_ff_15230:FAff port map(x=>p(364)(32),y=>p(365)(32),Cin=>p(366)(32),clock=>clock,reset=>reset,s=>p(373)(32),cout=>p(374)(33));
FA_ff_15231:FAff port map(x=>p(364)(33),y=>p(365)(33),Cin=>p(366)(33),clock=>clock,reset=>reset,s=>p(373)(33),cout=>p(374)(34));
FA_ff_15232:FAff port map(x=>p(364)(34),y=>p(365)(34),Cin=>p(366)(34),clock=>clock,reset=>reset,s=>p(373)(34),cout=>p(374)(35));
FA_ff_15233:FAff port map(x=>p(364)(35),y=>p(365)(35),Cin=>p(366)(35),clock=>clock,reset=>reset,s=>p(373)(35),cout=>p(374)(36));
FA_ff_15234:FAff port map(x=>p(364)(36),y=>p(365)(36),Cin=>p(366)(36),clock=>clock,reset=>reset,s=>p(373)(36),cout=>p(374)(37));
FA_ff_15235:FAff port map(x=>p(364)(37),y=>p(365)(37),Cin=>p(366)(37),clock=>clock,reset=>reset,s=>p(373)(37),cout=>p(374)(38));
FA_ff_15236:FAff port map(x=>p(364)(38),y=>p(365)(38),Cin=>p(366)(38),clock=>clock,reset=>reset,s=>p(373)(38),cout=>p(374)(39));
FA_ff_15237:FAff port map(x=>p(364)(39),y=>p(365)(39),Cin=>p(366)(39),clock=>clock,reset=>reset,s=>p(373)(39),cout=>p(374)(40));
FA_ff_15238:FAff port map(x=>p(364)(40),y=>p(365)(40),Cin=>p(366)(40),clock=>clock,reset=>reset,s=>p(373)(40),cout=>p(374)(41));
FA_ff_15239:FAff port map(x=>p(364)(41),y=>p(365)(41),Cin=>p(366)(41),clock=>clock,reset=>reset,s=>p(373)(41),cout=>p(374)(42));
FA_ff_15240:FAff port map(x=>p(364)(42),y=>p(365)(42),Cin=>p(366)(42),clock=>clock,reset=>reset,s=>p(373)(42),cout=>p(374)(43));
FA_ff_15241:FAff port map(x=>p(364)(43),y=>p(365)(43),Cin=>p(366)(43),clock=>clock,reset=>reset,s=>p(373)(43),cout=>p(374)(44));
FA_ff_15242:FAff port map(x=>p(364)(44),y=>p(365)(44),Cin=>p(366)(44),clock=>clock,reset=>reset,s=>p(373)(44),cout=>p(374)(45));
FA_ff_15243:FAff port map(x=>p(364)(45),y=>p(365)(45),Cin=>p(366)(45),clock=>clock,reset=>reset,s=>p(373)(45),cout=>p(374)(46));
FA_ff_15244:FAff port map(x=>p(364)(46),y=>p(365)(46),Cin=>p(366)(46),clock=>clock,reset=>reset,s=>p(373)(46),cout=>p(374)(47));
FA_ff_15245:FAff port map(x=>p(364)(47),y=>p(365)(47),Cin=>p(366)(47),clock=>clock,reset=>reset,s=>p(373)(47),cout=>p(374)(48));
FA_ff_15246:FAff port map(x=>p(364)(48),y=>p(365)(48),Cin=>p(366)(48),clock=>clock,reset=>reset,s=>p(373)(48),cout=>p(374)(49));
FA_ff_15247:FAff port map(x=>p(364)(49),y=>p(365)(49),Cin=>p(366)(49),clock=>clock,reset=>reset,s=>p(373)(49),cout=>p(374)(50));
FA_ff_15248:FAff port map(x=>p(364)(50),y=>p(365)(50),Cin=>p(366)(50),clock=>clock,reset=>reset,s=>p(373)(50),cout=>p(374)(51));
FA_ff_15249:FAff port map(x=>p(364)(51),y=>p(365)(51),Cin=>p(366)(51),clock=>clock,reset=>reset,s=>p(373)(51),cout=>p(374)(52));
FA_ff_15250:FAff port map(x=>p(364)(52),y=>p(365)(52),Cin=>p(366)(52),clock=>clock,reset=>reset,s=>p(373)(52),cout=>p(374)(53));
FA_ff_15251:FAff port map(x=>p(364)(53),y=>p(365)(53),Cin=>p(366)(53),clock=>clock,reset=>reset,s=>p(373)(53),cout=>p(374)(54));
FA_ff_15252:FAff port map(x=>p(364)(54),y=>p(365)(54),Cin=>p(366)(54),clock=>clock,reset=>reset,s=>p(373)(54),cout=>p(374)(55));
FA_ff_15253:FAff port map(x=>p(364)(55),y=>p(365)(55),Cin=>p(366)(55),clock=>clock,reset=>reset,s=>p(373)(55),cout=>p(374)(56));
FA_ff_15254:FAff port map(x=>p(364)(56),y=>p(365)(56),Cin=>p(366)(56),clock=>clock,reset=>reset,s=>p(373)(56),cout=>p(374)(57));
FA_ff_15255:FAff port map(x=>p(364)(57),y=>p(365)(57),Cin=>p(366)(57),clock=>clock,reset=>reset,s=>p(373)(57),cout=>p(374)(58));
FA_ff_15256:FAff port map(x=>p(364)(58),y=>p(365)(58),Cin=>p(366)(58),clock=>clock,reset=>reset,s=>p(373)(58),cout=>p(374)(59));
FA_ff_15257:FAff port map(x=>p(364)(59),y=>p(365)(59),Cin=>p(366)(59),clock=>clock,reset=>reset,s=>p(373)(59),cout=>p(374)(60));
FA_ff_15258:FAff port map(x=>p(364)(60),y=>p(365)(60),Cin=>p(366)(60),clock=>clock,reset=>reset,s=>p(373)(60),cout=>p(374)(61));
FA_ff_15259:FAff port map(x=>p(364)(61),y=>p(365)(61),Cin=>p(366)(61),clock=>clock,reset=>reset,s=>p(373)(61),cout=>p(374)(62));
FA_ff_15260:FAff port map(x=>p(364)(62),y=>p(365)(62),Cin=>p(366)(62),clock=>clock,reset=>reset,s=>p(373)(62),cout=>p(374)(63));
FA_ff_15261:FAff port map(x=>p(364)(63),y=>p(365)(63),Cin=>p(366)(63),clock=>clock,reset=>reset,s=>p(373)(63),cout=>p(374)(64));
FA_ff_15262:FAff port map(x=>p(364)(64),y=>p(365)(64),Cin=>p(366)(64),clock=>clock,reset=>reset,s=>p(373)(64),cout=>p(374)(65));
FA_ff_15263:FAff port map(x=>p(364)(65),y=>p(365)(65),Cin=>p(366)(65),clock=>clock,reset=>reset,s=>p(373)(65),cout=>p(374)(66));
FA_ff_15264:FAff port map(x=>p(364)(66),y=>p(365)(66),Cin=>p(366)(66),clock=>clock,reset=>reset,s=>p(373)(66),cout=>p(374)(67));
FA_ff_15265:FAff port map(x=>p(364)(67),y=>p(365)(67),Cin=>p(366)(67),clock=>clock,reset=>reset,s=>p(373)(67),cout=>p(374)(68));
FA_ff_15266:FAff port map(x=>p(364)(68),y=>p(365)(68),Cin=>p(366)(68),clock=>clock,reset=>reset,s=>p(373)(68),cout=>p(374)(69));
FA_ff_15267:FAff port map(x=>p(364)(69),y=>p(365)(69),Cin=>p(366)(69),clock=>clock,reset=>reset,s=>p(373)(69),cout=>p(374)(70));
FA_ff_15268:FAff port map(x=>p(364)(70),y=>p(365)(70),Cin=>p(366)(70),clock=>clock,reset=>reset,s=>p(373)(70),cout=>p(374)(71));
FA_ff_15269:FAff port map(x=>p(364)(71),y=>p(365)(71),Cin=>p(366)(71),clock=>clock,reset=>reset,s=>p(373)(71),cout=>p(374)(72));
FA_ff_15270:FAff port map(x=>p(364)(72),y=>p(365)(72),Cin=>p(366)(72),clock=>clock,reset=>reset,s=>p(373)(72),cout=>p(374)(73));
FA_ff_15271:FAff port map(x=>p(364)(73),y=>p(365)(73),Cin=>p(366)(73),clock=>clock,reset=>reset,s=>p(373)(73),cout=>p(374)(74));
FA_ff_15272:FAff port map(x=>p(364)(74),y=>p(365)(74),Cin=>p(366)(74),clock=>clock,reset=>reset,s=>p(373)(74),cout=>p(374)(75));
FA_ff_15273:FAff port map(x=>p(364)(75),y=>p(365)(75),Cin=>p(366)(75),clock=>clock,reset=>reset,s=>p(373)(75),cout=>p(374)(76));
FA_ff_15274:FAff port map(x=>p(364)(76),y=>p(365)(76),Cin=>p(366)(76),clock=>clock,reset=>reset,s=>p(373)(76),cout=>p(374)(77));
FA_ff_15275:FAff port map(x=>p(364)(77),y=>p(365)(77),Cin=>p(366)(77),clock=>clock,reset=>reset,s=>p(373)(77),cout=>p(374)(78));
FA_ff_15276:FAff port map(x=>p(364)(78),y=>p(365)(78),Cin=>p(366)(78),clock=>clock,reset=>reset,s=>p(373)(78),cout=>p(374)(79));
FA_ff_15277:FAff port map(x=>p(364)(79),y=>p(365)(79),Cin=>p(366)(79),clock=>clock,reset=>reset,s=>p(373)(79),cout=>p(374)(80));
FA_ff_15278:FAff port map(x=>p(364)(80),y=>p(365)(80),Cin=>p(366)(80),clock=>clock,reset=>reset,s=>p(373)(80),cout=>p(374)(81));
FA_ff_15279:FAff port map(x=>p(364)(81),y=>p(365)(81),Cin=>p(366)(81),clock=>clock,reset=>reset,s=>p(373)(81),cout=>p(374)(82));
FA_ff_15280:FAff port map(x=>p(364)(82),y=>p(365)(82),Cin=>p(366)(82),clock=>clock,reset=>reset,s=>p(373)(82),cout=>p(374)(83));
FA_ff_15281:FAff port map(x=>p(364)(83),y=>p(365)(83),Cin=>p(366)(83),clock=>clock,reset=>reset,s=>p(373)(83),cout=>p(374)(84));
FA_ff_15282:FAff port map(x=>p(364)(84),y=>p(365)(84),Cin=>p(366)(84),clock=>clock,reset=>reset,s=>p(373)(84),cout=>p(374)(85));
FA_ff_15283:FAff port map(x=>p(364)(85),y=>p(365)(85),Cin=>p(366)(85),clock=>clock,reset=>reset,s=>p(373)(85),cout=>p(374)(86));
FA_ff_15284:FAff port map(x=>p(364)(86),y=>p(365)(86),Cin=>p(366)(86),clock=>clock,reset=>reset,s=>p(373)(86),cout=>p(374)(87));
FA_ff_15285:FAff port map(x=>p(364)(87),y=>p(365)(87),Cin=>p(366)(87),clock=>clock,reset=>reset,s=>p(373)(87),cout=>p(374)(88));
FA_ff_15286:FAff port map(x=>p(364)(88),y=>p(365)(88),Cin=>p(366)(88),clock=>clock,reset=>reset,s=>p(373)(88),cout=>p(374)(89));
FA_ff_15287:FAff port map(x=>p(364)(89),y=>p(365)(89),Cin=>p(366)(89),clock=>clock,reset=>reset,s=>p(373)(89),cout=>p(374)(90));
FA_ff_15288:FAff port map(x=>p(364)(90),y=>p(365)(90),Cin=>p(366)(90),clock=>clock,reset=>reset,s=>p(373)(90),cout=>p(374)(91));
FA_ff_15289:FAff port map(x=>p(364)(91),y=>p(365)(91),Cin=>p(366)(91),clock=>clock,reset=>reset,s=>p(373)(91),cout=>p(374)(92));
FA_ff_15290:FAff port map(x=>p(364)(92),y=>p(365)(92),Cin=>p(366)(92),clock=>clock,reset=>reset,s=>p(373)(92),cout=>p(374)(93));
FA_ff_15291:FAff port map(x=>p(364)(93),y=>p(365)(93),Cin=>p(366)(93),clock=>clock,reset=>reset,s=>p(373)(93),cout=>p(374)(94));
FA_ff_15292:FAff port map(x=>p(364)(94),y=>p(365)(94),Cin=>p(366)(94),clock=>clock,reset=>reset,s=>p(373)(94),cout=>p(374)(95));
FA_ff_15293:FAff port map(x=>p(364)(95),y=>p(365)(95),Cin=>p(366)(95),clock=>clock,reset=>reset,s=>p(373)(95),cout=>p(374)(96));
FA_ff_15294:FAff port map(x=>p(364)(96),y=>p(365)(96),Cin=>p(366)(96),clock=>clock,reset=>reset,s=>p(373)(96),cout=>p(374)(97));
FA_ff_15295:FAff port map(x=>p(364)(97),y=>p(365)(97),Cin=>p(366)(97),clock=>clock,reset=>reset,s=>p(373)(97),cout=>p(374)(98));
FA_ff_15296:FAff port map(x=>p(364)(98),y=>p(365)(98),Cin=>p(366)(98),clock=>clock,reset=>reset,s=>p(373)(98),cout=>p(374)(99));
FA_ff_15297:FAff port map(x=>p(364)(99),y=>p(365)(99),Cin=>p(366)(99),clock=>clock,reset=>reset,s=>p(373)(99),cout=>p(374)(100));
FA_ff_15298:FAff port map(x=>p(364)(100),y=>p(365)(100),Cin=>p(366)(100),clock=>clock,reset=>reset,s=>p(373)(100),cout=>p(374)(101));
FA_ff_15299:FAff port map(x=>p(364)(101),y=>p(365)(101),Cin=>p(366)(101),clock=>clock,reset=>reset,s=>p(373)(101),cout=>p(374)(102));
FA_ff_15300:FAff port map(x=>p(364)(102),y=>p(365)(102),Cin=>p(366)(102),clock=>clock,reset=>reset,s=>p(373)(102),cout=>p(374)(103));
FA_ff_15301:FAff port map(x=>p(364)(103),y=>p(365)(103),Cin=>p(366)(103),clock=>clock,reset=>reset,s=>p(373)(103),cout=>p(374)(104));
FA_ff_15302:FAff port map(x=>p(364)(104),y=>p(365)(104),Cin=>p(366)(104),clock=>clock,reset=>reset,s=>p(373)(104),cout=>p(374)(105));
FA_ff_15303:FAff port map(x=>p(364)(105),y=>p(365)(105),Cin=>p(366)(105),clock=>clock,reset=>reset,s=>p(373)(105),cout=>p(374)(106));
FA_ff_15304:FAff port map(x=>p(364)(106),y=>p(365)(106),Cin=>p(366)(106),clock=>clock,reset=>reset,s=>p(373)(106),cout=>p(374)(107));
FA_ff_15305:FAff port map(x=>p(364)(107),y=>p(365)(107),Cin=>p(366)(107),clock=>clock,reset=>reset,s=>p(373)(107),cout=>p(374)(108));
FA_ff_15306:FAff port map(x=>p(364)(108),y=>p(365)(108),Cin=>p(366)(108),clock=>clock,reset=>reset,s=>p(373)(108),cout=>p(374)(109));
FA_ff_15307:FAff port map(x=>p(364)(109),y=>p(365)(109),Cin=>p(366)(109),clock=>clock,reset=>reset,s=>p(373)(109),cout=>p(374)(110));
FA_ff_15308:FAff port map(x=>p(364)(110),y=>p(365)(110),Cin=>p(366)(110),clock=>clock,reset=>reset,s=>p(373)(110),cout=>p(374)(111));
FA_ff_15309:FAff port map(x=>p(364)(111),y=>p(365)(111),Cin=>p(366)(111),clock=>clock,reset=>reset,s=>p(373)(111),cout=>p(374)(112));
FA_ff_15310:FAff port map(x=>p(364)(112),y=>p(365)(112),Cin=>p(366)(112),clock=>clock,reset=>reset,s=>p(373)(112),cout=>p(374)(113));
FA_ff_15311:FAff port map(x=>p(364)(113),y=>p(365)(113),Cin=>p(366)(113),clock=>clock,reset=>reset,s=>p(373)(113),cout=>p(374)(114));
FA_ff_15312:FAff port map(x=>p(364)(114),y=>p(365)(114),Cin=>p(366)(114),clock=>clock,reset=>reset,s=>p(373)(114),cout=>p(374)(115));
FA_ff_15313:FAff port map(x=>p(364)(115),y=>p(365)(115),Cin=>p(366)(115),clock=>clock,reset=>reset,s=>p(373)(115),cout=>p(374)(116));
FA_ff_15314:FAff port map(x=>p(364)(116),y=>p(365)(116),Cin=>p(366)(116),clock=>clock,reset=>reset,s=>p(373)(116),cout=>p(374)(117));
FA_ff_15315:FAff port map(x=>p(364)(117),y=>p(365)(117),Cin=>p(366)(117),clock=>clock,reset=>reset,s=>p(373)(117),cout=>p(374)(118));
FA_ff_15316:FAff port map(x=>p(364)(118),y=>p(365)(118),Cin=>p(366)(118),clock=>clock,reset=>reset,s=>p(373)(118),cout=>p(374)(119));
FA_ff_15317:FAff port map(x=>p(364)(119),y=>p(365)(119),Cin=>p(366)(119),clock=>clock,reset=>reset,s=>p(373)(119),cout=>p(374)(120));
FA_ff_15318:FAff port map(x=>p(364)(120),y=>p(365)(120),Cin=>p(366)(120),clock=>clock,reset=>reset,s=>p(373)(120),cout=>p(374)(121));
FA_ff_15319:FAff port map(x=>p(364)(121),y=>p(365)(121),Cin=>p(366)(121),clock=>clock,reset=>reset,s=>p(373)(121),cout=>p(374)(122));
FA_ff_15320:FAff port map(x=>p(364)(122),y=>p(365)(122),Cin=>p(366)(122),clock=>clock,reset=>reset,s=>p(373)(122),cout=>p(374)(123));
FA_ff_15321:FAff port map(x=>p(364)(123),y=>p(365)(123),Cin=>p(366)(123),clock=>clock,reset=>reset,s=>p(373)(123),cout=>p(374)(124));
FA_ff_15322:FAff port map(x=>p(364)(124),y=>p(365)(124),Cin=>p(366)(124),clock=>clock,reset=>reset,s=>p(373)(124),cout=>p(374)(125));
FA_ff_15323:FAff port map(x=>p(364)(125),y=>p(365)(125),Cin=>p(366)(125),clock=>clock,reset=>reset,s=>p(373)(125),cout=>p(374)(126));
FA_ff_15324:FAff port map(x=>p(364)(126),y=>p(365)(126),Cin=>p(366)(126),clock=>clock,reset=>reset,s=>p(373)(126),cout=>p(374)(127));
FA_ff_15325:FAff port map(x=>p(364)(127),y=>p(365)(127),Cin=>p(366)(127),clock=>clock,reset=>reset,s=>p(373)(127),cout=>p(374)(128));
FA_ff_15326:FAff port map(x=>p(364)(128),y=>p(365)(128),Cin=>p(366)(128),clock=>clock,reset=>reset,s=>p(373)(128),cout=>p(374)(129));
FA_ff_15327:FAff port map(x=>p(364)(129),y=>p(365)(129),Cin=>p(366)(129),clock=>clock,reset=>reset,s=>p(373)(129),cout=>p(374)(130));
FA_ff_15328:FAff port map(x=>p(364)(130),y=>p(365)(130),Cin=>p(366)(130),clock=>clock,reset=>reset,s=>p(373)(130),cout=>p(374)(131));
FA_ff_15329:FAff port map(x=>p(364)(131),y=>p(365)(131),Cin=>p(366)(131),clock=>clock,reset=>reset,s=>p(373)(131),cout=>p(374)(132));
HA_ff_105:HAff port map(x=>p(367)(0),y=>p(369)(0),clock=>clock,reset=>reset,s=>p(375)(0),c=>p(376)(1));
FA_ff_15330:FAff port map(x=>p(367)(1),y=>p(368)(1),Cin=>p(369)(1),clock=>clock,reset=>reset,s=>p(375)(1),cout=>p(376)(2));
FA_ff_15331:FAff port map(x=>p(367)(2),y=>p(368)(2),Cin=>p(369)(2),clock=>clock,reset=>reset,s=>p(375)(2),cout=>p(376)(3));
FA_ff_15332:FAff port map(x=>p(367)(3),y=>p(368)(3),Cin=>p(369)(3),clock=>clock,reset=>reset,s=>p(375)(3),cout=>p(376)(4));
FA_ff_15333:FAff port map(x=>p(367)(4),y=>p(368)(4),Cin=>p(369)(4),clock=>clock,reset=>reset,s=>p(375)(4),cout=>p(376)(5));
FA_ff_15334:FAff port map(x=>p(367)(5),y=>p(368)(5),Cin=>p(369)(5),clock=>clock,reset=>reset,s=>p(375)(5),cout=>p(376)(6));
FA_ff_15335:FAff port map(x=>p(367)(6),y=>p(368)(6),Cin=>p(369)(6),clock=>clock,reset=>reset,s=>p(375)(6),cout=>p(376)(7));
FA_ff_15336:FAff port map(x=>p(367)(7),y=>p(368)(7),Cin=>p(369)(7),clock=>clock,reset=>reset,s=>p(375)(7),cout=>p(376)(8));
FA_ff_15337:FAff port map(x=>p(367)(8),y=>p(368)(8),Cin=>p(369)(8),clock=>clock,reset=>reset,s=>p(375)(8),cout=>p(376)(9));
FA_ff_15338:FAff port map(x=>p(367)(9),y=>p(368)(9),Cin=>p(369)(9),clock=>clock,reset=>reset,s=>p(375)(9),cout=>p(376)(10));
FA_ff_15339:FAff port map(x=>p(367)(10),y=>p(368)(10),Cin=>p(369)(10),clock=>clock,reset=>reset,s=>p(375)(10),cout=>p(376)(11));
FA_ff_15340:FAff port map(x=>p(367)(11),y=>p(368)(11),Cin=>p(369)(11),clock=>clock,reset=>reset,s=>p(375)(11),cout=>p(376)(12));
FA_ff_15341:FAff port map(x=>p(367)(12),y=>p(368)(12),Cin=>p(369)(12),clock=>clock,reset=>reset,s=>p(375)(12),cout=>p(376)(13));
FA_ff_15342:FAff port map(x=>p(367)(13),y=>p(368)(13),Cin=>p(369)(13),clock=>clock,reset=>reset,s=>p(375)(13),cout=>p(376)(14));
FA_ff_15343:FAff port map(x=>p(367)(14),y=>p(368)(14),Cin=>p(369)(14),clock=>clock,reset=>reset,s=>p(375)(14),cout=>p(376)(15));
FA_ff_15344:FAff port map(x=>p(367)(15),y=>p(368)(15),Cin=>p(369)(15),clock=>clock,reset=>reset,s=>p(375)(15),cout=>p(376)(16));
FA_ff_15345:FAff port map(x=>p(367)(16),y=>p(368)(16),Cin=>p(369)(16),clock=>clock,reset=>reset,s=>p(375)(16),cout=>p(376)(17));
FA_ff_15346:FAff port map(x=>p(367)(17),y=>p(368)(17),Cin=>p(369)(17),clock=>clock,reset=>reset,s=>p(375)(17),cout=>p(376)(18));
FA_ff_15347:FAff port map(x=>p(367)(18),y=>p(368)(18),Cin=>p(369)(18),clock=>clock,reset=>reset,s=>p(375)(18),cout=>p(376)(19));
FA_ff_15348:FAff port map(x=>p(367)(19),y=>p(368)(19),Cin=>p(369)(19),clock=>clock,reset=>reset,s=>p(375)(19),cout=>p(376)(20));
FA_ff_15349:FAff port map(x=>p(367)(20),y=>p(368)(20),Cin=>p(369)(20),clock=>clock,reset=>reset,s=>p(375)(20),cout=>p(376)(21));
FA_ff_15350:FAff port map(x=>p(367)(21),y=>p(368)(21),Cin=>p(369)(21),clock=>clock,reset=>reset,s=>p(375)(21),cout=>p(376)(22));
FA_ff_15351:FAff port map(x=>p(367)(22),y=>p(368)(22),Cin=>p(369)(22),clock=>clock,reset=>reset,s=>p(375)(22),cout=>p(376)(23));
FA_ff_15352:FAff port map(x=>p(367)(23),y=>p(368)(23),Cin=>p(369)(23),clock=>clock,reset=>reset,s=>p(375)(23),cout=>p(376)(24));
FA_ff_15353:FAff port map(x=>p(367)(24),y=>p(368)(24),Cin=>p(369)(24),clock=>clock,reset=>reset,s=>p(375)(24),cout=>p(376)(25));
FA_ff_15354:FAff port map(x=>p(367)(25),y=>p(368)(25),Cin=>p(369)(25),clock=>clock,reset=>reset,s=>p(375)(25),cout=>p(376)(26));
FA_ff_15355:FAff port map(x=>p(367)(26),y=>p(368)(26),Cin=>p(369)(26),clock=>clock,reset=>reset,s=>p(375)(26),cout=>p(376)(27));
FA_ff_15356:FAff port map(x=>p(367)(27),y=>p(368)(27),Cin=>p(369)(27),clock=>clock,reset=>reset,s=>p(375)(27),cout=>p(376)(28));
FA_ff_15357:FAff port map(x=>p(367)(28),y=>p(368)(28),Cin=>p(369)(28),clock=>clock,reset=>reset,s=>p(375)(28),cout=>p(376)(29));
FA_ff_15358:FAff port map(x=>p(367)(29),y=>p(368)(29),Cin=>p(369)(29),clock=>clock,reset=>reset,s=>p(375)(29),cout=>p(376)(30));
FA_ff_15359:FAff port map(x=>p(367)(30),y=>p(368)(30),Cin=>p(369)(30),clock=>clock,reset=>reset,s=>p(375)(30),cout=>p(376)(31));
FA_ff_15360:FAff port map(x=>p(367)(31),y=>p(368)(31),Cin=>p(369)(31),clock=>clock,reset=>reset,s=>p(375)(31),cout=>p(376)(32));
FA_ff_15361:FAff port map(x=>p(367)(32),y=>p(368)(32),Cin=>p(369)(32),clock=>clock,reset=>reset,s=>p(375)(32),cout=>p(376)(33));
FA_ff_15362:FAff port map(x=>p(367)(33),y=>p(368)(33),Cin=>p(369)(33),clock=>clock,reset=>reset,s=>p(375)(33),cout=>p(376)(34));
FA_ff_15363:FAff port map(x=>p(367)(34),y=>p(368)(34),Cin=>p(369)(34),clock=>clock,reset=>reset,s=>p(375)(34),cout=>p(376)(35));
FA_ff_15364:FAff port map(x=>p(367)(35),y=>p(368)(35),Cin=>p(369)(35),clock=>clock,reset=>reset,s=>p(375)(35),cout=>p(376)(36));
FA_ff_15365:FAff port map(x=>p(367)(36),y=>p(368)(36),Cin=>p(369)(36),clock=>clock,reset=>reset,s=>p(375)(36),cout=>p(376)(37));
FA_ff_15366:FAff port map(x=>p(367)(37),y=>p(368)(37),Cin=>p(369)(37),clock=>clock,reset=>reset,s=>p(375)(37),cout=>p(376)(38));
FA_ff_15367:FAff port map(x=>p(367)(38),y=>p(368)(38),Cin=>p(369)(38),clock=>clock,reset=>reset,s=>p(375)(38),cout=>p(376)(39));
FA_ff_15368:FAff port map(x=>p(367)(39),y=>p(368)(39),Cin=>p(369)(39),clock=>clock,reset=>reset,s=>p(375)(39),cout=>p(376)(40));
FA_ff_15369:FAff port map(x=>p(367)(40),y=>p(368)(40),Cin=>p(369)(40),clock=>clock,reset=>reset,s=>p(375)(40),cout=>p(376)(41));
FA_ff_15370:FAff port map(x=>p(367)(41),y=>p(368)(41),Cin=>p(369)(41),clock=>clock,reset=>reset,s=>p(375)(41),cout=>p(376)(42));
FA_ff_15371:FAff port map(x=>p(367)(42),y=>p(368)(42),Cin=>p(369)(42),clock=>clock,reset=>reset,s=>p(375)(42),cout=>p(376)(43));
FA_ff_15372:FAff port map(x=>p(367)(43),y=>p(368)(43),Cin=>p(369)(43),clock=>clock,reset=>reset,s=>p(375)(43),cout=>p(376)(44));
FA_ff_15373:FAff port map(x=>p(367)(44),y=>p(368)(44),Cin=>p(369)(44),clock=>clock,reset=>reset,s=>p(375)(44),cout=>p(376)(45));
FA_ff_15374:FAff port map(x=>p(367)(45),y=>p(368)(45),Cin=>p(369)(45),clock=>clock,reset=>reset,s=>p(375)(45),cout=>p(376)(46));
FA_ff_15375:FAff port map(x=>p(367)(46),y=>p(368)(46),Cin=>p(369)(46),clock=>clock,reset=>reset,s=>p(375)(46),cout=>p(376)(47));
FA_ff_15376:FAff port map(x=>p(367)(47),y=>p(368)(47),Cin=>p(369)(47),clock=>clock,reset=>reset,s=>p(375)(47),cout=>p(376)(48));
FA_ff_15377:FAff port map(x=>p(367)(48),y=>p(368)(48),Cin=>p(369)(48),clock=>clock,reset=>reset,s=>p(375)(48),cout=>p(376)(49));
FA_ff_15378:FAff port map(x=>p(367)(49),y=>p(368)(49),Cin=>p(369)(49),clock=>clock,reset=>reset,s=>p(375)(49),cout=>p(376)(50));
FA_ff_15379:FAff port map(x=>p(367)(50),y=>p(368)(50),Cin=>p(369)(50),clock=>clock,reset=>reset,s=>p(375)(50),cout=>p(376)(51));
FA_ff_15380:FAff port map(x=>p(367)(51),y=>p(368)(51),Cin=>p(369)(51),clock=>clock,reset=>reset,s=>p(375)(51),cout=>p(376)(52));
FA_ff_15381:FAff port map(x=>p(367)(52),y=>p(368)(52),Cin=>p(369)(52),clock=>clock,reset=>reset,s=>p(375)(52),cout=>p(376)(53));
FA_ff_15382:FAff port map(x=>p(367)(53),y=>p(368)(53),Cin=>p(369)(53),clock=>clock,reset=>reset,s=>p(375)(53),cout=>p(376)(54));
FA_ff_15383:FAff port map(x=>p(367)(54),y=>p(368)(54),Cin=>p(369)(54),clock=>clock,reset=>reset,s=>p(375)(54),cout=>p(376)(55));
FA_ff_15384:FAff port map(x=>p(367)(55),y=>p(368)(55),Cin=>p(369)(55),clock=>clock,reset=>reset,s=>p(375)(55),cout=>p(376)(56));
FA_ff_15385:FAff port map(x=>p(367)(56),y=>p(368)(56),Cin=>p(369)(56),clock=>clock,reset=>reset,s=>p(375)(56),cout=>p(376)(57));
FA_ff_15386:FAff port map(x=>p(367)(57),y=>p(368)(57),Cin=>p(369)(57),clock=>clock,reset=>reset,s=>p(375)(57),cout=>p(376)(58));
FA_ff_15387:FAff port map(x=>p(367)(58),y=>p(368)(58),Cin=>p(369)(58),clock=>clock,reset=>reset,s=>p(375)(58),cout=>p(376)(59));
FA_ff_15388:FAff port map(x=>p(367)(59),y=>p(368)(59),Cin=>p(369)(59),clock=>clock,reset=>reset,s=>p(375)(59),cout=>p(376)(60));
FA_ff_15389:FAff port map(x=>p(367)(60),y=>p(368)(60),Cin=>p(369)(60),clock=>clock,reset=>reset,s=>p(375)(60),cout=>p(376)(61));
FA_ff_15390:FAff port map(x=>p(367)(61),y=>p(368)(61),Cin=>p(369)(61),clock=>clock,reset=>reset,s=>p(375)(61),cout=>p(376)(62));
FA_ff_15391:FAff port map(x=>p(367)(62),y=>p(368)(62),Cin=>p(369)(62),clock=>clock,reset=>reset,s=>p(375)(62),cout=>p(376)(63));
FA_ff_15392:FAff port map(x=>p(367)(63),y=>p(368)(63),Cin=>p(369)(63),clock=>clock,reset=>reset,s=>p(375)(63),cout=>p(376)(64));
FA_ff_15393:FAff port map(x=>p(367)(64),y=>p(368)(64),Cin=>p(369)(64),clock=>clock,reset=>reset,s=>p(375)(64),cout=>p(376)(65));
FA_ff_15394:FAff port map(x=>p(367)(65),y=>p(368)(65),Cin=>p(369)(65),clock=>clock,reset=>reset,s=>p(375)(65),cout=>p(376)(66));
FA_ff_15395:FAff port map(x=>p(367)(66),y=>p(368)(66),Cin=>p(369)(66),clock=>clock,reset=>reset,s=>p(375)(66),cout=>p(376)(67));
FA_ff_15396:FAff port map(x=>p(367)(67),y=>p(368)(67),Cin=>p(369)(67),clock=>clock,reset=>reset,s=>p(375)(67),cout=>p(376)(68));
FA_ff_15397:FAff port map(x=>p(367)(68),y=>p(368)(68),Cin=>p(369)(68),clock=>clock,reset=>reset,s=>p(375)(68),cout=>p(376)(69));
FA_ff_15398:FAff port map(x=>p(367)(69),y=>p(368)(69),Cin=>p(369)(69),clock=>clock,reset=>reset,s=>p(375)(69),cout=>p(376)(70));
FA_ff_15399:FAff port map(x=>p(367)(70),y=>p(368)(70),Cin=>p(369)(70),clock=>clock,reset=>reset,s=>p(375)(70),cout=>p(376)(71));
FA_ff_15400:FAff port map(x=>p(367)(71),y=>p(368)(71),Cin=>p(369)(71),clock=>clock,reset=>reset,s=>p(375)(71),cout=>p(376)(72));
FA_ff_15401:FAff port map(x=>p(367)(72),y=>p(368)(72),Cin=>p(369)(72),clock=>clock,reset=>reset,s=>p(375)(72),cout=>p(376)(73));
FA_ff_15402:FAff port map(x=>p(367)(73),y=>p(368)(73),Cin=>p(369)(73),clock=>clock,reset=>reset,s=>p(375)(73),cout=>p(376)(74));
FA_ff_15403:FAff port map(x=>p(367)(74),y=>p(368)(74),Cin=>p(369)(74),clock=>clock,reset=>reset,s=>p(375)(74),cout=>p(376)(75));
FA_ff_15404:FAff port map(x=>p(367)(75),y=>p(368)(75),Cin=>p(369)(75),clock=>clock,reset=>reset,s=>p(375)(75),cout=>p(376)(76));
FA_ff_15405:FAff port map(x=>p(367)(76),y=>p(368)(76),Cin=>p(369)(76),clock=>clock,reset=>reset,s=>p(375)(76),cout=>p(376)(77));
FA_ff_15406:FAff port map(x=>p(367)(77),y=>p(368)(77),Cin=>p(369)(77),clock=>clock,reset=>reset,s=>p(375)(77),cout=>p(376)(78));
FA_ff_15407:FAff port map(x=>p(367)(78),y=>p(368)(78),Cin=>p(369)(78),clock=>clock,reset=>reset,s=>p(375)(78),cout=>p(376)(79));
FA_ff_15408:FAff port map(x=>p(367)(79),y=>p(368)(79),Cin=>p(369)(79),clock=>clock,reset=>reset,s=>p(375)(79),cout=>p(376)(80));
FA_ff_15409:FAff port map(x=>p(367)(80),y=>p(368)(80),Cin=>p(369)(80),clock=>clock,reset=>reset,s=>p(375)(80),cout=>p(376)(81));
FA_ff_15410:FAff port map(x=>p(367)(81),y=>p(368)(81),Cin=>p(369)(81),clock=>clock,reset=>reset,s=>p(375)(81),cout=>p(376)(82));
FA_ff_15411:FAff port map(x=>p(367)(82),y=>p(368)(82),Cin=>p(369)(82),clock=>clock,reset=>reset,s=>p(375)(82),cout=>p(376)(83));
FA_ff_15412:FAff port map(x=>p(367)(83),y=>p(368)(83),Cin=>p(369)(83),clock=>clock,reset=>reset,s=>p(375)(83),cout=>p(376)(84));
FA_ff_15413:FAff port map(x=>p(367)(84),y=>p(368)(84),Cin=>p(369)(84),clock=>clock,reset=>reset,s=>p(375)(84),cout=>p(376)(85));
FA_ff_15414:FAff port map(x=>p(367)(85),y=>p(368)(85),Cin=>p(369)(85),clock=>clock,reset=>reset,s=>p(375)(85),cout=>p(376)(86));
FA_ff_15415:FAff port map(x=>p(367)(86),y=>p(368)(86),Cin=>p(369)(86),clock=>clock,reset=>reset,s=>p(375)(86),cout=>p(376)(87));
FA_ff_15416:FAff port map(x=>p(367)(87),y=>p(368)(87),Cin=>p(369)(87),clock=>clock,reset=>reset,s=>p(375)(87),cout=>p(376)(88));
FA_ff_15417:FAff port map(x=>p(367)(88),y=>p(368)(88),Cin=>p(369)(88),clock=>clock,reset=>reset,s=>p(375)(88),cout=>p(376)(89));
FA_ff_15418:FAff port map(x=>p(367)(89),y=>p(368)(89),Cin=>p(369)(89),clock=>clock,reset=>reset,s=>p(375)(89),cout=>p(376)(90));
FA_ff_15419:FAff port map(x=>p(367)(90),y=>p(368)(90),Cin=>p(369)(90),clock=>clock,reset=>reset,s=>p(375)(90),cout=>p(376)(91));
FA_ff_15420:FAff port map(x=>p(367)(91),y=>p(368)(91),Cin=>p(369)(91),clock=>clock,reset=>reset,s=>p(375)(91),cout=>p(376)(92));
FA_ff_15421:FAff port map(x=>p(367)(92),y=>p(368)(92),Cin=>p(369)(92),clock=>clock,reset=>reset,s=>p(375)(92),cout=>p(376)(93));
FA_ff_15422:FAff port map(x=>p(367)(93),y=>p(368)(93),Cin=>p(369)(93),clock=>clock,reset=>reset,s=>p(375)(93),cout=>p(376)(94));
FA_ff_15423:FAff port map(x=>p(367)(94),y=>p(368)(94),Cin=>p(369)(94),clock=>clock,reset=>reset,s=>p(375)(94),cout=>p(376)(95));
FA_ff_15424:FAff port map(x=>p(367)(95),y=>p(368)(95),Cin=>p(369)(95),clock=>clock,reset=>reset,s=>p(375)(95),cout=>p(376)(96));
FA_ff_15425:FAff port map(x=>p(367)(96),y=>p(368)(96),Cin=>p(369)(96),clock=>clock,reset=>reset,s=>p(375)(96),cout=>p(376)(97));
FA_ff_15426:FAff port map(x=>p(367)(97),y=>p(368)(97),Cin=>p(369)(97),clock=>clock,reset=>reset,s=>p(375)(97),cout=>p(376)(98));
FA_ff_15427:FAff port map(x=>p(367)(98),y=>p(368)(98),Cin=>p(369)(98),clock=>clock,reset=>reset,s=>p(375)(98),cout=>p(376)(99));
FA_ff_15428:FAff port map(x=>p(367)(99),y=>p(368)(99),Cin=>p(369)(99),clock=>clock,reset=>reset,s=>p(375)(99),cout=>p(376)(100));
FA_ff_15429:FAff port map(x=>p(367)(100),y=>p(368)(100),Cin=>p(369)(100),clock=>clock,reset=>reset,s=>p(375)(100),cout=>p(376)(101));
FA_ff_15430:FAff port map(x=>p(367)(101),y=>p(368)(101),Cin=>p(369)(101),clock=>clock,reset=>reset,s=>p(375)(101),cout=>p(376)(102));
FA_ff_15431:FAff port map(x=>p(367)(102),y=>p(368)(102),Cin=>p(369)(102),clock=>clock,reset=>reset,s=>p(375)(102),cout=>p(376)(103));
FA_ff_15432:FAff port map(x=>p(367)(103),y=>p(368)(103),Cin=>p(369)(103),clock=>clock,reset=>reset,s=>p(375)(103),cout=>p(376)(104));
FA_ff_15433:FAff port map(x=>p(367)(104),y=>p(368)(104),Cin=>p(369)(104),clock=>clock,reset=>reset,s=>p(375)(104),cout=>p(376)(105));
FA_ff_15434:FAff port map(x=>p(367)(105),y=>p(368)(105),Cin=>p(369)(105),clock=>clock,reset=>reset,s=>p(375)(105),cout=>p(376)(106));
FA_ff_15435:FAff port map(x=>p(367)(106),y=>p(368)(106),Cin=>p(369)(106),clock=>clock,reset=>reset,s=>p(375)(106),cout=>p(376)(107));
FA_ff_15436:FAff port map(x=>p(367)(107),y=>p(368)(107),Cin=>p(369)(107),clock=>clock,reset=>reset,s=>p(375)(107),cout=>p(376)(108));
FA_ff_15437:FAff port map(x=>p(367)(108),y=>p(368)(108),Cin=>p(369)(108),clock=>clock,reset=>reset,s=>p(375)(108),cout=>p(376)(109));
FA_ff_15438:FAff port map(x=>p(367)(109),y=>p(368)(109),Cin=>p(369)(109),clock=>clock,reset=>reset,s=>p(375)(109),cout=>p(376)(110));
FA_ff_15439:FAff port map(x=>p(367)(110),y=>p(368)(110),Cin=>p(369)(110),clock=>clock,reset=>reset,s=>p(375)(110),cout=>p(376)(111));
FA_ff_15440:FAff port map(x=>p(367)(111),y=>p(368)(111),Cin=>p(369)(111),clock=>clock,reset=>reset,s=>p(375)(111),cout=>p(376)(112));
FA_ff_15441:FAff port map(x=>p(367)(112),y=>p(368)(112),Cin=>p(369)(112),clock=>clock,reset=>reset,s=>p(375)(112),cout=>p(376)(113));
FA_ff_15442:FAff port map(x=>p(367)(113),y=>p(368)(113),Cin=>p(369)(113),clock=>clock,reset=>reset,s=>p(375)(113),cout=>p(376)(114));
FA_ff_15443:FAff port map(x=>p(367)(114),y=>p(368)(114),Cin=>p(369)(114),clock=>clock,reset=>reset,s=>p(375)(114),cout=>p(376)(115));
FA_ff_15444:FAff port map(x=>p(367)(115),y=>p(368)(115),Cin=>p(369)(115),clock=>clock,reset=>reset,s=>p(375)(115),cout=>p(376)(116));
FA_ff_15445:FAff port map(x=>p(367)(116),y=>p(368)(116),Cin=>p(369)(116),clock=>clock,reset=>reset,s=>p(375)(116),cout=>p(376)(117));
FA_ff_15446:FAff port map(x=>p(367)(117),y=>p(368)(117),Cin=>p(369)(117),clock=>clock,reset=>reset,s=>p(375)(117),cout=>p(376)(118));
FA_ff_15447:FAff port map(x=>p(367)(118),y=>p(368)(118),Cin=>p(369)(118),clock=>clock,reset=>reset,s=>p(375)(118),cout=>p(376)(119));
FA_ff_15448:FAff port map(x=>p(367)(119),y=>p(368)(119),Cin=>p(369)(119),clock=>clock,reset=>reset,s=>p(375)(119),cout=>p(376)(120));
FA_ff_15449:FAff port map(x=>p(367)(120),y=>p(368)(120),Cin=>p(369)(120),clock=>clock,reset=>reset,s=>p(375)(120),cout=>p(376)(121));
FA_ff_15450:FAff port map(x=>p(367)(121),y=>p(368)(121),Cin=>p(369)(121),clock=>clock,reset=>reset,s=>p(375)(121),cout=>p(376)(122));
FA_ff_15451:FAff port map(x=>p(367)(122),y=>p(368)(122),Cin=>p(369)(122),clock=>clock,reset=>reset,s=>p(375)(122),cout=>p(376)(123));
FA_ff_15452:FAff port map(x=>p(367)(123),y=>p(368)(123),Cin=>p(369)(123),clock=>clock,reset=>reset,s=>p(375)(123),cout=>p(376)(124));
FA_ff_15453:FAff port map(x=>p(367)(124),y=>p(368)(124),Cin=>p(369)(124),clock=>clock,reset=>reset,s=>p(375)(124),cout=>p(376)(125));
FA_ff_15454:FAff port map(x=>p(367)(125),y=>p(368)(125),Cin=>p(369)(125),clock=>clock,reset=>reset,s=>p(375)(125),cout=>p(376)(126));
FA_ff_15455:FAff port map(x=>p(367)(126),y=>p(368)(126),Cin=>p(369)(126),clock=>clock,reset=>reset,s=>p(375)(126),cout=>p(376)(127));
FA_ff_15456:FAff port map(x=>p(367)(127),y=>p(368)(127),Cin=>p(369)(127),clock=>clock,reset=>reset,s=>p(375)(127),cout=>p(376)(128));
FA_ff_15457:FAff port map(x=>p(367)(128),y=>p(368)(128),Cin=>p(369)(128),clock=>clock,reset=>reset,s=>p(375)(128),cout=>p(376)(129));
FA_ff_15458:FAff port map(x=>p(367)(129),y=>p(368)(129),Cin=>p(369)(129),clock=>clock,reset=>reset,s=>p(375)(129),cout=>p(376)(130));
FA_ff_15459:FAff port map(x=>p(367)(130),y=>p(368)(130),Cin=>p(369)(130),clock=>clock,reset=>reset,s=>p(375)(130),cout=>p(376)(131));
FA_ff_15460:FAff port map(x=>p(367)(131),y=>p(368)(131),Cin=>p(369)(131),clock=>clock,reset=>reset,s=>p(375)(131),cout=>p(376)(132));
p(375)(132)<=p(368)(132);
p(377)(0)<=p(371)(0);
HA_ff_106:HAff port map(x=>p(371)(1),y=>p(372)(1),clock=>clock,reset=>reset,s=>p(377)(1),c=>p(378)(2));
FA_ff_15461:FAff port map(x=>p(370)(2),y=>p(371)(2),Cin=>p(372)(2),clock=>clock,reset=>reset,s=>p(377)(2),cout=>p(378)(3));
FA_ff_15462:FAff port map(x=>p(370)(3),y=>p(371)(3),Cin=>p(372)(3),clock=>clock,reset=>reset,s=>p(377)(3),cout=>p(378)(4));
FA_ff_15463:FAff port map(x=>p(370)(4),y=>p(371)(4),Cin=>p(372)(4),clock=>clock,reset=>reset,s=>p(377)(4),cout=>p(378)(5));
FA_ff_15464:FAff port map(x=>p(370)(5),y=>p(371)(5),Cin=>p(372)(5),clock=>clock,reset=>reset,s=>p(377)(5),cout=>p(378)(6));
FA_ff_15465:FAff port map(x=>p(370)(6),y=>p(371)(6),Cin=>p(372)(6),clock=>clock,reset=>reset,s=>p(377)(6),cout=>p(378)(7));
FA_ff_15466:FAff port map(x=>p(370)(7),y=>p(371)(7),Cin=>p(372)(7),clock=>clock,reset=>reset,s=>p(377)(7),cout=>p(378)(8));
FA_ff_15467:FAff port map(x=>p(370)(8),y=>p(371)(8),Cin=>p(372)(8),clock=>clock,reset=>reset,s=>p(377)(8),cout=>p(378)(9));
FA_ff_15468:FAff port map(x=>p(370)(9),y=>p(371)(9),Cin=>p(372)(9),clock=>clock,reset=>reset,s=>p(377)(9),cout=>p(378)(10));
FA_ff_15469:FAff port map(x=>p(370)(10),y=>p(371)(10),Cin=>p(372)(10),clock=>clock,reset=>reset,s=>p(377)(10),cout=>p(378)(11));
FA_ff_15470:FAff port map(x=>p(370)(11),y=>p(371)(11),Cin=>p(372)(11),clock=>clock,reset=>reset,s=>p(377)(11),cout=>p(378)(12));
FA_ff_15471:FAff port map(x=>p(370)(12),y=>p(371)(12),Cin=>p(372)(12),clock=>clock,reset=>reset,s=>p(377)(12),cout=>p(378)(13));
FA_ff_15472:FAff port map(x=>p(370)(13),y=>p(371)(13),Cin=>p(372)(13),clock=>clock,reset=>reset,s=>p(377)(13),cout=>p(378)(14));
FA_ff_15473:FAff port map(x=>p(370)(14),y=>p(371)(14),Cin=>p(372)(14),clock=>clock,reset=>reset,s=>p(377)(14),cout=>p(378)(15));
FA_ff_15474:FAff port map(x=>p(370)(15),y=>p(371)(15),Cin=>p(372)(15),clock=>clock,reset=>reset,s=>p(377)(15),cout=>p(378)(16));
FA_ff_15475:FAff port map(x=>p(370)(16),y=>p(371)(16),Cin=>p(372)(16),clock=>clock,reset=>reset,s=>p(377)(16),cout=>p(378)(17));
FA_ff_15476:FAff port map(x=>p(370)(17),y=>p(371)(17),Cin=>p(372)(17),clock=>clock,reset=>reset,s=>p(377)(17),cout=>p(378)(18));
FA_ff_15477:FAff port map(x=>p(370)(18),y=>p(371)(18),Cin=>p(372)(18),clock=>clock,reset=>reset,s=>p(377)(18),cout=>p(378)(19));
FA_ff_15478:FAff port map(x=>p(370)(19),y=>p(371)(19),Cin=>p(372)(19),clock=>clock,reset=>reset,s=>p(377)(19),cout=>p(378)(20));
FA_ff_15479:FAff port map(x=>p(370)(20),y=>p(371)(20),Cin=>p(372)(20),clock=>clock,reset=>reset,s=>p(377)(20),cout=>p(378)(21));
FA_ff_15480:FAff port map(x=>p(370)(21),y=>p(371)(21),Cin=>p(372)(21),clock=>clock,reset=>reset,s=>p(377)(21),cout=>p(378)(22));
FA_ff_15481:FAff port map(x=>p(370)(22),y=>p(371)(22),Cin=>p(372)(22),clock=>clock,reset=>reset,s=>p(377)(22),cout=>p(378)(23));
FA_ff_15482:FAff port map(x=>p(370)(23),y=>p(371)(23),Cin=>p(372)(23),clock=>clock,reset=>reset,s=>p(377)(23),cout=>p(378)(24));
FA_ff_15483:FAff port map(x=>p(370)(24),y=>p(371)(24),Cin=>p(372)(24),clock=>clock,reset=>reset,s=>p(377)(24),cout=>p(378)(25));
FA_ff_15484:FAff port map(x=>p(370)(25),y=>p(371)(25),Cin=>p(372)(25),clock=>clock,reset=>reset,s=>p(377)(25),cout=>p(378)(26));
FA_ff_15485:FAff port map(x=>p(370)(26),y=>p(371)(26),Cin=>p(372)(26),clock=>clock,reset=>reset,s=>p(377)(26),cout=>p(378)(27));
FA_ff_15486:FAff port map(x=>p(370)(27),y=>p(371)(27),Cin=>p(372)(27),clock=>clock,reset=>reset,s=>p(377)(27),cout=>p(378)(28));
FA_ff_15487:FAff port map(x=>p(370)(28),y=>p(371)(28),Cin=>p(372)(28),clock=>clock,reset=>reset,s=>p(377)(28),cout=>p(378)(29));
FA_ff_15488:FAff port map(x=>p(370)(29),y=>p(371)(29),Cin=>p(372)(29),clock=>clock,reset=>reset,s=>p(377)(29),cout=>p(378)(30));
FA_ff_15489:FAff port map(x=>p(370)(30),y=>p(371)(30),Cin=>p(372)(30),clock=>clock,reset=>reset,s=>p(377)(30),cout=>p(378)(31));
FA_ff_15490:FAff port map(x=>p(370)(31),y=>p(371)(31),Cin=>p(372)(31),clock=>clock,reset=>reset,s=>p(377)(31),cout=>p(378)(32));
FA_ff_15491:FAff port map(x=>p(370)(32),y=>p(371)(32),Cin=>p(372)(32),clock=>clock,reset=>reset,s=>p(377)(32),cout=>p(378)(33));
FA_ff_15492:FAff port map(x=>p(370)(33),y=>p(371)(33),Cin=>p(372)(33),clock=>clock,reset=>reset,s=>p(377)(33),cout=>p(378)(34));
FA_ff_15493:FAff port map(x=>p(370)(34),y=>p(371)(34),Cin=>p(372)(34),clock=>clock,reset=>reset,s=>p(377)(34),cout=>p(378)(35));
FA_ff_15494:FAff port map(x=>p(370)(35),y=>p(371)(35),Cin=>p(372)(35),clock=>clock,reset=>reset,s=>p(377)(35),cout=>p(378)(36));
FA_ff_15495:FAff port map(x=>p(370)(36),y=>p(371)(36),Cin=>p(372)(36),clock=>clock,reset=>reset,s=>p(377)(36),cout=>p(378)(37));
FA_ff_15496:FAff port map(x=>p(370)(37),y=>p(371)(37),Cin=>p(372)(37),clock=>clock,reset=>reset,s=>p(377)(37),cout=>p(378)(38));
FA_ff_15497:FAff port map(x=>p(370)(38),y=>p(371)(38),Cin=>p(372)(38),clock=>clock,reset=>reset,s=>p(377)(38),cout=>p(378)(39));
FA_ff_15498:FAff port map(x=>p(370)(39),y=>p(371)(39),Cin=>p(372)(39),clock=>clock,reset=>reset,s=>p(377)(39),cout=>p(378)(40));
FA_ff_15499:FAff port map(x=>p(370)(40),y=>p(371)(40),Cin=>p(372)(40),clock=>clock,reset=>reset,s=>p(377)(40),cout=>p(378)(41));
FA_ff_15500:FAff port map(x=>p(370)(41),y=>p(371)(41),Cin=>p(372)(41),clock=>clock,reset=>reset,s=>p(377)(41),cout=>p(378)(42));
FA_ff_15501:FAff port map(x=>p(370)(42),y=>p(371)(42),Cin=>p(372)(42),clock=>clock,reset=>reset,s=>p(377)(42),cout=>p(378)(43));
FA_ff_15502:FAff port map(x=>p(370)(43),y=>p(371)(43),Cin=>p(372)(43),clock=>clock,reset=>reset,s=>p(377)(43),cout=>p(378)(44));
FA_ff_15503:FAff port map(x=>p(370)(44),y=>p(371)(44),Cin=>p(372)(44),clock=>clock,reset=>reset,s=>p(377)(44),cout=>p(378)(45));
FA_ff_15504:FAff port map(x=>p(370)(45),y=>p(371)(45),Cin=>p(372)(45),clock=>clock,reset=>reset,s=>p(377)(45),cout=>p(378)(46));
FA_ff_15505:FAff port map(x=>p(370)(46),y=>p(371)(46),Cin=>p(372)(46),clock=>clock,reset=>reset,s=>p(377)(46),cout=>p(378)(47));
FA_ff_15506:FAff port map(x=>p(370)(47),y=>p(371)(47),Cin=>p(372)(47),clock=>clock,reset=>reset,s=>p(377)(47),cout=>p(378)(48));
FA_ff_15507:FAff port map(x=>p(370)(48),y=>p(371)(48),Cin=>p(372)(48),clock=>clock,reset=>reset,s=>p(377)(48),cout=>p(378)(49));
FA_ff_15508:FAff port map(x=>p(370)(49),y=>p(371)(49),Cin=>p(372)(49),clock=>clock,reset=>reset,s=>p(377)(49),cout=>p(378)(50));
FA_ff_15509:FAff port map(x=>p(370)(50),y=>p(371)(50),Cin=>p(372)(50),clock=>clock,reset=>reset,s=>p(377)(50),cout=>p(378)(51));
FA_ff_15510:FAff port map(x=>p(370)(51),y=>p(371)(51),Cin=>p(372)(51),clock=>clock,reset=>reset,s=>p(377)(51),cout=>p(378)(52));
FA_ff_15511:FAff port map(x=>p(370)(52),y=>p(371)(52),Cin=>p(372)(52),clock=>clock,reset=>reset,s=>p(377)(52),cout=>p(378)(53));
FA_ff_15512:FAff port map(x=>p(370)(53),y=>p(371)(53),Cin=>p(372)(53),clock=>clock,reset=>reset,s=>p(377)(53),cout=>p(378)(54));
FA_ff_15513:FAff port map(x=>p(370)(54),y=>p(371)(54),Cin=>p(372)(54),clock=>clock,reset=>reset,s=>p(377)(54),cout=>p(378)(55));
FA_ff_15514:FAff port map(x=>p(370)(55),y=>p(371)(55),Cin=>p(372)(55),clock=>clock,reset=>reset,s=>p(377)(55),cout=>p(378)(56));
FA_ff_15515:FAff port map(x=>p(370)(56),y=>p(371)(56),Cin=>p(372)(56),clock=>clock,reset=>reset,s=>p(377)(56),cout=>p(378)(57));
FA_ff_15516:FAff port map(x=>p(370)(57),y=>p(371)(57),Cin=>p(372)(57),clock=>clock,reset=>reset,s=>p(377)(57),cout=>p(378)(58));
FA_ff_15517:FAff port map(x=>p(370)(58),y=>p(371)(58),Cin=>p(372)(58),clock=>clock,reset=>reset,s=>p(377)(58),cout=>p(378)(59));
FA_ff_15518:FAff port map(x=>p(370)(59),y=>p(371)(59),Cin=>p(372)(59),clock=>clock,reset=>reset,s=>p(377)(59),cout=>p(378)(60));
FA_ff_15519:FAff port map(x=>p(370)(60),y=>p(371)(60),Cin=>p(372)(60),clock=>clock,reset=>reset,s=>p(377)(60),cout=>p(378)(61));
FA_ff_15520:FAff port map(x=>p(370)(61),y=>p(371)(61),Cin=>p(372)(61),clock=>clock,reset=>reset,s=>p(377)(61),cout=>p(378)(62));
FA_ff_15521:FAff port map(x=>p(370)(62),y=>p(371)(62),Cin=>p(372)(62),clock=>clock,reset=>reset,s=>p(377)(62),cout=>p(378)(63));
FA_ff_15522:FAff port map(x=>p(370)(63),y=>p(371)(63),Cin=>p(372)(63),clock=>clock,reset=>reset,s=>p(377)(63),cout=>p(378)(64));
FA_ff_15523:FAff port map(x=>p(370)(64),y=>p(371)(64),Cin=>p(372)(64),clock=>clock,reset=>reset,s=>p(377)(64),cout=>p(378)(65));
FA_ff_15524:FAff port map(x=>p(370)(65),y=>p(371)(65),Cin=>p(372)(65),clock=>clock,reset=>reset,s=>p(377)(65),cout=>p(378)(66));
FA_ff_15525:FAff port map(x=>p(370)(66),y=>p(371)(66),Cin=>p(372)(66),clock=>clock,reset=>reset,s=>p(377)(66),cout=>p(378)(67));
FA_ff_15526:FAff port map(x=>p(370)(67),y=>p(371)(67),Cin=>p(372)(67),clock=>clock,reset=>reset,s=>p(377)(67),cout=>p(378)(68));
FA_ff_15527:FAff port map(x=>p(370)(68),y=>p(371)(68),Cin=>p(372)(68),clock=>clock,reset=>reset,s=>p(377)(68),cout=>p(378)(69));
FA_ff_15528:FAff port map(x=>p(370)(69),y=>p(371)(69),Cin=>p(372)(69),clock=>clock,reset=>reset,s=>p(377)(69),cout=>p(378)(70));
FA_ff_15529:FAff port map(x=>p(370)(70),y=>p(371)(70),Cin=>p(372)(70),clock=>clock,reset=>reset,s=>p(377)(70),cout=>p(378)(71));
FA_ff_15530:FAff port map(x=>p(370)(71),y=>p(371)(71),Cin=>p(372)(71),clock=>clock,reset=>reset,s=>p(377)(71),cout=>p(378)(72));
FA_ff_15531:FAff port map(x=>p(370)(72),y=>p(371)(72),Cin=>p(372)(72),clock=>clock,reset=>reset,s=>p(377)(72),cout=>p(378)(73));
FA_ff_15532:FAff port map(x=>p(370)(73),y=>p(371)(73),Cin=>p(372)(73),clock=>clock,reset=>reset,s=>p(377)(73),cout=>p(378)(74));
FA_ff_15533:FAff port map(x=>p(370)(74),y=>p(371)(74),Cin=>p(372)(74),clock=>clock,reset=>reset,s=>p(377)(74),cout=>p(378)(75));
FA_ff_15534:FAff port map(x=>p(370)(75),y=>p(371)(75),Cin=>p(372)(75),clock=>clock,reset=>reset,s=>p(377)(75),cout=>p(378)(76));
FA_ff_15535:FAff port map(x=>p(370)(76),y=>p(371)(76),Cin=>p(372)(76),clock=>clock,reset=>reset,s=>p(377)(76),cout=>p(378)(77));
FA_ff_15536:FAff port map(x=>p(370)(77),y=>p(371)(77),Cin=>p(372)(77),clock=>clock,reset=>reset,s=>p(377)(77),cout=>p(378)(78));
FA_ff_15537:FAff port map(x=>p(370)(78),y=>p(371)(78),Cin=>p(372)(78),clock=>clock,reset=>reset,s=>p(377)(78),cout=>p(378)(79));
FA_ff_15538:FAff port map(x=>p(370)(79),y=>p(371)(79),Cin=>p(372)(79),clock=>clock,reset=>reset,s=>p(377)(79),cout=>p(378)(80));
FA_ff_15539:FAff port map(x=>p(370)(80),y=>p(371)(80),Cin=>p(372)(80),clock=>clock,reset=>reset,s=>p(377)(80),cout=>p(378)(81));
FA_ff_15540:FAff port map(x=>p(370)(81),y=>p(371)(81),Cin=>p(372)(81),clock=>clock,reset=>reset,s=>p(377)(81),cout=>p(378)(82));
FA_ff_15541:FAff port map(x=>p(370)(82),y=>p(371)(82),Cin=>p(372)(82),clock=>clock,reset=>reset,s=>p(377)(82),cout=>p(378)(83));
FA_ff_15542:FAff port map(x=>p(370)(83),y=>p(371)(83),Cin=>p(372)(83),clock=>clock,reset=>reset,s=>p(377)(83),cout=>p(378)(84));
FA_ff_15543:FAff port map(x=>p(370)(84),y=>p(371)(84),Cin=>p(372)(84),clock=>clock,reset=>reset,s=>p(377)(84),cout=>p(378)(85));
FA_ff_15544:FAff port map(x=>p(370)(85),y=>p(371)(85),Cin=>p(372)(85),clock=>clock,reset=>reset,s=>p(377)(85),cout=>p(378)(86));
FA_ff_15545:FAff port map(x=>p(370)(86),y=>p(371)(86),Cin=>p(372)(86),clock=>clock,reset=>reset,s=>p(377)(86),cout=>p(378)(87));
FA_ff_15546:FAff port map(x=>p(370)(87),y=>p(371)(87),Cin=>p(372)(87),clock=>clock,reset=>reset,s=>p(377)(87),cout=>p(378)(88));
FA_ff_15547:FAff port map(x=>p(370)(88),y=>p(371)(88),Cin=>p(372)(88),clock=>clock,reset=>reset,s=>p(377)(88),cout=>p(378)(89));
FA_ff_15548:FAff port map(x=>p(370)(89),y=>p(371)(89),Cin=>p(372)(89),clock=>clock,reset=>reset,s=>p(377)(89),cout=>p(378)(90));
FA_ff_15549:FAff port map(x=>p(370)(90),y=>p(371)(90),Cin=>p(372)(90),clock=>clock,reset=>reset,s=>p(377)(90),cout=>p(378)(91));
FA_ff_15550:FAff port map(x=>p(370)(91),y=>p(371)(91),Cin=>p(372)(91),clock=>clock,reset=>reset,s=>p(377)(91),cout=>p(378)(92));
FA_ff_15551:FAff port map(x=>p(370)(92),y=>p(371)(92),Cin=>p(372)(92),clock=>clock,reset=>reset,s=>p(377)(92),cout=>p(378)(93));
FA_ff_15552:FAff port map(x=>p(370)(93),y=>p(371)(93),Cin=>p(372)(93),clock=>clock,reset=>reset,s=>p(377)(93),cout=>p(378)(94));
FA_ff_15553:FAff port map(x=>p(370)(94),y=>p(371)(94),Cin=>p(372)(94),clock=>clock,reset=>reset,s=>p(377)(94),cout=>p(378)(95));
FA_ff_15554:FAff port map(x=>p(370)(95),y=>p(371)(95),Cin=>p(372)(95),clock=>clock,reset=>reset,s=>p(377)(95),cout=>p(378)(96));
FA_ff_15555:FAff port map(x=>p(370)(96),y=>p(371)(96),Cin=>p(372)(96),clock=>clock,reset=>reset,s=>p(377)(96),cout=>p(378)(97));
FA_ff_15556:FAff port map(x=>p(370)(97),y=>p(371)(97),Cin=>p(372)(97),clock=>clock,reset=>reset,s=>p(377)(97),cout=>p(378)(98));
FA_ff_15557:FAff port map(x=>p(370)(98),y=>p(371)(98),Cin=>p(372)(98),clock=>clock,reset=>reset,s=>p(377)(98),cout=>p(378)(99));
FA_ff_15558:FAff port map(x=>p(370)(99),y=>p(371)(99),Cin=>p(372)(99),clock=>clock,reset=>reset,s=>p(377)(99),cout=>p(378)(100));
FA_ff_15559:FAff port map(x=>p(370)(100),y=>p(371)(100),Cin=>p(372)(100),clock=>clock,reset=>reset,s=>p(377)(100),cout=>p(378)(101));
FA_ff_15560:FAff port map(x=>p(370)(101),y=>p(371)(101),Cin=>p(372)(101),clock=>clock,reset=>reset,s=>p(377)(101),cout=>p(378)(102));
FA_ff_15561:FAff port map(x=>p(370)(102),y=>p(371)(102),Cin=>p(372)(102),clock=>clock,reset=>reset,s=>p(377)(102),cout=>p(378)(103));
FA_ff_15562:FAff port map(x=>p(370)(103),y=>p(371)(103),Cin=>p(372)(103),clock=>clock,reset=>reset,s=>p(377)(103),cout=>p(378)(104));
FA_ff_15563:FAff port map(x=>p(370)(104),y=>p(371)(104),Cin=>p(372)(104),clock=>clock,reset=>reset,s=>p(377)(104),cout=>p(378)(105));
FA_ff_15564:FAff port map(x=>p(370)(105),y=>p(371)(105),Cin=>p(372)(105),clock=>clock,reset=>reset,s=>p(377)(105),cout=>p(378)(106));
FA_ff_15565:FAff port map(x=>p(370)(106),y=>p(371)(106),Cin=>p(372)(106),clock=>clock,reset=>reset,s=>p(377)(106),cout=>p(378)(107));
FA_ff_15566:FAff port map(x=>p(370)(107),y=>p(371)(107),Cin=>p(372)(107),clock=>clock,reset=>reset,s=>p(377)(107),cout=>p(378)(108));
FA_ff_15567:FAff port map(x=>p(370)(108),y=>p(371)(108),Cin=>p(372)(108),clock=>clock,reset=>reset,s=>p(377)(108),cout=>p(378)(109));
FA_ff_15568:FAff port map(x=>p(370)(109),y=>p(371)(109),Cin=>p(372)(109),clock=>clock,reset=>reset,s=>p(377)(109),cout=>p(378)(110));
FA_ff_15569:FAff port map(x=>p(370)(110),y=>p(371)(110),Cin=>p(372)(110),clock=>clock,reset=>reset,s=>p(377)(110),cout=>p(378)(111));
FA_ff_15570:FAff port map(x=>p(370)(111),y=>p(371)(111),Cin=>p(372)(111),clock=>clock,reset=>reset,s=>p(377)(111),cout=>p(378)(112));
FA_ff_15571:FAff port map(x=>p(370)(112),y=>p(371)(112),Cin=>p(372)(112),clock=>clock,reset=>reset,s=>p(377)(112),cout=>p(378)(113));
FA_ff_15572:FAff port map(x=>p(370)(113),y=>p(371)(113),Cin=>p(372)(113),clock=>clock,reset=>reset,s=>p(377)(113),cout=>p(378)(114));
FA_ff_15573:FAff port map(x=>p(370)(114),y=>p(371)(114),Cin=>p(372)(114),clock=>clock,reset=>reset,s=>p(377)(114),cout=>p(378)(115));
FA_ff_15574:FAff port map(x=>p(370)(115),y=>p(371)(115),Cin=>p(372)(115),clock=>clock,reset=>reset,s=>p(377)(115),cout=>p(378)(116));
FA_ff_15575:FAff port map(x=>p(370)(116),y=>p(371)(116),Cin=>p(372)(116),clock=>clock,reset=>reset,s=>p(377)(116),cout=>p(378)(117));
FA_ff_15576:FAff port map(x=>p(370)(117),y=>p(371)(117),Cin=>p(372)(117),clock=>clock,reset=>reset,s=>p(377)(117),cout=>p(378)(118));
FA_ff_15577:FAff port map(x=>p(370)(118),y=>p(371)(118),Cin=>p(372)(118),clock=>clock,reset=>reset,s=>p(377)(118),cout=>p(378)(119));
FA_ff_15578:FAff port map(x=>p(370)(119),y=>p(371)(119),Cin=>p(372)(119),clock=>clock,reset=>reset,s=>p(377)(119),cout=>p(378)(120));
FA_ff_15579:FAff port map(x=>p(370)(120),y=>p(371)(120),Cin=>p(372)(120),clock=>clock,reset=>reset,s=>p(377)(120),cout=>p(378)(121));
FA_ff_15580:FAff port map(x=>p(370)(121),y=>p(371)(121),Cin=>p(372)(121),clock=>clock,reset=>reset,s=>p(377)(121),cout=>p(378)(122));
FA_ff_15581:FAff port map(x=>p(370)(122),y=>p(371)(122),Cin=>p(372)(122),clock=>clock,reset=>reset,s=>p(377)(122),cout=>p(378)(123));
FA_ff_15582:FAff port map(x=>p(370)(123),y=>p(371)(123),Cin=>p(372)(123),clock=>clock,reset=>reset,s=>p(377)(123),cout=>p(378)(124));
FA_ff_15583:FAff port map(x=>p(370)(124),y=>p(371)(124),Cin=>p(372)(124),clock=>clock,reset=>reset,s=>p(377)(124),cout=>p(378)(125));
FA_ff_15584:FAff port map(x=>p(370)(125),y=>p(371)(125),Cin=>p(372)(125),clock=>clock,reset=>reset,s=>p(377)(125),cout=>p(378)(126));
FA_ff_15585:FAff port map(x=>p(370)(126),y=>p(371)(126),Cin=>p(372)(126),clock=>clock,reset=>reset,s=>p(377)(126),cout=>p(378)(127));
FA_ff_15586:FAff port map(x=>p(370)(127),y=>p(371)(127),Cin=>p(372)(127),clock=>clock,reset=>reset,s=>p(377)(127),cout=>p(378)(128));
FA_ff_15587:FAff port map(x=>p(370)(128),y=>p(371)(128),Cin=>p(372)(128),clock=>clock,reset=>reset,s=>p(377)(128),cout=>p(378)(129));
FA_ff_15588:FAff port map(x=>p(370)(129),y=>p(371)(129),Cin=>p(372)(129),clock=>clock,reset=>reset,s=>p(377)(129),cout=>p(378)(130));
FA_ff_15589:FAff port map(x=>p(370)(130),y=>p(371)(130),Cin=>p(372)(130),clock=>clock,reset=>reset,s=>p(377)(130),cout=>p(378)(131));
FA_ff_15590:FAff port map(x=>p(370)(131),y=>p(371)(131),Cin=>p(372)(131),clock=>clock,reset=>reset,s=>p(377)(131),cout=>p(378)(132));
HA_ff_107:HAff port map(x=>p(370)(132),y=>p(372)(132),clock=>clock,reset=>reset,s=>p(377)(132),c=>p(378)(133));
p(379)(0)<=p(373)(0);
p(379)(1)<=p(373)(1);
p(379)(2)<=p(373)(2);
p(379)(3)<=p(373)(3);
p(379)(4)<=p(373)(4);
p(379)(5)<=p(373)(5);
p(379)(6)<=p(373)(6);
p(379)(7)<=p(373)(7);
p(379)(8)<=p(373)(8);
p(379)(9)<=p(373)(9);
p(379)(10)<=p(373)(10);
p(379)(11)<=p(373)(11);
p(379)(12)<=p(373)(12);
p(379)(13)<=p(373)(13);
p(379)(14)<=p(373)(14);
p(379)(15)<=p(373)(15);
p(379)(16)<=p(373)(16);
p(379)(17)<=p(373)(17);
p(379)(18)<=p(373)(18);
p(379)(19)<=p(373)(19);
p(379)(20)<=p(373)(20);
p(379)(21)<=p(373)(21);
p(379)(22)<=p(373)(22);
p(379)(23)<=p(373)(23);
p(379)(24)<=p(373)(24);
p(379)(25)<=p(373)(25);
p(379)(26)<=p(373)(26);
p(379)(27)<=p(373)(27);
p(379)(28)<=p(373)(28);
p(379)(29)<=p(373)(29);
p(379)(30)<=p(373)(30);
p(379)(31)<=p(373)(31);
p(379)(32)<=p(373)(32);
p(379)(33)<=p(373)(33);
p(379)(34)<=p(373)(34);
p(379)(35)<=p(373)(35);
p(379)(36)<=p(373)(36);
p(379)(37)<=p(373)(37);
p(379)(38)<=p(373)(38);
p(379)(39)<=p(373)(39);
p(379)(40)<=p(373)(40);
p(379)(41)<=p(373)(41);
p(379)(42)<=p(373)(42);
p(379)(43)<=p(373)(43);
p(379)(44)<=p(373)(44);
p(379)(45)<=p(373)(45);
p(379)(46)<=p(373)(46);
p(379)(47)<=p(373)(47);
p(379)(48)<=p(373)(48);
p(379)(49)<=p(373)(49);
p(379)(50)<=p(373)(50);
p(379)(51)<=p(373)(51);
p(379)(52)<=p(373)(52);
p(379)(53)<=p(373)(53);
p(379)(54)<=p(373)(54);
p(379)(55)<=p(373)(55);
p(379)(56)<=p(373)(56);
p(379)(57)<=p(373)(57);
p(379)(58)<=p(373)(58);
p(379)(59)<=p(373)(59);
p(379)(60)<=p(373)(60);
p(379)(61)<=p(373)(61);
p(379)(62)<=p(373)(62);
p(379)(63)<=p(373)(63);
p(379)(64)<=p(373)(64);
p(379)(65)<=p(373)(65);
p(379)(66)<=p(373)(66);
p(379)(67)<=p(373)(67);
p(379)(68)<=p(373)(68);
p(379)(69)<=p(373)(69);
p(379)(70)<=p(373)(70);
p(379)(71)<=p(373)(71);
p(379)(72)<=p(373)(72);
p(379)(73)<=p(373)(73);
p(379)(74)<=p(373)(74);
p(379)(75)<=p(373)(75);
p(379)(76)<=p(373)(76);
p(379)(77)<=p(373)(77);
p(379)(78)<=p(373)(78);
p(379)(79)<=p(373)(79);
p(379)(80)<=p(373)(80);
p(379)(81)<=p(373)(81);
p(379)(82)<=p(373)(82);
p(379)(83)<=p(373)(83);
p(379)(84)<=p(373)(84);
p(379)(85)<=p(373)(85);
p(379)(86)<=p(373)(86);
p(379)(87)<=p(373)(87);
p(379)(88)<=p(373)(88);
p(379)(89)<=p(373)(89);
p(379)(90)<=p(373)(90);
p(379)(91)<=p(373)(91);
p(379)(92)<=p(373)(92);
p(379)(93)<=p(373)(93);
p(379)(94)<=p(373)(94);
p(379)(95)<=p(373)(95);
p(379)(96)<=p(373)(96);
p(379)(97)<=p(373)(97);
p(379)(98)<=p(373)(98);
p(379)(99)<=p(373)(99);
p(379)(100)<=p(373)(100);
p(379)(101)<=p(373)(101);
p(379)(102)<=p(373)(102);
p(379)(103)<=p(373)(103);
p(379)(104)<=p(373)(104);
p(379)(105)<=p(373)(105);
p(379)(106)<=p(373)(106);
p(379)(107)<=p(373)(107);
p(379)(108)<=p(373)(108);
p(379)(109)<=p(373)(109);
p(379)(110)<=p(373)(110);
p(379)(111)<=p(373)(111);
p(379)(112)<=p(373)(112);
p(379)(113)<=p(373)(113);
p(379)(114)<=p(373)(114);
p(379)(115)<=p(373)(115);
p(379)(116)<=p(373)(116);
p(379)(117)<=p(373)(117);
p(379)(118)<=p(373)(118);
p(379)(119)<=p(373)(119);
p(379)(120)<=p(373)(120);
p(379)(121)<=p(373)(121);
p(379)(122)<=p(373)(122);
p(379)(123)<=p(373)(123);
p(379)(124)<=p(373)(124);
p(379)(125)<=p(373)(125);
p(379)(126)<=p(373)(126);
p(379)(127)<=p(373)(127);
p(379)(128)<=p(373)(128);
p(379)(129)<=p(373)(129);
p(379)(130)<=p(373)(130);
p(379)(131)<=p(373)(131);
p(379)(132)<=p(373)(132);
p(379)(133)<=p(373)(133);
p(379)(134)<=p(373)(134);
p(380)(0)<=p(374)(0);
p(380)(1)<=p(374)(1);
p(380)(2)<=p(374)(2);
p(380)(3)<=p(374)(3);
p(380)(4)<=p(374)(4);
p(380)(5)<=p(374)(5);
p(380)(6)<=p(374)(6);
p(380)(7)<=p(374)(7);
p(380)(8)<=p(374)(8);
p(380)(9)<=p(374)(9);
p(380)(10)<=p(374)(10);
p(380)(11)<=p(374)(11);
p(380)(12)<=p(374)(12);
p(380)(13)<=p(374)(13);
p(380)(14)<=p(374)(14);
p(380)(15)<=p(374)(15);
p(380)(16)<=p(374)(16);
p(380)(17)<=p(374)(17);
p(380)(18)<=p(374)(18);
p(380)(19)<=p(374)(19);
p(380)(20)<=p(374)(20);
p(380)(21)<=p(374)(21);
p(380)(22)<=p(374)(22);
p(380)(23)<=p(374)(23);
p(380)(24)<=p(374)(24);
p(380)(25)<=p(374)(25);
p(380)(26)<=p(374)(26);
p(380)(27)<=p(374)(27);
p(380)(28)<=p(374)(28);
p(380)(29)<=p(374)(29);
p(380)(30)<=p(374)(30);
p(380)(31)<=p(374)(31);
p(380)(32)<=p(374)(32);
p(380)(33)<=p(374)(33);
p(380)(34)<=p(374)(34);
p(380)(35)<=p(374)(35);
p(380)(36)<=p(374)(36);
p(380)(37)<=p(374)(37);
p(380)(38)<=p(374)(38);
p(380)(39)<=p(374)(39);
p(380)(40)<=p(374)(40);
p(380)(41)<=p(374)(41);
p(380)(42)<=p(374)(42);
p(380)(43)<=p(374)(43);
p(380)(44)<=p(374)(44);
p(380)(45)<=p(374)(45);
p(380)(46)<=p(374)(46);
p(380)(47)<=p(374)(47);
p(380)(48)<=p(374)(48);
p(380)(49)<=p(374)(49);
p(380)(50)<=p(374)(50);
p(380)(51)<=p(374)(51);
p(380)(52)<=p(374)(52);
p(380)(53)<=p(374)(53);
p(380)(54)<=p(374)(54);
p(380)(55)<=p(374)(55);
p(380)(56)<=p(374)(56);
p(380)(57)<=p(374)(57);
p(380)(58)<=p(374)(58);
p(380)(59)<=p(374)(59);
p(380)(60)<=p(374)(60);
p(380)(61)<=p(374)(61);
p(380)(62)<=p(374)(62);
p(380)(63)<=p(374)(63);
p(380)(64)<=p(374)(64);
p(380)(65)<=p(374)(65);
p(380)(66)<=p(374)(66);
p(380)(67)<=p(374)(67);
p(380)(68)<=p(374)(68);
p(380)(69)<=p(374)(69);
p(380)(70)<=p(374)(70);
p(380)(71)<=p(374)(71);
p(380)(72)<=p(374)(72);
p(380)(73)<=p(374)(73);
p(380)(74)<=p(374)(74);
p(380)(75)<=p(374)(75);
p(380)(76)<=p(374)(76);
p(380)(77)<=p(374)(77);
p(380)(78)<=p(374)(78);
p(380)(79)<=p(374)(79);
p(380)(80)<=p(374)(80);
p(380)(81)<=p(374)(81);
p(380)(82)<=p(374)(82);
p(380)(83)<=p(374)(83);
p(380)(84)<=p(374)(84);
p(380)(85)<=p(374)(85);
p(380)(86)<=p(374)(86);
p(380)(87)<=p(374)(87);
p(380)(88)<=p(374)(88);
p(380)(89)<=p(374)(89);
p(380)(90)<=p(374)(90);
p(380)(91)<=p(374)(91);
p(380)(92)<=p(374)(92);
p(380)(93)<=p(374)(93);
p(380)(94)<=p(374)(94);
p(380)(95)<=p(374)(95);
p(380)(96)<=p(374)(96);
p(380)(97)<=p(374)(97);
p(380)(98)<=p(374)(98);
p(380)(99)<=p(374)(99);
p(380)(100)<=p(374)(100);
p(380)(101)<=p(374)(101);
p(380)(102)<=p(374)(102);
p(380)(103)<=p(374)(103);
p(380)(104)<=p(374)(104);
p(380)(105)<=p(374)(105);
p(380)(106)<=p(374)(106);
p(380)(107)<=p(374)(107);
p(380)(108)<=p(374)(108);
p(380)(109)<=p(374)(109);
p(380)(110)<=p(374)(110);
p(380)(111)<=p(374)(111);
p(380)(112)<=p(374)(112);
p(380)(113)<=p(374)(113);
p(380)(114)<=p(374)(114);
p(380)(115)<=p(374)(115);
p(380)(116)<=p(374)(116);
p(380)(117)<=p(374)(117);
p(380)(118)<=p(374)(118);
p(380)(119)<=p(374)(119);
p(380)(120)<=p(374)(120);
p(380)(121)<=p(374)(121);
p(380)(122)<=p(374)(122);
p(380)(123)<=p(374)(123);
p(380)(124)<=p(374)(124);
p(380)(125)<=p(374)(125);
p(380)(126)<=p(374)(126);
p(380)(127)<=p(374)(127);
p(380)(128)<=p(374)(128);
p(380)(129)<=p(374)(129);
p(380)(130)<=p(374)(130);
p(380)(131)<=p(374)(131);
p(380)(132)<=p(374)(132);
p(380)(133)<=p(374)(133);
p(380)(134)<=p(374)(134);
HA_ff_108:HAff port map(x=>p(375)(0),y=>p(377)(0),clock=>clock,reset=>reset,s=>p(381)(0),c=>p(382)(1));
FA_ff_15591:FAff port map(x=>p(375)(1),y=>p(376)(1),Cin=>p(377)(1),clock=>clock,reset=>reset,s=>p(381)(1),cout=>p(382)(2));
FA_ff_15592:FAff port map(x=>p(375)(2),y=>p(376)(2),Cin=>p(377)(2),clock=>clock,reset=>reset,s=>p(381)(2),cout=>p(382)(3));
FA_ff_15593:FAff port map(x=>p(375)(3),y=>p(376)(3),Cin=>p(377)(3),clock=>clock,reset=>reset,s=>p(381)(3),cout=>p(382)(4));
FA_ff_15594:FAff port map(x=>p(375)(4),y=>p(376)(4),Cin=>p(377)(4),clock=>clock,reset=>reset,s=>p(381)(4),cout=>p(382)(5));
FA_ff_15595:FAff port map(x=>p(375)(5),y=>p(376)(5),Cin=>p(377)(5),clock=>clock,reset=>reset,s=>p(381)(5),cout=>p(382)(6));
FA_ff_15596:FAff port map(x=>p(375)(6),y=>p(376)(6),Cin=>p(377)(6),clock=>clock,reset=>reset,s=>p(381)(6),cout=>p(382)(7));
FA_ff_15597:FAff port map(x=>p(375)(7),y=>p(376)(7),Cin=>p(377)(7),clock=>clock,reset=>reset,s=>p(381)(7),cout=>p(382)(8));
FA_ff_15598:FAff port map(x=>p(375)(8),y=>p(376)(8),Cin=>p(377)(8),clock=>clock,reset=>reset,s=>p(381)(8),cout=>p(382)(9));
FA_ff_15599:FAff port map(x=>p(375)(9),y=>p(376)(9),Cin=>p(377)(9),clock=>clock,reset=>reset,s=>p(381)(9),cout=>p(382)(10));
FA_ff_15600:FAff port map(x=>p(375)(10),y=>p(376)(10),Cin=>p(377)(10),clock=>clock,reset=>reset,s=>p(381)(10),cout=>p(382)(11));
FA_ff_15601:FAff port map(x=>p(375)(11),y=>p(376)(11),Cin=>p(377)(11),clock=>clock,reset=>reset,s=>p(381)(11),cout=>p(382)(12));
FA_ff_15602:FAff port map(x=>p(375)(12),y=>p(376)(12),Cin=>p(377)(12),clock=>clock,reset=>reset,s=>p(381)(12),cout=>p(382)(13));
FA_ff_15603:FAff port map(x=>p(375)(13),y=>p(376)(13),Cin=>p(377)(13),clock=>clock,reset=>reset,s=>p(381)(13),cout=>p(382)(14));
FA_ff_15604:FAff port map(x=>p(375)(14),y=>p(376)(14),Cin=>p(377)(14),clock=>clock,reset=>reset,s=>p(381)(14),cout=>p(382)(15));
FA_ff_15605:FAff port map(x=>p(375)(15),y=>p(376)(15),Cin=>p(377)(15),clock=>clock,reset=>reset,s=>p(381)(15),cout=>p(382)(16));
FA_ff_15606:FAff port map(x=>p(375)(16),y=>p(376)(16),Cin=>p(377)(16),clock=>clock,reset=>reset,s=>p(381)(16),cout=>p(382)(17));
FA_ff_15607:FAff port map(x=>p(375)(17),y=>p(376)(17),Cin=>p(377)(17),clock=>clock,reset=>reset,s=>p(381)(17),cout=>p(382)(18));
FA_ff_15608:FAff port map(x=>p(375)(18),y=>p(376)(18),Cin=>p(377)(18),clock=>clock,reset=>reset,s=>p(381)(18),cout=>p(382)(19));
FA_ff_15609:FAff port map(x=>p(375)(19),y=>p(376)(19),Cin=>p(377)(19),clock=>clock,reset=>reset,s=>p(381)(19),cout=>p(382)(20));
FA_ff_15610:FAff port map(x=>p(375)(20),y=>p(376)(20),Cin=>p(377)(20),clock=>clock,reset=>reset,s=>p(381)(20),cout=>p(382)(21));
FA_ff_15611:FAff port map(x=>p(375)(21),y=>p(376)(21),Cin=>p(377)(21),clock=>clock,reset=>reset,s=>p(381)(21),cout=>p(382)(22));
FA_ff_15612:FAff port map(x=>p(375)(22),y=>p(376)(22),Cin=>p(377)(22),clock=>clock,reset=>reset,s=>p(381)(22),cout=>p(382)(23));
FA_ff_15613:FAff port map(x=>p(375)(23),y=>p(376)(23),Cin=>p(377)(23),clock=>clock,reset=>reset,s=>p(381)(23),cout=>p(382)(24));
FA_ff_15614:FAff port map(x=>p(375)(24),y=>p(376)(24),Cin=>p(377)(24),clock=>clock,reset=>reset,s=>p(381)(24),cout=>p(382)(25));
FA_ff_15615:FAff port map(x=>p(375)(25),y=>p(376)(25),Cin=>p(377)(25),clock=>clock,reset=>reset,s=>p(381)(25),cout=>p(382)(26));
FA_ff_15616:FAff port map(x=>p(375)(26),y=>p(376)(26),Cin=>p(377)(26),clock=>clock,reset=>reset,s=>p(381)(26),cout=>p(382)(27));
FA_ff_15617:FAff port map(x=>p(375)(27),y=>p(376)(27),Cin=>p(377)(27),clock=>clock,reset=>reset,s=>p(381)(27),cout=>p(382)(28));
FA_ff_15618:FAff port map(x=>p(375)(28),y=>p(376)(28),Cin=>p(377)(28),clock=>clock,reset=>reset,s=>p(381)(28),cout=>p(382)(29));
FA_ff_15619:FAff port map(x=>p(375)(29),y=>p(376)(29),Cin=>p(377)(29),clock=>clock,reset=>reset,s=>p(381)(29),cout=>p(382)(30));
FA_ff_15620:FAff port map(x=>p(375)(30),y=>p(376)(30),Cin=>p(377)(30),clock=>clock,reset=>reset,s=>p(381)(30),cout=>p(382)(31));
FA_ff_15621:FAff port map(x=>p(375)(31),y=>p(376)(31),Cin=>p(377)(31),clock=>clock,reset=>reset,s=>p(381)(31),cout=>p(382)(32));
FA_ff_15622:FAff port map(x=>p(375)(32),y=>p(376)(32),Cin=>p(377)(32),clock=>clock,reset=>reset,s=>p(381)(32),cout=>p(382)(33));
FA_ff_15623:FAff port map(x=>p(375)(33),y=>p(376)(33),Cin=>p(377)(33),clock=>clock,reset=>reset,s=>p(381)(33),cout=>p(382)(34));
FA_ff_15624:FAff port map(x=>p(375)(34),y=>p(376)(34),Cin=>p(377)(34),clock=>clock,reset=>reset,s=>p(381)(34),cout=>p(382)(35));
FA_ff_15625:FAff port map(x=>p(375)(35),y=>p(376)(35),Cin=>p(377)(35),clock=>clock,reset=>reset,s=>p(381)(35),cout=>p(382)(36));
FA_ff_15626:FAff port map(x=>p(375)(36),y=>p(376)(36),Cin=>p(377)(36),clock=>clock,reset=>reset,s=>p(381)(36),cout=>p(382)(37));
FA_ff_15627:FAff port map(x=>p(375)(37),y=>p(376)(37),Cin=>p(377)(37),clock=>clock,reset=>reset,s=>p(381)(37),cout=>p(382)(38));
FA_ff_15628:FAff port map(x=>p(375)(38),y=>p(376)(38),Cin=>p(377)(38),clock=>clock,reset=>reset,s=>p(381)(38),cout=>p(382)(39));
FA_ff_15629:FAff port map(x=>p(375)(39),y=>p(376)(39),Cin=>p(377)(39),clock=>clock,reset=>reset,s=>p(381)(39),cout=>p(382)(40));
FA_ff_15630:FAff port map(x=>p(375)(40),y=>p(376)(40),Cin=>p(377)(40),clock=>clock,reset=>reset,s=>p(381)(40),cout=>p(382)(41));
FA_ff_15631:FAff port map(x=>p(375)(41),y=>p(376)(41),Cin=>p(377)(41),clock=>clock,reset=>reset,s=>p(381)(41),cout=>p(382)(42));
FA_ff_15632:FAff port map(x=>p(375)(42),y=>p(376)(42),Cin=>p(377)(42),clock=>clock,reset=>reset,s=>p(381)(42),cout=>p(382)(43));
FA_ff_15633:FAff port map(x=>p(375)(43),y=>p(376)(43),Cin=>p(377)(43),clock=>clock,reset=>reset,s=>p(381)(43),cout=>p(382)(44));
FA_ff_15634:FAff port map(x=>p(375)(44),y=>p(376)(44),Cin=>p(377)(44),clock=>clock,reset=>reset,s=>p(381)(44),cout=>p(382)(45));
FA_ff_15635:FAff port map(x=>p(375)(45),y=>p(376)(45),Cin=>p(377)(45),clock=>clock,reset=>reset,s=>p(381)(45),cout=>p(382)(46));
FA_ff_15636:FAff port map(x=>p(375)(46),y=>p(376)(46),Cin=>p(377)(46),clock=>clock,reset=>reset,s=>p(381)(46),cout=>p(382)(47));
FA_ff_15637:FAff port map(x=>p(375)(47),y=>p(376)(47),Cin=>p(377)(47),clock=>clock,reset=>reset,s=>p(381)(47),cout=>p(382)(48));
FA_ff_15638:FAff port map(x=>p(375)(48),y=>p(376)(48),Cin=>p(377)(48),clock=>clock,reset=>reset,s=>p(381)(48),cout=>p(382)(49));
FA_ff_15639:FAff port map(x=>p(375)(49),y=>p(376)(49),Cin=>p(377)(49),clock=>clock,reset=>reset,s=>p(381)(49),cout=>p(382)(50));
FA_ff_15640:FAff port map(x=>p(375)(50),y=>p(376)(50),Cin=>p(377)(50),clock=>clock,reset=>reset,s=>p(381)(50),cout=>p(382)(51));
FA_ff_15641:FAff port map(x=>p(375)(51),y=>p(376)(51),Cin=>p(377)(51),clock=>clock,reset=>reset,s=>p(381)(51),cout=>p(382)(52));
FA_ff_15642:FAff port map(x=>p(375)(52),y=>p(376)(52),Cin=>p(377)(52),clock=>clock,reset=>reset,s=>p(381)(52),cout=>p(382)(53));
FA_ff_15643:FAff port map(x=>p(375)(53),y=>p(376)(53),Cin=>p(377)(53),clock=>clock,reset=>reset,s=>p(381)(53),cout=>p(382)(54));
FA_ff_15644:FAff port map(x=>p(375)(54),y=>p(376)(54),Cin=>p(377)(54),clock=>clock,reset=>reset,s=>p(381)(54),cout=>p(382)(55));
FA_ff_15645:FAff port map(x=>p(375)(55),y=>p(376)(55),Cin=>p(377)(55),clock=>clock,reset=>reset,s=>p(381)(55),cout=>p(382)(56));
FA_ff_15646:FAff port map(x=>p(375)(56),y=>p(376)(56),Cin=>p(377)(56),clock=>clock,reset=>reset,s=>p(381)(56),cout=>p(382)(57));
FA_ff_15647:FAff port map(x=>p(375)(57),y=>p(376)(57),Cin=>p(377)(57),clock=>clock,reset=>reset,s=>p(381)(57),cout=>p(382)(58));
FA_ff_15648:FAff port map(x=>p(375)(58),y=>p(376)(58),Cin=>p(377)(58),clock=>clock,reset=>reset,s=>p(381)(58),cout=>p(382)(59));
FA_ff_15649:FAff port map(x=>p(375)(59),y=>p(376)(59),Cin=>p(377)(59),clock=>clock,reset=>reset,s=>p(381)(59),cout=>p(382)(60));
FA_ff_15650:FAff port map(x=>p(375)(60),y=>p(376)(60),Cin=>p(377)(60),clock=>clock,reset=>reset,s=>p(381)(60),cout=>p(382)(61));
FA_ff_15651:FAff port map(x=>p(375)(61),y=>p(376)(61),Cin=>p(377)(61),clock=>clock,reset=>reset,s=>p(381)(61),cout=>p(382)(62));
FA_ff_15652:FAff port map(x=>p(375)(62),y=>p(376)(62),Cin=>p(377)(62),clock=>clock,reset=>reset,s=>p(381)(62),cout=>p(382)(63));
FA_ff_15653:FAff port map(x=>p(375)(63),y=>p(376)(63),Cin=>p(377)(63),clock=>clock,reset=>reset,s=>p(381)(63),cout=>p(382)(64));
FA_ff_15654:FAff port map(x=>p(375)(64),y=>p(376)(64),Cin=>p(377)(64),clock=>clock,reset=>reset,s=>p(381)(64),cout=>p(382)(65));
FA_ff_15655:FAff port map(x=>p(375)(65),y=>p(376)(65),Cin=>p(377)(65),clock=>clock,reset=>reset,s=>p(381)(65),cout=>p(382)(66));
FA_ff_15656:FAff port map(x=>p(375)(66),y=>p(376)(66),Cin=>p(377)(66),clock=>clock,reset=>reset,s=>p(381)(66),cout=>p(382)(67));
FA_ff_15657:FAff port map(x=>p(375)(67),y=>p(376)(67),Cin=>p(377)(67),clock=>clock,reset=>reset,s=>p(381)(67),cout=>p(382)(68));
FA_ff_15658:FAff port map(x=>p(375)(68),y=>p(376)(68),Cin=>p(377)(68),clock=>clock,reset=>reset,s=>p(381)(68),cout=>p(382)(69));
FA_ff_15659:FAff port map(x=>p(375)(69),y=>p(376)(69),Cin=>p(377)(69),clock=>clock,reset=>reset,s=>p(381)(69),cout=>p(382)(70));
FA_ff_15660:FAff port map(x=>p(375)(70),y=>p(376)(70),Cin=>p(377)(70),clock=>clock,reset=>reset,s=>p(381)(70),cout=>p(382)(71));
FA_ff_15661:FAff port map(x=>p(375)(71),y=>p(376)(71),Cin=>p(377)(71),clock=>clock,reset=>reset,s=>p(381)(71),cout=>p(382)(72));
FA_ff_15662:FAff port map(x=>p(375)(72),y=>p(376)(72),Cin=>p(377)(72),clock=>clock,reset=>reset,s=>p(381)(72),cout=>p(382)(73));
FA_ff_15663:FAff port map(x=>p(375)(73),y=>p(376)(73),Cin=>p(377)(73),clock=>clock,reset=>reset,s=>p(381)(73),cout=>p(382)(74));
FA_ff_15664:FAff port map(x=>p(375)(74),y=>p(376)(74),Cin=>p(377)(74),clock=>clock,reset=>reset,s=>p(381)(74),cout=>p(382)(75));
FA_ff_15665:FAff port map(x=>p(375)(75),y=>p(376)(75),Cin=>p(377)(75),clock=>clock,reset=>reset,s=>p(381)(75),cout=>p(382)(76));
FA_ff_15666:FAff port map(x=>p(375)(76),y=>p(376)(76),Cin=>p(377)(76),clock=>clock,reset=>reset,s=>p(381)(76),cout=>p(382)(77));
FA_ff_15667:FAff port map(x=>p(375)(77),y=>p(376)(77),Cin=>p(377)(77),clock=>clock,reset=>reset,s=>p(381)(77),cout=>p(382)(78));
FA_ff_15668:FAff port map(x=>p(375)(78),y=>p(376)(78),Cin=>p(377)(78),clock=>clock,reset=>reset,s=>p(381)(78),cout=>p(382)(79));
FA_ff_15669:FAff port map(x=>p(375)(79),y=>p(376)(79),Cin=>p(377)(79),clock=>clock,reset=>reset,s=>p(381)(79),cout=>p(382)(80));
FA_ff_15670:FAff port map(x=>p(375)(80),y=>p(376)(80),Cin=>p(377)(80),clock=>clock,reset=>reset,s=>p(381)(80),cout=>p(382)(81));
FA_ff_15671:FAff port map(x=>p(375)(81),y=>p(376)(81),Cin=>p(377)(81),clock=>clock,reset=>reset,s=>p(381)(81),cout=>p(382)(82));
FA_ff_15672:FAff port map(x=>p(375)(82),y=>p(376)(82),Cin=>p(377)(82),clock=>clock,reset=>reset,s=>p(381)(82),cout=>p(382)(83));
FA_ff_15673:FAff port map(x=>p(375)(83),y=>p(376)(83),Cin=>p(377)(83),clock=>clock,reset=>reset,s=>p(381)(83),cout=>p(382)(84));
FA_ff_15674:FAff port map(x=>p(375)(84),y=>p(376)(84),Cin=>p(377)(84),clock=>clock,reset=>reset,s=>p(381)(84),cout=>p(382)(85));
FA_ff_15675:FAff port map(x=>p(375)(85),y=>p(376)(85),Cin=>p(377)(85),clock=>clock,reset=>reset,s=>p(381)(85),cout=>p(382)(86));
FA_ff_15676:FAff port map(x=>p(375)(86),y=>p(376)(86),Cin=>p(377)(86),clock=>clock,reset=>reset,s=>p(381)(86),cout=>p(382)(87));
FA_ff_15677:FAff port map(x=>p(375)(87),y=>p(376)(87),Cin=>p(377)(87),clock=>clock,reset=>reset,s=>p(381)(87),cout=>p(382)(88));
FA_ff_15678:FAff port map(x=>p(375)(88),y=>p(376)(88),Cin=>p(377)(88),clock=>clock,reset=>reset,s=>p(381)(88),cout=>p(382)(89));
FA_ff_15679:FAff port map(x=>p(375)(89),y=>p(376)(89),Cin=>p(377)(89),clock=>clock,reset=>reset,s=>p(381)(89),cout=>p(382)(90));
FA_ff_15680:FAff port map(x=>p(375)(90),y=>p(376)(90),Cin=>p(377)(90),clock=>clock,reset=>reset,s=>p(381)(90),cout=>p(382)(91));
FA_ff_15681:FAff port map(x=>p(375)(91),y=>p(376)(91),Cin=>p(377)(91),clock=>clock,reset=>reset,s=>p(381)(91),cout=>p(382)(92));
FA_ff_15682:FAff port map(x=>p(375)(92),y=>p(376)(92),Cin=>p(377)(92),clock=>clock,reset=>reset,s=>p(381)(92),cout=>p(382)(93));
FA_ff_15683:FAff port map(x=>p(375)(93),y=>p(376)(93),Cin=>p(377)(93),clock=>clock,reset=>reset,s=>p(381)(93),cout=>p(382)(94));
FA_ff_15684:FAff port map(x=>p(375)(94),y=>p(376)(94),Cin=>p(377)(94),clock=>clock,reset=>reset,s=>p(381)(94),cout=>p(382)(95));
FA_ff_15685:FAff port map(x=>p(375)(95),y=>p(376)(95),Cin=>p(377)(95),clock=>clock,reset=>reset,s=>p(381)(95),cout=>p(382)(96));
FA_ff_15686:FAff port map(x=>p(375)(96),y=>p(376)(96),Cin=>p(377)(96),clock=>clock,reset=>reset,s=>p(381)(96),cout=>p(382)(97));
FA_ff_15687:FAff port map(x=>p(375)(97),y=>p(376)(97),Cin=>p(377)(97),clock=>clock,reset=>reset,s=>p(381)(97),cout=>p(382)(98));
FA_ff_15688:FAff port map(x=>p(375)(98),y=>p(376)(98),Cin=>p(377)(98),clock=>clock,reset=>reset,s=>p(381)(98),cout=>p(382)(99));
FA_ff_15689:FAff port map(x=>p(375)(99),y=>p(376)(99),Cin=>p(377)(99),clock=>clock,reset=>reset,s=>p(381)(99),cout=>p(382)(100));
FA_ff_15690:FAff port map(x=>p(375)(100),y=>p(376)(100),Cin=>p(377)(100),clock=>clock,reset=>reset,s=>p(381)(100),cout=>p(382)(101));
FA_ff_15691:FAff port map(x=>p(375)(101),y=>p(376)(101),Cin=>p(377)(101),clock=>clock,reset=>reset,s=>p(381)(101),cout=>p(382)(102));
FA_ff_15692:FAff port map(x=>p(375)(102),y=>p(376)(102),Cin=>p(377)(102),clock=>clock,reset=>reset,s=>p(381)(102),cout=>p(382)(103));
FA_ff_15693:FAff port map(x=>p(375)(103),y=>p(376)(103),Cin=>p(377)(103),clock=>clock,reset=>reset,s=>p(381)(103),cout=>p(382)(104));
FA_ff_15694:FAff port map(x=>p(375)(104),y=>p(376)(104),Cin=>p(377)(104),clock=>clock,reset=>reset,s=>p(381)(104),cout=>p(382)(105));
FA_ff_15695:FAff port map(x=>p(375)(105),y=>p(376)(105),Cin=>p(377)(105),clock=>clock,reset=>reset,s=>p(381)(105),cout=>p(382)(106));
FA_ff_15696:FAff port map(x=>p(375)(106),y=>p(376)(106),Cin=>p(377)(106),clock=>clock,reset=>reset,s=>p(381)(106),cout=>p(382)(107));
FA_ff_15697:FAff port map(x=>p(375)(107),y=>p(376)(107),Cin=>p(377)(107),clock=>clock,reset=>reset,s=>p(381)(107),cout=>p(382)(108));
FA_ff_15698:FAff port map(x=>p(375)(108),y=>p(376)(108),Cin=>p(377)(108),clock=>clock,reset=>reset,s=>p(381)(108),cout=>p(382)(109));
FA_ff_15699:FAff port map(x=>p(375)(109),y=>p(376)(109),Cin=>p(377)(109),clock=>clock,reset=>reset,s=>p(381)(109),cout=>p(382)(110));
FA_ff_15700:FAff port map(x=>p(375)(110),y=>p(376)(110),Cin=>p(377)(110),clock=>clock,reset=>reset,s=>p(381)(110),cout=>p(382)(111));
FA_ff_15701:FAff port map(x=>p(375)(111),y=>p(376)(111),Cin=>p(377)(111),clock=>clock,reset=>reset,s=>p(381)(111),cout=>p(382)(112));
FA_ff_15702:FAff port map(x=>p(375)(112),y=>p(376)(112),Cin=>p(377)(112),clock=>clock,reset=>reset,s=>p(381)(112),cout=>p(382)(113));
FA_ff_15703:FAff port map(x=>p(375)(113),y=>p(376)(113),Cin=>p(377)(113),clock=>clock,reset=>reset,s=>p(381)(113),cout=>p(382)(114));
FA_ff_15704:FAff port map(x=>p(375)(114),y=>p(376)(114),Cin=>p(377)(114),clock=>clock,reset=>reset,s=>p(381)(114),cout=>p(382)(115));
FA_ff_15705:FAff port map(x=>p(375)(115),y=>p(376)(115),Cin=>p(377)(115),clock=>clock,reset=>reset,s=>p(381)(115),cout=>p(382)(116));
FA_ff_15706:FAff port map(x=>p(375)(116),y=>p(376)(116),Cin=>p(377)(116),clock=>clock,reset=>reset,s=>p(381)(116),cout=>p(382)(117));
FA_ff_15707:FAff port map(x=>p(375)(117),y=>p(376)(117),Cin=>p(377)(117),clock=>clock,reset=>reset,s=>p(381)(117),cout=>p(382)(118));
FA_ff_15708:FAff port map(x=>p(375)(118),y=>p(376)(118),Cin=>p(377)(118),clock=>clock,reset=>reset,s=>p(381)(118),cout=>p(382)(119));
FA_ff_15709:FAff port map(x=>p(375)(119),y=>p(376)(119),Cin=>p(377)(119),clock=>clock,reset=>reset,s=>p(381)(119),cout=>p(382)(120));
FA_ff_15710:FAff port map(x=>p(375)(120),y=>p(376)(120),Cin=>p(377)(120),clock=>clock,reset=>reset,s=>p(381)(120),cout=>p(382)(121));
FA_ff_15711:FAff port map(x=>p(375)(121),y=>p(376)(121),Cin=>p(377)(121),clock=>clock,reset=>reset,s=>p(381)(121),cout=>p(382)(122));
FA_ff_15712:FAff port map(x=>p(375)(122),y=>p(376)(122),Cin=>p(377)(122),clock=>clock,reset=>reset,s=>p(381)(122),cout=>p(382)(123));
FA_ff_15713:FAff port map(x=>p(375)(123),y=>p(376)(123),Cin=>p(377)(123),clock=>clock,reset=>reset,s=>p(381)(123),cout=>p(382)(124));
FA_ff_15714:FAff port map(x=>p(375)(124),y=>p(376)(124),Cin=>p(377)(124),clock=>clock,reset=>reset,s=>p(381)(124),cout=>p(382)(125));
FA_ff_15715:FAff port map(x=>p(375)(125),y=>p(376)(125),Cin=>p(377)(125),clock=>clock,reset=>reset,s=>p(381)(125),cout=>p(382)(126));
FA_ff_15716:FAff port map(x=>p(375)(126),y=>p(376)(126),Cin=>p(377)(126),clock=>clock,reset=>reset,s=>p(381)(126),cout=>p(382)(127));
FA_ff_15717:FAff port map(x=>p(375)(127),y=>p(376)(127),Cin=>p(377)(127),clock=>clock,reset=>reset,s=>p(381)(127),cout=>p(382)(128));
FA_ff_15718:FAff port map(x=>p(375)(128),y=>p(376)(128),Cin=>p(377)(128),clock=>clock,reset=>reset,s=>p(381)(128),cout=>p(382)(129));
FA_ff_15719:FAff port map(x=>p(375)(129),y=>p(376)(129),Cin=>p(377)(129),clock=>clock,reset=>reset,s=>p(381)(129),cout=>p(382)(130));
FA_ff_15720:FAff port map(x=>p(375)(130),y=>p(376)(130),Cin=>p(377)(130),clock=>clock,reset=>reset,s=>p(381)(130),cout=>p(382)(131));
FA_ff_15721:FAff port map(x=>p(375)(131),y=>p(376)(131),Cin=>p(377)(131),clock=>clock,reset=>reset,s=>p(381)(131),cout=>p(382)(132));
FA_ff_15722:FAff port map(x=>p(375)(132),y=>p(376)(132),Cin=>p(377)(132),clock=>clock,reset=>reset,s=>p(381)(132),cout=>p(382)(133));
p(383)(0)<=p(379)(0);
p(383)(1)<=p(379)(1);
FA_ff_15723:FAff port map(x=>p(378)(2),y=>p(379)(2),Cin=>p(380)(2),clock=>clock,reset=>reset,s=>p(383)(2),cout=>p(384)(3));
FA_ff_15724:FAff port map(x=>p(378)(3),y=>p(379)(3),Cin=>p(380)(3),clock=>clock,reset=>reset,s=>p(383)(3),cout=>p(384)(4));
FA_ff_15725:FAff port map(x=>p(378)(4),y=>p(379)(4),Cin=>p(380)(4),clock=>clock,reset=>reset,s=>p(383)(4),cout=>p(384)(5));
FA_ff_15726:FAff port map(x=>p(378)(5),y=>p(379)(5),Cin=>p(380)(5),clock=>clock,reset=>reset,s=>p(383)(5),cout=>p(384)(6));
FA_ff_15727:FAff port map(x=>p(378)(6),y=>p(379)(6),Cin=>p(380)(6),clock=>clock,reset=>reset,s=>p(383)(6),cout=>p(384)(7));
FA_ff_15728:FAff port map(x=>p(378)(7),y=>p(379)(7),Cin=>p(380)(7),clock=>clock,reset=>reset,s=>p(383)(7),cout=>p(384)(8));
FA_ff_15729:FAff port map(x=>p(378)(8),y=>p(379)(8),Cin=>p(380)(8),clock=>clock,reset=>reset,s=>p(383)(8),cout=>p(384)(9));
FA_ff_15730:FAff port map(x=>p(378)(9),y=>p(379)(9),Cin=>p(380)(9),clock=>clock,reset=>reset,s=>p(383)(9),cout=>p(384)(10));
FA_ff_15731:FAff port map(x=>p(378)(10),y=>p(379)(10),Cin=>p(380)(10),clock=>clock,reset=>reset,s=>p(383)(10),cout=>p(384)(11));
FA_ff_15732:FAff port map(x=>p(378)(11),y=>p(379)(11),Cin=>p(380)(11),clock=>clock,reset=>reset,s=>p(383)(11),cout=>p(384)(12));
FA_ff_15733:FAff port map(x=>p(378)(12),y=>p(379)(12),Cin=>p(380)(12),clock=>clock,reset=>reset,s=>p(383)(12),cout=>p(384)(13));
FA_ff_15734:FAff port map(x=>p(378)(13),y=>p(379)(13),Cin=>p(380)(13),clock=>clock,reset=>reset,s=>p(383)(13),cout=>p(384)(14));
FA_ff_15735:FAff port map(x=>p(378)(14),y=>p(379)(14),Cin=>p(380)(14),clock=>clock,reset=>reset,s=>p(383)(14),cout=>p(384)(15));
FA_ff_15736:FAff port map(x=>p(378)(15),y=>p(379)(15),Cin=>p(380)(15),clock=>clock,reset=>reset,s=>p(383)(15),cout=>p(384)(16));
FA_ff_15737:FAff port map(x=>p(378)(16),y=>p(379)(16),Cin=>p(380)(16),clock=>clock,reset=>reset,s=>p(383)(16),cout=>p(384)(17));
FA_ff_15738:FAff port map(x=>p(378)(17),y=>p(379)(17),Cin=>p(380)(17),clock=>clock,reset=>reset,s=>p(383)(17),cout=>p(384)(18));
FA_ff_15739:FAff port map(x=>p(378)(18),y=>p(379)(18),Cin=>p(380)(18),clock=>clock,reset=>reset,s=>p(383)(18),cout=>p(384)(19));
FA_ff_15740:FAff port map(x=>p(378)(19),y=>p(379)(19),Cin=>p(380)(19),clock=>clock,reset=>reset,s=>p(383)(19),cout=>p(384)(20));
FA_ff_15741:FAff port map(x=>p(378)(20),y=>p(379)(20),Cin=>p(380)(20),clock=>clock,reset=>reset,s=>p(383)(20),cout=>p(384)(21));
FA_ff_15742:FAff port map(x=>p(378)(21),y=>p(379)(21),Cin=>p(380)(21),clock=>clock,reset=>reset,s=>p(383)(21),cout=>p(384)(22));
FA_ff_15743:FAff port map(x=>p(378)(22),y=>p(379)(22),Cin=>p(380)(22),clock=>clock,reset=>reset,s=>p(383)(22),cout=>p(384)(23));
FA_ff_15744:FAff port map(x=>p(378)(23),y=>p(379)(23),Cin=>p(380)(23),clock=>clock,reset=>reset,s=>p(383)(23),cout=>p(384)(24));
FA_ff_15745:FAff port map(x=>p(378)(24),y=>p(379)(24),Cin=>p(380)(24),clock=>clock,reset=>reset,s=>p(383)(24),cout=>p(384)(25));
FA_ff_15746:FAff port map(x=>p(378)(25),y=>p(379)(25),Cin=>p(380)(25),clock=>clock,reset=>reset,s=>p(383)(25),cout=>p(384)(26));
FA_ff_15747:FAff port map(x=>p(378)(26),y=>p(379)(26),Cin=>p(380)(26),clock=>clock,reset=>reset,s=>p(383)(26),cout=>p(384)(27));
FA_ff_15748:FAff port map(x=>p(378)(27),y=>p(379)(27),Cin=>p(380)(27),clock=>clock,reset=>reset,s=>p(383)(27),cout=>p(384)(28));
FA_ff_15749:FAff port map(x=>p(378)(28),y=>p(379)(28),Cin=>p(380)(28),clock=>clock,reset=>reset,s=>p(383)(28),cout=>p(384)(29));
FA_ff_15750:FAff port map(x=>p(378)(29),y=>p(379)(29),Cin=>p(380)(29),clock=>clock,reset=>reset,s=>p(383)(29),cout=>p(384)(30));
FA_ff_15751:FAff port map(x=>p(378)(30),y=>p(379)(30),Cin=>p(380)(30),clock=>clock,reset=>reset,s=>p(383)(30),cout=>p(384)(31));
FA_ff_15752:FAff port map(x=>p(378)(31),y=>p(379)(31),Cin=>p(380)(31),clock=>clock,reset=>reset,s=>p(383)(31),cout=>p(384)(32));
FA_ff_15753:FAff port map(x=>p(378)(32),y=>p(379)(32),Cin=>p(380)(32),clock=>clock,reset=>reset,s=>p(383)(32),cout=>p(384)(33));
FA_ff_15754:FAff port map(x=>p(378)(33),y=>p(379)(33),Cin=>p(380)(33),clock=>clock,reset=>reset,s=>p(383)(33),cout=>p(384)(34));
FA_ff_15755:FAff port map(x=>p(378)(34),y=>p(379)(34),Cin=>p(380)(34),clock=>clock,reset=>reset,s=>p(383)(34),cout=>p(384)(35));
FA_ff_15756:FAff port map(x=>p(378)(35),y=>p(379)(35),Cin=>p(380)(35),clock=>clock,reset=>reset,s=>p(383)(35),cout=>p(384)(36));
FA_ff_15757:FAff port map(x=>p(378)(36),y=>p(379)(36),Cin=>p(380)(36),clock=>clock,reset=>reset,s=>p(383)(36),cout=>p(384)(37));
FA_ff_15758:FAff port map(x=>p(378)(37),y=>p(379)(37),Cin=>p(380)(37),clock=>clock,reset=>reset,s=>p(383)(37),cout=>p(384)(38));
FA_ff_15759:FAff port map(x=>p(378)(38),y=>p(379)(38),Cin=>p(380)(38),clock=>clock,reset=>reset,s=>p(383)(38),cout=>p(384)(39));
FA_ff_15760:FAff port map(x=>p(378)(39),y=>p(379)(39),Cin=>p(380)(39),clock=>clock,reset=>reset,s=>p(383)(39),cout=>p(384)(40));
FA_ff_15761:FAff port map(x=>p(378)(40),y=>p(379)(40),Cin=>p(380)(40),clock=>clock,reset=>reset,s=>p(383)(40),cout=>p(384)(41));
FA_ff_15762:FAff port map(x=>p(378)(41),y=>p(379)(41),Cin=>p(380)(41),clock=>clock,reset=>reset,s=>p(383)(41),cout=>p(384)(42));
FA_ff_15763:FAff port map(x=>p(378)(42),y=>p(379)(42),Cin=>p(380)(42),clock=>clock,reset=>reset,s=>p(383)(42),cout=>p(384)(43));
FA_ff_15764:FAff port map(x=>p(378)(43),y=>p(379)(43),Cin=>p(380)(43),clock=>clock,reset=>reset,s=>p(383)(43),cout=>p(384)(44));
FA_ff_15765:FAff port map(x=>p(378)(44),y=>p(379)(44),Cin=>p(380)(44),clock=>clock,reset=>reset,s=>p(383)(44),cout=>p(384)(45));
FA_ff_15766:FAff port map(x=>p(378)(45),y=>p(379)(45),Cin=>p(380)(45),clock=>clock,reset=>reset,s=>p(383)(45),cout=>p(384)(46));
FA_ff_15767:FAff port map(x=>p(378)(46),y=>p(379)(46),Cin=>p(380)(46),clock=>clock,reset=>reset,s=>p(383)(46),cout=>p(384)(47));
FA_ff_15768:FAff port map(x=>p(378)(47),y=>p(379)(47),Cin=>p(380)(47),clock=>clock,reset=>reset,s=>p(383)(47),cout=>p(384)(48));
FA_ff_15769:FAff port map(x=>p(378)(48),y=>p(379)(48),Cin=>p(380)(48),clock=>clock,reset=>reset,s=>p(383)(48),cout=>p(384)(49));
FA_ff_15770:FAff port map(x=>p(378)(49),y=>p(379)(49),Cin=>p(380)(49),clock=>clock,reset=>reset,s=>p(383)(49),cout=>p(384)(50));
FA_ff_15771:FAff port map(x=>p(378)(50),y=>p(379)(50),Cin=>p(380)(50),clock=>clock,reset=>reset,s=>p(383)(50),cout=>p(384)(51));
FA_ff_15772:FAff port map(x=>p(378)(51),y=>p(379)(51),Cin=>p(380)(51),clock=>clock,reset=>reset,s=>p(383)(51),cout=>p(384)(52));
FA_ff_15773:FAff port map(x=>p(378)(52),y=>p(379)(52),Cin=>p(380)(52),clock=>clock,reset=>reset,s=>p(383)(52),cout=>p(384)(53));
FA_ff_15774:FAff port map(x=>p(378)(53),y=>p(379)(53),Cin=>p(380)(53),clock=>clock,reset=>reset,s=>p(383)(53),cout=>p(384)(54));
FA_ff_15775:FAff port map(x=>p(378)(54),y=>p(379)(54),Cin=>p(380)(54),clock=>clock,reset=>reset,s=>p(383)(54),cout=>p(384)(55));
FA_ff_15776:FAff port map(x=>p(378)(55),y=>p(379)(55),Cin=>p(380)(55),clock=>clock,reset=>reset,s=>p(383)(55),cout=>p(384)(56));
FA_ff_15777:FAff port map(x=>p(378)(56),y=>p(379)(56),Cin=>p(380)(56),clock=>clock,reset=>reset,s=>p(383)(56),cout=>p(384)(57));
FA_ff_15778:FAff port map(x=>p(378)(57),y=>p(379)(57),Cin=>p(380)(57),clock=>clock,reset=>reset,s=>p(383)(57),cout=>p(384)(58));
FA_ff_15779:FAff port map(x=>p(378)(58),y=>p(379)(58),Cin=>p(380)(58),clock=>clock,reset=>reset,s=>p(383)(58),cout=>p(384)(59));
FA_ff_15780:FAff port map(x=>p(378)(59),y=>p(379)(59),Cin=>p(380)(59),clock=>clock,reset=>reset,s=>p(383)(59),cout=>p(384)(60));
FA_ff_15781:FAff port map(x=>p(378)(60),y=>p(379)(60),Cin=>p(380)(60),clock=>clock,reset=>reset,s=>p(383)(60),cout=>p(384)(61));
FA_ff_15782:FAff port map(x=>p(378)(61),y=>p(379)(61),Cin=>p(380)(61),clock=>clock,reset=>reset,s=>p(383)(61),cout=>p(384)(62));
FA_ff_15783:FAff port map(x=>p(378)(62),y=>p(379)(62),Cin=>p(380)(62),clock=>clock,reset=>reset,s=>p(383)(62),cout=>p(384)(63));
FA_ff_15784:FAff port map(x=>p(378)(63),y=>p(379)(63),Cin=>p(380)(63),clock=>clock,reset=>reset,s=>p(383)(63),cout=>p(384)(64));
FA_ff_15785:FAff port map(x=>p(378)(64),y=>p(379)(64),Cin=>p(380)(64),clock=>clock,reset=>reset,s=>p(383)(64),cout=>p(384)(65));
FA_ff_15786:FAff port map(x=>p(378)(65),y=>p(379)(65),Cin=>p(380)(65),clock=>clock,reset=>reset,s=>p(383)(65),cout=>p(384)(66));
FA_ff_15787:FAff port map(x=>p(378)(66),y=>p(379)(66),Cin=>p(380)(66),clock=>clock,reset=>reset,s=>p(383)(66),cout=>p(384)(67));
FA_ff_15788:FAff port map(x=>p(378)(67),y=>p(379)(67),Cin=>p(380)(67),clock=>clock,reset=>reset,s=>p(383)(67),cout=>p(384)(68));
FA_ff_15789:FAff port map(x=>p(378)(68),y=>p(379)(68),Cin=>p(380)(68),clock=>clock,reset=>reset,s=>p(383)(68),cout=>p(384)(69));
FA_ff_15790:FAff port map(x=>p(378)(69),y=>p(379)(69),Cin=>p(380)(69),clock=>clock,reset=>reset,s=>p(383)(69),cout=>p(384)(70));
FA_ff_15791:FAff port map(x=>p(378)(70),y=>p(379)(70),Cin=>p(380)(70),clock=>clock,reset=>reset,s=>p(383)(70),cout=>p(384)(71));
FA_ff_15792:FAff port map(x=>p(378)(71),y=>p(379)(71),Cin=>p(380)(71),clock=>clock,reset=>reset,s=>p(383)(71),cout=>p(384)(72));
FA_ff_15793:FAff port map(x=>p(378)(72),y=>p(379)(72),Cin=>p(380)(72),clock=>clock,reset=>reset,s=>p(383)(72),cout=>p(384)(73));
FA_ff_15794:FAff port map(x=>p(378)(73),y=>p(379)(73),Cin=>p(380)(73),clock=>clock,reset=>reset,s=>p(383)(73),cout=>p(384)(74));
FA_ff_15795:FAff port map(x=>p(378)(74),y=>p(379)(74),Cin=>p(380)(74),clock=>clock,reset=>reset,s=>p(383)(74),cout=>p(384)(75));
FA_ff_15796:FAff port map(x=>p(378)(75),y=>p(379)(75),Cin=>p(380)(75),clock=>clock,reset=>reset,s=>p(383)(75),cout=>p(384)(76));
FA_ff_15797:FAff port map(x=>p(378)(76),y=>p(379)(76),Cin=>p(380)(76),clock=>clock,reset=>reset,s=>p(383)(76),cout=>p(384)(77));
FA_ff_15798:FAff port map(x=>p(378)(77),y=>p(379)(77),Cin=>p(380)(77),clock=>clock,reset=>reset,s=>p(383)(77),cout=>p(384)(78));
FA_ff_15799:FAff port map(x=>p(378)(78),y=>p(379)(78),Cin=>p(380)(78),clock=>clock,reset=>reset,s=>p(383)(78),cout=>p(384)(79));
FA_ff_15800:FAff port map(x=>p(378)(79),y=>p(379)(79),Cin=>p(380)(79),clock=>clock,reset=>reset,s=>p(383)(79),cout=>p(384)(80));
FA_ff_15801:FAff port map(x=>p(378)(80),y=>p(379)(80),Cin=>p(380)(80),clock=>clock,reset=>reset,s=>p(383)(80),cout=>p(384)(81));
FA_ff_15802:FAff port map(x=>p(378)(81),y=>p(379)(81),Cin=>p(380)(81),clock=>clock,reset=>reset,s=>p(383)(81),cout=>p(384)(82));
FA_ff_15803:FAff port map(x=>p(378)(82),y=>p(379)(82),Cin=>p(380)(82),clock=>clock,reset=>reset,s=>p(383)(82),cout=>p(384)(83));
FA_ff_15804:FAff port map(x=>p(378)(83),y=>p(379)(83),Cin=>p(380)(83),clock=>clock,reset=>reset,s=>p(383)(83),cout=>p(384)(84));
FA_ff_15805:FAff port map(x=>p(378)(84),y=>p(379)(84),Cin=>p(380)(84),clock=>clock,reset=>reset,s=>p(383)(84),cout=>p(384)(85));
FA_ff_15806:FAff port map(x=>p(378)(85),y=>p(379)(85),Cin=>p(380)(85),clock=>clock,reset=>reset,s=>p(383)(85),cout=>p(384)(86));
FA_ff_15807:FAff port map(x=>p(378)(86),y=>p(379)(86),Cin=>p(380)(86),clock=>clock,reset=>reset,s=>p(383)(86),cout=>p(384)(87));
FA_ff_15808:FAff port map(x=>p(378)(87),y=>p(379)(87),Cin=>p(380)(87),clock=>clock,reset=>reset,s=>p(383)(87),cout=>p(384)(88));
FA_ff_15809:FAff port map(x=>p(378)(88),y=>p(379)(88),Cin=>p(380)(88),clock=>clock,reset=>reset,s=>p(383)(88),cout=>p(384)(89));
FA_ff_15810:FAff port map(x=>p(378)(89),y=>p(379)(89),Cin=>p(380)(89),clock=>clock,reset=>reset,s=>p(383)(89),cout=>p(384)(90));
FA_ff_15811:FAff port map(x=>p(378)(90),y=>p(379)(90),Cin=>p(380)(90),clock=>clock,reset=>reset,s=>p(383)(90),cout=>p(384)(91));
FA_ff_15812:FAff port map(x=>p(378)(91),y=>p(379)(91),Cin=>p(380)(91),clock=>clock,reset=>reset,s=>p(383)(91),cout=>p(384)(92));
FA_ff_15813:FAff port map(x=>p(378)(92),y=>p(379)(92),Cin=>p(380)(92),clock=>clock,reset=>reset,s=>p(383)(92),cout=>p(384)(93));
FA_ff_15814:FAff port map(x=>p(378)(93),y=>p(379)(93),Cin=>p(380)(93),clock=>clock,reset=>reset,s=>p(383)(93),cout=>p(384)(94));
FA_ff_15815:FAff port map(x=>p(378)(94),y=>p(379)(94),Cin=>p(380)(94),clock=>clock,reset=>reset,s=>p(383)(94),cout=>p(384)(95));
FA_ff_15816:FAff port map(x=>p(378)(95),y=>p(379)(95),Cin=>p(380)(95),clock=>clock,reset=>reset,s=>p(383)(95),cout=>p(384)(96));
FA_ff_15817:FAff port map(x=>p(378)(96),y=>p(379)(96),Cin=>p(380)(96),clock=>clock,reset=>reset,s=>p(383)(96),cout=>p(384)(97));
FA_ff_15818:FAff port map(x=>p(378)(97),y=>p(379)(97),Cin=>p(380)(97),clock=>clock,reset=>reset,s=>p(383)(97),cout=>p(384)(98));
FA_ff_15819:FAff port map(x=>p(378)(98),y=>p(379)(98),Cin=>p(380)(98),clock=>clock,reset=>reset,s=>p(383)(98),cout=>p(384)(99));
FA_ff_15820:FAff port map(x=>p(378)(99),y=>p(379)(99),Cin=>p(380)(99),clock=>clock,reset=>reset,s=>p(383)(99),cout=>p(384)(100));
FA_ff_15821:FAff port map(x=>p(378)(100),y=>p(379)(100),Cin=>p(380)(100),clock=>clock,reset=>reset,s=>p(383)(100),cout=>p(384)(101));
FA_ff_15822:FAff port map(x=>p(378)(101),y=>p(379)(101),Cin=>p(380)(101),clock=>clock,reset=>reset,s=>p(383)(101),cout=>p(384)(102));
FA_ff_15823:FAff port map(x=>p(378)(102),y=>p(379)(102),Cin=>p(380)(102),clock=>clock,reset=>reset,s=>p(383)(102),cout=>p(384)(103));
FA_ff_15824:FAff port map(x=>p(378)(103),y=>p(379)(103),Cin=>p(380)(103),clock=>clock,reset=>reset,s=>p(383)(103),cout=>p(384)(104));
FA_ff_15825:FAff port map(x=>p(378)(104),y=>p(379)(104),Cin=>p(380)(104),clock=>clock,reset=>reset,s=>p(383)(104),cout=>p(384)(105));
FA_ff_15826:FAff port map(x=>p(378)(105),y=>p(379)(105),Cin=>p(380)(105),clock=>clock,reset=>reset,s=>p(383)(105),cout=>p(384)(106));
FA_ff_15827:FAff port map(x=>p(378)(106),y=>p(379)(106),Cin=>p(380)(106),clock=>clock,reset=>reset,s=>p(383)(106),cout=>p(384)(107));
FA_ff_15828:FAff port map(x=>p(378)(107),y=>p(379)(107),Cin=>p(380)(107),clock=>clock,reset=>reset,s=>p(383)(107),cout=>p(384)(108));
FA_ff_15829:FAff port map(x=>p(378)(108),y=>p(379)(108),Cin=>p(380)(108),clock=>clock,reset=>reset,s=>p(383)(108),cout=>p(384)(109));
FA_ff_15830:FAff port map(x=>p(378)(109),y=>p(379)(109),Cin=>p(380)(109),clock=>clock,reset=>reset,s=>p(383)(109),cout=>p(384)(110));
FA_ff_15831:FAff port map(x=>p(378)(110),y=>p(379)(110),Cin=>p(380)(110),clock=>clock,reset=>reset,s=>p(383)(110),cout=>p(384)(111));
FA_ff_15832:FAff port map(x=>p(378)(111),y=>p(379)(111),Cin=>p(380)(111),clock=>clock,reset=>reset,s=>p(383)(111),cout=>p(384)(112));
FA_ff_15833:FAff port map(x=>p(378)(112),y=>p(379)(112),Cin=>p(380)(112),clock=>clock,reset=>reset,s=>p(383)(112),cout=>p(384)(113));
FA_ff_15834:FAff port map(x=>p(378)(113),y=>p(379)(113),Cin=>p(380)(113),clock=>clock,reset=>reset,s=>p(383)(113),cout=>p(384)(114));
FA_ff_15835:FAff port map(x=>p(378)(114),y=>p(379)(114),Cin=>p(380)(114),clock=>clock,reset=>reset,s=>p(383)(114),cout=>p(384)(115));
FA_ff_15836:FAff port map(x=>p(378)(115),y=>p(379)(115),Cin=>p(380)(115),clock=>clock,reset=>reset,s=>p(383)(115),cout=>p(384)(116));
FA_ff_15837:FAff port map(x=>p(378)(116),y=>p(379)(116),Cin=>p(380)(116),clock=>clock,reset=>reset,s=>p(383)(116),cout=>p(384)(117));
FA_ff_15838:FAff port map(x=>p(378)(117),y=>p(379)(117),Cin=>p(380)(117),clock=>clock,reset=>reset,s=>p(383)(117),cout=>p(384)(118));
FA_ff_15839:FAff port map(x=>p(378)(118),y=>p(379)(118),Cin=>p(380)(118),clock=>clock,reset=>reset,s=>p(383)(118),cout=>p(384)(119));
FA_ff_15840:FAff port map(x=>p(378)(119),y=>p(379)(119),Cin=>p(380)(119),clock=>clock,reset=>reset,s=>p(383)(119),cout=>p(384)(120));
FA_ff_15841:FAff port map(x=>p(378)(120),y=>p(379)(120),Cin=>p(380)(120),clock=>clock,reset=>reset,s=>p(383)(120),cout=>p(384)(121));
FA_ff_15842:FAff port map(x=>p(378)(121),y=>p(379)(121),Cin=>p(380)(121),clock=>clock,reset=>reset,s=>p(383)(121),cout=>p(384)(122));
FA_ff_15843:FAff port map(x=>p(378)(122),y=>p(379)(122),Cin=>p(380)(122),clock=>clock,reset=>reset,s=>p(383)(122),cout=>p(384)(123));
FA_ff_15844:FAff port map(x=>p(378)(123),y=>p(379)(123),Cin=>p(380)(123),clock=>clock,reset=>reset,s=>p(383)(123),cout=>p(384)(124));
FA_ff_15845:FAff port map(x=>p(378)(124),y=>p(379)(124),Cin=>p(380)(124),clock=>clock,reset=>reset,s=>p(383)(124),cout=>p(384)(125));
FA_ff_15846:FAff port map(x=>p(378)(125),y=>p(379)(125),Cin=>p(380)(125),clock=>clock,reset=>reset,s=>p(383)(125),cout=>p(384)(126));
FA_ff_15847:FAff port map(x=>p(378)(126),y=>p(379)(126),Cin=>p(380)(126),clock=>clock,reset=>reset,s=>p(383)(126),cout=>p(384)(127));
FA_ff_15848:FAff port map(x=>p(378)(127),y=>p(379)(127),Cin=>p(380)(127),clock=>clock,reset=>reset,s=>p(383)(127),cout=>p(384)(128));
FA_ff_15849:FAff port map(x=>p(378)(128),y=>p(379)(128),Cin=>p(380)(128),clock=>clock,reset=>reset,s=>p(383)(128),cout=>p(384)(129));
FA_ff_15850:FAff port map(x=>p(378)(129),y=>p(379)(129),Cin=>p(380)(129),clock=>clock,reset=>reset,s=>p(383)(129),cout=>p(384)(130));
FA_ff_15851:FAff port map(x=>p(378)(130),y=>p(379)(130),Cin=>p(380)(130),clock=>clock,reset=>reset,s=>p(383)(130),cout=>p(384)(131));
FA_ff_15852:FAff port map(x=>p(378)(131),y=>p(379)(131),Cin=>p(380)(131),clock=>clock,reset=>reset,s=>p(383)(131),cout=>p(384)(132));
HA_ff_109:HAff port map(x=>p(378)(132),y=>p(380)(132),clock=>clock,reset=>reset,s=>p(383)(132),c=>p(384)(133));
p(383)(133)<=p(378)(133);
HA_ff_110:HAff port map(x=>p(381)(0),y=>p(383)(0),clock=>clock,reset=>reset,s=>p(385)(0),c=>p(386)(1));
FA_ff_15853:FAff port map(x=>p(381)(1),y=>p(382)(1),Cin=>p(383)(1),clock=>clock,reset=>reset,s=>p(385)(1),cout=>p(386)(2));
FA_ff_15854:FAff port map(x=>p(381)(2),y=>p(382)(2),Cin=>p(383)(2),clock=>clock,reset=>reset,s=>p(385)(2),cout=>p(386)(3));
FA_ff_15855:FAff port map(x=>p(381)(3),y=>p(382)(3),Cin=>p(383)(3),clock=>clock,reset=>reset,s=>p(385)(3),cout=>p(386)(4));
FA_ff_15856:FAff port map(x=>p(381)(4),y=>p(382)(4),Cin=>p(383)(4),clock=>clock,reset=>reset,s=>p(385)(4),cout=>p(386)(5));
FA_ff_15857:FAff port map(x=>p(381)(5),y=>p(382)(5),Cin=>p(383)(5),clock=>clock,reset=>reset,s=>p(385)(5),cout=>p(386)(6));
FA_ff_15858:FAff port map(x=>p(381)(6),y=>p(382)(6),Cin=>p(383)(6),clock=>clock,reset=>reset,s=>p(385)(6),cout=>p(386)(7));
FA_ff_15859:FAff port map(x=>p(381)(7),y=>p(382)(7),Cin=>p(383)(7),clock=>clock,reset=>reset,s=>p(385)(7),cout=>p(386)(8));
FA_ff_15860:FAff port map(x=>p(381)(8),y=>p(382)(8),Cin=>p(383)(8),clock=>clock,reset=>reset,s=>p(385)(8),cout=>p(386)(9));
FA_ff_15861:FAff port map(x=>p(381)(9),y=>p(382)(9),Cin=>p(383)(9),clock=>clock,reset=>reset,s=>p(385)(9),cout=>p(386)(10));
FA_ff_15862:FAff port map(x=>p(381)(10),y=>p(382)(10),Cin=>p(383)(10),clock=>clock,reset=>reset,s=>p(385)(10),cout=>p(386)(11));
FA_ff_15863:FAff port map(x=>p(381)(11),y=>p(382)(11),Cin=>p(383)(11),clock=>clock,reset=>reset,s=>p(385)(11),cout=>p(386)(12));
FA_ff_15864:FAff port map(x=>p(381)(12),y=>p(382)(12),Cin=>p(383)(12),clock=>clock,reset=>reset,s=>p(385)(12),cout=>p(386)(13));
FA_ff_15865:FAff port map(x=>p(381)(13),y=>p(382)(13),Cin=>p(383)(13),clock=>clock,reset=>reset,s=>p(385)(13),cout=>p(386)(14));
FA_ff_15866:FAff port map(x=>p(381)(14),y=>p(382)(14),Cin=>p(383)(14),clock=>clock,reset=>reset,s=>p(385)(14),cout=>p(386)(15));
FA_ff_15867:FAff port map(x=>p(381)(15),y=>p(382)(15),Cin=>p(383)(15),clock=>clock,reset=>reset,s=>p(385)(15),cout=>p(386)(16));
FA_ff_15868:FAff port map(x=>p(381)(16),y=>p(382)(16),Cin=>p(383)(16),clock=>clock,reset=>reset,s=>p(385)(16),cout=>p(386)(17));
FA_ff_15869:FAff port map(x=>p(381)(17),y=>p(382)(17),Cin=>p(383)(17),clock=>clock,reset=>reset,s=>p(385)(17),cout=>p(386)(18));
FA_ff_15870:FAff port map(x=>p(381)(18),y=>p(382)(18),Cin=>p(383)(18),clock=>clock,reset=>reset,s=>p(385)(18),cout=>p(386)(19));
FA_ff_15871:FAff port map(x=>p(381)(19),y=>p(382)(19),Cin=>p(383)(19),clock=>clock,reset=>reset,s=>p(385)(19),cout=>p(386)(20));
FA_ff_15872:FAff port map(x=>p(381)(20),y=>p(382)(20),Cin=>p(383)(20),clock=>clock,reset=>reset,s=>p(385)(20),cout=>p(386)(21));
FA_ff_15873:FAff port map(x=>p(381)(21),y=>p(382)(21),Cin=>p(383)(21),clock=>clock,reset=>reset,s=>p(385)(21),cout=>p(386)(22));
FA_ff_15874:FAff port map(x=>p(381)(22),y=>p(382)(22),Cin=>p(383)(22),clock=>clock,reset=>reset,s=>p(385)(22),cout=>p(386)(23));
FA_ff_15875:FAff port map(x=>p(381)(23),y=>p(382)(23),Cin=>p(383)(23),clock=>clock,reset=>reset,s=>p(385)(23),cout=>p(386)(24));
FA_ff_15876:FAff port map(x=>p(381)(24),y=>p(382)(24),Cin=>p(383)(24),clock=>clock,reset=>reset,s=>p(385)(24),cout=>p(386)(25));
FA_ff_15877:FAff port map(x=>p(381)(25),y=>p(382)(25),Cin=>p(383)(25),clock=>clock,reset=>reset,s=>p(385)(25),cout=>p(386)(26));
FA_ff_15878:FAff port map(x=>p(381)(26),y=>p(382)(26),Cin=>p(383)(26),clock=>clock,reset=>reset,s=>p(385)(26),cout=>p(386)(27));
FA_ff_15879:FAff port map(x=>p(381)(27),y=>p(382)(27),Cin=>p(383)(27),clock=>clock,reset=>reset,s=>p(385)(27),cout=>p(386)(28));
FA_ff_15880:FAff port map(x=>p(381)(28),y=>p(382)(28),Cin=>p(383)(28),clock=>clock,reset=>reset,s=>p(385)(28),cout=>p(386)(29));
FA_ff_15881:FAff port map(x=>p(381)(29),y=>p(382)(29),Cin=>p(383)(29),clock=>clock,reset=>reset,s=>p(385)(29),cout=>p(386)(30));
FA_ff_15882:FAff port map(x=>p(381)(30),y=>p(382)(30),Cin=>p(383)(30),clock=>clock,reset=>reset,s=>p(385)(30),cout=>p(386)(31));
FA_ff_15883:FAff port map(x=>p(381)(31),y=>p(382)(31),Cin=>p(383)(31),clock=>clock,reset=>reset,s=>p(385)(31),cout=>p(386)(32));
FA_ff_15884:FAff port map(x=>p(381)(32),y=>p(382)(32),Cin=>p(383)(32),clock=>clock,reset=>reset,s=>p(385)(32),cout=>p(386)(33));
FA_ff_15885:FAff port map(x=>p(381)(33),y=>p(382)(33),Cin=>p(383)(33),clock=>clock,reset=>reset,s=>p(385)(33),cout=>p(386)(34));
FA_ff_15886:FAff port map(x=>p(381)(34),y=>p(382)(34),Cin=>p(383)(34),clock=>clock,reset=>reset,s=>p(385)(34),cout=>p(386)(35));
FA_ff_15887:FAff port map(x=>p(381)(35),y=>p(382)(35),Cin=>p(383)(35),clock=>clock,reset=>reset,s=>p(385)(35),cout=>p(386)(36));
FA_ff_15888:FAff port map(x=>p(381)(36),y=>p(382)(36),Cin=>p(383)(36),clock=>clock,reset=>reset,s=>p(385)(36),cout=>p(386)(37));
FA_ff_15889:FAff port map(x=>p(381)(37),y=>p(382)(37),Cin=>p(383)(37),clock=>clock,reset=>reset,s=>p(385)(37),cout=>p(386)(38));
FA_ff_15890:FAff port map(x=>p(381)(38),y=>p(382)(38),Cin=>p(383)(38),clock=>clock,reset=>reset,s=>p(385)(38),cout=>p(386)(39));
FA_ff_15891:FAff port map(x=>p(381)(39),y=>p(382)(39),Cin=>p(383)(39),clock=>clock,reset=>reset,s=>p(385)(39),cout=>p(386)(40));
FA_ff_15892:FAff port map(x=>p(381)(40),y=>p(382)(40),Cin=>p(383)(40),clock=>clock,reset=>reset,s=>p(385)(40),cout=>p(386)(41));
FA_ff_15893:FAff port map(x=>p(381)(41),y=>p(382)(41),Cin=>p(383)(41),clock=>clock,reset=>reset,s=>p(385)(41),cout=>p(386)(42));
FA_ff_15894:FAff port map(x=>p(381)(42),y=>p(382)(42),Cin=>p(383)(42),clock=>clock,reset=>reset,s=>p(385)(42),cout=>p(386)(43));
FA_ff_15895:FAff port map(x=>p(381)(43),y=>p(382)(43),Cin=>p(383)(43),clock=>clock,reset=>reset,s=>p(385)(43),cout=>p(386)(44));
FA_ff_15896:FAff port map(x=>p(381)(44),y=>p(382)(44),Cin=>p(383)(44),clock=>clock,reset=>reset,s=>p(385)(44),cout=>p(386)(45));
FA_ff_15897:FAff port map(x=>p(381)(45),y=>p(382)(45),Cin=>p(383)(45),clock=>clock,reset=>reset,s=>p(385)(45),cout=>p(386)(46));
FA_ff_15898:FAff port map(x=>p(381)(46),y=>p(382)(46),Cin=>p(383)(46),clock=>clock,reset=>reset,s=>p(385)(46),cout=>p(386)(47));
FA_ff_15899:FAff port map(x=>p(381)(47),y=>p(382)(47),Cin=>p(383)(47),clock=>clock,reset=>reset,s=>p(385)(47),cout=>p(386)(48));
FA_ff_15900:FAff port map(x=>p(381)(48),y=>p(382)(48),Cin=>p(383)(48),clock=>clock,reset=>reset,s=>p(385)(48),cout=>p(386)(49));
FA_ff_15901:FAff port map(x=>p(381)(49),y=>p(382)(49),Cin=>p(383)(49),clock=>clock,reset=>reset,s=>p(385)(49),cout=>p(386)(50));
FA_ff_15902:FAff port map(x=>p(381)(50),y=>p(382)(50),Cin=>p(383)(50),clock=>clock,reset=>reset,s=>p(385)(50),cout=>p(386)(51));
FA_ff_15903:FAff port map(x=>p(381)(51),y=>p(382)(51),Cin=>p(383)(51),clock=>clock,reset=>reset,s=>p(385)(51),cout=>p(386)(52));
FA_ff_15904:FAff port map(x=>p(381)(52),y=>p(382)(52),Cin=>p(383)(52),clock=>clock,reset=>reset,s=>p(385)(52),cout=>p(386)(53));
FA_ff_15905:FAff port map(x=>p(381)(53),y=>p(382)(53),Cin=>p(383)(53),clock=>clock,reset=>reset,s=>p(385)(53),cout=>p(386)(54));
FA_ff_15906:FAff port map(x=>p(381)(54),y=>p(382)(54),Cin=>p(383)(54),clock=>clock,reset=>reset,s=>p(385)(54),cout=>p(386)(55));
FA_ff_15907:FAff port map(x=>p(381)(55),y=>p(382)(55),Cin=>p(383)(55),clock=>clock,reset=>reset,s=>p(385)(55),cout=>p(386)(56));
FA_ff_15908:FAff port map(x=>p(381)(56),y=>p(382)(56),Cin=>p(383)(56),clock=>clock,reset=>reset,s=>p(385)(56),cout=>p(386)(57));
FA_ff_15909:FAff port map(x=>p(381)(57),y=>p(382)(57),Cin=>p(383)(57),clock=>clock,reset=>reset,s=>p(385)(57),cout=>p(386)(58));
FA_ff_15910:FAff port map(x=>p(381)(58),y=>p(382)(58),Cin=>p(383)(58),clock=>clock,reset=>reset,s=>p(385)(58),cout=>p(386)(59));
FA_ff_15911:FAff port map(x=>p(381)(59),y=>p(382)(59),Cin=>p(383)(59),clock=>clock,reset=>reset,s=>p(385)(59),cout=>p(386)(60));
FA_ff_15912:FAff port map(x=>p(381)(60),y=>p(382)(60),Cin=>p(383)(60),clock=>clock,reset=>reset,s=>p(385)(60),cout=>p(386)(61));
FA_ff_15913:FAff port map(x=>p(381)(61),y=>p(382)(61),Cin=>p(383)(61),clock=>clock,reset=>reset,s=>p(385)(61),cout=>p(386)(62));
FA_ff_15914:FAff port map(x=>p(381)(62),y=>p(382)(62),Cin=>p(383)(62),clock=>clock,reset=>reset,s=>p(385)(62),cout=>p(386)(63));
FA_ff_15915:FAff port map(x=>p(381)(63),y=>p(382)(63),Cin=>p(383)(63),clock=>clock,reset=>reset,s=>p(385)(63),cout=>p(386)(64));
FA_ff_15916:FAff port map(x=>p(381)(64),y=>p(382)(64),Cin=>p(383)(64),clock=>clock,reset=>reset,s=>p(385)(64),cout=>p(386)(65));
FA_ff_15917:FAff port map(x=>p(381)(65),y=>p(382)(65),Cin=>p(383)(65),clock=>clock,reset=>reset,s=>p(385)(65),cout=>p(386)(66));
FA_ff_15918:FAff port map(x=>p(381)(66),y=>p(382)(66),Cin=>p(383)(66),clock=>clock,reset=>reset,s=>p(385)(66),cout=>p(386)(67));
FA_ff_15919:FAff port map(x=>p(381)(67),y=>p(382)(67),Cin=>p(383)(67),clock=>clock,reset=>reset,s=>p(385)(67),cout=>p(386)(68));
FA_ff_15920:FAff port map(x=>p(381)(68),y=>p(382)(68),Cin=>p(383)(68),clock=>clock,reset=>reset,s=>p(385)(68),cout=>p(386)(69));
FA_ff_15921:FAff port map(x=>p(381)(69),y=>p(382)(69),Cin=>p(383)(69),clock=>clock,reset=>reset,s=>p(385)(69),cout=>p(386)(70));
FA_ff_15922:FAff port map(x=>p(381)(70),y=>p(382)(70),Cin=>p(383)(70),clock=>clock,reset=>reset,s=>p(385)(70),cout=>p(386)(71));
FA_ff_15923:FAff port map(x=>p(381)(71),y=>p(382)(71),Cin=>p(383)(71),clock=>clock,reset=>reset,s=>p(385)(71),cout=>p(386)(72));
FA_ff_15924:FAff port map(x=>p(381)(72),y=>p(382)(72),Cin=>p(383)(72),clock=>clock,reset=>reset,s=>p(385)(72),cout=>p(386)(73));
FA_ff_15925:FAff port map(x=>p(381)(73),y=>p(382)(73),Cin=>p(383)(73),clock=>clock,reset=>reset,s=>p(385)(73),cout=>p(386)(74));
FA_ff_15926:FAff port map(x=>p(381)(74),y=>p(382)(74),Cin=>p(383)(74),clock=>clock,reset=>reset,s=>p(385)(74),cout=>p(386)(75));
FA_ff_15927:FAff port map(x=>p(381)(75),y=>p(382)(75),Cin=>p(383)(75),clock=>clock,reset=>reset,s=>p(385)(75),cout=>p(386)(76));
FA_ff_15928:FAff port map(x=>p(381)(76),y=>p(382)(76),Cin=>p(383)(76),clock=>clock,reset=>reset,s=>p(385)(76),cout=>p(386)(77));
FA_ff_15929:FAff port map(x=>p(381)(77),y=>p(382)(77),Cin=>p(383)(77),clock=>clock,reset=>reset,s=>p(385)(77),cout=>p(386)(78));
FA_ff_15930:FAff port map(x=>p(381)(78),y=>p(382)(78),Cin=>p(383)(78),clock=>clock,reset=>reset,s=>p(385)(78),cout=>p(386)(79));
FA_ff_15931:FAff port map(x=>p(381)(79),y=>p(382)(79),Cin=>p(383)(79),clock=>clock,reset=>reset,s=>p(385)(79),cout=>p(386)(80));
FA_ff_15932:FAff port map(x=>p(381)(80),y=>p(382)(80),Cin=>p(383)(80),clock=>clock,reset=>reset,s=>p(385)(80),cout=>p(386)(81));
FA_ff_15933:FAff port map(x=>p(381)(81),y=>p(382)(81),Cin=>p(383)(81),clock=>clock,reset=>reset,s=>p(385)(81),cout=>p(386)(82));
FA_ff_15934:FAff port map(x=>p(381)(82),y=>p(382)(82),Cin=>p(383)(82),clock=>clock,reset=>reset,s=>p(385)(82),cout=>p(386)(83));
FA_ff_15935:FAff port map(x=>p(381)(83),y=>p(382)(83),Cin=>p(383)(83),clock=>clock,reset=>reset,s=>p(385)(83),cout=>p(386)(84));
FA_ff_15936:FAff port map(x=>p(381)(84),y=>p(382)(84),Cin=>p(383)(84),clock=>clock,reset=>reset,s=>p(385)(84),cout=>p(386)(85));
FA_ff_15937:FAff port map(x=>p(381)(85),y=>p(382)(85),Cin=>p(383)(85),clock=>clock,reset=>reset,s=>p(385)(85),cout=>p(386)(86));
FA_ff_15938:FAff port map(x=>p(381)(86),y=>p(382)(86),Cin=>p(383)(86),clock=>clock,reset=>reset,s=>p(385)(86),cout=>p(386)(87));
FA_ff_15939:FAff port map(x=>p(381)(87),y=>p(382)(87),Cin=>p(383)(87),clock=>clock,reset=>reset,s=>p(385)(87),cout=>p(386)(88));
FA_ff_15940:FAff port map(x=>p(381)(88),y=>p(382)(88),Cin=>p(383)(88),clock=>clock,reset=>reset,s=>p(385)(88),cout=>p(386)(89));
FA_ff_15941:FAff port map(x=>p(381)(89),y=>p(382)(89),Cin=>p(383)(89),clock=>clock,reset=>reset,s=>p(385)(89),cout=>p(386)(90));
FA_ff_15942:FAff port map(x=>p(381)(90),y=>p(382)(90),Cin=>p(383)(90),clock=>clock,reset=>reset,s=>p(385)(90),cout=>p(386)(91));
FA_ff_15943:FAff port map(x=>p(381)(91),y=>p(382)(91),Cin=>p(383)(91),clock=>clock,reset=>reset,s=>p(385)(91),cout=>p(386)(92));
FA_ff_15944:FAff port map(x=>p(381)(92),y=>p(382)(92),Cin=>p(383)(92),clock=>clock,reset=>reset,s=>p(385)(92),cout=>p(386)(93));
FA_ff_15945:FAff port map(x=>p(381)(93),y=>p(382)(93),Cin=>p(383)(93),clock=>clock,reset=>reset,s=>p(385)(93),cout=>p(386)(94));
FA_ff_15946:FAff port map(x=>p(381)(94),y=>p(382)(94),Cin=>p(383)(94),clock=>clock,reset=>reset,s=>p(385)(94),cout=>p(386)(95));
FA_ff_15947:FAff port map(x=>p(381)(95),y=>p(382)(95),Cin=>p(383)(95),clock=>clock,reset=>reset,s=>p(385)(95),cout=>p(386)(96));
FA_ff_15948:FAff port map(x=>p(381)(96),y=>p(382)(96),Cin=>p(383)(96),clock=>clock,reset=>reset,s=>p(385)(96),cout=>p(386)(97));
FA_ff_15949:FAff port map(x=>p(381)(97),y=>p(382)(97),Cin=>p(383)(97),clock=>clock,reset=>reset,s=>p(385)(97),cout=>p(386)(98));
FA_ff_15950:FAff port map(x=>p(381)(98),y=>p(382)(98),Cin=>p(383)(98),clock=>clock,reset=>reset,s=>p(385)(98),cout=>p(386)(99));
FA_ff_15951:FAff port map(x=>p(381)(99),y=>p(382)(99),Cin=>p(383)(99),clock=>clock,reset=>reset,s=>p(385)(99),cout=>p(386)(100));
FA_ff_15952:FAff port map(x=>p(381)(100),y=>p(382)(100),Cin=>p(383)(100),clock=>clock,reset=>reset,s=>p(385)(100),cout=>p(386)(101));
FA_ff_15953:FAff port map(x=>p(381)(101),y=>p(382)(101),Cin=>p(383)(101),clock=>clock,reset=>reset,s=>p(385)(101),cout=>p(386)(102));
FA_ff_15954:FAff port map(x=>p(381)(102),y=>p(382)(102),Cin=>p(383)(102),clock=>clock,reset=>reset,s=>p(385)(102),cout=>p(386)(103));
FA_ff_15955:FAff port map(x=>p(381)(103),y=>p(382)(103),Cin=>p(383)(103),clock=>clock,reset=>reset,s=>p(385)(103),cout=>p(386)(104));
FA_ff_15956:FAff port map(x=>p(381)(104),y=>p(382)(104),Cin=>p(383)(104),clock=>clock,reset=>reset,s=>p(385)(104),cout=>p(386)(105));
FA_ff_15957:FAff port map(x=>p(381)(105),y=>p(382)(105),Cin=>p(383)(105),clock=>clock,reset=>reset,s=>p(385)(105),cout=>p(386)(106));
FA_ff_15958:FAff port map(x=>p(381)(106),y=>p(382)(106),Cin=>p(383)(106),clock=>clock,reset=>reset,s=>p(385)(106),cout=>p(386)(107));
FA_ff_15959:FAff port map(x=>p(381)(107),y=>p(382)(107),Cin=>p(383)(107),clock=>clock,reset=>reset,s=>p(385)(107),cout=>p(386)(108));
FA_ff_15960:FAff port map(x=>p(381)(108),y=>p(382)(108),Cin=>p(383)(108),clock=>clock,reset=>reset,s=>p(385)(108),cout=>p(386)(109));
FA_ff_15961:FAff port map(x=>p(381)(109),y=>p(382)(109),Cin=>p(383)(109),clock=>clock,reset=>reset,s=>p(385)(109),cout=>p(386)(110));
FA_ff_15962:FAff port map(x=>p(381)(110),y=>p(382)(110),Cin=>p(383)(110),clock=>clock,reset=>reset,s=>p(385)(110),cout=>p(386)(111));
FA_ff_15963:FAff port map(x=>p(381)(111),y=>p(382)(111),Cin=>p(383)(111),clock=>clock,reset=>reset,s=>p(385)(111),cout=>p(386)(112));
FA_ff_15964:FAff port map(x=>p(381)(112),y=>p(382)(112),Cin=>p(383)(112),clock=>clock,reset=>reset,s=>p(385)(112),cout=>p(386)(113));
FA_ff_15965:FAff port map(x=>p(381)(113),y=>p(382)(113),Cin=>p(383)(113),clock=>clock,reset=>reset,s=>p(385)(113),cout=>p(386)(114));
FA_ff_15966:FAff port map(x=>p(381)(114),y=>p(382)(114),Cin=>p(383)(114),clock=>clock,reset=>reset,s=>p(385)(114),cout=>p(386)(115));
FA_ff_15967:FAff port map(x=>p(381)(115),y=>p(382)(115),Cin=>p(383)(115),clock=>clock,reset=>reset,s=>p(385)(115),cout=>p(386)(116));
FA_ff_15968:FAff port map(x=>p(381)(116),y=>p(382)(116),Cin=>p(383)(116),clock=>clock,reset=>reset,s=>p(385)(116),cout=>p(386)(117));
FA_ff_15969:FAff port map(x=>p(381)(117),y=>p(382)(117),Cin=>p(383)(117),clock=>clock,reset=>reset,s=>p(385)(117),cout=>p(386)(118));
FA_ff_15970:FAff port map(x=>p(381)(118),y=>p(382)(118),Cin=>p(383)(118),clock=>clock,reset=>reset,s=>p(385)(118),cout=>p(386)(119));
FA_ff_15971:FAff port map(x=>p(381)(119),y=>p(382)(119),Cin=>p(383)(119),clock=>clock,reset=>reset,s=>p(385)(119),cout=>p(386)(120));
FA_ff_15972:FAff port map(x=>p(381)(120),y=>p(382)(120),Cin=>p(383)(120),clock=>clock,reset=>reset,s=>p(385)(120),cout=>p(386)(121));
FA_ff_15973:FAff port map(x=>p(381)(121),y=>p(382)(121),Cin=>p(383)(121),clock=>clock,reset=>reset,s=>p(385)(121),cout=>p(386)(122));
FA_ff_15974:FAff port map(x=>p(381)(122),y=>p(382)(122),Cin=>p(383)(122),clock=>clock,reset=>reset,s=>p(385)(122),cout=>p(386)(123));
FA_ff_15975:FAff port map(x=>p(381)(123),y=>p(382)(123),Cin=>p(383)(123),clock=>clock,reset=>reset,s=>p(385)(123),cout=>p(386)(124));
FA_ff_15976:FAff port map(x=>p(381)(124),y=>p(382)(124),Cin=>p(383)(124),clock=>clock,reset=>reset,s=>p(385)(124),cout=>p(386)(125));
FA_ff_15977:FAff port map(x=>p(381)(125),y=>p(382)(125),Cin=>p(383)(125),clock=>clock,reset=>reset,s=>p(385)(125),cout=>p(386)(126));
FA_ff_15978:FAff port map(x=>p(381)(126),y=>p(382)(126),Cin=>p(383)(126),clock=>clock,reset=>reset,s=>p(385)(126),cout=>p(386)(127));
FA_ff_15979:FAff port map(x=>p(381)(127),y=>p(382)(127),Cin=>p(383)(127),clock=>clock,reset=>reset,s=>p(385)(127),cout=>p(386)(128));
FA_ff_15980:FAff port map(x=>p(381)(128),y=>p(382)(128),Cin=>p(383)(128),clock=>clock,reset=>reset,s=>p(385)(128),cout=>p(386)(129));
FA_ff_15981:FAff port map(x=>p(381)(129),y=>p(382)(129),Cin=>p(383)(129),clock=>clock,reset=>reset,s=>p(385)(129),cout=>p(386)(130));
FA_ff_15982:FAff port map(x=>p(381)(130),y=>p(382)(130),Cin=>p(383)(130),clock=>clock,reset=>reset,s=>p(385)(130),cout=>p(386)(131));
FA_ff_15983:FAff port map(x=>p(381)(131),y=>p(382)(131),Cin=>p(383)(131),clock=>clock,reset=>reset,s=>p(385)(131),cout=>p(386)(132));
FA_ff_15984:FAff port map(x=>p(381)(132),y=>p(382)(132),Cin=>p(383)(132),clock=>clock,reset=>reset,s=>p(385)(132),cout=>p(386)(133));
HA_ff_111:HAff port map(x=>p(382)(133),y=>p(383)(133),clock=>clock,reset=>reset,s=>p(385)(133),c=>p(386)(134));
p(387)(0)<=p(384)(0);
p(387)(1)<=p(384)(1);
p(387)(2)<=p(384)(2);
p(387)(3)<=p(384)(3);
p(387)(4)<=p(384)(4);
p(387)(5)<=p(384)(5);
p(387)(6)<=p(384)(6);
p(387)(7)<=p(384)(7);
p(387)(8)<=p(384)(8);
p(387)(9)<=p(384)(9);
p(387)(10)<=p(384)(10);
p(387)(11)<=p(384)(11);
p(387)(12)<=p(384)(12);
p(387)(13)<=p(384)(13);
p(387)(14)<=p(384)(14);
p(387)(15)<=p(384)(15);
p(387)(16)<=p(384)(16);
p(387)(17)<=p(384)(17);
p(387)(18)<=p(384)(18);
p(387)(19)<=p(384)(19);
p(387)(20)<=p(384)(20);
p(387)(21)<=p(384)(21);
p(387)(22)<=p(384)(22);
p(387)(23)<=p(384)(23);
p(387)(24)<=p(384)(24);
p(387)(25)<=p(384)(25);
p(387)(26)<=p(384)(26);
p(387)(27)<=p(384)(27);
p(387)(28)<=p(384)(28);
p(387)(29)<=p(384)(29);
p(387)(30)<=p(384)(30);
p(387)(31)<=p(384)(31);
p(387)(32)<=p(384)(32);
p(387)(33)<=p(384)(33);
p(387)(34)<=p(384)(34);
p(387)(35)<=p(384)(35);
p(387)(36)<=p(384)(36);
p(387)(37)<=p(384)(37);
p(387)(38)<=p(384)(38);
p(387)(39)<=p(384)(39);
p(387)(40)<=p(384)(40);
p(387)(41)<=p(384)(41);
p(387)(42)<=p(384)(42);
p(387)(43)<=p(384)(43);
p(387)(44)<=p(384)(44);
p(387)(45)<=p(384)(45);
p(387)(46)<=p(384)(46);
p(387)(47)<=p(384)(47);
p(387)(48)<=p(384)(48);
p(387)(49)<=p(384)(49);
p(387)(50)<=p(384)(50);
p(387)(51)<=p(384)(51);
p(387)(52)<=p(384)(52);
p(387)(53)<=p(384)(53);
p(387)(54)<=p(384)(54);
p(387)(55)<=p(384)(55);
p(387)(56)<=p(384)(56);
p(387)(57)<=p(384)(57);
p(387)(58)<=p(384)(58);
p(387)(59)<=p(384)(59);
p(387)(60)<=p(384)(60);
p(387)(61)<=p(384)(61);
p(387)(62)<=p(384)(62);
p(387)(63)<=p(384)(63);
p(387)(64)<=p(384)(64);
p(387)(65)<=p(384)(65);
p(387)(66)<=p(384)(66);
p(387)(67)<=p(384)(67);
p(387)(68)<=p(384)(68);
p(387)(69)<=p(384)(69);
p(387)(70)<=p(384)(70);
p(387)(71)<=p(384)(71);
p(387)(72)<=p(384)(72);
p(387)(73)<=p(384)(73);
p(387)(74)<=p(384)(74);
p(387)(75)<=p(384)(75);
p(387)(76)<=p(384)(76);
p(387)(77)<=p(384)(77);
p(387)(78)<=p(384)(78);
p(387)(79)<=p(384)(79);
p(387)(80)<=p(384)(80);
p(387)(81)<=p(384)(81);
p(387)(82)<=p(384)(82);
p(387)(83)<=p(384)(83);
p(387)(84)<=p(384)(84);
p(387)(85)<=p(384)(85);
p(387)(86)<=p(384)(86);
p(387)(87)<=p(384)(87);
p(387)(88)<=p(384)(88);
p(387)(89)<=p(384)(89);
p(387)(90)<=p(384)(90);
p(387)(91)<=p(384)(91);
p(387)(92)<=p(384)(92);
p(387)(93)<=p(384)(93);
p(387)(94)<=p(384)(94);
p(387)(95)<=p(384)(95);
p(387)(96)<=p(384)(96);
p(387)(97)<=p(384)(97);
p(387)(98)<=p(384)(98);
p(387)(99)<=p(384)(99);
p(387)(100)<=p(384)(100);
p(387)(101)<=p(384)(101);
p(387)(102)<=p(384)(102);
p(387)(103)<=p(384)(103);
p(387)(104)<=p(384)(104);
p(387)(105)<=p(384)(105);
p(387)(106)<=p(384)(106);
p(387)(107)<=p(384)(107);
p(387)(108)<=p(384)(108);
p(387)(109)<=p(384)(109);
p(387)(110)<=p(384)(110);
p(387)(111)<=p(384)(111);
p(387)(112)<=p(384)(112);
p(387)(113)<=p(384)(113);
p(387)(114)<=p(384)(114);
p(387)(115)<=p(384)(115);
p(387)(116)<=p(384)(116);
p(387)(117)<=p(384)(117);
p(387)(118)<=p(384)(118);
p(387)(119)<=p(384)(119);
p(387)(120)<=p(384)(120);
p(387)(121)<=p(384)(121);
p(387)(122)<=p(384)(122);
p(387)(123)<=p(384)(123);
p(387)(124)<=p(384)(124);
p(387)(125)<=p(384)(125);
p(387)(126)<=p(384)(126);
p(387)(127)<=p(384)(127);
p(387)(128)<=p(384)(128);
p(387)(129)<=p(384)(129);
p(387)(130)<=p(384)(130);
p(387)(131)<=p(384)(131);
p(387)(132)<=p(384)(132);
p(387)(133)<=p(384)(133);
p(387)(134)<=p(384)(134);
p(388)(0)<=p(385)(0);
HA_ff_112:HAff port map(x=>p(385)(1),y=>p(386)(1),clock=>clock,reset=>reset,s=>p(388)(1),c=>p(389)(2));
HA_ff_113:HAff port map(x=>p(385)(2),y=>p(386)(2),clock=>clock,reset=>reset,s=>p(388)(2),c=>p(389)(3));
FA_ff_15985:FAff port map(x=>p(385)(3),y=>p(386)(3),Cin=>p(387)(3),clock=>clock,reset=>reset,s=>p(388)(3),cout=>p(389)(4));
FA_ff_15986:FAff port map(x=>p(385)(4),y=>p(386)(4),Cin=>p(387)(4),clock=>clock,reset=>reset,s=>p(388)(4),cout=>p(389)(5));
FA_ff_15987:FAff port map(x=>p(385)(5),y=>p(386)(5),Cin=>p(387)(5),clock=>clock,reset=>reset,s=>p(388)(5),cout=>p(389)(6));
FA_ff_15988:FAff port map(x=>p(385)(6),y=>p(386)(6),Cin=>p(387)(6),clock=>clock,reset=>reset,s=>p(388)(6),cout=>p(389)(7));
FA_ff_15989:FAff port map(x=>p(385)(7),y=>p(386)(7),Cin=>p(387)(7),clock=>clock,reset=>reset,s=>p(388)(7),cout=>p(389)(8));
FA_ff_15990:FAff port map(x=>p(385)(8),y=>p(386)(8),Cin=>p(387)(8),clock=>clock,reset=>reset,s=>p(388)(8),cout=>p(389)(9));
FA_ff_15991:FAff port map(x=>p(385)(9),y=>p(386)(9),Cin=>p(387)(9),clock=>clock,reset=>reset,s=>p(388)(9),cout=>p(389)(10));
FA_ff_15992:FAff port map(x=>p(385)(10),y=>p(386)(10),Cin=>p(387)(10),clock=>clock,reset=>reset,s=>p(388)(10),cout=>p(389)(11));
FA_ff_15993:FAff port map(x=>p(385)(11),y=>p(386)(11),Cin=>p(387)(11),clock=>clock,reset=>reset,s=>p(388)(11),cout=>p(389)(12));
FA_ff_15994:FAff port map(x=>p(385)(12),y=>p(386)(12),Cin=>p(387)(12),clock=>clock,reset=>reset,s=>p(388)(12),cout=>p(389)(13));
FA_ff_15995:FAff port map(x=>p(385)(13),y=>p(386)(13),Cin=>p(387)(13),clock=>clock,reset=>reset,s=>p(388)(13),cout=>p(389)(14));
FA_ff_15996:FAff port map(x=>p(385)(14),y=>p(386)(14),Cin=>p(387)(14),clock=>clock,reset=>reset,s=>p(388)(14),cout=>p(389)(15));
FA_ff_15997:FAff port map(x=>p(385)(15),y=>p(386)(15),Cin=>p(387)(15),clock=>clock,reset=>reset,s=>p(388)(15),cout=>p(389)(16));
FA_ff_15998:FAff port map(x=>p(385)(16),y=>p(386)(16),Cin=>p(387)(16),clock=>clock,reset=>reset,s=>p(388)(16),cout=>p(389)(17));
FA_ff_15999:FAff port map(x=>p(385)(17),y=>p(386)(17),Cin=>p(387)(17),clock=>clock,reset=>reset,s=>p(388)(17),cout=>p(389)(18));
FA_ff_16000:FAff port map(x=>p(385)(18),y=>p(386)(18),Cin=>p(387)(18),clock=>clock,reset=>reset,s=>p(388)(18),cout=>p(389)(19));
FA_ff_16001:FAff port map(x=>p(385)(19),y=>p(386)(19),Cin=>p(387)(19),clock=>clock,reset=>reset,s=>p(388)(19),cout=>p(389)(20));
FA_ff_16002:FAff port map(x=>p(385)(20),y=>p(386)(20),Cin=>p(387)(20),clock=>clock,reset=>reset,s=>p(388)(20),cout=>p(389)(21));
FA_ff_16003:FAff port map(x=>p(385)(21),y=>p(386)(21),Cin=>p(387)(21),clock=>clock,reset=>reset,s=>p(388)(21),cout=>p(389)(22));
FA_ff_16004:FAff port map(x=>p(385)(22),y=>p(386)(22),Cin=>p(387)(22),clock=>clock,reset=>reset,s=>p(388)(22),cout=>p(389)(23));
FA_ff_16005:FAff port map(x=>p(385)(23),y=>p(386)(23),Cin=>p(387)(23),clock=>clock,reset=>reset,s=>p(388)(23),cout=>p(389)(24));
FA_ff_16006:FAff port map(x=>p(385)(24),y=>p(386)(24),Cin=>p(387)(24),clock=>clock,reset=>reset,s=>p(388)(24),cout=>p(389)(25));
FA_ff_16007:FAff port map(x=>p(385)(25),y=>p(386)(25),Cin=>p(387)(25),clock=>clock,reset=>reset,s=>p(388)(25),cout=>p(389)(26));
FA_ff_16008:FAff port map(x=>p(385)(26),y=>p(386)(26),Cin=>p(387)(26),clock=>clock,reset=>reset,s=>p(388)(26),cout=>p(389)(27));
FA_ff_16009:FAff port map(x=>p(385)(27),y=>p(386)(27),Cin=>p(387)(27),clock=>clock,reset=>reset,s=>p(388)(27),cout=>p(389)(28));
FA_ff_16010:FAff port map(x=>p(385)(28),y=>p(386)(28),Cin=>p(387)(28),clock=>clock,reset=>reset,s=>p(388)(28),cout=>p(389)(29));
FA_ff_16011:FAff port map(x=>p(385)(29),y=>p(386)(29),Cin=>p(387)(29),clock=>clock,reset=>reset,s=>p(388)(29),cout=>p(389)(30));
FA_ff_16012:FAff port map(x=>p(385)(30),y=>p(386)(30),Cin=>p(387)(30),clock=>clock,reset=>reset,s=>p(388)(30),cout=>p(389)(31));
FA_ff_16013:FAff port map(x=>p(385)(31),y=>p(386)(31),Cin=>p(387)(31),clock=>clock,reset=>reset,s=>p(388)(31),cout=>p(389)(32));
FA_ff_16014:FAff port map(x=>p(385)(32),y=>p(386)(32),Cin=>p(387)(32),clock=>clock,reset=>reset,s=>p(388)(32),cout=>p(389)(33));
FA_ff_16015:FAff port map(x=>p(385)(33),y=>p(386)(33),Cin=>p(387)(33),clock=>clock,reset=>reset,s=>p(388)(33),cout=>p(389)(34));
FA_ff_16016:FAff port map(x=>p(385)(34),y=>p(386)(34),Cin=>p(387)(34),clock=>clock,reset=>reset,s=>p(388)(34),cout=>p(389)(35));
FA_ff_16017:FAff port map(x=>p(385)(35),y=>p(386)(35),Cin=>p(387)(35),clock=>clock,reset=>reset,s=>p(388)(35),cout=>p(389)(36));
FA_ff_16018:FAff port map(x=>p(385)(36),y=>p(386)(36),Cin=>p(387)(36),clock=>clock,reset=>reset,s=>p(388)(36),cout=>p(389)(37));
FA_ff_16019:FAff port map(x=>p(385)(37),y=>p(386)(37),Cin=>p(387)(37),clock=>clock,reset=>reset,s=>p(388)(37),cout=>p(389)(38));
FA_ff_16020:FAff port map(x=>p(385)(38),y=>p(386)(38),Cin=>p(387)(38),clock=>clock,reset=>reset,s=>p(388)(38),cout=>p(389)(39));
FA_ff_16021:FAff port map(x=>p(385)(39),y=>p(386)(39),Cin=>p(387)(39),clock=>clock,reset=>reset,s=>p(388)(39),cout=>p(389)(40));
FA_ff_16022:FAff port map(x=>p(385)(40),y=>p(386)(40),Cin=>p(387)(40),clock=>clock,reset=>reset,s=>p(388)(40),cout=>p(389)(41));
FA_ff_16023:FAff port map(x=>p(385)(41),y=>p(386)(41),Cin=>p(387)(41),clock=>clock,reset=>reset,s=>p(388)(41),cout=>p(389)(42));
FA_ff_16024:FAff port map(x=>p(385)(42),y=>p(386)(42),Cin=>p(387)(42),clock=>clock,reset=>reset,s=>p(388)(42),cout=>p(389)(43));
FA_ff_16025:FAff port map(x=>p(385)(43),y=>p(386)(43),Cin=>p(387)(43),clock=>clock,reset=>reset,s=>p(388)(43),cout=>p(389)(44));
FA_ff_16026:FAff port map(x=>p(385)(44),y=>p(386)(44),Cin=>p(387)(44),clock=>clock,reset=>reset,s=>p(388)(44),cout=>p(389)(45));
FA_ff_16027:FAff port map(x=>p(385)(45),y=>p(386)(45),Cin=>p(387)(45),clock=>clock,reset=>reset,s=>p(388)(45),cout=>p(389)(46));
FA_ff_16028:FAff port map(x=>p(385)(46),y=>p(386)(46),Cin=>p(387)(46),clock=>clock,reset=>reset,s=>p(388)(46),cout=>p(389)(47));
FA_ff_16029:FAff port map(x=>p(385)(47),y=>p(386)(47),Cin=>p(387)(47),clock=>clock,reset=>reset,s=>p(388)(47),cout=>p(389)(48));
FA_ff_16030:FAff port map(x=>p(385)(48),y=>p(386)(48),Cin=>p(387)(48),clock=>clock,reset=>reset,s=>p(388)(48),cout=>p(389)(49));
FA_ff_16031:FAff port map(x=>p(385)(49),y=>p(386)(49),Cin=>p(387)(49),clock=>clock,reset=>reset,s=>p(388)(49),cout=>p(389)(50));
FA_ff_16032:FAff port map(x=>p(385)(50),y=>p(386)(50),Cin=>p(387)(50),clock=>clock,reset=>reset,s=>p(388)(50),cout=>p(389)(51));
FA_ff_16033:FAff port map(x=>p(385)(51),y=>p(386)(51),Cin=>p(387)(51),clock=>clock,reset=>reset,s=>p(388)(51),cout=>p(389)(52));
FA_ff_16034:FAff port map(x=>p(385)(52),y=>p(386)(52),Cin=>p(387)(52),clock=>clock,reset=>reset,s=>p(388)(52),cout=>p(389)(53));
FA_ff_16035:FAff port map(x=>p(385)(53),y=>p(386)(53),Cin=>p(387)(53),clock=>clock,reset=>reset,s=>p(388)(53),cout=>p(389)(54));
FA_ff_16036:FAff port map(x=>p(385)(54),y=>p(386)(54),Cin=>p(387)(54),clock=>clock,reset=>reset,s=>p(388)(54),cout=>p(389)(55));
FA_ff_16037:FAff port map(x=>p(385)(55),y=>p(386)(55),Cin=>p(387)(55),clock=>clock,reset=>reset,s=>p(388)(55),cout=>p(389)(56));
FA_ff_16038:FAff port map(x=>p(385)(56),y=>p(386)(56),Cin=>p(387)(56),clock=>clock,reset=>reset,s=>p(388)(56),cout=>p(389)(57));
FA_ff_16039:FAff port map(x=>p(385)(57),y=>p(386)(57),Cin=>p(387)(57),clock=>clock,reset=>reset,s=>p(388)(57),cout=>p(389)(58));
FA_ff_16040:FAff port map(x=>p(385)(58),y=>p(386)(58),Cin=>p(387)(58),clock=>clock,reset=>reset,s=>p(388)(58),cout=>p(389)(59));
FA_ff_16041:FAff port map(x=>p(385)(59),y=>p(386)(59),Cin=>p(387)(59),clock=>clock,reset=>reset,s=>p(388)(59),cout=>p(389)(60));
FA_ff_16042:FAff port map(x=>p(385)(60),y=>p(386)(60),Cin=>p(387)(60),clock=>clock,reset=>reset,s=>p(388)(60),cout=>p(389)(61));
FA_ff_16043:FAff port map(x=>p(385)(61),y=>p(386)(61),Cin=>p(387)(61),clock=>clock,reset=>reset,s=>p(388)(61),cout=>p(389)(62));
FA_ff_16044:FAff port map(x=>p(385)(62),y=>p(386)(62),Cin=>p(387)(62),clock=>clock,reset=>reset,s=>p(388)(62),cout=>p(389)(63));
FA_ff_16045:FAff port map(x=>p(385)(63),y=>p(386)(63),Cin=>p(387)(63),clock=>clock,reset=>reset,s=>p(388)(63),cout=>p(389)(64));
FA_ff_16046:FAff port map(x=>p(385)(64),y=>p(386)(64),Cin=>p(387)(64),clock=>clock,reset=>reset,s=>p(388)(64),cout=>p(389)(65));
FA_ff_16047:FAff port map(x=>p(385)(65),y=>p(386)(65),Cin=>p(387)(65),clock=>clock,reset=>reset,s=>p(388)(65),cout=>p(389)(66));
FA_ff_16048:FAff port map(x=>p(385)(66),y=>p(386)(66),Cin=>p(387)(66),clock=>clock,reset=>reset,s=>p(388)(66),cout=>p(389)(67));
FA_ff_16049:FAff port map(x=>p(385)(67),y=>p(386)(67),Cin=>p(387)(67),clock=>clock,reset=>reset,s=>p(388)(67),cout=>p(389)(68));
FA_ff_16050:FAff port map(x=>p(385)(68),y=>p(386)(68),Cin=>p(387)(68),clock=>clock,reset=>reset,s=>p(388)(68),cout=>p(389)(69));
FA_ff_16051:FAff port map(x=>p(385)(69),y=>p(386)(69),Cin=>p(387)(69),clock=>clock,reset=>reset,s=>p(388)(69),cout=>p(389)(70));
FA_ff_16052:FAff port map(x=>p(385)(70),y=>p(386)(70),Cin=>p(387)(70),clock=>clock,reset=>reset,s=>p(388)(70),cout=>p(389)(71));
FA_ff_16053:FAff port map(x=>p(385)(71),y=>p(386)(71),Cin=>p(387)(71),clock=>clock,reset=>reset,s=>p(388)(71),cout=>p(389)(72));
FA_ff_16054:FAff port map(x=>p(385)(72),y=>p(386)(72),Cin=>p(387)(72),clock=>clock,reset=>reset,s=>p(388)(72),cout=>p(389)(73));
FA_ff_16055:FAff port map(x=>p(385)(73),y=>p(386)(73),Cin=>p(387)(73),clock=>clock,reset=>reset,s=>p(388)(73),cout=>p(389)(74));
FA_ff_16056:FAff port map(x=>p(385)(74),y=>p(386)(74),Cin=>p(387)(74),clock=>clock,reset=>reset,s=>p(388)(74),cout=>p(389)(75));
FA_ff_16057:FAff port map(x=>p(385)(75),y=>p(386)(75),Cin=>p(387)(75),clock=>clock,reset=>reset,s=>p(388)(75),cout=>p(389)(76));
FA_ff_16058:FAff port map(x=>p(385)(76),y=>p(386)(76),Cin=>p(387)(76),clock=>clock,reset=>reset,s=>p(388)(76),cout=>p(389)(77));
FA_ff_16059:FAff port map(x=>p(385)(77),y=>p(386)(77),Cin=>p(387)(77),clock=>clock,reset=>reset,s=>p(388)(77),cout=>p(389)(78));
FA_ff_16060:FAff port map(x=>p(385)(78),y=>p(386)(78),Cin=>p(387)(78),clock=>clock,reset=>reset,s=>p(388)(78),cout=>p(389)(79));
FA_ff_16061:FAff port map(x=>p(385)(79),y=>p(386)(79),Cin=>p(387)(79),clock=>clock,reset=>reset,s=>p(388)(79),cout=>p(389)(80));
FA_ff_16062:FAff port map(x=>p(385)(80),y=>p(386)(80),Cin=>p(387)(80),clock=>clock,reset=>reset,s=>p(388)(80),cout=>p(389)(81));
FA_ff_16063:FAff port map(x=>p(385)(81),y=>p(386)(81),Cin=>p(387)(81),clock=>clock,reset=>reset,s=>p(388)(81),cout=>p(389)(82));
FA_ff_16064:FAff port map(x=>p(385)(82),y=>p(386)(82),Cin=>p(387)(82),clock=>clock,reset=>reset,s=>p(388)(82),cout=>p(389)(83));
FA_ff_16065:FAff port map(x=>p(385)(83),y=>p(386)(83),Cin=>p(387)(83),clock=>clock,reset=>reset,s=>p(388)(83),cout=>p(389)(84));
FA_ff_16066:FAff port map(x=>p(385)(84),y=>p(386)(84),Cin=>p(387)(84),clock=>clock,reset=>reset,s=>p(388)(84),cout=>p(389)(85));
FA_ff_16067:FAff port map(x=>p(385)(85),y=>p(386)(85),Cin=>p(387)(85),clock=>clock,reset=>reset,s=>p(388)(85),cout=>p(389)(86));
FA_ff_16068:FAff port map(x=>p(385)(86),y=>p(386)(86),Cin=>p(387)(86),clock=>clock,reset=>reset,s=>p(388)(86),cout=>p(389)(87));
FA_ff_16069:FAff port map(x=>p(385)(87),y=>p(386)(87),Cin=>p(387)(87),clock=>clock,reset=>reset,s=>p(388)(87),cout=>p(389)(88));
FA_ff_16070:FAff port map(x=>p(385)(88),y=>p(386)(88),Cin=>p(387)(88),clock=>clock,reset=>reset,s=>p(388)(88),cout=>p(389)(89));
FA_ff_16071:FAff port map(x=>p(385)(89),y=>p(386)(89),Cin=>p(387)(89),clock=>clock,reset=>reset,s=>p(388)(89),cout=>p(389)(90));
FA_ff_16072:FAff port map(x=>p(385)(90),y=>p(386)(90),Cin=>p(387)(90),clock=>clock,reset=>reset,s=>p(388)(90),cout=>p(389)(91));
FA_ff_16073:FAff port map(x=>p(385)(91),y=>p(386)(91),Cin=>p(387)(91),clock=>clock,reset=>reset,s=>p(388)(91),cout=>p(389)(92));
FA_ff_16074:FAff port map(x=>p(385)(92),y=>p(386)(92),Cin=>p(387)(92),clock=>clock,reset=>reset,s=>p(388)(92),cout=>p(389)(93));
FA_ff_16075:FAff port map(x=>p(385)(93),y=>p(386)(93),Cin=>p(387)(93),clock=>clock,reset=>reset,s=>p(388)(93),cout=>p(389)(94));
FA_ff_16076:FAff port map(x=>p(385)(94),y=>p(386)(94),Cin=>p(387)(94),clock=>clock,reset=>reset,s=>p(388)(94),cout=>p(389)(95));
FA_ff_16077:FAff port map(x=>p(385)(95),y=>p(386)(95),Cin=>p(387)(95),clock=>clock,reset=>reset,s=>p(388)(95),cout=>p(389)(96));
FA_ff_16078:FAff port map(x=>p(385)(96),y=>p(386)(96),Cin=>p(387)(96),clock=>clock,reset=>reset,s=>p(388)(96),cout=>p(389)(97));
FA_ff_16079:FAff port map(x=>p(385)(97),y=>p(386)(97),Cin=>p(387)(97),clock=>clock,reset=>reset,s=>p(388)(97),cout=>p(389)(98));
FA_ff_16080:FAff port map(x=>p(385)(98),y=>p(386)(98),Cin=>p(387)(98),clock=>clock,reset=>reset,s=>p(388)(98),cout=>p(389)(99));
FA_ff_16081:FAff port map(x=>p(385)(99),y=>p(386)(99),Cin=>p(387)(99),clock=>clock,reset=>reset,s=>p(388)(99),cout=>p(389)(100));
FA_ff_16082:FAff port map(x=>p(385)(100),y=>p(386)(100),Cin=>p(387)(100),clock=>clock,reset=>reset,s=>p(388)(100),cout=>p(389)(101));
FA_ff_16083:FAff port map(x=>p(385)(101),y=>p(386)(101),Cin=>p(387)(101),clock=>clock,reset=>reset,s=>p(388)(101),cout=>p(389)(102));
FA_ff_16084:FAff port map(x=>p(385)(102),y=>p(386)(102),Cin=>p(387)(102),clock=>clock,reset=>reset,s=>p(388)(102),cout=>p(389)(103));
FA_ff_16085:FAff port map(x=>p(385)(103),y=>p(386)(103),Cin=>p(387)(103),clock=>clock,reset=>reset,s=>p(388)(103),cout=>p(389)(104));
FA_ff_16086:FAff port map(x=>p(385)(104),y=>p(386)(104),Cin=>p(387)(104),clock=>clock,reset=>reset,s=>p(388)(104),cout=>p(389)(105));
FA_ff_16087:FAff port map(x=>p(385)(105),y=>p(386)(105),Cin=>p(387)(105),clock=>clock,reset=>reset,s=>p(388)(105),cout=>p(389)(106));
FA_ff_16088:FAff port map(x=>p(385)(106),y=>p(386)(106),Cin=>p(387)(106),clock=>clock,reset=>reset,s=>p(388)(106),cout=>p(389)(107));
FA_ff_16089:FAff port map(x=>p(385)(107),y=>p(386)(107),Cin=>p(387)(107),clock=>clock,reset=>reset,s=>p(388)(107),cout=>p(389)(108));
FA_ff_16090:FAff port map(x=>p(385)(108),y=>p(386)(108),Cin=>p(387)(108),clock=>clock,reset=>reset,s=>p(388)(108),cout=>p(389)(109));
FA_ff_16091:FAff port map(x=>p(385)(109),y=>p(386)(109),Cin=>p(387)(109),clock=>clock,reset=>reset,s=>p(388)(109),cout=>p(389)(110));
FA_ff_16092:FAff port map(x=>p(385)(110),y=>p(386)(110),Cin=>p(387)(110),clock=>clock,reset=>reset,s=>p(388)(110),cout=>p(389)(111));
FA_ff_16093:FAff port map(x=>p(385)(111),y=>p(386)(111),Cin=>p(387)(111),clock=>clock,reset=>reset,s=>p(388)(111),cout=>p(389)(112));
FA_ff_16094:FAff port map(x=>p(385)(112),y=>p(386)(112),Cin=>p(387)(112),clock=>clock,reset=>reset,s=>p(388)(112),cout=>p(389)(113));
FA_ff_16095:FAff port map(x=>p(385)(113),y=>p(386)(113),Cin=>p(387)(113),clock=>clock,reset=>reset,s=>p(388)(113),cout=>p(389)(114));
FA_ff_16096:FAff port map(x=>p(385)(114),y=>p(386)(114),Cin=>p(387)(114),clock=>clock,reset=>reset,s=>p(388)(114),cout=>p(389)(115));
FA_ff_16097:FAff port map(x=>p(385)(115),y=>p(386)(115),Cin=>p(387)(115),clock=>clock,reset=>reset,s=>p(388)(115),cout=>p(389)(116));
FA_ff_16098:FAff port map(x=>p(385)(116),y=>p(386)(116),Cin=>p(387)(116),clock=>clock,reset=>reset,s=>p(388)(116),cout=>p(389)(117));
FA_ff_16099:FAff port map(x=>p(385)(117),y=>p(386)(117),Cin=>p(387)(117),clock=>clock,reset=>reset,s=>p(388)(117),cout=>p(389)(118));
FA_ff_16100:FAff port map(x=>p(385)(118),y=>p(386)(118),Cin=>p(387)(118),clock=>clock,reset=>reset,s=>p(388)(118),cout=>p(389)(119));
FA_ff_16101:FAff port map(x=>p(385)(119),y=>p(386)(119),Cin=>p(387)(119),clock=>clock,reset=>reset,s=>p(388)(119),cout=>p(389)(120));
FA_ff_16102:FAff port map(x=>p(385)(120),y=>p(386)(120),Cin=>p(387)(120),clock=>clock,reset=>reset,s=>p(388)(120),cout=>p(389)(121));
FA_ff_16103:FAff port map(x=>p(385)(121),y=>p(386)(121),Cin=>p(387)(121),clock=>clock,reset=>reset,s=>p(388)(121),cout=>p(389)(122));
FA_ff_16104:FAff port map(x=>p(385)(122),y=>p(386)(122),Cin=>p(387)(122),clock=>clock,reset=>reset,s=>p(388)(122),cout=>p(389)(123));
FA_ff_16105:FAff port map(x=>p(385)(123),y=>p(386)(123),Cin=>p(387)(123),clock=>clock,reset=>reset,s=>p(388)(123),cout=>p(389)(124));
FA_ff_16106:FAff port map(x=>p(385)(124),y=>p(386)(124),Cin=>p(387)(124),clock=>clock,reset=>reset,s=>p(388)(124),cout=>p(389)(125));
FA_ff_16107:FAff port map(x=>p(385)(125),y=>p(386)(125),Cin=>p(387)(125),clock=>clock,reset=>reset,s=>p(388)(125),cout=>p(389)(126));
FA_ff_16108:FAff port map(x=>p(385)(126),y=>p(386)(126),Cin=>p(387)(126),clock=>clock,reset=>reset,s=>p(388)(126),cout=>p(389)(127));
FA_ff_16109:FAff port map(x=>p(385)(127),y=>p(386)(127),Cin=>p(387)(127),clock=>clock,reset=>reset,s=>p(388)(127),cout=>p(389)(128));
FA_ff_16110:FAff port map(x=>p(385)(128),y=>p(386)(128),Cin=>p(387)(128),clock=>clock,reset=>reset,s=>p(388)(128),cout=>p(389)(129));
FA_ff_16111:FAff port map(x=>p(385)(129),y=>p(386)(129),Cin=>p(387)(129),clock=>clock,reset=>reset,s=>p(388)(129),cout=>p(389)(130));
FA_ff_16112:FAff port map(x=>p(385)(130),y=>p(386)(130),Cin=>p(387)(130),clock=>clock,reset=>reset,s=>p(388)(130),cout=>p(389)(131));
FA_ff_16113:FAff port map(x=>p(385)(131),y=>p(386)(131),Cin=>p(387)(131),clock=>clock,reset=>reset,s=>p(388)(131),cout=>p(389)(132));
FA_ff_16114:FAff port map(x=>p(385)(132),y=>p(386)(132),Cin=>p(387)(132),clock=>clock,reset=>reset,s=>p(388)(132),cout=>p(389)(133));
FA_ff_16115:FAff port map(x=>p(385)(133),y=>p(386)(133),Cin=>p(387)(133),clock=>clock,reset=>reset,s=>p(388)(133),cout=>p(389)(134));
p(388)(134)<=p(386)(134);
res(0)<=p(388)(0);
res(1)<=p(388)(1);
add1(0)<=p(388)(2);
add2(0)<=p(389)(2);
add1(1)<=p(388)(3);
add2(1)<=p(389)(3);
add1(2)<=p(388)(4);
add2(2)<=p(389)(4);
add1(3)<=p(388)(5);
add2(3)<=p(389)(5);
add1(4)<=p(388)(6);
add2(4)<=p(389)(6);
add1(5)<=p(388)(7);
add2(5)<=p(389)(7);
add1(6)<=p(388)(8);
add2(6)<=p(389)(8);
add1(7)<=p(388)(9);
add2(7)<=p(389)(9);
add1(8)<=p(388)(10);
add2(8)<=p(389)(10);
add1(9)<=p(388)(11);
add2(9)<=p(389)(11);
add1(10)<=p(388)(12);
add2(10)<=p(389)(12);
add1(11)<=p(388)(13);
add2(11)<=p(389)(13);
add1(12)<=p(388)(14);
add2(12)<=p(389)(14);
add1(13)<=p(388)(15);
add2(13)<=p(389)(15);
add1(14)<=p(388)(16);
add2(14)<=p(389)(16);
add1(15)<=p(388)(17);
add2(15)<=p(389)(17);
add1(16)<=p(388)(18);
add2(16)<=p(389)(18);
add1(17)<=p(388)(19);
add2(17)<=p(389)(19);
add1(18)<=p(388)(20);
add2(18)<=p(389)(20);
add1(19)<=p(388)(21);
add2(19)<=p(389)(21);
add1(20)<=p(388)(22);
add2(20)<=p(389)(22);
add1(21)<=p(388)(23);
add2(21)<=p(389)(23);
add1(22)<=p(388)(24);
add2(22)<=p(389)(24);
add1(23)<=p(388)(25);
add2(23)<=p(389)(25);
add1(24)<=p(388)(26);
add2(24)<=p(389)(26);
add1(25)<=p(388)(27);
add2(25)<=p(389)(27);
add1(26)<=p(388)(28);
add2(26)<=p(389)(28);
add1(27)<=p(388)(29);
add2(27)<=p(389)(29);
add1(28)<=p(388)(30);
add2(28)<=p(389)(30);
add1(29)<=p(388)(31);
add2(29)<=p(389)(31);
add1(30)<=p(388)(32);
add2(30)<=p(389)(32);
add1(31)<=p(388)(33);
add2(31)<=p(389)(33);
add1(32)<=p(388)(34);
add2(32)<=p(389)(34);
add1(33)<=p(388)(35);
add2(33)<=p(389)(35);
add1(34)<=p(388)(36);
add2(34)<=p(389)(36);
add1(35)<=p(388)(37);
add2(35)<=p(389)(37);
add1(36)<=p(388)(38);
add2(36)<=p(389)(38);
add1(37)<=p(388)(39);
add2(37)<=p(389)(39);
add1(38)<=p(388)(40);
add2(38)<=p(389)(40);
add1(39)<=p(388)(41);
add2(39)<=p(389)(41);
add1(40)<=p(388)(42);
add2(40)<=p(389)(42);
add1(41)<=p(388)(43);
add2(41)<=p(389)(43);
add1(42)<=p(388)(44);
add2(42)<=p(389)(44);
add1(43)<=p(388)(45);
add2(43)<=p(389)(45);
add1(44)<=p(388)(46);
add2(44)<=p(389)(46);
add1(45)<=p(388)(47);
add2(45)<=p(389)(47);
add1(46)<=p(388)(48);
add2(46)<=p(389)(48);
add1(47)<=p(388)(49);
add2(47)<=p(389)(49);
add1(48)<=p(388)(50);
add2(48)<=p(389)(50);
add1(49)<=p(388)(51);
add2(49)<=p(389)(51);
add1(50)<=p(388)(52);
add2(50)<=p(389)(52);
add1(51)<=p(388)(53);
add2(51)<=p(389)(53);
add1(52)<=p(388)(54);
add2(52)<=p(389)(54);
add1(53)<=p(388)(55);
add2(53)<=p(389)(55);
add1(54)<=p(388)(56);
add2(54)<=p(389)(56);
add1(55)<=p(388)(57);
add2(55)<=p(389)(57);
add1(56)<=p(388)(58);
add2(56)<=p(389)(58);
add1(57)<=p(388)(59);
add2(57)<=p(389)(59);
add1(58)<=p(388)(60);
add2(58)<=p(389)(60);
add1(59)<=p(388)(61);
add2(59)<=p(389)(61);
add1(60)<=p(388)(62);
add2(60)<=p(389)(62);
add1(61)<=p(388)(63);
add2(61)<=p(389)(63);
add1(62)<=p(388)(64);
add2(62)<=p(389)(64);
add1(63)<=p(388)(65);
add2(63)<=p(389)(65);
add1(64)<=p(388)(66);
add2(64)<=p(389)(66);
add1(65)<=p(388)(67);
add2(65)<=p(389)(67);
add1(66)<=p(388)(68);
add2(66)<=p(389)(68);
add1(67)<=p(388)(69);
add2(67)<=p(389)(69);
add1(68)<=p(388)(70);
add2(68)<=p(389)(70);
add1(69)<=p(388)(71);
add2(69)<=p(389)(71);
add1(70)<=p(388)(72);
add2(70)<=p(389)(72);
add1(71)<=p(388)(73);
add2(71)<=p(389)(73);
add1(72)<=p(388)(74);
add2(72)<=p(389)(74);
add1(73)<=p(388)(75);
add2(73)<=p(389)(75);
add1(74)<=p(388)(76);
add2(74)<=p(389)(76);
add1(75)<=p(388)(77);
add2(75)<=p(389)(77);
add1(76)<=p(388)(78);
add2(76)<=p(389)(78);
add1(77)<=p(388)(79);
add2(77)<=p(389)(79);
add1(78)<=p(388)(80);
add2(78)<=p(389)(80);
add1(79)<=p(388)(81);
add2(79)<=p(389)(81);
add1(80)<=p(388)(82);
add2(80)<=p(389)(82);
add1(81)<=p(388)(83);
add2(81)<=p(389)(83);
add1(82)<=p(388)(84);
add2(82)<=p(389)(84);
add1(83)<=p(388)(85);
add2(83)<=p(389)(85);
add1(84)<=p(388)(86);
add2(84)<=p(389)(86);
add1(85)<=p(388)(87);
add2(85)<=p(389)(87);
add1(86)<=p(388)(88);
add2(86)<=p(389)(88);
add1(87)<=p(388)(89);
add2(87)<=p(389)(89);
add1(88)<=p(388)(90);
add2(88)<=p(389)(90);
add1(89)<=p(388)(91);
add2(89)<=p(389)(91);
add1(90)<=p(388)(92);
add2(90)<=p(389)(92);
add1(91)<=p(388)(93);
add2(91)<=p(389)(93);
add1(92)<=p(388)(94);
add2(92)<=p(389)(94);
add1(93)<=p(388)(95);
add2(93)<=p(389)(95);
add1(94)<=p(388)(96);
add2(94)<=p(389)(96);
add1(95)<=p(388)(97);
add2(95)<=p(389)(97);
add1(96)<=p(388)(98);
add2(96)<=p(389)(98);
add1(97)<=p(388)(99);
add2(97)<=p(389)(99);
add1(98)<=p(388)(100);
add2(98)<=p(389)(100);
add1(99)<=p(388)(101);
add2(99)<=p(389)(101);
add1(100)<=p(388)(102);
add2(100)<=p(389)(102);
add1(101)<=p(388)(103);
add2(101)<=p(389)(103);
add1(102)<=p(388)(104);
add2(102)<=p(389)(104);
add1(103)<=p(388)(105);
add2(103)<=p(389)(105);
add1(104)<=p(388)(106);
add2(104)<=p(389)(106);
add1(105)<=p(388)(107);
add2(105)<=p(389)(107);
add1(106)<=p(388)(108);
add2(106)<=p(389)(108);
add1(107)<=p(388)(109);
add2(107)<=p(389)(109);
add1(108)<=p(388)(110);
add2(108)<=p(389)(110);
add1(109)<=p(388)(111);
add2(109)<=p(389)(111);
add1(110)<=p(388)(112);
add2(110)<=p(389)(112);
add1(111)<=p(388)(113);
add2(111)<=p(389)(113);
add1(112)<=p(388)(114);
add2(112)<=p(389)(114);
add1(113)<=p(388)(115);
add2(113)<=p(389)(115);
add1(114)<=p(388)(116);
add2(114)<=p(389)(116);
add1(115)<=p(388)(117);
add2(115)<=p(389)(117);
add1(116)<=p(388)(118);
add2(116)<=p(389)(118);
add1(117)<=p(388)(119);
add2(117)<=p(389)(119);
add1(118)<=p(388)(120);
add2(118)<=p(389)(120);
add1(119)<=p(388)(121);
add2(119)<=p(389)(121);
add1(120)<=p(388)(122);
add2(120)<=p(389)(122);
add1(121)<=p(388)(123);
add2(121)<=p(389)(123);
add1(122)<=p(388)(124);
add2(122)<=p(389)(124);
add1(123)<=p(388)(125);
add2(123)<=p(389)(125);
add1(124)<=p(388)(126);
add2(124)<=p(389)(126);
add1(125)<=p(388)(127);
add2(125)<=p(389)(127);
add1(126)<=p(388)(128);
add2(126)<=p(389)(128);
add1(127)<=p(388)(129);
add2(127)<=p(389)(129);
add1(128)<=p(388)(130);
add2(128)<=p(389)(130);
add1(129)<=p(388)(131);
add2(129)<=p(389)(131);
add1(130)<=p(388)(132);
add2(130)<=p(389)(132);
add1(131)<=p(388)(133);
add2(131)<=p(389)(133);
add1(132)<=p(388)(134);
add2(132)<=p(389)(134);
end architecture behavioural;