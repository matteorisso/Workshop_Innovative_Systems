library verilog;
use verilog.vl_types.all;
entity globals_sv is
end globals_sv;
