
module SNPS_CLOCK_GATE_HIGH_avr_pooling_fsm ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(ENCLK) );
endmodule


module avr_pooling_unrolled ( clk, rst_fsm, start, done, en, size_1, size_2, 
        pool_sel, d_0, d_1, d_2, d_3, d_4, d_5, d_6, d_7, o_pool_1, o_pool_2, 
        o_pool_3, o_pool_4 );
  input [4:0] size_1;
  input [4:0] size_2;
  input [15:0] d_0;
  input [15:0] d_1;
  input [15:0] d_2;
  input [15:0] d_3;
  input [15:0] d_4;
  input [15:0] d_5;
  input [15:0] d_6;
  input [15:0] d_7;
  output [15:0] o_pool_1;
  output [15:0] o_pool_2;
  output [15:0] o_pool_3;
  output [15:0] o_pool_4;
  input clk, rst_fsm, start, done, en, pool_sel;
  wire   pool_ld_h, pool_rst_cnt_r, pool_rst_cnt_c, pool_tc, pool_en_cnt,
         pool_rst_cnt, pool_sync_clr, pool_sel0, pool_pool_cnt_0_,
         pool_pool_cnt_1_, pool_pool_interface_mux_0_n9,
         pool_pool_interface_mux_0_n8, pool_pool_interface_mux_0_n7,
         pool_pool_interface_mux_0_n6, pool_pool_interface_mux_0_n5,
         pool_pool_interface_mux_0_n4, pool_pool_interface_mux_0_n3,
         pool_pool_interface_mux_0_n2, pool_pool_interface_mux_0_n1,
         pool_pool_interface_mux_0_n33, pool_pool_interface_mux_0_n32,
         pool_pool_interface_mux_0_n31, pool_pool_interface_mux_0_n30,
         pool_pool_interface_mux_0_n29, pool_pool_interface_mux_0_n28,
         pool_pool_interface_mux_0_n27, pool_pool_interface_mux_0_n26,
         pool_pool_interface_mux_0_n25, pool_pool_interface_mux_0_n24,
         pool_pool_interface_mux_0_n23, pool_pool_interface_mux_0_n22,
         pool_pool_interface_mux_0_n21, pool_pool_interface_mux_0_n20,
         pool_pool_interface_mux_0_n19, pool_pool_interface_mux_0_n18,
         pool_pool_interface_mux_1_n57, pool_pool_interface_mux_1_n56,
         pool_pool_interface_mux_1_n55, pool_pool_interface_mux_1_n54,
         pool_pool_interface_mux_1_n53, pool_pool_interface_mux_1_n52,
         pool_pool_interface_mux_1_n51, pool_pool_interface_mux_1_n50,
         pool_pool_interface_mux_1_n49, pool_pool_interface_mux_1_n48,
         pool_pool_interface_mux_1_n47, pool_pool_interface_mux_1_n46,
         pool_pool_interface_mux_1_n45, pool_pool_interface_mux_1_n44,
         pool_pool_interface_mux_1_n43, pool_pool_interface_mux_1_n42,
         pool_pool_interface_mux_1_n9, pool_pool_interface_mux_1_n8,
         pool_pool_interface_mux_1_n7, pool_pool_interface_mux_1_n6,
         pool_pool_interface_mux_1_n5, pool_pool_interface_mux_1_n4,
         pool_pool_interface_mux_1_n3, pool_pool_interface_mux_1_n2,
         pool_pool_interface_mux_1_n1, pool_pool_interface_mux_2_n57,
         pool_pool_interface_mux_2_n56, pool_pool_interface_mux_2_n55,
         pool_pool_interface_mux_2_n54, pool_pool_interface_mux_2_n53,
         pool_pool_interface_mux_2_n52, pool_pool_interface_mux_2_n51,
         pool_pool_interface_mux_2_n50, pool_pool_interface_mux_2_n49,
         pool_pool_interface_mux_2_n48, pool_pool_interface_mux_2_n47,
         pool_pool_interface_mux_2_n46, pool_pool_interface_mux_2_n45,
         pool_pool_interface_mux_2_n44, pool_pool_interface_mux_2_n43,
         pool_pool_interface_mux_2_n42, pool_pool_interface_mux_2_n9,
         pool_pool_interface_mux_2_n8, pool_pool_interface_mux_2_n7,
         pool_pool_interface_mux_2_n6, pool_pool_interface_mux_2_n5,
         pool_pool_interface_mux_2_n4, pool_pool_interface_mux_2_n3,
         pool_pool_interface_mux_2_n2, pool_pool_interface_mux_2_n1,
         pool_pool_interface_mux_3_n57, pool_pool_interface_mux_3_n56,
         pool_pool_interface_mux_3_n55, pool_pool_interface_mux_3_n54,
         pool_pool_interface_mux_3_n53, pool_pool_interface_mux_3_n52,
         pool_pool_interface_mux_3_n51, pool_pool_interface_mux_3_n50,
         pool_pool_interface_mux_3_n49, pool_pool_interface_mux_3_n48,
         pool_pool_interface_mux_3_n47, pool_pool_interface_mux_3_n46,
         pool_pool_interface_mux_3_n45, pool_pool_interface_mux_3_n44,
         pool_pool_interface_mux_3_n43, pool_pool_interface_mux_3_n42,
         pool_pool_interface_mux_3_n9, pool_pool_interface_mux_3_n8,
         pool_pool_interface_mux_3_n7, pool_pool_interface_mux_3_n6,
         pool_pool_interface_mux_3_n5, pool_pool_interface_mux_3_n4,
         pool_pool_interface_mux_3_n3, pool_pool_interface_mux_3_n2,
         pool_pool_interface_mux_3_n1, pool_pool_pe_b_n7, pool_pool_pe_b_n6,
         pool_pool_pe_b_n1, pool_pool_pe_b_n5, pool_pool_pe_b_n4,
         pool_pool_pe_b_n3, pool_pool_pe_b_n2, pool_pool_pe_b_peij_0_0_n14,
         pool_pool_pe_b_peij_0_0_n12, pool_pool_pe_b_peij_0_0_n11,
         pool_pool_pe_b_peij_0_0_n10, pool_pool_pe_b_peij_0_0_n9,
         pool_pool_pe_b_peij_0_0_n8, pool_pool_pe_b_peij_0_0_n7,
         pool_pool_pe_b_peij_0_0_n6, pool_pool_pe_b_peij_0_0_n5,
         pool_pool_pe_b_peij_0_0_n4, pool_pool_pe_b_peij_0_0_n3,
         pool_pool_pe_b_peij_0_0_n2, pool_pool_pe_b_peij_0_0_n1,
         pool_pool_pe_b_peij_0_0_q_k, pool_pool_pe_b_peij_0_0_gck,
         pool_pool_pe_b_peij_0_0_add_c_out,
         pool_pool_pe_b_peij_0_0_add_fai_0_n3,
         pool_pool_pe_b_peij_0_0_add_fai_0_n2,
         pool_pool_pe_b_peij_0_0_add_fai_1_n5,
         pool_pool_pe_b_peij_0_0_add_fai_1_n4,
         pool_pool_pe_b_peij_0_0_add_fai_2_n5,
         pool_pool_pe_b_peij_0_0_add_fai_2_n4,
         pool_pool_pe_b_peij_0_0_add_fai_3_n5,
         pool_pool_pe_b_peij_0_0_add_fai_3_n4,
         pool_pool_pe_b_peij_0_0_add_fai_4_n5,
         pool_pool_pe_b_peij_0_0_add_fai_4_n4,
         pool_pool_pe_b_peij_0_0_add_fai_5_n5,
         pool_pool_pe_b_peij_0_0_add_fai_5_n4,
         pool_pool_pe_b_peij_0_0_add_fai_6_n5,
         pool_pool_pe_b_peij_0_0_add_fai_6_n4,
         pool_pool_pe_b_peij_0_0_add_fai_7_n5,
         pool_pool_pe_b_peij_0_0_add_fai_7_n4,
         pool_pool_pe_b_peij_0_0_add_fai_8_n5,
         pool_pool_pe_b_peij_0_0_add_fai_8_n4,
         pool_pool_pe_b_peij_0_0_add_fai_9_n5,
         pool_pool_pe_b_peij_0_0_add_fai_9_n4,
         pool_pool_pe_b_peij_0_0_add_fai_10_n5,
         pool_pool_pe_b_peij_0_0_add_fai_10_n4, pool_pool_pe_b_peij_0_1_n14,
         pool_pool_pe_b_peij_0_1_n12, pool_pool_pe_b_peij_0_1_n11,
         pool_pool_pe_b_peij_0_1_n10, pool_pool_pe_b_peij_0_1_n9,
         pool_pool_pe_b_peij_0_1_n8, pool_pool_pe_b_peij_0_1_n7,
         pool_pool_pe_b_peij_0_1_n6, pool_pool_pe_b_peij_0_1_n5,
         pool_pool_pe_b_peij_0_1_n4, pool_pool_pe_b_peij_0_1_n3,
         pool_pool_pe_b_peij_0_1_n2, pool_pool_pe_b_peij_0_1_n1,
         pool_pool_pe_b_peij_0_1_q_k, pool_pool_pe_b_peij_0_1_gck,
         pool_pool_pe_b_peij_0_1_add_c_out,
         pool_pool_pe_b_peij_0_1_add_fai_0_n5,
         pool_pool_pe_b_peij_0_1_add_fai_0_n4,
         pool_pool_pe_b_peij_0_1_add_fai_1_n5,
         pool_pool_pe_b_peij_0_1_add_fai_1_n4,
         pool_pool_pe_b_peij_0_1_add_fai_2_n5,
         pool_pool_pe_b_peij_0_1_add_fai_2_n4,
         pool_pool_pe_b_peij_0_1_add_fai_3_n5,
         pool_pool_pe_b_peij_0_1_add_fai_3_n4,
         pool_pool_pe_b_peij_0_1_add_fai_4_n5,
         pool_pool_pe_b_peij_0_1_add_fai_4_n4,
         pool_pool_pe_b_peij_0_1_add_fai_5_n5,
         pool_pool_pe_b_peij_0_1_add_fai_5_n4,
         pool_pool_pe_b_peij_0_1_add_fai_6_n5,
         pool_pool_pe_b_peij_0_1_add_fai_6_n4,
         pool_pool_pe_b_peij_0_1_add_fai_7_n5,
         pool_pool_pe_b_peij_0_1_add_fai_7_n4,
         pool_pool_pe_b_peij_0_1_add_fai_8_n5,
         pool_pool_pe_b_peij_0_1_add_fai_8_n4,
         pool_pool_pe_b_peij_0_1_add_fai_9_n5,
         pool_pool_pe_b_peij_0_1_add_fai_9_n4,
         pool_pool_pe_b_peij_0_1_add_fai_10_n5,
         pool_pool_pe_b_peij_0_1_add_fai_10_n4, pool_pool_pe_b_peij_0_2_n14,
         pool_pool_pe_b_peij_0_2_n12, pool_pool_pe_b_peij_0_2_n11,
         pool_pool_pe_b_peij_0_2_n10, pool_pool_pe_b_peij_0_2_n9,
         pool_pool_pe_b_peij_0_2_n8, pool_pool_pe_b_peij_0_2_n7,
         pool_pool_pe_b_peij_0_2_n6, pool_pool_pe_b_peij_0_2_n5,
         pool_pool_pe_b_peij_0_2_n4, pool_pool_pe_b_peij_0_2_n3,
         pool_pool_pe_b_peij_0_2_n2, pool_pool_pe_b_peij_0_2_n1,
         pool_pool_pe_b_peij_0_2_q_k, pool_pool_pe_b_peij_0_2_gck,
         pool_pool_pe_b_peij_0_2_add_c_out,
         pool_pool_pe_b_peij_0_2_add_fai_0_n5,
         pool_pool_pe_b_peij_0_2_add_fai_0_n4,
         pool_pool_pe_b_peij_0_2_add_fai_1_n5,
         pool_pool_pe_b_peij_0_2_add_fai_1_n4,
         pool_pool_pe_b_peij_0_2_add_fai_2_n5,
         pool_pool_pe_b_peij_0_2_add_fai_2_n4,
         pool_pool_pe_b_peij_0_2_add_fai_3_n5,
         pool_pool_pe_b_peij_0_2_add_fai_3_n4,
         pool_pool_pe_b_peij_0_2_add_fai_4_n5,
         pool_pool_pe_b_peij_0_2_add_fai_4_n4,
         pool_pool_pe_b_peij_0_2_add_fai_5_n5,
         pool_pool_pe_b_peij_0_2_add_fai_5_n4,
         pool_pool_pe_b_peij_0_2_add_fai_6_n5,
         pool_pool_pe_b_peij_0_2_add_fai_6_n4,
         pool_pool_pe_b_peij_0_2_add_fai_7_n5,
         pool_pool_pe_b_peij_0_2_add_fai_7_n4,
         pool_pool_pe_b_peij_0_2_add_fai_8_n5,
         pool_pool_pe_b_peij_0_2_add_fai_8_n4,
         pool_pool_pe_b_peij_0_2_add_fai_9_n5,
         pool_pool_pe_b_peij_0_2_add_fai_9_n4,
         pool_pool_pe_b_peij_0_2_add_fai_10_n5,
         pool_pool_pe_b_peij_0_2_add_fai_10_n4, pool_pool_pe_b_peij_0_3_n14,
         pool_pool_pe_b_peij_0_3_n12, pool_pool_pe_b_peij_0_3_n11,
         pool_pool_pe_b_peij_0_3_n10, pool_pool_pe_b_peij_0_3_n9,
         pool_pool_pe_b_peij_0_3_n8, pool_pool_pe_b_peij_0_3_n7,
         pool_pool_pe_b_peij_0_3_n6, pool_pool_pe_b_peij_0_3_n5,
         pool_pool_pe_b_peij_0_3_n4, pool_pool_pe_b_peij_0_3_n3,
         pool_pool_pe_b_peij_0_3_n2, pool_pool_pe_b_peij_0_3_n1,
         pool_pool_pe_b_peij_0_3_q_k, pool_pool_pe_b_peij_0_3_gck,
         pool_pool_pe_b_peij_0_3_add_c_out,
         pool_pool_pe_b_peij_0_3_add_fai_0_n5,
         pool_pool_pe_b_peij_0_3_add_fai_0_n4,
         pool_pool_pe_b_peij_0_3_add_fai_1_n5,
         pool_pool_pe_b_peij_0_3_add_fai_1_n4,
         pool_pool_pe_b_peij_0_3_add_fai_2_n5,
         pool_pool_pe_b_peij_0_3_add_fai_2_n4,
         pool_pool_pe_b_peij_0_3_add_fai_3_n5,
         pool_pool_pe_b_peij_0_3_add_fai_3_n4,
         pool_pool_pe_b_peij_0_3_add_fai_4_n5,
         pool_pool_pe_b_peij_0_3_add_fai_4_n4,
         pool_pool_pe_b_peij_0_3_add_fai_5_n5,
         pool_pool_pe_b_peij_0_3_add_fai_5_n4,
         pool_pool_pe_b_peij_0_3_add_fai_6_n5,
         pool_pool_pe_b_peij_0_3_add_fai_6_n4,
         pool_pool_pe_b_peij_0_3_add_fai_7_n5,
         pool_pool_pe_b_peij_0_3_add_fai_7_n4,
         pool_pool_pe_b_peij_0_3_add_fai_8_n5,
         pool_pool_pe_b_peij_0_3_add_fai_8_n4,
         pool_pool_pe_b_peij_0_3_add_fai_9_n5,
         pool_pool_pe_b_peij_0_3_add_fai_9_n4,
         pool_pool_pe_b_peij_0_3_add_fai_10_n5,
         pool_pool_pe_b_peij_0_3_add_fai_10_n4, pool_pool_pe_b_peij_1_0_n14,
         pool_pool_pe_b_peij_1_0_n12, pool_pool_pe_b_peij_1_0_n11,
         pool_pool_pe_b_peij_1_0_n10, pool_pool_pe_b_peij_1_0_n9,
         pool_pool_pe_b_peij_1_0_n8, pool_pool_pe_b_peij_1_0_n7,
         pool_pool_pe_b_peij_1_0_n6, pool_pool_pe_b_peij_1_0_n5,
         pool_pool_pe_b_peij_1_0_n4, pool_pool_pe_b_peij_1_0_n3,
         pool_pool_pe_b_peij_1_0_n2, pool_pool_pe_b_peij_1_0_n1,
         pool_pool_pe_b_peij_1_0_q_k, pool_pool_pe_b_peij_1_0_gck,
         pool_pool_pe_b_peij_1_0_add_c_out,
         pool_pool_pe_b_peij_1_0_add_fai_0_n5,
         pool_pool_pe_b_peij_1_0_add_fai_0_n4,
         pool_pool_pe_b_peij_1_0_add_fai_1_n5,
         pool_pool_pe_b_peij_1_0_add_fai_1_n4,
         pool_pool_pe_b_peij_1_0_add_fai_2_n5,
         pool_pool_pe_b_peij_1_0_add_fai_2_n4,
         pool_pool_pe_b_peij_1_0_add_fai_3_n5,
         pool_pool_pe_b_peij_1_0_add_fai_3_n4,
         pool_pool_pe_b_peij_1_0_add_fai_4_n5,
         pool_pool_pe_b_peij_1_0_add_fai_4_n4,
         pool_pool_pe_b_peij_1_0_add_fai_5_n5,
         pool_pool_pe_b_peij_1_0_add_fai_5_n4,
         pool_pool_pe_b_peij_1_0_add_fai_6_n5,
         pool_pool_pe_b_peij_1_0_add_fai_6_n4,
         pool_pool_pe_b_peij_1_0_add_fai_7_n5,
         pool_pool_pe_b_peij_1_0_add_fai_7_n4,
         pool_pool_pe_b_peij_1_0_add_fai_8_n5,
         pool_pool_pe_b_peij_1_0_add_fai_8_n4,
         pool_pool_pe_b_peij_1_0_add_fai_9_n5,
         pool_pool_pe_b_peij_1_0_add_fai_9_n4,
         pool_pool_pe_b_peij_1_0_add_fai_10_n5,
         pool_pool_pe_b_peij_1_0_add_fai_10_n4, pool_pool_pe_b_peij_1_1_n14,
         pool_pool_pe_b_peij_1_1_n12, pool_pool_pe_b_peij_1_1_n11,
         pool_pool_pe_b_peij_1_1_n10, pool_pool_pe_b_peij_1_1_n9,
         pool_pool_pe_b_peij_1_1_n8, pool_pool_pe_b_peij_1_1_n7,
         pool_pool_pe_b_peij_1_1_n6, pool_pool_pe_b_peij_1_1_n5,
         pool_pool_pe_b_peij_1_1_n4, pool_pool_pe_b_peij_1_1_n3,
         pool_pool_pe_b_peij_1_1_n2, pool_pool_pe_b_peij_1_1_n1,
         pool_pool_pe_b_peij_1_1_q_k, pool_pool_pe_b_peij_1_1_gck,
         pool_pool_pe_b_peij_1_1_add_c_out,
         pool_pool_pe_b_peij_1_1_add_fai_0_n5,
         pool_pool_pe_b_peij_1_1_add_fai_0_n4,
         pool_pool_pe_b_peij_1_1_add_fai_1_n5,
         pool_pool_pe_b_peij_1_1_add_fai_1_n4,
         pool_pool_pe_b_peij_1_1_add_fai_2_n5,
         pool_pool_pe_b_peij_1_1_add_fai_2_n4,
         pool_pool_pe_b_peij_1_1_add_fai_3_n5,
         pool_pool_pe_b_peij_1_1_add_fai_3_n4,
         pool_pool_pe_b_peij_1_1_add_fai_4_n5,
         pool_pool_pe_b_peij_1_1_add_fai_4_n4,
         pool_pool_pe_b_peij_1_1_add_fai_5_n5,
         pool_pool_pe_b_peij_1_1_add_fai_5_n4,
         pool_pool_pe_b_peij_1_1_add_fai_6_n5,
         pool_pool_pe_b_peij_1_1_add_fai_6_n4,
         pool_pool_pe_b_peij_1_1_add_fai_7_n5,
         pool_pool_pe_b_peij_1_1_add_fai_7_n4,
         pool_pool_pe_b_peij_1_1_add_fai_8_n5,
         pool_pool_pe_b_peij_1_1_add_fai_8_n4,
         pool_pool_pe_b_peij_1_1_add_fai_9_n5,
         pool_pool_pe_b_peij_1_1_add_fai_9_n4,
         pool_pool_pe_b_peij_1_1_add_fai_10_n5,
         pool_pool_pe_b_peij_1_1_add_fai_10_n4, pool_pool_pe_b_peij_1_2_n14,
         pool_pool_pe_b_peij_1_2_n12, pool_pool_pe_b_peij_1_2_n11,
         pool_pool_pe_b_peij_1_2_n10, pool_pool_pe_b_peij_1_2_n9,
         pool_pool_pe_b_peij_1_2_n8, pool_pool_pe_b_peij_1_2_n7,
         pool_pool_pe_b_peij_1_2_n6, pool_pool_pe_b_peij_1_2_n5,
         pool_pool_pe_b_peij_1_2_n4, pool_pool_pe_b_peij_1_2_n3,
         pool_pool_pe_b_peij_1_2_n2, pool_pool_pe_b_peij_1_2_n1,
         pool_pool_pe_b_peij_1_2_q_k, pool_pool_pe_b_peij_1_2_gck,
         pool_pool_pe_b_peij_1_2_add_c_out,
         pool_pool_pe_b_peij_1_2_add_fai_0_n5,
         pool_pool_pe_b_peij_1_2_add_fai_0_n4,
         pool_pool_pe_b_peij_1_2_add_fai_1_n5,
         pool_pool_pe_b_peij_1_2_add_fai_1_n4,
         pool_pool_pe_b_peij_1_2_add_fai_2_n5,
         pool_pool_pe_b_peij_1_2_add_fai_2_n4,
         pool_pool_pe_b_peij_1_2_add_fai_3_n5,
         pool_pool_pe_b_peij_1_2_add_fai_3_n4,
         pool_pool_pe_b_peij_1_2_add_fai_4_n5,
         pool_pool_pe_b_peij_1_2_add_fai_4_n4,
         pool_pool_pe_b_peij_1_2_add_fai_5_n5,
         pool_pool_pe_b_peij_1_2_add_fai_5_n4,
         pool_pool_pe_b_peij_1_2_add_fai_6_n5,
         pool_pool_pe_b_peij_1_2_add_fai_6_n4,
         pool_pool_pe_b_peij_1_2_add_fai_7_n5,
         pool_pool_pe_b_peij_1_2_add_fai_7_n4,
         pool_pool_pe_b_peij_1_2_add_fai_8_n5,
         pool_pool_pe_b_peij_1_2_add_fai_8_n4,
         pool_pool_pe_b_peij_1_2_add_fai_9_n5,
         pool_pool_pe_b_peij_1_2_add_fai_9_n4,
         pool_pool_pe_b_peij_1_2_add_fai_10_n5,
         pool_pool_pe_b_peij_1_2_add_fai_10_n4, pool_pool_pe_b_peij_1_3_n14,
         pool_pool_pe_b_peij_1_3_n12, pool_pool_pe_b_peij_1_3_n11,
         pool_pool_pe_b_peij_1_3_n10, pool_pool_pe_b_peij_1_3_n9,
         pool_pool_pe_b_peij_1_3_n8, pool_pool_pe_b_peij_1_3_n7,
         pool_pool_pe_b_peij_1_3_n6, pool_pool_pe_b_peij_1_3_n5,
         pool_pool_pe_b_peij_1_3_n4, pool_pool_pe_b_peij_1_3_n3,
         pool_pool_pe_b_peij_1_3_n2, pool_pool_pe_b_peij_1_3_n1,
         pool_pool_pe_b_peij_1_3_q_k, pool_pool_pe_b_peij_1_3_gck,
         pool_pool_pe_b_peij_1_3_add_c_out,
         pool_pool_pe_b_peij_1_3_add_fai_0_n5,
         pool_pool_pe_b_peij_1_3_add_fai_0_n4,
         pool_pool_pe_b_peij_1_3_add_fai_1_n5,
         pool_pool_pe_b_peij_1_3_add_fai_1_n4,
         pool_pool_pe_b_peij_1_3_add_fai_2_n5,
         pool_pool_pe_b_peij_1_3_add_fai_2_n4,
         pool_pool_pe_b_peij_1_3_add_fai_3_n5,
         pool_pool_pe_b_peij_1_3_add_fai_3_n4,
         pool_pool_pe_b_peij_1_3_add_fai_4_n5,
         pool_pool_pe_b_peij_1_3_add_fai_4_n4,
         pool_pool_pe_b_peij_1_3_add_fai_5_n5,
         pool_pool_pe_b_peij_1_3_add_fai_5_n4,
         pool_pool_pe_b_peij_1_3_add_fai_6_n5,
         pool_pool_pe_b_peij_1_3_add_fai_6_n4,
         pool_pool_pe_b_peij_1_3_add_fai_7_n5,
         pool_pool_pe_b_peij_1_3_add_fai_7_n4,
         pool_pool_pe_b_peij_1_3_add_fai_8_n5,
         pool_pool_pe_b_peij_1_3_add_fai_8_n4,
         pool_pool_pe_b_peij_1_3_add_fai_9_n5,
         pool_pool_pe_b_peij_1_3_add_fai_9_n4,
         pool_pool_pe_b_peij_1_3_add_fai_10_n5,
         pool_pool_pe_b_peij_1_3_add_fai_10_n4, pool_pool_pe_b_peij_2_0_n14,
         pool_pool_pe_b_peij_2_0_n12, pool_pool_pe_b_peij_2_0_n11,
         pool_pool_pe_b_peij_2_0_n10, pool_pool_pe_b_peij_2_0_n9,
         pool_pool_pe_b_peij_2_0_n8, pool_pool_pe_b_peij_2_0_n7,
         pool_pool_pe_b_peij_2_0_n6, pool_pool_pe_b_peij_2_0_n5,
         pool_pool_pe_b_peij_2_0_n4, pool_pool_pe_b_peij_2_0_n3,
         pool_pool_pe_b_peij_2_0_n2, pool_pool_pe_b_peij_2_0_n1,
         pool_pool_pe_b_peij_2_0_q_k, pool_pool_pe_b_peij_2_0_gck,
         pool_pool_pe_b_peij_2_0_add_c_out,
         pool_pool_pe_b_peij_2_0_add_fai_0_n5,
         pool_pool_pe_b_peij_2_0_add_fai_0_n4,
         pool_pool_pe_b_peij_2_0_add_fai_1_n5,
         pool_pool_pe_b_peij_2_0_add_fai_1_n4,
         pool_pool_pe_b_peij_2_0_add_fai_2_n5,
         pool_pool_pe_b_peij_2_0_add_fai_2_n4,
         pool_pool_pe_b_peij_2_0_add_fai_3_n5,
         pool_pool_pe_b_peij_2_0_add_fai_3_n4,
         pool_pool_pe_b_peij_2_0_add_fai_4_n5,
         pool_pool_pe_b_peij_2_0_add_fai_4_n4,
         pool_pool_pe_b_peij_2_0_add_fai_5_n5,
         pool_pool_pe_b_peij_2_0_add_fai_5_n4,
         pool_pool_pe_b_peij_2_0_add_fai_6_n5,
         pool_pool_pe_b_peij_2_0_add_fai_6_n4,
         pool_pool_pe_b_peij_2_0_add_fai_7_n5,
         pool_pool_pe_b_peij_2_0_add_fai_7_n4,
         pool_pool_pe_b_peij_2_0_add_fai_8_n5,
         pool_pool_pe_b_peij_2_0_add_fai_8_n4,
         pool_pool_pe_b_peij_2_0_add_fai_9_n5,
         pool_pool_pe_b_peij_2_0_add_fai_9_n4,
         pool_pool_pe_b_peij_2_0_add_fai_10_n5,
         pool_pool_pe_b_peij_2_0_add_fai_10_n4, pool_pool_pe_b_peij_2_1_n14,
         pool_pool_pe_b_peij_2_1_n12, pool_pool_pe_b_peij_2_1_n11,
         pool_pool_pe_b_peij_2_1_n10, pool_pool_pe_b_peij_2_1_n9,
         pool_pool_pe_b_peij_2_1_n8, pool_pool_pe_b_peij_2_1_n7,
         pool_pool_pe_b_peij_2_1_n6, pool_pool_pe_b_peij_2_1_n5,
         pool_pool_pe_b_peij_2_1_n4, pool_pool_pe_b_peij_2_1_n3,
         pool_pool_pe_b_peij_2_1_n2, pool_pool_pe_b_peij_2_1_n1,
         pool_pool_pe_b_peij_2_1_q_k, pool_pool_pe_b_peij_2_1_gck,
         pool_pool_pe_b_peij_2_1_add_c_out,
         pool_pool_pe_b_peij_2_1_add_fai_0_n5,
         pool_pool_pe_b_peij_2_1_add_fai_0_n4,
         pool_pool_pe_b_peij_2_1_add_fai_1_n5,
         pool_pool_pe_b_peij_2_1_add_fai_1_n4,
         pool_pool_pe_b_peij_2_1_add_fai_2_n5,
         pool_pool_pe_b_peij_2_1_add_fai_2_n4,
         pool_pool_pe_b_peij_2_1_add_fai_3_n5,
         pool_pool_pe_b_peij_2_1_add_fai_3_n4,
         pool_pool_pe_b_peij_2_1_add_fai_4_n5,
         pool_pool_pe_b_peij_2_1_add_fai_4_n4,
         pool_pool_pe_b_peij_2_1_add_fai_5_n5,
         pool_pool_pe_b_peij_2_1_add_fai_5_n4,
         pool_pool_pe_b_peij_2_1_add_fai_6_n5,
         pool_pool_pe_b_peij_2_1_add_fai_6_n4,
         pool_pool_pe_b_peij_2_1_add_fai_7_n5,
         pool_pool_pe_b_peij_2_1_add_fai_7_n4,
         pool_pool_pe_b_peij_2_1_add_fai_8_n5,
         pool_pool_pe_b_peij_2_1_add_fai_8_n4,
         pool_pool_pe_b_peij_2_1_add_fai_9_n5,
         pool_pool_pe_b_peij_2_1_add_fai_9_n4,
         pool_pool_pe_b_peij_2_1_add_fai_10_n5,
         pool_pool_pe_b_peij_2_1_add_fai_10_n4, pool_pool_pe_b_peij_2_2_n14,
         pool_pool_pe_b_peij_2_2_n12, pool_pool_pe_b_peij_2_2_n11,
         pool_pool_pe_b_peij_2_2_n10, pool_pool_pe_b_peij_2_2_n9,
         pool_pool_pe_b_peij_2_2_n8, pool_pool_pe_b_peij_2_2_n7,
         pool_pool_pe_b_peij_2_2_n6, pool_pool_pe_b_peij_2_2_n5,
         pool_pool_pe_b_peij_2_2_n4, pool_pool_pe_b_peij_2_2_n3,
         pool_pool_pe_b_peij_2_2_n2, pool_pool_pe_b_peij_2_2_n1,
         pool_pool_pe_b_peij_2_2_q_k, pool_pool_pe_b_peij_2_2_gck,
         pool_pool_pe_b_peij_2_2_add_c_out,
         pool_pool_pe_b_peij_2_2_add_fai_0_n5,
         pool_pool_pe_b_peij_2_2_add_fai_0_n4,
         pool_pool_pe_b_peij_2_2_add_fai_1_n5,
         pool_pool_pe_b_peij_2_2_add_fai_1_n4,
         pool_pool_pe_b_peij_2_2_add_fai_2_n5,
         pool_pool_pe_b_peij_2_2_add_fai_2_n4,
         pool_pool_pe_b_peij_2_2_add_fai_3_n5,
         pool_pool_pe_b_peij_2_2_add_fai_3_n4,
         pool_pool_pe_b_peij_2_2_add_fai_4_n5,
         pool_pool_pe_b_peij_2_2_add_fai_4_n4,
         pool_pool_pe_b_peij_2_2_add_fai_5_n5,
         pool_pool_pe_b_peij_2_2_add_fai_5_n4,
         pool_pool_pe_b_peij_2_2_add_fai_6_n5,
         pool_pool_pe_b_peij_2_2_add_fai_6_n4,
         pool_pool_pe_b_peij_2_2_add_fai_7_n5,
         pool_pool_pe_b_peij_2_2_add_fai_7_n4,
         pool_pool_pe_b_peij_2_2_add_fai_8_n5,
         pool_pool_pe_b_peij_2_2_add_fai_8_n4,
         pool_pool_pe_b_peij_2_2_add_fai_9_n5,
         pool_pool_pe_b_peij_2_2_add_fai_9_n4,
         pool_pool_pe_b_peij_2_2_add_fai_10_n5,
         pool_pool_pe_b_peij_2_2_add_fai_10_n4, pool_pool_pe_b_peij_2_3_n14,
         pool_pool_pe_b_peij_2_3_n12, pool_pool_pe_b_peij_2_3_n11,
         pool_pool_pe_b_peij_2_3_n10, pool_pool_pe_b_peij_2_3_n9,
         pool_pool_pe_b_peij_2_3_n8, pool_pool_pe_b_peij_2_3_n7,
         pool_pool_pe_b_peij_2_3_n6, pool_pool_pe_b_peij_2_3_n5,
         pool_pool_pe_b_peij_2_3_n4, pool_pool_pe_b_peij_2_3_n3,
         pool_pool_pe_b_peij_2_3_n2, pool_pool_pe_b_peij_2_3_n1,
         pool_pool_pe_b_peij_2_3_q_k, pool_pool_pe_b_peij_2_3_gck,
         pool_pool_pe_b_peij_2_3_add_c_out,
         pool_pool_pe_b_peij_2_3_add_fai_0_n5,
         pool_pool_pe_b_peij_2_3_add_fai_0_n4,
         pool_pool_pe_b_peij_2_3_add_fai_1_n5,
         pool_pool_pe_b_peij_2_3_add_fai_1_n4,
         pool_pool_pe_b_peij_2_3_add_fai_2_n5,
         pool_pool_pe_b_peij_2_3_add_fai_2_n4,
         pool_pool_pe_b_peij_2_3_add_fai_3_n5,
         pool_pool_pe_b_peij_2_3_add_fai_3_n4,
         pool_pool_pe_b_peij_2_3_add_fai_4_n5,
         pool_pool_pe_b_peij_2_3_add_fai_4_n4,
         pool_pool_pe_b_peij_2_3_add_fai_5_n5,
         pool_pool_pe_b_peij_2_3_add_fai_5_n4,
         pool_pool_pe_b_peij_2_3_add_fai_6_n5,
         pool_pool_pe_b_peij_2_3_add_fai_6_n4,
         pool_pool_pe_b_peij_2_3_add_fai_7_n5,
         pool_pool_pe_b_peij_2_3_add_fai_7_n4,
         pool_pool_pe_b_peij_2_3_add_fai_8_n5,
         pool_pool_pe_b_peij_2_3_add_fai_8_n4,
         pool_pool_pe_b_peij_2_3_add_fai_9_n5,
         pool_pool_pe_b_peij_2_3_add_fai_9_n4,
         pool_pool_pe_b_peij_2_3_add_fai_10_n5,
         pool_pool_pe_b_peij_2_3_add_fai_10_n4, pool_pool_pe_b_peij_3_0_n14,
         pool_pool_pe_b_peij_3_0_n12, pool_pool_pe_b_peij_3_0_n11,
         pool_pool_pe_b_peij_3_0_n10, pool_pool_pe_b_peij_3_0_n9,
         pool_pool_pe_b_peij_3_0_n8, pool_pool_pe_b_peij_3_0_n7,
         pool_pool_pe_b_peij_3_0_n6, pool_pool_pe_b_peij_3_0_n5,
         pool_pool_pe_b_peij_3_0_n4, pool_pool_pe_b_peij_3_0_n3,
         pool_pool_pe_b_peij_3_0_n2, pool_pool_pe_b_peij_3_0_n1,
         pool_pool_pe_b_peij_3_0_q_k, pool_pool_pe_b_peij_3_0_gck,
         pool_pool_pe_b_peij_3_0_add_c_out,
         pool_pool_pe_b_peij_3_0_add_fai_0_n5,
         pool_pool_pe_b_peij_3_0_add_fai_0_n4,
         pool_pool_pe_b_peij_3_0_add_fai_1_n5,
         pool_pool_pe_b_peij_3_0_add_fai_1_n4,
         pool_pool_pe_b_peij_3_0_add_fai_2_n5,
         pool_pool_pe_b_peij_3_0_add_fai_2_n4,
         pool_pool_pe_b_peij_3_0_add_fai_3_n5,
         pool_pool_pe_b_peij_3_0_add_fai_3_n4,
         pool_pool_pe_b_peij_3_0_add_fai_4_n5,
         pool_pool_pe_b_peij_3_0_add_fai_4_n4,
         pool_pool_pe_b_peij_3_0_add_fai_5_n5,
         pool_pool_pe_b_peij_3_0_add_fai_5_n4,
         pool_pool_pe_b_peij_3_0_add_fai_6_n5,
         pool_pool_pe_b_peij_3_0_add_fai_6_n4,
         pool_pool_pe_b_peij_3_0_add_fai_7_n5,
         pool_pool_pe_b_peij_3_0_add_fai_7_n4,
         pool_pool_pe_b_peij_3_0_add_fai_8_n5,
         pool_pool_pe_b_peij_3_0_add_fai_8_n4,
         pool_pool_pe_b_peij_3_0_add_fai_9_n5,
         pool_pool_pe_b_peij_3_0_add_fai_9_n4,
         pool_pool_pe_b_peij_3_0_add_fai_10_n5,
         pool_pool_pe_b_peij_3_0_add_fai_10_n4, pool_pool_pe_b_peij_3_1_n14,
         pool_pool_pe_b_peij_3_1_n12, pool_pool_pe_b_peij_3_1_n11,
         pool_pool_pe_b_peij_3_1_n10, pool_pool_pe_b_peij_3_1_n9,
         pool_pool_pe_b_peij_3_1_n8, pool_pool_pe_b_peij_3_1_n7,
         pool_pool_pe_b_peij_3_1_n6, pool_pool_pe_b_peij_3_1_n5,
         pool_pool_pe_b_peij_3_1_n4, pool_pool_pe_b_peij_3_1_n3,
         pool_pool_pe_b_peij_3_1_n2, pool_pool_pe_b_peij_3_1_n1,
         pool_pool_pe_b_peij_3_1_q_k, pool_pool_pe_b_peij_3_1_gck,
         pool_pool_pe_b_peij_3_1_add_c_out,
         pool_pool_pe_b_peij_3_1_add_fai_0_n5,
         pool_pool_pe_b_peij_3_1_add_fai_0_n4,
         pool_pool_pe_b_peij_3_1_add_fai_1_n5,
         pool_pool_pe_b_peij_3_1_add_fai_1_n4,
         pool_pool_pe_b_peij_3_1_add_fai_2_n5,
         pool_pool_pe_b_peij_3_1_add_fai_2_n4,
         pool_pool_pe_b_peij_3_1_add_fai_3_n5,
         pool_pool_pe_b_peij_3_1_add_fai_3_n4,
         pool_pool_pe_b_peij_3_1_add_fai_4_n5,
         pool_pool_pe_b_peij_3_1_add_fai_4_n4,
         pool_pool_pe_b_peij_3_1_add_fai_5_n5,
         pool_pool_pe_b_peij_3_1_add_fai_5_n4,
         pool_pool_pe_b_peij_3_1_add_fai_6_n5,
         pool_pool_pe_b_peij_3_1_add_fai_6_n4,
         pool_pool_pe_b_peij_3_1_add_fai_7_n5,
         pool_pool_pe_b_peij_3_1_add_fai_7_n4,
         pool_pool_pe_b_peij_3_1_add_fai_8_n5,
         pool_pool_pe_b_peij_3_1_add_fai_8_n4,
         pool_pool_pe_b_peij_3_1_add_fai_9_n5,
         pool_pool_pe_b_peij_3_1_add_fai_9_n4,
         pool_pool_pe_b_peij_3_1_add_fai_10_n5,
         pool_pool_pe_b_peij_3_1_add_fai_10_n4, pool_pool_pe_b_peij_3_2_n14,
         pool_pool_pe_b_peij_3_2_n12, pool_pool_pe_b_peij_3_2_n11,
         pool_pool_pe_b_peij_3_2_n10, pool_pool_pe_b_peij_3_2_n9,
         pool_pool_pe_b_peij_3_2_n8, pool_pool_pe_b_peij_3_2_n7,
         pool_pool_pe_b_peij_3_2_n6, pool_pool_pe_b_peij_3_2_n5,
         pool_pool_pe_b_peij_3_2_n4, pool_pool_pe_b_peij_3_2_n3,
         pool_pool_pe_b_peij_3_2_n2, pool_pool_pe_b_peij_3_2_n1,
         pool_pool_pe_b_peij_3_2_q_k, pool_pool_pe_b_peij_3_2_gck,
         pool_pool_pe_b_peij_3_2_add_c_out,
         pool_pool_pe_b_peij_3_2_add_fai_0_n5,
         pool_pool_pe_b_peij_3_2_add_fai_0_n4,
         pool_pool_pe_b_peij_3_2_add_fai_1_n5,
         pool_pool_pe_b_peij_3_2_add_fai_1_n4,
         pool_pool_pe_b_peij_3_2_add_fai_2_n5,
         pool_pool_pe_b_peij_3_2_add_fai_2_n4,
         pool_pool_pe_b_peij_3_2_add_fai_3_n5,
         pool_pool_pe_b_peij_3_2_add_fai_3_n4,
         pool_pool_pe_b_peij_3_2_add_fai_4_n5,
         pool_pool_pe_b_peij_3_2_add_fai_4_n4,
         pool_pool_pe_b_peij_3_2_add_fai_5_n5,
         pool_pool_pe_b_peij_3_2_add_fai_5_n4,
         pool_pool_pe_b_peij_3_2_add_fai_6_n5,
         pool_pool_pe_b_peij_3_2_add_fai_6_n4,
         pool_pool_pe_b_peij_3_2_add_fai_7_n5,
         pool_pool_pe_b_peij_3_2_add_fai_7_n4,
         pool_pool_pe_b_peij_3_2_add_fai_8_n5,
         pool_pool_pe_b_peij_3_2_add_fai_8_n4,
         pool_pool_pe_b_peij_3_2_add_fai_9_n5,
         pool_pool_pe_b_peij_3_2_add_fai_9_n4,
         pool_pool_pe_b_peij_3_2_add_fai_10_n5,
         pool_pool_pe_b_peij_3_2_add_fai_10_n4, pool_pool_pe_b_peij_3_3_n14,
         pool_pool_pe_b_peij_3_3_n12, pool_pool_pe_b_peij_3_3_n11,
         pool_pool_pe_b_peij_3_3_n10, pool_pool_pe_b_peij_3_3_n9,
         pool_pool_pe_b_peij_3_3_n8, pool_pool_pe_b_peij_3_3_n7,
         pool_pool_pe_b_peij_3_3_n6, pool_pool_pe_b_peij_3_3_n5,
         pool_pool_pe_b_peij_3_3_n4, pool_pool_pe_b_peij_3_3_n3,
         pool_pool_pe_b_peij_3_3_n2, pool_pool_pe_b_peij_3_3_n1,
         pool_pool_pe_b_peij_3_3_q_k, pool_pool_pe_b_peij_3_3_gck,
         pool_pool_pe_b_peij_3_3_add_c_out,
         pool_pool_pe_b_peij_3_3_add_fai_0_n5,
         pool_pool_pe_b_peij_3_3_add_fai_0_n4,
         pool_pool_pe_b_peij_3_3_add_fai_1_n5,
         pool_pool_pe_b_peij_3_3_add_fai_1_n4,
         pool_pool_pe_b_peij_3_3_add_fai_2_n5,
         pool_pool_pe_b_peij_3_3_add_fai_2_n4,
         pool_pool_pe_b_peij_3_3_add_fai_3_n5,
         pool_pool_pe_b_peij_3_3_add_fai_3_n4,
         pool_pool_pe_b_peij_3_3_add_fai_4_n5,
         pool_pool_pe_b_peij_3_3_add_fai_4_n4,
         pool_pool_pe_b_peij_3_3_add_fai_5_n5,
         pool_pool_pe_b_peij_3_3_add_fai_5_n4,
         pool_pool_pe_b_peij_3_3_add_fai_6_n5,
         pool_pool_pe_b_peij_3_3_add_fai_6_n4,
         pool_pool_pe_b_peij_3_3_add_fai_7_n5,
         pool_pool_pe_b_peij_3_3_add_fai_7_n4,
         pool_pool_pe_b_peij_3_3_add_fai_8_n5,
         pool_pool_pe_b_peij_3_3_add_fai_8_n4,
         pool_pool_pe_b_peij_3_3_add_fai_9_n5,
         pool_pool_pe_b_peij_3_3_add_fai_9_n4,
         pool_pool_pe_b_peij_3_3_add_fai_10_n5,
         pool_pool_pe_b_peij_3_3_add_fai_10_n4, pool_pool_count_n12,
         pool_pool_count_n10, pool_pool_count_n9, pool_pool_count_n7,
         pool_pool_count_n4, pool_pool_count_n3, pool_pool_count_n2,
         pool_pool_count_n1, pool_pool_count_n18, pool_pool_count_n17,
         pool_pool_count_n15, pool_pool_count_n13, pool_pool_count_n11,
         pool_pool_count_n8, pool_pool_count_n6, pool_pool_count_n5,
         pool_pool_shift_row0_n4, pool_pool_shift_row0_n3,
         pool_pool_shift_row0_n2, pool_pool_shift_row0_n1,
         pool_pool_shift_row0_n12, pool_pool_shift_row0_n11,
         pool_pool_shift_row0_n10, pool_pool_shift_row0_n9,
         pool_pool_shift_row0_n8, pool_pool_shift_row0_n7,
         pool_pool_shift_row0_n6, pool_pool_shift_row0_n5,
         pool_pool_shift_row1_n20, pool_pool_shift_row1_n19,
         pool_pool_shift_row1_n18, pool_pool_shift_row1_n17,
         pool_pool_shift_row1_n16, pool_pool_shift_row1_n15,
         pool_pool_shift_row1_n14, pool_pool_shift_row1_n13,
         pool_pool_shift_row1_n4, pool_pool_shift_row1_n3,
         pool_pool_shift_row1_n2, pool_pool_shift_row1_n1,
         pool_pool_shift_row2_n20, pool_pool_shift_row2_n19,
         pool_pool_shift_row2_n18, pool_pool_shift_row2_n17,
         pool_pool_shift_row2_n16, pool_pool_shift_row2_n15,
         pool_pool_shift_row2_n14, pool_pool_shift_row2_n13,
         pool_pool_shift_row2_n4, pool_pool_shift_row2_n3,
         pool_pool_shift_row2_n2, pool_pool_shift_row2_n1,
         pool_pool_shift_row3_n20, pool_pool_shift_row3_n19,
         pool_pool_shift_row3_n18, pool_pool_shift_row3_n17,
         pool_pool_shift_row3_n16, pool_pool_shift_row3_n15,
         pool_pool_shift_row3_n14, pool_pool_shift_row3_n13,
         pool_pool_shift_row3_n4, pool_pool_shift_row3_n3,
         pool_pool_shift_row3_n2, pool_pool_shift_row3_n1, pool_fsm_n18,
         pool_fsm_n17, pool_fsm_n10, pool_fsm_n5, pool_fsm_n4, pool_fsm_n2,
         pool_fsm_n19, pool_fsm_n16, pool_fsm_n15, pool_fsm_n14, pool_fsm_n13,
         pool_fsm_n12, pool_fsm_n11, pool_fsm_n9, pool_fsm_n8, pool_fsm_n6,
         pool_fsm_net424, pool_fsm_N31, pool_fsm_N29, pool_fsm_N28,
         pool_fsm_N11, pool_fsm_current_state_0_, pool_fsm_current_state_1_,
         pool_fsm_current_state_2_, pool_gate_clk_n31, pool_gate_clk_n30,
         pool_gate_clk_n29, pool_gate_clk_n28, pool_gate_clk_n14,
         pool_gate_clk_n7, pool_gate_clk_n5, pool_gate_clk_n4,
         pool_gate_clk_n3, pool_gate_clk_n2, pool_gate_clk_n1,
         pool_gate_clk_n27, pool_gate_clk_n26, pool_gate_clk_n25,
         pool_gate_clk_n24, pool_gate_clk_n23, pool_gate_clk_n22,
         pool_gate_clk_n21, pool_gate_clk_n20, pool_gate_clk_n19,
         pool_gate_clk_n18, pool_gate_clk_n17, pool_gate_clk_n16,
         pool_gate_clk_n15, pool_gate_clk_n10, pool_gate_clk_n9,
         pool_gate_clk_n8, pool_gate_clk_n6, pool_gate_clk_del_tc_r_1,
         pool_gate_clk_N45, pool_gate_clk_del_tc_r, pool_gate_clk_cnt_r_out_0_,
         pool_gate_clk_cnt_r_out_1_, pool_gate_clk_tc_c,
         pool_gate_clk_cnt_c_out_0_, pool_gate_clk_cnt_c_out_1_,
         pool_gate_clk_del_1_tc, pool_gate_clk_del_0_tc, pool_gate_clk_N18,
         pool_gate_clk_N13, pool_gate_clk_dec_out_0_, pool_gate_clk_dec_out_1_,
         pool_gate_clk_dec_out_2_, pool_gate_clk_pool_size_1_,
         pool_gate_clk_pool_size_2_, pool_gate_clk_pool_size_3_,
         pool_gate_clk_pool_size_4_, pool_gate_clk_N0,
         pool_gate_clk_mux_pool_n6, pool_gate_clk_mux_pool_n11,
         pool_gate_clk_mux_pool_n10, pool_gate_clk_mux_pool_n9,
         pool_gate_clk_mux_pool_n8, pool_gate_clk_mux_pool_n7,
         pool_gate_clk_mux_cmask_n1, pool_gate_clk_mux_rmask_n1;
  wire   [3:0] pool_ckg_cmask;
  wire   [3:0] pool_ckg_rmask;
  wire   [175:0] pool_pool_pe_b_o_data;
  wire   [63:0] pool_pool_pe_b_i_data;
  wire   [15:0] pool_pool_pe_b_int_pe_en;
  wire   [10:0] pool_pool_pe_b_peij_0_0_d_acc;
  wire   [2:0] pool_pool_pe_b_peij_0_0_sgnext;
  wire   [10:0] pool_pool_pe_b_peij_0_0_add_notb;
  wire   [10:1] pool_pool_pe_b_peij_0_0_add_cprop;
  wire   [10:0] pool_pool_pe_b_peij_0_1_d_acc;
  wire   [2:0] pool_pool_pe_b_peij_0_1_sgnext;
  wire   [10:0] pool_pool_pe_b_peij_0_1_add_notb;
  wire   [10:1] pool_pool_pe_b_peij_0_1_add_cprop;
  wire   [10:0] pool_pool_pe_b_peij_0_2_d_acc;
  wire   [2:0] pool_pool_pe_b_peij_0_2_sgnext;
  wire   [10:0] pool_pool_pe_b_peij_0_2_add_notb;
  wire   [10:1] pool_pool_pe_b_peij_0_2_add_cprop;
  wire   [10:0] pool_pool_pe_b_peij_0_3_d_acc;
  wire   [2:0] pool_pool_pe_b_peij_0_3_sgnext;
  wire   [10:0] pool_pool_pe_b_peij_0_3_add_notb;
  wire   [10:1] pool_pool_pe_b_peij_0_3_add_cprop;
  wire   [10:0] pool_pool_pe_b_peij_1_0_d_acc;
  wire   [2:0] pool_pool_pe_b_peij_1_0_sgnext;
  wire   [10:0] pool_pool_pe_b_peij_1_0_add_notb;
  wire   [10:1] pool_pool_pe_b_peij_1_0_add_cprop;
  wire   [10:0] pool_pool_pe_b_peij_1_1_d_acc;
  wire   [2:0] pool_pool_pe_b_peij_1_1_sgnext;
  wire   [10:0] pool_pool_pe_b_peij_1_1_add_notb;
  wire   [10:1] pool_pool_pe_b_peij_1_1_add_cprop;
  wire   [10:0] pool_pool_pe_b_peij_1_2_d_acc;
  wire   [2:0] pool_pool_pe_b_peij_1_2_sgnext;
  wire   [10:0] pool_pool_pe_b_peij_1_2_add_notb;
  wire   [10:1] pool_pool_pe_b_peij_1_2_add_cprop;
  wire   [10:0] pool_pool_pe_b_peij_1_3_d_acc;
  wire   [2:0] pool_pool_pe_b_peij_1_3_sgnext;
  wire   [10:0] pool_pool_pe_b_peij_1_3_add_notb;
  wire   [10:1] pool_pool_pe_b_peij_1_3_add_cprop;
  wire   [10:0] pool_pool_pe_b_peij_2_0_d_acc;
  wire   [2:0] pool_pool_pe_b_peij_2_0_sgnext;
  wire   [10:0] pool_pool_pe_b_peij_2_0_add_notb;
  wire   [10:1] pool_pool_pe_b_peij_2_0_add_cprop;
  wire   [10:0] pool_pool_pe_b_peij_2_1_d_acc;
  wire   [2:0] pool_pool_pe_b_peij_2_1_sgnext;
  wire   [10:0] pool_pool_pe_b_peij_2_1_add_notb;
  wire   [10:1] pool_pool_pe_b_peij_2_1_add_cprop;
  wire   [10:0] pool_pool_pe_b_peij_2_2_d_acc;
  wire   [2:0] pool_pool_pe_b_peij_2_2_sgnext;
  wire   [10:0] pool_pool_pe_b_peij_2_2_add_notb;
  wire   [10:1] pool_pool_pe_b_peij_2_2_add_cprop;
  wire   [10:0] pool_pool_pe_b_peij_2_3_d_acc;
  wire   [2:0] pool_pool_pe_b_peij_2_3_sgnext;
  wire   [10:0] pool_pool_pe_b_peij_2_3_add_notb;
  wire   [10:1] pool_pool_pe_b_peij_2_3_add_cprop;
  wire   [10:0] pool_pool_pe_b_peij_3_0_d_acc;
  wire   [2:0] pool_pool_pe_b_peij_3_0_sgnext;
  wire   [10:0] pool_pool_pe_b_peij_3_0_add_notb;
  wire   [10:1] pool_pool_pe_b_peij_3_0_add_cprop;
  wire   [10:0] pool_pool_pe_b_peij_3_1_d_acc;
  wire   [2:0] pool_pool_pe_b_peij_3_1_sgnext;
  wire   [10:0] pool_pool_pe_b_peij_3_1_add_notb;
  wire   [10:1] pool_pool_pe_b_peij_3_1_add_cprop;
  wire   [10:0] pool_pool_pe_b_peij_3_2_d_acc;
  wire   [2:0] pool_pool_pe_b_peij_3_2_sgnext;
  wire   [10:0] pool_pool_pe_b_peij_3_2_add_notb;
  wire   [10:1] pool_pool_pe_b_peij_3_2_add_cprop;
  wire   [10:0] pool_pool_pe_b_peij_3_3_d_acc;
  wire   [2:0] pool_pool_pe_b_peij_3_3_sgnext;
  wire   [10:0] pool_pool_pe_b_peij_3_3_add_notb;
  wire   [10:1] pool_pool_pe_b_peij_3_3_add_cprop;
  wire   [1:0] pool_fsm_next_state;
  assign o_pool_1[15] = 1'b0;
  assign o_pool_1[11] = 1'b0;
  assign o_pool_1[7] = 1'b0;
  assign o_pool_1[3] = 1'b0;
  assign o_pool_4[15] = 1'b0;
  assign o_pool_4[11] = 1'b0;
  assign o_pool_4[7] = 1'b0;
  assign o_pool_4[3] = 1'b0;
  assign o_pool_3[15] = 1'b0;
  assign o_pool_3[11] = 1'b0;
  assign o_pool_3[7] = 1'b0;
  assign o_pool_3[3] = 1'b0;
  assign o_pool_2[15] = 1'b0;
  assign o_pool_2[11] = 1'b0;
  assign o_pool_2[7] = 1'b0;
  assign o_pool_2[3] = 1'b0;

  INV_X2 pool_pool_interface_mux_0_U41 ( .A(pool_pool_interface_mux_0_n33), 
        .ZN(pool_pool_pe_b_i_data[48]) );
  INV_X2 pool_pool_interface_mux_0_U40 ( .A(pool_pool_interface_mux_0_n32), 
        .ZN(pool_pool_pe_b_i_data[58]) );
  INV_X2 pool_pool_interface_mux_0_U39 ( .A(pool_pool_interface_mux_0_n31), 
        .ZN(pool_pool_pe_b_i_data[59]) );
  INV_X2 pool_pool_interface_mux_0_U38 ( .A(pool_pool_interface_mux_0_n30), 
        .ZN(pool_pool_pe_b_i_data[60]) );
  INV_X2 pool_pool_interface_mux_0_U37 ( .A(pool_pool_interface_mux_0_n29), 
        .ZN(pool_pool_pe_b_i_data[61]) );
  INV_X2 pool_pool_interface_mux_0_U36 ( .A(pool_pool_interface_mux_0_n28), 
        .ZN(pool_pool_pe_b_i_data[62]) );
  INV_X2 pool_pool_interface_mux_0_U35 ( .A(pool_pool_interface_mux_0_n27), 
        .ZN(pool_pool_pe_b_i_data[63]) );
  INV_X2 pool_pool_interface_mux_0_U34 ( .A(pool_pool_interface_mux_0_n26), 
        .ZN(pool_pool_pe_b_i_data[49]) );
  INV_X2 pool_pool_interface_mux_0_U33 ( .A(pool_pool_interface_mux_0_n25), 
        .ZN(pool_pool_pe_b_i_data[50]) );
  INV_X2 pool_pool_interface_mux_0_U32 ( .A(pool_pool_interface_mux_0_n24), 
        .ZN(pool_pool_pe_b_i_data[51]) );
  INV_X2 pool_pool_interface_mux_0_U31 ( .A(pool_pool_interface_mux_0_n23), 
        .ZN(pool_pool_pe_b_i_data[52]) );
  INV_X2 pool_pool_interface_mux_0_U30 ( .A(pool_pool_interface_mux_0_n22), 
        .ZN(pool_pool_pe_b_i_data[53]) );
  INV_X2 pool_pool_interface_mux_0_U29 ( .A(pool_pool_interface_mux_0_n21), 
        .ZN(pool_pool_pe_b_i_data[54]) );
  INV_X2 pool_pool_interface_mux_0_U28 ( .A(pool_pool_interface_mux_0_n20), 
        .ZN(pool_pool_pe_b_i_data[55]) );
  INV_X2 pool_pool_interface_mux_0_U27 ( .A(pool_pool_interface_mux_0_n19), 
        .ZN(pool_pool_pe_b_i_data[56]) );
  INV_X2 pool_pool_interface_mux_0_U26 ( .A(pool_pool_interface_mux_0_n18), 
        .ZN(pool_pool_pe_b_i_data[57]) );
  CLKBUF_X3 pool_pool_interface_mux_0_U25 ( .A(pool_pool_interface_mux_0_n2), 
        .Z(pool_pool_interface_mux_0_n9) );
  CLKBUF_X3 pool_pool_interface_mux_0_U24 ( .A(pool_pool_interface_mux_0_n2), 
        .Z(pool_pool_interface_mux_0_n8) );
  CLKBUF_X3 pool_pool_interface_mux_0_U23 ( .A(pool_pool_interface_mux_0_n1), 
        .Z(pool_pool_interface_mux_0_n7) );
  CLKBUF_X3 pool_pool_interface_mux_0_U22 ( .A(pool_pool_interface_mux_0_n1), 
        .Z(pool_pool_interface_mux_0_n6) );
  CLKBUF_X3 pool_pool_interface_mux_0_U21 ( .A(pool_pool_interface_mux_0_n1), 
        .Z(pool_pool_interface_mux_0_n5) );
  INV_X1 pool_pool_interface_mux_0_U20 ( .A(pool_pool_interface_mux_0_n9), 
        .ZN(pool_pool_interface_mux_0_n4) );
  CLKBUF_X3 pool_pool_interface_mux_0_U19 ( .A(pool_sel0), .Z(
        pool_pool_interface_mux_0_n2) );
  CLKBUF_X3 pool_pool_interface_mux_0_U18 ( .A(pool_sel0), .Z(
        pool_pool_interface_mux_0_n1) );
  INV_X4 pool_pool_interface_mux_0_U17 ( .A(pool_pool_interface_mux_0_n9), 
        .ZN(pool_pool_interface_mux_0_n3) );
  AOI22_X2 pool_pool_interface_mux_0_U16 ( .A1(d_0[0]), .A2(
        pool_pool_interface_mux_0_n3), .B1(d_4[0]), .B2(
        pool_pool_interface_mux_0_n8), .ZN(pool_pool_interface_mux_0_n33) );
  AOI22_X2 pool_pool_interface_mux_0_U15 ( .A1(d_0[10]), .A2(
        pool_pool_interface_mux_0_n3), .B1(d_4[10]), .B2(
        pool_pool_interface_mux_0_n8), .ZN(pool_pool_interface_mux_0_n32) );
  AOI22_X2 pool_pool_interface_mux_0_U14 ( .A1(d_0[11]), .A2(
        pool_pool_interface_mux_0_n3), .B1(d_4[11]), .B2(
        pool_pool_interface_mux_0_n8), .ZN(pool_pool_interface_mux_0_n31) );
  AOI22_X2 pool_pool_interface_mux_0_U13 ( .A1(d_0[12]), .A2(
        pool_pool_interface_mux_0_n3), .B1(d_4[12]), .B2(
        pool_pool_interface_mux_0_n7), .ZN(pool_pool_interface_mux_0_n30) );
  AOI22_X2 pool_pool_interface_mux_0_U12 ( .A1(d_0[13]), .A2(
        pool_pool_interface_mux_0_n3), .B1(d_4[13]), .B2(
        pool_pool_interface_mux_0_n7), .ZN(pool_pool_interface_mux_0_n29) );
  AOI22_X2 pool_pool_interface_mux_0_U11 ( .A1(d_0[14]), .A2(
        pool_pool_interface_mux_0_n3), .B1(d_4[14]), .B2(
        pool_pool_interface_mux_0_n7), .ZN(pool_pool_interface_mux_0_n28) );
  AOI22_X2 pool_pool_interface_mux_0_U10 ( .A1(d_0[15]), .A2(
        pool_pool_interface_mux_0_n3), .B1(d_4[15]), .B2(
        pool_pool_interface_mux_0_n6), .ZN(pool_pool_interface_mux_0_n27) );
  AOI22_X2 pool_pool_interface_mux_0_U9 ( .A1(d_0[1]), .A2(
        pool_pool_interface_mux_0_n3), .B1(d_4[1]), .B2(
        pool_pool_interface_mux_0_n6), .ZN(pool_pool_interface_mux_0_n26) );
  AOI22_X2 pool_pool_interface_mux_0_U8 ( .A1(d_0[2]), .A2(
        pool_pool_interface_mux_0_n3), .B1(d_4[2]), .B2(
        pool_pool_interface_mux_0_n6), .ZN(pool_pool_interface_mux_0_n25) );
  AOI22_X2 pool_pool_interface_mux_0_U7 ( .A1(d_0[3]), .A2(
        pool_pool_interface_mux_0_n3), .B1(d_4[3]), .B2(
        pool_pool_interface_mux_0_n6), .ZN(pool_pool_interface_mux_0_n24) );
  AOI22_X2 pool_pool_interface_mux_0_U6 ( .A1(d_0[4]), .A2(
        pool_pool_interface_mux_0_n3), .B1(d_4[4]), .B2(
        pool_pool_interface_mux_0_n5), .ZN(pool_pool_interface_mux_0_n23) );
  AOI22_X2 pool_pool_interface_mux_0_U5 ( .A1(d_0[5]), .A2(
        pool_pool_interface_mux_0_n3), .B1(d_4[5]), .B2(
        pool_pool_interface_mux_0_n7), .ZN(pool_pool_interface_mux_0_n22) );
  AOI22_X2 pool_pool_interface_mux_0_U4 ( .A1(d_0[6]), .A2(
        pool_pool_interface_mux_0_n4), .B1(d_4[6]), .B2(
        pool_pool_interface_mux_0_n5), .ZN(pool_pool_interface_mux_0_n21) );
  AOI22_X2 pool_pool_interface_mux_0_U3 ( .A1(d_0[7]), .A2(
        pool_pool_interface_mux_0_n4), .B1(d_4[7]), .B2(
        pool_pool_interface_mux_0_n5), .ZN(pool_pool_interface_mux_0_n20) );
  AOI22_X2 pool_pool_interface_mux_0_U2 ( .A1(d_0[8]), .A2(
        pool_pool_interface_mux_0_n4), .B1(d_4[8]), .B2(
        pool_pool_interface_mux_0_n5), .ZN(pool_pool_interface_mux_0_n19) );
  AOI22_X2 pool_pool_interface_mux_0_U1 ( .A1(d_0[9]), .A2(
        pool_pool_interface_mux_0_n4), .B1(pool_pool_interface_mux_0_n8), .B2(
        d_4[9]), .ZN(pool_pool_interface_mux_0_n18) );
  INV_X2 pool_pool_interface_mux_1_U41 ( .A(pool_pool_interface_mux_1_n42), 
        .ZN(pool_pool_pe_b_i_data[32]) );
  INV_X2 pool_pool_interface_mux_1_U40 ( .A(pool_pool_interface_mux_1_n43), 
        .ZN(pool_pool_pe_b_i_data[42]) );
  INV_X2 pool_pool_interface_mux_1_U39 ( .A(pool_pool_interface_mux_1_n44), 
        .ZN(pool_pool_pe_b_i_data[43]) );
  INV_X2 pool_pool_interface_mux_1_U38 ( .A(pool_pool_interface_mux_1_n45), 
        .ZN(pool_pool_pe_b_i_data[44]) );
  INV_X2 pool_pool_interface_mux_1_U37 ( .A(pool_pool_interface_mux_1_n46), 
        .ZN(pool_pool_pe_b_i_data[45]) );
  INV_X2 pool_pool_interface_mux_1_U36 ( .A(pool_pool_interface_mux_1_n47), 
        .ZN(pool_pool_pe_b_i_data[46]) );
  INV_X2 pool_pool_interface_mux_1_U35 ( .A(pool_pool_interface_mux_1_n48), 
        .ZN(pool_pool_pe_b_i_data[47]) );
  INV_X2 pool_pool_interface_mux_1_U34 ( .A(pool_pool_interface_mux_1_n49), 
        .ZN(pool_pool_pe_b_i_data[33]) );
  INV_X2 pool_pool_interface_mux_1_U33 ( .A(pool_pool_interface_mux_1_n50), 
        .ZN(pool_pool_pe_b_i_data[34]) );
  INV_X2 pool_pool_interface_mux_1_U32 ( .A(pool_pool_interface_mux_1_n51), 
        .ZN(pool_pool_pe_b_i_data[35]) );
  INV_X2 pool_pool_interface_mux_1_U31 ( .A(pool_pool_interface_mux_1_n52), 
        .ZN(pool_pool_pe_b_i_data[36]) );
  INV_X2 pool_pool_interface_mux_1_U30 ( .A(pool_pool_interface_mux_1_n53), 
        .ZN(pool_pool_pe_b_i_data[37]) );
  INV_X2 pool_pool_interface_mux_1_U29 ( .A(pool_pool_interface_mux_1_n54), 
        .ZN(pool_pool_pe_b_i_data[38]) );
  INV_X2 pool_pool_interface_mux_1_U28 ( .A(pool_pool_interface_mux_1_n55), 
        .ZN(pool_pool_pe_b_i_data[39]) );
  INV_X2 pool_pool_interface_mux_1_U27 ( .A(pool_pool_interface_mux_1_n56), 
        .ZN(pool_pool_pe_b_i_data[40]) );
  INV_X2 pool_pool_interface_mux_1_U26 ( .A(pool_pool_interface_mux_1_n57), 
        .ZN(pool_pool_pe_b_i_data[41]) );
  CLKBUF_X3 pool_pool_interface_mux_1_U25 ( .A(pool_pool_interface_mux_1_n2), 
        .Z(pool_pool_interface_mux_1_n9) );
  CLKBUF_X3 pool_pool_interface_mux_1_U24 ( .A(pool_pool_interface_mux_1_n2), 
        .Z(pool_pool_interface_mux_1_n8) );
  CLKBUF_X3 pool_pool_interface_mux_1_U23 ( .A(pool_pool_interface_mux_1_n1), 
        .Z(pool_pool_interface_mux_1_n7) );
  CLKBUF_X3 pool_pool_interface_mux_1_U22 ( .A(pool_pool_interface_mux_1_n1), 
        .Z(pool_pool_interface_mux_1_n6) );
  CLKBUF_X3 pool_pool_interface_mux_1_U21 ( .A(pool_pool_interface_mux_1_n1), 
        .Z(pool_pool_interface_mux_1_n5) );
  INV_X1 pool_pool_interface_mux_1_U20 ( .A(pool_pool_interface_mux_1_n9), 
        .ZN(pool_pool_interface_mux_1_n4) );
  CLKBUF_X3 pool_pool_interface_mux_1_U19 ( .A(pool_sel0), .Z(
        pool_pool_interface_mux_1_n2) );
  CLKBUF_X3 pool_pool_interface_mux_1_U18 ( .A(pool_sel0), .Z(
        pool_pool_interface_mux_1_n1) );
  INV_X4 pool_pool_interface_mux_1_U17 ( .A(pool_pool_interface_mux_1_n9), 
        .ZN(pool_pool_interface_mux_1_n3) );
  AOI22_X2 pool_pool_interface_mux_1_U16 ( .A1(d_1[0]), .A2(
        pool_pool_interface_mux_1_n3), .B1(d_5[0]), .B2(
        pool_pool_interface_mux_1_n8), .ZN(pool_pool_interface_mux_1_n42) );
  AOI22_X2 pool_pool_interface_mux_1_U15 ( .A1(d_1[10]), .A2(
        pool_pool_interface_mux_1_n3), .B1(d_5[10]), .B2(
        pool_pool_interface_mux_1_n8), .ZN(pool_pool_interface_mux_1_n43) );
  AOI22_X2 pool_pool_interface_mux_1_U14 ( .A1(d_1[11]), .A2(
        pool_pool_interface_mux_1_n3), .B1(d_5[11]), .B2(
        pool_pool_interface_mux_1_n8), .ZN(pool_pool_interface_mux_1_n44) );
  AOI22_X2 pool_pool_interface_mux_1_U13 ( .A1(d_1[12]), .A2(
        pool_pool_interface_mux_1_n3), .B1(d_5[12]), .B2(
        pool_pool_interface_mux_1_n7), .ZN(pool_pool_interface_mux_1_n45) );
  AOI22_X2 pool_pool_interface_mux_1_U12 ( .A1(d_1[13]), .A2(
        pool_pool_interface_mux_1_n3), .B1(d_5[13]), .B2(
        pool_pool_interface_mux_1_n7), .ZN(pool_pool_interface_mux_1_n46) );
  AOI22_X2 pool_pool_interface_mux_1_U11 ( .A1(d_1[14]), .A2(
        pool_pool_interface_mux_1_n3), .B1(d_5[14]), .B2(
        pool_pool_interface_mux_1_n7), .ZN(pool_pool_interface_mux_1_n47) );
  AOI22_X2 pool_pool_interface_mux_1_U10 ( .A1(d_1[15]), .A2(
        pool_pool_interface_mux_1_n3), .B1(d_5[15]), .B2(
        pool_pool_interface_mux_1_n6), .ZN(pool_pool_interface_mux_1_n48) );
  AOI22_X2 pool_pool_interface_mux_1_U9 ( .A1(d_1[1]), .A2(
        pool_pool_interface_mux_1_n3), .B1(d_5[1]), .B2(
        pool_pool_interface_mux_1_n6), .ZN(pool_pool_interface_mux_1_n49) );
  AOI22_X2 pool_pool_interface_mux_1_U8 ( .A1(d_1[2]), .A2(
        pool_pool_interface_mux_1_n3), .B1(d_5[2]), .B2(
        pool_pool_interface_mux_1_n6), .ZN(pool_pool_interface_mux_1_n50) );
  AOI22_X2 pool_pool_interface_mux_1_U7 ( .A1(d_1[3]), .A2(
        pool_pool_interface_mux_1_n3), .B1(d_5[3]), .B2(
        pool_pool_interface_mux_1_n6), .ZN(pool_pool_interface_mux_1_n51) );
  AOI22_X2 pool_pool_interface_mux_1_U6 ( .A1(d_1[4]), .A2(
        pool_pool_interface_mux_1_n3), .B1(d_5[4]), .B2(
        pool_pool_interface_mux_1_n5), .ZN(pool_pool_interface_mux_1_n52) );
  AOI22_X2 pool_pool_interface_mux_1_U5 ( .A1(d_1[5]), .A2(
        pool_pool_interface_mux_1_n3), .B1(d_5[5]), .B2(
        pool_pool_interface_mux_1_n7), .ZN(pool_pool_interface_mux_1_n53) );
  AOI22_X2 pool_pool_interface_mux_1_U4 ( .A1(d_1[6]), .A2(
        pool_pool_interface_mux_1_n4), .B1(d_5[6]), .B2(
        pool_pool_interface_mux_1_n5), .ZN(pool_pool_interface_mux_1_n54) );
  AOI22_X2 pool_pool_interface_mux_1_U3 ( .A1(d_1[7]), .A2(
        pool_pool_interface_mux_1_n4), .B1(d_5[7]), .B2(
        pool_pool_interface_mux_1_n5), .ZN(pool_pool_interface_mux_1_n55) );
  AOI22_X2 pool_pool_interface_mux_1_U2 ( .A1(d_1[8]), .A2(
        pool_pool_interface_mux_1_n4), .B1(d_5[8]), .B2(
        pool_pool_interface_mux_1_n5), .ZN(pool_pool_interface_mux_1_n56) );
  AOI22_X2 pool_pool_interface_mux_1_U1 ( .A1(d_1[9]), .A2(
        pool_pool_interface_mux_1_n4), .B1(pool_pool_interface_mux_1_n8), .B2(
        d_5[9]), .ZN(pool_pool_interface_mux_1_n57) );
  INV_X2 pool_pool_interface_mux_2_U41 ( .A(pool_pool_interface_mux_2_n42), 
        .ZN(pool_pool_pe_b_i_data[16]) );
  INV_X2 pool_pool_interface_mux_2_U40 ( .A(pool_pool_interface_mux_2_n43), 
        .ZN(pool_pool_pe_b_i_data[26]) );
  INV_X2 pool_pool_interface_mux_2_U39 ( .A(pool_pool_interface_mux_2_n44), 
        .ZN(pool_pool_pe_b_i_data[27]) );
  INV_X2 pool_pool_interface_mux_2_U38 ( .A(pool_pool_interface_mux_2_n45), 
        .ZN(pool_pool_pe_b_i_data[28]) );
  INV_X2 pool_pool_interface_mux_2_U37 ( .A(pool_pool_interface_mux_2_n46), 
        .ZN(pool_pool_pe_b_i_data[29]) );
  INV_X2 pool_pool_interface_mux_2_U36 ( .A(pool_pool_interface_mux_2_n47), 
        .ZN(pool_pool_pe_b_i_data[30]) );
  INV_X2 pool_pool_interface_mux_2_U35 ( .A(pool_pool_interface_mux_2_n48), 
        .ZN(pool_pool_pe_b_i_data[31]) );
  INV_X2 pool_pool_interface_mux_2_U34 ( .A(pool_pool_interface_mux_2_n49), 
        .ZN(pool_pool_pe_b_i_data[17]) );
  INV_X2 pool_pool_interface_mux_2_U33 ( .A(pool_pool_interface_mux_2_n50), 
        .ZN(pool_pool_pe_b_i_data[18]) );
  INV_X2 pool_pool_interface_mux_2_U32 ( .A(pool_pool_interface_mux_2_n51), 
        .ZN(pool_pool_pe_b_i_data[19]) );
  INV_X2 pool_pool_interface_mux_2_U31 ( .A(pool_pool_interface_mux_2_n52), 
        .ZN(pool_pool_pe_b_i_data[20]) );
  INV_X2 pool_pool_interface_mux_2_U30 ( .A(pool_pool_interface_mux_2_n53), 
        .ZN(pool_pool_pe_b_i_data[21]) );
  INV_X2 pool_pool_interface_mux_2_U29 ( .A(pool_pool_interface_mux_2_n54), 
        .ZN(pool_pool_pe_b_i_data[22]) );
  INV_X2 pool_pool_interface_mux_2_U28 ( .A(pool_pool_interface_mux_2_n55), 
        .ZN(pool_pool_pe_b_i_data[23]) );
  INV_X2 pool_pool_interface_mux_2_U27 ( .A(pool_pool_interface_mux_2_n56), 
        .ZN(pool_pool_pe_b_i_data[24]) );
  INV_X2 pool_pool_interface_mux_2_U26 ( .A(pool_pool_interface_mux_2_n57), 
        .ZN(pool_pool_pe_b_i_data[25]) );
  CLKBUF_X3 pool_pool_interface_mux_2_U25 ( .A(pool_pool_interface_mux_2_n2), 
        .Z(pool_pool_interface_mux_2_n9) );
  CLKBUF_X3 pool_pool_interface_mux_2_U24 ( .A(pool_pool_interface_mux_2_n2), 
        .Z(pool_pool_interface_mux_2_n8) );
  CLKBUF_X3 pool_pool_interface_mux_2_U23 ( .A(pool_pool_interface_mux_2_n1), 
        .Z(pool_pool_interface_mux_2_n7) );
  CLKBUF_X3 pool_pool_interface_mux_2_U22 ( .A(pool_pool_interface_mux_2_n1), 
        .Z(pool_pool_interface_mux_2_n6) );
  CLKBUF_X3 pool_pool_interface_mux_2_U21 ( .A(pool_pool_interface_mux_2_n1), 
        .Z(pool_pool_interface_mux_2_n5) );
  INV_X1 pool_pool_interface_mux_2_U20 ( .A(pool_pool_interface_mux_2_n9), 
        .ZN(pool_pool_interface_mux_2_n4) );
  CLKBUF_X3 pool_pool_interface_mux_2_U19 ( .A(pool_sel0), .Z(
        pool_pool_interface_mux_2_n2) );
  CLKBUF_X3 pool_pool_interface_mux_2_U18 ( .A(pool_sel0), .Z(
        pool_pool_interface_mux_2_n1) );
  INV_X4 pool_pool_interface_mux_2_U17 ( .A(pool_pool_interface_mux_2_n9), 
        .ZN(pool_pool_interface_mux_2_n3) );
  AOI22_X2 pool_pool_interface_mux_2_U16 ( .A1(d_2[0]), .A2(
        pool_pool_interface_mux_2_n3), .B1(d_6[0]), .B2(
        pool_pool_interface_mux_2_n8), .ZN(pool_pool_interface_mux_2_n42) );
  AOI22_X2 pool_pool_interface_mux_2_U15 ( .A1(d_2[10]), .A2(
        pool_pool_interface_mux_2_n3), .B1(d_6[10]), .B2(
        pool_pool_interface_mux_2_n8), .ZN(pool_pool_interface_mux_2_n43) );
  AOI22_X2 pool_pool_interface_mux_2_U14 ( .A1(d_2[11]), .A2(
        pool_pool_interface_mux_2_n3), .B1(d_6[11]), .B2(
        pool_pool_interface_mux_2_n8), .ZN(pool_pool_interface_mux_2_n44) );
  AOI22_X2 pool_pool_interface_mux_2_U13 ( .A1(d_2[12]), .A2(
        pool_pool_interface_mux_2_n3), .B1(d_6[12]), .B2(
        pool_pool_interface_mux_2_n7), .ZN(pool_pool_interface_mux_2_n45) );
  AOI22_X2 pool_pool_interface_mux_2_U12 ( .A1(d_2[13]), .A2(
        pool_pool_interface_mux_2_n3), .B1(d_6[13]), .B2(
        pool_pool_interface_mux_2_n7), .ZN(pool_pool_interface_mux_2_n46) );
  AOI22_X2 pool_pool_interface_mux_2_U11 ( .A1(d_2[14]), .A2(
        pool_pool_interface_mux_2_n3), .B1(d_6[14]), .B2(
        pool_pool_interface_mux_2_n7), .ZN(pool_pool_interface_mux_2_n47) );
  AOI22_X2 pool_pool_interface_mux_2_U10 ( .A1(d_2[15]), .A2(
        pool_pool_interface_mux_2_n3), .B1(d_6[15]), .B2(
        pool_pool_interface_mux_2_n6), .ZN(pool_pool_interface_mux_2_n48) );
  AOI22_X2 pool_pool_interface_mux_2_U9 ( .A1(d_2[1]), .A2(
        pool_pool_interface_mux_2_n3), .B1(d_6[1]), .B2(
        pool_pool_interface_mux_2_n6), .ZN(pool_pool_interface_mux_2_n49) );
  AOI22_X2 pool_pool_interface_mux_2_U8 ( .A1(d_2[2]), .A2(
        pool_pool_interface_mux_2_n3), .B1(d_6[2]), .B2(
        pool_pool_interface_mux_2_n6), .ZN(pool_pool_interface_mux_2_n50) );
  AOI22_X2 pool_pool_interface_mux_2_U7 ( .A1(d_2[3]), .A2(
        pool_pool_interface_mux_2_n3), .B1(d_6[3]), .B2(
        pool_pool_interface_mux_2_n6), .ZN(pool_pool_interface_mux_2_n51) );
  AOI22_X2 pool_pool_interface_mux_2_U6 ( .A1(d_2[4]), .A2(
        pool_pool_interface_mux_2_n3), .B1(d_6[4]), .B2(
        pool_pool_interface_mux_2_n5), .ZN(pool_pool_interface_mux_2_n52) );
  AOI22_X2 pool_pool_interface_mux_2_U5 ( .A1(d_2[5]), .A2(
        pool_pool_interface_mux_2_n3), .B1(d_6[5]), .B2(
        pool_pool_interface_mux_2_n7), .ZN(pool_pool_interface_mux_2_n53) );
  AOI22_X2 pool_pool_interface_mux_2_U4 ( .A1(d_2[6]), .A2(
        pool_pool_interface_mux_2_n4), .B1(d_6[6]), .B2(
        pool_pool_interface_mux_2_n5), .ZN(pool_pool_interface_mux_2_n54) );
  AOI22_X2 pool_pool_interface_mux_2_U3 ( .A1(d_2[7]), .A2(
        pool_pool_interface_mux_2_n4), .B1(d_6[7]), .B2(
        pool_pool_interface_mux_2_n5), .ZN(pool_pool_interface_mux_2_n55) );
  AOI22_X2 pool_pool_interface_mux_2_U2 ( .A1(d_2[8]), .A2(
        pool_pool_interface_mux_2_n4), .B1(d_6[8]), .B2(
        pool_pool_interface_mux_2_n5), .ZN(pool_pool_interface_mux_2_n56) );
  AOI22_X2 pool_pool_interface_mux_2_U1 ( .A1(d_2[9]), .A2(
        pool_pool_interface_mux_2_n4), .B1(pool_pool_interface_mux_2_n8), .B2(
        d_6[9]), .ZN(pool_pool_interface_mux_2_n57) );
  INV_X2 pool_pool_interface_mux_3_U41 ( .A(pool_pool_interface_mux_3_n42), 
        .ZN(pool_pool_pe_b_i_data[0]) );
  INV_X2 pool_pool_interface_mux_3_U40 ( .A(pool_pool_interface_mux_3_n43), 
        .ZN(pool_pool_pe_b_i_data[10]) );
  INV_X2 pool_pool_interface_mux_3_U39 ( .A(pool_pool_interface_mux_3_n44), 
        .ZN(pool_pool_pe_b_i_data[11]) );
  INV_X2 pool_pool_interface_mux_3_U38 ( .A(pool_pool_interface_mux_3_n45), 
        .ZN(pool_pool_pe_b_i_data[12]) );
  INV_X2 pool_pool_interface_mux_3_U37 ( .A(pool_pool_interface_mux_3_n46), 
        .ZN(pool_pool_pe_b_i_data[13]) );
  INV_X2 pool_pool_interface_mux_3_U36 ( .A(pool_pool_interface_mux_3_n47), 
        .ZN(pool_pool_pe_b_i_data[14]) );
  INV_X2 pool_pool_interface_mux_3_U35 ( .A(pool_pool_interface_mux_3_n48), 
        .ZN(pool_pool_pe_b_i_data[15]) );
  INV_X2 pool_pool_interface_mux_3_U34 ( .A(pool_pool_interface_mux_3_n49), 
        .ZN(pool_pool_pe_b_i_data[1]) );
  INV_X2 pool_pool_interface_mux_3_U33 ( .A(pool_pool_interface_mux_3_n50), 
        .ZN(pool_pool_pe_b_i_data[2]) );
  INV_X2 pool_pool_interface_mux_3_U32 ( .A(pool_pool_interface_mux_3_n51), 
        .ZN(pool_pool_pe_b_i_data[3]) );
  INV_X2 pool_pool_interface_mux_3_U31 ( .A(pool_pool_interface_mux_3_n52), 
        .ZN(pool_pool_pe_b_i_data[4]) );
  INV_X2 pool_pool_interface_mux_3_U30 ( .A(pool_pool_interface_mux_3_n53), 
        .ZN(pool_pool_pe_b_i_data[5]) );
  INV_X2 pool_pool_interface_mux_3_U29 ( .A(pool_pool_interface_mux_3_n54), 
        .ZN(pool_pool_pe_b_i_data[6]) );
  INV_X2 pool_pool_interface_mux_3_U28 ( .A(pool_pool_interface_mux_3_n55), 
        .ZN(pool_pool_pe_b_i_data[7]) );
  INV_X2 pool_pool_interface_mux_3_U27 ( .A(pool_pool_interface_mux_3_n56), 
        .ZN(pool_pool_pe_b_i_data[8]) );
  INV_X2 pool_pool_interface_mux_3_U26 ( .A(pool_pool_interface_mux_3_n57), 
        .ZN(pool_pool_pe_b_i_data[9]) );
  CLKBUF_X3 pool_pool_interface_mux_3_U25 ( .A(pool_pool_interface_mux_3_n2), 
        .Z(pool_pool_interface_mux_3_n9) );
  CLKBUF_X3 pool_pool_interface_mux_3_U24 ( .A(pool_pool_interface_mux_3_n2), 
        .Z(pool_pool_interface_mux_3_n8) );
  CLKBUF_X3 pool_pool_interface_mux_3_U23 ( .A(pool_pool_interface_mux_3_n1), 
        .Z(pool_pool_interface_mux_3_n7) );
  CLKBUF_X3 pool_pool_interface_mux_3_U22 ( .A(pool_pool_interface_mux_3_n1), 
        .Z(pool_pool_interface_mux_3_n6) );
  CLKBUF_X3 pool_pool_interface_mux_3_U21 ( .A(pool_pool_interface_mux_3_n1), 
        .Z(pool_pool_interface_mux_3_n5) );
  INV_X1 pool_pool_interface_mux_3_U20 ( .A(pool_pool_interface_mux_3_n9), 
        .ZN(pool_pool_interface_mux_3_n4) );
  CLKBUF_X3 pool_pool_interface_mux_3_U19 ( .A(pool_sel0), .Z(
        pool_pool_interface_mux_3_n2) );
  CLKBUF_X3 pool_pool_interface_mux_3_U18 ( .A(pool_sel0), .Z(
        pool_pool_interface_mux_3_n1) );
  INV_X4 pool_pool_interface_mux_3_U17 ( .A(pool_pool_interface_mux_3_n9), 
        .ZN(pool_pool_interface_mux_3_n3) );
  AOI22_X2 pool_pool_interface_mux_3_U16 ( .A1(d_3[0]), .A2(
        pool_pool_interface_mux_3_n3), .B1(d_7[0]), .B2(
        pool_pool_interface_mux_3_n8), .ZN(pool_pool_interface_mux_3_n42) );
  AOI22_X2 pool_pool_interface_mux_3_U15 ( .A1(d_3[10]), .A2(
        pool_pool_interface_mux_3_n3), .B1(d_7[10]), .B2(
        pool_pool_interface_mux_3_n8), .ZN(pool_pool_interface_mux_3_n43) );
  AOI22_X2 pool_pool_interface_mux_3_U14 ( .A1(d_3[11]), .A2(
        pool_pool_interface_mux_3_n3), .B1(d_7[11]), .B2(
        pool_pool_interface_mux_3_n8), .ZN(pool_pool_interface_mux_3_n44) );
  AOI22_X2 pool_pool_interface_mux_3_U13 ( .A1(d_3[12]), .A2(
        pool_pool_interface_mux_3_n3), .B1(d_7[12]), .B2(
        pool_pool_interface_mux_3_n7), .ZN(pool_pool_interface_mux_3_n45) );
  AOI22_X2 pool_pool_interface_mux_3_U12 ( .A1(d_3[13]), .A2(
        pool_pool_interface_mux_3_n3), .B1(d_7[13]), .B2(
        pool_pool_interface_mux_3_n7), .ZN(pool_pool_interface_mux_3_n46) );
  AOI22_X2 pool_pool_interface_mux_3_U11 ( .A1(d_3[14]), .A2(
        pool_pool_interface_mux_3_n3), .B1(d_7[14]), .B2(
        pool_pool_interface_mux_3_n7), .ZN(pool_pool_interface_mux_3_n47) );
  AOI22_X2 pool_pool_interface_mux_3_U10 ( .A1(d_3[15]), .A2(
        pool_pool_interface_mux_3_n3), .B1(d_7[15]), .B2(
        pool_pool_interface_mux_3_n6), .ZN(pool_pool_interface_mux_3_n48) );
  AOI22_X2 pool_pool_interface_mux_3_U9 ( .A1(d_3[1]), .A2(
        pool_pool_interface_mux_3_n3), .B1(d_7[1]), .B2(
        pool_pool_interface_mux_3_n6), .ZN(pool_pool_interface_mux_3_n49) );
  AOI22_X2 pool_pool_interface_mux_3_U8 ( .A1(d_3[2]), .A2(
        pool_pool_interface_mux_3_n3), .B1(d_7[2]), .B2(
        pool_pool_interface_mux_3_n6), .ZN(pool_pool_interface_mux_3_n50) );
  AOI22_X2 pool_pool_interface_mux_3_U7 ( .A1(d_3[3]), .A2(
        pool_pool_interface_mux_3_n3), .B1(d_7[3]), .B2(
        pool_pool_interface_mux_3_n6), .ZN(pool_pool_interface_mux_3_n51) );
  AOI22_X2 pool_pool_interface_mux_3_U6 ( .A1(d_3[4]), .A2(
        pool_pool_interface_mux_3_n3), .B1(d_7[4]), .B2(
        pool_pool_interface_mux_3_n5), .ZN(pool_pool_interface_mux_3_n52) );
  AOI22_X2 pool_pool_interface_mux_3_U5 ( .A1(d_3[5]), .A2(
        pool_pool_interface_mux_3_n3), .B1(d_7[5]), .B2(
        pool_pool_interface_mux_3_n7), .ZN(pool_pool_interface_mux_3_n53) );
  AOI22_X2 pool_pool_interface_mux_3_U4 ( .A1(d_3[6]), .A2(
        pool_pool_interface_mux_3_n4), .B1(d_7[6]), .B2(
        pool_pool_interface_mux_3_n5), .ZN(pool_pool_interface_mux_3_n54) );
  AOI22_X2 pool_pool_interface_mux_3_U3 ( .A1(d_3[7]), .A2(
        pool_pool_interface_mux_3_n4), .B1(d_7[7]), .B2(
        pool_pool_interface_mux_3_n5), .ZN(pool_pool_interface_mux_3_n55) );
  AOI22_X2 pool_pool_interface_mux_3_U2 ( .A1(d_3[8]), .A2(
        pool_pool_interface_mux_3_n4), .B1(d_7[8]), .B2(
        pool_pool_interface_mux_3_n5), .ZN(pool_pool_interface_mux_3_n56) );
  AOI22_X2 pool_pool_interface_mux_3_U1 ( .A1(d_3[9]), .A2(
        pool_pool_interface_mux_3_n4), .B1(pool_pool_interface_mux_3_n8), .B2(
        d_7[9]), .ZN(pool_pool_interface_mux_3_n57) );
  INV_X2 pool_pool_pe_b_U23 ( .A(en), .ZN(pool_pool_pe_b_n7) );
  CLKBUF_X3 pool_pool_pe_b_U22 ( .A(pool_ld_h), .Z(pool_pool_pe_b_n6) );
  CLKBUF_X3 pool_pool_pe_b_U21 ( .A(pool_ld_h), .Z(pool_pool_pe_b_n1) );
  OR2_X2 pool_pool_pe_b_U20 ( .A1(pool_ckg_rmask[3]), .A2(pool_pool_pe_b_n7), 
        .ZN(pool_pool_pe_b_n5) );
  NOR2_X2 pool_pool_pe_b_U19 ( .A1(pool_ckg_cmask[3]), .A2(pool_pool_pe_b_n5), 
        .ZN(pool_pool_pe_b_int_pe_en[15]) );
  NOR2_X2 pool_pool_pe_b_U18 ( .A1(pool_ckg_cmask[2]), .A2(pool_pool_pe_b_n5), 
        .ZN(pool_pool_pe_b_int_pe_en[14]) );
  NOR2_X2 pool_pool_pe_b_U17 ( .A1(pool_ckg_cmask[1]), .A2(pool_pool_pe_b_n5), 
        .ZN(pool_pool_pe_b_int_pe_en[13]) );
  NOR2_X2 pool_pool_pe_b_U16 ( .A1(pool_ckg_cmask[0]), .A2(pool_pool_pe_b_n5), 
        .ZN(pool_pool_pe_b_int_pe_en[12]) );
  OR2_X2 pool_pool_pe_b_U15 ( .A1(pool_ckg_rmask[2]), .A2(pool_pool_pe_b_n7), 
        .ZN(pool_pool_pe_b_n4) );
  NOR2_X2 pool_pool_pe_b_U14 ( .A1(pool_ckg_cmask[3]), .A2(pool_pool_pe_b_n4), 
        .ZN(pool_pool_pe_b_int_pe_en[11]) );
  NOR2_X2 pool_pool_pe_b_U13 ( .A1(pool_ckg_cmask[2]), .A2(pool_pool_pe_b_n4), 
        .ZN(pool_pool_pe_b_int_pe_en[10]) );
  NOR2_X2 pool_pool_pe_b_U12 ( .A1(pool_ckg_cmask[1]), .A2(pool_pool_pe_b_n4), 
        .ZN(pool_pool_pe_b_int_pe_en[9]) );
  NOR2_X2 pool_pool_pe_b_U11 ( .A1(pool_ckg_cmask[0]), .A2(pool_pool_pe_b_n4), 
        .ZN(pool_pool_pe_b_int_pe_en[8]) );
  OR2_X2 pool_pool_pe_b_U10 ( .A1(pool_ckg_rmask[1]), .A2(pool_pool_pe_b_n7), 
        .ZN(pool_pool_pe_b_n3) );
  NOR2_X2 pool_pool_pe_b_U9 ( .A1(pool_ckg_cmask[3]), .A2(pool_pool_pe_b_n3), 
        .ZN(pool_pool_pe_b_int_pe_en[7]) );
  NOR2_X2 pool_pool_pe_b_U8 ( .A1(pool_ckg_cmask[2]), .A2(pool_pool_pe_b_n3), 
        .ZN(pool_pool_pe_b_int_pe_en[6]) );
  NOR2_X2 pool_pool_pe_b_U7 ( .A1(pool_ckg_cmask[1]), .A2(pool_pool_pe_b_n3), 
        .ZN(pool_pool_pe_b_int_pe_en[5]) );
  NOR2_X2 pool_pool_pe_b_U6 ( .A1(pool_ckg_cmask[0]), .A2(pool_pool_pe_b_n3), 
        .ZN(pool_pool_pe_b_int_pe_en[4]) );
  OR2_X2 pool_pool_pe_b_U5 ( .A1(pool_ckg_rmask[0]), .A2(pool_pool_pe_b_n7), 
        .ZN(pool_pool_pe_b_n2) );
  NOR2_X2 pool_pool_pe_b_U4 ( .A1(pool_ckg_cmask[3]), .A2(pool_pool_pe_b_n2), 
        .ZN(pool_pool_pe_b_int_pe_en[3]) );
  NOR2_X2 pool_pool_pe_b_U3 ( .A1(pool_ckg_cmask[2]), .A2(pool_pool_pe_b_n2), 
        .ZN(pool_pool_pe_b_int_pe_en[2]) );
  NOR2_X2 pool_pool_pe_b_U2 ( .A1(pool_ckg_cmask[1]), .A2(pool_pool_pe_b_n2), 
        .ZN(pool_pool_pe_b_int_pe_en[1]) );
  NOR2_X2 pool_pool_pe_b_U1 ( .A1(pool_ckg_cmask[0]), .A2(pool_pool_pe_b_n2), 
        .ZN(pool_pool_pe_b_int_pe_en[0]) );
  INV_X2 pool_pool_pe_b_peij_0_0_U21 ( .A(pool_sync_clr), .ZN(
        pool_pool_pe_b_peij_0_0_n14) );
  INV_X1 pool_pool_pe_b_peij_0_0_U18 ( .A(pool_pool_pe_b_n1), .ZN(
        pool_pool_pe_b_peij_0_0_n12) );
  AND2_X1 pool_pool_pe_b_peij_0_0_U13 ( .A1(pool_pool_pe_b_peij_0_0_d_acc[0]), 
        .A2(pool_pool_pe_b_peij_0_0_n14), .ZN(pool_pool_pe_b_peij_0_0_n11) );
  AND2_X1 pool_pool_pe_b_peij_0_0_U12 ( .A1(pool_pool_pe_b_peij_0_0_d_acc[1]), 
        .A2(pool_pool_pe_b_peij_0_0_n14), .ZN(pool_pool_pe_b_peij_0_0_n10) );
  AND2_X1 pool_pool_pe_b_peij_0_0_U11 ( .A1(pool_pool_pe_b_peij_0_0_d_acc[2]), 
        .A2(pool_pool_pe_b_peij_0_0_n14), .ZN(pool_pool_pe_b_peij_0_0_n9) );
  AND2_X1 pool_pool_pe_b_peij_0_0_U10 ( .A1(pool_pool_pe_b_peij_0_0_d_acc[3]), 
        .A2(pool_pool_pe_b_peij_0_0_n14), .ZN(pool_pool_pe_b_peij_0_0_n8) );
  AND2_X1 pool_pool_pe_b_peij_0_0_U9 ( .A1(pool_pool_pe_b_peij_0_0_d_acc[4]), 
        .A2(pool_pool_pe_b_peij_0_0_n14), .ZN(pool_pool_pe_b_peij_0_0_n7) );
  AND2_X1 pool_pool_pe_b_peij_0_0_U8 ( .A1(pool_pool_pe_b_peij_0_0_d_acc[5]), 
        .A2(pool_pool_pe_b_peij_0_0_n14), .ZN(pool_pool_pe_b_peij_0_0_n6) );
  AND2_X1 pool_pool_pe_b_peij_0_0_U7 ( .A1(pool_pool_pe_b_peij_0_0_d_acc[6]), 
        .A2(pool_pool_pe_b_peij_0_0_n14), .ZN(pool_pool_pe_b_peij_0_0_n5) );
  AND2_X1 pool_pool_pe_b_peij_0_0_U6 ( .A1(pool_pool_pe_b_peij_0_0_d_acc[7]), 
        .A2(pool_pool_pe_b_peij_0_0_n14), .ZN(pool_pool_pe_b_peij_0_0_n4) );
  AND2_X1 pool_pool_pe_b_peij_0_0_U5 ( .A1(pool_pool_pe_b_peij_0_0_d_acc[8]), 
        .A2(pool_pool_pe_b_peij_0_0_n14), .ZN(pool_pool_pe_b_peij_0_0_n3) );
  AND2_X1 pool_pool_pe_b_peij_0_0_U4 ( .A1(pool_pool_pe_b_peij_0_0_d_acc[9]), 
        .A2(pool_pool_pe_b_peij_0_0_n14), .ZN(pool_pool_pe_b_peij_0_0_n2) );
  AND2_X1 pool_pool_pe_b_peij_0_0_U3 ( .A1(pool_pool_pe_b_peij_0_0_d_acc[10]), 
        .A2(pool_pool_pe_b_peij_0_0_n14), .ZN(pool_pool_pe_b_peij_0_0_n1) );
  DFFR_X1 pool_pool_pe_b_peij_0_0_q_acc_reg_10_ ( .D(
        pool_pool_pe_b_peij_0_0_n1), .CK(pool_pool_pe_b_peij_0_0_gck), .RN(
        pool_pool_pe_b_peij_0_0_n12), .Q(pool_pool_pe_b_o_data[175]) );
  DFFR_X1 pool_pool_pe_b_peij_0_0_q_acc_reg_9_ ( .D(pool_pool_pe_b_peij_0_0_n2), .CK(pool_pool_pe_b_peij_0_0_gck), .RN(pool_pool_pe_b_peij_0_0_n12), .Q(
        pool_pool_pe_b_o_data[174]) );
  DFFR_X1 pool_pool_pe_b_peij_0_0_q_acc_reg_8_ ( .D(pool_pool_pe_b_peij_0_0_n3), .CK(pool_pool_pe_b_peij_0_0_gck), .RN(pool_pool_pe_b_peij_0_0_n12), .Q(
        pool_pool_pe_b_o_data[173]) );
  DFFR_X1 pool_pool_pe_b_peij_0_0_q_acc_reg_7_ ( .D(pool_pool_pe_b_peij_0_0_n4), .CK(pool_pool_pe_b_peij_0_0_gck), .RN(pool_pool_pe_b_peij_0_0_n12), .Q(
        pool_pool_pe_b_o_data[172]) );
  DFFR_X1 pool_pool_pe_b_peij_0_0_q_acc_reg_6_ ( .D(pool_pool_pe_b_peij_0_0_n5), .CK(pool_pool_pe_b_peij_0_0_gck), .RN(pool_pool_pe_b_peij_0_0_n12), .Q(
        pool_pool_pe_b_o_data[171]) );
  DFFR_X1 pool_pool_pe_b_peij_0_0_q_acc_reg_5_ ( .D(pool_pool_pe_b_peij_0_0_n6), .CK(pool_pool_pe_b_peij_0_0_gck), .RN(pool_pool_pe_b_peij_0_0_n12), .Q(
        pool_pool_pe_b_o_data[170]) );
  DFFR_X1 pool_pool_pe_b_peij_0_0_q_acc_reg_4_ ( .D(pool_pool_pe_b_peij_0_0_n7), .CK(pool_pool_pe_b_peij_0_0_gck), .RN(pool_pool_pe_b_peij_0_0_n12), .Q(
        pool_pool_pe_b_o_data[169]) );
  DFFR_X1 pool_pool_pe_b_peij_0_0_q_acc_reg_3_ ( .D(pool_pool_pe_b_peij_0_0_n8), .CK(pool_pool_pe_b_peij_0_0_gck), .RN(pool_pool_pe_b_peij_0_0_n12), .Q(
        pool_pool_pe_b_o_data[168]) );
  DFFR_X1 pool_pool_pe_b_peij_0_0_q_acc_reg_2_ ( .D(pool_pool_pe_b_peij_0_0_n9), .CK(pool_pool_pe_b_peij_0_0_gck), .RN(pool_pool_pe_b_peij_0_0_n12), .Q(
        pool_pool_pe_b_o_data[167]) );
  DFFR_X1 pool_pool_pe_b_peij_0_0_q_acc_reg_1_ ( .D(
        pool_pool_pe_b_peij_0_0_n10), .CK(pool_pool_pe_b_peij_0_0_gck), .RN(
        pool_pool_pe_b_peij_0_0_n12), .Q(pool_pool_pe_b_o_data[166]) );
  DFFR_X1 pool_pool_pe_b_peij_0_0_q_acc_reg_0_ ( .D(
        pool_pool_pe_b_peij_0_0_n11), .CK(pool_pool_pe_b_peij_0_0_gck), .RN(
        pool_pool_pe_b_peij_0_0_n12), .Q(pool_pool_pe_b_o_data[165]) );
  AND3_X2 pool_pool_pe_b_peij_0_0_U20 ( .A1(pool_pool_pe_b_int_pe_en[15]), 
        .A2(clk), .A3(1'b1), .ZN(pool_pool_pe_b_peij_0_0_gck) );
  SDFFR_X1 pool_pool_pe_b_peij_0_0_q_k_reg ( .D(1'b0), .SI(
        pool_pool_pe_b_peij_0_0_n14), .SE(1'b0), .CK(
        pool_pool_pe_b_peij_0_0_gck), .RN(pool_pool_pe_b_peij_0_0_n12), .Q(
        pool_pool_pe_b_peij_0_0_q_k) );
  XOR2_X1 pool_pool_pe_b_peij_0_0_add_U11 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_0_q_k), .Z(pool_pool_pe_b_peij_0_0_add_notb[0])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_0_add_U10 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_0_q_k), .Z(pool_pool_pe_b_peij_0_0_add_notb[10])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_0_add_U9 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_0_q_k), .Z(pool_pool_pe_b_peij_0_0_add_notb[1])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_0_add_U8 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_0_q_k), .Z(pool_pool_pe_b_peij_0_0_add_notb[2])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_0_add_U7 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_0_q_k), .Z(pool_pool_pe_b_peij_0_0_add_notb[3])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_0_add_U6 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_0_q_k), .Z(pool_pool_pe_b_peij_0_0_add_notb[4])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_0_add_U5 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_0_q_k), .Z(pool_pool_pe_b_peij_0_0_add_notb[5])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_0_add_U4 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_0_q_k), .Z(pool_pool_pe_b_peij_0_0_add_notb[6])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_0_add_U3 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_0_q_k), .Z(pool_pool_pe_b_peij_0_0_add_notb[7])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_0_add_U2 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_0_q_k), .Z(pool_pool_pe_b_peij_0_0_add_notb[8])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_0_add_U1 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_0_q_k), .Z(pool_pool_pe_b_peij_0_0_add_notb[9])
         );
  INV_X2 pool_pool_pe_b_peij_0_0_add_fai_0_U2 ( .A(
        pool_pool_pe_b_peij_0_0_add_fai_0_n3), .ZN(
        pool_pool_pe_b_peij_0_0_add_cprop[1]) );
  XOR2_X1 pool_pool_pe_b_peij_0_0_add_fai_0_U4 ( .A(pool_pool_pe_b_o_data[165]), .B(pool_pool_pe_b_peij_0_0_add_notb[0]), .Z(
        pool_pool_pe_b_peij_0_0_add_fai_0_n2) );
  XOR2_X1 pool_pool_pe_b_peij_0_0_add_fai_0_U3 ( .A(
        pool_pool_pe_b_peij_0_0_q_k), .B(pool_pool_pe_b_peij_0_0_add_fai_0_n2), 
        .Z(pool_pool_pe_b_peij_0_0_d_acc[0]) );
  AOI22_X2 pool_pool_pe_b_peij_0_0_add_fai_0_U1 ( .A1(
        pool_pool_pe_b_peij_0_0_add_notb[0]), .A2(pool_pool_pe_b_o_data[165]), 
        .B1(pool_pool_pe_b_peij_0_0_add_fai_0_n2), .B2(
        pool_pool_pe_b_peij_0_0_q_k), .ZN(pool_pool_pe_b_peij_0_0_add_fai_0_n3) );
  INV_X2 pool_pool_pe_b_peij_0_0_add_fai_1_U2 ( .A(
        pool_pool_pe_b_peij_0_0_add_fai_1_n4), .ZN(
        pool_pool_pe_b_peij_0_0_add_cprop[2]) );
  XOR2_X1 pool_pool_pe_b_peij_0_0_add_fai_1_U4 ( .A(pool_pool_pe_b_o_data[166]), .B(pool_pool_pe_b_peij_0_0_add_notb[1]), .Z(
        pool_pool_pe_b_peij_0_0_add_fai_1_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_0_add_fai_1_U3 ( .A(
        pool_pool_pe_b_peij_0_0_add_cprop[1]), .B(
        pool_pool_pe_b_peij_0_0_add_fai_1_n5), .Z(
        pool_pool_pe_b_peij_0_0_d_acc[1]) );
  AOI22_X2 pool_pool_pe_b_peij_0_0_add_fai_1_U1 ( .A1(
        pool_pool_pe_b_peij_0_0_add_notb[1]), .A2(pool_pool_pe_b_o_data[166]), 
        .B1(pool_pool_pe_b_peij_0_0_add_fai_1_n5), .B2(
        pool_pool_pe_b_peij_0_0_add_cprop[1]), .ZN(
        pool_pool_pe_b_peij_0_0_add_fai_1_n4) );
  INV_X2 pool_pool_pe_b_peij_0_0_add_fai_2_U2 ( .A(
        pool_pool_pe_b_peij_0_0_add_fai_2_n4), .ZN(
        pool_pool_pe_b_peij_0_0_add_cprop[3]) );
  XOR2_X1 pool_pool_pe_b_peij_0_0_add_fai_2_U4 ( .A(pool_pool_pe_b_o_data[167]), .B(pool_pool_pe_b_peij_0_0_add_notb[2]), .Z(
        pool_pool_pe_b_peij_0_0_add_fai_2_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_0_add_fai_2_U3 ( .A(
        pool_pool_pe_b_peij_0_0_add_cprop[2]), .B(
        pool_pool_pe_b_peij_0_0_add_fai_2_n5), .Z(
        pool_pool_pe_b_peij_0_0_d_acc[2]) );
  AOI22_X2 pool_pool_pe_b_peij_0_0_add_fai_2_U1 ( .A1(
        pool_pool_pe_b_peij_0_0_add_notb[2]), .A2(pool_pool_pe_b_o_data[167]), 
        .B1(pool_pool_pe_b_peij_0_0_add_fai_2_n5), .B2(
        pool_pool_pe_b_peij_0_0_add_cprop[2]), .ZN(
        pool_pool_pe_b_peij_0_0_add_fai_2_n4) );
  INV_X2 pool_pool_pe_b_peij_0_0_add_fai_3_U2 ( .A(
        pool_pool_pe_b_peij_0_0_add_fai_3_n4), .ZN(
        pool_pool_pe_b_peij_0_0_add_cprop[4]) );
  XOR2_X1 pool_pool_pe_b_peij_0_0_add_fai_3_U4 ( .A(pool_pool_pe_b_o_data[168]), .B(pool_pool_pe_b_peij_0_0_add_notb[3]), .Z(
        pool_pool_pe_b_peij_0_0_add_fai_3_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_0_add_fai_3_U3 ( .A(
        pool_pool_pe_b_peij_0_0_add_cprop[3]), .B(
        pool_pool_pe_b_peij_0_0_add_fai_3_n5), .Z(
        pool_pool_pe_b_peij_0_0_d_acc[3]) );
  AOI22_X2 pool_pool_pe_b_peij_0_0_add_fai_3_U1 ( .A1(
        pool_pool_pe_b_peij_0_0_add_notb[3]), .A2(pool_pool_pe_b_o_data[168]), 
        .B1(pool_pool_pe_b_peij_0_0_add_fai_3_n5), .B2(
        pool_pool_pe_b_peij_0_0_add_cprop[3]), .ZN(
        pool_pool_pe_b_peij_0_0_add_fai_3_n4) );
  INV_X2 pool_pool_pe_b_peij_0_0_add_fai_4_U2 ( .A(
        pool_pool_pe_b_peij_0_0_add_fai_4_n4), .ZN(
        pool_pool_pe_b_peij_0_0_add_cprop[5]) );
  XOR2_X1 pool_pool_pe_b_peij_0_0_add_fai_4_U4 ( .A(pool_pool_pe_b_o_data[169]), .B(pool_pool_pe_b_peij_0_0_add_notb[4]), .Z(
        pool_pool_pe_b_peij_0_0_add_fai_4_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_0_add_fai_4_U3 ( .A(
        pool_pool_pe_b_peij_0_0_add_cprop[4]), .B(
        pool_pool_pe_b_peij_0_0_add_fai_4_n5), .Z(
        pool_pool_pe_b_peij_0_0_d_acc[4]) );
  AOI22_X2 pool_pool_pe_b_peij_0_0_add_fai_4_U1 ( .A1(
        pool_pool_pe_b_peij_0_0_add_notb[4]), .A2(pool_pool_pe_b_o_data[169]), 
        .B1(pool_pool_pe_b_peij_0_0_add_fai_4_n5), .B2(
        pool_pool_pe_b_peij_0_0_add_cprop[4]), .ZN(
        pool_pool_pe_b_peij_0_0_add_fai_4_n4) );
  INV_X2 pool_pool_pe_b_peij_0_0_add_fai_5_U2 ( .A(
        pool_pool_pe_b_peij_0_0_add_fai_5_n4), .ZN(
        pool_pool_pe_b_peij_0_0_add_cprop[6]) );
  XOR2_X1 pool_pool_pe_b_peij_0_0_add_fai_5_U4 ( .A(pool_pool_pe_b_o_data[170]), .B(pool_pool_pe_b_peij_0_0_add_notb[5]), .Z(
        pool_pool_pe_b_peij_0_0_add_fai_5_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_0_add_fai_5_U3 ( .A(
        pool_pool_pe_b_peij_0_0_add_cprop[5]), .B(
        pool_pool_pe_b_peij_0_0_add_fai_5_n5), .Z(
        pool_pool_pe_b_peij_0_0_d_acc[5]) );
  AOI22_X2 pool_pool_pe_b_peij_0_0_add_fai_5_U1 ( .A1(
        pool_pool_pe_b_peij_0_0_add_notb[5]), .A2(pool_pool_pe_b_o_data[170]), 
        .B1(pool_pool_pe_b_peij_0_0_add_fai_5_n5), .B2(
        pool_pool_pe_b_peij_0_0_add_cprop[5]), .ZN(
        pool_pool_pe_b_peij_0_0_add_fai_5_n4) );
  INV_X2 pool_pool_pe_b_peij_0_0_add_fai_6_U2 ( .A(
        pool_pool_pe_b_peij_0_0_add_fai_6_n4), .ZN(
        pool_pool_pe_b_peij_0_0_add_cprop[7]) );
  XOR2_X1 pool_pool_pe_b_peij_0_0_add_fai_6_U4 ( .A(pool_pool_pe_b_o_data[171]), .B(pool_pool_pe_b_peij_0_0_add_notb[6]), .Z(
        pool_pool_pe_b_peij_0_0_add_fai_6_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_0_add_fai_6_U3 ( .A(
        pool_pool_pe_b_peij_0_0_add_cprop[6]), .B(
        pool_pool_pe_b_peij_0_0_add_fai_6_n5), .Z(
        pool_pool_pe_b_peij_0_0_d_acc[6]) );
  AOI22_X2 pool_pool_pe_b_peij_0_0_add_fai_6_U1 ( .A1(
        pool_pool_pe_b_peij_0_0_add_notb[6]), .A2(pool_pool_pe_b_o_data[171]), 
        .B1(pool_pool_pe_b_peij_0_0_add_fai_6_n5), .B2(
        pool_pool_pe_b_peij_0_0_add_cprop[6]), .ZN(
        pool_pool_pe_b_peij_0_0_add_fai_6_n4) );
  INV_X2 pool_pool_pe_b_peij_0_0_add_fai_7_U2 ( .A(
        pool_pool_pe_b_peij_0_0_add_fai_7_n4), .ZN(
        pool_pool_pe_b_peij_0_0_add_cprop[8]) );
  XOR2_X1 pool_pool_pe_b_peij_0_0_add_fai_7_U4 ( .A(pool_pool_pe_b_o_data[172]), .B(pool_pool_pe_b_peij_0_0_add_notb[7]), .Z(
        pool_pool_pe_b_peij_0_0_add_fai_7_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_0_add_fai_7_U3 ( .A(
        pool_pool_pe_b_peij_0_0_add_cprop[7]), .B(
        pool_pool_pe_b_peij_0_0_add_fai_7_n5), .Z(
        pool_pool_pe_b_peij_0_0_d_acc[7]) );
  AOI22_X2 pool_pool_pe_b_peij_0_0_add_fai_7_U1 ( .A1(
        pool_pool_pe_b_peij_0_0_add_notb[7]), .A2(pool_pool_pe_b_o_data[172]), 
        .B1(pool_pool_pe_b_peij_0_0_add_fai_7_n5), .B2(
        pool_pool_pe_b_peij_0_0_add_cprop[7]), .ZN(
        pool_pool_pe_b_peij_0_0_add_fai_7_n4) );
  INV_X2 pool_pool_pe_b_peij_0_0_add_fai_8_U2 ( .A(
        pool_pool_pe_b_peij_0_0_add_fai_8_n4), .ZN(
        pool_pool_pe_b_peij_0_0_add_cprop[9]) );
  XOR2_X1 pool_pool_pe_b_peij_0_0_add_fai_8_U4 ( .A(pool_pool_pe_b_o_data[173]), .B(pool_pool_pe_b_peij_0_0_add_notb[8]), .Z(
        pool_pool_pe_b_peij_0_0_add_fai_8_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_0_add_fai_8_U3 ( .A(
        pool_pool_pe_b_peij_0_0_add_cprop[8]), .B(
        pool_pool_pe_b_peij_0_0_add_fai_8_n5), .Z(
        pool_pool_pe_b_peij_0_0_d_acc[8]) );
  AOI22_X2 pool_pool_pe_b_peij_0_0_add_fai_8_U1 ( .A1(
        pool_pool_pe_b_peij_0_0_add_notb[8]), .A2(pool_pool_pe_b_o_data[173]), 
        .B1(pool_pool_pe_b_peij_0_0_add_fai_8_n5), .B2(
        pool_pool_pe_b_peij_0_0_add_cprop[8]), .ZN(
        pool_pool_pe_b_peij_0_0_add_fai_8_n4) );
  INV_X2 pool_pool_pe_b_peij_0_0_add_fai_9_U2 ( .A(
        pool_pool_pe_b_peij_0_0_add_fai_9_n4), .ZN(
        pool_pool_pe_b_peij_0_0_add_cprop[10]) );
  XOR2_X1 pool_pool_pe_b_peij_0_0_add_fai_9_U4 ( .A(pool_pool_pe_b_o_data[174]), .B(pool_pool_pe_b_peij_0_0_add_notb[9]), .Z(
        pool_pool_pe_b_peij_0_0_add_fai_9_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_0_add_fai_9_U3 ( .A(
        pool_pool_pe_b_peij_0_0_add_cprop[9]), .B(
        pool_pool_pe_b_peij_0_0_add_fai_9_n5), .Z(
        pool_pool_pe_b_peij_0_0_d_acc[9]) );
  AOI22_X2 pool_pool_pe_b_peij_0_0_add_fai_9_U1 ( .A1(
        pool_pool_pe_b_peij_0_0_add_notb[9]), .A2(pool_pool_pe_b_o_data[174]), 
        .B1(pool_pool_pe_b_peij_0_0_add_fai_9_n5), .B2(
        pool_pool_pe_b_peij_0_0_add_cprop[9]), .ZN(
        pool_pool_pe_b_peij_0_0_add_fai_9_n4) );
  INV_X2 pool_pool_pe_b_peij_0_0_add_fai_10_U2 ( .A(
        pool_pool_pe_b_peij_0_0_add_fai_10_n4), .ZN(
        pool_pool_pe_b_peij_0_0_add_c_out) );
  XOR2_X1 pool_pool_pe_b_peij_0_0_add_fai_10_U4 ( .A(
        pool_pool_pe_b_o_data[175]), .B(pool_pool_pe_b_peij_0_0_add_notb[10]), 
        .Z(pool_pool_pe_b_peij_0_0_add_fai_10_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_0_add_fai_10_U3 ( .A(
        pool_pool_pe_b_peij_0_0_add_cprop[10]), .B(
        pool_pool_pe_b_peij_0_0_add_fai_10_n5), .Z(
        pool_pool_pe_b_peij_0_0_d_acc[10]) );
  AOI22_X2 pool_pool_pe_b_peij_0_0_add_fai_10_U1 ( .A1(
        pool_pool_pe_b_peij_0_0_add_notb[10]), .A2(pool_pool_pe_b_o_data[175]), 
        .B1(pool_pool_pe_b_peij_0_0_add_fai_10_n5), .B2(
        pool_pool_pe_b_peij_0_0_add_cprop[10]), .ZN(
        pool_pool_pe_b_peij_0_0_add_fai_10_n4) );
  INV_X2 pool_pool_pe_b_peij_0_1_U21 ( .A(pool_sync_clr), .ZN(
        pool_pool_pe_b_peij_0_1_n14) );
  INV_X1 pool_pool_pe_b_peij_0_1_U18 ( .A(pool_pool_pe_b_n6), .ZN(
        pool_pool_pe_b_peij_0_1_n12) );
  AND2_X1 pool_pool_pe_b_peij_0_1_U13 ( .A1(pool_pool_pe_b_peij_0_1_d_acc[0]), 
        .A2(pool_pool_pe_b_peij_0_1_n14), .ZN(pool_pool_pe_b_peij_0_1_n11) );
  AND2_X1 pool_pool_pe_b_peij_0_1_U12 ( .A1(pool_pool_pe_b_peij_0_1_d_acc[1]), 
        .A2(pool_pool_pe_b_peij_0_1_n14), .ZN(pool_pool_pe_b_peij_0_1_n10) );
  AND2_X1 pool_pool_pe_b_peij_0_1_U11 ( .A1(pool_pool_pe_b_peij_0_1_d_acc[2]), 
        .A2(pool_pool_pe_b_peij_0_1_n14), .ZN(pool_pool_pe_b_peij_0_1_n9) );
  AND2_X1 pool_pool_pe_b_peij_0_1_U10 ( .A1(pool_pool_pe_b_peij_0_1_d_acc[3]), 
        .A2(pool_pool_pe_b_peij_0_1_n14), .ZN(pool_pool_pe_b_peij_0_1_n8) );
  AND2_X1 pool_pool_pe_b_peij_0_1_U9 ( .A1(pool_pool_pe_b_peij_0_1_d_acc[4]), 
        .A2(pool_pool_pe_b_peij_0_1_n14), .ZN(pool_pool_pe_b_peij_0_1_n7) );
  AND2_X1 pool_pool_pe_b_peij_0_1_U8 ( .A1(pool_pool_pe_b_peij_0_1_d_acc[5]), 
        .A2(pool_pool_pe_b_peij_0_1_n14), .ZN(pool_pool_pe_b_peij_0_1_n6) );
  AND2_X1 pool_pool_pe_b_peij_0_1_U7 ( .A1(pool_pool_pe_b_peij_0_1_d_acc[6]), 
        .A2(pool_pool_pe_b_peij_0_1_n14), .ZN(pool_pool_pe_b_peij_0_1_n5) );
  AND2_X1 pool_pool_pe_b_peij_0_1_U6 ( .A1(pool_pool_pe_b_peij_0_1_d_acc[7]), 
        .A2(pool_pool_pe_b_peij_0_1_n14), .ZN(pool_pool_pe_b_peij_0_1_n4) );
  AND2_X1 pool_pool_pe_b_peij_0_1_U5 ( .A1(pool_pool_pe_b_peij_0_1_d_acc[8]), 
        .A2(pool_pool_pe_b_peij_0_1_n14), .ZN(pool_pool_pe_b_peij_0_1_n3) );
  AND2_X1 pool_pool_pe_b_peij_0_1_U4 ( .A1(pool_pool_pe_b_peij_0_1_d_acc[9]), 
        .A2(pool_pool_pe_b_peij_0_1_n14), .ZN(pool_pool_pe_b_peij_0_1_n2) );
  AND2_X1 pool_pool_pe_b_peij_0_1_U3 ( .A1(pool_pool_pe_b_peij_0_1_d_acc[10]), 
        .A2(pool_pool_pe_b_peij_0_1_n14), .ZN(pool_pool_pe_b_peij_0_1_n1) );
  DFFR_X1 pool_pool_pe_b_peij_0_1_q_acc_reg_10_ ( .D(
        pool_pool_pe_b_peij_0_1_n1), .CK(pool_pool_pe_b_peij_0_1_gck), .RN(
        pool_pool_pe_b_peij_0_1_n12), .Q(pool_pool_pe_b_o_data[164]) );
  DFFR_X1 pool_pool_pe_b_peij_0_1_q_acc_reg_9_ ( .D(pool_pool_pe_b_peij_0_1_n2), .CK(pool_pool_pe_b_peij_0_1_gck), .RN(pool_pool_pe_b_peij_0_1_n12), .Q(
        pool_pool_pe_b_o_data[163]) );
  DFFR_X1 pool_pool_pe_b_peij_0_1_q_acc_reg_8_ ( .D(pool_pool_pe_b_peij_0_1_n3), .CK(pool_pool_pe_b_peij_0_1_gck), .RN(pool_pool_pe_b_peij_0_1_n12), .Q(
        pool_pool_pe_b_o_data[162]) );
  DFFR_X1 pool_pool_pe_b_peij_0_1_q_acc_reg_7_ ( .D(pool_pool_pe_b_peij_0_1_n4), .CK(pool_pool_pe_b_peij_0_1_gck), .RN(pool_pool_pe_b_peij_0_1_n12), .Q(
        pool_pool_pe_b_o_data[161]) );
  DFFR_X1 pool_pool_pe_b_peij_0_1_q_acc_reg_6_ ( .D(pool_pool_pe_b_peij_0_1_n5), .CK(pool_pool_pe_b_peij_0_1_gck), .RN(pool_pool_pe_b_peij_0_1_n12), .Q(
        pool_pool_pe_b_o_data[160]) );
  DFFR_X1 pool_pool_pe_b_peij_0_1_q_acc_reg_5_ ( .D(pool_pool_pe_b_peij_0_1_n6), .CK(pool_pool_pe_b_peij_0_1_gck), .RN(pool_pool_pe_b_peij_0_1_n12), .Q(
        pool_pool_pe_b_o_data[159]) );
  DFFR_X1 pool_pool_pe_b_peij_0_1_q_acc_reg_4_ ( .D(pool_pool_pe_b_peij_0_1_n7), .CK(pool_pool_pe_b_peij_0_1_gck), .RN(pool_pool_pe_b_peij_0_1_n12), .Q(
        pool_pool_pe_b_o_data[158]) );
  DFFR_X1 pool_pool_pe_b_peij_0_1_q_acc_reg_3_ ( .D(pool_pool_pe_b_peij_0_1_n8), .CK(pool_pool_pe_b_peij_0_1_gck), .RN(pool_pool_pe_b_peij_0_1_n12), .Q(
        pool_pool_pe_b_o_data[157]) );
  DFFR_X1 pool_pool_pe_b_peij_0_1_q_acc_reg_2_ ( .D(pool_pool_pe_b_peij_0_1_n9), .CK(pool_pool_pe_b_peij_0_1_gck), .RN(pool_pool_pe_b_peij_0_1_n12), .Q(
        pool_pool_pe_b_o_data[156]) );
  DFFR_X1 pool_pool_pe_b_peij_0_1_q_acc_reg_1_ ( .D(
        pool_pool_pe_b_peij_0_1_n10), .CK(pool_pool_pe_b_peij_0_1_gck), .RN(
        pool_pool_pe_b_peij_0_1_n12), .Q(pool_pool_pe_b_o_data[155]) );
  DFFR_X1 pool_pool_pe_b_peij_0_1_q_acc_reg_0_ ( .D(
        pool_pool_pe_b_peij_0_1_n11), .CK(pool_pool_pe_b_peij_0_1_gck), .RN(
        pool_pool_pe_b_peij_0_1_n12), .Q(pool_pool_pe_b_o_data[154]) );
  AND3_X2 pool_pool_pe_b_peij_0_1_U20 ( .A1(pool_pool_pe_b_int_pe_en[14]), 
        .A2(clk), .A3(1'b1), .ZN(pool_pool_pe_b_peij_0_1_gck) );
  SDFFR_X1 pool_pool_pe_b_peij_0_1_q_k_reg ( .D(1'b0), .SI(
        pool_pool_pe_b_peij_0_1_n14), .SE(1'b0), .CK(
        pool_pool_pe_b_peij_0_1_gck), .RN(pool_pool_pe_b_peij_0_1_n12), .Q(
        pool_pool_pe_b_peij_0_1_q_k) );
  XOR2_X1 pool_pool_pe_b_peij_0_1_add_U11 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_1_q_k), .Z(pool_pool_pe_b_peij_0_1_add_notb[0])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_1_add_U10 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_1_q_k), .Z(pool_pool_pe_b_peij_0_1_add_notb[10])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_1_add_U9 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_1_q_k), .Z(pool_pool_pe_b_peij_0_1_add_notb[1])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_1_add_U8 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_1_q_k), .Z(pool_pool_pe_b_peij_0_1_add_notb[2])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_1_add_U7 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_1_q_k), .Z(pool_pool_pe_b_peij_0_1_add_notb[3])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_1_add_U6 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_1_q_k), .Z(pool_pool_pe_b_peij_0_1_add_notb[4])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_1_add_U5 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_1_q_k), .Z(pool_pool_pe_b_peij_0_1_add_notb[5])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_1_add_U4 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_1_q_k), .Z(pool_pool_pe_b_peij_0_1_add_notb[6])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_1_add_U3 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_1_q_k), .Z(pool_pool_pe_b_peij_0_1_add_notb[7])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_1_add_U2 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_1_q_k), .Z(pool_pool_pe_b_peij_0_1_add_notb[8])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_1_add_U1 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_1_q_k), .Z(pool_pool_pe_b_peij_0_1_add_notb[9])
         );
  INV_X2 pool_pool_pe_b_peij_0_1_add_fai_0_U2 ( .A(
        pool_pool_pe_b_peij_0_1_add_fai_0_n4), .ZN(
        pool_pool_pe_b_peij_0_1_add_cprop[1]) );
  XOR2_X1 pool_pool_pe_b_peij_0_1_add_fai_0_U4 ( .A(pool_pool_pe_b_o_data[154]), .B(pool_pool_pe_b_peij_0_1_add_notb[0]), .Z(
        pool_pool_pe_b_peij_0_1_add_fai_0_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_1_add_fai_0_U3 ( .A(
        pool_pool_pe_b_peij_0_1_q_k), .B(pool_pool_pe_b_peij_0_1_add_fai_0_n5), 
        .Z(pool_pool_pe_b_peij_0_1_d_acc[0]) );
  AOI22_X2 pool_pool_pe_b_peij_0_1_add_fai_0_U1 ( .A1(
        pool_pool_pe_b_peij_0_1_add_notb[0]), .A2(pool_pool_pe_b_o_data[154]), 
        .B1(pool_pool_pe_b_peij_0_1_add_fai_0_n5), .B2(
        pool_pool_pe_b_peij_0_1_q_k), .ZN(pool_pool_pe_b_peij_0_1_add_fai_0_n4) );
  INV_X2 pool_pool_pe_b_peij_0_1_add_fai_1_U2 ( .A(
        pool_pool_pe_b_peij_0_1_add_fai_1_n4), .ZN(
        pool_pool_pe_b_peij_0_1_add_cprop[2]) );
  XOR2_X1 pool_pool_pe_b_peij_0_1_add_fai_1_U4 ( .A(pool_pool_pe_b_o_data[155]), .B(pool_pool_pe_b_peij_0_1_add_notb[1]), .Z(
        pool_pool_pe_b_peij_0_1_add_fai_1_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_1_add_fai_1_U3 ( .A(
        pool_pool_pe_b_peij_0_1_add_cprop[1]), .B(
        pool_pool_pe_b_peij_0_1_add_fai_1_n5), .Z(
        pool_pool_pe_b_peij_0_1_d_acc[1]) );
  AOI22_X2 pool_pool_pe_b_peij_0_1_add_fai_1_U1 ( .A1(
        pool_pool_pe_b_peij_0_1_add_notb[1]), .A2(pool_pool_pe_b_o_data[155]), 
        .B1(pool_pool_pe_b_peij_0_1_add_fai_1_n5), .B2(
        pool_pool_pe_b_peij_0_1_add_cprop[1]), .ZN(
        pool_pool_pe_b_peij_0_1_add_fai_1_n4) );
  INV_X2 pool_pool_pe_b_peij_0_1_add_fai_2_U2 ( .A(
        pool_pool_pe_b_peij_0_1_add_fai_2_n4), .ZN(
        pool_pool_pe_b_peij_0_1_add_cprop[3]) );
  XOR2_X1 pool_pool_pe_b_peij_0_1_add_fai_2_U4 ( .A(pool_pool_pe_b_o_data[156]), .B(pool_pool_pe_b_peij_0_1_add_notb[2]), .Z(
        pool_pool_pe_b_peij_0_1_add_fai_2_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_1_add_fai_2_U3 ( .A(
        pool_pool_pe_b_peij_0_1_add_cprop[2]), .B(
        pool_pool_pe_b_peij_0_1_add_fai_2_n5), .Z(
        pool_pool_pe_b_peij_0_1_d_acc[2]) );
  AOI22_X2 pool_pool_pe_b_peij_0_1_add_fai_2_U1 ( .A1(
        pool_pool_pe_b_peij_0_1_add_notb[2]), .A2(pool_pool_pe_b_o_data[156]), 
        .B1(pool_pool_pe_b_peij_0_1_add_fai_2_n5), .B2(
        pool_pool_pe_b_peij_0_1_add_cprop[2]), .ZN(
        pool_pool_pe_b_peij_0_1_add_fai_2_n4) );
  INV_X2 pool_pool_pe_b_peij_0_1_add_fai_3_U2 ( .A(
        pool_pool_pe_b_peij_0_1_add_fai_3_n4), .ZN(
        pool_pool_pe_b_peij_0_1_add_cprop[4]) );
  XOR2_X1 pool_pool_pe_b_peij_0_1_add_fai_3_U4 ( .A(pool_pool_pe_b_o_data[157]), .B(pool_pool_pe_b_peij_0_1_add_notb[3]), .Z(
        pool_pool_pe_b_peij_0_1_add_fai_3_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_1_add_fai_3_U3 ( .A(
        pool_pool_pe_b_peij_0_1_add_cprop[3]), .B(
        pool_pool_pe_b_peij_0_1_add_fai_3_n5), .Z(
        pool_pool_pe_b_peij_0_1_d_acc[3]) );
  AOI22_X2 pool_pool_pe_b_peij_0_1_add_fai_3_U1 ( .A1(
        pool_pool_pe_b_peij_0_1_add_notb[3]), .A2(pool_pool_pe_b_o_data[157]), 
        .B1(pool_pool_pe_b_peij_0_1_add_fai_3_n5), .B2(
        pool_pool_pe_b_peij_0_1_add_cprop[3]), .ZN(
        pool_pool_pe_b_peij_0_1_add_fai_3_n4) );
  INV_X2 pool_pool_pe_b_peij_0_1_add_fai_4_U2 ( .A(
        pool_pool_pe_b_peij_0_1_add_fai_4_n4), .ZN(
        pool_pool_pe_b_peij_0_1_add_cprop[5]) );
  XOR2_X1 pool_pool_pe_b_peij_0_1_add_fai_4_U4 ( .A(pool_pool_pe_b_o_data[158]), .B(pool_pool_pe_b_peij_0_1_add_notb[4]), .Z(
        pool_pool_pe_b_peij_0_1_add_fai_4_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_1_add_fai_4_U3 ( .A(
        pool_pool_pe_b_peij_0_1_add_cprop[4]), .B(
        pool_pool_pe_b_peij_0_1_add_fai_4_n5), .Z(
        pool_pool_pe_b_peij_0_1_d_acc[4]) );
  AOI22_X2 pool_pool_pe_b_peij_0_1_add_fai_4_U1 ( .A1(
        pool_pool_pe_b_peij_0_1_add_notb[4]), .A2(pool_pool_pe_b_o_data[158]), 
        .B1(pool_pool_pe_b_peij_0_1_add_fai_4_n5), .B2(
        pool_pool_pe_b_peij_0_1_add_cprop[4]), .ZN(
        pool_pool_pe_b_peij_0_1_add_fai_4_n4) );
  INV_X2 pool_pool_pe_b_peij_0_1_add_fai_5_U2 ( .A(
        pool_pool_pe_b_peij_0_1_add_fai_5_n4), .ZN(
        pool_pool_pe_b_peij_0_1_add_cprop[6]) );
  XOR2_X1 pool_pool_pe_b_peij_0_1_add_fai_5_U4 ( .A(pool_pool_pe_b_o_data[159]), .B(pool_pool_pe_b_peij_0_1_add_notb[5]), .Z(
        pool_pool_pe_b_peij_0_1_add_fai_5_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_1_add_fai_5_U3 ( .A(
        pool_pool_pe_b_peij_0_1_add_cprop[5]), .B(
        pool_pool_pe_b_peij_0_1_add_fai_5_n5), .Z(
        pool_pool_pe_b_peij_0_1_d_acc[5]) );
  AOI22_X2 pool_pool_pe_b_peij_0_1_add_fai_5_U1 ( .A1(
        pool_pool_pe_b_peij_0_1_add_notb[5]), .A2(pool_pool_pe_b_o_data[159]), 
        .B1(pool_pool_pe_b_peij_0_1_add_fai_5_n5), .B2(
        pool_pool_pe_b_peij_0_1_add_cprop[5]), .ZN(
        pool_pool_pe_b_peij_0_1_add_fai_5_n4) );
  INV_X2 pool_pool_pe_b_peij_0_1_add_fai_6_U2 ( .A(
        pool_pool_pe_b_peij_0_1_add_fai_6_n4), .ZN(
        pool_pool_pe_b_peij_0_1_add_cprop[7]) );
  XOR2_X1 pool_pool_pe_b_peij_0_1_add_fai_6_U4 ( .A(pool_pool_pe_b_o_data[160]), .B(pool_pool_pe_b_peij_0_1_add_notb[6]), .Z(
        pool_pool_pe_b_peij_0_1_add_fai_6_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_1_add_fai_6_U3 ( .A(
        pool_pool_pe_b_peij_0_1_add_cprop[6]), .B(
        pool_pool_pe_b_peij_0_1_add_fai_6_n5), .Z(
        pool_pool_pe_b_peij_0_1_d_acc[6]) );
  AOI22_X2 pool_pool_pe_b_peij_0_1_add_fai_6_U1 ( .A1(
        pool_pool_pe_b_peij_0_1_add_notb[6]), .A2(pool_pool_pe_b_o_data[160]), 
        .B1(pool_pool_pe_b_peij_0_1_add_fai_6_n5), .B2(
        pool_pool_pe_b_peij_0_1_add_cprop[6]), .ZN(
        pool_pool_pe_b_peij_0_1_add_fai_6_n4) );
  INV_X2 pool_pool_pe_b_peij_0_1_add_fai_7_U2 ( .A(
        pool_pool_pe_b_peij_0_1_add_fai_7_n4), .ZN(
        pool_pool_pe_b_peij_0_1_add_cprop[8]) );
  XOR2_X1 pool_pool_pe_b_peij_0_1_add_fai_7_U4 ( .A(pool_pool_pe_b_o_data[161]), .B(pool_pool_pe_b_peij_0_1_add_notb[7]), .Z(
        pool_pool_pe_b_peij_0_1_add_fai_7_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_1_add_fai_7_U3 ( .A(
        pool_pool_pe_b_peij_0_1_add_cprop[7]), .B(
        pool_pool_pe_b_peij_0_1_add_fai_7_n5), .Z(
        pool_pool_pe_b_peij_0_1_d_acc[7]) );
  AOI22_X2 pool_pool_pe_b_peij_0_1_add_fai_7_U1 ( .A1(
        pool_pool_pe_b_peij_0_1_add_notb[7]), .A2(pool_pool_pe_b_o_data[161]), 
        .B1(pool_pool_pe_b_peij_0_1_add_fai_7_n5), .B2(
        pool_pool_pe_b_peij_0_1_add_cprop[7]), .ZN(
        pool_pool_pe_b_peij_0_1_add_fai_7_n4) );
  INV_X2 pool_pool_pe_b_peij_0_1_add_fai_8_U2 ( .A(
        pool_pool_pe_b_peij_0_1_add_fai_8_n4), .ZN(
        pool_pool_pe_b_peij_0_1_add_cprop[9]) );
  XOR2_X1 pool_pool_pe_b_peij_0_1_add_fai_8_U4 ( .A(pool_pool_pe_b_o_data[162]), .B(pool_pool_pe_b_peij_0_1_add_notb[8]), .Z(
        pool_pool_pe_b_peij_0_1_add_fai_8_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_1_add_fai_8_U3 ( .A(
        pool_pool_pe_b_peij_0_1_add_cprop[8]), .B(
        pool_pool_pe_b_peij_0_1_add_fai_8_n5), .Z(
        pool_pool_pe_b_peij_0_1_d_acc[8]) );
  AOI22_X2 pool_pool_pe_b_peij_0_1_add_fai_8_U1 ( .A1(
        pool_pool_pe_b_peij_0_1_add_notb[8]), .A2(pool_pool_pe_b_o_data[162]), 
        .B1(pool_pool_pe_b_peij_0_1_add_fai_8_n5), .B2(
        pool_pool_pe_b_peij_0_1_add_cprop[8]), .ZN(
        pool_pool_pe_b_peij_0_1_add_fai_8_n4) );
  INV_X2 pool_pool_pe_b_peij_0_1_add_fai_9_U2 ( .A(
        pool_pool_pe_b_peij_0_1_add_fai_9_n4), .ZN(
        pool_pool_pe_b_peij_0_1_add_cprop[10]) );
  XOR2_X1 pool_pool_pe_b_peij_0_1_add_fai_9_U4 ( .A(pool_pool_pe_b_o_data[163]), .B(pool_pool_pe_b_peij_0_1_add_notb[9]), .Z(
        pool_pool_pe_b_peij_0_1_add_fai_9_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_1_add_fai_9_U3 ( .A(
        pool_pool_pe_b_peij_0_1_add_cprop[9]), .B(
        pool_pool_pe_b_peij_0_1_add_fai_9_n5), .Z(
        pool_pool_pe_b_peij_0_1_d_acc[9]) );
  AOI22_X2 pool_pool_pe_b_peij_0_1_add_fai_9_U1 ( .A1(
        pool_pool_pe_b_peij_0_1_add_notb[9]), .A2(pool_pool_pe_b_o_data[163]), 
        .B1(pool_pool_pe_b_peij_0_1_add_fai_9_n5), .B2(
        pool_pool_pe_b_peij_0_1_add_cprop[9]), .ZN(
        pool_pool_pe_b_peij_0_1_add_fai_9_n4) );
  INV_X2 pool_pool_pe_b_peij_0_1_add_fai_10_U2 ( .A(
        pool_pool_pe_b_peij_0_1_add_fai_10_n4), .ZN(
        pool_pool_pe_b_peij_0_1_add_c_out) );
  XOR2_X1 pool_pool_pe_b_peij_0_1_add_fai_10_U4 ( .A(
        pool_pool_pe_b_o_data[164]), .B(pool_pool_pe_b_peij_0_1_add_notb[10]), 
        .Z(pool_pool_pe_b_peij_0_1_add_fai_10_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_1_add_fai_10_U3 ( .A(
        pool_pool_pe_b_peij_0_1_add_cprop[10]), .B(
        pool_pool_pe_b_peij_0_1_add_fai_10_n5), .Z(
        pool_pool_pe_b_peij_0_1_d_acc[10]) );
  AOI22_X2 pool_pool_pe_b_peij_0_1_add_fai_10_U1 ( .A1(
        pool_pool_pe_b_peij_0_1_add_notb[10]), .A2(pool_pool_pe_b_o_data[164]), 
        .B1(pool_pool_pe_b_peij_0_1_add_fai_10_n5), .B2(
        pool_pool_pe_b_peij_0_1_add_cprop[10]), .ZN(
        pool_pool_pe_b_peij_0_1_add_fai_10_n4) );
  INV_X2 pool_pool_pe_b_peij_0_2_U21 ( .A(pool_sync_clr), .ZN(
        pool_pool_pe_b_peij_0_2_n14) );
  INV_X1 pool_pool_pe_b_peij_0_2_U18 ( .A(pool_pool_pe_b_n6), .ZN(
        pool_pool_pe_b_peij_0_2_n12) );
  AND2_X1 pool_pool_pe_b_peij_0_2_U13 ( .A1(pool_pool_pe_b_peij_0_2_d_acc[0]), 
        .A2(pool_pool_pe_b_peij_0_2_n14), .ZN(pool_pool_pe_b_peij_0_2_n11) );
  AND2_X1 pool_pool_pe_b_peij_0_2_U12 ( .A1(pool_pool_pe_b_peij_0_2_d_acc[1]), 
        .A2(pool_pool_pe_b_peij_0_2_n14), .ZN(pool_pool_pe_b_peij_0_2_n10) );
  AND2_X1 pool_pool_pe_b_peij_0_2_U11 ( .A1(pool_pool_pe_b_peij_0_2_d_acc[2]), 
        .A2(pool_pool_pe_b_peij_0_2_n14), .ZN(pool_pool_pe_b_peij_0_2_n9) );
  AND2_X1 pool_pool_pe_b_peij_0_2_U10 ( .A1(pool_pool_pe_b_peij_0_2_d_acc[3]), 
        .A2(pool_pool_pe_b_peij_0_2_n14), .ZN(pool_pool_pe_b_peij_0_2_n8) );
  AND2_X1 pool_pool_pe_b_peij_0_2_U9 ( .A1(pool_pool_pe_b_peij_0_2_d_acc[4]), 
        .A2(pool_pool_pe_b_peij_0_2_n14), .ZN(pool_pool_pe_b_peij_0_2_n7) );
  AND2_X1 pool_pool_pe_b_peij_0_2_U8 ( .A1(pool_pool_pe_b_peij_0_2_d_acc[5]), 
        .A2(pool_pool_pe_b_peij_0_2_n14), .ZN(pool_pool_pe_b_peij_0_2_n6) );
  AND2_X1 pool_pool_pe_b_peij_0_2_U7 ( .A1(pool_pool_pe_b_peij_0_2_d_acc[6]), 
        .A2(pool_pool_pe_b_peij_0_2_n14), .ZN(pool_pool_pe_b_peij_0_2_n5) );
  AND2_X1 pool_pool_pe_b_peij_0_2_U6 ( .A1(pool_pool_pe_b_peij_0_2_d_acc[7]), 
        .A2(pool_pool_pe_b_peij_0_2_n14), .ZN(pool_pool_pe_b_peij_0_2_n4) );
  AND2_X1 pool_pool_pe_b_peij_0_2_U5 ( .A1(pool_pool_pe_b_peij_0_2_d_acc[8]), 
        .A2(pool_pool_pe_b_peij_0_2_n14), .ZN(pool_pool_pe_b_peij_0_2_n3) );
  AND2_X1 pool_pool_pe_b_peij_0_2_U4 ( .A1(pool_pool_pe_b_peij_0_2_d_acc[9]), 
        .A2(pool_pool_pe_b_peij_0_2_n14), .ZN(pool_pool_pe_b_peij_0_2_n2) );
  AND2_X1 pool_pool_pe_b_peij_0_2_U3 ( .A1(pool_pool_pe_b_peij_0_2_d_acc[10]), 
        .A2(pool_pool_pe_b_peij_0_2_n14), .ZN(pool_pool_pe_b_peij_0_2_n1) );
  DFFR_X1 pool_pool_pe_b_peij_0_2_q_acc_reg_10_ ( .D(
        pool_pool_pe_b_peij_0_2_n1), .CK(pool_pool_pe_b_peij_0_2_gck), .RN(
        pool_pool_pe_b_peij_0_2_n12), .Q(pool_pool_pe_b_o_data[153]) );
  DFFR_X1 pool_pool_pe_b_peij_0_2_q_acc_reg_9_ ( .D(pool_pool_pe_b_peij_0_2_n2), .CK(pool_pool_pe_b_peij_0_2_gck), .RN(pool_pool_pe_b_peij_0_2_n12), .Q(
        pool_pool_pe_b_o_data[152]) );
  DFFR_X1 pool_pool_pe_b_peij_0_2_q_acc_reg_8_ ( .D(pool_pool_pe_b_peij_0_2_n3), .CK(pool_pool_pe_b_peij_0_2_gck), .RN(pool_pool_pe_b_peij_0_2_n12), .Q(
        pool_pool_pe_b_o_data[151]) );
  DFFR_X1 pool_pool_pe_b_peij_0_2_q_acc_reg_7_ ( .D(pool_pool_pe_b_peij_0_2_n4), .CK(pool_pool_pe_b_peij_0_2_gck), .RN(pool_pool_pe_b_peij_0_2_n12), .Q(
        pool_pool_pe_b_o_data[150]) );
  DFFR_X1 pool_pool_pe_b_peij_0_2_q_acc_reg_6_ ( .D(pool_pool_pe_b_peij_0_2_n5), .CK(pool_pool_pe_b_peij_0_2_gck), .RN(pool_pool_pe_b_peij_0_2_n12), .Q(
        pool_pool_pe_b_o_data[149]) );
  DFFR_X1 pool_pool_pe_b_peij_0_2_q_acc_reg_5_ ( .D(pool_pool_pe_b_peij_0_2_n6), .CK(pool_pool_pe_b_peij_0_2_gck), .RN(pool_pool_pe_b_peij_0_2_n12), .Q(
        pool_pool_pe_b_o_data[148]) );
  DFFR_X1 pool_pool_pe_b_peij_0_2_q_acc_reg_4_ ( .D(pool_pool_pe_b_peij_0_2_n7), .CK(pool_pool_pe_b_peij_0_2_gck), .RN(pool_pool_pe_b_peij_0_2_n12), .Q(
        pool_pool_pe_b_o_data[147]) );
  DFFR_X1 pool_pool_pe_b_peij_0_2_q_acc_reg_3_ ( .D(pool_pool_pe_b_peij_0_2_n8), .CK(pool_pool_pe_b_peij_0_2_gck), .RN(pool_pool_pe_b_peij_0_2_n12), .Q(
        pool_pool_pe_b_o_data[146]) );
  DFFR_X1 pool_pool_pe_b_peij_0_2_q_acc_reg_2_ ( .D(pool_pool_pe_b_peij_0_2_n9), .CK(pool_pool_pe_b_peij_0_2_gck), .RN(pool_pool_pe_b_peij_0_2_n12), .Q(
        pool_pool_pe_b_o_data[145]) );
  DFFR_X1 pool_pool_pe_b_peij_0_2_q_acc_reg_1_ ( .D(
        pool_pool_pe_b_peij_0_2_n10), .CK(pool_pool_pe_b_peij_0_2_gck), .RN(
        pool_pool_pe_b_peij_0_2_n12), .Q(pool_pool_pe_b_o_data[144]) );
  DFFR_X1 pool_pool_pe_b_peij_0_2_q_acc_reg_0_ ( .D(
        pool_pool_pe_b_peij_0_2_n11), .CK(pool_pool_pe_b_peij_0_2_gck), .RN(
        pool_pool_pe_b_peij_0_2_n12), .Q(pool_pool_pe_b_o_data[143]) );
  AND3_X2 pool_pool_pe_b_peij_0_2_U20 ( .A1(pool_pool_pe_b_int_pe_en[13]), 
        .A2(clk), .A3(1'b1), .ZN(pool_pool_pe_b_peij_0_2_gck) );
  SDFFR_X1 pool_pool_pe_b_peij_0_2_q_k_reg ( .D(1'b0), .SI(
        pool_pool_pe_b_peij_0_2_n14), .SE(1'b0), .CK(
        pool_pool_pe_b_peij_0_2_gck), .RN(pool_pool_pe_b_peij_0_2_n12), .Q(
        pool_pool_pe_b_peij_0_2_q_k) );
  XOR2_X1 pool_pool_pe_b_peij_0_2_add_U11 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_2_q_k), .Z(pool_pool_pe_b_peij_0_2_add_notb[0])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_2_add_U10 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_2_q_k), .Z(pool_pool_pe_b_peij_0_2_add_notb[10])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_2_add_U9 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_2_q_k), .Z(pool_pool_pe_b_peij_0_2_add_notb[1])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_2_add_U8 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_2_q_k), .Z(pool_pool_pe_b_peij_0_2_add_notb[2])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_2_add_U7 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_2_q_k), .Z(pool_pool_pe_b_peij_0_2_add_notb[3])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_2_add_U6 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_2_q_k), .Z(pool_pool_pe_b_peij_0_2_add_notb[4])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_2_add_U5 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_2_q_k), .Z(pool_pool_pe_b_peij_0_2_add_notb[5])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_2_add_U4 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_2_q_k), .Z(pool_pool_pe_b_peij_0_2_add_notb[6])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_2_add_U3 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_2_q_k), .Z(pool_pool_pe_b_peij_0_2_add_notb[7])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_2_add_U2 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_2_q_k), .Z(pool_pool_pe_b_peij_0_2_add_notb[8])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_2_add_U1 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_2_q_k), .Z(pool_pool_pe_b_peij_0_2_add_notb[9])
         );
  INV_X2 pool_pool_pe_b_peij_0_2_add_fai_0_U2 ( .A(
        pool_pool_pe_b_peij_0_2_add_fai_0_n4), .ZN(
        pool_pool_pe_b_peij_0_2_add_cprop[1]) );
  XOR2_X1 pool_pool_pe_b_peij_0_2_add_fai_0_U4 ( .A(pool_pool_pe_b_o_data[143]), .B(pool_pool_pe_b_peij_0_2_add_notb[0]), .Z(
        pool_pool_pe_b_peij_0_2_add_fai_0_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_2_add_fai_0_U3 ( .A(
        pool_pool_pe_b_peij_0_2_q_k), .B(pool_pool_pe_b_peij_0_2_add_fai_0_n5), 
        .Z(pool_pool_pe_b_peij_0_2_d_acc[0]) );
  AOI22_X2 pool_pool_pe_b_peij_0_2_add_fai_0_U1 ( .A1(
        pool_pool_pe_b_peij_0_2_add_notb[0]), .A2(pool_pool_pe_b_o_data[143]), 
        .B1(pool_pool_pe_b_peij_0_2_add_fai_0_n5), .B2(
        pool_pool_pe_b_peij_0_2_q_k), .ZN(pool_pool_pe_b_peij_0_2_add_fai_0_n4) );
  INV_X2 pool_pool_pe_b_peij_0_2_add_fai_1_U2 ( .A(
        pool_pool_pe_b_peij_0_2_add_fai_1_n4), .ZN(
        pool_pool_pe_b_peij_0_2_add_cprop[2]) );
  XOR2_X1 pool_pool_pe_b_peij_0_2_add_fai_1_U4 ( .A(pool_pool_pe_b_o_data[144]), .B(pool_pool_pe_b_peij_0_2_add_notb[1]), .Z(
        pool_pool_pe_b_peij_0_2_add_fai_1_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_2_add_fai_1_U3 ( .A(
        pool_pool_pe_b_peij_0_2_add_cprop[1]), .B(
        pool_pool_pe_b_peij_0_2_add_fai_1_n5), .Z(
        pool_pool_pe_b_peij_0_2_d_acc[1]) );
  AOI22_X2 pool_pool_pe_b_peij_0_2_add_fai_1_U1 ( .A1(
        pool_pool_pe_b_peij_0_2_add_notb[1]), .A2(pool_pool_pe_b_o_data[144]), 
        .B1(pool_pool_pe_b_peij_0_2_add_fai_1_n5), .B2(
        pool_pool_pe_b_peij_0_2_add_cprop[1]), .ZN(
        pool_pool_pe_b_peij_0_2_add_fai_1_n4) );
  INV_X2 pool_pool_pe_b_peij_0_2_add_fai_2_U2 ( .A(
        pool_pool_pe_b_peij_0_2_add_fai_2_n4), .ZN(
        pool_pool_pe_b_peij_0_2_add_cprop[3]) );
  XOR2_X1 pool_pool_pe_b_peij_0_2_add_fai_2_U4 ( .A(pool_pool_pe_b_o_data[145]), .B(pool_pool_pe_b_peij_0_2_add_notb[2]), .Z(
        pool_pool_pe_b_peij_0_2_add_fai_2_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_2_add_fai_2_U3 ( .A(
        pool_pool_pe_b_peij_0_2_add_cprop[2]), .B(
        pool_pool_pe_b_peij_0_2_add_fai_2_n5), .Z(
        pool_pool_pe_b_peij_0_2_d_acc[2]) );
  AOI22_X2 pool_pool_pe_b_peij_0_2_add_fai_2_U1 ( .A1(
        pool_pool_pe_b_peij_0_2_add_notb[2]), .A2(pool_pool_pe_b_o_data[145]), 
        .B1(pool_pool_pe_b_peij_0_2_add_fai_2_n5), .B2(
        pool_pool_pe_b_peij_0_2_add_cprop[2]), .ZN(
        pool_pool_pe_b_peij_0_2_add_fai_2_n4) );
  INV_X2 pool_pool_pe_b_peij_0_2_add_fai_3_U2 ( .A(
        pool_pool_pe_b_peij_0_2_add_fai_3_n4), .ZN(
        pool_pool_pe_b_peij_0_2_add_cprop[4]) );
  XOR2_X1 pool_pool_pe_b_peij_0_2_add_fai_3_U4 ( .A(pool_pool_pe_b_o_data[146]), .B(pool_pool_pe_b_peij_0_2_add_notb[3]), .Z(
        pool_pool_pe_b_peij_0_2_add_fai_3_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_2_add_fai_3_U3 ( .A(
        pool_pool_pe_b_peij_0_2_add_cprop[3]), .B(
        pool_pool_pe_b_peij_0_2_add_fai_3_n5), .Z(
        pool_pool_pe_b_peij_0_2_d_acc[3]) );
  AOI22_X2 pool_pool_pe_b_peij_0_2_add_fai_3_U1 ( .A1(
        pool_pool_pe_b_peij_0_2_add_notb[3]), .A2(pool_pool_pe_b_o_data[146]), 
        .B1(pool_pool_pe_b_peij_0_2_add_fai_3_n5), .B2(
        pool_pool_pe_b_peij_0_2_add_cprop[3]), .ZN(
        pool_pool_pe_b_peij_0_2_add_fai_3_n4) );
  INV_X2 pool_pool_pe_b_peij_0_2_add_fai_4_U2 ( .A(
        pool_pool_pe_b_peij_0_2_add_fai_4_n4), .ZN(
        pool_pool_pe_b_peij_0_2_add_cprop[5]) );
  XOR2_X1 pool_pool_pe_b_peij_0_2_add_fai_4_U4 ( .A(pool_pool_pe_b_o_data[147]), .B(pool_pool_pe_b_peij_0_2_add_notb[4]), .Z(
        pool_pool_pe_b_peij_0_2_add_fai_4_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_2_add_fai_4_U3 ( .A(
        pool_pool_pe_b_peij_0_2_add_cprop[4]), .B(
        pool_pool_pe_b_peij_0_2_add_fai_4_n5), .Z(
        pool_pool_pe_b_peij_0_2_d_acc[4]) );
  AOI22_X2 pool_pool_pe_b_peij_0_2_add_fai_4_U1 ( .A1(
        pool_pool_pe_b_peij_0_2_add_notb[4]), .A2(pool_pool_pe_b_o_data[147]), 
        .B1(pool_pool_pe_b_peij_0_2_add_fai_4_n5), .B2(
        pool_pool_pe_b_peij_0_2_add_cprop[4]), .ZN(
        pool_pool_pe_b_peij_0_2_add_fai_4_n4) );
  INV_X2 pool_pool_pe_b_peij_0_2_add_fai_5_U2 ( .A(
        pool_pool_pe_b_peij_0_2_add_fai_5_n4), .ZN(
        pool_pool_pe_b_peij_0_2_add_cprop[6]) );
  XOR2_X1 pool_pool_pe_b_peij_0_2_add_fai_5_U4 ( .A(pool_pool_pe_b_o_data[148]), .B(pool_pool_pe_b_peij_0_2_add_notb[5]), .Z(
        pool_pool_pe_b_peij_0_2_add_fai_5_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_2_add_fai_5_U3 ( .A(
        pool_pool_pe_b_peij_0_2_add_cprop[5]), .B(
        pool_pool_pe_b_peij_0_2_add_fai_5_n5), .Z(
        pool_pool_pe_b_peij_0_2_d_acc[5]) );
  AOI22_X2 pool_pool_pe_b_peij_0_2_add_fai_5_U1 ( .A1(
        pool_pool_pe_b_peij_0_2_add_notb[5]), .A2(pool_pool_pe_b_o_data[148]), 
        .B1(pool_pool_pe_b_peij_0_2_add_fai_5_n5), .B2(
        pool_pool_pe_b_peij_0_2_add_cprop[5]), .ZN(
        pool_pool_pe_b_peij_0_2_add_fai_5_n4) );
  INV_X2 pool_pool_pe_b_peij_0_2_add_fai_6_U2 ( .A(
        pool_pool_pe_b_peij_0_2_add_fai_6_n4), .ZN(
        pool_pool_pe_b_peij_0_2_add_cprop[7]) );
  XOR2_X1 pool_pool_pe_b_peij_0_2_add_fai_6_U4 ( .A(pool_pool_pe_b_o_data[149]), .B(pool_pool_pe_b_peij_0_2_add_notb[6]), .Z(
        pool_pool_pe_b_peij_0_2_add_fai_6_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_2_add_fai_6_U3 ( .A(
        pool_pool_pe_b_peij_0_2_add_cprop[6]), .B(
        pool_pool_pe_b_peij_0_2_add_fai_6_n5), .Z(
        pool_pool_pe_b_peij_0_2_d_acc[6]) );
  AOI22_X2 pool_pool_pe_b_peij_0_2_add_fai_6_U1 ( .A1(
        pool_pool_pe_b_peij_0_2_add_notb[6]), .A2(pool_pool_pe_b_o_data[149]), 
        .B1(pool_pool_pe_b_peij_0_2_add_fai_6_n5), .B2(
        pool_pool_pe_b_peij_0_2_add_cprop[6]), .ZN(
        pool_pool_pe_b_peij_0_2_add_fai_6_n4) );
  INV_X2 pool_pool_pe_b_peij_0_2_add_fai_7_U2 ( .A(
        pool_pool_pe_b_peij_0_2_add_fai_7_n4), .ZN(
        pool_pool_pe_b_peij_0_2_add_cprop[8]) );
  XOR2_X1 pool_pool_pe_b_peij_0_2_add_fai_7_U4 ( .A(pool_pool_pe_b_o_data[150]), .B(pool_pool_pe_b_peij_0_2_add_notb[7]), .Z(
        pool_pool_pe_b_peij_0_2_add_fai_7_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_2_add_fai_7_U3 ( .A(
        pool_pool_pe_b_peij_0_2_add_cprop[7]), .B(
        pool_pool_pe_b_peij_0_2_add_fai_7_n5), .Z(
        pool_pool_pe_b_peij_0_2_d_acc[7]) );
  AOI22_X2 pool_pool_pe_b_peij_0_2_add_fai_7_U1 ( .A1(
        pool_pool_pe_b_peij_0_2_add_notb[7]), .A2(pool_pool_pe_b_o_data[150]), 
        .B1(pool_pool_pe_b_peij_0_2_add_fai_7_n5), .B2(
        pool_pool_pe_b_peij_0_2_add_cprop[7]), .ZN(
        pool_pool_pe_b_peij_0_2_add_fai_7_n4) );
  INV_X2 pool_pool_pe_b_peij_0_2_add_fai_8_U2 ( .A(
        pool_pool_pe_b_peij_0_2_add_fai_8_n4), .ZN(
        pool_pool_pe_b_peij_0_2_add_cprop[9]) );
  XOR2_X1 pool_pool_pe_b_peij_0_2_add_fai_8_U4 ( .A(pool_pool_pe_b_o_data[151]), .B(pool_pool_pe_b_peij_0_2_add_notb[8]), .Z(
        pool_pool_pe_b_peij_0_2_add_fai_8_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_2_add_fai_8_U3 ( .A(
        pool_pool_pe_b_peij_0_2_add_cprop[8]), .B(
        pool_pool_pe_b_peij_0_2_add_fai_8_n5), .Z(
        pool_pool_pe_b_peij_0_2_d_acc[8]) );
  AOI22_X2 pool_pool_pe_b_peij_0_2_add_fai_8_U1 ( .A1(
        pool_pool_pe_b_peij_0_2_add_notb[8]), .A2(pool_pool_pe_b_o_data[151]), 
        .B1(pool_pool_pe_b_peij_0_2_add_fai_8_n5), .B2(
        pool_pool_pe_b_peij_0_2_add_cprop[8]), .ZN(
        pool_pool_pe_b_peij_0_2_add_fai_8_n4) );
  INV_X2 pool_pool_pe_b_peij_0_2_add_fai_9_U2 ( .A(
        pool_pool_pe_b_peij_0_2_add_fai_9_n4), .ZN(
        pool_pool_pe_b_peij_0_2_add_cprop[10]) );
  XOR2_X1 pool_pool_pe_b_peij_0_2_add_fai_9_U4 ( .A(pool_pool_pe_b_o_data[152]), .B(pool_pool_pe_b_peij_0_2_add_notb[9]), .Z(
        pool_pool_pe_b_peij_0_2_add_fai_9_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_2_add_fai_9_U3 ( .A(
        pool_pool_pe_b_peij_0_2_add_cprop[9]), .B(
        pool_pool_pe_b_peij_0_2_add_fai_9_n5), .Z(
        pool_pool_pe_b_peij_0_2_d_acc[9]) );
  AOI22_X2 pool_pool_pe_b_peij_0_2_add_fai_9_U1 ( .A1(
        pool_pool_pe_b_peij_0_2_add_notb[9]), .A2(pool_pool_pe_b_o_data[152]), 
        .B1(pool_pool_pe_b_peij_0_2_add_fai_9_n5), .B2(
        pool_pool_pe_b_peij_0_2_add_cprop[9]), .ZN(
        pool_pool_pe_b_peij_0_2_add_fai_9_n4) );
  INV_X2 pool_pool_pe_b_peij_0_2_add_fai_10_U2 ( .A(
        pool_pool_pe_b_peij_0_2_add_fai_10_n4), .ZN(
        pool_pool_pe_b_peij_0_2_add_c_out) );
  XOR2_X1 pool_pool_pe_b_peij_0_2_add_fai_10_U4 ( .A(
        pool_pool_pe_b_o_data[153]), .B(pool_pool_pe_b_peij_0_2_add_notb[10]), 
        .Z(pool_pool_pe_b_peij_0_2_add_fai_10_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_2_add_fai_10_U3 ( .A(
        pool_pool_pe_b_peij_0_2_add_cprop[10]), .B(
        pool_pool_pe_b_peij_0_2_add_fai_10_n5), .Z(
        pool_pool_pe_b_peij_0_2_d_acc[10]) );
  AOI22_X2 pool_pool_pe_b_peij_0_2_add_fai_10_U1 ( .A1(
        pool_pool_pe_b_peij_0_2_add_notb[10]), .A2(pool_pool_pe_b_o_data[153]), 
        .B1(pool_pool_pe_b_peij_0_2_add_fai_10_n5), .B2(
        pool_pool_pe_b_peij_0_2_add_cprop[10]), .ZN(
        pool_pool_pe_b_peij_0_2_add_fai_10_n4) );
  INV_X2 pool_pool_pe_b_peij_0_3_U21 ( .A(pool_sync_clr), .ZN(
        pool_pool_pe_b_peij_0_3_n14) );
  INV_X1 pool_pool_pe_b_peij_0_3_U18 ( .A(pool_pool_pe_b_n6), .ZN(
        pool_pool_pe_b_peij_0_3_n12) );
  AND2_X1 pool_pool_pe_b_peij_0_3_U13 ( .A1(pool_pool_pe_b_peij_0_3_d_acc[0]), 
        .A2(pool_pool_pe_b_peij_0_3_n14), .ZN(pool_pool_pe_b_peij_0_3_n11) );
  AND2_X1 pool_pool_pe_b_peij_0_3_U12 ( .A1(pool_pool_pe_b_peij_0_3_d_acc[1]), 
        .A2(pool_pool_pe_b_peij_0_3_n14), .ZN(pool_pool_pe_b_peij_0_3_n10) );
  AND2_X1 pool_pool_pe_b_peij_0_3_U11 ( .A1(pool_pool_pe_b_peij_0_3_d_acc[2]), 
        .A2(pool_pool_pe_b_peij_0_3_n14), .ZN(pool_pool_pe_b_peij_0_3_n9) );
  AND2_X1 pool_pool_pe_b_peij_0_3_U10 ( .A1(pool_pool_pe_b_peij_0_3_d_acc[3]), 
        .A2(pool_pool_pe_b_peij_0_3_n14), .ZN(pool_pool_pe_b_peij_0_3_n8) );
  AND2_X1 pool_pool_pe_b_peij_0_3_U9 ( .A1(pool_pool_pe_b_peij_0_3_d_acc[4]), 
        .A2(pool_pool_pe_b_peij_0_3_n14), .ZN(pool_pool_pe_b_peij_0_3_n7) );
  AND2_X1 pool_pool_pe_b_peij_0_3_U8 ( .A1(pool_pool_pe_b_peij_0_3_d_acc[5]), 
        .A2(pool_pool_pe_b_peij_0_3_n14), .ZN(pool_pool_pe_b_peij_0_3_n6) );
  AND2_X1 pool_pool_pe_b_peij_0_3_U7 ( .A1(pool_pool_pe_b_peij_0_3_d_acc[6]), 
        .A2(pool_pool_pe_b_peij_0_3_n14), .ZN(pool_pool_pe_b_peij_0_3_n5) );
  AND2_X1 pool_pool_pe_b_peij_0_3_U6 ( .A1(pool_pool_pe_b_peij_0_3_d_acc[7]), 
        .A2(pool_pool_pe_b_peij_0_3_n14), .ZN(pool_pool_pe_b_peij_0_3_n4) );
  AND2_X1 pool_pool_pe_b_peij_0_3_U5 ( .A1(pool_pool_pe_b_peij_0_3_d_acc[8]), 
        .A2(pool_pool_pe_b_peij_0_3_n14), .ZN(pool_pool_pe_b_peij_0_3_n3) );
  AND2_X1 pool_pool_pe_b_peij_0_3_U4 ( .A1(pool_pool_pe_b_peij_0_3_d_acc[9]), 
        .A2(pool_pool_pe_b_peij_0_3_n14), .ZN(pool_pool_pe_b_peij_0_3_n2) );
  AND2_X1 pool_pool_pe_b_peij_0_3_U3 ( .A1(pool_pool_pe_b_peij_0_3_d_acc[10]), 
        .A2(pool_pool_pe_b_peij_0_3_n14), .ZN(pool_pool_pe_b_peij_0_3_n1) );
  DFFR_X1 pool_pool_pe_b_peij_0_3_q_acc_reg_10_ ( .D(
        pool_pool_pe_b_peij_0_3_n1), .CK(pool_pool_pe_b_peij_0_3_gck), .RN(
        pool_pool_pe_b_peij_0_3_n12), .Q(pool_pool_pe_b_o_data[142]) );
  DFFR_X1 pool_pool_pe_b_peij_0_3_q_acc_reg_9_ ( .D(pool_pool_pe_b_peij_0_3_n2), .CK(pool_pool_pe_b_peij_0_3_gck), .RN(pool_pool_pe_b_peij_0_3_n12), .Q(
        pool_pool_pe_b_o_data[141]) );
  DFFR_X1 pool_pool_pe_b_peij_0_3_q_acc_reg_8_ ( .D(pool_pool_pe_b_peij_0_3_n3), .CK(pool_pool_pe_b_peij_0_3_gck), .RN(pool_pool_pe_b_peij_0_3_n12), .Q(
        pool_pool_pe_b_o_data[140]) );
  DFFR_X1 pool_pool_pe_b_peij_0_3_q_acc_reg_7_ ( .D(pool_pool_pe_b_peij_0_3_n4), .CK(pool_pool_pe_b_peij_0_3_gck), .RN(pool_pool_pe_b_peij_0_3_n12), .Q(
        pool_pool_pe_b_o_data[139]) );
  DFFR_X1 pool_pool_pe_b_peij_0_3_q_acc_reg_6_ ( .D(pool_pool_pe_b_peij_0_3_n5), .CK(pool_pool_pe_b_peij_0_3_gck), .RN(pool_pool_pe_b_peij_0_3_n12), .Q(
        pool_pool_pe_b_o_data[138]) );
  DFFR_X1 pool_pool_pe_b_peij_0_3_q_acc_reg_5_ ( .D(pool_pool_pe_b_peij_0_3_n6), .CK(pool_pool_pe_b_peij_0_3_gck), .RN(pool_pool_pe_b_peij_0_3_n12), .Q(
        pool_pool_pe_b_o_data[137]) );
  DFFR_X1 pool_pool_pe_b_peij_0_3_q_acc_reg_4_ ( .D(pool_pool_pe_b_peij_0_3_n7), .CK(pool_pool_pe_b_peij_0_3_gck), .RN(pool_pool_pe_b_peij_0_3_n12), .Q(
        pool_pool_pe_b_o_data[136]) );
  DFFR_X1 pool_pool_pe_b_peij_0_3_q_acc_reg_3_ ( .D(pool_pool_pe_b_peij_0_3_n8), .CK(pool_pool_pe_b_peij_0_3_gck), .RN(pool_pool_pe_b_peij_0_3_n12), .Q(
        pool_pool_pe_b_o_data[135]) );
  DFFR_X1 pool_pool_pe_b_peij_0_3_q_acc_reg_2_ ( .D(pool_pool_pe_b_peij_0_3_n9), .CK(pool_pool_pe_b_peij_0_3_gck), .RN(pool_pool_pe_b_peij_0_3_n12), .Q(
        pool_pool_pe_b_o_data[134]) );
  DFFR_X1 pool_pool_pe_b_peij_0_3_q_acc_reg_1_ ( .D(
        pool_pool_pe_b_peij_0_3_n10), .CK(pool_pool_pe_b_peij_0_3_gck), .RN(
        pool_pool_pe_b_peij_0_3_n12), .Q(pool_pool_pe_b_o_data[133]) );
  DFFR_X1 pool_pool_pe_b_peij_0_3_q_acc_reg_0_ ( .D(
        pool_pool_pe_b_peij_0_3_n11), .CK(pool_pool_pe_b_peij_0_3_gck), .RN(
        pool_pool_pe_b_peij_0_3_n12), .Q(pool_pool_pe_b_o_data[132]) );
  AND3_X2 pool_pool_pe_b_peij_0_3_U20 ( .A1(pool_pool_pe_b_int_pe_en[12]), 
        .A2(clk), .A3(1'b1), .ZN(pool_pool_pe_b_peij_0_3_gck) );
  SDFFR_X1 pool_pool_pe_b_peij_0_3_q_k_reg ( .D(1'b0), .SI(
        pool_pool_pe_b_peij_0_3_n14), .SE(1'b0), .CK(
        pool_pool_pe_b_peij_0_3_gck), .RN(pool_pool_pe_b_peij_0_3_n12), .Q(
        pool_pool_pe_b_peij_0_3_q_k) );
  XOR2_X1 pool_pool_pe_b_peij_0_3_add_U11 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_3_q_k), .Z(pool_pool_pe_b_peij_0_3_add_notb[0])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_3_add_U10 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_3_q_k), .Z(pool_pool_pe_b_peij_0_3_add_notb[10])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_3_add_U9 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_3_q_k), .Z(pool_pool_pe_b_peij_0_3_add_notb[1])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_3_add_U8 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_3_q_k), .Z(pool_pool_pe_b_peij_0_3_add_notb[2])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_3_add_U7 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_3_q_k), .Z(pool_pool_pe_b_peij_0_3_add_notb[3])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_3_add_U6 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_3_q_k), .Z(pool_pool_pe_b_peij_0_3_add_notb[4])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_3_add_U5 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_3_q_k), .Z(pool_pool_pe_b_peij_0_3_add_notb[5])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_3_add_U4 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_3_q_k), .Z(pool_pool_pe_b_peij_0_3_add_notb[6])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_3_add_U3 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_3_q_k), .Z(pool_pool_pe_b_peij_0_3_add_notb[7])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_3_add_U2 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_3_q_k), .Z(pool_pool_pe_b_peij_0_3_add_notb[8])
         );
  XOR2_X1 pool_pool_pe_b_peij_0_3_add_U1 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_0_3_q_k), .Z(pool_pool_pe_b_peij_0_3_add_notb[9])
         );
  INV_X2 pool_pool_pe_b_peij_0_3_add_fai_0_U2 ( .A(
        pool_pool_pe_b_peij_0_3_add_fai_0_n4), .ZN(
        pool_pool_pe_b_peij_0_3_add_cprop[1]) );
  XOR2_X1 pool_pool_pe_b_peij_0_3_add_fai_0_U4 ( .A(pool_pool_pe_b_o_data[132]), .B(pool_pool_pe_b_peij_0_3_add_notb[0]), .Z(
        pool_pool_pe_b_peij_0_3_add_fai_0_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_3_add_fai_0_U3 ( .A(
        pool_pool_pe_b_peij_0_3_q_k), .B(pool_pool_pe_b_peij_0_3_add_fai_0_n5), 
        .Z(pool_pool_pe_b_peij_0_3_d_acc[0]) );
  AOI22_X2 pool_pool_pe_b_peij_0_3_add_fai_0_U1 ( .A1(
        pool_pool_pe_b_peij_0_3_add_notb[0]), .A2(pool_pool_pe_b_o_data[132]), 
        .B1(pool_pool_pe_b_peij_0_3_add_fai_0_n5), .B2(
        pool_pool_pe_b_peij_0_3_q_k), .ZN(pool_pool_pe_b_peij_0_3_add_fai_0_n4) );
  INV_X2 pool_pool_pe_b_peij_0_3_add_fai_1_U2 ( .A(
        pool_pool_pe_b_peij_0_3_add_fai_1_n4), .ZN(
        pool_pool_pe_b_peij_0_3_add_cprop[2]) );
  XOR2_X1 pool_pool_pe_b_peij_0_3_add_fai_1_U4 ( .A(pool_pool_pe_b_o_data[133]), .B(pool_pool_pe_b_peij_0_3_add_notb[1]), .Z(
        pool_pool_pe_b_peij_0_3_add_fai_1_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_3_add_fai_1_U3 ( .A(
        pool_pool_pe_b_peij_0_3_add_cprop[1]), .B(
        pool_pool_pe_b_peij_0_3_add_fai_1_n5), .Z(
        pool_pool_pe_b_peij_0_3_d_acc[1]) );
  AOI22_X2 pool_pool_pe_b_peij_0_3_add_fai_1_U1 ( .A1(
        pool_pool_pe_b_peij_0_3_add_notb[1]), .A2(pool_pool_pe_b_o_data[133]), 
        .B1(pool_pool_pe_b_peij_0_3_add_fai_1_n5), .B2(
        pool_pool_pe_b_peij_0_3_add_cprop[1]), .ZN(
        pool_pool_pe_b_peij_0_3_add_fai_1_n4) );
  INV_X2 pool_pool_pe_b_peij_0_3_add_fai_2_U2 ( .A(
        pool_pool_pe_b_peij_0_3_add_fai_2_n4), .ZN(
        pool_pool_pe_b_peij_0_3_add_cprop[3]) );
  XOR2_X1 pool_pool_pe_b_peij_0_3_add_fai_2_U4 ( .A(pool_pool_pe_b_o_data[134]), .B(pool_pool_pe_b_peij_0_3_add_notb[2]), .Z(
        pool_pool_pe_b_peij_0_3_add_fai_2_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_3_add_fai_2_U3 ( .A(
        pool_pool_pe_b_peij_0_3_add_cprop[2]), .B(
        pool_pool_pe_b_peij_0_3_add_fai_2_n5), .Z(
        pool_pool_pe_b_peij_0_3_d_acc[2]) );
  AOI22_X2 pool_pool_pe_b_peij_0_3_add_fai_2_U1 ( .A1(
        pool_pool_pe_b_peij_0_3_add_notb[2]), .A2(pool_pool_pe_b_o_data[134]), 
        .B1(pool_pool_pe_b_peij_0_3_add_fai_2_n5), .B2(
        pool_pool_pe_b_peij_0_3_add_cprop[2]), .ZN(
        pool_pool_pe_b_peij_0_3_add_fai_2_n4) );
  INV_X2 pool_pool_pe_b_peij_0_3_add_fai_3_U2 ( .A(
        pool_pool_pe_b_peij_0_3_add_fai_3_n4), .ZN(
        pool_pool_pe_b_peij_0_3_add_cprop[4]) );
  XOR2_X1 pool_pool_pe_b_peij_0_3_add_fai_3_U4 ( .A(pool_pool_pe_b_o_data[135]), .B(pool_pool_pe_b_peij_0_3_add_notb[3]), .Z(
        pool_pool_pe_b_peij_0_3_add_fai_3_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_3_add_fai_3_U3 ( .A(
        pool_pool_pe_b_peij_0_3_add_cprop[3]), .B(
        pool_pool_pe_b_peij_0_3_add_fai_3_n5), .Z(
        pool_pool_pe_b_peij_0_3_d_acc[3]) );
  AOI22_X2 pool_pool_pe_b_peij_0_3_add_fai_3_U1 ( .A1(
        pool_pool_pe_b_peij_0_3_add_notb[3]), .A2(pool_pool_pe_b_o_data[135]), 
        .B1(pool_pool_pe_b_peij_0_3_add_fai_3_n5), .B2(
        pool_pool_pe_b_peij_0_3_add_cprop[3]), .ZN(
        pool_pool_pe_b_peij_0_3_add_fai_3_n4) );
  INV_X2 pool_pool_pe_b_peij_0_3_add_fai_4_U2 ( .A(
        pool_pool_pe_b_peij_0_3_add_fai_4_n4), .ZN(
        pool_pool_pe_b_peij_0_3_add_cprop[5]) );
  XOR2_X1 pool_pool_pe_b_peij_0_3_add_fai_4_U4 ( .A(pool_pool_pe_b_o_data[136]), .B(pool_pool_pe_b_peij_0_3_add_notb[4]), .Z(
        pool_pool_pe_b_peij_0_3_add_fai_4_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_3_add_fai_4_U3 ( .A(
        pool_pool_pe_b_peij_0_3_add_cprop[4]), .B(
        pool_pool_pe_b_peij_0_3_add_fai_4_n5), .Z(
        pool_pool_pe_b_peij_0_3_d_acc[4]) );
  AOI22_X2 pool_pool_pe_b_peij_0_3_add_fai_4_U1 ( .A1(
        pool_pool_pe_b_peij_0_3_add_notb[4]), .A2(pool_pool_pe_b_o_data[136]), 
        .B1(pool_pool_pe_b_peij_0_3_add_fai_4_n5), .B2(
        pool_pool_pe_b_peij_0_3_add_cprop[4]), .ZN(
        pool_pool_pe_b_peij_0_3_add_fai_4_n4) );
  INV_X2 pool_pool_pe_b_peij_0_3_add_fai_5_U2 ( .A(
        pool_pool_pe_b_peij_0_3_add_fai_5_n4), .ZN(
        pool_pool_pe_b_peij_0_3_add_cprop[6]) );
  XOR2_X1 pool_pool_pe_b_peij_0_3_add_fai_5_U4 ( .A(pool_pool_pe_b_o_data[137]), .B(pool_pool_pe_b_peij_0_3_add_notb[5]), .Z(
        pool_pool_pe_b_peij_0_3_add_fai_5_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_3_add_fai_5_U3 ( .A(
        pool_pool_pe_b_peij_0_3_add_cprop[5]), .B(
        pool_pool_pe_b_peij_0_3_add_fai_5_n5), .Z(
        pool_pool_pe_b_peij_0_3_d_acc[5]) );
  AOI22_X2 pool_pool_pe_b_peij_0_3_add_fai_5_U1 ( .A1(
        pool_pool_pe_b_peij_0_3_add_notb[5]), .A2(pool_pool_pe_b_o_data[137]), 
        .B1(pool_pool_pe_b_peij_0_3_add_fai_5_n5), .B2(
        pool_pool_pe_b_peij_0_3_add_cprop[5]), .ZN(
        pool_pool_pe_b_peij_0_3_add_fai_5_n4) );
  INV_X2 pool_pool_pe_b_peij_0_3_add_fai_6_U2 ( .A(
        pool_pool_pe_b_peij_0_3_add_fai_6_n4), .ZN(
        pool_pool_pe_b_peij_0_3_add_cprop[7]) );
  XOR2_X1 pool_pool_pe_b_peij_0_3_add_fai_6_U4 ( .A(pool_pool_pe_b_o_data[138]), .B(pool_pool_pe_b_peij_0_3_add_notb[6]), .Z(
        pool_pool_pe_b_peij_0_3_add_fai_6_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_3_add_fai_6_U3 ( .A(
        pool_pool_pe_b_peij_0_3_add_cprop[6]), .B(
        pool_pool_pe_b_peij_0_3_add_fai_6_n5), .Z(
        pool_pool_pe_b_peij_0_3_d_acc[6]) );
  AOI22_X2 pool_pool_pe_b_peij_0_3_add_fai_6_U1 ( .A1(
        pool_pool_pe_b_peij_0_3_add_notb[6]), .A2(pool_pool_pe_b_o_data[138]), 
        .B1(pool_pool_pe_b_peij_0_3_add_fai_6_n5), .B2(
        pool_pool_pe_b_peij_0_3_add_cprop[6]), .ZN(
        pool_pool_pe_b_peij_0_3_add_fai_6_n4) );
  INV_X2 pool_pool_pe_b_peij_0_3_add_fai_7_U2 ( .A(
        pool_pool_pe_b_peij_0_3_add_fai_7_n4), .ZN(
        pool_pool_pe_b_peij_0_3_add_cprop[8]) );
  XOR2_X1 pool_pool_pe_b_peij_0_3_add_fai_7_U4 ( .A(pool_pool_pe_b_o_data[139]), .B(pool_pool_pe_b_peij_0_3_add_notb[7]), .Z(
        pool_pool_pe_b_peij_0_3_add_fai_7_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_3_add_fai_7_U3 ( .A(
        pool_pool_pe_b_peij_0_3_add_cprop[7]), .B(
        pool_pool_pe_b_peij_0_3_add_fai_7_n5), .Z(
        pool_pool_pe_b_peij_0_3_d_acc[7]) );
  AOI22_X2 pool_pool_pe_b_peij_0_3_add_fai_7_U1 ( .A1(
        pool_pool_pe_b_peij_0_3_add_notb[7]), .A2(pool_pool_pe_b_o_data[139]), 
        .B1(pool_pool_pe_b_peij_0_3_add_fai_7_n5), .B2(
        pool_pool_pe_b_peij_0_3_add_cprop[7]), .ZN(
        pool_pool_pe_b_peij_0_3_add_fai_7_n4) );
  INV_X2 pool_pool_pe_b_peij_0_3_add_fai_8_U2 ( .A(
        pool_pool_pe_b_peij_0_3_add_fai_8_n4), .ZN(
        pool_pool_pe_b_peij_0_3_add_cprop[9]) );
  XOR2_X1 pool_pool_pe_b_peij_0_3_add_fai_8_U4 ( .A(pool_pool_pe_b_o_data[140]), .B(pool_pool_pe_b_peij_0_3_add_notb[8]), .Z(
        pool_pool_pe_b_peij_0_3_add_fai_8_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_3_add_fai_8_U3 ( .A(
        pool_pool_pe_b_peij_0_3_add_cprop[8]), .B(
        pool_pool_pe_b_peij_0_3_add_fai_8_n5), .Z(
        pool_pool_pe_b_peij_0_3_d_acc[8]) );
  AOI22_X2 pool_pool_pe_b_peij_0_3_add_fai_8_U1 ( .A1(
        pool_pool_pe_b_peij_0_3_add_notb[8]), .A2(pool_pool_pe_b_o_data[140]), 
        .B1(pool_pool_pe_b_peij_0_3_add_fai_8_n5), .B2(
        pool_pool_pe_b_peij_0_3_add_cprop[8]), .ZN(
        pool_pool_pe_b_peij_0_3_add_fai_8_n4) );
  INV_X2 pool_pool_pe_b_peij_0_3_add_fai_9_U2 ( .A(
        pool_pool_pe_b_peij_0_3_add_fai_9_n4), .ZN(
        pool_pool_pe_b_peij_0_3_add_cprop[10]) );
  XOR2_X1 pool_pool_pe_b_peij_0_3_add_fai_9_U4 ( .A(pool_pool_pe_b_o_data[141]), .B(pool_pool_pe_b_peij_0_3_add_notb[9]), .Z(
        pool_pool_pe_b_peij_0_3_add_fai_9_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_3_add_fai_9_U3 ( .A(
        pool_pool_pe_b_peij_0_3_add_cprop[9]), .B(
        pool_pool_pe_b_peij_0_3_add_fai_9_n5), .Z(
        pool_pool_pe_b_peij_0_3_d_acc[9]) );
  AOI22_X2 pool_pool_pe_b_peij_0_3_add_fai_9_U1 ( .A1(
        pool_pool_pe_b_peij_0_3_add_notb[9]), .A2(pool_pool_pe_b_o_data[141]), 
        .B1(pool_pool_pe_b_peij_0_3_add_fai_9_n5), .B2(
        pool_pool_pe_b_peij_0_3_add_cprop[9]), .ZN(
        pool_pool_pe_b_peij_0_3_add_fai_9_n4) );
  INV_X2 pool_pool_pe_b_peij_0_3_add_fai_10_U2 ( .A(
        pool_pool_pe_b_peij_0_3_add_fai_10_n4), .ZN(
        pool_pool_pe_b_peij_0_3_add_c_out) );
  XOR2_X1 pool_pool_pe_b_peij_0_3_add_fai_10_U4 ( .A(
        pool_pool_pe_b_o_data[142]), .B(pool_pool_pe_b_peij_0_3_add_notb[10]), 
        .Z(pool_pool_pe_b_peij_0_3_add_fai_10_n5) );
  XOR2_X1 pool_pool_pe_b_peij_0_3_add_fai_10_U3 ( .A(
        pool_pool_pe_b_peij_0_3_add_cprop[10]), .B(
        pool_pool_pe_b_peij_0_3_add_fai_10_n5), .Z(
        pool_pool_pe_b_peij_0_3_d_acc[10]) );
  AOI22_X2 pool_pool_pe_b_peij_0_3_add_fai_10_U1 ( .A1(
        pool_pool_pe_b_peij_0_3_add_notb[10]), .A2(pool_pool_pe_b_o_data[142]), 
        .B1(pool_pool_pe_b_peij_0_3_add_fai_10_n5), .B2(
        pool_pool_pe_b_peij_0_3_add_cprop[10]), .ZN(
        pool_pool_pe_b_peij_0_3_add_fai_10_n4) );
  INV_X2 pool_pool_pe_b_peij_1_0_U21 ( .A(pool_sync_clr), .ZN(
        pool_pool_pe_b_peij_1_0_n14) );
  INV_X1 pool_pool_pe_b_peij_1_0_U18 ( .A(pool_pool_pe_b_n6), .ZN(
        pool_pool_pe_b_peij_1_0_n12) );
  AND2_X1 pool_pool_pe_b_peij_1_0_U13 ( .A1(pool_pool_pe_b_peij_1_0_d_acc[0]), 
        .A2(pool_pool_pe_b_peij_1_0_n14), .ZN(pool_pool_pe_b_peij_1_0_n11) );
  AND2_X1 pool_pool_pe_b_peij_1_0_U12 ( .A1(pool_pool_pe_b_peij_1_0_d_acc[1]), 
        .A2(pool_pool_pe_b_peij_1_0_n14), .ZN(pool_pool_pe_b_peij_1_0_n10) );
  AND2_X1 pool_pool_pe_b_peij_1_0_U11 ( .A1(pool_pool_pe_b_peij_1_0_d_acc[2]), 
        .A2(pool_pool_pe_b_peij_1_0_n14), .ZN(pool_pool_pe_b_peij_1_0_n9) );
  AND2_X1 pool_pool_pe_b_peij_1_0_U10 ( .A1(pool_pool_pe_b_peij_1_0_d_acc[3]), 
        .A2(pool_pool_pe_b_peij_1_0_n14), .ZN(pool_pool_pe_b_peij_1_0_n8) );
  AND2_X1 pool_pool_pe_b_peij_1_0_U9 ( .A1(pool_pool_pe_b_peij_1_0_d_acc[4]), 
        .A2(pool_pool_pe_b_peij_1_0_n14), .ZN(pool_pool_pe_b_peij_1_0_n7) );
  AND2_X1 pool_pool_pe_b_peij_1_0_U8 ( .A1(pool_pool_pe_b_peij_1_0_d_acc[5]), 
        .A2(pool_pool_pe_b_peij_1_0_n14), .ZN(pool_pool_pe_b_peij_1_0_n6) );
  AND2_X1 pool_pool_pe_b_peij_1_0_U7 ( .A1(pool_pool_pe_b_peij_1_0_d_acc[6]), 
        .A2(pool_pool_pe_b_peij_1_0_n14), .ZN(pool_pool_pe_b_peij_1_0_n5) );
  AND2_X1 pool_pool_pe_b_peij_1_0_U6 ( .A1(pool_pool_pe_b_peij_1_0_d_acc[7]), 
        .A2(pool_pool_pe_b_peij_1_0_n14), .ZN(pool_pool_pe_b_peij_1_0_n4) );
  AND2_X1 pool_pool_pe_b_peij_1_0_U5 ( .A1(pool_pool_pe_b_peij_1_0_d_acc[8]), 
        .A2(pool_pool_pe_b_peij_1_0_n14), .ZN(pool_pool_pe_b_peij_1_0_n3) );
  AND2_X1 pool_pool_pe_b_peij_1_0_U4 ( .A1(pool_pool_pe_b_peij_1_0_d_acc[9]), 
        .A2(pool_pool_pe_b_peij_1_0_n14), .ZN(pool_pool_pe_b_peij_1_0_n2) );
  AND2_X1 pool_pool_pe_b_peij_1_0_U3 ( .A1(pool_pool_pe_b_peij_1_0_d_acc[10]), 
        .A2(pool_pool_pe_b_peij_1_0_n14), .ZN(pool_pool_pe_b_peij_1_0_n1) );
  DFFR_X1 pool_pool_pe_b_peij_1_0_q_acc_reg_10_ ( .D(
        pool_pool_pe_b_peij_1_0_n1), .CK(pool_pool_pe_b_peij_1_0_gck), .RN(
        pool_pool_pe_b_peij_1_0_n12), .Q(pool_pool_pe_b_o_data[131]) );
  DFFR_X1 pool_pool_pe_b_peij_1_0_q_acc_reg_9_ ( .D(pool_pool_pe_b_peij_1_0_n2), .CK(pool_pool_pe_b_peij_1_0_gck), .RN(pool_pool_pe_b_peij_1_0_n12), .Q(
        pool_pool_pe_b_o_data[130]) );
  DFFR_X1 pool_pool_pe_b_peij_1_0_q_acc_reg_8_ ( .D(pool_pool_pe_b_peij_1_0_n3), .CK(pool_pool_pe_b_peij_1_0_gck), .RN(pool_pool_pe_b_peij_1_0_n12), .Q(
        pool_pool_pe_b_o_data[129]) );
  DFFR_X1 pool_pool_pe_b_peij_1_0_q_acc_reg_7_ ( .D(pool_pool_pe_b_peij_1_0_n4), .CK(pool_pool_pe_b_peij_1_0_gck), .RN(pool_pool_pe_b_peij_1_0_n12), .Q(
        pool_pool_pe_b_o_data[128]) );
  DFFR_X1 pool_pool_pe_b_peij_1_0_q_acc_reg_6_ ( .D(pool_pool_pe_b_peij_1_0_n5), .CK(pool_pool_pe_b_peij_1_0_gck), .RN(pool_pool_pe_b_peij_1_0_n12), .Q(
        pool_pool_pe_b_o_data[127]) );
  DFFR_X1 pool_pool_pe_b_peij_1_0_q_acc_reg_5_ ( .D(pool_pool_pe_b_peij_1_0_n6), .CK(pool_pool_pe_b_peij_1_0_gck), .RN(pool_pool_pe_b_peij_1_0_n12), .Q(
        pool_pool_pe_b_o_data[126]) );
  DFFR_X1 pool_pool_pe_b_peij_1_0_q_acc_reg_4_ ( .D(pool_pool_pe_b_peij_1_0_n7), .CK(pool_pool_pe_b_peij_1_0_gck), .RN(pool_pool_pe_b_peij_1_0_n12), .Q(
        pool_pool_pe_b_o_data[125]) );
  DFFR_X1 pool_pool_pe_b_peij_1_0_q_acc_reg_3_ ( .D(pool_pool_pe_b_peij_1_0_n8), .CK(pool_pool_pe_b_peij_1_0_gck), .RN(pool_pool_pe_b_peij_1_0_n12), .Q(
        pool_pool_pe_b_o_data[124]) );
  DFFR_X1 pool_pool_pe_b_peij_1_0_q_acc_reg_2_ ( .D(pool_pool_pe_b_peij_1_0_n9), .CK(pool_pool_pe_b_peij_1_0_gck), .RN(pool_pool_pe_b_peij_1_0_n12), .Q(
        pool_pool_pe_b_o_data[123]) );
  DFFR_X1 pool_pool_pe_b_peij_1_0_q_acc_reg_1_ ( .D(
        pool_pool_pe_b_peij_1_0_n10), .CK(pool_pool_pe_b_peij_1_0_gck), .RN(
        pool_pool_pe_b_peij_1_0_n12), .Q(pool_pool_pe_b_o_data[122]) );
  DFFR_X1 pool_pool_pe_b_peij_1_0_q_acc_reg_0_ ( .D(
        pool_pool_pe_b_peij_1_0_n11), .CK(pool_pool_pe_b_peij_1_0_gck), .RN(
        pool_pool_pe_b_peij_1_0_n12), .Q(pool_pool_pe_b_o_data[121]) );
  AND3_X2 pool_pool_pe_b_peij_1_0_U20 ( .A1(pool_pool_pe_b_int_pe_en[11]), 
        .A2(clk), .A3(1'b1), .ZN(pool_pool_pe_b_peij_1_0_gck) );
  SDFFR_X1 pool_pool_pe_b_peij_1_0_q_k_reg ( .D(1'b0), .SI(
        pool_pool_pe_b_peij_1_0_n14), .SE(1'b0), .CK(
        pool_pool_pe_b_peij_1_0_gck), .RN(pool_pool_pe_b_peij_1_0_n12), .Q(
        pool_pool_pe_b_peij_1_0_q_k) );
  XOR2_X1 pool_pool_pe_b_peij_1_0_add_U11 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_0_q_k), .Z(pool_pool_pe_b_peij_1_0_add_notb[0])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_0_add_U10 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_0_q_k), .Z(pool_pool_pe_b_peij_1_0_add_notb[10])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_0_add_U9 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_0_q_k), .Z(pool_pool_pe_b_peij_1_0_add_notb[1])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_0_add_U8 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_0_q_k), .Z(pool_pool_pe_b_peij_1_0_add_notb[2])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_0_add_U7 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_0_q_k), .Z(pool_pool_pe_b_peij_1_0_add_notb[3])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_0_add_U6 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_0_q_k), .Z(pool_pool_pe_b_peij_1_0_add_notb[4])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_0_add_U5 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_0_q_k), .Z(pool_pool_pe_b_peij_1_0_add_notb[5])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_0_add_U4 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_0_q_k), .Z(pool_pool_pe_b_peij_1_0_add_notb[6])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_0_add_U3 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_0_q_k), .Z(pool_pool_pe_b_peij_1_0_add_notb[7])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_0_add_U2 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_0_q_k), .Z(pool_pool_pe_b_peij_1_0_add_notb[8])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_0_add_U1 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_0_q_k), .Z(pool_pool_pe_b_peij_1_0_add_notb[9])
         );
  INV_X2 pool_pool_pe_b_peij_1_0_add_fai_0_U2 ( .A(
        pool_pool_pe_b_peij_1_0_add_fai_0_n4), .ZN(
        pool_pool_pe_b_peij_1_0_add_cprop[1]) );
  XOR2_X1 pool_pool_pe_b_peij_1_0_add_fai_0_U4 ( .A(pool_pool_pe_b_o_data[121]), .B(pool_pool_pe_b_peij_1_0_add_notb[0]), .Z(
        pool_pool_pe_b_peij_1_0_add_fai_0_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_0_add_fai_0_U3 ( .A(
        pool_pool_pe_b_peij_1_0_q_k), .B(pool_pool_pe_b_peij_1_0_add_fai_0_n5), 
        .Z(pool_pool_pe_b_peij_1_0_d_acc[0]) );
  AOI22_X2 pool_pool_pe_b_peij_1_0_add_fai_0_U1 ( .A1(
        pool_pool_pe_b_peij_1_0_add_notb[0]), .A2(pool_pool_pe_b_o_data[121]), 
        .B1(pool_pool_pe_b_peij_1_0_add_fai_0_n5), .B2(
        pool_pool_pe_b_peij_1_0_q_k), .ZN(pool_pool_pe_b_peij_1_0_add_fai_0_n4) );
  INV_X2 pool_pool_pe_b_peij_1_0_add_fai_1_U2 ( .A(
        pool_pool_pe_b_peij_1_0_add_fai_1_n4), .ZN(
        pool_pool_pe_b_peij_1_0_add_cprop[2]) );
  XOR2_X1 pool_pool_pe_b_peij_1_0_add_fai_1_U4 ( .A(pool_pool_pe_b_o_data[122]), .B(pool_pool_pe_b_peij_1_0_add_notb[1]), .Z(
        pool_pool_pe_b_peij_1_0_add_fai_1_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_0_add_fai_1_U3 ( .A(
        pool_pool_pe_b_peij_1_0_add_cprop[1]), .B(
        pool_pool_pe_b_peij_1_0_add_fai_1_n5), .Z(
        pool_pool_pe_b_peij_1_0_d_acc[1]) );
  AOI22_X2 pool_pool_pe_b_peij_1_0_add_fai_1_U1 ( .A1(
        pool_pool_pe_b_peij_1_0_add_notb[1]), .A2(pool_pool_pe_b_o_data[122]), 
        .B1(pool_pool_pe_b_peij_1_0_add_fai_1_n5), .B2(
        pool_pool_pe_b_peij_1_0_add_cprop[1]), .ZN(
        pool_pool_pe_b_peij_1_0_add_fai_1_n4) );
  INV_X2 pool_pool_pe_b_peij_1_0_add_fai_2_U2 ( .A(
        pool_pool_pe_b_peij_1_0_add_fai_2_n4), .ZN(
        pool_pool_pe_b_peij_1_0_add_cprop[3]) );
  XOR2_X1 pool_pool_pe_b_peij_1_0_add_fai_2_U4 ( .A(pool_pool_pe_b_o_data[123]), .B(pool_pool_pe_b_peij_1_0_add_notb[2]), .Z(
        pool_pool_pe_b_peij_1_0_add_fai_2_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_0_add_fai_2_U3 ( .A(
        pool_pool_pe_b_peij_1_0_add_cprop[2]), .B(
        pool_pool_pe_b_peij_1_0_add_fai_2_n5), .Z(
        pool_pool_pe_b_peij_1_0_d_acc[2]) );
  AOI22_X2 pool_pool_pe_b_peij_1_0_add_fai_2_U1 ( .A1(
        pool_pool_pe_b_peij_1_0_add_notb[2]), .A2(pool_pool_pe_b_o_data[123]), 
        .B1(pool_pool_pe_b_peij_1_0_add_fai_2_n5), .B2(
        pool_pool_pe_b_peij_1_0_add_cprop[2]), .ZN(
        pool_pool_pe_b_peij_1_0_add_fai_2_n4) );
  INV_X2 pool_pool_pe_b_peij_1_0_add_fai_3_U2 ( .A(
        pool_pool_pe_b_peij_1_0_add_fai_3_n4), .ZN(
        pool_pool_pe_b_peij_1_0_add_cprop[4]) );
  XOR2_X1 pool_pool_pe_b_peij_1_0_add_fai_3_U4 ( .A(pool_pool_pe_b_o_data[124]), .B(pool_pool_pe_b_peij_1_0_add_notb[3]), .Z(
        pool_pool_pe_b_peij_1_0_add_fai_3_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_0_add_fai_3_U3 ( .A(
        pool_pool_pe_b_peij_1_0_add_cprop[3]), .B(
        pool_pool_pe_b_peij_1_0_add_fai_3_n5), .Z(
        pool_pool_pe_b_peij_1_0_d_acc[3]) );
  AOI22_X2 pool_pool_pe_b_peij_1_0_add_fai_3_U1 ( .A1(
        pool_pool_pe_b_peij_1_0_add_notb[3]), .A2(pool_pool_pe_b_o_data[124]), 
        .B1(pool_pool_pe_b_peij_1_0_add_fai_3_n5), .B2(
        pool_pool_pe_b_peij_1_0_add_cprop[3]), .ZN(
        pool_pool_pe_b_peij_1_0_add_fai_3_n4) );
  INV_X2 pool_pool_pe_b_peij_1_0_add_fai_4_U2 ( .A(
        pool_pool_pe_b_peij_1_0_add_fai_4_n4), .ZN(
        pool_pool_pe_b_peij_1_0_add_cprop[5]) );
  XOR2_X1 pool_pool_pe_b_peij_1_0_add_fai_4_U4 ( .A(pool_pool_pe_b_o_data[125]), .B(pool_pool_pe_b_peij_1_0_add_notb[4]), .Z(
        pool_pool_pe_b_peij_1_0_add_fai_4_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_0_add_fai_4_U3 ( .A(
        pool_pool_pe_b_peij_1_0_add_cprop[4]), .B(
        pool_pool_pe_b_peij_1_0_add_fai_4_n5), .Z(
        pool_pool_pe_b_peij_1_0_d_acc[4]) );
  AOI22_X2 pool_pool_pe_b_peij_1_0_add_fai_4_U1 ( .A1(
        pool_pool_pe_b_peij_1_0_add_notb[4]), .A2(pool_pool_pe_b_o_data[125]), 
        .B1(pool_pool_pe_b_peij_1_0_add_fai_4_n5), .B2(
        pool_pool_pe_b_peij_1_0_add_cprop[4]), .ZN(
        pool_pool_pe_b_peij_1_0_add_fai_4_n4) );
  INV_X2 pool_pool_pe_b_peij_1_0_add_fai_5_U2 ( .A(
        pool_pool_pe_b_peij_1_0_add_fai_5_n4), .ZN(
        pool_pool_pe_b_peij_1_0_add_cprop[6]) );
  XOR2_X1 pool_pool_pe_b_peij_1_0_add_fai_5_U4 ( .A(pool_pool_pe_b_o_data[126]), .B(pool_pool_pe_b_peij_1_0_add_notb[5]), .Z(
        pool_pool_pe_b_peij_1_0_add_fai_5_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_0_add_fai_5_U3 ( .A(
        pool_pool_pe_b_peij_1_0_add_cprop[5]), .B(
        pool_pool_pe_b_peij_1_0_add_fai_5_n5), .Z(
        pool_pool_pe_b_peij_1_0_d_acc[5]) );
  AOI22_X2 pool_pool_pe_b_peij_1_0_add_fai_5_U1 ( .A1(
        pool_pool_pe_b_peij_1_0_add_notb[5]), .A2(pool_pool_pe_b_o_data[126]), 
        .B1(pool_pool_pe_b_peij_1_0_add_fai_5_n5), .B2(
        pool_pool_pe_b_peij_1_0_add_cprop[5]), .ZN(
        pool_pool_pe_b_peij_1_0_add_fai_5_n4) );
  INV_X2 pool_pool_pe_b_peij_1_0_add_fai_6_U2 ( .A(
        pool_pool_pe_b_peij_1_0_add_fai_6_n4), .ZN(
        pool_pool_pe_b_peij_1_0_add_cprop[7]) );
  XOR2_X1 pool_pool_pe_b_peij_1_0_add_fai_6_U4 ( .A(pool_pool_pe_b_o_data[127]), .B(pool_pool_pe_b_peij_1_0_add_notb[6]), .Z(
        pool_pool_pe_b_peij_1_0_add_fai_6_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_0_add_fai_6_U3 ( .A(
        pool_pool_pe_b_peij_1_0_add_cprop[6]), .B(
        pool_pool_pe_b_peij_1_0_add_fai_6_n5), .Z(
        pool_pool_pe_b_peij_1_0_d_acc[6]) );
  AOI22_X2 pool_pool_pe_b_peij_1_0_add_fai_6_U1 ( .A1(
        pool_pool_pe_b_peij_1_0_add_notb[6]), .A2(pool_pool_pe_b_o_data[127]), 
        .B1(pool_pool_pe_b_peij_1_0_add_fai_6_n5), .B2(
        pool_pool_pe_b_peij_1_0_add_cprop[6]), .ZN(
        pool_pool_pe_b_peij_1_0_add_fai_6_n4) );
  INV_X2 pool_pool_pe_b_peij_1_0_add_fai_7_U2 ( .A(
        pool_pool_pe_b_peij_1_0_add_fai_7_n4), .ZN(
        pool_pool_pe_b_peij_1_0_add_cprop[8]) );
  XOR2_X1 pool_pool_pe_b_peij_1_0_add_fai_7_U4 ( .A(pool_pool_pe_b_o_data[128]), .B(pool_pool_pe_b_peij_1_0_add_notb[7]), .Z(
        pool_pool_pe_b_peij_1_0_add_fai_7_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_0_add_fai_7_U3 ( .A(
        pool_pool_pe_b_peij_1_0_add_cprop[7]), .B(
        pool_pool_pe_b_peij_1_0_add_fai_7_n5), .Z(
        pool_pool_pe_b_peij_1_0_d_acc[7]) );
  AOI22_X2 pool_pool_pe_b_peij_1_0_add_fai_7_U1 ( .A1(
        pool_pool_pe_b_peij_1_0_add_notb[7]), .A2(pool_pool_pe_b_o_data[128]), 
        .B1(pool_pool_pe_b_peij_1_0_add_fai_7_n5), .B2(
        pool_pool_pe_b_peij_1_0_add_cprop[7]), .ZN(
        pool_pool_pe_b_peij_1_0_add_fai_7_n4) );
  INV_X2 pool_pool_pe_b_peij_1_0_add_fai_8_U2 ( .A(
        pool_pool_pe_b_peij_1_0_add_fai_8_n4), .ZN(
        pool_pool_pe_b_peij_1_0_add_cprop[9]) );
  XOR2_X1 pool_pool_pe_b_peij_1_0_add_fai_8_U4 ( .A(pool_pool_pe_b_o_data[129]), .B(pool_pool_pe_b_peij_1_0_add_notb[8]), .Z(
        pool_pool_pe_b_peij_1_0_add_fai_8_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_0_add_fai_8_U3 ( .A(
        pool_pool_pe_b_peij_1_0_add_cprop[8]), .B(
        pool_pool_pe_b_peij_1_0_add_fai_8_n5), .Z(
        pool_pool_pe_b_peij_1_0_d_acc[8]) );
  AOI22_X2 pool_pool_pe_b_peij_1_0_add_fai_8_U1 ( .A1(
        pool_pool_pe_b_peij_1_0_add_notb[8]), .A2(pool_pool_pe_b_o_data[129]), 
        .B1(pool_pool_pe_b_peij_1_0_add_fai_8_n5), .B2(
        pool_pool_pe_b_peij_1_0_add_cprop[8]), .ZN(
        pool_pool_pe_b_peij_1_0_add_fai_8_n4) );
  INV_X2 pool_pool_pe_b_peij_1_0_add_fai_9_U2 ( .A(
        pool_pool_pe_b_peij_1_0_add_fai_9_n4), .ZN(
        pool_pool_pe_b_peij_1_0_add_cprop[10]) );
  XOR2_X1 pool_pool_pe_b_peij_1_0_add_fai_9_U4 ( .A(pool_pool_pe_b_o_data[130]), .B(pool_pool_pe_b_peij_1_0_add_notb[9]), .Z(
        pool_pool_pe_b_peij_1_0_add_fai_9_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_0_add_fai_9_U3 ( .A(
        pool_pool_pe_b_peij_1_0_add_cprop[9]), .B(
        pool_pool_pe_b_peij_1_0_add_fai_9_n5), .Z(
        pool_pool_pe_b_peij_1_0_d_acc[9]) );
  AOI22_X2 pool_pool_pe_b_peij_1_0_add_fai_9_U1 ( .A1(
        pool_pool_pe_b_peij_1_0_add_notb[9]), .A2(pool_pool_pe_b_o_data[130]), 
        .B1(pool_pool_pe_b_peij_1_0_add_fai_9_n5), .B2(
        pool_pool_pe_b_peij_1_0_add_cprop[9]), .ZN(
        pool_pool_pe_b_peij_1_0_add_fai_9_n4) );
  INV_X2 pool_pool_pe_b_peij_1_0_add_fai_10_U2 ( .A(
        pool_pool_pe_b_peij_1_0_add_fai_10_n4), .ZN(
        pool_pool_pe_b_peij_1_0_add_c_out) );
  XOR2_X1 pool_pool_pe_b_peij_1_0_add_fai_10_U4 ( .A(
        pool_pool_pe_b_o_data[131]), .B(pool_pool_pe_b_peij_1_0_add_notb[10]), 
        .Z(pool_pool_pe_b_peij_1_0_add_fai_10_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_0_add_fai_10_U3 ( .A(
        pool_pool_pe_b_peij_1_0_add_cprop[10]), .B(
        pool_pool_pe_b_peij_1_0_add_fai_10_n5), .Z(
        pool_pool_pe_b_peij_1_0_d_acc[10]) );
  AOI22_X2 pool_pool_pe_b_peij_1_0_add_fai_10_U1 ( .A1(
        pool_pool_pe_b_peij_1_0_add_notb[10]), .A2(pool_pool_pe_b_o_data[131]), 
        .B1(pool_pool_pe_b_peij_1_0_add_fai_10_n5), .B2(
        pool_pool_pe_b_peij_1_0_add_cprop[10]), .ZN(
        pool_pool_pe_b_peij_1_0_add_fai_10_n4) );
  INV_X2 pool_pool_pe_b_peij_1_1_U21 ( .A(pool_sync_clr), .ZN(
        pool_pool_pe_b_peij_1_1_n14) );
  INV_X1 pool_pool_pe_b_peij_1_1_U18 ( .A(pool_pool_pe_b_n1), .ZN(
        pool_pool_pe_b_peij_1_1_n12) );
  AND2_X1 pool_pool_pe_b_peij_1_1_U13 ( .A1(pool_pool_pe_b_peij_1_1_d_acc[0]), 
        .A2(pool_pool_pe_b_peij_1_1_n14), .ZN(pool_pool_pe_b_peij_1_1_n11) );
  AND2_X1 pool_pool_pe_b_peij_1_1_U12 ( .A1(pool_pool_pe_b_peij_1_1_d_acc[1]), 
        .A2(pool_pool_pe_b_peij_1_1_n14), .ZN(pool_pool_pe_b_peij_1_1_n10) );
  AND2_X1 pool_pool_pe_b_peij_1_1_U11 ( .A1(pool_pool_pe_b_peij_1_1_d_acc[2]), 
        .A2(pool_pool_pe_b_peij_1_1_n14), .ZN(pool_pool_pe_b_peij_1_1_n9) );
  AND2_X1 pool_pool_pe_b_peij_1_1_U10 ( .A1(pool_pool_pe_b_peij_1_1_d_acc[3]), 
        .A2(pool_pool_pe_b_peij_1_1_n14), .ZN(pool_pool_pe_b_peij_1_1_n8) );
  AND2_X1 pool_pool_pe_b_peij_1_1_U9 ( .A1(pool_pool_pe_b_peij_1_1_d_acc[4]), 
        .A2(pool_pool_pe_b_peij_1_1_n14), .ZN(pool_pool_pe_b_peij_1_1_n7) );
  AND2_X1 pool_pool_pe_b_peij_1_1_U8 ( .A1(pool_pool_pe_b_peij_1_1_d_acc[5]), 
        .A2(pool_pool_pe_b_peij_1_1_n14), .ZN(pool_pool_pe_b_peij_1_1_n6) );
  AND2_X1 pool_pool_pe_b_peij_1_1_U7 ( .A1(pool_pool_pe_b_peij_1_1_d_acc[6]), 
        .A2(pool_pool_pe_b_peij_1_1_n14), .ZN(pool_pool_pe_b_peij_1_1_n5) );
  AND2_X1 pool_pool_pe_b_peij_1_1_U6 ( .A1(pool_pool_pe_b_peij_1_1_d_acc[7]), 
        .A2(pool_pool_pe_b_peij_1_1_n14), .ZN(pool_pool_pe_b_peij_1_1_n4) );
  AND2_X1 pool_pool_pe_b_peij_1_1_U5 ( .A1(pool_pool_pe_b_peij_1_1_d_acc[8]), 
        .A2(pool_pool_pe_b_peij_1_1_n14), .ZN(pool_pool_pe_b_peij_1_1_n3) );
  AND2_X1 pool_pool_pe_b_peij_1_1_U4 ( .A1(pool_pool_pe_b_peij_1_1_d_acc[9]), 
        .A2(pool_pool_pe_b_peij_1_1_n14), .ZN(pool_pool_pe_b_peij_1_1_n2) );
  AND2_X1 pool_pool_pe_b_peij_1_1_U3 ( .A1(pool_pool_pe_b_peij_1_1_d_acc[10]), 
        .A2(pool_pool_pe_b_peij_1_1_n14), .ZN(pool_pool_pe_b_peij_1_1_n1) );
  DFFR_X1 pool_pool_pe_b_peij_1_1_q_acc_reg_10_ ( .D(
        pool_pool_pe_b_peij_1_1_n1), .CK(pool_pool_pe_b_peij_1_1_gck), .RN(
        pool_pool_pe_b_peij_1_1_n12), .Q(pool_pool_pe_b_o_data[120]) );
  DFFR_X1 pool_pool_pe_b_peij_1_1_q_acc_reg_9_ ( .D(pool_pool_pe_b_peij_1_1_n2), .CK(pool_pool_pe_b_peij_1_1_gck), .RN(pool_pool_pe_b_peij_1_1_n12), .Q(
        pool_pool_pe_b_o_data[119]) );
  DFFR_X1 pool_pool_pe_b_peij_1_1_q_acc_reg_8_ ( .D(pool_pool_pe_b_peij_1_1_n3), .CK(pool_pool_pe_b_peij_1_1_gck), .RN(pool_pool_pe_b_peij_1_1_n12), .Q(
        pool_pool_pe_b_o_data[118]) );
  DFFR_X1 pool_pool_pe_b_peij_1_1_q_acc_reg_7_ ( .D(pool_pool_pe_b_peij_1_1_n4), .CK(pool_pool_pe_b_peij_1_1_gck), .RN(pool_pool_pe_b_peij_1_1_n12), .Q(
        pool_pool_pe_b_o_data[117]) );
  DFFR_X1 pool_pool_pe_b_peij_1_1_q_acc_reg_6_ ( .D(pool_pool_pe_b_peij_1_1_n5), .CK(pool_pool_pe_b_peij_1_1_gck), .RN(pool_pool_pe_b_peij_1_1_n12), .Q(
        pool_pool_pe_b_o_data[116]) );
  DFFR_X1 pool_pool_pe_b_peij_1_1_q_acc_reg_5_ ( .D(pool_pool_pe_b_peij_1_1_n6), .CK(pool_pool_pe_b_peij_1_1_gck), .RN(pool_pool_pe_b_peij_1_1_n12), .Q(
        pool_pool_pe_b_o_data[115]) );
  DFFR_X1 pool_pool_pe_b_peij_1_1_q_acc_reg_4_ ( .D(pool_pool_pe_b_peij_1_1_n7), .CK(pool_pool_pe_b_peij_1_1_gck), .RN(pool_pool_pe_b_peij_1_1_n12), .Q(
        pool_pool_pe_b_o_data[114]) );
  DFFR_X1 pool_pool_pe_b_peij_1_1_q_acc_reg_3_ ( .D(pool_pool_pe_b_peij_1_1_n8), .CK(pool_pool_pe_b_peij_1_1_gck), .RN(pool_pool_pe_b_peij_1_1_n12), .Q(
        pool_pool_pe_b_o_data[113]) );
  DFFR_X1 pool_pool_pe_b_peij_1_1_q_acc_reg_2_ ( .D(pool_pool_pe_b_peij_1_1_n9), .CK(pool_pool_pe_b_peij_1_1_gck), .RN(pool_pool_pe_b_peij_1_1_n12), .Q(
        pool_pool_pe_b_o_data[112]) );
  DFFR_X1 pool_pool_pe_b_peij_1_1_q_acc_reg_1_ ( .D(
        pool_pool_pe_b_peij_1_1_n10), .CK(pool_pool_pe_b_peij_1_1_gck), .RN(
        pool_pool_pe_b_peij_1_1_n12), .Q(pool_pool_pe_b_o_data[111]) );
  DFFR_X1 pool_pool_pe_b_peij_1_1_q_acc_reg_0_ ( .D(
        pool_pool_pe_b_peij_1_1_n11), .CK(pool_pool_pe_b_peij_1_1_gck), .RN(
        pool_pool_pe_b_peij_1_1_n12), .Q(pool_pool_pe_b_o_data[110]) );
  AND3_X2 pool_pool_pe_b_peij_1_1_U20 ( .A1(pool_pool_pe_b_int_pe_en[10]), 
        .A2(clk), .A3(1'b1), .ZN(pool_pool_pe_b_peij_1_1_gck) );
  SDFFR_X1 pool_pool_pe_b_peij_1_1_q_k_reg ( .D(1'b0), .SI(
        pool_pool_pe_b_peij_1_1_n14), .SE(1'b0), .CK(
        pool_pool_pe_b_peij_1_1_gck), .RN(pool_pool_pe_b_peij_1_1_n12), .Q(
        pool_pool_pe_b_peij_1_1_q_k) );
  XOR2_X1 pool_pool_pe_b_peij_1_1_add_U11 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_1_q_k), .Z(pool_pool_pe_b_peij_1_1_add_notb[0])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_1_add_U10 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_1_q_k), .Z(pool_pool_pe_b_peij_1_1_add_notb[10])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_1_add_U9 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_1_q_k), .Z(pool_pool_pe_b_peij_1_1_add_notb[1])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_1_add_U8 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_1_q_k), .Z(pool_pool_pe_b_peij_1_1_add_notb[2])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_1_add_U7 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_1_q_k), .Z(pool_pool_pe_b_peij_1_1_add_notb[3])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_1_add_U6 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_1_q_k), .Z(pool_pool_pe_b_peij_1_1_add_notb[4])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_1_add_U5 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_1_q_k), .Z(pool_pool_pe_b_peij_1_1_add_notb[5])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_1_add_U4 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_1_q_k), .Z(pool_pool_pe_b_peij_1_1_add_notb[6])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_1_add_U3 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_1_q_k), .Z(pool_pool_pe_b_peij_1_1_add_notb[7])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_1_add_U2 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_1_q_k), .Z(pool_pool_pe_b_peij_1_1_add_notb[8])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_1_add_U1 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_1_q_k), .Z(pool_pool_pe_b_peij_1_1_add_notb[9])
         );
  INV_X2 pool_pool_pe_b_peij_1_1_add_fai_0_U2 ( .A(
        pool_pool_pe_b_peij_1_1_add_fai_0_n4), .ZN(
        pool_pool_pe_b_peij_1_1_add_cprop[1]) );
  XOR2_X1 pool_pool_pe_b_peij_1_1_add_fai_0_U4 ( .A(pool_pool_pe_b_o_data[110]), .B(pool_pool_pe_b_peij_1_1_add_notb[0]), .Z(
        pool_pool_pe_b_peij_1_1_add_fai_0_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_1_add_fai_0_U3 ( .A(
        pool_pool_pe_b_peij_1_1_q_k), .B(pool_pool_pe_b_peij_1_1_add_fai_0_n5), 
        .Z(pool_pool_pe_b_peij_1_1_d_acc[0]) );
  AOI22_X2 pool_pool_pe_b_peij_1_1_add_fai_0_U1 ( .A1(
        pool_pool_pe_b_peij_1_1_add_notb[0]), .A2(pool_pool_pe_b_o_data[110]), 
        .B1(pool_pool_pe_b_peij_1_1_add_fai_0_n5), .B2(
        pool_pool_pe_b_peij_1_1_q_k), .ZN(pool_pool_pe_b_peij_1_1_add_fai_0_n4) );
  INV_X2 pool_pool_pe_b_peij_1_1_add_fai_1_U2 ( .A(
        pool_pool_pe_b_peij_1_1_add_fai_1_n4), .ZN(
        pool_pool_pe_b_peij_1_1_add_cprop[2]) );
  XOR2_X1 pool_pool_pe_b_peij_1_1_add_fai_1_U4 ( .A(pool_pool_pe_b_o_data[111]), .B(pool_pool_pe_b_peij_1_1_add_notb[1]), .Z(
        pool_pool_pe_b_peij_1_1_add_fai_1_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_1_add_fai_1_U3 ( .A(
        pool_pool_pe_b_peij_1_1_add_cprop[1]), .B(
        pool_pool_pe_b_peij_1_1_add_fai_1_n5), .Z(
        pool_pool_pe_b_peij_1_1_d_acc[1]) );
  AOI22_X2 pool_pool_pe_b_peij_1_1_add_fai_1_U1 ( .A1(
        pool_pool_pe_b_peij_1_1_add_notb[1]), .A2(pool_pool_pe_b_o_data[111]), 
        .B1(pool_pool_pe_b_peij_1_1_add_fai_1_n5), .B2(
        pool_pool_pe_b_peij_1_1_add_cprop[1]), .ZN(
        pool_pool_pe_b_peij_1_1_add_fai_1_n4) );
  INV_X2 pool_pool_pe_b_peij_1_1_add_fai_2_U2 ( .A(
        pool_pool_pe_b_peij_1_1_add_fai_2_n4), .ZN(
        pool_pool_pe_b_peij_1_1_add_cprop[3]) );
  XOR2_X1 pool_pool_pe_b_peij_1_1_add_fai_2_U4 ( .A(pool_pool_pe_b_o_data[112]), .B(pool_pool_pe_b_peij_1_1_add_notb[2]), .Z(
        pool_pool_pe_b_peij_1_1_add_fai_2_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_1_add_fai_2_U3 ( .A(
        pool_pool_pe_b_peij_1_1_add_cprop[2]), .B(
        pool_pool_pe_b_peij_1_1_add_fai_2_n5), .Z(
        pool_pool_pe_b_peij_1_1_d_acc[2]) );
  AOI22_X2 pool_pool_pe_b_peij_1_1_add_fai_2_U1 ( .A1(
        pool_pool_pe_b_peij_1_1_add_notb[2]), .A2(pool_pool_pe_b_o_data[112]), 
        .B1(pool_pool_pe_b_peij_1_1_add_fai_2_n5), .B2(
        pool_pool_pe_b_peij_1_1_add_cprop[2]), .ZN(
        pool_pool_pe_b_peij_1_1_add_fai_2_n4) );
  INV_X2 pool_pool_pe_b_peij_1_1_add_fai_3_U2 ( .A(
        pool_pool_pe_b_peij_1_1_add_fai_3_n4), .ZN(
        pool_pool_pe_b_peij_1_1_add_cprop[4]) );
  XOR2_X1 pool_pool_pe_b_peij_1_1_add_fai_3_U4 ( .A(pool_pool_pe_b_o_data[113]), .B(pool_pool_pe_b_peij_1_1_add_notb[3]), .Z(
        pool_pool_pe_b_peij_1_1_add_fai_3_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_1_add_fai_3_U3 ( .A(
        pool_pool_pe_b_peij_1_1_add_cprop[3]), .B(
        pool_pool_pe_b_peij_1_1_add_fai_3_n5), .Z(
        pool_pool_pe_b_peij_1_1_d_acc[3]) );
  AOI22_X2 pool_pool_pe_b_peij_1_1_add_fai_3_U1 ( .A1(
        pool_pool_pe_b_peij_1_1_add_notb[3]), .A2(pool_pool_pe_b_o_data[113]), 
        .B1(pool_pool_pe_b_peij_1_1_add_fai_3_n5), .B2(
        pool_pool_pe_b_peij_1_1_add_cprop[3]), .ZN(
        pool_pool_pe_b_peij_1_1_add_fai_3_n4) );
  INV_X2 pool_pool_pe_b_peij_1_1_add_fai_4_U2 ( .A(
        pool_pool_pe_b_peij_1_1_add_fai_4_n4), .ZN(
        pool_pool_pe_b_peij_1_1_add_cprop[5]) );
  XOR2_X1 pool_pool_pe_b_peij_1_1_add_fai_4_U4 ( .A(pool_pool_pe_b_o_data[114]), .B(pool_pool_pe_b_peij_1_1_add_notb[4]), .Z(
        pool_pool_pe_b_peij_1_1_add_fai_4_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_1_add_fai_4_U3 ( .A(
        pool_pool_pe_b_peij_1_1_add_cprop[4]), .B(
        pool_pool_pe_b_peij_1_1_add_fai_4_n5), .Z(
        pool_pool_pe_b_peij_1_1_d_acc[4]) );
  AOI22_X2 pool_pool_pe_b_peij_1_1_add_fai_4_U1 ( .A1(
        pool_pool_pe_b_peij_1_1_add_notb[4]), .A2(pool_pool_pe_b_o_data[114]), 
        .B1(pool_pool_pe_b_peij_1_1_add_fai_4_n5), .B2(
        pool_pool_pe_b_peij_1_1_add_cprop[4]), .ZN(
        pool_pool_pe_b_peij_1_1_add_fai_4_n4) );
  INV_X2 pool_pool_pe_b_peij_1_1_add_fai_5_U2 ( .A(
        pool_pool_pe_b_peij_1_1_add_fai_5_n4), .ZN(
        pool_pool_pe_b_peij_1_1_add_cprop[6]) );
  XOR2_X1 pool_pool_pe_b_peij_1_1_add_fai_5_U4 ( .A(pool_pool_pe_b_o_data[115]), .B(pool_pool_pe_b_peij_1_1_add_notb[5]), .Z(
        pool_pool_pe_b_peij_1_1_add_fai_5_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_1_add_fai_5_U3 ( .A(
        pool_pool_pe_b_peij_1_1_add_cprop[5]), .B(
        pool_pool_pe_b_peij_1_1_add_fai_5_n5), .Z(
        pool_pool_pe_b_peij_1_1_d_acc[5]) );
  AOI22_X2 pool_pool_pe_b_peij_1_1_add_fai_5_U1 ( .A1(
        pool_pool_pe_b_peij_1_1_add_notb[5]), .A2(pool_pool_pe_b_o_data[115]), 
        .B1(pool_pool_pe_b_peij_1_1_add_fai_5_n5), .B2(
        pool_pool_pe_b_peij_1_1_add_cprop[5]), .ZN(
        pool_pool_pe_b_peij_1_1_add_fai_5_n4) );
  INV_X2 pool_pool_pe_b_peij_1_1_add_fai_6_U2 ( .A(
        pool_pool_pe_b_peij_1_1_add_fai_6_n4), .ZN(
        pool_pool_pe_b_peij_1_1_add_cprop[7]) );
  XOR2_X1 pool_pool_pe_b_peij_1_1_add_fai_6_U4 ( .A(pool_pool_pe_b_o_data[116]), .B(pool_pool_pe_b_peij_1_1_add_notb[6]), .Z(
        pool_pool_pe_b_peij_1_1_add_fai_6_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_1_add_fai_6_U3 ( .A(
        pool_pool_pe_b_peij_1_1_add_cprop[6]), .B(
        pool_pool_pe_b_peij_1_1_add_fai_6_n5), .Z(
        pool_pool_pe_b_peij_1_1_d_acc[6]) );
  AOI22_X2 pool_pool_pe_b_peij_1_1_add_fai_6_U1 ( .A1(
        pool_pool_pe_b_peij_1_1_add_notb[6]), .A2(pool_pool_pe_b_o_data[116]), 
        .B1(pool_pool_pe_b_peij_1_1_add_fai_6_n5), .B2(
        pool_pool_pe_b_peij_1_1_add_cprop[6]), .ZN(
        pool_pool_pe_b_peij_1_1_add_fai_6_n4) );
  INV_X2 pool_pool_pe_b_peij_1_1_add_fai_7_U2 ( .A(
        pool_pool_pe_b_peij_1_1_add_fai_7_n4), .ZN(
        pool_pool_pe_b_peij_1_1_add_cprop[8]) );
  XOR2_X1 pool_pool_pe_b_peij_1_1_add_fai_7_U4 ( .A(pool_pool_pe_b_o_data[117]), .B(pool_pool_pe_b_peij_1_1_add_notb[7]), .Z(
        pool_pool_pe_b_peij_1_1_add_fai_7_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_1_add_fai_7_U3 ( .A(
        pool_pool_pe_b_peij_1_1_add_cprop[7]), .B(
        pool_pool_pe_b_peij_1_1_add_fai_7_n5), .Z(
        pool_pool_pe_b_peij_1_1_d_acc[7]) );
  AOI22_X2 pool_pool_pe_b_peij_1_1_add_fai_7_U1 ( .A1(
        pool_pool_pe_b_peij_1_1_add_notb[7]), .A2(pool_pool_pe_b_o_data[117]), 
        .B1(pool_pool_pe_b_peij_1_1_add_fai_7_n5), .B2(
        pool_pool_pe_b_peij_1_1_add_cprop[7]), .ZN(
        pool_pool_pe_b_peij_1_1_add_fai_7_n4) );
  INV_X2 pool_pool_pe_b_peij_1_1_add_fai_8_U2 ( .A(
        pool_pool_pe_b_peij_1_1_add_fai_8_n4), .ZN(
        pool_pool_pe_b_peij_1_1_add_cprop[9]) );
  XOR2_X1 pool_pool_pe_b_peij_1_1_add_fai_8_U4 ( .A(pool_pool_pe_b_o_data[118]), .B(pool_pool_pe_b_peij_1_1_add_notb[8]), .Z(
        pool_pool_pe_b_peij_1_1_add_fai_8_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_1_add_fai_8_U3 ( .A(
        pool_pool_pe_b_peij_1_1_add_cprop[8]), .B(
        pool_pool_pe_b_peij_1_1_add_fai_8_n5), .Z(
        pool_pool_pe_b_peij_1_1_d_acc[8]) );
  AOI22_X2 pool_pool_pe_b_peij_1_1_add_fai_8_U1 ( .A1(
        pool_pool_pe_b_peij_1_1_add_notb[8]), .A2(pool_pool_pe_b_o_data[118]), 
        .B1(pool_pool_pe_b_peij_1_1_add_fai_8_n5), .B2(
        pool_pool_pe_b_peij_1_1_add_cprop[8]), .ZN(
        pool_pool_pe_b_peij_1_1_add_fai_8_n4) );
  INV_X2 pool_pool_pe_b_peij_1_1_add_fai_9_U2 ( .A(
        pool_pool_pe_b_peij_1_1_add_fai_9_n4), .ZN(
        pool_pool_pe_b_peij_1_1_add_cprop[10]) );
  XOR2_X1 pool_pool_pe_b_peij_1_1_add_fai_9_U4 ( .A(pool_pool_pe_b_o_data[119]), .B(pool_pool_pe_b_peij_1_1_add_notb[9]), .Z(
        pool_pool_pe_b_peij_1_1_add_fai_9_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_1_add_fai_9_U3 ( .A(
        pool_pool_pe_b_peij_1_1_add_cprop[9]), .B(
        pool_pool_pe_b_peij_1_1_add_fai_9_n5), .Z(
        pool_pool_pe_b_peij_1_1_d_acc[9]) );
  AOI22_X2 pool_pool_pe_b_peij_1_1_add_fai_9_U1 ( .A1(
        pool_pool_pe_b_peij_1_1_add_notb[9]), .A2(pool_pool_pe_b_o_data[119]), 
        .B1(pool_pool_pe_b_peij_1_1_add_fai_9_n5), .B2(
        pool_pool_pe_b_peij_1_1_add_cprop[9]), .ZN(
        pool_pool_pe_b_peij_1_1_add_fai_9_n4) );
  INV_X2 pool_pool_pe_b_peij_1_1_add_fai_10_U2 ( .A(
        pool_pool_pe_b_peij_1_1_add_fai_10_n4), .ZN(
        pool_pool_pe_b_peij_1_1_add_c_out) );
  XOR2_X1 pool_pool_pe_b_peij_1_1_add_fai_10_U4 ( .A(
        pool_pool_pe_b_o_data[120]), .B(pool_pool_pe_b_peij_1_1_add_notb[10]), 
        .Z(pool_pool_pe_b_peij_1_1_add_fai_10_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_1_add_fai_10_U3 ( .A(
        pool_pool_pe_b_peij_1_1_add_cprop[10]), .B(
        pool_pool_pe_b_peij_1_1_add_fai_10_n5), .Z(
        pool_pool_pe_b_peij_1_1_d_acc[10]) );
  AOI22_X2 pool_pool_pe_b_peij_1_1_add_fai_10_U1 ( .A1(
        pool_pool_pe_b_peij_1_1_add_notb[10]), .A2(pool_pool_pe_b_o_data[120]), 
        .B1(pool_pool_pe_b_peij_1_1_add_fai_10_n5), .B2(
        pool_pool_pe_b_peij_1_1_add_cprop[10]), .ZN(
        pool_pool_pe_b_peij_1_1_add_fai_10_n4) );
  INV_X2 pool_pool_pe_b_peij_1_2_U21 ( .A(pool_sync_clr), .ZN(
        pool_pool_pe_b_peij_1_2_n14) );
  INV_X1 pool_pool_pe_b_peij_1_2_U18 ( .A(pool_pool_pe_b_n1), .ZN(
        pool_pool_pe_b_peij_1_2_n12) );
  AND2_X1 pool_pool_pe_b_peij_1_2_U13 ( .A1(pool_pool_pe_b_peij_1_2_d_acc[0]), 
        .A2(pool_pool_pe_b_peij_1_2_n14), .ZN(pool_pool_pe_b_peij_1_2_n11) );
  AND2_X1 pool_pool_pe_b_peij_1_2_U12 ( .A1(pool_pool_pe_b_peij_1_2_d_acc[1]), 
        .A2(pool_pool_pe_b_peij_1_2_n14), .ZN(pool_pool_pe_b_peij_1_2_n10) );
  AND2_X1 pool_pool_pe_b_peij_1_2_U11 ( .A1(pool_pool_pe_b_peij_1_2_d_acc[2]), 
        .A2(pool_pool_pe_b_peij_1_2_n14), .ZN(pool_pool_pe_b_peij_1_2_n9) );
  AND2_X1 pool_pool_pe_b_peij_1_2_U10 ( .A1(pool_pool_pe_b_peij_1_2_d_acc[3]), 
        .A2(pool_pool_pe_b_peij_1_2_n14), .ZN(pool_pool_pe_b_peij_1_2_n8) );
  AND2_X1 pool_pool_pe_b_peij_1_2_U9 ( .A1(pool_pool_pe_b_peij_1_2_d_acc[4]), 
        .A2(pool_pool_pe_b_peij_1_2_n14), .ZN(pool_pool_pe_b_peij_1_2_n7) );
  AND2_X1 pool_pool_pe_b_peij_1_2_U8 ( .A1(pool_pool_pe_b_peij_1_2_d_acc[5]), 
        .A2(pool_pool_pe_b_peij_1_2_n14), .ZN(pool_pool_pe_b_peij_1_2_n6) );
  AND2_X1 pool_pool_pe_b_peij_1_2_U7 ( .A1(pool_pool_pe_b_peij_1_2_d_acc[6]), 
        .A2(pool_pool_pe_b_peij_1_2_n14), .ZN(pool_pool_pe_b_peij_1_2_n5) );
  AND2_X1 pool_pool_pe_b_peij_1_2_U6 ( .A1(pool_pool_pe_b_peij_1_2_d_acc[7]), 
        .A2(pool_pool_pe_b_peij_1_2_n14), .ZN(pool_pool_pe_b_peij_1_2_n4) );
  AND2_X1 pool_pool_pe_b_peij_1_2_U5 ( .A1(pool_pool_pe_b_peij_1_2_d_acc[8]), 
        .A2(pool_pool_pe_b_peij_1_2_n14), .ZN(pool_pool_pe_b_peij_1_2_n3) );
  AND2_X1 pool_pool_pe_b_peij_1_2_U4 ( .A1(pool_pool_pe_b_peij_1_2_d_acc[9]), 
        .A2(pool_pool_pe_b_peij_1_2_n14), .ZN(pool_pool_pe_b_peij_1_2_n2) );
  AND2_X1 pool_pool_pe_b_peij_1_2_U3 ( .A1(pool_pool_pe_b_peij_1_2_d_acc[10]), 
        .A2(pool_pool_pe_b_peij_1_2_n14), .ZN(pool_pool_pe_b_peij_1_2_n1) );
  DFFR_X1 pool_pool_pe_b_peij_1_2_q_acc_reg_10_ ( .D(
        pool_pool_pe_b_peij_1_2_n1), .CK(pool_pool_pe_b_peij_1_2_gck), .RN(
        pool_pool_pe_b_peij_1_2_n12), .Q(pool_pool_pe_b_o_data[109]) );
  DFFR_X1 pool_pool_pe_b_peij_1_2_q_acc_reg_9_ ( .D(pool_pool_pe_b_peij_1_2_n2), .CK(pool_pool_pe_b_peij_1_2_gck), .RN(pool_pool_pe_b_peij_1_2_n12), .Q(
        pool_pool_pe_b_o_data[108]) );
  DFFR_X1 pool_pool_pe_b_peij_1_2_q_acc_reg_8_ ( .D(pool_pool_pe_b_peij_1_2_n3), .CK(pool_pool_pe_b_peij_1_2_gck), .RN(pool_pool_pe_b_peij_1_2_n12), .Q(
        pool_pool_pe_b_o_data[107]) );
  DFFR_X1 pool_pool_pe_b_peij_1_2_q_acc_reg_7_ ( .D(pool_pool_pe_b_peij_1_2_n4), .CK(pool_pool_pe_b_peij_1_2_gck), .RN(pool_pool_pe_b_peij_1_2_n12), .Q(
        pool_pool_pe_b_o_data[106]) );
  DFFR_X1 pool_pool_pe_b_peij_1_2_q_acc_reg_6_ ( .D(pool_pool_pe_b_peij_1_2_n5), .CK(pool_pool_pe_b_peij_1_2_gck), .RN(pool_pool_pe_b_peij_1_2_n12), .Q(
        pool_pool_pe_b_o_data[105]) );
  DFFR_X1 pool_pool_pe_b_peij_1_2_q_acc_reg_5_ ( .D(pool_pool_pe_b_peij_1_2_n6), .CK(pool_pool_pe_b_peij_1_2_gck), .RN(pool_pool_pe_b_peij_1_2_n12), .Q(
        pool_pool_pe_b_o_data[104]) );
  DFFR_X1 pool_pool_pe_b_peij_1_2_q_acc_reg_4_ ( .D(pool_pool_pe_b_peij_1_2_n7), .CK(pool_pool_pe_b_peij_1_2_gck), .RN(pool_pool_pe_b_peij_1_2_n12), .Q(
        pool_pool_pe_b_o_data[103]) );
  DFFR_X1 pool_pool_pe_b_peij_1_2_q_acc_reg_3_ ( .D(pool_pool_pe_b_peij_1_2_n8), .CK(pool_pool_pe_b_peij_1_2_gck), .RN(pool_pool_pe_b_peij_1_2_n12), .Q(
        pool_pool_pe_b_o_data[102]) );
  DFFR_X1 pool_pool_pe_b_peij_1_2_q_acc_reg_2_ ( .D(pool_pool_pe_b_peij_1_2_n9), .CK(pool_pool_pe_b_peij_1_2_gck), .RN(pool_pool_pe_b_peij_1_2_n12), .Q(
        pool_pool_pe_b_o_data[101]) );
  DFFR_X1 pool_pool_pe_b_peij_1_2_q_acc_reg_1_ ( .D(
        pool_pool_pe_b_peij_1_2_n10), .CK(pool_pool_pe_b_peij_1_2_gck), .RN(
        pool_pool_pe_b_peij_1_2_n12), .Q(pool_pool_pe_b_o_data[100]) );
  DFFR_X1 pool_pool_pe_b_peij_1_2_q_acc_reg_0_ ( .D(
        pool_pool_pe_b_peij_1_2_n11), .CK(pool_pool_pe_b_peij_1_2_gck), .RN(
        pool_pool_pe_b_peij_1_2_n12), .Q(pool_pool_pe_b_o_data[99]) );
  AND3_X2 pool_pool_pe_b_peij_1_2_U20 ( .A1(pool_pool_pe_b_int_pe_en[9]), .A2(
        clk), .A3(1'b1), .ZN(pool_pool_pe_b_peij_1_2_gck) );
  SDFFR_X1 pool_pool_pe_b_peij_1_2_q_k_reg ( .D(1'b0), .SI(
        pool_pool_pe_b_peij_1_2_n14), .SE(1'b0), .CK(
        pool_pool_pe_b_peij_1_2_gck), .RN(pool_pool_pe_b_peij_1_2_n12), .Q(
        pool_pool_pe_b_peij_1_2_q_k) );
  XOR2_X1 pool_pool_pe_b_peij_1_2_add_U11 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_2_q_k), .Z(pool_pool_pe_b_peij_1_2_add_notb[0])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_2_add_U10 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_2_q_k), .Z(pool_pool_pe_b_peij_1_2_add_notb[10])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_2_add_U9 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_2_q_k), .Z(pool_pool_pe_b_peij_1_2_add_notb[1])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_2_add_U8 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_2_q_k), .Z(pool_pool_pe_b_peij_1_2_add_notb[2])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_2_add_U7 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_2_q_k), .Z(pool_pool_pe_b_peij_1_2_add_notb[3])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_2_add_U6 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_2_q_k), .Z(pool_pool_pe_b_peij_1_2_add_notb[4])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_2_add_U5 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_2_q_k), .Z(pool_pool_pe_b_peij_1_2_add_notb[5])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_2_add_U4 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_2_q_k), .Z(pool_pool_pe_b_peij_1_2_add_notb[6])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_2_add_U3 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_2_q_k), .Z(pool_pool_pe_b_peij_1_2_add_notb[7])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_2_add_U2 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_2_q_k), .Z(pool_pool_pe_b_peij_1_2_add_notb[8])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_2_add_U1 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_2_q_k), .Z(pool_pool_pe_b_peij_1_2_add_notb[9])
         );
  INV_X2 pool_pool_pe_b_peij_1_2_add_fai_0_U2 ( .A(
        pool_pool_pe_b_peij_1_2_add_fai_0_n4), .ZN(
        pool_pool_pe_b_peij_1_2_add_cprop[1]) );
  XOR2_X1 pool_pool_pe_b_peij_1_2_add_fai_0_U4 ( .A(pool_pool_pe_b_o_data[99]), 
        .B(pool_pool_pe_b_peij_1_2_add_notb[0]), .Z(
        pool_pool_pe_b_peij_1_2_add_fai_0_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_2_add_fai_0_U3 ( .A(
        pool_pool_pe_b_peij_1_2_q_k), .B(pool_pool_pe_b_peij_1_2_add_fai_0_n5), 
        .Z(pool_pool_pe_b_peij_1_2_d_acc[0]) );
  AOI22_X2 pool_pool_pe_b_peij_1_2_add_fai_0_U1 ( .A1(
        pool_pool_pe_b_peij_1_2_add_notb[0]), .A2(pool_pool_pe_b_o_data[99]), 
        .B1(pool_pool_pe_b_peij_1_2_add_fai_0_n5), .B2(
        pool_pool_pe_b_peij_1_2_q_k), .ZN(pool_pool_pe_b_peij_1_2_add_fai_0_n4) );
  INV_X2 pool_pool_pe_b_peij_1_2_add_fai_1_U2 ( .A(
        pool_pool_pe_b_peij_1_2_add_fai_1_n4), .ZN(
        pool_pool_pe_b_peij_1_2_add_cprop[2]) );
  XOR2_X1 pool_pool_pe_b_peij_1_2_add_fai_1_U4 ( .A(pool_pool_pe_b_o_data[100]), .B(pool_pool_pe_b_peij_1_2_add_notb[1]), .Z(
        pool_pool_pe_b_peij_1_2_add_fai_1_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_2_add_fai_1_U3 ( .A(
        pool_pool_pe_b_peij_1_2_add_cprop[1]), .B(
        pool_pool_pe_b_peij_1_2_add_fai_1_n5), .Z(
        pool_pool_pe_b_peij_1_2_d_acc[1]) );
  AOI22_X2 pool_pool_pe_b_peij_1_2_add_fai_1_U1 ( .A1(
        pool_pool_pe_b_peij_1_2_add_notb[1]), .A2(pool_pool_pe_b_o_data[100]), 
        .B1(pool_pool_pe_b_peij_1_2_add_fai_1_n5), .B2(
        pool_pool_pe_b_peij_1_2_add_cprop[1]), .ZN(
        pool_pool_pe_b_peij_1_2_add_fai_1_n4) );
  INV_X2 pool_pool_pe_b_peij_1_2_add_fai_2_U2 ( .A(
        pool_pool_pe_b_peij_1_2_add_fai_2_n4), .ZN(
        pool_pool_pe_b_peij_1_2_add_cprop[3]) );
  XOR2_X1 pool_pool_pe_b_peij_1_2_add_fai_2_U4 ( .A(pool_pool_pe_b_o_data[101]), .B(pool_pool_pe_b_peij_1_2_add_notb[2]), .Z(
        pool_pool_pe_b_peij_1_2_add_fai_2_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_2_add_fai_2_U3 ( .A(
        pool_pool_pe_b_peij_1_2_add_cprop[2]), .B(
        pool_pool_pe_b_peij_1_2_add_fai_2_n5), .Z(
        pool_pool_pe_b_peij_1_2_d_acc[2]) );
  AOI22_X2 pool_pool_pe_b_peij_1_2_add_fai_2_U1 ( .A1(
        pool_pool_pe_b_peij_1_2_add_notb[2]), .A2(pool_pool_pe_b_o_data[101]), 
        .B1(pool_pool_pe_b_peij_1_2_add_fai_2_n5), .B2(
        pool_pool_pe_b_peij_1_2_add_cprop[2]), .ZN(
        pool_pool_pe_b_peij_1_2_add_fai_2_n4) );
  INV_X2 pool_pool_pe_b_peij_1_2_add_fai_3_U2 ( .A(
        pool_pool_pe_b_peij_1_2_add_fai_3_n4), .ZN(
        pool_pool_pe_b_peij_1_2_add_cprop[4]) );
  XOR2_X1 pool_pool_pe_b_peij_1_2_add_fai_3_U4 ( .A(pool_pool_pe_b_o_data[102]), .B(pool_pool_pe_b_peij_1_2_add_notb[3]), .Z(
        pool_pool_pe_b_peij_1_2_add_fai_3_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_2_add_fai_3_U3 ( .A(
        pool_pool_pe_b_peij_1_2_add_cprop[3]), .B(
        pool_pool_pe_b_peij_1_2_add_fai_3_n5), .Z(
        pool_pool_pe_b_peij_1_2_d_acc[3]) );
  AOI22_X2 pool_pool_pe_b_peij_1_2_add_fai_3_U1 ( .A1(
        pool_pool_pe_b_peij_1_2_add_notb[3]), .A2(pool_pool_pe_b_o_data[102]), 
        .B1(pool_pool_pe_b_peij_1_2_add_fai_3_n5), .B2(
        pool_pool_pe_b_peij_1_2_add_cprop[3]), .ZN(
        pool_pool_pe_b_peij_1_2_add_fai_3_n4) );
  INV_X2 pool_pool_pe_b_peij_1_2_add_fai_4_U2 ( .A(
        pool_pool_pe_b_peij_1_2_add_fai_4_n4), .ZN(
        pool_pool_pe_b_peij_1_2_add_cprop[5]) );
  XOR2_X1 pool_pool_pe_b_peij_1_2_add_fai_4_U4 ( .A(pool_pool_pe_b_o_data[103]), .B(pool_pool_pe_b_peij_1_2_add_notb[4]), .Z(
        pool_pool_pe_b_peij_1_2_add_fai_4_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_2_add_fai_4_U3 ( .A(
        pool_pool_pe_b_peij_1_2_add_cprop[4]), .B(
        pool_pool_pe_b_peij_1_2_add_fai_4_n5), .Z(
        pool_pool_pe_b_peij_1_2_d_acc[4]) );
  AOI22_X2 pool_pool_pe_b_peij_1_2_add_fai_4_U1 ( .A1(
        pool_pool_pe_b_peij_1_2_add_notb[4]), .A2(pool_pool_pe_b_o_data[103]), 
        .B1(pool_pool_pe_b_peij_1_2_add_fai_4_n5), .B2(
        pool_pool_pe_b_peij_1_2_add_cprop[4]), .ZN(
        pool_pool_pe_b_peij_1_2_add_fai_4_n4) );
  INV_X2 pool_pool_pe_b_peij_1_2_add_fai_5_U2 ( .A(
        pool_pool_pe_b_peij_1_2_add_fai_5_n4), .ZN(
        pool_pool_pe_b_peij_1_2_add_cprop[6]) );
  XOR2_X1 pool_pool_pe_b_peij_1_2_add_fai_5_U4 ( .A(pool_pool_pe_b_o_data[104]), .B(pool_pool_pe_b_peij_1_2_add_notb[5]), .Z(
        pool_pool_pe_b_peij_1_2_add_fai_5_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_2_add_fai_5_U3 ( .A(
        pool_pool_pe_b_peij_1_2_add_cprop[5]), .B(
        pool_pool_pe_b_peij_1_2_add_fai_5_n5), .Z(
        pool_pool_pe_b_peij_1_2_d_acc[5]) );
  AOI22_X2 pool_pool_pe_b_peij_1_2_add_fai_5_U1 ( .A1(
        pool_pool_pe_b_peij_1_2_add_notb[5]), .A2(pool_pool_pe_b_o_data[104]), 
        .B1(pool_pool_pe_b_peij_1_2_add_fai_5_n5), .B2(
        pool_pool_pe_b_peij_1_2_add_cprop[5]), .ZN(
        pool_pool_pe_b_peij_1_2_add_fai_5_n4) );
  INV_X2 pool_pool_pe_b_peij_1_2_add_fai_6_U2 ( .A(
        pool_pool_pe_b_peij_1_2_add_fai_6_n4), .ZN(
        pool_pool_pe_b_peij_1_2_add_cprop[7]) );
  XOR2_X1 pool_pool_pe_b_peij_1_2_add_fai_6_U4 ( .A(pool_pool_pe_b_o_data[105]), .B(pool_pool_pe_b_peij_1_2_add_notb[6]), .Z(
        pool_pool_pe_b_peij_1_2_add_fai_6_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_2_add_fai_6_U3 ( .A(
        pool_pool_pe_b_peij_1_2_add_cprop[6]), .B(
        pool_pool_pe_b_peij_1_2_add_fai_6_n5), .Z(
        pool_pool_pe_b_peij_1_2_d_acc[6]) );
  AOI22_X2 pool_pool_pe_b_peij_1_2_add_fai_6_U1 ( .A1(
        pool_pool_pe_b_peij_1_2_add_notb[6]), .A2(pool_pool_pe_b_o_data[105]), 
        .B1(pool_pool_pe_b_peij_1_2_add_fai_6_n5), .B2(
        pool_pool_pe_b_peij_1_2_add_cprop[6]), .ZN(
        pool_pool_pe_b_peij_1_2_add_fai_6_n4) );
  INV_X2 pool_pool_pe_b_peij_1_2_add_fai_7_U2 ( .A(
        pool_pool_pe_b_peij_1_2_add_fai_7_n4), .ZN(
        pool_pool_pe_b_peij_1_2_add_cprop[8]) );
  XOR2_X1 pool_pool_pe_b_peij_1_2_add_fai_7_U4 ( .A(pool_pool_pe_b_o_data[106]), .B(pool_pool_pe_b_peij_1_2_add_notb[7]), .Z(
        pool_pool_pe_b_peij_1_2_add_fai_7_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_2_add_fai_7_U3 ( .A(
        pool_pool_pe_b_peij_1_2_add_cprop[7]), .B(
        pool_pool_pe_b_peij_1_2_add_fai_7_n5), .Z(
        pool_pool_pe_b_peij_1_2_d_acc[7]) );
  AOI22_X2 pool_pool_pe_b_peij_1_2_add_fai_7_U1 ( .A1(
        pool_pool_pe_b_peij_1_2_add_notb[7]), .A2(pool_pool_pe_b_o_data[106]), 
        .B1(pool_pool_pe_b_peij_1_2_add_fai_7_n5), .B2(
        pool_pool_pe_b_peij_1_2_add_cprop[7]), .ZN(
        pool_pool_pe_b_peij_1_2_add_fai_7_n4) );
  INV_X2 pool_pool_pe_b_peij_1_2_add_fai_8_U2 ( .A(
        pool_pool_pe_b_peij_1_2_add_fai_8_n4), .ZN(
        pool_pool_pe_b_peij_1_2_add_cprop[9]) );
  XOR2_X1 pool_pool_pe_b_peij_1_2_add_fai_8_U4 ( .A(pool_pool_pe_b_o_data[107]), .B(pool_pool_pe_b_peij_1_2_add_notb[8]), .Z(
        pool_pool_pe_b_peij_1_2_add_fai_8_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_2_add_fai_8_U3 ( .A(
        pool_pool_pe_b_peij_1_2_add_cprop[8]), .B(
        pool_pool_pe_b_peij_1_2_add_fai_8_n5), .Z(
        pool_pool_pe_b_peij_1_2_d_acc[8]) );
  AOI22_X2 pool_pool_pe_b_peij_1_2_add_fai_8_U1 ( .A1(
        pool_pool_pe_b_peij_1_2_add_notb[8]), .A2(pool_pool_pe_b_o_data[107]), 
        .B1(pool_pool_pe_b_peij_1_2_add_fai_8_n5), .B2(
        pool_pool_pe_b_peij_1_2_add_cprop[8]), .ZN(
        pool_pool_pe_b_peij_1_2_add_fai_8_n4) );
  INV_X2 pool_pool_pe_b_peij_1_2_add_fai_9_U2 ( .A(
        pool_pool_pe_b_peij_1_2_add_fai_9_n4), .ZN(
        pool_pool_pe_b_peij_1_2_add_cprop[10]) );
  XOR2_X1 pool_pool_pe_b_peij_1_2_add_fai_9_U4 ( .A(pool_pool_pe_b_o_data[108]), .B(pool_pool_pe_b_peij_1_2_add_notb[9]), .Z(
        pool_pool_pe_b_peij_1_2_add_fai_9_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_2_add_fai_9_U3 ( .A(
        pool_pool_pe_b_peij_1_2_add_cprop[9]), .B(
        pool_pool_pe_b_peij_1_2_add_fai_9_n5), .Z(
        pool_pool_pe_b_peij_1_2_d_acc[9]) );
  AOI22_X2 pool_pool_pe_b_peij_1_2_add_fai_9_U1 ( .A1(
        pool_pool_pe_b_peij_1_2_add_notb[9]), .A2(pool_pool_pe_b_o_data[108]), 
        .B1(pool_pool_pe_b_peij_1_2_add_fai_9_n5), .B2(
        pool_pool_pe_b_peij_1_2_add_cprop[9]), .ZN(
        pool_pool_pe_b_peij_1_2_add_fai_9_n4) );
  INV_X2 pool_pool_pe_b_peij_1_2_add_fai_10_U2 ( .A(
        pool_pool_pe_b_peij_1_2_add_fai_10_n4), .ZN(
        pool_pool_pe_b_peij_1_2_add_c_out) );
  XOR2_X1 pool_pool_pe_b_peij_1_2_add_fai_10_U4 ( .A(
        pool_pool_pe_b_o_data[109]), .B(pool_pool_pe_b_peij_1_2_add_notb[10]), 
        .Z(pool_pool_pe_b_peij_1_2_add_fai_10_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_2_add_fai_10_U3 ( .A(
        pool_pool_pe_b_peij_1_2_add_cprop[10]), .B(
        pool_pool_pe_b_peij_1_2_add_fai_10_n5), .Z(
        pool_pool_pe_b_peij_1_2_d_acc[10]) );
  AOI22_X2 pool_pool_pe_b_peij_1_2_add_fai_10_U1 ( .A1(
        pool_pool_pe_b_peij_1_2_add_notb[10]), .A2(pool_pool_pe_b_o_data[109]), 
        .B1(pool_pool_pe_b_peij_1_2_add_fai_10_n5), .B2(
        pool_pool_pe_b_peij_1_2_add_cprop[10]), .ZN(
        pool_pool_pe_b_peij_1_2_add_fai_10_n4) );
  INV_X2 pool_pool_pe_b_peij_1_3_U21 ( .A(pool_sync_clr), .ZN(
        pool_pool_pe_b_peij_1_3_n14) );
  INV_X1 pool_pool_pe_b_peij_1_3_U18 ( .A(pool_pool_pe_b_n1), .ZN(
        pool_pool_pe_b_peij_1_3_n12) );
  AND2_X1 pool_pool_pe_b_peij_1_3_U13 ( .A1(pool_pool_pe_b_peij_1_3_d_acc[0]), 
        .A2(pool_pool_pe_b_peij_1_3_n14), .ZN(pool_pool_pe_b_peij_1_3_n11) );
  AND2_X1 pool_pool_pe_b_peij_1_3_U12 ( .A1(pool_pool_pe_b_peij_1_3_d_acc[1]), 
        .A2(pool_pool_pe_b_peij_1_3_n14), .ZN(pool_pool_pe_b_peij_1_3_n10) );
  AND2_X1 pool_pool_pe_b_peij_1_3_U11 ( .A1(pool_pool_pe_b_peij_1_3_d_acc[2]), 
        .A2(pool_pool_pe_b_peij_1_3_n14), .ZN(pool_pool_pe_b_peij_1_3_n9) );
  AND2_X1 pool_pool_pe_b_peij_1_3_U10 ( .A1(pool_pool_pe_b_peij_1_3_d_acc[3]), 
        .A2(pool_pool_pe_b_peij_1_3_n14), .ZN(pool_pool_pe_b_peij_1_3_n8) );
  AND2_X1 pool_pool_pe_b_peij_1_3_U9 ( .A1(pool_pool_pe_b_peij_1_3_d_acc[4]), 
        .A2(pool_pool_pe_b_peij_1_3_n14), .ZN(pool_pool_pe_b_peij_1_3_n7) );
  AND2_X1 pool_pool_pe_b_peij_1_3_U8 ( .A1(pool_pool_pe_b_peij_1_3_d_acc[5]), 
        .A2(pool_pool_pe_b_peij_1_3_n14), .ZN(pool_pool_pe_b_peij_1_3_n6) );
  AND2_X1 pool_pool_pe_b_peij_1_3_U7 ( .A1(pool_pool_pe_b_peij_1_3_d_acc[6]), 
        .A2(pool_pool_pe_b_peij_1_3_n14), .ZN(pool_pool_pe_b_peij_1_3_n5) );
  AND2_X1 pool_pool_pe_b_peij_1_3_U6 ( .A1(pool_pool_pe_b_peij_1_3_d_acc[7]), 
        .A2(pool_pool_pe_b_peij_1_3_n14), .ZN(pool_pool_pe_b_peij_1_3_n4) );
  AND2_X1 pool_pool_pe_b_peij_1_3_U5 ( .A1(pool_pool_pe_b_peij_1_3_d_acc[8]), 
        .A2(pool_pool_pe_b_peij_1_3_n14), .ZN(pool_pool_pe_b_peij_1_3_n3) );
  AND2_X1 pool_pool_pe_b_peij_1_3_U4 ( .A1(pool_pool_pe_b_peij_1_3_d_acc[9]), 
        .A2(pool_pool_pe_b_peij_1_3_n14), .ZN(pool_pool_pe_b_peij_1_3_n2) );
  AND2_X1 pool_pool_pe_b_peij_1_3_U3 ( .A1(pool_pool_pe_b_peij_1_3_d_acc[10]), 
        .A2(pool_pool_pe_b_peij_1_3_n14), .ZN(pool_pool_pe_b_peij_1_3_n1) );
  DFFR_X1 pool_pool_pe_b_peij_1_3_q_acc_reg_10_ ( .D(
        pool_pool_pe_b_peij_1_3_n1), .CK(pool_pool_pe_b_peij_1_3_gck), .RN(
        pool_pool_pe_b_peij_1_3_n12), .Q(pool_pool_pe_b_o_data[98]) );
  DFFR_X1 pool_pool_pe_b_peij_1_3_q_acc_reg_9_ ( .D(pool_pool_pe_b_peij_1_3_n2), .CK(pool_pool_pe_b_peij_1_3_gck), .RN(pool_pool_pe_b_peij_1_3_n12), .Q(
        pool_pool_pe_b_o_data[97]) );
  DFFR_X1 pool_pool_pe_b_peij_1_3_q_acc_reg_8_ ( .D(pool_pool_pe_b_peij_1_3_n3), .CK(pool_pool_pe_b_peij_1_3_gck), .RN(pool_pool_pe_b_peij_1_3_n12), .Q(
        pool_pool_pe_b_o_data[96]) );
  DFFR_X1 pool_pool_pe_b_peij_1_3_q_acc_reg_7_ ( .D(pool_pool_pe_b_peij_1_3_n4), .CK(pool_pool_pe_b_peij_1_3_gck), .RN(pool_pool_pe_b_peij_1_3_n12), .Q(
        pool_pool_pe_b_o_data[95]) );
  DFFR_X1 pool_pool_pe_b_peij_1_3_q_acc_reg_6_ ( .D(pool_pool_pe_b_peij_1_3_n5), .CK(pool_pool_pe_b_peij_1_3_gck), .RN(pool_pool_pe_b_peij_1_3_n12), .Q(
        pool_pool_pe_b_o_data[94]) );
  DFFR_X1 pool_pool_pe_b_peij_1_3_q_acc_reg_5_ ( .D(pool_pool_pe_b_peij_1_3_n6), .CK(pool_pool_pe_b_peij_1_3_gck), .RN(pool_pool_pe_b_peij_1_3_n12), .Q(
        pool_pool_pe_b_o_data[93]) );
  DFFR_X1 pool_pool_pe_b_peij_1_3_q_acc_reg_4_ ( .D(pool_pool_pe_b_peij_1_3_n7), .CK(pool_pool_pe_b_peij_1_3_gck), .RN(pool_pool_pe_b_peij_1_3_n12), .Q(
        pool_pool_pe_b_o_data[92]) );
  DFFR_X1 pool_pool_pe_b_peij_1_3_q_acc_reg_3_ ( .D(pool_pool_pe_b_peij_1_3_n8), .CK(pool_pool_pe_b_peij_1_3_gck), .RN(pool_pool_pe_b_peij_1_3_n12), .Q(
        pool_pool_pe_b_o_data[91]) );
  DFFR_X1 pool_pool_pe_b_peij_1_3_q_acc_reg_2_ ( .D(pool_pool_pe_b_peij_1_3_n9), .CK(pool_pool_pe_b_peij_1_3_gck), .RN(pool_pool_pe_b_peij_1_3_n12), .Q(
        pool_pool_pe_b_o_data[90]) );
  DFFR_X1 pool_pool_pe_b_peij_1_3_q_acc_reg_1_ ( .D(
        pool_pool_pe_b_peij_1_3_n10), .CK(pool_pool_pe_b_peij_1_3_gck), .RN(
        pool_pool_pe_b_peij_1_3_n12), .Q(pool_pool_pe_b_o_data[89]) );
  DFFR_X1 pool_pool_pe_b_peij_1_3_q_acc_reg_0_ ( .D(
        pool_pool_pe_b_peij_1_3_n11), .CK(pool_pool_pe_b_peij_1_3_gck), .RN(
        pool_pool_pe_b_peij_1_3_n12), .Q(pool_pool_pe_b_o_data[88]) );
  AND3_X2 pool_pool_pe_b_peij_1_3_U20 ( .A1(pool_pool_pe_b_int_pe_en[8]), .A2(
        clk), .A3(1'b1), .ZN(pool_pool_pe_b_peij_1_3_gck) );
  SDFFR_X1 pool_pool_pe_b_peij_1_3_q_k_reg ( .D(1'b0), .SI(
        pool_pool_pe_b_peij_1_3_n14), .SE(1'b0), .CK(
        pool_pool_pe_b_peij_1_3_gck), .RN(pool_pool_pe_b_peij_1_3_n12), .Q(
        pool_pool_pe_b_peij_1_3_q_k) );
  XOR2_X1 pool_pool_pe_b_peij_1_3_add_U11 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_3_q_k), .Z(pool_pool_pe_b_peij_1_3_add_notb[0])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_3_add_U10 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_3_q_k), .Z(pool_pool_pe_b_peij_1_3_add_notb[10])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_3_add_U9 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_3_q_k), .Z(pool_pool_pe_b_peij_1_3_add_notb[1])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_3_add_U8 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_3_q_k), .Z(pool_pool_pe_b_peij_1_3_add_notb[2])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_3_add_U7 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_3_q_k), .Z(pool_pool_pe_b_peij_1_3_add_notb[3])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_3_add_U6 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_3_q_k), .Z(pool_pool_pe_b_peij_1_3_add_notb[4])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_3_add_U5 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_3_q_k), .Z(pool_pool_pe_b_peij_1_3_add_notb[5])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_3_add_U4 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_3_q_k), .Z(pool_pool_pe_b_peij_1_3_add_notb[6])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_3_add_U3 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_3_q_k), .Z(pool_pool_pe_b_peij_1_3_add_notb[7])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_3_add_U2 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_3_q_k), .Z(pool_pool_pe_b_peij_1_3_add_notb[8])
         );
  XOR2_X1 pool_pool_pe_b_peij_1_3_add_U1 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_1_3_q_k), .Z(pool_pool_pe_b_peij_1_3_add_notb[9])
         );
  INV_X2 pool_pool_pe_b_peij_1_3_add_fai_0_U2 ( .A(
        pool_pool_pe_b_peij_1_3_add_fai_0_n4), .ZN(
        pool_pool_pe_b_peij_1_3_add_cprop[1]) );
  XOR2_X1 pool_pool_pe_b_peij_1_3_add_fai_0_U4 ( .A(pool_pool_pe_b_o_data[88]), 
        .B(pool_pool_pe_b_peij_1_3_add_notb[0]), .Z(
        pool_pool_pe_b_peij_1_3_add_fai_0_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_3_add_fai_0_U3 ( .A(
        pool_pool_pe_b_peij_1_3_q_k), .B(pool_pool_pe_b_peij_1_3_add_fai_0_n5), 
        .Z(pool_pool_pe_b_peij_1_3_d_acc[0]) );
  AOI22_X2 pool_pool_pe_b_peij_1_3_add_fai_0_U1 ( .A1(
        pool_pool_pe_b_peij_1_3_add_notb[0]), .A2(pool_pool_pe_b_o_data[88]), 
        .B1(pool_pool_pe_b_peij_1_3_add_fai_0_n5), .B2(
        pool_pool_pe_b_peij_1_3_q_k), .ZN(pool_pool_pe_b_peij_1_3_add_fai_0_n4) );
  INV_X2 pool_pool_pe_b_peij_1_3_add_fai_1_U2 ( .A(
        pool_pool_pe_b_peij_1_3_add_fai_1_n4), .ZN(
        pool_pool_pe_b_peij_1_3_add_cprop[2]) );
  XOR2_X1 pool_pool_pe_b_peij_1_3_add_fai_1_U4 ( .A(pool_pool_pe_b_o_data[89]), 
        .B(pool_pool_pe_b_peij_1_3_add_notb[1]), .Z(
        pool_pool_pe_b_peij_1_3_add_fai_1_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_3_add_fai_1_U3 ( .A(
        pool_pool_pe_b_peij_1_3_add_cprop[1]), .B(
        pool_pool_pe_b_peij_1_3_add_fai_1_n5), .Z(
        pool_pool_pe_b_peij_1_3_d_acc[1]) );
  AOI22_X2 pool_pool_pe_b_peij_1_3_add_fai_1_U1 ( .A1(
        pool_pool_pe_b_peij_1_3_add_notb[1]), .A2(pool_pool_pe_b_o_data[89]), 
        .B1(pool_pool_pe_b_peij_1_3_add_fai_1_n5), .B2(
        pool_pool_pe_b_peij_1_3_add_cprop[1]), .ZN(
        pool_pool_pe_b_peij_1_3_add_fai_1_n4) );
  INV_X2 pool_pool_pe_b_peij_1_3_add_fai_2_U2 ( .A(
        pool_pool_pe_b_peij_1_3_add_fai_2_n4), .ZN(
        pool_pool_pe_b_peij_1_3_add_cprop[3]) );
  XOR2_X1 pool_pool_pe_b_peij_1_3_add_fai_2_U4 ( .A(pool_pool_pe_b_o_data[90]), 
        .B(pool_pool_pe_b_peij_1_3_add_notb[2]), .Z(
        pool_pool_pe_b_peij_1_3_add_fai_2_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_3_add_fai_2_U3 ( .A(
        pool_pool_pe_b_peij_1_3_add_cprop[2]), .B(
        pool_pool_pe_b_peij_1_3_add_fai_2_n5), .Z(
        pool_pool_pe_b_peij_1_3_d_acc[2]) );
  AOI22_X2 pool_pool_pe_b_peij_1_3_add_fai_2_U1 ( .A1(
        pool_pool_pe_b_peij_1_3_add_notb[2]), .A2(pool_pool_pe_b_o_data[90]), 
        .B1(pool_pool_pe_b_peij_1_3_add_fai_2_n5), .B2(
        pool_pool_pe_b_peij_1_3_add_cprop[2]), .ZN(
        pool_pool_pe_b_peij_1_3_add_fai_2_n4) );
  INV_X2 pool_pool_pe_b_peij_1_3_add_fai_3_U2 ( .A(
        pool_pool_pe_b_peij_1_3_add_fai_3_n4), .ZN(
        pool_pool_pe_b_peij_1_3_add_cprop[4]) );
  XOR2_X1 pool_pool_pe_b_peij_1_3_add_fai_3_U4 ( .A(pool_pool_pe_b_o_data[91]), 
        .B(pool_pool_pe_b_peij_1_3_add_notb[3]), .Z(
        pool_pool_pe_b_peij_1_3_add_fai_3_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_3_add_fai_3_U3 ( .A(
        pool_pool_pe_b_peij_1_3_add_cprop[3]), .B(
        pool_pool_pe_b_peij_1_3_add_fai_3_n5), .Z(
        pool_pool_pe_b_peij_1_3_d_acc[3]) );
  AOI22_X2 pool_pool_pe_b_peij_1_3_add_fai_3_U1 ( .A1(
        pool_pool_pe_b_peij_1_3_add_notb[3]), .A2(pool_pool_pe_b_o_data[91]), 
        .B1(pool_pool_pe_b_peij_1_3_add_fai_3_n5), .B2(
        pool_pool_pe_b_peij_1_3_add_cprop[3]), .ZN(
        pool_pool_pe_b_peij_1_3_add_fai_3_n4) );
  INV_X2 pool_pool_pe_b_peij_1_3_add_fai_4_U2 ( .A(
        pool_pool_pe_b_peij_1_3_add_fai_4_n4), .ZN(
        pool_pool_pe_b_peij_1_3_add_cprop[5]) );
  XOR2_X1 pool_pool_pe_b_peij_1_3_add_fai_4_U4 ( .A(pool_pool_pe_b_o_data[92]), 
        .B(pool_pool_pe_b_peij_1_3_add_notb[4]), .Z(
        pool_pool_pe_b_peij_1_3_add_fai_4_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_3_add_fai_4_U3 ( .A(
        pool_pool_pe_b_peij_1_3_add_cprop[4]), .B(
        pool_pool_pe_b_peij_1_3_add_fai_4_n5), .Z(
        pool_pool_pe_b_peij_1_3_d_acc[4]) );
  AOI22_X2 pool_pool_pe_b_peij_1_3_add_fai_4_U1 ( .A1(
        pool_pool_pe_b_peij_1_3_add_notb[4]), .A2(pool_pool_pe_b_o_data[92]), 
        .B1(pool_pool_pe_b_peij_1_3_add_fai_4_n5), .B2(
        pool_pool_pe_b_peij_1_3_add_cprop[4]), .ZN(
        pool_pool_pe_b_peij_1_3_add_fai_4_n4) );
  INV_X2 pool_pool_pe_b_peij_1_3_add_fai_5_U2 ( .A(
        pool_pool_pe_b_peij_1_3_add_fai_5_n4), .ZN(
        pool_pool_pe_b_peij_1_3_add_cprop[6]) );
  XOR2_X1 pool_pool_pe_b_peij_1_3_add_fai_5_U4 ( .A(pool_pool_pe_b_o_data[93]), 
        .B(pool_pool_pe_b_peij_1_3_add_notb[5]), .Z(
        pool_pool_pe_b_peij_1_3_add_fai_5_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_3_add_fai_5_U3 ( .A(
        pool_pool_pe_b_peij_1_3_add_cprop[5]), .B(
        pool_pool_pe_b_peij_1_3_add_fai_5_n5), .Z(
        pool_pool_pe_b_peij_1_3_d_acc[5]) );
  AOI22_X2 pool_pool_pe_b_peij_1_3_add_fai_5_U1 ( .A1(
        pool_pool_pe_b_peij_1_3_add_notb[5]), .A2(pool_pool_pe_b_o_data[93]), 
        .B1(pool_pool_pe_b_peij_1_3_add_fai_5_n5), .B2(
        pool_pool_pe_b_peij_1_3_add_cprop[5]), .ZN(
        pool_pool_pe_b_peij_1_3_add_fai_5_n4) );
  INV_X2 pool_pool_pe_b_peij_1_3_add_fai_6_U2 ( .A(
        pool_pool_pe_b_peij_1_3_add_fai_6_n4), .ZN(
        pool_pool_pe_b_peij_1_3_add_cprop[7]) );
  XOR2_X1 pool_pool_pe_b_peij_1_3_add_fai_6_U4 ( .A(pool_pool_pe_b_o_data[94]), 
        .B(pool_pool_pe_b_peij_1_3_add_notb[6]), .Z(
        pool_pool_pe_b_peij_1_3_add_fai_6_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_3_add_fai_6_U3 ( .A(
        pool_pool_pe_b_peij_1_3_add_cprop[6]), .B(
        pool_pool_pe_b_peij_1_3_add_fai_6_n5), .Z(
        pool_pool_pe_b_peij_1_3_d_acc[6]) );
  AOI22_X2 pool_pool_pe_b_peij_1_3_add_fai_6_U1 ( .A1(
        pool_pool_pe_b_peij_1_3_add_notb[6]), .A2(pool_pool_pe_b_o_data[94]), 
        .B1(pool_pool_pe_b_peij_1_3_add_fai_6_n5), .B2(
        pool_pool_pe_b_peij_1_3_add_cprop[6]), .ZN(
        pool_pool_pe_b_peij_1_3_add_fai_6_n4) );
  INV_X2 pool_pool_pe_b_peij_1_3_add_fai_7_U2 ( .A(
        pool_pool_pe_b_peij_1_3_add_fai_7_n4), .ZN(
        pool_pool_pe_b_peij_1_3_add_cprop[8]) );
  XOR2_X1 pool_pool_pe_b_peij_1_3_add_fai_7_U4 ( .A(pool_pool_pe_b_o_data[95]), 
        .B(pool_pool_pe_b_peij_1_3_add_notb[7]), .Z(
        pool_pool_pe_b_peij_1_3_add_fai_7_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_3_add_fai_7_U3 ( .A(
        pool_pool_pe_b_peij_1_3_add_cprop[7]), .B(
        pool_pool_pe_b_peij_1_3_add_fai_7_n5), .Z(
        pool_pool_pe_b_peij_1_3_d_acc[7]) );
  AOI22_X2 pool_pool_pe_b_peij_1_3_add_fai_7_U1 ( .A1(
        pool_pool_pe_b_peij_1_3_add_notb[7]), .A2(pool_pool_pe_b_o_data[95]), 
        .B1(pool_pool_pe_b_peij_1_3_add_fai_7_n5), .B2(
        pool_pool_pe_b_peij_1_3_add_cprop[7]), .ZN(
        pool_pool_pe_b_peij_1_3_add_fai_7_n4) );
  INV_X2 pool_pool_pe_b_peij_1_3_add_fai_8_U2 ( .A(
        pool_pool_pe_b_peij_1_3_add_fai_8_n4), .ZN(
        pool_pool_pe_b_peij_1_3_add_cprop[9]) );
  XOR2_X1 pool_pool_pe_b_peij_1_3_add_fai_8_U4 ( .A(pool_pool_pe_b_o_data[96]), 
        .B(pool_pool_pe_b_peij_1_3_add_notb[8]), .Z(
        pool_pool_pe_b_peij_1_3_add_fai_8_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_3_add_fai_8_U3 ( .A(
        pool_pool_pe_b_peij_1_3_add_cprop[8]), .B(
        pool_pool_pe_b_peij_1_3_add_fai_8_n5), .Z(
        pool_pool_pe_b_peij_1_3_d_acc[8]) );
  AOI22_X2 pool_pool_pe_b_peij_1_3_add_fai_8_U1 ( .A1(
        pool_pool_pe_b_peij_1_3_add_notb[8]), .A2(pool_pool_pe_b_o_data[96]), 
        .B1(pool_pool_pe_b_peij_1_3_add_fai_8_n5), .B2(
        pool_pool_pe_b_peij_1_3_add_cprop[8]), .ZN(
        pool_pool_pe_b_peij_1_3_add_fai_8_n4) );
  INV_X2 pool_pool_pe_b_peij_1_3_add_fai_9_U2 ( .A(
        pool_pool_pe_b_peij_1_3_add_fai_9_n4), .ZN(
        pool_pool_pe_b_peij_1_3_add_cprop[10]) );
  XOR2_X1 pool_pool_pe_b_peij_1_3_add_fai_9_U4 ( .A(pool_pool_pe_b_o_data[97]), 
        .B(pool_pool_pe_b_peij_1_3_add_notb[9]), .Z(
        pool_pool_pe_b_peij_1_3_add_fai_9_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_3_add_fai_9_U3 ( .A(
        pool_pool_pe_b_peij_1_3_add_cprop[9]), .B(
        pool_pool_pe_b_peij_1_3_add_fai_9_n5), .Z(
        pool_pool_pe_b_peij_1_3_d_acc[9]) );
  AOI22_X2 pool_pool_pe_b_peij_1_3_add_fai_9_U1 ( .A1(
        pool_pool_pe_b_peij_1_3_add_notb[9]), .A2(pool_pool_pe_b_o_data[97]), 
        .B1(pool_pool_pe_b_peij_1_3_add_fai_9_n5), .B2(
        pool_pool_pe_b_peij_1_3_add_cprop[9]), .ZN(
        pool_pool_pe_b_peij_1_3_add_fai_9_n4) );
  INV_X2 pool_pool_pe_b_peij_1_3_add_fai_10_U2 ( .A(
        pool_pool_pe_b_peij_1_3_add_fai_10_n4), .ZN(
        pool_pool_pe_b_peij_1_3_add_c_out) );
  XOR2_X1 pool_pool_pe_b_peij_1_3_add_fai_10_U4 ( .A(pool_pool_pe_b_o_data[98]), .B(pool_pool_pe_b_peij_1_3_add_notb[10]), .Z(
        pool_pool_pe_b_peij_1_3_add_fai_10_n5) );
  XOR2_X1 pool_pool_pe_b_peij_1_3_add_fai_10_U3 ( .A(
        pool_pool_pe_b_peij_1_3_add_cprop[10]), .B(
        pool_pool_pe_b_peij_1_3_add_fai_10_n5), .Z(
        pool_pool_pe_b_peij_1_3_d_acc[10]) );
  AOI22_X2 pool_pool_pe_b_peij_1_3_add_fai_10_U1 ( .A1(
        pool_pool_pe_b_peij_1_3_add_notb[10]), .A2(pool_pool_pe_b_o_data[98]), 
        .B1(pool_pool_pe_b_peij_1_3_add_fai_10_n5), .B2(
        pool_pool_pe_b_peij_1_3_add_cprop[10]), .ZN(
        pool_pool_pe_b_peij_1_3_add_fai_10_n4) );
  INV_X2 pool_pool_pe_b_peij_2_0_U21 ( .A(pool_sync_clr), .ZN(
        pool_pool_pe_b_peij_2_0_n14) );
  INV_X1 pool_pool_pe_b_peij_2_0_U18 ( .A(pool_pool_pe_b_n1), .ZN(
        pool_pool_pe_b_peij_2_0_n12) );
  AND2_X1 pool_pool_pe_b_peij_2_0_U13 ( .A1(pool_pool_pe_b_peij_2_0_d_acc[0]), 
        .A2(pool_pool_pe_b_peij_2_0_n14), .ZN(pool_pool_pe_b_peij_2_0_n11) );
  AND2_X1 pool_pool_pe_b_peij_2_0_U12 ( .A1(pool_pool_pe_b_peij_2_0_d_acc[1]), 
        .A2(pool_pool_pe_b_peij_2_0_n14), .ZN(pool_pool_pe_b_peij_2_0_n10) );
  AND2_X1 pool_pool_pe_b_peij_2_0_U11 ( .A1(pool_pool_pe_b_peij_2_0_d_acc[2]), 
        .A2(pool_pool_pe_b_peij_2_0_n14), .ZN(pool_pool_pe_b_peij_2_0_n9) );
  AND2_X1 pool_pool_pe_b_peij_2_0_U10 ( .A1(pool_pool_pe_b_peij_2_0_d_acc[3]), 
        .A2(pool_pool_pe_b_peij_2_0_n14), .ZN(pool_pool_pe_b_peij_2_0_n8) );
  AND2_X1 pool_pool_pe_b_peij_2_0_U9 ( .A1(pool_pool_pe_b_peij_2_0_d_acc[4]), 
        .A2(pool_pool_pe_b_peij_2_0_n14), .ZN(pool_pool_pe_b_peij_2_0_n7) );
  AND2_X1 pool_pool_pe_b_peij_2_0_U8 ( .A1(pool_pool_pe_b_peij_2_0_d_acc[5]), 
        .A2(pool_pool_pe_b_peij_2_0_n14), .ZN(pool_pool_pe_b_peij_2_0_n6) );
  AND2_X1 pool_pool_pe_b_peij_2_0_U7 ( .A1(pool_pool_pe_b_peij_2_0_d_acc[6]), 
        .A2(pool_pool_pe_b_peij_2_0_n14), .ZN(pool_pool_pe_b_peij_2_0_n5) );
  AND2_X1 pool_pool_pe_b_peij_2_0_U6 ( .A1(pool_pool_pe_b_peij_2_0_d_acc[7]), 
        .A2(pool_pool_pe_b_peij_2_0_n14), .ZN(pool_pool_pe_b_peij_2_0_n4) );
  AND2_X1 pool_pool_pe_b_peij_2_0_U5 ( .A1(pool_pool_pe_b_peij_2_0_d_acc[8]), 
        .A2(pool_pool_pe_b_peij_2_0_n14), .ZN(pool_pool_pe_b_peij_2_0_n3) );
  AND2_X1 pool_pool_pe_b_peij_2_0_U4 ( .A1(pool_pool_pe_b_peij_2_0_d_acc[9]), 
        .A2(pool_pool_pe_b_peij_2_0_n14), .ZN(pool_pool_pe_b_peij_2_0_n2) );
  AND2_X1 pool_pool_pe_b_peij_2_0_U3 ( .A1(pool_pool_pe_b_peij_2_0_d_acc[10]), 
        .A2(pool_pool_pe_b_peij_2_0_n14), .ZN(pool_pool_pe_b_peij_2_0_n1) );
  DFFR_X1 pool_pool_pe_b_peij_2_0_q_acc_reg_10_ ( .D(
        pool_pool_pe_b_peij_2_0_n1), .CK(pool_pool_pe_b_peij_2_0_gck), .RN(
        pool_pool_pe_b_peij_2_0_n12), .Q(pool_pool_pe_b_o_data[87]) );
  DFFR_X1 pool_pool_pe_b_peij_2_0_q_acc_reg_9_ ( .D(pool_pool_pe_b_peij_2_0_n2), .CK(pool_pool_pe_b_peij_2_0_gck), .RN(pool_pool_pe_b_peij_2_0_n12), .Q(
        pool_pool_pe_b_o_data[86]) );
  DFFR_X1 pool_pool_pe_b_peij_2_0_q_acc_reg_8_ ( .D(pool_pool_pe_b_peij_2_0_n3), .CK(pool_pool_pe_b_peij_2_0_gck), .RN(pool_pool_pe_b_peij_2_0_n12), .Q(
        pool_pool_pe_b_o_data[85]) );
  DFFR_X1 pool_pool_pe_b_peij_2_0_q_acc_reg_7_ ( .D(pool_pool_pe_b_peij_2_0_n4), .CK(pool_pool_pe_b_peij_2_0_gck), .RN(pool_pool_pe_b_peij_2_0_n12), .Q(
        pool_pool_pe_b_o_data[84]) );
  DFFR_X1 pool_pool_pe_b_peij_2_0_q_acc_reg_6_ ( .D(pool_pool_pe_b_peij_2_0_n5), .CK(pool_pool_pe_b_peij_2_0_gck), .RN(pool_pool_pe_b_peij_2_0_n12), .Q(
        pool_pool_pe_b_o_data[83]) );
  DFFR_X1 pool_pool_pe_b_peij_2_0_q_acc_reg_5_ ( .D(pool_pool_pe_b_peij_2_0_n6), .CK(pool_pool_pe_b_peij_2_0_gck), .RN(pool_pool_pe_b_peij_2_0_n12), .Q(
        pool_pool_pe_b_o_data[82]) );
  DFFR_X1 pool_pool_pe_b_peij_2_0_q_acc_reg_4_ ( .D(pool_pool_pe_b_peij_2_0_n7), .CK(pool_pool_pe_b_peij_2_0_gck), .RN(pool_pool_pe_b_peij_2_0_n12), .Q(
        pool_pool_pe_b_o_data[81]) );
  DFFR_X1 pool_pool_pe_b_peij_2_0_q_acc_reg_3_ ( .D(pool_pool_pe_b_peij_2_0_n8), .CK(pool_pool_pe_b_peij_2_0_gck), .RN(pool_pool_pe_b_peij_2_0_n12), .Q(
        pool_pool_pe_b_o_data[80]) );
  DFFR_X1 pool_pool_pe_b_peij_2_0_q_acc_reg_2_ ( .D(pool_pool_pe_b_peij_2_0_n9), .CK(pool_pool_pe_b_peij_2_0_gck), .RN(pool_pool_pe_b_peij_2_0_n12), .Q(
        pool_pool_pe_b_o_data[79]) );
  DFFR_X1 pool_pool_pe_b_peij_2_0_q_acc_reg_1_ ( .D(
        pool_pool_pe_b_peij_2_0_n10), .CK(pool_pool_pe_b_peij_2_0_gck), .RN(
        pool_pool_pe_b_peij_2_0_n12), .Q(pool_pool_pe_b_o_data[78]) );
  DFFR_X1 pool_pool_pe_b_peij_2_0_q_acc_reg_0_ ( .D(
        pool_pool_pe_b_peij_2_0_n11), .CK(pool_pool_pe_b_peij_2_0_gck), .RN(
        pool_pool_pe_b_peij_2_0_n12), .Q(pool_pool_pe_b_o_data[77]) );
  AND3_X2 pool_pool_pe_b_peij_2_0_U20 ( .A1(pool_pool_pe_b_int_pe_en[7]), .A2(
        clk), .A3(1'b1), .ZN(pool_pool_pe_b_peij_2_0_gck) );
  SDFFR_X1 pool_pool_pe_b_peij_2_0_q_k_reg ( .D(1'b0), .SI(
        pool_pool_pe_b_peij_2_0_n14), .SE(1'b0), .CK(
        pool_pool_pe_b_peij_2_0_gck), .RN(pool_pool_pe_b_peij_2_0_n12), .Q(
        pool_pool_pe_b_peij_2_0_q_k) );
  XOR2_X1 pool_pool_pe_b_peij_2_0_add_U11 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_0_q_k), .Z(pool_pool_pe_b_peij_2_0_add_notb[0])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_0_add_U10 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_0_q_k), .Z(pool_pool_pe_b_peij_2_0_add_notb[10])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_0_add_U9 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_0_q_k), .Z(pool_pool_pe_b_peij_2_0_add_notb[1])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_0_add_U8 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_0_q_k), .Z(pool_pool_pe_b_peij_2_0_add_notb[2])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_0_add_U7 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_0_q_k), .Z(pool_pool_pe_b_peij_2_0_add_notb[3])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_0_add_U6 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_0_q_k), .Z(pool_pool_pe_b_peij_2_0_add_notb[4])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_0_add_U5 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_0_q_k), .Z(pool_pool_pe_b_peij_2_0_add_notb[5])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_0_add_U4 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_0_q_k), .Z(pool_pool_pe_b_peij_2_0_add_notb[6])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_0_add_U3 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_0_q_k), .Z(pool_pool_pe_b_peij_2_0_add_notb[7])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_0_add_U2 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_0_q_k), .Z(pool_pool_pe_b_peij_2_0_add_notb[8])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_0_add_U1 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_0_q_k), .Z(pool_pool_pe_b_peij_2_0_add_notb[9])
         );
  INV_X2 pool_pool_pe_b_peij_2_0_add_fai_0_U2 ( .A(
        pool_pool_pe_b_peij_2_0_add_fai_0_n4), .ZN(
        pool_pool_pe_b_peij_2_0_add_cprop[1]) );
  XOR2_X1 pool_pool_pe_b_peij_2_0_add_fai_0_U4 ( .A(pool_pool_pe_b_o_data[77]), 
        .B(pool_pool_pe_b_peij_2_0_add_notb[0]), .Z(
        pool_pool_pe_b_peij_2_0_add_fai_0_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_0_add_fai_0_U3 ( .A(
        pool_pool_pe_b_peij_2_0_q_k), .B(pool_pool_pe_b_peij_2_0_add_fai_0_n5), 
        .Z(pool_pool_pe_b_peij_2_0_d_acc[0]) );
  AOI22_X2 pool_pool_pe_b_peij_2_0_add_fai_0_U1 ( .A1(
        pool_pool_pe_b_peij_2_0_add_notb[0]), .A2(pool_pool_pe_b_o_data[77]), 
        .B1(pool_pool_pe_b_peij_2_0_add_fai_0_n5), .B2(
        pool_pool_pe_b_peij_2_0_q_k), .ZN(pool_pool_pe_b_peij_2_0_add_fai_0_n4) );
  INV_X2 pool_pool_pe_b_peij_2_0_add_fai_1_U2 ( .A(
        pool_pool_pe_b_peij_2_0_add_fai_1_n4), .ZN(
        pool_pool_pe_b_peij_2_0_add_cprop[2]) );
  XOR2_X1 pool_pool_pe_b_peij_2_0_add_fai_1_U4 ( .A(pool_pool_pe_b_o_data[78]), 
        .B(pool_pool_pe_b_peij_2_0_add_notb[1]), .Z(
        pool_pool_pe_b_peij_2_0_add_fai_1_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_0_add_fai_1_U3 ( .A(
        pool_pool_pe_b_peij_2_0_add_cprop[1]), .B(
        pool_pool_pe_b_peij_2_0_add_fai_1_n5), .Z(
        pool_pool_pe_b_peij_2_0_d_acc[1]) );
  AOI22_X2 pool_pool_pe_b_peij_2_0_add_fai_1_U1 ( .A1(
        pool_pool_pe_b_peij_2_0_add_notb[1]), .A2(pool_pool_pe_b_o_data[78]), 
        .B1(pool_pool_pe_b_peij_2_0_add_fai_1_n5), .B2(
        pool_pool_pe_b_peij_2_0_add_cprop[1]), .ZN(
        pool_pool_pe_b_peij_2_0_add_fai_1_n4) );
  INV_X2 pool_pool_pe_b_peij_2_0_add_fai_2_U2 ( .A(
        pool_pool_pe_b_peij_2_0_add_fai_2_n4), .ZN(
        pool_pool_pe_b_peij_2_0_add_cprop[3]) );
  XOR2_X1 pool_pool_pe_b_peij_2_0_add_fai_2_U4 ( .A(pool_pool_pe_b_o_data[79]), 
        .B(pool_pool_pe_b_peij_2_0_add_notb[2]), .Z(
        pool_pool_pe_b_peij_2_0_add_fai_2_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_0_add_fai_2_U3 ( .A(
        pool_pool_pe_b_peij_2_0_add_cprop[2]), .B(
        pool_pool_pe_b_peij_2_0_add_fai_2_n5), .Z(
        pool_pool_pe_b_peij_2_0_d_acc[2]) );
  AOI22_X2 pool_pool_pe_b_peij_2_0_add_fai_2_U1 ( .A1(
        pool_pool_pe_b_peij_2_0_add_notb[2]), .A2(pool_pool_pe_b_o_data[79]), 
        .B1(pool_pool_pe_b_peij_2_0_add_fai_2_n5), .B2(
        pool_pool_pe_b_peij_2_0_add_cprop[2]), .ZN(
        pool_pool_pe_b_peij_2_0_add_fai_2_n4) );
  INV_X2 pool_pool_pe_b_peij_2_0_add_fai_3_U2 ( .A(
        pool_pool_pe_b_peij_2_0_add_fai_3_n4), .ZN(
        pool_pool_pe_b_peij_2_0_add_cprop[4]) );
  XOR2_X1 pool_pool_pe_b_peij_2_0_add_fai_3_U4 ( .A(pool_pool_pe_b_o_data[80]), 
        .B(pool_pool_pe_b_peij_2_0_add_notb[3]), .Z(
        pool_pool_pe_b_peij_2_0_add_fai_3_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_0_add_fai_3_U3 ( .A(
        pool_pool_pe_b_peij_2_0_add_cprop[3]), .B(
        pool_pool_pe_b_peij_2_0_add_fai_3_n5), .Z(
        pool_pool_pe_b_peij_2_0_d_acc[3]) );
  AOI22_X2 pool_pool_pe_b_peij_2_0_add_fai_3_U1 ( .A1(
        pool_pool_pe_b_peij_2_0_add_notb[3]), .A2(pool_pool_pe_b_o_data[80]), 
        .B1(pool_pool_pe_b_peij_2_0_add_fai_3_n5), .B2(
        pool_pool_pe_b_peij_2_0_add_cprop[3]), .ZN(
        pool_pool_pe_b_peij_2_0_add_fai_3_n4) );
  INV_X2 pool_pool_pe_b_peij_2_0_add_fai_4_U2 ( .A(
        pool_pool_pe_b_peij_2_0_add_fai_4_n4), .ZN(
        pool_pool_pe_b_peij_2_0_add_cprop[5]) );
  XOR2_X1 pool_pool_pe_b_peij_2_0_add_fai_4_U4 ( .A(pool_pool_pe_b_o_data[81]), 
        .B(pool_pool_pe_b_peij_2_0_add_notb[4]), .Z(
        pool_pool_pe_b_peij_2_0_add_fai_4_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_0_add_fai_4_U3 ( .A(
        pool_pool_pe_b_peij_2_0_add_cprop[4]), .B(
        pool_pool_pe_b_peij_2_0_add_fai_4_n5), .Z(
        pool_pool_pe_b_peij_2_0_d_acc[4]) );
  AOI22_X2 pool_pool_pe_b_peij_2_0_add_fai_4_U1 ( .A1(
        pool_pool_pe_b_peij_2_0_add_notb[4]), .A2(pool_pool_pe_b_o_data[81]), 
        .B1(pool_pool_pe_b_peij_2_0_add_fai_4_n5), .B2(
        pool_pool_pe_b_peij_2_0_add_cprop[4]), .ZN(
        pool_pool_pe_b_peij_2_0_add_fai_4_n4) );
  INV_X2 pool_pool_pe_b_peij_2_0_add_fai_5_U2 ( .A(
        pool_pool_pe_b_peij_2_0_add_fai_5_n4), .ZN(
        pool_pool_pe_b_peij_2_0_add_cprop[6]) );
  XOR2_X1 pool_pool_pe_b_peij_2_0_add_fai_5_U4 ( .A(pool_pool_pe_b_o_data[82]), 
        .B(pool_pool_pe_b_peij_2_0_add_notb[5]), .Z(
        pool_pool_pe_b_peij_2_0_add_fai_5_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_0_add_fai_5_U3 ( .A(
        pool_pool_pe_b_peij_2_0_add_cprop[5]), .B(
        pool_pool_pe_b_peij_2_0_add_fai_5_n5), .Z(
        pool_pool_pe_b_peij_2_0_d_acc[5]) );
  AOI22_X2 pool_pool_pe_b_peij_2_0_add_fai_5_U1 ( .A1(
        pool_pool_pe_b_peij_2_0_add_notb[5]), .A2(pool_pool_pe_b_o_data[82]), 
        .B1(pool_pool_pe_b_peij_2_0_add_fai_5_n5), .B2(
        pool_pool_pe_b_peij_2_0_add_cprop[5]), .ZN(
        pool_pool_pe_b_peij_2_0_add_fai_5_n4) );
  INV_X2 pool_pool_pe_b_peij_2_0_add_fai_6_U2 ( .A(
        pool_pool_pe_b_peij_2_0_add_fai_6_n4), .ZN(
        pool_pool_pe_b_peij_2_0_add_cprop[7]) );
  XOR2_X1 pool_pool_pe_b_peij_2_0_add_fai_6_U4 ( .A(pool_pool_pe_b_o_data[83]), 
        .B(pool_pool_pe_b_peij_2_0_add_notb[6]), .Z(
        pool_pool_pe_b_peij_2_0_add_fai_6_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_0_add_fai_6_U3 ( .A(
        pool_pool_pe_b_peij_2_0_add_cprop[6]), .B(
        pool_pool_pe_b_peij_2_0_add_fai_6_n5), .Z(
        pool_pool_pe_b_peij_2_0_d_acc[6]) );
  AOI22_X2 pool_pool_pe_b_peij_2_0_add_fai_6_U1 ( .A1(
        pool_pool_pe_b_peij_2_0_add_notb[6]), .A2(pool_pool_pe_b_o_data[83]), 
        .B1(pool_pool_pe_b_peij_2_0_add_fai_6_n5), .B2(
        pool_pool_pe_b_peij_2_0_add_cprop[6]), .ZN(
        pool_pool_pe_b_peij_2_0_add_fai_6_n4) );
  INV_X2 pool_pool_pe_b_peij_2_0_add_fai_7_U2 ( .A(
        pool_pool_pe_b_peij_2_0_add_fai_7_n4), .ZN(
        pool_pool_pe_b_peij_2_0_add_cprop[8]) );
  XOR2_X1 pool_pool_pe_b_peij_2_0_add_fai_7_U4 ( .A(pool_pool_pe_b_o_data[84]), 
        .B(pool_pool_pe_b_peij_2_0_add_notb[7]), .Z(
        pool_pool_pe_b_peij_2_0_add_fai_7_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_0_add_fai_7_U3 ( .A(
        pool_pool_pe_b_peij_2_0_add_cprop[7]), .B(
        pool_pool_pe_b_peij_2_0_add_fai_7_n5), .Z(
        pool_pool_pe_b_peij_2_0_d_acc[7]) );
  AOI22_X2 pool_pool_pe_b_peij_2_0_add_fai_7_U1 ( .A1(
        pool_pool_pe_b_peij_2_0_add_notb[7]), .A2(pool_pool_pe_b_o_data[84]), 
        .B1(pool_pool_pe_b_peij_2_0_add_fai_7_n5), .B2(
        pool_pool_pe_b_peij_2_0_add_cprop[7]), .ZN(
        pool_pool_pe_b_peij_2_0_add_fai_7_n4) );
  INV_X2 pool_pool_pe_b_peij_2_0_add_fai_8_U2 ( .A(
        pool_pool_pe_b_peij_2_0_add_fai_8_n4), .ZN(
        pool_pool_pe_b_peij_2_0_add_cprop[9]) );
  XOR2_X1 pool_pool_pe_b_peij_2_0_add_fai_8_U4 ( .A(pool_pool_pe_b_o_data[85]), 
        .B(pool_pool_pe_b_peij_2_0_add_notb[8]), .Z(
        pool_pool_pe_b_peij_2_0_add_fai_8_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_0_add_fai_8_U3 ( .A(
        pool_pool_pe_b_peij_2_0_add_cprop[8]), .B(
        pool_pool_pe_b_peij_2_0_add_fai_8_n5), .Z(
        pool_pool_pe_b_peij_2_0_d_acc[8]) );
  AOI22_X2 pool_pool_pe_b_peij_2_0_add_fai_8_U1 ( .A1(
        pool_pool_pe_b_peij_2_0_add_notb[8]), .A2(pool_pool_pe_b_o_data[85]), 
        .B1(pool_pool_pe_b_peij_2_0_add_fai_8_n5), .B2(
        pool_pool_pe_b_peij_2_0_add_cprop[8]), .ZN(
        pool_pool_pe_b_peij_2_0_add_fai_8_n4) );
  INV_X2 pool_pool_pe_b_peij_2_0_add_fai_9_U2 ( .A(
        pool_pool_pe_b_peij_2_0_add_fai_9_n4), .ZN(
        pool_pool_pe_b_peij_2_0_add_cprop[10]) );
  XOR2_X1 pool_pool_pe_b_peij_2_0_add_fai_9_U4 ( .A(pool_pool_pe_b_o_data[86]), 
        .B(pool_pool_pe_b_peij_2_0_add_notb[9]), .Z(
        pool_pool_pe_b_peij_2_0_add_fai_9_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_0_add_fai_9_U3 ( .A(
        pool_pool_pe_b_peij_2_0_add_cprop[9]), .B(
        pool_pool_pe_b_peij_2_0_add_fai_9_n5), .Z(
        pool_pool_pe_b_peij_2_0_d_acc[9]) );
  AOI22_X2 pool_pool_pe_b_peij_2_0_add_fai_9_U1 ( .A1(
        pool_pool_pe_b_peij_2_0_add_notb[9]), .A2(pool_pool_pe_b_o_data[86]), 
        .B1(pool_pool_pe_b_peij_2_0_add_fai_9_n5), .B2(
        pool_pool_pe_b_peij_2_0_add_cprop[9]), .ZN(
        pool_pool_pe_b_peij_2_0_add_fai_9_n4) );
  INV_X2 pool_pool_pe_b_peij_2_0_add_fai_10_U2 ( .A(
        pool_pool_pe_b_peij_2_0_add_fai_10_n4), .ZN(
        pool_pool_pe_b_peij_2_0_add_c_out) );
  XOR2_X1 pool_pool_pe_b_peij_2_0_add_fai_10_U4 ( .A(pool_pool_pe_b_o_data[87]), .B(pool_pool_pe_b_peij_2_0_add_notb[10]), .Z(
        pool_pool_pe_b_peij_2_0_add_fai_10_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_0_add_fai_10_U3 ( .A(
        pool_pool_pe_b_peij_2_0_add_cprop[10]), .B(
        pool_pool_pe_b_peij_2_0_add_fai_10_n5), .Z(
        pool_pool_pe_b_peij_2_0_d_acc[10]) );
  AOI22_X2 pool_pool_pe_b_peij_2_0_add_fai_10_U1 ( .A1(
        pool_pool_pe_b_peij_2_0_add_notb[10]), .A2(pool_pool_pe_b_o_data[87]), 
        .B1(pool_pool_pe_b_peij_2_0_add_fai_10_n5), .B2(
        pool_pool_pe_b_peij_2_0_add_cprop[10]), .ZN(
        pool_pool_pe_b_peij_2_0_add_fai_10_n4) );
  INV_X2 pool_pool_pe_b_peij_2_1_U21 ( .A(pool_sync_clr), .ZN(
        pool_pool_pe_b_peij_2_1_n14) );
  INV_X1 pool_pool_pe_b_peij_2_1_U18 ( .A(pool_pool_pe_b_n1), .ZN(
        pool_pool_pe_b_peij_2_1_n12) );
  AND2_X1 pool_pool_pe_b_peij_2_1_U13 ( .A1(pool_pool_pe_b_peij_2_1_d_acc[0]), 
        .A2(pool_pool_pe_b_peij_2_1_n14), .ZN(pool_pool_pe_b_peij_2_1_n11) );
  AND2_X1 pool_pool_pe_b_peij_2_1_U12 ( .A1(pool_pool_pe_b_peij_2_1_d_acc[1]), 
        .A2(pool_pool_pe_b_peij_2_1_n14), .ZN(pool_pool_pe_b_peij_2_1_n10) );
  AND2_X1 pool_pool_pe_b_peij_2_1_U11 ( .A1(pool_pool_pe_b_peij_2_1_d_acc[2]), 
        .A2(pool_pool_pe_b_peij_2_1_n14), .ZN(pool_pool_pe_b_peij_2_1_n9) );
  AND2_X1 pool_pool_pe_b_peij_2_1_U10 ( .A1(pool_pool_pe_b_peij_2_1_d_acc[3]), 
        .A2(pool_pool_pe_b_peij_2_1_n14), .ZN(pool_pool_pe_b_peij_2_1_n8) );
  AND2_X1 pool_pool_pe_b_peij_2_1_U9 ( .A1(pool_pool_pe_b_peij_2_1_d_acc[4]), 
        .A2(pool_pool_pe_b_peij_2_1_n14), .ZN(pool_pool_pe_b_peij_2_1_n7) );
  AND2_X1 pool_pool_pe_b_peij_2_1_U8 ( .A1(pool_pool_pe_b_peij_2_1_d_acc[5]), 
        .A2(pool_pool_pe_b_peij_2_1_n14), .ZN(pool_pool_pe_b_peij_2_1_n6) );
  AND2_X1 pool_pool_pe_b_peij_2_1_U7 ( .A1(pool_pool_pe_b_peij_2_1_d_acc[6]), 
        .A2(pool_pool_pe_b_peij_2_1_n14), .ZN(pool_pool_pe_b_peij_2_1_n5) );
  AND2_X1 pool_pool_pe_b_peij_2_1_U6 ( .A1(pool_pool_pe_b_peij_2_1_d_acc[7]), 
        .A2(pool_pool_pe_b_peij_2_1_n14), .ZN(pool_pool_pe_b_peij_2_1_n4) );
  AND2_X1 pool_pool_pe_b_peij_2_1_U5 ( .A1(pool_pool_pe_b_peij_2_1_d_acc[8]), 
        .A2(pool_pool_pe_b_peij_2_1_n14), .ZN(pool_pool_pe_b_peij_2_1_n3) );
  AND2_X1 pool_pool_pe_b_peij_2_1_U4 ( .A1(pool_pool_pe_b_peij_2_1_d_acc[9]), 
        .A2(pool_pool_pe_b_peij_2_1_n14), .ZN(pool_pool_pe_b_peij_2_1_n2) );
  AND2_X1 pool_pool_pe_b_peij_2_1_U3 ( .A1(pool_pool_pe_b_peij_2_1_d_acc[10]), 
        .A2(pool_pool_pe_b_peij_2_1_n14), .ZN(pool_pool_pe_b_peij_2_1_n1) );
  DFFR_X1 pool_pool_pe_b_peij_2_1_q_acc_reg_10_ ( .D(
        pool_pool_pe_b_peij_2_1_n1), .CK(pool_pool_pe_b_peij_2_1_gck), .RN(
        pool_pool_pe_b_peij_2_1_n12), .Q(pool_pool_pe_b_o_data[76]) );
  DFFR_X1 pool_pool_pe_b_peij_2_1_q_acc_reg_9_ ( .D(pool_pool_pe_b_peij_2_1_n2), .CK(pool_pool_pe_b_peij_2_1_gck), .RN(pool_pool_pe_b_peij_2_1_n12), .Q(
        pool_pool_pe_b_o_data[75]) );
  DFFR_X1 pool_pool_pe_b_peij_2_1_q_acc_reg_8_ ( .D(pool_pool_pe_b_peij_2_1_n3), .CK(pool_pool_pe_b_peij_2_1_gck), .RN(pool_pool_pe_b_peij_2_1_n12), .Q(
        pool_pool_pe_b_o_data[74]) );
  DFFR_X1 pool_pool_pe_b_peij_2_1_q_acc_reg_7_ ( .D(pool_pool_pe_b_peij_2_1_n4), .CK(pool_pool_pe_b_peij_2_1_gck), .RN(pool_pool_pe_b_peij_2_1_n12), .Q(
        pool_pool_pe_b_o_data[73]) );
  DFFR_X1 pool_pool_pe_b_peij_2_1_q_acc_reg_6_ ( .D(pool_pool_pe_b_peij_2_1_n5), .CK(pool_pool_pe_b_peij_2_1_gck), .RN(pool_pool_pe_b_peij_2_1_n12), .Q(
        pool_pool_pe_b_o_data[72]) );
  DFFR_X1 pool_pool_pe_b_peij_2_1_q_acc_reg_5_ ( .D(pool_pool_pe_b_peij_2_1_n6), .CK(pool_pool_pe_b_peij_2_1_gck), .RN(pool_pool_pe_b_peij_2_1_n12), .Q(
        pool_pool_pe_b_o_data[71]) );
  DFFR_X1 pool_pool_pe_b_peij_2_1_q_acc_reg_4_ ( .D(pool_pool_pe_b_peij_2_1_n7), .CK(pool_pool_pe_b_peij_2_1_gck), .RN(pool_pool_pe_b_peij_2_1_n12), .Q(
        pool_pool_pe_b_o_data[70]) );
  DFFR_X1 pool_pool_pe_b_peij_2_1_q_acc_reg_3_ ( .D(pool_pool_pe_b_peij_2_1_n8), .CK(pool_pool_pe_b_peij_2_1_gck), .RN(pool_pool_pe_b_peij_2_1_n12), .Q(
        pool_pool_pe_b_o_data[69]) );
  DFFR_X1 pool_pool_pe_b_peij_2_1_q_acc_reg_2_ ( .D(pool_pool_pe_b_peij_2_1_n9), .CK(pool_pool_pe_b_peij_2_1_gck), .RN(pool_pool_pe_b_peij_2_1_n12), .Q(
        pool_pool_pe_b_o_data[68]) );
  DFFR_X1 pool_pool_pe_b_peij_2_1_q_acc_reg_1_ ( .D(
        pool_pool_pe_b_peij_2_1_n10), .CK(pool_pool_pe_b_peij_2_1_gck), .RN(
        pool_pool_pe_b_peij_2_1_n12), .Q(pool_pool_pe_b_o_data[67]) );
  DFFR_X1 pool_pool_pe_b_peij_2_1_q_acc_reg_0_ ( .D(
        pool_pool_pe_b_peij_2_1_n11), .CK(pool_pool_pe_b_peij_2_1_gck), .RN(
        pool_pool_pe_b_peij_2_1_n12), .Q(pool_pool_pe_b_o_data[66]) );
  AND3_X2 pool_pool_pe_b_peij_2_1_U20 ( .A1(pool_pool_pe_b_int_pe_en[6]), .A2(
        clk), .A3(1'b1), .ZN(pool_pool_pe_b_peij_2_1_gck) );
  SDFFR_X1 pool_pool_pe_b_peij_2_1_q_k_reg ( .D(1'b0), .SI(
        pool_pool_pe_b_peij_2_1_n14), .SE(1'b0), .CK(
        pool_pool_pe_b_peij_2_1_gck), .RN(pool_pool_pe_b_peij_2_1_n12), .Q(
        pool_pool_pe_b_peij_2_1_q_k) );
  XOR2_X1 pool_pool_pe_b_peij_2_1_add_U11 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_1_q_k), .Z(pool_pool_pe_b_peij_2_1_add_notb[0])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_1_add_U10 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_1_q_k), .Z(pool_pool_pe_b_peij_2_1_add_notb[10])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_1_add_U9 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_1_q_k), .Z(pool_pool_pe_b_peij_2_1_add_notb[1])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_1_add_U8 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_1_q_k), .Z(pool_pool_pe_b_peij_2_1_add_notb[2])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_1_add_U7 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_1_q_k), .Z(pool_pool_pe_b_peij_2_1_add_notb[3])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_1_add_U6 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_1_q_k), .Z(pool_pool_pe_b_peij_2_1_add_notb[4])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_1_add_U5 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_1_q_k), .Z(pool_pool_pe_b_peij_2_1_add_notb[5])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_1_add_U4 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_1_q_k), .Z(pool_pool_pe_b_peij_2_1_add_notb[6])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_1_add_U3 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_1_q_k), .Z(pool_pool_pe_b_peij_2_1_add_notb[7])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_1_add_U2 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_1_q_k), .Z(pool_pool_pe_b_peij_2_1_add_notb[8])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_1_add_U1 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_1_q_k), .Z(pool_pool_pe_b_peij_2_1_add_notb[9])
         );
  INV_X2 pool_pool_pe_b_peij_2_1_add_fai_0_U2 ( .A(
        pool_pool_pe_b_peij_2_1_add_fai_0_n4), .ZN(
        pool_pool_pe_b_peij_2_1_add_cprop[1]) );
  XOR2_X1 pool_pool_pe_b_peij_2_1_add_fai_0_U4 ( .A(pool_pool_pe_b_o_data[66]), 
        .B(pool_pool_pe_b_peij_2_1_add_notb[0]), .Z(
        pool_pool_pe_b_peij_2_1_add_fai_0_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_1_add_fai_0_U3 ( .A(
        pool_pool_pe_b_peij_2_1_q_k), .B(pool_pool_pe_b_peij_2_1_add_fai_0_n5), 
        .Z(pool_pool_pe_b_peij_2_1_d_acc[0]) );
  AOI22_X2 pool_pool_pe_b_peij_2_1_add_fai_0_U1 ( .A1(
        pool_pool_pe_b_peij_2_1_add_notb[0]), .A2(pool_pool_pe_b_o_data[66]), 
        .B1(pool_pool_pe_b_peij_2_1_add_fai_0_n5), .B2(
        pool_pool_pe_b_peij_2_1_q_k), .ZN(pool_pool_pe_b_peij_2_1_add_fai_0_n4) );
  INV_X2 pool_pool_pe_b_peij_2_1_add_fai_1_U2 ( .A(
        pool_pool_pe_b_peij_2_1_add_fai_1_n4), .ZN(
        pool_pool_pe_b_peij_2_1_add_cprop[2]) );
  XOR2_X1 pool_pool_pe_b_peij_2_1_add_fai_1_U4 ( .A(pool_pool_pe_b_o_data[67]), 
        .B(pool_pool_pe_b_peij_2_1_add_notb[1]), .Z(
        pool_pool_pe_b_peij_2_1_add_fai_1_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_1_add_fai_1_U3 ( .A(
        pool_pool_pe_b_peij_2_1_add_cprop[1]), .B(
        pool_pool_pe_b_peij_2_1_add_fai_1_n5), .Z(
        pool_pool_pe_b_peij_2_1_d_acc[1]) );
  AOI22_X2 pool_pool_pe_b_peij_2_1_add_fai_1_U1 ( .A1(
        pool_pool_pe_b_peij_2_1_add_notb[1]), .A2(pool_pool_pe_b_o_data[67]), 
        .B1(pool_pool_pe_b_peij_2_1_add_fai_1_n5), .B2(
        pool_pool_pe_b_peij_2_1_add_cprop[1]), .ZN(
        pool_pool_pe_b_peij_2_1_add_fai_1_n4) );
  INV_X2 pool_pool_pe_b_peij_2_1_add_fai_2_U2 ( .A(
        pool_pool_pe_b_peij_2_1_add_fai_2_n4), .ZN(
        pool_pool_pe_b_peij_2_1_add_cprop[3]) );
  XOR2_X1 pool_pool_pe_b_peij_2_1_add_fai_2_U4 ( .A(pool_pool_pe_b_o_data[68]), 
        .B(pool_pool_pe_b_peij_2_1_add_notb[2]), .Z(
        pool_pool_pe_b_peij_2_1_add_fai_2_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_1_add_fai_2_U3 ( .A(
        pool_pool_pe_b_peij_2_1_add_cprop[2]), .B(
        pool_pool_pe_b_peij_2_1_add_fai_2_n5), .Z(
        pool_pool_pe_b_peij_2_1_d_acc[2]) );
  AOI22_X2 pool_pool_pe_b_peij_2_1_add_fai_2_U1 ( .A1(
        pool_pool_pe_b_peij_2_1_add_notb[2]), .A2(pool_pool_pe_b_o_data[68]), 
        .B1(pool_pool_pe_b_peij_2_1_add_fai_2_n5), .B2(
        pool_pool_pe_b_peij_2_1_add_cprop[2]), .ZN(
        pool_pool_pe_b_peij_2_1_add_fai_2_n4) );
  INV_X2 pool_pool_pe_b_peij_2_1_add_fai_3_U2 ( .A(
        pool_pool_pe_b_peij_2_1_add_fai_3_n4), .ZN(
        pool_pool_pe_b_peij_2_1_add_cprop[4]) );
  XOR2_X1 pool_pool_pe_b_peij_2_1_add_fai_3_U4 ( .A(pool_pool_pe_b_o_data[69]), 
        .B(pool_pool_pe_b_peij_2_1_add_notb[3]), .Z(
        pool_pool_pe_b_peij_2_1_add_fai_3_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_1_add_fai_3_U3 ( .A(
        pool_pool_pe_b_peij_2_1_add_cprop[3]), .B(
        pool_pool_pe_b_peij_2_1_add_fai_3_n5), .Z(
        pool_pool_pe_b_peij_2_1_d_acc[3]) );
  AOI22_X2 pool_pool_pe_b_peij_2_1_add_fai_3_U1 ( .A1(
        pool_pool_pe_b_peij_2_1_add_notb[3]), .A2(pool_pool_pe_b_o_data[69]), 
        .B1(pool_pool_pe_b_peij_2_1_add_fai_3_n5), .B2(
        pool_pool_pe_b_peij_2_1_add_cprop[3]), .ZN(
        pool_pool_pe_b_peij_2_1_add_fai_3_n4) );
  INV_X2 pool_pool_pe_b_peij_2_1_add_fai_4_U2 ( .A(
        pool_pool_pe_b_peij_2_1_add_fai_4_n4), .ZN(
        pool_pool_pe_b_peij_2_1_add_cprop[5]) );
  XOR2_X1 pool_pool_pe_b_peij_2_1_add_fai_4_U4 ( .A(pool_pool_pe_b_o_data[70]), 
        .B(pool_pool_pe_b_peij_2_1_add_notb[4]), .Z(
        pool_pool_pe_b_peij_2_1_add_fai_4_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_1_add_fai_4_U3 ( .A(
        pool_pool_pe_b_peij_2_1_add_cprop[4]), .B(
        pool_pool_pe_b_peij_2_1_add_fai_4_n5), .Z(
        pool_pool_pe_b_peij_2_1_d_acc[4]) );
  AOI22_X2 pool_pool_pe_b_peij_2_1_add_fai_4_U1 ( .A1(
        pool_pool_pe_b_peij_2_1_add_notb[4]), .A2(pool_pool_pe_b_o_data[70]), 
        .B1(pool_pool_pe_b_peij_2_1_add_fai_4_n5), .B2(
        pool_pool_pe_b_peij_2_1_add_cprop[4]), .ZN(
        pool_pool_pe_b_peij_2_1_add_fai_4_n4) );
  INV_X2 pool_pool_pe_b_peij_2_1_add_fai_5_U2 ( .A(
        pool_pool_pe_b_peij_2_1_add_fai_5_n4), .ZN(
        pool_pool_pe_b_peij_2_1_add_cprop[6]) );
  XOR2_X1 pool_pool_pe_b_peij_2_1_add_fai_5_U4 ( .A(pool_pool_pe_b_o_data[71]), 
        .B(pool_pool_pe_b_peij_2_1_add_notb[5]), .Z(
        pool_pool_pe_b_peij_2_1_add_fai_5_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_1_add_fai_5_U3 ( .A(
        pool_pool_pe_b_peij_2_1_add_cprop[5]), .B(
        pool_pool_pe_b_peij_2_1_add_fai_5_n5), .Z(
        pool_pool_pe_b_peij_2_1_d_acc[5]) );
  AOI22_X2 pool_pool_pe_b_peij_2_1_add_fai_5_U1 ( .A1(
        pool_pool_pe_b_peij_2_1_add_notb[5]), .A2(pool_pool_pe_b_o_data[71]), 
        .B1(pool_pool_pe_b_peij_2_1_add_fai_5_n5), .B2(
        pool_pool_pe_b_peij_2_1_add_cprop[5]), .ZN(
        pool_pool_pe_b_peij_2_1_add_fai_5_n4) );
  INV_X2 pool_pool_pe_b_peij_2_1_add_fai_6_U2 ( .A(
        pool_pool_pe_b_peij_2_1_add_fai_6_n4), .ZN(
        pool_pool_pe_b_peij_2_1_add_cprop[7]) );
  XOR2_X1 pool_pool_pe_b_peij_2_1_add_fai_6_U4 ( .A(pool_pool_pe_b_o_data[72]), 
        .B(pool_pool_pe_b_peij_2_1_add_notb[6]), .Z(
        pool_pool_pe_b_peij_2_1_add_fai_6_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_1_add_fai_6_U3 ( .A(
        pool_pool_pe_b_peij_2_1_add_cprop[6]), .B(
        pool_pool_pe_b_peij_2_1_add_fai_6_n5), .Z(
        pool_pool_pe_b_peij_2_1_d_acc[6]) );
  AOI22_X2 pool_pool_pe_b_peij_2_1_add_fai_6_U1 ( .A1(
        pool_pool_pe_b_peij_2_1_add_notb[6]), .A2(pool_pool_pe_b_o_data[72]), 
        .B1(pool_pool_pe_b_peij_2_1_add_fai_6_n5), .B2(
        pool_pool_pe_b_peij_2_1_add_cprop[6]), .ZN(
        pool_pool_pe_b_peij_2_1_add_fai_6_n4) );
  INV_X2 pool_pool_pe_b_peij_2_1_add_fai_7_U2 ( .A(
        pool_pool_pe_b_peij_2_1_add_fai_7_n4), .ZN(
        pool_pool_pe_b_peij_2_1_add_cprop[8]) );
  XOR2_X1 pool_pool_pe_b_peij_2_1_add_fai_7_U4 ( .A(pool_pool_pe_b_o_data[73]), 
        .B(pool_pool_pe_b_peij_2_1_add_notb[7]), .Z(
        pool_pool_pe_b_peij_2_1_add_fai_7_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_1_add_fai_7_U3 ( .A(
        pool_pool_pe_b_peij_2_1_add_cprop[7]), .B(
        pool_pool_pe_b_peij_2_1_add_fai_7_n5), .Z(
        pool_pool_pe_b_peij_2_1_d_acc[7]) );
  AOI22_X2 pool_pool_pe_b_peij_2_1_add_fai_7_U1 ( .A1(
        pool_pool_pe_b_peij_2_1_add_notb[7]), .A2(pool_pool_pe_b_o_data[73]), 
        .B1(pool_pool_pe_b_peij_2_1_add_fai_7_n5), .B2(
        pool_pool_pe_b_peij_2_1_add_cprop[7]), .ZN(
        pool_pool_pe_b_peij_2_1_add_fai_7_n4) );
  INV_X2 pool_pool_pe_b_peij_2_1_add_fai_8_U2 ( .A(
        pool_pool_pe_b_peij_2_1_add_fai_8_n4), .ZN(
        pool_pool_pe_b_peij_2_1_add_cprop[9]) );
  XOR2_X1 pool_pool_pe_b_peij_2_1_add_fai_8_U4 ( .A(pool_pool_pe_b_o_data[74]), 
        .B(pool_pool_pe_b_peij_2_1_add_notb[8]), .Z(
        pool_pool_pe_b_peij_2_1_add_fai_8_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_1_add_fai_8_U3 ( .A(
        pool_pool_pe_b_peij_2_1_add_cprop[8]), .B(
        pool_pool_pe_b_peij_2_1_add_fai_8_n5), .Z(
        pool_pool_pe_b_peij_2_1_d_acc[8]) );
  AOI22_X2 pool_pool_pe_b_peij_2_1_add_fai_8_U1 ( .A1(
        pool_pool_pe_b_peij_2_1_add_notb[8]), .A2(pool_pool_pe_b_o_data[74]), 
        .B1(pool_pool_pe_b_peij_2_1_add_fai_8_n5), .B2(
        pool_pool_pe_b_peij_2_1_add_cprop[8]), .ZN(
        pool_pool_pe_b_peij_2_1_add_fai_8_n4) );
  INV_X2 pool_pool_pe_b_peij_2_1_add_fai_9_U2 ( .A(
        pool_pool_pe_b_peij_2_1_add_fai_9_n4), .ZN(
        pool_pool_pe_b_peij_2_1_add_cprop[10]) );
  XOR2_X1 pool_pool_pe_b_peij_2_1_add_fai_9_U4 ( .A(pool_pool_pe_b_o_data[75]), 
        .B(pool_pool_pe_b_peij_2_1_add_notb[9]), .Z(
        pool_pool_pe_b_peij_2_1_add_fai_9_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_1_add_fai_9_U3 ( .A(
        pool_pool_pe_b_peij_2_1_add_cprop[9]), .B(
        pool_pool_pe_b_peij_2_1_add_fai_9_n5), .Z(
        pool_pool_pe_b_peij_2_1_d_acc[9]) );
  AOI22_X2 pool_pool_pe_b_peij_2_1_add_fai_9_U1 ( .A1(
        pool_pool_pe_b_peij_2_1_add_notb[9]), .A2(pool_pool_pe_b_o_data[75]), 
        .B1(pool_pool_pe_b_peij_2_1_add_fai_9_n5), .B2(
        pool_pool_pe_b_peij_2_1_add_cprop[9]), .ZN(
        pool_pool_pe_b_peij_2_1_add_fai_9_n4) );
  INV_X2 pool_pool_pe_b_peij_2_1_add_fai_10_U2 ( .A(
        pool_pool_pe_b_peij_2_1_add_fai_10_n4), .ZN(
        pool_pool_pe_b_peij_2_1_add_c_out) );
  XOR2_X1 pool_pool_pe_b_peij_2_1_add_fai_10_U4 ( .A(pool_pool_pe_b_o_data[76]), .B(pool_pool_pe_b_peij_2_1_add_notb[10]), .Z(
        pool_pool_pe_b_peij_2_1_add_fai_10_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_1_add_fai_10_U3 ( .A(
        pool_pool_pe_b_peij_2_1_add_cprop[10]), .B(
        pool_pool_pe_b_peij_2_1_add_fai_10_n5), .Z(
        pool_pool_pe_b_peij_2_1_d_acc[10]) );
  AOI22_X2 pool_pool_pe_b_peij_2_1_add_fai_10_U1 ( .A1(
        pool_pool_pe_b_peij_2_1_add_notb[10]), .A2(pool_pool_pe_b_o_data[76]), 
        .B1(pool_pool_pe_b_peij_2_1_add_fai_10_n5), .B2(
        pool_pool_pe_b_peij_2_1_add_cprop[10]), .ZN(
        pool_pool_pe_b_peij_2_1_add_fai_10_n4) );
  INV_X2 pool_pool_pe_b_peij_2_2_U21 ( .A(pool_sync_clr), .ZN(
        pool_pool_pe_b_peij_2_2_n14) );
  INV_X1 pool_pool_pe_b_peij_2_2_U18 ( .A(pool_pool_pe_b_n1), .ZN(
        pool_pool_pe_b_peij_2_2_n12) );
  AND2_X1 pool_pool_pe_b_peij_2_2_U13 ( .A1(pool_pool_pe_b_peij_2_2_d_acc[0]), 
        .A2(pool_pool_pe_b_peij_2_2_n14), .ZN(pool_pool_pe_b_peij_2_2_n11) );
  AND2_X1 pool_pool_pe_b_peij_2_2_U12 ( .A1(pool_pool_pe_b_peij_2_2_d_acc[1]), 
        .A2(pool_pool_pe_b_peij_2_2_n14), .ZN(pool_pool_pe_b_peij_2_2_n10) );
  AND2_X1 pool_pool_pe_b_peij_2_2_U11 ( .A1(pool_pool_pe_b_peij_2_2_d_acc[2]), 
        .A2(pool_pool_pe_b_peij_2_2_n14), .ZN(pool_pool_pe_b_peij_2_2_n9) );
  AND2_X1 pool_pool_pe_b_peij_2_2_U10 ( .A1(pool_pool_pe_b_peij_2_2_d_acc[3]), 
        .A2(pool_pool_pe_b_peij_2_2_n14), .ZN(pool_pool_pe_b_peij_2_2_n8) );
  AND2_X1 pool_pool_pe_b_peij_2_2_U9 ( .A1(pool_pool_pe_b_peij_2_2_d_acc[4]), 
        .A2(pool_pool_pe_b_peij_2_2_n14), .ZN(pool_pool_pe_b_peij_2_2_n7) );
  AND2_X1 pool_pool_pe_b_peij_2_2_U8 ( .A1(pool_pool_pe_b_peij_2_2_d_acc[5]), 
        .A2(pool_pool_pe_b_peij_2_2_n14), .ZN(pool_pool_pe_b_peij_2_2_n6) );
  AND2_X1 pool_pool_pe_b_peij_2_2_U7 ( .A1(pool_pool_pe_b_peij_2_2_d_acc[6]), 
        .A2(pool_pool_pe_b_peij_2_2_n14), .ZN(pool_pool_pe_b_peij_2_2_n5) );
  AND2_X1 pool_pool_pe_b_peij_2_2_U6 ( .A1(pool_pool_pe_b_peij_2_2_d_acc[7]), 
        .A2(pool_pool_pe_b_peij_2_2_n14), .ZN(pool_pool_pe_b_peij_2_2_n4) );
  AND2_X1 pool_pool_pe_b_peij_2_2_U5 ( .A1(pool_pool_pe_b_peij_2_2_d_acc[8]), 
        .A2(pool_pool_pe_b_peij_2_2_n14), .ZN(pool_pool_pe_b_peij_2_2_n3) );
  AND2_X1 pool_pool_pe_b_peij_2_2_U4 ( .A1(pool_pool_pe_b_peij_2_2_d_acc[9]), 
        .A2(pool_pool_pe_b_peij_2_2_n14), .ZN(pool_pool_pe_b_peij_2_2_n2) );
  AND2_X1 pool_pool_pe_b_peij_2_2_U3 ( .A1(pool_pool_pe_b_peij_2_2_d_acc[10]), 
        .A2(pool_pool_pe_b_peij_2_2_n14), .ZN(pool_pool_pe_b_peij_2_2_n1) );
  DFFR_X1 pool_pool_pe_b_peij_2_2_q_acc_reg_10_ ( .D(
        pool_pool_pe_b_peij_2_2_n1), .CK(pool_pool_pe_b_peij_2_2_gck), .RN(
        pool_pool_pe_b_peij_2_2_n12), .Q(pool_pool_pe_b_o_data[65]) );
  DFFR_X1 pool_pool_pe_b_peij_2_2_q_acc_reg_9_ ( .D(pool_pool_pe_b_peij_2_2_n2), .CK(pool_pool_pe_b_peij_2_2_gck), .RN(pool_pool_pe_b_peij_2_2_n12), .Q(
        pool_pool_pe_b_o_data[64]) );
  DFFR_X1 pool_pool_pe_b_peij_2_2_q_acc_reg_8_ ( .D(pool_pool_pe_b_peij_2_2_n3), .CK(pool_pool_pe_b_peij_2_2_gck), .RN(pool_pool_pe_b_peij_2_2_n12), .Q(
        pool_pool_pe_b_o_data[63]) );
  DFFR_X1 pool_pool_pe_b_peij_2_2_q_acc_reg_7_ ( .D(pool_pool_pe_b_peij_2_2_n4), .CK(pool_pool_pe_b_peij_2_2_gck), .RN(pool_pool_pe_b_peij_2_2_n12), .Q(
        pool_pool_pe_b_o_data[62]) );
  DFFR_X1 pool_pool_pe_b_peij_2_2_q_acc_reg_6_ ( .D(pool_pool_pe_b_peij_2_2_n5), .CK(pool_pool_pe_b_peij_2_2_gck), .RN(pool_pool_pe_b_peij_2_2_n12), .Q(
        pool_pool_pe_b_o_data[61]) );
  DFFR_X1 pool_pool_pe_b_peij_2_2_q_acc_reg_5_ ( .D(pool_pool_pe_b_peij_2_2_n6), .CK(pool_pool_pe_b_peij_2_2_gck), .RN(pool_pool_pe_b_peij_2_2_n12), .Q(
        pool_pool_pe_b_o_data[60]) );
  DFFR_X1 pool_pool_pe_b_peij_2_2_q_acc_reg_4_ ( .D(pool_pool_pe_b_peij_2_2_n7), .CK(pool_pool_pe_b_peij_2_2_gck), .RN(pool_pool_pe_b_peij_2_2_n12), .Q(
        pool_pool_pe_b_o_data[59]) );
  DFFR_X1 pool_pool_pe_b_peij_2_2_q_acc_reg_3_ ( .D(pool_pool_pe_b_peij_2_2_n8), .CK(pool_pool_pe_b_peij_2_2_gck), .RN(pool_pool_pe_b_peij_2_2_n12), .Q(
        pool_pool_pe_b_o_data[58]) );
  DFFR_X1 pool_pool_pe_b_peij_2_2_q_acc_reg_2_ ( .D(pool_pool_pe_b_peij_2_2_n9), .CK(pool_pool_pe_b_peij_2_2_gck), .RN(pool_pool_pe_b_peij_2_2_n12), .Q(
        pool_pool_pe_b_o_data[57]) );
  DFFR_X1 pool_pool_pe_b_peij_2_2_q_acc_reg_1_ ( .D(
        pool_pool_pe_b_peij_2_2_n10), .CK(pool_pool_pe_b_peij_2_2_gck), .RN(
        pool_pool_pe_b_peij_2_2_n12), .Q(pool_pool_pe_b_o_data[56]) );
  DFFR_X1 pool_pool_pe_b_peij_2_2_q_acc_reg_0_ ( .D(
        pool_pool_pe_b_peij_2_2_n11), .CK(pool_pool_pe_b_peij_2_2_gck), .RN(
        pool_pool_pe_b_peij_2_2_n12), .Q(pool_pool_pe_b_o_data[55]) );
  AND3_X2 pool_pool_pe_b_peij_2_2_U20 ( .A1(pool_pool_pe_b_int_pe_en[5]), .A2(
        clk), .A3(1'b1), .ZN(pool_pool_pe_b_peij_2_2_gck) );
  SDFFR_X1 pool_pool_pe_b_peij_2_2_q_k_reg ( .D(1'b0), .SI(
        pool_pool_pe_b_peij_2_2_n14), .SE(1'b0), .CK(
        pool_pool_pe_b_peij_2_2_gck), .RN(pool_pool_pe_b_peij_2_2_n12), .Q(
        pool_pool_pe_b_peij_2_2_q_k) );
  XOR2_X1 pool_pool_pe_b_peij_2_2_add_U11 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_2_q_k), .Z(pool_pool_pe_b_peij_2_2_add_notb[0])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_2_add_U10 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_2_q_k), .Z(pool_pool_pe_b_peij_2_2_add_notb[10])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_2_add_U9 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_2_q_k), .Z(pool_pool_pe_b_peij_2_2_add_notb[1])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_2_add_U8 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_2_q_k), .Z(pool_pool_pe_b_peij_2_2_add_notb[2])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_2_add_U7 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_2_q_k), .Z(pool_pool_pe_b_peij_2_2_add_notb[3])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_2_add_U6 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_2_q_k), .Z(pool_pool_pe_b_peij_2_2_add_notb[4])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_2_add_U5 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_2_q_k), .Z(pool_pool_pe_b_peij_2_2_add_notb[5])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_2_add_U4 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_2_q_k), .Z(pool_pool_pe_b_peij_2_2_add_notb[6])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_2_add_U3 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_2_q_k), .Z(pool_pool_pe_b_peij_2_2_add_notb[7])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_2_add_U2 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_2_q_k), .Z(pool_pool_pe_b_peij_2_2_add_notb[8])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_2_add_U1 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_2_q_k), .Z(pool_pool_pe_b_peij_2_2_add_notb[9])
         );
  INV_X2 pool_pool_pe_b_peij_2_2_add_fai_0_U2 ( .A(
        pool_pool_pe_b_peij_2_2_add_fai_0_n4), .ZN(
        pool_pool_pe_b_peij_2_2_add_cprop[1]) );
  XOR2_X1 pool_pool_pe_b_peij_2_2_add_fai_0_U4 ( .A(pool_pool_pe_b_o_data[55]), 
        .B(pool_pool_pe_b_peij_2_2_add_notb[0]), .Z(
        pool_pool_pe_b_peij_2_2_add_fai_0_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_2_add_fai_0_U3 ( .A(
        pool_pool_pe_b_peij_2_2_q_k), .B(pool_pool_pe_b_peij_2_2_add_fai_0_n5), 
        .Z(pool_pool_pe_b_peij_2_2_d_acc[0]) );
  AOI22_X2 pool_pool_pe_b_peij_2_2_add_fai_0_U1 ( .A1(
        pool_pool_pe_b_peij_2_2_add_notb[0]), .A2(pool_pool_pe_b_o_data[55]), 
        .B1(pool_pool_pe_b_peij_2_2_add_fai_0_n5), .B2(
        pool_pool_pe_b_peij_2_2_q_k), .ZN(pool_pool_pe_b_peij_2_2_add_fai_0_n4) );
  INV_X2 pool_pool_pe_b_peij_2_2_add_fai_1_U2 ( .A(
        pool_pool_pe_b_peij_2_2_add_fai_1_n4), .ZN(
        pool_pool_pe_b_peij_2_2_add_cprop[2]) );
  XOR2_X1 pool_pool_pe_b_peij_2_2_add_fai_1_U4 ( .A(pool_pool_pe_b_o_data[56]), 
        .B(pool_pool_pe_b_peij_2_2_add_notb[1]), .Z(
        pool_pool_pe_b_peij_2_2_add_fai_1_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_2_add_fai_1_U3 ( .A(
        pool_pool_pe_b_peij_2_2_add_cprop[1]), .B(
        pool_pool_pe_b_peij_2_2_add_fai_1_n5), .Z(
        pool_pool_pe_b_peij_2_2_d_acc[1]) );
  AOI22_X2 pool_pool_pe_b_peij_2_2_add_fai_1_U1 ( .A1(
        pool_pool_pe_b_peij_2_2_add_notb[1]), .A2(pool_pool_pe_b_o_data[56]), 
        .B1(pool_pool_pe_b_peij_2_2_add_fai_1_n5), .B2(
        pool_pool_pe_b_peij_2_2_add_cprop[1]), .ZN(
        pool_pool_pe_b_peij_2_2_add_fai_1_n4) );
  INV_X2 pool_pool_pe_b_peij_2_2_add_fai_2_U2 ( .A(
        pool_pool_pe_b_peij_2_2_add_fai_2_n4), .ZN(
        pool_pool_pe_b_peij_2_2_add_cprop[3]) );
  XOR2_X1 pool_pool_pe_b_peij_2_2_add_fai_2_U4 ( .A(pool_pool_pe_b_o_data[57]), 
        .B(pool_pool_pe_b_peij_2_2_add_notb[2]), .Z(
        pool_pool_pe_b_peij_2_2_add_fai_2_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_2_add_fai_2_U3 ( .A(
        pool_pool_pe_b_peij_2_2_add_cprop[2]), .B(
        pool_pool_pe_b_peij_2_2_add_fai_2_n5), .Z(
        pool_pool_pe_b_peij_2_2_d_acc[2]) );
  AOI22_X2 pool_pool_pe_b_peij_2_2_add_fai_2_U1 ( .A1(
        pool_pool_pe_b_peij_2_2_add_notb[2]), .A2(pool_pool_pe_b_o_data[57]), 
        .B1(pool_pool_pe_b_peij_2_2_add_fai_2_n5), .B2(
        pool_pool_pe_b_peij_2_2_add_cprop[2]), .ZN(
        pool_pool_pe_b_peij_2_2_add_fai_2_n4) );
  INV_X2 pool_pool_pe_b_peij_2_2_add_fai_3_U2 ( .A(
        pool_pool_pe_b_peij_2_2_add_fai_3_n4), .ZN(
        pool_pool_pe_b_peij_2_2_add_cprop[4]) );
  XOR2_X1 pool_pool_pe_b_peij_2_2_add_fai_3_U4 ( .A(pool_pool_pe_b_o_data[58]), 
        .B(pool_pool_pe_b_peij_2_2_add_notb[3]), .Z(
        pool_pool_pe_b_peij_2_2_add_fai_3_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_2_add_fai_3_U3 ( .A(
        pool_pool_pe_b_peij_2_2_add_cprop[3]), .B(
        pool_pool_pe_b_peij_2_2_add_fai_3_n5), .Z(
        pool_pool_pe_b_peij_2_2_d_acc[3]) );
  AOI22_X2 pool_pool_pe_b_peij_2_2_add_fai_3_U1 ( .A1(
        pool_pool_pe_b_peij_2_2_add_notb[3]), .A2(pool_pool_pe_b_o_data[58]), 
        .B1(pool_pool_pe_b_peij_2_2_add_fai_3_n5), .B2(
        pool_pool_pe_b_peij_2_2_add_cprop[3]), .ZN(
        pool_pool_pe_b_peij_2_2_add_fai_3_n4) );
  INV_X2 pool_pool_pe_b_peij_2_2_add_fai_4_U2 ( .A(
        pool_pool_pe_b_peij_2_2_add_fai_4_n4), .ZN(
        pool_pool_pe_b_peij_2_2_add_cprop[5]) );
  XOR2_X1 pool_pool_pe_b_peij_2_2_add_fai_4_U4 ( .A(pool_pool_pe_b_o_data[59]), 
        .B(pool_pool_pe_b_peij_2_2_add_notb[4]), .Z(
        pool_pool_pe_b_peij_2_2_add_fai_4_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_2_add_fai_4_U3 ( .A(
        pool_pool_pe_b_peij_2_2_add_cprop[4]), .B(
        pool_pool_pe_b_peij_2_2_add_fai_4_n5), .Z(
        pool_pool_pe_b_peij_2_2_d_acc[4]) );
  AOI22_X2 pool_pool_pe_b_peij_2_2_add_fai_4_U1 ( .A1(
        pool_pool_pe_b_peij_2_2_add_notb[4]), .A2(pool_pool_pe_b_o_data[59]), 
        .B1(pool_pool_pe_b_peij_2_2_add_fai_4_n5), .B2(
        pool_pool_pe_b_peij_2_2_add_cprop[4]), .ZN(
        pool_pool_pe_b_peij_2_2_add_fai_4_n4) );
  INV_X2 pool_pool_pe_b_peij_2_2_add_fai_5_U2 ( .A(
        pool_pool_pe_b_peij_2_2_add_fai_5_n4), .ZN(
        pool_pool_pe_b_peij_2_2_add_cprop[6]) );
  XOR2_X1 pool_pool_pe_b_peij_2_2_add_fai_5_U4 ( .A(pool_pool_pe_b_o_data[60]), 
        .B(pool_pool_pe_b_peij_2_2_add_notb[5]), .Z(
        pool_pool_pe_b_peij_2_2_add_fai_5_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_2_add_fai_5_U3 ( .A(
        pool_pool_pe_b_peij_2_2_add_cprop[5]), .B(
        pool_pool_pe_b_peij_2_2_add_fai_5_n5), .Z(
        pool_pool_pe_b_peij_2_2_d_acc[5]) );
  AOI22_X2 pool_pool_pe_b_peij_2_2_add_fai_5_U1 ( .A1(
        pool_pool_pe_b_peij_2_2_add_notb[5]), .A2(pool_pool_pe_b_o_data[60]), 
        .B1(pool_pool_pe_b_peij_2_2_add_fai_5_n5), .B2(
        pool_pool_pe_b_peij_2_2_add_cprop[5]), .ZN(
        pool_pool_pe_b_peij_2_2_add_fai_5_n4) );
  INV_X2 pool_pool_pe_b_peij_2_2_add_fai_6_U2 ( .A(
        pool_pool_pe_b_peij_2_2_add_fai_6_n4), .ZN(
        pool_pool_pe_b_peij_2_2_add_cprop[7]) );
  XOR2_X1 pool_pool_pe_b_peij_2_2_add_fai_6_U4 ( .A(pool_pool_pe_b_o_data[61]), 
        .B(pool_pool_pe_b_peij_2_2_add_notb[6]), .Z(
        pool_pool_pe_b_peij_2_2_add_fai_6_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_2_add_fai_6_U3 ( .A(
        pool_pool_pe_b_peij_2_2_add_cprop[6]), .B(
        pool_pool_pe_b_peij_2_2_add_fai_6_n5), .Z(
        pool_pool_pe_b_peij_2_2_d_acc[6]) );
  AOI22_X2 pool_pool_pe_b_peij_2_2_add_fai_6_U1 ( .A1(
        pool_pool_pe_b_peij_2_2_add_notb[6]), .A2(pool_pool_pe_b_o_data[61]), 
        .B1(pool_pool_pe_b_peij_2_2_add_fai_6_n5), .B2(
        pool_pool_pe_b_peij_2_2_add_cprop[6]), .ZN(
        pool_pool_pe_b_peij_2_2_add_fai_6_n4) );
  INV_X2 pool_pool_pe_b_peij_2_2_add_fai_7_U2 ( .A(
        pool_pool_pe_b_peij_2_2_add_fai_7_n4), .ZN(
        pool_pool_pe_b_peij_2_2_add_cprop[8]) );
  XOR2_X1 pool_pool_pe_b_peij_2_2_add_fai_7_U4 ( .A(pool_pool_pe_b_o_data[62]), 
        .B(pool_pool_pe_b_peij_2_2_add_notb[7]), .Z(
        pool_pool_pe_b_peij_2_2_add_fai_7_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_2_add_fai_7_U3 ( .A(
        pool_pool_pe_b_peij_2_2_add_cprop[7]), .B(
        pool_pool_pe_b_peij_2_2_add_fai_7_n5), .Z(
        pool_pool_pe_b_peij_2_2_d_acc[7]) );
  AOI22_X2 pool_pool_pe_b_peij_2_2_add_fai_7_U1 ( .A1(
        pool_pool_pe_b_peij_2_2_add_notb[7]), .A2(pool_pool_pe_b_o_data[62]), 
        .B1(pool_pool_pe_b_peij_2_2_add_fai_7_n5), .B2(
        pool_pool_pe_b_peij_2_2_add_cprop[7]), .ZN(
        pool_pool_pe_b_peij_2_2_add_fai_7_n4) );
  INV_X2 pool_pool_pe_b_peij_2_2_add_fai_8_U2 ( .A(
        pool_pool_pe_b_peij_2_2_add_fai_8_n4), .ZN(
        pool_pool_pe_b_peij_2_2_add_cprop[9]) );
  XOR2_X1 pool_pool_pe_b_peij_2_2_add_fai_8_U4 ( .A(pool_pool_pe_b_o_data[63]), 
        .B(pool_pool_pe_b_peij_2_2_add_notb[8]), .Z(
        pool_pool_pe_b_peij_2_2_add_fai_8_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_2_add_fai_8_U3 ( .A(
        pool_pool_pe_b_peij_2_2_add_cprop[8]), .B(
        pool_pool_pe_b_peij_2_2_add_fai_8_n5), .Z(
        pool_pool_pe_b_peij_2_2_d_acc[8]) );
  AOI22_X2 pool_pool_pe_b_peij_2_2_add_fai_8_U1 ( .A1(
        pool_pool_pe_b_peij_2_2_add_notb[8]), .A2(pool_pool_pe_b_o_data[63]), 
        .B1(pool_pool_pe_b_peij_2_2_add_fai_8_n5), .B2(
        pool_pool_pe_b_peij_2_2_add_cprop[8]), .ZN(
        pool_pool_pe_b_peij_2_2_add_fai_8_n4) );
  INV_X2 pool_pool_pe_b_peij_2_2_add_fai_9_U2 ( .A(
        pool_pool_pe_b_peij_2_2_add_fai_9_n4), .ZN(
        pool_pool_pe_b_peij_2_2_add_cprop[10]) );
  XOR2_X1 pool_pool_pe_b_peij_2_2_add_fai_9_U4 ( .A(pool_pool_pe_b_o_data[64]), 
        .B(pool_pool_pe_b_peij_2_2_add_notb[9]), .Z(
        pool_pool_pe_b_peij_2_2_add_fai_9_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_2_add_fai_9_U3 ( .A(
        pool_pool_pe_b_peij_2_2_add_cprop[9]), .B(
        pool_pool_pe_b_peij_2_2_add_fai_9_n5), .Z(
        pool_pool_pe_b_peij_2_2_d_acc[9]) );
  AOI22_X2 pool_pool_pe_b_peij_2_2_add_fai_9_U1 ( .A1(
        pool_pool_pe_b_peij_2_2_add_notb[9]), .A2(pool_pool_pe_b_o_data[64]), 
        .B1(pool_pool_pe_b_peij_2_2_add_fai_9_n5), .B2(
        pool_pool_pe_b_peij_2_2_add_cprop[9]), .ZN(
        pool_pool_pe_b_peij_2_2_add_fai_9_n4) );
  INV_X2 pool_pool_pe_b_peij_2_2_add_fai_10_U2 ( .A(
        pool_pool_pe_b_peij_2_2_add_fai_10_n4), .ZN(
        pool_pool_pe_b_peij_2_2_add_c_out) );
  XOR2_X1 pool_pool_pe_b_peij_2_2_add_fai_10_U4 ( .A(pool_pool_pe_b_o_data[65]), .B(pool_pool_pe_b_peij_2_2_add_notb[10]), .Z(
        pool_pool_pe_b_peij_2_2_add_fai_10_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_2_add_fai_10_U3 ( .A(
        pool_pool_pe_b_peij_2_2_add_cprop[10]), .B(
        pool_pool_pe_b_peij_2_2_add_fai_10_n5), .Z(
        pool_pool_pe_b_peij_2_2_d_acc[10]) );
  AOI22_X2 pool_pool_pe_b_peij_2_2_add_fai_10_U1 ( .A1(
        pool_pool_pe_b_peij_2_2_add_notb[10]), .A2(pool_pool_pe_b_o_data[65]), 
        .B1(pool_pool_pe_b_peij_2_2_add_fai_10_n5), .B2(
        pool_pool_pe_b_peij_2_2_add_cprop[10]), .ZN(
        pool_pool_pe_b_peij_2_2_add_fai_10_n4) );
  INV_X2 pool_pool_pe_b_peij_2_3_U21 ( .A(pool_sync_clr), .ZN(
        pool_pool_pe_b_peij_2_3_n14) );
  INV_X1 pool_pool_pe_b_peij_2_3_U18 ( .A(pool_pool_pe_b_n1), .ZN(
        pool_pool_pe_b_peij_2_3_n12) );
  AND2_X1 pool_pool_pe_b_peij_2_3_U13 ( .A1(pool_pool_pe_b_peij_2_3_d_acc[0]), 
        .A2(pool_pool_pe_b_peij_2_3_n14), .ZN(pool_pool_pe_b_peij_2_3_n11) );
  AND2_X1 pool_pool_pe_b_peij_2_3_U12 ( .A1(pool_pool_pe_b_peij_2_3_d_acc[1]), 
        .A2(pool_pool_pe_b_peij_2_3_n14), .ZN(pool_pool_pe_b_peij_2_3_n10) );
  AND2_X1 pool_pool_pe_b_peij_2_3_U11 ( .A1(pool_pool_pe_b_peij_2_3_d_acc[2]), 
        .A2(pool_pool_pe_b_peij_2_3_n14), .ZN(pool_pool_pe_b_peij_2_3_n9) );
  AND2_X1 pool_pool_pe_b_peij_2_3_U10 ( .A1(pool_pool_pe_b_peij_2_3_d_acc[3]), 
        .A2(pool_pool_pe_b_peij_2_3_n14), .ZN(pool_pool_pe_b_peij_2_3_n8) );
  AND2_X1 pool_pool_pe_b_peij_2_3_U9 ( .A1(pool_pool_pe_b_peij_2_3_d_acc[4]), 
        .A2(pool_pool_pe_b_peij_2_3_n14), .ZN(pool_pool_pe_b_peij_2_3_n7) );
  AND2_X1 pool_pool_pe_b_peij_2_3_U8 ( .A1(pool_pool_pe_b_peij_2_3_d_acc[5]), 
        .A2(pool_pool_pe_b_peij_2_3_n14), .ZN(pool_pool_pe_b_peij_2_3_n6) );
  AND2_X1 pool_pool_pe_b_peij_2_3_U7 ( .A1(pool_pool_pe_b_peij_2_3_d_acc[6]), 
        .A2(pool_pool_pe_b_peij_2_3_n14), .ZN(pool_pool_pe_b_peij_2_3_n5) );
  AND2_X1 pool_pool_pe_b_peij_2_3_U6 ( .A1(pool_pool_pe_b_peij_2_3_d_acc[7]), 
        .A2(pool_pool_pe_b_peij_2_3_n14), .ZN(pool_pool_pe_b_peij_2_3_n4) );
  AND2_X1 pool_pool_pe_b_peij_2_3_U5 ( .A1(pool_pool_pe_b_peij_2_3_d_acc[8]), 
        .A2(pool_pool_pe_b_peij_2_3_n14), .ZN(pool_pool_pe_b_peij_2_3_n3) );
  AND2_X1 pool_pool_pe_b_peij_2_3_U4 ( .A1(pool_pool_pe_b_peij_2_3_d_acc[9]), 
        .A2(pool_pool_pe_b_peij_2_3_n14), .ZN(pool_pool_pe_b_peij_2_3_n2) );
  AND2_X1 pool_pool_pe_b_peij_2_3_U3 ( .A1(pool_pool_pe_b_peij_2_3_d_acc[10]), 
        .A2(pool_pool_pe_b_peij_2_3_n14), .ZN(pool_pool_pe_b_peij_2_3_n1) );
  DFFR_X1 pool_pool_pe_b_peij_2_3_q_acc_reg_10_ ( .D(
        pool_pool_pe_b_peij_2_3_n1), .CK(pool_pool_pe_b_peij_2_3_gck), .RN(
        pool_pool_pe_b_peij_2_3_n12), .Q(pool_pool_pe_b_o_data[54]) );
  DFFR_X1 pool_pool_pe_b_peij_2_3_q_acc_reg_9_ ( .D(pool_pool_pe_b_peij_2_3_n2), .CK(pool_pool_pe_b_peij_2_3_gck), .RN(pool_pool_pe_b_peij_2_3_n12), .Q(
        pool_pool_pe_b_o_data[53]) );
  DFFR_X1 pool_pool_pe_b_peij_2_3_q_acc_reg_8_ ( .D(pool_pool_pe_b_peij_2_3_n3), .CK(pool_pool_pe_b_peij_2_3_gck), .RN(pool_pool_pe_b_peij_2_3_n12), .Q(
        pool_pool_pe_b_o_data[52]) );
  DFFR_X1 pool_pool_pe_b_peij_2_3_q_acc_reg_7_ ( .D(pool_pool_pe_b_peij_2_3_n4), .CK(pool_pool_pe_b_peij_2_3_gck), .RN(pool_pool_pe_b_peij_2_3_n12), .Q(
        pool_pool_pe_b_o_data[51]) );
  DFFR_X1 pool_pool_pe_b_peij_2_3_q_acc_reg_6_ ( .D(pool_pool_pe_b_peij_2_3_n5), .CK(pool_pool_pe_b_peij_2_3_gck), .RN(pool_pool_pe_b_peij_2_3_n12), .Q(
        pool_pool_pe_b_o_data[50]) );
  DFFR_X1 pool_pool_pe_b_peij_2_3_q_acc_reg_5_ ( .D(pool_pool_pe_b_peij_2_3_n6), .CK(pool_pool_pe_b_peij_2_3_gck), .RN(pool_pool_pe_b_peij_2_3_n12), .Q(
        pool_pool_pe_b_o_data[49]) );
  DFFR_X1 pool_pool_pe_b_peij_2_3_q_acc_reg_4_ ( .D(pool_pool_pe_b_peij_2_3_n7), .CK(pool_pool_pe_b_peij_2_3_gck), .RN(pool_pool_pe_b_peij_2_3_n12), .Q(
        pool_pool_pe_b_o_data[48]) );
  DFFR_X1 pool_pool_pe_b_peij_2_3_q_acc_reg_3_ ( .D(pool_pool_pe_b_peij_2_3_n8), .CK(pool_pool_pe_b_peij_2_3_gck), .RN(pool_pool_pe_b_peij_2_3_n12), .Q(
        pool_pool_pe_b_o_data[47]) );
  DFFR_X1 pool_pool_pe_b_peij_2_3_q_acc_reg_2_ ( .D(pool_pool_pe_b_peij_2_3_n9), .CK(pool_pool_pe_b_peij_2_3_gck), .RN(pool_pool_pe_b_peij_2_3_n12), .Q(
        pool_pool_pe_b_o_data[46]) );
  DFFR_X1 pool_pool_pe_b_peij_2_3_q_acc_reg_1_ ( .D(
        pool_pool_pe_b_peij_2_3_n10), .CK(pool_pool_pe_b_peij_2_3_gck), .RN(
        pool_pool_pe_b_peij_2_3_n12), .Q(pool_pool_pe_b_o_data[45]) );
  DFFR_X1 pool_pool_pe_b_peij_2_3_q_acc_reg_0_ ( .D(
        pool_pool_pe_b_peij_2_3_n11), .CK(pool_pool_pe_b_peij_2_3_gck), .RN(
        pool_pool_pe_b_peij_2_3_n12), .Q(pool_pool_pe_b_o_data[44]) );
  AND3_X2 pool_pool_pe_b_peij_2_3_U20 ( .A1(pool_pool_pe_b_int_pe_en[4]), .A2(
        clk), .A3(1'b1), .ZN(pool_pool_pe_b_peij_2_3_gck) );
  SDFFR_X1 pool_pool_pe_b_peij_2_3_q_k_reg ( .D(1'b0), .SI(
        pool_pool_pe_b_peij_2_3_n14), .SE(1'b0), .CK(
        pool_pool_pe_b_peij_2_3_gck), .RN(pool_pool_pe_b_peij_2_3_n12), .Q(
        pool_pool_pe_b_peij_2_3_q_k) );
  XOR2_X1 pool_pool_pe_b_peij_2_3_add_U11 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_3_q_k), .Z(pool_pool_pe_b_peij_2_3_add_notb[0])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_3_add_U10 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_3_q_k), .Z(pool_pool_pe_b_peij_2_3_add_notb[10])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_3_add_U9 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_3_q_k), .Z(pool_pool_pe_b_peij_2_3_add_notb[1])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_3_add_U8 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_3_q_k), .Z(pool_pool_pe_b_peij_2_3_add_notb[2])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_3_add_U7 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_3_q_k), .Z(pool_pool_pe_b_peij_2_3_add_notb[3])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_3_add_U6 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_3_q_k), .Z(pool_pool_pe_b_peij_2_3_add_notb[4])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_3_add_U5 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_3_q_k), .Z(pool_pool_pe_b_peij_2_3_add_notb[5])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_3_add_U4 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_3_q_k), .Z(pool_pool_pe_b_peij_2_3_add_notb[6])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_3_add_U3 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_3_q_k), .Z(pool_pool_pe_b_peij_2_3_add_notb[7])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_3_add_U2 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_3_q_k), .Z(pool_pool_pe_b_peij_2_3_add_notb[8])
         );
  XOR2_X1 pool_pool_pe_b_peij_2_3_add_U1 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_2_3_q_k), .Z(pool_pool_pe_b_peij_2_3_add_notb[9])
         );
  INV_X2 pool_pool_pe_b_peij_2_3_add_fai_0_U2 ( .A(
        pool_pool_pe_b_peij_2_3_add_fai_0_n4), .ZN(
        pool_pool_pe_b_peij_2_3_add_cprop[1]) );
  XOR2_X1 pool_pool_pe_b_peij_2_3_add_fai_0_U4 ( .A(pool_pool_pe_b_o_data[44]), 
        .B(pool_pool_pe_b_peij_2_3_add_notb[0]), .Z(
        pool_pool_pe_b_peij_2_3_add_fai_0_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_3_add_fai_0_U3 ( .A(
        pool_pool_pe_b_peij_2_3_q_k), .B(pool_pool_pe_b_peij_2_3_add_fai_0_n5), 
        .Z(pool_pool_pe_b_peij_2_3_d_acc[0]) );
  AOI22_X2 pool_pool_pe_b_peij_2_3_add_fai_0_U1 ( .A1(
        pool_pool_pe_b_peij_2_3_add_notb[0]), .A2(pool_pool_pe_b_o_data[44]), 
        .B1(pool_pool_pe_b_peij_2_3_add_fai_0_n5), .B2(
        pool_pool_pe_b_peij_2_3_q_k), .ZN(pool_pool_pe_b_peij_2_3_add_fai_0_n4) );
  INV_X2 pool_pool_pe_b_peij_2_3_add_fai_1_U2 ( .A(
        pool_pool_pe_b_peij_2_3_add_fai_1_n4), .ZN(
        pool_pool_pe_b_peij_2_3_add_cprop[2]) );
  XOR2_X1 pool_pool_pe_b_peij_2_3_add_fai_1_U4 ( .A(pool_pool_pe_b_o_data[45]), 
        .B(pool_pool_pe_b_peij_2_3_add_notb[1]), .Z(
        pool_pool_pe_b_peij_2_3_add_fai_1_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_3_add_fai_1_U3 ( .A(
        pool_pool_pe_b_peij_2_3_add_cprop[1]), .B(
        pool_pool_pe_b_peij_2_3_add_fai_1_n5), .Z(
        pool_pool_pe_b_peij_2_3_d_acc[1]) );
  AOI22_X2 pool_pool_pe_b_peij_2_3_add_fai_1_U1 ( .A1(
        pool_pool_pe_b_peij_2_3_add_notb[1]), .A2(pool_pool_pe_b_o_data[45]), 
        .B1(pool_pool_pe_b_peij_2_3_add_fai_1_n5), .B2(
        pool_pool_pe_b_peij_2_3_add_cprop[1]), .ZN(
        pool_pool_pe_b_peij_2_3_add_fai_1_n4) );
  INV_X2 pool_pool_pe_b_peij_2_3_add_fai_2_U2 ( .A(
        pool_pool_pe_b_peij_2_3_add_fai_2_n4), .ZN(
        pool_pool_pe_b_peij_2_3_add_cprop[3]) );
  XOR2_X1 pool_pool_pe_b_peij_2_3_add_fai_2_U4 ( .A(pool_pool_pe_b_o_data[46]), 
        .B(pool_pool_pe_b_peij_2_3_add_notb[2]), .Z(
        pool_pool_pe_b_peij_2_3_add_fai_2_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_3_add_fai_2_U3 ( .A(
        pool_pool_pe_b_peij_2_3_add_cprop[2]), .B(
        pool_pool_pe_b_peij_2_3_add_fai_2_n5), .Z(
        pool_pool_pe_b_peij_2_3_d_acc[2]) );
  AOI22_X2 pool_pool_pe_b_peij_2_3_add_fai_2_U1 ( .A1(
        pool_pool_pe_b_peij_2_3_add_notb[2]), .A2(pool_pool_pe_b_o_data[46]), 
        .B1(pool_pool_pe_b_peij_2_3_add_fai_2_n5), .B2(
        pool_pool_pe_b_peij_2_3_add_cprop[2]), .ZN(
        pool_pool_pe_b_peij_2_3_add_fai_2_n4) );
  INV_X2 pool_pool_pe_b_peij_2_3_add_fai_3_U2 ( .A(
        pool_pool_pe_b_peij_2_3_add_fai_3_n4), .ZN(
        pool_pool_pe_b_peij_2_3_add_cprop[4]) );
  XOR2_X1 pool_pool_pe_b_peij_2_3_add_fai_3_U4 ( .A(pool_pool_pe_b_o_data[47]), 
        .B(pool_pool_pe_b_peij_2_3_add_notb[3]), .Z(
        pool_pool_pe_b_peij_2_3_add_fai_3_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_3_add_fai_3_U3 ( .A(
        pool_pool_pe_b_peij_2_3_add_cprop[3]), .B(
        pool_pool_pe_b_peij_2_3_add_fai_3_n5), .Z(
        pool_pool_pe_b_peij_2_3_d_acc[3]) );
  AOI22_X2 pool_pool_pe_b_peij_2_3_add_fai_3_U1 ( .A1(
        pool_pool_pe_b_peij_2_3_add_notb[3]), .A2(pool_pool_pe_b_o_data[47]), 
        .B1(pool_pool_pe_b_peij_2_3_add_fai_3_n5), .B2(
        pool_pool_pe_b_peij_2_3_add_cprop[3]), .ZN(
        pool_pool_pe_b_peij_2_3_add_fai_3_n4) );
  INV_X2 pool_pool_pe_b_peij_2_3_add_fai_4_U2 ( .A(
        pool_pool_pe_b_peij_2_3_add_fai_4_n4), .ZN(
        pool_pool_pe_b_peij_2_3_add_cprop[5]) );
  XOR2_X1 pool_pool_pe_b_peij_2_3_add_fai_4_U4 ( .A(pool_pool_pe_b_o_data[48]), 
        .B(pool_pool_pe_b_peij_2_3_add_notb[4]), .Z(
        pool_pool_pe_b_peij_2_3_add_fai_4_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_3_add_fai_4_U3 ( .A(
        pool_pool_pe_b_peij_2_3_add_cprop[4]), .B(
        pool_pool_pe_b_peij_2_3_add_fai_4_n5), .Z(
        pool_pool_pe_b_peij_2_3_d_acc[4]) );
  AOI22_X2 pool_pool_pe_b_peij_2_3_add_fai_4_U1 ( .A1(
        pool_pool_pe_b_peij_2_3_add_notb[4]), .A2(pool_pool_pe_b_o_data[48]), 
        .B1(pool_pool_pe_b_peij_2_3_add_fai_4_n5), .B2(
        pool_pool_pe_b_peij_2_3_add_cprop[4]), .ZN(
        pool_pool_pe_b_peij_2_3_add_fai_4_n4) );
  INV_X2 pool_pool_pe_b_peij_2_3_add_fai_5_U2 ( .A(
        pool_pool_pe_b_peij_2_3_add_fai_5_n4), .ZN(
        pool_pool_pe_b_peij_2_3_add_cprop[6]) );
  XOR2_X1 pool_pool_pe_b_peij_2_3_add_fai_5_U4 ( .A(pool_pool_pe_b_o_data[49]), 
        .B(pool_pool_pe_b_peij_2_3_add_notb[5]), .Z(
        pool_pool_pe_b_peij_2_3_add_fai_5_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_3_add_fai_5_U3 ( .A(
        pool_pool_pe_b_peij_2_3_add_cprop[5]), .B(
        pool_pool_pe_b_peij_2_3_add_fai_5_n5), .Z(
        pool_pool_pe_b_peij_2_3_d_acc[5]) );
  AOI22_X2 pool_pool_pe_b_peij_2_3_add_fai_5_U1 ( .A1(
        pool_pool_pe_b_peij_2_3_add_notb[5]), .A2(pool_pool_pe_b_o_data[49]), 
        .B1(pool_pool_pe_b_peij_2_3_add_fai_5_n5), .B2(
        pool_pool_pe_b_peij_2_3_add_cprop[5]), .ZN(
        pool_pool_pe_b_peij_2_3_add_fai_5_n4) );
  INV_X2 pool_pool_pe_b_peij_2_3_add_fai_6_U2 ( .A(
        pool_pool_pe_b_peij_2_3_add_fai_6_n4), .ZN(
        pool_pool_pe_b_peij_2_3_add_cprop[7]) );
  XOR2_X1 pool_pool_pe_b_peij_2_3_add_fai_6_U4 ( .A(pool_pool_pe_b_o_data[50]), 
        .B(pool_pool_pe_b_peij_2_3_add_notb[6]), .Z(
        pool_pool_pe_b_peij_2_3_add_fai_6_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_3_add_fai_6_U3 ( .A(
        pool_pool_pe_b_peij_2_3_add_cprop[6]), .B(
        pool_pool_pe_b_peij_2_3_add_fai_6_n5), .Z(
        pool_pool_pe_b_peij_2_3_d_acc[6]) );
  AOI22_X2 pool_pool_pe_b_peij_2_3_add_fai_6_U1 ( .A1(
        pool_pool_pe_b_peij_2_3_add_notb[6]), .A2(pool_pool_pe_b_o_data[50]), 
        .B1(pool_pool_pe_b_peij_2_3_add_fai_6_n5), .B2(
        pool_pool_pe_b_peij_2_3_add_cprop[6]), .ZN(
        pool_pool_pe_b_peij_2_3_add_fai_6_n4) );
  INV_X2 pool_pool_pe_b_peij_2_3_add_fai_7_U2 ( .A(
        pool_pool_pe_b_peij_2_3_add_fai_7_n4), .ZN(
        pool_pool_pe_b_peij_2_3_add_cprop[8]) );
  XOR2_X1 pool_pool_pe_b_peij_2_3_add_fai_7_U4 ( .A(pool_pool_pe_b_o_data[51]), 
        .B(pool_pool_pe_b_peij_2_3_add_notb[7]), .Z(
        pool_pool_pe_b_peij_2_3_add_fai_7_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_3_add_fai_7_U3 ( .A(
        pool_pool_pe_b_peij_2_3_add_cprop[7]), .B(
        pool_pool_pe_b_peij_2_3_add_fai_7_n5), .Z(
        pool_pool_pe_b_peij_2_3_d_acc[7]) );
  AOI22_X2 pool_pool_pe_b_peij_2_3_add_fai_7_U1 ( .A1(
        pool_pool_pe_b_peij_2_3_add_notb[7]), .A2(pool_pool_pe_b_o_data[51]), 
        .B1(pool_pool_pe_b_peij_2_3_add_fai_7_n5), .B2(
        pool_pool_pe_b_peij_2_3_add_cprop[7]), .ZN(
        pool_pool_pe_b_peij_2_3_add_fai_7_n4) );
  INV_X2 pool_pool_pe_b_peij_2_3_add_fai_8_U2 ( .A(
        pool_pool_pe_b_peij_2_3_add_fai_8_n4), .ZN(
        pool_pool_pe_b_peij_2_3_add_cprop[9]) );
  XOR2_X1 pool_pool_pe_b_peij_2_3_add_fai_8_U4 ( .A(pool_pool_pe_b_o_data[52]), 
        .B(pool_pool_pe_b_peij_2_3_add_notb[8]), .Z(
        pool_pool_pe_b_peij_2_3_add_fai_8_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_3_add_fai_8_U3 ( .A(
        pool_pool_pe_b_peij_2_3_add_cprop[8]), .B(
        pool_pool_pe_b_peij_2_3_add_fai_8_n5), .Z(
        pool_pool_pe_b_peij_2_3_d_acc[8]) );
  AOI22_X2 pool_pool_pe_b_peij_2_3_add_fai_8_U1 ( .A1(
        pool_pool_pe_b_peij_2_3_add_notb[8]), .A2(pool_pool_pe_b_o_data[52]), 
        .B1(pool_pool_pe_b_peij_2_3_add_fai_8_n5), .B2(
        pool_pool_pe_b_peij_2_3_add_cprop[8]), .ZN(
        pool_pool_pe_b_peij_2_3_add_fai_8_n4) );
  INV_X2 pool_pool_pe_b_peij_2_3_add_fai_9_U2 ( .A(
        pool_pool_pe_b_peij_2_3_add_fai_9_n4), .ZN(
        pool_pool_pe_b_peij_2_3_add_cprop[10]) );
  XOR2_X1 pool_pool_pe_b_peij_2_3_add_fai_9_U4 ( .A(pool_pool_pe_b_o_data[53]), 
        .B(pool_pool_pe_b_peij_2_3_add_notb[9]), .Z(
        pool_pool_pe_b_peij_2_3_add_fai_9_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_3_add_fai_9_U3 ( .A(
        pool_pool_pe_b_peij_2_3_add_cprop[9]), .B(
        pool_pool_pe_b_peij_2_3_add_fai_9_n5), .Z(
        pool_pool_pe_b_peij_2_3_d_acc[9]) );
  AOI22_X2 pool_pool_pe_b_peij_2_3_add_fai_9_U1 ( .A1(
        pool_pool_pe_b_peij_2_3_add_notb[9]), .A2(pool_pool_pe_b_o_data[53]), 
        .B1(pool_pool_pe_b_peij_2_3_add_fai_9_n5), .B2(
        pool_pool_pe_b_peij_2_3_add_cprop[9]), .ZN(
        pool_pool_pe_b_peij_2_3_add_fai_9_n4) );
  INV_X2 pool_pool_pe_b_peij_2_3_add_fai_10_U2 ( .A(
        pool_pool_pe_b_peij_2_3_add_fai_10_n4), .ZN(
        pool_pool_pe_b_peij_2_3_add_c_out) );
  XOR2_X1 pool_pool_pe_b_peij_2_3_add_fai_10_U4 ( .A(pool_pool_pe_b_o_data[54]), .B(pool_pool_pe_b_peij_2_3_add_notb[10]), .Z(
        pool_pool_pe_b_peij_2_3_add_fai_10_n5) );
  XOR2_X1 pool_pool_pe_b_peij_2_3_add_fai_10_U3 ( .A(
        pool_pool_pe_b_peij_2_3_add_cprop[10]), .B(
        pool_pool_pe_b_peij_2_3_add_fai_10_n5), .Z(
        pool_pool_pe_b_peij_2_3_d_acc[10]) );
  AOI22_X2 pool_pool_pe_b_peij_2_3_add_fai_10_U1 ( .A1(
        pool_pool_pe_b_peij_2_3_add_notb[10]), .A2(pool_pool_pe_b_o_data[54]), 
        .B1(pool_pool_pe_b_peij_2_3_add_fai_10_n5), .B2(
        pool_pool_pe_b_peij_2_3_add_cprop[10]), .ZN(
        pool_pool_pe_b_peij_2_3_add_fai_10_n4) );
  INV_X2 pool_pool_pe_b_peij_3_0_U21 ( .A(pool_sync_clr), .ZN(
        pool_pool_pe_b_peij_3_0_n14) );
  INV_X1 pool_pool_pe_b_peij_3_0_U18 ( .A(pool_pool_pe_b_n1), .ZN(
        pool_pool_pe_b_peij_3_0_n12) );
  AND2_X1 pool_pool_pe_b_peij_3_0_U13 ( .A1(pool_pool_pe_b_peij_3_0_d_acc[0]), 
        .A2(pool_pool_pe_b_peij_3_0_n14), .ZN(pool_pool_pe_b_peij_3_0_n11) );
  AND2_X1 pool_pool_pe_b_peij_3_0_U12 ( .A1(pool_pool_pe_b_peij_3_0_d_acc[1]), 
        .A2(pool_pool_pe_b_peij_3_0_n14), .ZN(pool_pool_pe_b_peij_3_0_n10) );
  AND2_X1 pool_pool_pe_b_peij_3_0_U11 ( .A1(pool_pool_pe_b_peij_3_0_d_acc[2]), 
        .A2(pool_pool_pe_b_peij_3_0_n14), .ZN(pool_pool_pe_b_peij_3_0_n9) );
  AND2_X1 pool_pool_pe_b_peij_3_0_U10 ( .A1(pool_pool_pe_b_peij_3_0_d_acc[3]), 
        .A2(pool_pool_pe_b_peij_3_0_n14), .ZN(pool_pool_pe_b_peij_3_0_n8) );
  AND2_X1 pool_pool_pe_b_peij_3_0_U9 ( .A1(pool_pool_pe_b_peij_3_0_d_acc[4]), 
        .A2(pool_pool_pe_b_peij_3_0_n14), .ZN(pool_pool_pe_b_peij_3_0_n7) );
  AND2_X1 pool_pool_pe_b_peij_3_0_U8 ( .A1(pool_pool_pe_b_peij_3_0_d_acc[5]), 
        .A2(pool_pool_pe_b_peij_3_0_n14), .ZN(pool_pool_pe_b_peij_3_0_n6) );
  AND2_X1 pool_pool_pe_b_peij_3_0_U7 ( .A1(pool_pool_pe_b_peij_3_0_d_acc[6]), 
        .A2(pool_pool_pe_b_peij_3_0_n14), .ZN(pool_pool_pe_b_peij_3_0_n5) );
  AND2_X1 pool_pool_pe_b_peij_3_0_U6 ( .A1(pool_pool_pe_b_peij_3_0_d_acc[7]), 
        .A2(pool_pool_pe_b_peij_3_0_n14), .ZN(pool_pool_pe_b_peij_3_0_n4) );
  AND2_X1 pool_pool_pe_b_peij_3_0_U5 ( .A1(pool_pool_pe_b_peij_3_0_d_acc[8]), 
        .A2(pool_pool_pe_b_peij_3_0_n14), .ZN(pool_pool_pe_b_peij_3_0_n3) );
  AND2_X1 pool_pool_pe_b_peij_3_0_U4 ( .A1(pool_pool_pe_b_peij_3_0_d_acc[9]), 
        .A2(pool_pool_pe_b_peij_3_0_n14), .ZN(pool_pool_pe_b_peij_3_0_n2) );
  AND2_X1 pool_pool_pe_b_peij_3_0_U3 ( .A1(pool_pool_pe_b_peij_3_0_d_acc[10]), 
        .A2(pool_pool_pe_b_peij_3_0_n14), .ZN(pool_pool_pe_b_peij_3_0_n1) );
  DFFR_X1 pool_pool_pe_b_peij_3_0_q_acc_reg_10_ ( .D(
        pool_pool_pe_b_peij_3_0_n1), .CK(pool_pool_pe_b_peij_3_0_gck), .RN(
        pool_pool_pe_b_peij_3_0_n12), .Q(pool_pool_pe_b_o_data[43]) );
  DFFR_X1 pool_pool_pe_b_peij_3_0_q_acc_reg_9_ ( .D(pool_pool_pe_b_peij_3_0_n2), .CK(pool_pool_pe_b_peij_3_0_gck), .RN(pool_pool_pe_b_peij_3_0_n12), .Q(
        pool_pool_pe_b_o_data[42]) );
  DFFR_X1 pool_pool_pe_b_peij_3_0_q_acc_reg_8_ ( .D(pool_pool_pe_b_peij_3_0_n3), .CK(pool_pool_pe_b_peij_3_0_gck), .RN(pool_pool_pe_b_peij_3_0_n12), .Q(
        pool_pool_pe_b_o_data[41]) );
  DFFR_X1 pool_pool_pe_b_peij_3_0_q_acc_reg_7_ ( .D(pool_pool_pe_b_peij_3_0_n4), .CK(pool_pool_pe_b_peij_3_0_gck), .RN(pool_pool_pe_b_peij_3_0_n12), .Q(
        pool_pool_pe_b_o_data[40]) );
  DFFR_X1 pool_pool_pe_b_peij_3_0_q_acc_reg_6_ ( .D(pool_pool_pe_b_peij_3_0_n5), .CK(pool_pool_pe_b_peij_3_0_gck), .RN(pool_pool_pe_b_peij_3_0_n12), .Q(
        pool_pool_pe_b_o_data[39]) );
  DFFR_X1 pool_pool_pe_b_peij_3_0_q_acc_reg_5_ ( .D(pool_pool_pe_b_peij_3_0_n6), .CK(pool_pool_pe_b_peij_3_0_gck), .RN(pool_pool_pe_b_peij_3_0_n12), .Q(
        pool_pool_pe_b_o_data[38]) );
  DFFR_X1 pool_pool_pe_b_peij_3_0_q_acc_reg_4_ ( .D(pool_pool_pe_b_peij_3_0_n7), .CK(pool_pool_pe_b_peij_3_0_gck), .RN(pool_pool_pe_b_peij_3_0_n12), .Q(
        pool_pool_pe_b_o_data[37]) );
  DFFR_X1 pool_pool_pe_b_peij_3_0_q_acc_reg_3_ ( .D(pool_pool_pe_b_peij_3_0_n8), .CK(pool_pool_pe_b_peij_3_0_gck), .RN(pool_pool_pe_b_peij_3_0_n12), .Q(
        pool_pool_pe_b_o_data[36]) );
  DFFR_X1 pool_pool_pe_b_peij_3_0_q_acc_reg_2_ ( .D(pool_pool_pe_b_peij_3_0_n9), .CK(pool_pool_pe_b_peij_3_0_gck), .RN(pool_pool_pe_b_peij_3_0_n12), .Q(
        pool_pool_pe_b_o_data[35]) );
  DFFR_X1 pool_pool_pe_b_peij_3_0_q_acc_reg_1_ ( .D(
        pool_pool_pe_b_peij_3_0_n10), .CK(pool_pool_pe_b_peij_3_0_gck), .RN(
        pool_pool_pe_b_peij_3_0_n12), .Q(pool_pool_pe_b_o_data[34]) );
  DFFR_X1 pool_pool_pe_b_peij_3_0_q_acc_reg_0_ ( .D(
        pool_pool_pe_b_peij_3_0_n11), .CK(pool_pool_pe_b_peij_3_0_gck), .RN(
        pool_pool_pe_b_peij_3_0_n12), .Q(pool_pool_pe_b_o_data[33]) );
  AND3_X2 pool_pool_pe_b_peij_3_0_U20 ( .A1(pool_pool_pe_b_int_pe_en[3]), .A2(
        clk), .A3(1'b1), .ZN(pool_pool_pe_b_peij_3_0_gck) );
  SDFFR_X1 pool_pool_pe_b_peij_3_0_q_k_reg ( .D(1'b0), .SI(
        pool_pool_pe_b_peij_3_0_n14), .SE(1'b0), .CK(
        pool_pool_pe_b_peij_3_0_gck), .RN(pool_pool_pe_b_peij_3_0_n12), .Q(
        pool_pool_pe_b_peij_3_0_q_k) );
  XOR2_X1 pool_pool_pe_b_peij_3_0_add_U11 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_0_q_k), .Z(pool_pool_pe_b_peij_3_0_add_notb[0])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_0_add_U10 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_0_q_k), .Z(pool_pool_pe_b_peij_3_0_add_notb[10])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_0_add_U9 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_0_q_k), .Z(pool_pool_pe_b_peij_3_0_add_notb[1])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_0_add_U8 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_0_q_k), .Z(pool_pool_pe_b_peij_3_0_add_notb[2])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_0_add_U7 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_0_q_k), .Z(pool_pool_pe_b_peij_3_0_add_notb[3])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_0_add_U6 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_0_q_k), .Z(pool_pool_pe_b_peij_3_0_add_notb[4])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_0_add_U5 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_0_q_k), .Z(pool_pool_pe_b_peij_3_0_add_notb[5])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_0_add_U4 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_0_q_k), .Z(pool_pool_pe_b_peij_3_0_add_notb[6])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_0_add_U3 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_0_q_k), .Z(pool_pool_pe_b_peij_3_0_add_notb[7])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_0_add_U2 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_0_q_k), .Z(pool_pool_pe_b_peij_3_0_add_notb[8])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_0_add_U1 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_0_q_k), .Z(pool_pool_pe_b_peij_3_0_add_notb[9])
         );
  INV_X2 pool_pool_pe_b_peij_3_0_add_fai_0_U2 ( .A(
        pool_pool_pe_b_peij_3_0_add_fai_0_n4), .ZN(
        pool_pool_pe_b_peij_3_0_add_cprop[1]) );
  XOR2_X1 pool_pool_pe_b_peij_3_0_add_fai_0_U4 ( .A(pool_pool_pe_b_o_data[33]), 
        .B(pool_pool_pe_b_peij_3_0_add_notb[0]), .Z(
        pool_pool_pe_b_peij_3_0_add_fai_0_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_0_add_fai_0_U3 ( .A(
        pool_pool_pe_b_peij_3_0_q_k), .B(pool_pool_pe_b_peij_3_0_add_fai_0_n5), 
        .Z(pool_pool_pe_b_peij_3_0_d_acc[0]) );
  AOI22_X2 pool_pool_pe_b_peij_3_0_add_fai_0_U1 ( .A1(
        pool_pool_pe_b_peij_3_0_add_notb[0]), .A2(pool_pool_pe_b_o_data[33]), 
        .B1(pool_pool_pe_b_peij_3_0_add_fai_0_n5), .B2(
        pool_pool_pe_b_peij_3_0_q_k), .ZN(pool_pool_pe_b_peij_3_0_add_fai_0_n4) );
  INV_X2 pool_pool_pe_b_peij_3_0_add_fai_1_U2 ( .A(
        pool_pool_pe_b_peij_3_0_add_fai_1_n4), .ZN(
        pool_pool_pe_b_peij_3_0_add_cprop[2]) );
  XOR2_X1 pool_pool_pe_b_peij_3_0_add_fai_1_U4 ( .A(pool_pool_pe_b_o_data[34]), 
        .B(pool_pool_pe_b_peij_3_0_add_notb[1]), .Z(
        pool_pool_pe_b_peij_3_0_add_fai_1_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_0_add_fai_1_U3 ( .A(
        pool_pool_pe_b_peij_3_0_add_cprop[1]), .B(
        pool_pool_pe_b_peij_3_0_add_fai_1_n5), .Z(
        pool_pool_pe_b_peij_3_0_d_acc[1]) );
  AOI22_X2 pool_pool_pe_b_peij_3_0_add_fai_1_U1 ( .A1(
        pool_pool_pe_b_peij_3_0_add_notb[1]), .A2(pool_pool_pe_b_o_data[34]), 
        .B1(pool_pool_pe_b_peij_3_0_add_fai_1_n5), .B2(
        pool_pool_pe_b_peij_3_0_add_cprop[1]), .ZN(
        pool_pool_pe_b_peij_3_0_add_fai_1_n4) );
  INV_X2 pool_pool_pe_b_peij_3_0_add_fai_2_U2 ( .A(
        pool_pool_pe_b_peij_3_0_add_fai_2_n4), .ZN(
        pool_pool_pe_b_peij_3_0_add_cprop[3]) );
  XOR2_X1 pool_pool_pe_b_peij_3_0_add_fai_2_U4 ( .A(pool_pool_pe_b_o_data[35]), 
        .B(pool_pool_pe_b_peij_3_0_add_notb[2]), .Z(
        pool_pool_pe_b_peij_3_0_add_fai_2_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_0_add_fai_2_U3 ( .A(
        pool_pool_pe_b_peij_3_0_add_cprop[2]), .B(
        pool_pool_pe_b_peij_3_0_add_fai_2_n5), .Z(
        pool_pool_pe_b_peij_3_0_d_acc[2]) );
  AOI22_X2 pool_pool_pe_b_peij_3_0_add_fai_2_U1 ( .A1(
        pool_pool_pe_b_peij_3_0_add_notb[2]), .A2(pool_pool_pe_b_o_data[35]), 
        .B1(pool_pool_pe_b_peij_3_0_add_fai_2_n5), .B2(
        pool_pool_pe_b_peij_3_0_add_cprop[2]), .ZN(
        pool_pool_pe_b_peij_3_0_add_fai_2_n4) );
  INV_X2 pool_pool_pe_b_peij_3_0_add_fai_3_U2 ( .A(
        pool_pool_pe_b_peij_3_0_add_fai_3_n4), .ZN(
        pool_pool_pe_b_peij_3_0_add_cprop[4]) );
  XOR2_X1 pool_pool_pe_b_peij_3_0_add_fai_3_U4 ( .A(pool_pool_pe_b_o_data[36]), 
        .B(pool_pool_pe_b_peij_3_0_add_notb[3]), .Z(
        pool_pool_pe_b_peij_3_0_add_fai_3_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_0_add_fai_3_U3 ( .A(
        pool_pool_pe_b_peij_3_0_add_cprop[3]), .B(
        pool_pool_pe_b_peij_3_0_add_fai_3_n5), .Z(
        pool_pool_pe_b_peij_3_0_d_acc[3]) );
  AOI22_X2 pool_pool_pe_b_peij_3_0_add_fai_3_U1 ( .A1(
        pool_pool_pe_b_peij_3_0_add_notb[3]), .A2(pool_pool_pe_b_o_data[36]), 
        .B1(pool_pool_pe_b_peij_3_0_add_fai_3_n5), .B2(
        pool_pool_pe_b_peij_3_0_add_cprop[3]), .ZN(
        pool_pool_pe_b_peij_3_0_add_fai_3_n4) );
  INV_X2 pool_pool_pe_b_peij_3_0_add_fai_4_U2 ( .A(
        pool_pool_pe_b_peij_3_0_add_fai_4_n4), .ZN(
        pool_pool_pe_b_peij_3_0_add_cprop[5]) );
  XOR2_X1 pool_pool_pe_b_peij_3_0_add_fai_4_U4 ( .A(pool_pool_pe_b_o_data[37]), 
        .B(pool_pool_pe_b_peij_3_0_add_notb[4]), .Z(
        pool_pool_pe_b_peij_3_0_add_fai_4_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_0_add_fai_4_U3 ( .A(
        pool_pool_pe_b_peij_3_0_add_cprop[4]), .B(
        pool_pool_pe_b_peij_3_0_add_fai_4_n5), .Z(
        pool_pool_pe_b_peij_3_0_d_acc[4]) );
  AOI22_X2 pool_pool_pe_b_peij_3_0_add_fai_4_U1 ( .A1(
        pool_pool_pe_b_peij_3_0_add_notb[4]), .A2(pool_pool_pe_b_o_data[37]), 
        .B1(pool_pool_pe_b_peij_3_0_add_fai_4_n5), .B2(
        pool_pool_pe_b_peij_3_0_add_cprop[4]), .ZN(
        pool_pool_pe_b_peij_3_0_add_fai_4_n4) );
  INV_X2 pool_pool_pe_b_peij_3_0_add_fai_5_U2 ( .A(
        pool_pool_pe_b_peij_3_0_add_fai_5_n4), .ZN(
        pool_pool_pe_b_peij_3_0_add_cprop[6]) );
  XOR2_X1 pool_pool_pe_b_peij_3_0_add_fai_5_U4 ( .A(pool_pool_pe_b_o_data[38]), 
        .B(pool_pool_pe_b_peij_3_0_add_notb[5]), .Z(
        pool_pool_pe_b_peij_3_0_add_fai_5_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_0_add_fai_5_U3 ( .A(
        pool_pool_pe_b_peij_3_0_add_cprop[5]), .B(
        pool_pool_pe_b_peij_3_0_add_fai_5_n5), .Z(
        pool_pool_pe_b_peij_3_0_d_acc[5]) );
  AOI22_X2 pool_pool_pe_b_peij_3_0_add_fai_5_U1 ( .A1(
        pool_pool_pe_b_peij_3_0_add_notb[5]), .A2(pool_pool_pe_b_o_data[38]), 
        .B1(pool_pool_pe_b_peij_3_0_add_fai_5_n5), .B2(
        pool_pool_pe_b_peij_3_0_add_cprop[5]), .ZN(
        pool_pool_pe_b_peij_3_0_add_fai_5_n4) );
  INV_X2 pool_pool_pe_b_peij_3_0_add_fai_6_U2 ( .A(
        pool_pool_pe_b_peij_3_0_add_fai_6_n4), .ZN(
        pool_pool_pe_b_peij_3_0_add_cprop[7]) );
  XOR2_X1 pool_pool_pe_b_peij_3_0_add_fai_6_U4 ( .A(pool_pool_pe_b_o_data[39]), 
        .B(pool_pool_pe_b_peij_3_0_add_notb[6]), .Z(
        pool_pool_pe_b_peij_3_0_add_fai_6_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_0_add_fai_6_U3 ( .A(
        pool_pool_pe_b_peij_3_0_add_cprop[6]), .B(
        pool_pool_pe_b_peij_3_0_add_fai_6_n5), .Z(
        pool_pool_pe_b_peij_3_0_d_acc[6]) );
  AOI22_X2 pool_pool_pe_b_peij_3_0_add_fai_6_U1 ( .A1(
        pool_pool_pe_b_peij_3_0_add_notb[6]), .A2(pool_pool_pe_b_o_data[39]), 
        .B1(pool_pool_pe_b_peij_3_0_add_fai_6_n5), .B2(
        pool_pool_pe_b_peij_3_0_add_cprop[6]), .ZN(
        pool_pool_pe_b_peij_3_0_add_fai_6_n4) );
  INV_X2 pool_pool_pe_b_peij_3_0_add_fai_7_U2 ( .A(
        pool_pool_pe_b_peij_3_0_add_fai_7_n4), .ZN(
        pool_pool_pe_b_peij_3_0_add_cprop[8]) );
  XOR2_X1 pool_pool_pe_b_peij_3_0_add_fai_7_U4 ( .A(pool_pool_pe_b_o_data[40]), 
        .B(pool_pool_pe_b_peij_3_0_add_notb[7]), .Z(
        pool_pool_pe_b_peij_3_0_add_fai_7_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_0_add_fai_7_U3 ( .A(
        pool_pool_pe_b_peij_3_0_add_cprop[7]), .B(
        pool_pool_pe_b_peij_3_0_add_fai_7_n5), .Z(
        pool_pool_pe_b_peij_3_0_d_acc[7]) );
  AOI22_X2 pool_pool_pe_b_peij_3_0_add_fai_7_U1 ( .A1(
        pool_pool_pe_b_peij_3_0_add_notb[7]), .A2(pool_pool_pe_b_o_data[40]), 
        .B1(pool_pool_pe_b_peij_3_0_add_fai_7_n5), .B2(
        pool_pool_pe_b_peij_3_0_add_cprop[7]), .ZN(
        pool_pool_pe_b_peij_3_0_add_fai_7_n4) );
  INV_X2 pool_pool_pe_b_peij_3_0_add_fai_8_U2 ( .A(
        pool_pool_pe_b_peij_3_0_add_fai_8_n4), .ZN(
        pool_pool_pe_b_peij_3_0_add_cprop[9]) );
  XOR2_X1 pool_pool_pe_b_peij_3_0_add_fai_8_U4 ( .A(pool_pool_pe_b_o_data[41]), 
        .B(pool_pool_pe_b_peij_3_0_add_notb[8]), .Z(
        pool_pool_pe_b_peij_3_0_add_fai_8_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_0_add_fai_8_U3 ( .A(
        pool_pool_pe_b_peij_3_0_add_cprop[8]), .B(
        pool_pool_pe_b_peij_3_0_add_fai_8_n5), .Z(
        pool_pool_pe_b_peij_3_0_d_acc[8]) );
  AOI22_X2 pool_pool_pe_b_peij_3_0_add_fai_8_U1 ( .A1(
        pool_pool_pe_b_peij_3_0_add_notb[8]), .A2(pool_pool_pe_b_o_data[41]), 
        .B1(pool_pool_pe_b_peij_3_0_add_fai_8_n5), .B2(
        pool_pool_pe_b_peij_3_0_add_cprop[8]), .ZN(
        pool_pool_pe_b_peij_3_0_add_fai_8_n4) );
  INV_X2 pool_pool_pe_b_peij_3_0_add_fai_9_U2 ( .A(
        pool_pool_pe_b_peij_3_0_add_fai_9_n4), .ZN(
        pool_pool_pe_b_peij_3_0_add_cprop[10]) );
  XOR2_X1 pool_pool_pe_b_peij_3_0_add_fai_9_U4 ( .A(pool_pool_pe_b_o_data[42]), 
        .B(pool_pool_pe_b_peij_3_0_add_notb[9]), .Z(
        pool_pool_pe_b_peij_3_0_add_fai_9_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_0_add_fai_9_U3 ( .A(
        pool_pool_pe_b_peij_3_0_add_cprop[9]), .B(
        pool_pool_pe_b_peij_3_0_add_fai_9_n5), .Z(
        pool_pool_pe_b_peij_3_0_d_acc[9]) );
  AOI22_X2 pool_pool_pe_b_peij_3_0_add_fai_9_U1 ( .A1(
        pool_pool_pe_b_peij_3_0_add_notb[9]), .A2(pool_pool_pe_b_o_data[42]), 
        .B1(pool_pool_pe_b_peij_3_0_add_fai_9_n5), .B2(
        pool_pool_pe_b_peij_3_0_add_cprop[9]), .ZN(
        pool_pool_pe_b_peij_3_0_add_fai_9_n4) );
  INV_X2 pool_pool_pe_b_peij_3_0_add_fai_10_U2 ( .A(
        pool_pool_pe_b_peij_3_0_add_fai_10_n4), .ZN(
        pool_pool_pe_b_peij_3_0_add_c_out) );
  XOR2_X1 pool_pool_pe_b_peij_3_0_add_fai_10_U4 ( .A(pool_pool_pe_b_o_data[43]), .B(pool_pool_pe_b_peij_3_0_add_notb[10]), .Z(
        pool_pool_pe_b_peij_3_0_add_fai_10_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_0_add_fai_10_U3 ( .A(
        pool_pool_pe_b_peij_3_0_add_cprop[10]), .B(
        pool_pool_pe_b_peij_3_0_add_fai_10_n5), .Z(
        pool_pool_pe_b_peij_3_0_d_acc[10]) );
  AOI22_X2 pool_pool_pe_b_peij_3_0_add_fai_10_U1 ( .A1(
        pool_pool_pe_b_peij_3_0_add_notb[10]), .A2(pool_pool_pe_b_o_data[43]), 
        .B1(pool_pool_pe_b_peij_3_0_add_fai_10_n5), .B2(
        pool_pool_pe_b_peij_3_0_add_cprop[10]), .ZN(
        pool_pool_pe_b_peij_3_0_add_fai_10_n4) );
  INV_X2 pool_pool_pe_b_peij_3_1_U21 ( .A(pool_sync_clr), .ZN(
        pool_pool_pe_b_peij_3_1_n14) );
  INV_X1 pool_pool_pe_b_peij_3_1_U18 ( .A(pool_pool_pe_b_n1), .ZN(
        pool_pool_pe_b_peij_3_1_n12) );
  AND2_X1 pool_pool_pe_b_peij_3_1_U13 ( .A1(pool_pool_pe_b_peij_3_1_d_acc[0]), 
        .A2(pool_pool_pe_b_peij_3_1_n14), .ZN(pool_pool_pe_b_peij_3_1_n11) );
  AND2_X1 pool_pool_pe_b_peij_3_1_U12 ( .A1(pool_pool_pe_b_peij_3_1_d_acc[1]), 
        .A2(pool_pool_pe_b_peij_3_1_n14), .ZN(pool_pool_pe_b_peij_3_1_n10) );
  AND2_X1 pool_pool_pe_b_peij_3_1_U11 ( .A1(pool_pool_pe_b_peij_3_1_d_acc[2]), 
        .A2(pool_pool_pe_b_peij_3_1_n14), .ZN(pool_pool_pe_b_peij_3_1_n9) );
  AND2_X1 pool_pool_pe_b_peij_3_1_U10 ( .A1(pool_pool_pe_b_peij_3_1_d_acc[3]), 
        .A2(pool_pool_pe_b_peij_3_1_n14), .ZN(pool_pool_pe_b_peij_3_1_n8) );
  AND2_X1 pool_pool_pe_b_peij_3_1_U9 ( .A1(pool_pool_pe_b_peij_3_1_d_acc[4]), 
        .A2(pool_pool_pe_b_peij_3_1_n14), .ZN(pool_pool_pe_b_peij_3_1_n7) );
  AND2_X1 pool_pool_pe_b_peij_3_1_U8 ( .A1(pool_pool_pe_b_peij_3_1_d_acc[5]), 
        .A2(pool_pool_pe_b_peij_3_1_n14), .ZN(pool_pool_pe_b_peij_3_1_n6) );
  AND2_X1 pool_pool_pe_b_peij_3_1_U7 ( .A1(pool_pool_pe_b_peij_3_1_d_acc[6]), 
        .A2(pool_pool_pe_b_peij_3_1_n14), .ZN(pool_pool_pe_b_peij_3_1_n5) );
  AND2_X1 pool_pool_pe_b_peij_3_1_U6 ( .A1(pool_pool_pe_b_peij_3_1_d_acc[7]), 
        .A2(pool_pool_pe_b_peij_3_1_n14), .ZN(pool_pool_pe_b_peij_3_1_n4) );
  AND2_X1 pool_pool_pe_b_peij_3_1_U5 ( .A1(pool_pool_pe_b_peij_3_1_d_acc[8]), 
        .A2(pool_pool_pe_b_peij_3_1_n14), .ZN(pool_pool_pe_b_peij_3_1_n3) );
  AND2_X1 pool_pool_pe_b_peij_3_1_U4 ( .A1(pool_pool_pe_b_peij_3_1_d_acc[9]), 
        .A2(pool_pool_pe_b_peij_3_1_n14), .ZN(pool_pool_pe_b_peij_3_1_n2) );
  AND2_X1 pool_pool_pe_b_peij_3_1_U3 ( .A1(pool_pool_pe_b_peij_3_1_d_acc[10]), 
        .A2(pool_pool_pe_b_peij_3_1_n14), .ZN(pool_pool_pe_b_peij_3_1_n1) );
  DFFR_X1 pool_pool_pe_b_peij_3_1_q_acc_reg_10_ ( .D(
        pool_pool_pe_b_peij_3_1_n1), .CK(pool_pool_pe_b_peij_3_1_gck), .RN(
        pool_pool_pe_b_peij_3_1_n12), .Q(pool_pool_pe_b_o_data[32]) );
  DFFR_X1 pool_pool_pe_b_peij_3_1_q_acc_reg_9_ ( .D(pool_pool_pe_b_peij_3_1_n2), .CK(pool_pool_pe_b_peij_3_1_gck), .RN(pool_pool_pe_b_peij_3_1_n12), .Q(
        pool_pool_pe_b_o_data[31]) );
  DFFR_X1 pool_pool_pe_b_peij_3_1_q_acc_reg_8_ ( .D(pool_pool_pe_b_peij_3_1_n3), .CK(pool_pool_pe_b_peij_3_1_gck), .RN(pool_pool_pe_b_peij_3_1_n12), .Q(
        pool_pool_pe_b_o_data[30]) );
  DFFR_X1 pool_pool_pe_b_peij_3_1_q_acc_reg_7_ ( .D(pool_pool_pe_b_peij_3_1_n4), .CK(pool_pool_pe_b_peij_3_1_gck), .RN(pool_pool_pe_b_peij_3_1_n12), .Q(
        pool_pool_pe_b_o_data[29]) );
  DFFR_X1 pool_pool_pe_b_peij_3_1_q_acc_reg_6_ ( .D(pool_pool_pe_b_peij_3_1_n5), .CK(pool_pool_pe_b_peij_3_1_gck), .RN(pool_pool_pe_b_peij_3_1_n12), .Q(
        pool_pool_pe_b_o_data[28]) );
  DFFR_X1 pool_pool_pe_b_peij_3_1_q_acc_reg_5_ ( .D(pool_pool_pe_b_peij_3_1_n6), .CK(pool_pool_pe_b_peij_3_1_gck), .RN(pool_pool_pe_b_peij_3_1_n12), .Q(
        pool_pool_pe_b_o_data[27]) );
  DFFR_X1 pool_pool_pe_b_peij_3_1_q_acc_reg_4_ ( .D(pool_pool_pe_b_peij_3_1_n7), .CK(pool_pool_pe_b_peij_3_1_gck), .RN(pool_pool_pe_b_peij_3_1_n12), .Q(
        pool_pool_pe_b_o_data[26]) );
  DFFR_X1 pool_pool_pe_b_peij_3_1_q_acc_reg_3_ ( .D(pool_pool_pe_b_peij_3_1_n8), .CK(pool_pool_pe_b_peij_3_1_gck), .RN(pool_pool_pe_b_peij_3_1_n12), .Q(
        pool_pool_pe_b_o_data[25]) );
  DFFR_X1 pool_pool_pe_b_peij_3_1_q_acc_reg_2_ ( .D(pool_pool_pe_b_peij_3_1_n9), .CK(pool_pool_pe_b_peij_3_1_gck), .RN(pool_pool_pe_b_peij_3_1_n12), .Q(
        pool_pool_pe_b_o_data[24]) );
  DFFR_X1 pool_pool_pe_b_peij_3_1_q_acc_reg_1_ ( .D(
        pool_pool_pe_b_peij_3_1_n10), .CK(pool_pool_pe_b_peij_3_1_gck), .RN(
        pool_pool_pe_b_peij_3_1_n12), .Q(pool_pool_pe_b_o_data[23]) );
  DFFR_X1 pool_pool_pe_b_peij_3_1_q_acc_reg_0_ ( .D(
        pool_pool_pe_b_peij_3_1_n11), .CK(pool_pool_pe_b_peij_3_1_gck), .RN(
        pool_pool_pe_b_peij_3_1_n12), .Q(pool_pool_pe_b_o_data[22]) );
  AND3_X2 pool_pool_pe_b_peij_3_1_U20 ( .A1(pool_pool_pe_b_int_pe_en[2]), .A2(
        clk), .A3(1'b1), .ZN(pool_pool_pe_b_peij_3_1_gck) );
  SDFFR_X1 pool_pool_pe_b_peij_3_1_q_k_reg ( .D(1'b0), .SI(
        pool_pool_pe_b_peij_3_1_n14), .SE(1'b0), .CK(
        pool_pool_pe_b_peij_3_1_gck), .RN(pool_pool_pe_b_peij_3_1_n12), .Q(
        pool_pool_pe_b_peij_3_1_q_k) );
  XOR2_X1 pool_pool_pe_b_peij_3_1_add_U11 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_1_q_k), .Z(pool_pool_pe_b_peij_3_1_add_notb[0])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_1_add_U10 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_1_q_k), .Z(pool_pool_pe_b_peij_3_1_add_notb[10])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_1_add_U9 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_1_q_k), .Z(pool_pool_pe_b_peij_3_1_add_notb[1])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_1_add_U8 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_1_q_k), .Z(pool_pool_pe_b_peij_3_1_add_notb[2])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_1_add_U7 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_1_q_k), .Z(pool_pool_pe_b_peij_3_1_add_notb[3])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_1_add_U6 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_1_q_k), .Z(pool_pool_pe_b_peij_3_1_add_notb[4])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_1_add_U5 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_1_q_k), .Z(pool_pool_pe_b_peij_3_1_add_notb[5])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_1_add_U4 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_1_q_k), .Z(pool_pool_pe_b_peij_3_1_add_notb[6])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_1_add_U3 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_1_q_k), .Z(pool_pool_pe_b_peij_3_1_add_notb[7])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_1_add_U2 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_1_q_k), .Z(pool_pool_pe_b_peij_3_1_add_notb[8])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_1_add_U1 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_1_q_k), .Z(pool_pool_pe_b_peij_3_1_add_notb[9])
         );
  INV_X2 pool_pool_pe_b_peij_3_1_add_fai_0_U2 ( .A(
        pool_pool_pe_b_peij_3_1_add_fai_0_n4), .ZN(
        pool_pool_pe_b_peij_3_1_add_cprop[1]) );
  XOR2_X1 pool_pool_pe_b_peij_3_1_add_fai_0_U4 ( .A(pool_pool_pe_b_o_data[22]), 
        .B(pool_pool_pe_b_peij_3_1_add_notb[0]), .Z(
        pool_pool_pe_b_peij_3_1_add_fai_0_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_1_add_fai_0_U3 ( .A(
        pool_pool_pe_b_peij_3_1_q_k), .B(pool_pool_pe_b_peij_3_1_add_fai_0_n5), 
        .Z(pool_pool_pe_b_peij_3_1_d_acc[0]) );
  AOI22_X2 pool_pool_pe_b_peij_3_1_add_fai_0_U1 ( .A1(
        pool_pool_pe_b_peij_3_1_add_notb[0]), .A2(pool_pool_pe_b_o_data[22]), 
        .B1(pool_pool_pe_b_peij_3_1_add_fai_0_n5), .B2(
        pool_pool_pe_b_peij_3_1_q_k), .ZN(pool_pool_pe_b_peij_3_1_add_fai_0_n4) );
  INV_X2 pool_pool_pe_b_peij_3_1_add_fai_1_U2 ( .A(
        pool_pool_pe_b_peij_3_1_add_fai_1_n4), .ZN(
        pool_pool_pe_b_peij_3_1_add_cprop[2]) );
  XOR2_X1 pool_pool_pe_b_peij_3_1_add_fai_1_U4 ( .A(pool_pool_pe_b_o_data[23]), 
        .B(pool_pool_pe_b_peij_3_1_add_notb[1]), .Z(
        pool_pool_pe_b_peij_3_1_add_fai_1_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_1_add_fai_1_U3 ( .A(
        pool_pool_pe_b_peij_3_1_add_cprop[1]), .B(
        pool_pool_pe_b_peij_3_1_add_fai_1_n5), .Z(
        pool_pool_pe_b_peij_3_1_d_acc[1]) );
  AOI22_X2 pool_pool_pe_b_peij_3_1_add_fai_1_U1 ( .A1(
        pool_pool_pe_b_peij_3_1_add_notb[1]), .A2(pool_pool_pe_b_o_data[23]), 
        .B1(pool_pool_pe_b_peij_3_1_add_fai_1_n5), .B2(
        pool_pool_pe_b_peij_3_1_add_cprop[1]), .ZN(
        pool_pool_pe_b_peij_3_1_add_fai_1_n4) );
  INV_X2 pool_pool_pe_b_peij_3_1_add_fai_2_U2 ( .A(
        pool_pool_pe_b_peij_3_1_add_fai_2_n4), .ZN(
        pool_pool_pe_b_peij_3_1_add_cprop[3]) );
  XOR2_X1 pool_pool_pe_b_peij_3_1_add_fai_2_U4 ( .A(pool_pool_pe_b_o_data[24]), 
        .B(pool_pool_pe_b_peij_3_1_add_notb[2]), .Z(
        pool_pool_pe_b_peij_3_1_add_fai_2_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_1_add_fai_2_U3 ( .A(
        pool_pool_pe_b_peij_3_1_add_cprop[2]), .B(
        pool_pool_pe_b_peij_3_1_add_fai_2_n5), .Z(
        pool_pool_pe_b_peij_3_1_d_acc[2]) );
  AOI22_X2 pool_pool_pe_b_peij_3_1_add_fai_2_U1 ( .A1(
        pool_pool_pe_b_peij_3_1_add_notb[2]), .A2(pool_pool_pe_b_o_data[24]), 
        .B1(pool_pool_pe_b_peij_3_1_add_fai_2_n5), .B2(
        pool_pool_pe_b_peij_3_1_add_cprop[2]), .ZN(
        pool_pool_pe_b_peij_3_1_add_fai_2_n4) );
  INV_X2 pool_pool_pe_b_peij_3_1_add_fai_3_U2 ( .A(
        pool_pool_pe_b_peij_3_1_add_fai_3_n4), .ZN(
        pool_pool_pe_b_peij_3_1_add_cprop[4]) );
  XOR2_X1 pool_pool_pe_b_peij_3_1_add_fai_3_U4 ( .A(pool_pool_pe_b_o_data[25]), 
        .B(pool_pool_pe_b_peij_3_1_add_notb[3]), .Z(
        pool_pool_pe_b_peij_3_1_add_fai_3_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_1_add_fai_3_U3 ( .A(
        pool_pool_pe_b_peij_3_1_add_cprop[3]), .B(
        pool_pool_pe_b_peij_3_1_add_fai_3_n5), .Z(
        pool_pool_pe_b_peij_3_1_d_acc[3]) );
  AOI22_X2 pool_pool_pe_b_peij_3_1_add_fai_3_U1 ( .A1(
        pool_pool_pe_b_peij_3_1_add_notb[3]), .A2(pool_pool_pe_b_o_data[25]), 
        .B1(pool_pool_pe_b_peij_3_1_add_fai_3_n5), .B2(
        pool_pool_pe_b_peij_3_1_add_cprop[3]), .ZN(
        pool_pool_pe_b_peij_3_1_add_fai_3_n4) );
  INV_X2 pool_pool_pe_b_peij_3_1_add_fai_4_U2 ( .A(
        pool_pool_pe_b_peij_3_1_add_fai_4_n4), .ZN(
        pool_pool_pe_b_peij_3_1_add_cprop[5]) );
  XOR2_X1 pool_pool_pe_b_peij_3_1_add_fai_4_U4 ( .A(pool_pool_pe_b_o_data[26]), 
        .B(pool_pool_pe_b_peij_3_1_add_notb[4]), .Z(
        pool_pool_pe_b_peij_3_1_add_fai_4_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_1_add_fai_4_U3 ( .A(
        pool_pool_pe_b_peij_3_1_add_cprop[4]), .B(
        pool_pool_pe_b_peij_3_1_add_fai_4_n5), .Z(
        pool_pool_pe_b_peij_3_1_d_acc[4]) );
  AOI22_X2 pool_pool_pe_b_peij_3_1_add_fai_4_U1 ( .A1(
        pool_pool_pe_b_peij_3_1_add_notb[4]), .A2(pool_pool_pe_b_o_data[26]), 
        .B1(pool_pool_pe_b_peij_3_1_add_fai_4_n5), .B2(
        pool_pool_pe_b_peij_3_1_add_cprop[4]), .ZN(
        pool_pool_pe_b_peij_3_1_add_fai_4_n4) );
  INV_X2 pool_pool_pe_b_peij_3_1_add_fai_5_U2 ( .A(
        pool_pool_pe_b_peij_3_1_add_fai_5_n4), .ZN(
        pool_pool_pe_b_peij_3_1_add_cprop[6]) );
  XOR2_X1 pool_pool_pe_b_peij_3_1_add_fai_5_U4 ( .A(pool_pool_pe_b_o_data[27]), 
        .B(pool_pool_pe_b_peij_3_1_add_notb[5]), .Z(
        pool_pool_pe_b_peij_3_1_add_fai_5_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_1_add_fai_5_U3 ( .A(
        pool_pool_pe_b_peij_3_1_add_cprop[5]), .B(
        pool_pool_pe_b_peij_3_1_add_fai_5_n5), .Z(
        pool_pool_pe_b_peij_3_1_d_acc[5]) );
  AOI22_X2 pool_pool_pe_b_peij_3_1_add_fai_5_U1 ( .A1(
        pool_pool_pe_b_peij_3_1_add_notb[5]), .A2(pool_pool_pe_b_o_data[27]), 
        .B1(pool_pool_pe_b_peij_3_1_add_fai_5_n5), .B2(
        pool_pool_pe_b_peij_3_1_add_cprop[5]), .ZN(
        pool_pool_pe_b_peij_3_1_add_fai_5_n4) );
  INV_X2 pool_pool_pe_b_peij_3_1_add_fai_6_U2 ( .A(
        pool_pool_pe_b_peij_3_1_add_fai_6_n4), .ZN(
        pool_pool_pe_b_peij_3_1_add_cprop[7]) );
  XOR2_X1 pool_pool_pe_b_peij_3_1_add_fai_6_U4 ( .A(pool_pool_pe_b_o_data[28]), 
        .B(pool_pool_pe_b_peij_3_1_add_notb[6]), .Z(
        pool_pool_pe_b_peij_3_1_add_fai_6_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_1_add_fai_6_U3 ( .A(
        pool_pool_pe_b_peij_3_1_add_cprop[6]), .B(
        pool_pool_pe_b_peij_3_1_add_fai_6_n5), .Z(
        pool_pool_pe_b_peij_3_1_d_acc[6]) );
  AOI22_X2 pool_pool_pe_b_peij_3_1_add_fai_6_U1 ( .A1(
        pool_pool_pe_b_peij_3_1_add_notb[6]), .A2(pool_pool_pe_b_o_data[28]), 
        .B1(pool_pool_pe_b_peij_3_1_add_fai_6_n5), .B2(
        pool_pool_pe_b_peij_3_1_add_cprop[6]), .ZN(
        pool_pool_pe_b_peij_3_1_add_fai_6_n4) );
  INV_X2 pool_pool_pe_b_peij_3_1_add_fai_7_U2 ( .A(
        pool_pool_pe_b_peij_3_1_add_fai_7_n4), .ZN(
        pool_pool_pe_b_peij_3_1_add_cprop[8]) );
  XOR2_X1 pool_pool_pe_b_peij_3_1_add_fai_7_U4 ( .A(pool_pool_pe_b_o_data[29]), 
        .B(pool_pool_pe_b_peij_3_1_add_notb[7]), .Z(
        pool_pool_pe_b_peij_3_1_add_fai_7_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_1_add_fai_7_U3 ( .A(
        pool_pool_pe_b_peij_3_1_add_cprop[7]), .B(
        pool_pool_pe_b_peij_3_1_add_fai_7_n5), .Z(
        pool_pool_pe_b_peij_3_1_d_acc[7]) );
  AOI22_X2 pool_pool_pe_b_peij_3_1_add_fai_7_U1 ( .A1(
        pool_pool_pe_b_peij_3_1_add_notb[7]), .A2(pool_pool_pe_b_o_data[29]), 
        .B1(pool_pool_pe_b_peij_3_1_add_fai_7_n5), .B2(
        pool_pool_pe_b_peij_3_1_add_cprop[7]), .ZN(
        pool_pool_pe_b_peij_3_1_add_fai_7_n4) );
  INV_X2 pool_pool_pe_b_peij_3_1_add_fai_8_U2 ( .A(
        pool_pool_pe_b_peij_3_1_add_fai_8_n4), .ZN(
        pool_pool_pe_b_peij_3_1_add_cprop[9]) );
  XOR2_X1 pool_pool_pe_b_peij_3_1_add_fai_8_U4 ( .A(pool_pool_pe_b_o_data[30]), 
        .B(pool_pool_pe_b_peij_3_1_add_notb[8]), .Z(
        pool_pool_pe_b_peij_3_1_add_fai_8_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_1_add_fai_8_U3 ( .A(
        pool_pool_pe_b_peij_3_1_add_cprop[8]), .B(
        pool_pool_pe_b_peij_3_1_add_fai_8_n5), .Z(
        pool_pool_pe_b_peij_3_1_d_acc[8]) );
  AOI22_X2 pool_pool_pe_b_peij_3_1_add_fai_8_U1 ( .A1(
        pool_pool_pe_b_peij_3_1_add_notb[8]), .A2(pool_pool_pe_b_o_data[30]), 
        .B1(pool_pool_pe_b_peij_3_1_add_fai_8_n5), .B2(
        pool_pool_pe_b_peij_3_1_add_cprop[8]), .ZN(
        pool_pool_pe_b_peij_3_1_add_fai_8_n4) );
  INV_X2 pool_pool_pe_b_peij_3_1_add_fai_9_U2 ( .A(
        pool_pool_pe_b_peij_3_1_add_fai_9_n4), .ZN(
        pool_pool_pe_b_peij_3_1_add_cprop[10]) );
  XOR2_X1 pool_pool_pe_b_peij_3_1_add_fai_9_U4 ( .A(pool_pool_pe_b_o_data[31]), 
        .B(pool_pool_pe_b_peij_3_1_add_notb[9]), .Z(
        pool_pool_pe_b_peij_3_1_add_fai_9_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_1_add_fai_9_U3 ( .A(
        pool_pool_pe_b_peij_3_1_add_cprop[9]), .B(
        pool_pool_pe_b_peij_3_1_add_fai_9_n5), .Z(
        pool_pool_pe_b_peij_3_1_d_acc[9]) );
  AOI22_X2 pool_pool_pe_b_peij_3_1_add_fai_9_U1 ( .A1(
        pool_pool_pe_b_peij_3_1_add_notb[9]), .A2(pool_pool_pe_b_o_data[31]), 
        .B1(pool_pool_pe_b_peij_3_1_add_fai_9_n5), .B2(
        pool_pool_pe_b_peij_3_1_add_cprop[9]), .ZN(
        pool_pool_pe_b_peij_3_1_add_fai_9_n4) );
  INV_X2 pool_pool_pe_b_peij_3_1_add_fai_10_U2 ( .A(
        pool_pool_pe_b_peij_3_1_add_fai_10_n4), .ZN(
        pool_pool_pe_b_peij_3_1_add_c_out) );
  XOR2_X1 pool_pool_pe_b_peij_3_1_add_fai_10_U4 ( .A(pool_pool_pe_b_o_data[32]), .B(pool_pool_pe_b_peij_3_1_add_notb[10]), .Z(
        pool_pool_pe_b_peij_3_1_add_fai_10_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_1_add_fai_10_U3 ( .A(
        pool_pool_pe_b_peij_3_1_add_cprop[10]), .B(
        pool_pool_pe_b_peij_3_1_add_fai_10_n5), .Z(
        pool_pool_pe_b_peij_3_1_d_acc[10]) );
  AOI22_X2 pool_pool_pe_b_peij_3_1_add_fai_10_U1 ( .A1(
        pool_pool_pe_b_peij_3_1_add_notb[10]), .A2(pool_pool_pe_b_o_data[32]), 
        .B1(pool_pool_pe_b_peij_3_1_add_fai_10_n5), .B2(
        pool_pool_pe_b_peij_3_1_add_cprop[10]), .ZN(
        pool_pool_pe_b_peij_3_1_add_fai_10_n4) );
  INV_X2 pool_pool_pe_b_peij_3_2_U21 ( .A(pool_sync_clr), .ZN(
        pool_pool_pe_b_peij_3_2_n14) );
  INV_X1 pool_pool_pe_b_peij_3_2_U18 ( .A(pool_pool_pe_b_n1), .ZN(
        pool_pool_pe_b_peij_3_2_n12) );
  AND2_X1 pool_pool_pe_b_peij_3_2_U13 ( .A1(pool_pool_pe_b_peij_3_2_d_acc[0]), 
        .A2(pool_pool_pe_b_peij_3_2_n14), .ZN(pool_pool_pe_b_peij_3_2_n11) );
  AND2_X1 pool_pool_pe_b_peij_3_2_U12 ( .A1(pool_pool_pe_b_peij_3_2_d_acc[1]), 
        .A2(pool_pool_pe_b_peij_3_2_n14), .ZN(pool_pool_pe_b_peij_3_2_n10) );
  AND2_X1 pool_pool_pe_b_peij_3_2_U11 ( .A1(pool_pool_pe_b_peij_3_2_d_acc[2]), 
        .A2(pool_pool_pe_b_peij_3_2_n14), .ZN(pool_pool_pe_b_peij_3_2_n9) );
  AND2_X1 pool_pool_pe_b_peij_3_2_U10 ( .A1(pool_pool_pe_b_peij_3_2_d_acc[3]), 
        .A2(pool_pool_pe_b_peij_3_2_n14), .ZN(pool_pool_pe_b_peij_3_2_n8) );
  AND2_X1 pool_pool_pe_b_peij_3_2_U9 ( .A1(pool_pool_pe_b_peij_3_2_d_acc[4]), 
        .A2(pool_pool_pe_b_peij_3_2_n14), .ZN(pool_pool_pe_b_peij_3_2_n7) );
  AND2_X1 pool_pool_pe_b_peij_3_2_U8 ( .A1(pool_pool_pe_b_peij_3_2_d_acc[5]), 
        .A2(pool_pool_pe_b_peij_3_2_n14), .ZN(pool_pool_pe_b_peij_3_2_n6) );
  AND2_X1 pool_pool_pe_b_peij_3_2_U7 ( .A1(pool_pool_pe_b_peij_3_2_d_acc[6]), 
        .A2(pool_pool_pe_b_peij_3_2_n14), .ZN(pool_pool_pe_b_peij_3_2_n5) );
  AND2_X1 pool_pool_pe_b_peij_3_2_U6 ( .A1(pool_pool_pe_b_peij_3_2_d_acc[7]), 
        .A2(pool_pool_pe_b_peij_3_2_n14), .ZN(pool_pool_pe_b_peij_3_2_n4) );
  AND2_X1 pool_pool_pe_b_peij_3_2_U5 ( .A1(pool_pool_pe_b_peij_3_2_d_acc[8]), 
        .A2(pool_pool_pe_b_peij_3_2_n14), .ZN(pool_pool_pe_b_peij_3_2_n3) );
  AND2_X1 pool_pool_pe_b_peij_3_2_U4 ( .A1(pool_pool_pe_b_peij_3_2_d_acc[9]), 
        .A2(pool_pool_pe_b_peij_3_2_n14), .ZN(pool_pool_pe_b_peij_3_2_n2) );
  AND2_X1 pool_pool_pe_b_peij_3_2_U3 ( .A1(pool_pool_pe_b_peij_3_2_d_acc[10]), 
        .A2(pool_pool_pe_b_peij_3_2_n14), .ZN(pool_pool_pe_b_peij_3_2_n1) );
  DFFR_X1 pool_pool_pe_b_peij_3_2_q_acc_reg_10_ ( .D(
        pool_pool_pe_b_peij_3_2_n1), .CK(pool_pool_pe_b_peij_3_2_gck), .RN(
        pool_pool_pe_b_peij_3_2_n12), .Q(pool_pool_pe_b_o_data[21]) );
  DFFR_X1 pool_pool_pe_b_peij_3_2_q_acc_reg_9_ ( .D(pool_pool_pe_b_peij_3_2_n2), .CK(pool_pool_pe_b_peij_3_2_gck), .RN(pool_pool_pe_b_peij_3_2_n12), .Q(
        pool_pool_pe_b_o_data[20]) );
  DFFR_X1 pool_pool_pe_b_peij_3_2_q_acc_reg_8_ ( .D(pool_pool_pe_b_peij_3_2_n3), .CK(pool_pool_pe_b_peij_3_2_gck), .RN(pool_pool_pe_b_peij_3_2_n12), .Q(
        pool_pool_pe_b_o_data[19]) );
  DFFR_X1 pool_pool_pe_b_peij_3_2_q_acc_reg_7_ ( .D(pool_pool_pe_b_peij_3_2_n4), .CK(pool_pool_pe_b_peij_3_2_gck), .RN(pool_pool_pe_b_peij_3_2_n12), .Q(
        pool_pool_pe_b_o_data[18]) );
  DFFR_X1 pool_pool_pe_b_peij_3_2_q_acc_reg_6_ ( .D(pool_pool_pe_b_peij_3_2_n5), .CK(pool_pool_pe_b_peij_3_2_gck), .RN(pool_pool_pe_b_peij_3_2_n12), .Q(
        pool_pool_pe_b_o_data[17]) );
  DFFR_X1 pool_pool_pe_b_peij_3_2_q_acc_reg_5_ ( .D(pool_pool_pe_b_peij_3_2_n6), .CK(pool_pool_pe_b_peij_3_2_gck), .RN(pool_pool_pe_b_peij_3_2_n12), .Q(
        pool_pool_pe_b_o_data[16]) );
  DFFR_X1 pool_pool_pe_b_peij_3_2_q_acc_reg_4_ ( .D(pool_pool_pe_b_peij_3_2_n7), .CK(pool_pool_pe_b_peij_3_2_gck), .RN(pool_pool_pe_b_peij_3_2_n12), .Q(
        pool_pool_pe_b_o_data[15]) );
  DFFR_X1 pool_pool_pe_b_peij_3_2_q_acc_reg_3_ ( .D(pool_pool_pe_b_peij_3_2_n8), .CK(pool_pool_pe_b_peij_3_2_gck), .RN(pool_pool_pe_b_peij_3_2_n12), .Q(
        pool_pool_pe_b_o_data[14]) );
  DFFR_X1 pool_pool_pe_b_peij_3_2_q_acc_reg_2_ ( .D(pool_pool_pe_b_peij_3_2_n9), .CK(pool_pool_pe_b_peij_3_2_gck), .RN(pool_pool_pe_b_peij_3_2_n12), .Q(
        pool_pool_pe_b_o_data[13]) );
  DFFR_X1 pool_pool_pe_b_peij_3_2_q_acc_reg_1_ ( .D(
        pool_pool_pe_b_peij_3_2_n10), .CK(pool_pool_pe_b_peij_3_2_gck), .RN(
        pool_pool_pe_b_peij_3_2_n12), .Q(pool_pool_pe_b_o_data[12]) );
  DFFR_X1 pool_pool_pe_b_peij_3_2_q_acc_reg_0_ ( .D(
        pool_pool_pe_b_peij_3_2_n11), .CK(pool_pool_pe_b_peij_3_2_gck), .RN(
        pool_pool_pe_b_peij_3_2_n12), .Q(pool_pool_pe_b_o_data[11]) );
  AND3_X2 pool_pool_pe_b_peij_3_2_U20 ( .A1(pool_pool_pe_b_int_pe_en[1]), .A2(
        clk), .A3(1'b1), .ZN(pool_pool_pe_b_peij_3_2_gck) );
  SDFFR_X1 pool_pool_pe_b_peij_3_2_q_k_reg ( .D(1'b0), .SI(
        pool_pool_pe_b_peij_3_2_n14), .SE(1'b0), .CK(
        pool_pool_pe_b_peij_3_2_gck), .RN(pool_pool_pe_b_peij_3_2_n12), .Q(
        pool_pool_pe_b_peij_3_2_q_k) );
  XOR2_X1 pool_pool_pe_b_peij_3_2_add_U11 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_2_q_k), .Z(pool_pool_pe_b_peij_3_2_add_notb[0])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_2_add_U10 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_2_q_k), .Z(pool_pool_pe_b_peij_3_2_add_notb[10])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_2_add_U9 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_2_q_k), .Z(pool_pool_pe_b_peij_3_2_add_notb[1])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_2_add_U8 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_2_q_k), .Z(pool_pool_pe_b_peij_3_2_add_notb[2])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_2_add_U7 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_2_q_k), .Z(pool_pool_pe_b_peij_3_2_add_notb[3])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_2_add_U6 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_2_q_k), .Z(pool_pool_pe_b_peij_3_2_add_notb[4])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_2_add_U5 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_2_q_k), .Z(pool_pool_pe_b_peij_3_2_add_notb[5])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_2_add_U4 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_2_q_k), .Z(pool_pool_pe_b_peij_3_2_add_notb[6])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_2_add_U3 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_2_q_k), .Z(pool_pool_pe_b_peij_3_2_add_notb[7])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_2_add_U2 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_2_q_k), .Z(pool_pool_pe_b_peij_3_2_add_notb[8])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_2_add_U1 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_2_q_k), .Z(pool_pool_pe_b_peij_3_2_add_notb[9])
         );
  INV_X2 pool_pool_pe_b_peij_3_2_add_fai_0_U2 ( .A(
        pool_pool_pe_b_peij_3_2_add_fai_0_n4), .ZN(
        pool_pool_pe_b_peij_3_2_add_cprop[1]) );
  XOR2_X1 pool_pool_pe_b_peij_3_2_add_fai_0_U4 ( .A(pool_pool_pe_b_o_data[11]), 
        .B(pool_pool_pe_b_peij_3_2_add_notb[0]), .Z(
        pool_pool_pe_b_peij_3_2_add_fai_0_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_2_add_fai_0_U3 ( .A(
        pool_pool_pe_b_peij_3_2_q_k), .B(pool_pool_pe_b_peij_3_2_add_fai_0_n5), 
        .Z(pool_pool_pe_b_peij_3_2_d_acc[0]) );
  AOI22_X2 pool_pool_pe_b_peij_3_2_add_fai_0_U1 ( .A1(
        pool_pool_pe_b_peij_3_2_add_notb[0]), .A2(pool_pool_pe_b_o_data[11]), 
        .B1(pool_pool_pe_b_peij_3_2_add_fai_0_n5), .B2(
        pool_pool_pe_b_peij_3_2_q_k), .ZN(pool_pool_pe_b_peij_3_2_add_fai_0_n4) );
  INV_X2 pool_pool_pe_b_peij_3_2_add_fai_1_U2 ( .A(
        pool_pool_pe_b_peij_3_2_add_fai_1_n4), .ZN(
        pool_pool_pe_b_peij_3_2_add_cprop[2]) );
  XOR2_X1 pool_pool_pe_b_peij_3_2_add_fai_1_U4 ( .A(pool_pool_pe_b_o_data[12]), 
        .B(pool_pool_pe_b_peij_3_2_add_notb[1]), .Z(
        pool_pool_pe_b_peij_3_2_add_fai_1_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_2_add_fai_1_U3 ( .A(
        pool_pool_pe_b_peij_3_2_add_cprop[1]), .B(
        pool_pool_pe_b_peij_3_2_add_fai_1_n5), .Z(
        pool_pool_pe_b_peij_3_2_d_acc[1]) );
  AOI22_X2 pool_pool_pe_b_peij_3_2_add_fai_1_U1 ( .A1(
        pool_pool_pe_b_peij_3_2_add_notb[1]), .A2(pool_pool_pe_b_o_data[12]), 
        .B1(pool_pool_pe_b_peij_3_2_add_fai_1_n5), .B2(
        pool_pool_pe_b_peij_3_2_add_cprop[1]), .ZN(
        pool_pool_pe_b_peij_3_2_add_fai_1_n4) );
  INV_X2 pool_pool_pe_b_peij_3_2_add_fai_2_U2 ( .A(
        pool_pool_pe_b_peij_3_2_add_fai_2_n4), .ZN(
        pool_pool_pe_b_peij_3_2_add_cprop[3]) );
  XOR2_X1 pool_pool_pe_b_peij_3_2_add_fai_2_U4 ( .A(pool_pool_pe_b_o_data[13]), 
        .B(pool_pool_pe_b_peij_3_2_add_notb[2]), .Z(
        pool_pool_pe_b_peij_3_2_add_fai_2_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_2_add_fai_2_U3 ( .A(
        pool_pool_pe_b_peij_3_2_add_cprop[2]), .B(
        pool_pool_pe_b_peij_3_2_add_fai_2_n5), .Z(
        pool_pool_pe_b_peij_3_2_d_acc[2]) );
  AOI22_X2 pool_pool_pe_b_peij_3_2_add_fai_2_U1 ( .A1(
        pool_pool_pe_b_peij_3_2_add_notb[2]), .A2(pool_pool_pe_b_o_data[13]), 
        .B1(pool_pool_pe_b_peij_3_2_add_fai_2_n5), .B2(
        pool_pool_pe_b_peij_3_2_add_cprop[2]), .ZN(
        pool_pool_pe_b_peij_3_2_add_fai_2_n4) );
  INV_X2 pool_pool_pe_b_peij_3_2_add_fai_3_U2 ( .A(
        pool_pool_pe_b_peij_3_2_add_fai_3_n4), .ZN(
        pool_pool_pe_b_peij_3_2_add_cprop[4]) );
  XOR2_X1 pool_pool_pe_b_peij_3_2_add_fai_3_U4 ( .A(pool_pool_pe_b_o_data[14]), 
        .B(pool_pool_pe_b_peij_3_2_add_notb[3]), .Z(
        pool_pool_pe_b_peij_3_2_add_fai_3_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_2_add_fai_3_U3 ( .A(
        pool_pool_pe_b_peij_3_2_add_cprop[3]), .B(
        pool_pool_pe_b_peij_3_2_add_fai_3_n5), .Z(
        pool_pool_pe_b_peij_3_2_d_acc[3]) );
  AOI22_X2 pool_pool_pe_b_peij_3_2_add_fai_3_U1 ( .A1(
        pool_pool_pe_b_peij_3_2_add_notb[3]), .A2(pool_pool_pe_b_o_data[14]), 
        .B1(pool_pool_pe_b_peij_3_2_add_fai_3_n5), .B2(
        pool_pool_pe_b_peij_3_2_add_cprop[3]), .ZN(
        pool_pool_pe_b_peij_3_2_add_fai_3_n4) );
  INV_X2 pool_pool_pe_b_peij_3_2_add_fai_4_U2 ( .A(
        pool_pool_pe_b_peij_3_2_add_fai_4_n4), .ZN(
        pool_pool_pe_b_peij_3_2_add_cprop[5]) );
  XOR2_X1 pool_pool_pe_b_peij_3_2_add_fai_4_U4 ( .A(pool_pool_pe_b_o_data[15]), 
        .B(pool_pool_pe_b_peij_3_2_add_notb[4]), .Z(
        pool_pool_pe_b_peij_3_2_add_fai_4_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_2_add_fai_4_U3 ( .A(
        pool_pool_pe_b_peij_3_2_add_cprop[4]), .B(
        pool_pool_pe_b_peij_3_2_add_fai_4_n5), .Z(
        pool_pool_pe_b_peij_3_2_d_acc[4]) );
  AOI22_X2 pool_pool_pe_b_peij_3_2_add_fai_4_U1 ( .A1(
        pool_pool_pe_b_peij_3_2_add_notb[4]), .A2(pool_pool_pe_b_o_data[15]), 
        .B1(pool_pool_pe_b_peij_3_2_add_fai_4_n5), .B2(
        pool_pool_pe_b_peij_3_2_add_cprop[4]), .ZN(
        pool_pool_pe_b_peij_3_2_add_fai_4_n4) );
  INV_X2 pool_pool_pe_b_peij_3_2_add_fai_5_U2 ( .A(
        pool_pool_pe_b_peij_3_2_add_fai_5_n4), .ZN(
        pool_pool_pe_b_peij_3_2_add_cprop[6]) );
  XOR2_X1 pool_pool_pe_b_peij_3_2_add_fai_5_U4 ( .A(pool_pool_pe_b_o_data[16]), 
        .B(pool_pool_pe_b_peij_3_2_add_notb[5]), .Z(
        pool_pool_pe_b_peij_3_2_add_fai_5_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_2_add_fai_5_U3 ( .A(
        pool_pool_pe_b_peij_3_2_add_cprop[5]), .B(
        pool_pool_pe_b_peij_3_2_add_fai_5_n5), .Z(
        pool_pool_pe_b_peij_3_2_d_acc[5]) );
  AOI22_X2 pool_pool_pe_b_peij_3_2_add_fai_5_U1 ( .A1(
        pool_pool_pe_b_peij_3_2_add_notb[5]), .A2(pool_pool_pe_b_o_data[16]), 
        .B1(pool_pool_pe_b_peij_3_2_add_fai_5_n5), .B2(
        pool_pool_pe_b_peij_3_2_add_cprop[5]), .ZN(
        pool_pool_pe_b_peij_3_2_add_fai_5_n4) );
  INV_X2 pool_pool_pe_b_peij_3_2_add_fai_6_U2 ( .A(
        pool_pool_pe_b_peij_3_2_add_fai_6_n4), .ZN(
        pool_pool_pe_b_peij_3_2_add_cprop[7]) );
  XOR2_X1 pool_pool_pe_b_peij_3_2_add_fai_6_U4 ( .A(pool_pool_pe_b_o_data[17]), 
        .B(pool_pool_pe_b_peij_3_2_add_notb[6]), .Z(
        pool_pool_pe_b_peij_3_2_add_fai_6_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_2_add_fai_6_U3 ( .A(
        pool_pool_pe_b_peij_3_2_add_cprop[6]), .B(
        pool_pool_pe_b_peij_3_2_add_fai_6_n5), .Z(
        pool_pool_pe_b_peij_3_2_d_acc[6]) );
  AOI22_X2 pool_pool_pe_b_peij_3_2_add_fai_6_U1 ( .A1(
        pool_pool_pe_b_peij_3_2_add_notb[6]), .A2(pool_pool_pe_b_o_data[17]), 
        .B1(pool_pool_pe_b_peij_3_2_add_fai_6_n5), .B2(
        pool_pool_pe_b_peij_3_2_add_cprop[6]), .ZN(
        pool_pool_pe_b_peij_3_2_add_fai_6_n4) );
  INV_X2 pool_pool_pe_b_peij_3_2_add_fai_7_U2 ( .A(
        pool_pool_pe_b_peij_3_2_add_fai_7_n4), .ZN(
        pool_pool_pe_b_peij_3_2_add_cprop[8]) );
  XOR2_X1 pool_pool_pe_b_peij_3_2_add_fai_7_U4 ( .A(pool_pool_pe_b_o_data[18]), 
        .B(pool_pool_pe_b_peij_3_2_add_notb[7]), .Z(
        pool_pool_pe_b_peij_3_2_add_fai_7_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_2_add_fai_7_U3 ( .A(
        pool_pool_pe_b_peij_3_2_add_cprop[7]), .B(
        pool_pool_pe_b_peij_3_2_add_fai_7_n5), .Z(
        pool_pool_pe_b_peij_3_2_d_acc[7]) );
  AOI22_X2 pool_pool_pe_b_peij_3_2_add_fai_7_U1 ( .A1(
        pool_pool_pe_b_peij_3_2_add_notb[7]), .A2(pool_pool_pe_b_o_data[18]), 
        .B1(pool_pool_pe_b_peij_3_2_add_fai_7_n5), .B2(
        pool_pool_pe_b_peij_3_2_add_cprop[7]), .ZN(
        pool_pool_pe_b_peij_3_2_add_fai_7_n4) );
  INV_X2 pool_pool_pe_b_peij_3_2_add_fai_8_U2 ( .A(
        pool_pool_pe_b_peij_3_2_add_fai_8_n4), .ZN(
        pool_pool_pe_b_peij_3_2_add_cprop[9]) );
  XOR2_X1 pool_pool_pe_b_peij_3_2_add_fai_8_U4 ( .A(pool_pool_pe_b_o_data[19]), 
        .B(pool_pool_pe_b_peij_3_2_add_notb[8]), .Z(
        pool_pool_pe_b_peij_3_2_add_fai_8_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_2_add_fai_8_U3 ( .A(
        pool_pool_pe_b_peij_3_2_add_cprop[8]), .B(
        pool_pool_pe_b_peij_3_2_add_fai_8_n5), .Z(
        pool_pool_pe_b_peij_3_2_d_acc[8]) );
  AOI22_X2 pool_pool_pe_b_peij_3_2_add_fai_8_U1 ( .A1(
        pool_pool_pe_b_peij_3_2_add_notb[8]), .A2(pool_pool_pe_b_o_data[19]), 
        .B1(pool_pool_pe_b_peij_3_2_add_fai_8_n5), .B2(
        pool_pool_pe_b_peij_3_2_add_cprop[8]), .ZN(
        pool_pool_pe_b_peij_3_2_add_fai_8_n4) );
  INV_X2 pool_pool_pe_b_peij_3_2_add_fai_9_U2 ( .A(
        pool_pool_pe_b_peij_3_2_add_fai_9_n4), .ZN(
        pool_pool_pe_b_peij_3_2_add_cprop[10]) );
  XOR2_X1 pool_pool_pe_b_peij_3_2_add_fai_9_U4 ( .A(pool_pool_pe_b_o_data[20]), 
        .B(pool_pool_pe_b_peij_3_2_add_notb[9]), .Z(
        pool_pool_pe_b_peij_3_2_add_fai_9_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_2_add_fai_9_U3 ( .A(
        pool_pool_pe_b_peij_3_2_add_cprop[9]), .B(
        pool_pool_pe_b_peij_3_2_add_fai_9_n5), .Z(
        pool_pool_pe_b_peij_3_2_d_acc[9]) );
  AOI22_X2 pool_pool_pe_b_peij_3_2_add_fai_9_U1 ( .A1(
        pool_pool_pe_b_peij_3_2_add_notb[9]), .A2(pool_pool_pe_b_o_data[20]), 
        .B1(pool_pool_pe_b_peij_3_2_add_fai_9_n5), .B2(
        pool_pool_pe_b_peij_3_2_add_cprop[9]), .ZN(
        pool_pool_pe_b_peij_3_2_add_fai_9_n4) );
  INV_X2 pool_pool_pe_b_peij_3_2_add_fai_10_U2 ( .A(
        pool_pool_pe_b_peij_3_2_add_fai_10_n4), .ZN(
        pool_pool_pe_b_peij_3_2_add_c_out) );
  XOR2_X1 pool_pool_pe_b_peij_3_2_add_fai_10_U4 ( .A(pool_pool_pe_b_o_data[21]), .B(pool_pool_pe_b_peij_3_2_add_notb[10]), .Z(
        pool_pool_pe_b_peij_3_2_add_fai_10_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_2_add_fai_10_U3 ( .A(
        pool_pool_pe_b_peij_3_2_add_cprop[10]), .B(
        pool_pool_pe_b_peij_3_2_add_fai_10_n5), .Z(
        pool_pool_pe_b_peij_3_2_d_acc[10]) );
  AOI22_X2 pool_pool_pe_b_peij_3_2_add_fai_10_U1 ( .A1(
        pool_pool_pe_b_peij_3_2_add_notb[10]), .A2(pool_pool_pe_b_o_data[21]), 
        .B1(pool_pool_pe_b_peij_3_2_add_fai_10_n5), .B2(
        pool_pool_pe_b_peij_3_2_add_cprop[10]), .ZN(
        pool_pool_pe_b_peij_3_2_add_fai_10_n4) );
  INV_X2 pool_pool_pe_b_peij_3_3_U21 ( .A(pool_sync_clr), .ZN(
        pool_pool_pe_b_peij_3_3_n14) );
  INV_X1 pool_pool_pe_b_peij_3_3_U18 ( .A(pool_pool_pe_b_n1), .ZN(
        pool_pool_pe_b_peij_3_3_n12) );
  AND2_X1 pool_pool_pe_b_peij_3_3_U13 ( .A1(pool_pool_pe_b_peij_3_3_d_acc[0]), 
        .A2(pool_pool_pe_b_peij_3_3_n14), .ZN(pool_pool_pe_b_peij_3_3_n11) );
  AND2_X1 pool_pool_pe_b_peij_3_3_U12 ( .A1(pool_pool_pe_b_peij_3_3_d_acc[1]), 
        .A2(pool_pool_pe_b_peij_3_3_n14), .ZN(pool_pool_pe_b_peij_3_3_n10) );
  AND2_X1 pool_pool_pe_b_peij_3_3_U11 ( .A1(pool_pool_pe_b_peij_3_3_d_acc[2]), 
        .A2(pool_pool_pe_b_peij_3_3_n14), .ZN(pool_pool_pe_b_peij_3_3_n9) );
  AND2_X1 pool_pool_pe_b_peij_3_3_U10 ( .A1(pool_pool_pe_b_peij_3_3_d_acc[3]), 
        .A2(pool_pool_pe_b_peij_3_3_n14), .ZN(pool_pool_pe_b_peij_3_3_n8) );
  AND2_X1 pool_pool_pe_b_peij_3_3_U9 ( .A1(pool_pool_pe_b_peij_3_3_d_acc[4]), 
        .A2(pool_pool_pe_b_peij_3_3_n14), .ZN(pool_pool_pe_b_peij_3_3_n7) );
  AND2_X1 pool_pool_pe_b_peij_3_3_U8 ( .A1(pool_pool_pe_b_peij_3_3_d_acc[5]), 
        .A2(pool_pool_pe_b_peij_3_3_n14), .ZN(pool_pool_pe_b_peij_3_3_n6) );
  AND2_X1 pool_pool_pe_b_peij_3_3_U7 ( .A1(pool_pool_pe_b_peij_3_3_d_acc[6]), 
        .A2(pool_pool_pe_b_peij_3_3_n14), .ZN(pool_pool_pe_b_peij_3_3_n5) );
  AND2_X1 pool_pool_pe_b_peij_3_3_U6 ( .A1(pool_pool_pe_b_peij_3_3_d_acc[7]), 
        .A2(pool_pool_pe_b_peij_3_3_n14), .ZN(pool_pool_pe_b_peij_3_3_n4) );
  AND2_X1 pool_pool_pe_b_peij_3_3_U5 ( .A1(pool_pool_pe_b_peij_3_3_d_acc[8]), 
        .A2(pool_pool_pe_b_peij_3_3_n14), .ZN(pool_pool_pe_b_peij_3_3_n3) );
  AND2_X1 pool_pool_pe_b_peij_3_3_U4 ( .A1(pool_pool_pe_b_peij_3_3_d_acc[9]), 
        .A2(pool_pool_pe_b_peij_3_3_n14), .ZN(pool_pool_pe_b_peij_3_3_n2) );
  AND2_X1 pool_pool_pe_b_peij_3_3_U3 ( .A1(pool_pool_pe_b_peij_3_3_d_acc[10]), 
        .A2(pool_pool_pe_b_peij_3_3_n14), .ZN(pool_pool_pe_b_peij_3_3_n1) );
  DFFR_X1 pool_pool_pe_b_peij_3_3_q_acc_reg_10_ ( .D(
        pool_pool_pe_b_peij_3_3_n1), .CK(pool_pool_pe_b_peij_3_3_gck), .RN(
        pool_pool_pe_b_peij_3_3_n12), .Q(pool_pool_pe_b_o_data[10]) );
  DFFR_X1 pool_pool_pe_b_peij_3_3_q_acc_reg_9_ ( .D(pool_pool_pe_b_peij_3_3_n2), .CK(pool_pool_pe_b_peij_3_3_gck), .RN(pool_pool_pe_b_peij_3_3_n12), .Q(
        pool_pool_pe_b_o_data[9]) );
  DFFR_X1 pool_pool_pe_b_peij_3_3_q_acc_reg_8_ ( .D(pool_pool_pe_b_peij_3_3_n3), .CK(pool_pool_pe_b_peij_3_3_gck), .RN(pool_pool_pe_b_peij_3_3_n12), .Q(
        pool_pool_pe_b_o_data[8]) );
  DFFR_X1 pool_pool_pe_b_peij_3_3_q_acc_reg_7_ ( .D(pool_pool_pe_b_peij_3_3_n4), .CK(pool_pool_pe_b_peij_3_3_gck), .RN(pool_pool_pe_b_peij_3_3_n12), .Q(
        pool_pool_pe_b_o_data[7]) );
  DFFR_X1 pool_pool_pe_b_peij_3_3_q_acc_reg_6_ ( .D(pool_pool_pe_b_peij_3_3_n5), .CK(pool_pool_pe_b_peij_3_3_gck), .RN(pool_pool_pe_b_peij_3_3_n12), .Q(
        pool_pool_pe_b_o_data[6]) );
  DFFR_X1 pool_pool_pe_b_peij_3_3_q_acc_reg_5_ ( .D(pool_pool_pe_b_peij_3_3_n6), .CK(pool_pool_pe_b_peij_3_3_gck), .RN(pool_pool_pe_b_peij_3_3_n12), .Q(
        pool_pool_pe_b_o_data[5]) );
  DFFR_X1 pool_pool_pe_b_peij_3_3_q_acc_reg_4_ ( .D(pool_pool_pe_b_peij_3_3_n7), .CK(pool_pool_pe_b_peij_3_3_gck), .RN(pool_pool_pe_b_peij_3_3_n12), .Q(
        pool_pool_pe_b_o_data[4]) );
  DFFR_X1 pool_pool_pe_b_peij_3_3_q_acc_reg_3_ ( .D(pool_pool_pe_b_peij_3_3_n8), .CK(pool_pool_pe_b_peij_3_3_gck), .RN(pool_pool_pe_b_peij_3_3_n12), .Q(
        pool_pool_pe_b_o_data[3]) );
  DFFR_X1 pool_pool_pe_b_peij_3_3_q_acc_reg_2_ ( .D(pool_pool_pe_b_peij_3_3_n9), .CK(pool_pool_pe_b_peij_3_3_gck), .RN(pool_pool_pe_b_peij_3_3_n12), .Q(
        pool_pool_pe_b_o_data[2]) );
  DFFR_X1 pool_pool_pe_b_peij_3_3_q_acc_reg_1_ ( .D(
        pool_pool_pe_b_peij_3_3_n10), .CK(pool_pool_pe_b_peij_3_3_gck), .RN(
        pool_pool_pe_b_peij_3_3_n12), .Q(pool_pool_pe_b_o_data[1]) );
  DFFR_X1 pool_pool_pe_b_peij_3_3_q_acc_reg_0_ ( .D(
        pool_pool_pe_b_peij_3_3_n11), .CK(pool_pool_pe_b_peij_3_3_gck), .RN(
        pool_pool_pe_b_peij_3_3_n12), .Q(pool_pool_pe_b_o_data[0]) );
  AND3_X2 pool_pool_pe_b_peij_3_3_U20 ( .A1(pool_pool_pe_b_int_pe_en[0]), .A2(
        clk), .A3(1'b1), .ZN(pool_pool_pe_b_peij_3_3_gck) );
  SDFFR_X1 pool_pool_pe_b_peij_3_3_q_k_reg ( .D(1'b0), .SI(
        pool_pool_pe_b_peij_3_3_n14), .SE(1'b0), .CK(
        pool_pool_pe_b_peij_3_3_gck), .RN(pool_pool_pe_b_peij_3_3_n12), .Q(
        pool_pool_pe_b_peij_3_3_q_k) );
  XOR2_X1 pool_pool_pe_b_peij_3_3_add_U11 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_3_q_k), .Z(pool_pool_pe_b_peij_3_3_add_notb[0])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_3_add_U10 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_3_q_k), .Z(pool_pool_pe_b_peij_3_3_add_notb[10])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_3_add_U9 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_3_q_k), .Z(pool_pool_pe_b_peij_3_3_add_notb[1])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_3_add_U8 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_3_q_k), .Z(pool_pool_pe_b_peij_3_3_add_notb[2])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_3_add_U7 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_3_q_k), .Z(pool_pool_pe_b_peij_3_3_add_notb[3])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_3_add_U6 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_3_q_k), .Z(pool_pool_pe_b_peij_3_3_add_notb[4])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_3_add_U5 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_3_q_k), .Z(pool_pool_pe_b_peij_3_3_add_notb[5])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_3_add_U4 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_3_q_k), .Z(pool_pool_pe_b_peij_3_3_add_notb[6])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_3_add_U3 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_3_q_k), .Z(pool_pool_pe_b_peij_3_3_add_notb[7])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_3_add_U2 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_3_q_k), .Z(pool_pool_pe_b_peij_3_3_add_notb[8])
         );
  XOR2_X1 pool_pool_pe_b_peij_3_3_add_U1 ( .A(1'b0), .B(
        pool_pool_pe_b_peij_3_3_q_k), .Z(pool_pool_pe_b_peij_3_3_add_notb[9])
         );
  INV_X2 pool_pool_pe_b_peij_3_3_add_fai_0_U2 ( .A(
        pool_pool_pe_b_peij_3_3_add_fai_0_n4), .ZN(
        pool_pool_pe_b_peij_3_3_add_cprop[1]) );
  XOR2_X1 pool_pool_pe_b_peij_3_3_add_fai_0_U4 ( .A(pool_pool_pe_b_o_data[0]), 
        .B(pool_pool_pe_b_peij_3_3_add_notb[0]), .Z(
        pool_pool_pe_b_peij_3_3_add_fai_0_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_3_add_fai_0_U3 ( .A(
        pool_pool_pe_b_peij_3_3_q_k), .B(pool_pool_pe_b_peij_3_3_add_fai_0_n5), 
        .Z(pool_pool_pe_b_peij_3_3_d_acc[0]) );
  AOI22_X2 pool_pool_pe_b_peij_3_3_add_fai_0_U1 ( .A1(
        pool_pool_pe_b_peij_3_3_add_notb[0]), .A2(pool_pool_pe_b_o_data[0]), 
        .B1(pool_pool_pe_b_peij_3_3_add_fai_0_n5), .B2(
        pool_pool_pe_b_peij_3_3_q_k), .ZN(pool_pool_pe_b_peij_3_3_add_fai_0_n4) );
  INV_X2 pool_pool_pe_b_peij_3_3_add_fai_1_U2 ( .A(
        pool_pool_pe_b_peij_3_3_add_fai_1_n4), .ZN(
        pool_pool_pe_b_peij_3_3_add_cprop[2]) );
  XOR2_X1 pool_pool_pe_b_peij_3_3_add_fai_1_U4 ( .A(pool_pool_pe_b_o_data[1]), 
        .B(pool_pool_pe_b_peij_3_3_add_notb[1]), .Z(
        pool_pool_pe_b_peij_3_3_add_fai_1_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_3_add_fai_1_U3 ( .A(
        pool_pool_pe_b_peij_3_3_add_cprop[1]), .B(
        pool_pool_pe_b_peij_3_3_add_fai_1_n5), .Z(
        pool_pool_pe_b_peij_3_3_d_acc[1]) );
  AOI22_X2 pool_pool_pe_b_peij_3_3_add_fai_1_U1 ( .A1(
        pool_pool_pe_b_peij_3_3_add_notb[1]), .A2(pool_pool_pe_b_o_data[1]), 
        .B1(pool_pool_pe_b_peij_3_3_add_fai_1_n5), .B2(
        pool_pool_pe_b_peij_3_3_add_cprop[1]), .ZN(
        pool_pool_pe_b_peij_3_3_add_fai_1_n4) );
  INV_X2 pool_pool_pe_b_peij_3_3_add_fai_2_U2 ( .A(
        pool_pool_pe_b_peij_3_3_add_fai_2_n4), .ZN(
        pool_pool_pe_b_peij_3_3_add_cprop[3]) );
  XOR2_X1 pool_pool_pe_b_peij_3_3_add_fai_2_U4 ( .A(pool_pool_pe_b_o_data[2]), 
        .B(pool_pool_pe_b_peij_3_3_add_notb[2]), .Z(
        pool_pool_pe_b_peij_3_3_add_fai_2_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_3_add_fai_2_U3 ( .A(
        pool_pool_pe_b_peij_3_3_add_cprop[2]), .B(
        pool_pool_pe_b_peij_3_3_add_fai_2_n5), .Z(
        pool_pool_pe_b_peij_3_3_d_acc[2]) );
  AOI22_X2 pool_pool_pe_b_peij_3_3_add_fai_2_U1 ( .A1(
        pool_pool_pe_b_peij_3_3_add_notb[2]), .A2(pool_pool_pe_b_o_data[2]), 
        .B1(pool_pool_pe_b_peij_3_3_add_fai_2_n5), .B2(
        pool_pool_pe_b_peij_3_3_add_cprop[2]), .ZN(
        pool_pool_pe_b_peij_3_3_add_fai_2_n4) );
  INV_X2 pool_pool_pe_b_peij_3_3_add_fai_3_U2 ( .A(
        pool_pool_pe_b_peij_3_3_add_fai_3_n4), .ZN(
        pool_pool_pe_b_peij_3_3_add_cprop[4]) );
  XOR2_X1 pool_pool_pe_b_peij_3_3_add_fai_3_U4 ( .A(pool_pool_pe_b_o_data[3]), 
        .B(pool_pool_pe_b_peij_3_3_add_notb[3]), .Z(
        pool_pool_pe_b_peij_3_3_add_fai_3_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_3_add_fai_3_U3 ( .A(
        pool_pool_pe_b_peij_3_3_add_cprop[3]), .B(
        pool_pool_pe_b_peij_3_3_add_fai_3_n5), .Z(
        pool_pool_pe_b_peij_3_3_d_acc[3]) );
  AOI22_X2 pool_pool_pe_b_peij_3_3_add_fai_3_U1 ( .A1(
        pool_pool_pe_b_peij_3_3_add_notb[3]), .A2(pool_pool_pe_b_o_data[3]), 
        .B1(pool_pool_pe_b_peij_3_3_add_fai_3_n5), .B2(
        pool_pool_pe_b_peij_3_3_add_cprop[3]), .ZN(
        pool_pool_pe_b_peij_3_3_add_fai_3_n4) );
  INV_X2 pool_pool_pe_b_peij_3_3_add_fai_4_U2 ( .A(
        pool_pool_pe_b_peij_3_3_add_fai_4_n4), .ZN(
        pool_pool_pe_b_peij_3_3_add_cprop[5]) );
  XOR2_X1 pool_pool_pe_b_peij_3_3_add_fai_4_U4 ( .A(pool_pool_pe_b_o_data[4]), 
        .B(pool_pool_pe_b_peij_3_3_add_notb[4]), .Z(
        pool_pool_pe_b_peij_3_3_add_fai_4_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_3_add_fai_4_U3 ( .A(
        pool_pool_pe_b_peij_3_3_add_cprop[4]), .B(
        pool_pool_pe_b_peij_3_3_add_fai_4_n5), .Z(
        pool_pool_pe_b_peij_3_3_d_acc[4]) );
  AOI22_X2 pool_pool_pe_b_peij_3_3_add_fai_4_U1 ( .A1(
        pool_pool_pe_b_peij_3_3_add_notb[4]), .A2(pool_pool_pe_b_o_data[4]), 
        .B1(pool_pool_pe_b_peij_3_3_add_fai_4_n5), .B2(
        pool_pool_pe_b_peij_3_3_add_cprop[4]), .ZN(
        pool_pool_pe_b_peij_3_3_add_fai_4_n4) );
  INV_X2 pool_pool_pe_b_peij_3_3_add_fai_5_U2 ( .A(
        pool_pool_pe_b_peij_3_3_add_fai_5_n4), .ZN(
        pool_pool_pe_b_peij_3_3_add_cprop[6]) );
  XOR2_X1 pool_pool_pe_b_peij_3_3_add_fai_5_U4 ( .A(pool_pool_pe_b_o_data[5]), 
        .B(pool_pool_pe_b_peij_3_3_add_notb[5]), .Z(
        pool_pool_pe_b_peij_3_3_add_fai_5_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_3_add_fai_5_U3 ( .A(
        pool_pool_pe_b_peij_3_3_add_cprop[5]), .B(
        pool_pool_pe_b_peij_3_3_add_fai_5_n5), .Z(
        pool_pool_pe_b_peij_3_3_d_acc[5]) );
  AOI22_X2 pool_pool_pe_b_peij_3_3_add_fai_5_U1 ( .A1(
        pool_pool_pe_b_peij_3_3_add_notb[5]), .A2(pool_pool_pe_b_o_data[5]), 
        .B1(pool_pool_pe_b_peij_3_3_add_fai_5_n5), .B2(
        pool_pool_pe_b_peij_3_3_add_cprop[5]), .ZN(
        pool_pool_pe_b_peij_3_3_add_fai_5_n4) );
  INV_X2 pool_pool_pe_b_peij_3_3_add_fai_6_U2 ( .A(
        pool_pool_pe_b_peij_3_3_add_fai_6_n4), .ZN(
        pool_pool_pe_b_peij_3_3_add_cprop[7]) );
  XOR2_X1 pool_pool_pe_b_peij_3_3_add_fai_6_U4 ( .A(pool_pool_pe_b_o_data[6]), 
        .B(pool_pool_pe_b_peij_3_3_add_notb[6]), .Z(
        pool_pool_pe_b_peij_3_3_add_fai_6_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_3_add_fai_6_U3 ( .A(
        pool_pool_pe_b_peij_3_3_add_cprop[6]), .B(
        pool_pool_pe_b_peij_3_3_add_fai_6_n5), .Z(
        pool_pool_pe_b_peij_3_3_d_acc[6]) );
  AOI22_X2 pool_pool_pe_b_peij_3_3_add_fai_6_U1 ( .A1(
        pool_pool_pe_b_peij_3_3_add_notb[6]), .A2(pool_pool_pe_b_o_data[6]), 
        .B1(pool_pool_pe_b_peij_3_3_add_fai_6_n5), .B2(
        pool_pool_pe_b_peij_3_3_add_cprop[6]), .ZN(
        pool_pool_pe_b_peij_3_3_add_fai_6_n4) );
  INV_X2 pool_pool_pe_b_peij_3_3_add_fai_7_U2 ( .A(
        pool_pool_pe_b_peij_3_3_add_fai_7_n4), .ZN(
        pool_pool_pe_b_peij_3_3_add_cprop[8]) );
  XOR2_X1 pool_pool_pe_b_peij_3_3_add_fai_7_U4 ( .A(pool_pool_pe_b_o_data[7]), 
        .B(pool_pool_pe_b_peij_3_3_add_notb[7]), .Z(
        pool_pool_pe_b_peij_3_3_add_fai_7_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_3_add_fai_7_U3 ( .A(
        pool_pool_pe_b_peij_3_3_add_cprop[7]), .B(
        pool_pool_pe_b_peij_3_3_add_fai_7_n5), .Z(
        pool_pool_pe_b_peij_3_3_d_acc[7]) );
  AOI22_X2 pool_pool_pe_b_peij_3_3_add_fai_7_U1 ( .A1(
        pool_pool_pe_b_peij_3_3_add_notb[7]), .A2(pool_pool_pe_b_o_data[7]), 
        .B1(pool_pool_pe_b_peij_3_3_add_fai_7_n5), .B2(
        pool_pool_pe_b_peij_3_3_add_cprop[7]), .ZN(
        pool_pool_pe_b_peij_3_3_add_fai_7_n4) );
  INV_X2 pool_pool_pe_b_peij_3_3_add_fai_8_U2 ( .A(
        pool_pool_pe_b_peij_3_3_add_fai_8_n4), .ZN(
        pool_pool_pe_b_peij_3_3_add_cprop[9]) );
  XOR2_X1 pool_pool_pe_b_peij_3_3_add_fai_8_U4 ( .A(pool_pool_pe_b_o_data[8]), 
        .B(pool_pool_pe_b_peij_3_3_add_notb[8]), .Z(
        pool_pool_pe_b_peij_3_3_add_fai_8_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_3_add_fai_8_U3 ( .A(
        pool_pool_pe_b_peij_3_3_add_cprop[8]), .B(
        pool_pool_pe_b_peij_3_3_add_fai_8_n5), .Z(
        pool_pool_pe_b_peij_3_3_d_acc[8]) );
  AOI22_X2 pool_pool_pe_b_peij_3_3_add_fai_8_U1 ( .A1(
        pool_pool_pe_b_peij_3_3_add_notb[8]), .A2(pool_pool_pe_b_o_data[8]), 
        .B1(pool_pool_pe_b_peij_3_3_add_fai_8_n5), .B2(
        pool_pool_pe_b_peij_3_3_add_cprop[8]), .ZN(
        pool_pool_pe_b_peij_3_3_add_fai_8_n4) );
  INV_X2 pool_pool_pe_b_peij_3_3_add_fai_9_U2 ( .A(
        pool_pool_pe_b_peij_3_3_add_fai_9_n4), .ZN(
        pool_pool_pe_b_peij_3_3_add_cprop[10]) );
  XOR2_X1 pool_pool_pe_b_peij_3_3_add_fai_9_U4 ( .A(pool_pool_pe_b_o_data[9]), 
        .B(pool_pool_pe_b_peij_3_3_add_notb[9]), .Z(
        pool_pool_pe_b_peij_3_3_add_fai_9_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_3_add_fai_9_U3 ( .A(
        pool_pool_pe_b_peij_3_3_add_cprop[9]), .B(
        pool_pool_pe_b_peij_3_3_add_fai_9_n5), .Z(
        pool_pool_pe_b_peij_3_3_d_acc[9]) );
  AOI22_X2 pool_pool_pe_b_peij_3_3_add_fai_9_U1 ( .A1(
        pool_pool_pe_b_peij_3_3_add_notb[9]), .A2(pool_pool_pe_b_o_data[9]), 
        .B1(pool_pool_pe_b_peij_3_3_add_fai_9_n5), .B2(
        pool_pool_pe_b_peij_3_3_add_cprop[9]), .ZN(
        pool_pool_pe_b_peij_3_3_add_fai_9_n4) );
  INV_X2 pool_pool_pe_b_peij_3_3_add_fai_10_U2 ( .A(
        pool_pool_pe_b_peij_3_3_add_fai_10_n4), .ZN(
        pool_pool_pe_b_peij_3_3_add_c_out) );
  XOR2_X1 pool_pool_pe_b_peij_3_3_add_fai_10_U4 ( .A(pool_pool_pe_b_o_data[10]), .B(pool_pool_pe_b_peij_3_3_add_notb[10]), .Z(
        pool_pool_pe_b_peij_3_3_add_fai_10_n5) );
  XOR2_X1 pool_pool_pe_b_peij_3_3_add_fai_10_U3 ( .A(
        pool_pool_pe_b_peij_3_3_add_cprop[10]), .B(
        pool_pool_pe_b_peij_3_3_add_fai_10_n5), .Z(
        pool_pool_pe_b_peij_3_3_d_acc[10]) );
  AOI22_X2 pool_pool_pe_b_peij_3_3_add_fai_10_U1 ( .A1(
        pool_pool_pe_b_peij_3_3_add_notb[10]), .A2(pool_pool_pe_b_o_data[10]), 
        .B1(pool_pool_pe_b_peij_3_3_add_fai_10_n5), .B2(
        pool_pool_pe_b_peij_3_3_add_cprop[10]), .ZN(
        pool_pool_pe_b_peij_3_3_add_fai_10_n4) );
  INV_X2 pool_pool_count_U13 ( .A(1'b1), .ZN(pool_pool_count_n12) );
  INV_X2 pool_pool_count_U12 ( .A(pool_rst_cnt), .ZN(pool_pool_count_n10) );
  INV_X2 pool_pool_count_U8 ( .A(pool_pool_count_n13), .ZN(pool_pool_count_n9)
         );
  INV_X2 pool_pool_count_U6 ( .A(pool_pool_count_n8), .ZN(pool_pool_count_n3)
         );
  INV_X2 pool_pool_count_U5 ( .A(pool_pool_count_n11), .ZN(pool_pool_count_n1)
         );
  DFFR_X1 pool_pool_count_cnt_out_reg_1_ ( .D(pool_pool_count_n15), .CK(clk), 
        .RN(pool_pool_count_n10), .Q(pool_pool_cnt_1_), .QN(pool_pool_count_n7) );
  DFFR_X1 pool_pool_count_cnt_out_reg_0_ ( .D(pool_pool_count_n17), .CK(clk), 
        .RN(pool_pool_count_n10), .Q(pool_pool_cnt_0_), .QN(pool_pool_count_n2) );
  DFFR_X1 pool_pool_count_terminal_cnt_reg ( .D(pool_pool_count_n18), .CK(clk), 
        .RN(pool_pool_count_n10), .Q(pool_tc), .QN(pool_pool_count_n4) );
  NAND2_X2 pool_pool_count_U11 ( .A1(pool_en_cnt), .A2(pool_pool_count_n4), 
        .ZN(pool_pool_count_n6) );
  OAI22_X2 pool_pool_count_U10 ( .A1(pool_pool_count_n1), .A2(
        pool_pool_count_n6), .B1(pool_en_cnt), .B2(pool_pool_count_n4), .ZN(
        pool_pool_count_n18) );
  OAI22_X2 pool_pool_count_U9 ( .A1(pool_en_cnt), .A2(pool_pool_count_n2), 
        .B1(pool_pool_cnt_0_), .B2(pool_pool_count_n6), .ZN(
        pool_pool_count_n17) );
  OAI21_X2 pool_pool_count_U7 ( .B1(pool_pool_cnt_0_), .B2(pool_tc), .A(
        pool_en_cnt), .ZN(pool_pool_count_n8) );
  OR3_X4 pool_pool_count_U4 ( .A1(pool_pool_count_n6), .A2(pool_pool_cnt_1_), 
        .A3(pool_pool_count_n2), .ZN(pool_pool_count_n5) );
  OAI21_X2 pool_pool_count_U3 ( .B1(pool_pool_count_n3), .B2(
        pool_pool_count_n7), .A(pool_pool_count_n5), .ZN(pool_pool_count_n15)
         );
  XOR2_X1 pool_pool_count_U17 ( .A(pool_pool_cnt_1_), .B(1'b1), .Z(
        pool_pool_count_n13) );
  OAI33_X1 pool_pool_count_U14 ( .A1(pool_pool_count_n12), .A2(
        pool_pool_cnt_0_), .A3(pool_pool_count_n13), .B1(pool_pool_count_n2), 
        .B2(1'b1), .B3(pool_pool_count_n9), .ZN(pool_pool_count_n11) );
  INV_X2 pool_pool_shift_row0_U13 ( .A(pool_pool_pe_b_o_data[168]), .ZN(
        pool_pool_shift_row0_n4) );
  INV_X2 pool_pool_shift_row0_U12 ( .A(pool_pool_pe_b_o_data[135]), .ZN(
        pool_pool_shift_row0_n3) );
  INV_X2 pool_pool_shift_row0_U11 ( .A(pool_pool_pe_b_o_data[146]), .ZN(
        pool_pool_shift_row0_n2) );
  INV_X2 pool_pool_shift_row0_U10 ( .A(pool_pool_pe_b_o_data[157]), .ZN(
        pool_pool_shift_row0_n1) );
  XOR2_X1 pool_pool_shift_row0_U25 ( .A(pool_pool_pe_b_o_data[167]), .B(
        pool_pool_pe_b_o_data[166]), .Z(o_pool_1[12]) );
  XOR2_X1 pool_pool_shift_row0_U24 ( .A(pool_pool_shift_row0_n4), .B(
        pool_pool_shift_row0_n12), .Z(o_pool_1[13]) );
  XOR2_X1 pool_pool_shift_row0_U23 ( .A(pool_pool_pe_b_o_data[169]), .B(
        pool_pool_shift_row0_n11), .Z(o_pool_1[14]) );
  XOR2_X1 pool_pool_shift_row0_U22 ( .A(pool_pool_pe_b_o_data[156]), .B(
        pool_pool_pe_b_o_data[155]), .Z(o_pool_1[8]) );
  XOR2_X1 pool_pool_shift_row0_U21 ( .A(pool_pool_shift_row0_n1), .B(
        pool_pool_shift_row0_n10), .Z(o_pool_1[9]) );
  XOR2_X1 pool_pool_shift_row0_U20 ( .A(pool_pool_pe_b_o_data[158]), .B(
        pool_pool_shift_row0_n9), .Z(o_pool_1[10]) );
  XOR2_X1 pool_pool_shift_row0_U19 ( .A(pool_pool_pe_b_o_data[145]), .B(
        pool_pool_pe_b_o_data[144]), .Z(o_pool_1[4]) );
  XOR2_X1 pool_pool_shift_row0_U18 ( .A(pool_pool_shift_row0_n2), .B(
        pool_pool_shift_row0_n8), .Z(o_pool_1[5]) );
  XOR2_X1 pool_pool_shift_row0_U17 ( .A(pool_pool_pe_b_o_data[147]), .B(
        pool_pool_shift_row0_n7), .Z(o_pool_1[6]) );
  XOR2_X1 pool_pool_shift_row0_U16 ( .A(pool_pool_pe_b_o_data[134]), .B(
        pool_pool_pe_b_o_data[133]), .Z(o_pool_1[0]) );
  XOR2_X1 pool_pool_shift_row0_U15 ( .A(pool_pool_shift_row0_n3), .B(
        pool_pool_shift_row0_n6), .Z(o_pool_1[1]) );
  XOR2_X1 pool_pool_shift_row0_U14 ( .A(pool_pool_pe_b_o_data[136]), .B(
        pool_pool_shift_row0_n5), .Z(o_pool_1[2]) );
  NAND2_X2 pool_pool_shift_row0_U9 ( .A1(pool_pool_pe_b_o_data[167]), .A2(
        pool_pool_pe_b_o_data[166]), .ZN(pool_pool_shift_row0_n12) );
  NOR2_X2 pool_pool_shift_row0_U8 ( .A1(pool_pool_shift_row0_n12), .A2(
        pool_pool_shift_row0_n4), .ZN(pool_pool_shift_row0_n11) );
  NAND2_X2 pool_pool_shift_row0_U7 ( .A1(pool_pool_pe_b_o_data[156]), .A2(
        pool_pool_pe_b_o_data[155]), .ZN(pool_pool_shift_row0_n10) );
  NOR2_X2 pool_pool_shift_row0_U6 ( .A1(pool_pool_shift_row0_n10), .A2(
        pool_pool_shift_row0_n1), .ZN(pool_pool_shift_row0_n9) );
  NAND2_X2 pool_pool_shift_row0_U5 ( .A1(pool_pool_pe_b_o_data[145]), .A2(
        pool_pool_pe_b_o_data[144]), .ZN(pool_pool_shift_row0_n8) );
  NOR2_X2 pool_pool_shift_row0_U4 ( .A1(pool_pool_shift_row0_n8), .A2(
        pool_pool_shift_row0_n2), .ZN(pool_pool_shift_row0_n7) );
  NAND2_X2 pool_pool_shift_row0_U3 ( .A1(pool_pool_pe_b_o_data[134]), .A2(
        pool_pool_pe_b_o_data[133]), .ZN(pool_pool_shift_row0_n6) );
  NOR2_X2 pool_pool_shift_row0_U2 ( .A1(pool_pool_shift_row0_n6), .A2(
        pool_pool_shift_row0_n3), .ZN(pool_pool_shift_row0_n5) );
  INV_X2 pool_pool_shift_row1_U13 ( .A(pool_pool_pe_b_o_data[91]), .ZN(
        pool_pool_shift_row1_n4) );
  INV_X2 pool_pool_shift_row1_U12 ( .A(pool_pool_pe_b_o_data[102]), .ZN(
        pool_pool_shift_row1_n3) );
  INV_X2 pool_pool_shift_row1_U11 ( .A(pool_pool_pe_b_o_data[113]), .ZN(
        pool_pool_shift_row1_n2) );
  INV_X2 pool_pool_shift_row1_U10 ( .A(pool_pool_pe_b_o_data[124]), .ZN(
        pool_pool_shift_row1_n1) );
  XOR2_X1 pool_pool_shift_row1_U25 ( .A(pool_pool_pe_b_o_data[123]), .B(
        pool_pool_pe_b_o_data[122]), .Z(o_pool_2[12]) );
  XOR2_X1 pool_pool_shift_row1_U24 ( .A(pool_pool_shift_row1_n1), .B(
        pool_pool_shift_row1_n13), .Z(o_pool_2[13]) );
  XOR2_X1 pool_pool_shift_row1_U23 ( .A(pool_pool_pe_b_o_data[125]), .B(
        pool_pool_shift_row1_n14), .Z(o_pool_2[14]) );
  XOR2_X1 pool_pool_shift_row1_U22 ( .A(pool_pool_pe_b_o_data[112]), .B(
        pool_pool_pe_b_o_data[111]), .Z(o_pool_2[8]) );
  XOR2_X1 pool_pool_shift_row1_U21 ( .A(pool_pool_shift_row1_n2), .B(
        pool_pool_shift_row1_n15), .Z(o_pool_2[9]) );
  XOR2_X1 pool_pool_shift_row1_U20 ( .A(pool_pool_pe_b_o_data[114]), .B(
        pool_pool_shift_row1_n16), .Z(o_pool_2[10]) );
  XOR2_X1 pool_pool_shift_row1_U19 ( .A(pool_pool_pe_b_o_data[101]), .B(
        pool_pool_pe_b_o_data[100]), .Z(o_pool_2[4]) );
  XOR2_X1 pool_pool_shift_row1_U18 ( .A(pool_pool_shift_row1_n3), .B(
        pool_pool_shift_row1_n17), .Z(o_pool_2[5]) );
  XOR2_X1 pool_pool_shift_row1_U17 ( .A(pool_pool_pe_b_o_data[103]), .B(
        pool_pool_shift_row1_n18), .Z(o_pool_2[6]) );
  XOR2_X1 pool_pool_shift_row1_U16 ( .A(pool_pool_pe_b_o_data[90]), .B(
        pool_pool_pe_b_o_data[89]), .Z(o_pool_2[0]) );
  XOR2_X1 pool_pool_shift_row1_U15 ( .A(pool_pool_shift_row1_n4), .B(
        pool_pool_shift_row1_n19), .Z(o_pool_2[1]) );
  XOR2_X1 pool_pool_shift_row1_U14 ( .A(pool_pool_pe_b_o_data[92]), .B(
        pool_pool_shift_row1_n20), .Z(o_pool_2[2]) );
  NAND2_X2 pool_pool_shift_row1_U9 ( .A1(pool_pool_pe_b_o_data[123]), .A2(
        pool_pool_pe_b_o_data[122]), .ZN(pool_pool_shift_row1_n13) );
  NOR2_X2 pool_pool_shift_row1_U8 ( .A1(pool_pool_shift_row1_n13), .A2(
        pool_pool_shift_row1_n1), .ZN(pool_pool_shift_row1_n14) );
  NAND2_X2 pool_pool_shift_row1_U7 ( .A1(pool_pool_pe_b_o_data[112]), .A2(
        pool_pool_pe_b_o_data[111]), .ZN(pool_pool_shift_row1_n15) );
  NOR2_X2 pool_pool_shift_row1_U6 ( .A1(pool_pool_shift_row1_n15), .A2(
        pool_pool_shift_row1_n2), .ZN(pool_pool_shift_row1_n16) );
  NAND2_X2 pool_pool_shift_row1_U5 ( .A1(pool_pool_pe_b_o_data[101]), .A2(
        pool_pool_pe_b_o_data[100]), .ZN(pool_pool_shift_row1_n17) );
  NOR2_X2 pool_pool_shift_row1_U4 ( .A1(pool_pool_shift_row1_n17), .A2(
        pool_pool_shift_row1_n3), .ZN(pool_pool_shift_row1_n18) );
  NAND2_X2 pool_pool_shift_row1_U3 ( .A1(pool_pool_pe_b_o_data[90]), .A2(
        pool_pool_pe_b_o_data[89]), .ZN(pool_pool_shift_row1_n19) );
  NOR2_X2 pool_pool_shift_row1_U2 ( .A1(pool_pool_shift_row1_n19), .A2(
        pool_pool_shift_row1_n4), .ZN(pool_pool_shift_row1_n20) );
  INV_X2 pool_pool_shift_row2_U13 ( .A(pool_pool_pe_b_o_data[47]), .ZN(
        pool_pool_shift_row2_n4) );
  INV_X2 pool_pool_shift_row2_U12 ( .A(pool_pool_pe_b_o_data[58]), .ZN(
        pool_pool_shift_row2_n3) );
  INV_X2 pool_pool_shift_row2_U11 ( .A(pool_pool_pe_b_o_data[69]), .ZN(
        pool_pool_shift_row2_n2) );
  INV_X2 pool_pool_shift_row2_U10 ( .A(pool_pool_pe_b_o_data[80]), .ZN(
        pool_pool_shift_row2_n1) );
  XOR2_X1 pool_pool_shift_row2_U25 ( .A(pool_pool_pe_b_o_data[79]), .B(
        pool_pool_pe_b_o_data[78]), .Z(o_pool_3[12]) );
  XOR2_X1 pool_pool_shift_row2_U24 ( .A(pool_pool_shift_row2_n1), .B(
        pool_pool_shift_row2_n13), .Z(o_pool_3[13]) );
  XOR2_X1 pool_pool_shift_row2_U23 ( .A(pool_pool_pe_b_o_data[81]), .B(
        pool_pool_shift_row2_n14), .Z(o_pool_3[14]) );
  XOR2_X1 pool_pool_shift_row2_U22 ( .A(pool_pool_pe_b_o_data[68]), .B(
        pool_pool_pe_b_o_data[67]), .Z(o_pool_3[8]) );
  XOR2_X1 pool_pool_shift_row2_U21 ( .A(pool_pool_shift_row2_n2), .B(
        pool_pool_shift_row2_n15), .Z(o_pool_3[9]) );
  XOR2_X1 pool_pool_shift_row2_U20 ( .A(pool_pool_pe_b_o_data[70]), .B(
        pool_pool_shift_row2_n16), .Z(o_pool_3[10]) );
  XOR2_X1 pool_pool_shift_row2_U19 ( .A(pool_pool_pe_b_o_data[57]), .B(
        pool_pool_pe_b_o_data[56]), .Z(o_pool_3[4]) );
  XOR2_X1 pool_pool_shift_row2_U18 ( .A(pool_pool_shift_row2_n3), .B(
        pool_pool_shift_row2_n17), .Z(o_pool_3[5]) );
  XOR2_X1 pool_pool_shift_row2_U17 ( .A(pool_pool_pe_b_o_data[59]), .B(
        pool_pool_shift_row2_n18), .Z(o_pool_3[6]) );
  XOR2_X1 pool_pool_shift_row2_U16 ( .A(pool_pool_pe_b_o_data[46]), .B(
        pool_pool_pe_b_o_data[45]), .Z(o_pool_3[0]) );
  XOR2_X1 pool_pool_shift_row2_U15 ( .A(pool_pool_shift_row2_n4), .B(
        pool_pool_shift_row2_n19), .Z(o_pool_3[1]) );
  XOR2_X1 pool_pool_shift_row2_U14 ( .A(pool_pool_pe_b_o_data[48]), .B(
        pool_pool_shift_row2_n20), .Z(o_pool_3[2]) );
  NAND2_X2 pool_pool_shift_row2_U9 ( .A1(pool_pool_pe_b_o_data[79]), .A2(
        pool_pool_pe_b_o_data[78]), .ZN(pool_pool_shift_row2_n13) );
  NOR2_X2 pool_pool_shift_row2_U8 ( .A1(pool_pool_shift_row2_n13), .A2(
        pool_pool_shift_row2_n1), .ZN(pool_pool_shift_row2_n14) );
  NAND2_X2 pool_pool_shift_row2_U7 ( .A1(pool_pool_pe_b_o_data[68]), .A2(
        pool_pool_pe_b_o_data[67]), .ZN(pool_pool_shift_row2_n15) );
  NOR2_X2 pool_pool_shift_row2_U6 ( .A1(pool_pool_shift_row2_n15), .A2(
        pool_pool_shift_row2_n2), .ZN(pool_pool_shift_row2_n16) );
  NAND2_X2 pool_pool_shift_row2_U5 ( .A1(pool_pool_pe_b_o_data[57]), .A2(
        pool_pool_pe_b_o_data[56]), .ZN(pool_pool_shift_row2_n17) );
  NOR2_X2 pool_pool_shift_row2_U4 ( .A1(pool_pool_shift_row2_n17), .A2(
        pool_pool_shift_row2_n3), .ZN(pool_pool_shift_row2_n18) );
  NAND2_X2 pool_pool_shift_row2_U3 ( .A1(pool_pool_pe_b_o_data[46]), .A2(
        pool_pool_pe_b_o_data[45]), .ZN(pool_pool_shift_row2_n19) );
  NOR2_X2 pool_pool_shift_row2_U2 ( .A1(pool_pool_shift_row2_n19), .A2(
        pool_pool_shift_row2_n4), .ZN(pool_pool_shift_row2_n20) );
  INV_X2 pool_pool_shift_row3_U13 ( .A(pool_pool_pe_b_o_data[3]), .ZN(
        pool_pool_shift_row3_n4) );
  INV_X2 pool_pool_shift_row3_U12 ( .A(pool_pool_pe_b_o_data[14]), .ZN(
        pool_pool_shift_row3_n3) );
  INV_X2 pool_pool_shift_row3_U11 ( .A(pool_pool_pe_b_o_data[25]), .ZN(
        pool_pool_shift_row3_n2) );
  INV_X2 pool_pool_shift_row3_U10 ( .A(pool_pool_pe_b_o_data[36]), .ZN(
        pool_pool_shift_row3_n1) );
  XOR2_X1 pool_pool_shift_row3_U25 ( .A(pool_pool_pe_b_o_data[35]), .B(
        pool_pool_pe_b_o_data[34]), .Z(o_pool_4[12]) );
  XOR2_X1 pool_pool_shift_row3_U24 ( .A(pool_pool_shift_row3_n1), .B(
        pool_pool_shift_row3_n13), .Z(o_pool_4[13]) );
  XOR2_X1 pool_pool_shift_row3_U23 ( .A(pool_pool_pe_b_o_data[37]), .B(
        pool_pool_shift_row3_n14), .Z(o_pool_4[14]) );
  XOR2_X1 pool_pool_shift_row3_U22 ( .A(pool_pool_pe_b_o_data[24]), .B(
        pool_pool_pe_b_o_data[23]), .Z(o_pool_4[8]) );
  XOR2_X1 pool_pool_shift_row3_U21 ( .A(pool_pool_shift_row3_n2), .B(
        pool_pool_shift_row3_n15), .Z(o_pool_4[9]) );
  XOR2_X1 pool_pool_shift_row3_U20 ( .A(pool_pool_pe_b_o_data[26]), .B(
        pool_pool_shift_row3_n16), .Z(o_pool_4[10]) );
  XOR2_X1 pool_pool_shift_row3_U19 ( .A(pool_pool_pe_b_o_data[13]), .B(
        pool_pool_pe_b_o_data[12]), .Z(o_pool_4[4]) );
  XOR2_X1 pool_pool_shift_row3_U18 ( .A(pool_pool_shift_row3_n3), .B(
        pool_pool_shift_row3_n17), .Z(o_pool_4[5]) );
  XOR2_X1 pool_pool_shift_row3_U17 ( .A(pool_pool_pe_b_o_data[15]), .B(
        pool_pool_shift_row3_n18), .Z(o_pool_4[6]) );
  XOR2_X1 pool_pool_shift_row3_U16 ( .A(pool_pool_pe_b_o_data[2]), .B(
        pool_pool_pe_b_o_data[1]), .Z(o_pool_4[0]) );
  XOR2_X1 pool_pool_shift_row3_U15 ( .A(pool_pool_shift_row3_n4), .B(
        pool_pool_shift_row3_n19), .Z(o_pool_4[1]) );
  XOR2_X1 pool_pool_shift_row3_U14 ( .A(pool_pool_pe_b_o_data[4]), .B(
        pool_pool_shift_row3_n20), .Z(o_pool_4[2]) );
  NAND2_X2 pool_pool_shift_row3_U9 ( .A1(pool_pool_pe_b_o_data[35]), .A2(
        pool_pool_pe_b_o_data[34]), .ZN(pool_pool_shift_row3_n13) );
  NOR2_X2 pool_pool_shift_row3_U8 ( .A1(pool_pool_shift_row3_n13), .A2(
        pool_pool_shift_row3_n1), .ZN(pool_pool_shift_row3_n14) );
  NAND2_X2 pool_pool_shift_row3_U7 ( .A1(pool_pool_pe_b_o_data[24]), .A2(
        pool_pool_pe_b_o_data[23]), .ZN(pool_pool_shift_row3_n15) );
  NOR2_X2 pool_pool_shift_row3_U6 ( .A1(pool_pool_shift_row3_n15), .A2(
        pool_pool_shift_row3_n2), .ZN(pool_pool_shift_row3_n16) );
  NAND2_X2 pool_pool_shift_row3_U5 ( .A1(pool_pool_pe_b_o_data[13]), .A2(
        pool_pool_pe_b_o_data[12]), .ZN(pool_pool_shift_row3_n17) );
  NOR2_X2 pool_pool_shift_row3_U4 ( .A1(pool_pool_shift_row3_n17), .A2(
        pool_pool_shift_row3_n3), .ZN(pool_pool_shift_row3_n18) );
  NAND2_X2 pool_pool_shift_row3_U3 ( .A1(pool_pool_pe_b_o_data[2]), .A2(
        pool_pool_pe_b_o_data[1]), .ZN(pool_pool_shift_row3_n19) );
  NOR2_X2 pool_pool_shift_row3_U2 ( .A1(pool_pool_shift_row3_n19), .A2(
        pool_pool_shift_row3_n4), .ZN(pool_pool_shift_row3_n20) );
  INV_X2 pool_fsm_U27 ( .A(done), .ZN(pool_fsm_n18) );
  INV_X2 pool_fsm_U26 ( .A(rst_fsm), .ZN(pool_fsm_n17) );
  INV_X2 pool_fsm_U21 ( .A(pool_sync_clr), .ZN(pool_fsm_n10) );
  INV_X2 pool_fsm_U20 ( .A(pool_fsm_n11), .ZN(pool_rst_cnt) );
  INV_X2 pool_fsm_U19 ( .A(pool_fsm_n16), .ZN(pool_fsm_n5) );
  INV_X1 pool_fsm_U18 ( .A(pool_fsm_N11), .ZN(pool_fsm_n4) );
  INV_X1 pool_fsm_U17 ( .A(pool_fsm_n4), .ZN(pool_ld_h) );
  INV_X2 pool_fsm_U16 ( .A(pool_fsm_n19), .ZN(pool_fsm_n2) );
  INV_X1 pool_fsm_U3 ( .A(pool_fsm_n2), .ZN(pool_sel0) );
  SNPS_CLOCK_GATE_HIGH_avr_pooling_fsm pool_fsm_clk_gate_current_state_reg ( 
        .CLK(clk), .EN(pool_fsm_N31), .ENCLK(pool_fsm_net424), .TE(1'b0) );
  NAND3_X1 pool_fsm_U25 ( .A1(pool_fsm_n8), .A2(pool_fsm_n6), .A3(
        pool_fsm_current_state_0_), .ZN(pool_fsm_n12) );
  NAND3_X1 pool_fsm_U24 ( .A1(pool_fsm_n9), .A2(pool_fsm_n8), .A3(
        pool_fsm_current_state_2_), .ZN(pool_fsm_n15) );
  NAND3_X1 pool_fsm_U23 ( .A1(pool_fsm_n12), .A2(pool_fsm_n15), .A3(
        pool_fsm_n5), .ZN(pool_fsm_N29) );
  NAND3_X1 pool_fsm_U22 ( .A1(pool_sel0), .A2(pool_fsm_n18), .A3(pool_tc), 
        .ZN(pool_fsm_n13) );
  NOR3_X2 pool_fsm_U15 ( .A1(pool_fsm_current_state_1_), .A2(
        pool_fsm_current_state_2_), .A3(pool_fsm_current_state_0_), .ZN(
        pool_fsm_N11) );
  NOR3_X2 pool_fsm_U14 ( .A1(pool_fsm_n9), .A2(pool_fsm_current_state_2_), 
        .A3(pool_fsm_n8), .ZN(pool_fsm_n16) );
  NAND2_X2 pool_fsm_U13 ( .A1(pool_fsm_n4), .A2(pool_fsm_n15), .ZN(
        pool_sync_clr) );
  NOR2_X2 pool_fsm_U12 ( .A1(pool_fsm_n16), .A2(pool_sync_clr), .ZN(
        pool_fsm_n11) );
  NAND2_X2 pool_fsm_U11 ( .A1(pool_fsm_n12), .A2(pool_fsm_n11), .ZN(
        pool_fsm_N28) );
  OR2_X2 pool_fsm_U10 ( .A1(start), .A2(pool_fsm_n4), .ZN(pool_fsm_N31) );
  NOR3_X2 pool_fsm_U9 ( .A1(pool_fsm_current_state_0_), .A2(
        pool_fsm_current_state_2_), .A3(pool_fsm_n8), .ZN(pool_fsm_n19) );
  NAND2_X2 pool_fsm_U8 ( .A1(pool_fsm_n12), .A2(pool_fsm_n2), .ZN(pool_en_cnt)
         );
  AND2_X2 pool_fsm_U7 ( .A1(pool_tc), .A2(done), .ZN(pool_fsm_n14) );
  OAI21_X2 pool_fsm_U6 ( .B1(pool_fsm_n14), .B2(pool_fsm_n2), .A(pool_fsm_n10), 
        .ZN(pool_fsm_next_state[0]) );
  NAND2_X2 pool_fsm_U5 ( .A1(pool_fsm_n12), .A2(pool_fsm_n13), .ZN(
        pool_fsm_next_state[1]) );
  OR2_X2 pool_fsm_U4 ( .A1(pool_sel0), .A2(pool_fsm_N29), .ZN(pool_rst_cnt_c)
         );
  DLH_X1 pool_fsm_rst_cnt_r_reg ( .G(pool_fsm_N28), .D(pool_fsm_N29), .Q(
        pool_rst_cnt_r) );
  DFFR_X1 pool_fsm_current_state_reg_2_ ( .D(pool_fsm_n16), .CK(
        pool_fsm_net424), .RN(pool_fsm_n17), .Q(pool_fsm_current_state_2_), 
        .QN(pool_fsm_n6) );
  DFFR_X1 pool_fsm_current_state_reg_1_ ( .D(pool_fsm_next_state[1]), .CK(
        pool_fsm_net424), .RN(pool_fsm_n17), .Q(pool_fsm_current_state_1_), 
        .QN(pool_fsm_n8) );
  DFFR_X1 pool_fsm_current_state_reg_0_ ( .D(pool_fsm_next_state[0]), .CK(
        pool_fsm_net424), .RN(pool_fsm_n17), .Q(pool_fsm_current_state_0_), 
        .QN(pool_fsm_n9) );
  INV_X2 pool_gate_clk_U36 ( .A(pool_gate_clk_pool_size_2_), .ZN(
        pool_gate_clk_n31) );
  INV_X2 pool_gate_clk_U35 ( .A(pool_rst_cnt_r), .ZN(pool_gate_clk_n30) );
  INV_X2 pool_gate_clk_U34 ( .A(pool_rst_cnt_c), .ZN(pool_gate_clk_n29) );
  INV_X2 pool_gate_clk_U33 ( .A(pool_gate_clk_n20), .ZN(pool_gate_clk_n28) );
  INV_X2 pool_gate_clk_U32 ( .A(pool_gate_clk_n15), .ZN(pool_gate_clk_n14) );
  MUX2_X1 pool_gate_clk_U28 ( .A(1'b0), .B(pool_gate_clk_N13), .S(
        pool_gate_clk_N0), .Z(pool_gate_clk_dec_out_2_) );
  MUX2_X1 pool_gate_clk_U27 ( .A(1'b0), .B(pool_gate_clk_n31), .S(
        pool_gate_clk_N0), .Z(pool_gate_clk_dec_out_1_) );
  MUX2_X1 pool_gate_clk_U26 ( .A(1'b0), .B(pool_gate_clk_N18), .S(
        pool_gate_clk_N0), .Z(pool_gate_clk_dec_out_0_) );
  INV_X4 pool_gate_clk_U25 ( .A(pool_ld_h), .ZN(pool_gate_clk_n7) );
  INV_X1 pool_gate_clk_U24 ( .A(pool_gate_clk_n7), .ZN(pool_gate_clk_n5) );
  INV_X1 pool_gate_clk_U16 ( .A(pool_ld_h), .ZN(pool_gate_clk_n4) );
  AND2_X1 pool_gate_clk_U5 ( .A1(pool_gate_clk_del_tc_r), .A2(pool_gate_clk_n4), .ZN(pool_gate_clk_n3) );
  AND2_X1 pool_gate_clk_U4 ( .A1(pool_gate_clk_del_0_tc), .A2(pool_gate_clk_n4), .ZN(pool_gate_clk_n2) );
  AND2_X1 pool_gate_clk_U3 ( .A1(pool_gate_clk_n4), .A2(pool_tc), .ZN(
        pool_gate_clk_n1) );
  DFF_X1 pool_gate_clk_del_0_tc_reg ( .D(pool_gate_clk_n1), .CK(clk), .Q(
        pool_gate_clk_del_0_tc) );
  DFF_X1 pool_gate_clk_del_1_tc_reg ( .D(pool_gate_clk_n2), .CK(clk), .Q(
        pool_gate_clk_del_1_tc) );
  DFF_X1 pool_gate_clk_del_tc_r_1_reg ( .D(pool_gate_clk_n3), .CK(clk), .Q(
        pool_gate_clk_del_tc_r_1) );
  NOR2_X2 pool_gate_clk_U23 ( .A1(pool_gate_clk_pool_size_2_), .A2(
        pool_gate_clk_pool_size_1_), .ZN(pool_gate_clk_N13) );
  NAND2_X2 pool_gate_clk_U22 ( .A1(pool_gate_clk_pool_size_1_), .A2(
        pool_gate_clk_pool_size_2_), .ZN(pool_gate_clk_N18) );
  NOR3_X2 pool_gate_clk_U21 ( .A1(pool_gate_clk_cnt_r_out_0_), .A2(pool_ld_h), 
        .A3(pool_gate_clk_cnt_r_out_1_), .ZN(pool_gate_clk_N45) );
  NOR3_X2 pool_gate_clk_U20 ( .A1(pool_gate_clk_n5), .A2(
        pool_gate_clk_del_1_tc), .A3(pool_gate_clk_n29), .ZN(pool_gate_clk_n20) );
  AOI221_X2 pool_gate_clk_U19 ( .B1(pool_gate_clk_n8), .B2(pool_gate_clk_n7), 
        .C1(pool_gate_clk_pool_size_3_), .C2(pool_gate_clk_n5), .A(
        pool_gate_clk_n29), .ZN(pool_gate_clk_n23) );
  OAI22_X2 pool_gate_clk_U18 ( .A1(pool_gate_clk_n8), .A2(pool_gate_clk_n28), 
        .B1(pool_gate_clk_n20), .B2(pool_gate_clk_n23), .ZN(pool_gate_clk_n27)
         );
  NOR2_X2 pool_gate_clk_U17 ( .A1(pool_gate_clk_cnt_c_out_0_), .A2(
        pool_gate_clk_cnt_c_out_1_), .ZN(pool_gate_clk_tc_c) );
  AOI221_X2 pool_gate_clk_U15 ( .B1(pool_gate_clk_tc_c), .B2(pool_gate_clk_n7), 
        .C1(pool_gate_clk_pool_size_4_), .C2(pool_gate_clk_n5), .A(
        pool_gate_clk_n29), .ZN(pool_gate_clk_n21) );
  AOI21_X2 pool_gate_clk_U14 ( .B1(pool_gate_clk_cnt_c_out_0_), .B2(
        pool_gate_clk_n7), .A(pool_gate_clk_n20), .ZN(pool_gate_clk_n22) );
  OAI22_X2 pool_gate_clk_U13 ( .A1(pool_gate_clk_n20), .A2(pool_gate_clk_n21), 
        .B1(pool_gate_clk_n22), .B2(pool_gate_clk_n6), .ZN(pool_gate_clk_n26)
         );
  AOI211_X2 pool_gate_clk_U12 ( .C1(pool_gate_clk_tc_c), .C2(pool_tc), .A(
        pool_gate_clk_n5), .B(pool_gate_clk_n30), .ZN(pool_gate_clk_n15) );
  AOI221_X2 pool_gate_clk_U11 ( .B1(pool_gate_clk_n10), .B2(pool_gate_clk_n7), 
        .C1(pool_gate_clk_pool_size_3_), .C2(pool_gate_clk_n5), .A(
        pool_gate_clk_n30), .ZN(pool_gate_clk_n19) );
  OAI22_X2 pool_gate_clk_U10 ( .A1(pool_gate_clk_n10), .A2(pool_gate_clk_n14), 
        .B1(pool_gate_clk_n15), .B2(pool_gate_clk_n19), .ZN(pool_gate_clk_n25)
         );
  NOR3_X2 pool_gate_clk_U9 ( .A1(pool_gate_clk_cnt_r_out_0_), .A2(
        pool_gate_clk_n5), .A3(pool_gate_clk_cnt_r_out_1_), .ZN(
        pool_gate_clk_n18) );
  AOI211_X2 pool_gate_clk_U8 ( .C1(pool_gate_clk_pool_size_4_), .C2(
        pool_gate_clk_n5), .A(pool_gate_clk_n30), .B(pool_gate_clk_n18), .ZN(
        pool_gate_clk_n16) );
  AOI21_X2 pool_gate_clk_U7 ( .B1(pool_gate_clk_cnt_r_out_0_), .B2(
        pool_gate_clk_n7), .A(pool_gate_clk_n15), .ZN(pool_gate_clk_n17) );
  OAI22_X2 pool_gate_clk_U6 ( .A1(pool_gate_clk_n15), .A2(pool_gate_clk_n16), 
        .B1(pool_gate_clk_n17), .B2(pool_gate_clk_n9), .ZN(pool_gate_clk_n24)
         );
  DFF_X1 pool_gate_clk_del_tc_r_reg ( .D(pool_gate_clk_N45), .CK(clk), .Q(
        pool_gate_clk_del_tc_r) );
  DFF_X1 pool_gate_clk_cnt_r_out_reg_1_ ( .D(pool_gate_clk_n24), .CK(clk), .Q(
        pool_gate_clk_cnt_r_out_1_), .QN(pool_gate_clk_n9) );
  DFF_X1 pool_gate_clk_cnt_r_out_reg_0_ ( .D(pool_gate_clk_n25), .CK(clk), .Q(
        pool_gate_clk_cnt_r_out_0_), .QN(pool_gate_clk_n10) );
  DFF_X1 pool_gate_clk_cnt_c_out_reg_1_ ( .D(pool_gate_clk_n26), .CK(clk), .Q(
        pool_gate_clk_cnt_c_out_1_), .QN(pool_gate_clk_n6) );
  DFF_X1 pool_gate_clk_cnt_c_out_reg_0_ ( .D(pool_gate_clk_n27), .CK(clk), .Q(
        pool_gate_clk_cnt_c_out_0_), .QN(pool_gate_clk_n8) );
  INV_X2 pool_gate_clk_mux_pool_U11 ( .A(pool_sel), .ZN(
        pool_gate_clk_mux_pool_n6) );
  INV_X2 pool_gate_clk_mux_pool_U10 ( .A(pool_gate_clk_mux_pool_n11), .ZN(
        pool_gate_clk_N0) );
  INV_X2 pool_gate_clk_mux_pool_U9 ( .A(pool_gate_clk_mux_pool_n10), .ZN(
        pool_gate_clk_pool_size_1_) );
  INV_X2 pool_gate_clk_mux_pool_U8 ( .A(pool_gate_clk_mux_pool_n9), .ZN(
        pool_gate_clk_pool_size_2_) );
  INV_X2 pool_gate_clk_mux_pool_U7 ( .A(pool_gate_clk_mux_pool_n8), .ZN(
        pool_gate_clk_pool_size_3_) );
  INV_X2 pool_gate_clk_mux_pool_U6 ( .A(pool_gate_clk_mux_pool_n7), .ZN(
        pool_gate_clk_pool_size_4_) );
  AOI22_X2 pool_gate_clk_mux_pool_U5 ( .A1(size_1[0]), .A2(
        pool_gate_clk_mux_pool_n6), .B1(size_2[0]), .B2(pool_sel), .ZN(
        pool_gate_clk_mux_pool_n11) );
  AOI22_X2 pool_gate_clk_mux_pool_U4 ( .A1(size_1[1]), .A2(
        pool_gate_clk_mux_pool_n6), .B1(size_2[1]), .B2(pool_sel), .ZN(
        pool_gate_clk_mux_pool_n10) );
  AOI22_X2 pool_gate_clk_mux_pool_U3 ( .A1(size_1[2]), .A2(
        pool_gate_clk_mux_pool_n6), .B1(size_2[2]), .B2(pool_sel), .ZN(
        pool_gate_clk_mux_pool_n9) );
  AOI22_X2 pool_gate_clk_mux_pool_U2 ( .A1(size_1[3]), .A2(
        pool_gate_clk_mux_pool_n6), .B1(size_2[3]), .B2(pool_sel), .ZN(
        pool_gate_clk_mux_pool_n8) );
  AOI22_X2 pool_gate_clk_mux_pool_U1 ( .A1(size_1[4]), .A2(
        pool_gate_clk_mux_pool_n6), .B1(pool_sel), .B2(size_2[4]), .ZN(
        pool_gate_clk_mux_pool_n7) );
  INV_X2 pool_gate_clk_mux_cmask_U5 ( .A(pool_gate_clk_tc_c), .ZN(
        pool_gate_clk_mux_cmask_n1) );
  MUX2_X1 pool_gate_clk_mux_cmask_U4 ( .A(1'b0), .B(1'b0), .S(
        pool_gate_clk_mux_cmask_n1), .Z(pool_ckg_cmask[3]) );
  MUX2_X1 pool_gate_clk_mux_cmask_U3 ( .A(pool_gate_clk_dec_out_2_), .B(1'b0), 
        .S(pool_gate_clk_mux_cmask_n1), .Z(pool_ckg_cmask[2]) );
  MUX2_X1 pool_gate_clk_mux_cmask_U2 ( .A(pool_gate_clk_dec_out_1_), .B(1'b0), 
        .S(pool_gate_clk_mux_cmask_n1), .Z(pool_ckg_cmask[1]) );
  MUX2_X1 pool_gate_clk_mux_cmask_U1 ( .A(pool_gate_clk_dec_out_0_), .B(1'b0), 
        .S(pool_gate_clk_mux_cmask_n1), .Z(pool_ckg_cmask[0]) );
  INV_X2 pool_gate_clk_mux_rmask_U5 ( .A(pool_gate_clk_del_tc_r_1), .ZN(
        pool_gate_clk_mux_rmask_n1) );
  MUX2_X1 pool_gate_clk_mux_rmask_U4 ( .A(1'b0), .B(1'b0), .S(
        pool_gate_clk_mux_rmask_n1), .Z(pool_ckg_rmask[3]) );
  MUX2_X1 pool_gate_clk_mux_rmask_U3 ( .A(pool_gate_clk_dec_out_2_), .B(1'b0), 
        .S(pool_gate_clk_mux_rmask_n1), .Z(pool_ckg_rmask[2]) );
  MUX2_X1 pool_gate_clk_mux_rmask_U2 ( .A(pool_gate_clk_dec_out_1_), .B(1'b0), 
        .S(pool_gate_clk_mux_rmask_n1), .Z(pool_ckg_rmask[1]) );
  MUX2_X1 pool_gate_clk_mux_rmask_U1 ( .A(pool_gate_clk_dec_out_0_), .B(1'b0), 
        .S(pool_gate_clk_mux_rmask_n1), .Z(pool_ckg_rmask[0]) );
endmodule

