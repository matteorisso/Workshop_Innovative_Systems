library verilog;
use verilog.vl_types.all;
entity tb_pool is
end tb_pool;
