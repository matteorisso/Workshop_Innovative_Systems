
module dp ( ck, rst, i_acth, i_actv, i_weight, arv_CKG, arv_KSI, arv_L0, 
        arv_L1, arv_L2, arv_L3, arv_L4, ctrl_en_npu, ctrl_ldh_v_n, 
        ctrl_en_hmode, ctrl_en_vmode, ctrl_wr_pipe, ctrl_en_p, ctrl_wr_mem, 
        s_tc_hmode, s_tc_vmode, s_tc_res, s_tc_L1, s_tc_L2, s_tc_L3, s_tc_L0, 
        s_tc_L4, i_weight_addr, i_data_ev_odd_n, i_data_even_addr, 
        i_data_odd_addr, o_data_ev_odd_n, o_data_even_addr, o_data_odd_addr, 
        o_data_wr, o_data_wrh_l_n, o_data, o_data_relu );
  input [15:0] i_acth;
  input [15:0] i_actv;
  input [1:0] i_weight;
  input [2:0] arv_CKG;
  input [2:0] arv_KSI;
  input [3:0] arv_L0;
  input [3:0] arv_L1;
  input [3:0] arv_L2;
  input [3:0] arv_L3;
  input [3:0] arv_L4;
  output [8:0] i_weight_addr;
  output [9:0] i_data_even_addr;
  output [9:0] i_data_odd_addr;
  output [9:0] o_data_even_addr;
  output [9:0] o_data_odd_addr;
  output [7:0] o_data;
  output [15:0] o_data_relu;
  input ck, rst, ctrl_en_npu, ctrl_ldh_v_n, ctrl_en_hmode, ctrl_en_vmode,
         ctrl_wr_pipe, ctrl_en_p, ctrl_wr_mem;
  output s_tc_hmode, s_tc_vmode, s_tc_res, s_tc_L1, s_tc_L2, s_tc_L3, s_tc_L0,
         s_tc_L4, i_data_ev_odd_n, o_data_ev_odd_n, o_data_wr, o_data_wrh_l_n;
  wire   ps_ctrl_en_npu, ps_ctrl_ldh_v_n, ps_ctrl_wr_pipe, ps_ctrl_en_p,
         int_en_hmode, int_en_vmode, int_en_L1_ptr, int_en_L2_ptr,
         int_en_L4_ptr, int_L3_ptr_1_, int_c_i_en_weight_addr, int_c_i_en_even,
         int_c_i_en_odd, ps_int_s_tc_res, ps_int_s_tc_L2, ps_int_s_tc_L3,
         int_c_o_en_offs_even, int_c_o_en_base_odd, int_c_o_en_offs_odd,
         net2764, n4, n7, n9, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, wrap_act_buffer_inst_n1, wrap_act_buffer_inst_net4585,
         wrap_act_buffer_inst_act_buffer_inst_n196,
         wrap_act_buffer_inst_act_buffer_inst_n195,
         wrap_act_buffer_inst_act_buffer_inst_n194,
         wrap_act_buffer_inst_act_buffer_inst_n193,
         wrap_act_buffer_inst_act_buffer_inst_n192,
         wrap_act_buffer_inst_act_buffer_inst_n191,
         wrap_act_buffer_inst_act_buffer_inst_n190,
         wrap_act_buffer_inst_act_buffer_inst_n189,
         wrap_act_buffer_inst_act_buffer_inst_n188,
         wrap_act_buffer_inst_act_buffer_inst_n187,
         wrap_act_buffer_inst_act_buffer_inst_n186,
         wrap_act_buffer_inst_act_buffer_inst_n185,
         wrap_act_buffer_inst_act_buffer_inst_n184,
         wrap_act_buffer_inst_act_buffer_inst_n183,
         wrap_act_buffer_inst_act_buffer_inst_n182,
         wrap_act_buffer_inst_act_buffer_inst_n181,
         wrap_act_buffer_inst_act_buffer_inst_n180,
         wrap_act_buffer_inst_act_buffer_inst_n179,
         wrap_act_buffer_inst_act_buffer_inst_n178,
         wrap_act_buffer_inst_act_buffer_inst_n177,
         wrap_act_buffer_inst_act_buffer_inst_n176,
         wrap_act_buffer_inst_act_buffer_inst_n175,
         wrap_act_buffer_inst_act_buffer_inst_n174,
         wrap_act_buffer_inst_act_buffer_inst_n173,
         wrap_act_buffer_inst_act_buffer_inst_n172,
         wrap_act_buffer_inst_act_buffer_inst_n171,
         wrap_act_buffer_inst_act_buffer_inst_n170,
         wrap_act_buffer_inst_act_buffer_inst_n169,
         wrap_act_buffer_inst_act_buffer_inst_n168,
         wrap_act_buffer_inst_act_buffer_inst_n167,
         wrap_act_buffer_inst_act_buffer_inst_n166,
         wrap_act_buffer_inst_act_buffer_inst_n165,
         wrap_act_buffer_inst_act_buffer_inst_n164,
         wrap_act_buffer_inst_act_buffer_inst_n163,
         wrap_act_buffer_inst_act_buffer_inst_n162,
         wrap_act_buffer_inst_act_buffer_inst_n161,
         wrap_act_buffer_inst_act_buffer_inst_n160,
         wrap_act_buffer_inst_act_buffer_inst_n159,
         wrap_act_buffer_inst_act_buffer_inst_n9,
         wrap_act_buffer_inst_act_buffer_inst_n8,
         wrap_act_buffer_inst_act_buffer_inst_n7,
         wrap_act_buffer_inst_act_buffer_inst_n6,
         wrap_act_buffer_inst_act_buffer_inst_n5,
         wrap_act_buffer_inst_act_buffer_inst_n4,
         wrap_act_buffer_inst_act_buffer_inst_n3,
         wrap_act_buffer_inst_act_buffer_inst_n2,
         wrap_act_buffer_inst_act_buffer_inst_n1,
         wrap_act_buffer_inst_act_buffer_inst_n158,
         wrap_act_buffer_inst_act_buffer_inst_n157,
         wrap_act_buffer_inst_act_buffer_inst_n156,
         wrap_act_buffer_inst_act_buffer_inst_n155,
         wrap_act_buffer_inst_act_buffer_inst_n154,
         wrap_act_buffer_inst_act_buffer_inst_n153,
         wrap_act_buffer_inst_act_buffer_inst_n152,
         wrap_act_buffer_inst_act_buffer_inst_n151,
         wrap_act_buffer_inst_act_buffer_inst_n150,
         wrap_act_buffer_inst_act_buffer_inst_n149,
         wrap_act_buffer_inst_act_buffer_inst_n148,
         wrap_act_buffer_inst_act_buffer_inst_n147,
         wrap_act_buffer_inst_act_buffer_inst_n146,
         wrap_act_buffer_inst_act_buffer_inst_n145,
         wrap_act_buffer_inst_act_buffer_inst_n144,
         wrap_act_buffer_inst_act_buffer_inst_n143,
         wrap_act_buffer_inst_act_buffer_inst_n142,
         wrap_act_buffer_inst_act_buffer_inst_n141,
         wrap_act_buffer_inst_act_buffer_inst_n140,
         wrap_act_buffer_inst_act_buffer_inst_n139,
         wrap_act_buffer_inst_act_buffer_inst_n138,
         wrap_act_buffer_inst_act_buffer_inst_n137,
         wrap_act_buffer_inst_act_buffer_inst_n136,
         wrap_act_buffer_inst_act_buffer_inst_n135,
         wrap_act_buffer_inst_act_buffer_inst_n134,
         wrap_act_buffer_inst_act_buffer_inst_n133,
         wrap_act_buffer_inst_act_buffer_inst_n132,
         wrap_act_buffer_inst_act_buffer_inst_n131,
         wrap_act_buffer_inst_act_buffer_inst_n130,
         wrap_act_buffer_inst_act_buffer_inst_n129,
         wrap_act_buffer_inst_act_buffer_inst_n128,
         wrap_act_buffer_inst_act_buffer_inst_n127,
         wrap_act_buffer_inst_act_buffer_inst_n126,
         wrap_act_buffer_inst_act_buffer_inst_n125,
         wrap_act_buffer_inst_act_buffer_inst_n124,
         wrap_act_buffer_inst_act_buffer_inst_n123,
         wrap_act_buffer_inst_act_buffer_inst_n122,
         wrap_act_buffer_inst_act_buffer_inst_n121,
         wrap_act_buffer_inst_act_buffer_inst_n120,
         wrap_act_buffer_inst_act_buffer_inst_n119,
         wrap_act_buffer_inst_act_buffer_inst_n118,
         wrap_act_buffer_inst_act_buffer_inst_n117,
         wrap_act_buffer_inst_act_buffer_inst_n116,
         wrap_act_buffer_inst_act_buffer_inst_n115,
         wrap_act_buffer_inst_act_buffer_inst_n114,
         wrap_act_buffer_inst_act_buffer_inst_n113,
         wrap_act_buffer_inst_act_buffer_inst_n112,
         wrap_act_buffer_inst_act_buffer_inst_n111,
         wrap_act_buffer_inst_act_buffer_inst_n110,
         wrap_act_buffer_inst_act_buffer_inst_n109,
         wrap_act_buffer_inst_act_buffer_inst_n108,
         wrap_act_buffer_inst_act_buffer_inst_n107,
         wrap_act_buffer_inst_act_buffer_inst_n106,
         wrap_act_buffer_inst_act_buffer_inst_n105,
         wrap_act_buffer_inst_act_buffer_inst_n104,
         wrap_act_buffer_inst_act_buffer_inst_n103,
         wrap_act_buffer_inst_act_buffer_inst_n102,
         wrap_act_buffer_inst_act_buffer_inst_n101,
         wrap_act_buffer_inst_act_buffer_inst_n100,
         wrap_act_buffer_inst_act_buffer_inst_n99,
         wrap_act_buffer_inst_act_buffer_inst_n98,
         wrap_act_buffer_inst_act_buffer_inst_n97,
         wrap_act_buffer_inst_act_buffer_inst_n96,
         wrap_act_buffer_inst_act_buffer_inst_n95,
         wrap_act_buffer_inst_act_buffer_inst_n94,
         wrap_act_buffer_inst_act_buffer_inst_n93,
         wrap_act_buffer_inst_act_buffer_inst_n92,
         wrap_act_buffer_inst_act_buffer_inst_n91,
         wrap_act_buffer_inst_act_buffer_inst_n90,
         wrap_act_buffer_inst_act_buffer_inst_n89,
         wrap_act_buffer_inst_act_buffer_inst_n88,
         wrap_act_buffer_inst_act_buffer_inst_n87,
         wrap_act_buffer_inst_act_buffer_inst_n86,
         wrap_act_buffer_inst_act_buffer_inst_n85,
         wrap_act_buffer_inst_act_buffer_inst_n84,
         wrap_act_buffer_inst_act_buffer_inst_n83,
         wrap_act_buffer_inst_act_buffer_inst_n82,
         wrap_act_buffer_inst_act_buffer_inst_n81,
         wrap_act_buffer_inst_act_buffer_inst_n80,
         wrap_act_buffer_inst_act_buffer_inst_n79,
         wrap_act_buffer_inst_act_buffer_inst_n78,
         wrap_act_buffer_inst_act_buffer_inst_n77,
         wrap_act_buffer_inst_act_buffer_inst_n76,
         wrap_act_buffer_inst_act_buffer_inst_n75,
         wrap_act_buffer_inst_act_buffer_inst_n74,
         wrap_act_buffer_inst_act_buffer_inst_n73,
         wrap_act_buffer_inst_act_buffer_inst_n72,
         wrap_act_buffer_inst_act_buffer_inst_n71,
         wrap_act_buffer_inst_act_buffer_inst_n70,
         wrap_act_buffer_inst_act_buffer_inst_n69,
         wrap_act_buffer_inst_act_buffer_inst_n68,
         wrap_act_buffer_inst_act_buffer_inst_n67,
         wrap_act_buffer_inst_act_buffer_inst_n66,
         wrap_act_buffer_inst_act_buffer_inst_n65,
         wrap_act_buffer_inst_act_buffer_inst_n64,
         wrap_act_buffer_inst_act_buffer_inst_n63,
         wrap_act_buffer_inst_act_buffer_inst_n62,
         wrap_act_buffer_inst_act_buffer_inst_n61,
         wrap_act_buffer_inst_act_buffer_inst_n60,
         wrap_act_buffer_inst_act_buffer_inst_n59,
         wrap_act_buffer_inst_act_buffer_inst_n58,
         wrap_act_buffer_inst_act_buffer_inst_n57,
         wrap_act_buffer_inst_act_buffer_inst_n56,
         wrap_act_buffer_inst_act_buffer_inst_n55,
         wrap_act_buffer_inst_act_buffer_inst_n54,
         wrap_act_buffer_inst_act_buffer_inst_n53,
         wrap_act_buffer_inst_act_buffer_inst_n52,
         wrap_act_buffer_inst_act_buffer_inst_n51,
         wrap_act_buffer_inst_act_buffer_inst_n50,
         wrap_act_buffer_inst_act_buffer_inst_n49,
         wrap_act_buffer_inst_act_buffer_inst_n48,
         wrap_act_buffer_inst_act_buffer_inst_n47,
         wrap_act_buffer_inst_act_buffer_inst_n46,
         wrap_act_buffer_inst_act_buffer_inst_n45,
         wrap_act_buffer_inst_act_buffer_inst_n44,
         wrap_act_buffer_inst_act_buffer_inst_n43,
         wrap_act_buffer_inst_act_buffer_inst_n42,
         wrap_act_buffer_inst_act_buffer_inst_n41,
         wrap_act_buffer_inst_act_buffer_inst_n40,
         wrap_act_buffer_inst_act_buffer_inst_n39,
         wrap_act_buffer_inst_act_buffer_inst_n38,
         wrap_act_buffer_inst_act_buffer_inst_n37,
         wrap_act_buffer_inst_act_buffer_inst_n36,
         wrap_act_buffer_inst_act_buffer_inst_n35,
         wrap_act_buffer_inst_act_buffer_inst_n34,
         wrap_act_buffer_inst_act_buffer_inst_n33,
         wrap_act_buffer_inst_act_buffer_inst_n32,
         wrap_act_buffer_inst_act_buffer_inst_n31,
         wrap_act_buffer_inst_act_buffer_inst_n30,
         wrap_act_buffer_inst_act_buffer_inst_n29,
         wrap_act_buffer_inst_act_buffer_inst_n28,
         wrap_act_buffer_inst_act_buffer_inst_n27,
         wrap_act_buffer_inst_act_buffer_inst_n26,
         wrap_act_buffer_inst_act_buffer_inst_n25,
         wrap_act_buffer_inst_act_buffer_inst_n24,
         wrap_act_buffer_inst_act_buffer_inst_n23,
         wrap_act_buffer_inst_act_buffer_inst_n22,
         wrap_act_buffer_inst_act_buffer_inst_n21,
         wrap_act_buffer_inst_act_buffer_inst_n20,
         wrap_act_buffer_inst_act_buffer_inst_n19,
         wrap_act_buffer_inst_act_buffer_inst_n18,
         wrap_act_buffer_inst_act_buffer_inst_n17,
         wrap_act_buffer_inst_act_buffer_inst_n16,
         wrap_act_buffer_inst_act_buffer_inst_n15,
         wrap_act_buffer_inst_act_buffer_inst_n14,
         wrap_act_buffer_inst_act_buffer_inst_n13,
         wrap_act_buffer_inst_act_buffer_inst_n12,
         wrap_act_buffer_inst_act_buffer_inst_n11,
         wrap_act_buffer_inst_act_buffer_inst_n10,
         wrap_act_buffer_inst_act_buffer_inst_net4839,
         wrap_act_buffer_inst_act_buffer_inst_net4834,
         wrap_act_buffer_inst_act_buffer_inst_net4829,
         wrap_act_buffer_inst_act_buffer_inst_net4824,
         wrap_act_buffer_inst_act_buffer_inst_net4819,
         wrap_act_buffer_inst_act_buffer_inst_net4814,
         wrap_act_buffer_inst_act_buffer_inst_net4809,
         wrap_act_buffer_inst_act_buffer_inst_net4804,
         wrap_act_buffer_inst_act_buffer_inst_net4799,
         wrap_act_buffer_inst_act_buffer_inst_net4794,
         wrap_act_buffer_inst_act_buffer_inst_net4789,
         wrap_act_buffer_inst_act_buffer_inst_net4784,
         wrap_act_buffer_inst_act_buffer_inst_net4779,
         wrap_act_buffer_inst_act_buffer_inst_net4774,
         wrap_act_buffer_inst_act_buffer_inst_net4769,
         wrap_act_buffer_inst_act_buffer_inst_net4764,
         wrap_act_buffer_inst_act_buffer_inst_net4759,
         wrap_act_buffer_inst_act_buffer_inst_net4754,
         wrap_act_buffer_inst_act_buffer_inst_net4749,
         wrap_act_buffer_inst_act_buffer_inst_net4744,
         wrap_act_buffer_inst_act_buffer_inst_net4739,
         wrap_act_buffer_inst_act_buffer_inst_net4734,
         wrap_act_buffer_inst_act_buffer_inst_net4729,
         wrap_act_buffer_inst_act_buffer_inst_net4724,
         wrap_act_buffer_inst_act_buffer_inst_net4719,
         wrap_act_buffer_inst_act_buffer_inst_net4714,
         wrap_act_buffer_inst_act_buffer_inst_net4709,
         wrap_act_buffer_inst_act_buffer_inst_net4704,
         wrap_act_buffer_inst_act_buffer_inst_net4699,
         wrap_act_buffer_inst_act_buffer_inst_net4694,
         wrap_act_buffer_inst_act_buffer_inst_net4689,
         wrap_act_buffer_inst_act_buffer_inst_net4684,
         wrap_act_buffer_inst_act_buffer_inst_net4679,
         wrap_act_buffer_inst_act_buffer_inst_net4674,
         wrap_act_buffer_inst_act_buffer_inst_net4669,
         wrap_act_buffer_inst_act_buffer_inst_net4664,
         wrap_act_buffer_inst_act_buffer_inst_net4659,
         wrap_act_buffer_inst_act_buffer_inst_net4654,
         wrap_act_buffer_inst_act_buffer_inst_net4649,
         wrap_act_buffer_inst_act_buffer_inst_net4644,
         wrap_act_buffer_inst_act_buffer_inst_net4639,
         wrap_act_buffer_inst_act_buffer_inst_net4634,
         wrap_act_buffer_inst_act_buffer_inst_net4629,
         wrap_act_buffer_inst_act_buffer_inst_net4624,
         wrap_act_buffer_inst_act_buffer_inst_net4619,
         wrap_act_buffer_inst_act_buffer_inst_net4614,
         wrap_act_buffer_inst_act_buffer_inst_net4609,
         wrap_act_buffer_inst_act_buffer_inst_net4603,
         wrap_act_buffer_inst_act_buffer_inst_N162,
         wrap_act_buffer_inst_act_buffer_inst_N161,
         wrap_act_buffer_inst_act_buffer_inst_N160,
         wrap_act_buffer_inst_act_buffer_inst_N159,
         wrap_act_buffer_inst_act_buffer_inst_N158,
         wrap_act_buffer_inst_act_buffer_inst_N157,
         wrap_act_buffer_inst_act_buffer_inst_N156,
         wrap_act_buffer_inst_act_buffer_inst_N155,
         wrap_act_buffer_inst_act_buffer_inst_N154,
         wrap_act_buffer_inst_act_buffer_inst_N153,
         wrap_act_buffer_inst_act_buffer_inst_N152,
         wrap_act_buffer_inst_act_buffer_inst_N151,
         wrap_act_buffer_inst_act_buffer_inst_N150,
         wrap_act_buffer_inst_act_buffer_inst_N149,
         wrap_act_buffer_inst_act_buffer_inst_N148,
         wrap_act_buffer_inst_act_buffer_inst_N147,
         wrap_act_buffer_inst_act_buffer_inst_N146,
         wrap_act_buffer_inst_act_buffer_inst_N145,
         wrap_act_buffer_inst_act_buffer_inst_N144,
         wrap_act_buffer_inst_act_buffer_inst_N143,
         wrap_act_buffer_inst_act_buffer_inst_N142,
         wrap_act_buffer_inst_act_buffer_inst_N141,
         wrap_act_buffer_inst_act_buffer_inst_N140,
         wrap_act_buffer_inst_act_buffer_inst_N139,
         wrap_act_buffer_inst_act_buffer_inst_N138,
         wrap_act_buffer_inst_act_buffer_inst_N137,
         wrap_act_buffer_inst_act_buffer_inst_N136,
         wrap_act_buffer_inst_act_buffer_inst_N135,
         wrap_act_buffer_inst_act_buffer_inst_N134,
         wrap_act_buffer_inst_act_buffer_inst_N133,
         wrap_act_buffer_inst_act_buffer_inst_N132,
         wrap_act_buffer_inst_act_buffer_inst_N131,
         wrap_act_buffer_inst_act_buffer_inst_N130,
         wrap_act_buffer_inst_act_buffer_inst_N129,
         wrap_act_buffer_inst_act_buffer_inst_N128,
         wrap_act_buffer_inst_act_buffer_inst_N127,
         wrap_act_buffer_inst_act_buffer_inst_N126,
         wrap_act_buffer_inst_act_buffer_inst_N125,
         wrap_act_buffer_inst_act_buffer_inst_N124,
         wrap_act_buffer_inst_act_buffer_inst_N123,
         wrap_act_buffer_inst_act_buffer_inst_N122,
         wrap_act_buffer_inst_act_buffer_inst_N121,
         wrap_act_buffer_inst_act_buffer_inst_N120,
         wrap_act_buffer_inst_act_buffer_inst_N119,
         wrap_act_buffer_inst_act_buffer_inst_N118,
         wrap_act_buffer_inst_act_buffer_inst_N117,
         wrap_act_buffer_inst_act_buffer_inst_N116,
         wrap_act_buffer_inst_act_buffer_inst_N115,
         wrap_act_buffer_inst_act_if_inst_n312,
         wrap_act_buffer_inst_act_if_inst_n311,
         wrap_act_buffer_inst_act_if_inst_n310,
         wrap_act_buffer_inst_act_if_inst_n309,
         wrap_act_buffer_inst_act_if_inst_n308,
         wrap_act_buffer_inst_act_if_inst_n307,
         wrap_act_buffer_inst_act_if_inst_n306,
         wrap_act_buffer_inst_act_if_inst_n305,
         wrap_act_buffer_inst_act_if_inst_n304,
         wrap_act_buffer_inst_act_if_inst_n303,
         wrap_act_buffer_inst_act_if_inst_n302,
         wrap_act_buffer_inst_act_if_inst_n301,
         wrap_act_buffer_inst_act_if_inst_n300,
         wrap_act_buffer_inst_act_if_inst_n299,
         wrap_act_buffer_inst_act_if_inst_n298,
         wrap_act_buffer_inst_act_if_inst_n297,
         wrap_act_buffer_inst_act_if_inst_n296,
         wrap_act_buffer_inst_act_if_inst_n295,
         wrap_act_buffer_inst_act_if_inst_n294,
         wrap_act_buffer_inst_act_if_inst_n293,
         wrap_act_buffer_inst_act_if_inst_n292,
         wrap_act_buffer_inst_act_if_inst_n291,
         wrap_act_buffer_inst_act_if_inst_n290,
         wrap_act_buffer_inst_act_if_inst_n289,
         wrap_act_buffer_inst_act_if_inst_n288,
         wrap_act_buffer_inst_act_if_inst_n287,
         wrap_act_buffer_inst_act_if_inst_n286,
         wrap_act_buffer_inst_act_if_inst_n285,
         wrap_act_buffer_inst_act_if_inst_n284,
         wrap_act_buffer_inst_act_if_inst_n283,
         wrap_act_buffer_inst_act_if_inst_n282,
         wrap_act_buffer_inst_act_if_inst_n281,
         wrap_act_buffer_inst_act_if_inst_n280,
         wrap_act_buffer_inst_act_if_inst_n279,
         wrap_act_buffer_inst_act_if_inst_n278,
         wrap_act_buffer_inst_act_if_inst_n277,
         wrap_act_buffer_inst_act_if_inst_n276,
         wrap_act_buffer_inst_act_if_inst_n275,
         wrap_act_buffer_inst_act_if_inst_n274,
         wrap_act_buffer_inst_act_if_inst_n273,
         wrap_act_buffer_inst_act_if_inst_n272,
         wrap_act_buffer_inst_act_if_inst_n271,
         wrap_act_buffer_inst_act_if_inst_n270,
         wrap_act_buffer_inst_act_if_inst_n269,
         wrap_act_buffer_inst_act_if_inst_n268,
         wrap_act_buffer_inst_act_if_inst_n267,
         wrap_act_buffer_inst_act_if_inst_n266,
         wrap_act_buffer_inst_act_if_inst_n265,
         wrap_act_buffer_inst_act_if_inst_n264,
         wrap_act_buffer_inst_act_if_inst_n263,
         wrap_act_buffer_inst_act_if_inst_n262,
         wrap_act_buffer_inst_act_if_inst_n261,
         wrap_act_buffer_inst_act_if_inst_n260,
         wrap_act_buffer_inst_act_if_inst_n259,
         wrap_act_buffer_inst_act_if_inst_n258,
         wrap_act_buffer_inst_act_if_inst_n257,
         wrap_act_buffer_inst_act_if_inst_n256,
         wrap_act_buffer_inst_act_if_inst_n255,
         wrap_act_buffer_inst_act_if_inst_n254,
         wrap_act_buffer_inst_act_if_inst_n253,
         wrap_act_buffer_inst_act_if_inst_n252,
         wrap_act_buffer_inst_act_if_inst_n251,
         wrap_act_buffer_inst_act_if_inst_n250,
         wrap_act_buffer_inst_act_if_inst_n249,
         wrap_act_buffer_inst_act_if_inst_n248,
         wrap_act_buffer_inst_act_if_inst_n247,
         wrap_act_buffer_inst_act_if_inst_n246,
         wrap_act_buffer_inst_act_if_inst_n245,
         wrap_act_buffer_inst_act_if_inst_n244,
         wrap_act_buffer_inst_act_if_inst_n243,
         wrap_act_buffer_inst_act_if_inst_n242,
         wrap_act_buffer_inst_act_if_inst_n241,
         wrap_act_buffer_inst_act_if_inst_n240,
         wrap_act_buffer_inst_act_if_inst_n239,
         wrap_act_buffer_inst_act_if_inst_n238,
         wrap_act_buffer_inst_act_if_inst_n237,
         wrap_act_buffer_inst_act_if_inst_n236,
         wrap_act_buffer_inst_act_if_inst_n235,
         wrap_act_buffer_inst_act_if_inst_n234,
         wrap_act_buffer_inst_act_if_inst_n233,
         wrap_act_buffer_inst_act_if_inst_n232,
         wrap_act_buffer_inst_act_if_inst_n231,
         wrap_act_buffer_inst_act_if_inst_n230,
         wrap_act_buffer_inst_act_if_inst_n229,
         wrap_act_buffer_inst_act_if_inst_n228,
         wrap_act_buffer_inst_act_if_inst_n227,
         wrap_act_buffer_inst_act_if_inst_n226,
         wrap_act_buffer_inst_act_if_inst_n225,
         wrap_act_buffer_inst_act_if_inst_n224,
         wrap_act_buffer_inst_act_if_inst_n223,
         wrap_act_buffer_inst_act_if_inst_n222,
         wrap_act_buffer_inst_act_if_inst_n221,
         wrap_act_buffer_inst_act_if_inst_n220,
         wrap_act_buffer_inst_act_if_inst_n219,
         wrap_act_buffer_inst_act_if_inst_n218,
         wrap_act_buffer_inst_act_if_inst_n217,
         wrap_act_buffer_inst_act_if_inst_n216,
         wrap_act_buffer_inst_act_if_inst_n215,
         wrap_act_buffer_inst_act_if_inst_n214,
         wrap_act_buffer_inst_act_if_inst_n213,
         wrap_act_buffer_inst_act_if_inst_n212,
         wrap_act_buffer_inst_act_if_inst_n211,
         wrap_act_buffer_inst_act_if_inst_n210,
         wrap_act_buffer_inst_act_if_inst_n209,
         wrap_act_buffer_inst_act_if_inst_n208,
         wrap_act_buffer_inst_act_if_inst_n207,
         wrap_act_buffer_inst_act_if_inst_n206,
         wrap_act_buffer_inst_act_if_inst_n205,
         wrap_act_buffer_inst_act_if_inst_n204,
         wrap_act_buffer_inst_act_if_inst_n203,
         wrap_act_buffer_inst_act_if_inst_n202,
         wrap_act_buffer_inst_act_if_inst_n201,
         wrap_act_buffer_inst_act_if_inst_n200,
         wrap_act_buffer_inst_act_if_inst_n199,
         wrap_act_buffer_inst_act_if_inst_n198,
         wrap_act_buffer_inst_act_if_inst_n197,
         wrap_act_buffer_inst_act_if_inst_n196,
         wrap_act_buffer_inst_act_if_inst_n195,
         wrap_act_buffer_inst_act_if_inst_n194,
         wrap_act_buffer_inst_act_if_inst_n193,
         wrap_act_buffer_inst_act_if_inst_n192,
         wrap_act_buffer_inst_act_if_inst_n191,
         wrap_act_buffer_inst_act_if_inst_n190,
         wrap_act_buffer_inst_act_if_inst_n189,
         wrap_act_buffer_inst_act_if_inst_n188,
         wrap_act_buffer_inst_act_if_inst_n187,
         wrap_act_buffer_inst_act_if_inst_n186,
         wrap_act_buffer_inst_act_if_inst_n185,
         wrap_act_buffer_inst_act_if_inst_n184,
         wrap_act_buffer_inst_act_if_inst_n183,
         wrap_act_buffer_inst_act_if_inst_n182,
         wrap_act_buffer_inst_act_if_inst_n181,
         wrap_act_buffer_inst_act_if_inst_n180,
         wrap_act_buffer_inst_act_if_inst_n179,
         wrap_act_buffer_inst_act_if_inst_n178,
         wrap_act_buffer_inst_act_if_inst_n177,
         wrap_act_buffer_inst_act_if_inst_n176,
         wrap_act_buffer_inst_act_if_inst_n175,
         wrap_act_buffer_inst_act_if_inst_n174,
         wrap_act_buffer_inst_act_if_inst_n173,
         wrap_act_buffer_inst_act_if_inst_n172,
         wrap_act_buffer_inst_act_if_inst_n171,
         wrap_act_buffer_inst_act_if_inst_n170,
         wrap_act_buffer_inst_act_if_inst_n169,
         wrap_act_buffer_inst_act_if_inst_n168,
         wrap_act_buffer_inst_act_if_inst_n167,
         wrap_act_buffer_inst_act_if_inst_n166,
         wrap_act_buffer_inst_act_if_inst_n165,
         wrap_act_buffer_inst_act_if_inst_n164,
         wrap_act_buffer_inst_act_if_inst_n163,
         wrap_act_buffer_inst_act_if_inst_n162,
         wrap_act_buffer_inst_act_if_inst_n161,
         wrap_act_buffer_inst_act_if_inst_n160,
         wrap_act_buffer_inst_act_if_inst_n159,
         wrap_act_buffer_inst_act_if_inst_n158,
         wrap_act_buffer_inst_act_if_inst_n157,
         wrap_act_buffer_inst_act_if_inst_n156,
         wrap_act_buffer_inst_act_if_inst_n155,
         wrap_act_buffer_inst_act_if_inst_n154,
         wrap_act_buffer_inst_act_if_inst_n153,
         wrap_act_buffer_inst_act_if_inst_n152,
         wrap_act_buffer_inst_act_if_inst_n151,
         wrap_act_buffer_inst_act_if_inst_n150,
         wrap_act_buffer_inst_act_if_inst_n149,
         wrap_act_buffer_inst_act_if_inst_n148,
         wrap_act_buffer_inst_act_if_inst_n147,
         wrap_act_buffer_inst_act_if_inst_n146,
         wrap_act_buffer_inst_act_if_inst_n145,
         wrap_act_buffer_inst_act_if_inst_n144,
         wrap_act_buffer_inst_act_if_inst_n143,
         wrap_act_buffer_inst_act_if_inst_n142,
         wrap_act_buffer_inst_act_if_inst_n141,
         wrap_act_buffer_inst_act_if_inst_n140,
         wrap_act_buffer_inst_act_if_inst_n139,
         wrap_act_buffer_inst_act_if_inst_n138,
         wrap_act_buffer_inst_act_if_inst_n137,
         wrap_act_buffer_inst_act_if_inst_n136,
         wrap_act_buffer_inst_act_if_inst_n135,
         wrap_act_buffer_inst_act_if_inst_n134,
         wrap_act_buffer_inst_act_if_inst_n133,
         wrap_act_buffer_inst_act_if_inst_n132,
         wrap_act_buffer_inst_act_if_inst_n131,
         wrap_act_buffer_inst_act_if_inst_n130,
         wrap_act_buffer_inst_act_if_inst_n129,
         wrap_act_buffer_inst_act_if_inst_n128,
         wrap_act_buffer_inst_act_if_inst_n127,
         wrap_act_buffer_inst_act_if_inst_n126,
         wrap_act_buffer_inst_act_if_inst_n125,
         wrap_act_buffer_inst_act_if_inst_n124,
         wrap_act_buffer_inst_act_if_inst_n123,
         wrap_act_buffer_inst_act_if_inst_n122,
         wrap_act_buffer_inst_act_if_inst_n121,
         wrap_act_buffer_inst_act_if_inst_n120,
         wrap_act_buffer_inst_act_if_inst_n119,
         wrap_act_buffer_inst_act_if_inst_n118,
         wrap_act_buffer_inst_act_if_inst_n117,
         wrap_act_buffer_inst_act_if_inst_n116,
         wrap_act_buffer_inst_act_if_inst_n115,
         wrap_act_buffer_inst_act_if_inst_n114,
         wrap_act_buffer_inst_act_if_inst_n113,
         wrap_act_buffer_inst_act_if_inst_n112,
         wrap_act_buffer_inst_act_if_inst_n111,
         wrap_act_buffer_inst_act_if_inst_n110,
         wrap_act_buffer_inst_act_if_inst_n109,
         wrap_act_buffer_inst_act_if_inst_n108,
         wrap_act_buffer_inst_act_if_inst_n107,
         wrap_act_buffer_inst_act_if_inst_n106,
         wrap_act_buffer_inst_act_if_inst_n105,
         wrap_act_buffer_inst_act_if_inst_n104,
         wrap_act_buffer_inst_act_if_inst_n103,
         wrap_act_buffer_inst_act_if_inst_n102,
         wrap_act_buffer_inst_act_if_inst_n101,
         wrap_act_buffer_inst_act_if_inst_n100,
         wrap_act_buffer_inst_act_if_inst_n99,
         wrap_act_buffer_inst_act_if_inst_n98,
         wrap_act_buffer_inst_act_if_inst_n97,
         wrap_act_buffer_inst_act_if_inst_n96,
         wrap_act_buffer_inst_act_if_inst_n95,
         wrap_act_buffer_inst_act_if_inst_n94,
         wrap_act_buffer_inst_act_if_inst_n93,
         wrap_act_buffer_inst_act_if_inst_n92,
         wrap_act_buffer_inst_act_if_inst_n91,
         wrap_act_buffer_inst_act_if_inst_n90,
         wrap_act_buffer_inst_act_if_inst_n89,
         wrap_act_buffer_inst_act_if_inst_n88,
         wrap_act_buffer_inst_act_if_inst_n87,
         wrap_act_buffer_inst_act_if_inst_n86,
         wrap_act_buffer_inst_act_if_inst_n85,
         wrap_act_buffer_inst_act_if_inst_n84,
         wrap_act_buffer_inst_act_if_inst_n83,
         wrap_act_buffer_inst_act_if_inst_n82,
         wrap_act_buffer_inst_act_if_inst_n81,
         wrap_act_buffer_inst_act_if_inst_n80,
         wrap_act_buffer_inst_act_if_inst_n79,
         wrap_act_buffer_inst_act_if_inst_n78,
         wrap_act_buffer_inst_act_if_inst_n77,
         wrap_act_buffer_inst_act_if_inst_n76,
         wrap_act_buffer_inst_act_if_inst_n75,
         wrap_act_buffer_inst_act_if_inst_n74,
         wrap_act_buffer_inst_act_if_inst_n73,
         wrap_act_buffer_inst_act_if_inst_n72,
         wrap_act_buffer_inst_act_if_inst_n71,
         wrap_act_buffer_inst_act_if_inst_n70,
         wrap_act_buffer_inst_act_if_inst_n69,
         wrap_act_buffer_inst_act_if_inst_n68,
         wrap_act_buffer_inst_act_if_inst_n67,
         wrap_act_buffer_inst_act_if_inst_n66,
         wrap_act_buffer_inst_act_if_inst_n65,
         wrap_act_buffer_inst_act_if_inst_n64,
         wrap_act_buffer_inst_act_if_inst_n63,
         wrap_act_buffer_inst_act_if_inst_n62,
         wrap_act_buffer_inst_act_if_inst_n61,
         wrap_act_buffer_inst_act_if_inst_n60,
         wrap_act_buffer_inst_act_if_inst_n59,
         wrap_act_buffer_inst_act_if_inst_n58,
         wrap_act_buffer_inst_act_if_inst_n57,
         wrap_act_buffer_inst_act_if_inst_n56,
         wrap_act_buffer_inst_act_if_inst_n55,
         wrap_act_buffer_inst_act_if_inst_n54,
         wrap_act_buffer_inst_act_if_inst_n53,
         wrap_act_buffer_inst_act_if_inst_n52,
         wrap_act_buffer_inst_act_if_inst_n51,
         wrap_act_buffer_inst_act_if_inst_n50,
         wrap_act_buffer_inst_act_if_inst_n49,
         wrap_act_buffer_inst_act_if_inst_n48,
         wrap_act_buffer_inst_act_if_inst_n47,
         wrap_act_buffer_inst_act_if_inst_n46,
         wrap_act_buffer_inst_act_if_inst_n45,
         wrap_act_buffer_inst_act_if_inst_n44,
         wrap_act_buffer_inst_act_if_inst_n43,
         wrap_act_buffer_inst_act_if_inst_n42,
         wrap_act_buffer_inst_act_if_inst_n41,
         wrap_act_buffer_inst_act_if_inst_n40,
         wrap_act_buffer_inst_act_if_inst_n39,
         wrap_act_buffer_inst_act_if_inst_n2,
         wrap_act_buffer_inst_act_if_inst_n1,
         wrap_act_buffer_inst_act_if_inst_n38,
         wrap_act_buffer_inst_act_if_inst_n37,
         wrap_act_buffer_inst_act_if_inst_n36,
         wrap_act_buffer_inst_act_if_inst_n35,
         wrap_act_buffer_inst_act_if_inst_n34,
         wrap_act_buffer_inst_act_if_inst_n33,
         wrap_act_buffer_inst_act_if_inst_n32,
         wrap_act_buffer_inst_act_if_inst_n31,
         wrap_act_buffer_inst_act_if_inst_n30,
         wrap_act_buffer_inst_act_if_inst_n29,
         wrap_act_buffer_inst_act_if_inst_n28,
         wrap_act_buffer_inst_act_if_inst_n27,
         wrap_act_buffer_inst_act_if_inst_n26,
         wrap_act_buffer_inst_act_if_inst_n25,
         wrap_act_buffer_inst_act_if_inst_n24,
         wrap_act_buffer_inst_act_if_inst_n23,
         wrap_act_buffer_inst_act_if_inst_n22,
         wrap_act_buffer_inst_act_if_inst_n21,
         wrap_act_buffer_inst_act_if_inst_n20,
         wrap_act_buffer_inst_act_if_inst_n19,
         wrap_act_buffer_inst_act_if_inst_n18,
         wrap_act_buffer_inst_act_if_inst_n17,
         wrap_act_buffer_inst_act_if_inst_n16,
         wrap_act_buffer_inst_act_if_inst_n15,
         wrap_act_buffer_inst_act_if_inst_n14,
         wrap_act_buffer_inst_act_if_inst_n13,
         wrap_act_buffer_inst_act_if_inst_n12,
         wrap_act_buffer_inst_act_if_inst_n11,
         wrap_act_buffer_inst_act_if_inst_n10,
         wrap_act_buffer_inst_act_if_inst_n9,
         wrap_act_buffer_inst_act_if_inst_n8,
         wrap_act_buffer_inst_act_if_inst_n7,
         wrap_act_buffer_inst_act_if_inst_n6,
         wrap_act_buffer_inst_act_if_inst_n5,
         wrap_act_buffer_inst_act_if_inst_n4,
         wrap_act_buffer_inst_act_if_inst_n3, npu_inst_n143, npu_inst_n142,
         npu_inst_n141, npu_inst_n140, npu_inst_n139, npu_inst_n138,
         npu_inst_n137, npu_inst_n136, npu_inst_n135, npu_inst_n134,
         npu_inst_n133, npu_inst_n132, npu_inst_n131, npu_inst_n130,
         npu_inst_n129, npu_inst_n128, npu_inst_n127, npu_inst_n126,
         npu_inst_n125, npu_inst_n124, npu_inst_n123, npu_inst_n122,
         npu_inst_n121, npu_inst_n120, npu_inst_n119, npu_inst_n118,
         npu_inst_n117, npu_inst_n116, npu_inst_n115, npu_inst_n114,
         npu_inst_n113, npu_inst_n112, npu_inst_n111, npu_inst_n110,
         npu_inst_n109, npu_inst_n108, npu_inst_n107, npu_inst_n106,
         npu_inst_n105, npu_inst_n104, npu_inst_n103, npu_inst_n102,
         npu_inst_n101, npu_inst_n100, npu_inst_n99, npu_inst_n98,
         npu_inst_n97, npu_inst_n96, npu_inst_n95, npu_inst_n94, npu_inst_n93,
         npu_inst_n92, npu_inst_n91, npu_inst_n90, npu_inst_n89, npu_inst_n88,
         npu_inst_n87, npu_inst_n86, npu_inst_n85, npu_inst_n84, npu_inst_n83,
         npu_inst_n82, npu_inst_n81, npu_inst_n80, npu_inst_n79, npu_inst_n78,
         npu_inst_n77, npu_inst_n76, npu_inst_n75, npu_inst_n74, npu_inst_n73,
         npu_inst_n72, npu_inst_n71, npu_inst_n70, npu_inst_n69, npu_inst_n68,
         npu_inst_n67, npu_inst_n66, npu_inst_n65, npu_inst_n64, npu_inst_n63,
         npu_inst_n62, npu_inst_n61, npu_inst_n60, npu_inst_n59, npu_inst_n58,
         npu_inst_n57, npu_inst_n56, npu_inst_n55, npu_inst_n54, npu_inst_n53,
         npu_inst_n52, npu_inst_n51, npu_inst_n50, npu_inst_n49, npu_inst_n48,
         npu_inst_n47, npu_inst_n46, npu_inst_n45, npu_inst_n44, npu_inst_n43,
         npu_inst_n42, npu_inst_n41, npu_inst_n40, npu_inst_n39, npu_inst_n38,
         npu_inst_n37, npu_inst_n36, npu_inst_n35, npu_inst_n34, npu_inst_n33,
         npu_inst_n32, npu_inst_n31, npu_inst_n30, npu_inst_n29, npu_inst_n28,
         npu_inst_n27, npu_inst_n26, npu_inst_n25, npu_inst_n24, npu_inst_n23,
         npu_inst_n22, npu_inst_n21, npu_inst_n20, npu_inst_n19, npu_inst_n18,
         npu_inst_n17, npu_inst_n16, npu_inst_n15, npu_inst_n14, npu_inst_n13,
         npu_inst_n12, npu_inst_n11, npu_inst_n10, npu_inst_n9, npu_inst_n8,
         npu_inst_n7, npu_inst_n6, npu_inst_n5, npu_inst_n4, npu_inst_n3,
         npu_inst_n2, npu_inst_n1, npu_inst_int_data_x_7__7__0_,
         npu_inst_int_data_x_7__7__1_, npu_inst_int_data_x_7__6__0_,
         npu_inst_int_data_x_7__6__1_, npu_inst_int_data_x_7__5__0_,
         npu_inst_int_data_x_7__5__1_, npu_inst_int_data_x_7__4__0_,
         npu_inst_int_data_x_7__4__1_, npu_inst_int_data_x_7__3__0_,
         npu_inst_int_data_x_7__3__1_, npu_inst_int_data_x_7__2__0_,
         npu_inst_int_data_x_7__2__1_, npu_inst_int_data_x_7__1__0_,
         npu_inst_int_data_x_7__1__1_, npu_inst_int_data_x_6__7__0_,
         npu_inst_int_data_x_6__7__1_, npu_inst_int_data_x_6__6__0_,
         npu_inst_int_data_x_6__6__1_, npu_inst_int_data_x_6__5__0_,
         npu_inst_int_data_x_6__5__1_, npu_inst_int_data_x_6__4__0_,
         npu_inst_int_data_x_6__4__1_, npu_inst_int_data_x_6__3__0_,
         npu_inst_int_data_x_6__3__1_, npu_inst_int_data_x_6__2__0_,
         npu_inst_int_data_x_6__2__1_, npu_inst_int_data_x_6__1__0_,
         npu_inst_int_data_x_6__1__1_, npu_inst_int_data_x_5__7__0_,
         npu_inst_int_data_x_5__7__1_, npu_inst_int_data_x_5__6__0_,
         npu_inst_int_data_x_5__6__1_, npu_inst_int_data_x_5__5__0_,
         npu_inst_int_data_x_5__5__1_, npu_inst_int_data_x_5__4__0_,
         npu_inst_int_data_x_5__4__1_, npu_inst_int_data_x_5__3__0_,
         npu_inst_int_data_x_5__3__1_, npu_inst_int_data_x_5__2__0_,
         npu_inst_int_data_x_5__2__1_, npu_inst_int_data_x_5__1__0_,
         npu_inst_int_data_x_5__1__1_, npu_inst_int_data_x_4__7__0_,
         npu_inst_int_data_x_4__7__1_, npu_inst_int_data_x_4__6__0_,
         npu_inst_int_data_x_4__6__1_, npu_inst_int_data_x_4__5__0_,
         npu_inst_int_data_x_4__5__1_, npu_inst_int_data_x_4__4__0_,
         npu_inst_int_data_x_4__4__1_, npu_inst_int_data_x_4__3__0_,
         npu_inst_int_data_x_4__3__1_, npu_inst_int_data_x_4__2__0_,
         npu_inst_int_data_x_4__2__1_, npu_inst_int_data_x_4__1__0_,
         npu_inst_int_data_x_4__1__1_, npu_inst_int_data_x_3__7__0_,
         npu_inst_int_data_x_3__7__1_, npu_inst_int_data_x_3__6__0_,
         npu_inst_int_data_x_3__6__1_, npu_inst_int_data_x_3__5__0_,
         npu_inst_int_data_x_3__5__1_, npu_inst_int_data_x_3__4__0_,
         npu_inst_int_data_x_3__4__1_, npu_inst_int_data_x_3__3__0_,
         npu_inst_int_data_x_3__3__1_, npu_inst_int_data_x_3__2__0_,
         npu_inst_int_data_x_3__2__1_, npu_inst_int_data_x_3__1__0_,
         npu_inst_int_data_x_3__1__1_, npu_inst_int_data_x_2__7__0_,
         npu_inst_int_data_x_2__7__1_, npu_inst_int_data_x_2__6__0_,
         npu_inst_int_data_x_2__6__1_, npu_inst_int_data_x_2__5__0_,
         npu_inst_int_data_x_2__5__1_, npu_inst_int_data_x_2__4__0_,
         npu_inst_int_data_x_2__4__1_, npu_inst_int_data_x_2__3__0_,
         npu_inst_int_data_x_2__3__1_, npu_inst_int_data_x_2__2__0_,
         npu_inst_int_data_x_2__2__1_, npu_inst_int_data_x_2__1__0_,
         npu_inst_int_data_x_2__1__1_, npu_inst_int_data_x_1__7__0_,
         npu_inst_int_data_x_1__7__1_, npu_inst_int_data_x_1__6__0_,
         npu_inst_int_data_x_1__6__1_, npu_inst_int_data_x_1__5__0_,
         npu_inst_int_data_x_1__5__1_, npu_inst_int_data_x_1__4__0_,
         npu_inst_int_data_x_1__4__1_, npu_inst_int_data_x_1__3__0_,
         npu_inst_int_data_x_1__3__1_, npu_inst_int_data_x_1__2__0_,
         npu_inst_int_data_x_1__2__1_, npu_inst_int_data_x_1__1__0_,
         npu_inst_int_data_x_1__1__1_, npu_inst_int_data_x_0__7__0_,
         npu_inst_int_data_x_0__7__1_, npu_inst_int_data_x_0__6__0_,
         npu_inst_int_data_x_0__6__1_, npu_inst_int_data_x_0__5__0_,
         npu_inst_int_data_x_0__5__1_, npu_inst_int_data_x_0__4__0_,
         npu_inst_int_data_x_0__4__1_, npu_inst_int_data_x_0__3__0_,
         npu_inst_int_data_x_0__3__1_, npu_inst_int_data_x_0__2__0_,
         npu_inst_int_data_x_0__2__1_, npu_inst_int_data_x_0__1__0_,
         npu_inst_int_data_x_0__1__1_, npu_inst_int_data_y_7__7__0_,
         npu_inst_int_data_y_7__7__1_, npu_inst_int_data_y_7__6__0_,
         npu_inst_int_data_y_7__6__1_, npu_inst_int_data_y_7__5__0_,
         npu_inst_int_data_y_7__5__1_, npu_inst_int_data_y_7__4__0_,
         npu_inst_int_data_y_7__4__1_, npu_inst_int_data_y_7__3__0_,
         npu_inst_int_data_y_7__3__1_, npu_inst_int_data_y_7__2__0_,
         npu_inst_int_data_y_7__2__1_, npu_inst_int_data_y_7__1__0_,
         npu_inst_int_data_y_7__1__1_, npu_inst_int_data_y_7__0__0_,
         npu_inst_int_data_y_7__0__1_, npu_inst_int_data_y_6__7__0_,
         npu_inst_int_data_y_6__7__1_, npu_inst_int_data_y_6__6__0_,
         npu_inst_int_data_y_6__6__1_, npu_inst_int_data_y_6__5__0_,
         npu_inst_int_data_y_6__5__1_, npu_inst_int_data_y_6__4__0_,
         npu_inst_int_data_y_6__4__1_, npu_inst_int_data_y_6__3__0_,
         npu_inst_int_data_y_6__3__1_, npu_inst_int_data_y_6__2__0_,
         npu_inst_int_data_y_6__2__1_, npu_inst_int_data_y_6__1__0_,
         npu_inst_int_data_y_6__1__1_, npu_inst_int_data_y_6__0__0_,
         npu_inst_int_data_y_6__0__1_, npu_inst_int_data_y_5__7__0_,
         npu_inst_int_data_y_5__7__1_, npu_inst_int_data_y_5__6__0_,
         npu_inst_int_data_y_5__6__1_, npu_inst_int_data_y_5__5__0_,
         npu_inst_int_data_y_5__5__1_, npu_inst_int_data_y_5__4__0_,
         npu_inst_int_data_y_5__4__1_, npu_inst_int_data_y_5__3__0_,
         npu_inst_int_data_y_5__3__1_, npu_inst_int_data_y_5__2__0_,
         npu_inst_int_data_y_5__2__1_, npu_inst_int_data_y_5__1__0_,
         npu_inst_int_data_y_5__1__1_, npu_inst_int_data_y_5__0__0_,
         npu_inst_int_data_y_5__0__1_, npu_inst_int_data_y_4__7__0_,
         npu_inst_int_data_y_4__7__1_, npu_inst_int_data_y_4__6__0_,
         npu_inst_int_data_y_4__6__1_, npu_inst_int_data_y_4__5__0_,
         npu_inst_int_data_y_4__5__1_, npu_inst_int_data_y_4__4__0_,
         npu_inst_int_data_y_4__4__1_, npu_inst_int_data_y_4__3__0_,
         npu_inst_int_data_y_4__3__1_, npu_inst_int_data_y_4__2__0_,
         npu_inst_int_data_y_4__2__1_, npu_inst_int_data_y_4__1__0_,
         npu_inst_int_data_y_4__1__1_, npu_inst_int_data_y_4__0__0_,
         npu_inst_int_data_y_4__0__1_, npu_inst_int_data_y_3__7__0_,
         npu_inst_int_data_y_3__7__1_, npu_inst_int_data_y_3__6__0_,
         npu_inst_int_data_y_3__6__1_, npu_inst_int_data_y_3__5__0_,
         npu_inst_int_data_y_3__5__1_, npu_inst_int_data_y_3__4__0_,
         npu_inst_int_data_y_3__4__1_, npu_inst_int_data_y_3__3__0_,
         npu_inst_int_data_y_3__3__1_, npu_inst_int_data_y_3__2__0_,
         npu_inst_int_data_y_3__2__1_, npu_inst_int_data_y_3__1__0_,
         npu_inst_int_data_y_3__1__1_, npu_inst_int_data_y_3__0__0_,
         npu_inst_int_data_y_3__0__1_, npu_inst_int_data_y_2__7__0_,
         npu_inst_int_data_y_2__7__1_, npu_inst_int_data_y_2__6__0_,
         npu_inst_int_data_y_2__6__1_, npu_inst_int_data_y_2__5__0_,
         npu_inst_int_data_y_2__5__1_, npu_inst_int_data_y_2__4__0_,
         npu_inst_int_data_y_2__4__1_, npu_inst_int_data_y_2__3__0_,
         npu_inst_int_data_y_2__3__1_, npu_inst_int_data_y_2__2__0_,
         npu_inst_int_data_y_2__2__1_, npu_inst_int_data_y_2__1__0_,
         npu_inst_int_data_y_2__1__1_, npu_inst_int_data_y_2__0__0_,
         npu_inst_int_data_y_2__0__1_, npu_inst_int_data_y_1__7__0_,
         npu_inst_int_data_y_1__7__1_, npu_inst_int_data_y_1__6__0_,
         npu_inst_int_data_y_1__6__1_, npu_inst_int_data_y_1__5__0_,
         npu_inst_int_data_y_1__5__1_, npu_inst_int_data_y_1__4__0_,
         npu_inst_int_data_y_1__4__1_, npu_inst_int_data_y_1__3__0_,
         npu_inst_int_data_y_1__3__1_, npu_inst_int_data_y_1__2__0_,
         npu_inst_int_data_y_1__2__1_, npu_inst_int_data_y_1__1__0_,
         npu_inst_int_data_y_1__1__1_, npu_inst_int_data_y_1__0__0_,
         npu_inst_int_data_y_1__0__1_, npu_inst_int_data_res_7__7__0_,
         npu_inst_int_data_res_7__7__1_, npu_inst_int_data_res_7__7__2_,
         npu_inst_int_data_res_7__7__3_, npu_inst_int_data_res_7__7__4_,
         npu_inst_int_data_res_7__7__5_, npu_inst_int_data_res_7__7__6_,
         npu_inst_int_data_res_7__7__7_, npu_inst_int_data_res_7__6__0_,
         npu_inst_int_data_res_7__6__1_, npu_inst_int_data_res_7__6__2_,
         npu_inst_int_data_res_7__6__3_, npu_inst_int_data_res_7__6__4_,
         npu_inst_int_data_res_7__6__5_, npu_inst_int_data_res_7__6__6_,
         npu_inst_int_data_res_7__6__7_, npu_inst_int_data_res_7__5__0_,
         npu_inst_int_data_res_7__5__1_, npu_inst_int_data_res_7__5__2_,
         npu_inst_int_data_res_7__5__3_, npu_inst_int_data_res_7__5__4_,
         npu_inst_int_data_res_7__5__5_, npu_inst_int_data_res_7__5__6_,
         npu_inst_int_data_res_7__5__7_, npu_inst_int_data_res_7__4__0_,
         npu_inst_int_data_res_7__4__1_, npu_inst_int_data_res_7__4__2_,
         npu_inst_int_data_res_7__4__3_, npu_inst_int_data_res_7__4__4_,
         npu_inst_int_data_res_7__4__5_, npu_inst_int_data_res_7__4__6_,
         npu_inst_int_data_res_7__4__7_, npu_inst_int_data_res_7__3__0_,
         npu_inst_int_data_res_7__3__1_, npu_inst_int_data_res_7__3__2_,
         npu_inst_int_data_res_7__3__3_, npu_inst_int_data_res_7__3__4_,
         npu_inst_int_data_res_7__3__5_, npu_inst_int_data_res_7__3__6_,
         npu_inst_int_data_res_7__3__7_, npu_inst_int_data_res_7__2__0_,
         npu_inst_int_data_res_7__2__1_, npu_inst_int_data_res_7__2__2_,
         npu_inst_int_data_res_7__2__3_, npu_inst_int_data_res_7__2__4_,
         npu_inst_int_data_res_7__2__5_, npu_inst_int_data_res_7__2__6_,
         npu_inst_int_data_res_7__2__7_, npu_inst_int_data_res_7__1__0_,
         npu_inst_int_data_res_7__1__1_, npu_inst_int_data_res_7__1__2_,
         npu_inst_int_data_res_7__1__3_, npu_inst_int_data_res_7__1__4_,
         npu_inst_int_data_res_7__1__5_, npu_inst_int_data_res_7__1__6_,
         npu_inst_int_data_res_7__1__7_, npu_inst_int_data_res_7__0__0_,
         npu_inst_int_data_res_7__0__1_, npu_inst_int_data_res_7__0__2_,
         npu_inst_int_data_res_7__0__3_, npu_inst_int_data_res_7__0__4_,
         npu_inst_int_data_res_7__0__5_, npu_inst_int_data_res_7__0__6_,
         npu_inst_int_data_res_7__0__7_, npu_inst_int_data_res_6__7__0_,
         npu_inst_int_data_res_6__7__1_, npu_inst_int_data_res_6__7__2_,
         npu_inst_int_data_res_6__7__3_, npu_inst_int_data_res_6__7__4_,
         npu_inst_int_data_res_6__7__5_, npu_inst_int_data_res_6__7__6_,
         npu_inst_int_data_res_6__7__7_, npu_inst_int_data_res_6__6__0_,
         npu_inst_int_data_res_6__6__1_, npu_inst_int_data_res_6__6__2_,
         npu_inst_int_data_res_6__6__3_, npu_inst_int_data_res_6__6__4_,
         npu_inst_int_data_res_6__6__5_, npu_inst_int_data_res_6__6__6_,
         npu_inst_int_data_res_6__6__7_, npu_inst_int_data_res_6__5__0_,
         npu_inst_int_data_res_6__5__1_, npu_inst_int_data_res_6__5__2_,
         npu_inst_int_data_res_6__5__3_, npu_inst_int_data_res_6__5__4_,
         npu_inst_int_data_res_6__5__5_, npu_inst_int_data_res_6__5__6_,
         npu_inst_int_data_res_6__5__7_, npu_inst_int_data_res_6__4__0_,
         npu_inst_int_data_res_6__4__1_, npu_inst_int_data_res_6__4__2_,
         npu_inst_int_data_res_6__4__3_, npu_inst_int_data_res_6__4__4_,
         npu_inst_int_data_res_6__4__5_, npu_inst_int_data_res_6__4__6_,
         npu_inst_int_data_res_6__4__7_, npu_inst_int_data_res_6__3__0_,
         npu_inst_int_data_res_6__3__1_, npu_inst_int_data_res_6__3__2_,
         npu_inst_int_data_res_6__3__3_, npu_inst_int_data_res_6__3__4_,
         npu_inst_int_data_res_6__3__5_, npu_inst_int_data_res_6__3__6_,
         npu_inst_int_data_res_6__3__7_, npu_inst_int_data_res_6__2__0_,
         npu_inst_int_data_res_6__2__1_, npu_inst_int_data_res_6__2__2_,
         npu_inst_int_data_res_6__2__3_, npu_inst_int_data_res_6__2__4_,
         npu_inst_int_data_res_6__2__5_, npu_inst_int_data_res_6__2__6_,
         npu_inst_int_data_res_6__2__7_, npu_inst_int_data_res_6__1__0_,
         npu_inst_int_data_res_6__1__1_, npu_inst_int_data_res_6__1__2_,
         npu_inst_int_data_res_6__1__3_, npu_inst_int_data_res_6__1__4_,
         npu_inst_int_data_res_6__1__5_, npu_inst_int_data_res_6__1__6_,
         npu_inst_int_data_res_6__1__7_, npu_inst_int_data_res_6__0__0_,
         npu_inst_int_data_res_6__0__1_, npu_inst_int_data_res_6__0__2_,
         npu_inst_int_data_res_6__0__3_, npu_inst_int_data_res_6__0__4_,
         npu_inst_int_data_res_6__0__5_, npu_inst_int_data_res_6__0__6_,
         npu_inst_int_data_res_6__0__7_, npu_inst_int_data_res_5__7__0_,
         npu_inst_int_data_res_5__7__1_, npu_inst_int_data_res_5__7__2_,
         npu_inst_int_data_res_5__7__3_, npu_inst_int_data_res_5__7__4_,
         npu_inst_int_data_res_5__7__5_, npu_inst_int_data_res_5__7__6_,
         npu_inst_int_data_res_5__7__7_, npu_inst_int_data_res_5__6__0_,
         npu_inst_int_data_res_5__6__1_, npu_inst_int_data_res_5__6__2_,
         npu_inst_int_data_res_5__6__3_, npu_inst_int_data_res_5__6__4_,
         npu_inst_int_data_res_5__6__5_, npu_inst_int_data_res_5__6__6_,
         npu_inst_int_data_res_5__6__7_, npu_inst_int_data_res_5__5__0_,
         npu_inst_int_data_res_5__5__1_, npu_inst_int_data_res_5__5__2_,
         npu_inst_int_data_res_5__5__3_, npu_inst_int_data_res_5__5__4_,
         npu_inst_int_data_res_5__5__5_, npu_inst_int_data_res_5__5__6_,
         npu_inst_int_data_res_5__5__7_, npu_inst_int_data_res_5__4__0_,
         npu_inst_int_data_res_5__4__1_, npu_inst_int_data_res_5__4__2_,
         npu_inst_int_data_res_5__4__3_, npu_inst_int_data_res_5__4__4_,
         npu_inst_int_data_res_5__4__5_, npu_inst_int_data_res_5__4__6_,
         npu_inst_int_data_res_5__4__7_, npu_inst_int_data_res_5__3__0_,
         npu_inst_int_data_res_5__3__1_, npu_inst_int_data_res_5__3__2_,
         npu_inst_int_data_res_5__3__3_, npu_inst_int_data_res_5__3__4_,
         npu_inst_int_data_res_5__3__5_, npu_inst_int_data_res_5__3__6_,
         npu_inst_int_data_res_5__3__7_, npu_inst_int_data_res_5__2__0_,
         npu_inst_int_data_res_5__2__1_, npu_inst_int_data_res_5__2__2_,
         npu_inst_int_data_res_5__2__3_, npu_inst_int_data_res_5__2__4_,
         npu_inst_int_data_res_5__2__5_, npu_inst_int_data_res_5__2__6_,
         npu_inst_int_data_res_5__2__7_, npu_inst_int_data_res_5__1__0_,
         npu_inst_int_data_res_5__1__1_, npu_inst_int_data_res_5__1__2_,
         npu_inst_int_data_res_5__1__3_, npu_inst_int_data_res_5__1__4_,
         npu_inst_int_data_res_5__1__5_, npu_inst_int_data_res_5__1__6_,
         npu_inst_int_data_res_5__1__7_, npu_inst_int_data_res_5__0__0_,
         npu_inst_int_data_res_5__0__1_, npu_inst_int_data_res_5__0__2_,
         npu_inst_int_data_res_5__0__3_, npu_inst_int_data_res_5__0__4_,
         npu_inst_int_data_res_5__0__5_, npu_inst_int_data_res_5__0__6_,
         npu_inst_int_data_res_5__0__7_, npu_inst_int_data_res_4__7__0_,
         npu_inst_int_data_res_4__7__1_, npu_inst_int_data_res_4__7__2_,
         npu_inst_int_data_res_4__7__3_, npu_inst_int_data_res_4__7__4_,
         npu_inst_int_data_res_4__7__5_, npu_inst_int_data_res_4__7__6_,
         npu_inst_int_data_res_4__7__7_, npu_inst_int_data_res_4__6__0_,
         npu_inst_int_data_res_4__6__1_, npu_inst_int_data_res_4__6__2_,
         npu_inst_int_data_res_4__6__3_, npu_inst_int_data_res_4__6__4_,
         npu_inst_int_data_res_4__6__5_, npu_inst_int_data_res_4__6__6_,
         npu_inst_int_data_res_4__6__7_, npu_inst_int_data_res_4__5__0_,
         npu_inst_int_data_res_4__5__1_, npu_inst_int_data_res_4__5__2_,
         npu_inst_int_data_res_4__5__3_, npu_inst_int_data_res_4__5__4_,
         npu_inst_int_data_res_4__5__5_, npu_inst_int_data_res_4__5__6_,
         npu_inst_int_data_res_4__5__7_, npu_inst_int_data_res_4__4__0_,
         npu_inst_int_data_res_4__4__1_, npu_inst_int_data_res_4__4__2_,
         npu_inst_int_data_res_4__4__3_, npu_inst_int_data_res_4__4__4_,
         npu_inst_int_data_res_4__4__5_, npu_inst_int_data_res_4__4__6_,
         npu_inst_int_data_res_4__4__7_, npu_inst_int_data_res_4__3__0_,
         npu_inst_int_data_res_4__3__1_, npu_inst_int_data_res_4__3__2_,
         npu_inst_int_data_res_4__3__3_, npu_inst_int_data_res_4__3__4_,
         npu_inst_int_data_res_4__3__5_, npu_inst_int_data_res_4__3__6_,
         npu_inst_int_data_res_4__3__7_, npu_inst_int_data_res_4__2__0_,
         npu_inst_int_data_res_4__2__1_, npu_inst_int_data_res_4__2__2_,
         npu_inst_int_data_res_4__2__3_, npu_inst_int_data_res_4__2__4_,
         npu_inst_int_data_res_4__2__5_, npu_inst_int_data_res_4__2__6_,
         npu_inst_int_data_res_4__2__7_, npu_inst_int_data_res_4__1__0_,
         npu_inst_int_data_res_4__1__1_, npu_inst_int_data_res_4__1__2_,
         npu_inst_int_data_res_4__1__3_, npu_inst_int_data_res_4__1__4_,
         npu_inst_int_data_res_4__1__5_, npu_inst_int_data_res_4__1__6_,
         npu_inst_int_data_res_4__1__7_, npu_inst_int_data_res_4__0__0_,
         npu_inst_int_data_res_4__0__1_, npu_inst_int_data_res_4__0__2_,
         npu_inst_int_data_res_4__0__3_, npu_inst_int_data_res_4__0__4_,
         npu_inst_int_data_res_4__0__5_, npu_inst_int_data_res_4__0__6_,
         npu_inst_int_data_res_4__0__7_, npu_inst_int_data_res_3__7__0_,
         npu_inst_int_data_res_3__7__1_, npu_inst_int_data_res_3__7__2_,
         npu_inst_int_data_res_3__7__3_, npu_inst_int_data_res_3__7__4_,
         npu_inst_int_data_res_3__7__5_, npu_inst_int_data_res_3__7__6_,
         npu_inst_int_data_res_3__7__7_, npu_inst_int_data_res_3__6__0_,
         npu_inst_int_data_res_3__6__1_, npu_inst_int_data_res_3__6__2_,
         npu_inst_int_data_res_3__6__3_, npu_inst_int_data_res_3__6__4_,
         npu_inst_int_data_res_3__6__5_, npu_inst_int_data_res_3__6__6_,
         npu_inst_int_data_res_3__6__7_, npu_inst_int_data_res_3__5__0_,
         npu_inst_int_data_res_3__5__1_, npu_inst_int_data_res_3__5__2_,
         npu_inst_int_data_res_3__5__3_, npu_inst_int_data_res_3__5__4_,
         npu_inst_int_data_res_3__5__5_, npu_inst_int_data_res_3__5__6_,
         npu_inst_int_data_res_3__5__7_, npu_inst_int_data_res_3__4__0_,
         npu_inst_int_data_res_3__4__1_, npu_inst_int_data_res_3__4__2_,
         npu_inst_int_data_res_3__4__3_, npu_inst_int_data_res_3__4__4_,
         npu_inst_int_data_res_3__4__5_, npu_inst_int_data_res_3__4__6_,
         npu_inst_int_data_res_3__4__7_, npu_inst_int_data_res_3__3__0_,
         npu_inst_int_data_res_3__3__1_, npu_inst_int_data_res_3__3__2_,
         npu_inst_int_data_res_3__3__3_, npu_inst_int_data_res_3__3__4_,
         npu_inst_int_data_res_3__3__5_, npu_inst_int_data_res_3__3__6_,
         npu_inst_int_data_res_3__3__7_, npu_inst_int_data_res_3__2__0_,
         npu_inst_int_data_res_3__2__1_, npu_inst_int_data_res_3__2__2_,
         npu_inst_int_data_res_3__2__3_, npu_inst_int_data_res_3__2__4_,
         npu_inst_int_data_res_3__2__5_, npu_inst_int_data_res_3__2__6_,
         npu_inst_int_data_res_3__2__7_, npu_inst_int_data_res_3__1__0_,
         npu_inst_int_data_res_3__1__1_, npu_inst_int_data_res_3__1__2_,
         npu_inst_int_data_res_3__1__3_, npu_inst_int_data_res_3__1__4_,
         npu_inst_int_data_res_3__1__5_, npu_inst_int_data_res_3__1__6_,
         npu_inst_int_data_res_3__1__7_, npu_inst_int_data_res_3__0__0_,
         npu_inst_int_data_res_3__0__1_, npu_inst_int_data_res_3__0__2_,
         npu_inst_int_data_res_3__0__3_, npu_inst_int_data_res_3__0__4_,
         npu_inst_int_data_res_3__0__5_, npu_inst_int_data_res_3__0__6_,
         npu_inst_int_data_res_3__0__7_, npu_inst_int_data_res_2__7__0_,
         npu_inst_int_data_res_2__7__1_, npu_inst_int_data_res_2__7__2_,
         npu_inst_int_data_res_2__7__3_, npu_inst_int_data_res_2__7__4_,
         npu_inst_int_data_res_2__7__5_, npu_inst_int_data_res_2__7__6_,
         npu_inst_int_data_res_2__7__7_, npu_inst_int_data_res_2__6__0_,
         npu_inst_int_data_res_2__6__1_, npu_inst_int_data_res_2__6__2_,
         npu_inst_int_data_res_2__6__3_, npu_inst_int_data_res_2__6__4_,
         npu_inst_int_data_res_2__6__5_, npu_inst_int_data_res_2__6__6_,
         npu_inst_int_data_res_2__6__7_, npu_inst_int_data_res_2__5__0_,
         npu_inst_int_data_res_2__5__1_, npu_inst_int_data_res_2__5__2_,
         npu_inst_int_data_res_2__5__3_, npu_inst_int_data_res_2__5__4_,
         npu_inst_int_data_res_2__5__5_, npu_inst_int_data_res_2__5__6_,
         npu_inst_int_data_res_2__5__7_, npu_inst_int_data_res_2__4__0_,
         npu_inst_int_data_res_2__4__1_, npu_inst_int_data_res_2__4__2_,
         npu_inst_int_data_res_2__4__3_, npu_inst_int_data_res_2__4__4_,
         npu_inst_int_data_res_2__4__5_, npu_inst_int_data_res_2__4__6_,
         npu_inst_int_data_res_2__4__7_, npu_inst_int_data_res_2__3__0_,
         npu_inst_int_data_res_2__3__1_, npu_inst_int_data_res_2__3__2_,
         npu_inst_int_data_res_2__3__3_, npu_inst_int_data_res_2__3__4_,
         npu_inst_int_data_res_2__3__5_, npu_inst_int_data_res_2__3__6_,
         npu_inst_int_data_res_2__3__7_, npu_inst_int_data_res_2__2__0_,
         npu_inst_int_data_res_2__2__1_, npu_inst_int_data_res_2__2__2_,
         npu_inst_int_data_res_2__2__3_, npu_inst_int_data_res_2__2__4_,
         npu_inst_int_data_res_2__2__5_, npu_inst_int_data_res_2__2__6_,
         npu_inst_int_data_res_2__2__7_, npu_inst_int_data_res_2__1__0_,
         npu_inst_int_data_res_2__1__1_, npu_inst_int_data_res_2__1__2_,
         npu_inst_int_data_res_2__1__3_, npu_inst_int_data_res_2__1__4_,
         npu_inst_int_data_res_2__1__5_, npu_inst_int_data_res_2__1__6_,
         npu_inst_int_data_res_2__1__7_, npu_inst_int_data_res_2__0__0_,
         npu_inst_int_data_res_2__0__1_, npu_inst_int_data_res_2__0__2_,
         npu_inst_int_data_res_2__0__3_, npu_inst_int_data_res_2__0__4_,
         npu_inst_int_data_res_2__0__5_, npu_inst_int_data_res_2__0__6_,
         npu_inst_int_data_res_2__0__7_, npu_inst_int_data_res_1__7__0_,
         npu_inst_int_data_res_1__7__1_, npu_inst_int_data_res_1__7__2_,
         npu_inst_int_data_res_1__7__3_, npu_inst_int_data_res_1__7__4_,
         npu_inst_int_data_res_1__7__5_, npu_inst_int_data_res_1__7__6_,
         npu_inst_int_data_res_1__7__7_, npu_inst_int_data_res_1__6__0_,
         npu_inst_int_data_res_1__6__1_, npu_inst_int_data_res_1__6__2_,
         npu_inst_int_data_res_1__6__3_, npu_inst_int_data_res_1__6__4_,
         npu_inst_int_data_res_1__6__5_, npu_inst_int_data_res_1__6__6_,
         npu_inst_int_data_res_1__6__7_, npu_inst_int_data_res_1__5__0_,
         npu_inst_int_data_res_1__5__1_, npu_inst_int_data_res_1__5__2_,
         npu_inst_int_data_res_1__5__3_, npu_inst_int_data_res_1__5__4_,
         npu_inst_int_data_res_1__5__5_, npu_inst_int_data_res_1__5__6_,
         npu_inst_int_data_res_1__5__7_, npu_inst_int_data_res_1__4__0_,
         npu_inst_int_data_res_1__4__1_, npu_inst_int_data_res_1__4__2_,
         npu_inst_int_data_res_1__4__3_, npu_inst_int_data_res_1__4__4_,
         npu_inst_int_data_res_1__4__5_, npu_inst_int_data_res_1__4__6_,
         npu_inst_int_data_res_1__4__7_, npu_inst_int_data_res_1__3__0_,
         npu_inst_int_data_res_1__3__1_, npu_inst_int_data_res_1__3__2_,
         npu_inst_int_data_res_1__3__3_, npu_inst_int_data_res_1__3__4_,
         npu_inst_int_data_res_1__3__5_, npu_inst_int_data_res_1__3__6_,
         npu_inst_int_data_res_1__3__7_, npu_inst_int_data_res_1__2__0_,
         npu_inst_int_data_res_1__2__1_, npu_inst_int_data_res_1__2__2_,
         npu_inst_int_data_res_1__2__3_, npu_inst_int_data_res_1__2__4_,
         npu_inst_int_data_res_1__2__5_, npu_inst_int_data_res_1__2__6_,
         npu_inst_int_data_res_1__2__7_, npu_inst_int_data_res_1__1__0_,
         npu_inst_int_data_res_1__1__1_, npu_inst_int_data_res_1__1__2_,
         npu_inst_int_data_res_1__1__3_, npu_inst_int_data_res_1__1__4_,
         npu_inst_int_data_res_1__1__5_, npu_inst_int_data_res_1__1__6_,
         npu_inst_int_data_res_1__1__7_, npu_inst_int_data_res_1__0__0_,
         npu_inst_int_data_res_1__0__1_, npu_inst_int_data_res_1__0__2_,
         npu_inst_int_data_res_1__0__3_, npu_inst_int_data_res_1__0__4_,
         npu_inst_int_data_res_1__0__5_, npu_inst_int_data_res_1__0__6_,
         npu_inst_int_data_res_1__0__7_, npu_inst_pe_1_0_0_n118,
         npu_inst_pe_1_0_0_n117, npu_inst_pe_1_0_0_n116,
         npu_inst_pe_1_0_0_n115, npu_inst_pe_1_0_0_n114,
         npu_inst_pe_1_0_0_n113, npu_inst_pe_1_0_0_n112,
         npu_inst_pe_1_0_0_n111, npu_inst_pe_1_0_0_n110,
         npu_inst_pe_1_0_0_n109, npu_inst_pe_1_0_0_n108,
         npu_inst_pe_1_0_0_n107, npu_inst_pe_1_0_0_n106,
         npu_inst_pe_1_0_0_n105, npu_inst_pe_1_0_0_n104,
         npu_inst_pe_1_0_0_n103, npu_inst_pe_1_0_0_n102,
         npu_inst_pe_1_0_0_n101, npu_inst_pe_1_0_0_n100, npu_inst_pe_1_0_0_n99,
         npu_inst_pe_1_0_0_n98, npu_inst_pe_1_0_0_n36, npu_inst_pe_1_0_0_n35,
         npu_inst_pe_1_0_0_n34, npu_inst_pe_1_0_0_n33, npu_inst_pe_1_0_0_n32,
         npu_inst_pe_1_0_0_n31, npu_inst_pe_1_0_0_n30, npu_inst_pe_1_0_0_n29,
         npu_inst_pe_1_0_0_n28, npu_inst_pe_1_0_0_n25, npu_inst_pe_1_0_0_n24,
         npu_inst_pe_1_0_0_n23, npu_inst_pe_1_0_0_n22, npu_inst_pe_1_0_0_n21,
         npu_inst_pe_1_0_0_n20, npu_inst_pe_1_0_0_n19, npu_inst_pe_1_0_0_n18,
         npu_inst_pe_1_0_0_n17, npu_inst_pe_1_0_0_n16, npu_inst_pe_1_0_0_n15,
         npu_inst_pe_1_0_0_n14, npu_inst_pe_1_0_0_n13, npu_inst_pe_1_0_0_n12,
         npu_inst_pe_1_0_0_n11, npu_inst_pe_1_0_0_n10, npu_inst_pe_1_0_0_n9,
         npu_inst_pe_1_0_0_n8, npu_inst_pe_1_0_0_n7, npu_inst_pe_1_0_0_n6,
         npu_inst_pe_1_0_0_n5, npu_inst_pe_1_0_0_n4, npu_inst_pe_1_0_0_n3,
         npu_inst_pe_1_0_0_n2, npu_inst_pe_1_0_0_n1,
         npu_inst_pe_1_0_0_sub_67_carry_7_, npu_inst_pe_1_0_0_sub_67_carry_6_,
         npu_inst_pe_1_0_0_sub_67_carry_5_, npu_inst_pe_1_0_0_sub_67_carry_4_,
         npu_inst_pe_1_0_0_sub_67_carry_3_, npu_inst_pe_1_0_0_sub_67_carry_2_,
         npu_inst_pe_1_0_0_sub_67_carry_1_, npu_inst_pe_1_0_0_add_69_carry_7_,
         npu_inst_pe_1_0_0_add_69_carry_6_, npu_inst_pe_1_0_0_add_69_carry_5_,
         npu_inst_pe_1_0_0_add_69_carry_4_, npu_inst_pe_1_0_0_add_69_carry_3_,
         npu_inst_pe_1_0_0_add_69_carry_2_, npu_inst_pe_1_0_0_add_69_carry_1_,
         npu_inst_pe_1_0_0_n97, npu_inst_pe_1_0_0_n96, npu_inst_pe_1_0_0_n95,
         npu_inst_pe_1_0_0_n94, npu_inst_pe_1_0_0_n93, npu_inst_pe_1_0_0_n92,
         npu_inst_pe_1_0_0_n91, npu_inst_pe_1_0_0_n90, npu_inst_pe_1_0_0_n89,
         npu_inst_pe_1_0_0_n88, npu_inst_pe_1_0_0_n87, npu_inst_pe_1_0_0_n86,
         npu_inst_pe_1_0_0_n85, npu_inst_pe_1_0_0_n84, npu_inst_pe_1_0_0_n83,
         npu_inst_pe_1_0_0_n82, npu_inst_pe_1_0_0_n81, npu_inst_pe_1_0_0_n80,
         npu_inst_pe_1_0_0_n79, npu_inst_pe_1_0_0_n78, npu_inst_pe_1_0_0_n77,
         npu_inst_pe_1_0_0_n76, npu_inst_pe_1_0_0_n75, npu_inst_pe_1_0_0_n74,
         npu_inst_pe_1_0_0_n73, npu_inst_pe_1_0_0_n72, npu_inst_pe_1_0_0_n71,
         npu_inst_pe_1_0_0_n70, npu_inst_pe_1_0_0_n69, npu_inst_pe_1_0_0_n68,
         npu_inst_pe_1_0_0_n67, npu_inst_pe_1_0_0_n66, npu_inst_pe_1_0_0_n65,
         npu_inst_pe_1_0_0_n64, npu_inst_pe_1_0_0_n63, npu_inst_pe_1_0_0_n62,
         npu_inst_pe_1_0_0_n61, npu_inst_pe_1_0_0_n60, npu_inst_pe_1_0_0_n59,
         npu_inst_pe_1_0_0_n58, npu_inst_pe_1_0_0_n57, npu_inst_pe_1_0_0_n56,
         npu_inst_pe_1_0_0_n55, npu_inst_pe_1_0_0_n54, npu_inst_pe_1_0_0_n53,
         npu_inst_pe_1_0_0_n52, npu_inst_pe_1_0_0_n51, npu_inst_pe_1_0_0_n50,
         npu_inst_pe_1_0_0_n49, npu_inst_pe_1_0_0_n48, npu_inst_pe_1_0_0_n47,
         npu_inst_pe_1_0_0_n46, npu_inst_pe_1_0_0_n45, npu_inst_pe_1_0_0_n44,
         npu_inst_pe_1_0_0_n43, npu_inst_pe_1_0_0_n42, npu_inst_pe_1_0_0_n41,
         npu_inst_pe_1_0_0_n40, npu_inst_pe_1_0_0_n39, npu_inst_pe_1_0_0_n38,
         npu_inst_pe_1_0_0_n37, npu_inst_pe_1_0_0_n27, npu_inst_pe_1_0_0_n26,
         npu_inst_pe_1_0_0_net4568, npu_inst_pe_1_0_0_net4562,
         npu_inst_pe_1_0_0_N94, npu_inst_pe_1_0_0_N93, npu_inst_pe_1_0_0_N84,
         npu_inst_pe_1_0_0_N80, npu_inst_pe_1_0_0_N79, npu_inst_pe_1_0_0_N78,
         npu_inst_pe_1_0_0_N77, npu_inst_pe_1_0_0_N76, npu_inst_pe_1_0_0_N75,
         npu_inst_pe_1_0_0_N74, npu_inst_pe_1_0_0_N73, npu_inst_pe_1_0_0_N72,
         npu_inst_pe_1_0_0_N71, npu_inst_pe_1_0_0_N70, npu_inst_pe_1_0_0_N69,
         npu_inst_pe_1_0_0_N68, npu_inst_pe_1_0_0_N67, npu_inst_pe_1_0_0_N66,
         npu_inst_pe_1_0_0_N65, npu_inst_pe_1_0_0_int_q_acc_0_,
         npu_inst_pe_1_0_0_int_q_acc_1_, npu_inst_pe_1_0_0_int_q_acc_2_,
         npu_inst_pe_1_0_0_int_q_acc_3_, npu_inst_pe_1_0_0_int_q_acc_4_,
         npu_inst_pe_1_0_0_int_q_acc_5_, npu_inst_pe_1_0_0_int_q_acc_6_,
         npu_inst_pe_1_0_0_int_q_acc_7_, npu_inst_pe_1_0_0_int_data_0_,
         npu_inst_pe_1_0_0_int_data_1_, npu_inst_pe_1_0_0_int_q_weight_0_,
         npu_inst_pe_1_0_0_int_q_weight_1_,
         npu_inst_pe_1_0_0_int_q_reg_v_5__0_,
         npu_inst_pe_1_0_0_int_q_reg_v_5__1_,
         npu_inst_pe_1_0_0_int_q_reg_v_4__0_,
         npu_inst_pe_1_0_0_int_q_reg_v_4__1_,
         npu_inst_pe_1_0_0_int_q_reg_v_3__0_,
         npu_inst_pe_1_0_0_int_q_reg_v_3__1_,
         npu_inst_pe_1_0_0_int_q_reg_v_2__0_,
         npu_inst_pe_1_0_0_int_q_reg_v_2__1_,
         npu_inst_pe_1_0_0_int_q_reg_v_1__0_,
         npu_inst_pe_1_0_0_int_q_reg_v_1__1_,
         npu_inst_pe_1_0_0_int_q_reg_v_0__0_,
         npu_inst_pe_1_0_0_int_q_reg_v_0__1_,
         npu_inst_pe_1_0_0_int_q_reg_h_5__0_,
         npu_inst_pe_1_0_0_int_q_reg_h_5__1_,
         npu_inst_pe_1_0_0_int_q_reg_h_4__0_,
         npu_inst_pe_1_0_0_int_q_reg_h_4__1_,
         npu_inst_pe_1_0_0_int_q_reg_h_3__0_,
         npu_inst_pe_1_0_0_int_q_reg_h_3__1_,
         npu_inst_pe_1_0_0_int_q_reg_h_2__0_,
         npu_inst_pe_1_0_0_int_q_reg_h_2__1_,
         npu_inst_pe_1_0_0_int_q_reg_h_1__0_,
         npu_inst_pe_1_0_0_int_q_reg_h_1__1_,
         npu_inst_pe_1_0_0_int_q_reg_h_0__0_,
         npu_inst_pe_1_0_0_int_q_reg_h_0__1_, npu_inst_pe_1_0_0_o_data_v_0_,
         npu_inst_pe_1_0_0_o_data_v_1_, npu_inst_pe_1_0_0_o_data_h_0_,
         npu_inst_pe_1_0_0_o_data_h_1_, npu_inst_pe_1_0_1_n117,
         npu_inst_pe_1_0_1_n116, npu_inst_pe_1_0_1_n115,
         npu_inst_pe_1_0_1_n114, npu_inst_pe_1_0_1_n113,
         npu_inst_pe_1_0_1_n112, npu_inst_pe_1_0_1_n111,
         npu_inst_pe_1_0_1_n110, npu_inst_pe_1_0_1_n109,
         npu_inst_pe_1_0_1_n108, npu_inst_pe_1_0_1_n107,
         npu_inst_pe_1_0_1_n106, npu_inst_pe_1_0_1_n105,
         npu_inst_pe_1_0_1_n104, npu_inst_pe_1_0_1_n103,
         npu_inst_pe_1_0_1_n102, npu_inst_pe_1_0_1_n101,
         npu_inst_pe_1_0_1_n100, npu_inst_pe_1_0_1_n99, npu_inst_pe_1_0_1_n98,
         npu_inst_pe_1_0_1_n36, npu_inst_pe_1_0_1_n35, npu_inst_pe_1_0_1_n34,
         npu_inst_pe_1_0_1_n33, npu_inst_pe_1_0_1_n32, npu_inst_pe_1_0_1_n31,
         npu_inst_pe_1_0_1_n30, npu_inst_pe_1_0_1_n29, npu_inst_pe_1_0_1_n28,
         npu_inst_pe_1_0_1_n25, npu_inst_pe_1_0_1_n24, npu_inst_pe_1_0_1_n23,
         npu_inst_pe_1_0_1_n22, npu_inst_pe_1_0_1_n21, npu_inst_pe_1_0_1_n20,
         npu_inst_pe_1_0_1_n19, npu_inst_pe_1_0_1_n18, npu_inst_pe_1_0_1_n17,
         npu_inst_pe_1_0_1_n16, npu_inst_pe_1_0_1_n15, npu_inst_pe_1_0_1_n14,
         npu_inst_pe_1_0_1_n13, npu_inst_pe_1_0_1_n12, npu_inst_pe_1_0_1_n11,
         npu_inst_pe_1_0_1_n10, npu_inst_pe_1_0_1_n9, npu_inst_pe_1_0_1_n8,
         npu_inst_pe_1_0_1_n7, npu_inst_pe_1_0_1_n6, npu_inst_pe_1_0_1_n5,
         npu_inst_pe_1_0_1_n4, npu_inst_pe_1_0_1_n3, npu_inst_pe_1_0_1_n2,
         npu_inst_pe_1_0_1_n1, npu_inst_pe_1_0_1_sub_67_carry_7_,
         npu_inst_pe_1_0_1_sub_67_carry_6_, npu_inst_pe_1_0_1_sub_67_carry_5_,
         npu_inst_pe_1_0_1_sub_67_carry_4_, npu_inst_pe_1_0_1_sub_67_carry_3_,
         npu_inst_pe_1_0_1_sub_67_carry_2_, npu_inst_pe_1_0_1_sub_67_carry_1_,
         npu_inst_pe_1_0_1_add_69_carry_7_, npu_inst_pe_1_0_1_add_69_carry_6_,
         npu_inst_pe_1_0_1_add_69_carry_5_, npu_inst_pe_1_0_1_add_69_carry_4_,
         npu_inst_pe_1_0_1_add_69_carry_3_, npu_inst_pe_1_0_1_add_69_carry_2_,
         npu_inst_pe_1_0_1_add_69_carry_1_, npu_inst_pe_1_0_1_n97,
         npu_inst_pe_1_0_1_n96, npu_inst_pe_1_0_1_n95, npu_inst_pe_1_0_1_n94,
         npu_inst_pe_1_0_1_n93, npu_inst_pe_1_0_1_n92, npu_inst_pe_1_0_1_n91,
         npu_inst_pe_1_0_1_n90, npu_inst_pe_1_0_1_n89, npu_inst_pe_1_0_1_n88,
         npu_inst_pe_1_0_1_n87, npu_inst_pe_1_0_1_n86, npu_inst_pe_1_0_1_n85,
         npu_inst_pe_1_0_1_n84, npu_inst_pe_1_0_1_n83, npu_inst_pe_1_0_1_n82,
         npu_inst_pe_1_0_1_n81, npu_inst_pe_1_0_1_n80, npu_inst_pe_1_0_1_n79,
         npu_inst_pe_1_0_1_n78, npu_inst_pe_1_0_1_n77, npu_inst_pe_1_0_1_n76,
         npu_inst_pe_1_0_1_n75, npu_inst_pe_1_0_1_n74, npu_inst_pe_1_0_1_n73,
         npu_inst_pe_1_0_1_n72, npu_inst_pe_1_0_1_n71, npu_inst_pe_1_0_1_n70,
         npu_inst_pe_1_0_1_n69, npu_inst_pe_1_0_1_n68, npu_inst_pe_1_0_1_n67,
         npu_inst_pe_1_0_1_n66, npu_inst_pe_1_0_1_n65, npu_inst_pe_1_0_1_n64,
         npu_inst_pe_1_0_1_n63, npu_inst_pe_1_0_1_n62, npu_inst_pe_1_0_1_n61,
         npu_inst_pe_1_0_1_n60, npu_inst_pe_1_0_1_n59, npu_inst_pe_1_0_1_n58,
         npu_inst_pe_1_0_1_n57, npu_inst_pe_1_0_1_n56, npu_inst_pe_1_0_1_n55,
         npu_inst_pe_1_0_1_n54, npu_inst_pe_1_0_1_n53, npu_inst_pe_1_0_1_n52,
         npu_inst_pe_1_0_1_n51, npu_inst_pe_1_0_1_n50, npu_inst_pe_1_0_1_n49,
         npu_inst_pe_1_0_1_n48, npu_inst_pe_1_0_1_n47, npu_inst_pe_1_0_1_n46,
         npu_inst_pe_1_0_1_n45, npu_inst_pe_1_0_1_n44, npu_inst_pe_1_0_1_n43,
         npu_inst_pe_1_0_1_n42, npu_inst_pe_1_0_1_n41, npu_inst_pe_1_0_1_n40,
         npu_inst_pe_1_0_1_n39, npu_inst_pe_1_0_1_n38, npu_inst_pe_1_0_1_n37,
         npu_inst_pe_1_0_1_n27, npu_inst_pe_1_0_1_n26,
         npu_inst_pe_1_0_1_net4545, npu_inst_pe_1_0_1_net4539,
         npu_inst_pe_1_0_1_N94, npu_inst_pe_1_0_1_N93, npu_inst_pe_1_0_1_N84,
         npu_inst_pe_1_0_1_N80, npu_inst_pe_1_0_1_N79, npu_inst_pe_1_0_1_N78,
         npu_inst_pe_1_0_1_N77, npu_inst_pe_1_0_1_N76, npu_inst_pe_1_0_1_N75,
         npu_inst_pe_1_0_1_N74, npu_inst_pe_1_0_1_N73, npu_inst_pe_1_0_1_N72,
         npu_inst_pe_1_0_1_N71, npu_inst_pe_1_0_1_N70, npu_inst_pe_1_0_1_N69,
         npu_inst_pe_1_0_1_N68, npu_inst_pe_1_0_1_N67, npu_inst_pe_1_0_1_N66,
         npu_inst_pe_1_0_1_N65, npu_inst_pe_1_0_1_int_q_acc_0_,
         npu_inst_pe_1_0_1_int_q_acc_1_, npu_inst_pe_1_0_1_int_q_acc_2_,
         npu_inst_pe_1_0_1_int_q_acc_3_, npu_inst_pe_1_0_1_int_q_acc_4_,
         npu_inst_pe_1_0_1_int_q_acc_5_, npu_inst_pe_1_0_1_int_q_acc_6_,
         npu_inst_pe_1_0_1_int_q_acc_7_, npu_inst_pe_1_0_1_int_data_0_,
         npu_inst_pe_1_0_1_int_data_1_, npu_inst_pe_1_0_1_int_q_weight_0_,
         npu_inst_pe_1_0_1_int_q_weight_1_,
         npu_inst_pe_1_0_1_int_q_reg_v_5__0_,
         npu_inst_pe_1_0_1_int_q_reg_v_5__1_,
         npu_inst_pe_1_0_1_int_q_reg_v_4__0_,
         npu_inst_pe_1_0_1_int_q_reg_v_4__1_,
         npu_inst_pe_1_0_1_int_q_reg_v_3__0_,
         npu_inst_pe_1_0_1_int_q_reg_v_3__1_,
         npu_inst_pe_1_0_1_int_q_reg_v_2__0_,
         npu_inst_pe_1_0_1_int_q_reg_v_2__1_,
         npu_inst_pe_1_0_1_int_q_reg_v_1__0_,
         npu_inst_pe_1_0_1_int_q_reg_v_1__1_,
         npu_inst_pe_1_0_1_int_q_reg_v_0__0_,
         npu_inst_pe_1_0_1_int_q_reg_v_0__1_,
         npu_inst_pe_1_0_1_int_q_reg_h_5__0_,
         npu_inst_pe_1_0_1_int_q_reg_h_5__1_,
         npu_inst_pe_1_0_1_int_q_reg_h_4__0_,
         npu_inst_pe_1_0_1_int_q_reg_h_4__1_,
         npu_inst_pe_1_0_1_int_q_reg_h_3__0_,
         npu_inst_pe_1_0_1_int_q_reg_h_3__1_,
         npu_inst_pe_1_0_1_int_q_reg_h_2__0_,
         npu_inst_pe_1_0_1_int_q_reg_h_2__1_,
         npu_inst_pe_1_0_1_int_q_reg_h_1__0_,
         npu_inst_pe_1_0_1_int_q_reg_h_1__1_,
         npu_inst_pe_1_0_1_int_q_reg_h_0__0_,
         npu_inst_pe_1_0_1_int_q_reg_h_0__1_, npu_inst_pe_1_0_1_o_data_v_0_,
         npu_inst_pe_1_0_1_o_data_v_1_, npu_inst_pe_1_0_2_n118,
         npu_inst_pe_1_0_2_n117, npu_inst_pe_1_0_2_n116,
         npu_inst_pe_1_0_2_n115, npu_inst_pe_1_0_2_n114,
         npu_inst_pe_1_0_2_n113, npu_inst_pe_1_0_2_n112,
         npu_inst_pe_1_0_2_n111, npu_inst_pe_1_0_2_n110,
         npu_inst_pe_1_0_2_n109, npu_inst_pe_1_0_2_n108,
         npu_inst_pe_1_0_2_n107, npu_inst_pe_1_0_2_n106,
         npu_inst_pe_1_0_2_n105, npu_inst_pe_1_0_2_n104,
         npu_inst_pe_1_0_2_n103, npu_inst_pe_1_0_2_n102,
         npu_inst_pe_1_0_2_n101, npu_inst_pe_1_0_2_n100, npu_inst_pe_1_0_2_n99,
         npu_inst_pe_1_0_2_n98, npu_inst_pe_1_0_2_n36, npu_inst_pe_1_0_2_n35,
         npu_inst_pe_1_0_2_n34, npu_inst_pe_1_0_2_n33, npu_inst_pe_1_0_2_n32,
         npu_inst_pe_1_0_2_n31, npu_inst_pe_1_0_2_n30, npu_inst_pe_1_0_2_n29,
         npu_inst_pe_1_0_2_n28, npu_inst_pe_1_0_2_n25, npu_inst_pe_1_0_2_n24,
         npu_inst_pe_1_0_2_n23, npu_inst_pe_1_0_2_n22, npu_inst_pe_1_0_2_n21,
         npu_inst_pe_1_0_2_n20, npu_inst_pe_1_0_2_n19, npu_inst_pe_1_0_2_n18,
         npu_inst_pe_1_0_2_n17, npu_inst_pe_1_0_2_n16, npu_inst_pe_1_0_2_n15,
         npu_inst_pe_1_0_2_n14, npu_inst_pe_1_0_2_n13, npu_inst_pe_1_0_2_n12,
         npu_inst_pe_1_0_2_n11, npu_inst_pe_1_0_2_n10, npu_inst_pe_1_0_2_n9,
         npu_inst_pe_1_0_2_n8, npu_inst_pe_1_0_2_n7, npu_inst_pe_1_0_2_n6,
         npu_inst_pe_1_0_2_n5, npu_inst_pe_1_0_2_n4, npu_inst_pe_1_0_2_n3,
         npu_inst_pe_1_0_2_n2, npu_inst_pe_1_0_2_n1,
         npu_inst_pe_1_0_2_sub_67_carry_7_, npu_inst_pe_1_0_2_sub_67_carry_6_,
         npu_inst_pe_1_0_2_sub_67_carry_5_, npu_inst_pe_1_0_2_sub_67_carry_4_,
         npu_inst_pe_1_0_2_sub_67_carry_3_, npu_inst_pe_1_0_2_sub_67_carry_2_,
         npu_inst_pe_1_0_2_sub_67_carry_1_, npu_inst_pe_1_0_2_add_69_carry_7_,
         npu_inst_pe_1_0_2_add_69_carry_6_, npu_inst_pe_1_0_2_add_69_carry_5_,
         npu_inst_pe_1_0_2_add_69_carry_4_, npu_inst_pe_1_0_2_add_69_carry_3_,
         npu_inst_pe_1_0_2_add_69_carry_2_, npu_inst_pe_1_0_2_add_69_carry_1_,
         npu_inst_pe_1_0_2_n97, npu_inst_pe_1_0_2_n96, npu_inst_pe_1_0_2_n95,
         npu_inst_pe_1_0_2_n94, npu_inst_pe_1_0_2_n93, npu_inst_pe_1_0_2_n92,
         npu_inst_pe_1_0_2_n91, npu_inst_pe_1_0_2_n90, npu_inst_pe_1_0_2_n89,
         npu_inst_pe_1_0_2_n88, npu_inst_pe_1_0_2_n87, npu_inst_pe_1_0_2_n86,
         npu_inst_pe_1_0_2_n85, npu_inst_pe_1_0_2_n84, npu_inst_pe_1_0_2_n83,
         npu_inst_pe_1_0_2_n82, npu_inst_pe_1_0_2_n81, npu_inst_pe_1_0_2_n80,
         npu_inst_pe_1_0_2_n79, npu_inst_pe_1_0_2_n78, npu_inst_pe_1_0_2_n77,
         npu_inst_pe_1_0_2_n76, npu_inst_pe_1_0_2_n75, npu_inst_pe_1_0_2_n74,
         npu_inst_pe_1_0_2_n73, npu_inst_pe_1_0_2_n72, npu_inst_pe_1_0_2_n71,
         npu_inst_pe_1_0_2_n70, npu_inst_pe_1_0_2_n69, npu_inst_pe_1_0_2_n68,
         npu_inst_pe_1_0_2_n67, npu_inst_pe_1_0_2_n66, npu_inst_pe_1_0_2_n65,
         npu_inst_pe_1_0_2_n64, npu_inst_pe_1_0_2_n63, npu_inst_pe_1_0_2_n62,
         npu_inst_pe_1_0_2_n61, npu_inst_pe_1_0_2_n60, npu_inst_pe_1_0_2_n59,
         npu_inst_pe_1_0_2_n58, npu_inst_pe_1_0_2_n57, npu_inst_pe_1_0_2_n56,
         npu_inst_pe_1_0_2_n55, npu_inst_pe_1_0_2_n54, npu_inst_pe_1_0_2_n53,
         npu_inst_pe_1_0_2_n52, npu_inst_pe_1_0_2_n51, npu_inst_pe_1_0_2_n50,
         npu_inst_pe_1_0_2_n49, npu_inst_pe_1_0_2_n48, npu_inst_pe_1_0_2_n47,
         npu_inst_pe_1_0_2_n46, npu_inst_pe_1_0_2_n45, npu_inst_pe_1_0_2_n44,
         npu_inst_pe_1_0_2_n43, npu_inst_pe_1_0_2_n42, npu_inst_pe_1_0_2_n41,
         npu_inst_pe_1_0_2_n40, npu_inst_pe_1_0_2_n39, npu_inst_pe_1_0_2_n38,
         npu_inst_pe_1_0_2_n37, npu_inst_pe_1_0_2_n27, npu_inst_pe_1_0_2_n26,
         npu_inst_pe_1_0_2_net4522, npu_inst_pe_1_0_2_net4516,
         npu_inst_pe_1_0_2_N94, npu_inst_pe_1_0_2_N93, npu_inst_pe_1_0_2_N84,
         npu_inst_pe_1_0_2_N80, npu_inst_pe_1_0_2_N79, npu_inst_pe_1_0_2_N78,
         npu_inst_pe_1_0_2_N77, npu_inst_pe_1_0_2_N76, npu_inst_pe_1_0_2_N75,
         npu_inst_pe_1_0_2_N74, npu_inst_pe_1_0_2_N73, npu_inst_pe_1_0_2_N72,
         npu_inst_pe_1_0_2_N71, npu_inst_pe_1_0_2_N70, npu_inst_pe_1_0_2_N69,
         npu_inst_pe_1_0_2_N68, npu_inst_pe_1_0_2_N67, npu_inst_pe_1_0_2_N66,
         npu_inst_pe_1_0_2_N65, npu_inst_pe_1_0_2_int_q_acc_0_,
         npu_inst_pe_1_0_2_int_q_acc_1_, npu_inst_pe_1_0_2_int_q_acc_2_,
         npu_inst_pe_1_0_2_int_q_acc_3_, npu_inst_pe_1_0_2_int_q_acc_4_,
         npu_inst_pe_1_0_2_int_q_acc_5_, npu_inst_pe_1_0_2_int_q_acc_6_,
         npu_inst_pe_1_0_2_int_q_acc_7_, npu_inst_pe_1_0_2_int_data_0_,
         npu_inst_pe_1_0_2_int_data_1_, npu_inst_pe_1_0_2_int_q_weight_0_,
         npu_inst_pe_1_0_2_int_q_weight_1_,
         npu_inst_pe_1_0_2_int_q_reg_v_5__0_,
         npu_inst_pe_1_0_2_int_q_reg_v_5__1_,
         npu_inst_pe_1_0_2_int_q_reg_v_4__0_,
         npu_inst_pe_1_0_2_int_q_reg_v_4__1_,
         npu_inst_pe_1_0_2_int_q_reg_v_3__0_,
         npu_inst_pe_1_0_2_int_q_reg_v_3__1_,
         npu_inst_pe_1_0_2_int_q_reg_v_2__0_,
         npu_inst_pe_1_0_2_int_q_reg_v_2__1_,
         npu_inst_pe_1_0_2_int_q_reg_v_1__0_,
         npu_inst_pe_1_0_2_int_q_reg_v_1__1_,
         npu_inst_pe_1_0_2_int_q_reg_v_0__0_,
         npu_inst_pe_1_0_2_int_q_reg_v_0__1_,
         npu_inst_pe_1_0_2_int_q_reg_h_5__0_,
         npu_inst_pe_1_0_2_int_q_reg_h_5__1_,
         npu_inst_pe_1_0_2_int_q_reg_h_4__0_,
         npu_inst_pe_1_0_2_int_q_reg_h_4__1_,
         npu_inst_pe_1_0_2_int_q_reg_h_3__0_,
         npu_inst_pe_1_0_2_int_q_reg_h_3__1_,
         npu_inst_pe_1_0_2_int_q_reg_h_2__0_,
         npu_inst_pe_1_0_2_int_q_reg_h_2__1_,
         npu_inst_pe_1_0_2_int_q_reg_h_1__0_,
         npu_inst_pe_1_0_2_int_q_reg_h_1__1_,
         npu_inst_pe_1_0_2_int_q_reg_h_0__0_,
         npu_inst_pe_1_0_2_int_q_reg_h_0__1_, npu_inst_pe_1_0_2_o_data_v_0_,
         npu_inst_pe_1_0_2_o_data_v_1_, npu_inst_pe_1_0_3_n119,
         npu_inst_pe_1_0_3_n118, npu_inst_pe_1_0_3_n117,
         npu_inst_pe_1_0_3_n116, npu_inst_pe_1_0_3_n115,
         npu_inst_pe_1_0_3_n114, npu_inst_pe_1_0_3_n113,
         npu_inst_pe_1_0_3_n112, npu_inst_pe_1_0_3_n111,
         npu_inst_pe_1_0_3_n110, npu_inst_pe_1_0_3_n109,
         npu_inst_pe_1_0_3_n108, npu_inst_pe_1_0_3_n107,
         npu_inst_pe_1_0_3_n106, npu_inst_pe_1_0_3_n105,
         npu_inst_pe_1_0_3_n104, npu_inst_pe_1_0_3_n103,
         npu_inst_pe_1_0_3_n102, npu_inst_pe_1_0_3_n101,
         npu_inst_pe_1_0_3_n100, npu_inst_pe_1_0_3_n99, npu_inst_pe_1_0_3_n98,
         npu_inst_pe_1_0_3_n36, npu_inst_pe_1_0_3_n35, npu_inst_pe_1_0_3_n34,
         npu_inst_pe_1_0_3_n33, npu_inst_pe_1_0_3_n32, npu_inst_pe_1_0_3_n31,
         npu_inst_pe_1_0_3_n30, npu_inst_pe_1_0_3_n29, npu_inst_pe_1_0_3_n28,
         npu_inst_pe_1_0_3_n25, npu_inst_pe_1_0_3_n24, npu_inst_pe_1_0_3_n23,
         npu_inst_pe_1_0_3_n22, npu_inst_pe_1_0_3_n21, npu_inst_pe_1_0_3_n20,
         npu_inst_pe_1_0_3_n19, npu_inst_pe_1_0_3_n18, npu_inst_pe_1_0_3_n17,
         npu_inst_pe_1_0_3_n16, npu_inst_pe_1_0_3_n15, npu_inst_pe_1_0_3_n14,
         npu_inst_pe_1_0_3_n13, npu_inst_pe_1_0_3_n12, npu_inst_pe_1_0_3_n11,
         npu_inst_pe_1_0_3_n10, npu_inst_pe_1_0_3_n9, npu_inst_pe_1_0_3_n8,
         npu_inst_pe_1_0_3_n7, npu_inst_pe_1_0_3_n6, npu_inst_pe_1_0_3_n5,
         npu_inst_pe_1_0_3_n4, npu_inst_pe_1_0_3_n3, npu_inst_pe_1_0_3_n2,
         npu_inst_pe_1_0_3_n1, npu_inst_pe_1_0_3_sub_67_carry_7_,
         npu_inst_pe_1_0_3_sub_67_carry_6_, npu_inst_pe_1_0_3_sub_67_carry_5_,
         npu_inst_pe_1_0_3_sub_67_carry_4_, npu_inst_pe_1_0_3_sub_67_carry_3_,
         npu_inst_pe_1_0_3_sub_67_carry_2_, npu_inst_pe_1_0_3_sub_67_carry_1_,
         npu_inst_pe_1_0_3_add_69_carry_7_, npu_inst_pe_1_0_3_add_69_carry_6_,
         npu_inst_pe_1_0_3_add_69_carry_5_, npu_inst_pe_1_0_3_add_69_carry_4_,
         npu_inst_pe_1_0_3_add_69_carry_3_, npu_inst_pe_1_0_3_add_69_carry_2_,
         npu_inst_pe_1_0_3_add_69_carry_1_, npu_inst_pe_1_0_3_n97,
         npu_inst_pe_1_0_3_n96, npu_inst_pe_1_0_3_n95, npu_inst_pe_1_0_3_n94,
         npu_inst_pe_1_0_3_n93, npu_inst_pe_1_0_3_n92, npu_inst_pe_1_0_3_n91,
         npu_inst_pe_1_0_3_n90, npu_inst_pe_1_0_3_n89, npu_inst_pe_1_0_3_n88,
         npu_inst_pe_1_0_3_n87, npu_inst_pe_1_0_3_n86, npu_inst_pe_1_0_3_n85,
         npu_inst_pe_1_0_3_n84, npu_inst_pe_1_0_3_n83, npu_inst_pe_1_0_3_n82,
         npu_inst_pe_1_0_3_n81, npu_inst_pe_1_0_3_n80, npu_inst_pe_1_0_3_n79,
         npu_inst_pe_1_0_3_n78, npu_inst_pe_1_0_3_n77, npu_inst_pe_1_0_3_n76,
         npu_inst_pe_1_0_3_n75, npu_inst_pe_1_0_3_n74, npu_inst_pe_1_0_3_n73,
         npu_inst_pe_1_0_3_n72, npu_inst_pe_1_0_3_n71, npu_inst_pe_1_0_3_n70,
         npu_inst_pe_1_0_3_n69, npu_inst_pe_1_0_3_n68, npu_inst_pe_1_0_3_n67,
         npu_inst_pe_1_0_3_n66, npu_inst_pe_1_0_3_n65, npu_inst_pe_1_0_3_n64,
         npu_inst_pe_1_0_3_n63, npu_inst_pe_1_0_3_n62, npu_inst_pe_1_0_3_n61,
         npu_inst_pe_1_0_3_n60, npu_inst_pe_1_0_3_n59, npu_inst_pe_1_0_3_n58,
         npu_inst_pe_1_0_3_n57, npu_inst_pe_1_0_3_n56, npu_inst_pe_1_0_3_n55,
         npu_inst_pe_1_0_3_n54, npu_inst_pe_1_0_3_n53, npu_inst_pe_1_0_3_n52,
         npu_inst_pe_1_0_3_n51, npu_inst_pe_1_0_3_n50, npu_inst_pe_1_0_3_n49,
         npu_inst_pe_1_0_3_n48, npu_inst_pe_1_0_3_n47, npu_inst_pe_1_0_3_n46,
         npu_inst_pe_1_0_3_n45, npu_inst_pe_1_0_3_n44, npu_inst_pe_1_0_3_n43,
         npu_inst_pe_1_0_3_n42, npu_inst_pe_1_0_3_n41, npu_inst_pe_1_0_3_n40,
         npu_inst_pe_1_0_3_n39, npu_inst_pe_1_0_3_n38, npu_inst_pe_1_0_3_n37,
         npu_inst_pe_1_0_3_n27, npu_inst_pe_1_0_3_n26,
         npu_inst_pe_1_0_3_net4499, npu_inst_pe_1_0_3_net4493,
         npu_inst_pe_1_0_3_N94, npu_inst_pe_1_0_3_N93, npu_inst_pe_1_0_3_N84,
         npu_inst_pe_1_0_3_N80, npu_inst_pe_1_0_3_N79, npu_inst_pe_1_0_3_N78,
         npu_inst_pe_1_0_3_N77, npu_inst_pe_1_0_3_N76, npu_inst_pe_1_0_3_N75,
         npu_inst_pe_1_0_3_N74, npu_inst_pe_1_0_3_N73, npu_inst_pe_1_0_3_N72,
         npu_inst_pe_1_0_3_N71, npu_inst_pe_1_0_3_N70, npu_inst_pe_1_0_3_N69,
         npu_inst_pe_1_0_3_N68, npu_inst_pe_1_0_3_N67, npu_inst_pe_1_0_3_N66,
         npu_inst_pe_1_0_3_N65, npu_inst_pe_1_0_3_int_q_acc_0_,
         npu_inst_pe_1_0_3_int_q_acc_1_, npu_inst_pe_1_0_3_int_q_acc_2_,
         npu_inst_pe_1_0_3_int_q_acc_3_, npu_inst_pe_1_0_3_int_q_acc_4_,
         npu_inst_pe_1_0_3_int_q_acc_5_, npu_inst_pe_1_0_3_int_q_acc_6_,
         npu_inst_pe_1_0_3_int_q_acc_7_, npu_inst_pe_1_0_3_int_data_0_,
         npu_inst_pe_1_0_3_int_data_1_, npu_inst_pe_1_0_3_int_q_weight_0_,
         npu_inst_pe_1_0_3_int_q_weight_1_,
         npu_inst_pe_1_0_3_int_q_reg_v_5__0_,
         npu_inst_pe_1_0_3_int_q_reg_v_5__1_,
         npu_inst_pe_1_0_3_int_q_reg_v_4__0_,
         npu_inst_pe_1_0_3_int_q_reg_v_4__1_,
         npu_inst_pe_1_0_3_int_q_reg_v_3__0_,
         npu_inst_pe_1_0_3_int_q_reg_v_3__1_,
         npu_inst_pe_1_0_3_int_q_reg_v_2__0_,
         npu_inst_pe_1_0_3_int_q_reg_v_2__1_,
         npu_inst_pe_1_0_3_int_q_reg_v_1__0_,
         npu_inst_pe_1_0_3_int_q_reg_v_1__1_,
         npu_inst_pe_1_0_3_int_q_reg_v_0__0_,
         npu_inst_pe_1_0_3_int_q_reg_v_0__1_,
         npu_inst_pe_1_0_3_int_q_reg_h_5__0_,
         npu_inst_pe_1_0_3_int_q_reg_h_5__1_,
         npu_inst_pe_1_0_3_int_q_reg_h_4__0_,
         npu_inst_pe_1_0_3_int_q_reg_h_4__1_,
         npu_inst_pe_1_0_3_int_q_reg_h_3__0_,
         npu_inst_pe_1_0_3_int_q_reg_h_3__1_,
         npu_inst_pe_1_0_3_int_q_reg_h_2__0_,
         npu_inst_pe_1_0_3_int_q_reg_h_2__1_,
         npu_inst_pe_1_0_3_int_q_reg_h_1__0_,
         npu_inst_pe_1_0_3_int_q_reg_h_1__1_,
         npu_inst_pe_1_0_3_int_q_reg_h_0__0_,
         npu_inst_pe_1_0_3_int_q_reg_h_0__1_, npu_inst_pe_1_0_3_o_data_v_0_,
         npu_inst_pe_1_0_3_o_data_v_1_, npu_inst_pe_1_0_4_n118,
         npu_inst_pe_1_0_4_n117, npu_inst_pe_1_0_4_n116,
         npu_inst_pe_1_0_4_n115, npu_inst_pe_1_0_4_n114,
         npu_inst_pe_1_0_4_n113, npu_inst_pe_1_0_4_n112,
         npu_inst_pe_1_0_4_n111, npu_inst_pe_1_0_4_n110,
         npu_inst_pe_1_0_4_n109, npu_inst_pe_1_0_4_n108,
         npu_inst_pe_1_0_4_n107, npu_inst_pe_1_0_4_n106,
         npu_inst_pe_1_0_4_n105, npu_inst_pe_1_0_4_n104,
         npu_inst_pe_1_0_4_n103, npu_inst_pe_1_0_4_n102,
         npu_inst_pe_1_0_4_n101, npu_inst_pe_1_0_4_n100, npu_inst_pe_1_0_4_n99,
         npu_inst_pe_1_0_4_n98, npu_inst_pe_1_0_4_n36, npu_inst_pe_1_0_4_n35,
         npu_inst_pe_1_0_4_n34, npu_inst_pe_1_0_4_n33, npu_inst_pe_1_0_4_n32,
         npu_inst_pe_1_0_4_n31, npu_inst_pe_1_0_4_n30, npu_inst_pe_1_0_4_n29,
         npu_inst_pe_1_0_4_n28, npu_inst_pe_1_0_4_n25, npu_inst_pe_1_0_4_n24,
         npu_inst_pe_1_0_4_n23, npu_inst_pe_1_0_4_n22, npu_inst_pe_1_0_4_n21,
         npu_inst_pe_1_0_4_n20, npu_inst_pe_1_0_4_n19, npu_inst_pe_1_0_4_n18,
         npu_inst_pe_1_0_4_n17, npu_inst_pe_1_0_4_n16, npu_inst_pe_1_0_4_n15,
         npu_inst_pe_1_0_4_n14, npu_inst_pe_1_0_4_n13, npu_inst_pe_1_0_4_n12,
         npu_inst_pe_1_0_4_n11, npu_inst_pe_1_0_4_n10, npu_inst_pe_1_0_4_n9,
         npu_inst_pe_1_0_4_n8, npu_inst_pe_1_0_4_n7, npu_inst_pe_1_0_4_n6,
         npu_inst_pe_1_0_4_n5, npu_inst_pe_1_0_4_n4, npu_inst_pe_1_0_4_n3,
         npu_inst_pe_1_0_4_n2, npu_inst_pe_1_0_4_n1,
         npu_inst_pe_1_0_4_sub_67_carry_7_, npu_inst_pe_1_0_4_sub_67_carry_6_,
         npu_inst_pe_1_0_4_sub_67_carry_5_, npu_inst_pe_1_0_4_sub_67_carry_4_,
         npu_inst_pe_1_0_4_sub_67_carry_3_, npu_inst_pe_1_0_4_sub_67_carry_2_,
         npu_inst_pe_1_0_4_sub_67_carry_1_, npu_inst_pe_1_0_4_add_69_carry_7_,
         npu_inst_pe_1_0_4_add_69_carry_6_, npu_inst_pe_1_0_4_add_69_carry_5_,
         npu_inst_pe_1_0_4_add_69_carry_4_, npu_inst_pe_1_0_4_add_69_carry_3_,
         npu_inst_pe_1_0_4_add_69_carry_2_, npu_inst_pe_1_0_4_add_69_carry_1_,
         npu_inst_pe_1_0_4_n97, npu_inst_pe_1_0_4_n96, npu_inst_pe_1_0_4_n95,
         npu_inst_pe_1_0_4_n94, npu_inst_pe_1_0_4_n93, npu_inst_pe_1_0_4_n92,
         npu_inst_pe_1_0_4_n91, npu_inst_pe_1_0_4_n90, npu_inst_pe_1_0_4_n89,
         npu_inst_pe_1_0_4_n88, npu_inst_pe_1_0_4_n87, npu_inst_pe_1_0_4_n86,
         npu_inst_pe_1_0_4_n85, npu_inst_pe_1_0_4_n84, npu_inst_pe_1_0_4_n83,
         npu_inst_pe_1_0_4_n82, npu_inst_pe_1_0_4_n81, npu_inst_pe_1_0_4_n80,
         npu_inst_pe_1_0_4_n79, npu_inst_pe_1_0_4_n78, npu_inst_pe_1_0_4_n77,
         npu_inst_pe_1_0_4_n76, npu_inst_pe_1_0_4_n75, npu_inst_pe_1_0_4_n74,
         npu_inst_pe_1_0_4_n73, npu_inst_pe_1_0_4_n72, npu_inst_pe_1_0_4_n71,
         npu_inst_pe_1_0_4_n70, npu_inst_pe_1_0_4_n69, npu_inst_pe_1_0_4_n68,
         npu_inst_pe_1_0_4_n67, npu_inst_pe_1_0_4_n66, npu_inst_pe_1_0_4_n65,
         npu_inst_pe_1_0_4_n64, npu_inst_pe_1_0_4_n63, npu_inst_pe_1_0_4_n62,
         npu_inst_pe_1_0_4_n61, npu_inst_pe_1_0_4_n60, npu_inst_pe_1_0_4_n59,
         npu_inst_pe_1_0_4_n58, npu_inst_pe_1_0_4_n57, npu_inst_pe_1_0_4_n56,
         npu_inst_pe_1_0_4_n55, npu_inst_pe_1_0_4_n54, npu_inst_pe_1_0_4_n53,
         npu_inst_pe_1_0_4_n52, npu_inst_pe_1_0_4_n51, npu_inst_pe_1_0_4_n50,
         npu_inst_pe_1_0_4_n49, npu_inst_pe_1_0_4_n48, npu_inst_pe_1_0_4_n47,
         npu_inst_pe_1_0_4_n46, npu_inst_pe_1_0_4_n45, npu_inst_pe_1_0_4_n44,
         npu_inst_pe_1_0_4_n43, npu_inst_pe_1_0_4_n42, npu_inst_pe_1_0_4_n41,
         npu_inst_pe_1_0_4_n40, npu_inst_pe_1_0_4_n39, npu_inst_pe_1_0_4_n38,
         npu_inst_pe_1_0_4_n37, npu_inst_pe_1_0_4_n27, npu_inst_pe_1_0_4_n26,
         npu_inst_pe_1_0_4_net4476, npu_inst_pe_1_0_4_net4470,
         npu_inst_pe_1_0_4_N94, npu_inst_pe_1_0_4_N93, npu_inst_pe_1_0_4_N84,
         npu_inst_pe_1_0_4_N80, npu_inst_pe_1_0_4_N79, npu_inst_pe_1_0_4_N78,
         npu_inst_pe_1_0_4_N77, npu_inst_pe_1_0_4_N76, npu_inst_pe_1_0_4_N75,
         npu_inst_pe_1_0_4_N74, npu_inst_pe_1_0_4_N73, npu_inst_pe_1_0_4_N72,
         npu_inst_pe_1_0_4_N71, npu_inst_pe_1_0_4_N70, npu_inst_pe_1_0_4_N69,
         npu_inst_pe_1_0_4_N68, npu_inst_pe_1_0_4_N67, npu_inst_pe_1_0_4_N66,
         npu_inst_pe_1_0_4_N65, npu_inst_pe_1_0_4_int_q_acc_0_,
         npu_inst_pe_1_0_4_int_q_acc_1_, npu_inst_pe_1_0_4_int_q_acc_2_,
         npu_inst_pe_1_0_4_int_q_acc_3_, npu_inst_pe_1_0_4_int_q_acc_4_,
         npu_inst_pe_1_0_4_int_q_acc_5_, npu_inst_pe_1_0_4_int_q_acc_6_,
         npu_inst_pe_1_0_4_int_q_acc_7_, npu_inst_pe_1_0_4_int_data_0_,
         npu_inst_pe_1_0_4_int_data_1_, npu_inst_pe_1_0_4_int_q_weight_0_,
         npu_inst_pe_1_0_4_int_q_weight_1_,
         npu_inst_pe_1_0_4_int_q_reg_v_5__0_,
         npu_inst_pe_1_0_4_int_q_reg_v_5__1_,
         npu_inst_pe_1_0_4_int_q_reg_v_4__0_,
         npu_inst_pe_1_0_4_int_q_reg_v_4__1_,
         npu_inst_pe_1_0_4_int_q_reg_v_3__0_,
         npu_inst_pe_1_0_4_int_q_reg_v_3__1_,
         npu_inst_pe_1_0_4_int_q_reg_v_2__0_,
         npu_inst_pe_1_0_4_int_q_reg_v_2__1_,
         npu_inst_pe_1_0_4_int_q_reg_v_1__0_,
         npu_inst_pe_1_0_4_int_q_reg_v_1__1_,
         npu_inst_pe_1_0_4_int_q_reg_v_0__0_,
         npu_inst_pe_1_0_4_int_q_reg_v_0__1_,
         npu_inst_pe_1_0_4_int_q_reg_h_5__0_,
         npu_inst_pe_1_0_4_int_q_reg_h_5__1_,
         npu_inst_pe_1_0_4_int_q_reg_h_4__0_,
         npu_inst_pe_1_0_4_int_q_reg_h_4__1_,
         npu_inst_pe_1_0_4_int_q_reg_h_3__0_,
         npu_inst_pe_1_0_4_int_q_reg_h_3__1_,
         npu_inst_pe_1_0_4_int_q_reg_h_2__0_,
         npu_inst_pe_1_0_4_int_q_reg_h_2__1_,
         npu_inst_pe_1_0_4_int_q_reg_h_1__0_,
         npu_inst_pe_1_0_4_int_q_reg_h_1__1_,
         npu_inst_pe_1_0_4_int_q_reg_h_0__0_,
         npu_inst_pe_1_0_4_int_q_reg_h_0__1_, npu_inst_pe_1_0_4_o_data_v_0_,
         npu_inst_pe_1_0_4_o_data_v_1_, npu_inst_pe_1_0_5_n119,
         npu_inst_pe_1_0_5_n118, npu_inst_pe_1_0_5_n117,
         npu_inst_pe_1_0_5_n116, npu_inst_pe_1_0_5_n115,
         npu_inst_pe_1_0_5_n114, npu_inst_pe_1_0_5_n113,
         npu_inst_pe_1_0_5_n112, npu_inst_pe_1_0_5_n111,
         npu_inst_pe_1_0_5_n110, npu_inst_pe_1_0_5_n109,
         npu_inst_pe_1_0_5_n108, npu_inst_pe_1_0_5_n107,
         npu_inst_pe_1_0_5_n106, npu_inst_pe_1_0_5_n105,
         npu_inst_pe_1_0_5_n104, npu_inst_pe_1_0_5_n103,
         npu_inst_pe_1_0_5_n102, npu_inst_pe_1_0_5_n101,
         npu_inst_pe_1_0_5_n100, npu_inst_pe_1_0_5_n99, npu_inst_pe_1_0_5_n98,
         npu_inst_pe_1_0_5_n36, npu_inst_pe_1_0_5_n35, npu_inst_pe_1_0_5_n34,
         npu_inst_pe_1_0_5_n33, npu_inst_pe_1_0_5_n32, npu_inst_pe_1_0_5_n31,
         npu_inst_pe_1_0_5_n30, npu_inst_pe_1_0_5_n29, npu_inst_pe_1_0_5_n28,
         npu_inst_pe_1_0_5_n25, npu_inst_pe_1_0_5_n24, npu_inst_pe_1_0_5_n23,
         npu_inst_pe_1_0_5_n22, npu_inst_pe_1_0_5_n21, npu_inst_pe_1_0_5_n20,
         npu_inst_pe_1_0_5_n19, npu_inst_pe_1_0_5_n18, npu_inst_pe_1_0_5_n17,
         npu_inst_pe_1_0_5_n16, npu_inst_pe_1_0_5_n15, npu_inst_pe_1_0_5_n14,
         npu_inst_pe_1_0_5_n13, npu_inst_pe_1_0_5_n12, npu_inst_pe_1_0_5_n11,
         npu_inst_pe_1_0_5_n10, npu_inst_pe_1_0_5_n9, npu_inst_pe_1_0_5_n8,
         npu_inst_pe_1_0_5_n7, npu_inst_pe_1_0_5_n6, npu_inst_pe_1_0_5_n5,
         npu_inst_pe_1_0_5_n4, npu_inst_pe_1_0_5_n3, npu_inst_pe_1_0_5_n2,
         npu_inst_pe_1_0_5_n1, npu_inst_pe_1_0_5_sub_67_carry_7_,
         npu_inst_pe_1_0_5_sub_67_carry_6_, npu_inst_pe_1_0_5_sub_67_carry_5_,
         npu_inst_pe_1_0_5_sub_67_carry_4_, npu_inst_pe_1_0_5_sub_67_carry_3_,
         npu_inst_pe_1_0_5_sub_67_carry_2_, npu_inst_pe_1_0_5_sub_67_carry_1_,
         npu_inst_pe_1_0_5_add_69_carry_7_, npu_inst_pe_1_0_5_add_69_carry_6_,
         npu_inst_pe_1_0_5_add_69_carry_5_, npu_inst_pe_1_0_5_add_69_carry_4_,
         npu_inst_pe_1_0_5_add_69_carry_3_, npu_inst_pe_1_0_5_add_69_carry_2_,
         npu_inst_pe_1_0_5_add_69_carry_1_, npu_inst_pe_1_0_5_n97,
         npu_inst_pe_1_0_5_n96, npu_inst_pe_1_0_5_n95, npu_inst_pe_1_0_5_n94,
         npu_inst_pe_1_0_5_n93, npu_inst_pe_1_0_5_n92, npu_inst_pe_1_0_5_n91,
         npu_inst_pe_1_0_5_n90, npu_inst_pe_1_0_5_n89, npu_inst_pe_1_0_5_n88,
         npu_inst_pe_1_0_5_n87, npu_inst_pe_1_0_5_n86, npu_inst_pe_1_0_5_n85,
         npu_inst_pe_1_0_5_n84, npu_inst_pe_1_0_5_n83, npu_inst_pe_1_0_5_n82,
         npu_inst_pe_1_0_5_n81, npu_inst_pe_1_0_5_n80, npu_inst_pe_1_0_5_n79,
         npu_inst_pe_1_0_5_n78, npu_inst_pe_1_0_5_n77, npu_inst_pe_1_0_5_n76,
         npu_inst_pe_1_0_5_n75, npu_inst_pe_1_0_5_n74, npu_inst_pe_1_0_5_n73,
         npu_inst_pe_1_0_5_n72, npu_inst_pe_1_0_5_n71, npu_inst_pe_1_0_5_n70,
         npu_inst_pe_1_0_5_n69, npu_inst_pe_1_0_5_n68, npu_inst_pe_1_0_5_n67,
         npu_inst_pe_1_0_5_n66, npu_inst_pe_1_0_5_n65, npu_inst_pe_1_0_5_n64,
         npu_inst_pe_1_0_5_n63, npu_inst_pe_1_0_5_n62, npu_inst_pe_1_0_5_n61,
         npu_inst_pe_1_0_5_n60, npu_inst_pe_1_0_5_n59, npu_inst_pe_1_0_5_n58,
         npu_inst_pe_1_0_5_n57, npu_inst_pe_1_0_5_n56, npu_inst_pe_1_0_5_n55,
         npu_inst_pe_1_0_5_n54, npu_inst_pe_1_0_5_n53, npu_inst_pe_1_0_5_n52,
         npu_inst_pe_1_0_5_n51, npu_inst_pe_1_0_5_n50, npu_inst_pe_1_0_5_n49,
         npu_inst_pe_1_0_5_n48, npu_inst_pe_1_0_5_n47, npu_inst_pe_1_0_5_n46,
         npu_inst_pe_1_0_5_n45, npu_inst_pe_1_0_5_n44, npu_inst_pe_1_0_5_n43,
         npu_inst_pe_1_0_5_n42, npu_inst_pe_1_0_5_n41, npu_inst_pe_1_0_5_n40,
         npu_inst_pe_1_0_5_n39, npu_inst_pe_1_0_5_n38, npu_inst_pe_1_0_5_n37,
         npu_inst_pe_1_0_5_n27, npu_inst_pe_1_0_5_n26,
         npu_inst_pe_1_0_5_net4453, npu_inst_pe_1_0_5_net4447,
         npu_inst_pe_1_0_5_N94, npu_inst_pe_1_0_5_N93, npu_inst_pe_1_0_5_N84,
         npu_inst_pe_1_0_5_N80, npu_inst_pe_1_0_5_N79, npu_inst_pe_1_0_5_N78,
         npu_inst_pe_1_0_5_N77, npu_inst_pe_1_0_5_N76, npu_inst_pe_1_0_5_N75,
         npu_inst_pe_1_0_5_N74, npu_inst_pe_1_0_5_N73, npu_inst_pe_1_0_5_N72,
         npu_inst_pe_1_0_5_N71, npu_inst_pe_1_0_5_N70, npu_inst_pe_1_0_5_N69,
         npu_inst_pe_1_0_5_N68, npu_inst_pe_1_0_5_N67, npu_inst_pe_1_0_5_N66,
         npu_inst_pe_1_0_5_N65, npu_inst_pe_1_0_5_int_q_acc_0_,
         npu_inst_pe_1_0_5_int_q_acc_1_, npu_inst_pe_1_0_5_int_q_acc_2_,
         npu_inst_pe_1_0_5_int_q_acc_3_, npu_inst_pe_1_0_5_int_q_acc_4_,
         npu_inst_pe_1_0_5_int_q_acc_5_, npu_inst_pe_1_0_5_int_q_acc_6_,
         npu_inst_pe_1_0_5_int_q_acc_7_, npu_inst_pe_1_0_5_int_data_0_,
         npu_inst_pe_1_0_5_int_data_1_, npu_inst_pe_1_0_5_int_q_weight_0_,
         npu_inst_pe_1_0_5_int_q_weight_1_,
         npu_inst_pe_1_0_5_int_q_reg_v_5__0_,
         npu_inst_pe_1_0_5_int_q_reg_v_5__1_,
         npu_inst_pe_1_0_5_int_q_reg_v_4__0_,
         npu_inst_pe_1_0_5_int_q_reg_v_4__1_,
         npu_inst_pe_1_0_5_int_q_reg_v_3__0_,
         npu_inst_pe_1_0_5_int_q_reg_v_3__1_,
         npu_inst_pe_1_0_5_int_q_reg_v_2__0_,
         npu_inst_pe_1_0_5_int_q_reg_v_2__1_,
         npu_inst_pe_1_0_5_int_q_reg_v_1__0_,
         npu_inst_pe_1_0_5_int_q_reg_v_1__1_,
         npu_inst_pe_1_0_5_int_q_reg_v_0__0_,
         npu_inst_pe_1_0_5_int_q_reg_v_0__1_,
         npu_inst_pe_1_0_5_int_q_reg_h_5__0_,
         npu_inst_pe_1_0_5_int_q_reg_h_5__1_,
         npu_inst_pe_1_0_5_int_q_reg_h_4__0_,
         npu_inst_pe_1_0_5_int_q_reg_h_4__1_,
         npu_inst_pe_1_0_5_int_q_reg_h_3__0_,
         npu_inst_pe_1_0_5_int_q_reg_h_3__1_,
         npu_inst_pe_1_0_5_int_q_reg_h_2__0_,
         npu_inst_pe_1_0_5_int_q_reg_h_2__1_,
         npu_inst_pe_1_0_5_int_q_reg_h_1__0_,
         npu_inst_pe_1_0_5_int_q_reg_h_1__1_,
         npu_inst_pe_1_0_5_int_q_reg_h_0__0_,
         npu_inst_pe_1_0_5_int_q_reg_h_0__1_, npu_inst_pe_1_0_5_o_data_v_0_,
         npu_inst_pe_1_0_5_o_data_v_1_, npu_inst_pe_1_0_6_n119,
         npu_inst_pe_1_0_6_n118, npu_inst_pe_1_0_6_n117,
         npu_inst_pe_1_0_6_n116, npu_inst_pe_1_0_6_n115,
         npu_inst_pe_1_0_6_n114, npu_inst_pe_1_0_6_n113,
         npu_inst_pe_1_0_6_n112, npu_inst_pe_1_0_6_n111,
         npu_inst_pe_1_0_6_n110, npu_inst_pe_1_0_6_n109,
         npu_inst_pe_1_0_6_n108, npu_inst_pe_1_0_6_n107,
         npu_inst_pe_1_0_6_n106, npu_inst_pe_1_0_6_n105,
         npu_inst_pe_1_0_6_n104, npu_inst_pe_1_0_6_n103,
         npu_inst_pe_1_0_6_n102, npu_inst_pe_1_0_6_n101,
         npu_inst_pe_1_0_6_n100, npu_inst_pe_1_0_6_n99, npu_inst_pe_1_0_6_n98,
         npu_inst_pe_1_0_6_n36, npu_inst_pe_1_0_6_n35, npu_inst_pe_1_0_6_n34,
         npu_inst_pe_1_0_6_n33, npu_inst_pe_1_0_6_n32, npu_inst_pe_1_0_6_n31,
         npu_inst_pe_1_0_6_n30, npu_inst_pe_1_0_6_n29, npu_inst_pe_1_0_6_n28,
         npu_inst_pe_1_0_6_n25, npu_inst_pe_1_0_6_n24, npu_inst_pe_1_0_6_n23,
         npu_inst_pe_1_0_6_n22, npu_inst_pe_1_0_6_n21, npu_inst_pe_1_0_6_n20,
         npu_inst_pe_1_0_6_n19, npu_inst_pe_1_0_6_n18, npu_inst_pe_1_0_6_n17,
         npu_inst_pe_1_0_6_n16, npu_inst_pe_1_0_6_n15, npu_inst_pe_1_0_6_n14,
         npu_inst_pe_1_0_6_n13, npu_inst_pe_1_0_6_n12, npu_inst_pe_1_0_6_n11,
         npu_inst_pe_1_0_6_n10, npu_inst_pe_1_0_6_n9, npu_inst_pe_1_0_6_n8,
         npu_inst_pe_1_0_6_n7, npu_inst_pe_1_0_6_n6, npu_inst_pe_1_0_6_n5,
         npu_inst_pe_1_0_6_n4, npu_inst_pe_1_0_6_n3, npu_inst_pe_1_0_6_n2,
         npu_inst_pe_1_0_6_n1, npu_inst_pe_1_0_6_sub_67_carry_7_,
         npu_inst_pe_1_0_6_sub_67_carry_6_, npu_inst_pe_1_0_6_sub_67_carry_5_,
         npu_inst_pe_1_0_6_sub_67_carry_4_, npu_inst_pe_1_0_6_sub_67_carry_3_,
         npu_inst_pe_1_0_6_sub_67_carry_2_, npu_inst_pe_1_0_6_sub_67_carry_1_,
         npu_inst_pe_1_0_6_add_69_carry_7_, npu_inst_pe_1_0_6_add_69_carry_6_,
         npu_inst_pe_1_0_6_add_69_carry_5_, npu_inst_pe_1_0_6_add_69_carry_4_,
         npu_inst_pe_1_0_6_add_69_carry_3_, npu_inst_pe_1_0_6_add_69_carry_2_,
         npu_inst_pe_1_0_6_add_69_carry_1_, npu_inst_pe_1_0_6_n97,
         npu_inst_pe_1_0_6_n96, npu_inst_pe_1_0_6_n95, npu_inst_pe_1_0_6_n94,
         npu_inst_pe_1_0_6_n93, npu_inst_pe_1_0_6_n92, npu_inst_pe_1_0_6_n91,
         npu_inst_pe_1_0_6_n90, npu_inst_pe_1_0_6_n89, npu_inst_pe_1_0_6_n88,
         npu_inst_pe_1_0_6_n87, npu_inst_pe_1_0_6_n86, npu_inst_pe_1_0_6_n85,
         npu_inst_pe_1_0_6_n84, npu_inst_pe_1_0_6_n83, npu_inst_pe_1_0_6_n82,
         npu_inst_pe_1_0_6_n81, npu_inst_pe_1_0_6_n80, npu_inst_pe_1_0_6_n79,
         npu_inst_pe_1_0_6_n78, npu_inst_pe_1_0_6_n77, npu_inst_pe_1_0_6_n76,
         npu_inst_pe_1_0_6_n75, npu_inst_pe_1_0_6_n74, npu_inst_pe_1_0_6_n73,
         npu_inst_pe_1_0_6_n72, npu_inst_pe_1_0_6_n71, npu_inst_pe_1_0_6_n70,
         npu_inst_pe_1_0_6_n69, npu_inst_pe_1_0_6_n68, npu_inst_pe_1_0_6_n67,
         npu_inst_pe_1_0_6_n66, npu_inst_pe_1_0_6_n65, npu_inst_pe_1_0_6_n64,
         npu_inst_pe_1_0_6_n63, npu_inst_pe_1_0_6_n62, npu_inst_pe_1_0_6_n61,
         npu_inst_pe_1_0_6_n60, npu_inst_pe_1_0_6_n59, npu_inst_pe_1_0_6_n58,
         npu_inst_pe_1_0_6_n57, npu_inst_pe_1_0_6_n56, npu_inst_pe_1_0_6_n55,
         npu_inst_pe_1_0_6_n54, npu_inst_pe_1_0_6_n53, npu_inst_pe_1_0_6_n52,
         npu_inst_pe_1_0_6_n51, npu_inst_pe_1_0_6_n50, npu_inst_pe_1_0_6_n49,
         npu_inst_pe_1_0_6_n48, npu_inst_pe_1_0_6_n47, npu_inst_pe_1_0_6_n46,
         npu_inst_pe_1_0_6_n45, npu_inst_pe_1_0_6_n44, npu_inst_pe_1_0_6_n43,
         npu_inst_pe_1_0_6_n42, npu_inst_pe_1_0_6_n41, npu_inst_pe_1_0_6_n40,
         npu_inst_pe_1_0_6_n39, npu_inst_pe_1_0_6_n38, npu_inst_pe_1_0_6_n37,
         npu_inst_pe_1_0_6_n27, npu_inst_pe_1_0_6_n26,
         npu_inst_pe_1_0_6_net4430, npu_inst_pe_1_0_6_net4424,
         npu_inst_pe_1_0_6_N94, npu_inst_pe_1_0_6_N93, npu_inst_pe_1_0_6_N84,
         npu_inst_pe_1_0_6_N80, npu_inst_pe_1_0_6_N79, npu_inst_pe_1_0_6_N78,
         npu_inst_pe_1_0_6_N77, npu_inst_pe_1_0_6_N76, npu_inst_pe_1_0_6_N75,
         npu_inst_pe_1_0_6_N74, npu_inst_pe_1_0_6_N73, npu_inst_pe_1_0_6_N72,
         npu_inst_pe_1_0_6_N71, npu_inst_pe_1_0_6_N70, npu_inst_pe_1_0_6_N69,
         npu_inst_pe_1_0_6_N68, npu_inst_pe_1_0_6_N67, npu_inst_pe_1_0_6_N66,
         npu_inst_pe_1_0_6_N65, npu_inst_pe_1_0_6_int_q_acc_0_,
         npu_inst_pe_1_0_6_int_q_acc_1_, npu_inst_pe_1_0_6_int_q_acc_2_,
         npu_inst_pe_1_0_6_int_q_acc_3_, npu_inst_pe_1_0_6_int_q_acc_4_,
         npu_inst_pe_1_0_6_int_q_acc_5_, npu_inst_pe_1_0_6_int_q_acc_6_,
         npu_inst_pe_1_0_6_int_q_acc_7_, npu_inst_pe_1_0_6_int_data_0_,
         npu_inst_pe_1_0_6_int_data_1_, npu_inst_pe_1_0_6_int_q_weight_0_,
         npu_inst_pe_1_0_6_int_q_weight_1_,
         npu_inst_pe_1_0_6_int_q_reg_v_5__0_,
         npu_inst_pe_1_0_6_int_q_reg_v_5__1_,
         npu_inst_pe_1_0_6_int_q_reg_v_4__0_,
         npu_inst_pe_1_0_6_int_q_reg_v_4__1_,
         npu_inst_pe_1_0_6_int_q_reg_v_3__0_,
         npu_inst_pe_1_0_6_int_q_reg_v_3__1_,
         npu_inst_pe_1_0_6_int_q_reg_v_2__0_,
         npu_inst_pe_1_0_6_int_q_reg_v_2__1_,
         npu_inst_pe_1_0_6_int_q_reg_v_1__0_,
         npu_inst_pe_1_0_6_int_q_reg_v_1__1_,
         npu_inst_pe_1_0_6_int_q_reg_v_0__0_,
         npu_inst_pe_1_0_6_int_q_reg_v_0__1_,
         npu_inst_pe_1_0_6_int_q_reg_h_5__0_,
         npu_inst_pe_1_0_6_int_q_reg_h_5__1_,
         npu_inst_pe_1_0_6_int_q_reg_h_4__0_,
         npu_inst_pe_1_0_6_int_q_reg_h_4__1_,
         npu_inst_pe_1_0_6_int_q_reg_h_3__0_,
         npu_inst_pe_1_0_6_int_q_reg_h_3__1_,
         npu_inst_pe_1_0_6_int_q_reg_h_2__0_,
         npu_inst_pe_1_0_6_int_q_reg_h_2__1_,
         npu_inst_pe_1_0_6_int_q_reg_h_1__0_,
         npu_inst_pe_1_0_6_int_q_reg_h_1__1_,
         npu_inst_pe_1_0_6_int_q_reg_h_0__0_,
         npu_inst_pe_1_0_6_int_q_reg_h_0__1_, npu_inst_pe_1_0_6_o_data_v_0_,
         npu_inst_pe_1_0_6_o_data_v_1_, npu_inst_pe_1_0_7_n119,
         npu_inst_pe_1_0_7_n118, npu_inst_pe_1_0_7_n117,
         npu_inst_pe_1_0_7_n116, npu_inst_pe_1_0_7_n115,
         npu_inst_pe_1_0_7_n114, npu_inst_pe_1_0_7_n113,
         npu_inst_pe_1_0_7_n112, npu_inst_pe_1_0_7_n111,
         npu_inst_pe_1_0_7_n110, npu_inst_pe_1_0_7_n109,
         npu_inst_pe_1_0_7_n108, npu_inst_pe_1_0_7_n107,
         npu_inst_pe_1_0_7_n106, npu_inst_pe_1_0_7_n105,
         npu_inst_pe_1_0_7_n104, npu_inst_pe_1_0_7_n103,
         npu_inst_pe_1_0_7_n102, npu_inst_pe_1_0_7_n101,
         npu_inst_pe_1_0_7_n100, npu_inst_pe_1_0_7_n99, npu_inst_pe_1_0_7_n98,
         npu_inst_pe_1_0_7_n36, npu_inst_pe_1_0_7_n35, npu_inst_pe_1_0_7_n34,
         npu_inst_pe_1_0_7_n33, npu_inst_pe_1_0_7_n32, npu_inst_pe_1_0_7_n31,
         npu_inst_pe_1_0_7_n30, npu_inst_pe_1_0_7_n29, npu_inst_pe_1_0_7_n28,
         npu_inst_pe_1_0_7_n25, npu_inst_pe_1_0_7_n24, npu_inst_pe_1_0_7_n23,
         npu_inst_pe_1_0_7_n22, npu_inst_pe_1_0_7_n21, npu_inst_pe_1_0_7_n20,
         npu_inst_pe_1_0_7_n19, npu_inst_pe_1_0_7_n18, npu_inst_pe_1_0_7_n17,
         npu_inst_pe_1_0_7_n16, npu_inst_pe_1_0_7_n15, npu_inst_pe_1_0_7_n14,
         npu_inst_pe_1_0_7_n13, npu_inst_pe_1_0_7_n12, npu_inst_pe_1_0_7_n11,
         npu_inst_pe_1_0_7_n10, npu_inst_pe_1_0_7_n9, npu_inst_pe_1_0_7_n8,
         npu_inst_pe_1_0_7_n7, npu_inst_pe_1_0_7_n6, npu_inst_pe_1_0_7_n5,
         npu_inst_pe_1_0_7_n4, npu_inst_pe_1_0_7_n3, npu_inst_pe_1_0_7_n2,
         npu_inst_pe_1_0_7_n1, npu_inst_pe_1_0_7_sub_67_carry_7_,
         npu_inst_pe_1_0_7_sub_67_carry_6_, npu_inst_pe_1_0_7_sub_67_carry_5_,
         npu_inst_pe_1_0_7_sub_67_carry_4_, npu_inst_pe_1_0_7_sub_67_carry_3_,
         npu_inst_pe_1_0_7_sub_67_carry_2_, npu_inst_pe_1_0_7_sub_67_carry_1_,
         npu_inst_pe_1_0_7_add_69_carry_7_, npu_inst_pe_1_0_7_add_69_carry_6_,
         npu_inst_pe_1_0_7_add_69_carry_5_, npu_inst_pe_1_0_7_add_69_carry_4_,
         npu_inst_pe_1_0_7_add_69_carry_3_, npu_inst_pe_1_0_7_add_69_carry_2_,
         npu_inst_pe_1_0_7_add_69_carry_1_, npu_inst_pe_1_0_7_n97,
         npu_inst_pe_1_0_7_n96, npu_inst_pe_1_0_7_n95, npu_inst_pe_1_0_7_n94,
         npu_inst_pe_1_0_7_n93, npu_inst_pe_1_0_7_n92, npu_inst_pe_1_0_7_n91,
         npu_inst_pe_1_0_7_n90, npu_inst_pe_1_0_7_n89, npu_inst_pe_1_0_7_n88,
         npu_inst_pe_1_0_7_n87, npu_inst_pe_1_0_7_n86, npu_inst_pe_1_0_7_n85,
         npu_inst_pe_1_0_7_n84, npu_inst_pe_1_0_7_n83, npu_inst_pe_1_0_7_n82,
         npu_inst_pe_1_0_7_n81, npu_inst_pe_1_0_7_n80, npu_inst_pe_1_0_7_n79,
         npu_inst_pe_1_0_7_n78, npu_inst_pe_1_0_7_n77, npu_inst_pe_1_0_7_n76,
         npu_inst_pe_1_0_7_n75, npu_inst_pe_1_0_7_n74, npu_inst_pe_1_0_7_n73,
         npu_inst_pe_1_0_7_n72, npu_inst_pe_1_0_7_n71, npu_inst_pe_1_0_7_n70,
         npu_inst_pe_1_0_7_n69, npu_inst_pe_1_0_7_n68, npu_inst_pe_1_0_7_n67,
         npu_inst_pe_1_0_7_n66, npu_inst_pe_1_0_7_n65, npu_inst_pe_1_0_7_n64,
         npu_inst_pe_1_0_7_n63, npu_inst_pe_1_0_7_n62, npu_inst_pe_1_0_7_n61,
         npu_inst_pe_1_0_7_n60, npu_inst_pe_1_0_7_n59, npu_inst_pe_1_0_7_n58,
         npu_inst_pe_1_0_7_n57, npu_inst_pe_1_0_7_n56, npu_inst_pe_1_0_7_n55,
         npu_inst_pe_1_0_7_n54, npu_inst_pe_1_0_7_n53, npu_inst_pe_1_0_7_n52,
         npu_inst_pe_1_0_7_n51, npu_inst_pe_1_0_7_n50, npu_inst_pe_1_0_7_n49,
         npu_inst_pe_1_0_7_n48, npu_inst_pe_1_0_7_n47, npu_inst_pe_1_0_7_n46,
         npu_inst_pe_1_0_7_n45, npu_inst_pe_1_0_7_n44, npu_inst_pe_1_0_7_n43,
         npu_inst_pe_1_0_7_n42, npu_inst_pe_1_0_7_n41, npu_inst_pe_1_0_7_n40,
         npu_inst_pe_1_0_7_n39, npu_inst_pe_1_0_7_n38, npu_inst_pe_1_0_7_n37,
         npu_inst_pe_1_0_7_n27, npu_inst_pe_1_0_7_n26,
         npu_inst_pe_1_0_7_net4407, npu_inst_pe_1_0_7_net4401,
         npu_inst_pe_1_0_7_N94, npu_inst_pe_1_0_7_N93, npu_inst_pe_1_0_7_N84,
         npu_inst_pe_1_0_7_N80, npu_inst_pe_1_0_7_N79, npu_inst_pe_1_0_7_N78,
         npu_inst_pe_1_0_7_N77, npu_inst_pe_1_0_7_N76, npu_inst_pe_1_0_7_N75,
         npu_inst_pe_1_0_7_N74, npu_inst_pe_1_0_7_N73, npu_inst_pe_1_0_7_N72,
         npu_inst_pe_1_0_7_N71, npu_inst_pe_1_0_7_N70, npu_inst_pe_1_0_7_N69,
         npu_inst_pe_1_0_7_N68, npu_inst_pe_1_0_7_N67, npu_inst_pe_1_0_7_N66,
         npu_inst_pe_1_0_7_N65, npu_inst_pe_1_0_7_int_q_acc_0_,
         npu_inst_pe_1_0_7_int_q_acc_1_, npu_inst_pe_1_0_7_int_q_acc_2_,
         npu_inst_pe_1_0_7_int_q_acc_3_, npu_inst_pe_1_0_7_int_q_acc_4_,
         npu_inst_pe_1_0_7_int_q_acc_5_, npu_inst_pe_1_0_7_int_q_acc_6_,
         npu_inst_pe_1_0_7_int_q_acc_7_, npu_inst_pe_1_0_7_int_data_0_,
         npu_inst_pe_1_0_7_int_data_1_, npu_inst_pe_1_0_7_int_q_weight_0_,
         npu_inst_pe_1_0_7_int_q_weight_1_,
         npu_inst_pe_1_0_7_int_q_reg_v_5__0_,
         npu_inst_pe_1_0_7_int_q_reg_v_5__1_,
         npu_inst_pe_1_0_7_int_q_reg_v_4__0_,
         npu_inst_pe_1_0_7_int_q_reg_v_4__1_,
         npu_inst_pe_1_0_7_int_q_reg_v_3__0_,
         npu_inst_pe_1_0_7_int_q_reg_v_3__1_,
         npu_inst_pe_1_0_7_int_q_reg_v_2__0_,
         npu_inst_pe_1_0_7_int_q_reg_v_2__1_,
         npu_inst_pe_1_0_7_int_q_reg_v_1__0_,
         npu_inst_pe_1_0_7_int_q_reg_v_1__1_,
         npu_inst_pe_1_0_7_int_q_reg_v_0__0_,
         npu_inst_pe_1_0_7_int_q_reg_v_0__1_,
         npu_inst_pe_1_0_7_int_q_reg_h_5__0_,
         npu_inst_pe_1_0_7_int_q_reg_h_5__1_,
         npu_inst_pe_1_0_7_int_q_reg_h_4__0_,
         npu_inst_pe_1_0_7_int_q_reg_h_4__1_,
         npu_inst_pe_1_0_7_int_q_reg_h_3__0_,
         npu_inst_pe_1_0_7_int_q_reg_h_3__1_,
         npu_inst_pe_1_0_7_int_q_reg_h_2__0_,
         npu_inst_pe_1_0_7_int_q_reg_h_2__1_,
         npu_inst_pe_1_0_7_int_q_reg_h_1__0_,
         npu_inst_pe_1_0_7_int_q_reg_h_1__1_,
         npu_inst_pe_1_0_7_int_q_reg_h_0__0_,
         npu_inst_pe_1_0_7_int_q_reg_h_0__1_, npu_inst_pe_1_0_7_o_data_v_0_,
         npu_inst_pe_1_0_7_o_data_v_1_, npu_inst_pe_1_1_0_n119,
         npu_inst_pe_1_1_0_n118, npu_inst_pe_1_1_0_n117,
         npu_inst_pe_1_1_0_n116, npu_inst_pe_1_1_0_n115,
         npu_inst_pe_1_1_0_n114, npu_inst_pe_1_1_0_n113,
         npu_inst_pe_1_1_0_n112, npu_inst_pe_1_1_0_n111,
         npu_inst_pe_1_1_0_n110, npu_inst_pe_1_1_0_n109,
         npu_inst_pe_1_1_0_n108, npu_inst_pe_1_1_0_n107,
         npu_inst_pe_1_1_0_n106, npu_inst_pe_1_1_0_n105,
         npu_inst_pe_1_1_0_n104, npu_inst_pe_1_1_0_n103,
         npu_inst_pe_1_1_0_n102, npu_inst_pe_1_1_0_n101,
         npu_inst_pe_1_1_0_n100, npu_inst_pe_1_1_0_n99, npu_inst_pe_1_1_0_n98,
         npu_inst_pe_1_1_0_n36, npu_inst_pe_1_1_0_n35, npu_inst_pe_1_1_0_n34,
         npu_inst_pe_1_1_0_n33, npu_inst_pe_1_1_0_n32, npu_inst_pe_1_1_0_n31,
         npu_inst_pe_1_1_0_n30, npu_inst_pe_1_1_0_n29, npu_inst_pe_1_1_0_n28,
         npu_inst_pe_1_1_0_n25, npu_inst_pe_1_1_0_n24, npu_inst_pe_1_1_0_n23,
         npu_inst_pe_1_1_0_n22, npu_inst_pe_1_1_0_n21, npu_inst_pe_1_1_0_n20,
         npu_inst_pe_1_1_0_n19, npu_inst_pe_1_1_0_n18, npu_inst_pe_1_1_0_n17,
         npu_inst_pe_1_1_0_n16, npu_inst_pe_1_1_0_n15, npu_inst_pe_1_1_0_n14,
         npu_inst_pe_1_1_0_n13, npu_inst_pe_1_1_0_n12, npu_inst_pe_1_1_0_n11,
         npu_inst_pe_1_1_0_n10, npu_inst_pe_1_1_0_n9, npu_inst_pe_1_1_0_n8,
         npu_inst_pe_1_1_0_n7, npu_inst_pe_1_1_0_n6, npu_inst_pe_1_1_0_n5,
         npu_inst_pe_1_1_0_n4, npu_inst_pe_1_1_0_n3, npu_inst_pe_1_1_0_n2,
         npu_inst_pe_1_1_0_n1, npu_inst_pe_1_1_0_sub_67_carry_7_,
         npu_inst_pe_1_1_0_sub_67_carry_6_, npu_inst_pe_1_1_0_sub_67_carry_5_,
         npu_inst_pe_1_1_0_sub_67_carry_4_, npu_inst_pe_1_1_0_sub_67_carry_3_,
         npu_inst_pe_1_1_0_sub_67_carry_2_, npu_inst_pe_1_1_0_sub_67_carry_1_,
         npu_inst_pe_1_1_0_add_69_carry_7_, npu_inst_pe_1_1_0_add_69_carry_6_,
         npu_inst_pe_1_1_0_add_69_carry_5_, npu_inst_pe_1_1_0_add_69_carry_4_,
         npu_inst_pe_1_1_0_add_69_carry_3_, npu_inst_pe_1_1_0_add_69_carry_2_,
         npu_inst_pe_1_1_0_add_69_carry_1_, npu_inst_pe_1_1_0_n97,
         npu_inst_pe_1_1_0_n96, npu_inst_pe_1_1_0_n95, npu_inst_pe_1_1_0_n94,
         npu_inst_pe_1_1_0_n93, npu_inst_pe_1_1_0_n92, npu_inst_pe_1_1_0_n91,
         npu_inst_pe_1_1_0_n90, npu_inst_pe_1_1_0_n89, npu_inst_pe_1_1_0_n88,
         npu_inst_pe_1_1_0_n87, npu_inst_pe_1_1_0_n86, npu_inst_pe_1_1_0_n85,
         npu_inst_pe_1_1_0_n84, npu_inst_pe_1_1_0_n83, npu_inst_pe_1_1_0_n82,
         npu_inst_pe_1_1_0_n81, npu_inst_pe_1_1_0_n80, npu_inst_pe_1_1_0_n79,
         npu_inst_pe_1_1_0_n78, npu_inst_pe_1_1_0_n77, npu_inst_pe_1_1_0_n76,
         npu_inst_pe_1_1_0_n75, npu_inst_pe_1_1_0_n74, npu_inst_pe_1_1_0_n73,
         npu_inst_pe_1_1_0_n72, npu_inst_pe_1_1_0_n71, npu_inst_pe_1_1_0_n70,
         npu_inst_pe_1_1_0_n69, npu_inst_pe_1_1_0_n68, npu_inst_pe_1_1_0_n67,
         npu_inst_pe_1_1_0_n66, npu_inst_pe_1_1_0_n65, npu_inst_pe_1_1_0_n64,
         npu_inst_pe_1_1_0_n63, npu_inst_pe_1_1_0_n62, npu_inst_pe_1_1_0_n61,
         npu_inst_pe_1_1_0_n60, npu_inst_pe_1_1_0_n59, npu_inst_pe_1_1_0_n58,
         npu_inst_pe_1_1_0_n57, npu_inst_pe_1_1_0_n56, npu_inst_pe_1_1_0_n55,
         npu_inst_pe_1_1_0_n54, npu_inst_pe_1_1_0_n53, npu_inst_pe_1_1_0_n52,
         npu_inst_pe_1_1_0_n51, npu_inst_pe_1_1_0_n50, npu_inst_pe_1_1_0_n49,
         npu_inst_pe_1_1_0_n48, npu_inst_pe_1_1_0_n47, npu_inst_pe_1_1_0_n46,
         npu_inst_pe_1_1_0_n45, npu_inst_pe_1_1_0_n44, npu_inst_pe_1_1_0_n43,
         npu_inst_pe_1_1_0_n42, npu_inst_pe_1_1_0_n41, npu_inst_pe_1_1_0_n40,
         npu_inst_pe_1_1_0_n39, npu_inst_pe_1_1_0_n38, npu_inst_pe_1_1_0_n37,
         npu_inst_pe_1_1_0_n27, npu_inst_pe_1_1_0_n26,
         npu_inst_pe_1_1_0_net4384, npu_inst_pe_1_1_0_net4378,
         npu_inst_pe_1_1_0_N94, npu_inst_pe_1_1_0_N93, npu_inst_pe_1_1_0_N84,
         npu_inst_pe_1_1_0_N80, npu_inst_pe_1_1_0_N79, npu_inst_pe_1_1_0_N78,
         npu_inst_pe_1_1_0_N77, npu_inst_pe_1_1_0_N76, npu_inst_pe_1_1_0_N75,
         npu_inst_pe_1_1_0_N74, npu_inst_pe_1_1_0_N73, npu_inst_pe_1_1_0_N72,
         npu_inst_pe_1_1_0_N71, npu_inst_pe_1_1_0_N70, npu_inst_pe_1_1_0_N69,
         npu_inst_pe_1_1_0_N68, npu_inst_pe_1_1_0_N67, npu_inst_pe_1_1_0_N66,
         npu_inst_pe_1_1_0_N65, npu_inst_pe_1_1_0_int_q_acc_0_,
         npu_inst_pe_1_1_0_int_q_acc_1_, npu_inst_pe_1_1_0_int_q_acc_2_,
         npu_inst_pe_1_1_0_int_q_acc_3_, npu_inst_pe_1_1_0_int_q_acc_4_,
         npu_inst_pe_1_1_0_int_q_acc_5_, npu_inst_pe_1_1_0_int_q_acc_6_,
         npu_inst_pe_1_1_0_int_q_acc_7_, npu_inst_pe_1_1_0_int_data_0_,
         npu_inst_pe_1_1_0_int_data_1_, npu_inst_pe_1_1_0_int_q_weight_0_,
         npu_inst_pe_1_1_0_int_q_weight_1_,
         npu_inst_pe_1_1_0_int_q_reg_v_5__0_,
         npu_inst_pe_1_1_0_int_q_reg_v_5__1_,
         npu_inst_pe_1_1_0_int_q_reg_v_4__0_,
         npu_inst_pe_1_1_0_int_q_reg_v_4__1_,
         npu_inst_pe_1_1_0_int_q_reg_v_3__0_,
         npu_inst_pe_1_1_0_int_q_reg_v_3__1_,
         npu_inst_pe_1_1_0_int_q_reg_v_2__0_,
         npu_inst_pe_1_1_0_int_q_reg_v_2__1_,
         npu_inst_pe_1_1_0_int_q_reg_v_1__0_,
         npu_inst_pe_1_1_0_int_q_reg_v_1__1_,
         npu_inst_pe_1_1_0_int_q_reg_v_0__0_,
         npu_inst_pe_1_1_0_int_q_reg_v_0__1_,
         npu_inst_pe_1_1_0_int_q_reg_h_5__0_,
         npu_inst_pe_1_1_0_int_q_reg_h_5__1_,
         npu_inst_pe_1_1_0_int_q_reg_h_4__0_,
         npu_inst_pe_1_1_0_int_q_reg_h_4__1_,
         npu_inst_pe_1_1_0_int_q_reg_h_3__0_,
         npu_inst_pe_1_1_0_int_q_reg_h_3__1_,
         npu_inst_pe_1_1_0_int_q_reg_h_2__0_,
         npu_inst_pe_1_1_0_int_q_reg_h_2__1_,
         npu_inst_pe_1_1_0_int_q_reg_h_1__0_,
         npu_inst_pe_1_1_0_int_q_reg_h_1__1_,
         npu_inst_pe_1_1_0_int_q_reg_h_0__0_,
         npu_inst_pe_1_1_0_int_q_reg_h_0__1_, npu_inst_pe_1_1_0_o_data_h_0_,
         npu_inst_pe_1_1_0_o_data_h_1_, npu_inst_pe_1_1_1_n119,
         npu_inst_pe_1_1_1_n118, npu_inst_pe_1_1_1_n117,
         npu_inst_pe_1_1_1_n116, npu_inst_pe_1_1_1_n115,
         npu_inst_pe_1_1_1_n114, npu_inst_pe_1_1_1_n113,
         npu_inst_pe_1_1_1_n112, npu_inst_pe_1_1_1_n111,
         npu_inst_pe_1_1_1_n110, npu_inst_pe_1_1_1_n109,
         npu_inst_pe_1_1_1_n108, npu_inst_pe_1_1_1_n107,
         npu_inst_pe_1_1_1_n106, npu_inst_pe_1_1_1_n105,
         npu_inst_pe_1_1_1_n104, npu_inst_pe_1_1_1_n103,
         npu_inst_pe_1_1_1_n102, npu_inst_pe_1_1_1_n101,
         npu_inst_pe_1_1_1_n100, npu_inst_pe_1_1_1_n99, npu_inst_pe_1_1_1_n98,
         npu_inst_pe_1_1_1_n36, npu_inst_pe_1_1_1_n35, npu_inst_pe_1_1_1_n34,
         npu_inst_pe_1_1_1_n33, npu_inst_pe_1_1_1_n32, npu_inst_pe_1_1_1_n31,
         npu_inst_pe_1_1_1_n30, npu_inst_pe_1_1_1_n29, npu_inst_pe_1_1_1_n28,
         npu_inst_pe_1_1_1_n25, npu_inst_pe_1_1_1_n24, npu_inst_pe_1_1_1_n23,
         npu_inst_pe_1_1_1_n22, npu_inst_pe_1_1_1_n21, npu_inst_pe_1_1_1_n20,
         npu_inst_pe_1_1_1_n19, npu_inst_pe_1_1_1_n18, npu_inst_pe_1_1_1_n17,
         npu_inst_pe_1_1_1_n16, npu_inst_pe_1_1_1_n15, npu_inst_pe_1_1_1_n14,
         npu_inst_pe_1_1_1_n13, npu_inst_pe_1_1_1_n12, npu_inst_pe_1_1_1_n11,
         npu_inst_pe_1_1_1_n10, npu_inst_pe_1_1_1_n9, npu_inst_pe_1_1_1_n8,
         npu_inst_pe_1_1_1_n7, npu_inst_pe_1_1_1_n6, npu_inst_pe_1_1_1_n5,
         npu_inst_pe_1_1_1_n4, npu_inst_pe_1_1_1_n3, npu_inst_pe_1_1_1_n2,
         npu_inst_pe_1_1_1_n1, npu_inst_pe_1_1_1_sub_67_carry_7_,
         npu_inst_pe_1_1_1_sub_67_carry_6_, npu_inst_pe_1_1_1_sub_67_carry_5_,
         npu_inst_pe_1_1_1_sub_67_carry_4_, npu_inst_pe_1_1_1_sub_67_carry_3_,
         npu_inst_pe_1_1_1_sub_67_carry_2_, npu_inst_pe_1_1_1_sub_67_carry_1_,
         npu_inst_pe_1_1_1_add_69_carry_7_, npu_inst_pe_1_1_1_add_69_carry_6_,
         npu_inst_pe_1_1_1_add_69_carry_5_, npu_inst_pe_1_1_1_add_69_carry_4_,
         npu_inst_pe_1_1_1_add_69_carry_3_, npu_inst_pe_1_1_1_add_69_carry_2_,
         npu_inst_pe_1_1_1_add_69_carry_1_, npu_inst_pe_1_1_1_n97,
         npu_inst_pe_1_1_1_n96, npu_inst_pe_1_1_1_n95, npu_inst_pe_1_1_1_n94,
         npu_inst_pe_1_1_1_n93, npu_inst_pe_1_1_1_n92, npu_inst_pe_1_1_1_n91,
         npu_inst_pe_1_1_1_n90, npu_inst_pe_1_1_1_n89, npu_inst_pe_1_1_1_n88,
         npu_inst_pe_1_1_1_n87, npu_inst_pe_1_1_1_n86, npu_inst_pe_1_1_1_n85,
         npu_inst_pe_1_1_1_n84, npu_inst_pe_1_1_1_n83, npu_inst_pe_1_1_1_n82,
         npu_inst_pe_1_1_1_n81, npu_inst_pe_1_1_1_n80, npu_inst_pe_1_1_1_n79,
         npu_inst_pe_1_1_1_n78, npu_inst_pe_1_1_1_n77, npu_inst_pe_1_1_1_n76,
         npu_inst_pe_1_1_1_n75, npu_inst_pe_1_1_1_n74, npu_inst_pe_1_1_1_n73,
         npu_inst_pe_1_1_1_n72, npu_inst_pe_1_1_1_n71, npu_inst_pe_1_1_1_n70,
         npu_inst_pe_1_1_1_n69, npu_inst_pe_1_1_1_n68, npu_inst_pe_1_1_1_n67,
         npu_inst_pe_1_1_1_n66, npu_inst_pe_1_1_1_n65, npu_inst_pe_1_1_1_n64,
         npu_inst_pe_1_1_1_n63, npu_inst_pe_1_1_1_n62, npu_inst_pe_1_1_1_n61,
         npu_inst_pe_1_1_1_n60, npu_inst_pe_1_1_1_n59, npu_inst_pe_1_1_1_n58,
         npu_inst_pe_1_1_1_n57, npu_inst_pe_1_1_1_n56, npu_inst_pe_1_1_1_n55,
         npu_inst_pe_1_1_1_n54, npu_inst_pe_1_1_1_n53, npu_inst_pe_1_1_1_n52,
         npu_inst_pe_1_1_1_n51, npu_inst_pe_1_1_1_n50, npu_inst_pe_1_1_1_n49,
         npu_inst_pe_1_1_1_n48, npu_inst_pe_1_1_1_n47, npu_inst_pe_1_1_1_n46,
         npu_inst_pe_1_1_1_n45, npu_inst_pe_1_1_1_n44, npu_inst_pe_1_1_1_n43,
         npu_inst_pe_1_1_1_n42, npu_inst_pe_1_1_1_n41, npu_inst_pe_1_1_1_n40,
         npu_inst_pe_1_1_1_n39, npu_inst_pe_1_1_1_n38, npu_inst_pe_1_1_1_n37,
         npu_inst_pe_1_1_1_n27, npu_inst_pe_1_1_1_n26,
         npu_inst_pe_1_1_1_net4361, npu_inst_pe_1_1_1_net4355,
         npu_inst_pe_1_1_1_N94, npu_inst_pe_1_1_1_N93, npu_inst_pe_1_1_1_N84,
         npu_inst_pe_1_1_1_N80, npu_inst_pe_1_1_1_N79, npu_inst_pe_1_1_1_N78,
         npu_inst_pe_1_1_1_N77, npu_inst_pe_1_1_1_N76, npu_inst_pe_1_1_1_N75,
         npu_inst_pe_1_1_1_N74, npu_inst_pe_1_1_1_N73, npu_inst_pe_1_1_1_N72,
         npu_inst_pe_1_1_1_N71, npu_inst_pe_1_1_1_N70, npu_inst_pe_1_1_1_N69,
         npu_inst_pe_1_1_1_N68, npu_inst_pe_1_1_1_N67, npu_inst_pe_1_1_1_N66,
         npu_inst_pe_1_1_1_N65, npu_inst_pe_1_1_1_int_q_acc_0_,
         npu_inst_pe_1_1_1_int_q_acc_1_, npu_inst_pe_1_1_1_int_q_acc_2_,
         npu_inst_pe_1_1_1_int_q_acc_3_, npu_inst_pe_1_1_1_int_q_acc_4_,
         npu_inst_pe_1_1_1_int_q_acc_5_, npu_inst_pe_1_1_1_int_q_acc_6_,
         npu_inst_pe_1_1_1_int_q_acc_7_, npu_inst_pe_1_1_1_int_data_0_,
         npu_inst_pe_1_1_1_int_data_1_, npu_inst_pe_1_1_1_int_q_weight_0_,
         npu_inst_pe_1_1_1_int_q_weight_1_,
         npu_inst_pe_1_1_1_int_q_reg_v_5__0_,
         npu_inst_pe_1_1_1_int_q_reg_v_5__1_,
         npu_inst_pe_1_1_1_int_q_reg_v_4__0_,
         npu_inst_pe_1_1_1_int_q_reg_v_4__1_,
         npu_inst_pe_1_1_1_int_q_reg_v_3__0_,
         npu_inst_pe_1_1_1_int_q_reg_v_3__1_,
         npu_inst_pe_1_1_1_int_q_reg_v_2__0_,
         npu_inst_pe_1_1_1_int_q_reg_v_2__1_,
         npu_inst_pe_1_1_1_int_q_reg_v_1__0_,
         npu_inst_pe_1_1_1_int_q_reg_v_1__1_,
         npu_inst_pe_1_1_1_int_q_reg_v_0__0_,
         npu_inst_pe_1_1_1_int_q_reg_v_0__1_,
         npu_inst_pe_1_1_1_int_q_reg_h_5__0_,
         npu_inst_pe_1_1_1_int_q_reg_h_5__1_,
         npu_inst_pe_1_1_1_int_q_reg_h_4__0_,
         npu_inst_pe_1_1_1_int_q_reg_h_4__1_,
         npu_inst_pe_1_1_1_int_q_reg_h_3__0_,
         npu_inst_pe_1_1_1_int_q_reg_h_3__1_,
         npu_inst_pe_1_1_1_int_q_reg_h_2__0_,
         npu_inst_pe_1_1_1_int_q_reg_h_2__1_,
         npu_inst_pe_1_1_1_int_q_reg_h_1__0_,
         npu_inst_pe_1_1_1_int_q_reg_h_1__1_,
         npu_inst_pe_1_1_1_int_q_reg_h_0__0_,
         npu_inst_pe_1_1_1_int_q_reg_h_0__1_, npu_inst_pe_1_1_2_n119,
         npu_inst_pe_1_1_2_n118, npu_inst_pe_1_1_2_n117,
         npu_inst_pe_1_1_2_n116, npu_inst_pe_1_1_2_n115,
         npu_inst_pe_1_1_2_n114, npu_inst_pe_1_1_2_n113,
         npu_inst_pe_1_1_2_n112, npu_inst_pe_1_1_2_n111,
         npu_inst_pe_1_1_2_n110, npu_inst_pe_1_1_2_n109,
         npu_inst_pe_1_1_2_n108, npu_inst_pe_1_1_2_n107,
         npu_inst_pe_1_1_2_n106, npu_inst_pe_1_1_2_n105,
         npu_inst_pe_1_1_2_n104, npu_inst_pe_1_1_2_n103,
         npu_inst_pe_1_1_2_n102, npu_inst_pe_1_1_2_n101,
         npu_inst_pe_1_1_2_n100, npu_inst_pe_1_1_2_n99, npu_inst_pe_1_1_2_n98,
         npu_inst_pe_1_1_2_n36, npu_inst_pe_1_1_2_n35, npu_inst_pe_1_1_2_n34,
         npu_inst_pe_1_1_2_n33, npu_inst_pe_1_1_2_n32, npu_inst_pe_1_1_2_n31,
         npu_inst_pe_1_1_2_n30, npu_inst_pe_1_1_2_n29, npu_inst_pe_1_1_2_n28,
         npu_inst_pe_1_1_2_n25, npu_inst_pe_1_1_2_n24, npu_inst_pe_1_1_2_n23,
         npu_inst_pe_1_1_2_n22, npu_inst_pe_1_1_2_n21, npu_inst_pe_1_1_2_n20,
         npu_inst_pe_1_1_2_n19, npu_inst_pe_1_1_2_n18, npu_inst_pe_1_1_2_n17,
         npu_inst_pe_1_1_2_n16, npu_inst_pe_1_1_2_n15, npu_inst_pe_1_1_2_n14,
         npu_inst_pe_1_1_2_n13, npu_inst_pe_1_1_2_n12, npu_inst_pe_1_1_2_n11,
         npu_inst_pe_1_1_2_n10, npu_inst_pe_1_1_2_n9, npu_inst_pe_1_1_2_n8,
         npu_inst_pe_1_1_2_n7, npu_inst_pe_1_1_2_n6, npu_inst_pe_1_1_2_n5,
         npu_inst_pe_1_1_2_n4, npu_inst_pe_1_1_2_n3, npu_inst_pe_1_1_2_n2,
         npu_inst_pe_1_1_2_n1, npu_inst_pe_1_1_2_sub_67_carry_7_,
         npu_inst_pe_1_1_2_sub_67_carry_6_, npu_inst_pe_1_1_2_sub_67_carry_5_,
         npu_inst_pe_1_1_2_sub_67_carry_4_, npu_inst_pe_1_1_2_sub_67_carry_3_,
         npu_inst_pe_1_1_2_sub_67_carry_2_, npu_inst_pe_1_1_2_sub_67_carry_1_,
         npu_inst_pe_1_1_2_add_69_carry_7_, npu_inst_pe_1_1_2_add_69_carry_6_,
         npu_inst_pe_1_1_2_add_69_carry_5_, npu_inst_pe_1_1_2_add_69_carry_4_,
         npu_inst_pe_1_1_2_add_69_carry_3_, npu_inst_pe_1_1_2_add_69_carry_2_,
         npu_inst_pe_1_1_2_add_69_carry_1_, npu_inst_pe_1_1_2_n97,
         npu_inst_pe_1_1_2_n96, npu_inst_pe_1_1_2_n95, npu_inst_pe_1_1_2_n94,
         npu_inst_pe_1_1_2_n93, npu_inst_pe_1_1_2_n92, npu_inst_pe_1_1_2_n91,
         npu_inst_pe_1_1_2_n90, npu_inst_pe_1_1_2_n89, npu_inst_pe_1_1_2_n88,
         npu_inst_pe_1_1_2_n87, npu_inst_pe_1_1_2_n86, npu_inst_pe_1_1_2_n85,
         npu_inst_pe_1_1_2_n84, npu_inst_pe_1_1_2_n83, npu_inst_pe_1_1_2_n82,
         npu_inst_pe_1_1_2_n81, npu_inst_pe_1_1_2_n80, npu_inst_pe_1_1_2_n79,
         npu_inst_pe_1_1_2_n78, npu_inst_pe_1_1_2_n77, npu_inst_pe_1_1_2_n76,
         npu_inst_pe_1_1_2_n75, npu_inst_pe_1_1_2_n74, npu_inst_pe_1_1_2_n73,
         npu_inst_pe_1_1_2_n72, npu_inst_pe_1_1_2_n71, npu_inst_pe_1_1_2_n70,
         npu_inst_pe_1_1_2_n69, npu_inst_pe_1_1_2_n68, npu_inst_pe_1_1_2_n67,
         npu_inst_pe_1_1_2_n66, npu_inst_pe_1_1_2_n65, npu_inst_pe_1_1_2_n64,
         npu_inst_pe_1_1_2_n63, npu_inst_pe_1_1_2_n62, npu_inst_pe_1_1_2_n61,
         npu_inst_pe_1_1_2_n60, npu_inst_pe_1_1_2_n59, npu_inst_pe_1_1_2_n58,
         npu_inst_pe_1_1_2_n57, npu_inst_pe_1_1_2_n56, npu_inst_pe_1_1_2_n55,
         npu_inst_pe_1_1_2_n54, npu_inst_pe_1_1_2_n53, npu_inst_pe_1_1_2_n52,
         npu_inst_pe_1_1_2_n51, npu_inst_pe_1_1_2_n50, npu_inst_pe_1_1_2_n49,
         npu_inst_pe_1_1_2_n48, npu_inst_pe_1_1_2_n47, npu_inst_pe_1_1_2_n46,
         npu_inst_pe_1_1_2_n45, npu_inst_pe_1_1_2_n44, npu_inst_pe_1_1_2_n43,
         npu_inst_pe_1_1_2_n42, npu_inst_pe_1_1_2_n41, npu_inst_pe_1_1_2_n40,
         npu_inst_pe_1_1_2_n39, npu_inst_pe_1_1_2_n38, npu_inst_pe_1_1_2_n37,
         npu_inst_pe_1_1_2_n27, npu_inst_pe_1_1_2_n26,
         npu_inst_pe_1_1_2_net4338, npu_inst_pe_1_1_2_net4332,
         npu_inst_pe_1_1_2_N94, npu_inst_pe_1_1_2_N93, npu_inst_pe_1_1_2_N84,
         npu_inst_pe_1_1_2_N80, npu_inst_pe_1_1_2_N79, npu_inst_pe_1_1_2_N78,
         npu_inst_pe_1_1_2_N77, npu_inst_pe_1_1_2_N76, npu_inst_pe_1_1_2_N75,
         npu_inst_pe_1_1_2_N74, npu_inst_pe_1_1_2_N73, npu_inst_pe_1_1_2_N72,
         npu_inst_pe_1_1_2_N71, npu_inst_pe_1_1_2_N70, npu_inst_pe_1_1_2_N69,
         npu_inst_pe_1_1_2_N68, npu_inst_pe_1_1_2_N67, npu_inst_pe_1_1_2_N66,
         npu_inst_pe_1_1_2_N65, npu_inst_pe_1_1_2_int_q_acc_0_,
         npu_inst_pe_1_1_2_int_q_acc_1_, npu_inst_pe_1_1_2_int_q_acc_2_,
         npu_inst_pe_1_1_2_int_q_acc_3_, npu_inst_pe_1_1_2_int_q_acc_4_,
         npu_inst_pe_1_1_2_int_q_acc_5_, npu_inst_pe_1_1_2_int_q_acc_6_,
         npu_inst_pe_1_1_2_int_q_acc_7_, npu_inst_pe_1_1_2_int_data_0_,
         npu_inst_pe_1_1_2_int_data_1_, npu_inst_pe_1_1_2_int_q_weight_0_,
         npu_inst_pe_1_1_2_int_q_weight_1_,
         npu_inst_pe_1_1_2_int_q_reg_v_5__0_,
         npu_inst_pe_1_1_2_int_q_reg_v_5__1_,
         npu_inst_pe_1_1_2_int_q_reg_v_4__0_,
         npu_inst_pe_1_1_2_int_q_reg_v_4__1_,
         npu_inst_pe_1_1_2_int_q_reg_v_3__0_,
         npu_inst_pe_1_1_2_int_q_reg_v_3__1_,
         npu_inst_pe_1_1_2_int_q_reg_v_2__0_,
         npu_inst_pe_1_1_2_int_q_reg_v_2__1_,
         npu_inst_pe_1_1_2_int_q_reg_v_1__0_,
         npu_inst_pe_1_1_2_int_q_reg_v_1__1_,
         npu_inst_pe_1_1_2_int_q_reg_v_0__0_,
         npu_inst_pe_1_1_2_int_q_reg_v_0__1_,
         npu_inst_pe_1_1_2_int_q_reg_h_5__0_,
         npu_inst_pe_1_1_2_int_q_reg_h_5__1_,
         npu_inst_pe_1_1_2_int_q_reg_h_4__0_,
         npu_inst_pe_1_1_2_int_q_reg_h_4__1_,
         npu_inst_pe_1_1_2_int_q_reg_h_3__0_,
         npu_inst_pe_1_1_2_int_q_reg_h_3__1_,
         npu_inst_pe_1_1_2_int_q_reg_h_2__0_,
         npu_inst_pe_1_1_2_int_q_reg_h_2__1_,
         npu_inst_pe_1_1_2_int_q_reg_h_1__0_,
         npu_inst_pe_1_1_2_int_q_reg_h_1__1_,
         npu_inst_pe_1_1_2_int_q_reg_h_0__0_,
         npu_inst_pe_1_1_2_int_q_reg_h_0__1_, npu_inst_pe_1_1_3_n119,
         npu_inst_pe_1_1_3_n118, npu_inst_pe_1_1_3_n117,
         npu_inst_pe_1_1_3_n116, npu_inst_pe_1_1_3_n115,
         npu_inst_pe_1_1_3_n114, npu_inst_pe_1_1_3_n113,
         npu_inst_pe_1_1_3_n112, npu_inst_pe_1_1_3_n111,
         npu_inst_pe_1_1_3_n110, npu_inst_pe_1_1_3_n109,
         npu_inst_pe_1_1_3_n108, npu_inst_pe_1_1_3_n107,
         npu_inst_pe_1_1_3_n106, npu_inst_pe_1_1_3_n105,
         npu_inst_pe_1_1_3_n104, npu_inst_pe_1_1_3_n103,
         npu_inst_pe_1_1_3_n102, npu_inst_pe_1_1_3_n101,
         npu_inst_pe_1_1_3_n100, npu_inst_pe_1_1_3_n99, npu_inst_pe_1_1_3_n98,
         npu_inst_pe_1_1_3_n36, npu_inst_pe_1_1_3_n35, npu_inst_pe_1_1_3_n34,
         npu_inst_pe_1_1_3_n33, npu_inst_pe_1_1_3_n32, npu_inst_pe_1_1_3_n31,
         npu_inst_pe_1_1_3_n30, npu_inst_pe_1_1_3_n29, npu_inst_pe_1_1_3_n28,
         npu_inst_pe_1_1_3_n25, npu_inst_pe_1_1_3_n24, npu_inst_pe_1_1_3_n23,
         npu_inst_pe_1_1_3_n22, npu_inst_pe_1_1_3_n21, npu_inst_pe_1_1_3_n20,
         npu_inst_pe_1_1_3_n19, npu_inst_pe_1_1_3_n18, npu_inst_pe_1_1_3_n17,
         npu_inst_pe_1_1_3_n16, npu_inst_pe_1_1_3_n15, npu_inst_pe_1_1_3_n14,
         npu_inst_pe_1_1_3_n13, npu_inst_pe_1_1_3_n12, npu_inst_pe_1_1_3_n11,
         npu_inst_pe_1_1_3_n10, npu_inst_pe_1_1_3_n9, npu_inst_pe_1_1_3_n8,
         npu_inst_pe_1_1_3_n7, npu_inst_pe_1_1_3_n6, npu_inst_pe_1_1_3_n5,
         npu_inst_pe_1_1_3_n4, npu_inst_pe_1_1_3_n3, npu_inst_pe_1_1_3_n2,
         npu_inst_pe_1_1_3_n1, npu_inst_pe_1_1_3_sub_67_carry_7_,
         npu_inst_pe_1_1_3_sub_67_carry_6_, npu_inst_pe_1_1_3_sub_67_carry_5_,
         npu_inst_pe_1_1_3_sub_67_carry_4_, npu_inst_pe_1_1_3_sub_67_carry_3_,
         npu_inst_pe_1_1_3_sub_67_carry_2_, npu_inst_pe_1_1_3_sub_67_carry_1_,
         npu_inst_pe_1_1_3_add_69_carry_7_, npu_inst_pe_1_1_3_add_69_carry_6_,
         npu_inst_pe_1_1_3_add_69_carry_5_, npu_inst_pe_1_1_3_add_69_carry_4_,
         npu_inst_pe_1_1_3_add_69_carry_3_, npu_inst_pe_1_1_3_add_69_carry_2_,
         npu_inst_pe_1_1_3_add_69_carry_1_, npu_inst_pe_1_1_3_n97,
         npu_inst_pe_1_1_3_n96, npu_inst_pe_1_1_3_n95, npu_inst_pe_1_1_3_n94,
         npu_inst_pe_1_1_3_n93, npu_inst_pe_1_1_3_n92, npu_inst_pe_1_1_3_n91,
         npu_inst_pe_1_1_3_n90, npu_inst_pe_1_1_3_n89, npu_inst_pe_1_1_3_n88,
         npu_inst_pe_1_1_3_n87, npu_inst_pe_1_1_3_n86, npu_inst_pe_1_1_3_n85,
         npu_inst_pe_1_1_3_n84, npu_inst_pe_1_1_3_n83, npu_inst_pe_1_1_3_n82,
         npu_inst_pe_1_1_3_n81, npu_inst_pe_1_1_3_n80, npu_inst_pe_1_1_3_n79,
         npu_inst_pe_1_1_3_n78, npu_inst_pe_1_1_3_n77, npu_inst_pe_1_1_3_n76,
         npu_inst_pe_1_1_3_n75, npu_inst_pe_1_1_3_n74, npu_inst_pe_1_1_3_n73,
         npu_inst_pe_1_1_3_n72, npu_inst_pe_1_1_3_n71, npu_inst_pe_1_1_3_n70,
         npu_inst_pe_1_1_3_n69, npu_inst_pe_1_1_3_n68, npu_inst_pe_1_1_3_n67,
         npu_inst_pe_1_1_3_n66, npu_inst_pe_1_1_3_n65, npu_inst_pe_1_1_3_n64,
         npu_inst_pe_1_1_3_n63, npu_inst_pe_1_1_3_n62, npu_inst_pe_1_1_3_n61,
         npu_inst_pe_1_1_3_n60, npu_inst_pe_1_1_3_n59, npu_inst_pe_1_1_3_n58,
         npu_inst_pe_1_1_3_n57, npu_inst_pe_1_1_3_n56, npu_inst_pe_1_1_3_n55,
         npu_inst_pe_1_1_3_n54, npu_inst_pe_1_1_3_n53, npu_inst_pe_1_1_3_n52,
         npu_inst_pe_1_1_3_n51, npu_inst_pe_1_1_3_n50, npu_inst_pe_1_1_3_n49,
         npu_inst_pe_1_1_3_n48, npu_inst_pe_1_1_3_n47, npu_inst_pe_1_1_3_n46,
         npu_inst_pe_1_1_3_n45, npu_inst_pe_1_1_3_n44, npu_inst_pe_1_1_3_n43,
         npu_inst_pe_1_1_3_n42, npu_inst_pe_1_1_3_n41, npu_inst_pe_1_1_3_n40,
         npu_inst_pe_1_1_3_n39, npu_inst_pe_1_1_3_n38, npu_inst_pe_1_1_3_n37,
         npu_inst_pe_1_1_3_n27, npu_inst_pe_1_1_3_n26,
         npu_inst_pe_1_1_3_net4315, npu_inst_pe_1_1_3_net4309,
         npu_inst_pe_1_1_3_N94, npu_inst_pe_1_1_3_N93, npu_inst_pe_1_1_3_N84,
         npu_inst_pe_1_1_3_N80, npu_inst_pe_1_1_3_N79, npu_inst_pe_1_1_3_N78,
         npu_inst_pe_1_1_3_N77, npu_inst_pe_1_1_3_N76, npu_inst_pe_1_1_3_N75,
         npu_inst_pe_1_1_3_N74, npu_inst_pe_1_1_3_N73, npu_inst_pe_1_1_3_N72,
         npu_inst_pe_1_1_3_N71, npu_inst_pe_1_1_3_N70, npu_inst_pe_1_1_3_N69,
         npu_inst_pe_1_1_3_N68, npu_inst_pe_1_1_3_N67, npu_inst_pe_1_1_3_N66,
         npu_inst_pe_1_1_3_N65, npu_inst_pe_1_1_3_int_q_acc_0_,
         npu_inst_pe_1_1_3_int_q_acc_1_, npu_inst_pe_1_1_3_int_q_acc_2_,
         npu_inst_pe_1_1_3_int_q_acc_3_, npu_inst_pe_1_1_3_int_q_acc_4_,
         npu_inst_pe_1_1_3_int_q_acc_5_, npu_inst_pe_1_1_3_int_q_acc_6_,
         npu_inst_pe_1_1_3_int_q_acc_7_, npu_inst_pe_1_1_3_int_data_0_,
         npu_inst_pe_1_1_3_int_data_1_, npu_inst_pe_1_1_3_int_q_weight_0_,
         npu_inst_pe_1_1_3_int_q_weight_1_,
         npu_inst_pe_1_1_3_int_q_reg_v_5__0_,
         npu_inst_pe_1_1_3_int_q_reg_v_5__1_,
         npu_inst_pe_1_1_3_int_q_reg_v_4__0_,
         npu_inst_pe_1_1_3_int_q_reg_v_4__1_,
         npu_inst_pe_1_1_3_int_q_reg_v_3__0_,
         npu_inst_pe_1_1_3_int_q_reg_v_3__1_,
         npu_inst_pe_1_1_3_int_q_reg_v_2__0_,
         npu_inst_pe_1_1_3_int_q_reg_v_2__1_,
         npu_inst_pe_1_1_3_int_q_reg_v_1__0_,
         npu_inst_pe_1_1_3_int_q_reg_v_1__1_,
         npu_inst_pe_1_1_3_int_q_reg_v_0__0_,
         npu_inst_pe_1_1_3_int_q_reg_v_0__1_,
         npu_inst_pe_1_1_3_int_q_reg_h_5__0_,
         npu_inst_pe_1_1_3_int_q_reg_h_5__1_,
         npu_inst_pe_1_1_3_int_q_reg_h_4__0_,
         npu_inst_pe_1_1_3_int_q_reg_h_4__1_,
         npu_inst_pe_1_1_3_int_q_reg_h_3__0_,
         npu_inst_pe_1_1_3_int_q_reg_h_3__1_,
         npu_inst_pe_1_1_3_int_q_reg_h_2__0_,
         npu_inst_pe_1_1_3_int_q_reg_h_2__1_,
         npu_inst_pe_1_1_3_int_q_reg_h_1__0_,
         npu_inst_pe_1_1_3_int_q_reg_h_1__1_,
         npu_inst_pe_1_1_3_int_q_reg_h_0__0_,
         npu_inst_pe_1_1_3_int_q_reg_h_0__1_, npu_inst_pe_1_1_4_n119,
         npu_inst_pe_1_1_4_n118, npu_inst_pe_1_1_4_n117,
         npu_inst_pe_1_1_4_n116, npu_inst_pe_1_1_4_n115,
         npu_inst_pe_1_1_4_n114, npu_inst_pe_1_1_4_n113,
         npu_inst_pe_1_1_4_n112, npu_inst_pe_1_1_4_n111,
         npu_inst_pe_1_1_4_n110, npu_inst_pe_1_1_4_n109,
         npu_inst_pe_1_1_4_n108, npu_inst_pe_1_1_4_n107,
         npu_inst_pe_1_1_4_n106, npu_inst_pe_1_1_4_n105,
         npu_inst_pe_1_1_4_n104, npu_inst_pe_1_1_4_n103,
         npu_inst_pe_1_1_4_n102, npu_inst_pe_1_1_4_n101,
         npu_inst_pe_1_1_4_n100, npu_inst_pe_1_1_4_n99, npu_inst_pe_1_1_4_n98,
         npu_inst_pe_1_1_4_n36, npu_inst_pe_1_1_4_n35, npu_inst_pe_1_1_4_n34,
         npu_inst_pe_1_1_4_n33, npu_inst_pe_1_1_4_n32, npu_inst_pe_1_1_4_n31,
         npu_inst_pe_1_1_4_n30, npu_inst_pe_1_1_4_n29, npu_inst_pe_1_1_4_n28,
         npu_inst_pe_1_1_4_n25, npu_inst_pe_1_1_4_n24, npu_inst_pe_1_1_4_n23,
         npu_inst_pe_1_1_4_n22, npu_inst_pe_1_1_4_n21, npu_inst_pe_1_1_4_n20,
         npu_inst_pe_1_1_4_n19, npu_inst_pe_1_1_4_n18, npu_inst_pe_1_1_4_n17,
         npu_inst_pe_1_1_4_n16, npu_inst_pe_1_1_4_n15, npu_inst_pe_1_1_4_n14,
         npu_inst_pe_1_1_4_n13, npu_inst_pe_1_1_4_n12, npu_inst_pe_1_1_4_n11,
         npu_inst_pe_1_1_4_n10, npu_inst_pe_1_1_4_n9, npu_inst_pe_1_1_4_n8,
         npu_inst_pe_1_1_4_n7, npu_inst_pe_1_1_4_n6, npu_inst_pe_1_1_4_n5,
         npu_inst_pe_1_1_4_n4, npu_inst_pe_1_1_4_n3, npu_inst_pe_1_1_4_n2,
         npu_inst_pe_1_1_4_n1, npu_inst_pe_1_1_4_sub_67_carry_7_,
         npu_inst_pe_1_1_4_sub_67_carry_6_, npu_inst_pe_1_1_4_sub_67_carry_5_,
         npu_inst_pe_1_1_4_sub_67_carry_4_, npu_inst_pe_1_1_4_sub_67_carry_3_,
         npu_inst_pe_1_1_4_sub_67_carry_2_, npu_inst_pe_1_1_4_sub_67_carry_1_,
         npu_inst_pe_1_1_4_add_69_carry_7_, npu_inst_pe_1_1_4_add_69_carry_6_,
         npu_inst_pe_1_1_4_add_69_carry_5_, npu_inst_pe_1_1_4_add_69_carry_4_,
         npu_inst_pe_1_1_4_add_69_carry_3_, npu_inst_pe_1_1_4_add_69_carry_2_,
         npu_inst_pe_1_1_4_add_69_carry_1_, npu_inst_pe_1_1_4_n97,
         npu_inst_pe_1_1_4_n96, npu_inst_pe_1_1_4_n95, npu_inst_pe_1_1_4_n94,
         npu_inst_pe_1_1_4_n93, npu_inst_pe_1_1_4_n92, npu_inst_pe_1_1_4_n91,
         npu_inst_pe_1_1_4_n90, npu_inst_pe_1_1_4_n89, npu_inst_pe_1_1_4_n88,
         npu_inst_pe_1_1_4_n87, npu_inst_pe_1_1_4_n86, npu_inst_pe_1_1_4_n85,
         npu_inst_pe_1_1_4_n84, npu_inst_pe_1_1_4_n83, npu_inst_pe_1_1_4_n82,
         npu_inst_pe_1_1_4_n81, npu_inst_pe_1_1_4_n80, npu_inst_pe_1_1_4_n79,
         npu_inst_pe_1_1_4_n78, npu_inst_pe_1_1_4_n77, npu_inst_pe_1_1_4_n76,
         npu_inst_pe_1_1_4_n75, npu_inst_pe_1_1_4_n74, npu_inst_pe_1_1_4_n73,
         npu_inst_pe_1_1_4_n72, npu_inst_pe_1_1_4_n71, npu_inst_pe_1_1_4_n70,
         npu_inst_pe_1_1_4_n69, npu_inst_pe_1_1_4_n68, npu_inst_pe_1_1_4_n67,
         npu_inst_pe_1_1_4_n66, npu_inst_pe_1_1_4_n65, npu_inst_pe_1_1_4_n64,
         npu_inst_pe_1_1_4_n63, npu_inst_pe_1_1_4_n62, npu_inst_pe_1_1_4_n61,
         npu_inst_pe_1_1_4_n60, npu_inst_pe_1_1_4_n59, npu_inst_pe_1_1_4_n58,
         npu_inst_pe_1_1_4_n57, npu_inst_pe_1_1_4_n56, npu_inst_pe_1_1_4_n55,
         npu_inst_pe_1_1_4_n54, npu_inst_pe_1_1_4_n53, npu_inst_pe_1_1_4_n52,
         npu_inst_pe_1_1_4_n51, npu_inst_pe_1_1_4_n50, npu_inst_pe_1_1_4_n49,
         npu_inst_pe_1_1_4_n48, npu_inst_pe_1_1_4_n47, npu_inst_pe_1_1_4_n46,
         npu_inst_pe_1_1_4_n45, npu_inst_pe_1_1_4_n44, npu_inst_pe_1_1_4_n43,
         npu_inst_pe_1_1_4_n42, npu_inst_pe_1_1_4_n41, npu_inst_pe_1_1_4_n40,
         npu_inst_pe_1_1_4_n39, npu_inst_pe_1_1_4_n38, npu_inst_pe_1_1_4_n37,
         npu_inst_pe_1_1_4_n27, npu_inst_pe_1_1_4_n26,
         npu_inst_pe_1_1_4_net4292, npu_inst_pe_1_1_4_net4286,
         npu_inst_pe_1_1_4_N94, npu_inst_pe_1_1_4_N93, npu_inst_pe_1_1_4_N84,
         npu_inst_pe_1_1_4_N80, npu_inst_pe_1_1_4_N79, npu_inst_pe_1_1_4_N78,
         npu_inst_pe_1_1_4_N77, npu_inst_pe_1_1_4_N76, npu_inst_pe_1_1_4_N75,
         npu_inst_pe_1_1_4_N74, npu_inst_pe_1_1_4_N73, npu_inst_pe_1_1_4_N72,
         npu_inst_pe_1_1_4_N71, npu_inst_pe_1_1_4_N70, npu_inst_pe_1_1_4_N69,
         npu_inst_pe_1_1_4_N68, npu_inst_pe_1_1_4_N67, npu_inst_pe_1_1_4_N66,
         npu_inst_pe_1_1_4_N65, npu_inst_pe_1_1_4_int_q_acc_0_,
         npu_inst_pe_1_1_4_int_q_acc_1_, npu_inst_pe_1_1_4_int_q_acc_2_,
         npu_inst_pe_1_1_4_int_q_acc_3_, npu_inst_pe_1_1_4_int_q_acc_4_,
         npu_inst_pe_1_1_4_int_q_acc_5_, npu_inst_pe_1_1_4_int_q_acc_6_,
         npu_inst_pe_1_1_4_int_q_acc_7_, npu_inst_pe_1_1_4_int_data_0_,
         npu_inst_pe_1_1_4_int_data_1_, npu_inst_pe_1_1_4_int_q_weight_0_,
         npu_inst_pe_1_1_4_int_q_weight_1_,
         npu_inst_pe_1_1_4_int_q_reg_v_5__0_,
         npu_inst_pe_1_1_4_int_q_reg_v_5__1_,
         npu_inst_pe_1_1_4_int_q_reg_v_4__0_,
         npu_inst_pe_1_1_4_int_q_reg_v_4__1_,
         npu_inst_pe_1_1_4_int_q_reg_v_3__0_,
         npu_inst_pe_1_1_4_int_q_reg_v_3__1_,
         npu_inst_pe_1_1_4_int_q_reg_v_2__0_,
         npu_inst_pe_1_1_4_int_q_reg_v_2__1_,
         npu_inst_pe_1_1_4_int_q_reg_v_1__0_,
         npu_inst_pe_1_1_4_int_q_reg_v_1__1_,
         npu_inst_pe_1_1_4_int_q_reg_v_0__0_,
         npu_inst_pe_1_1_4_int_q_reg_v_0__1_,
         npu_inst_pe_1_1_4_int_q_reg_h_5__0_,
         npu_inst_pe_1_1_4_int_q_reg_h_5__1_,
         npu_inst_pe_1_1_4_int_q_reg_h_4__0_,
         npu_inst_pe_1_1_4_int_q_reg_h_4__1_,
         npu_inst_pe_1_1_4_int_q_reg_h_3__0_,
         npu_inst_pe_1_1_4_int_q_reg_h_3__1_,
         npu_inst_pe_1_1_4_int_q_reg_h_2__0_,
         npu_inst_pe_1_1_4_int_q_reg_h_2__1_,
         npu_inst_pe_1_1_4_int_q_reg_h_1__0_,
         npu_inst_pe_1_1_4_int_q_reg_h_1__1_,
         npu_inst_pe_1_1_4_int_q_reg_h_0__0_,
         npu_inst_pe_1_1_4_int_q_reg_h_0__1_, npu_inst_pe_1_1_5_n119,
         npu_inst_pe_1_1_5_n118, npu_inst_pe_1_1_5_n117,
         npu_inst_pe_1_1_5_n116, npu_inst_pe_1_1_5_n115,
         npu_inst_pe_1_1_5_n114, npu_inst_pe_1_1_5_n113,
         npu_inst_pe_1_1_5_n112, npu_inst_pe_1_1_5_n111,
         npu_inst_pe_1_1_5_n110, npu_inst_pe_1_1_5_n109,
         npu_inst_pe_1_1_5_n108, npu_inst_pe_1_1_5_n107,
         npu_inst_pe_1_1_5_n106, npu_inst_pe_1_1_5_n105,
         npu_inst_pe_1_1_5_n104, npu_inst_pe_1_1_5_n103,
         npu_inst_pe_1_1_5_n102, npu_inst_pe_1_1_5_n101,
         npu_inst_pe_1_1_5_n100, npu_inst_pe_1_1_5_n99, npu_inst_pe_1_1_5_n98,
         npu_inst_pe_1_1_5_n36, npu_inst_pe_1_1_5_n35, npu_inst_pe_1_1_5_n34,
         npu_inst_pe_1_1_5_n33, npu_inst_pe_1_1_5_n32, npu_inst_pe_1_1_5_n31,
         npu_inst_pe_1_1_5_n30, npu_inst_pe_1_1_5_n29, npu_inst_pe_1_1_5_n28,
         npu_inst_pe_1_1_5_n25, npu_inst_pe_1_1_5_n24, npu_inst_pe_1_1_5_n23,
         npu_inst_pe_1_1_5_n22, npu_inst_pe_1_1_5_n21, npu_inst_pe_1_1_5_n20,
         npu_inst_pe_1_1_5_n19, npu_inst_pe_1_1_5_n18, npu_inst_pe_1_1_5_n17,
         npu_inst_pe_1_1_5_n16, npu_inst_pe_1_1_5_n15, npu_inst_pe_1_1_5_n14,
         npu_inst_pe_1_1_5_n13, npu_inst_pe_1_1_5_n12, npu_inst_pe_1_1_5_n11,
         npu_inst_pe_1_1_5_n10, npu_inst_pe_1_1_5_n9, npu_inst_pe_1_1_5_n8,
         npu_inst_pe_1_1_5_n7, npu_inst_pe_1_1_5_n6, npu_inst_pe_1_1_5_n5,
         npu_inst_pe_1_1_5_n4, npu_inst_pe_1_1_5_n3, npu_inst_pe_1_1_5_n2,
         npu_inst_pe_1_1_5_n1, npu_inst_pe_1_1_5_sub_67_carry_7_,
         npu_inst_pe_1_1_5_sub_67_carry_6_, npu_inst_pe_1_1_5_sub_67_carry_5_,
         npu_inst_pe_1_1_5_sub_67_carry_4_, npu_inst_pe_1_1_5_sub_67_carry_3_,
         npu_inst_pe_1_1_5_sub_67_carry_2_, npu_inst_pe_1_1_5_sub_67_carry_1_,
         npu_inst_pe_1_1_5_add_69_carry_7_, npu_inst_pe_1_1_5_add_69_carry_6_,
         npu_inst_pe_1_1_5_add_69_carry_5_, npu_inst_pe_1_1_5_add_69_carry_4_,
         npu_inst_pe_1_1_5_add_69_carry_3_, npu_inst_pe_1_1_5_add_69_carry_2_,
         npu_inst_pe_1_1_5_add_69_carry_1_, npu_inst_pe_1_1_5_n97,
         npu_inst_pe_1_1_5_n96, npu_inst_pe_1_1_5_n95, npu_inst_pe_1_1_5_n94,
         npu_inst_pe_1_1_5_n93, npu_inst_pe_1_1_5_n92, npu_inst_pe_1_1_5_n91,
         npu_inst_pe_1_1_5_n90, npu_inst_pe_1_1_5_n89, npu_inst_pe_1_1_5_n88,
         npu_inst_pe_1_1_5_n87, npu_inst_pe_1_1_5_n86, npu_inst_pe_1_1_5_n85,
         npu_inst_pe_1_1_5_n84, npu_inst_pe_1_1_5_n83, npu_inst_pe_1_1_5_n82,
         npu_inst_pe_1_1_5_n81, npu_inst_pe_1_1_5_n80, npu_inst_pe_1_1_5_n79,
         npu_inst_pe_1_1_5_n78, npu_inst_pe_1_1_5_n77, npu_inst_pe_1_1_5_n76,
         npu_inst_pe_1_1_5_n75, npu_inst_pe_1_1_5_n74, npu_inst_pe_1_1_5_n73,
         npu_inst_pe_1_1_5_n72, npu_inst_pe_1_1_5_n71, npu_inst_pe_1_1_5_n70,
         npu_inst_pe_1_1_5_n69, npu_inst_pe_1_1_5_n68, npu_inst_pe_1_1_5_n67,
         npu_inst_pe_1_1_5_n66, npu_inst_pe_1_1_5_n65, npu_inst_pe_1_1_5_n64,
         npu_inst_pe_1_1_5_n63, npu_inst_pe_1_1_5_n62, npu_inst_pe_1_1_5_n61,
         npu_inst_pe_1_1_5_n60, npu_inst_pe_1_1_5_n59, npu_inst_pe_1_1_5_n58,
         npu_inst_pe_1_1_5_n57, npu_inst_pe_1_1_5_n56, npu_inst_pe_1_1_5_n55,
         npu_inst_pe_1_1_5_n54, npu_inst_pe_1_1_5_n53, npu_inst_pe_1_1_5_n52,
         npu_inst_pe_1_1_5_n51, npu_inst_pe_1_1_5_n50, npu_inst_pe_1_1_5_n49,
         npu_inst_pe_1_1_5_n48, npu_inst_pe_1_1_5_n47, npu_inst_pe_1_1_5_n46,
         npu_inst_pe_1_1_5_n45, npu_inst_pe_1_1_5_n44, npu_inst_pe_1_1_5_n43,
         npu_inst_pe_1_1_5_n42, npu_inst_pe_1_1_5_n41, npu_inst_pe_1_1_5_n40,
         npu_inst_pe_1_1_5_n39, npu_inst_pe_1_1_5_n38, npu_inst_pe_1_1_5_n37,
         npu_inst_pe_1_1_5_n27, npu_inst_pe_1_1_5_n26,
         npu_inst_pe_1_1_5_net4269, npu_inst_pe_1_1_5_net4263,
         npu_inst_pe_1_1_5_N94, npu_inst_pe_1_1_5_N93, npu_inst_pe_1_1_5_N84,
         npu_inst_pe_1_1_5_N80, npu_inst_pe_1_1_5_N79, npu_inst_pe_1_1_5_N78,
         npu_inst_pe_1_1_5_N77, npu_inst_pe_1_1_5_N76, npu_inst_pe_1_1_5_N75,
         npu_inst_pe_1_1_5_N74, npu_inst_pe_1_1_5_N73, npu_inst_pe_1_1_5_N72,
         npu_inst_pe_1_1_5_N71, npu_inst_pe_1_1_5_N70, npu_inst_pe_1_1_5_N69,
         npu_inst_pe_1_1_5_N68, npu_inst_pe_1_1_5_N67, npu_inst_pe_1_1_5_N66,
         npu_inst_pe_1_1_5_N65, npu_inst_pe_1_1_5_int_q_acc_0_,
         npu_inst_pe_1_1_5_int_q_acc_1_, npu_inst_pe_1_1_5_int_q_acc_2_,
         npu_inst_pe_1_1_5_int_q_acc_3_, npu_inst_pe_1_1_5_int_q_acc_4_,
         npu_inst_pe_1_1_5_int_q_acc_5_, npu_inst_pe_1_1_5_int_q_acc_6_,
         npu_inst_pe_1_1_5_int_q_acc_7_, npu_inst_pe_1_1_5_int_data_0_,
         npu_inst_pe_1_1_5_int_data_1_, npu_inst_pe_1_1_5_int_q_weight_0_,
         npu_inst_pe_1_1_5_int_q_weight_1_,
         npu_inst_pe_1_1_5_int_q_reg_v_5__0_,
         npu_inst_pe_1_1_5_int_q_reg_v_5__1_,
         npu_inst_pe_1_1_5_int_q_reg_v_4__0_,
         npu_inst_pe_1_1_5_int_q_reg_v_4__1_,
         npu_inst_pe_1_1_5_int_q_reg_v_3__0_,
         npu_inst_pe_1_1_5_int_q_reg_v_3__1_,
         npu_inst_pe_1_1_5_int_q_reg_v_2__0_,
         npu_inst_pe_1_1_5_int_q_reg_v_2__1_,
         npu_inst_pe_1_1_5_int_q_reg_v_1__0_,
         npu_inst_pe_1_1_5_int_q_reg_v_1__1_,
         npu_inst_pe_1_1_5_int_q_reg_v_0__0_,
         npu_inst_pe_1_1_5_int_q_reg_v_0__1_,
         npu_inst_pe_1_1_5_int_q_reg_h_5__0_,
         npu_inst_pe_1_1_5_int_q_reg_h_5__1_,
         npu_inst_pe_1_1_5_int_q_reg_h_4__0_,
         npu_inst_pe_1_1_5_int_q_reg_h_4__1_,
         npu_inst_pe_1_1_5_int_q_reg_h_3__0_,
         npu_inst_pe_1_1_5_int_q_reg_h_3__1_,
         npu_inst_pe_1_1_5_int_q_reg_h_2__0_,
         npu_inst_pe_1_1_5_int_q_reg_h_2__1_,
         npu_inst_pe_1_1_5_int_q_reg_h_1__0_,
         npu_inst_pe_1_1_5_int_q_reg_h_1__1_,
         npu_inst_pe_1_1_5_int_q_reg_h_0__0_,
         npu_inst_pe_1_1_5_int_q_reg_h_0__1_, npu_inst_pe_1_1_6_n119,
         npu_inst_pe_1_1_6_n118, npu_inst_pe_1_1_6_n117,
         npu_inst_pe_1_1_6_n116, npu_inst_pe_1_1_6_n115,
         npu_inst_pe_1_1_6_n114, npu_inst_pe_1_1_6_n113,
         npu_inst_pe_1_1_6_n112, npu_inst_pe_1_1_6_n111,
         npu_inst_pe_1_1_6_n110, npu_inst_pe_1_1_6_n109,
         npu_inst_pe_1_1_6_n108, npu_inst_pe_1_1_6_n107,
         npu_inst_pe_1_1_6_n106, npu_inst_pe_1_1_6_n105,
         npu_inst_pe_1_1_6_n104, npu_inst_pe_1_1_6_n103,
         npu_inst_pe_1_1_6_n102, npu_inst_pe_1_1_6_n101,
         npu_inst_pe_1_1_6_n100, npu_inst_pe_1_1_6_n99, npu_inst_pe_1_1_6_n98,
         npu_inst_pe_1_1_6_n36, npu_inst_pe_1_1_6_n35, npu_inst_pe_1_1_6_n34,
         npu_inst_pe_1_1_6_n33, npu_inst_pe_1_1_6_n32, npu_inst_pe_1_1_6_n31,
         npu_inst_pe_1_1_6_n30, npu_inst_pe_1_1_6_n29, npu_inst_pe_1_1_6_n28,
         npu_inst_pe_1_1_6_n25, npu_inst_pe_1_1_6_n24, npu_inst_pe_1_1_6_n23,
         npu_inst_pe_1_1_6_n22, npu_inst_pe_1_1_6_n21, npu_inst_pe_1_1_6_n20,
         npu_inst_pe_1_1_6_n19, npu_inst_pe_1_1_6_n18, npu_inst_pe_1_1_6_n17,
         npu_inst_pe_1_1_6_n16, npu_inst_pe_1_1_6_n15, npu_inst_pe_1_1_6_n14,
         npu_inst_pe_1_1_6_n13, npu_inst_pe_1_1_6_n12, npu_inst_pe_1_1_6_n11,
         npu_inst_pe_1_1_6_n10, npu_inst_pe_1_1_6_n9, npu_inst_pe_1_1_6_n8,
         npu_inst_pe_1_1_6_n7, npu_inst_pe_1_1_6_n6, npu_inst_pe_1_1_6_n5,
         npu_inst_pe_1_1_6_n4, npu_inst_pe_1_1_6_n3, npu_inst_pe_1_1_6_n2,
         npu_inst_pe_1_1_6_n1, npu_inst_pe_1_1_6_sub_67_carry_7_,
         npu_inst_pe_1_1_6_sub_67_carry_6_, npu_inst_pe_1_1_6_sub_67_carry_5_,
         npu_inst_pe_1_1_6_sub_67_carry_4_, npu_inst_pe_1_1_6_sub_67_carry_3_,
         npu_inst_pe_1_1_6_sub_67_carry_2_, npu_inst_pe_1_1_6_sub_67_carry_1_,
         npu_inst_pe_1_1_6_add_69_carry_7_, npu_inst_pe_1_1_6_add_69_carry_6_,
         npu_inst_pe_1_1_6_add_69_carry_5_, npu_inst_pe_1_1_6_add_69_carry_4_,
         npu_inst_pe_1_1_6_add_69_carry_3_, npu_inst_pe_1_1_6_add_69_carry_2_,
         npu_inst_pe_1_1_6_add_69_carry_1_, npu_inst_pe_1_1_6_n97,
         npu_inst_pe_1_1_6_n96, npu_inst_pe_1_1_6_n95, npu_inst_pe_1_1_6_n94,
         npu_inst_pe_1_1_6_n93, npu_inst_pe_1_1_6_n92, npu_inst_pe_1_1_6_n91,
         npu_inst_pe_1_1_6_n90, npu_inst_pe_1_1_6_n89, npu_inst_pe_1_1_6_n88,
         npu_inst_pe_1_1_6_n87, npu_inst_pe_1_1_6_n86, npu_inst_pe_1_1_6_n85,
         npu_inst_pe_1_1_6_n84, npu_inst_pe_1_1_6_n83, npu_inst_pe_1_1_6_n82,
         npu_inst_pe_1_1_6_n81, npu_inst_pe_1_1_6_n80, npu_inst_pe_1_1_6_n79,
         npu_inst_pe_1_1_6_n78, npu_inst_pe_1_1_6_n77, npu_inst_pe_1_1_6_n76,
         npu_inst_pe_1_1_6_n75, npu_inst_pe_1_1_6_n74, npu_inst_pe_1_1_6_n73,
         npu_inst_pe_1_1_6_n72, npu_inst_pe_1_1_6_n71, npu_inst_pe_1_1_6_n70,
         npu_inst_pe_1_1_6_n69, npu_inst_pe_1_1_6_n68, npu_inst_pe_1_1_6_n67,
         npu_inst_pe_1_1_6_n66, npu_inst_pe_1_1_6_n65, npu_inst_pe_1_1_6_n64,
         npu_inst_pe_1_1_6_n63, npu_inst_pe_1_1_6_n62, npu_inst_pe_1_1_6_n61,
         npu_inst_pe_1_1_6_n60, npu_inst_pe_1_1_6_n59, npu_inst_pe_1_1_6_n58,
         npu_inst_pe_1_1_6_n57, npu_inst_pe_1_1_6_n56, npu_inst_pe_1_1_6_n55,
         npu_inst_pe_1_1_6_n54, npu_inst_pe_1_1_6_n53, npu_inst_pe_1_1_6_n52,
         npu_inst_pe_1_1_6_n51, npu_inst_pe_1_1_6_n50, npu_inst_pe_1_1_6_n49,
         npu_inst_pe_1_1_6_n48, npu_inst_pe_1_1_6_n47, npu_inst_pe_1_1_6_n46,
         npu_inst_pe_1_1_6_n45, npu_inst_pe_1_1_6_n44, npu_inst_pe_1_1_6_n43,
         npu_inst_pe_1_1_6_n42, npu_inst_pe_1_1_6_n41, npu_inst_pe_1_1_6_n40,
         npu_inst_pe_1_1_6_n39, npu_inst_pe_1_1_6_n38, npu_inst_pe_1_1_6_n37,
         npu_inst_pe_1_1_6_n27, npu_inst_pe_1_1_6_n26,
         npu_inst_pe_1_1_6_net4246, npu_inst_pe_1_1_6_net4240,
         npu_inst_pe_1_1_6_N94, npu_inst_pe_1_1_6_N93, npu_inst_pe_1_1_6_N84,
         npu_inst_pe_1_1_6_N80, npu_inst_pe_1_1_6_N79, npu_inst_pe_1_1_6_N78,
         npu_inst_pe_1_1_6_N77, npu_inst_pe_1_1_6_N76, npu_inst_pe_1_1_6_N75,
         npu_inst_pe_1_1_6_N74, npu_inst_pe_1_1_6_N73, npu_inst_pe_1_1_6_N72,
         npu_inst_pe_1_1_6_N71, npu_inst_pe_1_1_6_N70, npu_inst_pe_1_1_6_N69,
         npu_inst_pe_1_1_6_N68, npu_inst_pe_1_1_6_N67, npu_inst_pe_1_1_6_N66,
         npu_inst_pe_1_1_6_N65, npu_inst_pe_1_1_6_int_q_acc_0_,
         npu_inst_pe_1_1_6_int_q_acc_1_, npu_inst_pe_1_1_6_int_q_acc_2_,
         npu_inst_pe_1_1_6_int_q_acc_3_, npu_inst_pe_1_1_6_int_q_acc_4_,
         npu_inst_pe_1_1_6_int_q_acc_5_, npu_inst_pe_1_1_6_int_q_acc_6_,
         npu_inst_pe_1_1_6_int_q_acc_7_, npu_inst_pe_1_1_6_int_data_0_,
         npu_inst_pe_1_1_6_int_data_1_, npu_inst_pe_1_1_6_int_q_weight_0_,
         npu_inst_pe_1_1_6_int_q_weight_1_,
         npu_inst_pe_1_1_6_int_q_reg_v_5__0_,
         npu_inst_pe_1_1_6_int_q_reg_v_5__1_,
         npu_inst_pe_1_1_6_int_q_reg_v_4__0_,
         npu_inst_pe_1_1_6_int_q_reg_v_4__1_,
         npu_inst_pe_1_1_6_int_q_reg_v_3__0_,
         npu_inst_pe_1_1_6_int_q_reg_v_3__1_,
         npu_inst_pe_1_1_6_int_q_reg_v_2__0_,
         npu_inst_pe_1_1_6_int_q_reg_v_2__1_,
         npu_inst_pe_1_1_6_int_q_reg_v_1__0_,
         npu_inst_pe_1_1_6_int_q_reg_v_1__1_,
         npu_inst_pe_1_1_6_int_q_reg_v_0__0_,
         npu_inst_pe_1_1_6_int_q_reg_v_0__1_,
         npu_inst_pe_1_1_6_int_q_reg_h_5__0_,
         npu_inst_pe_1_1_6_int_q_reg_h_5__1_,
         npu_inst_pe_1_1_6_int_q_reg_h_4__0_,
         npu_inst_pe_1_1_6_int_q_reg_h_4__1_,
         npu_inst_pe_1_1_6_int_q_reg_h_3__0_,
         npu_inst_pe_1_1_6_int_q_reg_h_3__1_,
         npu_inst_pe_1_1_6_int_q_reg_h_2__0_,
         npu_inst_pe_1_1_6_int_q_reg_h_2__1_,
         npu_inst_pe_1_1_6_int_q_reg_h_1__0_,
         npu_inst_pe_1_1_6_int_q_reg_h_1__1_,
         npu_inst_pe_1_1_6_int_q_reg_h_0__0_,
         npu_inst_pe_1_1_6_int_q_reg_h_0__1_, npu_inst_pe_1_1_7_n119,
         npu_inst_pe_1_1_7_n118, npu_inst_pe_1_1_7_n117,
         npu_inst_pe_1_1_7_n116, npu_inst_pe_1_1_7_n115,
         npu_inst_pe_1_1_7_n114, npu_inst_pe_1_1_7_n113,
         npu_inst_pe_1_1_7_n112, npu_inst_pe_1_1_7_n111,
         npu_inst_pe_1_1_7_n110, npu_inst_pe_1_1_7_n109,
         npu_inst_pe_1_1_7_n108, npu_inst_pe_1_1_7_n107,
         npu_inst_pe_1_1_7_n106, npu_inst_pe_1_1_7_n105,
         npu_inst_pe_1_1_7_n104, npu_inst_pe_1_1_7_n103,
         npu_inst_pe_1_1_7_n102, npu_inst_pe_1_1_7_n101,
         npu_inst_pe_1_1_7_n100, npu_inst_pe_1_1_7_n99, npu_inst_pe_1_1_7_n98,
         npu_inst_pe_1_1_7_n36, npu_inst_pe_1_1_7_n35, npu_inst_pe_1_1_7_n34,
         npu_inst_pe_1_1_7_n33, npu_inst_pe_1_1_7_n32, npu_inst_pe_1_1_7_n31,
         npu_inst_pe_1_1_7_n30, npu_inst_pe_1_1_7_n29, npu_inst_pe_1_1_7_n28,
         npu_inst_pe_1_1_7_n25, npu_inst_pe_1_1_7_n24, npu_inst_pe_1_1_7_n23,
         npu_inst_pe_1_1_7_n22, npu_inst_pe_1_1_7_n21, npu_inst_pe_1_1_7_n20,
         npu_inst_pe_1_1_7_n19, npu_inst_pe_1_1_7_n18, npu_inst_pe_1_1_7_n17,
         npu_inst_pe_1_1_7_n16, npu_inst_pe_1_1_7_n15, npu_inst_pe_1_1_7_n14,
         npu_inst_pe_1_1_7_n13, npu_inst_pe_1_1_7_n12, npu_inst_pe_1_1_7_n11,
         npu_inst_pe_1_1_7_n10, npu_inst_pe_1_1_7_n9, npu_inst_pe_1_1_7_n8,
         npu_inst_pe_1_1_7_n7, npu_inst_pe_1_1_7_n6, npu_inst_pe_1_1_7_n5,
         npu_inst_pe_1_1_7_n4, npu_inst_pe_1_1_7_n3, npu_inst_pe_1_1_7_n2,
         npu_inst_pe_1_1_7_n1, npu_inst_pe_1_1_7_sub_67_carry_7_,
         npu_inst_pe_1_1_7_sub_67_carry_6_, npu_inst_pe_1_1_7_sub_67_carry_5_,
         npu_inst_pe_1_1_7_sub_67_carry_4_, npu_inst_pe_1_1_7_sub_67_carry_3_,
         npu_inst_pe_1_1_7_sub_67_carry_2_, npu_inst_pe_1_1_7_sub_67_carry_1_,
         npu_inst_pe_1_1_7_add_69_carry_7_, npu_inst_pe_1_1_7_add_69_carry_6_,
         npu_inst_pe_1_1_7_add_69_carry_5_, npu_inst_pe_1_1_7_add_69_carry_4_,
         npu_inst_pe_1_1_7_add_69_carry_3_, npu_inst_pe_1_1_7_add_69_carry_2_,
         npu_inst_pe_1_1_7_add_69_carry_1_, npu_inst_pe_1_1_7_n97,
         npu_inst_pe_1_1_7_n96, npu_inst_pe_1_1_7_n95, npu_inst_pe_1_1_7_n94,
         npu_inst_pe_1_1_7_n93, npu_inst_pe_1_1_7_n92, npu_inst_pe_1_1_7_n91,
         npu_inst_pe_1_1_7_n90, npu_inst_pe_1_1_7_n89, npu_inst_pe_1_1_7_n88,
         npu_inst_pe_1_1_7_n87, npu_inst_pe_1_1_7_n86, npu_inst_pe_1_1_7_n85,
         npu_inst_pe_1_1_7_n84, npu_inst_pe_1_1_7_n83, npu_inst_pe_1_1_7_n82,
         npu_inst_pe_1_1_7_n81, npu_inst_pe_1_1_7_n80, npu_inst_pe_1_1_7_n79,
         npu_inst_pe_1_1_7_n78, npu_inst_pe_1_1_7_n77, npu_inst_pe_1_1_7_n76,
         npu_inst_pe_1_1_7_n75, npu_inst_pe_1_1_7_n74, npu_inst_pe_1_1_7_n73,
         npu_inst_pe_1_1_7_n72, npu_inst_pe_1_1_7_n71, npu_inst_pe_1_1_7_n70,
         npu_inst_pe_1_1_7_n69, npu_inst_pe_1_1_7_n68, npu_inst_pe_1_1_7_n67,
         npu_inst_pe_1_1_7_n66, npu_inst_pe_1_1_7_n65, npu_inst_pe_1_1_7_n64,
         npu_inst_pe_1_1_7_n63, npu_inst_pe_1_1_7_n62, npu_inst_pe_1_1_7_n61,
         npu_inst_pe_1_1_7_n60, npu_inst_pe_1_1_7_n59, npu_inst_pe_1_1_7_n58,
         npu_inst_pe_1_1_7_n57, npu_inst_pe_1_1_7_n56, npu_inst_pe_1_1_7_n55,
         npu_inst_pe_1_1_7_n54, npu_inst_pe_1_1_7_n53, npu_inst_pe_1_1_7_n52,
         npu_inst_pe_1_1_7_n51, npu_inst_pe_1_1_7_n50, npu_inst_pe_1_1_7_n49,
         npu_inst_pe_1_1_7_n48, npu_inst_pe_1_1_7_n47, npu_inst_pe_1_1_7_n46,
         npu_inst_pe_1_1_7_n45, npu_inst_pe_1_1_7_n44, npu_inst_pe_1_1_7_n43,
         npu_inst_pe_1_1_7_n42, npu_inst_pe_1_1_7_n41, npu_inst_pe_1_1_7_n40,
         npu_inst_pe_1_1_7_n39, npu_inst_pe_1_1_7_n38, npu_inst_pe_1_1_7_n37,
         npu_inst_pe_1_1_7_n27, npu_inst_pe_1_1_7_n26,
         npu_inst_pe_1_1_7_net4223, npu_inst_pe_1_1_7_net4217,
         npu_inst_pe_1_1_7_N94, npu_inst_pe_1_1_7_N93, npu_inst_pe_1_1_7_N84,
         npu_inst_pe_1_1_7_N80, npu_inst_pe_1_1_7_N79, npu_inst_pe_1_1_7_N78,
         npu_inst_pe_1_1_7_N77, npu_inst_pe_1_1_7_N76, npu_inst_pe_1_1_7_N75,
         npu_inst_pe_1_1_7_N74, npu_inst_pe_1_1_7_N73, npu_inst_pe_1_1_7_N72,
         npu_inst_pe_1_1_7_N71, npu_inst_pe_1_1_7_N70, npu_inst_pe_1_1_7_N69,
         npu_inst_pe_1_1_7_N68, npu_inst_pe_1_1_7_N67, npu_inst_pe_1_1_7_N66,
         npu_inst_pe_1_1_7_N65, npu_inst_pe_1_1_7_int_q_acc_0_,
         npu_inst_pe_1_1_7_int_q_acc_1_, npu_inst_pe_1_1_7_int_q_acc_2_,
         npu_inst_pe_1_1_7_int_q_acc_3_, npu_inst_pe_1_1_7_int_q_acc_4_,
         npu_inst_pe_1_1_7_int_q_acc_5_, npu_inst_pe_1_1_7_int_q_acc_6_,
         npu_inst_pe_1_1_7_int_q_acc_7_, npu_inst_pe_1_1_7_int_data_0_,
         npu_inst_pe_1_1_7_int_data_1_, npu_inst_pe_1_1_7_int_q_weight_0_,
         npu_inst_pe_1_1_7_int_q_weight_1_,
         npu_inst_pe_1_1_7_int_q_reg_v_5__0_,
         npu_inst_pe_1_1_7_int_q_reg_v_5__1_,
         npu_inst_pe_1_1_7_int_q_reg_v_4__0_,
         npu_inst_pe_1_1_7_int_q_reg_v_4__1_,
         npu_inst_pe_1_1_7_int_q_reg_v_3__0_,
         npu_inst_pe_1_1_7_int_q_reg_v_3__1_,
         npu_inst_pe_1_1_7_int_q_reg_v_2__0_,
         npu_inst_pe_1_1_7_int_q_reg_v_2__1_,
         npu_inst_pe_1_1_7_int_q_reg_v_1__0_,
         npu_inst_pe_1_1_7_int_q_reg_v_1__1_,
         npu_inst_pe_1_1_7_int_q_reg_v_0__0_,
         npu_inst_pe_1_1_7_int_q_reg_v_0__1_,
         npu_inst_pe_1_1_7_int_q_reg_h_5__0_,
         npu_inst_pe_1_1_7_int_q_reg_h_5__1_,
         npu_inst_pe_1_1_7_int_q_reg_h_4__0_,
         npu_inst_pe_1_1_7_int_q_reg_h_4__1_,
         npu_inst_pe_1_1_7_int_q_reg_h_3__0_,
         npu_inst_pe_1_1_7_int_q_reg_h_3__1_,
         npu_inst_pe_1_1_7_int_q_reg_h_2__0_,
         npu_inst_pe_1_1_7_int_q_reg_h_2__1_,
         npu_inst_pe_1_1_7_int_q_reg_h_1__0_,
         npu_inst_pe_1_1_7_int_q_reg_h_1__1_,
         npu_inst_pe_1_1_7_int_q_reg_h_0__0_,
         npu_inst_pe_1_1_7_int_q_reg_h_0__1_, npu_inst_pe_1_2_0_n118,
         npu_inst_pe_1_2_0_n117, npu_inst_pe_1_2_0_n116,
         npu_inst_pe_1_2_0_n115, npu_inst_pe_1_2_0_n114,
         npu_inst_pe_1_2_0_n113, npu_inst_pe_1_2_0_n112,
         npu_inst_pe_1_2_0_n111, npu_inst_pe_1_2_0_n110,
         npu_inst_pe_1_2_0_n109, npu_inst_pe_1_2_0_n108,
         npu_inst_pe_1_2_0_n107, npu_inst_pe_1_2_0_n106,
         npu_inst_pe_1_2_0_n105, npu_inst_pe_1_2_0_n104,
         npu_inst_pe_1_2_0_n103, npu_inst_pe_1_2_0_n102,
         npu_inst_pe_1_2_0_n101, npu_inst_pe_1_2_0_n100, npu_inst_pe_1_2_0_n99,
         npu_inst_pe_1_2_0_n98, npu_inst_pe_1_2_0_n36, npu_inst_pe_1_2_0_n35,
         npu_inst_pe_1_2_0_n34, npu_inst_pe_1_2_0_n33, npu_inst_pe_1_2_0_n32,
         npu_inst_pe_1_2_0_n31, npu_inst_pe_1_2_0_n30, npu_inst_pe_1_2_0_n29,
         npu_inst_pe_1_2_0_n28, npu_inst_pe_1_2_0_n25, npu_inst_pe_1_2_0_n24,
         npu_inst_pe_1_2_0_n23, npu_inst_pe_1_2_0_n22, npu_inst_pe_1_2_0_n21,
         npu_inst_pe_1_2_0_n20, npu_inst_pe_1_2_0_n19, npu_inst_pe_1_2_0_n18,
         npu_inst_pe_1_2_0_n17, npu_inst_pe_1_2_0_n16, npu_inst_pe_1_2_0_n15,
         npu_inst_pe_1_2_0_n14, npu_inst_pe_1_2_0_n13, npu_inst_pe_1_2_0_n12,
         npu_inst_pe_1_2_0_n11, npu_inst_pe_1_2_0_n10, npu_inst_pe_1_2_0_n9,
         npu_inst_pe_1_2_0_n8, npu_inst_pe_1_2_0_n7, npu_inst_pe_1_2_0_n6,
         npu_inst_pe_1_2_0_n5, npu_inst_pe_1_2_0_n4, npu_inst_pe_1_2_0_n3,
         npu_inst_pe_1_2_0_n2, npu_inst_pe_1_2_0_n1,
         npu_inst_pe_1_2_0_sub_67_carry_7_, npu_inst_pe_1_2_0_sub_67_carry_6_,
         npu_inst_pe_1_2_0_sub_67_carry_5_, npu_inst_pe_1_2_0_sub_67_carry_4_,
         npu_inst_pe_1_2_0_sub_67_carry_3_, npu_inst_pe_1_2_0_sub_67_carry_2_,
         npu_inst_pe_1_2_0_sub_67_carry_1_, npu_inst_pe_1_2_0_add_69_carry_7_,
         npu_inst_pe_1_2_0_add_69_carry_6_, npu_inst_pe_1_2_0_add_69_carry_5_,
         npu_inst_pe_1_2_0_add_69_carry_4_, npu_inst_pe_1_2_0_add_69_carry_3_,
         npu_inst_pe_1_2_0_add_69_carry_2_, npu_inst_pe_1_2_0_add_69_carry_1_,
         npu_inst_pe_1_2_0_n97, npu_inst_pe_1_2_0_n96, npu_inst_pe_1_2_0_n95,
         npu_inst_pe_1_2_0_n94, npu_inst_pe_1_2_0_n93, npu_inst_pe_1_2_0_n92,
         npu_inst_pe_1_2_0_n91, npu_inst_pe_1_2_0_n90, npu_inst_pe_1_2_0_n89,
         npu_inst_pe_1_2_0_n88, npu_inst_pe_1_2_0_n87, npu_inst_pe_1_2_0_n86,
         npu_inst_pe_1_2_0_n85, npu_inst_pe_1_2_0_n84, npu_inst_pe_1_2_0_n83,
         npu_inst_pe_1_2_0_n82, npu_inst_pe_1_2_0_n81, npu_inst_pe_1_2_0_n80,
         npu_inst_pe_1_2_0_n79, npu_inst_pe_1_2_0_n78, npu_inst_pe_1_2_0_n77,
         npu_inst_pe_1_2_0_n76, npu_inst_pe_1_2_0_n75, npu_inst_pe_1_2_0_n74,
         npu_inst_pe_1_2_0_n73, npu_inst_pe_1_2_0_n72, npu_inst_pe_1_2_0_n71,
         npu_inst_pe_1_2_0_n70, npu_inst_pe_1_2_0_n69, npu_inst_pe_1_2_0_n68,
         npu_inst_pe_1_2_0_n67, npu_inst_pe_1_2_0_n66, npu_inst_pe_1_2_0_n65,
         npu_inst_pe_1_2_0_n64, npu_inst_pe_1_2_0_n63, npu_inst_pe_1_2_0_n62,
         npu_inst_pe_1_2_0_n61, npu_inst_pe_1_2_0_n60, npu_inst_pe_1_2_0_n59,
         npu_inst_pe_1_2_0_n58, npu_inst_pe_1_2_0_n57, npu_inst_pe_1_2_0_n56,
         npu_inst_pe_1_2_0_n55, npu_inst_pe_1_2_0_n54, npu_inst_pe_1_2_0_n53,
         npu_inst_pe_1_2_0_n52, npu_inst_pe_1_2_0_n51, npu_inst_pe_1_2_0_n50,
         npu_inst_pe_1_2_0_n49, npu_inst_pe_1_2_0_n48, npu_inst_pe_1_2_0_n47,
         npu_inst_pe_1_2_0_n46, npu_inst_pe_1_2_0_n45, npu_inst_pe_1_2_0_n44,
         npu_inst_pe_1_2_0_n43, npu_inst_pe_1_2_0_n42, npu_inst_pe_1_2_0_n41,
         npu_inst_pe_1_2_0_n40, npu_inst_pe_1_2_0_n39, npu_inst_pe_1_2_0_n38,
         npu_inst_pe_1_2_0_n37, npu_inst_pe_1_2_0_n27, npu_inst_pe_1_2_0_n26,
         npu_inst_pe_1_2_0_net4200, npu_inst_pe_1_2_0_net4194,
         npu_inst_pe_1_2_0_N94, npu_inst_pe_1_2_0_N93, npu_inst_pe_1_2_0_N84,
         npu_inst_pe_1_2_0_N80, npu_inst_pe_1_2_0_N79, npu_inst_pe_1_2_0_N78,
         npu_inst_pe_1_2_0_N77, npu_inst_pe_1_2_0_N76, npu_inst_pe_1_2_0_N75,
         npu_inst_pe_1_2_0_N74, npu_inst_pe_1_2_0_N73, npu_inst_pe_1_2_0_N72,
         npu_inst_pe_1_2_0_N71, npu_inst_pe_1_2_0_N70, npu_inst_pe_1_2_0_N69,
         npu_inst_pe_1_2_0_N68, npu_inst_pe_1_2_0_N67, npu_inst_pe_1_2_0_N66,
         npu_inst_pe_1_2_0_N65, npu_inst_pe_1_2_0_int_q_acc_0_,
         npu_inst_pe_1_2_0_int_q_acc_1_, npu_inst_pe_1_2_0_int_q_acc_2_,
         npu_inst_pe_1_2_0_int_q_acc_3_, npu_inst_pe_1_2_0_int_q_acc_4_,
         npu_inst_pe_1_2_0_int_q_acc_5_, npu_inst_pe_1_2_0_int_q_acc_6_,
         npu_inst_pe_1_2_0_int_q_acc_7_, npu_inst_pe_1_2_0_int_data_0_,
         npu_inst_pe_1_2_0_int_data_1_, npu_inst_pe_1_2_0_int_q_weight_0_,
         npu_inst_pe_1_2_0_int_q_weight_1_,
         npu_inst_pe_1_2_0_int_q_reg_v_5__0_,
         npu_inst_pe_1_2_0_int_q_reg_v_5__1_,
         npu_inst_pe_1_2_0_int_q_reg_v_4__0_,
         npu_inst_pe_1_2_0_int_q_reg_v_4__1_,
         npu_inst_pe_1_2_0_int_q_reg_v_3__0_,
         npu_inst_pe_1_2_0_int_q_reg_v_3__1_,
         npu_inst_pe_1_2_0_int_q_reg_v_2__0_,
         npu_inst_pe_1_2_0_int_q_reg_v_2__1_,
         npu_inst_pe_1_2_0_int_q_reg_v_1__0_,
         npu_inst_pe_1_2_0_int_q_reg_v_1__1_,
         npu_inst_pe_1_2_0_int_q_reg_v_0__0_,
         npu_inst_pe_1_2_0_int_q_reg_v_0__1_,
         npu_inst_pe_1_2_0_int_q_reg_h_5__0_,
         npu_inst_pe_1_2_0_int_q_reg_h_5__1_,
         npu_inst_pe_1_2_0_int_q_reg_h_4__0_,
         npu_inst_pe_1_2_0_int_q_reg_h_4__1_,
         npu_inst_pe_1_2_0_int_q_reg_h_3__0_,
         npu_inst_pe_1_2_0_int_q_reg_h_3__1_,
         npu_inst_pe_1_2_0_int_q_reg_h_2__0_,
         npu_inst_pe_1_2_0_int_q_reg_h_2__1_,
         npu_inst_pe_1_2_0_int_q_reg_h_1__0_,
         npu_inst_pe_1_2_0_int_q_reg_h_1__1_,
         npu_inst_pe_1_2_0_int_q_reg_h_0__0_,
         npu_inst_pe_1_2_0_int_q_reg_h_0__1_, npu_inst_pe_1_2_0_o_data_h_0_,
         npu_inst_pe_1_2_0_o_data_h_1_, npu_inst_pe_1_2_1_n119,
         npu_inst_pe_1_2_1_n118, npu_inst_pe_1_2_1_n117,
         npu_inst_pe_1_2_1_n116, npu_inst_pe_1_2_1_n115,
         npu_inst_pe_1_2_1_n114, npu_inst_pe_1_2_1_n113,
         npu_inst_pe_1_2_1_n112, npu_inst_pe_1_2_1_n111,
         npu_inst_pe_1_2_1_n110, npu_inst_pe_1_2_1_n109,
         npu_inst_pe_1_2_1_n108, npu_inst_pe_1_2_1_n107,
         npu_inst_pe_1_2_1_n106, npu_inst_pe_1_2_1_n105,
         npu_inst_pe_1_2_1_n104, npu_inst_pe_1_2_1_n103,
         npu_inst_pe_1_2_1_n102, npu_inst_pe_1_2_1_n101,
         npu_inst_pe_1_2_1_n100, npu_inst_pe_1_2_1_n99, npu_inst_pe_1_2_1_n98,
         npu_inst_pe_1_2_1_n36, npu_inst_pe_1_2_1_n35, npu_inst_pe_1_2_1_n34,
         npu_inst_pe_1_2_1_n33, npu_inst_pe_1_2_1_n32, npu_inst_pe_1_2_1_n31,
         npu_inst_pe_1_2_1_n30, npu_inst_pe_1_2_1_n29, npu_inst_pe_1_2_1_n28,
         npu_inst_pe_1_2_1_n25, npu_inst_pe_1_2_1_n24, npu_inst_pe_1_2_1_n23,
         npu_inst_pe_1_2_1_n22, npu_inst_pe_1_2_1_n21, npu_inst_pe_1_2_1_n20,
         npu_inst_pe_1_2_1_n19, npu_inst_pe_1_2_1_n18, npu_inst_pe_1_2_1_n17,
         npu_inst_pe_1_2_1_n16, npu_inst_pe_1_2_1_n15, npu_inst_pe_1_2_1_n14,
         npu_inst_pe_1_2_1_n13, npu_inst_pe_1_2_1_n12, npu_inst_pe_1_2_1_n11,
         npu_inst_pe_1_2_1_n10, npu_inst_pe_1_2_1_n9, npu_inst_pe_1_2_1_n8,
         npu_inst_pe_1_2_1_n7, npu_inst_pe_1_2_1_n6, npu_inst_pe_1_2_1_n5,
         npu_inst_pe_1_2_1_n4, npu_inst_pe_1_2_1_n3, npu_inst_pe_1_2_1_n2,
         npu_inst_pe_1_2_1_n1, npu_inst_pe_1_2_1_sub_67_carry_7_,
         npu_inst_pe_1_2_1_sub_67_carry_6_, npu_inst_pe_1_2_1_sub_67_carry_5_,
         npu_inst_pe_1_2_1_sub_67_carry_4_, npu_inst_pe_1_2_1_sub_67_carry_3_,
         npu_inst_pe_1_2_1_sub_67_carry_2_, npu_inst_pe_1_2_1_sub_67_carry_1_,
         npu_inst_pe_1_2_1_add_69_carry_7_, npu_inst_pe_1_2_1_add_69_carry_6_,
         npu_inst_pe_1_2_1_add_69_carry_5_, npu_inst_pe_1_2_1_add_69_carry_4_,
         npu_inst_pe_1_2_1_add_69_carry_3_, npu_inst_pe_1_2_1_add_69_carry_2_,
         npu_inst_pe_1_2_1_add_69_carry_1_, npu_inst_pe_1_2_1_n97,
         npu_inst_pe_1_2_1_n96, npu_inst_pe_1_2_1_n95, npu_inst_pe_1_2_1_n94,
         npu_inst_pe_1_2_1_n93, npu_inst_pe_1_2_1_n92, npu_inst_pe_1_2_1_n91,
         npu_inst_pe_1_2_1_n90, npu_inst_pe_1_2_1_n89, npu_inst_pe_1_2_1_n88,
         npu_inst_pe_1_2_1_n87, npu_inst_pe_1_2_1_n86, npu_inst_pe_1_2_1_n85,
         npu_inst_pe_1_2_1_n84, npu_inst_pe_1_2_1_n83, npu_inst_pe_1_2_1_n82,
         npu_inst_pe_1_2_1_n81, npu_inst_pe_1_2_1_n80, npu_inst_pe_1_2_1_n79,
         npu_inst_pe_1_2_1_n78, npu_inst_pe_1_2_1_n77, npu_inst_pe_1_2_1_n76,
         npu_inst_pe_1_2_1_n75, npu_inst_pe_1_2_1_n74, npu_inst_pe_1_2_1_n73,
         npu_inst_pe_1_2_1_n72, npu_inst_pe_1_2_1_n71, npu_inst_pe_1_2_1_n70,
         npu_inst_pe_1_2_1_n69, npu_inst_pe_1_2_1_n68, npu_inst_pe_1_2_1_n67,
         npu_inst_pe_1_2_1_n66, npu_inst_pe_1_2_1_n65, npu_inst_pe_1_2_1_n64,
         npu_inst_pe_1_2_1_n63, npu_inst_pe_1_2_1_n62, npu_inst_pe_1_2_1_n61,
         npu_inst_pe_1_2_1_n60, npu_inst_pe_1_2_1_n59, npu_inst_pe_1_2_1_n58,
         npu_inst_pe_1_2_1_n57, npu_inst_pe_1_2_1_n56, npu_inst_pe_1_2_1_n55,
         npu_inst_pe_1_2_1_n54, npu_inst_pe_1_2_1_n53, npu_inst_pe_1_2_1_n52,
         npu_inst_pe_1_2_1_n51, npu_inst_pe_1_2_1_n50, npu_inst_pe_1_2_1_n49,
         npu_inst_pe_1_2_1_n48, npu_inst_pe_1_2_1_n47, npu_inst_pe_1_2_1_n46,
         npu_inst_pe_1_2_1_n45, npu_inst_pe_1_2_1_n44, npu_inst_pe_1_2_1_n43,
         npu_inst_pe_1_2_1_n42, npu_inst_pe_1_2_1_n41, npu_inst_pe_1_2_1_n40,
         npu_inst_pe_1_2_1_n39, npu_inst_pe_1_2_1_n38, npu_inst_pe_1_2_1_n37,
         npu_inst_pe_1_2_1_n27, npu_inst_pe_1_2_1_n26,
         npu_inst_pe_1_2_1_net4177, npu_inst_pe_1_2_1_net4171,
         npu_inst_pe_1_2_1_N94, npu_inst_pe_1_2_1_N93, npu_inst_pe_1_2_1_N84,
         npu_inst_pe_1_2_1_N80, npu_inst_pe_1_2_1_N79, npu_inst_pe_1_2_1_N78,
         npu_inst_pe_1_2_1_N77, npu_inst_pe_1_2_1_N76, npu_inst_pe_1_2_1_N75,
         npu_inst_pe_1_2_1_N74, npu_inst_pe_1_2_1_N73, npu_inst_pe_1_2_1_N72,
         npu_inst_pe_1_2_1_N71, npu_inst_pe_1_2_1_N70, npu_inst_pe_1_2_1_N69,
         npu_inst_pe_1_2_1_N68, npu_inst_pe_1_2_1_N67, npu_inst_pe_1_2_1_N66,
         npu_inst_pe_1_2_1_N65, npu_inst_pe_1_2_1_int_q_acc_0_,
         npu_inst_pe_1_2_1_int_q_acc_1_, npu_inst_pe_1_2_1_int_q_acc_2_,
         npu_inst_pe_1_2_1_int_q_acc_3_, npu_inst_pe_1_2_1_int_q_acc_4_,
         npu_inst_pe_1_2_1_int_q_acc_5_, npu_inst_pe_1_2_1_int_q_acc_6_,
         npu_inst_pe_1_2_1_int_q_acc_7_, npu_inst_pe_1_2_1_int_data_0_,
         npu_inst_pe_1_2_1_int_data_1_, npu_inst_pe_1_2_1_int_q_weight_0_,
         npu_inst_pe_1_2_1_int_q_weight_1_,
         npu_inst_pe_1_2_1_int_q_reg_v_5__0_,
         npu_inst_pe_1_2_1_int_q_reg_v_5__1_,
         npu_inst_pe_1_2_1_int_q_reg_v_4__0_,
         npu_inst_pe_1_2_1_int_q_reg_v_4__1_,
         npu_inst_pe_1_2_1_int_q_reg_v_3__0_,
         npu_inst_pe_1_2_1_int_q_reg_v_3__1_,
         npu_inst_pe_1_2_1_int_q_reg_v_2__0_,
         npu_inst_pe_1_2_1_int_q_reg_v_2__1_,
         npu_inst_pe_1_2_1_int_q_reg_v_1__0_,
         npu_inst_pe_1_2_1_int_q_reg_v_1__1_,
         npu_inst_pe_1_2_1_int_q_reg_v_0__0_,
         npu_inst_pe_1_2_1_int_q_reg_v_0__1_,
         npu_inst_pe_1_2_1_int_q_reg_h_5__0_,
         npu_inst_pe_1_2_1_int_q_reg_h_5__1_,
         npu_inst_pe_1_2_1_int_q_reg_h_4__0_,
         npu_inst_pe_1_2_1_int_q_reg_h_4__1_,
         npu_inst_pe_1_2_1_int_q_reg_h_3__0_,
         npu_inst_pe_1_2_1_int_q_reg_h_3__1_,
         npu_inst_pe_1_2_1_int_q_reg_h_2__0_,
         npu_inst_pe_1_2_1_int_q_reg_h_2__1_,
         npu_inst_pe_1_2_1_int_q_reg_h_1__0_,
         npu_inst_pe_1_2_1_int_q_reg_h_1__1_,
         npu_inst_pe_1_2_1_int_q_reg_h_0__0_,
         npu_inst_pe_1_2_1_int_q_reg_h_0__1_, npu_inst_pe_1_2_2_n119,
         npu_inst_pe_1_2_2_n118, npu_inst_pe_1_2_2_n117,
         npu_inst_pe_1_2_2_n116, npu_inst_pe_1_2_2_n115,
         npu_inst_pe_1_2_2_n114, npu_inst_pe_1_2_2_n113,
         npu_inst_pe_1_2_2_n112, npu_inst_pe_1_2_2_n111,
         npu_inst_pe_1_2_2_n110, npu_inst_pe_1_2_2_n109,
         npu_inst_pe_1_2_2_n108, npu_inst_pe_1_2_2_n107,
         npu_inst_pe_1_2_2_n106, npu_inst_pe_1_2_2_n105,
         npu_inst_pe_1_2_2_n104, npu_inst_pe_1_2_2_n103,
         npu_inst_pe_1_2_2_n102, npu_inst_pe_1_2_2_n101,
         npu_inst_pe_1_2_2_n100, npu_inst_pe_1_2_2_n99, npu_inst_pe_1_2_2_n98,
         npu_inst_pe_1_2_2_n36, npu_inst_pe_1_2_2_n35, npu_inst_pe_1_2_2_n34,
         npu_inst_pe_1_2_2_n33, npu_inst_pe_1_2_2_n32, npu_inst_pe_1_2_2_n31,
         npu_inst_pe_1_2_2_n30, npu_inst_pe_1_2_2_n29, npu_inst_pe_1_2_2_n28,
         npu_inst_pe_1_2_2_n25, npu_inst_pe_1_2_2_n24, npu_inst_pe_1_2_2_n23,
         npu_inst_pe_1_2_2_n22, npu_inst_pe_1_2_2_n21, npu_inst_pe_1_2_2_n20,
         npu_inst_pe_1_2_2_n19, npu_inst_pe_1_2_2_n18, npu_inst_pe_1_2_2_n17,
         npu_inst_pe_1_2_2_n16, npu_inst_pe_1_2_2_n15, npu_inst_pe_1_2_2_n14,
         npu_inst_pe_1_2_2_n13, npu_inst_pe_1_2_2_n12, npu_inst_pe_1_2_2_n11,
         npu_inst_pe_1_2_2_n10, npu_inst_pe_1_2_2_n9, npu_inst_pe_1_2_2_n8,
         npu_inst_pe_1_2_2_n7, npu_inst_pe_1_2_2_n6, npu_inst_pe_1_2_2_n5,
         npu_inst_pe_1_2_2_n4, npu_inst_pe_1_2_2_n3, npu_inst_pe_1_2_2_n2,
         npu_inst_pe_1_2_2_n1, npu_inst_pe_1_2_2_sub_67_carry_7_,
         npu_inst_pe_1_2_2_sub_67_carry_6_, npu_inst_pe_1_2_2_sub_67_carry_5_,
         npu_inst_pe_1_2_2_sub_67_carry_4_, npu_inst_pe_1_2_2_sub_67_carry_3_,
         npu_inst_pe_1_2_2_sub_67_carry_2_, npu_inst_pe_1_2_2_sub_67_carry_1_,
         npu_inst_pe_1_2_2_add_69_carry_7_, npu_inst_pe_1_2_2_add_69_carry_6_,
         npu_inst_pe_1_2_2_add_69_carry_5_, npu_inst_pe_1_2_2_add_69_carry_4_,
         npu_inst_pe_1_2_2_add_69_carry_3_, npu_inst_pe_1_2_2_add_69_carry_2_,
         npu_inst_pe_1_2_2_add_69_carry_1_, npu_inst_pe_1_2_2_n97,
         npu_inst_pe_1_2_2_n96, npu_inst_pe_1_2_2_n95, npu_inst_pe_1_2_2_n94,
         npu_inst_pe_1_2_2_n93, npu_inst_pe_1_2_2_n92, npu_inst_pe_1_2_2_n91,
         npu_inst_pe_1_2_2_n90, npu_inst_pe_1_2_2_n89, npu_inst_pe_1_2_2_n88,
         npu_inst_pe_1_2_2_n87, npu_inst_pe_1_2_2_n86, npu_inst_pe_1_2_2_n85,
         npu_inst_pe_1_2_2_n84, npu_inst_pe_1_2_2_n83, npu_inst_pe_1_2_2_n82,
         npu_inst_pe_1_2_2_n81, npu_inst_pe_1_2_2_n80, npu_inst_pe_1_2_2_n79,
         npu_inst_pe_1_2_2_n78, npu_inst_pe_1_2_2_n77, npu_inst_pe_1_2_2_n76,
         npu_inst_pe_1_2_2_n75, npu_inst_pe_1_2_2_n74, npu_inst_pe_1_2_2_n73,
         npu_inst_pe_1_2_2_n72, npu_inst_pe_1_2_2_n71, npu_inst_pe_1_2_2_n70,
         npu_inst_pe_1_2_2_n69, npu_inst_pe_1_2_2_n68, npu_inst_pe_1_2_2_n67,
         npu_inst_pe_1_2_2_n66, npu_inst_pe_1_2_2_n65, npu_inst_pe_1_2_2_n64,
         npu_inst_pe_1_2_2_n63, npu_inst_pe_1_2_2_n62, npu_inst_pe_1_2_2_n61,
         npu_inst_pe_1_2_2_n60, npu_inst_pe_1_2_2_n59, npu_inst_pe_1_2_2_n58,
         npu_inst_pe_1_2_2_n57, npu_inst_pe_1_2_2_n56, npu_inst_pe_1_2_2_n55,
         npu_inst_pe_1_2_2_n54, npu_inst_pe_1_2_2_n53, npu_inst_pe_1_2_2_n52,
         npu_inst_pe_1_2_2_n51, npu_inst_pe_1_2_2_n50, npu_inst_pe_1_2_2_n49,
         npu_inst_pe_1_2_2_n48, npu_inst_pe_1_2_2_n47, npu_inst_pe_1_2_2_n46,
         npu_inst_pe_1_2_2_n45, npu_inst_pe_1_2_2_n44, npu_inst_pe_1_2_2_n43,
         npu_inst_pe_1_2_2_n42, npu_inst_pe_1_2_2_n41, npu_inst_pe_1_2_2_n40,
         npu_inst_pe_1_2_2_n39, npu_inst_pe_1_2_2_n38, npu_inst_pe_1_2_2_n37,
         npu_inst_pe_1_2_2_n27, npu_inst_pe_1_2_2_n26,
         npu_inst_pe_1_2_2_net4154, npu_inst_pe_1_2_2_net4148,
         npu_inst_pe_1_2_2_N94, npu_inst_pe_1_2_2_N93, npu_inst_pe_1_2_2_N84,
         npu_inst_pe_1_2_2_N80, npu_inst_pe_1_2_2_N79, npu_inst_pe_1_2_2_N78,
         npu_inst_pe_1_2_2_N77, npu_inst_pe_1_2_2_N76, npu_inst_pe_1_2_2_N75,
         npu_inst_pe_1_2_2_N74, npu_inst_pe_1_2_2_N73, npu_inst_pe_1_2_2_N72,
         npu_inst_pe_1_2_2_N71, npu_inst_pe_1_2_2_N70, npu_inst_pe_1_2_2_N69,
         npu_inst_pe_1_2_2_N68, npu_inst_pe_1_2_2_N67, npu_inst_pe_1_2_2_N66,
         npu_inst_pe_1_2_2_N65, npu_inst_pe_1_2_2_int_q_acc_0_,
         npu_inst_pe_1_2_2_int_q_acc_1_, npu_inst_pe_1_2_2_int_q_acc_2_,
         npu_inst_pe_1_2_2_int_q_acc_3_, npu_inst_pe_1_2_2_int_q_acc_4_,
         npu_inst_pe_1_2_2_int_q_acc_5_, npu_inst_pe_1_2_2_int_q_acc_6_,
         npu_inst_pe_1_2_2_int_q_acc_7_, npu_inst_pe_1_2_2_int_data_0_,
         npu_inst_pe_1_2_2_int_data_1_, npu_inst_pe_1_2_2_int_q_weight_0_,
         npu_inst_pe_1_2_2_int_q_weight_1_,
         npu_inst_pe_1_2_2_int_q_reg_v_5__0_,
         npu_inst_pe_1_2_2_int_q_reg_v_5__1_,
         npu_inst_pe_1_2_2_int_q_reg_v_4__0_,
         npu_inst_pe_1_2_2_int_q_reg_v_4__1_,
         npu_inst_pe_1_2_2_int_q_reg_v_3__0_,
         npu_inst_pe_1_2_2_int_q_reg_v_3__1_,
         npu_inst_pe_1_2_2_int_q_reg_v_2__0_,
         npu_inst_pe_1_2_2_int_q_reg_v_2__1_,
         npu_inst_pe_1_2_2_int_q_reg_v_1__0_,
         npu_inst_pe_1_2_2_int_q_reg_v_1__1_,
         npu_inst_pe_1_2_2_int_q_reg_v_0__0_,
         npu_inst_pe_1_2_2_int_q_reg_v_0__1_,
         npu_inst_pe_1_2_2_int_q_reg_h_5__0_,
         npu_inst_pe_1_2_2_int_q_reg_h_5__1_,
         npu_inst_pe_1_2_2_int_q_reg_h_4__0_,
         npu_inst_pe_1_2_2_int_q_reg_h_4__1_,
         npu_inst_pe_1_2_2_int_q_reg_h_3__0_,
         npu_inst_pe_1_2_2_int_q_reg_h_3__1_,
         npu_inst_pe_1_2_2_int_q_reg_h_2__0_,
         npu_inst_pe_1_2_2_int_q_reg_h_2__1_,
         npu_inst_pe_1_2_2_int_q_reg_h_1__0_,
         npu_inst_pe_1_2_2_int_q_reg_h_1__1_,
         npu_inst_pe_1_2_2_int_q_reg_h_0__0_,
         npu_inst_pe_1_2_2_int_q_reg_h_0__1_, npu_inst_pe_1_2_3_n119,
         npu_inst_pe_1_2_3_n118, npu_inst_pe_1_2_3_n117,
         npu_inst_pe_1_2_3_n116, npu_inst_pe_1_2_3_n115,
         npu_inst_pe_1_2_3_n114, npu_inst_pe_1_2_3_n113,
         npu_inst_pe_1_2_3_n112, npu_inst_pe_1_2_3_n111,
         npu_inst_pe_1_2_3_n110, npu_inst_pe_1_2_3_n109,
         npu_inst_pe_1_2_3_n108, npu_inst_pe_1_2_3_n107,
         npu_inst_pe_1_2_3_n106, npu_inst_pe_1_2_3_n105,
         npu_inst_pe_1_2_3_n104, npu_inst_pe_1_2_3_n103,
         npu_inst_pe_1_2_3_n102, npu_inst_pe_1_2_3_n101,
         npu_inst_pe_1_2_3_n100, npu_inst_pe_1_2_3_n99, npu_inst_pe_1_2_3_n98,
         npu_inst_pe_1_2_3_n36, npu_inst_pe_1_2_3_n35, npu_inst_pe_1_2_3_n34,
         npu_inst_pe_1_2_3_n33, npu_inst_pe_1_2_3_n32, npu_inst_pe_1_2_3_n31,
         npu_inst_pe_1_2_3_n30, npu_inst_pe_1_2_3_n29, npu_inst_pe_1_2_3_n28,
         npu_inst_pe_1_2_3_n25, npu_inst_pe_1_2_3_n24, npu_inst_pe_1_2_3_n23,
         npu_inst_pe_1_2_3_n22, npu_inst_pe_1_2_3_n21, npu_inst_pe_1_2_3_n20,
         npu_inst_pe_1_2_3_n19, npu_inst_pe_1_2_3_n18, npu_inst_pe_1_2_3_n17,
         npu_inst_pe_1_2_3_n16, npu_inst_pe_1_2_3_n15, npu_inst_pe_1_2_3_n14,
         npu_inst_pe_1_2_3_n13, npu_inst_pe_1_2_3_n12, npu_inst_pe_1_2_3_n11,
         npu_inst_pe_1_2_3_n10, npu_inst_pe_1_2_3_n9, npu_inst_pe_1_2_3_n8,
         npu_inst_pe_1_2_3_n7, npu_inst_pe_1_2_3_n6, npu_inst_pe_1_2_3_n5,
         npu_inst_pe_1_2_3_n4, npu_inst_pe_1_2_3_n3, npu_inst_pe_1_2_3_n2,
         npu_inst_pe_1_2_3_n1, npu_inst_pe_1_2_3_sub_67_carry_7_,
         npu_inst_pe_1_2_3_sub_67_carry_6_, npu_inst_pe_1_2_3_sub_67_carry_5_,
         npu_inst_pe_1_2_3_sub_67_carry_4_, npu_inst_pe_1_2_3_sub_67_carry_3_,
         npu_inst_pe_1_2_3_sub_67_carry_2_, npu_inst_pe_1_2_3_sub_67_carry_1_,
         npu_inst_pe_1_2_3_add_69_carry_7_, npu_inst_pe_1_2_3_add_69_carry_6_,
         npu_inst_pe_1_2_3_add_69_carry_5_, npu_inst_pe_1_2_3_add_69_carry_4_,
         npu_inst_pe_1_2_3_add_69_carry_3_, npu_inst_pe_1_2_3_add_69_carry_2_,
         npu_inst_pe_1_2_3_add_69_carry_1_, npu_inst_pe_1_2_3_n97,
         npu_inst_pe_1_2_3_n96, npu_inst_pe_1_2_3_n95, npu_inst_pe_1_2_3_n94,
         npu_inst_pe_1_2_3_n93, npu_inst_pe_1_2_3_n92, npu_inst_pe_1_2_3_n91,
         npu_inst_pe_1_2_3_n90, npu_inst_pe_1_2_3_n89, npu_inst_pe_1_2_3_n88,
         npu_inst_pe_1_2_3_n87, npu_inst_pe_1_2_3_n86, npu_inst_pe_1_2_3_n85,
         npu_inst_pe_1_2_3_n84, npu_inst_pe_1_2_3_n83, npu_inst_pe_1_2_3_n82,
         npu_inst_pe_1_2_3_n81, npu_inst_pe_1_2_3_n80, npu_inst_pe_1_2_3_n79,
         npu_inst_pe_1_2_3_n78, npu_inst_pe_1_2_3_n77, npu_inst_pe_1_2_3_n76,
         npu_inst_pe_1_2_3_n75, npu_inst_pe_1_2_3_n74, npu_inst_pe_1_2_3_n73,
         npu_inst_pe_1_2_3_n72, npu_inst_pe_1_2_3_n71, npu_inst_pe_1_2_3_n70,
         npu_inst_pe_1_2_3_n69, npu_inst_pe_1_2_3_n68, npu_inst_pe_1_2_3_n67,
         npu_inst_pe_1_2_3_n66, npu_inst_pe_1_2_3_n65, npu_inst_pe_1_2_3_n64,
         npu_inst_pe_1_2_3_n63, npu_inst_pe_1_2_3_n62, npu_inst_pe_1_2_3_n61,
         npu_inst_pe_1_2_3_n60, npu_inst_pe_1_2_3_n59, npu_inst_pe_1_2_3_n58,
         npu_inst_pe_1_2_3_n57, npu_inst_pe_1_2_3_n56, npu_inst_pe_1_2_3_n55,
         npu_inst_pe_1_2_3_n54, npu_inst_pe_1_2_3_n53, npu_inst_pe_1_2_3_n52,
         npu_inst_pe_1_2_3_n51, npu_inst_pe_1_2_3_n50, npu_inst_pe_1_2_3_n49,
         npu_inst_pe_1_2_3_n48, npu_inst_pe_1_2_3_n47, npu_inst_pe_1_2_3_n46,
         npu_inst_pe_1_2_3_n45, npu_inst_pe_1_2_3_n44, npu_inst_pe_1_2_3_n43,
         npu_inst_pe_1_2_3_n42, npu_inst_pe_1_2_3_n41, npu_inst_pe_1_2_3_n40,
         npu_inst_pe_1_2_3_n39, npu_inst_pe_1_2_3_n38, npu_inst_pe_1_2_3_n37,
         npu_inst_pe_1_2_3_n27, npu_inst_pe_1_2_3_n26,
         npu_inst_pe_1_2_3_net4131, npu_inst_pe_1_2_3_net4125,
         npu_inst_pe_1_2_3_N94, npu_inst_pe_1_2_3_N93, npu_inst_pe_1_2_3_N84,
         npu_inst_pe_1_2_3_N80, npu_inst_pe_1_2_3_N79, npu_inst_pe_1_2_3_N78,
         npu_inst_pe_1_2_3_N77, npu_inst_pe_1_2_3_N76, npu_inst_pe_1_2_3_N75,
         npu_inst_pe_1_2_3_N74, npu_inst_pe_1_2_3_N73, npu_inst_pe_1_2_3_N72,
         npu_inst_pe_1_2_3_N71, npu_inst_pe_1_2_3_N70, npu_inst_pe_1_2_3_N69,
         npu_inst_pe_1_2_3_N68, npu_inst_pe_1_2_3_N67, npu_inst_pe_1_2_3_N66,
         npu_inst_pe_1_2_3_N65, npu_inst_pe_1_2_3_int_q_acc_0_,
         npu_inst_pe_1_2_3_int_q_acc_1_, npu_inst_pe_1_2_3_int_q_acc_2_,
         npu_inst_pe_1_2_3_int_q_acc_3_, npu_inst_pe_1_2_3_int_q_acc_4_,
         npu_inst_pe_1_2_3_int_q_acc_5_, npu_inst_pe_1_2_3_int_q_acc_6_,
         npu_inst_pe_1_2_3_int_q_acc_7_, npu_inst_pe_1_2_3_int_data_0_,
         npu_inst_pe_1_2_3_int_data_1_, npu_inst_pe_1_2_3_int_q_weight_0_,
         npu_inst_pe_1_2_3_int_q_weight_1_,
         npu_inst_pe_1_2_3_int_q_reg_v_5__0_,
         npu_inst_pe_1_2_3_int_q_reg_v_5__1_,
         npu_inst_pe_1_2_3_int_q_reg_v_4__0_,
         npu_inst_pe_1_2_3_int_q_reg_v_4__1_,
         npu_inst_pe_1_2_3_int_q_reg_v_3__0_,
         npu_inst_pe_1_2_3_int_q_reg_v_3__1_,
         npu_inst_pe_1_2_3_int_q_reg_v_2__0_,
         npu_inst_pe_1_2_3_int_q_reg_v_2__1_,
         npu_inst_pe_1_2_3_int_q_reg_v_1__0_,
         npu_inst_pe_1_2_3_int_q_reg_v_1__1_,
         npu_inst_pe_1_2_3_int_q_reg_v_0__0_,
         npu_inst_pe_1_2_3_int_q_reg_v_0__1_,
         npu_inst_pe_1_2_3_int_q_reg_h_5__0_,
         npu_inst_pe_1_2_3_int_q_reg_h_5__1_,
         npu_inst_pe_1_2_3_int_q_reg_h_4__0_,
         npu_inst_pe_1_2_3_int_q_reg_h_4__1_,
         npu_inst_pe_1_2_3_int_q_reg_h_3__0_,
         npu_inst_pe_1_2_3_int_q_reg_h_3__1_,
         npu_inst_pe_1_2_3_int_q_reg_h_2__0_,
         npu_inst_pe_1_2_3_int_q_reg_h_2__1_,
         npu_inst_pe_1_2_3_int_q_reg_h_1__0_,
         npu_inst_pe_1_2_3_int_q_reg_h_1__1_,
         npu_inst_pe_1_2_3_int_q_reg_h_0__0_,
         npu_inst_pe_1_2_3_int_q_reg_h_0__1_, npu_inst_pe_1_2_4_n119,
         npu_inst_pe_1_2_4_n118, npu_inst_pe_1_2_4_n117,
         npu_inst_pe_1_2_4_n116, npu_inst_pe_1_2_4_n115,
         npu_inst_pe_1_2_4_n114, npu_inst_pe_1_2_4_n113,
         npu_inst_pe_1_2_4_n112, npu_inst_pe_1_2_4_n111,
         npu_inst_pe_1_2_4_n110, npu_inst_pe_1_2_4_n109,
         npu_inst_pe_1_2_4_n108, npu_inst_pe_1_2_4_n107,
         npu_inst_pe_1_2_4_n106, npu_inst_pe_1_2_4_n105,
         npu_inst_pe_1_2_4_n104, npu_inst_pe_1_2_4_n103,
         npu_inst_pe_1_2_4_n102, npu_inst_pe_1_2_4_n101,
         npu_inst_pe_1_2_4_n100, npu_inst_pe_1_2_4_n99, npu_inst_pe_1_2_4_n98,
         npu_inst_pe_1_2_4_n36, npu_inst_pe_1_2_4_n35, npu_inst_pe_1_2_4_n34,
         npu_inst_pe_1_2_4_n33, npu_inst_pe_1_2_4_n32, npu_inst_pe_1_2_4_n31,
         npu_inst_pe_1_2_4_n30, npu_inst_pe_1_2_4_n29, npu_inst_pe_1_2_4_n28,
         npu_inst_pe_1_2_4_n25, npu_inst_pe_1_2_4_n24, npu_inst_pe_1_2_4_n23,
         npu_inst_pe_1_2_4_n22, npu_inst_pe_1_2_4_n21, npu_inst_pe_1_2_4_n20,
         npu_inst_pe_1_2_4_n19, npu_inst_pe_1_2_4_n18, npu_inst_pe_1_2_4_n17,
         npu_inst_pe_1_2_4_n16, npu_inst_pe_1_2_4_n15, npu_inst_pe_1_2_4_n14,
         npu_inst_pe_1_2_4_n13, npu_inst_pe_1_2_4_n12, npu_inst_pe_1_2_4_n11,
         npu_inst_pe_1_2_4_n10, npu_inst_pe_1_2_4_n9, npu_inst_pe_1_2_4_n8,
         npu_inst_pe_1_2_4_n7, npu_inst_pe_1_2_4_n6, npu_inst_pe_1_2_4_n5,
         npu_inst_pe_1_2_4_n4, npu_inst_pe_1_2_4_n3, npu_inst_pe_1_2_4_n2,
         npu_inst_pe_1_2_4_n1, npu_inst_pe_1_2_4_sub_67_carry_7_,
         npu_inst_pe_1_2_4_sub_67_carry_6_, npu_inst_pe_1_2_4_sub_67_carry_5_,
         npu_inst_pe_1_2_4_sub_67_carry_4_, npu_inst_pe_1_2_4_sub_67_carry_3_,
         npu_inst_pe_1_2_4_sub_67_carry_2_, npu_inst_pe_1_2_4_sub_67_carry_1_,
         npu_inst_pe_1_2_4_add_69_carry_7_, npu_inst_pe_1_2_4_add_69_carry_6_,
         npu_inst_pe_1_2_4_add_69_carry_5_, npu_inst_pe_1_2_4_add_69_carry_4_,
         npu_inst_pe_1_2_4_add_69_carry_3_, npu_inst_pe_1_2_4_add_69_carry_2_,
         npu_inst_pe_1_2_4_add_69_carry_1_, npu_inst_pe_1_2_4_n97,
         npu_inst_pe_1_2_4_n96, npu_inst_pe_1_2_4_n95, npu_inst_pe_1_2_4_n94,
         npu_inst_pe_1_2_4_n93, npu_inst_pe_1_2_4_n92, npu_inst_pe_1_2_4_n91,
         npu_inst_pe_1_2_4_n90, npu_inst_pe_1_2_4_n89, npu_inst_pe_1_2_4_n88,
         npu_inst_pe_1_2_4_n87, npu_inst_pe_1_2_4_n86, npu_inst_pe_1_2_4_n85,
         npu_inst_pe_1_2_4_n84, npu_inst_pe_1_2_4_n83, npu_inst_pe_1_2_4_n82,
         npu_inst_pe_1_2_4_n81, npu_inst_pe_1_2_4_n80, npu_inst_pe_1_2_4_n79,
         npu_inst_pe_1_2_4_n78, npu_inst_pe_1_2_4_n77, npu_inst_pe_1_2_4_n76,
         npu_inst_pe_1_2_4_n75, npu_inst_pe_1_2_4_n74, npu_inst_pe_1_2_4_n73,
         npu_inst_pe_1_2_4_n72, npu_inst_pe_1_2_4_n71, npu_inst_pe_1_2_4_n70,
         npu_inst_pe_1_2_4_n69, npu_inst_pe_1_2_4_n68, npu_inst_pe_1_2_4_n67,
         npu_inst_pe_1_2_4_n66, npu_inst_pe_1_2_4_n65, npu_inst_pe_1_2_4_n64,
         npu_inst_pe_1_2_4_n63, npu_inst_pe_1_2_4_n62, npu_inst_pe_1_2_4_n61,
         npu_inst_pe_1_2_4_n60, npu_inst_pe_1_2_4_n59, npu_inst_pe_1_2_4_n58,
         npu_inst_pe_1_2_4_n57, npu_inst_pe_1_2_4_n56, npu_inst_pe_1_2_4_n55,
         npu_inst_pe_1_2_4_n54, npu_inst_pe_1_2_4_n53, npu_inst_pe_1_2_4_n52,
         npu_inst_pe_1_2_4_n51, npu_inst_pe_1_2_4_n50, npu_inst_pe_1_2_4_n49,
         npu_inst_pe_1_2_4_n48, npu_inst_pe_1_2_4_n47, npu_inst_pe_1_2_4_n46,
         npu_inst_pe_1_2_4_n45, npu_inst_pe_1_2_4_n44, npu_inst_pe_1_2_4_n43,
         npu_inst_pe_1_2_4_n42, npu_inst_pe_1_2_4_n41, npu_inst_pe_1_2_4_n40,
         npu_inst_pe_1_2_4_n39, npu_inst_pe_1_2_4_n38, npu_inst_pe_1_2_4_n37,
         npu_inst_pe_1_2_4_n27, npu_inst_pe_1_2_4_n26,
         npu_inst_pe_1_2_4_net4108, npu_inst_pe_1_2_4_net4102,
         npu_inst_pe_1_2_4_N94, npu_inst_pe_1_2_4_N93, npu_inst_pe_1_2_4_N84,
         npu_inst_pe_1_2_4_N80, npu_inst_pe_1_2_4_N79, npu_inst_pe_1_2_4_N78,
         npu_inst_pe_1_2_4_N77, npu_inst_pe_1_2_4_N76, npu_inst_pe_1_2_4_N75,
         npu_inst_pe_1_2_4_N74, npu_inst_pe_1_2_4_N73, npu_inst_pe_1_2_4_N72,
         npu_inst_pe_1_2_4_N71, npu_inst_pe_1_2_4_N70, npu_inst_pe_1_2_4_N69,
         npu_inst_pe_1_2_4_N68, npu_inst_pe_1_2_4_N67, npu_inst_pe_1_2_4_N66,
         npu_inst_pe_1_2_4_N65, npu_inst_pe_1_2_4_int_q_acc_0_,
         npu_inst_pe_1_2_4_int_q_acc_1_, npu_inst_pe_1_2_4_int_q_acc_2_,
         npu_inst_pe_1_2_4_int_q_acc_3_, npu_inst_pe_1_2_4_int_q_acc_4_,
         npu_inst_pe_1_2_4_int_q_acc_5_, npu_inst_pe_1_2_4_int_q_acc_6_,
         npu_inst_pe_1_2_4_int_q_acc_7_, npu_inst_pe_1_2_4_int_data_0_,
         npu_inst_pe_1_2_4_int_data_1_, npu_inst_pe_1_2_4_int_q_weight_0_,
         npu_inst_pe_1_2_4_int_q_weight_1_,
         npu_inst_pe_1_2_4_int_q_reg_v_5__0_,
         npu_inst_pe_1_2_4_int_q_reg_v_5__1_,
         npu_inst_pe_1_2_4_int_q_reg_v_4__0_,
         npu_inst_pe_1_2_4_int_q_reg_v_4__1_,
         npu_inst_pe_1_2_4_int_q_reg_v_3__0_,
         npu_inst_pe_1_2_4_int_q_reg_v_3__1_,
         npu_inst_pe_1_2_4_int_q_reg_v_2__0_,
         npu_inst_pe_1_2_4_int_q_reg_v_2__1_,
         npu_inst_pe_1_2_4_int_q_reg_v_1__0_,
         npu_inst_pe_1_2_4_int_q_reg_v_1__1_,
         npu_inst_pe_1_2_4_int_q_reg_v_0__0_,
         npu_inst_pe_1_2_4_int_q_reg_v_0__1_,
         npu_inst_pe_1_2_4_int_q_reg_h_5__0_,
         npu_inst_pe_1_2_4_int_q_reg_h_5__1_,
         npu_inst_pe_1_2_4_int_q_reg_h_4__0_,
         npu_inst_pe_1_2_4_int_q_reg_h_4__1_,
         npu_inst_pe_1_2_4_int_q_reg_h_3__0_,
         npu_inst_pe_1_2_4_int_q_reg_h_3__1_,
         npu_inst_pe_1_2_4_int_q_reg_h_2__0_,
         npu_inst_pe_1_2_4_int_q_reg_h_2__1_,
         npu_inst_pe_1_2_4_int_q_reg_h_1__0_,
         npu_inst_pe_1_2_4_int_q_reg_h_1__1_,
         npu_inst_pe_1_2_4_int_q_reg_h_0__0_,
         npu_inst_pe_1_2_4_int_q_reg_h_0__1_, npu_inst_pe_1_2_5_n119,
         npu_inst_pe_1_2_5_n118, npu_inst_pe_1_2_5_n117,
         npu_inst_pe_1_2_5_n116, npu_inst_pe_1_2_5_n115,
         npu_inst_pe_1_2_5_n114, npu_inst_pe_1_2_5_n113,
         npu_inst_pe_1_2_5_n112, npu_inst_pe_1_2_5_n111,
         npu_inst_pe_1_2_5_n110, npu_inst_pe_1_2_5_n109,
         npu_inst_pe_1_2_5_n108, npu_inst_pe_1_2_5_n107,
         npu_inst_pe_1_2_5_n106, npu_inst_pe_1_2_5_n105,
         npu_inst_pe_1_2_5_n104, npu_inst_pe_1_2_5_n103,
         npu_inst_pe_1_2_5_n102, npu_inst_pe_1_2_5_n101,
         npu_inst_pe_1_2_5_n100, npu_inst_pe_1_2_5_n99, npu_inst_pe_1_2_5_n98,
         npu_inst_pe_1_2_5_n36, npu_inst_pe_1_2_5_n35, npu_inst_pe_1_2_5_n34,
         npu_inst_pe_1_2_5_n33, npu_inst_pe_1_2_5_n32, npu_inst_pe_1_2_5_n31,
         npu_inst_pe_1_2_5_n30, npu_inst_pe_1_2_5_n29, npu_inst_pe_1_2_5_n28,
         npu_inst_pe_1_2_5_n25, npu_inst_pe_1_2_5_n24, npu_inst_pe_1_2_5_n23,
         npu_inst_pe_1_2_5_n22, npu_inst_pe_1_2_5_n21, npu_inst_pe_1_2_5_n20,
         npu_inst_pe_1_2_5_n19, npu_inst_pe_1_2_5_n18, npu_inst_pe_1_2_5_n17,
         npu_inst_pe_1_2_5_n16, npu_inst_pe_1_2_5_n15, npu_inst_pe_1_2_5_n14,
         npu_inst_pe_1_2_5_n13, npu_inst_pe_1_2_5_n12, npu_inst_pe_1_2_5_n11,
         npu_inst_pe_1_2_5_n10, npu_inst_pe_1_2_5_n9, npu_inst_pe_1_2_5_n8,
         npu_inst_pe_1_2_5_n7, npu_inst_pe_1_2_5_n6, npu_inst_pe_1_2_5_n5,
         npu_inst_pe_1_2_5_n4, npu_inst_pe_1_2_5_n3, npu_inst_pe_1_2_5_n2,
         npu_inst_pe_1_2_5_n1, npu_inst_pe_1_2_5_sub_67_carry_7_,
         npu_inst_pe_1_2_5_sub_67_carry_6_, npu_inst_pe_1_2_5_sub_67_carry_5_,
         npu_inst_pe_1_2_5_sub_67_carry_4_, npu_inst_pe_1_2_5_sub_67_carry_3_,
         npu_inst_pe_1_2_5_sub_67_carry_2_, npu_inst_pe_1_2_5_sub_67_carry_1_,
         npu_inst_pe_1_2_5_add_69_carry_7_, npu_inst_pe_1_2_5_add_69_carry_6_,
         npu_inst_pe_1_2_5_add_69_carry_5_, npu_inst_pe_1_2_5_add_69_carry_4_,
         npu_inst_pe_1_2_5_add_69_carry_3_, npu_inst_pe_1_2_5_add_69_carry_2_,
         npu_inst_pe_1_2_5_add_69_carry_1_, npu_inst_pe_1_2_5_n97,
         npu_inst_pe_1_2_5_n96, npu_inst_pe_1_2_5_n95, npu_inst_pe_1_2_5_n94,
         npu_inst_pe_1_2_5_n93, npu_inst_pe_1_2_5_n92, npu_inst_pe_1_2_5_n91,
         npu_inst_pe_1_2_5_n90, npu_inst_pe_1_2_5_n89, npu_inst_pe_1_2_5_n88,
         npu_inst_pe_1_2_5_n87, npu_inst_pe_1_2_5_n86, npu_inst_pe_1_2_5_n85,
         npu_inst_pe_1_2_5_n84, npu_inst_pe_1_2_5_n83, npu_inst_pe_1_2_5_n82,
         npu_inst_pe_1_2_5_n81, npu_inst_pe_1_2_5_n80, npu_inst_pe_1_2_5_n79,
         npu_inst_pe_1_2_5_n78, npu_inst_pe_1_2_5_n77, npu_inst_pe_1_2_5_n76,
         npu_inst_pe_1_2_5_n75, npu_inst_pe_1_2_5_n74, npu_inst_pe_1_2_5_n73,
         npu_inst_pe_1_2_5_n72, npu_inst_pe_1_2_5_n71, npu_inst_pe_1_2_5_n70,
         npu_inst_pe_1_2_5_n69, npu_inst_pe_1_2_5_n68, npu_inst_pe_1_2_5_n67,
         npu_inst_pe_1_2_5_n66, npu_inst_pe_1_2_5_n65, npu_inst_pe_1_2_5_n64,
         npu_inst_pe_1_2_5_n63, npu_inst_pe_1_2_5_n62, npu_inst_pe_1_2_5_n61,
         npu_inst_pe_1_2_5_n60, npu_inst_pe_1_2_5_n59, npu_inst_pe_1_2_5_n58,
         npu_inst_pe_1_2_5_n57, npu_inst_pe_1_2_5_n56, npu_inst_pe_1_2_5_n55,
         npu_inst_pe_1_2_5_n54, npu_inst_pe_1_2_5_n53, npu_inst_pe_1_2_5_n52,
         npu_inst_pe_1_2_5_n51, npu_inst_pe_1_2_5_n50, npu_inst_pe_1_2_5_n49,
         npu_inst_pe_1_2_5_n48, npu_inst_pe_1_2_5_n47, npu_inst_pe_1_2_5_n46,
         npu_inst_pe_1_2_5_n45, npu_inst_pe_1_2_5_n44, npu_inst_pe_1_2_5_n43,
         npu_inst_pe_1_2_5_n42, npu_inst_pe_1_2_5_n41, npu_inst_pe_1_2_5_n40,
         npu_inst_pe_1_2_5_n39, npu_inst_pe_1_2_5_n38, npu_inst_pe_1_2_5_n37,
         npu_inst_pe_1_2_5_n27, npu_inst_pe_1_2_5_n26,
         npu_inst_pe_1_2_5_net4085, npu_inst_pe_1_2_5_net4079,
         npu_inst_pe_1_2_5_N94, npu_inst_pe_1_2_5_N93, npu_inst_pe_1_2_5_N84,
         npu_inst_pe_1_2_5_N80, npu_inst_pe_1_2_5_N79, npu_inst_pe_1_2_5_N78,
         npu_inst_pe_1_2_5_N77, npu_inst_pe_1_2_5_N76, npu_inst_pe_1_2_5_N75,
         npu_inst_pe_1_2_5_N74, npu_inst_pe_1_2_5_N73, npu_inst_pe_1_2_5_N72,
         npu_inst_pe_1_2_5_N71, npu_inst_pe_1_2_5_N70, npu_inst_pe_1_2_5_N69,
         npu_inst_pe_1_2_5_N68, npu_inst_pe_1_2_5_N67, npu_inst_pe_1_2_5_N66,
         npu_inst_pe_1_2_5_N65, npu_inst_pe_1_2_5_int_q_acc_0_,
         npu_inst_pe_1_2_5_int_q_acc_1_, npu_inst_pe_1_2_5_int_q_acc_2_,
         npu_inst_pe_1_2_5_int_q_acc_3_, npu_inst_pe_1_2_5_int_q_acc_4_,
         npu_inst_pe_1_2_5_int_q_acc_5_, npu_inst_pe_1_2_5_int_q_acc_6_,
         npu_inst_pe_1_2_5_int_q_acc_7_, npu_inst_pe_1_2_5_int_data_0_,
         npu_inst_pe_1_2_5_int_data_1_, npu_inst_pe_1_2_5_int_q_weight_0_,
         npu_inst_pe_1_2_5_int_q_weight_1_,
         npu_inst_pe_1_2_5_int_q_reg_v_5__0_,
         npu_inst_pe_1_2_5_int_q_reg_v_5__1_,
         npu_inst_pe_1_2_5_int_q_reg_v_4__0_,
         npu_inst_pe_1_2_5_int_q_reg_v_4__1_,
         npu_inst_pe_1_2_5_int_q_reg_v_3__0_,
         npu_inst_pe_1_2_5_int_q_reg_v_3__1_,
         npu_inst_pe_1_2_5_int_q_reg_v_2__0_,
         npu_inst_pe_1_2_5_int_q_reg_v_2__1_,
         npu_inst_pe_1_2_5_int_q_reg_v_1__0_,
         npu_inst_pe_1_2_5_int_q_reg_v_1__1_,
         npu_inst_pe_1_2_5_int_q_reg_v_0__0_,
         npu_inst_pe_1_2_5_int_q_reg_v_0__1_,
         npu_inst_pe_1_2_5_int_q_reg_h_5__0_,
         npu_inst_pe_1_2_5_int_q_reg_h_5__1_,
         npu_inst_pe_1_2_5_int_q_reg_h_4__0_,
         npu_inst_pe_1_2_5_int_q_reg_h_4__1_,
         npu_inst_pe_1_2_5_int_q_reg_h_3__0_,
         npu_inst_pe_1_2_5_int_q_reg_h_3__1_,
         npu_inst_pe_1_2_5_int_q_reg_h_2__0_,
         npu_inst_pe_1_2_5_int_q_reg_h_2__1_,
         npu_inst_pe_1_2_5_int_q_reg_h_1__0_,
         npu_inst_pe_1_2_5_int_q_reg_h_1__1_,
         npu_inst_pe_1_2_5_int_q_reg_h_0__0_,
         npu_inst_pe_1_2_5_int_q_reg_h_0__1_, npu_inst_pe_1_2_6_n119,
         npu_inst_pe_1_2_6_n118, npu_inst_pe_1_2_6_n117,
         npu_inst_pe_1_2_6_n116, npu_inst_pe_1_2_6_n115,
         npu_inst_pe_1_2_6_n114, npu_inst_pe_1_2_6_n113,
         npu_inst_pe_1_2_6_n112, npu_inst_pe_1_2_6_n111,
         npu_inst_pe_1_2_6_n110, npu_inst_pe_1_2_6_n109,
         npu_inst_pe_1_2_6_n108, npu_inst_pe_1_2_6_n107,
         npu_inst_pe_1_2_6_n106, npu_inst_pe_1_2_6_n105,
         npu_inst_pe_1_2_6_n104, npu_inst_pe_1_2_6_n103,
         npu_inst_pe_1_2_6_n102, npu_inst_pe_1_2_6_n101,
         npu_inst_pe_1_2_6_n100, npu_inst_pe_1_2_6_n99, npu_inst_pe_1_2_6_n98,
         npu_inst_pe_1_2_6_n36, npu_inst_pe_1_2_6_n35, npu_inst_pe_1_2_6_n34,
         npu_inst_pe_1_2_6_n33, npu_inst_pe_1_2_6_n32, npu_inst_pe_1_2_6_n31,
         npu_inst_pe_1_2_6_n30, npu_inst_pe_1_2_6_n29, npu_inst_pe_1_2_6_n28,
         npu_inst_pe_1_2_6_n25, npu_inst_pe_1_2_6_n24, npu_inst_pe_1_2_6_n23,
         npu_inst_pe_1_2_6_n22, npu_inst_pe_1_2_6_n21, npu_inst_pe_1_2_6_n20,
         npu_inst_pe_1_2_6_n19, npu_inst_pe_1_2_6_n18, npu_inst_pe_1_2_6_n17,
         npu_inst_pe_1_2_6_n16, npu_inst_pe_1_2_6_n15, npu_inst_pe_1_2_6_n14,
         npu_inst_pe_1_2_6_n13, npu_inst_pe_1_2_6_n12, npu_inst_pe_1_2_6_n11,
         npu_inst_pe_1_2_6_n10, npu_inst_pe_1_2_6_n9, npu_inst_pe_1_2_6_n8,
         npu_inst_pe_1_2_6_n7, npu_inst_pe_1_2_6_n6, npu_inst_pe_1_2_6_n5,
         npu_inst_pe_1_2_6_n4, npu_inst_pe_1_2_6_n3, npu_inst_pe_1_2_6_n2,
         npu_inst_pe_1_2_6_n1, npu_inst_pe_1_2_6_sub_67_carry_7_,
         npu_inst_pe_1_2_6_sub_67_carry_6_, npu_inst_pe_1_2_6_sub_67_carry_5_,
         npu_inst_pe_1_2_6_sub_67_carry_4_, npu_inst_pe_1_2_6_sub_67_carry_3_,
         npu_inst_pe_1_2_6_sub_67_carry_2_, npu_inst_pe_1_2_6_sub_67_carry_1_,
         npu_inst_pe_1_2_6_add_69_carry_7_, npu_inst_pe_1_2_6_add_69_carry_6_,
         npu_inst_pe_1_2_6_add_69_carry_5_, npu_inst_pe_1_2_6_add_69_carry_4_,
         npu_inst_pe_1_2_6_add_69_carry_3_, npu_inst_pe_1_2_6_add_69_carry_2_,
         npu_inst_pe_1_2_6_add_69_carry_1_, npu_inst_pe_1_2_6_n97,
         npu_inst_pe_1_2_6_n96, npu_inst_pe_1_2_6_n95, npu_inst_pe_1_2_6_n94,
         npu_inst_pe_1_2_6_n93, npu_inst_pe_1_2_6_n92, npu_inst_pe_1_2_6_n91,
         npu_inst_pe_1_2_6_n90, npu_inst_pe_1_2_6_n89, npu_inst_pe_1_2_6_n88,
         npu_inst_pe_1_2_6_n87, npu_inst_pe_1_2_6_n86, npu_inst_pe_1_2_6_n85,
         npu_inst_pe_1_2_6_n84, npu_inst_pe_1_2_6_n83, npu_inst_pe_1_2_6_n82,
         npu_inst_pe_1_2_6_n81, npu_inst_pe_1_2_6_n80, npu_inst_pe_1_2_6_n79,
         npu_inst_pe_1_2_6_n78, npu_inst_pe_1_2_6_n77, npu_inst_pe_1_2_6_n76,
         npu_inst_pe_1_2_6_n75, npu_inst_pe_1_2_6_n74, npu_inst_pe_1_2_6_n73,
         npu_inst_pe_1_2_6_n72, npu_inst_pe_1_2_6_n71, npu_inst_pe_1_2_6_n70,
         npu_inst_pe_1_2_6_n69, npu_inst_pe_1_2_6_n68, npu_inst_pe_1_2_6_n67,
         npu_inst_pe_1_2_6_n66, npu_inst_pe_1_2_6_n65, npu_inst_pe_1_2_6_n64,
         npu_inst_pe_1_2_6_n63, npu_inst_pe_1_2_6_n62, npu_inst_pe_1_2_6_n61,
         npu_inst_pe_1_2_6_n60, npu_inst_pe_1_2_6_n59, npu_inst_pe_1_2_6_n58,
         npu_inst_pe_1_2_6_n57, npu_inst_pe_1_2_6_n56, npu_inst_pe_1_2_6_n55,
         npu_inst_pe_1_2_6_n54, npu_inst_pe_1_2_6_n53, npu_inst_pe_1_2_6_n52,
         npu_inst_pe_1_2_6_n51, npu_inst_pe_1_2_6_n50, npu_inst_pe_1_2_6_n49,
         npu_inst_pe_1_2_6_n48, npu_inst_pe_1_2_6_n47, npu_inst_pe_1_2_6_n46,
         npu_inst_pe_1_2_6_n45, npu_inst_pe_1_2_6_n44, npu_inst_pe_1_2_6_n43,
         npu_inst_pe_1_2_6_n42, npu_inst_pe_1_2_6_n41, npu_inst_pe_1_2_6_n40,
         npu_inst_pe_1_2_6_n39, npu_inst_pe_1_2_6_n38, npu_inst_pe_1_2_6_n37,
         npu_inst_pe_1_2_6_n27, npu_inst_pe_1_2_6_n26,
         npu_inst_pe_1_2_6_net4062, npu_inst_pe_1_2_6_net4056,
         npu_inst_pe_1_2_6_N94, npu_inst_pe_1_2_6_N93, npu_inst_pe_1_2_6_N84,
         npu_inst_pe_1_2_6_N80, npu_inst_pe_1_2_6_N79, npu_inst_pe_1_2_6_N78,
         npu_inst_pe_1_2_6_N77, npu_inst_pe_1_2_6_N76, npu_inst_pe_1_2_6_N75,
         npu_inst_pe_1_2_6_N74, npu_inst_pe_1_2_6_N73, npu_inst_pe_1_2_6_N72,
         npu_inst_pe_1_2_6_N71, npu_inst_pe_1_2_6_N70, npu_inst_pe_1_2_6_N69,
         npu_inst_pe_1_2_6_N68, npu_inst_pe_1_2_6_N67, npu_inst_pe_1_2_6_N66,
         npu_inst_pe_1_2_6_N65, npu_inst_pe_1_2_6_int_q_acc_0_,
         npu_inst_pe_1_2_6_int_q_acc_1_, npu_inst_pe_1_2_6_int_q_acc_2_,
         npu_inst_pe_1_2_6_int_q_acc_3_, npu_inst_pe_1_2_6_int_q_acc_4_,
         npu_inst_pe_1_2_6_int_q_acc_5_, npu_inst_pe_1_2_6_int_q_acc_6_,
         npu_inst_pe_1_2_6_int_q_acc_7_, npu_inst_pe_1_2_6_int_data_0_,
         npu_inst_pe_1_2_6_int_data_1_, npu_inst_pe_1_2_6_int_q_weight_0_,
         npu_inst_pe_1_2_6_int_q_weight_1_,
         npu_inst_pe_1_2_6_int_q_reg_v_5__0_,
         npu_inst_pe_1_2_6_int_q_reg_v_5__1_,
         npu_inst_pe_1_2_6_int_q_reg_v_4__0_,
         npu_inst_pe_1_2_6_int_q_reg_v_4__1_,
         npu_inst_pe_1_2_6_int_q_reg_v_3__0_,
         npu_inst_pe_1_2_6_int_q_reg_v_3__1_,
         npu_inst_pe_1_2_6_int_q_reg_v_2__0_,
         npu_inst_pe_1_2_6_int_q_reg_v_2__1_,
         npu_inst_pe_1_2_6_int_q_reg_v_1__0_,
         npu_inst_pe_1_2_6_int_q_reg_v_1__1_,
         npu_inst_pe_1_2_6_int_q_reg_v_0__0_,
         npu_inst_pe_1_2_6_int_q_reg_v_0__1_,
         npu_inst_pe_1_2_6_int_q_reg_h_5__0_,
         npu_inst_pe_1_2_6_int_q_reg_h_5__1_,
         npu_inst_pe_1_2_6_int_q_reg_h_4__0_,
         npu_inst_pe_1_2_6_int_q_reg_h_4__1_,
         npu_inst_pe_1_2_6_int_q_reg_h_3__0_,
         npu_inst_pe_1_2_6_int_q_reg_h_3__1_,
         npu_inst_pe_1_2_6_int_q_reg_h_2__0_,
         npu_inst_pe_1_2_6_int_q_reg_h_2__1_,
         npu_inst_pe_1_2_6_int_q_reg_h_1__0_,
         npu_inst_pe_1_2_6_int_q_reg_h_1__1_,
         npu_inst_pe_1_2_6_int_q_reg_h_0__0_,
         npu_inst_pe_1_2_6_int_q_reg_h_0__1_, npu_inst_pe_1_2_7_n119,
         npu_inst_pe_1_2_7_n118, npu_inst_pe_1_2_7_n117,
         npu_inst_pe_1_2_7_n116, npu_inst_pe_1_2_7_n115,
         npu_inst_pe_1_2_7_n114, npu_inst_pe_1_2_7_n113,
         npu_inst_pe_1_2_7_n112, npu_inst_pe_1_2_7_n111,
         npu_inst_pe_1_2_7_n110, npu_inst_pe_1_2_7_n109,
         npu_inst_pe_1_2_7_n108, npu_inst_pe_1_2_7_n107,
         npu_inst_pe_1_2_7_n106, npu_inst_pe_1_2_7_n105,
         npu_inst_pe_1_2_7_n104, npu_inst_pe_1_2_7_n103,
         npu_inst_pe_1_2_7_n102, npu_inst_pe_1_2_7_n101,
         npu_inst_pe_1_2_7_n100, npu_inst_pe_1_2_7_n99, npu_inst_pe_1_2_7_n98,
         npu_inst_pe_1_2_7_n36, npu_inst_pe_1_2_7_n35, npu_inst_pe_1_2_7_n34,
         npu_inst_pe_1_2_7_n33, npu_inst_pe_1_2_7_n32, npu_inst_pe_1_2_7_n31,
         npu_inst_pe_1_2_7_n30, npu_inst_pe_1_2_7_n29, npu_inst_pe_1_2_7_n28,
         npu_inst_pe_1_2_7_n25, npu_inst_pe_1_2_7_n24, npu_inst_pe_1_2_7_n23,
         npu_inst_pe_1_2_7_n22, npu_inst_pe_1_2_7_n21, npu_inst_pe_1_2_7_n20,
         npu_inst_pe_1_2_7_n19, npu_inst_pe_1_2_7_n18, npu_inst_pe_1_2_7_n17,
         npu_inst_pe_1_2_7_n16, npu_inst_pe_1_2_7_n15, npu_inst_pe_1_2_7_n14,
         npu_inst_pe_1_2_7_n13, npu_inst_pe_1_2_7_n12, npu_inst_pe_1_2_7_n11,
         npu_inst_pe_1_2_7_n10, npu_inst_pe_1_2_7_n9, npu_inst_pe_1_2_7_n8,
         npu_inst_pe_1_2_7_n7, npu_inst_pe_1_2_7_n6, npu_inst_pe_1_2_7_n5,
         npu_inst_pe_1_2_7_n4, npu_inst_pe_1_2_7_n3, npu_inst_pe_1_2_7_n2,
         npu_inst_pe_1_2_7_n1, npu_inst_pe_1_2_7_sub_67_carry_7_,
         npu_inst_pe_1_2_7_sub_67_carry_6_, npu_inst_pe_1_2_7_sub_67_carry_5_,
         npu_inst_pe_1_2_7_sub_67_carry_4_, npu_inst_pe_1_2_7_sub_67_carry_3_,
         npu_inst_pe_1_2_7_sub_67_carry_2_, npu_inst_pe_1_2_7_sub_67_carry_1_,
         npu_inst_pe_1_2_7_add_69_carry_7_, npu_inst_pe_1_2_7_add_69_carry_6_,
         npu_inst_pe_1_2_7_add_69_carry_5_, npu_inst_pe_1_2_7_add_69_carry_4_,
         npu_inst_pe_1_2_7_add_69_carry_3_, npu_inst_pe_1_2_7_add_69_carry_2_,
         npu_inst_pe_1_2_7_add_69_carry_1_, npu_inst_pe_1_2_7_n97,
         npu_inst_pe_1_2_7_n96, npu_inst_pe_1_2_7_n95, npu_inst_pe_1_2_7_n94,
         npu_inst_pe_1_2_7_n93, npu_inst_pe_1_2_7_n92, npu_inst_pe_1_2_7_n91,
         npu_inst_pe_1_2_7_n90, npu_inst_pe_1_2_7_n89, npu_inst_pe_1_2_7_n88,
         npu_inst_pe_1_2_7_n87, npu_inst_pe_1_2_7_n86, npu_inst_pe_1_2_7_n85,
         npu_inst_pe_1_2_7_n84, npu_inst_pe_1_2_7_n83, npu_inst_pe_1_2_7_n82,
         npu_inst_pe_1_2_7_n81, npu_inst_pe_1_2_7_n80, npu_inst_pe_1_2_7_n79,
         npu_inst_pe_1_2_7_n78, npu_inst_pe_1_2_7_n77, npu_inst_pe_1_2_7_n76,
         npu_inst_pe_1_2_7_n75, npu_inst_pe_1_2_7_n74, npu_inst_pe_1_2_7_n73,
         npu_inst_pe_1_2_7_n72, npu_inst_pe_1_2_7_n71, npu_inst_pe_1_2_7_n70,
         npu_inst_pe_1_2_7_n69, npu_inst_pe_1_2_7_n68, npu_inst_pe_1_2_7_n67,
         npu_inst_pe_1_2_7_n66, npu_inst_pe_1_2_7_n65, npu_inst_pe_1_2_7_n64,
         npu_inst_pe_1_2_7_n63, npu_inst_pe_1_2_7_n62, npu_inst_pe_1_2_7_n61,
         npu_inst_pe_1_2_7_n60, npu_inst_pe_1_2_7_n59, npu_inst_pe_1_2_7_n58,
         npu_inst_pe_1_2_7_n57, npu_inst_pe_1_2_7_n56, npu_inst_pe_1_2_7_n55,
         npu_inst_pe_1_2_7_n54, npu_inst_pe_1_2_7_n53, npu_inst_pe_1_2_7_n52,
         npu_inst_pe_1_2_7_n51, npu_inst_pe_1_2_7_n50, npu_inst_pe_1_2_7_n49,
         npu_inst_pe_1_2_7_n48, npu_inst_pe_1_2_7_n47, npu_inst_pe_1_2_7_n46,
         npu_inst_pe_1_2_7_n45, npu_inst_pe_1_2_7_n44, npu_inst_pe_1_2_7_n43,
         npu_inst_pe_1_2_7_n42, npu_inst_pe_1_2_7_n41, npu_inst_pe_1_2_7_n40,
         npu_inst_pe_1_2_7_n39, npu_inst_pe_1_2_7_n38, npu_inst_pe_1_2_7_n37,
         npu_inst_pe_1_2_7_n27, npu_inst_pe_1_2_7_n26,
         npu_inst_pe_1_2_7_net4039, npu_inst_pe_1_2_7_net4033,
         npu_inst_pe_1_2_7_N94, npu_inst_pe_1_2_7_N93, npu_inst_pe_1_2_7_N84,
         npu_inst_pe_1_2_7_N80, npu_inst_pe_1_2_7_N79, npu_inst_pe_1_2_7_N78,
         npu_inst_pe_1_2_7_N77, npu_inst_pe_1_2_7_N76, npu_inst_pe_1_2_7_N75,
         npu_inst_pe_1_2_7_N74, npu_inst_pe_1_2_7_N73, npu_inst_pe_1_2_7_N72,
         npu_inst_pe_1_2_7_N71, npu_inst_pe_1_2_7_N70, npu_inst_pe_1_2_7_N69,
         npu_inst_pe_1_2_7_N68, npu_inst_pe_1_2_7_N67, npu_inst_pe_1_2_7_N66,
         npu_inst_pe_1_2_7_N65, npu_inst_pe_1_2_7_int_q_acc_0_,
         npu_inst_pe_1_2_7_int_q_acc_1_, npu_inst_pe_1_2_7_int_q_acc_2_,
         npu_inst_pe_1_2_7_int_q_acc_3_, npu_inst_pe_1_2_7_int_q_acc_4_,
         npu_inst_pe_1_2_7_int_q_acc_5_, npu_inst_pe_1_2_7_int_q_acc_6_,
         npu_inst_pe_1_2_7_int_q_acc_7_, npu_inst_pe_1_2_7_int_data_0_,
         npu_inst_pe_1_2_7_int_data_1_, npu_inst_pe_1_2_7_int_q_weight_0_,
         npu_inst_pe_1_2_7_int_q_weight_1_,
         npu_inst_pe_1_2_7_int_q_reg_v_5__0_,
         npu_inst_pe_1_2_7_int_q_reg_v_5__1_,
         npu_inst_pe_1_2_7_int_q_reg_v_4__0_,
         npu_inst_pe_1_2_7_int_q_reg_v_4__1_,
         npu_inst_pe_1_2_7_int_q_reg_v_3__0_,
         npu_inst_pe_1_2_7_int_q_reg_v_3__1_,
         npu_inst_pe_1_2_7_int_q_reg_v_2__0_,
         npu_inst_pe_1_2_7_int_q_reg_v_2__1_,
         npu_inst_pe_1_2_7_int_q_reg_v_1__0_,
         npu_inst_pe_1_2_7_int_q_reg_v_1__1_,
         npu_inst_pe_1_2_7_int_q_reg_v_0__0_,
         npu_inst_pe_1_2_7_int_q_reg_v_0__1_,
         npu_inst_pe_1_2_7_int_q_reg_h_5__0_,
         npu_inst_pe_1_2_7_int_q_reg_h_5__1_,
         npu_inst_pe_1_2_7_int_q_reg_h_4__0_,
         npu_inst_pe_1_2_7_int_q_reg_h_4__1_,
         npu_inst_pe_1_2_7_int_q_reg_h_3__0_,
         npu_inst_pe_1_2_7_int_q_reg_h_3__1_,
         npu_inst_pe_1_2_7_int_q_reg_h_2__0_,
         npu_inst_pe_1_2_7_int_q_reg_h_2__1_,
         npu_inst_pe_1_2_7_int_q_reg_h_1__0_,
         npu_inst_pe_1_2_7_int_q_reg_h_1__1_,
         npu_inst_pe_1_2_7_int_q_reg_h_0__0_,
         npu_inst_pe_1_2_7_int_q_reg_h_0__1_, npu_inst_pe_1_3_0_n119,
         npu_inst_pe_1_3_0_n118, npu_inst_pe_1_3_0_n117,
         npu_inst_pe_1_3_0_n116, npu_inst_pe_1_3_0_n115,
         npu_inst_pe_1_3_0_n114, npu_inst_pe_1_3_0_n113,
         npu_inst_pe_1_3_0_n112, npu_inst_pe_1_3_0_n111,
         npu_inst_pe_1_3_0_n110, npu_inst_pe_1_3_0_n109,
         npu_inst_pe_1_3_0_n108, npu_inst_pe_1_3_0_n107,
         npu_inst_pe_1_3_0_n106, npu_inst_pe_1_3_0_n105,
         npu_inst_pe_1_3_0_n104, npu_inst_pe_1_3_0_n103,
         npu_inst_pe_1_3_0_n102, npu_inst_pe_1_3_0_n101,
         npu_inst_pe_1_3_0_n100, npu_inst_pe_1_3_0_n99, npu_inst_pe_1_3_0_n98,
         npu_inst_pe_1_3_0_n36, npu_inst_pe_1_3_0_n35, npu_inst_pe_1_3_0_n34,
         npu_inst_pe_1_3_0_n33, npu_inst_pe_1_3_0_n32, npu_inst_pe_1_3_0_n31,
         npu_inst_pe_1_3_0_n30, npu_inst_pe_1_3_0_n29, npu_inst_pe_1_3_0_n28,
         npu_inst_pe_1_3_0_n25, npu_inst_pe_1_3_0_n24, npu_inst_pe_1_3_0_n23,
         npu_inst_pe_1_3_0_n22, npu_inst_pe_1_3_0_n21, npu_inst_pe_1_3_0_n20,
         npu_inst_pe_1_3_0_n19, npu_inst_pe_1_3_0_n18, npu_inst_pe_1_3_0_n17,
         npu_inst_pe_1_3_0_n16, npu_inst_pe_1_3_0_n15, npu_inst_pe_1_3_0_n14,
         npu_inst_pe_1_3_0_n13, npu_inst_pe_1_3_0_n12, npu_inst_pe_1_3_0_n11,
         npu_inst_pe_1_3_0_n10, npu_inst_pe_1_3_0_n9, npu_inst_pe_1_3_0_n8,
         npu_inst_pe_1_3_0_n7, npu_inst_pe_1_3_0_n6, npu_inst_pe_1_3_0_n5,
         npu_inst_pe_1_3_0_n4, npu_inst_pe_1_3_0_n3, npu_inst_pe_1_3_0_n2,
         npu_inst_pe_1_3_0_n1, npu_inst_pe_1_3_0_sub_67_carry_7_,
         npu_inst_pe_1_3_0_sub_67_carry_6_, npu_inst_pe_1_3_0_sub_67_carry_5_,
         npu_inst_pe_1_3_0_sub_67_carry_4_, npu_inst_pe_1_3_0_sub_67_carry_3_,
         npu_inst_pe_1_3_0_sub_67_carry_2_, npu_inst_pe_1_3_0_sub_67_carry_1_,
         npu_inst_pe_1_3_0_add_69_carry_7_, npu_inst_pe_1_3_0_add_69_carry_6_,
         npu_inst_pe_1_3_0_add_69_carry_5_, npu_inst_pe_1_3_0_add_69_carry_4_,
         npu_inst_pe_1_3_0_add_69_carry_3_, npu_inst_pe_1_3_0_add_69_carry_2_,
         npu_inst_pe_1_3_0_add_69_carry_1_, npu_inst_pe_1_3_0_n97,
         npu_inst_pe_1_3_0_n96, npu_inst_pe_1_3_0_n95, npu_inst_pe_1_3_0_n94,
         npu_inst_pe_1_3_0_n93, npu_inst_pe_1_3_0_n92, npu_inst_pe_1_3_0_n91,
         npu_inst_pe_1_3_0_n90, npu_inst_pe_1_3_0_n89, npu_inst_pe_1_3_0_n88,
         npu_inst_pe_1_3_0_n87, npu_inst_pe_1_3_0_n86, npu_inst_pe_1_3_0_n85,
         npu_inst_pe_1_3_0_n84, npu_inst_pe_1_3_0_n83, npu_inst_pe_1_3_0_n82,
         npu_inst_pe_1_3_0_n81, npu_inst_pe_1_3_0_n80, npu_inst_pe_1_3_0_n79,
         npu_inst_pe_1_3_0_n78, npu_inst_pe_1_3_0_n77, npu_inst_pe_1_3_0_n76,
         npu_inst_pe_1_3_0_n75, npu_inst_pe_1_3_0_n74, npu_inst_pe_1_3_0_n73,
         npu_inst_pe_1_3_0_n72, npu_inst_pe_1_3_0_n71, npu_inst_pe_1_3_0_n70,
         npu_inst_pe_1_3_0_n69, npu_inst_pe_1_3_0_n68, npu_inst_pe_1_3_0_n67,
         npu_inst_pe_1_3_0_n66, npu_inst_pe_1_3_0_n65, npu_inst_pe_1_3_0_n64,
         npu_inst_pe_1_3_0_n63, npu_inst_pe_1_3_0_n62, npu_inst_pe_1_3_0_n61,
         npu_inst_pe_1_3_0_n60, npu_inst_pe_1_3_0_n59, npu_inst_pe_1_3_0_n58,
         npu_inst_pe_1_3_0_n57, npu_inst_pe_1_3_0_n56, npu_inst_pe_1_3_0_n55,
         npu_inst_pe_1_3_0_n54, npu_inst_pe_1_3_0_n53, npu_inst_pe_1_3_0_n52,
         npu_inst_pe_1_3_0_n51, npu_inst_pe_1_3_0_n50, npu_inst_pe_1_3_0_n49,
         npu_inst_pe_1_3_0_n48, npu_inst_pe_1_3_0_n47, npu_inst_pe_1_3_0_n46,
         npu_inst_pe_1_3_0_n45, npu_inst_pe_1_3_0_n44, npu_inst_pe_1_3_0_n43,
         npu_inst_pe_1_3_0_n42, npu_inst_pe_1_3_0_n41, npu_inst_pe_1_3_0_n40,
         npu_inst_pe_1_3_0_n39, npu_inst_pe_1_3_0_n38, npu_inst_pe_1_3_0_n37,
         npu_inst_pe_1_3_0_n27, npu_inst_pe_1_3_0_n26,
         npu_inst_pe_1_3_0_net4016, npu_inst_pe_1_3_0_net4010,
         npu_inst_pe_1_3_0_N94, npu_inst_pe_1_3_0_N93, npu_inst_pe_1_3_0_N84,
         npu_inst_pe_1_3_0_N80, npu_inst_pe_1_3_0_N79, npu_inst_pe_1_3_0_N78,
         npu_inst_pe_1_3_0_N77, npu_inst_pe_1_3_0_N76, npu_inst_pe_1_3_0_N75,
         npu_inst_pe_1_3_0_N74, npu_inst_pe_1_3_0_N73, npu_inst_pe_1_3_0_N72,
         npu_inst_pe_1_3_0_N71, npu_inst_pe_1_3_0_N70, npu_inst_pe_1_3_0_N69,
         npu_inst_pe_1_3_0_N68, npu_inst_pe_1_3_0_N67, npu_inst_pe_1_3_0_N66,
         npu_inst_pe_1_3_0_N65, npu_inst_pe_1_3_0_int_q_acc_0_,
         npu_inst_pe_1_3_0_int_q_acc_1_, npu_inst_pe_1_3_0_int_q_acc_2_,
         npu_inst_pe_1_3_0_int_q_acc_3_, npu_inst_pe_1_3_0_int_q_acc_4_,
         npu_inst_pe_1_3_0_int_q_acc_5_, npu_inst_pe_1_3_0_int_q_acc_6_,
         npu_inst_pe_1_3_0_int_q_acc_7_, npu_inst_pe_1_3_0_int_data_0_,
         npu_inst_pe_1_3_0_int_data_1_, npu_inst_pe_1_3_0_int_q_weight_0_,
         npu_inst_pe_1_3_0_int_q_weight_1_,
         npu_inst_pe_1_3_0_int_q_reg_v_5__0_,
         npu_inst_pe_1_3_0_int_q_reg_v_5__1_,
         npu_inst_pe_1_3_0_int_q_reg_v_4__0_,
         npu_inst_pe_1_3_0_int_q_reg_v_4__1_,
         npu_inst_pe_1_3_0_int_q_reg_v_3__0_,
         npu_inst_pe_1_3_0_int_q_reg_v_3__1_,
         npu_inst_pe_1_3_0_int_q_reg_v_2__0_,
         npu_inst_pe_1_3_0_int_q_reg_v_2__1_,
         npu_inst_pe_1_3_0_int_q_reg_v_1__0_,
         npu_inst_pe_1_3_0_int_q_reg_v_1__1_,
         npu_inst_pe_1_3_0_int_q_reg_v_0__0_,
         npu_inst_pe_1_3_0_int_q_reg_v_0__1_,
         npu_inst_pe_1_3_0_int_q_reg_h_5__0_,
         npu_inst_pe_1_3_0_int_q_reg_h_5__1_,
         npu_inst_pe_1_3_0_int_q_reg_h_4__0_,
         npu_inst_pe_1_3_0_int_q_reg_h_4__1_,
         npu_inst_pe_1_3_0_int_q_reg_h_3__0_,
         npu_inst_pe_1_3_0_int_q_reg_h_3__1_,
         npu_inst_pe_1_3_0_int_q_reg_h_2__0_,
         npu_inst_pe_1_3_0_int_q_reg_h_2__1_,
         npu_inst_pe_1_3_0_int_q_reg_h_1__0_,
         npu_inst_pe_1_3_0_int_q_reg_h_1__1_,
         npu_inst_pe_1_3_0_int_q_reg_h_0__0_,
         npu_inst_pe_1_3_0_int_q_reg_h_0__1_, npu_inst_pe_1_3_0_o_data_h_0_,
         npu_inst_pe_1_3_0_o_data_h_1_, npu_inst_pe_1_3_1_n119,
         npu_inst_pe_1_3_1_n118, npu_inst_pe_1_3_1_n117,
         npu_inst_pe_1_3_1_n116, npu_inst_pe_1_3_1_n115,
         npu_inst_pe_1_3_1_n114, npu_inst_pe_1_3_1_n113,
         npu_inst_pe_1_3_1_n112, npu_inst_pe_1_3_1_n111,
         npu_inst_pe_1_3_1_n110, npu_inst_pe_1_3_1_n109,
         npu_inst_pe_1_3_1_n108, npu_inst_pe_1_3_1_n107,
         npu_inst_pe_1_3_1_n106, npu_inst_pe_1_3_1_n105,
         npu_inst_pe_1_3_1_n104, npu_inst_pe_1_3_1_n103,
         npu_inst_pe_1_3_1_n102, npu_inst_pe_1_3_1_n101,
         npu_inst_pe_1_3_1_n100, npu_inst_pe_1_3_1_n99, npu_inst_pe_1_3_1_n98,
         npu_inst_pe_1_3_1_n36, npu_inst_pe_1_3_1_n35, npu_inst_pe_1_3_1_n34,
         npu_inst_pe_1_3_1_n33, npu_inst_pe_1_3_1_n32, npu_inst_pe_1_3_1_n31,
         npu_inst_pe_1_3_1_n30, npu_inst_pe_1_3_1_n29, npu_inst_pe_1_3_1_n28,
         npu_inst_pe_1_3_1_n25, npu_inst_pe_1_3_1_n24, npu_inst_pe_1_3_1_n23,
         npu_inst_pe_1_3_1_n22, npu_inst_pe_1_3_1_n21, npu_inst_pe_1_3_1_n20,
         npu_inst_pe_1_3_1_n19, npu_inst_pe_1_3_1_n18, npu_inst_pe_1_3_1_n17,
         npu_inst_pe_1_3_1_n16, npu_inst_pe_1_3_1_n15, npu_inst_pe_1_3_1_n14,
         npu_inst_pe_1_3_1_n13, npu_inst_pe_1_3_1_n12, npu_inst_pe_1_3_1_n11,
         npu_inst_pe_1_3_1_n10, npu_inst_pe_1_3_1_n9, npu_inst_pe_1_3_1_n8,
         npu_inst_pe_1_3_1_n7, npu_inst_pe_1_3_1_n6, npu_inst_pe_1_3_1_n5,
         npu_inst_pe_1_3_1_n4, npu_inst_pe_1_3_1_n3, npu_inst_pe_1_3_1_n2,
         npu_inst_pe_1_3_1_n1, npu_inst_pe_1_3_1_sub_67_carry_7_,
         npu_inst_pe_1_3_1_sub_67_carry_6_, npu_inst_pe_1_3_1_sub_67_carry_5_,
         npu_inst_pe_1_3_1_sub_67_carry_4_, npu_inst_pe_1_3_1_sub_67_carry_3_,
         npu_inst_pe_1_3_1_sub_67_carry_2_, npu_inst_pe_1_3_1_sub_67_carry_1_,
         npu_inst_pe_1_3_1_add_69_carry_7_, npu_inst_pe_1_3_1_add_69_carry_6_,
         npu_inst_pe_1_3_1_add_69_carry_5_, npu_inst_pe_1_3_1_add_69_carry_4_,
         npu_inst_pe_1_3_1_add_69_carry_3_, npu_inst_pe_1_3_1_add_69_carry_2_,
         npu_inst_pe_1_3_1_add_69_carry_1_, npu_inst_pe_1_3_1_n97,
         npu_inst_pe_1_3_1_n96, npu_inst_pe_1_3_1_n95, npu_inst_pe_1_3_1_n94,
         npu_inst_pe_1_3_1_n93, npu_inst_pe_1_3_1_n92, npu_inst_pe_1_3_1_n91,
         npu_inst_pe_1_3_1_n90, npu_inst_pe_1_3_1_n89, npu_inst_pe_1_3_1_n88,
         npu_inst_pe_1_3_1_n87, npu_inst_pe_1_3_1_n86, npu_inst_pe_1_3_1_n85,
         npu_inst_pe_1_3_1_n84, npu_inst_pe_1_3_1_n83, npu_inst_pe_1_3_1_n82,
         npu_inst_pe_1_3_1_n81, npu_inst_pe_1_3_1_n80, npu_inst_pe_1_3_1_n79,
         npu_inst_pe_1_3_1_n78, npu_inst_pe_1_3_1_n77, npu_inst_pe_1_3_1_n76,
         npu_inst_pe_1_3_1_n75, npu_inst_pe_1_3_1_n74, npu_inst_pe_1_3_1_n73,
         npu_inst_pe_1_3_1_n72, npu_inst_pe_1_3_1_n71, npu_inst_pe_1_3_1_n70,
         npu_inst_pe_1_3_1_n69, npu_inst_pe_1_3_1_n68, npu_inst_pe_1_3_1_n67,
         npu_inst_pe_1_3_1_n66, npu_inst_pe_1_3_1_n65, npu_inst_pe_1_3_1_n64,
         npu_inst_pe_1_3_1_n63, npu_inst_pe_1_3_1_n62, npu_inst_pe_1_3_1_n61,
         npu_inst_pe_1_3_1_n60, npu_inst_pe_1_3_1_n59, npu_inst_pe_1_3_1_n58,
         npu_inst_pe_1_3_1_n57, npu_inst_pe_1_3_1_n56, npu_inst_pe_1_3_1_n55,
         npu_inst_pe_1_3_1_n54, npu_inst_pe_1_3_1_n53, npu_inst_pe_1_3_1_n52,
         npu_inst_pe_1_3_1_n51, npu_inst_pe_1_3_1_n50, npu_inst_pe_1_3_1_n49,
         npu_inst_pe_1_3_1_n48, npu_inst_pe_1_3_1_n47, npu_inst_pe_1_3_1_n46,
         npu_inst_pe_1_3_1_n45, npu_inst_pe_1_3_1_n44, npu_inst_pe_1_3_1_n43,
         npu_inst_pe_1_3_1_n42, npu_inst_pe_1_3_1_n41, npu_inst_pe_1_3_1_n40,
         npu_inst_pe_1_3_1_n39, npu_inst_pe_1_3_1_n38, npu_inst_pe_1_3_1_n37,
         npu_inst_pe_1_3_1_n27, npu_inst_pe_1_3_1_n26,
         npu_inst_pe_1_3_1_net3993, npu_inst_pe_1_3_1_net3987,
         npu_inst_pe_1_3_1_N94, npu_inst_pe_1_3_1_N93, npu_inst_pe_1_3_1_N84,
         npu_inst_pe_1_3_1_N80, npu_inst_pe_1_3_1_N79, npu_inst_pe_1_3_1_N78,
         npu_inst_pe_1_3_1_N77, npu_inst_pe_1_3_1_N76, npu_inst_pe_1_3_1_N75,
         npu_inst_pe_1_3_1_N74, npu_inst_pe_1_3_1_N73, npu_inst_pe_1_3_1_N72,
         npu_inst_pe_1_3_1_N71, npu_inst_pe_1_3_1_N70, npu_inst_pe_1_3_1_N69,
         npu_inst_pe_1_3_1_N68, npu_inst_pe_1_3_1_N67, npu_inst_pe_1_3_1_N66,
         npu_inst_pe_1_3_1_N65, npu_inst_pe_1_3_1_int_q_acc_0_,
         npu_inst_pe_1_3_1_int_q_acc_1_, npu_inst_pe_1_3_1_int_q_acc_2_,
         npu_inst_pe_1_3_1_int_q_acc_3_, npu_inst_pe_1_3_1_int_q_acc_4_,
         npu_inst_pe_1_3_1_int_q_acc_5_, npu_inst_pe_1_3_1_int_q_acc_6_,
         npu_inst_pe_1_3_1_int_q_acc_7_, npu_inst_pe_1_3_1_int_data_0_,
         npu_inst_pe_1_3_1_int_data_1_, npu_inst_pe_1_3_1_int_q_weight_0_,
         npu_inst_pe_1_3_1_int_q_weight_1_,
         npu_inst_pe_1_3_1_int_q_reg_v_5__0_,
         npu_inst_pe_1_3_1_int_q_reg_v_5__1_,
         npu_inst_pe_1_3_1_int_q_reg_v_4__0_,
         npu_inst_pe_1_3_1_int_q_reg_v_4__1_,
         npu_inst_pe_1_3_1_int_q_reg_v_3__0_,
         npu_inst_pe_1_3_1_int_q_reg_v_3__1_,
         npu_inst_pe_1_3_1_int_q_reg_v_2__0_,
         npu_inst_pe_1_3_1_int_q_reg_v_2__1_,
         npu_inst_pe_1_3_1_int_q_reg_v_1__0_,
         npu_inst_pe_1_3_1_int_q_reg_v_1__1_,
         npu_inst_pe_1_3_1_int_q_reg_v_0__0_,
         npu_inst_pe_1_3_1_int_q_reg_v_0__1_,
         npu_inst_pe_1_3_1_int_q_reg_h_5__0_,
         npu_inst_pe_1_3_1_int_q_reg_h_5__1_,
         npu_inst_pe_1_3_1_int_q_reg_h_4__0_,
         npu_inst_pe_1_3_1_int_q_reg_h_4__1_,
         npu_inst_pe_1_3_1_int_q_reg_h_3__0_,
         npu_inst_pe_1_3_1_int_q_reg_h_3__1_,
         npu_inst_pe_1_3_1_int_q_reg_h_2__0_,
         npu_inst_pe_1_3_1_int_q_reg_h_2__1_,
         npu_inst_pe_1_3_1_int_q_reg_h_1__0_,
         npu_inst_pe_1_3_1_int_q_reg_h_1__1_,
         npu_inst_pe_1_3_1_int_q_reg_h_0__0_,
         npu_inst_pe_1_3_1_int_q_reg_h_0__1_, npu_inst_pe_1_3_2_n119,
         npu_inst_pe_1_3_2_n118, npu_inst_pe_1_3_2_n117,
         npu_inst_pe_1_3_2_n116, npu_inst_pe_1_3_2_n115,
         npu_inst_pe_1_3_2_n114, npu_inst_pe_1_3_2_n113,
         npu_inst_pe_1_3_2_n112, npu_inst_pe_1_3_2_n111,
         npu_inst_pe_1_3_2_n110, npu_inst_pe_1_3_2_n109,
         npu_inst_pe_1_3_2_n108, npu_inst_pe_1_3_2_n107,
         npu_inst_pe_1_3_2_n106, npu_inst_pe_1_3_2_n105,
         npu_inst_pe_1_3_2_n104, npu_inst_pe_1_3_2_n103,
         npu_inst_pe_1_3_2_n102, npu_inst_pe_1_3_2_n101,
         npu_inst_pe_1_3_2_n100, npu_inst_pe_1_3_2_n99, npu_inst_pe_1_3_2_n98,
         npu_inst_pe_1_3_2_n36, npu_inst_pe_1_3_2_n35, npu_inst_pe_1_3_2_n34,
         npu_inst_pe_1_3_2_n33, npu_inst_pe_1_3_2_n32, npu_inst_pe_1_3_2_n31,
         npu_inst_pe_1_3_2_n30, npu_inst_pe_1_3_2_n29, npu_inst_pe_1_3_2_n28,
         npu_inst_pe_1_3_2_n25, npu_inst_pe_1_3_2_n24, npu_inst_pe_1_3_2_n23,
         npu_inst_pe_1_3_2_n22, npu_inst_pe_1_3_2_n21, npu_inst_pe_1_3_2_n20,
         npu_inst_pe_1_3_2_n19, npu_inst_pe_1_3_2_n18, npu_inst_pe_1_3_2_n17,
         npu_inst_pe_1_3_2_n16, npu_inst_pe_1_3_2_n15, npu_inst_pe_1_3_2_n14,
         npu_inst_pe_1_3_2_n13, npu_inst_pe_1_3_2_n12, npu_inst_pe_1_3_2_n11,
         npu_inst_pe_1_3_2_n10, npu_inst_pe_1_3_2_n9, npu_inst_pe_1_3_2_n8,
         npu_inst_pe_1_3_2_n7, npu_inst_pe_1_3_2_n6, npu_inst_pe_1_3_2_n5,
         npu_inst_pe_1_3_2_n4, npu_inst_pe_1_3_2_n3, npu_inst_pe_1_3_2_n2,
         npu_inst_pe_1_3_2_n1, npu_inst_pe_1_3_2_sub_67_carry_7_,
         npu_inst_pe_1_3_2_sub_67_carry_6_, npu_inst_pe_1_3_2_sub_67_carry_5_,
         npu_inst_pe_1_3_2_sub_67_carry_4_, npu_inst_pe_1_3_2_sub_67_carry_3_,
         npu_inst_pe_1_3_2_sub_67_carry_2_, npu_inst_pe_1_3_2_sub_67_carry_1_,
         npu_inst_pe_1_3_2_add_69_carry_7_, npu_inst_pe_1_3_2_add_69_carry_6_,
         npu_inst_pe_1_3_2_add_69_carry_5_, npu_inst_pe_1_3_2_add_69_carry_4_,
         npu_inst_pe_1_3_2_add_69_carry_3_, npu_inst_pe_1_3_2_add_69_carry_2_,
         npu_inst_pe_1_3_2_add_69_carry_1_, npu_inst_pe_1_3_2_n97,
         npu_inst_pe_1_3_2_n96, npu_inst_pe_1_3_2_n95, npu_inst_pe_1_3_2_n94,
         npu_inst_pe_1_3_2_n93, npu_inst_pe_1_3_2_n92, npu_inst_pe_1_3_2_n91,
         npu_inst_pe_1_3_2_n90, npu_inst_pe_1_3_2_n89, npu_inst_pe_1_3_2_n88,
         npu_inst_pe_1_3_2_n87, npu_inst_pe_1_3_2_n86, npu_inst_pe_1_3_2_n85,
         npu_inst_pe_1_3_2_n84, npu_inst_pe_1_3_2_n83, npu_inst_pe_1_3_2_n82,
         npu_inst_pe_1_3_2_n81, npu_inst_pe_1_3_2_n80, npu_inst_pe_1_3_2_n79,
         npu_inst_pe_1_3_2_n78, npu_inst_pe_1_3_2_n77, npu_inst_pe_1_3_2_n76,
         npu_inst_pe_1_3_2_n75, npu_inst_pe_1_3_2_n74, npu_inst_pe_1_3_2_n73,
         npu_inst_pe_1_3_2_n72, npu_inst_pe_1_3_2_n71, npu_inst_pe_1_3_2_n70,
         npu_inst_pe_1_3_2_n69, npu_inst_pe_1_3_2_n68, npu_inst_pe_1_3_2_n67,
         npu_inst_pe_1_3_2_n66, npu_inst_pe_1_3_2_n65, npu_inst_pe_1_3_2_n64,
         npu_inst_pe_1_3_2_n63, npu_inst_pe_1_3_2_n62, npu_inst_pe_1_3_2_n61,
         npu_inst_pe_1_3_2_n60, npu_inst_pe_1_3_2_n59, npu_inst_pe_1_3_2_n58,
         npu_inst_pe_1_3_2_n57, npu_inst_pe_1_3_2_n56, npu_inst_pe_1_3_2_n55,
         npu_inst_pe_1_3_2_n54, npu_inst_pe_1_3_2_n53, npu_inst_pe_1_3_2_n52,
         npu_inst_pe_1_3_2_n51, npu_inst_pe_1_3_2_n50, npu_inst_pe_1_3_2_n49,
         npu_inst_pe_1_3_2_n48, npu_inst_pe_1_3_2_n47, npu_inst_pe_1_3_2_n46,
         npu_inst_pe_1_3_2_n45, npu_inst_pe_1_3_2_n44, npu_inst_pe_1_3_2_n43,
         npu_inst_pe_1_3_2_n42, npu_inst_pe_1_3_2_n41, npu_inst_pe_1_3_2_n40,
         npu_inst_pe_1_3_2_n39, npu_inst_pe_1_3_2_n38, npu_inst_pe_1_3_2_n37,
         npu_inst_pe_1_3_2_n27, npu_inst_pe_1_3_2_n26,
         npu_inst_pe_1_3_2_net3970, npu_inst_pe_1_3_2_net3964,
         npu_inst_pe_1_3_2_N94, npu_inst_pe_1_3_2_N93, npu_inst_pe_1_3_2_N84,
         npu_inst_pe_1_3_2_N80, npu_inst_pe_1_3_2_N79, npu_inst_pe_1_3_2_N78,
         npu_inst_pe_1_3_2_N77, npu_inst_pe_1_3_2_N76, npu_inst_pe_1_3_2_N75,
         npu_inst_pe_1_3_2_N74, npu_inst_pe_1_3_2_N73, npu_inst_pe_1_3_2_N72,
         npu_inst_pe_1_3_2_N71, npu_inst_pe_1_3_2_N70, npu_inst_pe_1_3_2_N69,
         npu_inst_pe_1_3_2_N68, npu_inst_pe_1_3_2_N67, npu_inst_pe_1_3_2_N66,
         npu_inst_pe_1_3_2_N65, npu_inst_pe_1_3_2_int_q_acc_0_,
         npu_inst_pe_1_3_2_int_q_acc_1_, npu_inst_pe_1_3_2_int_q_acc_2_,
         npu_inst_pe_1_3_2_int_q_acc_3_, npu_inst_pe_1_3_2_int_q_acc_4_,
         npu_inst_pe_1_3_2_int_q_acc_5_, npu_inst_pe_1_3_2_int_q_acc_6_,
         npu_inst_pe_1_3_2_int_q_acc_7_, npu_inst_pe_1_3_2_int_data_0_,
         npu_inst_pe_1_3_2_int_data_1_, npu_inst_pe_1_3_2_int_q_weight_0_,
         npu_inst_pe_1_3_2_int_q_weight_1_,
         npu_inst_pe_1_3_2_int_q_reg_v_5__0_,
         npu_inst_pe_1_3_2_int_q_reg_v_5__1_,
         npu_inst_pe_1_3_2_int_q_reg_v_4__0_,
         npu_inst_pe_1_3_2_int_q_reg_v_4__1_,
         npu_inst_pe_1_3_2_int_q_reg_v_3__0_,
         npu_inst_pe_1_3_2_int_q_reg_v_3__1_,
         npu_inst_pe_1_3_2_int_q_reg_v_2__0_,
         npu_inst_pe_1_3_2_int_q_reg_v_2__1_,
         npu_inst_pe_1_3_2_int_q_reg_v_1__0_,
         npu_inst_pe_1_3_2_int_q_reg_v_1__1_,
         npu_inst_pe_1_3_2_int_q_reg_v_0__0_,
         npu_inst_pe_1_3_2_int_q_reg_v_0__1_,
         npu_inst_pe_1_3_2_int_q_reg_h_5__0_,
         npu_inst_pe_1_3_2_int_q_reg_h_5__1_,
         npu_inst_pe_1_3_2_int_q_reg_h_4__0_,
         npu_inst_pe_1_3_2_int_q_reg_h_4__1_,
         npu_inst_pe_1_3_2_int_q_reg_h_3__0_,
         npu_inst_pe_1_3_2_int_q_reg_h_3__1_,
         npu_inst_pe_1_3_2_int_q_reg_h_2__0_,
         npu_inst_pe_1_3_2_int_q_reg_h_2__1_,
         npu_inst_pe_1_3_2_int_q_reg_h_1__0_,
         npu_inst_pe_1_3_2_int_q_reg_h_1__1_,
         npu_inst_pe_1_3_2_int_q_reg_h_0__0_,
         npu_inst_pe_1_3_2_int_q_reg_h_0__1_, npu_inst_pe_1_3_3_n119,
         npu_inst_pe_1_3_3_n118, npu_inst_pe_1_3_3_n117,
         npu_inst_pe_1_3_3_n116, npu_inst_pe_1_3_3_n115,
         npu_inst_pe_1_3_3_n114, npu_inst_pe_1_3_3_n113,
         npu_inst_pe_1_3_3_n112, npu_inst_pe_1_3_3_n111,
         npu_inst_pe_1_3_3_n110, npu_inst_pe_1_3_3_n109,
         npu_inst_pe_1_3_3_n108, npu_inst_pe_1_3_3_n107,
         npu_inst_pe_1_3_3_n106, npu_inst_pe_1_3_3_n105,
         npu_inst_pe_1_3_3_n104, npu_inst_pe_1_3_3_n103,
         npu_inst_pe_1_3_3_n102, npu_inst_pe_1_3_3_n101,
         npu_inst_pe_1_3_3_n100, npu_inst_pe_1_3_3_n99, npu_inst_pe_1_3_3_n98,
         npu_inst_pe_1_3_3_n36, npu_inst_pe_1_3_3_n35, npu_inst_pe_1_3_3_n34,
         npu_inst_pe_1_3_3_n33, npu_inst_pe_1_3_3_n32, npu_inst_pe_1_3_3_n31,
         npu_inst_pe_1_3_3_n30, npu_inst_pe_1_3_3_n29, npu_inst_pe_1_3_3_n28,
         npu_inst_pe_1_3_3_n25, npu_inst_pe_1_3_3_n24, npu_inst_pe_1_3_3_n23,
         npu_inst_pe_1_3_3_n22, npu_inst_pe_1_3_3_n21, npu_inst_pe_1_3_3_n20,
         npu_inst_pe_1_3_3_n19, npu_inst_pe_1_3_3_n18, npu_inst_pe_1_3_3_n17,
         npu_inst_pe_1_3_3_n16, npu_inst_pe_1_3_3_n15, npu_inst_pe_1_3_3_n14,
         npu_inst_pe_1_3_3_n13, npu_inst_pe_1_3_3_n12, npu_inst_pe_1_3_3_n11,
         npu_inst_pe_1_3_3_n10, npu_inst_pe_1_3_3_n9, npu_inst_pe_1_3_3_n8,
         npu_inst_pe_1_3_3_n7, npu_inst_pe_1_3_3_n6, npu_inst_pe_1_3_3_n5,
         npu_inst_pe_1_3_3_n4, npu_inst_pe_1_3_3_n3, npu_inst_pe_1_3_3_n2,
         npu_inst_pe_1_3_3_n1, npu_inst_pe_1_3_3_sub_67_carry_7_,
         npu_inst_pe_1_3_3_sub_67_carry_6_, npu_inst_pe_1_3_3_sub_67_carry_5_,
         npu_inst_pe_1_3_3_sub_67_carry_4_, npu_inst_pe_1_3_3_sub_67_carry_3_,
         npu_inst_pe_1_3_3_sub_67_carry_2_, npu_inst_pe_1_3_3_sub_67_carry_1_,
         npu_inst_pe_1_3_3_add_69_carry_7_, npu_inst_pe_1_3_3_add_69_carry_6_,
         npu_inst_pe_1_3_3_add_69_carry_5_, npu_inst_pe_1_3_3_add_69_carry_4_,
         npu_inst_pe_1_3_3_add_69_carry_3_, npu_inst_pe_1_3_3_add_69_carry_2_,
         npu_inst_pe_1_3_3_add_69_carry_1_, npu_inst_pe_1_3_3_n97,
         npu_inst_pe_1_3_3_n96, npu_inst_pe_1_3_3_n95, npu_inst_pe_1_3_3_n94,
         npu_inst_pe_1_3_3_n93, npu_inst_pe_1_3_3_n92, npu_inst_pe_1_3_3_n91,
         npu_inst_pe_1_3_3_n90, npu_inst_pe_1_3_3_n89, npu_inst_pe_1_3_3_n88,
         npu_inst_pe_1_3_3_n87, npu_inst_pe_1_3_3_n86, npu_inst_pe_1_3_3_n85,
         npu_inst_pe_1_3_3_n84, npu_inst_pe_1_3_3_n83, npu_inst_pe_1_3_3_n82,
         npu_inst_pe_1_3_3_n81, npu_inst_pe_1_3_3_n80, npu_inst_pe_1_3_3_n79,
         npu_inst_pe_1_3_3_n78, npu_inst_pe_1_3_3_n77, npu_inst_pe_1_3_3_n76,
         npu_inst_pe_1_3_3_n75, npu_inst_pe_1_3_3_n74, npu_inst_pe_1_3_3_n73,
         npu_inst_pe_1_3_3_n72, npu_inst_pe_1_3_3_n71, npu_inst_pe_1_3_3_n70,
         npu_inst_pe_1_3_3_n69, npu_inst_pe_1_3_3_n68, npu_inst_pe_1_3_3_n67,
         npu_inst_pe_1_3_3_n66, npu_inst_pe_1_3_3_n65, npu_inst_pe_1_3_3_n64,
         npu_inst_pe_1_3_3_n63, npu_inst_pe_1_3_3_n62, npu_inst_pe_1_3_3_n61,
         npu_inst_pe_1_3_3_n60, npu_inst_pe_1_3_3_n59, npu_inst_pe_1_3_3_n58,
         npu_inst_pe_1_3_3_n57, npu_inst_pe_1_3_3_n56, npu_inst_pe_1_3_3_n55,
         npu_inst_pe_1_3_3_n54, npu_inst_pe_1_3_3_n53, npu_inst_pe_1_3_3_n52,
         npu_inst_pe_1_3_3_n51, npu_inst_pe_1_3_3_n50, npu_inst_pe_1_3_3_n49,
         npu_inst_pe_1_3_3_n48, npu_inst_pe_1_3_3_n47, npu_inst_pe_1_3_3_n46,
         npu_inst_pe_1_3_3_n45, npu_inst_pe_1_3_3_n44, npu_inst_pe_1_3_3_n43,
         npu_inst_pe_1_3_3_n42, npu_inst_pe_1_3_3_n41, npu_inst_pe_1_3_3_n40,
         npu_inst_pe_1_3_3_n39, npu_inst_pe_1_3_3_n38, npu_inst_pe_1_3_3_n37,
         npu_inst_pe_1_3_3_n27, npu_inst_pe_1_3_3_n26,
         npu_inst_pe_1_3_3_net3947, npu_inst_pe_1_3_3_net3941,
         npu_inst_pe_1_3_3_N94, npu_inst_pe_1_3_3_N93, npu_inst_pe_1_3_3_N84,
         npu_inst_pe_1_3_3_N80, npu_inst_pe_1_3_3_N79, npu_inst_pe_1_3_3_N78,
         npu_inst_pe_1_3_3_N77, npu_inst_pe_1_3_3_N76, npu_inst_pe_1_3_3_N75,
         npu_inst_pe_1_3_3_N74, npu_inst_pe_1_3_3_N73, npu_inst_pe_1_3_3_N72,
         npu_inst_pe_1_3_3_N71, npu_inst_pe_1_3_3_N70, npu_inst_pe_1_3_3_N69,
         npu_inst_pe_1_3_3_N68, npu_inst_pe_1_3_3_N67, npu_inst_pe_1_3_3_N66,
         npu_inst_pe_1_3_3_N65, npu_inst_pe_1_3_3_int_q_acc_0_,
         npu_inst_pe_1_3_3_int_q_acc_1_, npu_inst_pe_1_3_3_int_q_acc_2_,
         npu_inst_pe_1_3_3_int_q_acc_3_, npu_inst_pe_1_3_3_int_q_acc_4_,
         npu_inst_pe_1_3_3_int_q_acc_5_, npu_inst_pe_1_3_3_int_q_acc_6_,
         npu_inst_pe_1_3_3_int_q_acc_7_, npu_inst_pe_1_3_3_int_data_0_,
         npu_inst_pe_1_3_3_int_data_1_, npu_inst_pe_1_3_3_int_q_weight_0_,
         npu_inst_pe_1_3_3_int_q_weight_1_,
         npu_inst_pe_1_3_3_int_q_reg_v_5__0_,
         npu_inst_pe_1_3_3_int_q_reg_v_5__1_,
         npu_inst_pe_1_3_3_int_q_reg_v_4__0_,
         npu_inst_pe_1_3_3_int_q_reg_v_4__1_,
         npu_inst_pe_1_3_3_int_q_reg_v_3__0_,
         npu_inst_pe_1_3_3_int_q_reg_v_3__1_,
         npu_inst_pe_1_3_3_int_q_reg_v_2__0_,
         npu_inst_pe_1_3_3_int_q_reg_v_2__1_,
         npu_inst_pe_1_3_3_int_q_reg_v_1__0_,
         npu_inst_pe_1_3_3_int_q_reg_v_1__1_,
         npu_inst_pe_1_3_3_int_q_reg_v_0__0_,
         npu_inst_pe_1_3_3_int_q_reg_v_0__1_,
         npu_inst_pe_1_3_3_int_q_reg_h_5__0_,
         npu_inst_pe_1_3_3_int_q_reg_h_5__1_,
         npu_inst_pe_1_3_3_int_q_reg_h_4__0_,
         npu_inst_pe_1_3_3_int_q_reg_h_4__1_,
         npu_inst_pe_1_3_3_int_q_reg_h_3__0_,
         npu_inst_pe_1_3_3_int_q_reg_h_3__1_,
         npu_inst_pe_1_3_3_int_q_reg_h_2__0_,
         npu_inst_pe_1_3_3_int_q_reg_h_2__1_,
         npu_inst_pe_1_3_3_int_q_reg_h_1__0_,
         npu_inst_pe_1_3_3_int_q_reg_h_1__1_,
         npu_inst_pe_1_3_3_int_q_reg_h_0__0_,
         npu_inst_pe_1_3_3_int_q_reg_h_0__1_, npu_inst_pe_1_3_4_n118,
         npu_inst_pe_1_3_4_n117, npu_inst_pe_1_3_4_n116,
         npu_inst_pe_1_3_4_n115, npu_inst_pe_1_3_4_n114,
         npu_inst_pe_1_3_4_n113, npu_inst_pe_1_3_4_n112,
         npu_inst_pe_1_3_4_n111, npu_inst_pe_1_3_4_n110,
         npu_inst_pe_1_3_4_n109, npu_inst_pe_1_3_4_n108,
         npu_inst_pe_1_3_4_n107, npu_inst_pe_1_3_4_n106,
         npu_inst_pe_1_3_4_n105, npu_inst_pe_1_3_4_n104,
         npu_inst_pe_1_3_4_n103, npu_inst_pe_1_3_4_n102,
         npu_inst_pe_1_3_4_n101, npu_inst_pe_1_3_4_n100, npu_inst_pe_1_3_4_n99,
         npu_inst_pe_1_3_4_n98, npu_inst_pe_1_3_4_n36, npu_inst_pe_1_3_4_n35,
         npu_inst_pe_1_3_4_n34, npu_inst_pe_1_3_4_n33, npu_inst_pe_1_3_4_n32,
         npu_inst_pe_1_3_4_n31, npu_inst_pe_1_3_4_n30, npu_inst_pe_1_3_4_n29,
         npu_inst_pe_1_3_4_n28, npu_inst_pe_1_3_4_n25, npu_inst_pe_1_3_4_n24,
         npu_inst_pe_1_3_4_n23, npu_inst_pe_1_3_4_n22, npu_inst_pe_1_3_4_n21,
         npu_inst_pe_1_3_4_n20, npu_inst_pe_1_3_4_n19, npu_inst_pe_1_3_4_n18,
         npu_inst_pe_1_3_4_n17, npu_inst_pe_1_3_4_n16, npu_inst_pe_1_3_4_n15,
         npu_inst_pe_1_3_4_n14, npu_inst_pe_1_3_4_n13, npu_inst_pe_1_3_4_n12,
         npu_inst_pe_1_3_4_n11, npu_inst_pe_1_3_4_n10, npu_inst_pe_1_3_4_n9,
         npu_inst_pe_1_3_4_n8, npu_inst_pe_1_3_4_n7, npu_inst_pe_1_3_4_n6,
         npu_inst_pe_1_3_4_n5, npu_inst_pe_1_3_4_n4, npu_inst_pe_1_3_4_n3,
         npu_inst_pe_1_3_4_n2, npu_inst_pe_1_3_4_n1,
         npu_inst_pe_1_3_4_sub_67_carry_7_, npu_inst_pe_1_3_4_sub_67_carry_6_,
         npu_inst_pe_1_3_4_sub_67_carry_5_, npu_inst_pe_1_3_4_sub_67_carry_4_,
         npu_inst_pe_1_3_4_sub_67_carry_3_, npu_inst_pe_1_3_4_sub_67_carry_2_,
         npu_inst_pe_1_3_4_sub_67_carry_1_, npu_inst_pe_1_3_4_add_69_carry_7_,
         npu_inst_pe_1_3_4_add_69_carry_6_, npu_inst_pe_1_3_4_add_69_carry_5_,
         npu_inst_pe_1_3_4_add_69_carry_4_, npu_inst_pe_1_3_4_add_69_carry_3_,
         npu_inst_pe_1_3_4_add_69_carry_2_, npu_inst_pe_1_3_4_add_69_carry_1_,
         npu_inst_pe_1_3_4_n97, npu_inst_pe_1_3_4_n96, npu_inst_pe_1_3_4_n95,
         npu_inst_pe_1_3_4_n94, npu_inst_pe_1_3_4_n93, npu_inst_pe_1_3_4_n92,
         npu_inst_pe_1_3_4_n91, npu_inst_pe_1_3_4_n90, npu_inst_pe_1_3_4_n89,
         npu_inst_pe_1_3_4_n88, npu_inst_pe_1_3_4_n87, npu_inst_pe_1_3_4_n86,
         npu_inst_pe_1_3_4_n85, npu_inst_pe_1_3_4_n84, npu_inst_pe_1_3_4_n83,
         npu_inst_pe_1_3_4_n82, npu_inst_pe_1_3_4_n81, npu_inst_pe_1_3_4_n80,
         npu_inst_pe_1_3_4_n79, npu_inst_pe_1_3_4_n78, npu_inst_pe_1_3_4_n77,
         npu_inst_pe_1_3_4_n76, npu_inst_pe_1_3_4_n75, npu_inst_pe_1_3_4_n74,
         npu_inst_pe_1_3_4_n73, npu_inst_pe_1_3_4_n72, npu_inst_pe_1_3_4_n71,
         npu_inst_pe_1_3_4_n70, npu_inst_pe_1_3_4_n69, npu_inst_pe_1_3_4_n68,
         npu_inst_pe_1_3_4_n67, npu_inst_pe_1_3_4_n66, npu_inst_pe_1_3_4_n65,
         npu_inst_pe_1_3_4_n64, npu_inst_pe_1_3_4_n63, npu_inst_pe_1_3_4_n62,
         npu_inst_pe_1_3_4_n61, npu_inst_pe_1_3_4_n60, npu_inst_pe_1_3_4_n59,
         npu_inst_pe_1_3_4_n58, npu_inst_pe_1_3_4_n57, npu_inst_pe_1_3_4_n56,
         npu_inst_pe_1_3_4_n55, npu_inst_pe_1_3_4_n54, npu_inst_pe_1_3_4_n53,
         npu_inst_pe_1_3_4_n52, npu_inst_pe_1_3_4_n51, npu_inst_pe_1_3_4_n50,
         npu_inst_pe_1_3_4_n49, npu_inst_pe_1_3_4_n48, npu_inst_pe_1_3_4_n47,
         npu_inst_pe_1_3_4_n46, npu_inst_pe_1_3_4_n45, npu_inst_pe_1_3_4_n44,
         npu_inst_pe_1_3_4_n43, npu_inst_pe_1_3_4_n42, npu_inst_pe_1_3_4_n41,
         npu_inst_pe_1_3_4_n40, npu_inst_pe_1_3_4_n39, npu_inst_pe_1_3_4_n38,
         npu_inst_pe_1_3_4_n37, npu_inst_pe_1_3_4_n27, npu_inst_pe_1_3_4_n26,
         npu_inst_pe_1_3_4_net3924, npu_inst_pe_1_3_4_net3918,
         npu_inst_pe_1_3_4_N94, npu_inst_pe_1_3_4_N93, npu_inst_pe_1_3_4_N84,
         npu_inst_pe_1_3_4_N80, npu_inst_pe_1_3_4_N79, npu_inst_pe_1_3_4_N78,
         npu_inst_pe_1_3_4_N77, npu_inst_pe_1_3_4_N76, npu_inst_pe_1_3_4_N75,
         npu_inst_pe_1_3_4_N74, npu_inst_pe_1_3_4_N73, npu_inst_pe_1_3_4_N72,
         npu_inst_pe_1_3_4_N71, npu_inst_pe_1_3_4_N70, npu_inst_pe_1_3_4_N69,
         npu_inst_pe_1_3_4_N68, npu_inst_pe_1_3_4_N67, npu_inst_pe_1_3_4_N66,
         npu_inst_pe_1_3_4_N65, npu_inst_pe_1_3_4_int_q_acc_0_,
         npu_inst_pe_1_3_4_int_q_acc_1_, npu_inst_pe_1_3_4_int_q_acc_2_,
         npu_inst_pe_1_3_4_int_q_acc_3_, npu_inst_pe_1_3_4_int_q_acc_4_,
         npu_inst_pe_1_3_4_int_q_acc_5_, npu_inst_pe_1_3_4_int_q_acc_6_,
         npu_inst_pe_1_3_4_int_q_acc_7_, npu_inst_pe_1_3_4_int_data_0_,
         npu_inst_pe_1_3_4_int_data_1_, npu_inst_pe_1_3_4_int_q_weight_0_,
         npu_inst_pe_1_3_4_int_q_weight_1_,
         npu_inst_pe_1_3_4_int_q_reg_v_5__0_,
         npu_inst_pe_1_3_4_int_q_reg_v_5__1_,
         npu_inst_pe_1_3_4_int_q_reg_v_4__0_,
         npu_inst_pe_1_3_4_int_q_reg_v_4__1_,
         npu_inst_pe_1_3_4_int_q_reg_v_3__0_,
         npu_inst_pe_1_3_4_int_q_reg_v_3__1_,
         npu_inst_pe_1_3_4_int_q_reg_v_2__0_,
         npu_inst_pe_1_3_4_int_q_reg_v_2__1_,
         npu_inst_pe_1_3_4_int_q_reg_v_1__0_,
         npu_inst_pe_1_3_4_int_q_reg_v_1__1_,
         npu_inst_pe_1_3_4_int_q_reg_v_0__0_,
         npu_inst_pe_1_3_4_int_q_reg_v_0__1_,
         npu_inst_pe_1_3_4_int_q_reg_h_5__0_,
         npu_inst_pe_1_3_4_int_q_reg_h_5__1_,
         npu_inst_pe_1_3_4_int_q_reg_h_4__0_,
         npu_inst_pe_1_3_4_int_q_reg_h_4__1_,
         npu_inst_pe_1_3_4_int_q_reg_h_3__0_,
         npu_inst_pe_1_3_4_int_q_reg_h_3__1_,
         npu_inst_pe_1_3_4_int_q_reg_h_2__0_,
         npu_inst_pe_1_3_4_int_q_reg_h_2__1_,
         npu_inst_pe_1_3_4_int_q_reg_h_1__0_,
         npu_inst_pe_1_3_4_int_q_reg_h_1__1_,
         npu_inst_pe_1_3_4_int_q_reg_h_0__0_,
         npu_inst_pe_1_3_4_int_q_reg_h_0__1_, npu_inst_pe_1_3_5_n119,
         npu_inst_pe_1_3_5_n118, npu_inst_pe_1_3_5_n117,
         npu_inst_pe_1_3_5_n116, npu_inst_pe_1_3_5_n115,
         npu_inst_pe_1_3_5_n114, npu_inst_pe_1_3_5_n113,
         npu_inst_pe_1_3_5_n112, npu_inst_pe_1_3_5_n111,
         npu_inst_pe_1_3_5_n110, npu_inst_pe_1_3_5_n109,
         npu_inst_pe_1_3_5_n108, npu_inst_pe_1_3_5_n107,
         npu_inst_pe_1_3_5_n106, npu_inst_pe_1_3_5_n105,
         npu_inst_pe_1_3_5_n104, npu_inst_pe_1_3_5_n103,
         npu_inst_pe_1_3_5_n102, npu_inst_pe_1_3_5_n101,
         npu_inst_pe_1_3_5_n100, npu_inst_pe_1_3_5_n99, npu_inst_pe_1_3_5_n98,
         npu_inst_pe_1_3_5_n36, npu_inst_pe_1_3_5_n35, npu_inst_pe_1_3_5_n34,
         npu_inst_pe_1_3_5_n33, npu_inst_pe_1_3_5_n32, npu_inst_pe_1_3_5_n31,
         npu_inst_pe_1_3_5_n30, npu_inst_pe_1_3_5_n29, npu_inst_pe_1_3_5_n28,
         npu_inst_pe_1_3_5_n25, npu_inst_pe_1_3_5_n24, npu_inst_pe_1_3_5_n23,
         npu_inst_pe_1_3_5_n22, npu_inst_pe_1_3_5_n21, npu_inst_pe_1_3_5_n20,
         npu_inst_pe_1_3_5_n19, npu_inst_pe_1_3_5_n18, npu_inst_pe_1_3_5_n17,
         npu_inst_pe_1_3_5_n16, npu_inst_pe_1_3_5_n15, npu_inst_pe_1_3_5_n14,
         npu_inst_pe_1_3_5_n13, npu_inst_pe_1_3_5_n12, npu_inst_pe_1_3_5_n11,
         npu_inst_pe_1_3_5_n10, npu_inst_pe_1_3_5_n9, npu_inst_pe_1_3_5_n8,
         npu_inst_pe_1_3_5_n7, npu_inst_pe_1_3_5_n6, npu_inst_pe_1_3_5_n5,
         npu_inst_pe_1_3_5_n4, npu_inst_pe_1_3_5_n3, npu_inst_pe_1_3_5_n2,
         npu_inst_pe_1_3_5_n1, npu_inst_pe_1_3_5_sub_67_carry_7_,
         npu_inst_pe_1_3_5_sub_67_carry_6_, npu_inst_pe_1_3_5_sub_67_carry_5_,
         npu_inst_pe_1_3_5_sub_67_carry_4_, npu_inst_pe_1_3_5_sub_67_carry_3_,
         npu_inst_pe_1_3_5_sub_67_carry_2_, npu_inst_pe_1_3_5_sub_67_carry_1_,
         npu_inst_pe_1_3_5_add_69_carry_7_, npu_inst_pe_1_3_5_add_69_carry_6_,
         npu_inst_pe_1_3_5_add_69_carry_5_, npu_inst_pe_1_3_5_add_69_carry_4_,
         npu_inst_pe_1_3_5_add_69_carry_3_, npu_inst_pe_1_3_5_add_69_carry_2_,
         npu_inst_pe_1_3_5_add_69_carry_1_, npu_inst_pe_1_3_5_n97,
         npu_inst_pe_1_3_5_n96, npu_inst_pe_1_3_5_n95, npu_inst_pe_1_3_5_n94,
         npu_inst_pe_1_3_5_n93, npu_inst_pe_1_3_5_n92, npu_inst_pe_1_3_5_n91,
         npu_inst_pe_1_3_5_n90, npu_inst_pe_1_3_5_n89, npu_inst_pe_1_3_5_n88,
         npu_inst_pe_1_3_5_n87, npu_inst_pe_1_3_5_n86, npu_inst_pe_1_3_5_n85,
         npu_inst_pe_1_3_5_n84, npu_inst_pe_1_3_5_n83, npu_inst_pe_1_3_5_n82,
         npu_inst_pe_1_3_5_n81, npu_inst_pe_1_3_5_n80, npu_inst_pe_1_3_5_n79,
         npu_inst_pe_1_3_5_n78, npu_inst_pe_1_3_5_n77, npu_inst_pe_1_3_5_n76,
         npu_inst_pe_1_3_5_n75, npu_inst_pe_1_3_5_n74, npu_inst_pe_1_3_5_n73,
         npu_inst_pe_1_3_5_n72, npu_inst_pe_1_3_5_n71, npu_inst_pe_1_3_5_n70,
         npu_inst_pe_1_3_5_n69, npu_inst_pe_1_3_5_n68, npu_inst_pe_1_3_5_n67,
         npu_inst_pe_1_3_5_n66, npu_inst_pe_1_3_5_n65, npu_inst_pe_1_3_5_n64,
         npu_inst_pe_1_3_5_n63, npu_inst_pe_1_3_5_n62, npu_inst_pe_1_3_5_n61,
         npu_inst_pe_1_3_5_n60, npu_inst_pe_1_3_5_n59, npu_inst_pe_1_3_5_n58,
         npu_inst_pe_1_3_5_n57, npu_inst_pe_1_3_5_n56, npu_inst_pe_1_3_5_n55,
         npu_inst_pe_1_3_5_n54, npu_inst_pe_1_3_5_n53, npu_inst_pe_1_3_5_n52,
         npu_inst_pe_1_3_5_n51, npu_inst_pe_1_3_5_n50, npu_inst_pe_1_3_5_n49,
         npu_inst_pe_1_3_5_n48, npu_inst_pe_1_3_5_n47, npu_inst_pe_1_3_5_n46,
         npu_inst_pe_1_3_5_n45, npu_inst_pe_1_3_5_n44, npu_inst_pe_1_3_5_n43,
         npu_inst_pe_1_3_5_n42, npu_inst_pe_1_3_5_n41, npu_inst_pe_1_3_5_n40,
         npu_inst_pe_1_3_5_n39, npu_inst_pe_1_3_5_n38, npu_inst_pe_1_3_5_n37,
         npu_inst_pe_1_3_5_n27, npu_inst_pe_1_3_5_n26,
         npu_inst_pe_1_3_5_net3901, npu_inst_pe_1_3_5_net3895,
         npu_inst_pe_1_3_5_N94, npu_inst_pe_1_3_5_N93, npu_inst_pe_1_3_5_N84,
         npu_inst_pe_1_3_5_N80, npu_inst_pe_1_3_5_N79, npu_inst_pe_1_3_5_N78,
         npu_inst_pe_1_3_5_N77, npu_inst_pe_1_3_5_N76, npu_inst_pe_1_3_5_N75,
         npu_inst_pe_1_3_5_N74, npu_inst_pe_1_3_5_N73, npu_inst_pe_1_3_5_N72,
         npu_inst_pe_1_3_5_N71, npu_inst_pe_1_3_5_N70, npu_inst_pe_1_3_5_N69,
         npu_inst_pe_1_3_5_N68, npu_inst_pe_1_3_5_N67, npu_inst_pe_1_3_5_N66,
         npu_inst_pe_1_3_5_N65, npu_inst_pe_1_3_5_int_q_acc_0_,
         npu_inst_pe_1_3_5_int_q_acc_1_, npu_inst_pe_1_3_5_int_q_acc_2_,
         npu_inst_pe_1_3_5_int_q_acc_3_, npu_inst_pe_1_3_5_int_q_acc_4_,
         npu_inst_pe_1_3_5_int_q_acc_5_, npu_inst_pe_1_3_5_int_q_acc_6_,
         npu_inst_pe_1_3_5_int_q_acc_7_, npu_inst_pe_1_3_5_int_data_0_,
         npu_inst_pe_1_3_5_int_data_1_, npu_inst_pe_1_3_5_int_q_weight_0_,
         npu_inst_pe_1_3_5_int_q_weight_1_,
         npu_inst_pe_1_3_5_int_q_reg_v_5__0_,
         npu_inst_pe_1_3_5_int_q_reg_v_5__1_,
         npu_inst_pe_1_3_5_int_q_reg_v_4__0_,
         npu_inst_pe_1_3_5_int_q_reg_v_4__1_,
         npu_inst_pe_1_3_5_int_q_reg_v_3__0_,
         npu_inst_pe_1_3_5_int_q_reg_v_3__1_,
         npu_inst_pe_1_3_5_int_q_reg_v_2__0_,
         npu_inst_pe_1_3_5_int_q_reg_v_2__1_,
         npu_inst_pe_1_3_5_int_q_reg_v_1__0_,
         npu_inst_pe_1_3_5_int_q_reg_v_1__1_,
         npu_inst_pe_1_3_5_int_q_reg_v_0__0_,
         npu_inst_pe_1_3_5_int_q_reg_v_0__1_,
         npu_inst_pe_1_3_5_int_q_reg_h_5__0_,
         npu_inst_pe_1_3_5_int_q_reg_h_5__1_,
         npu_inst_pe_1_3_5_int_q_reg_h_4__0_,
         npu_inst_pe_1_3_5_int_q_reg_h_4__1_,
         npu_inst_pe_1_3_5_int_q_reg_h_3__0_,
         npu_inst_pe_1_3_5_int_q_reg_h_3__1_,
         npu_inst_pe_1_3_5_int_q_reg_h_2__0_,
         npu_inst_pe_1_3_5_int_q_reg_h_2__1_,
         npu_inst_pe_1_3_5_int_q_reg_h_1__0_,
         npu_inst_pe_1_3_5_int_q_reg_h_1__1_,
         npu_inst_pe_1_3_5_int_q_reg_h_0__0_,
         npu_inst_pe_1_3_5_int_q_reg_h_0__1_, npu_inst_pe_1_3_6_n119,
         npu_inst_pe_1_3_6_n118, npu_inst_pe_1_3_6_n117,
         npu_inst_pe_1_3_6_n116, npu_inst_pe_1_3_6_n115,
         npu_inst_pe_1_3_6_n114, npu_inst_pe_1_3_6_n113,
         npu_inst_pe_1_3_6_n112, npu_inst_pe_1_3_6_n111,
         npu_inst_pe_1_3_6_n110, npu_inst_pe_1_3_6_n109,
         npu_inst_pe_1_3_6_n108, npu_inst_pe_1_3_6_n107,
         npu_inst_pe_1_3_6_n106, npu_inst_pe_1_3_6_n105,
         npu_inst_pe_1_3_6_n104, npu_inst_pe_1_3_6_n103,
         npu_inst_pe_1_3_6_n102, npu_inst_pe_1_3_6_n101,
         npu_inst_pe_1_3_6_n100, npu_inst_pe_1_3_6_n99, npu_inst_pe_1_3_6_n98,
         npu_inst_pe_1_3_6_n36, npu_inst_pe_1_3_6_n35, npu_inst_pe_1_3_6_n34,
         npu_inst_pe_1_3_6_n33, npu_inst_pe_1_3_6_n32, npu_inst_pe_1_3_6_n31,
         npu_inst_pe_1_3_6_n30, npu_inst_pe_1_3_6_n29, npu_inst_pe_1_3_6_n28,
         npu_inst_pe_1_3_6_n25, npu_inst_pe_1_3_6_n24, npu_inst_pe_1_3_6_n23,
         npu_inst_pe_1_3_6_n22, npu_inst_pe_1_3_6_n21, npu_inst_pe_1_3_6_n20,
         npu_inst_pe_1_3_6_n19, npu_inst_pe_1_3_6_n18, npu_inst_pe_1_3_6_n17,
         npu_inst_pe_1_3_6_n16, npu_inst_pe_1_3_6_n15, npu_inst_pe_1_3_6_n14,
         npu_inst_pe_1_3_6_n13, npu_inst_pe_1_3_6_n12, npu_inst_pe_1_3_6_n11,
         npu_inst_pe_1_3_6_n10, npu_inst_pe_1_3_6_n9, npu_inst_pe_1_3_6_n8,
         npu_inst_pe_1_3_6_n7, npu_inst_pe_1_3_6_n6, npu_inst_pe_1_3_6_n5,
         npu_inst_pe_1_3_6_n4, npu_inst_pe_1_3_6_n3, npu_inst_pe_1_3_6_n2,
         npu_inst_pe_1_3_6_n1, npu_inst_pe_1_3_6_sub_67_carry_7_,
         npu_inst_pe_1_3_6_sub_67_carry_6_, npu_inst_pe_1_3_6_sub_67_carry_5_,
         npu_inst_pe_1_3_6_sub_67_carry_4_, npu_inst_pe_1_3_6_sub_67_carry_3_,
         npu_inst_pe_1_3_6_sub_67_carry_2_, npu_inst_pe_1_3_6_sub_67_carry_1_,
         npu_inst_pe_1_3_6_add_69_carry_7_, npu_inst_pe_1_3_6_add_69_carry_6_,
         npu_inst_pe_1_3_6_add_69_carry_5_, npu_inst_pe_1_3_6_add_69_carry_4_,
         npu_inst_pe_1_3_6_add_69_carry_3_, npu_inst_pe_1_3_6_add_69_carry_2_,
         npu_inst_pe_1_3_6_add_69_carry_1_, npu_inst_pe_1_3_6_n97,
         npu_inst_pe_1_3_6_n96, npu_inst_pe_1_3_6_n95, npu_inst_pe_1_3_6_n94,
         npu_inst_pe_1_3_6_n93, npu_inst_pe_1_3_6_n92, npu_inst_pe_1_3_6_n91,
         npu_inst_pe_1_3_6_n90, npu_inst_pe_1_3_6_n89, npu_inst_pe_1_3_6_n88,
         npu_inst_pe_1_3_6_n87, npu_inst_pe_1_3_6_n86, npu_inst_pe_1_3_6_n85,
         npu_inst_pe_1_3_6_n84, npu_inst_pe_1_3_6_n83, npu_inst_pe_1_3_6_n82,
         npu_inst_pe_1_3_6_n81, npu_inst_pe_1_3_6_n80, npu_inst_pe_1_3_6_n79,
         npu_inst_pe_1_3_6_n78, npu_inst_pe_1_3_6_n77, npu_inst_pe_1_3_6_n76,
         npu_inst_pe_1_3_6_n75, npu_inst_pe_1_3_6_n74, npu_inst_pe_1_3_6_n73,
         npu_inst_pe_1_3_6_n72, npu_inst_pe_1_3_6_n71, npu_inst_pe_1_3_6_n70,
         npu_inst_pe_1_3_6_n69, npu_inst_pe_1_3_6_n68, npu_inst_pe_1_3_6_n67,
         npu_inst_pe_1_3_6_n66, npu_inst_pe_1_3_6_n65, npu_inst_pe_1_3_6_n64,
         npu_inst_pe_1_3_6_n63, npu_inst_pe_1_3_6_n62, npu_inst_pe_1_3_6_n61,
         npu_inst_pe_1_3_6_n60, npu_inst_pe_1_3_6_n59, npu_inst_pe_1_3_6_n58,
         npu_inst_pe_1_3_6_n57, npu_inst_pe_1_3_6_n56, npu_inst_pe_1_3_6_n55,
         npu_inst_pe_1_3_6_n54, npu_inst_pe_1_3_6_n53, npu_inst_pe_1_3_6_n52,
         npu_inst_pe_1_3_6_n51, npu_inst_pe_1_3_6_n50, npu_inst_pe_1_3_6_n49,
         npu_inst_pe_1_3_6_n48, npu_inst_pe_1_3_6_n47, npu_inst_pe_1_3_6_n46,
         npu_inst_pe_1_3_6_n45, npu_inst_pe_1_3_6_n44, npu_inst_pe_1_3_6_n43,
         npu_inst_pe_1_3_6_n42, npu_inst_pe_1_3_6_n41, npu_inst_pe_1_3_6_n40,
         npu_inst_pe_1_3_6_n39, npu_inst_pe_1_3_6_n38, npu_inst_pe_1_3_6_n37,
         npu_inst_pe_1_3_6_n27, npu_inst_pe_1_3_6_n26,
         npu_inst_pe_1_3_6_net3878, npu_inst_pe_1_3_6_net3872,
         npu_inst_pe_1_3_6_N94, npu_inst_pe_1_3_6_N93, npu_inst_pe_1_3_6_N84,
         npu_inst_pe_1_3_6_N80, npu_inst_pe_1_3_6_N79, npu_inst_pe_1_3_6_N78,
         npu_inst_pe_1_3_6_N77, npu_inst_pe_1_3_6_N76, npu_inst_pe_1_3_6_N75,
         npu_inst_pe_1_3_6_N74, npu_inst_pe_1_3_6_N73, npu_inst_pe_1_3_6_N72,
         npu_inst_pe_1_3_6_N71, npu_inst_pe_1_3_6_N70, npu_inst_pe_1_3_6_N69,
         npu_inst_pe_1_3_6_N68, npu_inst_pe_1_3_6_N67, npu_inst_pe_1_3_6_N66,
         npu_inst_pe_1_3_6_N65, npu_inst_pe_1_3_6_int_q_acc_0_,
         npu_inst_pe_1_3_6_int_q_acc_1_, npu_inst_pe_1_3_6_int_q_acc_2_,
         npu_inst_pe_1_3_6_int_q_acc_3_, npu_inst_pe_1_3_6_int_q_acc_4_,
         npu_inst_pe_1_3_6_int_q_acc_5_, npu_inst_pe_1_3_6_int_q_acc_6_,
         npu_inst_pe_1_3_6_int_q_acc_7_, npu_inst_pe_1_3_6_int_data_0_,
         npu_inst_pe_1_3_6_int_data_1_, npu_inst_pe_1_3_6_int_q_weight_0_,
         npu_inst_pe_1_3_6_int_q_weight_1_,
         npu_inst_pe_1_3_6_int_q_reg_v_5__0_,
         npu_inst_pe_1_3_6_int_q_reg_v_5__1_,
         npu_inst_pe_1_3_6_int_q_reg_v_4__0_,
         npu_inst_pe_1_3_6_int_q_reg_v_4__1_,
         npu_inst_pe_1_3_6_int_q_reg_v_3__0_,
         npu_inst_pe_1_3_6_int_q_reg_v_3__1_,
         npu_inst_pe_1_3_6_int_q_reg_v_2__0_,
         npu_inst_pe_1_3_6_int_q_reg_v_2__1_,
         npu_inst_pe_1_3_6_int_q_reg_v_1__0_,
         npu_inst_pe_1_3_6_int_q_reg_v_1__1_,
         npu_inst_pe_1_3_6_int_q_reg_v_0__0_,
         npu_inst_pe_1_3_6_int_q_reg_v_0__1_,
         npu_inst_pe_1_3_6_int_q_reg_h_5__0_,
         npu_inst_pe_1_3_6_int_q_reg_h_5__1_,
         npu_inst_pe_1_3_6_int_q_reg_h_4__0_,
         npu_inst_pe_1_3_6_int_q_reg_h_4__1_,
         npu_inst_pe_1_3_6_int_q_reg_h_3__0_,
         npu_inst_pe_1_3_6_int_q_reg_h_3__1_,
         npu_inst_pe_1_3_6_int_q_reg_h_2__0_,
         npu_inst_pe_1_3_6_int_q_reg_h_2__1_,
         npu_inst_pe_1_3_6_int_q_reg_h_1__0_,
         npu_inst_pe_1_3_6_int_q_reg_h_1__1_,
         npu_inst_pe_1_3_6_int_q_reg_h_0__0_,
         npu_inst_pe_1_3_6_int_q_reg_h_0__1_, npu_inst_pe_1_3_7_n119,
         npu_inst_pe_1_3_7_n118, npu_inst_pe_1_3_7_n117,
         npu_inst_pe_1_3_7_n116, npu_inst_pe_1_3_7_n115,
         npu_inst_pe_1_3_7_n114, npu_inst_pe_1_3_7_n113,
         npu_inst_pe_1_3_7_n112, npu_inst_pe_1_3_7_n111,
         npu_inst_pe_1_3_7_n110, npu_inst_pe_1_3_7_n109,
         npu_inst_pe_1_3_7_n108, npu_inst_pe_1_3_7_n107,
         npu_inst_pe_1_3_7_n106, npu_inst_pe_1_3_7_n105,
         npu_inst_pe_1_3_7_n104, npu_inst_pe_1_3_7_n103,
         npu_inst_pe_1_3_7_n102, npu_inst_pe_1_3_7_n101,
         npu_inst_pe_1_3_7_n100, npu_inst_pe_1_3_7_n99, npu_inst_pe_1_3_7_n98,
         npu_inst_pe_1_3_7_n36, npu_inst_pe_1_3_7_n35, npu_inst_pe_1_3_7_n34,
         npu_inst_pe_1_3_7_n33, npu_inst_pe_1_3_7_n32, npu_inst_pe_1_3_7_n31,
         npu_inst_pe_1_3_7_n30, npu_inst_pe_1_3_7_n29, npu_inst_pe_1_3_7_n28,
         npu_inst_pe_1_3_7_n25, npu_inst_pe_1_3_7_n24, npu_inst_pe_1_3_7_n23,
         npu_inst_pe_1_3_7_n22, npu_inst_pe_1_3_7_n21, npu_inst_pe_1_3_7_n20,
         npu_inst_pe_1_3_7_n19, npu_inst_pe_1_3_7_n18, npu_inst_pe_1_3_7_n17,
         npu_inst_pe_1_3_7_n16, npu_inst_pe_1_3_7_n15, npu_inst_pe_1_3_7_n14,
         npu_inst_pe_1_3_7_n13, npu_inst_pe_1_3_7_n12, npu_inst_pe_1_3_7_n11,
         npu_inst_pe_1_3_7_n10, npu_inst_pe_1_3_7_n9, npu_inst_pe_1_3_7_n8,
         npu_inst_pe_1_3_7_n7, npu_inst_pe_1_3_7_n6, npu_inst_pe_1_3_7_n5,
         npu_inst_pe_1_3_7_n4, npu_inst_pe_1_3_7_n3, npu_inst_pe_1_3_7_n2,
         npu_inst_pe_1_3_7_n1, npu_inst_pe_1_3_7_sub_67_carry_7_,
         npu_inst_pe_1_3_7_sub_67_carry_6_, npu_inst_pe_1_3_7_sub_67_carry_5_,
         npu_inst_pe_1_3_7_sub_67_carry_4_, npu_inst_pe_1_3_7_sub_67_carry_3_,
         npu_inst_pe_1_3_7_sub_67_carry_2_, npu_inst_pe_1_3_7_sub_67_carry_1_,
         npu_inst_pe_1_3_7_add_69_carry_7_, npu_inst_pe_1_3_7_add_69_carry_6_,
         npu_inst_pe_1_3_7_add_69_carry_5_, npu_inst_pe_1_3_7_add_69_carry_4_,
         npu_inst_pe_1_3_7_add_69_carry_3_, npu_inst_pe_1_3_7_add_69_carry_2_,
         npu_inst_pe_1_3_7_add_69_carry_1_, npu_inst_pe_1_3_7_n97,
         npu_inst_pe_1_3_7_n96, npu_inst_pe_1_3_7_n95, npu_inst_pe_1_3_7_n94,
         npu_inst_pe_1_3_7_n93, npu_inst_pe_1_3_7_n92, npu_inst_pe_1_3_7_n91,
         npu_inst_pe_1_3_7_n90, npu_inst_pe_1_3_7_n89, npu_inst_pe_1_3_7_n88,
         npu_inst_pe_1_3_7_n87, npu_inst_pe_1_3_7_n86, npu_inst_pe_1_3_7_n85,
         npu_inst_pe_1_3_7_n84, npu_inst_pe_1_3_7_n83, npu_inst_pe_1_3_7_n82,
         npu_inst_pe_1_3_7_n81, npu_inst_pe_1_3_7_n80, npu_inst_pe_1_3_7_n79,
         npu_inst_pe_1_3_7_n78, npu_inst_pe_1_3_7_n77, npu_inst_pe_1_3_7_n76,
         npu_inst_pe_1_3_7_n75, npu_inst_pe_1_3_7_n74, npu_inst_pe_1_3_7_n73,
         npu_inst_pe_1_3_7_n72, npu_inst_pe_1_3_7_n71, npu_inst_pe_1_3_7_n70,
         npu_inst_pe_1_3_7_n69, npu_inst_pe_1_3_7_n68, npu_inst_pe_1_3_7_n67,
         npu_inst_pe_1_3_7_n66, npu_inst_pe_1_3_7_n65, npu_inst_pe_1_3_7_n64,
         npu_inst_pe_1_3_7_n63, npu_inst_pe_1_3_7_n62, npu_inst_pe_1_3_7_n61,
         npu_inst_pe_1_3_7_n60, npu_inst_pe_1_3_7_n59, npu_inst_pe_1_3_7_n58,
         npu_inst_pe_1_3_7_n57, npu_inst_pe_1_3_7_n56, npu_inst_pe_1_3_7_n55,
         npu_inst_pe_1_3_7_n54, npu_inst_pe_1_3_7_n53, npu_inst_pe_1_3_7_n52,
         npu_inst_pe_1_3_7_n51, npu_inst_pe_1_3_7_n50, npu_inst_pe_1_3_7_n49,
         npu_inst_pe_1_3_7_n48, npu_inst_pe_1_3_7_n47, npu_inst_pe_1_3_7_n46,
         npu_inst_pe_1_3_7_n45, npu_inst_pe_1_3_7_n44, npu_inst_pe_1_3_7_n43,
         npu_inst_pe_1_3_7_n42, npu_inst_pe_1_3_7_n41, npu_inst_pe_1_3_7_n40,
         npu_inst_pe_1_3_7_n39, npu_inst_pe_1_3_7_n38, npu_inst_pe_1_3_7_n37,
         npu_inst_pe_1_3_7_n27, npu_inst_pe_1_3_7_n26,
         npu_inst_pe_1_3_7_net3855, npu_inst_pe_1_3_7_net3849,
         npu_inst_pe_1_3_7_N94, npu_inst_pe_1_3_7_N93, npu_inst_pe_1_3_7_N84,
         npu_inst_pe_1_3_7_N80, npu_inst_pe_1_3_7_N79, npu_inst_pe_1_3_7_N78,
         npu_inst_pe_1_3_7_N77, npu_inst_pe_1_3_7_N76, npu_inst_pe_1_3_7_N75,
         npu_inst_pe_1_3_7_N74, npu_inst_pe_1_3_7_N73, npu_inst_pe_1_3_7_N72,
         npu_inst_pe_1_3_7_N71, npu_inst_pe_1_3_7_N70, npu_inst_pe_1_3_7_N69,
         npu_inst_pe_1_3_7_N68, npu_inst_pe_1_3_7_N67, npu_inst_pe_1_3_7_N66,
         npu_inst_pe_1_3_7_N65, npu_inst_pe_1_3_7_int_q_acc_0_,
         npu_inst_pe_1_3_7_int_q_acc_1_, npu_inst_pe_1_3_7_int_q_acc_2_,
         npu_inst_pe_1_3_7_int_q_acc_3_, npu_inst_pe_1_3_7_int_q_acc_4_,
         npu_inst_pe_1_3_7_int_q_acc_5_, npu_inst_pe_1_3_7_int_q_acc_6_,
         npu_inst_pe_1_3_7_int_q_acc_7_, npu_inst_pe_1_3_7_int_data_0_,
         npu_inst_pe_1_3_7_int_data_1_, npu_inst_pe_1_3_7_int_q_weight_0_,
         npu_inst_pe_1_3_7_int_q_weight_1_,
         npu_inst_pe_1_3_7_int_q_reg_v_5__0_,
         npu_inst_pe_1_3_7_int_q_reg_v_5__1_,
         npu_inst_pe_1_3_7_int_q_reg_v_4__0_,
         npu_inst_pe_1_3_7_int_q_reg_v_4__1_,
         npu_inst_pe_1_3_7_int_q_reg_v_3__0_,
         npu_inst_pe_1_3_7_int_q_reg_v_3__1_,
         npu_inst_pe_1_3_7_int_q_reg_v_2__0_,
         npu_inst_pe_1_3_7_int_q_reg_v_2__1_,
         npu_inst_pe_1_3_7_int_q_reg_v_1__0_,
         npu_inst_pe_1_3_7_int_q_reg_v_1__1_,
         npu_inst_pe_1_3_7_int_q_reg_v_0__0_,
         npu_inst_pe_1_3_7_int_q_reg_v_0__1_,
         npu_inst_pe_1_3_7_int_q_reg_h_5__0_,
         npu_inst_pe_1_3_7_int_q_reg_h_5__1_,
         npu_inst_pe_1_3_7_int_q_reg_h_4__0_,
         npu_inst_pe_1_3_7_int_q_reg_h_4__1_,
         npu_inst_pe_1_3_7_int_q_reg_h_3__0_,
         npu_inst_pe_1_3_7_int_q_reg_h_3__1_,
         npu_inst_pe_1_3_7_int_q_reg_h_2__0_,
         npu_inst_pe_1_3_7_int_q_reg_h_2__1_,
         npu_inst_pe_1_3_7_int_q_reg_h_1__0_,
         npu_inst_pe_1_3_7_int_q_reg_h_1__1_,
         npu_inst_pe_1_3_7_int_q_reg_h_0__0_,
         npu_inst_pe_1_3_7_int_q_reg_h_0__1_, npu_inst_pe_1_4_0_n119,
         npu_inst_pe_1_4_0_n118, npu_inst_pe_1_4_0_n117,
         npu_inst_pe_1_4_0_n116, npu_inst_pe_1_4_0_n115,
         npu_inst_pe_1_4_0_n114, npu_inst_pe_1_4_0_n113,
         npu_inst_pe_1_4_0_n112, npu_inst_pe_1_4_0_n111,
         npu_inst_pe_1_4_0_n110, npu_inst_pe_1_4_0_n109,
         npu_inst_pe_1_4_0_n108, npu_inst_pe_1_4_0_n107,
         npu_inst_pe_1_4_0_n106, npu_inst_pe_1_4_0_n105,
         npu_inst_pe_1_4_0_n104, npu_inst_pe_1_4_0_n103,
         npu_inst_pe_1_4_0_n102, npu_inst_pe_1_4_0_n101,
         npu_inst_pe_1_4_0_n100, npu_inst_pe_1_4_0_n99, npu_inst_pe_1_4_0_n98,
         npu_inst_pe_1_4_0_n36, npu_inst_pe_1_4_0_n35, npu_inst_pe_1_4_0_n34,
         npu_inst_pe_1_4_0_n33, npu_inst_pe_1_4_0_n32, npu_inst_pe_1_4_0_n31,
         npu_inst_pe_1_4_0_n30, npu_inst_pe_1_4_0_n29, npu_inst_pe_1_4_0_n28,
         npu_inst_pe_1_4_0_n25, npu_inst_pe_1_4_0_n24, npu_inst_pe_1_4_0_n23,
         npu_inst_pe_1_4_0_n22, npu_inst_pe_1_4_0_n21, npu_inst_pe_1_4_0_n20,
         npu_inst_pe_1_4_0_n19, npu_inst_pe_1_4_0_n18, npu_inst_pe_1_4_0_n17,
         npu_inst_pe_1_4_0_n16, npu_inst_pe_1_4_0_n15, npu_inst_pe_1_4_0_n14,
         npu_inst_pe_1_4_0_n13, npu_inst_pe_1_4_0_n12, npu_inst_pe_1_4_0_n11,
         npu_inst_pe_1_4_0_n10, npu_inst_pe_1_4_0_n9, npu_inst_pe_1_4_0_n8,
         npu_inst_pe_1_4_0_n7, npu_inst_pe_1_4_0_n6, npu_inst_pe_1_4_0_n5,
         npu_inst_pe_1_4_0_n4, npu_inst_pe_1_4_0_n3, npu_inst_pe_1_4_0_n2,
         npu_inst_pe_1_4_0_n1, npu_inst_pe_1_4_0_sub_67_carry_7_,
         npu_inst_pe_1_4_0_sub_67_carry_6_, npu_inst_pe_1_4_0_sub_67_carry_5_,
         npu_inst_pe_1_4_0_sub_67_carry_4_, npu_inst_pe_1_4_0_sub_67_carry_3_,
         npu_inst_pe_1_4_0_sub_67_carry_2_, npu_inst_pe_1_4_0_sub_67_carry_1_,
         npu_inst_pe_1_4_0_add_69_carry_7_, npu_inst_pe_1_4_0_add_69_carry_6_,
         npu_inst_pe_1_4_0_add_69_carry_5_, npu_inst_pe_1_4_0_add_69_carry_4_,
         npu_inst_pe_1_4_0_add_69_carry_3_, npu_inst_pe_1_4_0_add_69_carry_2_,
         npu_inst_pe_1_4_0_add_69_carry_1_, npu_inst_pe_1_4_0_n97,
         npu_inst_pe_1_4_0_n96, npu_inst_pe_1_4_0_n95, npu_inst_pe_1_4_0_n94,
         npu_inst_pe_1_4_0_n93, npu_inst_pe_1_4_0_n92, npu_inst_pe_1_4_0_n91,
         npu_inst_pe_1_4_0_n90, npu_inst_pe_1_4_0_n89, npu_inst_pe_1_4_0_n88,
         npu_inst_pe_1_4_0_n87, npu_inst_pe_1_4_0_n86, npu_inst_pe_1_4_0_n85,
         npu_inst_pe_1_4_0_n84, npu_inst_pe_1_4_0_n83, npu_inst_pe_1_4_0_n82,
         npu_inst_pe_1_4_0_n81, npu_inst_pe_1_4_0_n80, npu_inst_pe_1_4_0_n79,
         npu_inst_pe_1_4_0_n78, npu_inst_pe_1_4_0_n77, npu_inst_pe_1_4_0_n76,
         npu_inst_pe_1_4_0_n75, npu_inst_pe_1_4_0_n74, npu_inst_pe_1_4_0_n73,
         npu_inst_pe_1_4_0_n72, npu_inst_pe_1_4_0_n71, npu_inst_pe_1_4_0_n70,
         npu_inst_pe_1_4_0_n69, npu_inst_pe_1_4_0_n68, npu_inst_pe_1_4_0_n67,
         npu_inst_pe_1_4_0_n66, npu_inst_pe_1_4_0_n65, npu_inst_pe_1_4_0_n64,
         npu_inst_pe_1_4_0_n63, npu_inst_pe_1_4_0_n62, npu_inst_pe_1_4_0_n61,
         npu_inst_pe_1_4_0_n60, npu_inst_pe_1_4_0_n59, npu_inst_pe_1_4_0_n58,
         npu_inst_pe_1_4_0_n57, npu_inst_pe_1_4_0_n56, npu_inst_pe_1_4_0_n55,
         npu_inst_pe_1_4_0_n54, npu_inst_pe_1_4_0_n53, npu_inst_pe_1_4_0_n52,
         npu_inst_pe_1_4_0_n51, npu_inst_pe_1_4_0_n50, npu_inst_pe_1_4_0_n49,
         npu_inst_pe_1_4_0_n48, npu_inst_pe_1_4_0_n47, npu_inst_pe_1_4_0_n46,
         npu_inst_pe_1_4_0_n45, npu_inst_pe_1_4_0_n44, npu_inst_pe_1_4_0_n43,
         npu_inst_pe_1_4_0_n42, npu_inst_pe_1_4_0_n41, npu_inst_pe_1_4_0_n40,
         npu_inst_pe_1_4_0_n39, npu_inst_pe_1_4_0_n38, npu_inst_pe_1_4_0_n37,
         npu_inst_pe_1_4_0_n27, npu_inst_pe_1_4_0_n26,
         npu_inst_pe_1_4_0_net3832, npu_inst_pe_1_4_0_net3826,
         npu_inst_pe_1_4_0_N94, npu_inst_pe_1_4_0_N93, npu_inst_pe_1_4_0_N84,
         npu_inst_pe_1_4_0_N80, npu_inst_pe_1_4_0_N79, npu_inst_pe_1_4_0_N78,
         npu_inst_pe_1_4_0_N77, npu_inst_pe_1_4_0_N76, npu_inst_pe_1_4_0_N75,
         npu_inst_pe_1_4_0_N74, npu_inst_pe_1_4_0_N73, npu_inst_pe_1_4_0_N72,
         npu_inst_pe_1_4_0_N71, npu_inst_pe_1_4_0_N70, npu_inst_pe_1_4_0_N69,
         npu_inst_pe_1_4_0_N68, npu_inst_pe_1_4_0_N67, npu_inst_pe_1_4_0_N66,
         npu_inst_pe_1_4_0_N65, npu_inst_pe_1_4_0_int_q_acc_0_,
         npu_inst_pe_1_4_0_int_q_acc_1_, npu_inst_pe_1_4_0_int_q_acc_2_,
         npu_inst_pe_1_4_0_int_q_acc_3_, npu_inst_pe_1_4_0_int_q_acc_4_,
         npu_inst_pe_1_4_0_int_q_acc_5_, npu_inst_pe_1_4_0_int_q_acc_6_,
         npu_inst_pe_1_4_0_int_q_acc_7_, npu_inst_pe_1_4_0_int_data_0_,
         npu_inst_pe_1_4_0_int_data_1_, npu_inst_pe_1_4_0_int_q_weight_0_,
         npu_inst_pe_1_4_0_int_q_weight_1_,
         npu_inst_pe_1_4_0_int_q_reg_v_5__0_,
         npu_inst_pe_1_4_0_int_q_reg_v_5__1_,
         npu_inst_pe_1_4_0_int_q_reg_v_4__0_,
         npu_inst_pe_1_4_0_int_q_reg_v_4__1_,
         npu_inst_pe_1_4_0_int_q_reg_v_3__0_,
         npu_inst_pe_1_4_0_int_q_reg_v_3__1_,
         npu_inst_pe_1_4_0_int_q_reg_v_2__0_,
         npu_inst_pe_1_4_0_int_q_reg_v_2__1_,
         npu_inst_pe_1_4_0_int_q_reg_v_1__0_,
         npu_inst_pe_1_4_0_int_q_reg_v_1__1_,
         npu_inst_pe_1_4_0_int_q_reg_v_0__0_,
         npu_inst_pe_1_4_0_int_q_reg_v_0__1_,
         npu_inst_pe_1_4_0_int_q_reg_h_5__0_,
         npu_inst_pe_1_4_0_int_q_reg_h_5__1_,
         npu_inst_pe_1_4_0_int_q_reg_h_4__0_,
         npu_inst_pe_1_4_0_int_q_reg_h_4__1_,
         npu_inst_pe_1_4_0_int_q_reg_h_3__0_,
         npu_inst_pe_1_4_0_int_q_reg_h_3__1_,
         npu_inst_pe_1_4_0_int_q_reg_h_2__0_,
         npu_inst_pe_1_4_0_int_q_reg_h_2__1_,
         npu_inst_pe_1_4_0_int_q_reg_h_1__0_,
         npu_inst_pe_1_4_0_int_q_reg_h_1__1_,
         npu_inst_pe_1_4_0_int_q_reg_h_0__0_,
         npu_inst_pe_1_4_0_int_q_reg_h_0__1_, npu_inst_pe_1_4_0_o_data_h_0_,
         npu_inst_pe_1_4_0_o_data_h_1_, npu_inst_pe_1_4_1_n119,
         npu_inst_pe_1_4_1_n118, npu_inst_pe_1_4_1_n117,
         npu_inst_pe_1_4_1_n116, npu_inst_pe_1_4_1_n115,
         npu_inst_pe_1_4_1_n114, npu_inst_pe_1_4_1_n113,
         npu_inst_pe_1_4_1_n112, npu_inst_pe_1_4_1_n111,
         npu_inst_pe_1_4_1_n110, npu_inst_pe_1_4_1_n109,
         npu_inst_pe_1_4_1_n108, npu_inst_pe_1_4_1_n107,
         npu_inst_pe_1_4_1_n106, npu_inst_pe_1_4_1_n105,
         npu_inst_pe_1_4_1_n104, npu_inst_pe_1_4_1_n103,
         npu_inst_pe_1_4_1_n102, npu_inst_pe_1_4_1_n101,
         npu_inst_pe_1_4_1_n100, npu_inst_pe_1_4_1_n99, npu_inst_pe_1_4_1_n98,
         npu_inst_pe_1_4_1_n36, npu_inst_pe_1_4_1_n35, npu_inst_pe_1_4_1_n34,
         npu_inst_pe_1_4_1_n33, npu_inst_pe_1_4_1_n32, npu_inst_pe_1_4_1_n31,
         npu_inst_pe_1_4_1_n30, npu_inst_pe_1_4_1_n29, npu_inst_pe_1_4_1_n28,
         npu_inst_pe_1_4_1_n25, npu_inst_pe_1_4_1_n24, npu_inst_pe_1_4_1_n23,
         npu_inst_pe_1_4_1_n22, npu_inst_pe_1_4_1_n21, npu_inst_pe_1_4_1_n20,
         npu_inst_pe_1_4_1_n19, npu_inst_pe_1_4_1_n18, npu_inst_pe_1_4_1_n17,
         npu_inst_pe_1_4_1_n16, npu_inst_pe_1_4_1_n15, npu_inst_pe_1_4_1_n14,
         npu_inst_pe_1_4_1_n13, npu_inst_pe_1_4_1_n12, npu_inst_pe_1_4_1_n11,
         npu_inst_pe_1_4_1_n10, npu_inst_pe_1_4_1_n9, npu_inst_pe_1_4_1_n8,
         npu_inst_pe_1_4_1_n7, npu_inst_pe_1_4_1_n6, npu_inst_pe_1_4_1_n5,
         npu_inst_pe_1_4_1_n4, npu_inst_pe_1_4_1_n3, npu_inst_pe_1_4_1_n2,
         npu_inst_pe_1_4_1_n1, npu_inst_pe_1_4_1_sub_67_carry_7_,
         npu_inst_pe_1_4_1_sub_67_carry_6_, npu_inst_pe_1_4_1_sub_67_carry_5_,
         npu_inst_pe_1_4_1_sub_67_carry_4_, npu_inst_pe_1_4_1_sub_67_carry_3_,
         npu_inst_pe_1_4_1_sub_67_carry_2_, npu_inst_pe_1_4_1_sub_67_carry_1_,
         npu_inst_pe_1_4_1_add_69_carry_7_, npu_inst_pe_1_4_1_add_69_carry_6_,
         npu_inst_pe_1_4_1_add_69_carry_5_, npu_inst_pe_1_4_1_add_69_carry_4_,
         npu_inst_pe_1_4_1_add_69_carry_3_, npu_inst_pe_1_4_1_add_69_carry_2_,
         npu_inst_pe_1_4_1_add_69_carry_1_, npu_inst_pe_1_4_1_n97,
         npu_inst_pe_1_4_1_n96, npu_inst_pe_1_4_1_n95, npu_inst_pe_1_4_1_n94,
         npu_inst_pe_1_4_1_n93, npu_inst_pe_1_4_1_n92, npu_inst_pe_1_4_1_n91,
         npu_inst_pe_1_4_1_n90, npu_inst_pe_1_4_1_n89, npu_inst_pe_1_4_1_n88,
         npu_inst_pe_1_4_1_n87, npu_inst_pe_1_4_1_n86, npu_inst_pe_1_4_1_n85,
         npu_inst_pe_1_4_1_n84, npu_inst_pe_1_4_1_n83, npu_inst_pe_1_4_1_n82,
         npu_inst_pe_1_4_1_n81, npu_inst_pe_1_4_1_n80, npu_inst_pe_1_4_1_n79,
         npu_inst_pe_1_4_1_n78, npu_inst_pe_1_4_1_n77, npu_inst_pe_1_4_1_n76,
         npu_inst_pe_1_4_1_n75, npu_inst_pe_1_4_1_n74, npu_inst_pe_1_4_1_n73,
         npu_inst_pe_1_4_1_n72, npu_inst_pe_1_4_1_n71, npu_inst_pe_1_4_1_n70,
         npu_inst_pe_1_4_1_n69, npu_inst_pe_1_4_1_n68, npu_inst_pe_1_4_1_n67,
         npu_inst_pe_1_4_1_n66, npu_inst_pe_1_4_1_n65, npu_inst_pe_1_4_1_n64,
         npu_inst_pe_1_4_1_n63, npu_inst_pe_1_4_1_n62, npu_inst_pe_1_4_1_n61,
         npu_inst_pe_1_4_1_n60, npu_inst_pe_1_4_1_n59, npu_inst_pe_1_4_1_n58,
         npu_inst_pe_1_4_1_n57, npu_inst_pe_1_4_1_n56, npu_inst_pe_1_4_1_n55,
         npu_inst_pe_1_4_1_n54, npu_inst_pe_1_4_1_n53, npu_inst_pe_1_4_1_n52,
         npu_inst_pe_1_4_1_n51, npu_inst_pe_1_4_1_n50, npu_inst_pe_1_4_1_n49,
         npu_inst_pe_1_4_1_n48, npu_inst_pe_1_4_1_n47, npu_inst_pe_1_4_1_n46,
         npu_inst_pe_1_4_1_n45, npu_inst_pe_1_4_1_n44, npu_inst_pe_1_4_1_n43,
         npu_inst_pe_1_4_1_n42, npu_inst_pe_1_4_1_n41, npu_inst_pe_1_4_1_n40,
         npu_inst_pe_1_4_1_n39, npu_inst_pe_1_4_1_n38, npu_inst_pe_1_4_1_n37,
         npu_inst_pe_1_4_1_n27, npu_inst_pe_1_4_1_n26,
         npu_inst_pe_1_4_1_net3809, npu_inst_pe_1_4_1_net3803,
         npu_inst_pe_1_4_1_N94, npu_inst_pe_1_4_1_N93, npu_inst_pe_1_4_1_N84,
         npu_inst_pe_1_4_1_N80, npu_inst_pe_1_4_1_N79, npu_inst_pe_1_4_1_N78,
         npu_inst_pe_1_4_1_N77, npu_inst_pe_1_4_1_N76, npu_inst_pe_1_4_1_N75,
         npu_inst_pe_1_4_1_N74, npu_inst_pe_1_4_1_N73, npu_inst_pe_1_4_1_N72,
         npu_inst_pe_1_4_1_N71, npu_inst_pe_1_4_1_N70, npu_inst_pe_1_4_1_N69,
         npu_inst_pe_1_4_1_N68, npu_inst_pe_1_4_1_N67, npu_inst_pe_1_4_1_N66,
         npu_inst_pe_1_4_1_N65, npu_inst_pe_1_4_1_int_q_acc_0_,
         npu_inst_pe_1_4_1_int_q_acc_1_, npu_inst_pe_1_4_1_int_q_acc_2_,
         npu_inst_pe_1_4_1_int_q_acc_3_, npu_inst_pe_1_4_1_int_q_acc_4_,
         npu_inst_pe_1_4_1_int_q_acc_5_, npu_inst_pe_1_4_1_int_q_acc_6_,
         npu_inst_pe_1_4_1_int_q_acc_7_, npu_inst_pe_1_4_1_int_data_0_,
         npu_inst_pe_1_4_1_int_data_1_, npu_inst_pe_1_4_1_int_q_weight_0_,
         npu_inst_pe_1_4_1_int_q_weight_1_,
         npu_inst_pe_1_4_1_int_q_reg_v_5__0_,
         npu_inst_pe_1_4_1_int_q_reg_v_5__1_,
         npu_inst_pe_1_4_1_int_q_reg_v_4__0_,
         npu_inst_pe_1_4_1_int_q_reg_v_4__1_,
         npu_inst_pe_1_4_1_int_q_reg_v_3__0_,
         npu_inst_pe_1_4_1_int_q_reg_v_3__1_,
         npu_inst_pe_1_4_1_int_q_reg_v_2__0_,
         npu_inst_pe_1_4_1_int_q_reg_v_2__1_,
         npu_inst_pe_1_4_1_int_q_reg_v_1__0_,
         npu_inst_pe_1_4_1_int_q_reg_v_1__1_,
         npu_inst_pe_1_4_1_int_q_reg_v_0__0_,
         npu_inst_pe_1_4_1_int_q_reg_v_0__1_,
         npu_inst_pe_1_4_1_int_q_reg_h_5__0_,
         npu_inst_pe_1_4_1_int_q_reg_h_5__1_,
         npu_inst_pe_1_4_1_int_q_reg_h_4__0_,
         npu_inst_pe_1_4_1_int_q_reg_h_4__1_,
         npu_inst_pe_1_4_1_int_q_reg_h_3__0_,
         npu_inst_pe_1_4_1_int_q_reg_h_3__1_,
         npu_inst_pe_1_4_1_int_q_reg_h_2__0_,
         npu_inst_pe_1_4_1_int_q_reg_h_2__1_,
         npu_inst_pe_1_4_1_int_q_reg_h_1__0_,
         npu_inst_pe_1_4_1_int_q_reg_h_1__1_,
         npu_inst_pe_1_4_1_int_q_reg_h_0__0_,
         npu_inst_pe_1_4_1_int_q_reg_h_0__1_, npu_inst_pe_1_4_2_n119,
         npu_inst_pe_1_4_2_n118, npu_inst_pe_1_4_2_n117,
         npu_inst_pe_1_4_2_n116, npu_inst_pe_1_4_2_n115,
         npu_inst_pe_1_4_2_n114, npu_inst_pe_1_4_2_n113,
         npu_inst_pe_1_4_2_n112, npu_inst_pe_1_4_2_n111,
         npu_inst_pe_1_4_2_n110, npu_inst_pe_1_4_2_n109,
         npu_inst_pe_1_4_2_n108, npu_inst_pe_1_4_2_n107,
         npu_inst_pe_1_4_2_n106, npu_inst_pe_1_4_2_n105,
         npu_inst_pe_1_4_2_n104, npu_inst_pe_1_4_2_n103,
         npu_inst_pe_1_4_2_n102, npu_inst_pe_1_4_2_n101,
         npu_inst_pe_1_4_2_n100, npu_inst_pe_1_4_2_n99, npu_inst_pe_1_4_2_n98,
         npu_inst_pe_1_4_2_n36, npu_inst_pe_1_4_2_n35, npu_inst_pe_1_4_2_n34,
         npu_inst_pe_1_4_2_n33, npu_inst_pe_1_4_2_n32, npu_inst_pe_1_4_2_n31,
         npu_inst_pe_1_4_2_n30, npu_inst_pe_1_4_2_n29, npu_inst_pe_1_4_2_n28,
         npu_inst_pe_1_4_2_n25, npu_inst_pe_1_4_2_n24, npu_inst_pe_1_4_2_n23,
         npu_inst_pe_1_4_2_n22, npu_inst_pe_1_4_2_n21, npu_inst_pe_1_4_2_n20,
         npu_inst_pe_1_4_2_n19, npu_inst_pe_1_4_2_n18, npu_inst_pe_1_4_2_n17,
         npu_inst_pe_1_4_2_n16, npu_inst_pe_1_4_2_n15, npu_inst_pe_1_4_2_n14,
         npu_inst_pe_1_4_2_n13, npu_inst_pe_1_4_2_n12, npu_inst_pe_1_4_2_n11,
         npu_inst_pe_1_4_2_n10, npu_inst_pe_1_4_2_n9, npu_inst_pe_1_4_2_n8,
         npu_inst_pe_1_4_2_n7, npu_inst_pe_1_4_2_n6, npu_inst_pe_1_4_2_n5,
         npu_inst_pe_1_4_2_n4, npu_inst_pe_1_4_2_n3, npu_inst_pe_1_4_2_n2,
         npu_inst_pe_1_4_2_n1, npu_inst_pe_1_4_2_sub_67_carry_7_,
         npu_inst_pe_1_4_2_sub_67_carry_6_, npu_inst_pe_1_4_2_sub_67_carry_5_,
         npu_inst_pe_1_4_2_sub_67_carry_4_, npu_inst_pe_1_4_2_sub_67_carry_3_,
         npu_inst_pe_1_4_2_sub_67_carry_2_, npu_inst_pe_1_4_2_sub_67_carry_1_,
         npu_inst_pe_1_4_2_add_69_carry_7_, npu_inst_pe_1_4_2_add_69_carry_6_,
         npu_inst_pe_1_4_2_add_69_carry_5_, npu_inst_pe_1_4_2_add_69_carry_4_,
         npu_inst_pe_1_4_2_add_69_carry_3_, npu_inst_pe_1_4_2_add_69_carry_2_,
         npu_inst_pe_1_4_2_add_69_carry_1_, npu_inst_pe_1_4_2_n97,
         npu_inst_pe_1_4_2_n96, npu_inst_pe_1_4_2_n95, npu_inst_pe_1_4_2_n94,
         npu_inst_pe_1_4_2_n93, npu_inst_pe_1_4_2_n92, npu_inst_pe_1_4_2_n91,
         npu_inst_pe_1_4_2_n90, npu_inst_pe_1_4_2_n89, npu_inst_pe_1_4_2_n88,
         npu_inst_pe_1_4_2_n87, npu_inst_pe_1_4_2_n86, npu_inst_pe_1_4_2_n85,
         npu_inst_pe_1_4_2_n84, npu_inst_pe_1_4_2_n83, npu_inst_pe_1_4_2_n82,
         npu_inst_pe_1_4_2_n81, npu_inst_pe_1_4_2_n80, npu_inst_pe_1_4_2_n79,
         npu_inst_pe_1_4_2_n78, npu_inst_pe_1_4_2_n77, npu_inst_pe_1_4_2_n76,
         npu_inst_pe_1_4_2_n75, npu_inst_pe_1_4_2_n74, npu_inst_pe_1_4_2_n73,
         npu_inst_pe_1_4_2_n72, npu_inst_pe_1_4_2_n71, npu_inst_pe_1_4_2_n70,
         npu_inst_pe_1_4_2_n69, npu_inst_pe_1_4_2_n68, npu_inst_pe_1_4_2_n67,
         npu_inst_pe_1_4_2_n66, npu_inst_pe_1_4_2_n65, npu_inst_pe_1_4_2_n64,
         npu_inst_pe_1_4_2_n63, npu_inst_pe_1_4_2_n62, npu_inst_pe_1_4_2_n61,
         npu_inst_pe_1_4_2_n60, npu_inst_pe_1_4_2_n59, npu_inst_pe_1_4_2_n58,
         npu_inst_pe_1_4_2_n57, npu_inst_pe_1_4_2_n56, npu_inst_pe_1_4_2_n55,
         npu_inst_pe_1_4_2_n54, npu_inst_pe_1_4_2_n53, npu_inst_pe_1_4_2_n52,
         npu_inst_pe_1_4_2_n51, npu_inst_pe_1_4_2_n50, npu_inst_pe_1_4_2_n49,
         npu_inst_pe_1_4_2_n48, npu_inst_pe_1_4_2_n47, npu_inst_pe_1_4_2_n46,
         npu_inst_pe_1_4_2_n45, npu_inst_pe_1_4_2_n44, npu_inst_pe_1_4_2_n43,
         npu_inst_pe_1_4_2_n42, npu_inst_pe_1_4_2_n41, npu_inst_pe_1_4_2_n40,
         npu_inst_pe_1_4_2_n39, npu_inst_pe_1_4_2_n38, npu_inst_pe_1_4_2_n37,
         npu_inst_pe_1_4_2_n27, npu_inst_pe_1_4_2_n26,
         npu_inst_pe_1_4_2_net3786, npu_inst_pe_1_4_2_net3780,
         npu_inst_pe_1_4_2_N94, npu_inst_pe_1_4_2_N93, npu_inst_pe_1_4_2_N84,
         npu_inst_pe_1_4_2_N80, npu_inst_pe_1_4_2_N79, npu_inst_pe_1_4_2_N78,
         npu_inst_pe_1_4_2_N77, npu_inst_pe_1_4_2_N76, npu_inst_pe_1_4_2_N75,
         npu_inst_pe_1_4_2_N74, npu_inst_pe_1_4_2_N73, npu_inst_pe_1_4_2_N72,
         npu_inst_pe_1_4_2_N71, npu_inst_pe_1_4_2_N70, npu_inst_pe_1_4_2_N69,
         npu_inst_pe_1_4_2_N68, npu_inst_pe_1_4_2_N67, npu_inst_pe_1_4_2_N66,
         npu_inst_pe_1_4_2_N65, npu_inst_pe_1_4_2_int_q_acc_0_,
         npu_inst_pe_1_4_2_int_q_acc_1_, npu_inst_pe_1_4_2_int_q_acc_2_,
         npu_inst_pe_1_4_2_int_q_acc_3_, npu_inst_pe_1_4_2_int_q_acc_4_,
         npu_inst_pe_1_4_2_int_q_acc_5_, npu_inst_pe_1_4_2_int_q_acc_6_,
         npu_inst_pe_1_4_2_int_q_acc_7_, npu_inst_pe_1_4_2_int_data_0_,
         npu_inst_pe_1_4_2_int_data_1_, npu_inst_pe_1_4_2_int_q_weight_0_,
         npu_inst_pe_1_4_2_int_q_weight_1_,
         npu_inst_pe_1_4_2_int_q_reg_v_5__0_,
         npu_inst_pe_1_4_2_int_q_reg_v_5__1_,
         npu_inst_pe_1_4_2_int_q_reg_v_4__0_,
         npu_inst_pe_1_4_2_int_q_reg_v_4__1_,
         npu_inst_pe_1_4_2_int_q_reg_v_3__0_,
         npu_inst_pe_1_4_2_int_q_reg_v_3__1_,
         npu_inst_pe_1_4_2_int_q_reg_v_2__0_,
         npu_inst_pe_1_4_2_int_q_reg_v_2__1_,
         npu_inst_pe_1_4_2_int_q_reg_v_1__0_,
         npu_inst_pe_1_4_2_int_q_reg_v_1__1_,
         npu_inst_pe_1_4_2_int_q_reg_v_0__0_,
         npu_inst_pe_1_4_2_int_q_reg_v_0__1_,
         npu_inst_pe_1_4_2_int_q_reg_h_5__0_,
         npu_inst_pe_1_4_2_int_q_reg_h_5__1_,
         npu_inst_pe_1_4_2_int_q_reg_h_4__0_,
         npu_inst_pe_1_4_2_int_q_reg_h_4__1_,
         npu_inst_pe_1_4_2_int_q_reg_h_3__0_,
         npu_inst_pe_1_4_2_int_q_reg_h_3__1_,
         npu_inst_pe_1_4_2_int_q_reg_h_2__0_,
         npu_inst_pe_1_4_2_int_q_reg_h_2__1_,
         npu_inst_pe_1_4_2_int_q_reg_h_1__0_,
         npu_inst_pe_1_4_2_int_q_reg_h_1__1_,
         npu_inst_pe_1_4_2_int_q_reg_h_0__0_,
         npu_inst_pe_1_4_2_int_q_reg_h_0__1_, npu_inst_pe_1_4_3_n119,
         npu_inst_pe_1_4_3_n118, npu_inst_pe_1_4_3_n117,
         npu_inst_pe_1_4_3_n116, npu_inst_pe_1_4_3_n115,
         npu_inst_pe_1_4_3_n114, npu_inst_pe_1_4_3_n113,
         npu_inst_pe_1_4_3_n112, npu_inst_pe_1_4_3_n111,
         npu_inst_pe_1_4_3_n110, npu_inst_pe_1_4_3_n109,
         npu_inst_pe_1_4_3_n108, npu_inst_pe_1_4_3_n107,
         npu_inst_pe_1_4_3_n106, npu_inst_pe_1_4_3_n105,
         npu_inst_pe_1_4_3_n104, npu_inst_pe_1_4_3_n103,
         npu_inst_pe_1_4_3_n102, npu_inst_pe_1_4_3_n101,
         npu_inst_pe_1_4_3_n100, npu_inst_pe_1_4_3_n99, npu_inst_pe_1_4_3_n98,
         npu_inst_pe_1_4_3_n36, npu_inst_pe_1_4_3_n35, npu_inst_pe_1_4_3_n34,
         npu_inst_pe_1_4_3_n33, npu_inst_pe_1_4_3_n32, npu_inst_pe_1_4_3_n31,
         npu_inst_pe_1_4_3_n30, npu_inst_pe_1_4_3_n29, npu_inst_pe_1_4_3_n28,
         npu_inst_pe_1_4_3_n25, npu_inst_pe_1_4_3_n24, npu_inst_pe_1_4_3_n23,
         npu_inst_pe_1_4_3_n22, npu_inst_pe_1_4_3_n21, npu_inst_pe_1_4_3_n20,
         npu_inst_pe_1_4_3_n19, npu_inst_pe_1_4_3_n18, npu_inst_pe_1_4_3_n17,
         npu_inst_pe_1_4_3_n16, npu_inst_pe_1_4_3_n15, npu_inst_pe_1_4_3_n14,
         npu_inst_pe_1_4_3_n13, npu_inst_pe_1_4_3_n12, npu_inst_pe_1_4_3_n11,
         npu_inst_pe_1_4_3_n10, npu_inst_pe_1_4_3_n9, npu_inst_pe_1_4_3_n8,
         npu_inst_pe_1_4_3_n7, npu_inst_pe_1_4_3_n6, npu_inst_pe_1_4_3_n5,
         npu_inst_pe_1_4_3_n4, npu_inst_pe_1_4_3_n3, npu_inst_pe_1_4_3_n2,
         npu_inst_pe_1_4_3_n1, npu_inst_pe_1_4_3_sub_67_carry_7_,
         npu_inst_pe_1_4_3_sub_67_carry_6_, npu_inst_pe_1_4_3_sub_67_carry_5_,
         npu_inst_pe_1_4_3_sub_67_carry_4_, npu_inst_pe_1_4_3_sub_67_carry_3_,
         npu_inst_pe_1_4_3_sub_67_carry_2_, npu_inst_pe_1_4_3_sub_67_carry_1_,
         npu_inst_pe_1_4_3_add_69_carry_7_, npu_inst_pe_1_4_3_add_69_carry_6_,
         npu_inst_pe_1_4_3_add_69_carry_5_, npu_inst_pe_1_4_3_add_69_carry_4_,
         npu_inst_pe_1_4_3_add_69_carry_3_, npu_inst_pe_1_4_3_add_69_carry_2_,
         npu_inst_pe_1_4_3_add_69_carry_1_, npu_inst_pe_1_4_3_n97,
         npu_inst_pe_1_4_3_n96, npu_inst_pe_1_4_3_n95, npu_inst_pe_1_4_3_n94,
         npu_inst_pe_1_4_3_n93, npu_inst_pe_1_4_3_n92, npu_inst_pe_1_4_3_n91,
         npu_inst_pe_1_4_3_n90, npu_inst_pe_1_4_3_n89, npu_inst_pe_1_4_3_n88,
         npu_inst_pe_1_4_3_n87, npu_inst_pe_1_4_3_n86, npu_inst_pe_1_4_3_n85,
         npu_inst_pe_1_4_3_n84, npu_inst_pe_1_4_3_n83, npu_inst_pe_1_4_3_n82,
         npu_inst_pe_1_4_3_n81, npu_inst_pe_1_4_3_n80, npu_inst_pe_1_4_3_n79,
         npu_inst_pe_1_4_3_n78, npu_inst_pe_1_4_3_n77, npu_inst_pe_1_4_3_n76,
         npu_inst_pe_1_4_3_n75, npu_inst_pe_1_4_3_n74, npu_inst_pe_1_4_3_n73,
         npu_inst_pe_1_4_3_n72, npu_inst_pe_1_4_3_n71, npu_inst_pe_1_4_3_n70,
         npu_inst_pe_1_4_3_n69, npu_inst_pe_1_4_3_n68, npu_inst_pe_1_4_3_n67,
         npu_inst_pe_1_4_3_n66, npu_inst_pe_1_4_3_n65, npu_inst_pe_1_4_3_n64,
         npu_inst_pe_1_4_3_n63, npu_inst_pe_1_4_3_n62, npu_inst_pe_1_4_3_n61,
         npu_inst_pe_1_4_3_n60, npu_inst_pe_1_4_3_n59, npu_inst_pe_1_4_3_n58,
         npu_inst_pe_1_4_3_n57, npu_inst_pe_1_4_3_n56, npu_inst_pe_1_4_3_n55,
         npu_inst_pe_1_4_3_n54, npu_inst_pe_1_4_3_n53, npu_inst_pe_1_4_3_n52,
         npu_inst_pe_1_4_3_n51, npu_inst_pe_1_4_3_n50, npu_inst_pe_1_4_3_n49,
         npu_inst_pe_1_4_3_n48, npu_inst_pe_1_4_3_n47, npu_inst_pe_1_4_3_n46,
         npu_inst_pe_1_4_3_n45, npu_inst_pe_1_4_3_n44, npu_inst_pe_1_4_3_n43,
         npu_inst_pe_1_4_3_n42, npu_inst_pe_1_4_3_n41, npu_inst_pe_1_4_3_n40,
         npu_inst_pe_1_4_3_n39, npu_inst_pe_1_4_3_n38, npu_inst_pe_1_4_3_n37,
         npu_inst_pe_1_4_3_n27, npu_inst_pe_1_4_3_n26,
         npu_inst_pe_1_4_3_net3763, npu_inst_pe_1_4_3_net3757,
         npu_inst_pe_1_4_3_N94, npu_inst_pe_1_4_3_N93, npu_inst_pe_1_4_3_N84,
         npu_inst_pe_1_4_3_N80, npu_inst_pe_1_4_3_N79, npu_inst_pe_1_4_3_N78,
         npu_inst_pe_1_4_3_N77, npu_inst_pe_1_4_3_N76, npu_inst_pe_1_4_3_N75,
         npu_inst_pe_1_4_3_N74, npu_inst_pe_1_4_3_N73, npu_inst_pe_1_4_3_N72,
         npu_inst_pe_1_4_3_N71, npu_inst_pe_1_4_3_N70, npu_inst_pe_1_4_3_N69,
         npu_inst_pe_1_4_3_N68, npu_inst_pe_1_4_3_N67, npu_inst_pe_1_4_3_N66,
         npu_inst_pe_1_4_3_N65, npu_inst_pe_1_4_3_int_q_acc_0_,
         npu_inst_pe_1_4_3_int_q_acc_1_, npu_inst_pe_1_4_3_int_q_acc_2_,
         npu_inst_pe_1_4_3_int_q_acc_3_, npu_inst_pe_1_4_3_int_q_acc_4_,
         npu_inst_pe_1_4_3_int_q_acc_5_, npu_inst_pe_1_4_3_int_q_acc_6_,
         npu_inst_pe_1_4_3_int_q_acc_7_, npu_inst_pe_1_4_3_int_data_0_,
         npu_inst_pe_1_4_3_int_data_1_, npu_inst_pe_1_4_3_int_q_weight_0_,
         npu_inst_pe_1_4_3_int_q_weight_1_,
         npu_inst_pe_1_4_3_int_q_reg_v_5__0_,
         npu_inst_pe_1_4_3_int_q_reg_v_5__1_,
         npu_inst_pe_1_4_3_int_q_reg_v_4__0_,
         npu_inst_pe_1_4_3_int_q_reg_v_4__1_,
         npu_inst_pe_1_4_3_int_q_reg_v_3__0_,
         npu_inst_pe_1_4_3_int_q_reg_v_3__1_,
         npu_inst_pe_1_4_3_int_q_reg_v_2__0_,
         npu_inst_pe_1_4_3_int_q_reg_v_2__1_,
         npu_inst_pe_1_4_3_int_q_reg_v_1__0_,
         npu_inst_pe_1_4_3_int_q_reg_v_1__1_,
         npu_inst_pe_1_4_3_int_q_reg_v_0__0_,
         npu_inst_pe_1_4_3_int_q_reg_v_0__1_,
         npu_inst_pe_1_4_3_int_q_reg_h_5__0_,
         npu_inst_pe_1_4_3_int_q_reg_h_5__1_,
         npu_inst_pe_1_4_3_int_q_reg_h_4__0_,
         npu_inst_pe_1_4_3_int_q_reg_h_4__1_,
         npu_inst_pe_1_4_3_int_q_reg_h_3__0_,
         npu_inst_pe_1_4_3_int_q_reg_h_3__1_,
         npu_inst_pe_1_4_3_int_q_reg_h_2__0_,
         npu_inst_pe_1_4_3_int_q_reg_h_2__1_,
         npu_inst_pe_1_4_3_int_q_reg_h_1__0_,
         npu_inst_pe_1_4_3_int_q_reg_h_1__1_,
         npu_inst_pe_1_4_3_int_q_reg_h_0__0_,
         npu_inst_pe_1_4_3_int_q_reg_h_0__1_, npu_inst_pe_1_4_4_n119,
         npu_inst_pe_1_4_4_n118, npu_inst_pe_1_4_4_n117,
         npu_inst_pe_1_4_4_n116, npu_inst_pe_1_4_4_n115,
         npu_inst_pe_1_4_4_n114, npu_inst_pe_1_4_4_n113,
         npu_inst_pe_1_4_4_n112, npu_inst_pe_1_4_4_n111,
         npu_inst_pe_1_4_4_n110, npu_inst_pe_1_4_4_n109,
         npu_inst_pe_1_4_4_n108, npu_inst_pe_1_4_4_n107,
         npu_inst_pe_1_4_4_n106, npu_inst_pe_1_4_4_n105,
         npu_inst_pe_1_4_4_n104, npu_inst_pe_1_4_4_n103,
         npu_inst_pe_1_4_4_n102, npu_inst_pe_1_4_4_n101,
         npu_inst_pe_1_4_4_n100, npu_inst_pe_1_4_4_n99, npu_inst_pe_1_4_4_n98,
         npu_inst_pe_1_4_4_n36, npu_inst_pe_1_4_4_n35, npu_inst_pe_1_4_4_n34,
         npu_inst_pe_1_4_4_n33, npu_inst_pe_1_4_4_n32, npu_inst_pe_1_4_4_n31,
         npu_inst_pe_1_4_4_n30, npu_inst_pe_1_4_4_n29, npu_inst_pe_1_4_4_n28,
         npu_inst_pe_1_4_4_n25, npu_inst_pe_1_4_4_n24, npu_inst_pe_1_4_4_n23,
         npu_inst_pe_1_4_4_n22, npu_inst_pe_1_4_4_n21, npu_inst_pe_1_4_4_n20,
         npu_inst_pe_1_4_4_n19, npu_inst_pe_1_4_4_n18, npu_inst_pe_1_4_4_n17,
         npu_inst_pe_1_4_4_n16, npu_inst_pe_1_4_4_n15, npu_inst_pe_1_4_4_n14,
         npu_inst_pe_1_4_4_n13, npu_inst_pe_1_4_4_n12, npu_inst_pe_1_4_4_n11,
         npu_inst_pe_1_4_4_n10, npu_inst_pe_1_4_4_n9, npu_inst_pe_1_4_4_n8,
         npu_inst_pe_1_4_4_n7, npu_inst_pe_1_4_4_n6, npu_inst_pe_1_4_4_n5,
         npu_inst_pe_1_4_4_n4, npu_inst_pe_1_4_4_n3, npu_inst_pe_1_4_4_n2,
         npu_inst_pe_1_4_4_n1, npu_inst_pe_1_4_4_sub_67_carry_7_,
         npu_inst_pe_1_4_4_sub_67_carry_6_, npu_inst_pe_1_4_4_sub_67_carry_5_,
         npu_inst_pe_1_4_4_sub_67_carry_4_, npu_inst_pe_1_4_4_sub_67_carry_3_,
         npu_inst_pe_1_4_4_sub_67_carry_2_, npu_inst_pe_1_4_4_sub_67_carry_1_,
         npu_inst_pe_1_4_4_add_69_carry_7_, npu_inst_pe_1_4_4_add_69_carry_6_,
         npu_inst_pe_1_4_4_add_69_carry_5_, npu_inst_pe_1_4_4_add_69_carry_4_,
         npu_inst_pe_1_4_4_add_69_carry_3_, npu_inst_pe_1_4_4_add_69_carry_2_,
         npu_inst_pe_1_4_4_add_69_carry_1_, npu_inst_pe_1_4_4_n97,
         npu_inst_pe_1_4_4_n96, npu_inst_pe_1_4_4_n95, npu_inst_pe_1_4_4_n94,
         npu_inst_pe_1_4_4_n93, npu_inst_pe_1_4_4_n92, npu_inst_pe_1_4_4_n91,
         npu_inst_pe_1_4_4_n90, npu_inst_pe_1_4_4_n89, npu_inst_pe_1_4_4_n88,
         npu_inst_pe_1_4_4_n87, npu_inst_pe_1_4_4_n86, npu_inst_pe_1_4_4_n85,
         npu_inst_pe_1_4_4_n84, npu_inst_pe_1_4_4_n83, npu_inst_pe_1_4_4_n82,
         npu_inst_pe_1_4_4_n81, npu_inst_pe_1_4_4_n80, npu_inst_pe_1_4_4_n79,
         npu_inst_pe_1_4_4_n78, npu_inst_pe_1_4_4_n77, npu_inst_pe_1_4_4_n76,
         npu_inst_pe_1_4_4_n75, npu_inst_pe_1_4_4_n74, npu_inst_pe_1_4_4_n73,
         npu_inst_pe_1_4_4_n72, npu_inst_pe_1_4_4_n71, npu_inst_pe_1_4_4_n70,
         npu_inst_pe_1_4_4_n69, npu_inst_pe_1_4_4_n68, npu_inst_pe_1_4_4_n67,
         npu_inst_pe_1_4_4_n66, npu_inst_pe_1_4_4_n65, npu_inst_pe_1_4_4_n64,
         npu_inst_pe_1_4_4_n63, npu_inst_pe_1_4_4_n62, npu_inst_pe_1_4_4_n61,
         npu_inst_pe_1_4_4_n60, npu_inst_pe_1_4_4_n59, npu_inst_pe_1_4_4_n58,
         npu_inst_pe_1_4_4_n57, npu_inst_pe_1_4_4_n56, npu_inst_pe_1_4_4_n55,
         npu_inst_pe_1_4_4_n54, npu_inst_pe_1_4_4_n53, npu_inst_pe_1_4_4_n52,
         npu_inst_pe_1_4_4_n51, npu_inst_pe_1_4_4_n50, npu_inst_pe_1_4_4_n49,
         npu_inst_pe_1_4_4_n48, npu_inst_pe_1_4_4_n47, npu_inst_pe_1_4_4_n46,
         npu_inst_pe_1_4_4_n45, npu_inst_pe_1_4_4_n44, npu_inst_pe_1_4_4_n43,
         npu_inst_pe_1_4_4_n42, npu_inst_pe_1_4_4_n41, npu_inst_pe_1_4_4_n40,
         npu_inst_pe_1_4_4_n39, npu_inst_pe_1_4_4_n38, npu_inst_pe_1_4_4_n37,
         npu_inst_pe_1_4_4_n27, npu_inst_pe_1_4_4_n26,
         npu_inst_pe_1_4_4_net3740, npu_inst_pe_1_4_4_net3734,
         npu_inst_pe_1_4_4_N94, npu_inst_pe_1_4_4_N93, npu_inst_pe_1_4_4_N84,
         npu_inst_pe_1_4_4_N80, npu_inst_pe_1_4_4_N79, npu_inst_pe_1_4_4_N78,
         npu_inst_pe_1_4_4_N77, npu_inst_pe_1_4_4_N76, npu_inst_pe_1_4_4_N75,
         npu_inst_pe_1_4_4_N74, npu_inst_pe_1_4_4_N73, npu_inst_pe_1_4_4_N72,
         npu_inst_pe_1_4_4_N71, npu_inst_pe_1_4_4_N70, npu_inst_pe_1_4_4_N69,
         npu_inst_pe_1_4_4_N68, npu_inst_pe_1_4_4_N67, npu_inst_pe_1_4_4_N66,
         npu_inst_pe_1_4_4_N65, npu_inst_pe_1_4_4_int_q_acc_0_,
         npu_inst_pe_1_4_4_int_q_acc_1_, npu_inst_pe_1_4_4_int_q_acc_2_,
         npu_inst_pe_1_4_4_int_q_acc_3_, npu_inst_pe_1_4_4_int_q_acc_4_,
         npu_inst_pe_1_4_4_int_q_acc_5_, npu_inst_pe_1_4_4_int_q_acc_6_,
         npu_inst_pe_1_4_4_int_q_acc_7_, npu_inst_pe_1_4_4_int_data_0_,
         npu_inst_pe_1_4_4_int_data_1_, npu_inst_pe_1_4_4_int_q_weight_0_,
         npu_inst_pe_1_4_4_int_q_weight_1_,
         npu_inst_pe_1_4_4_int_q_reg_v_5__0_,
         npu_inst_pe_1_4_4_int_q_reg_v_5__1_,
         npu_inst_pe_1_4_4_int_q_reg_v_4__0_,
         npu_inst_pe_1_4_4_int_q_reg_v_4__1_,
         npu_inst_pe_1_4_4_int_q_reg_v_3__0_,
         npu_inst_pe_1_4_4_int_q_reg_v_3__1_,
         npu_inst_pe_1_4_4_int_q_reg_v_2__0_,
         npu_inst_pe_1_4_4_int_q_reg_v_2__1_,
         npu_inst_pe_1_4_4_int_q_reg_v_1__0_,
         npu_inst_pe_1_4_4_int_q_reg_v_1__1_,
         npu_inst_pe_1_4_4_int_q_reg_v_0__0_,
         npu_inst_pe_1_4_4_int_q_reg_v_0__1_,
         npu_inst_pe_1_4_4_int_q_reg_h_5__0_,
         npu_inst_pe_1_4_4_int_q_reg_h_5__1_,
         npu_inst_pe_1_4_4_int_q_reg_h_4__0_,
         npu_inst_pe_1_4_4_int_q_reg_h_4__1_,
         npu_inst_pe_1_4_4_int_q_reg_h_3__0_,
         npu_inst_pe_1_4_4_int_q_reg_h_3__1_,
         npu_inst_pe_1_4_4_int_q_reg_h_2__0_,
         npu_inst_pe_1_4_4_int_q_reg_h_2__1_,
         npu_inst_pe_1_4_4_int_q_reg_h_1__0_,
         npu_inst_pe_1_4_4_int_q_reg_h_1__1_,
         npu_inst_pe_1_4_4_int_q_reg_h_0__0_,
         npu_inst_pe_1_4_4_int_q_reg_h_0__1_, npu_inst_pe_1_4_5_n119,
         npu_inst_pe_1_4_5_n118, npu_inst_pe_1_4_5_n117,
         npu_inst_pe_1_4_5_n116, npu_inst_pe_1_4_5_n115,
         npu_inst_pe_1_4_5_n114, npu_inst_pe_1_4_5_n113,
         npu_inst_pe_1_4_5_n112, npu_inst_pe_1_4_5_n111,
         npu_inst_pe_1_4_5_n110, npu_inst_pe_1_4_5_n109,
         npu_inst_pe_1_4_5_n108, npu_inst_pe_1_4_5_n107,
         npu_inst_pe_1_4_5_n106, npu_inst_pe_1_4_5_n105,
         npu_inst_pe_1_4_5_n104, npu_inst_pe_1_4_5_n103,
         npu_inst_pe_1_4_5_n102, npu_inst_pe_1_4_5_n101,
         npu_inst_pe_1_4_5_n100, npu_inst_pe_1_4_5_n99, npu_inst_pe_1_4_5_n98,
         npu_inst_pe_1_4_5_n36, npu_inst_pe_1_4_5_n35, npu_inst_pe_1_4_5_n34,
         npu_inst_pe_1_4_5_n33, npu_inst_pe_1_4_5_n32, npu_inst_pe_1_4_5_n31,
         npu_inst_pe_1_4_5_n30, npu_inst_pe_1_4_5_n29, npu_inst_pe_1_4_5_n28,
         npu_inst_pe_1_4_5_n25, npu_inst_pe_1_4_5_n24, npu_inst_pe_1_4_5_n23,
         npu_inst_pe_1_4_5_n22, npu_inst_pe_1_4_5_n21, npu_inst_pe_1_4_5_n20,
         npu_inst_pe_1_4_5_n19, npu_inst_pe_1_4_5_n18, npu_inst_pe_1_4_5_n17,
         npu_inst_pe_1_4_5_n16, npu_inst_pe_1_4_5_n15, npu_inst_pe_1_4_5_n14,
         npu_inst_pe_1_4_5_n13, npu_inst_pe_1_4_5_n12, npu_inst_pe_1_4_5_n11,
         npu_inst_pe_1_4_5_n10, npu_inst_pe_1_4_5_n9, npu_inst_pe_1_4_5_n8,
         npu_inst_pe_1_4_5_n7, npu_inst_pe_1_4_5_n6, npu_inst_pe_1_4_5_n5,
         npu_inst_pe_1_4_5_n4, npu_inst_pe_1_4_5_n3, npu_inst_pe_1_4_5_n2,
         npu_inst_pe_1_4_5_n1, npu_inst_pe_1_4_5_sub_67_carry_7_,
         npu_inst_pe_1_4_5_sub_67_carry_6_, npu_inst_pe_1_4_5_sub_67_carry_5_,
         npu_inst_pe_1_4_5_sub_67_carry_4_, npu_inst_pe_1_4_5_sub_67_carry_3_,
         npu_inst_pe_1_4_5_sub_67_carry_2_, npu_inst_pe_1_4_5_sub_67_carry_1_,
         npu_inst_pe_1_4_5_add_69_carry_7_, npu_inst_pe_1_4_5_add_69_carry_6_,
         npu_inst_pe_1_4_5_add_69_carry_5_, npu_inst_pe_1_4_5_add_69_carry_4_,
         npu_inst_pe_1_4_5_add_69_carry_3_, npu_inst_pe_1_4_5_add_69_carry_2_,
         npu_inst_pe_1_4_5_add_69_carry_1_, npu_inst_pe_1_4_5_n97,
         npu_inst_pe_1_4_5_n96, npu_inst_pe_1_4_5_n95, npu_inst_pe_1_4_5_n94,
         npu_inst_pe_1_4_5_n93, npu_inst_pe_1_4_5_n92, npu_inst_pe_1_4_5_n91,
         npu_inst_pe_1_4_5_n90, npu_inst_pe_1_4_5_n89, npu_inst_pe_1_4_5_n88,
         npu_inst_pe_1_4_5_n87, npu_inst_pe_1_4_5_n86, npu_inst_pe_1_4_5_n85,
         npu_inst_pe_1_4_5_n84, npu_inst_pe_1_4_5_n83, npu_inst_pe_1_4_5_n82,
         npu_inst_pe_1_4_5_n81, npu_inst_pe_1_4_5_n80, npu_inst_pe_1_4_5_n79,
         npu_inst_pe_1_4_5_n78, npu_inst_pe_1_4_5_n77, npu_inst_pe_1_4_5_n76,
         npu_inst_pe_1_4_5_n75, npu_inst_pe_1_4_5_n74, npu_inst_pe_1_4_5_n73,
         npu_inst_pe_1_4_5_n72, npu_inst_pe_1_4_5_n71, npu_inst_pe_1_4_5_n70,
         npu_inst_pe_1_4_5_n69, npu_inst_pe_1_4_5_n68, npu_inst_pe_1_4_5_n67,
         npu_inst_pe_1_4_5_n66, npu_inst_pe_1_4_5_n65, npu_inst_pe_1_4_5_n64,
         npu_inst_pe_1_4_5_n63, npu_inst_pe_1_4_5_n62, npu_inst_pe_1_4_5_n61,
         npu_inst_pe_1_4_5_n60, npu_inst_pe_1_4_5_n59, npu_inst_pe_1_4_5_n58,
         npu_inst_pe_1_4_5_n57, npu_inst_pe_1_4_5_n56, npu_inst_pe_1_4_5_n55,
         npu_inst_pe_1_4_5_n54, npu_inst_pe_1_4_5_n53, npu_inst_pe_1_4_5_n52,
         npu_inst_pe_1_4_5_n51, npu_inst_pe_1_4_5_n50, npu_inst_pe_1_4_5_n49,
         npu_inst_pe_1_4_5_n48, npu_inst_pe_1_4_5_n47, npu_inst_pe_1_4_5_n46,
         npu_inst_pe_1_4_5_n45, npu_inst_pe_1_4_5_n44, npu_inst_pe_1_4_5_n43,
         npu_inst_pe_1_4_5_n42, npu_inst_pe_1_4_5_n41, npu_inst_pe_1_4_5_n40,
         npu_inst_pe_1_4_5_n39, npu_inst_pe_1_4_5_n38, npu_inst_pe_1_4_5_n37,
         npu_inst_pe_1_4_5_n27, npu_inst_pe_1_4_5_n26,
         npu_inst_pe_1_4_5_net3717, npu_inst_pe_1_4_5_net3711,
         npu_inst_pe_1_4_5_N94, npu_inst_pe_1_4_5_N93, npu_inst_pe_1_4_5_N84,
         npu_inst_pe_1_4_5_N80, npu_inst_pe_1_4_5_N79, npu_inst_pe_1_4_5_N78,
         npu_inst_pe_1_4_5_N77, npu_inst_pe_1_4_5_N76, npu_inst_pe_1_4_5_N75,
         npu_inst_pe_1_4_5_N74, npu_inst_pe_1_4_5_N73, npu_inst_pe_1_4_5_N72,
         npu_inst_pe_1_4_5_N71, npu_inst_pe_1_4_5_N70, npu_inst_pe_1_4_5_N69,
         npu_inst_pe_1_4_5_N68, npu_inst_pe_1_4_5_N67, npu_inst_pe_1_4_5_N66,
         npu_inst_pe_1_4_5_N65, npu_inst_pe_1_4_5_int_q_acc_0_,
         npu_inst_pe_1_4_5_int_q_acc_1_, npu_inst_pe_1_4_5_int_q_acc_2_,
         npu_inst_pe_1_4_5_int_q_acc_3_, npu_inst_pe_1_4_5_int_q_acc_4_,
         npu_inst_pe_1_4_5_int_q_acc_5_, npu_inst_pe_1_4_5_int_q_acc_6_,
         npu_inst_pe_1_4_5_int_q_acc_7_, npu_inst_pe_1_4_5_int_data_0_,
         npu_inst_pe_1_4_5_int_data_1_, npu_inst_pe_1_4_5_int_q_weight_0_,
         npu_inst_pe_1_4_5_int_q_weight_1_,
         npu_inst_pe_1_4_5_int_q_reg_v_5__0_,
         npu_inst_pe_1_4_5_int_q_reg_v_5__1_,
         npu_inst_pe_1_4_5_int_q_reg_v_4__0_,
         npu_inst_pe_1_4_5_int_q_reg_v_4__1_,
         npu_inst_pe_1_4_5_int_q_reg_v_3__0_,
         npu_inst_pe_1_4_5_int_q_reg_v_3__1_,
         npu_inst_pe_1_4_5_int_q_reg_v_2__0_,
         npu_inst_pe_1_4_5_int_q_reg_v_2__1_,
         npu_inst_pe_1_4_5_int_q_reg_v_1__0_,
         npu_inst_pe_1_4_5_int_q_reg_v_1__1_,
         npu_inst_pe_1_4_5_int_q_reg_v_0__0_,
         npu_inst_pe_1_4_5_int_q_reg_v_0__1_,
         npu_inst_pe_1_4_5_int_q_reg_h_5__0_,
         npu_inst_pe_1_4_5_int_q_reg_h_5__1_,
         npu_inst_pe_1_4_5_int_q_reg_h_4__0_,
         npu_inst_pe_1_4_5_int_q_reg_h_4__1_,
         npu_inst_pe_1_4_5_int_q_reg_h_3__0_,
         npu_inst_pe_1_4_5_int_q_reg_h_3__1_,
         npu_inst_pe_1_4_5_int_q_reg_h_2__0_,
         npu_inst_pe_1_4_5_int_q_reg_h_2__1_,
         npu_inst_pe_1_4_5_int_q_reg_h_1__0_,
         npu_inst_pe_1_4_5_int_q_reg_h_1__1_,
         npu_inst_pe_1_4_5_int_q_reg_h_0__0_,
         npu_inst_pe_1_4_5_int_q_reg_h_0__1_, npu_inst_pe_1_4_6_n119,
         npu_inst_pe_1_4_6_n118, npu_inst_pe_1_4_6_n117,
         npu_inst_pe_1_4_6_n116, npu_inst_pe_1_4_6_n115,
         npu_inst_pe_1_4_6_n114, npu_inst_pe_1_4_6_n113,
         npu_inst_pe_1_4_6_n112, npu_inst_pe_1_4_6_n111,
         npu_inst_pe_1_4_6_n110, npu_inst_pe_1_4_6_n109,
         npu_inst_pe_1_4_6_n108, npu_inst_pe_1_4_6_n107,
         npu_inst_pe_1_4_6_n106, npu_inst_pe_1_4_6_n105,
         npu_inst_pe_1_4_6_n104, npu_inst_pe_1_4_6_n103,
         npu_inst_pe_1_4_6_n102, npu_inst_pe_1_4_6_n101,
         npu_inst_pe_1_4_6_n100, npu_inst_pe_1_4_6_n99, npu_inst_pe_1_4_6_n98,
         npu_inst_pe_1_4_6_n36, npu_inst_pe_1_4_6_n35, npu_inst_pe_1_4_6_n34,
         npu_inst_pe_1_4_6_n33, npu_inst_pe_1_4_6_n32, npu_inst_pe_1_4_6_n31,
         npu_inst_pe_1_4_6_n30, npu_inst_pe_1_4_6_n29, npu_inst_pe_1_4_6_n28,
         npu_inst_pe_1_4_6_n25, npu_inst_pe_1_4_6_n24, npu_inst_pe_1_4_6_n23,
         npu_inst_pe_1_4_6_n22, npu_inst_pe_1_4_6_n21, npu_inst_pe_1_4_6_n20,
         npu_inst_pe_1_4_6_n19, npu_inst_pe_1_4_6_n18, npu_inst_pe_1_4_6_n17,
         npu_inst_pe_1_4_6_n16, npu_inst_pe_1_4_6_n15, npu_inst_pe_1_4_6_n14,
         npu_inst_pe_1_4_6_n13, npu_inst_pe_1_4_6_n12, npu_inst_pe_1_4_6_n11,
         npu_inst_pe_1_4_6_n10, npu_inst_pe_1_4_6_n9, npu_inst_pe_1_4_6_n8,
         npu_inst_pe_1_4_6_n7, npu_inst_pe_1_4_6_n6, npu_inst_pe_1_4_6_n5,
         npu_inst_pe_1_4_6_n4, npu_inst_pe_1_4_6_n3, npu_inst_pe_1_4_6_n2,
         npu_inst_pe_1_4_6_n1, npu_inst_pe_1_4_6_sub_67_carry_7_,
         npu_inst_pe_1_4_6_sub_67_carry_6_, npu_inst_pe_1_4_6_sub_67_carry_5_,
         npu_inst_pe_1_4_6_sub_67_carry_4_, npu_inst_pe_1_4_6_sub_67_carry_3_,
         npu_inst_pe_1_4_6_sub_67_carry_2_, npu_inst_pe_1_4_6_sub_67_carry_1_,
         npu_inst_pe_1_4_6_add_69_carry_7_, npu_inst_pe_1_4_6_add_69_carry_6_,
         npu_inst_pe_1_4_6_add_69_carry_5_, npu_inst_pe_1_4_6_add_69_carry_4_,
         npu_inst_pe_1_4_6_add_69_carry_3_, npu_inst_pe_1_4_6_add_69_carry_2_,
         npu_inst_pe_1_4_6_add_69_carry_1_, npu_inst_pe_1_4_6_n97,
         npu_inst_pe_1_4_6_n96, npu_inst_pe_1_4_6_n95, npu_inst_pe_1_4_6_n94,
         npu_inst_pe_1_4_6_n93, npu_inst_pe_1_4_6_n92, npu_inst_pe_1_4_6_n91,
         npu_inst_pe_1_4_6_n90, npu_inst_pe_1_4_6_n89, npu_inst_pe_1_4_6_n88,
         npu_inst_pe_1_4_6_n87, npu_inst_pe_1_4_6_n86, npu_inst_pe_1_4_6_n85,
         npu_inst_pe_1_4_6_n84, npu_inst_pe_1_4_6_n83, npu_inst_pe_1_4_6_n82,
         npu_inst_pe_1_4_6_n81, npu_inst_pe_1_4_6_n80, npu_inst_pe_1_4_6_n79,
         npu_inst_pe_1_4_6_n78, npu_inst_pe_1_4_6_n77, npu_inst_pe_1_4_6_n76,
         npu_inst_pe_1_4_6_n75, npu_inst_pe_1_4_6_n74, npu_inst_pe_1_4_6_n73,
         npu_inst_pe_1_4_6_n72, npu_inst_pe_1_4_6_n71, npu_inst_pe_1_4_6_n70,
         npu_inst_pe_1_4_6_n69, npu_inst_pe_1_4_6_n68, npu_inst_pe_1_4_6_n67,
         npu_inst_pe_1_4_6_n66, npu_inst_pe_1_4_6_n65, npu_inst_pe_1_4_6_n64,
         npu_inst_pe_1_4_6_n63, npu_inst_pe_1_4_6_n62, npu_inst_pe_1_4_6_n61,
         npu_inst_pe_1_4_6_n60, npu_inst_pe_1_4_6_n59, npu_inst_pe_1_4_6_n58,
         npu_inst_pe_1_4_6_n57, npu_inst_pe_1_4_6_n56, npu_inst_pe_1_4_6_n55,
         npu_inst_pe_1_4_6_n54, npu_inst_pe_1_4_6_n53, npu_inst_pe_1_4_6_n52,
         npu_inst_pe_1_4_6_n51, npu_inst_pe_1_4_6_n50, npu_inst_pe_1_4_6_n49,
         npu_inst_pe_1_4_6_n48, npu_inst_pe_1_4_6_n47, npu_inst_pe_1_4_6_n46,
         npu_inst_pe_1_4_6_n45, npu_inst_pe_1_4_6_n44, npu_inst_pe_1_4_6_n43,
         npu_inst_pe_1_4_6_n42, npu_inst_pe_1_4_6_n41, npu_inst_pe_1_4_6_n40,
         npu_inst_pe_1_4_6_n39, npu_inst_pe_1_4_6_n38, npu_inst_pe_1_4_6_n37,
         npu_inst_pe_1_4_6_n27, npu_inst_pe_1_4_6_n26,
         npu_inst_pe_1_4_6_net3694, npu_inst_pe_1_4_6_net3688,
         npu_inst_pe_1_4_6_N94, npu_inst_pe_1_4_6_N93, npu_inst_pe_1_4_6_N84,
         npu_inst_pe_1_4_6_N80, npu_inst_pe_1_4_6_N79, npu_inst_pe_1_4_6_N78,
         npu_inst_pe_1_4_6_N77, npu_inst_pe_1_4_6_N76, npu_inst_pe_1_4_6_N75,
         npu_inst_pe_1_4_6_N74, npu_inst_pe_1_4_6_N73, npu_inst_pe_1_4_6_N72,
         npu_inst_pe_1_4_6_N71, npu_inst_pe_1_4_6_N70, npu_inst_pe_1_4_6_N69,
         npu_inst_pe_1_4_6_N68, npu_inst_pe_1_4_6_N67, npu_inst_pe_1_4_6_N66,
         npu_inst_pe_1_4_6_N65, npu_inst_pe_1_4_6_int_q_acc_0_,
         npu_inst_pe_1_4_6_int_q_acc_1_, npu_inst_pe_1_4_6_int_q_acc_2_,
         npu_inst_pe_1_4_6_int_q_acc_3_, npu_inst_pe_1_4_6_int_q_acc_4_,
         npu_inst_pe_1_4_6_int_q_acc_5_, npu_inst_pe_1_4_6_int_q_acc_6_,
         npu_inst_pe_1_4_6_int_q_acc_7_, npu_inst_pe_1_4_6_int_data_0_,
         npu_inst_pe_1_4_6_int_data_1_, npu_inst_pe_1_4_6_int_q_weight_0_,
         npu_inst_pe_1_4_6_int_q_weight_1_,
         npu_inst_pe_1_4_6_int_q_reg_v_5__0_,
         npu_inst_pe_1_4_6_int_q_reg_v_5__1_,
         npu_inst_pe_1_4_6_int_q_reg_v_4__0_,
         npu_inst_pe_1_4_6_int_q_reg_v_4__1_,
         npu_inst_pe_1_4_6_int_q_reg_v_3__0_,
         npu_inst_pe_1_4_6_int_q_reg_v_3__1_,
         npu_inst_pe_1_4_6_int_q_reg_v_2__0_,
         npu_inst_pe_1_4_6_int_q_reg_v_2__1_,
         npu_inst_pe_1_4_6_int_q_reg_v_1__0_,
         npu_inst_pe_1_4_6_int_q_reg_v_1__1_,
         npu_inst_pe_1_4_6_int_q_reg_v_0__0_,
         npu_inst_pe_1_4_6_int_q_reg_v_0__1_,
         npu_inst_pe_1_4_6_int_q_reg_h_5__0_,
         npu_inst_pe_1_4_6_int_q_reg_h_5__1_,
         npu_inst_pe_1_4_6_int_q_reg_h_4__0_,
         npu_inst_pe_1_4_6_int_q_reg_h_4__1_,
         npu_inst_pe_1_4_6_int_q_reg_h_3__0_,
         npu_inst_pe_1_4_6_int_q_reg_h_3__1_,
         npu_inst_pe_1_4_6_int_q_reg_h_2__0_,
         npu_inst_pe_1_4_6_int_q_reg_h_2__1_,
         npu_inst_pe_1_4_6_int_q_reg_h_1__0_,
         npu_inst_pe_1_4_6_int_q_reg_h_1__1_,
         npu_inst_pe_1_4_6_int_q_reg_h_0__0_,
         npu_inst_pe_1_4_6_int_q_reg_h_0__1_, npu_inst_pe_1_4_7_n119,
         npu_inst_pe_1_4_7_n118, npu_inst_pe_1_4_7_n117,
         npu_inst_pe_1_4_7_n116, npu_inst_pe_1_4_7_n115,
         npu_inst_pe_1_4_7_n114, npu_inst_pe_1_4_7_n113,
         npu_inst_pe_1_4_7_n112, npu_inst_pe_1_4_7_n111,
         npu_inst_pe_1_4_7_n110, npu_inst_pe_1_4_7_n109,
         npu_inst_pe_1_4_7_n108, npu_inst_pe_1_4_7_n107,
         npu_inst_pe_1_4_7_n106, npu_inst_pe_1_4_7_n105,
         npu_inst_pe_1_4_7_n104, npu_inst_pe_1_4_7_n103,
         npu_inst_pe_1_4_7_n102, npu_inst_pe_1_4_7_n101,
         npu_inst_pe_1_4_7_n100, npu_inst_pe_1_4_7_n99, npu_inst_pe_1_4_7_n98,
         npu_inst_pe_1_4_7_n36, npu_inst_pe_1_4_7_n35, npu_inst_pe_1_4_7_n34,
         npu_inst_pe_1_4_7_n33, npu_inst_pe_1_4_7_n32, npu_inst_pe_1_4_7_n31,
         npu_inst_pe_1_4_7_n30, npu_inst_pe_1_4_7_n29, npu_inst_pe_1_4_7_n28,
         npu_inst_pe_1_4_7_n25, npu_inst_pe_1_4_7_n24, npu_inst_pe_1_4_7_n23,
         npu_inst_pe_1_4_7_n22, npu_inst_pe_1_4_7_n21, npu_inst_pe_1_4_7_n20,
         npu_inst_pe_1_4_7_n19, npu_inst_pe_1_4_7_n18, npu_inst_pe_1_4_7_n17,
         npu_inst_pe_1_4_7_n16, npu_inst_pe_1_4_7_n15, npu_inst_pe_1_4_7_n14,
         npu_inst_pe_1_4_7_n13, npu_inst_pe_1_4_7_n12, npu_inst_pe_1_4_7_n11,
         npu_inst_pe_1_4_7_n10, npu_inst_pe_1_4_7_n9, npu_inst_pe_1_4_7_n8,
         npu_inst_pe_1_4_7_n7, npu_inst_pe_1_4_7_n6, npu_inst_pe_1_4_7_n5,
         npu_inst_pe_1_4_7_n4, npu_inst_pe_1_4_7_n3, npu_inst_pe_1_4_7_n2,
         npu_inst_pe_1_4_7_n1, npu_inst_pe_1_4_7_sub_67_carry_7_,
         npu_inst_pe_1_4_7_sub_67_carry_6_, npu_inst_pe_1_4_7_sub_67_carry_5_,
         npu_inst_pe_1_4_7_sub_67_carry_4_, npu_inst_pe_1_4_7_sub_67_carry_3_,
         npu_inst_pe_1_4_7_sub_67_carry_2_, npu_inst_pe_1_4_7_sub_67_carry_1_,
         npu_inst_pe_1_4_7_add_69_carry_7_, npu_inst_pe_1_4_7_add_69_carry_6_,
         npu_inst_pe_1_4_7_add_69_carry_5_, npu_inst_pe_1_4_7_add_69_carry_4_,
         npu_inst_pe_1_4_7_add_69_carry_3_, npu_inst_pe_1_4_7_add_69_carry_2_,
         npu_inst_pe_1_4_7_add_69_carry_1_, npu_inst_pe_1_4_7_n97,
         npu_inst_pe_1_4_7_n96, npu_inst_pe_1_4_7_n95, npu_inst_pe_1_4_7_n94,
         npu_inst_pe_1_4_7_n93, npu_inst_pe_1_4_7_n92, npu_inst_pe_1_4_7_n91,
         npu_inst_pe_1_4_7_n90, npu_inst_pe_1_4_7_n89, npu_inst_pe_1_4_7_n88,
         npu_inst_pe_1_4_7_n87, npu_inst_pe_1_4_7_n86, npu_inst_pe_1_4_7_n85,
         npu_inst_pe_1_4_7_n84, npu_inst_pe_1_4_7_n83, npu_inst_pe_1_4_7_n82,
         npu_inst_pe_1_4_7_n81, npu_inst_pe_1_4_7_n80, npu_inst_pe_1_4_7_n79,
         npu_inst_pe_1_4_7_n78, npu_inst_pe_1_4_7_n77, npu_inst_pe_1_4_7_n76,
         npu_inst_pe_1_4_7_n75, npu_inst_pe_1_4_7_n74, npu_inst_pe_1_4_7_n73,
         npu_inst_pe_1_4_7_n72, npu_inst_pe_1_4_7_n71, npu_inst_pe_1_4_7_n70,
         npu_inst_pe_1_4_7_n69, npu_inst_pe_1_4_7_n68, npu_inst_pe_1_4_7_n67,
         npu_inst_pe_1_4_7_n66, npu_inst_pe_1_4_7_n65, npu_inst_pe_1_4_7_n64,
         npu_inst_pe_1_4_7_n63, npu_inst_pe_1_4_7_n62, npu_inst_pe_1_4_7_n61,
         npu_inst_pe_1_4_7_n60, npu_inst_pe_1_4_7_n59, npu_inst_pe_1_4_7_n58,
         npu_inst_pe_1_4_7_n57, npu_inst_pe_1_4_7_n56, npu_inst_pe_1_4_7_n55,
         npu_inst_pe_1_4_7_n54, npu_inst_pe_1_4_7_n53, npu_inst_pe_1_4_7_n52,
         npu_inst_pe_1_4_7_n51, npu_inst_pe_1_4_7_n50, npu_inst_pe_1_4_7_n49,
         npu_inst_pe_1_4_7_n48, npu_inst_pe_1_4_7_n47, npu_inst_pe_1_4_7_n46,
         npu_inst_pe_1_4_7_n45, npu_inst_pe_1_4_7_n44, npu_inst_pe_1_4_7_n43,
         npu_inst_pe_1_4_7_n42, npu_inst_pe_1_4_7_n41, npu_inst_pe_1_4_7_n40,
         npu_inst_pe_1_4_7_n39, npu_inst_pe_1_4_7_n38, npu_inst_pe_1_4_7_n37,
         npu_inst_pe_1_4_7_n27, npu_inst_pe_1_4_7_n26,
         npu_inst_pe_1_4_7_net3671, npu_inst_pe_1_4_7_net3665,
         npu_inst_pe_1_4_7_N94, npu_inst_pe_1_4_7_N93, npu_inst_pe_1_4_7_N84,
         npu_inst_pe_1_4_7_N80, npu_inst_pe_1_4_7_N79, npu_inst_pe_1_4_7_N78,
         npu_inst_pe_1_4_7_N77, npu_inst_pe_1_4_7_N76, npu_inst_pe_1_4_7_N75,
         npu_inst_pe_1_4_7_N74, npu_inst_pe_1_4_7_N73, npu_inst_pe_1_4_7_N72,
         npu_inst_pe_1_4_7_N71, npu_inst_pe_1_4_7_N70, npu_inst_pe_1_4_7_N69,
         npu_inst_pe_1_4_7_N68, npu_inst_pe_1_4_7_N67, npu_inst_pe_1_4_7_N66,
         npu_inst_pe_1_4_7_N65, npu_inst_pe_1_4_7_int_q_acc_0_,
         npu_inst_pe_1_4_7_int_q_acc_1_, npu_inst_pe_1_4_7_int_q_acc_2_,
         npu_inst_pe_1_4_7_int_q_acc_3_, npu_inst_pe_1_4_7_int_q_acc_4_,
         npu_inst_pe_1_4_7_int_q_acc_5_, npu_inst_pe_1_4_7_int_q_acc_6_,
         npu_inst_pe_1_4_7_int_q_acc_7_, npu_inst_pe_1_4_7_int_data_0_,
         npu_inst_pe_1_4_7_int_data_1_, npu_inst_pe_1_4_7_int_q_weight_0_,
         npu_inst_pe_1_4_7_int_q_weight_1_,
         npu_inst_pe_1_4_7_int_q_reg_v_5__0_,
         npu_inst_pe_1_4_7_int_q_reg_v_5__1_,
         npu_inst_pe_1_4_7_int_q_reg_v_4__0_,
         npu_inst_pe_1_4_7_int_q_reg_v_4__1_,
         npu_inst_pe_1_4_7_int_q_reg_v_3__0_,
         npu_inst_pe_1_4_7_int_q_reg_v_3__1_,
         npu_inst_pe_1_4_7_int_q_reg_v_2__0_,
         npu_inst_pe_1_4_7_int_q_reg_v_2__1_,
         npu_inst_pe_1_4_7_int_q_reg_v_1__0_,
         npu_inst_pe_1_4_7_int_q_reg_v_1__1_,
         npu_inst_pe_1_4_7_int_q_reg_v_0__0_,
         npu_inst_pe_1_4_7_int_q_reg_v_0__1_,
         npu_inst_pe_1_4_7_int_q_reg_h_5__0_,
         npu_inst_pe_1_4_7_int_q_reg_h_5__1_,
         npu_inst_pe_1_4_7_int_q_reg_h_4__0_,
         npu_inst_pe_1_4_7_int_q_reg_h_4__1_,
         npu_inst_pe_1_4_7_int_q_reg_h_3__0_,
         npu_inst_pe_1_4_7_int_q_reg_h_3__1_,
         npu_inst_pe_1_4_7_int_q_reg_h_2__0_,
         npu_inst_pe_1_4_7_int_q_reg_h_2__1_,
         npu_inst_pe_1_4_7_int_q_reg_h_1__0_,
         npu_inst_pe_1_4_7_int_q_reg_h_1__1_,
         npu_inst_pe_1_4_7_int_q_reg_h_0__0_,
         npu_inst_pe_1_4_7_int_q_reg_h_0__1_, npu_inst_pe_1_5_0_n118,
         npu_inst_pe_1_5_0_n117, npu_inst_pe_1_5_0_n116,
         npu_inst_pe_1_5_0_n115, npu_inst_pe_1_5_0_n114,
         npu_inst_pe_1_5_0_n113, npu_inst_pe_1_5_0_n112,
         npu_inst_pe_1_5_0_n111, npu_inst_pe_1_5_0_n110,
         npu_inst_pe_1_5_0_n109, npu_inst_pe_1_5_0_n108,
         npu_inst_pe_1_5_0_n107, npu_inst_pe_1_5_0_n106,
         npu_inst_pe_1_5_0_n105, npu_inst_pe_1_5_0_n104,
         npu_inst_pe_1_5_0_n103, npu_inst_pe_1_5_0_n102,
         npu_inst_pe_1_5_0_n101, npu_inst_pe_1_5_0_n100, npu_inst_pe_1_5_0_n99,
         npu_inst_pe_1_5_0_n98, npu_inst_pe_1_5_0_n36, npu_inst_pe_1_5_0_n35,
         npu_inst_pe_1_5_0_n34, npu_inst_pe_1_5_0_n33, npu_inst_pe_1_5_0_n32,
         npu_inst_pe_1_5_0_n31, npu_inst_pe_1_5_0_n30, npu_inst_pe_1_5_0_n29,
         npu_inst_pe_1_5_0_n28, npu_inst_pe_1_5_0_n25, npu_inst_pe_1_5_0_n24,
         npu_inst_pe_1_5_0_n23, npu_inst_pe_1_5_0_n22, npu_inst_pe_1_5_0_n21,
         npu_inst_pe_1_5_0_n20, npu_inst_pe_1_5_0_n19, npu_inst_pe_1_5_0_n18,
         npu_inst_pe_1_5_0_n17, npu_inst_pe_1_5_0_n16, npu_inst_pe_1_5_0_n15,
         npu_inst_pe_1_5_0_n14, npu_inst_pe_1_5_0_n13, npu_inst_pe_1_5_0_n12,
         npu_inst_pe_1_5_0_n11, npu_inst_pe_1_5_0_n10, npu_inst_pe_1_5_0_n9,
         npu_inst_pe_1_5_0_n8, npu_inst_pe_1_5_0_n7, npu_inst_pe_1_5_0_n6,
         npu_inst_pe_1_5_0_n5, npu_inst_pe_1_5_0_n4, npu_inst_pe_1_5_0_n3,
         npu_inst_pe_1_5_0_n2, npu_inst_pe_1_5_0_n1,
         npu_inst_pe_1_5_0_sub_67_carry_7_, npu_inst_pe_1_5_0_sub_67_carry_6_,
         npu_inst_pe_1_5_0_sub_67_carry_5_, npu_inst_pe_1_5_0_sub_67_carry_4_,
         npu_inst_pe_1_5_0_sub_67_carry_3_, npu_inst_pe_1_5_0_sub_67_carry_2_,
         npu_inst_pe_1_5_0_sub_67_carry_1_, npu_inst_pe_1_5_0_add_69_carry_7_,
         npu_inst_pe_1_5_0_add_69_carry_6_, npu_inst_pe_1_5_0_add_69_carry_5_,
         npu_inst_pe_1_5_0_add_69_carry_4_, npu_inst_pe_1_5_0_add_69_carry_3_,
         npu_inst_pe_1_5_0_add_69_carry_2_, npu_inst_pe_1_5_0_add_69_carry_1_,
         npu_inst_pe_1_5_0_n97, npu_inst_pe_1_5_0_n96, npu_inst_pe_1_5_0_n95,
         npu_inst_pe_1_5_0_n94, npu_inst_pe_1_5_0_n93, npu_inst_pe_1_5_0_n92,
         npu_inst_pe_1_5_0_n91, npu_inst_pe_1_5_0_n90, npu_inst_pe_1_5_0_n89,
         npu_inst_pe_1_5_0_n88, npu_inst_pe_1_5_0_n87, npu_inst_pe_1_5_0_n86,
         npu_inst_pe_1_5_0_n85, npu_inst_pe_1_5_0_n84, npu_inst_pe_1_5_0_n83,
         npu_inst_pe_1_5_0_n82, npu_inst_pe_1_5_0_n81, npu_inst_pe_1_5_0_n80,
         npu_inst_pe_1_5_0_n79, npu_inst_pe_1_5_0_n78, npu_inst_pe_1_5_0_n77,
         npu_inst_pe_1_5_0_n76, npu_inst_pe_1_5_0_n75, npu_inst_pe_1_5_0_n74,
         npu_inst_pe_1_5_0_n73, npu_inst_pe_1_5_0_n72, npu_inst_pe_1_5_0_n71,
         npu_inst_pe_1_5_0_n70, npu_inst_pe_1_5_0_n69, npu_inst_pe_1_5_0_n68,
         npu_inst_pe_1_5_0_n67, npu_inst_pe_1_5_0_n66, npu_inst_pe_1_5_0_n65,
         npu_inst_pe_1_5_0_n64, npu_inst_pe_1_5_0_n63, npu_inst_pe_1_5_0_n62,
         npu_inst_pe_1_5_0_n61, npu_inst_pe_1_5_0_n60, npu_inst_pe_1_5_0_n59,
         npu_inst_pe_1_5_0_n58, npu_inst_pe_1_5_0_n57, npu_inst_pe_1_5_0_n56,
         npu_inst_pe_1_5_0_n55, npu_inst_pe_1_5_0_n54, npu_inst_pe_1_5_0_n53,
         npu_inst_pe_1_5_0_n52, npu_inst_pe_1_5_0_n51, npu_inst_pe_1_5_0_n50,
         npu_inst_pe_1_5_0_n49, npu_inst_pe_1_5_0_n48, npu_inst_pe_1_5_0_n47,
         npu_inst_pe_1_5_0_n46, npu_inst_pe_1_5_0_n45, npu_inst_pe_1_5_0_n44,
         npu_inst_pe_1_5_0_n43, npu_inst_pe_1_5_0_n42, npu_inst_pe_1_5_0_n41,
         npu_inst_pe_1_5_0_n40, npu_inst_pe_1_5_0_n39, npu_inst_pe_1_5_0_n38,
         npu_inst_pe_1_5_0_n37, npu_inst_pe_1_5_0_n27, npu_inst_pe_1_5_0_n26,
         npu_inst_pe_1_5_0_net3648, npu_inst_pe_1_5_0_net3642,
         npu_inst_pe_1_5_0_N94, npu_inst_pe_1_5_0_N93, npu_inst_pe_1_5_0_N84,
         npu_inst_pe_1_5_0_N80, npu_inst_pe_1_5_0_N79, npu_inst_pe_1_5_0_N78,
         npu_inst_pe_1_5_0_N77, npu_inst_pe_1_5_0_N76, npu_inst_pe_1_5_0_N75,
         npu_inst_pe_1_5_0_N74, npu_inst_pe_1_5_0_N73, npu_inst_pe_1_5_0_N72,
         npu_inst_pe_1_5_0_N71, npu_inst_pe_1_5_0_N70, npu_inst_pe_1_5_0_N69,
         npu_inst_pe_1_5_0_N68, npu_inst_pe_1_5_0_N67, npu_inst_pe_1_5_0_N66,
         npu_inst_pe_1_5_0_N65, npu_inst_pe_1_5_0_int_q_acc_0_,
         npu_inst_pe_1_5_0_int_q_acc_1_, npu_inst_pe_1_5_0_int_q_acc_2_,
         npu_inst_pe_1_5_0_int_q_acc_3_, npu_inst_pe_1_5_0_int_q_acc_4_,
         npu_inst_pe_1_5_0_int_q_acc_5_, npu_inst_pe_1_5_0_int_q_acc_6_,
         npu_inst_pe_1_5_0_int_q_acc_7_, npu_inst_pe_1_5_0_int_data_0_,
         npu_inst_pe_1_5_0_int_data_1_, npu_inst_pe_1_5_0_int_q_weight_0_,
         npu_inst_pe_1_5_0_int_q_weight_1_,
         npu_inst_pe_1_5_0_int_q_reg_v_5__0_,
         npu_inst_pe_1_5_0_int_q_reg_v_5__1_,
         npu_inst_pe_1_5_0_int_q_reg_v_4__0_,
         npu_inst_pe_1_5_0_int_q_reg_v_4__1_,
         npu_inst_pe_1_5_0_int_q_reg_v_3__0_,
         npu_inst_pe_1_5_0_int_q_reg_v_3__1_,
         npu_inst_pe_1_5_0_int_q_reg_v_2__0_,
         npu_inst_pe_1_5_0_int_q_reg_v_2__1_,
         npu_inst_pe_1_5_0_int_q_reg_v_1__0_,
         npu_inst_pe_1_5_0_int_q_reg_v_1__1_,
         npu_inst_pe_1_5_0_int_q_reg_v_0__0_,
         npu_inst_pe_1_5_0_int_q_reg_v_0__1_,
         npu_inst_pe_1_5_0_int_q_reg_h_5__0_,
         npu_inst_pe_1_5_0_int_q_reg_h_5__1_,
         npu_inst_pe_1_5_0_int_q_reg_h_4__0_,
         npu_inst_pe_1_5_0_int_q_reg_h_4__1_,
         npu_inst_pe_1_5_0_int_q_reg_h_3__0_,
         npu_inst_pe_1_5_0_int_q_reg_h_3__1_,
         npu_inst_pe_1_5_0_int_q_reg_h_2__0_,
         npu_inst_pe_1_5_0_int_q_reg_h_2__1_,
         npu_inst_pe_1_5_0_int_q_reg_h_1__0_,
         npu_inst_pe_1_5_0_int_q_reg_h_1__1_,
         npu_inst_pe_1_5_0_int_q_reg_h_0__0_,
         npu_inst_pe_1_5_0_int_q_reg_h_0__1_, npu_inst_pe_1_5_0_o_data_h_0_,
         npu_inst_pe_1_5_0_o_data_h_1_, npu_inst_pe_1_5_1_n119,
         npu_inst_pe_1_5_1_n118, npu_inst_pe_1_5_1_n117,
         npu_inst_pe_1_5_1_n116, npu_inst_pe_1_5_1_n115,
         npu_inst_pe_1_5_1_n114, npu_inst_pe_1_5_1_n113,
         npu_inst_pe_1_5_1_n112, npu_inst_pe_1_5_1_n111,
         npu_inst_pe_1_5_1_n110, npu_inst_pe_1_5_1_n109,
         npu_inst_pe_1_5_1_n108, npu_inst_pe_1_5_1_n107,
         npu_inst_pe_1_5_1_n106, npu_inst_pe_1_5_1_n105,
         npu_inst_pe_1_5_1_n104, npu_inst_pe_1_5_1_n103,
         npu_inst_pe_1_5_1_n102, npu_inst_pe_1_5_1_n101,
         npu_inst_pe_1_5_1_n100, npu_inst_pe_1_5_1_n99, npu_inst_pe_1_5_1_n98,
         npu_inst_pe_1_5_1_n36, npu_inst_pe_1_5_1_n35, npu_inst_pe_1_5_1_n34,
         npu_inst_pe_1_5_1_n33, npu_inst_pe_1_5_1_n32, npu_inst_pe_1_5_1_n31,
         npu_inst_pe_1_5_1_n30, npu_inst_pe_1_5_1_n29, npu_inst_pe_1_5_1_n28,
         npu_inst_pe_1_5_1_n25, npu_inst_pe_1_5_1_n24, npu_inst_pe_1_5_1_n23,
         npu_inst_pe_1_5_1_n22, npu_inst_pe_1_5_1_n21, npu_inst_pe_1_5_1_n20,
         npu_inst_pe_1_5_1_n19, npu_inst_pe_1_5_1_n18, npu_inst_pe_1_5_1_n17,
         npu_inst_pe_1_5_1_n16, npu_inst_pe_1_5_1_n15, npu_inst_pe_1_5_1_n14,
         npu_inst_pe_1_5_1_n13, npu_inst_pe_1_5_1_n12, npu_inst_pe_1_5_1_n11,
         npu_inst_pe_1_5_1_n10, npu_inst_pe_1_5_1_n9, npu_inst_pe_1_5_1_n8,
         npu_inst_pe_1_5_1_n7, npu_inst_pe_1_5_1_n6, npu_inst_pe_1_5_1_n5,
         npu_inst_pe_1_5_1_n4, npu_inst_pe_1_5_1_n3, npu_inst_pe_1_5_1_n2,
         npu_inst_pe_1_5_1_n1, npu_inst_pe_1_5_1_sub_67_carry_7_,
         npu_inst_pe_1_5_1_sub_67_carry_6_, npu_inst_pe_1_5_1_sub_67_carry_5_,
         npu_inst_pe_1_5_1_sub_67_carry_4_, npu_inst_pe_1_5_1_sub_67_carry_3_,
         npu_inst_pe_1_5_1_sub_67_carry_2_, npu_inst_pe_1_5_1_sub_67_carry_1_,
         npu_inst_pe_1_5_1_add_69_carry_7_, npu_inst_pe_1_5_1_add_69_carry_6_,
         npu_inst_pe_1_5_1_add_69_carry_5_, npu_inst_pe_1_5_1_add_69_carry_4_,
         npu_inst_pe_1_5_1_add_69_carry_3_, npu_inst_pe_1_5_1_add_69_carry_2_,
         npu_inst_pe_1_5_1_add_69_carry_1_, npu_inst_pe_1_5_1_n97,
         npu_inst_pe_1_5_1_n96, npu_inst_pe_1_5_1_n95, npu_inst_pe_1_5_1_n94,
         npu_inst_pe_1_5_1_n93, npu_inst_pe_1_5_1_n92, npu_inst_pe_1_5_1_n91,
         npu_inst_pe_1_5_1_n90, npu_inst_pe_1_5_1_n89, npu_inst_pe_1_5_1_n88,
         npu_inst_pe_1_5_1_n87, npu_inst_pe_1_5_1_n86, npu_inst_pe_1_5_1_n85,
         npu_inst_pe_1_5_1_n84, npu_inst_pe_1_5_1_n83, npu_inst_pe_1_5_1_n82,
         npu_inst_pe_1_5_1_n81, npu_inst_pe_1_5_1_n80, npu_inst_pe_1_5_1_n79,
         npu_inst_pe_1_5_1_n78, npu_inst_pe_1_5_1_n77, npu_inst_pe_1_5_1_n76,
         npu_inst_pe_1_5_1_n75, npu_inst_pe_1_5_1_n74, npu_inst_pe_1_5_1_n73,
         npu_inst_pe_1_5_1_n72, npu_inst_pe_1_5_1_n71, npu_inst_pe_1_5_1_n70,
         npu_inst_pe_1_5_1_n69, npu_inst_pe_1_5_1_n68, npu_inst_pe_1_5_1_n67,
         npu_inst_pe_1_5_1_n66, npu_inst_pe_1_5_1_n65, npu_inst_pe_1_5_1_n64,
         npu_inst_pe_1_5_1_n63, npu_inst_pe_1_5_1_n62, npu_inst_pe_1_5_1_n61,
         npu_inst_pe_1_5_1_n60, npu_inst_pe_1_5_1_n59, npu_inst_pe_1_5_1_n58,
         npu_inst_pe_1_5_1_n57, npu_inst_pe_1_5_1_n56, npu_inst_pe_1_5_1_n55,
         npu_inst_pe_1_5_1_n54, npu_inst_pe_1_5_1_n53, npu_inst_pe_1_5_1_n52,
         npu_inst_pe_1_5_1_n51, npu_inst_pe_1_5_1_n50, npu_inst_pe_1_5_1_n49,
         npu_inst_pe_1_5_1_n48, npu_inst_pe_1_5_1_n47, npu_inst_pe_1_5_1_n46,
         npu_inst_pe_1_5_1_n45, npu_inst_pe_1_5_1_n44, npu_inst_pe_1_5_1_n43,
         npu_inst_pe_1_5_1_n42, npu_inst_pe_1_5_1_n41, npu_inst_pe_1_5_1_n40,
         npu_inst_pe_1_5_1_n39, npu_inst_pe_1_5_1_n38, npu_inst_pe_1_5_1_n37,
         npu_inst_pe_1_5_1_n27, npu_inst_pe_1_5_1_n26,
         npu_inst_pe_1_5_1_net3625, npu_inst_pe_1_5_1_net3619,
         npu_inst_pe_1_5_1_N94, npu_inst_pe_1_5_1_N93, npu_inst_pe_1_5_1_N84,
         npu_inst_pe_1_5_1_N80, npu_inst_pe_1_5_1_N79, npu_inst_pe_1_5_1_N78,
         npu_inst_pe_1_5_1_N77, npu_inst_pe_1_5_1_N76, npu_inst_pe_1_5_1_N75,
         npu_inst_pe_1_5_1_N74, npu_inst_pe_1_5_1_N73, npu_inst_pe_1_5_1_N72,
         npu_inst_pe_1_5_1_N71, npu_inst_pe_1_5_1_N70, npu_inst_pe_1_5_1_N69,
         npu_inst_pe_1_5_1_N68, npu_inst_pe_1_5_1_N67, npu_inst_pe_1_5_1_N66,
         npu_inst_pe_1_5_1_N65, npu_inst_pe_1_5_1_int_q_acc_0_,
         npu_inst_pe_1_5_1_int_q_acc_1_, npu_inst_pe_1_5_1_int_q_acc_2_,
         npu_inst_pe_1_5_1_int_q_acc_3_, npu_inst_pe_1_5_1_int_q_acc_4_,
         npu_inst_pe_1_5_1_int_q_acc_5_, npu_inst_pe_1_5_1_int_q_acc_6_,
         npu_inst_pe_1_5_1_int_q_acc_7_, npu_inst_pe_1_5_1_int_data_0_,
         npu_inst_pe_1_5_1_int_data_1_, npu_inst_pe_1_5_1_int_q_weight_0_,
         npu_inst_pe_1_5_1_int_q_weight_1_,
         npu_inst_pe_1_5_1_int_q_reg_v_5__0_,
         npu_inst_pe_1_5_1_int_q_reg_v_5__1_,
         npu_inst_pe_1_5_1_int_q_reg_v_4__0_,
         npu_inst_pe_1_5_1_int_q_reg_v_4__1_,
         npu_inst_pe_1_5_1_int_q_reg_v_3__0_,
         npu_inst_pe_1_5_1_int_q_reg_v_3__1_,
         npu_inst_pe_1_5_1_int_q_reg_v_2__0_,
         npu_inst_pe_1_5_1_int_q_reg_v_2__1_,
         npu_inst_pe_1_5_1_int_q_reg_v_1__0_,
         npu_inst_pe_1_5_1_int_q_reg_v_1__1_,
         npu_inst_pe_1_5_1_int_q_reg_v_0__0_,
         npu_inst_pe_1_5_1_int_q_reg_v_0__1_,
         npu_inst_pe_1_5_1_int_q_reg_h_5__0_,
         npu_inst_pe_1_5_1_int_q_reg_h_5__1_,
         npu_inst_pe_1_5_1_int_q_reg_h_4__0_,
         npu_inst_pe_1_5_1_int_q_reg_h_4__1_,
         npu_inst_pe_1_5_1_int_q_reg_h_3__0_,
         npu_inst_pe_1_5_1_int_q_reg_h_3__1_,
         npu_inst_pe_1_5_1_int_q_reg_h_2__0_,
         npu_inst_pe_1_5_1_int_q_reg_h_2__1_,
         npu_inst_pe_1_5_1_int_q_reg_h_1__0_,
         npu_inst_pe_1_5_1_int_q_reg_h_1__1_,
         npu_inst_pe_1_5_1_int_q_reg_h_0__0_,
         npu_inst_pe_1_5_1_int_q_reg_h_0__1_, npu_inst_pe_1_5_2_n119,
         npu_inst_pe_1_5_2_n118, npu_inst_pe_1_5_2_n117,
         npu_inst_pe_1_5_2_n116, npu_inst_pe_1_5_2_n115,
         npu_inst_pe_1_5_2_n114, npu_inst_pe_1_5_2_n113,
         npu_inst_pe_1_5_2_n112, npu_inst_pe_1_5_2_n111,
         npu_inst_pe_1_5_2_n110, npu_inst_pe_1_5_2_n109,
         npu_inst_pe_1_5_2_n108, npu_inst_pe_1_5_2_n107,
         npu_inst_pe_1_5_2_n106, npu_inst_pe_1_5_2_n105,
         npu_inst_pe_1_5_2_n104, npu_inst_pe_1_5_2_n103,
         npu_inst_pe_1_5_2_n102, npu_inst_pe_1_5_2_n101,
         npu_inst_pe_1_5_2_n100, npu_inst_pe_1_5_2_n99, npu_inst_pe_1_5_2_n98,
         npu_inst_pe_1_5_2_n36, npu_inst_pe_1_5_2_n35, npu_inst_pe_1_5_2_n34,
         npu_inst_pe_1_5_2_n33, npu_inst_pe_1_5_2_n32, npu_inst_pe_1_5_2_n31,
         npu_inst_pe_1_5_2_n30, npu_inst_pe_1_5_2_n29, npu_inst_pe_1_5_2_n28,
         npu_inst_pe_1_5_2_n25, npu_inst_pe_1_5_2_n24, npu_inst_pe_1_5_2_n23,
         npu_inst_pe_1_5_2_n22, npu_inst_pe_1_5_2_n21, npu_inst_pe_1_5_2_n20,
         npu_inst_pe_1_5_2_n19, npu_inst_pe_1_5_2_n18, npu_inst_pe_1_5_2_n17,
         npu_inst_pe_1_5_2_n16, npu_inst_pe_1_5_2_n15, npu_inst_pe_1_5_2_n14,
         npu_inst_pe_1_5_2_n13, npu_inst_pe_1_5_2_n12, npu_inst_pe_1_5_2_n11,
         npu_inst_pe_1_5_2_n10, npu_inst_pe_1_5_2_n9, npu_inst_pe_1_5_2_n8,
         npu_inst_pe_1_5_2_n7, npu_inst_pe_1_5_2_n6, npu_inst_pe_1_5_2_n5,
         npu_inst_pe_1_5_2_n4, npu_inst_pe_1_5_2_n3, npu_inst_pe_1_5_2_n2,
         npu_inst_pe_1_5_2_n1, npu_inst_pe_1_5_2_sub_67_carry_7_,
         npu_inst_pe_1_5_2_sub_67_carry_6_, npu_inst_pe_1_5_2_sub_67_carry_5_,
         npu_inst_pe_1_5_2_sub_67_carry_4_, npu_inst_pe_1_5_2_sub_67_carry_3_,
         npu_inst_pe_1_5_2_sub_67_carry_2_, npu_inst_pe_1_5_2_sub_67_carry_1_,
         npu_inst_pe_1_5_2_add_69_carry_7_, npu_inst_pe_1_5_2_add_69_carry_6_,
         npu_inst_pe_1_5_2_add_69_carry_5_, npu_inst_pe_1_5_2_add_69_carry_4_,
         npu_inst_pe_1_5_2_add_69_carry_3_, npu_inst_pe_1_5_2_add_69_carry_2_,
         npu_inst_pe_1_5_2_add_69_carry_1_, npu_inst_pe_1_5_2_n97,
         npu_inst_pe_1_5_2_n96, npu_inst_pe_1_5_2_n95, npu_inst_pe_1_5_2_n94,
         npu_inst_pe_1_5_2_n93, npu_inst_pe_1_5_2_n92, npu_inst_pe_1_5_2_n91,
         npu_inst_pe_1_5_2_n90, npu_inst_pe_1_5_2_n89, npu_inst_pe_1_5_2_n88,
         npu_inst_pe_1_5_2_n87, npu_inst_pe_1_5_2_n86, npu_inst_pe_1_5_2_n85,
         npu_inst_pe_1_5_2_n84, npu_inst_pe_1_5_2_n83, npu_inst_pe_1_5_2_n82,
         npu_inst_pe_1_5_2_n81, npu_inst_pe_1_5_2_n80, npu_inst_pe_1_5_2_n79,
         npu_inst_pe_1_5_2_n78, npu_inst_pe_1_5_2_n77, npu_inst_pe_1_5_2_n76,
         npu_inst_pe_1_5_2_n75, npu_inst_pe_1_5_2_n74, npu_inst_pe_1_5_2_n73,
         npu_inst_pe_1_5_2_n72, npu_inst_pe_1_5_2_n71, npu_inst_pe_1_5_2_n70,
         npu_inst_pe_1_5_2_n69, npu_inst_pe_1_5_2_n68, npu_inst_pe_1_5_2_n67,
         npu_inst_pe_1_5_2_n66, npu_inst_pe_1_5_2_n65, npu_inst_pe_1_5_2_n64,
         npu_inst_pe_1_5_2_n63, npu_inst_pe_1_5_2_n62, npu_inst_pe_1_5_2_n61,
         npu_inst_pe_1_5_2_n60, npu_inst_pe_1_5_2_n59, npu_inst_pe_1_5_2_n58,
         npu_inst_pe_1_5_2_n57, npu_inst_pe_1_5_2_n56, npu_inst_pe_1_5_2_n55,
         npu_inst_pe_1_5_2_n54, npu_inst_pe_1_5_2_n53, npu_inst_pe_1_5_2_n52,
         npu_inst_pe_1_5_2_n51, npu_inst_pe_1_5_2_n50, npu_inst_pe_1_5_2_n49,
         npu_inst_pe_1_5_2_n48, npu_inst_pe_1_5_2_n47, npu_inst_pe_1_5_2_n46,
         npu_inst_pe_1_5_2_n45, npu_inst_pe_1_5_2_n44, npu_inst_pe_1_5_2_n43,
         npu_inst_pe_1_5_2_n42, npu_inst_pe_1_5_2_n41, npu_inst_pe_1_5_2_n40,
         npu_inst_pe_1_5_2_n39, npu_inst_pe_1_5_2_n38, npu_inst_pe_1_5_2_n37,
         npu_inst_pe_1_5_2_n27, npu_inst_pe_1_5_2_n26,
         npu_inst_pe_1_5_2_net3602, npu_inst_pe_1_5_2_net3596,
         npu_inst_pe_1_5_2_N94, npu_inst_pe_1_5_2_N93, npu_inst_pe_1_5_2_N84,
         npu_inst_pe_1_5_2_N80, npu_inst_pe_1_5_2_N79, npu_inst_pe_1_5_2_N78,
         npu_inst_pe_1_5_2_N77, npu_inst_pe_1_5_2_N76, npu_inst_pe_1_5_2_N75,
         npu_inst_pe_1_5_2_N74, npu_inst_pe_1_5_2_N73, npu_inst_pe_1_5_2_N72,
         npu_inst_pe_1_5_2_N71, npu_inst_pe_1_5_2_N70, npu_inst_pe_1_5_2_N69,
         npu_inst_pe_1_5_2_N68, npu_inst_pe_1_5_2_N67, npu_inst_pe_1_5_2_N66,
         npu_inst_pe_1_5_2_N65, npu_inst_pe_1_5_2_int_q_acc_0_,
         npu_inst_pe_1_5_2_int_q_acc_1_, npu_inst_pe_1_5_2_int_q_acc_2_,
         npu_inst_pe_1_5_2_int_q_acc_3_, npu_inst_pe_1_5_2_int_q_acc_4_,
         npu_inst_pe_1_5_2_int_q_acc_5_, npu_inst_pe_1_5_2_int_q_acc_6_,
         npu_inst_pe_1_5_2_int_q_acc_7_, npu_inst_pe_1_5_2_int_data_0_,
         npu_inst_pe_1_5_2_int_data_1_, npu_inst_pe_1_5_2_int_q_weight_0_,
         npu_inst_pe_1_5_2_int_q_weight_1_,
         npu_inst_pe_1_5_2_int_q_reg_v_5__0_,
         npu_inst_pe_1_5_2_int_q_reg_v_5__1_,
         npu_inst_pe_1_5_2_int_q_reg_v_4__0_,
         npu_inst_pe_1_5_2_int_q_reg_v_4__1_,
         npu_inst_pe_1_5_2_int_q_reg_v_3__0_,
         npu_inst_pe_1_5_2_int_q_reg_v_3__1_,
         npu_inst_pe_1_5_2_int_q_reg_v_2__0_,
         npu_inst_pe_1_5_2_int_q_reg_v_2__1_,
         npu_inst_pe_1_5_2_int_q_reg_v_1__0_,
         npu_inst_pe_1_5_2_int_q_reg_v_1__1_,
         npu_inst_pe_1_5_2_int_q_reg_v_0__0_,
         npu_inst_pe_1_5_2_int_q_reg_v_0__1_,
         npu_inst_pe_1_5_2_int_q_reg_h_5__0_,
         npu_inst_pe_1_5_2_int_q_reg_h_5__1_,
         npu_inst_pe_1_5_2_int_q_reg_h_4__0_,
         npu_inst_pe_1_5_2_int_q_reg_h_4__1_,
         npu_inst_pe_1_5_2_int_q_reg_h_3__0_,
         npu_inst_pe_1_5_2_int_q_reg_h_3__1_,
         npu_inst_pe_1_5_2_int_q_reg_h_2__0_,
         npu_inst_pe_1_5_2_int_q_reg_h_2__1_,
         npu_inst_pe_1_5_2_int_q_reg_h_1__0_,
         npu_inst_pe_1_5_2_int_q_reg_h_1__1_,
         npu_inst_pe_1_5_2_int_q_reg_h_0__0_,
         npu_inst_pe_1_5_2_int_q_reg_h_0__1_, npu_inst_pe_1_5_3_n119,
         npu_inst_pe_1_5_3_n118, npu_inst_pe_1_5_3_n117,
         npu_inst_pe_1_5_3_n116, npu_inst_pe_1_5_3_n115,
         npu_inst_pe_1_5_3_n114, npu_inst_pe_1_5_3_n113,
         npu_inst_pe_1_5_3_n112, npu_inst_pe_1_5_3_n111,
         npu_inst_pe_1_5_3_n110, npu_inst_pe_1_5_3_n109,
         npu_inst_pe_1_5_3_n108, npu_inst_pe_1_5_3_n107,
         npu_inst_pe_1_5_3_n106, npu_inst_pe_1_5_3_n105,
         npu_inst_pe_1_5_3_n104, npu_inst_pe_1_5_3_n103,
         npu_inst_pe_1_5_3_n102, npu_inst_pe_1_5_3_n101,
         npu_inst_pe_1_5_3_n100, npu_inst_pe_1_5_3_n99, npu_inst_pe_1_5_3_n98,
         npu_inst_pe_1_5_3_n36, npu_inst_pe_1_5_3_n35, npu_inst_pe_1_5_3_n34,
         npu_inst_pe_1_5_3_n33, npu_inst_pe_1_5_3_n32, npu_inst_pe_1_5_3_n31,
         npu_inst_pe_1_5_3_n30, npu_inst_pe_1_5_3_n29, npu_inst_pe_1_5_3_n28,
         npu_inst_pe_1_5_3_n25, npu_inst_pe_1_5_3_n24, npu_inst_pe_1_5_3_n23,
         npu_inst_pe_1_5_3_n22, npu_inst_pe_1_5_3_n21, npu_inst_pe_1_5_3_n20,
         npu_inst_pe_1_5_3_n19, npu_inst_pe_1_5_3_n18, npu_inst_pe_1_5_3_n17,
         npu_inst_pe_1_5_3_n16, npu_inst_pe_1_5_3_n15, npu_inst_pe_1_5_3_n14,
         npu_inst_pe_1_5_3_n13, npu_inst_pe_1_5_3_n12, npu_inst_pe_1_5_3_n11,
         npu_inst_pe_1_5_3_n10, npu_inst_pe_1_5_3_n9, npu_inst_pe_1_5_3_n8,
         npu_inst_pe_1_5_3_n7, npu_inst_pe_1_5_3_n6, npu_inst_pe_1_5_3_n5,
         npu_inst_pe_1_5_3_n4, npu_inst_pe_1_5_3_n3, npu_inst_pe_1_5_3_n2,
         npu_inst_pe_1_5_3_n1, npu_inst_pe_1_5_3_sub_67_carry_7_,
         npu_inst_pe_1_5_3_sub_67_carry_6_, npu_inst_pe_1_5_3_sub_67_carry_5_,
         npu_inst_pe_1_5_3_sub_67_carry_4_, npu_inst_pe_1_5_3_sub_67_carry_3_,
         npu_inst_pe_1_5_3_sub_67_carry_2_, npu_inst_pe_1_5_3_sub_67_carry_1_,
         npu_inst_pe_1_5_3_add_69_carry_7_, npu_inst_pe_1_5_3_add_69_carry_6_,
         npu_inst_pe_1_5_3_add_69_carry_5_, npu_inst_pe_1_5_3_add_69_carry_4_,
         npu_inst_pe_1_5_3_add_69_carry_3_, npu_inst_pe_1_5_3_add_69_carry_2_,
         npu_inst_pe_1_5_3_add_69_carry_1_, npu_inst_pe_1_5_3_n97,
         npu_inst_pe_1_5_3_n96, npu_inst_pe_1_5_3_n95, npu_inst_pe_1_5_3_n94,
         npu_inst_pe_1_5_3_n93, npu_inst_pe_1_5_3_n92, npu_inst_pe_1_5_3_n91,
         npu_inst_pe_1_5_3_n90, npu_inst_pe_1_5_3_n89, npu_inst_pe_1_5_3_n88,
         npu_inst_pe_1_5_3_n87, npu_inst_pe_1_5_3_n86, npu_inst_pe_1_5_3_n85,
         npu_inst_pe_1_5_3_n84, npu_inst_pe_1_5_3_n83, npu_inst_pe_1_5_3_n82,
         npu_inst_pe_1_5_3_n81, npu_inst_pe_1_5_3_n80, npu_inst_pe_1_5_3_n79,
         npu_inst_pe_1_5_3_n78, npu_inst_pe_1_5_3_n77, npu_inst_pe_1_5_3_n76,
         npu_inst_pe_1_5_3_n75, npu_inst_pe_1_5_3_n74, npu_inst_pe_1_5_3_n73,
         npu_inst_pe_1_5_3_n72, npu_inst_pe_1_5_3_n71, npu_inst_pe_1_5_3_n70,
         npu_inst_pe_1_5_3_n69, npu_inst_pe_1_5_3_n68, npu_inst_pe_1_5_3_n67,
         npu_inst_pe_1_5_3_n66, npu_inst_pe_1_5_3_n65, npu_inst_pe_1_5_3_n64,
         npu_inst_pe_1_5_3_n63, npu_inst_pe_1_5_3_n62, npu_inst_pe_1_5_3_n61,
         npu_inst_pe_1_5_3_n60, npu_inst_pe_1_5_3_n59, npu_inst_pe_1_5_3_n58,
         npu_inst_pe_1_5_3_n57, npu_inst_pe_1_5_3_n56, npu_inst_pe_1_5_3_n55,
         npu_inst_pe_1_5_3_n54, npu_inst_pe_1_5_3_n53, npu_inst_pe_1_5_3_n52,
         npu_inst_pe_1_5_3_n51, npu_inst_pe_1_5_3_n50, npu_inst_pe_1_5_3_n49,
         npu_inst_pe_1_5_3_n48, npu_inst_pe_1_5_3_n47, npu_inst_pe_1_5_3_n46,
         npu_inst_pe_1_5_3_n45, npu_inst_pe_1_5_3_n44, npu_inst_pe_1_5_3_n43,
         npu_inst_pe_1_5_3_n42, npu_inst_pe_1_5_3_n41, npu_inst_pe_1_5_3_n40,
         npu_inst_pe_1_5_3_n39, npu_inst_pe_1_5_3_n38, npu_inst_pe_1_5_3_n37,
         npu_inst_pe_1_5_3_n27, npu_inst_pe_1_5_3_n26,
         npu_inst_pe_1_5_3_net3579, npu_inst_pe_1_5_3_net3573,
         npu_inst_pe_1_5_3_N94, npu_inst_pe_1_5_3_N93, npu_inst_pe_1_5_3_N84,
         npu_inst_pe_1_5_3_N80, npu_inst_pe_1_5_3_N79, npu_inst_pe_1_5_3_N78,
         npu_inst_pe_1_5_3_N77, npu_inst_pe_1_5_3_N76, npu_inst_pe_1_5_3_N75,
         npu_inst_pe_1_5_3_N74, npu_inst_pe_1_5_3_N73, npu_inst_pe_1_5_3_N72,
         npu_inst_pe_1_5_3_N71, npu_inst_pe_1_5_3_N70, npu_inst_pe_1_5_3_N69,
         npu_inst_pe_1_5_3_N68, npu_inst_pe_1_5_3_N67, npu_inst_pe_1_5_3_N66,
         npu_inst_pe_1_5_3_N65, npu_inst_pe_1_5_3_int_q_acc_0_,
         npu_inst_pe_1_5_3_int_q_acc_1_, npu_inst_pe_1_5_3_int_q_acc_2_,
         npu_inst_pe_1_5_3_int_q_acc_3_, npu_inst_pe_1_5_3_int_q_acc_4_,
         npu_inst_pe_1_5_3_int_q_acc_5_, npu_inst_pe_1_5_3_int_q_acc_6_,
         npu_inst_pe_1_5_3_int_q_acc_7_, npu_inst_pe_1_5_3_int_data_0_,
         npu_inst_pe_1_5_3_int_data_1_, npu_inst_pe_1_5_3_int_q_weight_0_,
         npu_inst_pe_1_5_3_int_q_weight_1_,
         npu_inst_pe_1_5_3_int_q_reg_v_5__0_,
         npu_inst_pe_1_5_3_int_q_reg_v_5__1_,
         npu_inst_pe_1_5_3_int_q_reg_v_4__0_,
         npu_inst_pe_1_5_3_int_q_reg_v_4__1_,
         npu_inst_pe_1_5_3_int_q_reg_v_3__0_,
         npu_inst_pe_1_5_3_int_q_reg_v_3__1_,
         npu_inst_pe_1_5_3_int_q_reg_v_2__0_,
         npu_inst_pe_1_5_3_int_q_reg_v_2__1_,
         npu_inst_pe_1_5_3_int_q_reg_v_1__0_,
         npu_inst_pe_1_5_3_int_q_reg_v_1__1_,
         npu_inst_pe_1_5_3_int_q_reg_v_0__0_,
         npu_inst_pe_1_5_3_int_q_reg_v_0__1_,
         npu_inst_pe_1_5_3_int_q_reg_h_5__0_,
         npu_inst_pe_1_5_3_int_q_reg_h_5__1_,
         npu_inst_pe_1_5_3_int_q_reg_h_4__0_,
         npu_inst_pe_1_5_3_int_q_reg_h_4__1_,
         npu_inst_pe_1_5_3_int_q_reg_h_3__0_,
         npu_inst_pe_1_5_3_int_q_reg_h_3__1_,
         npu_inst_pe_1_5_3_int_q_reg_h_2__0_,
         npu_inst_pe_1_5_3_int_q_reg_h_2__1_,
         npu_inst_pe_1_5_3_int_q_reg_h_1__0_,
         npu_inst_pe_1_5_3_int_q_reg_h_1__1_,
         npu_inst_pe_1_5_3_int_q_reg_h_0__0_,
         npu_inst_pe_1_5_3_int_q_reg_h_0__1_, npu_inst_pe_1_5_4_n119,
         npu_inst_pe_1_5_4_n118, npu_inst_pe_1_5_4_n117,
         npu_inst_pe_1_5_4_n116, npu_inst_pe_1_5_4_n115,
         npu_inst_pe_1_5_4_n114, npu_inst_pe_1_5_4_n113,
         npu_inst_pe_1_5_4_n112, npu_inst_pe_1_5_4_n111,
         npu_inst_pe_1_5_4_n110, npu_inst_pe_1_5_4_n109,
         npu_inst_pe_1_5_4_n108, npu_inst_pe_1_5_4_n107,
         npu_inst_pe_1_5_4_n106, npu_inst_pe_1_5_4_n105,
         npu_inst_pe_1_5_4_n104, npu_inst_pe_1_5_4_n103,
         npu_inst_pe_1_5_4_n102, npu_inst_pe_1_5_4_n101,
         npu_inst_pe_1_5_4_n100, npu_inst_pe_1_5_4_n99, npu_inst_pe_1_5_4_n98,
         npu_inst_pe_1_5_4_n36, npu_inst_pe_1_5_4_n35, npu_inst_pe_1_5_4_n34,
         npu_inst_pe_1_5_4_n33, npu_inst_pe_1_5_4_n32, npu_inst_pe_1_5_4_n31,
         npu_inst_pe_1_5_4_n30, npu_inst_pe_1_5_4_n29, npu_inst_pe_1_5_4_n28,
         npu_inst_pe_1_5_4_n25, npu_inst_pe_1_5_4_n24, npu_inst_pe_1_5_4_n23,
         npu_inst_pe_1_5_4_n22, npu_inst_pe_1_5_4_n21, npu_inst_pe_1_5_4_n20,
         npu_inst_pe_1_5_4_n19, npu_inst_pe_1_5_4_n18, npu_inst_pe_1_5_4_n17,
         npu_inst_pe_1_5_4_n16, npu_inst_pe_1_5_4_n15, npu_inst_pe_1_5_4_n14,
         npu_inst_pe_1_5_4_n13, npu_inst_pe_1_5_4_n12, npu_inst_pe_1_5_4_n11,
         npu_inst_pe_1_5_4_n10, npu_inst_pe_1_5_4_n9, npu_inst_pe_1_5_4_n8,
         npu_inst_pe_1_5_4_n7, npu_inst_pe_1_5_4_n6, npu_inst_pe_1_5_4_n5,
         npu_inst_pe_1_5_4_n4, npu_inst_pe_1_5_4_n3, npu_inst_pe_1_5_4_n2,
         npu_inst_pe_1_5_4_n1, npu_inst_pe_1_5_4_sub_67_carry_7_,
         npu_inst_pe_1_5_4_sub_67_carry_6_, npu_inst_pe_1_5_4_sub_67_carry_5_,
         npu_inst_pe_1_5_4_sub_67_carry_4_, npu_inst_pe_1_5_4_sub_67_carry_3_,
         npu_inst_pe_1_5_4_sub_67_carry_2_, npu_inst_pe_1_5_4_sub_67_carry_1_,
         npu_inst_pe_1_5_4_add_69_carry_7_, npu_inst_pe_1_5_4_add_69_carry_6_,
         npu_inst_pe_1_5_4_add_69_carry_5_, npu_inst_pe_1_5_4_add_69_carry_4_,
         npu_inst_pe_1_5_4_add_69_carry_3_, npu_inst_pe_1_5_4_add_69_carry_2_,
         npu_inst_pe_1_5_4_add_69_carry_1_, npu_inst_pe_1_5_4_n97,
         npu_inst_pe_1_5_4_n96, npu_inst_pe_1_5_4_n95, npu_inst_pe_1_5_4_n94,
         npu_inst_pe_1_5_4_n93, npu_inst_pe_1_5_4_n92, npu_inst_pe_1_5_4_n91,
         npu_inst_pe_1_5_4_n90, npu_inst_pe_1_5_4_n89, npu_inst_pe_1_5_4_n88,
         npu_inst_pe_1_5_4_n87, npu_inst_pe_1_5_4_n86, npu_inst_pe_1_5_4_n85,
         npu_inst_pe_1_5_4_n84, npu_inst_pe_1_5_4_n83, npu_inst_pe_1_5_4_n82,
         npu_inst_pe_1_5_4_n81, npu_inst_pe_1_5_4_n80, npu_inst_pe_1_5_4_n79,
         npu_inst_pe_1_5_4_n78, npu_inst_pe_1_5_4_n77, npu_inst_pe_1_5_4_n76,
         npu_inst_pe_1_5_4_n75, npu_inst_pe_1_5_4_n74, npu_inst_pe_1_5_4_n73,
         npu_inst_pe_1_5_4_n72, npu_inst_pe_1_5_4_n71, npu_inst_pe_1_5_4_n70,
         npu_inst_pe_1_5_4_n69, npu_inst_pe_1_5_4_n68, npu_inst_pe_1_5_4_n67,
         npu_inst_pe_1_5_4_n66, npu_inst_pe_1_5_4_n65, npu_inst_pe_1_5_4_n64,
         npu_inst_pe_1_5_4_n63, npu_inst_pe_1_5_4_n62, npu_inst_pe_1_5_4_n61,
         npu_inst_pe_1_5_4_n60, npu_inst_pe_1_5_4_n59, npu_inst_pe_1_5_4_n58,
         npu_inst_pe_1_5_4_n57, npu_inst_pe_1_5_4_n56, npu_inst_pe_1_5_4_n55,
         npu_inst_pe_1_5_4_n54, npu_inst_pe_1_5_4_n53, npu_inst_pe_1_5_4_n52,
         npu_inst_pe_1_5_4_n51, npu_inst_pe_1_5_4_n50, npu_inst_pe_1_5_4_n49,
         npu_inst_pe_1_5_4_n48, npu_inst_pe_1_5_4_n47, npu_inst_pe_1_5_4_n46,
         npu_inst_pe_1_5_4_n45, npu_inst_pe_1_5_4_n44, npu_inst_pe_1_5_4_n43,
         npu_inst_pe_1_5_4_n42, npu_inst_pe_1_5_4_n41, npu_inst_pe_1_5_4_n40,
         npu_inst_pe_1_5_4_n39, npu_inst_pe_1_5_4_n38, npu_inst_pe_1_5_4_n37,
         npu_inst_pe_1_5_4_n27, npu_inst_pe_1_5_4_n26,
         npu_inst_pe_1_5_4_net3556, npu_inst_pe_1_5_4_net3550,
         npu_inst_pe_1_5_4_N94, npu_inst_pe_1_5_4_N93, npu_inst_pe_1_5_4_N84,
         npu_inst_pe_1_5_4_N80, npu_inst_pe_1_5_4_N79, npu_inst_pe_1_5_4_N78,
         npu_inst_pe_1_5_4_N77, npu_inst_pe_1_5_4_N76, npu_inst_pe_1_5_4_N75,
         npu_inst_pe_1_5_4_N74, npu_inst_pe_1_5_4_N73, npu_inst_pe_1_5_4_N72,
         npu_inst_pe_1_5_4_N71, npu_inst_pe_1_5_4_N70, npu_inst_pe_1_5_4_N69,
         npu_inst_pe_1_5_4_N68, npu_inst_pe_1_5_4_N67, npu_inst_pe_1_5_4_N66,
         npu_inst_pe_1_5_4_N65, npu_inst_pe_1_5_4_int_q_acc_0_,
         npu_inst_pe_1_5_4_int_q_acc_1_, npu_inst_pe_1_5_4_int_q_acc_2_,
         npu_inst_pe_1_5_4_int_q_acc_3_, npu_inst_pe_1_5_4_int_q_acc_4_,
         npu_inst_pe_1_5_4_int_q_acc_5_, npu_inst_pe_1_5_4_int_q_acc_6_,
         npu_inst_pe_1_5_4_int_q_acc_7_, npu_inst_pe_1_5_4_int_data_0_,
         npu_inst_pe_1_5_4_int_data_1_, npu_inst_pe_1_5_4_int_q_weight_0_,
         npu_inst_pe_1_5_4_int_q_weight_1_,
         npu_inst_pe_1_5_4_int_q_reg_v_5__0_,
         npu_inst_pe_1_5_4_int_q_reg_v_5__1_,
         npu_inst_pe_1_5_4_int_q_reg_v_4__0_,
         npu_inst_pe_1_5_4_int_q_reg_v_4__1_,
         npu_inst_pe_1_5_4_int_q_reg_v_3__0_,
         npu_inst_pe_1_5_4_int_q_reg_v_3__1_,
         npu_inst_pe_1_5_4_int_q_reg_v_2__0_,
         npu_inst_pe_1_5_4_int_q_reg_v_2__1_,
         npu_inst_pe_1_5_4_int_q_reg_v_1__0_,
         npu_inst_pe_1_5_4_int_q_reg_v_1__1_,
         npu_inst_pe_1_5_4_int_q_reg_v_0__0_,
         npu_inst_pe_1_5_4_int_q_reg_v_0__1_,
         npu_inst_pe_1_5_4_int_q_reg_h_5__0_,
         npu_inst_pe_1_5_4_int_q_reg_h_5__1_,
         npu_inst_pe_1_5_4_int_q_reg_h_4__0_,
         npu_inst_pe_1_5_4_int_q_reg_h_4__1_,
         npu_inst_pe_1_5_4_int_q_reg_h_3__0_,
         npu_inst_pe_1_5_4_int_q_reg_h_3__1_,
         npu_inst_pe_1_5_4_int_q_reg_h_2__0_,
         npu_inst_pe_1_5_4_int_q_reg_h_2__1_,
         npu_inst_pe_1_5_4_int_q_reg_h_1__0_,
         npu_inst_pe_1_5_4_int_q_reg_h_1__1_,
         npu_inst_pe_1_5_4_int_q_reg_h_0__0_,
         npu_inst_pe_1_5_4_int_q_reg_h_0__1_, npu_inst_pe_1_5_5_n119,
         npu_inst_pe_1_5_5_n118, npu_inst_pe_1_5_5_n117,
         npu_inst_pe_1_5_5_n116, npu_inst_pe_1_5_5_n115,
         npu_inst_pe_1_5_5_n114, npu_inst_pe_1_5_5_n113,
         npu_inst_pe_1_5_5_n112, npu_inst_pe_1_5_5_n111,
         npu_inst_pe_1_5_5_n110, npu_inst_pe_1_5_5_n109,
         npu_inst_pe_1_5_5_n108, npu_inst_pe_1_5_5_n107,
         npu_inst_pe_1_5_5_n106, npu_inst_pe_1_5_5_n105,
         npu_inst_pe_1_5_5_n104, npu_inst_pe_1_5_5_n103,
         npu_inst_pe_1_5_5_n102, npu_inst_pe_1_5_5_n101,
         npu_inst_pe_1_5_5_n100, npu_inst_pe_1_5_5_n99, npu_inst_pe_1_5_5_n98,
         npu_inst_pe_1_5_5_n36, npu_inst_pe_1_5_5_n35, npu_inst_pe_1_5_5_n34,
         npu_inst_pe_1_5_5_n33, npu_inst_pe_1_5_5_n32, npu_inst_pe_1_5_5_n31,
         npu_inst_pe_1_5_5_n30, npu_inst_pe_1_5_5_n29, npu_inst_pe_1_5_5_n28,
         npu_inst_pe_1_5_5_n25, npu_inst_pe_1_5_5_n24, npu_inst_pe_1_5_5_n23,
         npu_inst_pe_1_5_5_n22, npu_inst_pe_1_5_5_n21, npu_inst_pe_1_5_5_n20,
         npu_inst_pe_1_5_5_n19, npu_inst_pe_1_5_5_n18, npu_inst_pe_1_5_5_n17,
         npu_inst_pe_1_5_5_n16, npu_inst_pe_1_5_5_n15, npu_inst_pe_1_5_5_n14,
         npu_inst_pe_1_5_5_n13, npu_inst_pe_1_5_5_n12, npu_inst_pe_1_5_5_n11,
         npu_inst_pe_1_5_5_n10, npu_inst_pe_1_5_5_n9, npu_inst_pe_1_5_5_n8,
         npu_inst_pe_1_5_5_n7, npu_inst_pe_1_5_5_n6, npu_inst_pe_1_5_5_n5,
         npu_inst_pe_1_5_5_n4, npu_inst_pe_1_5_5_n3, npu_inst_pe_1_5_5_n2,
         npu_inst_pe_1_5_5_n1, npu_inst_pe_1_5_5_sub_67_carry_7_,
         npu_inst_pe_1_5_5_sub_67_carry_6_, npu_inst_pe_1_5_5_sub_67_carry_5_,
         npu_inst_pe_1_5_5_sub_67_carry_4_, npu_inst_pe_1_5_5_sub_67_carry_3_,
         npu_inst_pe_1_5_5_sub_67_carry_2_, npu_inst_pe_1_5_5_sub_67_carry_1_,
         npu_inst_pe_1_5_5_add_69_carry_7_, npu_inst_pe_1_5_5_add_69_carry_6_,
         npu_inst_pe_1_5_5_add_69_carry_5_, npu_inst_pe_1_5_5_add_69_carry_4_,
         npu_inst_pe_1_5_5_add_69_carry_3_, npu_inst_pe_1_5_5_add_69_carry_2_,
         npu_inst_pe_1_5_5_add_69_carry_1_, npu_inst_pe_1_5_5_n97,
         npu_inst_pe_1_5_5_n96, npu_inst_pe_1_5_5_n95, npu_inst_pe_1_5_5_n94,
         npu_inst_pe_1_5_5_n93, npu_inst_pe_1_5_5_n92, npu_inst_pe_1_5_5_n91,
         npu_inst_pe_1_5_5_n90, npu_inst_pe_1_5_5_n89, npu_inst_pe_1_5_5_n88,
         npu_inst_pe_1_5_5_n87, npu_inst_pe_1_5_5_n86, npu_inst_pe_1_5_5_n85,
         npu_inst_pe_1_5_5_n84, npu_inst_pe_1_5_5_n83, npu_inst_pe_1_5_5_n82,
         npu_inst_pe_1_5_5_n81, npu_inst_pe_1_5_5_n80, npu_inst_pe_1_5_5_n79,
         npu_inst_pe_1_5_5_n78, npu_inst_pe_1_5_5_n77, npu_inst_pe_1_5_5_n76,
         npu_inst_pe_1_5_5_n75, npu_inst_pe_1_5_5_n74, npu_inst_pe_1_5_5_n73,
         npu_inst_pe_1_5_5_n72, npu_inst_pe_1_5_5_n71, npu_inst_pe_1_5_5_n70,
         npu_inst_pe_1_5_5_n69, npu_inst_pe_1_5_5_n68, npu_inst_pe_1_5_5_n67,
         npu_inst_pe_1_5_5_n66, npu_inst_pe_1_5_5_n65, npu_inst_pe_1_5_5_n64,
         npu_inst_pe_1_5_5_n63, npu_inst_pe_1_5_5_n62, npu_inst_pe_1_5_5_n61,
         npu_inst_pe_1_5_5_n60, npu_inst_pe_1_5_5_n59, npu_inst_pe_1_5_5_n58,
         npu_inst_pe_1_5_5_n57, npu_inst_pe_1_5_5_n56, npu_inst_pe_1_5_5_n55,
         npu_inst_pe_1_5_5_n54, npu_inst_pe_1_5_5_n53, npu_inst_pe_1_5_5_n52,
         npu_inst_pe_1_5_5_n51, npu_inst_pe_1_5_5_n50, npu_inst_pe_1_5_5_n49,
         npu_inst_pe_1_5_5_n48, npu_inst_pe_1_5_5_n47, npu_inst_pe_1_5_5_n46,
         npu_inst_pe_1_5_5_n45, npu_inst_pe_1_5_5_n44, npu_inst_pe_1_5_5_n43,
         npu_inst_pe_1_5_5_n42, npu_inst_pe_1_5_5_n41, npu_inst_pe_1_5_5_n40,
         npu_inst_pe_1_5_5_n39, npu_inst_pe_1_5_5_n38, npu_inst_pe_1_5_5_n37,
         npu_inst_pe_1_5_5_n27, npu_inst_pe_1_5_5_n26,
         npu_inst_pe_1_5_5_net3533, npu_inst_pe_1_5_5_net3527,
         npu_inst_pe_1_5_5_N94, npu_inst_pe_1_5_5_N93, npu_inst_pe_1_5_5_N84,
         npu_inst_pe_1_5_5_N80, npu_inst_pe_1_5_5_N79, npu_inst_pe_1_5_5_N78,
         npu_inst_pe_1_5_5_N77, npu_inst_pe_1_5_5_N76, npu_inst_pe_1_5_5_N75,
         npu_inst_pe_1_5_5_N74, npu_inst_pe_1_5_5_N73, npu_inst_pe_1_5_5_N72,
         npu_inst_pe_1_5_5_N71, npu_inst_pe_1_5_5_N70, npu_inst_pe_1_5_5_N69,
         npu_inst_pe_1_5_5_N68, npu_inst_pe_1_5_5_N67, npu_inst_pe_1_5_5_N66,
         npu_inst_pe_1_5_5_N65, npu_inst_pe_1_5_5_int_q_acc_0_,
         npu_inst_pe_1_5_5_int_q_acc_1_, npu_inst_pe_1_5_5_int_q_acc_2_,
         npu_inst_pe_1_5_5_int_q_acc_3_, npu_inst_pe_1_5_5_int_q_acc_4_,
         npu_inst_pe_1_5_5_int_q_acc_5_, npu_inst_pe_1_5_5_int_q_acc_6_,
         npu_inst_pe_1_5_5_int_q_acc_7_, npu_inst_pe_1_5_5_int_data_0_,
         npu_inst_pe_1_5_5_int_data_1_, npu_inst_pe_1_5_5_int_q_weight_0_,
         npu_inst_pe_1_5_5_int_q_weight_1_,
         npu_inst_pe_1_5_5_int_q_reg_v_5__0_,
         npu_inst_pe_1_5_5_int_q_reg_v_5__1_,
         npu_inst_pe_1_5_5_int_q_reg_v_4__0_,
         npu_inst_pe_1_5_5_int_q_reg_v_4__1_,
         npu_inst_pe_1_5_5_int_q_reg_v_3__0_,
         npu_inst_pe_1_5_5_int_q_reg_v_3__1_,
         npu_inst_pe_1_5_5_int_q_reg_v_2__0_,
         npu_inst_pe_1_5_5_int_q_reg_v_2__1_,
         npu_inst_pe_1_5_5_int_q_reg_v_1__0_,
         npu_inst_pe_1_5_5_int_q_reg_v_1__1_,
         npu_inst_pe_1_5_5_int_q_reg_v_0__0_,
         npu_inst_pe_1_5_5_int_q_reg_v_0__1_,
         npu_inst_pe_1_5_5_int_q_reg_h_5__0_,
         npu_inst_pe_1_5_5_int_q_reg_h_5__1_,
         npu_inst_pe_1_5_5_int_q_reg_h_4__0_,
         npu_inst_pe_1_5_5_int_q_reg_h_4__1_,
         npu_inst_pe_1_5_5_int_q_reg_h_3__0_,
         npu_inst_pe_1_5_5_int_q_reg_h_3__1_,
         npu_inst_pe_1_5_5_int_q_reg_h_2__0_,
         npu_inst_pe_1_5_5_int_q_reg_h_2__1_,
         npu_inst_pe_1_5_5_int_q_reg_h_1__0_,
         npu_inst_pe_1_5_5_int_q_reg_h_1__1_,
         npu_inst_pe_1_5_5_int_q_reg_h_0__0_,
         npu_inst_pe_1_5_5_int_q_reg_h_0__1_, npu_inst_pe_1_5_6_n119,
         npu_inst_pe_1_5_6_n118, npu_inst_pe_1_5_6_n117,
         npu_inst_pe_1_5_6_n116, npu_inst_pe_1_5_6_n115,
         npu_inst_pe_1_5_6_n114, npu_inst_pe_1_5_6_n113,
         npu_inst_pe_1_5_6_n112, npu_inst_pe_1_5_6_n111,
         npu_inst_pe_1_5_6_n110, npu_inst_pe_1_5_6_n109,
         npu_inst_pe_1_5_6_n108, npu_inst_pe_1_5_6_n107,
         npu_inst_pe_1_5_6_n106, npu_inst_pe_1_5_6_n105,
         npu_inst_pe_1_5_6_n104, npu_inst_pe_1_5_6_n103,
         npu_inst_pe_1_5_6_n102, npu_inst_pe_1_5_6_n101,
         npu_inst_pe_1_5_6_n100, npu_inst_pe_1_5_6_n99, npu_inst_pe_1_5_6_n98,
         npu_inst_pe_1_5_6_n36, npu_inst_pe_1_5_6_n35, npu_inst_pe_1_5_6_n34,
         npu_inst_pe_1_5_6_n33, npu_inst_pe_1_5_6_n32, npu_inst_pe_1_5_6_n31,
         npu_inst_pe_1_5_6_n30, npu_inst_pe_1_5_6_n29, npu_inst_pe_1_5_6_n28,
         npu_inst_pe_1_5_6_n25, npu_inst_pe_1_5_6_n24, npu_inst_pe_1_5_6_n23,
         npu_inst_pe_1_5_6_n22, npu_inst_pe_1_5_6_n21, npu_inst_pe_1_5_6_n20,
         npu_inst_pe_1_5_6_n19, npu_inst_pe_1_5_6_n18, npu_inst_pe_1_5_6_n17,
         npu_inst_pe_1_5_6_n16, npu_inst_pe_1_5_6_n15, npu_inst_pe_1_5_6_n14,
         npu_inst_pe_1_5_6_n13, npu_inst_pe_1_5_6_n12, npu_inst_pe_1_5_6_n11,
         npu_inst_pe_1_5_6_n10, npu_inst_pe_1_5_6_n9, npu_inst_pe_1_5_6_n8,
         npu_inst_pe_1_5_6_n7, npu_inst_pe_1_5_6_n6, npu_inst_pe_1_5_6_n5,
         npu_inst_pe_1_5_6_n4, npu_inst_pe_1_5_6_n3, npu_inst_pe_1_5_6_n2,
         npu_inst_pe_1_5_6_n1, npu_inst_pe_1_5_6_sub_67_carry_7_,
         npu_inst_pe_1_5_6_sub_67_carry_6_, npu_inst_pe_1_5_6_sub_67_carry_5_,
         npu_inst_pe_1_5_6_sub_67_carry_4_, npu_inst_pe_1_5_6_sub_67_carry_3_,
         npu_inst_pe_1_5_6_sub_67_carry_2_, npu_inst_pe_1_5_6_sub_67_carry_1_,
         npu_inst_pe_1_5_6_add_69_carry_7_, npu_inst_pe_1_5_6_add_69_carry_6_,
         npu_inst_pe_1_5_6_add_69_carry_5_, npu_inst_pe_1_5_6_add_69_carry_4_,
         npu_inst_pe_1_5_6_add_69_carry_3_, npu_inst_pe_1_5_6_add_69_carry_2_,
         npu_inst_pe_1_5_6_add_69_carry_1_, npu_inst_pe_1_5_6_n97,
         npu_inst_pe_1_5_6_n96, npu_inst_pe_1_5_6_n95, npu_inst_pe_1_5_6_n94,
         npu_inst_pe_1_5_6_n93, npu_inst_pe_1_5_6_n92, npu_inst_pe_1_5_6_n91,
         npu_inst_pe_1_5_6_n90, npu_inst_pe_1_5_6_n89, npu_inst_pe_1_5_6_n88,
         npu_inst_pe_1_5_6_n87, npu_inst_pe_1_5_6_n86, npu_inst_pe_1_5_6_n85,
         npu_inst_pe_1_5_6_n84, npu_inst_pe_1_5_6_n83, npu_inst_pe_1_5_6_n82,
         npu_inst_pe_1_5_6_n81, npu_inst_pe_1_5_6_n80, npu_inst_pe_1_5_6_n79,
         npu_inst_pe_1_5_6_n78, npu_inst_pe_1_5_6_n77, npu_inst_pe_1_5_6_n76,
         npu_inst_pe_1_5_6_n75, npu_inst_pe_1_5_6_n74, npu_inst_pe_1_5_6_n73,
         npu_inst_pe_1_5_6_n72, npu_inst_pe_1_5_6_n71, npu_inst_pe_1_5_6_n70,
         npu_inst_pe_1_5_6_n69, npu_inst_pe_1_5_6_n68, npu_inst_pe_1_5_6_n67,
         npu_inst_pe_1_5_6_n66, npu_inst_pe_1_5_6_n65, npu_inst_pe_1_5_6_n64,
         npu_inst_pe_1_5_6_n63, npu_inst_pe_1_5_6_n62, npu_inst_pe_1_5_6_n61,
         npu_inst_pe_1_5_6_n60, npu_inst_pe_1_5_6_n59, npu_inst_pe_1_5_6_n58,
         npu_inst_pe_1_5_6_n57, npu_inst_pe_1_5_6_n56, npu_inst_pe_1_5_6_n55,
         npu_inst_pe_1_5_6_n54, npu_inst_pe_1_5_6_n53, npu_inst_pe_1_5_6_n52,
         npu_inst_pe_1_5_6_n51, npu_inst_pe_1_5_6_n50, npu_inst_pe_1_5_6_n49,
         npu_inst_pe_1_5_6_n48, npu_inst_pe_1_5_6_n47, npu_inst_pe_1_5_6_n46,
         npu_inst_pe_1_5_6_n45, npu_inst_pe_1_5_6_n44, npu_inst_pe_1_5_6_n43,
         npu_inst_pe_1_5_6_n42, npu_inst_pe_1_5_6_n41, npu_inst_pe_1_5_6_n40,
         npu_inst_pe_1_5_6_n39, npu_inst_pe_1_5_6_n38, npu_inst_pe_1_5_6_n37,
         npu_inst_pe_1_5_6_n27, npu_inst_pe_1_5_6_n26,
         npu_inst_pe_1_5_6_net3510, npu_inst_pe_1_5_6_net3504,
         npu_inst_pe_1_5_6_N94, npu_inst_pe_1_5_6_N93, npu_inst_pe_1_5_6_N84,
         npu_inst_pe_1_5_6_N80, npu_inst_pe_1_5_6_N79, npu_inst_pe_1_5_6_N78,
         npu_inst_pe_1_5_6_N77, npu_inst_pe_1_5_6_N76, npu_inst_pe_1_5_6_N75,
         npu_inst_pe_1_5_6_N74, npu_inst_pe_1_5_6_N73, npu_inst_pe_1_5_6_N72,
         npu_inst_pe_1_5_6_N71, npu_inst_pe_1_5_6_N70, npu_inst_pe_1_5_6_N69,
         npu_inst_pe_1_5_6_N68, npu_inst_pe_1_5_6_N67, npu_inst_pe_1_5_6_N66,
         npu_inst_pe_1_5_6_N65, npu_inst_pe_1_5_6_int_q_acc_0_,
         npu_inst_pe_1_5_6_int_q_acc_1_, npu_inst_pe_1_5_6_int_q_acc_2_,
         npu_inst_pe_1_5_6_int_q_acc_3_, npu_inst_pe_1_5_6_int_q_acc_4_,
         npu_inst_pe_1_5_6_int_q_acc_5_, npu_inst_pe_1_5_6_int_q_acc_6_,
         npu_inst_pe_1_5_6_int_q_acc_7_, npu_inst_pe_1_5_6_int_data_0_,
         npu_inst_pe_1_5_6_int_data_1_, npu_inst_pe_1_5_6_int_q_weight_0_,
         npu_inst_pe_1_5_6_int_q_weight_1_,
         npu_inst_pe_1_5_6_int_q_reg_v_5__0_,
         npu_inst_pe_1_5_6_int_q_reg_v_5__1_,
         npu_inst_pe_1_5_6_int_q_reg_v_4__0_,
         npu_inst_pe_1_5_6_int_q_reg_v_4__1_,
         npu_inst_pe_1_5_6_int_q_reg_v_3__0_,
         npu_inst_pe_1_5_6_int_q_reg_v_3__1_,
         npu_inst_pe_1_5_6_int_q_reg_v_2__0_,
         npu_inst_pe_1_5_6_int_q_reg_v_2__1_,
         npu_inst_pe_1_5_6_int_q_reg_v_1__0_,
         npu_inst_pe_1_5_6_int_q_reg_v_1__1_,
         npu_inst_pe_1_5_6_int_q_reg_v_0__0_,
         npu_inst_pe_1_5_6_int_q_reg_v_0__1_,
         npu_inst_pe_1_5_6_int_q_reg_h_5__0_,
         npu_inst_pe_1_5_6_int_q_reg_h_5__1_,
         npu_inst_pe_1_5_6_int_q_reg_h_4__0_,
         npu_inst_pe_1_5_6_int_q_reg_h_4__1_,
         npu_inst_pe_1_5_6_int_q_reg_h_3__0_,
         npu_inst_pe_1_5_6_int_q_reg_h_3__1_,
         npu_inst_pe_1_5_6_int_q_reg_h_2__0_,
         npu_inst_pe_1_5_6_int_q_reg_h_2__1_,
         npu_inst_pe_1_5_6_int_q_reg_h_1__0_,
         npu_inst_pe_1_5_6_int_q_reg_h_1__1_,
         npu_inst_pe_1_5_6_int_q_reg_h_0__0_,
         npu_inst_pe_1_5_6_int_q_reg_h_0__1_, npu_inst_pe_1_5_7_n119,
         npu_inst_pe_1_5_7_n118, npu_inst_pe_1_5_7_n117,
         npu_inst_pe_1_5_7_n116, npu_inst_pe_1_5_7_n115,
         npu_inst_pe_1_5_7_n114, npu_inst_pe_1_5_7_n113,
         npu_inst_pe_1_5_7_n112, npu_inst_pe_1_5_7_n111,
         npu_inst_pe_1_5_7_n110, npu_inst_pe_1_5_7_n109,
         npu_inst_pe_1_5_7_n108, npu_inst_pe_1_5_7_n107,
         npu_inst_pe_1_5_7_n106, npu_inst_pe_1_5_7_n105,
         npu_inst_pe_1_5_7_n104, npu_inst_pe_1_5_7_n103,
         npu_inst_pe_1_5_7_n102, npu_inst_pe_1_5_7_n101,
         npu_inst_pe_1_5_7_n100, npu_inst_pe_1_5_7_n99, npu_inst_pe_1_5_7_n98,
         npu_inst_pe_1_5_7_n36, npu_inst_pe_1_5_7_n35, npu_inst_pe_1_5_7_n34,
         npu_inst_pe_1_5_7_n33, npu_inst_pe_1_5_7_n32, npu_inst_pe_1_5_7_n31,
         npu_inst_pe_1_5_7_n30, npu_inst_pe_1_5_7_n29, npu_inst_pe_1_5_7_n28,
         npu_inst_pe_1_5_7_n25, npu_inst_pe_1_5_7_n24, npu_inst_pe_1_5_7_n23,
         npu_inst_pe_1_5_7_n22, npu_inst_pe_1_5_7_n21, npu_inst_pe_1_5_7_n20,
         npu_inst_pe_1_5_7_n19, npu_inst_pe_1_5_7_n18, npu_inst_pe_1_5_7_n17,
         npu_inst_pe_1_5_7_n16, npu_inst_pe_1_5_7_n15, npu_inst_pe_1_5_7_n14,
         npu_inst_pe_1_5_7_n13, npu_inst_pe_1_5_7_n12, npu_inst_pe_1_5_7_n11,
         npu_inst_pe_1_5_7_n10, npu_inst_pe_1_5_7_n9, npu_inst_pe_1_5_7_n8,
         npu_inst_pe_1_5_7_n7, npu_inst_pe_1_5_7_n6, npu_inst_pe_1_5_7_n5,
         npu_inst_pe_1_5_7_n4, npu_inst_pe_1_5_7_n3, npu_inst_pe_1_5_7_n2,
         npu_inst_pe_1_5_7_n1, npu_inst_pe_1_5_7_sub_67_carry_7_,
         npu_inst_pe_1_5_7_sub_67_carry_6_, npu_inst_pe_1_5_7_sub_67_carry_5_,
         npu_inst_pe_1_5_7_sub_67_carry_4_, npu_inst_pe_1_5_7_sub_67_carry_3_,
         npu_inst_pe_1_5_7_sub_67_carry_2_, npu_inst_pe_1_5_7_sub_67_carry_1_,
         npu_inst_pe_1_5_7_add_69_carry_7_, npu_inst_pe_1_5_7_add_69_carry_6_,
         npu_inst_pe_1_5_7_add_69_carry_5_, npu_inst_pe_1_5_7_add_69_carry_4_,
         npu_inst_pe_1_5_7_add_69_carry_3_, npu_inst_pe_1_5_7_add_69_carry_2_,
         npu_inst_pe_1_5_7_add_69_carry_1_, npu_inst_pe_1_5_7_n97,
         npu_inst_pe_1_5_7_n96, npu_inst_pe_1_5_7_n95, npu_inst_pe_1_5_7_n94,
         npu_inst_pe_1_5_7_n93, npu_inst_pe_1_5_7_n92, npu_inst_pe_1_5_7_n91,
         npu_inst_pe_1_5_7_n90, npu_inst_pe_1_5_7_n89, npu_inst_pe_1_5_7_n88,
         npu_inst_pe_1_5_7_n87, npu_inst_pe_1_5_7_n86, npu_inst_pe_1_5_7_n85,
         npu_inst_pe_1_5_7_n84, npu_inst_pe_1_5_7_n83, npu_inst_pe_1_5_7_n82,
         npu_inst_pe_1_5_7_n81, npu_inst_pe_1_5_7_n80, npu_inst_pe_1_5_7_n79,
         npu_inst_pe_1_5_7_n78, npu_inst_pe_1_5_7_n77, npu_inst_pe_1_5_7_n76,
         npu_inst_pe_1_5_7_n75, npu_inst_pe_1_5_7_n74, npu_inst_pe_1_5_7_n73,
         npu_inst_pe_1_5_7_n72, npu_inst_pe_1_5_7_n71, npu_inst_pe_1_5_7_n70,
         npu_inst_pe_1_5_7_n69, npu_inst_pe_1_5_7_n68, npu_inst_pe_1_5_7_n67,
         npu_inst_pe_1_5_7_n66, npu_inst_pe_1_5_7_n65, npu_inst_pe_1_5_7_n64,
         npu_inst_pe_1_5_7_n63, npu_inst_pe_1_5_7_n62, npu_inst_pe_1_5_7_n61,
         npu_inst_pe_1_5_7_n60, npu_inst_pe_1_5_7_n59, npu_inst_pe_1_5_7_n58,
         npu_inst_pe_1_5_7_n57, npu_inst_pe_1_5_7_n56, npu_inst_pe_1_5_7_n55,
         npu_inst_pe_1_5_7_n54, npu_inst_pe_1_5_7_n53, npu_inst_pe_1_5_7_n52,
         npu_inst_pe_1_5_7_n51, npu_inst_pe_1_5_7_n50, npu_inst_pe_1_5_7_n49,
         npu_inst_pe_1_5_7_n48, npu_inst_pe_1_5_7_n47, npu_inst_pe_1_5_7_n46,
         npu_inst_pe_1_5_7_n45, npu_inst_pe_1_5_7_n44, npu_inst_pe_1_5_7_n43,
         npu_inst_pe_1_5_7_n42, npu_inst_pe_1_5_7_n41, npu_inst_pe_1_5_7_n40,
         npu_inst_pe_1_5_7_n39, npu_inst_pe_1_5_7_n38, npu_inst_pe_1_5_7_n37,
         npu_inst_pe_1_5_7_n27, npu_inst_pe_1_5_7_n26,
         npu_inst_pe_1_5_7_net3487, npu_inst_pe_1_5_7_net3481,
         npu_inst_pe_1_5_7_N94, npu_inst_pe_1_5_7_N93, npu_inst_pe_1_5_7_N84,
         npu_inst_pe_1_5_7_N80, npu_inst_pe_1_5_7_N79, npu_inst_pe_1_5_7_N78,
         npu_inst_pe_1_5_7_N77, npu_inst_pe_1_5_7_N76, npu_inst_pe_1_5_7_N75,
         npu_inst_pe_1_5_7_N74, npu_inst_pe_1_5_7_N73, npu_inst_pe_1_5_7_N72,
         npu_inst_pe_1_5_7_N71, npu_inst_pe_1_5_7_N70, npu_inst_pe_1_5_7_N69,
         npu_inst_pe_1_5_7_N68, npu_inst_pe_1_5_7_N67, npu_inst_pe_1_5_7_N66,
         npu_inst_pe_1_5_7_N65, npu_inst_pe_1_5_7_int_q_acc_0_,
         npu_inst_pe_1_5_7_int_q_acc_1_, npu_inst_pe_1_5_7_int_q_acc_2_,
         npu_inst_pe_1_5_7_int_q_acc_3_, npu_inst_pe_1_5_7_int_q_acc_4_,
         npu_inst_pe_1_5_7_int_q_acc_5_, npu_inst_pe_1_5_7_int_q_acc_6_,
         npu_inst_pe_1_5_7_int_q_acc_7_, npu_inst_pe_1_5_7_int_data_0_,
         npu_inst_pe_1_5_7_int_data_1_, npu_inst_pe_1_5_7_int_q_weight_0_,
         npu_inst_pe_1_5_7_int_q_weight_1_,
         npu_inst_pe_1_5_7_int_q_reg_v_5__0_,
         npu_inst_pe_1_5_7_int_q_reg_v_5__1_,
         npu_inst_pe_1_5_7_int_q_reg_v_4__0_,
         npu_inst_pe_1_5_7_int_q_reg_v_4__1_,
         npu_inst_pe_1_5_7_int_q_reg_v_3__0_,
         npu_inst_pe_1_5_7_int_q_reg_v_3__1_,
         npu_inst_pe_1_5_7_int_q_reg_v_2__0_,
         npu_inst_pe_1_5_7_int_q_reg_v_2__1_,
         npu_inst_pe_1_5_7_int_q_reg_v_1__0_,
         npu_inst_pe_1_5_7_int_q_reg_v_1__1_,
         npu_inst_pe_1_5_7_int_q_reg_v_0__0_,
         npu_inst_pe_1_5_7_int_q_reg_v_0__1_,
         npu_inst_pe_1_5_7_int_q_reg_h_5__0_,
         npu_inst_pe_1_5_7_int_q_reg_h_5__1_,
         npu_inst_pe_1_5_7_int_q_reg_h_4__0_,
         npu_inst_pe_1_5_7_int_q_reg_h_4__1_,
         npu_inst_pe_1_5_7_int_q_reg_h_3__0_,
         npu_inst_pe_1_5_7_int_q_reg_h_3__1_,
         npu_inst_pe_1_5_7_int_q_reg_h_2__0_,
         npu_inst_pe_1_5_7_int_q_reg_h_2__1_,
         npu_inst_pe_1_5_7_int_q_reg_h_1__0_,
         npu_inst_pe_1_5_7_int_q_reg_h_1__1_,
         npu_inst_pe_1_5_7_int_q_reg_h_0__0_,
         npu_inst_pe_1_5_7_int_q_reg_h_0__1_, npu_inst_pe_1_6_0_n119,
         npu_inst_pe_1_6_0_n118, npu_inst_pe_1_6_0_n117,
         npu_inst_pe_1_6_0_n116, npu_inst_pe_1_6_0_n115,
         npu_inst_pe_1_6_0_n114, npu_inst_pe_1_6_0_n113,
         npu_inst_pe_1_6_0_n112, npu_inst_pe_1_6_0_n111,
         npu_inst_pe_1_6_0_n110, npu_inst_pe_1_6_0_n109,
         npu_inst_pe_1_6_0_n108, npu_inst_pe_1_6_0_n107,
         npu_inst_pe_1_6_0_n106, npu_inst_pe_1_6_0_n105,
         npu_inst_pe_1_6_0_n104, npu_inst_pe_1_6_0_n103,
         npu_inst_pe_1_6_0_n102, npu_inst_pe_1_6_0_n101,
         npu_inst_pe_1_6_0_n100, npu_inst_pe_1_6_0_n99, npu_inst_pe_1_6_0_n98,
         npu_inst_pe_1_6_0_n36, npu_inst_pe_1_6_0_n35, npu_inst_pe_1_6_0_n34,
         npu_inst_pe_1_6_0_n33, npu_inst_pe_1_6_0_n32, npu_inst_pe_1_6_0_n31,
         npu_inst_pe_1_6_0_n30, npu_inst_pe_1_6_0_n29, npu_inst_pe_1_6_0_n28,
         npu_inst_pe_1_6_0_n25, npu_inst_pe_1_6_0_n24, npu_inst_pe_1_6_0_n23,
         npu_inst_pe_1_6_0_n22, npu_inst_pe_1_6_0_n21, npu_inst_pe_1_6_0_n20,
         npu_inst_pe_1_6_0_n19, npu_inst_pe_1_6_0_n18, npu_inst_pe_1_6_0_n17,
         npu_inst_pe_1_6_0_n16, npu_inst_pe_1_6_0_n15, npu_inst_pe_1_6_0_n14,
         npu_inst_pe_1_6_0_n13, npu_inst_pe_1_6_0_n12, npu_inst_pe_1_6_0_n11,
         npu_inst_pe_1_6_0_n10, npu_inst_pe_1_6_0_n9, npu_inst_pe_1_6_0_n8,
         npu_inst_pe_1_6_0_n7, npu_inst_pe_1_6_0_n6, npu_inst_pe_1_6_0_n5,
         npu_inst_pe_1_6_0_n4, npu_inst_pe_1_6_0_n3, npu_inst_pe_1_6_0_n2,
         npu_inst_pe_1_6_0_n1, npu_inst_pe_1_6_0_sub_67_carry_7_,
         npu_inst_pe_1_6_0_sub_67_carry_6_, npu_inst_pe_1_6_0_sub_67_carry_5_,
         npu_inst_pe_1_6_0_sub_67_carry_4_, npu_inst_pe_1_6_0_sub_67_carry_3_,
         npu_inst_pe_1_6_0_sub_67_carry_2_, npu_inst_pe_1_6_0_sub_67_carry_1_,
         npu_inst_pe_1_6_0_add_69_carry_7_, npu_inst_pe_1_6_0_add_69_carry_6_,
         npu_inst_pe_1_6_0_add_69_carry_5_, npu_inst_pe_1_6_0_add_69_carry_4_,
         npu_inst_pe_1_6_0_add_69_carry_3_, npu_inst_pe_1_6_0_add_69_carry_2_,
         npu_inst_pe_1_6_0_add_69_carry_1_, npu_inst_pe_1_6_0_n97,
         npu_inst_pe_1_6_0_n96, npu_inst_pe_1_6_0_n95, npu_inst_pe_1_6_0_n94,
         npu_inst_pe_1_6_0_n93, npu_inst_pe_1_6_0_n92, npu_inst_pe_1_6_0_n91,
         npu_inst_pe_1_6_0_n90, npu_inst_pe_1_6_0_n89, npu_inst_pe_1_6_0_n88,
         npu_inst_pe_1_6_0_n87, npu_inst_pe_1_6_0_n86, npu_inst_pe_1_6_0_n85,
         npu_inst_pe_1_6_0_n84, npu_inst_pe_1_6_0_n83, npu_inst_pe_1_6_0_n82,
         npu_inst_pe_1_6_0_n81, npu_inst_pe_1_6_0_n80, npu_inst_pe_1_6_0_n79,
         npu_inst_pe_1_6_0_n78, npu_inst_pe_1_6_0_n77, npu_inst_pe_1_6_0_n76,
         npu_inst_pe_1_6_0_n75, npu_inst_pe_1_6_0_n74, npu_inst_pe_1_6_0_n73,
         npu_inst_pe_1_6_0_n72, npu_inst_pe_1_6_0_n71, npu_inst_pe_1_6_0_n70,
         npu_inst_pe_1_6_0_n69, npu_inst_pe_1_6_0_n68, npu_inst_pe_1_6_0_n67,
         npu_inst_pe_1_6_0_n66, npu_inst_pe_1_6_0_n65, npu_inst_pe_1_6_0_n64,
         npu_inst_pe_1_6_0_n63, npu_inst_pe_1_6_0_n62, npu_inst_pe_1_6_0_n61,
         npu_inst_pe_1_6_0_n60, npu_inst_pe_1_6_0_n59, npu_inst_pe_1_6_0_n58,
         npu_inst_pe_1_6_0_n57, npu_inst_pe_1_6_0_n56, npu_inst_pe_1_6_0_n55,
         npu_inst_pe_1_6_0_n54, npu_inst_pe_1_6_0_n53, npu_inst_pe_1_6_0_n52,
         npu_inst_pe_1_6_0_n51, npu_inst_pe_1_6_0_n50, npu_inst_pe_1_6_0_n49,
         npu_inst_pe_1_6_0_n48, npu_inst_pe_1_6_0_n47, npu_inst_pe_1_6_0_n46,
         npu_inst_pe_1_6_0_n45, npu_inst_pe_1_6_0_n44, npu_inst_pe_1_6_0_n43,
         npu_inst_pe_1_6_0_n42, npu_inst_pe_1_6_0_n41, npu_inst_pe_1_6_0_n40,
         npu_inst_pe_1_6_0_n39, npu_inst_pe_1_6_0_n38, npu_inst_pe_1_6_0_n37,
         npu_inst_pe_1_6_0_n27, npu_inst_pe_1_6_0_n26,
         npu_inst_pe_1_6_0_net3464, npu_inst_pe_1_6_0_net3458,
         npu_inst_pe_1_6_0_N94, npu_inst_pe_1_6_0_N93, npu_inst_pe_1_6_0_N84,
         npu_inst_pe_1_6_0_N80, npu_inst_pe_1_6_0_N79, npu_inst_pe_1_6_0_N78,
         npu_inst_pe_1_6_0_N77, npu_inst_pe_1_6_0_N76, npu_inst_pe_1_6_0_N75,
         npu_inst_pe_1_6_0_N74, npu_inst_pe_1_6_0_N73, npu_inst_pe_1_6_0_N72,
         npu_inst_pe_1_6_0_N71, npu_inst_pe_1_6_0_N70, npu_inst_pe_1_6_0_N69,
         npu_inst_pe_1_6_0_N68, npu_inst_pe_1_6_0_N67, npu_inst_pe_1_6_0_N66,
         npu_inst_pe_1_6_0_N65, npu_inst_pe_1_6_0_int_q_acc_0_,
         npu_inst_pe_1_6_0_int_q_acc_1_, npu_inst_pe_1_6_0_int_q_acc_2_,
         npu_inst_pe_1_6_0_int_q_acc_3_, npu_inst_pe_1_6_0_int_q_acc_4_,
         npu_inst_pe_1_6_0_int_q_acc_5_, npu_inst_pe_1_6_0_int_q_acc_6_,
         npu_inst_pe_1_6_0_int_q_acc_7_, npu_inst_pe_1_6_0_int_data_0_,
         npu_inst_pe_1_6_0_int_data_1_, npu_inst_pe_1_6_0_int_q_weight_0_,
         npu_inst_pe_1_6_0_int_q_weight_1_,
         npu_inst_pe_1_6_0_int_q_reg_v_5__0_,
         npu_inst_pe_1_6_0_int_q_reg_v_5__1_,
         npu_inst_pe_1_6_0_int_q_reg_v_4__0_,
         npu_inst_pe_1_6_0_int_q_reg_v_4__1_,
         npu_inst_pe_1_6_0_int_q_reg_v_3__0_,
         npu_inst_pe_1_6_0_int_q_reg_v_3__1_,
         npu_inst_pe_1_6_0_int_q_reg_v_2__0_,
         npu_inst_pe_1_6_0_int_q_reg_v_2__1_,
         npu_inst_pe_1_6_0_int_q_reg_v_1__0_,
         npu_inst_pe_1_6_0_int_q_reg_v_1__1_,
         npu_inst_pe_1_6_0_int_q_reg_v_0__0_,
         npu_inst_pe_1_6_0_int_q_reg_v_0__1_,
         npu_inst_pe_1_6_0_int_q_reg_h_5__0_,
         npu_inst_pe_1_6_0_int_q_reg_h_5__1_,
         npu_inst_pe_1_6_0_int_q_reg_h_4__0_,
         npu_inst_pe_1_6_0_int_q_reg_h_4__1_,
         npu_inst_pe_1_6_0_int_q_reg_h_3__0_,
         npu_inst_pe_1_6_0_int_q_reg_h_3__1_,
         npu_inst_pe_1_6_0_int_q_reg_h_2__0_,
         npu_inst_pe_1_6_0_int_q_reg_h_2__1_,
         npu_inst_pe_1_6_0_int_q_reg_h_1__0_,
         npu_inst_pe_1_6_0_int_q_reg_h_1__1_,
         npu_inst_pe_1_6_0_int_q_reg_h_0__0_,
         npu_inst_pe_1_6_0_int_q_reg_h_0__1_, npu_inst_pe_1_6_0_o_data_h_0_,
         npu_inst_pe_1_6_0_o_data_h_1_, npu_inst_pe_1_6_1_n119,
         npu_inst_pe_1_6_1_n118, npu_inst_pe_1_6_1_n117,
         npu_inst_pe_1_6_1_n116, npu_inst_pe_1_6_1_n115,
         npu_inst_pe_1_6_1_n114, npu_inst_pe_1_6_1_n113,
         npu_inst_pe_1_6_1_n112, npu_inst_pe_1_6_1_n111,
         npu_inst_pe_1_6_1_n110, npu_inst_pe_1_6_1_n109,
         npu_inst_pe_1_6_1_n108, npu_inst_pe_1_6_1_n107,
         npu_inst_pe_1_6_1_n106, npu_inst_pe_1_6_1_n105,
         npu_inst_pe_1_6_1_n104, npu_inst_pe_1_6_1_n103,
         npu_inst_pe_1_6_1_n102, npu_inst_pe_1_6_1_n101,
         npu_inst_pe_1_6_1_n100, npu_inst_pe_1_6_1_n99, npu_inst_pe_1_6_1_n98,
         npu_inst_pe_1_6_1_n36, npu_inst_pe_1_6_1_n35, npu_inst_pe_1_6_1_n34,
         npu_inst_pe_1_6_1_n33, npu_inst_pe_1_6_1_n32, npu_inst_pe_1_6_1_n31,
         npu_inst_pe_1_6_1_n30, npu_inst_pe_1_6_1_n29, npu_inst_pe_1_6_1_n28,
         npu_inst_pe_1_6_1_n25, npu_inst_pe_1_6_1_n24, npu_inst_pe_1_6_1_n23,
         npu_inst_pe_1_6_1_n22, npu_inst_pe_1_6_1_n21, npu_inst_pe_1_6_1_n20,
         npu_inst_pe_1_6_1_n19, npu_inst_pe_1_6_1_n18, npu_inst_pe_1_6_1_n17,
         npu_inst_pe_1_6_1_n16, npu_inst_pe_1_6_1_n15, npu_inst_pe_1_6_1_n14,
         npu_inst_pe_1_6_1_n13, npu_inst_pe_1_6_1_n12, npu_inst_pe_1_6_1_n11,
         npu_inst_pe_1_6_1_n10, npu_inst_pe_1_6_1_n9, npu_inst_pe_1_6_1_n8,
         npu_inst_pe_1_6_1_n7, npu_inst_pe_1_6_1_n6, npu_inst_pe_1_6_1_n5,
         npu_inst_pe_1_6_1_n4, npu_inst_pe_1_6_1_n3, npu_inst_pe_1_6_1_n2,
         npu_inst_pe_1_6_1_n1, npu_inst_pe_1_6_1_sub_67_carry_7_,
         npu_inst_pe_1_6_1_sub_67_carry_6_, npu_inst_pe_1_6_1_sub_67_carry_5_,
         npu_inst_pe_1_6_1_sub_67_carry_4_, npu_inst_pe_1_6_1_sub_67_carry_3_,
         npu_inst_pe_1_6_1_sub_67_carry_2_, npu_inst_pe_1_6_1_sub_67_carry_1_,
         npu_inst_pe_1_6_1_add_69_carry_7_, npu_inst_pe_1_6_1_add_69_carry_6_,
         npu_inst_pe_1_6_1_add_69_carry_5_, npu_inst_pe_1_6_1_add_69_carry_4_,
         npu_inst_pe_1_6_1_add_69_carry_3_, npu_inst_pe_1_6_1_add_69_carry_2_,
         npu_inst_pe_1_6_1_add_69_carry_1_, npu_inst_pe_1_6_1_n97,
         npu_inst_pe_1_6_1_n96, npu_inst_pe_1_6_1_n95, npu_inst_pe_1_6_1_n94,
         npu_inst_pe_1_6_1_n93, npu_inst_pe_1_6_1_n92, npu_inst_pe_1_6_1_n91,
         npu_inst_pe_1_6_1_n90, npu_inst_pe_1_6_1_n89, npu_inst_pe_1_6_1_n88,
         npu_inst_pe_1_6_1_n87, npu_inst_pe_1_6_1_n86, npu_inst_pe_1_6_1_n85,
         npu_inst_pe_1_6_1_n84, npu_inst_pe_1_6_1_n83, npu_inst_pe_1_6_1_n82,
         npu_inst_pe_1_6_1_n81, npu_inst_pe_1_6_1_n80, npu_inst_pe_1_6_1_n79,
         npu_inst_pe_1_6_1_n78, npu_inst_pe_1_6_1_n77, npu_inst_pe_1_6_1_n76,
         npu_inst_pe_1_6_1_n75, npu_inst_pe_1_6_1_n74, npu_inst_pe_1_6_1_n73,
         npu_inst_pe_1_6_1_n72, npu_inst_pe_1_6_1_n71, npu_inst_pe_1_6_1_n70,
         npu_inst_pe_1_6_1_n69, npu_inst_pe_1_6_1_n68, npu_inst_pe_1_6_1_n67,
         npu_inst_pe_1_6_1_n66, npu_inst_pe_1_6_1_n65, npu_inst_pe_1_6_1_n64,
         npu_inst_pe_1_6_1_n63, npu_inst_pe_1_6_1_n62, npu_inst_pe_1_6_1_n61,
         npu_inst_pe_1_6_1_n60, npu_inst_pe_1_6_1_n59, npu_inst_pe_1_6_1_n58,
         npu_inst_pe_1_6_1_n57, npu_inst_pe_1_6_1_n56, npu_inst_pe_1_6_1_n55,
         npu_inst_pe_1_6_1_n54, npu_inst_pe_1_6_1_n53, npu_inst_pe_1_6_1_n52,
         npu_inst_pe_1_6_1_n51, npu_inst_pe_1_6_1_n50, npu_inst_pe_1_6_1_n49,
         npu_inst_pe_1_6_1_n48, npu_inst_pe_1_6_1_n47, npu_inst_pe_1_6_1_n46,
         npu_inst_pe_1_6_1_n45, npu_inst_pe_1_6_1_n44, npu_inst_pe_1_6_1_n43,
         npu_inst_pe_1_6_1_n42, npu_inst_pe_1_6_1_n41, npu_inst_pe_1_6_1_n40,
         npu_inst_pe_1_6_1_n39, npu_inst_pe_1_6_1_n38, npu_inst_pe_1_6_1_n37,
         npu_inst_pe_1_6_1_n27, npu_inst_pe_1_6_1_n26,
         npu_inst_pe_1_6_1_net3441, npu_inst_pe_1_6_1_net3435,
         npu_inst_pe_1_6_1_N94, npu_inst_pe_1_6_1_N93, npu_inst_pe_1_6_1_N84,
         npu_inst_pe_1_6_1_N80, npu_inst_pe_1_6_1_N79, npu_inst_pe_1_6_1_N78,
         npu_inst_pe_1_6_1_N77, npu_inst_pe_1_6_1_N76, npu_inst_pe_1_6_1_N75,
         npu_inst_pe_1_6_1_N74, npu_inst_pe_1_6_1_N73, npu_inst_pe_1_6_1_N72,
         npu_inst_pe_1_6_1_N71, npu_inst_pe_1_6_1_N70, npu_inst_pe_1_6_1_N69,
         npu_inst_pe_1_6_1_N68, npu_inst_pe_1_6_1_N67, npu_inst_pe_1_6_1_N66,
         npu_inst_pe_1_6_1_N65, npu_inst_pe_1_6_1_int_q_acc_0_,
         npu_inst_pe_1_6_1_int_q_acc_1_, npu_inst_pe_1_6_1_int_q_acc_2_,
         npu_inst_pe_1_6_1_int_q_acc_3_, npu_inst_pe_1_6_1_int_q_acc_4_,
         npu_inst_pe_1_6_1_int_q_acc_5_, npu_inst_pe_1_6_1_int_q_acc_6_,
         npu_inst_pe_1_6_1_int_q_acc_7_, npu_inst_pe_1_6_1_int_data_0_,
         npu_inst_pe_1_6_1_int_data_1_, npu_inst_pe_1_6_1_int_q_weight_0_,
         npu_inst_pe_1_6_1_int_q_weight_1_,
         npu_inst_pe_1_6_1_int_q_reg_v_5__0_,
         npu_inst_pe_1_6_1_int_q_reg_v_5__1_,
         npu_inst_pe_1_6_1_int_q_reg_v_4__0_,
         npu_inst_pe_1_6_1_int_q_reg_v_4__1_,
         npu_inst_pe_1_6_1_int_q_reg_v_3__0_,
         npu_inst_pe_1_6_1_int_q_reg_v_3__1_,
         npu_inst_pe_1_6_1_int_q_reg_v_2__0_,
         npu_inst_pe_1_6_1_int_q_reg_v_2__1_,
         npu_inst_pe_1_6_1_int_q_reg_v_1__0_,
         npu_inst_pe_1_6_1_int_q_reg_v_1__1_,
         npu_inst_pe_1_6_1_int_q_reg_v_0__0_,
         npu_inst_pe_1_6_1_int_q_reg_v_0__1_,
         npu_inst_pe_1_6_1_int_q_reg_h_5__0_,
         npu_inst_pe_1_6_1_int_q_reg_h_5__1_,
         npu_inst_pe_1_6_1_int_q_reg_h_4__0_,
         npu_inst_pe_1_6_1_int_q_reg_h_4__1_,
         npu_inst_pe_1_6_1_int_q_reg_h_3__0_,
         npu_inst_pe_1_6_1_int_q_reg_h_3__1_,
         npu_inst_pe_1_6_1_int_q_reg_h_2__0_,
         npu_inst_pe_1_6_1_int_q_reg_h_2__1_,
         npu_inst_pe_1_6_1_int_q_reg_h_1__0_,
         npu_inst_pe_1_6_1_int_q_reg_h_1__1_,
         npu_inst_pe_1_6_1_int_q_reg_h_0__0_,
         npu_inst_pe_1_6_1_int_q_reg_h_0__1_, npu_inst_pe_1_6_2_n119,
         npu_inst_pe_1_6_2_n118, npu_inst_pe_1_6_2_n117,
         npu_inst_pe_1_6_2_n116, npu_inst_pe_1_6_2_n115,
         npu_inst_pe_1_6_2_n114, npu_inst_pe_1_6_2_n113,
         npu_inst_pe_1_6_2_n112, npu_inst_pe_1_6_2_n111,
         npu_inst_pe_1_6_2_n110, npu_inst_pe_1_6_2_n109,
         npu_inst_pe_1_6_2_n108, npu_inst_pe_1_6_2_n107,
         npu_inst_pe_1_6_2_n106, npu_inst_pe_1_6_2_n105,
         npu_inst_pe_1_6_2_n104, npu_inst_pe_1_6_2_n103,
         npu_inst_pe_1_6_2_n102, npu_inst_pe_1_6_2_n101,
         npu_inst_pe_1_6_2_n100, npu_inst_pe_1_6_2_n99, npu_inst_pe_1_6_2_n98,
         npu_inst_pe_1_6_2_n36, npu_inst_pe_1_6_2_n35, npu_inst_pe_1_6_2_n34,
         npu_inst_pe_1_6_2_n33, npu_inst_pe_1_6_2_n32, npu_inst_pe_1_6_2_n31,
         npu_inst_pe_1_6_2_n30, npu_inst_pe_1_6_2_n29, npu_inst_pe_1_6_2_n28,
         npu_inst_pe_1_6_2_n25, npu_inst_pe_1_6_2_n24, npu_inst_pe_1_6_2_n23,
         npu_inst_pe_1_6_2_n22, npu_inst_pe_1_6_2_n21, npu_inst_pe_1_6_2_n20,
         npu_inst_pe_1_6_2_n19, npu_inst_pe_1_6_2_n18, npu_inst_pe_1_6_2_n17,
         npu_inst_pe_1_6_2_n16, npu_inst_pe_1_6_2_n15, npu_inst_pe_1_6_2_n14,
         npu_inst_pe_1_6_2_n13, npu_inst_pe_1_6_2_n12, npu_inst_pe_1_6_2_n11,
         npu_inst_pe_1_6_2_n10, npu_inst_pe_1_6_2_n9, npu_inst_pe_1_6_2_n8,
         npu_inst_pe_1_6_2_n7, npu_inst_pe_1_6_2_n6, npu_inst_pe_1_6_2_n5,
         npu_inst_pe_1_6_2_n4, npu_inst_pe_1_6_2_n3, npu_inst_pe_1_6_2_n2,
         npu_inst_pe_1_6_2_n1, npu_inst_pe_1_6_2_sub_67_carry_7_,
         npu_inst_pe_1_6_2_sub_67_carry_6_, npu_inst_pe_1_6_2_sub_67_carry_5_,
         npu_inst_pe_1_6_2_sub_67_carry_4_, npu_inst_pe_1_6_2_sub_67_carry_3_,
         npu_inst_pe_1_6_2_sub_67_carry_2_, npu_inst_pe_1_6_2_sub_67_carry_1_,
         npu_inst_pe_1_6_2_add_69_carry_7_, npu_inst_pe_1_6_2_add_69_carry_6_,
         npu_inst_pe_1_6_2_add_69_carry_5_, npu_inst_pe_1_6_2_add_69_carry_4_,
         npu_inst_pe_1_6_2_add_69_carry_3_, npu_inst_pe_1_6_2_add_69_carry_2_,
         npu_inst_pe_1_6_2_add_69_carry_1_, npu_inst_pe_1_6_2_n97,
         npu_inst_pe_1_6_2_n96, npu_inst_pe_1_6_2_n95, npu_inst_pe_1_6_2_n94,
         npu_inst_pe_1_6_2_n93, npu_inst_pe_1_6_2_n92, npu_inst_pe_1_6_2_n91,
         npu_inst_pe_1_6_2_n90, npu_inst_pe_1_6_2_n89, npu_inst_pe_1_6_2_n88,
         npu_inst_pe_1_6_2_n87, npu_inst_pe_1_6_2_n86, npu_inst_pe_1_6_2_n85,
         npu_inst_pe_1_6_2_n84, npu_inst_pe_1_6_2_n83, npu_inst_pe_1_6_2_n82,
         npu_inst_pe_1_6_2_n81, npu_inst_pe_1_6_2_n80, npu_inst_pe_1_6_2_n79,
         npu_inst_pe_1_6_2_n78, npu_inst_pe_1_6_2_n77, npu_inst_pe_1_6_2_n76,
         npu_inst_pe_1_6_2_n75, npu_inst_pe_1_6_2_n74, npu_inst_pe_1_6_2_n73,
         npu_inst_pe_1_6_2_n72, npu_inst_pe_1_6_2_n71, npu_inst_pe_1_6_2_n70,
         npu_inst_pe_1_6_2_n69, npu_inst_pe_1_6_2_n68, npu_inst_pe_1_6_2_n67,
         npu_inst_pe_1_6_2_n66, npu_inst_pe_1_6_2_n65, npu_inst_pe_1_6_2_n64,
         npu_inst_pe_1_6_2_n63, npu_inst_pe_1_6_2_n62, npu_inst_pe_1_6_2_n61,
         npu_inst_pe_1_6_2_n60, npu_inst_pe_1_6_2_n59, npu_inst_pe_1_6_2_n58,
         npu_inst_pe_1_6_2_n57, npu_inst_pe_1_6_2_n56, npu_inst_pe_1_6_2_n55,
         npu_inst_pe_1_6_2_n54, npu_inst_pe_1_6_2_n53, npu_inst_pe_1_6_2_n52,
         npu_inst_pe_1_6_2_n51, npu_inst_pe_1_6_2_n50, npu_inst_pe_1_6_2_n49,
         npu_inst_pe_1_6_2_n48, npu_inst_pe_1_6_2_n47, npu_inst_pe_1_6_2_n46,
         npu_inst_pe_1_6_2_n45, npu_inst_pe_1_6_2_n44, npu_inst_pe_1_6_2_n43,
         npu_inst_pe_1_6_2_n42, npu_inst_pe_1_6_2_n41, npu_inst_pe_1_6_2_n40,
         npu_inst_pe_1_6_2_n39, npu_inst_pe_1_6_2_n38, npu_inst_pe_1_6_2_n37,
         npu_inst_pe_1_6_2_n27, npu_inst_pe_1_6_2_n26,
         npu_inst_pe_1_6_2_net3418, npu_inst_pe_1_6_2_net3412,
         npu_inst_pe_1_6_2_N94, npu_inst_pe_1_6_2_N93, npu_inst_pe_1_6_2_N84,
         npu_inst_pe_1_6_2_N80, npu_inst_pe_1_6_2_N79, npu_inst_pe_1_6_2_N78,
         npu_inst_pe_1_6_2_N77, npu_inst_pe_1_6_2_N76, npu_inst_pe_1_6_2_N75,
         npu_inst_pe_1_6_2_N74, npu_inst_pe_1_6_2_N73, npu_inst_pe_1_6_2_N72,
         npu_inst_pe_1_6_2_N71, npu_inst_pe_1_6_2_N70, npu_inst_pe_1_6_2_N69,
         npu_inst_pe_1_6_2_N68, npu_inst_pe_1_6_2_N67, npu_inst_pe_1_6_2_N66,
         npu_inst_pe_1_6_2_N65, npu_inst_pe_1_6_2_int_q_acc_0_,
         npu_inst_pe_1_6_2_int_q_acc_1_, npu_inst_pe_1_6_2_int_q_acc_2_,
         npu_inst_pe_1_6_2_int_q_acc_3_, npu_inst_pe_1_6_2_int_q_acc_4_,
         npu_inst_pe_1_6_2_int_q_acc_5_, npu_inst_pe_1_6_2_int_q_acc_6_,
         npu_inst_pe_1_6_2_int_q_acc_7_, npu_inst_pe_1_6_2_int_data_0_,
         npu_inst_pe_1_6_2_int_data_1_, npu_inst_pe_1_6_2_int_q_weight_0_,
         npu_inst_pe_1_6_2_int_q_weight_1_,
         npu_inst_pe_1_6_2_int_q_reg_v_5__0_,
         npu_inst_pe_1_6_2_int_q_reg_v_5__1_,
         npu_inst_pe_1_6_2_int_q_reg_v_4__0_,
         npu_inst_pe_1_6_2_int_q_reg_v_4__1_,
         npu_inst_pe_1_6_2_int_q_reg_v_3__0_,
         npu_inst_pe_1_6_2_int_q_reg_v_3__1_,
         npu_inst_pe_1_6_2_int_q_reg_v_2__0_,
         npu_inst_pe_1_6_2_int_q_reg_v_2__1_,
         npu_inst_pe_1_6_2_int_q_reg_v_1__0_,
         npu_inst_pe_1_6_2_int_q_reg_v_1__1_,
         npu_inst_pe_1_6_2_int_q_reg_v_0__0_,
         npu_inst_pe_1_6_2_int_q_reg_v_0__1_,
         npu_inst_pe_1_6_2_int_q_reg_h_5__0_,
         npu_inst_pe_1_6_2_int_q_reg_h_5__1_,
         npu_inst_pe_1_6_2_int_q_reg_h_4__0_,
         npu_inst_pe_1_6_2_int_q_reg_h_4__1_,
         npu_inst_pe_1_6_2_int_q_reg_h_3__0_,
         npu_inst_pe_1_6_2_int_q_reg_h_3__1_,
         npu_inst_pe_1_6_2_int_q_reg_h_2__0_,
         npu_inst_pe_1_6_2_int_q_reg_h_2__1_,
         npu_inst_pe_1_6_2_int_q_reg_h_1__0_,
         npu_inst_pe_1_6_2_int_q_reg_h_1__1_,
         npu_inst_pe_1_6_2_int_q_reg_h_0__0_,
         npu_inst_pe_1_6_2_int_q_reg_h_0__1_, npu_inst_pe_1_6_3_n119,
         npu_inst_pe_1_6_3_n118, npu_inst_pe_1_6_3_n117,
         npu_inst_pe_1_6_3_n116, npu_inst_pe_1_6_3_n115,
         npu_inst_pe_1_6_3_n114, npu_inst_pe_1_6_3_n113,
         npu_inst_pe_1_6_3_n112, npu_inst_pe_1_6_3_n111,
         npu_inst_pe_1_6_3_n110, npu_inst_pe_1_6_3_n109,
         npu_inst_pe_1_6_3_n108, npu_inst_pe_1_6_3_n107,
         npu_inst_pe_1_6_3_n106, npu_inst_pe_1_6_3_n105,
         npu_inst_pe_1_6_3_n104, npu_inst_pe_1_6_3_n103,
         npu_inst_pe_1_6_3_n102, npu_inst_pe_1_6_3_n101,
         npu_inst_pe_1_6_3_n100, npu_inst_pe_1_6_3_n99, npu_inst_pe_1_6_3_n98,
         npu_inst_pe_1_6_3_n36, npu_inst_pe_1_6_3_n35, npu_inst_pe_1_6_3_n34,
         npu_inst_pe_1_6_3_n33, npu_inst_pe_1_6_3_n32, npu_inst_pe_1_6_3_n31,
         npu_inst_pe_1_6_3_n30, npu_inst_pe_1_6_3_n29, npu_inst_pe_1_6_3_n28,
         npu_inst_pe_1_6_3_n25, npu_inst_pe_1_6_3_n24, npu_inst_pe_1_6_3_n23,
         npu_inst_pe_1_6_3_n22, npu_inst_pe_1_6_3_n21, npu_inst_pe_1_6_3_n20,
         npu_inst_pe_1_6_3_n19, npu_inst_pe_1_6_3_n18, npu_inst_pe_1_6_3_n17,
         npu_inst_pe_1_6_3_n16, npu_inst_pe_1_6_3_n15, npu_inst_pe_1_6_3_n14,
         npu_inst_pe_1_6_3_n13, npu_inst_pe_1_6_3_n12, npu_inst_pe_1_6_3_n11,
         npu_inst_pe_1_6_3_n10, npu_inst_pe_1_6_3_n9, npu_inst_pe_1_6_3_n8,
         npu_inst_pe_1_6_3_n7, npu_inst_pe_1_6_3_n6, npu_inst_pe_1_6_3_n5,
         npu_inst_pe_1_6_3_n4, npu_inst_pe_1_6_3_n3, npu_inst_pe_1_6_3_n2,
         npu_inst_pe_1_6_3_n1, npu_inst_pe_1_6_3_sub_67_carry_7_,
         npu_inst_pe_1_6_3_sub_67_carry_6_, npu_inst_pe_1_6_3_sub_67_carry_5_,
         npu_inst_pe_1_6_3_sub_67_carry_4_, npu_inst_pe_1_6_3_sub_67_carry_3_,
         npu_inst_pe_1_6_3_sub_67_carry_2_, npu_inst_pe_1_6_3_sub_67_carry_1_,
         npu_inst_pe_1_6_3_add_69_carry_7_, npu_inst_pe_1_6_3_add_69_carry_6_,
         npu_inst_pe_1_6_3_add_69_carry_5_, npu_inst_pe_1_6_3_add_69_carry_4_,
         npu_inst_pe_1_6_3_add_69_carry_3_, npu_inst_pe_1_6_3_add_69_carry_2_,
         npu_inst_pe_1_6_3_add_69_carry_1_, npu_inst_pe_1_6_3_n97,
         npu_inst_pe_1_6_3_n96, npu_inst_pe_1_6_3_n95, npu_inst_pe_1_6_3_n94,
         npu_inst_pe_1_6_3_n93, npu_inst_pe_1_6_3_n92, npu_inst_pe_1_6_3_n91,
         npu_inst_pe_1_6_3_n90, npu_inst_pe_1_6_3_n89, npu_inst_pe_1_6_3_n88,
         npu_inst_pe_1_6_3_n87, npu_inst_pe_1_6_3_n86, npu_inst_pe_1_6_3_n85,
         npu_inst_pe_1_6_3_n84, npu_inst_pe_1_6_3_n83, npu_inst_pe_1_6_3_n82,
         npu_inst_pe_1_6_3_n81, npu_inst_pe_1_6_3_n80, npu_inst_pe_1_6_3_n79,
         npu_inst_pe_1_6_3_n78, npu_inst_pe_1_6_3_n77, npu_inst_pe_1_6_3_n76,
         npu_inst_pe_1_6_3_n75, npu_inst_pe_1_6_3_n74, npu_inst_pe_1_6_3_n73,
         npu_inst_pe_1_6_3_n72, npu_inst_pe_1_6_3_n71, npu_inst_pe_1_6_3_n70,
         npu_inst_pe_1_6_3_n69, npu_inst_pe_1_6_3_n68, npu_inst_pe_1_6_3_n67,
         npu_inst_pe_1_6_3_n66, npu_inst_pe_1_6_3_n65, npu_inst_pe_1_6_3_n64,
         npu_inst_pe_1_6_3_n63, npu_inst_pe_1_6_3_n62, npu_inst_pe_1_6_3_n61,
         npu_inst_pe_1_6_3_n60, npu_inst_pe_1_6_3_n59, npu_inst_pe_1_6_3_n58,
         npu_inst_pe_1_6_3_n57, npu_inst_pe_1_6_3_n56, npu_inst_pe_1_6_3_n55,
         npu_inst_pe_1_6_3_n54, npu_inst_pe_1_6_3_n53, npu_inst_pe_1_6_3_n52,
         npu_inst_pe_1_6_3_n51, npu_inst_pe_1_6_3_n50, npu_inst_pe_1_6_3_n49,
         npu_inst_pe_1_6_3_n48, npu_inst_pe_1_6_3_n47, npu_inst_pe_1_6_3_n46,
         npu_inst_pe_1_6_3_n45, npu_inst_pe_1_6_3_n44, npu_inst_pe_1_6_3_n43,
         npu_inst_pe_1_6_3_n42, npu_inst_pe_1_6_3_n41, npu_inst_pe_1_6_3_n40,
         npu_inst_pe_1_6_3_n39, npu_inst_pe_1_6_3_n38, npu_inst_pe_1_6_3_n37,
         npu_inst_pe_1_6_3_n27, npu_inst_pe_1_6_3_n26,
         npu_inst_pe_1_6_3_net3395, npu_inst_pe_1_6_3_net3389,
         npu_inst_pe_1_6_3_N94, npu_inst_pe_1_6_3_N93, npu_inst_pe_1_6_3_N84,
         npu_inst_pe_1_6_3_N80, npu_inst_pe_1_6_3_N79, npu_inst_pe_1_6_3_N78,
         npu_inst_pe_1_6_3_N77, npu_inst_pe_1_6_3_N76, npu_inst_pe_1_6_3_N75,
         npu_inst_pe_1_6_3_N74, npu_inst_pe_1_6_3_N73, npu_inst_pe_1_6_3_N72,
         npu_inst_pe_1_6_3_N71, npu_inst_pe_1_6_3_N70, npu_inst_pe_1_6_3_N69,
         npu_inst_pe_1_6_3_N68, npu_inst_pe_1_6_3_N67, npu_inst_pe_1_6_3_N66,
         npu_inst_pe_1_6_3_N65, npu_inst_pe_1_6_3_int_q_acc_0_,
         npu_inst_pe_1_6_3_int_q_acc_1_, npu_inst_pe_1_6_3_int_q_acc_2_,
         npu_inst_pe_1_6_3_int_q_acc_3_, npu_inst_pe_1_6_3_int_q_acc_4_,
         npu_inst_pe_1_6_3_int_q_acc_5_, npu_inst_pe_1_6_3_int_q_acc_6_,
         npu_inst_pe_1_6_3_int_q_acc_7_, npu_inst_pe_1_6_3_int_data_0_,
         npu_inst_pe_1_6_3_int_data_1_, npu_inst_pe_1_6_3_int_q_weight_0_,
         npu_inst_pe_1_6_3_int_q_weight_1_,
         npu_inst_pe_1_6_3_int_q_reg_v_5__0_,
         npu_inst_pe_1_6_3_int_q_reg_v_5__1_,
         npu_inst_pe_1_6_3_int_q_reg_v_4__0_,
         npu_inst_pe_1_6_3_int_q_reg_v_4__1_,
         npu_inst_pe_1_6_3_int_q_reg_v_3__0_,
         npu_inst_pe_1_6_3_int_q_reg_v_3__1_,
         npu_inst_pe_1_6_3_int_q_reg_v_2__0_,
         npu_inst_pe_1_6_3_int_q_reg_v_2__1_,
         npu_inst_pe_1_6_3_int_q_reg_v_1__0_,
         npu_inst_pe_1_6_3_int_q_reg_v_1__1_,
         npu_inst_pe_1_6_3_int_q_reg_v_0__0_,
         npu_inst_pe_1_6_3_int_q_reg_v_0__1_,
         npu_inst_pe_1_6_3_int_q_reg_h_5__0_,
         npu_inst_pe_1_6_3_int_q_reg_h_5__1_,
         npu_inst_pe_1_6_3_int_q_reg_h_4__0_,
         npu_inst_pe_1_6_3_int_q_reg_h_4__1_,
         npu_inst_pe_1_6_3_int_q_reg_h_3__0_,
         npu_inst_pe_1_6_3_int_q_reg_h_3__1_,
         npu_inst_pe_1_6_3_int_q_reg_h_2__0_,
         npu_inst_pe_1_6_3_int_q_reg_h_2__1_,
         npu_inst_pe_1_6_3_int_q_reg_h_1__0_,
         npu_inst_pe_1_6_3_int_q_reg_h_1__1_,
         npu_inst_pe_1_6_3_int_q_reg_h_0__0_,
         npu_inst_pe_1_6_3_int_q_reg_h_0__1_, npu_inst_pe_1_6_4_n118,
         npu_inst_pe_1_6_4_n117, npu_inst_pe_1_6_4_n116,
         npu_inst_pe_1_6_4_n115, npu_inst_pe_1_6_4_n114,
         npu_inst_pe_1_6_4_n113, npu_inst_pe_1_6_4_n112,
         npu_inst_pe_1_6_4_n111, npu_inst_pe_1_6_4_n110,
         npu_inst_pe_1_6_4_n109, npu_inst_pe_1_6_4_n108,
         npu_inst_pe_1_6_4_n107, npu_inst_pe_1_6_4_n106,
         npu_inst_pe_1_6_4_n105, npu_inst_pe_1_6_4_n104,
         npu_inst_pe_1_6_4_n103, npu_inst_pe_1_6_4_n102,
         npu_inst_pe_1_6_4_n101, npu_inst_pe_1_6_4_n100, npu_inst_pe_1_6_4_n99,
         npu_inst_pe_1_6_4_n98, npu_inst_pe_1_6_4_n36, npu_inst_pe_1_6_4_n35,
         npu_inst_pe_1_6_4_n34, npu_inst_pe_1_6_4_n33, npu_inst_pe_1_6_4_n32,
         npu_inst_pe_1_6_4_n31, npu_inst_pe_1_6_4_n30, npu_inst_pe_1_6_4_n29,
         npu_inst_pe_1_6_4_n28, npu_inst_pe_1_6_4_n25, npu_inst_pe_1_6_4_n24,
         npu_inst_pe_1_6_4_n23, npu_inst_pe_1_6_4_n22, npu_inst_pe_1_6_4_n21,
         npu_inst_pe_1_6_4_n20, npu_inst_pe_1_6_4_n19, npu_inst_pe_1_6_4_n18,
         npu_inst_pe_1_6_4_n17, npu_inst_pe_1_6_4_n16, npu_inst_pe_1_6_4_n15,
         npu_inst_pe_1_6_4_n14, npu_inst_pe_1_6_4_n13, npu_inst_pe_1_6_4_n12,
         npu_inst_pe_1_6_4_n11, npu_inst_pe_1_6_4_n10, npu_inst_pe_1_6_4_n9,
         npu_inst_pe_1_6_4_n8, npu_inst_pe_1_6_4_n7, npu_inst_pe_1_6_4_n6,
         npu_inst_pe_1_6_4_n5, npu_inst_pe_1_6_4_n4, npu_inst_pe_1_6_4_n3,
         npu_inst_pe_1_6_4_n2, npu_inst_pe_1_6_4_n1,
         npu_inst_pe_1_6_4_sub_67_carry_7_, npu_inst_pe_1_6_4_sub_67_carry_6_,
         npu_inst_pe_1_6_4_sub_67_carry_5_, npu_inst_pe_1_6_4_sub_67_carry_4_,
         npu_inst_pe_1_6_4_sub_67_carry_3_, npu_inst_pe_1_6_4_sub_67_carry_2_,
         npu_inst_pe_1_6_4_sub_67_carry_1_, npu_inst_pe_1_6_4_add_69_carry_7_,
         npu_inst_pe_1_6_4_add_69_carry_6_, npu_inst_pe_1_6_4_add_69_carry_5_,
         npu_inst_pe_1_6_4_add_69_carry_4_, npu_inst_pe_1_6_4_add_69_carry_3_,
         npu_inst_pe_1_6_4_add_69_carry_2_, npu_inst_pe_1_6_4_add_69_carry_1_,
         npu_inst_pe_1_6_4_n97, npu_inst_pe_1_6_4_n96, npu_inst_pe_1_6_4_n95,
         npu_inst_pe_1_6_4_n94, npu_inst_pe_1_6_4_n93, npu_inst_pe_1_6_4_n92,
         npu_inst_pe_1_6_4_n91, npu_inst_pe_1_6_4_n90, npu_inst_pe_1_6_4_n89,
         npu_inst_pe_1_6_4_n88, npu_inst_pe_1_6_4_n87, npu_inst_pe_1_6_4_n86,
         npu_inst_pe_1_6_4_n85, npu_inst_pe_1_6_4_n84, npu_inst_pe_1_6_4_n83,
         npu_inst_pe_1_6_4_n82, npu_inst_pe_1_6_4_n81, npu_inst_pe_1_6_4_n80,
         npu_inst_pe_1_6_4_n79, npu_inst_pe_1_6_4_n78, npu_inst_pe_1_6_4_n77,
         npu_inst_pe_1_6_4_n76, npu_inst_pe_1_6_4_n75, npu_inst_pe_1_6_4_n74,
         npu_inst_pe_1_6_4_n73, npu_inst_pe_1_6_4_n72, npu_inst_pe_1_6_4_n71,
         npu_inst_pe_1_6_4_n70, npu_inst_pe_1_6_4_n69, npu_inst_pe_1_6_4_n68,
         npu_inst_pe_1_6_4_n67, npu_inst_pe_1_6_4_n66, npu_inst_pe_1_6_4_n65,
         npu_inst_pe_1_6_4_n64, npu_inst_pe_1_6_4_n63, npu_inst_pe_1_6_4_n62,
         npu_inst_pe_1_6_4_n61, npu_inst_pe_1_6_4_n60, npu_inst_pe_1_6_4_n59,
         npu_inst_pe_1_6_4_n58, npu_inst_pe_1_6_4_n57, npu_inst_pe_1_6_4_n56,
         npu_inst_pe_1_6_4_n55, npu_inst_pe_1_6_4_n54, npu_inst_pe_1_6_4_n53,
         npu_inst_pe_1_6_4_n52, npu_inst_pe_1_6_4_n51, npu_inst_pe_1_6_4_n50,
         npu_inst_pe_1_6_4_n49, npu_inst_pe_1_6_4_n48, npu_inst_pe_1_6_4_n47,
         npu_inst_pe_1_6_4_n46, npu_inst_pe_1_6_4_n45, npu_inst_pe_1_6_4_n44,
         npu_inst_pe_1_6_4_n43, npu_inst_pe_1_6_4_n42, npu_inst_pe_1_6_4_n41,
         npu_inst_pe_1_6_4_n40, npu_inst_pe_1_6_4_n39, npu_inst_pe_1_6_4_n38,
         npu_inst_pe_1_6_4_n37, npu_inst_pe_1_6_4_n27, npu_inst_pe_1_6_4_n26,
         npu_inst_pe_1_6_4_net3372, npu_inst_pe_1_6_4_net3366,
         npu_inst_pe_1_6_4_N94, npu_inst_pe_1_6_4_N93, npu_inst_pe_1_6_4_N84,
         npu_inst_pe_1_6_4_N80, npu_inst_pe_1_6_4_N79, npu_inst_pe_1_6_4_N78,
         npu_inst_pe_1_6_4_N77, npu_inst_pe_1_6_4_N76, npu_inst_pe_1_6_4_N75,
         npu_inst_pe_1_6_4_N74, npu_inst_pe_1_6_4_N73, npu_inst_pe_1_6_4_N72,
         npu_inst_pe_1_6_4_N71, npu_inst_pe_1_6_4_N70, npu_inst_pe_1_6_4_N69,
         npu_inst_pe_1_6_4_N68, npu_inst_pe_1_6_4_N67, npu_inst_pe_1_6_4_N66,
         npu_inst_pe_1_6_4_N65, npu_inst_pe_1_6_4_int_q_acc_0_,
         npu_inst_pe_1_6_4_int_q_acc_1_, npu_inst_pe_1_6_4_int_q_acc_2_,
         npu_inst_pe_1_6_4_int_q_acc_3_, npu_inst_pe_1_6_4_int_q_acc_4_,
         npu_inst_pe_1_6_4_int_q_acc_5_, npu_inst_pe_1_6_4_int_q_acc_6_,
         npu_inst_pe_1_6_4_int_q_acc_7_, npu_inst_pe_1_6_4_int_data_0_,
         npu_inst_pe_1_6_4_int_data_1_, npu_inst_pe_1_6_4_int_q_weight_0_,
         npu_inst_pe_1_6_4_int_q_weight_1_,
         npu_inst_pe_1_6_4_int_q_reg_v_5__0_,
         npu_inst_pe_1_6_4_int_q_reg_v_5__1_,
         npu_inst_pe_1_6_4_int_q_reg_v_4__0_,
         npu_inst_pe_1_6_4_int_q_reg_v_4__1_,
         npu_inst_pe_1_6_4_int_q_reg_v_3__0_,
         npu_inst_pe_1_6_4_int_q_reg_v_3__1_,
         npu_inst_pe_1_6_4_int_q_reg_v_2__0_,
         npu_inst_pe_1_6_4_int_q_reg_v_2__1_,
         npu_inst_pe_1_6_4_int_q_reg_v_1__0_,
         npu_inst_pe_1_6_4_int_q_reg_v_1__1_,
         npu_inst_pe_1_6_4_int_q_reg_v_0__0_,
         npu_inst_pe_1_6_4_int_q_reg_v_0__1_,
         npu_inst_pe_1_6_4_int_q_reg_h_5__0_,
         npu_inst_pe_1_6_4_int_q_reg_h_5__1_,
         npu_inst_pe_1_6_4_int_q_reg_h_4__0_,
         npu_inst_pe_1_6_4_int_q_reg_h_4__1_,
         npu_inst_pe_1_6_4_int_q_reg_h_3__0_,
         npu_inst_pe_1_6_4_int_q_reg_h_3__1_,
         npu_inst_pe_1_6_4_int_q_reg_h_2__0_,
         npu_inst_pe_1_6_4_int_q_reg_h_2__1_,
         npu_inst_pe_1_6_4_int_q_reg_h_1__0_,
         npu_inst_pe_1_6_4_int_q_reg_h_1__1_,
         npu_inst_pe_1_6_4_int_q_reg_h_0__0_,
         npu_inst_pe_1_6_4_int_q_reg_h_0__1_, npu_inst_pe_1_6_5_n119,
         npu_inst_pe_1_6_5_n118, npu_inst_pe_1_6_5_n117,
         npu_inst_pe_1_6_5_n116, npu_inst_pe_1_6_5_n115,
         npu_inst_pe_1_6_5_n114, npu_inst_pe_1_6_5_n113,
         npu_inst_pe_1_6_5_n112, npu_inst_pe_1_6_5_n111,
         npu_inst_pe_1_6_5_n110, npu_inst_pe_1_6_5_n109,
         npu_inst_pe_1_6_5_n108, npu_inst_pe_1_6_5_n107,
         npu_inst_pe_1_6_5_n106, npu_inst_pe_1_6_5_n105,
         npu_inst_pe_1_6_5_n104, npu_inst_pe_1_6_5_n103,
         npu_inst_pe_1_6_5_n102, npu_inst_pe_1_6_5_n101,
         npu_inst_pe_1_6_5_n100, npu_inst_pe_1_6_5_n99, npu_inst_pe_1_6_5_n98,
         npu_inst_pe_1_6_5_n36, npu_inst_pe_1_6_5_n35, npu_inst_pe_1_6_5_n34,
         npu_inst_pe_1_6_5_n33, npu_inst_pe_1_6_5_n32, npu_inst_pe_1_6_5_n31,
         npu_inst_pe_1_6_5_n30, npu_inst_pe_1_6_5_n29, npu_inst_pe_1_6_5_n28,
         npu_inst_pe_1_6_5_n25, npu_inst_pe_1_6_5_n24, npu_inst_pe_1_6_5_n23,
         npu_inst_pe_1_6_5_n22, npu_inst_pe_1_6_5_n21, npu_inst_pe_1_6_5_n20,
         npu_inst_pe_1_6_5_n19, npu_inst_pe_1_6_5_n18, npu_inst_pe_1_6_5_n17,
         npu_inst_pe_1_6_5_n16, npu_inst_pe_1_6_5_n15, npu_inst_pe_1_6_5_n14,
         npu_inst_pe_1_6_5_n13, npu_inst_pe_1_6_5_n12, npu_inst_pe_1_6_5_n11,
         npu_inst_pe_1_6_5_n10, npu_inst_pe_1_6_5_n9, npu_inst_pe_1_6_5_n8,
         npu_inst_pe_1_6_5_n7, npu_inst_pe_1_6_5_n6, npu_inst_pe_1_6_5_n5,
         npu_inst_pe_1_6_5_n4, npu_inst_pe_1_6_5_n3, npu_inst_pe_1_6_5_n2,
         npu_inst_pe_1_6_5_n1, npu_inst_pe_1_6_5_sub_67_carry_7_,
         npu_inst_pe_1_6_5_sub_67_carry_6_, npu_inst_pe_1_6_5_sub_67_carry_5_,
         npu_inst_pe_1_6_5_sub_67_carry_4_, npu_inst_pe_1_6_5_sub_67_carry_3_,
         npu_inst_pe_1_6_5_sub_67_carry_2_, npu_inst_pe_1_6_5_sub_67_carry_1_,
         npu_inst_pe_1_6_5_add_69_carry_7_, npu_inst_pe_1_6_5_add_69_carry_6_,
         npu_inst_pe_1_6_5_add_69_carry_5_, npu_inst_pe_1_6_5_add_69_carry_4_,
         npu_inst_pe_1_6_5_add_69_carry_3_, npu_inst_pe_1_6_5_add_69_carry_2_,
         npu_inst_pe_1_6_5_add_69_carry_1_, npu_inst_pe_1_6_5_n97,
         npu_inst_pe_1_6_5_n96, npu_inst_pe_1_6_5_n95, npu_inst_pe_1_6_5_n94,
         npu_inst_pe_1_6_5_n93, npu_inst_pe_1_6_5_n92, npu_inst_pe_1_6_5_n91,
         npu_inst_pe_1_6_5_n90, npu_inst_pe_1_6_5_n89, npu_inst_pe_1_6_5_n88,
         npu_inst_pe_1_6_5_n87, npu_inst_pe_1_6_5_n86, npu_inst_pe_1_6_5_n85,
         npu_inst_pe_1_6_5_n84, npu_inst_pe_1_6_5_n83, npu_inst_pe_1_6_5_n82,
         npu_inst_pe_1_6_5_n81, npu_inst_pe_1_6_5_n80, npu_inst_pe_1_6_5_n79,
         npu_inst_pe_1_6_5_n78, npu_inst_pe_1_6_5_n77, npu_inst_pe_1_6_5_n76,
         npu_inst_pe_1_6_5_n75, npu_inst_pe_1_6_5_n74, npu_inst_pe_1_6_5_n73,
         npu_inst_pe_1_6_5_n72, npu_inst_pe_1_6_5_n71, npu_inst_pe_1_6_5_n70,
         npu_inst_pe_1_6_5_n69, npu_inst_pe_1_6_5_n68, npu_inst_pe_1_6_5_n67,
         npu_inst_pe_1_6_5_n66, npu_inst_pe_1_6_5_n65, npu_inst_pe_1_6_5_n64,
         npu_inst_pe_1_6_5_n63, npu_inst_pe_1_6_5_n62, npu_inst_pe_1_6_5_n61,
         npu_inst_pe_1_6_5_n60, npu_inst_pe_1_6_5_n59, npu_inst_pe_1_6_5_n58,
         npu_inst_pe_1_6_5_n57, npu_inst_pe_1_6_5_n56, npu_inst_pe_1_6_5_n55,
         npu_inst_pe_1_6_5_n54, npu_inst_pe_1_6_5_n53, npu_inst_pe_1_6_5_n52,
         npu_inst_pe_1_6_5_n51, npu_inst_pe_1_6_5_n50, npu_inst_pe_1_6_5_n49,
         npu_inst_pe_1_6_5_n48, npu_inst_pe_1_6_5_n47, npu_inst_pe_1_6_5_n46,
         npu_inst_pe_1_6_5_n45, npu_inst_pe_1_6_5_n44, npu_inst_pe_1_6_5_n43,
         npu_inst_pe_1_6_5_n42, npu_inst_pe_1_6_5_n41, npu_inst_pe_1_6_5_n40,
         npu_inst_pe_1_6_5_n39, npu_inst_pe_1_6_5_n38, npu_inst_pe_1_6_5_n37,
         npu_inst_pe_1_6_5_n27, npu_inst_pe_1_6_5_n26,
         npu_inst_pe_1_6_5_net3349, npu_inst_pe_1_6_5_net3343,
         npu_inst_pe_1_6_5_N94, npu_inst_pe_1_6_5_N93, npu_inst_pe_1_6_5_N84,
         npu_inst_pe_1_6_5_N80, npu_inst_pe_1_6_5_N79, npu_inst_pe_1_6_5_N78,
         npu_inst_pe_1_6_5_N77, npu_inst_pe_1_6_5_N76, npu_inst_pe_1_6_5_N75,
         npu_inst_pe_1_6_5_N74, npu_inst_pe_1_6_5_N73, npu_inst_pe_1_6_5_N72,
         npu_inst_pe_1_6_5_N71, npu_inst_pe_1_6_5_N70, npu_inst_pe_1_6_5_N69,
         npu_inst_pe_1_6_5_N68, npu_inst_pe_1_6_5_N67, npu_inst_pe_1_6_5_N66,
         npu_inst_pe_1_6_5_N65, npu_inst_pe_1_6_5_int_q_acc_0_,
         npu_inst_pe_1_6_5_int_q_acc_1_, npu_inst_pe_1_6_5_int_q_acc_2_,
         npu_inst_pe_1_6_5_int_q_acc_3_, npu_inst_pe_1_6_5_int_q_acc_4_,
         npu_inst_pe_1_6_5_int_q_acc_5_, npu_inst_pe_1_6_5_int_q_acc_6_,
         npu_inst_pe_1_6_5_int_q_acc_7_, npu_inst_pe_1_6_5_int_data_0_,
         npu_inst_pe_1_6_5_int_data_1_, npu_inst_pe_1_6_5_int_q_weight_0_,
         npu_inst_pe_1_6_5_int_q_weight_1_,
         npu_inst_pe_1_6_5_int_q_reg_v_5__0_,
         npu_inst_pe_1_6_5_int_q_reg_v_5__1_,
         npu_inst_pe_1_6_5_int_q_reg_v_4__0_,
         npu_inst_pe_1_6_5_int_q_reg_v_4__1_,
         npu_inst_pe_1_6_5_int_q_reg_v_3__0_,
         npu_inst_pe_1_6_5_int_q_reg_v_3__1_,
         npu_inst_pe_1_6_5_int_q_reg_v_2__0_,
         npu_inst_pe_1_6_5_int_q_reg_v_2__1_,
         npu_inst_pe_1_6_5_int_q_reg_v_1__0_,
         npu_inst_pe_1_6_5_int_q_reg_v_1__1_,
         npu_inst_pe_1_6_5_int_q_reg_v_0__0_,
         npu_inst_pe_1_6_5_int_q_reg_v_0__1_,
         npu_inst_pe_1_6_5_int_q_reg_h_5__0_,
         npu_inst_pe_1_6_5_int_q_reg_h_5__1_,
         npu_inst_pe_1_6_5_int_q_reg_h_4__0_,
         npu_inst_pe_1_6_5_int_q_reg_h_4__1_,
         npu_inst_pe_1_6_5_int_q_reg_h_3__0_,
         npu_inst_pe_1_6_5_int_q_reg_h_3__1_,
         npu_inst_pe_1_6_5_int_q_reg_h_2__0_,
         npu_inst_pe_1_6_5_int_q_reg_h_2__1_,
         npu_inst_pe_1_6_5_int_q_reg_h_1__0_,
         npu_inst_pe_1_6_5_int_q_reg_h_1__1_,
         npu_inst_pe_1_6_5_int_q_reg_h_0__0_,
         npu_inst_pe_1_6_5_int_q_reg_h_0__1_, npu_inst_pe_1_6_6_n119,
         npu_inst_pe_1_6_6_n118, npu_inst_pe_1_6_6_n117,
         npu_inst_pe_1_6_6_n116, npu_inst_pe_1_6_6_n115,
         npu_inst_pe_1_6_6_n114, npu_inst_pe_1_6_6_n113,
         npu_inst_pe_1_6_6_n112, npu_inst_pe_1_6_6_n111,
         npu_inst_pe_1_6_6_n110, npu_inst_pe_1_6_6_n109,
         npu_inst_pe_1_6_6_n108, npu_inst_pe_1_6_6_n107,
         npu_inst_pe_1_6_6_n106, npu_inst_pe_1_6_6_n105,
         npu_inst_pe_1_6_6_n104, npu_inst_pe_1_6_6_n103,
         npu_inst_pe_1_6_6_n102, npu_inst_pe_1_6_6_n101,
         npu_inst_pe_1_6_6_n100, npu_inst_pe_1_6_6_n99, npu_inst_pe_1_6_6_n98,
         npu_inst_pe_1_6_6_n36, npu_inst_pe_1_6_6_n35, npu_inst_pe_1_6_6_n34,
         npu_inst_pe_1_6_6_n33, npu_inst_pe_1_6_6_n32, npu_inst_pe_1_6_6_n31,
         npu_inst_pe_1_6_6_n30, npu_inst_pe_1_6_6_n29, npu_inst_pe_1_6_6_n28,
         npu_inst_pe_1_6_6_n25, npu_inst_pe_1_6_6_n24, npu_inst_pe_1_6_6_n23,
         npu_inst_pe_1_6_6_n22, npu_inst_pe_1_6_6_n21, npu_inst_pe_1_6_6_n20,
         npu_inst_pe_1_6_6_n19, npu_inst_pe_1_6_6_n18, npu_inst_pe_1_6_6_n17,
         npu_inst_pe_1_6_6_n16, npu_inst_pe_1_6_6_n15, npu_inst_pe_1_6_6_n14,
         npu_inst_pe_1_6_6_n13, npu_inst_pe_1_6_6_n12, npu_inst_pe_1_6_6_n11,
         npu_inst_pe_1_6_6_n10, npu_inst_pe_1_6_6_n9, npu_inst_pe_1_6_6_n8,
         npu_inst_pe_1_6_6_n7, npu_inst_pe_1_6_6_n6, npu_inst_pe_1_6_6_n5,
         npu_inst_pe_1_6_6_n4, npu_inst_pe_1_6_6_n3, npu_inst_pe_1_6_6_n2,
         npu_inst_pe_1_6_6_n1, npu_inst_pe_1_6_6_sub_67_carry_7_,
         npu_inst_pe_1_6_6_sub_67_carry_6_, npu_inst_pe_1_6_6_sub_67_carry_5_,
         npu_inst_pe_1_6_6_sub_67_carry_4_, npu_inst_pe_1_6_6_sub_67_carry_3_,
         npu_inst_pe_1_6_6_sub_67_carry_2_, npu_inst_pe_1_6_6_sub_67_carry_1_,
         npu_inst_pe_1_6_6_add_69_carry_7_, npu_inst_pe_1_6_6_add_69_carry_6_,
         npu_inst_pe_1_6_6_add_69_carry_5_, npu_inst_pe_1_6_6_add_69_carry_4_,
         npu_inst_pe_1_6_6_add_69_carry_3_, npu_inst_pe_1_6_6_add_69_carry_2_,
         npu_inst_pe_1_6_6_add_69_carry_1_, npu_inst_pe_1_6_6_n97,
         npu_inst_pe_1_6_6_n96, npu_inst_pe_1_6_6_n95, npu_inst_pe_1_6_6_n94,
         npu_inst_pe_1_6_6_n93, npu_inst_pe_1_6_6_n92, npu_inst_pe_1_6_6_n91,
         npu_inst_pe_1_6_6_n90, npu_inst_pe_1_6_6_n89, npu_inst_pe_1_6_6_n88,
         npu_inst_pe_1_6_6_n87, npu_inst_pe_1_6_6_n86, npu_inst_pe_1_6_6_n85,
         npu_inst_pe_1_6_6_n84, npu_inst_pe_1_6_6_n83, npu_inst_pe_1_6_6_n82,
         npu_inst_pe_1_6_6_n81, npu_inst_pe_1_6_6_n80, npu_inst_pe_1_6_6_n79,
         npu_inst_pe_1_6_6_n78, npu_inst_pe_1_6_6_n77, npu_inst_pe_1_6_6_n76,
         npu_inst_pe_1_6_6_n75, npu_inst_pe_1_6_6_n74, npu_inst_pe_1_6_6_n73,
         npu_inst_pe_1_6_6_n72, npu_inst_pe_1_6_6_n71, npu_inst_pe_1_6_6_n70,
         npu_inst_pe_1_6_6_n69, npu_inst_pe_1_6_6_n68, npu_inst_pe_1_6_6_n67,
         npu_inst_pe_1_6_6_n66, npu_inst_pe_1_6_6_n65, npu_inst_pe_1_6_6_n64,
         npu_inst_pe_1_6_6_n63, npu_inst_pe_1_6_6_n62, npu_inst_pe_1_6_6_n61,
         npu_inst_pe_1_6_6_n60, npu_inst_pe_1_6_6_n59, npu_inst_pe_1_6_6_n58,
         npu_inst_pe_1_6_6_n57, npu_inst_pe_1_6_6_n56, npu_inst_pe_1_6_6_n55,
         npu_inst_pe_1_6_6_n54, npu_inst_pe_1_6_6_n53, npu_inst_pe_1_6_6_n52,
         npu_inst_pe_1_6_6_n51, npu_inst_pe_1_6_6_n50, npu_inst_pe_1_6_6_n49,
         npu_inst_pe_1_6_6_n48, npu_inst_pe_1_6_6_n47, npu_inst_pe_1_6_6_n46,
         npu_inst_pe_1_6_6_n45, npu_inst_pe_1_6_6_n44, npu_inst_pe_1_6_6_n43,
         npu_inst_pe_1_6_6_n42, npu_inst_pe_1_6_6_n41, npu_inst_pe_1_6_6_n40,
         npu_inst_pe_1_6_6_n39, npu_inst_pe_1_6_6_n38, npu_inst_pe_1_6_6_n37,
         npu_inst_pe_1_6_6_n27, npu_inst_pe_1_6_6_n26,
         npu_inst_pe_1_6_6_net3326, npu_inst_pe_1_6_6_net3320,
         npu_inst_pe_1_6_6_N94, npu_inst_pe_1_6_6_N93, npu_inst_pe_1_6_6_N84,
         npu_inst_pe_1_6_6_N80, npu_inst_pe_1_6_6_N79, npu_inst_pe_1_6_6_N78,
         npu_inst_pe_1_6_6_N77, npu_inst_pe_1_6_6_N76, npu_inst_pe_1_6_6_N75,
         npu_inst_pe_1_6_6_N74, npu_inst_pe_1_6_6_N73, npu_inst_pe_1_6_6_N72,
         npu_inst_pe_1_6_6_N71, npu_inst_pe_1_6_6_N70, npu_inst_pe_1_6_6_N69,
         npu_inst_pe_1_6_6_N68, npu_inst_pe_1_6_6_N67, npu_inst_pe_1_6_6_N66,
         npu_inst_pe_1_6_6_N65, npu_inst_pe_1_6_6_int_q_acc_0_,
         npu_inst_pe_1_6_6_int_q_acc_1_, npu_inst_pe_1_6_6_int_q_acc_2_,
         npu_inst_pe_1_6_6_int_q_acc_3_, npu_inst_pe_1_6_6_int_q_acc_4_,
         npu_inst_pe_1_6_6_int_q_acc_5_, npu_inst_pe_1_6_6_int_q_acc_6_,
         npu_inst_pe_1_6_6_int_q_acc_7_, npu_inst_pe_1_6_6_int_data_0_,
         npu_inst_pe_1_6_6_int_data_1_, npu_inst_pe_1_6_6_int_q_weight_0_,
         npu_inst_pe_1_6_6_int_q_weight_1_,
         npu_inst_pe_1_6_6_int_q_reg_v_5__0_,
         npu_inst_pe_1_6_6_int_q_reg_v_5__1_,
         npu_inst_pe_1_6_6_int_q_reg_v_4__0_,
         npu_inst_pe_1_6_6_int_q_reg_v_4__1_,
         npu_inst_pe_1_6_6_int_q_reg_v_3__0_,
         npu_inst_pe_1_6_6_int_q_reg_v_3__1_,
         npu_inst_pe_1_6_6_int_q_reg_v_2__0_,
         npu_inst_pe_1_6_6_int_q_reg_v_2__1_,
         npu_inst_pe_1_6_6_int_q_reg_v_1__0_,
         npu_inst_pe_1_6_6_int_q_reg_v_1__1_,
         npu_inst_pe_1_6_6_int_q_reg_v_0__0_,
         npu_inst_pe_1_6_6_int_q_reg_v_0__1_,
         npu_inst_pe_1_6_6_int_q_reg_h_5__0_,
         npu_inst_pe_1_6_6_int_q_reg_h_5__1_,
         npu_inst_pe_1_6_6_int_q_reg_h_4__0_,
         npu_inst_pe_1_6_6_int_q_reg_h_4__1_,
         npu_inst_pe_1_6_6_int_q_reg_h_3__0_,
         npu_inst_pe_1_6_6_int_q_reg_h_3__1_,
         npu_inst_pe_1_6_6_int_q_reg_h_2__0_,
         npu_inst_pe_1_6_6_int_q_reg_h_2__1_,
         npu_inst_pe_1_6_6_int_q_reg_h_1__0_,
         npu_inst_pe_1_6_6_int_q_reg_h_1__1_,
         npu_inst_pe_1_6_6_int_q_reg_h_0__0_,
         npu_inst_pe_1_6_6_int_q_reg_h_0__1_, npu_inst_pe_1_6_7_n119,
         npu_inst_pe_1_6_7_n118, npu_inst_pe_1_6_7_n117,
         npu_inst_pe_1_6_7_n116, npu_inst_pe_1_6_7_n115,
         npu_inst_pe_1_6_7_n114, npu_inst_pe_1_6_7_n113,
         npu_inst_pe_1_6_7_n112, npu_inst_pe_1_6_7_n111,
         npu_inst_pe_1_6_7_n110, npu_inst_pe_1_6_7_n109,
         npu_inst_pe_1_6_7_n108, npu_inst_pe_1_6_7_n107,
         npu_inst_pe_1_6_7_n106, npu_inst_pe_1_6_7_n105,
         npu_inst_pe_1_6_7_n104, npu_inst_pe_1_6_7_n103,
         npu_inst_pe_1_6_7_n102, npu_inst_pe_1_6_7_n101,
         npu_inst_pe_1_6_7_n100, npu_inst_pe_1_6_7_n99, npu_inst_pe_1_6_7_n98,
         npu_inst_pe_1_6_7_n36, npu_inst_pe_1_6_7_n35, npu_inst_pe_1_6_7_n34,
         npu_inst_pe_1_6_7_n33, npu_inst_pe_1_6_7_n32, npu_inst_pe_1_6_7_n31,
         npu_inst_pe_1_6_7_n30, npu_inst_pe_1_6_7_n29, npu_inst_pe_1_6_7_n28,
         npu_inst_pe_1_6_7_n25, npu_inst_pe_1_6_7_n24, npu_inst_pe_1_6_7_n23,
         npu_inst_pe_1_6_7_n22, npu_inst_pe_1_6_7_n21, npu_inst_pe_1_6_7_n20,
         npu_inst_pe_1_6_7_n19, npu_inst_pe_1_6_7_n18, npu_inst_pe_1_6_7_n17,
         npu_inst_pe_1_6_7_n16, npu_inst_pe_1_6_7_n15, npu_inst_pe_1_6_7_n14,
         npu_inst_pe_1_6_7_n13, npu_inst_pe_1_6_7_n12, npu_inst_pe_1_6_7_n11,
         npu_inst_pe_1_6_7_n10, npu_inst_pe_1_6_7_n9, npu_inst_pe_1_6_7_n8,
         npu_inst_pe_1_6_7_n7, npu_inst_pe_1_6_7_n6, npu_inst_pe_1_6_7_n5,
         npu_inst_pe_1_6_7_n4, npu_inst_pe_1_6_7_n3, npu_inst_pe_1_6_7_n2,
         npu_inst_pe_1_6_7_n1, npu_inst_pe_1_6_7_sub_67_carry_7_,
         npu_inst_pe_1_6_7_sub_67_carry_6_, npu_inst_pe_1_6_7_sub_67_carry_5_,
         npu_inst_pe_1_6_7_sub_67_carry_4_, npu_inst_pe_1_6_7_sub_67_carry_3_,
         npu_inst_pe_1_6_7_sub_67_carry_2_, npu_inst_pe_1_6_7_sub_67_carry_1_,
         npu_inst_pe_1_6_7_add_69_carry_7_, npu_inst_pe_1_6_7_add_69_carry_6_,
         npu_inst_pe_1_6_7_add_69_carry_5_, npu_inst_pe_1_6_7_add_69_carry_4_,
         npu_inst_pe_1_6_7_add_69_carry_3_, npu_inst_pe_1_6_7_add_69_carry_2_,
         npu_inst_pe_1_6_7_add_69_carry_1_, npu_inst_pe_1_6_7_n97,
         npu_inst_pe_1_6_7_n96, npu_inst_pe_1_6_7_n95, npu_inst_pe_1_6_7_n94,
         npu_inst_pe_1_6_7_n93, npu_inst_pe_1_6_7_n92, npu_inst_pe_1_6_7_n91,
         npu_inst_pe_1_6_7_n90, npu_inst_pe_1_6_7_n89, npu_inst_pe_1_6_7_n88,
         npu_inst_pe_1_6_7_n87, npu_inst_pe_1_6_7_n86, npu_inst_pe_1_6_7_n85,
         npu_inst_pe_1_6_7_n84, npu_inst_pe_1_6_7_n83, npu_inst_pe_1_6_7_n82,
         npu_inst_pe_1_6_7_n81, npu_inst_pe_1_6_7_n80, npu_inst_pe_1_6_7_n79,
         npu_inst_pe_1_6_7_n78, npu_inst_pe_1_6_7_n77, npu_inst_pe_1_6_7_n76,
         npu_inst_pe_1_6_7_n75, npu_inst_pe_1_6_7_n74, npu_inst_pe_1_6_7_n73,
         npu_inst_pe_1_6_7_n72, npu_inst_pe_1_6_7_n71, npu_inst_pe_1_6_7_n70,
         npu_inst_pe_1_6_7_n69, npu_inst_pe_1_6_7_n68, npu_inst_pe_1_6_7_n67,
         npu_inst_pe_1_6_7_n66, npu_inst_pe_1_6_7_n65, npu_inst_pe_1_6_7_n64,
         npu_inst_pe_1_6_7_n63, npu_inst_pe_1_6_7_n62, npu_inst_pe_1_6_7_n61,
         npu_inst_pe_1_6_7_n60, npu_inst_pe_1_6_7_n59, npu_inst_pe_1_6_7_n58,
         npu_inst_pe_1_6_7_n57, npu_inst_pe_1_6_7_n56, npu_inst_pe_1_6_7_n55,
         npu_inst_pe_1_6_7_n54, npu_inst_pe_1_6_7_n53, npu_inst_pe_1_6_7_n52,
         npu_inst_pe_1_6_7_n51, npu_inst_pe_1_6_7_n50, npu_inst_pe_1_6_7_n49,
         npu_inst_pe_1_6_7_n48, npu_inst_pe_1_6_7_n47, npu_inst_pe_1_6_7_n46,
         npu_inst_pe_1_6_7_n45, npu_inst_pe_1_6_7_n44, npu_inst_pe_1_6_7_n43,
         npu_inst_pe_1_6_7_n42, npu_inst_pe_1_6_7_n41, npu_inst_pe_1_6_7_n40,
         npu_inst_pe_1_6_7_n39, npu_inst_pe_1_6_7_n38, npu_inst_pe_1_6_7_n37,
         npu_inst_pe_1_6_7_n27, npu_inst_pe_1_6_7_n26,
         npu_inst_pe_1_6_7_net3303, npu_inst_pe_1_6_7_net3297,
         npu_inst_pe_1_6_7_N94, npu_inst_pe_1_6_7_N93, npu_inst_pe_1_6_7_N84,
         npu_inst_pe_1_6_7_N80, npu_inst_pe_1_6_7_N79, npu_inst_pe_1_6_7_N78,
         npu_inst_pe_1_6_7_N77, npu_inst_pe_1_6_7_N76, npu_inst_pe_1_6_7_N75,
         npu_inst_pe_1_6_7_N74, npu_inst_pe_1_6_7_N73, npu_inst_pe_1_6_7_N72,
         npu_inst_pe_1_6_7_N71, npu_inst_pe_1_6_7_N70, npu_inst_pe_1_6_7_N69,
         npu_inst_pe_1_6_7_N68, npu_inst_pe_1_6_7_N67, npu_inst_pe_1_6_7_N66,
         npu_inst_pe_1_6_7_N65, npu_inst_pe_1_6_7_int_q_acc_0_,
         npu_inst_pe_1_6_7_int_q_acc_1_, npu_inst_pe_1_6_7_int_q_acc_2_,
         npu_inst_pe_1_6_7_int_q_acc_3_, npu_inst_pe_1_6_7_int_q_acc_4_,
         npu_inst_pe_1_6_7_int_q_acc_5_, npu_inst_pe_1_6_7_int_q_acc_6_,
         npu_inst_pe_1_6_7_int_q_acc_7_, npu_inst_pe_1_6_7_int_data_0_,
         npu_inst_pe_1_6_7_int_data_1_, npu_inst_pe_1_6_7_int_q_weight_0_,
         npu_inst_pe_1_6_7_int_q_weight_1_,
         npu_inst_pe_1_6_7_int_q_reg_v_5__0_,
         npu_inst_pe_1_6_7_int_q_reg_v_5__1_,
         npu_inst_pe_1_6_7_int_q_reg_v_4__0_,
         npu_inst_pe_1_6_7_int_q_reg_v_4__1_,
         npu_inst_pe_1_6_7_int_q_reg_v_3__0_,
         npu_inst_pe_1_6_7_int_q_reg_v_3__1_,
         npu_inst_pe_1_6_7_int_q_reg_v_2__0_,
         npu_inst_pe_1_6_7_int_q_reg_v_2__1_,
         npu_inst_pe_1_6_7_int_q_reg_v_1__0_,
         npu_inst_pe_1_6_7_int_q_reg_v_1__1_,
         npu_inst_pe_1_6_7_int_q_reg_v_0__0_,
         npu_inst_pe_1_6_7_int_q_reg_v_0__1_,
         npu_inst_pe_1_6_7_int_q_reg_h_5__0_,
         npu_inst_pe_1_6_7_int_q_reg_h_5__1_,
         npu_inst_pe_1_6_7_int_q_reg_h_4__0_,
         npu_inst_pe_1_6_7_int_q_reg_h_4__1_,
         npu_inst_pe_1_6_7_int_q_reg_h_3__0_,
         npu_inst_pe_1_6_7_int_q_reg_h_3__1_,
         npu_inst_pe_1_6_7_int_q_reg_h_2__0_,
         npu_inst_pe_1_6_7_int_q_reg_h_2__1_,
         npu_inst_pe_1_6_7_int_q_reg_h_1__0_,
         npu_inst_pe_1_6_7_int_q_reg_h_1__1_,
         npu_inst_pe_1_6_7_int_q_reg_h_0__0_,
         npu_inst_pe_1_6_7_int_q_reg_h_0__1_, npu_inst_pe_1_7_0_n119,
         npu_inst_pe_1_7_0_n118, npu_inst_pe_1_7_0_n117,
         npu_inst_pe_1_7_0_n116, npu_inst_pe_1_7_0_n115,
         npu_inst_pe_1_7_0_n114, npu_inst_pe_1_7_0_n113,
         npu_inst_pe_1_7_0_n112, npu_inst_pe_1_7_0_n111,
         npu_inst_pe_1_7_0_n110, npu_inst_pe_1_7_0_n109,
         npu_inst_pe_1_7_0_n108, npu_inst_pe_1_7_0_n107,
         npu_inst_pe_1_7_0_n106, npu_inst_pe_1_7_0_n105,
         npu_inst_pe_1_7_0_n104, npu_inst_pe_1_7_0_n103,
         npu_inst_pe_1_7_0_n102, npu_inst_pe_1_7_0_n101,
         npu_inst_pe_1_7_0_n100, npu_inst_pe_1_7_0_n99, npu_inst_pe_1_7_0_n98,
         npu_inst_pe_1_7_0_n36, npu_inst_pe_1_7_0_n35, npu_inst_pe_1_7_0_n34,
         npu_inst_pe_1_7_0_n33, npu_inst_pe_1_7_0_n32, npu_inst_pe_1_7_0_n31,
         npu_inst_pe_1_7_0_n30, npu_inst_pe_1_7_0_n29, npu_inst_pe_1_7_0_n28,
         npu_inst_pe_1_7_0_n25, npu_inst_pe_1_7_0_n24, npu_inst_pe_1_7_0_n23,
         npu_inst_pe_1_7_0_n22, npu_inst_pe_1_7_0_n21, npu_inst_pe_1_7_0_n20,
         npu_inst_pe_1_7_0_n19, npu_inst_pe_1_7_0_n18, npu_inst_pe_1_7_0_n17,
         npu_inst_pe_1_7_0_n16, npu_inst_pe_1_7_0_n15, npu_inst_pe_1_7_0_n14,
         npu_inst_pe_1_7_0_n13, npu_inst_pe_1_7_0_n12, npu_inst_pe_1_7_0_n11,
         npu_inst_pe_1_7_0_n10, npu_inst_pe_1_7_0_n9, npu_inst_pe_1_7_0_n8,
         npu_inst_pe_1_7_0_n7, npu_inst_pe_1_7_0_n6, npu_inst_pe_1_7_0_n5,
         npu_inst_pe_1_7_0_n4, npu_inst_pe_1_7_0_n3, npu_inst_pe_1_7_0_n2,
         npu_inst_pe_1_7_0_n1, npu_inst_pe_1_7_0_sub_67_carry_7_,
         npu_inst_pe_1_7_0_sub_67_carry_6_, npu_inst_pe_1_7_0_sub_67_carry_5_,
         npu_inst_pe_1_7_0_sub_67_carry_4_, npu_inst_pe_1_7_0_sub_67_carry_3_,
         npu_inst_pe_1_7_0_sub_67_carry_2_, npu_inst_pe_1_7_0_sub_67_carry_1_,
         npu_inst_pe_1_7_0_add_69_carry_7_, npu_inst_pe_1_7_0_add_69_carry_6_,
         npu_inst_pe_1_7_0_add_69_carry_5_, npu_inst_pe_1_7_0_add_69_carry_4_,
         npu_inst_pe_1_7_0_add_69_carry_3_, npu_inst_pe_1_7_0_add_69_carry_2_,
         npu_inst_pe_1_7_0_add_69_carry_1_, npu_inst_pe_1_7_0_n97,
         npu_inst_pe_1_7_0_n96, npu_inst_pe_1_7_0_n95, npu_inst_pe_1_7_0_n94,
         npu_inst_pe_1_7_0_n93, npu_inst_pe_1_7_0_n92, npu_inst_pe_1_7_0_n91,
         npu_inst_pe_1_7_0_n90, npu_inst_pe_1_7_0_n89, npu_inst_pe_1_7_0_n88,
         npu_inst_pe_1_7_0_n87, npu_inst_pe_1_7_0_n86, npu_inst_pe_1_7_0_n85,
         npu_inst_pe_1_7_0_n84, npu_inst_pe_1_7_0_n83, npu_inst_pe_1_7_0_n82,
         npu_inst_pe_1_7_0_n81, npu_inst_pe_1_7_0_n80, npu_inst_pe_1_7_0_n79,
         npu_inst_pe_1_7_0_n78, npu_inst_pe_1_7_0_n77, npu_inst_pe_1_7_0_n76,
         npu_inst_pe_1_7_0_n75, npu_inst_pe_1_7_0_n74, npu_inst_pe_1_7_0_n73,
         npu_inst_pe_1_7_0_n72, npu_inst_pe_1_7_0_n71, npu_inst_pe_1_7_0_n70,
         npu_inst_pe_1_7_0_n69, npu_inst_pe_1_7_0_n68, npu_inst_pe_1_7_0_n67,
         npu_inst_pe_1_7_0_n66, npu_inst_pe_1_7_0_n65, npu_inst_pe_1_7_0_n64,
         npu_inst_pe_1_7_0_n63, npu_inst_pe_1_7_0_n62, npu_inst_pe_1_7_0_n61,
         npu_inst_pe_1_7_0_n60, npu_inst_pe_1_7_0_n59, npu_inst_pe_1_7_0_n58,
         npu_inst_pe_1_7_0_n57, npu_inst_pe_1_7_0_n56, npu_inst_pe_1_7_0_n55,
         npu_inst_pe_1_7_0_n54, npu_inst_pe_1_7_0_n53, npu_inst_pe_1_7_0_n52,
         npu_inst_pe_1_7_0_n51, npu_inst_pe_1_7_0_n50, npu_inst_pe_1_7_0_n49,
         npu_inst_pe_1_7_0_n48, npu_inst_pe_1_7_0_n47, npu_inst_pe_1_7_0_n46,
         npu_inst_pe_1_7_0_n45, npu_inst_pe_1_7_0_n44, npu_inst_pe_1_7_0_n43,
         npu_inst_pe_1_7_0_n42, npu_inst_pe_1_7_0_n41, npu_inst_pe_1_7_0_n40,
         npu_inst_pe_1_7_0_n39, npu_inst_pe_1_7_0_n38, npu_inst_pe_1_7_0_n37,
         npu_inst_pe_1_7_0_n27, npu_inst_pe_1_7_0_n26,
         npu_inst_pe_1_7_0_net3280, npu_inst_pe_1_7_0_net3274,
         npu_inst_pe_1_7_0_N94, npu_inst_pe_1_7_0_N93, npu_inst_pe_1_7_0_N84,
         npu_inst_pe_1_7_0_N80, npu_inst_pe_1_7_0_N79, npu_inst_pe_1_7_0_N78,
         npu_inst_pe_1_7_0_N77, npu_inst_pe_1_7_0_N76, npu_inst_pe_1_7_0_N75,
         npu_inst_pe_1_7_0_N74, npu_inst_pe_1_7_0_N73, npu_inst_pe_1_7_0_N72,
         npu_inst_pe_1_7_0_N71, npu_inst_pe_1_7_0_N70, npu_inst_pe_1_7_0_N69,
         npu_inst_pe_1_7_0_N68, npu_inst_pe_1_7_0_N67, npu_inst_pe_1_7_0_N66,
         npu_inst_pe_1_7_0_N65, npu_inst_pe_1_7_0_int_q_acc_0_,
         npu_inst_pe_1_7_0_int_q_acc_1_, npu_inst_pe_1_7_0_int_q_acc_2_,
         npu_inst_pe_1_7_0_int_q_acc_3_, npu_inst_pe_1_7_0_int_q_acc_4_,
         npu_inst_pe_1_7_0_int_q_acc_5_, npu_inst_pe_1_7_0_int_q_acc_6_,
         npu_inst_pe_1_7_0_int_q_acc_7_, npu_inst_pe_1_7_0_int_data_0_,
         npu_inst_pe_1_7_0_int_data_1_, npu_inst_pe_1_7_0_int_q_weight_0_,
         npu_inst_pe_1_7_0_int_q_weight_1_,
         npu_inst_pe_1_7_0_int_q_reg_v_5__0_,
         npu_inst_pe_1_7_0_int_q_reg_v_5__1_,
         npu_inst_pe_1_7_0_int_q_reg_v_4__0_,
         npu_inst_pe_1_7_0_int_q_reg_v_4__1_,
         npu_inst_pe_1_7_0_int_q_reg_v_3__0_,
         npu_inst_pe_1_7_0_int_q_reg_v_3__1_,
         npu_inst_pe_1_7_0_int_q_reg_v_2__0_,
         npu_inst_pe_1_7_0_int_q_reg_v_2__1_,
         npu_inst_pe_1_7_0_int_q_reg_v_1__0_,
         npu_inst_pe_1_7_0_int_q_reg_v_1__1_,
         npu_inst_pe_1_7_0_int_q_reg_v_0__0_,
         npu_inst_pe_1_7_0_int_q_reg_v_0__1_,
         npu_inst_pe_1_7_0_int_q_reg_h_5__0_,
         npu_inst_pe_1_7_0_int_q_reg_h_5__1_,
         npu_inst_pe_1_7_0_int_q_reg_h_4__0_,
         npu_inst_pe_1_7_0_int_q_reg_h_4__1_,
         npu_inst_pe_1_7_0_int_q_reg_h_3__0_,
         npu_inst_pe_1_7_0_int_q_reg_h_3__1_,
         npu_inst_pe_1_7_0_int_q_reg_h_2__0_,
         npu_inst_pe_1_7_0_int_q_reg_h_2__1_,
         npu_inst_pe_1_7_0_int_q_reg_h_1__0_,
         npu_inst_pe_1_7_0_int_q_reg_h_1__1_,
         npu_inst_pe_1_7_0_int_q_reg_h_0__0_,
         npu_inst_pe_1_7_0_int_q_reg_h_0__1_, npu_inst_pe_1_7_0_o_data_h_0_,
         npu_inst_pe_1_7_0_o_data_h_1_, npu_inst_pe_1_7_1_n119,
         npu_inst_pe_1_7_1_n118, npu_inst_pe_1_7_1_n117,
         npu_inst_pe_1_7_1_n116, npu_inst_pe_1_7_1_n115,
         npu_inst_pe_1_7_1_n114, npu_inst_pe_1_7_1_n113,
         npu_inst_pe_1_7_1_n112, npu_inst_pe_1_7_1_n111,
         npu_inst_pe_1_7_1_n110, npu_inst_pe_1_7_1_n109,
         npu_inst_pe_1_7_1_n108, npu_inst_pe_1_7_1_n107,
         npu_inst_pe_1_7_1_n106, npu_inst_pe_1_7_1_n105,
         npu_inst_pe_1_7_1_n104, npu_inst_pe_1_7_1_n103,
         npu_inst_pe_1_7_1_n102, npu_inst_pe_1_7_1_n101,
         npu_inst_pe_1_7_1_n100, npu_inst_pe_1_7_1_n99, npu_inst_pe_1_7_1_n98,
         npu_inst_pe_1_7_1_n36, npu_inst_pe_1_7_1_n35, npu_inst_pe_1_7_1_n34,
         npu_inst_pe_1_7_1_n33, npu_inst_pe_1_7_1_n32, npu_inst_pe_1_7_1_n31,
         npu_inst_pe_1_7_1_n30, npu_inst_pe_1_7_1_n29, npu_inst_pe_1_7_1_n28,
         npu_inst_pe_1_7_1_n25, npu_inst_pe_1_7_1_n24, npu_inst_pe_1_7_1_n23,
         npu_inst_pe_1_7_1_n22, npu_inst_pe_1_7_1_n21, npu_inst_pe_1_7_1_n20,
         npu_inst_pe_1_7_1_n19, npu_inst_pe_1_7_1_n18, npu_inst_pe_1_7_1_n17,
         npu_inst_pe_1_7_1_n16, npu_inst_pe_1_7_1_n15, npu_inst_pe_1_7_1_n14,
         npu_inst_pe_1_7_1_n13, npu_inst_pe_1_7_1_n12, npu_inst_pe_1_7_1_n11,
         npu_inst_pe_1_7_1_n10, npu_inst_pe_1_7_1_n9, npu_inst_pe_1_7_1_n8,
         npu_inst_pe_1_7_1_n7, npu_inst_pe_1_7_1_n6, npu_inst_pe_1_7_1_n5,
         npu_inst_pe_1_7_1_n4, npu_inst_pe_1_7_1_n3, npu_inst_pe_1_7_1_n2,
         npu_inst_pe_1_7_1_n1, npu_inst_pe_1_7_1_sub_67_carry_7_,
         npu_inst_pe_1_7_1_sub_67_carry_6_, npu_inst_pe_1_7_1_sub_67_carry_5_,
         npu_inst_pe_1_7_1_sub_67_carry_4_, npu_inst_pe_1_7_1_sub_67_carry_3_,
         npu_inst_pe_1_7_1_sub_67_carry_2_, npu_inst_pe_1_7_1_sub_67_carry_1_,
         npu_inst_pe_1_7_1_add_69_carry_7_, npu_inst_pe_1_7_1_add_69_carry_6_,
         npu_inst_pe_1_7_1_add_69_carry_5_, npu_inst_pe_1_7_1_add_69_carry_4_,
         npu_inst_pe_1_7_1_add_69_carry_3_, npu_inst_pe_1_7_1_add_69_carry_2_,
         npu_inst_pe_1_7_1_add_69_carry_1_, npu_inst_pe_1_7_1_n97,
         npu_inst_pe_1_7_1_n96, npu_inst_pe_1_7_1_n95, npu_inst_pe_1_7_1_n94,
         npu_inst_pe_1_7_1_n93, npu_inst_pe_1_7_1_n92, npu_inst_pe_1_7_1_n91,
         npu_inst_pe_1_7_1_n90, npu_inst_pe_1_7_1_n89, npu_inst_pe_1_7_1_n88,
         npu_inst_pe_1_7_1_n87, npu_inst_pe_1_7_1_n86, npu_inst_pe_1_7_1_n85,
         npu_inst_pe_1_7_1_n84, npu_inst_pe_1_7_1_n83, npu_inst_pe_1_7_1_n82,
         npu_inst_pe_1_7_1_n81, npu_inst_pe_1_7_1_n80, npu_inst_pe_1_7_1_n79,
         npu_inst_pe_1_7_1_n78, npu_inst_pe_1_7_1_n77, npu_inst_pe_1_7_1_n76,
         npu_inst_pe_1_7_1_n75, npu_inst_pe_1_7_1_n74, npu_inst_pe_1_7_1_n73,
         npu_inst_pe_1_7_1_n72, npu_inst_pe_1_7_1_n71, npu_inst_pe_1_7_1_n70,
         npu_inst_pe_1_7_1_n69, npu_inst_pe_1_7_1_n68, npu_inst_pe_1_7_1_n67,
         npu_inst_pe_1_7_1_n66, npu_inst_pe_1_7_1_n65, npu_inst_pe_1_7_1_n64,
         npu_inst_pe_1_7_1_n63, npu_inst_pe_1_7_1_n62, npu_inst_pe_1_7_1_n61,
         npu_inst_pe_1_7_1_n60, npu_inst_pe_1_7_1_n59, npu_inst_pe_1_7_1_n58,
         npu_inst_pe_1_7_1_n57, npu_inst_pe_1_7_1_n56, npu_inst_pe_1_7_1_n55,
         npu_inst_pe_1_7_1_n54, npu_inst_pe_1_7_1_n53, npu_inst_pe_1_7_1_n52,
         npu_inst_pe_1_7_1_n51, npu_inst_pe_1_7_1_n50, npu_inst_pe_1_7_1_n49,
         npu_inst_pe_1_7_1_n48, npu_inst_pe_1_7_1_n47, npu_inst_pe_1_7_1_n46,
         npu_inst_pe_1_7_1_n45, npu_inst_pe_1_7_1_n44, npu_inst_pe_1_7_1_n43,
         npu_inst_pe_1_7_1_n42, npu_inst_pe_1_7_1_n41, npu_inst_pe_1_7_1_n40,
         npu_inst_pe_1_7_1_n39, npu_inst_pe_1_7_1_n38, npu_inst_pe_1_7_1_n37,
         npu_inst_pe_1_7_1_n27, npu_inst_pe_1_7_1_n26,
         npu_inst_pe_1_7_1_net3257, npu_inst_pe_1_7_1_net3251,
         npu_inst_pe_1_7_1_N94, npu_inst_pe_1_7_1_N93, npu_inst_pe_1_7_1_N84,
         npu_inst_pe_1_7_1_N80, npu_inst_pe_1_7_1_N79, npu_inst_pe_1_7_1_N78,
         npu_inst_pe_1_7_1_N77, npu_inst_pe_1_7_1_N76, npu_inst_pe_1_7_1_N75,
         npu_inst_pe_1_7_1_N74, npu_inst_pe_1_7_1_N73, npu_inst_pe_1_7_1_N72,
         npu_inst_pe_1_7_1_N71, npu_inst_pe_1_7_1_N70, npu_inst_pe_1_7_1_N69,
         npu_inst_pe_1_7_1_N68, npu_inst_pe_1_7_1_N67, npu_inst_pe_1_7_1_N66,
         npu_inst_pe_1_7_1_N65, npu_inst_pe_1_7_1_int_q_acc_0_,
         npu_inst_pe_1_7_1_int_q_acc_1_, npu_inst_pe_1_7_1_int_q_acc_2_,
         npu_inst_pe_1_7_1_int_q_acc_3_, npu_inst_pe_1_7_1_int_q_acc_4_,
         npu_inst_pe_1_7_1_int_q_acc_5_, npu_inst_pe_1_7_1_int_q_acc_6_,
         npu_inst_pe_1_7_1_int_q_acc_7_, npu_inst_pe_1_7_1_int_data_0_,
         npu_inst_pe_1_7_1_int_data_1_, npu_inst_pe_1_7_1_int_q_weight_0_,
         npu_inst_pe_1_7_1_int_q_weight_1_,
         npu_inst_pe_1_7_1_int_q_reg_v_5__0_,
         npu_inst_pe_1_7_1_int_q_reg_v_5__1_,
         npu_inst_pe_1_7_1_int_q_reg_v_4__0_,
         npu_inst_pe_1_7_1_int_q_reg_v_4__1_,
         npu_inst_pe_1_7_1_int_q_reg_v_3__0_,
         npu_inst_pe_1_7_1_int_q_reg_v_3__1_,
         npu_inst_pe_1_7_1_int_q_reg_v_2__0_,
         npu_inst_pe_1_7_1_int_q_reg_v_2__1_,
         npu_inst_pe_1_7_1_int_q_reg_v_1__0_,
         npu_inst_pe_1_7_1_int_q_reg_v_1__1_,
         npu_inst_pe_1_7_1_int_q_reg_v_0__0_,
         npu_inst_pe_1_7_1_int_q_reg_v_0__1_,
         npu_inst_pe_1_7_1_int_q_reg_h_5__0_,
         npu_inst_pe_1_7_1_int_q_reg_h_5__1_,
         npu_inst_pe_1_7_1_int_q_reg_h_4__0_,
         npu_inst_pe_1_7_1_int_q_reg_h_4__1_,
         npu_inst_pe_1_7_1_int_q_reg_h_3__0_,
         npu_inst_pe_1_7_1_int_q_reg_h_3__1_,
         npu_inst_pe_1_7_1_int_q_reg_h_2__0_,
         npu_inst_pe_1_7_1_int_q_reg_h_2__1_,
         npu_inst_pe_1_7_1_int_q_reg_h_1__0_,
         npu_inst_pe_1_7_1_int_q_reg_h_1__1_,
         npu_inst_pe_1_7_1_int_q_reg_h_0__0_,
         npu_inst_pe_1_7_1_int_q_reg_h_0__1_, npu_inst_pe_1_7_2_n119,
         npu_inst_pe_1_7_2_n118, npu_inst_pe_1_7_2_n117,
         npu_inst_pe_1_7_2_n116, npu_inst_pe_1_7_2_n115,
         npu_inst_pe_1_7_2_n114, npu_inst_pe_1_7_2_n113,
         npu_inst_pe_1_7_2_n112, npu_inst_pe_1_7_2_n111,
         npu_inst_pe_1_7_2_n110, npu_inst_pe_1_7_2_n109,
         npu_inst_pe_1_7_2_n108, npu_inst_pe_1_7_2_n107,
         npu_inst_pe_1_7_2_n106, npu_inst_pe_1_7_2_n105,
         npu_inst_pe_1_7_2_n104, npu_inst_pe_1_7_2_n103,
         npu_inst_pe_1_7_2_n102, npu_inst_pe_1_7_2_n101,
         npu_inst_pe_1_7_2_n100, npu_inst_pe_1_7_2_n99, npu_inst_pe_1_7_2_n98,
         npu_inst_pe_1_7_2_n36, npu_inst_pe_1_7_2_n35, npu_inst_pe_1_7_2_n34,
         npu_inst_pe_1_7_2_n33, npu_inst_pe_1_7_2_n32, npu_inst_pe_1_7_2_n31,
         npu_inst_pe_1_7_2_n30, npu_inst_pe_1_7_2_n29, npu_inst_pe_1_7_2_n28,
         npu_inst_pe_1_7_2_n25, npu_inst_pe_1_7_2_n24, npu_inst_pe_1_7_2_n23,
         npu_inst_pe_1_7_2_n22, npu_inst_pe_1_7_2_n21, npu_inst_pe_1_7_2_n20,
         npu_inst_pe_1_7_2_n19, npu_inst_pe_1_7_2_n18, npu_inst_pe_1_7_2_n17,
         npu_inst_pe_1_7_2_n16, npu_inst_pe_1_7_2_n15, npu_inst_pe_1_7_2_n14,
         npu_inst_pe_1_7_2_n13, npu_inst_pe_1_7_2_n12, npu_inst_pe_1_7_2_n11,
         npu_inst_pe_1_7_2_n10, npu_inst_pe_1_7_2_n9, npu_inst_pe_1_7_2_n8,
         npu_inst_pe_1_7_2_n7, npu_inst_pe_1_7_2_n6, npu_inst_pe_1_7_2_n5,
         npu_inst_pe_1_7_2_n4, npu_inst_pe_1_7_2_n3, npu_inst_pe_1_7_2_n2,
         npu_inst_pe_1_7_2_n1, npu_inst_pe_1_7_2_sub_67_carry_7_,
         npu_inst_pe_1_7_2_sub_67_carry_6_, npu_inst_pe_1_7_2_sub_67_carry_5_,
         npu_inst_pe_1_7_2_sub_67_carry_4_, npu_inst_pe_1_7_2_sub_67_carry_3_,
         npu_inst_pe_1_7_2_sub_67_carry_2_, npu_inst_pe_1_7_2_sub_67_carry_1_,
         npu_inst_pe_1_7_2_add_69_carry_7_, npu_inst_pe_1_7_2_add_69_carry_6_,
         npu_inst_pe_1_7_2_add_69_carry_5_, npu_inst_pe_1_7_2_add_69_carry_4_,
         npu_inst_pe_1_7_2_add_69_carry_3_, npu_inst_pe_1_7_2_add_69_carry_2_,
         npu_inst_pe_1_7_2_add_69_carry_1_, npu_inst_pe_1_7_2_n97,
         npu_inst_pe_1_7_2_n96, npu_inst_pe_1_7_2_n95, npu_inst_pe_1_7_2_n94,
         npu_inst_pe_1_7_2_n93, npu_inst_pe_1_7_2_n92, npu_inst_pe_1_7_2_n91,
         npu_inst_pe_1_7_2_n90, npu_inst_pe_1_7_2_n89, npu_inst_pe_1_7_2_n88,
         npu_inst_pe_1_7_2_n87, npu_inst_pe_1_7_2_n86, npu_inst_pe_1_7_2_n85,
         npu_inst_pe_1_7_2_n84, npu_inst_pe_1_7_2_n83, npu_inst_pe_1_7_2_n82,
         npu_inst_pe_1_7_2_n81, npu_inst_pe_1_7_2_n80, npu_inst_pe_1_7_2_n79,
         npu_inst_pe_1_7_2_n78, npu_inst_pe_1_7_2_n77, npu_inst_pe_1_7_2_n76,
         npu_inst_pe_1_7_2_n75, npu_inst_pe_1_7_2_n74, npu_inst_pe_1_7_2_n73,
         npu_inst_pe_1_7_2_n72, npu_inst_pe_1_7_2_n71, npu_inst_pe_1_7_2_n70,
         npu_inst_pe_1_7_2_n69, npu_inst_pe_1_7_2_n68, npu_inst_pe_1_7_2_n67,
         npu_inst_pe_1_7_2_n66, npu_inst_pe_1_7_2_n65, npu_inst_pe_1_7_2_n64,
         npu_inst_pe_1_7_2_n63, npu_inst_pe_1_7_2_n62, npu_inst_pe_1_7_2_n61,
         npu_inst_pe_1_7_2_n60, npu_inst_pe_1_7_2_n59, npu_inst_pe_1_7_2_n58,
         npu_inst_pe_1_7_2_n57, npu_inst_pe_1_7_2_n56, npu_inst_pe_1_7_2_n55,
         npu_inst_pe_1_7_2_n54, npu_inst_pe_1_7_2_n53, npu_inst_pe_1_7_2_n52,
         npu_inst_pe_1_7_2_n51, npu_inst_pe_1_7_2_n50, npu_inst_pe_1_7_2_n49,
         npu_inst_pe_1_7_2_n48, npu_inst_pe_1_7_2_n47, npu_inst_pe_1_7_2_n46,
         npu_inst_pe_1_7_2_n45, npu_inst_pe_1_7_2_n44, npu_inst_pe_1_7_2_n43,
         npu_inst_pe_1_7_2_n42, npu_inst_pe_1_7_2_n41, npu_inst_pe_1_7_2_n40,
         npu_inst_pe_1_7_2_n39, npu_inst_pe_1_7_2_n38, npu_inst_pe_1_7_2_n37,
         npu_inst_pe_1_7_2_n27, npu_inst_pe_1_7_2_n26,
         npu_inst_pe_1_7_2_net3234, npu_inst_pe_1_7_2_net3228,
         npu_inst_pe_1_7_2_N94, npu_inst_pe_1_7_2_N93, npu_inst_pe_1_7_2_N84,
         npu_inst_pe_1_7_2_N80, npu_inst_pe_1_7_2_N79, npu_inst_pe_1_7_2_N78,
         npu_inst_pe_1_7_2_N77, npu_inst_pe_1_7_2_N76, npu_inst_pe_1_7_2_N75,
         npu_inst_pe_1_7_2_N74, npu_inst_pe_1_7_2_N73, npu_inst_pe_1_7_2_N72,
         npu_inst_pe_1_7_2_N71, npu_inst_pe_1_7_2_N70, npu_inst_pe_1_7_2_N69,
         npu_inst_pe_1_7_2_N68, npu_inst_pe_1_7_2_N67, npu_inst_pe_1_7_2_N66,
         npu_inst_pe_1_7_2_N65, npu_inst_pe_1_7_2_int_q_acc_0_,
         npu_inst_pe_1_7_2_int_q_acc_1_, npu_inst_pe_1_7_2_int_q_acc_2_,
         npu_inst_pe_1_7_2_int_q_acc_3_, npu_inst_pe_1_7_2_int_q_acc_4_,
         npu_inst_pe_1_7_2_int_q_acc_5_, npu_inst_pe_1_7_2_int_q_acc_6_,
         npu_inst_pe_1_7_2_int_q_acc_7_, npu_inst_pe_1_7_2_int_data_0_,
         npu_inst_pe_1_7_2_int_data_1_, npu_inst_pe_1_7_2_int_q_weight_0_,
         npu_inst_pe_1_7_2_int_q_weight_1_,
         npu_inst_pe_1_7_2_int_q_reg_v_5__0_,
         npu_inst_pe_1_7_2_int_q_reg_v_5__1_,
         npu_inst_pe_1_7_2_int_q_reg_v_4__0_,
         npu_inst_pe_1_7_2_int_q_reg_v_4__1_,
         npu_inst_pe_1_7_2_int_q_reg_v_3__0_,
         npu_inst_pe_1_7_2_int_q_reg_v_3__1_,
         npu_inst_pe_1_7_2_int_q_reg_v_2__0_,
         npu_inst_pe_1_7_2_int_q_reg_v_2__1_,
         npu_inst_pe_1_7_2_int_q_reg_v_1__0_,
         npu_inst_pe_1_7_2_int_q_reg_v_1__1_,
         npu_inst_pe_1_7_2_int_q_reg_v_0__0_,
         npu_inst_pe_1_7_2_int_q_reg_v_0__1_,
         npu_inst_pe_1_7_2_int_q_reg_h_5__0_,
         npu_inst_pe_1_7_2_int_q_reg_h_5__1_,
         npu_inst_pe_1_7_2_int_q_reg_h_4__0_,
         npu_inst_pe_1_7_2_int_q_reg_h_4__1_,
         npu_inst_pe_1_7_2_int_q_reg_h_3__0_,
         npu_inst_pe_1_7_2_int_q_reg_h_3__1_,
         npu_inst_pe_1_7_2_int_q_reg_h_2__0_,
         npu_inst_pe_1_7_2_int_q_reg_h_2__1_,
         npu_inst_pe_1_7_2_int_q_reg_h_1__0_,
         npu_inst_pe_1_7_2_int_q_reg_h_1__1_,
         npu_inst_pe_1_7_2_int_q_reg_h_0__0_,
         npu_inst_pe_1_7_2_int_q_reg_h_0__1_, npu_inst_pe_1_7_3_n119,
         npu_inst_pe_1_7_3_n118, npu_inst_pe_1_7_3_n117,
         npu_inst_pe_1_7_3_n116, npu_inst_pe_1_7_3_n115,
         npu_inst_pe_1_7_3_n114, npu_inst_pe_1_7_3_n113,
         npu_inst_pe_1_7_3_n112, npu_inst_pe_1_7_3_n111,
         npu_inst_pe_1_7_3_n110, npu_inst_pe_1_7_3_n109,
         npu_inst_pe_1_7_3_n108, npu_inst_pe_1_7_3_n107,
         npu_inst_pe_1_7_3_n106, npu_inst_pe_1_7_3_n105,
         npu_inst_pe_1_7_3_n104, npu_inst_pe_1_7_3_n103,
         npu_inst_pe_1_7_3_n102, npu_inst_pe_1_7_3_n101,
         npu_inst_pe_1_7_3_n100, npu_inst_pe_1_7_3_n99, npu_inst_pe_1_7_3_n98,
         npu_inst_pe_1_7_3_n36, npu_inst_pe_1_7_3_n35, npu_inst_pe_1_7_3_n34,
         npu_inst_pe_1_7_3_n33, npu_inst_pe_1_7_3_n32, npu_inst_pe_1_7_3_n31,
         npu_inst_pe_1_7_3_n30, npu_inst_pe_1_7_3_n29, npu_inst_pe_1_7_3_n28,
         npu_inst_pe_1_7_3_n25, npu_inst_pe_1_7_3_n24, npu_inst_pe_1_7_3_n23,
         npu_inst_pe_1_7_3_n22, npu_inst_pe_1_7_3_n21, npu_inst_pe_1_7_3_n20,
         npu_inst_pe_1_7_3_n19, npu_inst_pe_1_7_3_n18, npu_inst_pe_1_7_3_n17,
         npu_inst_pe_1_7_3_n16, npu_inst_pe_1_7_3_n15, npu_inst_pe_1_7_3_n14,
         npu_inst_pe_1_7_3_n13, npu_inst_pe_1_7_3_n12, npu_inst_pe_1_7_3_n11,
         npu_inst_pe_1_7_3_n10, npu_inst_pe_1_7_3_n9, npu_inst_pe_1_7_3_n8,
         npu_inst_pe_1_7_3_n7, npu_inst_pe_1_7_3_n6, npu_inst_pe_1_7_3_n5,
         npu_inst_pe_1_7_3_n4, npu_inst_pe_1_7_3_n3, npu_inst_pe_1_7_3_n2,
         npu_inst_pe_1_7_3_n1, npu_inst_pe_1_7_3_sub_67_carry_7_,
         npu_inst_pe_1_7_3_sub_67_carry_6_, npu_inst_pe_1_7_3_sub_67_carry_5_,
         npu_inst_pe_1_7_3_sub_67_carry_4_, npu_inst_pe_1_7_3_sub_67_carry_3_,
         npu_inst_pe_1_7_3_sub_67_carry_2_, npu_inst_pe_1_7_3_sub_67_carry_1_,
         npu_inst_pe_1_7_3_add_69_carry_7_, npu_inst_pe_1_7_3_add_69_carry_6_,
         npu_inst_pe_1_7_3_add_69_carry_5_, npu_inst_pe_1_7_3_add_69_carry_4_,
         npu_inst_pe_1_7_3_add_69_carry_3_, npu_inst_pe_1_7_3_add_69_carry_2_,
         npu_inst_pe_1_7_3_add_69_carry_1_, npu_inst_pe_1_7_3_n97,
         npu_inst_pe_1_7_3_n96, npu_inst_pe_1_7_3_n95, npu_inst_pe_1_7_3_n94,
         npu_inst_pe_1_7_3_n93, npu_inst_pe_1_7_3_n92, npu_inst_pe_1_7_3_n91,
         npu_inst_pe_1_7_3_n90, npu_inst_pe_1_7_3_n89, npu_inst_pe_1_7_3_n88,
         npu_inst_pe_1_7_3_n87, npu_inst_pe_1_7_3_n86, npu_inst_pe_1_7_3_n85,
         npu_inst_pe_1_7_3_n84, npu_inst_pe_1_7_3_n83, npu_inst_pe_1_7_3_n82,
         npu_inst_pe_1_7_3_n81, npu_inst_pe_1_7_3_n80, npu_inst_pe_1_7_3_n79,
         npu_inst_pe_1_7_3_n78, npu_inst_pe_1_7_3_n77, npu_inst_pe_1_7_3_n76,
         npu_inst_pe_1_7_3_n75, npu_inst_pe_1_7_3_n74, npu_inst_pe_1_7_3_n73,
         npu_inst_pe_1_7_3_n72, npu_inst_pe_1_7_3_n71, npu_inst_pe_1_7_3_n70,
         npu_inst_pe_1_7_3_n69, npu_inst_pe_1_7_3_n68, npu_inst_pe_1_7_3_n67,
         npu_inst_pe_1_7_3_n66, npu_inst_pe_1_7_3_n65, npu_inst_pe_1_7_3_n64,
         npu_inst_pe_1_7_3_n63, npu_inst_pe_1_7_3_n62, npu_inst_pe_1_7_3_n61,
         npu_inst_pe_1_7_3_n60, npu_inst_pe_1_7_3_n59, npu_inst_pe_1_7_3_n58,
         npu_inst_pe_1_7_3_n57, npu_inst_pe_1_7_3_n56, npu_inst_pe_1_7_3_n55,
         npu_inst_pe_1_7_3_n54, npu_inst_pe_1_7_3_n53, npu_inst_pe_1_7_3_n52,
         npu_inst_pe_1_7_3_n51, npu_inst_pe_1_7_3_n50, npu_inst_pe_1_7_3_n49,
         npu_inst_pe_1_7_3_n48, npu_inst_pe_1_7_3_n47, npu_inst_pe_1_7_3_n46,
         npu_inst_pe_1_7_3_n45, npu_inst_pe_1_7_3_n44, npu_inst_pe_1_7_3_n43,
         npu_inst_pe_1_7_3_n42, npu_inst_pe_1_7_3_n41, npu_inst_pe_1_7_3_n40,
         npu_inst_pe_1_7_3_n39, npu_inst_pe_1_7_3_n38, npu_inst_pe_1_7_3_n37,
         npu_inst_pe_1_7_3_n27, npu_inst_pe_1_7_3_n26,
         npu_inst_pe_1_7_3_net3211, npu_inst_pe_1_7_3_net3205,
         npu_inst_pe_1_7_3_N94, npu_inst_pe_1_7_3_N93, npu_inst_pe_1_7_3_N84,
         npu_inst_pe_1_7_3_N80, npu_inst_pe_1_7_3_N79, npu_inst_pe_1_7_3_N78,
         npu_inst_pe_1_7_3_N77, npu_inst_pe_1_7_3_N76, npu_inst_pe_1_7_3_N75,
         npu_inst_pe_1_7_3_N74, npu_inst_pe_1_7_3_N73, npu_inst_pe_1_7_3_N72,
         npu_inst_pe_1_7_3_N71, npu_inst_pe_1_7_3_N70, npu_inst_pe_1_7_3_N69,
         npu_inst_pe_1_7_3_N68, npu_inst_pe_1_7_3_N67, npu_inst_pe_1_7_3_N66,
         npu_inst_pe_1_7_3_N65, npu_inst_pe_1_7_3_int_q_acc_0_,
         npu_inst_pe_1_7_3_int_q_acc_1_, npu_inst_pe_1_7_3_int_q_acc_2_,
         npu_inst_pe_1_7_3_int_q_acc_3_, npu_inst_pe_1_7_3_int_q_acc_4_,
         npu_inst_pe_1_7_3_int_q_acc_5_, npu_inst_pe_1_7_3_int_q_acc_6_,
         npu_inst_pe_1_7_3_int_q_acc_7_, npu_inst_pe_1_7_3_int_data_0_,
         npu_inst_pe_1_7_3_int_data_1_, npu_inst_pe_1_7_3_int_q_weight_0_,
         npu_inst_pe_1_7_3_int_q_weight_1_,
         npu_inst_pe_1_7_3_int_q_reg_v_5__0_,
         npu_inst_pe_1_7_3_int_q_reg_v_5__1_,
         npu_inst_pe_1_7_3_int_q_reg_v_4__0_,
         npu_inst_pe_1_7_3_int_q_reg_v_4__1_,
         npu_inst_pe_1_7_3_int_q_reg_v_3__0_,
         npu_inst_pe_1_7_3_int_q_reg_v_3__1_,
         npu_inst_pe_1_7_3_int_q_reg_v_2__0_,
         npu_inst_pe_1_7_3_int_q_reg_v_2__1_,
         npu_inst_pe_1_7_3_int_q_reg_v_1__0_,
         npu_inst_pe_1_7_3_int_q_reg_v_1__1_,
         npu_inst_pe_1_7_3_int_q_reg_v_0__0_,
         npu_inst_pe_1_7_3_int_q_reg_v_0__1_,
         npu_inst_pe_1_7_3_int_q_reg_h_5__0_,
         npu_inst_pe_1_7_3_int_q_reg_h_5__1_,
         npu_inst_pe_1_7_3_int_q_reg_h_4__0_,
         npu_inst_pe_1_7_3_int_q_reg_h_4__1_,
         npu_inst_pe_1_7_3_int_q_reg_h_3__0_,
         npu_inst_pe_1_7_3_int_q_reg_h_3__1_,
         npu_inst_pe_1_7_3_int_q_reg_h_2__0_,
         npu_inst_pe_1_7_3_int_q_reg_h_2__1_,
         npu_inst_pe_1_7_3_int_q_reg_h_1__0_,
         npu_inst_pe_1_7_3_int_q_reg_h_1__1_,
         npu_inst_pe_1_7_3_int_q_reg_h_0__0_,
         npu_inst_pe_1_7_3_int_q_reg_h_0__1_, npu_inst_pe_1_7_4_n119,
         npu_inst_pe_1_7_4_n118, npu_inst_pe_1_7_4_n117,
         npu_inst_pe_1_7_4_n116, npu_inst_pe_1_7_4_n115,
         npu_inst_pe_1_7_4_n114, npu_inst_pe_1_7_4_n113,
         npu_inst_pe_1_7_4_n112, npu_inst_pe_1_7_4_n111,
         npu_inst_pe_1_7_4_n110, npu_inst_pe_1_7_4_n109,
         npu_inst_pe_1_7_4_n108, npu_inst_pe_1_7_4_n107,
         npu_inst_pe_1_7_4_n106, npu_inst_pe_1_7_4_n105,
         npu_inst_pe_1_7_4_n104, npu_inst_pe_1_7_4_n103,
         npu_inst_pe_1_7_4_n102, npu_inst_pe_1_7_4_n101,
         npu_inst_pe_1_7_4_n100, npu_inst_pe_1_7_4_n99, npu_inst_pe_1_7_4_n98,
         npu_inst_pe_1_7_4_n36, npu_inst_pe_1_7_4_n35, npu_inst_pe_1_7_4_n34,
         npu_inst_pe_1_7_4_n33, npu_inst_pe_1_7_4_n32, npu_inst_pe_1_7_4_n31,
         npu_inst_pe_1_7_4_n30, npu_inst_pe_1_7_4_n29, npu_inst_pe_1_7_4_n28,
         npu_inst_pe_1_7_4_n25, npu_inst_pe_1_7_4_n24, npu_inst_pe_1_7_4_n23,
         npu_inst_pe_1_7_4_n22, npu_inst_pe_1_7_4_n21, npu_inst_pe_1_7_4_n20,
         npu_inst_pe_1_7_4_n19, npu_inst_pe_1_7_4_n18, npu_inst_pe_1_7_4_n17,
         npu_inst_pe_1_7_4_n16, npu_inst_pe_1_7_4_n15, npu_inst_pe_1_7_4_n14,
         npu_inst_pe_1_7_4_n13, npu_inst_pe_1_7_4_n12, npu_inst_pe_1_7_4_n11,
         npu_inst_pe_1_7_4_n10, npu_inst_pe_1_7_4_n9, npu_inst_pe_1_7_4_n8,
         npu_inst_pe_1_7_4_n7, npu_inst_pe_1_7_4_n6, npu_inst_pe_1_7_4_n5,
         npu_inst_pe_1_7_4_n4, npu_inst_pe_1_7_4_n3, npu_inst_pe_1_7_4_n2,
         npu_inst_pe_1_7_4_n1, npu_inst_pe_1_7_4_sub_67_carry_7_,
         npu_inst_pe_1_7_4_sub_67_carry_6_, npu_inst_pe_1_7_4_sub_67_carry_5_,
         npu_inst_pe_1_7_4_sub_67_carry_4_, npu_inst_pe_1_7_4_sub_67_carry_3_,
         npu_inst_pe_1_7_4_sub_67_carry_2_, npu_inst_pe_1_7_4_sub_67_carry_1_,
         npu_inst_pe_1_7_4_add_69_carry_7_, npu_inst_pe_1_7_4_add_69_carry_6_,
         npu_inst_pe_1_7_4_add_69_carry_5_, npu_inst_pe_1_7_4_add_69_carry_4_,
         npu_inst_pe_1_7_4_add_69_carry_3_, npu_inst_pe_1_7_4_add_69_carry_2_,
         npu_inst_pe_1_7_4_add_69_carry_1_, npu_inst_pe_1_7_4_n97,
         npu_inst_pe_1_7_4_n96, npu_inst_pe_1_7_4_n95, npu_inst_pe_1_7_4_n94,
         npu_inst_pe_1_7_4_n93, npu_inst_pe_1_7_4_n92, npu_inst_pe_1_7_4_n91,
         npu_inst_pe_1_7_4_n90, npu_inst_pe_1_7_4_n89, npu_inst_pe_1_7_4_n88,
         npu_inst_pe_1_7_4_n87, npu_inst_pe_1_7_4_n86, npu_inst_pe_1_7_4_n85,
         npu_inst_pe_1_7_4_n84, npu_inst_pe_1_7_4_n83, npu_inst_pe_1_7_4_n82,
         npu_inst_pe_1_7_4_n81, npu_inst_pe_1_7_4_n80, npu_inst_pe_1_7_4_n79,
         npu_inst_pe_1_7_4_n78, npu_inst_pe_1_7_4_n77, npu_inst_pe_1_7_4_n76,
         npu_inst_pe_1_7_4_n75, npu_inst_pe_1_7_4_n74, npu_inst_pe_1_7_4_n73,
         npu_inst_pe_1_7_4_n72, npu_inst_pe_1_7_4_n71, npu_inst_pe_1_7_4_n70,
         npu_inst_pe_1_7_4_n69, npu_inst_pe_1_7_4_n68, npu_inst_pe_1_7_4_n67,
         npu_inst_pe_1_7_4_n66, npu_inst_pe_1_7_4_n65, npu_inst_pe_1_7_4_n64,
         npu_inst_pe_1_7_4_n63, npu_inst_pe_1_7_4_n62, npu_inst_pe_1_7_4_n61,
         npu_inst_pe_1_7_4_n60, npu_inst_pe_1_7_4_n59, npu_inst_pe_1_7_4_n58,
         npu_inst_pe_1_7_4_n57, npu_inst_pe_1_7_4_n56, npu_inst_pe_1_7_4_n55,
         npu_inst_pe_1_7_4_n54, npu_inst_pe_1_7_4_n53, npu_inst_pe_1_7_4_n52,
         npu_inst_pe_1_7_4_n51, npu_inst_pe_1_7_4_n50, npu_inst_pe_1_7_4_n49,
         npu_inst_pe_1_7_4_n48, npu_inst_pe_1_7_4_n47, npu_inst_pe_1_7_4_n46,
         npu_inst_pe_1_7_4_n45, npu_inst_pe_1_7_4_n44, npu_inst_pe_1_7_4_n43,
         npu_inst_pe_1_7_4_n42, npu_inst_pe_1_7_4_n41, npu_inst_pe_1_7_4_n40,
         npu_inst_pe_1_7_4_n39, npu_inst_pe_1_7_4_n38, npu_inst_pe_1_7_4_n37,
         npu_inst_pe_1_7_4_n27, npu_inst_pe_1_7_4_n26,
         npu_inst_pe_1_7_4_net3188, npu_inst_pe_1_7_4_net3182,
         npu_inst_pe_1_7_4_N94, npu_inst_pe_1_7_4_N93, npu_inst_pe_1_7_4_N84,
         npu_inst_pe_1_7_4_N80, npu_inst_pe_1_7_4_N79, npu_inst_pe_1_7_4_N78,
         npu_inst_pe_1_7_4_N77, npu_inst_pe_1_7_4_N76, npu_inst_pe_1_7_4_N75,
         npu_inst_pe_1_7_4_N74, npu_inst_pe_1_7_4_N73, npu_inst_pe_1_7_4_N72,
         npu_inst_pe_1_7_4_N71, npu_inst_pe_1_7_4_N70, npu_inst_pe_1_7_4_N69,
         npu_inst_pe_1_7_4_N68, npu_inst_pe_1_7_4_N67, npu_inst_pe_1_7_4_N66,
         npu_inst_pe_1_7_4_N65, npu_inst_pe_1_7_4_int_q_acc_0_,
         npu_inst_pe_1_7_4_int_q_acc_1_, npu_inst_pe_1_7_4_int_q_acc_2_,
         npu_inst_pe_1_7_4_int_q_acc_3_, npu_inst_pe_1_7_4_int_q_acc_4_,
         npu_inst_pe_1_7_4_int_q_acc_5_, npu_inst_pe_1_7_4_int_q_acc_6_,
         npu_inst_pe_1_7_4_int_q_acc_7_, npu_inst_pe_1_7_4_int_data_0_,
         npu_inst_pe_1_7_4_int_data_1_, npu_inst_pe_1_7_4_int_q_weight_0_,
         npu_inst_pe_1_7_4_int_q_weight_1_,
         npu_inst_pe_1_7_4_int_q_reg_v_5__0_,
         npu_inst_pe_1_7_4_int_q_reg_v_5__1_,
         npu_inst_pe_1_7_4_int_q_reg_v_4__0_,
         npu_inst_pe_1_7_4_int_q_reg_v_4__1_,
         npu_inst_pe_1_7_4_int_q_reg_v_3__0_,
         npu_inst_pe_1_7_4_int_q_reg_v_3__1_,
         npu_inst_pe_1_7_4_int_q_reg_v_2__0_,
         npu_inst_pe_1_7_4_int_q_reg_v_2__1_,
         npu_inst_pe_1_7_4_int_q_reg_v_1__0_,
         npu_inst_pe_1_7_4_int_q_reg_v_1__1_,
         npu_inst_pe_1_7_4_int_q_reg_v_0__0_,
         npu_inst_pe_1_7_4_int_q_reg_v_0__1_,
         npu_inst_pe_1_7_4_int_q_reg_h_5__0_,
         npu_inst_pe_1_7_4_int_q_reg_h_5__1_,
         npu_inst_pe_1_7_4_int_q_reg_h_4__0_,
         npu_inst_pe_1_7_4_int_q_reg_h_4__1_,
         npu_inst_pe_1_7_4_int_q_reg_h_3__0_,
         npu_inst_pe_1_7_4_int_q_reg_h_3__1_,
         npu_inst_pe_1_7_4_int_q_reg_h_2__0_,
         npu_inst_pe_1_7_4_int_q_reg_h_2__1_,
         npu_inst_pe_1_7_4_int_q_reg_h_1__0_,
         npu_inst_pe_1_7_4_int_q_reg_h_1__1_,
         npu_inst_pe_1_7_4_int_q_reg_h_0__0_,
         npu_inst_pe_1_7_4_int_q_reg_h_0__1_, npu_inst_pe_1_7_5_n119,
         npu_inst_pe_1_7_5_n118, npu_inst_pe_1_7_5_n117,
         npu_inst_pe_1_7_5_n116, npu_inst_pe_1_7_5_n115,
         npu_inst_pe_1_7_5_n114, npu_inst_pe_1_7_5_n113,
         npu_inst_pe_1_7_5_n112, npu_inst_pe_1_7_5_n111,
         npu_inst_pe_1_7_5_n110, npu_inst_pe_1_7_5_n109,
         npu_inst_pe_1_7_5_n108, npu_inst_pe_1_7_5_n107,
         npu_inst_pe_1_7_5_n106, npu_inst_pe_1_7_5_n105,
         npu_inst_pe_1_7_5_n104, npu_inst_pe_1_7_5_n103,
         npu_inst_pe_1_7_5_n102, npu_inst_pe_1_7_5_n101,
         npu_inst_pe_1_7_5_n100, npu_inst_pe_1_7_5_n99, npu_inst_pe_1_7_5_n98,
         npu_inst_pe_1_7_5_n36, npu_inst_pe_1_7_5_n35, npu_inst_pe_1_7_5_n34,
         npu_inst_pe_1_7_5_n33, npu_inst_pe_1_7_5_n32, npu_inst_pe_1_7_5_n31,
         npu_inst_pe_1_7_5_n30, npu_inst_pe_1_7_5_n29, npu_inst_pe_1_7_5_n28,
         npu_inst_pe_1_7_5_n25, npu_inst_pe_1_7_5_n24, npu_inst_pe_1_7_5_n23,
         npu_inst_pe_1_7_5_n22, npu_inst_pe_1_7_5_n21, npu_inst_pe_1_7_5_n20,
         npu_inst_pe_1_7_5_n19, npu_inst_pe_1_7_5_n18, npu_inst_pe_1_7_5_n17,
         npu_inst_pe_1_7_5_n16, npu_inst_pe_1_7_5_n15, npu_inst_pe_1_7_5_n14,
         npu_inst_pe_1_7_5_n13, npu_inst_pe_1_7_5_n12, npu_inst_pe_1_7_5_n11,
         npu_inst_pe_1_7_5_n10, npu_inst_pe_1_7_5_n9, npu_inst_pe_1_7_5_n8,
         npu_inst_pe_1_7_5_n7, npu_inst_pe_1_7_5_n6, npu_inst_pe_1_7_5_n5,
         npu_inst_pe_1_7_5_n4, npu_inst_pe_1_7_5_n3, npu_inst_pe_1_7_5_n2,
         npu_inst_pe_1_7_5_n1, npu_inst_pe_1_7_5_sub_67_carry_7_,
         npu_inst_pe_1_7_5_sub_67_carry_6_, npu_inst_pe_1_7_5_sub_67_carry_5_,
         npu_inst_pe_1_7_5_sub_67_carry_4_, npu_inst_pe_1_7_5_sub_67_carry_3_,
         npu_inst_pe_1_7_5_sub_67_carry_2_, npu_inst_pe_1_7_5_sub_67_carry_1_,
         npu_inst_pe_1_7_5_add_69_carry_7_, npu_inst_pe_1_7_5_add_69_carry_6_,
         npu_inst_pe_1_7_5_add_69_carry_5_, npu_inst_pe_1_7_5_add_69_carry_4_,
         npu_inst_pe_1_7_5_add_69_carry_3_, npu_inst_pe_1_7_5_add_69_carry_2_,
         npu_inst_pe_1_7_5_add_69_carry_1_, npu_inst_pe_1_7_5_n97,
         npu_inst_pe_1_7_5_n96, npu_inst_pe_1_7_5_n95, npu_inst_pe_1_7_5_n94,
         npu_inst_pe_1_7_5_n93, npu_inst_pe_1_7_5_n92, npu_inst_pe_1_7_5_n91,
         npu_inst_pe_1_7_5_n90, npu_inst_pe_1_7_5_n89, npu_inst_pe_1_7_5_n88,
         npu_inst_pe_1_7_5_n87, npu_inst_pe_1_7_5_n86, npu_inst_pe_1_7_5_n85,
         npu_inst_pe_1_7_5_n84, npu_inst_pe_1_7_5_n83, npu_inst_pe_1_7_5_n82,
         npu_inst_pe_1_7_5_n81, npu_inst_pe_1_7_5_n80, npu_inst_pe_1_7_5_n79,
         npu_inst_pe_1_7_5_n78, npu_inst_pe_1_7_5_n77, npu_inst_pe_1_7_5_n76,
         npu_inst_pe_1_7_5_n75, npu_inst_pe_1_7_5_n74, npu_inst_pe_1_7_5_n73,
         npu_inst_pe_1_7_5_n72, npu_inst_pe_1_7_5_n71, npu_inst_pe_1_7_5_n70,
         npu_inst_pe_1_7_5_n69, npu_inst_pe_1_7_5_n68, npu_inst_pe_1_7_5_n67,
         npu_inst_pe_1_7_5_n66, npu_inst_pe_1_7_5_n65, npu_inst_pe_1_7_5_n64,
         npu_inst_pe_1_7_5_n63, npu_inst_pe_1_7_5_n62, npu_inst_pe_1_7_5_n61,
         npu_inst_pe_1_7_5_n60, npu_inst_pe_1_7_5_n59, npu_inst_pe_1_7_5_n58,
         npu_inst_pe_1_7_5_n57, npu_inst_pe_1_7_5_n56, npu_inst_pe_1_7_5_n55,
         npu_inst_pe_1_7_5_n54, npu_inst_pe_1_7_5_n53, npu_inst_pe_1_7_5_n52,
         npu_inst_pe_1_7_5_n51, npu_inst_pe_1_7_5_n50, npu_inst_pe_1_7_5_n49,
         npu_inst_pe_1_7_5_n48, npu_inst_pe_1_7_5_n47, npu_inst_pe_1_7_5_n46,
         npu_inst_pe_1_7_5_n45, npu_inst_pe_1_7_5_n44, npu_inst_pe_1_7_5_n43,
         npu_inst_pe_1_7_5_n42, npu_inst_pe_1_7_5_n41, npu_inst_pe_1_7_5_n40,
         npu_inst_pe_1_7_5_n39, npu_inst_pe_1_7_5_n38, npu_inst_pe_1_7_5_n37,
         npu_inst_pe_1_7_5_n27, npu_inst_pe_1_7_5_n26,
         npu_inst_pe_1_7_5_net3165, npu_inst_pe_1_7_5_net3159,
         npu_inst_pe_1_7_5_N94, npu_inst_pe_1_7_5_N93, npu_inst_pe_1_7_5_N84,
         npu_inst_pe_1_7_5_N80, npu_inst_pe_1_7_5_N79, npu_inst_pe_1_7_5_N78,
         npu_inst_pe_1_7_5_N77, npu_inst_pe_1_7_5_N76, npu_inst_pe_1_7_5_N75,
         npu_inst_pe_1_7_5_N74, npu_inst_pe_1_7_5_N73, npu_inst_pe_1_7_5_N72,
         npu_inst_pe_1_7_5_N71, npu_inst_pe_1_7_5_N70, npu_inst_pe_1_7_5_N69,
         npu_inst_pe_1_7_5_N68, npu_inst_pe_1_7_5_N67, npu_inst_pe_1_7_5_N66,
         npu_inst_pe_1_7_5_N65, npu_inst_pe_1_7_5_int_q_acc_0_,
         npu_inst_pe_1_7_5_int_q_acc_1_, npu_inst_pe_1_7_5_int_q_acc_2_,
         npu_inst_pe_1_7_5_int_q_acc_3_, npu_inst_pe_1_7_5_int_q_acc_4_,
         npu_inst_pe_1_7_5_int_q_acc_5_, npu_inst_pe_1_7_5_int_q_acc_6_,
         npu_inst_pe_1_7_5_int_q_acc_7_, npu_inst_pe_1_7_5_int_data_0_,
         npu_inst_pe_1_7_5_int_data_1_, npu_inst_pe_1_7_5_int_q_weight_0_,
         npu_inst_pe_1_7_5_int_q_weight_1_,
         npu_inst_pe_1_7_5_int_q_reg_v_5__0_,
         npu_inst_pe_1_7_5_int_q_reg_v_5__1_,
         npu_inst_pe_1_7_5_int_q_reg_v_4__0_,
         npu_inst_pe_1_7_5_int_q_reg_v_4__1_,
         npu_inst_pe_1_7_5_int_q_reg_v_3__0_,
         npu_inst_pe_1_7_5_int_q_reg_v_3__1_,
         npu_inst_pe_1_7_5_int_q_reg_v_2__0_,
         npu_inst_pe_1_7_5_int_q_reg_v_2__1_,
         npu_inst_pe_1_7_5_int_q_reg_v_1__0_,
         npu_inst_pe_1_7_5_int_q_reg_v_1__1_,
         npu_inst_pe_1_7_5_int_q_reg_v_0__0_,
         npu_inst_pe_1_7_5_int_q_reg_v_0__1_,
         npu_inst_pe_1_7_5_int_q_reg_h_5__0_,
         npu_inst_pe_1_7_5_int_q_reg_h_5__1_,
         npu_inst_pe_1_7_5_int_q_reg_h_4__0_,
         npu_inst_pe_1_7_5_int_q_reg_h_4__1_,
         npu_inst_pe_1_7_5_int_q_reg_h_3__0_,
         npu_inst_pe_1_7_5_int_q_reg_h_3__1_,
         npu_inst_pe_1_7_5_int_q_reg_h_2__0_,
         npu_inst_pe_1_7_5_int_q_reg_h_2__1_,
         npu_inst_pe_1_7_5_int_q_reg_h_1__0_,
         npu_inst_pe_1_7_5_int_q_reg_h_1__1_,
         npu_inst_pe_1_7_5_int_q_reg_h_0__0_,
         npu_inst_pe_1_7_5_int_q_reg_h_0__1_, npu_inst_pe_1_7_6_n119,
         npu_inst_pe_1_7_6_n118, npu_inst_pe_1_7_6_n117,
         npu_inst_pe_1_7_6_n116, npu_inst_pe_1_7_6_n115,
         npu_inst_pe_1_7_6_n114, npu_inst_pe_1_7_6_n113,
         npu_inst_pe_1_7_6_n112, npu_inst_pe_1_7_6_n111,
         npu_inst_pe_1_7_6_n110, npu_inst_pe_1_7_6_n109,
         npu_inst_pe_1_7_6_n108, npu_inst_pe_1_7_6_n107,
         npu_inst_pe_1_7_6_n106, npu_inst_pe_1_7_6_n105,
         npu_inst_pe_1_7_6_n104, npu_inst_pe_1_7_6_n103,
         npu_inst_pe_1_7_6_n102, npu_inst_pe_1_7_6_n101,
         npu_inst_pe_1_7_6_n100, npu_inst_pe_1_7_6_n99, npu_inst_pe_1_7_6_n98,
         npu_inst_pe_1_7_6_n36, npu_inst_pe_1_7_6_n35, npu_inst_pe_1_7_6_n34,
         npu_inst_pe_1_7_6_n33, npu_inst_pe_1_7_6_n32, npu_inst_pe_1_7_6_n31,
         npu_inst_pe_1_7_6_n30, npu_inst_pe_1_7_6_n29, npu_inst_pe_1_7_6_n28,
         npu_inst_pe_1_7_6_n25, npu_inst_pe_1_7_6_n24, npu_inst_pe_1_7_6_n23,
         npu_inst_pe_1_7_6_n22, npu_inst_pe_1_7_6_n21, npu_inst_pe_1_7_6_n20,
         npu_inst_pe_1_7_6_n19, npu_inst_pe_1_7_6_n18, npu_inst_pe_1_7_6_n17,
         npu_inst_pe_1_7_6_n16, npu_inst_pe_1_7_6_n15, npu_inst_pe_1_7_6_n14,
         npu_inst_pe_1_7_6_n13, npu_inst_pe_1_7_6_n12, npu_inst_pe_1_7_6_n11,
         npu_inst_pe_1_7_6_n10, npu_inst_pe_1_7_6_n9, npu_inst_pe_1_7_6_n8,
         npu_inst_pe_1_7_6_n7, npu_inst_pe_1_7_6_n6, npu_inst_pe_1_7_6_n5,
         npu_inst_pe_1_7_6_n4, npu_inst_pe_1_7_6_n3, npu_inst_pe_1_7_6_n2,
         npu_inst_pe_1_7_6_n1, npu_inst_pe_1_7_6_sub_67_carry_7_,
         npu_inst_pe_1_7_6_sub_67_carry_6_, npu_inst_pe_1_7_6_sub_67_carry_5_,
         npu_inst_pe_1_7_6_sub_67_carry_4_, npu_inst_pe_1_7_6_sub_67_carry_3_,
         npu_inst_pe_1_7_6_sub_67_carry_2_, npu_inst_pe_1_7_6_sub_67_carry_1_,
         npu_inst_pe_1_7_6_add_69_carry_7_, npu_inst_pe_1_7_6_add_69_carry_6_,
         npu_inst_pe_1_7_6_add_69_carry_5_, npu_inst_pe_1_7_6_add_69_carry_4_,
         npu_inst_pe_1_7_6_add_69_carry_3_, npu_inst_pe_1_7_6_add_69_carry_2_,
         npu_inst_pe_1_7_6_add_69_carry_1_, npu_inst_pe_1_7_6_n97,
         npu_inst_pe_1_7_6_n96, npu_inst_pe_1_7_6_n95, npu_inst_pe_1_7_6_n94,
         npu_inst_pe_1_7_6_n93, npu_inst_pe_1_7_6_n92, npu_inst_pe_1_7_6_n91,
         npu_inst_pe_1_7_6_n90, npu_inst_pe_1_7_6_n89, npu_inst_pe_1_7_6_n88,
         npu_inst_pe_1_7_6_n87, npu_inst_pe_1_7_6_n86, npu_inst_pe_1_7_6_n85,
         npu_inst_pe_1_7_6_n84, npu_inst_pe_1_7_6_n83, npu_inst_pe_1_7_6_n82,
         npu_inst_pe_1_7_6_n81, npu_inst_pe_1_7_6_n80, npu_inst_pe_1_7_6_n79,
         npu_inst_pe_1_7_6_n78, npu_inst_pe_1_7_6_n77, npu_inst_pe_1_7_6_n76,
         npu_inst_pe_1_7_6_n75, npu_inst_pe_1_7_6_n74, npu_inst_pe_1_7_6_n73,
         npu_inst_pe_1_7_6_n72, npu_inst_pe_1_7_6_n71, npu_inst_pe_1_7_6_n70,
         npu_inst_pe_1_7_6_n69, npu_inst_pe_1_7_6_n68, npu_inst_pe_1_7_6_n67,
         npu_inst_pe_1_7_6_n66, npu_inst_pe_1_7_6_n65, npu_inst_pe_1_7_6_n64,
         npu_inst_pe_1_7_6_n63, npu_inst_pe_1_7_6_n62, npu_inst_pe_1_7_6_n61,
         npu_inst_pe_1_7_6_n60, npu_inst_pe_1_7_6_n59, npu_inst_pe_1_7_6_n58,
         npu_inst_pe_1_7_6_n57, npu_inst_pe_1_7_6_n56, npu_inst_pe_1_7_6_n55,
         npu_inst_pe_1_7_6_n54, npu_inst_pe_1_7_6_n53, npu_inst_pe_1_7_6_n52,
         npu_inst_pe_1_7_6_n51, npu_inst_pe_1_7_6_n50, npu_inst_pe_1_7_6_n49,
         npu_inst_pe_1_7_6_n48, npu_inst_pe_1_7_6_n47, npu_inst_pe_1_7_6_n46,
         npu_inst_pe_1_7_6_n45, npu_inst_pe_1_7_6_n44, npu_inst_pe_1_7_6_n43,
         npu_inst_pe_1_7_6_n42, npu_inst_pe_1_7_6_n41, npu_inst_pe_1_7_6_n40,
         npu_inst_pe_1_7_6_n39, npu_inst_pe_1_7_6_n38, npu_inst_pe_1_7_6_n37,
         npu_inst_pe_1_7_6_n27, npu_inst_pe_1_7_6_n26,
         npu_inst_pe_1_7_6_net3142, npu_inst_pe_1_7_6_net3136,
         npu_inst_pe_1_7_6_N94, npu_inst_pe_1_7_6_N93, npu_inst_pe_1_7_6_N84,
         npu_inst_pe_1_7_6_N80, npu_inst_pe_1_7_6_N79, npu_inst_pe_1_7_6_N78,
         npu_inst_pe_1_7_6_N77, npu_inst_pe_1_7_6_N76, npu_inst_pe_1_7_6_N75,
         npu_inst_pe_1_7_6_N74, npu_inst_pe_1_7_6_N73, npu_inst_pe_1_7_6_N72,
         npu_inst_pe_1_7_6_N71, npu_inst_pe_1_7_6_N70, npu_inst_pe_1_7_6_N69,
         npu_inst_pe_1_7_6_N68, npu_inst_pe_1_7_6_N67, npu_inst_pe_1_7_6_N66,
         npu_inst_pe_1_7_6_N65, npu_inst_pe_1_7_6_int_q_acc_0_,
         npu_inst_pe_1_7_6_int_q_acc_1_, npu_inst_pe_1_7_6_int_q_acc_2_,
         npu_inst_pe_1_7_6_int_q_acc_3_, npu_inst_pe_1_7_6_int_q_acc_4_,
         npu_inst_pe_1_7_6_int_q_acc_5_, npu_inst_pe_1_7_6_int_q_acc_6_,
         npu_inst_pe_1_7_6_int_q_acc_7_, npu_inst_pe_1_7_6_int_data_0_,
         npu_inst_pe_1_7_6_int_data_1_, npu_inst_pe_1_7_6_int_q_weight_0_,
         npu_inst_pe_1_7_6_int_q_weight_1_,
         npu_inst_pe_1_7_6_int_q_reg_v_5__0_,
         npu_inst_pe_1_7_6_int_q_reg_v_5__1_,
         npu_inst_pe_1_7_6_int_q_reg_v_4__0_,
         npu_inst_pe_1_7_6_int_q_reg_v_4__1_,
         npu_inst_pe_1_7_6_int_q_reg_v_3__0_,
         npu_inst_pe_1_7_6_int_q_reg_v_3__1_,
         npu_inst_pe_1_7_6_int_q_reg_v_2__0_,
         npu_inst_pe_1_7_6_int_q_reg_v_2__1_,
         npu_inst_pe_1_7_6_int_q_reg_v_1__0_,
         npu_inst_pe_1_7_6_int_q_reg_v_1__1_,
         npu_inst_pe_1_7_6_int_q_reg_v_0__0_,
         npu_inst_pe_1_7_6_int_q_reg_v_0__1_,
         npu_inst_pe_1_7_6_int_q_reg_h_5__0_,
         npu_inst_pe_1_7_6_int_q_reg_h_5__1_,
         npu_inst_pe_1_7_6_int_q_reg_h_4__0_,
         npu_inst_pe_1_7_6_int_q_reg_h_4__1_,
         npu_inst_pe_1_7_6_int_q_reg_h_3__0_,
         npu_inst_pe_1_7_6_int_q_reg_h_3__1_,
         npu_inst_pe_1_7_6_int_q_reg_h_2__0_,
         npu_inst_pe_1_7_6_int_q_reg_h_2__1_,
         npu_inst_pe_1_7_6_int_q_reg_h_1__0_,
         npu_inst_pe_1_7_6_int_q_reg_h_1__1_,
         npu_inst_pe_1_7_6_int_q_reg_h_0__0_,
         npu_inst_pe_1_7_6_int_q_reg_h_0__1_, npu_inst_pe_1_7_7_n119,
         npu_inst_pe_1_7_7_n118, npu_inst_pe_1_7_7_n117,
         npu_inst_pe_1_7_7_n116, npu_inst_pe_1_7_7_n115,
         npu_inst_pe_1_7_7_n114, npu_inst_pe_1_7_7_n113,
         npu_inst_pe_1_7_7_n112, npu_inst_pe_1_7_7_n111,
         npu_inst_pe_1_7_7_n110, npu_inst_pe_1_7_7_n109,
         npu_inst_pe_1_7_7_n108, npu_inst_pe_1_7_7_n107,
         npu_inst_pe_1_7_7_n106, npu_inst_pe_1_7_7_n105,
         npu_inst_pe_1_7_7_n104, npu_inst_pe_1_7_7_n103,
         npu_inst_pe_1_7_7_n102, npu_inst_pe_1_7_7_n101,
         npu_inst_pe_1_7_7_n100, npu_inst_pe_1_7_7_n99, npu_inst_pe_1_7_7_n98,
         npu_inst_pe_1_7_7_n36, npu_inst_pe_1_7_7_n35, npu_inst_pe_1_7_7_n34,
         npu_inst_pe_1_7_7_n33, npu_inst_pe_1_7_7_n32, npu_inst_pe_1_7_7_n31,
         npu_inst_pe_1_7_7_n30, npu_inst_pe_1_7_7_n29, npu_inst_pe_1_7_7_n28,
         npu_inst_pe_1_7_7_n25, npu_inst_pe_1_7_7_n24, npu_inst_pe_1_7_7_n23,
         npu_inst_pe_1_7_7_n22, npu_inst_pe_1_7_7_n21, npu_inst_pe_1_7_7_n20,
         npu_inst_pe_1_7_7_n19, npu_inst_pe_1_7_7_n18, npu_inst_pe_1_7_7_n17,
         npu_inst_pe_1_7_7_n16, npu_inst_pe_1_7_7_n15, npu_inst_pe_1_7_7_n14,
         npu_inst_pe_1_7_7_n13, npu_inst_pe_1_7_7_n12, npu_inst_pe_1_7_7_n11,
         npu_inst_pe_1_7_7_n10, npu_inst_pe_1_7_7_n9, npu_inst_pe_1_7_7_n8,
         npu_inst_pe_1_7_7_n7, npu_inst_pe_1_7_7_n6, npu_inst_pe_1_7_7_n5,
         npu_inst_pe_1_7_7_n4, npu_inst_pe_1_7_7_n3, npu_inst_pe_1_7_7_n2,
         npu_inst_pe_1_7_7_n1, npu_inst_pe_1_7_7_sub_67_carry_7_,
         npu_inst_pe_1_7_7_sub_67_carry_6_, npu_inst_pe_1_7_7_sub_67_carry_5_,
         npu_inst_pe_1_7_7_sub_67_carry_4_, npu_inst_pe_1_7_7_sub_67_carry_3_,
         npu_inst_pe_1_7_7_sub_67_carry_2_, npu_inst_pe_1_7_7_sub_67_carry_1_,
         npu_inst_pe_1_7_7_add_69_carry_7_, npu_inst_pe_1_7_7_add_69_carry_6_,
         npu_inst_pe_1_7_7_add_69_carry_5_, npu_inst_pe_1_7_7_add_69_carry_4_,
         npu_inst_pe_1_7_7_add_69_carry_3_, npu_inst_pe_1_7_7_add_69_carry_2_,
         npu_inst_pe_1_7_7_add_69_carry_1_, npu_inst_pe_1_7_7_n97,
         npu_inst_pe_1_7_7_n96, npu_inst_pe_1_7_7_n95, npu_inst_pe_1_7_7_n94,
         npu_inst_pe_1_7_7_n93, npu_inst_pe_1_7_7_n92, npu_inst_pe_1_7_7_n91,
         npu_inst_pe_1_7_7_n90, npu_inst_pe_1_7_7_n89, npu_inst_pe_1_7_7_n88,
         npu_inst_pe_1_7_7_n87, npu_inst_pe_1_7_7_n86, npu_inst_pe_1_7_7_n85,
         npu_inst_pe_1_7_7_n84, npu_inst_pe_1_7_7_n83, npu_inst_pe_1_7_7_n82,
         npu_inst_pe_1_7_7_n81, npu_inst_pe_1_7_7_n80, npu_inst_pe_1_7_7_n79,
         npu_inst_pe_1_7_7_n78, npu_inst_pe_1_7_7_n77, npu_inst_pe_1_7_7_n76,
         npu_inst_pe_1_7_7_n75, npu_inst_pe_1_7_7_n74, npu_inst_pe_1_7_7_n73,
         npu_inst_pe_1_7_7_n72, npu_inst_pe_1_7_7_n71, npu_inst_pe_1_7_7_n70,
         npu_inst_pe_1_7_7_n69, npu_inst_pe_1_7_7_n68, npu_inst_pe_1_7_7_n67,
         npu_inst_pe_1_7_7_n66, npu_inst_pe_1_7_7_n65, npu_inst_pe_1_7_7_n64,
         npu_inst_pe_1_7_7_n63, npu_inst_pe_1_7_7_n62, npu_inst_pe_1_7_7_n61,
         npu_inst_pe_1_7_7_n60, npu_inst_pe_1_7_7_n59, npu_inst_pe_1_7_7_n58,
         npu_inst_pe_1_7_7_n57, npu_inst_pe_1_7_7_n56, npu_inst_pe_1_7_7_n55,
         npu_inst_pe_1_7_7_n54, npu_inst_pe_1_7_7_n53, npu_inst_pe_1_7_7_n52,
         npu_inst_pe_1_7_7_n51, npu_inst_pe_1_7_7_n50, npu_inst_pe_1_7_7_n49,
         npu_inst_pe_1_7_7_n48, npu_inst_pe_1_7_7_n47, npu_inst_pe_1_7_7_n46,
         npu_inst_pe_1_7_7_n45, npu_inst_pe_1_7_7_n44, npu_inst_pe_1_7_7_n43,
         npu_inst_pe_1_7_7_n42, npu_inst_pe_1_7_7_n41, npu_inst_pe_1_7_7_n40,
         npu_inst_pe_1_7_7_n39, npu_inst_pe_1_7_7_n38, npu_inst_pe_1_7_7_n37,
         npu_inst_pe_1_7_7_n27, npu_inst_pe_1_7_7_n26,
         npu_inst_pe_1_7_7_net3119, npu_inst_pe_1_7_7_net3113,
         npu_inst_pe_1_7_7_N94, npu_inst_pe_1_7_7_N93, npu_inst_pe_1_7_7_N84,
         npu_inst_pe_1_7_7_N80, npu_inst_pe_1_7_7_N79, npu_inst_pe_1_7_7_N78,
         npu_inst_pe_1_7_7_N77, npu_inst_pe_1_7_7_N76, npu_inst_pe_1_7_7_N75,
         npu_inst_pe_1_7_7_N74, npu_inst_pe_1_7_7_N73, npu_inst_pe_1_7_7_N72,
         npu_inst_pe_1_7_7_N71, npu_inst_pe_1_7_7_N70, npu_inst_pe_1_7_7_N69,
         npu_inst_pe_1_7_7_N68, npu_inst_pe_1_7_7_N67, npu_inst_pe_1_7_7_N66,
         npu_inst_pe_1_7_7_N65, npu_inst_pe_1_7_7_int_q_acc_0_,
         npu_inst_pe_1_7_7_int_q_acc_1_, npu_inst_pe_1_7_7_int_q_acc_2_,
         npu_inst_pe_1_7_7_int_q_acc_3_, npu_inst_pe_1_7_7_int_q_acc_4_,
         npu_inst_pe_1_7_7_int_q_acc_5_, npu_inst_pe_1_7_7_int_q_acc_6_,
         npu_inst_pe_1_7_7_int_q_acc_7_, npu_inst_pe_1_7_7_int_data_0_,
         npu_inst_pe_1_7_7_int_data_1_, npu_inst_pe_1_7_7_int_q_weight_0_,
         npu_inst_pe_1_7_7_int_q_weight_1_,
         npu_inst_pe_1_7_7_int_q_reg_v_5__0_,
         npu_inst_pe_1_7_7_int_q_reg_v_5__1_,
         npu_inst_pe_1_7_7_int_q_reg_v_4__0_,
         npu_inst_pe_1_7_7_int_q_reg_v_4__1_,
         npu_inst_pe_1_7_7_int_q_reg_v_3__0_,
         npu_inst_pe_1_7_7_int_q_reg_v_3__1_,
         npu_inst_pe_1_7_7_int_q_reg_v_2__0_,
         npu_inst_pe_1_7_7_int_q_reg_v_2__1_,
         npu_inst_pe_1_7_7_int_q_reg_v_1__0_,
         npu_inst_pe_1_7_7_int_q_reg_v_1__1_,
         npu_inst_pe_1_7_7_int_q_reg_v_0__0_,
         npu_inst_pe_1_7_7_int_q_reg_v_0__1_,
         npu_inst_pe_1_7_7_int_q_reg_h_5__0_,
         npu_inst_pe_1_7_7_int_q_reg_h_5__1_,
         npu_inst_pe_1_7_7_int_q_reg_h_4__0_,
         npu_inst_pe_1_7_7_int_q_reg_h_4__1_,
         npu_inst_pe_1_7_7_int_q_reg_h_3__0_,
         npu_inst_pe_1_7_7_int_q_reg_h_3__1_,
         npu_inst_pe_1_7_7_int_q_reg_h_2__0_,
         npu_inst_pe_1_7_7_int_q_reg_h_2__1_,
         npu_inst_pe_1_7_7_int_q_reg_h_1__0_,
         npu_inst_pe_1_7_7_int_q_reg_h_1__1_,
         npu_inst_pe_1_7_7_int_q_reg_h_0__0_,
         npu_inst_pe_1_7_7_int_q_reg_h_0__1_, qrelu_i_0_n3, qrelu_i_0_n2,
         qrelu_i_0_n1, qrelu_i_0_n6, qrelu_i_0_n5, qrelu_i_0_n4, qrelu_i_1_n9,
         qrelu_i_1_n8, qrelu_i_1_n7, qrelu_i_1_n3, qrelu_i_1_n2, qrelu_i_1_n1,
         qrelu_i_2_n9, qrelu_i_2_n8, qrelu_i_2_n7, qrelu_i_2_n3, qrelu_i_2_n2,
         qrelu_i_2_n1, qrelu_i_3_n9, qrelu_i_3_n8, qrelu_i_3_n7, qrelu_i_3_n3,
         qrelu_i_3_n2, qrelu_i_3_n1, qrelu_i_4_n9, qrelu_i_4_n8, qrelu_i_4_n7,
         qrelu_i_4_n3, qrelu_i_4_n2, qrelu_i_4_n1, qrelu_i_5_n9, qrelu_i_5_n8,
         qrelu_i_5_n7, qrelu_i_5_n3, qrelu_i_5_n2, qrelu_i_5_n1, qrelu_i_6_n9,
         qrelu_i_6_n8, qrelu_i_6_n7, qrelu_i_6_n3, qrelu_i_6_n2, qrelu_i_6_n1,
         qrelu_i_7_n9, qrelu_i_7_n8, qrelu_i_7_n7, qrelu_i_7_n3, qrelu_i_7_n2,
         qrelu_i_7_n1, p_unit_i_0_n17, p_unit_i_0_n16, p_unit_i_0_n12,
         p_unit_i_0_n11, p_unit_i_0_n7, p_unit_i_0_n6, p_unit_i_0_n5,
         p_unit_i_0_n4, p_unit_i_0_n3, p_unit_i_0_n2, p_unit_i_0_n1,
         p_unit_i_0_n15, p_unit_i_0_n14, p_unit_i_0_n13, p_unit_i_0_n10,
         p_unit_i_0_n9, p_unit_i_0_n8, p_unit_i_0_net3095, p_unit_i_0_N7,
         p_unit_i_0_N6, p_unit_i_0_N5, p_unit_i_0_N3, p_unit_i_0_N2,
         p_unit_i_0_int_ps1_0_, p_unit_i_0_int_ps1_1_, p_unit_i_0_int_ps1_2_,
         p_unit_i_0_int_ps0_0_, p_unit_i_0_int_ps0_1_, p_unit_i_0_int_ps0_2_,
         p_unit_i_1_n17, p_unit_i_1_n16, p_unit_i_1_n12, p_unit_i_1_n11,
         p_unit_i_1_n7, p_unit_i_1_n6, p_unit_i_1_n5, p_unit_i_1_n4,
         p_unit_i_1_n3, p_unit_i_1_n2, p_unit_i_1_n1, p_unit_i_1_n15,
         p_unit_i_1_n14, p_unit_i_1_n13, p_unit_i_1_n10, p_unit_i_1_n9,
         p_unit_i_1_n8, p_unit_i_1_net3077, p_unit_i_1_N7, p_unit_i_1_N6,
         p_unit_i_1_N5, p_unit_i_1_N3, p_unit_i_1_N2, p_unit_i_1_int_ps1_0_,
         p_unit_i_1_int_ps1_1_, p_unit_i_1_int_ps1_2_, p_unit_i_1_int_ps0_0_,
         p_unit_i_1_int_ps0_1_, p_unit_i_1_int_ps0_2_, p_unit_i_2_n17,
         p_unit_i_2_n16, p_unit_i_2_n12, p_unit_i_2_n11, p_unit_i_2_n7,
         p_unit_i_2_n6, p_unit_i_2_n5, p_unit_i_2_n4, p_unit_i_2_n3,
         p_unit_i_2_n2, p_unit_i_2_n1, p_unit_i_2_n15, p_unit_i_2_n14,
         p_unit_i_2_n13, p_unit_i_2_n10, p_unit_i_2_n9, p_unit_i_2_n8,
         p_unit_i_2_net3059, p_unit_i_2_N7, p_unit_i_2_N6, p_unit_i_2_N5,
         p_unit_i_2_N3, p_unit_i_2_N2, p_unit_i_2_int_ps1_0_,
         p_unit_i_2_int_ps1_1_, p_unit_i_2_int_ps1_2_, p_unit_i_2_int_ps0_0_,
         p_unit_i_2_int_ps0_1_, p_unit_i_2_int_ps0_2_, p_unit_i_3_n17,
         p_unit_i_3_n16, p_unit_i_3_n12, p_unit_i_3_n11, p_unit_i_3_n7,
         p_unit_i_3_n6, p_unit_i_3_n5, p_unit_i_3_n4, p_unit_i_3_n3,
         p_unit_i_3_n2, p_unit_i_3_n1, p_unit_i_3_n15, p_unit_i_3_n14,
         p_unit_i_3_n13, p_unit_i_3_n10, p_unit_i_3_n9, p_unit_i_3_n8,
         p_unit_i_3_net3041, p_unit_i_3_N7, p_unit_i_3_N6, p_unit_i_3_N5,
         p_unit_i_3_N3, p_unit_i_3_N2, p_unit_i_3_int_ps1_0_,
         p_unit_i_3_int_ps1_1_, p_unit_i_3_int_ps1_2_, p_unit_i_3_int_ps0_0_,
         p_unit_i_3_int_ps0_1_, p_unit_i_3_int_ps0_2_, round_i_0_n2,
         round_i_0_n1, round_i_0_n3, round_i_1_n4, round_i_1_n2, round_i_1_n1,
         round_i_2_n4, round_i_2_n2, round_i_2_n1, round_i_3_n4, round_i_3_n2,
         round_i_3_n1, hmode_cnt_inst_n12, hmode_cnt_inst_n6,
         hmode_cnt_inst_n4, hmode_cnt_inst_n2, hmode_cnt_inst_n1,
         hmode_cnt_inst_n11, hmode_cnt_inst_n10, hmode_cnt_inst_n9,
         hmode_cnt_inst_n8, hmode_cnt_inst_n7, hmode_cnt_inst_n5,
         hmode_cnt_inst_net3023, hmode_cnt_inst_N12, hmode_cnt_inst_N10,
         vmode_cnt_inst_n12, vmode_cnt_inst_n6, vmode_cnt_inst_n4,
         vmode_cnt_inst_n2, vmode_cnt_inst_n1, vmode_cnt_inst_n11,
         vmode_cnt_inst_n10, vmode_cnt_inst_n9, vmode_cnt_inst_n8,
         vmode_cnt_inst_n7, vmode_cnt_inst_n5, vmode_cnt_inst_net3005,
         vmode_cnt_inst_N12, vmode_cnt_inst_N10, vmode_cnt_inst_q_0_,
         vmode_cnt_inst_q_1_, vmode_cnt_inst_q_2_, res_cnt_inst_n2,
         res_cnt_inst_n1, res_cnt_inst_n14, res_cnt_inst_n13, res_cnt_inst_n12,
         res_cnt_inst_n11, res_cnt_inst_n10, res_cnt_inst_n9, res_cnt_inst_n8,
         res_cnt_inst_n7, res_cnt_inst_n5, res_cnt_inst_net2987,
         res_cnt_inst_N12, res_cnt_inst_N10, res_cnt_inst_q_0_,
         res_cnt_inst_q_1_, res_cnt_inst_q_2_, i_data_npu_cnt_inst_n4,
         i_data_npu_cnt_inst_n2, i_data_npu_cnt_inst_n1,
         i_data_npu_cnt_inst_n19, i_data_npu_cnt_inst_n18,
         i_data_npu_cnt_inst_n17, i_data_npu_cnt_inst_n16,
         i_data_npu_cnt_inst_n15, i_data_npu_cnt_inst_n14,
         i_data_npu_cnt_inst_n13, i_data_npu_cnt_inst_n12,
         i_data_npu_cnt_inst_n11, i_data_npu_cnt_inst_n10,
         i_data_npu_cnt_inst_n9, i_data_npu_cnt_inst_n8,
         i_data_npu_cnt_inst_n5, i_data_npu_cnt_inst_net2969,
         i_data_npu_cnt_inst_N14, i_data_npu_cnt_inst_N13,
         i_data_npu_cnt_inst_N11, i_data_npu_cnt_inst_q_3_,
         i_data_L2_cnt_inst_n4, i_data_L2_cnt_inst_n2, i_data_L2_cnt_inst_n1,
         i_data_L2_cnt_inst_n19, i_data_L2_cnt_inst_n18,
         i_data_L2_cnt_inst_n17, i_data_L2_cnt_inst_n16,
         i_data_L2_cnt_inst_n15, i_data_L2_cnt_inst_n14,
         i_data_L2_cnt_inst_n13, i_data_L2_cnt_inst_n12,
         i_data_L2_cnt_inst_n11, i_data_L2_cnt_inst_n10, i_data_L2_cnt_inst_n9,
         i_data_L2_cnt_inst_n8, i_data_L2_cnt_inst_n5,
         i_data_L2_cnt_inst_net2951, i_data_L2_cnt_inst_N14,
         i_data_L2_cnt_inst_N13, i_data_L2_cnt_inst_N11,
         i_data_L2_cnt_inst_q_0_, i_data_L2_cnt_inst_q_1_,
         i_data_L2_cnt_inst_q_2_, i_data_L2_cnt_inst_q_3_,
         i_data_L3_cnt_inst_n4, i_data_L3_cnt_inst_n2, i_data_L3_cnt_inst_n1,
         i_data_L3_cnt_inst_n19, i_data_L3_cnt_inst_n18,
         i_data_L3_cnt_inst_n17, i_data_L3_cnt_inst_n16,
         i_data_L3_cnt_inst_n15, i_data_L3_cnt_inst_n14,
         i_data_L3_cnt_inst_n13, i_data_L3_cnt_inst_n12,
         i_data_L3_cnt_inst_n11, i_data_L3_cnt_inst_n10, i_data_L3_cnt_inst_n9,
         i_data_L3_cnt_inst_n8, i_data_L3_cnt_inst_n5,
         i_data_L3_cnt_inst_net2933, i_data_L3_cnt_inst_N14,
         i_data_L3_cnt_inst_N13, i_data_L3_cnt_inst_N11,
         i_data_L3_cnt_inst_q_2_, i_data_L3_cnt_inst_q_3_, L0_cnt_inst_n4,
         L0_cnt_inst_n2, L0_cnt_inst_n1, L0_cnt_inst_n19, L0_cnt_inst_n18,
         L0_cnt_inst_n17, L0_cnt_inst_n16, L0_cnt_inst_n15, L0_cnt_inst_n14,
         L0_cnt_inst_n13, L0_cnt_inst_n12, L0_cnt_inst_n11, L0_cnt_inst_n10,
         L0_cnt_inst_n9, L0_cnt_inst_n8, L0_cnt_inst_n5, L0_cnt_inst_net2915,
         L0_cnt_inst_N14, L0_cnt_inst_N13, L0_cnt_inst_N11, L0_cnt_inst_q_3_,
         L4_cnt_inst_n4, L4_cnt_inst_n2, L4_cnt_inst_n1, L4_cnt_inst_n19,
         L4_cnt_inst_n18, L4_cnt_inst_n17, L4_cnt_inst_n16, L4_cnt_inst_n15,
         L4_cnt_inst_n14, L4_cnt_inst_n13, L4_cnt_inst_n12, L4_cnt_inst_n11,
         L4_cnt_inst_n10, L4_cnt_inst_n9, L4_cnt_inst_n8, L4_cnt_inst_n5,
         L4_cnt_inst_net2897, L4_cnt_inst_N14, L4_cnt_inst_N13,
         L4_cnt_inst_N11, L4_cnt_inst_q_0_, L4_cnt_inst_q_1_, L4_cnt_inst_q_2_,
         L4_cnt_inst_q_3_, i_weight_addr_gen_inst_n26,
         i_weight_addr_gen_inst_n25, i_weight_addr_gen_inst_n24,
         i_weight_addr_gen_inst_n23, i_weight_addr_gen_inst_n22,
         i_weight_addr_gen_inst_n21, i_weight_addr_gen_inst_n20,
         i_weight_addr_gen_inst_n19, i_weight_addr_gen_inst_n17,
         i_weight_addr_gen_inst_n8, i_weight_addr_gen_inst_n7,
         i_weight_addr_gen_inst_n6, i_weight_addr_gen_inst_n5,
         i_weight_addr_gen_inst_n40, i_weight_addr_gen_inst_n39,
         i_weight_addr_gen_inst_n38, i_weight_addr_gen_inst_n37,
         i_weight_addr_gen_inst_n36, i_weight_addr_gen_inst_n35,
         i_weight_addr_gen_inst_n34, i_weight_addr_gen_inst_n33,
         i_weight_addr_gen_inst_n32, i_weight_addr_gen_inst_n31,
         i_weight_addr_gen_inst_n30, i_weight_addr_gen_inst_net2880,
         i_weight_addr_gen_inst_net2874, i_weight_addr_gen_inst_N60,
         i_weight_addr_gen_inst_N59, i_weight_addr_gen_inst_N58,
         i_weight_addr_gen_inst_N57, i_weight_addr_gen_inst_N56,
         i_weight_addr_gen_inst_N55, i_weight_addr_gen_inst_N54,
         i_weight_addr_gen_inst_N53, i_weight_addr_gen_inst_N52,
         i_weight_addr_gen_inst_N51, i_weight_addr_gen_inst_N37,
         i_weight_addr_gen_inst_N27, i_weight_addr_gen_inst_N26,
         i_weight_addr_gen_inst_N25, i_weight_addr_gen_inst_N24,
         i_weight_addr_gen_inst_N23, i_weight_addr_gen_inst_N22,
         i_weight_addr_gen_inst_N21, i_weight_addr_gen_inst_N20,
         i_weight_addr_gen_inst_N19, i_weight_addr_gen_inst_N18,
         i_weight_addr_gen_inst_N17, i_weight_addr_gen_inst_N16,
         i_weight_addr_gen_inst_N15, i_weight_addr_gen_inst_N14,
         i_weight_addr_gen_inst_N13, i_weight_addr_gen_inst_N12,
         i_weight_addr_gen_inst_N11, i_weight_addr_gen_inst_N10,
         i_weight_addr_gen_inst_int_offs_addr_0_,
         i_weight_addr_gen_inst_int_offs_addr_1_,
         i_weight_addr_gen_inst_int_offs_addr_2_,
         i_weight_addr_gen_inst_int_offs_addr_3_,
         i_weight_addr_gen_inst_int_offs_addr_4_,
         i_weight_addr_gen_inst_int_offs_addr_5_,
         i_weight_addr_gen_inst_int_offs_addr_6_,
         i_weight_addr_gen_inst_int_offs_addr_7_,
         i_weight_addr_gen_inst_int_offs_addr_8_,
         i_weight_addr_gen_inst_int_base_addr_0_,
         i_weight_addr_gen_inst_int_base_addr_1_,
         i_weight_addr_gen_inst_int_base_addr_2_,
         i_weight_addr_gen_inst_int_base_addr_3_,
         i_weight_addr_gen_inst_int_base_addr_4_,
         i_weight_addr_gen_inst_int_base_addr_5_,
         i_weight_addr_gen_inst_int_base_addr_6_,
         i_weight_addr_gen_inst_int_base_addr_7_,
         i_weight_addr_gen_inst_int_base_addr_8_,
         i_weight_addr_gen_inst_add_60_n1, i_weight_addr_gen_inst_add_45_n2,
         i_weight_addr_gen_inst_add_43_n2, i_weight_addr_gen_inst_add_31_n1,
         i_data_even_addr_gen_inst_n28, i_data_even_addr_gen_inst_n27,
         i_data_even_addr_gen_inst_n26, i_data_even_addr_gen_inst_n25,
         i_data_even_addr_gen_inst_n24, i_data_even_addr_gen_inst_n23,
         i_data_even_addr_gen_inst_n22, i_data_even_addr_gen_inst_n21,
         i_data_even_addr_gen_inst_n20, i_data_even_addr_gen_inst_n18,
         i_data_even_addr_gen_inst_n8, i_data_even_addr_gen_inst_n7,
         i_data_even_addr_gen_inst_n6, i_data_even_addr_gen_inst_n5,
         i_data_even_addr_gen_inst_n43, i_data_even_addr_gen_inst_n42,
         i_data_even_addr_gen_inst_n41, i_data_even_addr_gen_inst_n40,
         i_data_even_addr_gen_inst_n39, i_data_even_addr_gen_inst_n38,
         i_data_even_addr_gen_inst_n37, i_data_even_addr_gen_inst_n36,
         i_data_even_addr_gen_inst_n35, i_data_even_addr_gen_inst_n34,
         i_data_even_addr_gen_inst_n33, i_data_even_addr_gen_inst_n32,
         i_data_even_addr_gen_inst_net2857, i_data_even_addr_gen_inst_net2851,
         i_data_even_addr_gen_inst_N65, i_data_even_addr_gen_inst_N64,
         i_data_even_addr_gen_inst_N63, i_data_even_addr_gen_inst_N62,
         i_data_even_addr_gen_inst_N61, i_data_even_addr_gen_inst_N60,
         i_data_even_addr_gen_inst_N59, i_data_even_addr_gen_inst_N58,
         i_data_even_addr_gen_inst_N57, i_data_even_addr_gen_inst_N56,
         i_data_even_addr_gen_inst_N55, i_data_even_addr_gen_inst_N40,
         i_data_even_addr_gen_inst_N29, i_data_even_addr_gen_inst_N28,
         i_data_even_addr_gen_inst_N27, i_data_even_addr_gen_inst_N26,
         i_data_even_addr_gen_inst_N25, i_data_even_addr_gen_inst_N24,
         i_data_even_addr_gen_inst_N23, i_data_even_addr_gen_inst_N22,
         i_data_even_addr_gen_inst_N21, i_data_even_addr_gen_inst_N20,
         i_data_even_addr_gen_inst_N19, i_data_even_addr_gen_inst_N18,
         i_data_even_addr_gen_inst_N17, i_data_even_addr_gen_inst_N16,
         i_data_even_addr_gen_inst_N15, i_data_even_addr_gen_inst_N14,
         i_data_even_addr_gen_inst_N13, i_data_even_addr_gen_inst_N12,
         i_data_even_addr_gen_inst_N11, i_data_even_addr_gen_inst_N10,
         i_data_even_addr_gen_inst_int_offs_addr_0_,
         i_data_even_addr_gen_inst_int_offs_addr_1_,
         i_data_even_addr_gen_inst_int_offs_addr_2_,
         i_data_even_addr_gen_inst_int_offs_addr_3_,
         i_data_even_addr_gen_inst_int_offs_addr_4_,
         i_data_even_addr_gen_inst_int_offs_addr_5_,
         i_data_even_addr_gen_inst_int_offs_addr_6_,
         i_data_even_addr_gen_inst_int_offs_addr_7_,
         i_data_even_addr_gen_inst_int_offs_addr_8_,
         i_data_even_addr_gen_inst_int_offs_addr_9_,
         i_data_even_addr_gen_inst_int_base_addr_0_,
         i_data_even_addr_gen_inst_int_base_addr_1_,
         i_data_even_addr_gen_inst_int_base_addr_2_,
         i_data_even_addr_gen_inst_int_base_addr_3_,
         i_data_even_addr_gen_inst_int_base_addr_4_,
         i_data_even_addr_gen_inst_int_base_addr_5_,
         i_data_even_addr_gen_inst_int_base_addr_6_,
         i_data_even_addr_gen_inst_int_base_addr_7_,
         i_data_even_addr_gen_inst_int_base_addr_8_,
         i_data_even_addr_gen_inst_int_base_addr_9_,
         i_data_even_addr_gen_inst_add_60_n1,
         i_data_even_addr_gen_inst_add_45_n2,
         i_data_even_addr_gen_inst_add_43_n2,
         i_data_even_addr_gen_inst_add_31_n2, i_data_odd_addr_gen_inst_n28,
         i_data_odd_addr_gen_inst_n27, i_data_odd_addr_gen_inst_n26,
         i_data_odd_addr_gen_inst_n25, i_data_odd_addr_gen_inst_n24,
         i_data_odd_addr_gen_inst_n23, i_data_odd_addr_gen_inst_n22,
         i_data_odd_addr_gen_inst_n21, i_data_odd_addr_gen_inst_n20,
         i_data_odd_addr_gen_inst_n18, i_data_odd_addr_gen_inst_n8,
         i_data_odd_addr_gen_inst_n7, i_data_odd_addr_gen_inst_n6,
         i_data_odd_addr_gen_inst_n5, i_data_odd_addr_gen_inst_n43,
         i_data_odd_addr_gen_inst_n42, i_data_odd_addr_gen_inst_n41,
         i_data_odd_addr_gen_inst_n40, i_data_odd_addr_gen_inst_n39,
         i_data_odd_addr_gen_inst_n38, i_data_odd_addr_gen_inst_n37,
         i_data_odd_addr_gen_inst_n36, i_data_odd_addr_gen_inst_n35,
         i_data_odd_addr_gen_inst_n34, i_data_odd_addr_gen_inst_n33,
         i_data_odd_addr_gen_inst_n32, i_data_odd_addr_gen_inst_net2834,
         i_data_odd_addr_gen_inst_net2828, i_data_odd_addr_gen_inst_N65,
         i_data_odd_addr_gen_inst_N64, i_data_odd_addr_gen_inst_N63,
         i_data_odd_addr_gen_inst_N62, i_data_odd_addr_gen_inst_N61,
         i_data_odd_addr_gen_inst_N60, i_data_odd_addr_gen_inst_N59,
         i_data_odd_addr_gen_inst_N58, i_data_odd_addr_gen_inst_N57,
         i_data_odd_addr_gen_inst_N56, i_data_odd_addr_gen_inst_N55,
         i_data_odd_addr_gen_inst_N40, i_data_odd_addr_gen_inst_N29,
         i_data_odd_addr_gen_inst_N28, i_data_odd_addr_gen_inst_N27,
         i_data_odd_addr_gen_inst_N26, i_data_odd_addr_gen_inst_N25,
         i_data_odd_addr_gen_inst_N24, i_data_odd_addr_gen_inst_N23,
         i_data_odd_addr_gen_inst_N22, i_data_odd_addr_gen_inst_N21,
         i_data_odd_addr_gen_inst_N20, i_data_odd_addr_gen_inst_N19,
         i_data_odd_addr_gen_inst_N18, i_data_odd_addr_gen_inst_N17,
         i_data_odd_addr_gen_inst_N16, i_data_odd_addr_gen_inst_N15,
         i_data_odd_addr_gen_inst_N14, i_data_odd_addr_gen_inst_N13,
         i_data_odd_addr_gen_inst_N12, i_data_odd_addr_gen_inst_N11,
         i_data_odd_addr_gen_inst_N10,
         i_data_odd_addr_gen_inst_int_offs_addr_0_,
         i_data_odd_addr_gen_inst_int_offs_addr_1_,
         i_data_odd_addr_gen_inst_int_offs_addr_2_,
         i_data_odd_addr_gen_inst_int_offs_addr_3_,
         i_data_odd_addr_gen_inst_int_offs_addr_4_,
         i_data_odd_addr_gen_inst_int_offs_addr_5_,
         i_data_odd_addr_gen_inst_int_offs_addr_6_,
         i_data_odd_addr_gen_inst_int_offs_addr_7_,
         i_data_odd_addr_gen_inst_int_offs_addr_8_,
         i_data_odd_addr_gen_inst_int_offs_addr_9_,
         i_data_odd_addr_gen_inst_int_base_addr_0_,
         i_data_odd_addr_gen_inst_int_base_addr_1_,
         i_data_odd_addr_gen_inst_int_base_addr_2_,
         i_data_odd_addr_gen_inst_int_base_addr_3_,
         i_data_odd_addr_gen_inst_int_base_addr_4_,
         i_data_odd_addr_gen_inst_int_base_addr_5_,
         i_data_odd_addr_gen_inst_int_base_addr_6_,
         i_data_odd_addr_gen_inst_int_base_addr_7_,
         i_data_odd_addr_gen_inst_int_base_addr_8_,
         i_data_odd_addr_gen_inst_int_base_addr_9_,
         i_data_odd_addr_gen_inst_add_60_n1,
         i_data_odd_addr_gen_inst_add_45_n2,
         i_data_odd_addr_gen_inst_add_43_n2,
         i_data_odd_addr_gen_inst_add_31_n2, o_data_even_addr_gen_inst_n28,
         o_data_even_addr_gen_inst_n27, o_data_even_addr_gen_inst_n26,
         o_data_even_addr_gen_inst_n25, o_data_even_addr_gen_inst_n24,
         o_data_even_addr_gen_inst_n23, o_data_even_addr_gen_inst_n22,
         o_data_even_addr_gen_inst_n21, o_data_even_addr_gen_inst_n20,
         o_data_even_addr_gen_inst_n18, o_data_even_addr_gen_inst_n8,
         o_data_even_addr_gen_inst_n7, o_data_even_addr_gen_inst_n6,
         o_data_even_addr_gen_inst_n5, o_data_even_addr_gen_inst_n43,
         o_data_even_addr_gen_inst_n42, o_data_even_addr_gen_inst_n41,
         o_data_even_addr_gen_inst_n40, o_data_even_addr_gen_inst_n39,
         o_data_even_addr_gen_inst_n38, o_data_even_addr_gen_inst_n37,
         o_data_even_addr_gen_inst_n36, o_data_even_addr_gen_inst_n35,
         o_data_even_addr_gen_inst_n34, o_data_even_addr_gen_inst_n33,
         o_data_even_addr_gen_inst_n32, o_data_even_addr_gen_inst_net2811,
         o_data_even_addr_gen_inst_net2805, o_data_even_addr_gen_inst_N65,
         o_data_even_addr_gen_inst_N64, o_data_even_addr_gen_inst_N63,
         o_data_even_addr_gen_inst_N62, o_data_even_addr_gen_inst_N61,
         o_data_even_addr_gen_inst_N60, o_data_even_addr_gen_inst_N59,
         o_data_even_addr_gen_inst_N58, o_data_even_addr_gen_inst_N57,
         o_data_even_addr_gen_inst_N56, o_data_even_addr_gen_inst_N55,
         o_data_even_addr_gen_inst_N40, o_data_even_addr_gen_inst_N29,
         o_data_even_addr_gen_inst_N28, o_data_even_addr_gen_inst_N27,
         o_data_even_addr_gen_inst_N26, o_data_even_addr_gen_inst_N25,
         o_data_even_addr_gen_inst_N24, o_data_even_addr_gen_inst_N23,
         o_data_even_addr_gen_inst_N22, o_data_even_addr_gen_inst_N21,
         o_data_even_addr_gen_inst_N20, o_data_even_addr_gen_inst_N19,
         o_data_even_addr_gen_inst_N18, o_data_even_addr_gen_inst_N17,
         o_data_even_addr_gen_inst_N16, o_data_even_addr_gen_inst_N15,
         o_data_even_addr_gen_inst_N14, o_data_even_addr_gen_inst_N13,
         o_data_even_addr_gen_inst_N12, o_data_even_addr_gen_inst_N11,
         o_data_even_addr_gen_inst_N10,
         o_data_even_addr_gen_inst_int_offs_addr_0_,
         o_data_even_addr_gen_inst_int_offs_addr_1_,
         o_data_even_addr_gen_inst_int_offs_addr_2_,
         o_data_even_addr_gen_inst_int_offs_addr_3_,
         o_data_even_addr_gen_inst_int_offs_addr_4_,
         o_data_even_addr_gen_inst_int_offs_addr_5_,
         o_data_even_addr_gen_inst_int_offs_addr_6_,
         o_data_even_addr_gen_inst_int_offs_addr_7_,
         o_data_even_addr_gen_inst_int_offs_addr_8_,
         o_data_even_addr_gen_inst_int_offs_addr_9_,
         o_data_even_addr_gen_inst_int_base_addr_0_,
         o_data_even_addr_gen_inst_int_base_addr_1_,
         o_data_even_addr_gen_inst_int_base_addr_2_,
         o_data_even_addr_gen_inst_int_base_addr_3_,
         o_data_even_addr_gen_inst_int_base_addr_4_,
         o_data_even_addr_gen_inst_int_base_addr_5_,
         o_data_even_addr_gen_inst_int_base_addr_6_,
         o_data_even_addr_gen_inst_int_base_addr_7_,
         o_data_even_addr_gen_inst_int_base_addr_8_,
         o_data_even_addr_gen_inst_int_base_addr_9_,
         o_data_even_addr_gen_inst_add_60_n1,
         o_data_even_addr_gen_inst_add_45_n2,
         o_data_even_addr_gen_inst_add_43_n2,
         o_data_even_addr_gen_inst_add_31_n1, o_data_odd_addr_gen_inst_n28,
         o_data_odd_addr_gen_inst_n27, o_data_odd_addr_gen_inst_n26,
         o_data_odd_addr_gen_inst_n25, o_data_odd_addr_gen_inst_n24,
         o_data_odd_addr_gen_inst_n23, o_data_odd_addr_gen_inst_n22,
         o_data_odd_addr_gen_inst_n21, o_data_odd_addr_gen_inst_n20,
         o_data_odd_addr_gen_inst_n18, o_data_odd_addr_gen_inst_n8,
         o_data_odd_addr_gen_inst_n7, o_data_odd_addr_gen_inst_n6,
         o_data_odd_addr_gen_inst_n5, o_data_odd_addr_gen_inst_n43,
         o_data_odd_addr_gen_inst_n42, o_data_odd_addr_gen_inst_n41,
         o_data_odd_addr_gen_inst_n40, o_data_odd_addr_gen_inst_n39,
         o_data_odd_addr_gen_inst_n38, o_data_odd_addr_gen_inst_n37,
         o_data_odd_addr_gen_inst_n36, o_data_odd_addr_gen_inst_n35,
         o_data_odd_addr_gen_inst_n34, o_data_odd_addr_gen_inst_n33,
         o_data_odd_addr_gen_inst_n32, o_data_odd_addr_gen_inst_net2788,
         o_data_odd_addr_gen_inst_net2782, o_data_odd_addr_gen_inst_N65,
         o_data_odd_addr_gen_inst_N64, o_data_odd_addr_gen_inst_N63,
         o_data_odd_addr_gen_inst_N62, o_data_odd_addr_gen_inst_N61,
         o_data_odd_addr_gen_inst_N60, o_data_odd_addr_gen_inst_N59,
         o_data_odd_addr_gen_inst_N58, o_data_odd_addr_gen_inst_N57,
         o_data_odd_addr_gen_inst_N56, o_data_odd_addr_gen_inst_N55,
         o_data_odd_addr_gen_inst_N40, o_data_odd_addr_gen_inst_N29,
         o_data_odd_addr_gen_inst_N28, o_data_odd_addr_gen_inst_N27,
         o_data_odd_addr_gen_inst_N26, o_data_odd_addr_gen_inst_N25,
         o_data_odd_addr_gen_inst_N24, o_data_odd_addr_gen_inst_N23,
         o_data_odd_addr_gen_inst_N22, o_data_odd_addr_gen_inst_N21,
         o_data_odd_addr_gen_inst_N20, o_data_odd_addr_gen_inst_N19,
         o_data_odd_addr_gen_inst_N18, o_data_odd_addr_gen_inst_N17,
         o_data_odd_addr_gen_inst_N16, o_data_odd_addr_gen_inst_N15,
         o_data_odd_addr_gen_inst_N14, o_data_odd_addr_gen_inst_N13,
         o_data_odd_addr_gen_inst_N12, o_data_odd_addr_gen_inst_N11,
         o_data_odd_addr_gen_inst_N10,
         o_data_odd_addr_gen_inst_int_offs_addr_0_,
         o_data_odd_addr_gen_inst_int_offs_addr_1_,
         o_data_odd_addr_gen_inst_int_offs_addr_2_,
         o_data_odd_addr_gen_inst_int_offs_addr_3_,
         o_data_odd_addr_gen_inst_int_offs_addr_4_,
         o_data_odd_addr_gen_inst_int_offs_addr_5_,
         o_data_odd_addr_gen_inst_int_offs_addr_6_,
         o_data_odd_addr_gen_inst_int_offs_addr_7_,
         o_data_odd_addr_gen_inst_int_offs_addr_8_,
         o_data_odd_addr_gen_inst_int_offs_addr_9_,
         o_data_odd_addr_gen_inst_int_base_addr_0_,
         o_data_odd_addr_gen_inst_int_base_addr_1_,
         o_data_odd_addr_gen_inst_int_base_addr_2_,
         o_data_odd_addr_gen_inst_int_base_addr_3_,
         o_data_odd_addr_gen_inst_int_base_addr_4_,
         o_data_odd_addr_gen_inst_int_base_addr_5_,
         o_data_odd_addr_gen_inst_int_base_addr_6_,
         o_data_odd_addr_gen_inst_int_base_addr_7_,
         o_data_odd_addr_gen_inst_int_base_addr_8_,
         o_data_odd_addr_gen_inst_int_base_addr_9_,
         o_data_odd_addr_gen_inst_add_60_n1,
         o_data_odd_addr_gen_inst_add_45_n2,
         o_data_odd_addr_gen_inst_add_43_n2,
         o_data_odd_addr_gen_inst_add_31_n1;
  wire   [2:0] ps_int_hmode_cnt;
  wire   [15:0] int_i_data_h_npu;
  wire   [15:0] int_i_data_v_npu;
  wire   [2:0] ps_int_L0_ptr;
  wire   [2:0] int_L0_ptr;
  wire   [2:0] int_L1_ptr;
  wire   [2:0] int_hmode_cnt;
  wire   [1:7] int_ckg_rmask;
  wire   [1:7] int_ckg_cmask;
  wire   [63:0] int_o_data_npu;
  wire   [15:0] int_o_data_p;
  wire   [2:0] int_arv_res;
  wire   [2:0] int_d_tc;
  wire   [4:0] int_c_o_inc_value_offs;
  wire   [3:2] add_538_carry;
  wire   [7:0] wrap_act_buffer_inst_int_i_data_if8;
  wire   [7:0] wrap_act_buffer_inst_int_i_data_if7;
  wire   [7:0] wrap_act_buffer_inst_int_i_data_if6;
  wire   [7:0] wrap_act_buffer_inst_int_i_data_if5;
  wire   [7:0] wrap_act_buffer_inst_int_i_data_if4;
  wire   [7:0] wrap_act_buffer_inst_int_i_data_if3;
  wire   [7:0] wrap_act_buffer_inst_int_i_data_if2;
  wire   [7:0] wrap_act_buffer_inst_int_i_data_if1;
  wire   [47:0] wrap_act_buffer_inst_act_buffer_inst_int_data8;
  wire   [47:0] wrap_act_buffer_inst_act_buffer_inst_int_data7;
  wire   [47:0] wrap_act_buffer_inst_act_buffer_inst_int_data6;
  wire   [47:0] wrap_act_buffer_inst_act_buffer_inst_int_data5;
  wire   [47:0] wrap_act_buffer_inst_act_buffer_inst_int_data4;
  wire   [47:0] wrap_act_buffer_inst_act_buffer_inst_int_data3;
  wire   [47:0] wrap_act_buffer_inst_act_buffer_inst_int_data2;
  wire   [47:0] wrap_act_buffer_inst_act_buffer_inst_int_data1;
  wire   [7:0] wrap_act_buffer_inst_act_if_inst_int_data8;
  wire   [7:0] wrap_act_buffer_inst_act_if_inst_int_data7;
  wire   [7:0] wrap_act_buffer_inst_act_if_inst_int_data6;
  wire   [7:0] wrap_act_buffer_inst_act_if_inst_int_data5;
  wire   [7:0] wrap_act_buffer_inst_act_if_inst_int_data4;
  wire   [7:0] wrap_act_buffer_inst_act_if_inst_int_data3;
  wire   [7:0] wrap_act_buffer_inst_act_if_inst_int_data2;
  wire   [7:0] wrap_act_buffer_inst_act_if_inst_int_data1;
  wire   [63:0] npu_inst_int_ckg;
  wire   [8:2] i_weight_addr_gen_inst_add_60_carry;
  wire   [8:2] i_weight_addr_gen_inst_add_45_carry;
  wire   [8:2] i_weight_addr_gen_inst_add_43_carry;
  wire   [8:2] i_weight_addr_gen_inst_add_31_carry;
  wire   [9:2] i_data_even_addr_gen_inst_add_60_carry;
  wire   [9:2] i_data_even_addr_gen_inst_add_45_carry;
  wire   [9:2] i_data_even_addr_gen_inst_add_43_carry;
  wire   [9:2] i_data_even_addr_gen_inst_add_31_carry;
  wire   [9:2] i_data_odd_addr_gen_inst_add_60_carry;
  wire   [9:2] i_data_odd_addr_gen_inst_add_45_carry;
  wire   [9:2] i_data_odd_addr_gen_inst_add_43_carry;
  wire   [9:2] i_data_odd_addr_gen_inst_add_31_carry;
  wire   [9:2] o_data_even_addr_gen_inst_add_60_carry;
  wire   [9:2] o_data_even_addr_gen_inst_add_45_carry;
  wire   [9:2] o_data_even_addr_gen_inst_add_43_carry;
  wire   [9:2] o_data_even_addr_gen_inst_add_31_carry;
  wire   [9:2] o_data_odd_addr_gen_inst_add_60_carry;
  wire   [9:2] o_data_odd_addr_gen_inst_add_45_carry;
  wire   [9:2] o_data_odd_addr_gen_inst_add_43_carry;
  wire   [9:2] o_data_odd_addr_gen_inst_add_31_carry;

  DFFR_X1 ps_ctrl_wr_mem_reg ( .D(ctrl_wr_mem), .CK(ck), .RN(n31), .Q(
        o_data_wr), .QN(n4) );
  DFFR_X1 int_q_tc_reg_2_ ( .D(int_d_tc[2]), .CK(net2764), .RN(n31), .Q(
        s_tc_L2), .QN(n7) );
  DFFR_X1 int_q_tc_reg_1_ ( .D(int_d_tc[1]), .CK(net2764), .RN(n31), .Q(
        s_tc_L3), .QN(n9) );
  DFFR_X1 int_q_tc_reg_0_ ( .D(int_d_tc[0]), .CK(net2764), .RN(n31), .Q(
        s_tc_L4) );
  DFFR_X1 ps_int_s_tc_res_reg ( .D(s_tc_res), .CK(ck), .RN(n32), .Q(
        ps_int_s_tc_res) );
  NAND3_X1 U54 ( .A1(n41), .A2(n37), .A3(n42), .ZN(n26) );
  HA_X1 add_538_U1_1_1 ( .A(arv_L4[1]), .B(arv_L4[0]), .CO(add_538_carry[2]), 
        .S(int_c_o_inc_value_offs[1]) );
  HA_X1 add_538_U1_1_2 ( .A(arv_L4[2]), .B(add_538_carry[2]), .CO(
        add_538_carry[3]), .S(int_c_o_inc_value_offs[2]) );
  HA_X1 add_538_U1_1_3 ( .A(arv_L4[3]), .B(add_538_carry[3]), .CO(
        int_c_o_inc_value_offs[4]), .S(int_c_o_inc_value_offs[3]) );
  DFFR_X1 ps_int_hmode_cnt_reg_1_ ( .D(int_hmode_cnt[1]), .CK(ck), .RN(n32), 
        .Q(ps_int_hmode_cnt[1]) );
  DFFR_X1 ps_int_hmode_cnt_reg_2_ ( .D(int_hmode_cnt[2]), .CK(ck), .RN(n31), 
        .Q(ps_int_hmode_cnt[2]) );
  DFFR_X1 ps_int_L0_ptr_reg_1_ ( .D(int_L0_ptr[1]), .CK(ck), .RN(n32), .Q(
        ps_int_L0_ptr[1]) );
  DFFR_X1 ps_int_s_tc_L3_reg ( .D(s_tc_L3), .CK(ck), .RN(n31), .Q(
        ps_int_s_tc_L3) );
  DFFR_X1 ps_int_hmode_cnt_reg_0_ ( .D(int_hmode_cnt[0]), .CK(ck), .RN(n32), 
        .Q(ps_int_hmode_cnt[0]) );
  DFFR_X1 ps_int_L0_ptr_reg_2_ ( .D(int_L0_ptr[2]), .CK(ck), .RN(n32), .Q(
        ps_int_L0_ptr[2]) );
  DFFR_X1 ps_int_s_tc_L2_reg ( .D(s_tc_L2), .CK(ck), .RN(n32), .Q(
        ps_int_s_tc_L2) );
  DFFR_X1 ps_int_L0_ptr_reg_0_ ( .D(int_L0_ptr[0]), .CK(ck), .RN(n32), .Q(
        ps_int_L0_ptr[0]) );
  DFFR_X1 int_o_data_wrh_l_n_reg ( .D(n30), .CK(ck), .RN(n32), .Q(
        o_data_wrh_l_n) );
  DFFR_X1 int_o_data_ev_odd_n_reg ( .D(n35), .CK(ck), .RN(n32), .Q(
        o_data_ev_odd_n) );
  DFFR_X1 ps_ctrl_en_p_reg ( .D(ctrl_en_p), .CK(ck), .RN(n32), .Q(ps_ctrl_en_p) );
  DFFR_X1 ps_ctrl_wr_pipe_reg ( .D(ctrl_wr_pipe), .CK(ck), .RN(n32), .Q(
        ps_ctrl_wr_pipe) );
  DFFR_X1 ps_ctrl_en_npu_reg ( .D(ctrl_en_npu), .CK(ck), .RN(n32), .Q(
        ps_ctrl_en_npu) );
  DFFR_X1 ps_ctrl_ldh_v_n_reg ( .D(ctrl_ldh_v_n), .CK(ck), .RN(n32), .Q(
        ps_ctrl_ldh_v_n) );
  INV_X1 U55 ( .A(n29), .ZN(n33) );
  AND2_X1 U56 ( .A1(int_d_tc[1]), .A2(n33), .ZN(int_en_L4_ptr) );
  NOR3_X1 U57 ( .A1(n42), .A2(n41), .A3(n24), .ZN(n22) );
  INV_X1 U58 ( .A(n27), .ZN(n39) );
  NOR2_X1 U59 ( .A1(n34), .A2(n29), .ZN(int_c_i_en_odd) );
  NAND2_X1 U60 ( .A1(n23), .A2(int_arv_res[1]), .ZN(int_ckg_rmask[6]) );
  INV_X1 U61 ( .A(n23), .ZN(n40) );
  AOI21_X1 U62 ( .B1(n37), .B2(n42), .A(n28), .ZN(n25) );
  NAND2_X1 U63 ( .A1(int_d_tc[2]), .A2(int_en_L2_ptr), .ZN(n29) );
  INV_X1 U64 ( .A(s_tc_res), .ZN(n36) );
  INV_X1 U65 ( .A(n28), .ZN(n38) );
  AND2_X1 U66 ( .A1(s_tc_L1), .A2(int_en_L1_ptr), .ZN(int_en_L2_ptr) );
  INV_X1 U67 ( .A(n19), .ZN(n43) );
  NOR3_X1 U68 ( .A1(n36), .A2(n7), .A3(n9), .ZN(int_c_i_en_weight_addr) );
  OAI21_X1 U69 ( .B1(arv_CKG[1]), .B2(n9), .A(n27), .ZN(int_ckg_cmask[6]) );
  NOR2_X1 U70 ( .A1(n22), .A2(n9), .ZN(int_ckg_cmask[7]) );
  NOR2_X1 U71 ( .A1(n25), .A2(n9), .ZN(int_ckg_cmask[3]) );
  NOR2_X1 U72 ( .A1(n38), .A2(n9), .ZN(int_ckg_cmask[2]) );
  NOR2_X1 U73 ( .A1(n26), .A2(n9), .ZN(int_ckg_cmask[1]) );
  NOR2_X1 U74 ( .A1(i_data_ev_odd_n), .A2(n29), .ZN(int_c_i_en_even) );
  OAI21_X1 U75 ( .B1(arv_CKG[1]), .B2(arv_CKG[0]), .A(arv_CKG[2]), .ZN(n24) );
  NOR2_X1 U76 ( .A1(n22), .A2(n7), .ZN(int_ckg_rmask[7]) );
  NOR2_X1 U77 ( .A1(n25), .A2(n7), .ZN(int_ckg_rmask[3]) );
  NOR2_X1 U78 ( .A1(n7), .A2(n38), .ZN(int_ckg_rmask[2]) );
  NOR2_X1 U79 ( .A1(n7), .A2(n26), .ZN(int_ckg_rmask[1]) );
  NOR2_X1 U80 ( .A1(arv_CKG[1]), .A2(arv_CKG[2]), .ZN(n28) );
  INV_X1 U81 ( .A(arv_L4[0]), .ZN(int_c_o_inc_value_offs[0]) );
  NAND2_X1 U82 ( .A1(s_tc_L2), .A2(n41), .ZN(int_arv_res[1]) );
  INV_X1 U83 ( .A(arv_CKG[0]), .ZN(n42) );
  NAND2_X1 U84 ( .A1(s_tc_L2), .A2(n24), .ZN(n23) );
  NAND2_X1 U85 ( .A1(s_tc_L2), .A2(n42), .ZN(int_arv_res[0]) );
  NAND2_X1 U86 ( .A1(s_tc_L2), .A2(n37), .ZN(int_arv_res[2]) );
  NAND2_X1 U87 ( .A1(s_tc_L3), .A2(n24), .ZN(n27) );
  INV_X1 U88 ( .A(arv_CKG[1]), .ZN(n41) );
  INV_X1 U89 ( .A(arv_CKG[2]), .ZN(n37) );
  AND2_X1 U90 ( .A1(ctrl_ldh_v_n), .A2(s_tc_L0), .ZN(int_en_L1_ptr) );
  NOR2_X1 U91 ( .A1(arv_CKG[2]), .A2(n9), .ZN(int_ckg_cmask[4]) );
  NOR2_X1 U92 ( .A1(arv_CKG[2]), .A2(n7), .ZN(int_ckg_rmask[4]) );
  AND2_X1 U93 ( .A1(ps_int_s_tc_L3), .A2(n43), .ZN(int_c_o_en_base_odd) );
  NAND2_X1 U94 ( .A1(ps_int_s_tc_res), .A2(ps_int_s_tc_L2), .ZN(n19) );
  INV_X1 U95 ( .A(i_data_ev_odd_n), .ZN(n34) );
  OAI21_X1 U96 ( .B1(n19), .B2(n34), .A(n20), .ZN(n30) );
  NAND2_X1 U97 ( .A1(o_data_wrh_l_n), .A2(n19), .ZN(n20) );
  NOR2_X1 U98 ( .A1(o_data_ev_odd_n), .A2(n4), .ZN(int_c_o_en_offs_even) );
  AND2_X1 U99 ( .A1(o_data_ev_odd_n), .A2(o_data_wr), .ZN(int_c_o_en_offs_odd)
         );
  NAND2_X1 U100 ( .A1(n36), .A2(n21), .ZN(int_en_vmode) );
  NAND2_X1 U101 ( .A1(s_tc_L0), .A2(ctrl_en_vmode), .ZN(n21) );
  INV_X1 U102 ( .A(n18), .ZN(n35) );
  AOI22_X1 U103 ( .A1(n43), .A2(int_L3_ptr_1_), .B1(n19), .B2(o_data_ev_odd_n), 
        .ZN(n18) );
  AND2_X1 U104 ( .A1(ctrl_en_hmode), .A2(s_tc_L0), .ZN(int_en_hmode) );
  INV_X1 U105 ( .A(rst), .ZN(n31) );
  INV_X1 U106 ( .A(rst), .ZN(n32) );
  INV_X1 wrap_act_buffer_inst_U2 ( .A(rst), .ZN(wrap_act_buffer_inst_n1) );
  DFFR_X1 wrap_act_buffer_inst_int_i_data_v_npu_reg_0_ ( .D(i_actv[0]), .CK(
        wrap_act_buffer_inst_net4585), .RN(wrap_act_buffer_inst_n1), .Q(
        int_i_data_v_npu[0]) );
  DFFR_X1 wrap_act_buffer_inst_int_i_data_v_npu_reg_1_ ( .D(i_actv[1]), .CK(
        wrap_act_buffer_inst_net4585), .RN(wrap_act_buffer_inst_n1), .Q(
        int_i_data_v_npu[1]) );
  DFFR_X1 wrap_act_buffer_inst_int_i_data_v_npu_reg_2_ ( .D(i_actv[2]), .CK(
        wrap_act_buffer_inst_net4585), .RN(wrap_act_buffer_inst_n1), .Q(
        int_i_data_v_npu[2]) );
  DFFR_X1 wrap_act_buffer_inst_int_i_data_v_npu_reg_3_ ( .D(i_actv[3]), .CK(
        wrap_act_buffer_inst_net4585), .RN(wrap_act_buffer_inst_n1), .Q(
        int_i_data_v_npu[3]) );
  DFFR_X1 wrap_act_buffer_inst_int_i_data_v_npu_reg_4_ ( .D(i_actv[4]), .CK(
        wrap_act_buffer_inst_net4585), .RN(wrap_act_buffer_inst_n1), .Q(
        int_i_data_v_npu[4]) );
  DFFR_X1 wrap_act_buffer_inst_int_i_data_v_npu_reg_5_ ( .D(i_actv[5]), .CK(
        wrap_act_buffer_inst_net4585), .RN(wrap_act_buffer_inst_n1), .Q(
        int_i_data_v_npu[5]) );
  DFFR_X1 wrap_act_buffer_inst_int_i_data_v_npu_reg_6_ ( .D(i_actv[6]), .CK(
        wrap_act_buffer_inst_net4585), .RN(wrap_act_buffer_inst_n1), .Q(
        int_i_data_v_npu[6]) );
  DFFR_X1 wrap_act_buffer_inst_int_i_data_v_npu_reg_7_ ( .D(i_actv[7]), .CK(
        wrap_act_buffer_inst_net4585), .RN(wrap_act_buffer_inst_n1), .Q(
        int_i_data_v_npu[7]) );
  DFFR_X1 wrap_act_buffer_inst_int_i_data_v_npu_reg_8_ ( .D(i_actv[8]), .CK(
        wrap_act_buffer_inst_net4585), .RN(wrap_act_buffer_inst_n1), .Q(
        int_i_data_v_npu[8]) );
  DFFR_X1 wrap_act_buffer_inst_int_i_data_v_npu_reg_9_ ( .D(i_actv[9]), .CK(
        wrap_act_buffer_inst_net4585), .RN(wrap_act_buffer_inst_n1), .Q(
        int_i_data_v_npu[9]) );
  DFFR_X1 wrap_act_buffer_inst_int_i_data_v_npu_reg_10_ ( .D(i_actv[10]), .CK(
        wrap_act_buffer_inst_net4585), .RN(wrap_act_buffer_inst_n1), .Q(
        int_i_data_v_npu[10]) );
  DFFR_X1 wrap_act_buffer_inst_int_i_data_v_npu_reg_11_ ( .D(i_actv[11]), .CK(
        wrap_act_buffer_inst_net4585), .RN(wrap_act_buffer_inst_n1), .Q(
        int_i_data_v_npu[11]) );
  DFFR_X1 wrap_act_buffer_inst_int_i_data_v_npu_reg_12_ ( .D(i_actv[12]), .CK(
        wrap_act_buffer_inst_net4585), .RN(wrap_act_buffer_inst_n1), .Q(
        int_i_data_v_npu[12]) );
  DFFR_X1 wrap_act_buffer_inst_int_i_data_v_npu_reg_13_ ( .D(i_actv[13]), .CK(
        wrap_act_buffer_inst_net4585), .RN(wrap_act_buffer_inst_n1), .Q(
        int_i_data_v_npu[13]) );
  DFFR_X1 wrap_act_buffer_inst_int_i_data_v_npu_reg_14_ ( .D(i_actv[14]), .CK(
        wrap_act_buffer_inst_net4585), .RN(wrap_act_buffer_inst_n1), .Q(
        int_i_data_v_npu[14]) );
  DFFR_X1 wrap_act_buffer_inst_int_i_data_v_npu_reg_15_ ( .D(i_actv[15]), .CK(
        wrap_act_buffer_inst_net4585), .RN(wrap_act_buffer_inst_n1), .Q(
        int_i_data_v_npu[15]) );
  INV_X1 wrap_act_buffer_inst_act_buffer_inst_U309 ( .A(ps_int_L0_ptr[0]), 
        .ZN(wrap_act_buffer_inst_act_buffer_inst_n192) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U308 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n12), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n188) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U307 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n13), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n182) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U306 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n14), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n176) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U305 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n15), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n170) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U304 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n16), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n164) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U303 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n17), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n9) );
  INV_X1 wrap_act_buffer_inst_act_buffer_inst_U302 ( .A(int_L1_ptr[2]), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n191) );
  INV_X1 wrap_act_buffer_inst_act_buffer_inst_U301 ( .A(int_L1_ptr[1]), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n190) );
  INV_X1 wrap_act_buffer_inst_act_buffer_inst_U300 ( .A(int_L1_ptr[0]), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n189) );
  INV_X1 wrap_act_buffer_inst_act_buffer_inst_U299 ( .A(int_L0_ptr[0]), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n194) );
  INV_X1 wrap_act_buffer_inst_act_buffer_inst_U298 ( .A(int_L0_ptr[2]), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n196) );
  INV_X1 wrap_act_buffer_inst_act_buffer_inst_U297 ( .A(int_L0_ptr[1]), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n195) );
  NAND4_X1 wrap_act_buffer_inst_act_buffer_inst_U296 ( .A1(ctrl_ldh_v_n), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n194), .A3(
        wrap_act_buffer_inst_act_buffer_inst_n195), .A4(
        wrap_act_buffer_inst_act_buffer_inst_n196), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n145) );
  NAND4_X1 wrap_act_buffer_inst_act_buffer_inst_U295 ( .A1(int_L0_ptr[1]), 
        .A2(ctrl_ldh_v_n), .A3(wrap_act_buffer_inst_act_buffer_inst_n194), 
        .A4(wrap_act_buffer_inst_act_buffer_inst_n196), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n147) );
  NAND4_X1 wrap_act_buffer_inst_act_buffer_inst_U294 ( .A1(int_L0_ptr[2]), 
        .A2(ctrl_ldh_v_n), .A3(wrap_act_buffer_inst_act_buffer_inst_n194), 
        .A4(wrap_act_buffer_inst_act_buffer_inst_n195), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n149) );
  NAND4_X1 wrap_act_buffer_inst_act_buffer_inst_U293 ( .A1(int_L0_ptr[2]), 
        .A2(int_L0_ptr[0]), .A3(ctrl_ldh_v_n), .A4(
        wrap_act_buffer_inst_act_buffer_inst_n195), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n150) );
  NAND4_X1 wrap_act_buffer_inst_act_buffer_inst_U292 ( .A1(int_L0_ptr[1]), 
        .A2(int_L0_ptr[0]), .A3(ctrl_ldh_v_n), .A4(
        wrap_act_buffer_inst_act_buffer_inst_n196), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n148) );
  NAND4_X1 wrap_act_buffer_inst_act_buffer_inst_U291 ( .A1(int_L0_ptr[0]), 
        .A2(ctrl_ldh_v_n), .A3(wrap_act_buffer_inst_act_buffer_inst_n195), 
        .A4(wrap_act_buffer_inst_act_buffer_inst_n196), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n146) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U290 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[43]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n165), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[27]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n159), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[35]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n4), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n136) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U289 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[19]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n183), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[3]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n177), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[11]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n171), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n137) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U288 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n136), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n137), .ZN(
        wrap_act_buffer_inst_int_i_data_if1[3]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U287 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[43]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n165), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[27]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n159), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[35]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n4), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n120) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U286 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[19]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n183), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[3]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n177), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[11]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n171), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n121) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U285 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n120), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n121), .ZN(
        wrap_act_buffer_inst_int_i_data_if2[3]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U284 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[19]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n185), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[3]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n179), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[11]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n173), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n73) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U283 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[43]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n167), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[27]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n161), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[35]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n6), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n72) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U282 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n72), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n73), .ZN(
        wrap_act_buffer_inst_int_i_data_if5[3]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U281 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[19]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n184), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[3]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n178), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[11]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n172), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n105) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U280 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[43]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n166), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[27]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n160), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[35]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n5), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n104) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U279 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n104), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n105), .ZN(
        wrap_act_buffer_inst_int_i_data_if3[3]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U278 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[19]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n185), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[3]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n179), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[11]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n173), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n89) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U277 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[43]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n167), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[27]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n161), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[35]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n6), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n88) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U276 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n88), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n89), .ZN(
        wrap_act_buffer_inst_int_i_data_if4[3]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U275 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[21]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n183), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[5]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n177), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[13]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n171), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n133) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U274 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[45]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n165), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[29]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n159), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[37]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n4), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n132) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U273 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n132), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n133), .ZN(
        wrap_act_buffer_inst_int_i_data_if1[5]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U272 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[21]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n184), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[5]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n178), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[13]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n172), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n117) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U264 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[45]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n166), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[29]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n160), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[37]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n5), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n116) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U263 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n116), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n117), .ZN(
        wrap_act_buffer_inst_int_i_data_if2[5]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U262 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[21]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n184), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[5]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n178), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[13]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n172), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n101) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U261 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[45]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n166), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[29]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n160), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[37]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n5), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n100) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U260 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n100), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n101), .ZN(
        wrap_act_buffer_inst_int_i_data_if3[5]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U259 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[21]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n185), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[5]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n179), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[13]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n173), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n85) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U258 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[45]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n167), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[29]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n161), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[37]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n6), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n84) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U257 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n84), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n85), .ZN(
        wrap_act_buffer_inst_int_i_data_if4[5]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U256 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[47]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n165), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[31]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n159), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[39]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n4), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n128) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U255 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[23]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n183), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[7]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n177), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[15]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n171), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n129) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U254 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n128), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n129), .ZN(
        wrap_act_buffer_inst_int_i_data_if1[7]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U253 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[23]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n184), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[7]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n178), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[15]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n172), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n113) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U252 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[47]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n166), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[31]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n160), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[39]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n5), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n112) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U251 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n112), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n113), .ZN(
        wrap_act_buffer_inst_int_i_data_if2[7]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U250 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[23]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n184), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[7]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n178), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[15]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n172), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n97) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U249 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[47]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n166), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[31]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n160), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[39]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n5), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n96) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U248 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n96), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n97), .ZN(
        wrap_act_buffer_inst_int_i_data_if3[7]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U247 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[23]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n185), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[7]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n179), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[15]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n173), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n81) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U246 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[47]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n167), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[31]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n161), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[39]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n6), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n80) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U245 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n80), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n81), .ZN(
        wrap_act_buffer_inst_int_i_data_if4[7]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U244 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[41]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n165), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[25]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n159), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[33]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n4), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n140) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U243 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[17]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n183), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[1]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n177), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[9]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n171), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n141) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U242 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n140), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n141), .ZN(
        wrap_act_buffer_inst_int_i_data_if1[1]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U241 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[41]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n165), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[25]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n159), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[33]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n4), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n124) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U240 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[17]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n183), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[1]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n177), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[9]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n171), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n125) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U239 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n124), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n125), .ZN(
        wrap_act_buffer_inst_int_i_data_if2[1]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U238 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[17]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n185), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[1]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n179), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[9]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n173), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n77) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U237 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[41]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n167), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[25]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n161), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[33]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n6), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n76) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U236 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n76), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n77), .ZN(
        wrap_act_buffer_inst_int_i_data_if5[1]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U235 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[17]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n184), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[1]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n178), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[9]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n172), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n109) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U234 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[41]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n166), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[25]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n160), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[33]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n5), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n108) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U233 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n108), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n109), .ZN(
        wrap_act_buffer_inst_int_i_data_if3[1]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U232 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[17]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n185), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[1]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n179), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[9]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n173), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n93) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U231 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[41]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n167), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[25]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n161), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[33]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n6), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n92) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U230 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n92), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n93), .ZN(
        wrap_act_buffer_inst_int_i_data_if4[1]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U229 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[42]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n165), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[26]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n159), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[34]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n4), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n138) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U228 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[18]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n183), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[2]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n177), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[10]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n171), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n139) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U227 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n138), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n139), .ZN(
        wrap_act_buffer_inst_int_i_data_if1[2]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U226 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[42]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n165), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[26]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n159), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[34]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n4), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n122) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U225 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[18]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n183), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[2]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n177), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[10]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n171), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n123) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U224 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n122), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n123), .ZN(
        wrap_act_buffer_inst_int_i_data_if2[2]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U223 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[18]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n185), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[2]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n179), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[10]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n173), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n75) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U222 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[42]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n167), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[26]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n161), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[34]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n6), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n74) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U221 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n74), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n75), .ZN(
        wrap_act_buffer_inst_int_i_data_if5[2]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U220 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[18]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n184), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[2]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n178), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[10]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n172), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n107) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U219 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[42]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n166), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[26]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n160), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[34]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n5), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n106) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U218 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n106), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n107), .ZN(
        wrap_act_buffer_inst_int_i_data_if3[2]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U217 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[18]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n185), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[2]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n179), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[10]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n173), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n91) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U216 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[42]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n167), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[26]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n161), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[34]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n6), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n90) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U215 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n90), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n91), .ZN(
        wrap_act_buffer_inst_int_i_data_if4[2]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U214 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[20]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n183), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[4]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n177), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[12]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n171), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n135) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U213 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[44]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n165), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[28]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n159), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[36]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n4), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n134) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U212 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n134), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n135), .ZN(
        wrap_act_buffer_inst_int_i_data_if1[4]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U211 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[20]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n184), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[4]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n178), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[12]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n172), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n119) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U210 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[44]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n166), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[28]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n160), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[36]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n5), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n118) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U209 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n118), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n119), .ZN(
        wrap_act_buffer_inst_int_i_data_if2[4]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U208 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[20]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n184), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[4]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n178), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[12]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n172), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n103) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U207 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[44]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n166), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[28]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n160), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[36]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n5), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n102) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U206 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n102), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n103), .ZN(
        wrap_act_buffer_inst_int_i_data_if3[4]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U205 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[20]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n185), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[4]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n179), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[12]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n173), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n87) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U204 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[44]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n167), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[28]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n161), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[36]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n6), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n86) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U203 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n86), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n87), .ZN(
        wrap_act_buffer_inst_int_i_data_if4[4]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U202 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[46]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n165), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[30]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n159), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[38]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n4), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n130) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U201 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[22]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n183), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[6]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n177), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[14]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n171), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n131) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U200 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n130), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n131), .ZN(
        wrap_act_buffer_inst_int_i_data_if1[6]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U199 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[22]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n184), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[6]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n178), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[14]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n172), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n115) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U198 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[46]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n166), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[30]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n160), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[38]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n5), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n114) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U197 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n114), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n115), .ZN(
        wrap_act_buffer_inst_int_i_data_if2[6]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U196 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[22]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n184), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[6]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n178), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[14]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n172), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n99) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U195 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[46]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n166), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[30]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n160), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[38]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n5), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n98) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U194 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n98), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n99), .ZN(
        wrap_act_buffer_inst_int_i_data_if3[6]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U193 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[22]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n185), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[6]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n179), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[14]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n173), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n83) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U192 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[46]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n167), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[30]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n161), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[38]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n6), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n82) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U191 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n82), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n83), .ZN(
        wrap_act_buffer_inst_int_i_data_if4[6]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U190 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[40]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n165), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[24]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n159), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[32]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n4), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n142) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U189 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[16]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n183), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[0]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n177), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[8]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n171), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n143) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U188 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n142), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n143), .ZN(
        wrap_act_buffer_inst_int_i_data_if1[0]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U187 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[40]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n165), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[24]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n159), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[32]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n4), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n126) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U186 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[16]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n183), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[0]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n177), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[8]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n171), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n127) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U185 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n126), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n127), .ZN(
        wrap_act_buffer_inst_int_i_data_if2[0]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U184 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[16]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n185), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[0]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n179), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[8]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n173), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n79) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U183 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[40]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n167), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[24]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n161), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[32]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n6), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n78) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U182 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n78), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n79), .ZN(
        wrap_act_buffer_inst_int_i_data_if5[0]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U181 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[16]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n185), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[0]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n179), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[8]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n173), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n95) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U180 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[40]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n167), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[24]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n161), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[32]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n6), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n94) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U179 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n94), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n95), .ZN(
        wrap_act_buffer_inst_int_i_data_if4[0]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U178 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[16]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n184), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[0]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n178), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[8]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n172), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n111) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U177 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[40]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n166), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[24]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n160), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[32]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n5), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n110) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U176 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n110), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n111), .ZN(
        wrap_act_buffer_inst_int_i_data_if3[0]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U175 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[19]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n186), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[3]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n180), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[11]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n174), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n57) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U174 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[43]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n168), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[27]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n162), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[35]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n7), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n56) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U173 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n56), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n57), .ZN(
        wrap_act_buffer_inst_int_i_data_if6[3]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U172 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[19]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n187), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[3]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n181), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[11]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n175), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n41) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U171 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[43]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n169), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[27]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n163), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[35]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n8), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n40) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U170 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n40), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n41), .ZN(
        wrap_act_buffer_inst_int_i_data_if7[3]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U169 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[19]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n187), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[3]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n181), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[11]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n175), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n25) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U168 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[43]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n169), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[27]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n163), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[35]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n8), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n24) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U167 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n24), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n25), .ZN(
        wrap_act_buffer_inst_int_i_data_if8[3]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U166 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[21]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n186), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[5]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n180), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[13]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n174), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n69) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U165 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[45]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n168), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[29]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n162), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[37]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n7), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n68) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U164 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n68), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n69), .ZN(
        wrap_act_buffer_inst_int_i_data_if5[5]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U163 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[21]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n186), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[5]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n180), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[13]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n174), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n53) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U162 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[45]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n168), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[29]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n162), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[37]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n7), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n52) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U161 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n52), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n53), .ZN(
        wrap_act_buffer_inst_int_i_data_if6[5]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U160 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[21]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n188), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[5]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n182), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[13]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n176), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n21) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U159 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[45]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n170), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[29]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n164), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[37]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n9), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n20) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U158 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n20), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n21), .ZN(
        wrap_act_buffer_inst_int_i_data_if8[5]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U157 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[21]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n187), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[5]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n181), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[13]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n175), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n37) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U156 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[45]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n169), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[29]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n163), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[37]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n8), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n36) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U155 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n36), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n37), .ZN(
        wrap_act_buffer_inst_int_i_data_if7[5]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U154 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[23]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n186), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[7]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n180), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[15]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n174), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n65) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U153 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[47]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n168), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[31]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n162), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[39]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n7), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n64) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U152 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n64), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n65), .ZN(
        wrap_act_buffer_inst_int_i_data_if5[7]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U151 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[23]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n186), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[7]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n180), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[15]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n174), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n49) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U150 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[47]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n168), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[31]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n162), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[39]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n7), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n48) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U149 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n48), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n49), .ZN(
        wrap_act_buffer_inst_int_i_data_if6[7]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U148 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[47]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n170), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[31]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n164), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[39]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n9), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n10) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U147 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[23]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n188), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[7]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n182), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[15]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n176), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n11) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U146 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n10), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n11), .ZN(
        wrap_act_buffer_inst_int_i_data_if8[7]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U145 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[23]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n187), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[7]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n181), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[15]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n175), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n33) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U144 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[47]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n169), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[31]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n163), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[39]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n8), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n32) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U143 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n32), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n33), .ZN(
        wrap_act_buffer_inst_int_i_data_if7[7]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U142 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[17]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n186), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[1]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n180), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[9]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n174), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n61) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U141 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[41]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n168), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[25]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n162), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[33]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n7), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n60) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U140 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n60), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n61), .ZN(
        wrap_act_buffer_inst_int_i_data_if6[1]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U139 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[17]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n187), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[1]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n181), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[9]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n175), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n29) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U138 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[41]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n169), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[25]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n163), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[33]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n8), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n28) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U137 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n28), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n29), .ZN(
        wrap_act_buffer_inst_int_i_data_if8[1]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U136 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[17]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n187), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[1]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n181), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[9]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n175), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n45) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U135 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[41]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n169), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[25]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n163), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[33]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n8), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n44) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U134 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n44), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n45), .ZN(
        wrap_act_buffer_inst_int_i_data_if7[1]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U133 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[18]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n186), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[2]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n180), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[10]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n174), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n59) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U132 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[42]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n168), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[26]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n162), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[34]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n7), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n58) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U131 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n58), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n59), .ZN(
        wrap_act_buffer_inst_int_i_data_if6[2]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U130 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[18]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n187), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[2]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n181), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[10]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n175), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n43) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U129 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[42]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n169), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[26]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n163), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[34]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n8), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n42) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U128 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n42), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n43), .ZN(
        wrap_act_buffer_inst_int_i_data_if7[2]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U127 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[18]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n187), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[2]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n181), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[10]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n175), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n27) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U126 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[42]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n169), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[26]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n163), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[34]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n8), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n26) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U125 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n26), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n27), .ZN(
        wrap_act_buffer_inst_int_i_data_if8[2]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U124 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[20]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n186), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[4]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n180), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[12]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n174), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n71) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U123 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[44]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n168), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[28]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n162), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[36]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n7), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n70) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U122 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n70), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n71), .ZN(
        wrap_act_buffer_inst_int_i_data_if5[4]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U121 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[20]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n186), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[4]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n180), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[12]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n174), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n55) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U120 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[44]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n168), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[28]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n162), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[36]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n7), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n54) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U119 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n54), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n55), .ZN(
        wrap_act_buffer_inst_int_i_data_if6[4]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U118 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[20]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n188), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[4]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n182), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[12]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n176), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n23) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U117 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[44]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n170), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[28]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n164), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[36]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n9), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n22) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U116 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n22), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n23), .ZN(
        wrap_act_buffer_inst_int_i_data_if8[4]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U115 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[20]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n187), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[4]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n181), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[12]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n175), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n39) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U114 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[44]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n169), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[28]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n163), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[36]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n8), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n38) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U113 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n38), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n39), .ZN(
        wrap_act_buffer_inst_int_i_data_if7[4]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U112 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[22]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n186), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[6]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n180), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[14]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n174), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n67) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U111 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[46]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n168), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[30]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n162), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[38]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n7), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n66) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U110 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n66), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n67), .ZN(
        wrap_act_buffer_inst_int_i_data_if5[6]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U109 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[22]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n186), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[6]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n180), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[14]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n174), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n51) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U108 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[46]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n168), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[30]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n162), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[38]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n7), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n50) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U107 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n50), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n51), .ZN(
        wrap_act_buffer_inst_int_i_data_if6[6]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U106 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[46]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n170), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[30]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n164), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[38]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n9), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n18) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U105 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[22]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n188), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[6]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n182), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[14]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n176), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n19) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U104 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n18), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n19), .ZN(
        wrap_act_buffer_inst_int_i_data_if8[6]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U103 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[22]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n187), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[6]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n181), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[14]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n175), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n35) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U102 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[46]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n169), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[30]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n163), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[38]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n8), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n34) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U101 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n34), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n35), .ZN(
        wrap_act_buffer_inst_int_i_data_if7[6]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U100 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[16]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n186), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[0]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n180), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[8]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n174), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n63) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U99 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[40]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n168), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[24]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n162), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[32]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n7), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n62) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U98 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n62), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n63), .ZN(
        wrap_act_buffer_inst_int_i_data_if6[0]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U97 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[16]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n187), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[0]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n181), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[8]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n175), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n31) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U96 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[40]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n169), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[24]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n163), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[32]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n8), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n30) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U95 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n30), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n31), .ZN(
        wrap_act_buffer_inst_int_i_data_if8[0]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U94 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[16]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n187), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[0]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n181), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[8]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n175), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n47) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U93 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[40]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n169), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[24]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n163), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[32]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n8), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n46) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U92 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n46), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n47), .ZN(
        wrap_act_buffer_inst_int_i_data_if7[0]) );
  INV_X1 wrap_act_buffer_inst_act_buffer_inst_U91 ( .A(ps_int_L0_ptr[1]), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n193) );
  AND2_X1 wrap_act_buffer_inst_act_buffer_inst_U90 ( .A1(ps_int_L0_ptr[2]), 
        .A2(wrap_act_buffer_inst_act_buffer_inst_n192), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n14) );
  AND2_X1 wrap_act_buffer_inst_act_buffer_inst_U89 ( .A1(ps_int_L0_ptr[2]), 
        .A2(ps_int_L0_ptr[0]), .ZN(wrap_act_buffer_inst_act_buffer_inst_n13)
         );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U88 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n193), .A2(ps_int_L0_ptr[0]), 
        .ZN(wrap_act_buffer_inst_act_buffer_inst_n16) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U87 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n145), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n157), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N120) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U86 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n145), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n151), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N156) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U85 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n145), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n152), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N150) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U84 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n145), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n153), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N144) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U83 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n145), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n154), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N138) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U82 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n145), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n155), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N132) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U81 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n145), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n156), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N126) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U80 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n147), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n151), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N154) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U79 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n147), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n152), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N148) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U78 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n147), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n153), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N142) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U77 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n147), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n154), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N136) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U76 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n147), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n155), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N130) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U75 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n147), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n156), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N124) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U74 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n147), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n157), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N118) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U73 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n149), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n151), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N152) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U72 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n149), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n152), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N146) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U71 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n149), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n153), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N140) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U70 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n149), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n154), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N134) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U69 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n149), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n155), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N128) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U68 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n149), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n156), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N122) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U67 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n149), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n157), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N116) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U66 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n150), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n151), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N151) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U65 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n148), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n151), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N153) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U64 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n150), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n152), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N145) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U63 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n148), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n152), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N147) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U62 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n150), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n153), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N139) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U61 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n148), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n153), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N141) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U60 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n150), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n154), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N133) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U59 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n148), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n154), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N135) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U58 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n150), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n155), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N127) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U57 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n148), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n155), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N129) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U56 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n150), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n156), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N121) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U55 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n148), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n156), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N123) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U54 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n150), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n157), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N115) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U53 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n148), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n157), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N117) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U52 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n146), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n151), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N155) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U51 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n146), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n152), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N149) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U50 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n146), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n153), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N143) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U49 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n146), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n154), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N137) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U48 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n146), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n155), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N131) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U47 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n146), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n156), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N125) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U46 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n146), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n157), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N119) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U45 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n144), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n150), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N157) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U44 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n144), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n149), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N158) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U43 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n144), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n148), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N159) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U42 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n144), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n147), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N160) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U41 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n144), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n146), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N161) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U40 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n144), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n145), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N162) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U39 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n15), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n165) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U38 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n15), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n167) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U37 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n15), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n168) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U36 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n15), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n166) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U35 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n14), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n171) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U34 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n17), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n4) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U33 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n17), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n6) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U32 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n17), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n7) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U31 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n17), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n5) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U30 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n17), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n8) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U29 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n13), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n177) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U28 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n13), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n179) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U27 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n13), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n178) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U26 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n16), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n159) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U25 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n16), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n161) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U24 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n16), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n160) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U23 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n193), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n192), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n12) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U22 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n15), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n169) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U21 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n14), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n173) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U20 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n14), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n174) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U19 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n14), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n172) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U18 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n14), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n175) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U17 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n13), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n180) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U16 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n13), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n181) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U15 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n16), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n162) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U14 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n16), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n163) );
  AND4_X1 wrap_act_buffer_inst_act_buffer_inst_U13 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n144), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n151), .A3(
        wrap_act_buffer_inst_act_buffer_inst_n152), .A4(
        wrap_act_buffer_inst_act_buffer_inst_n153), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n158) );
  NAND4_X1 wrap_act_buffer_inst_act_buffer_inst_U12 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n155), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n154), .A3(
        wrap_act_buffer_inst_act_buffer_inst_n156), .A4(
        wrap_act_buffer_inst_act_buffer_inst_n158), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n157) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U11 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n12), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n183) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U10 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n12), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n185) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U9 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n12), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n186) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U8 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n12), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n184) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U7 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n12), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n187) );
  INV_X8 wrap_act_buffer_inst_act_buffer_inst_U6 ( .A(rst), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n3) );
  INV_X8 wrap_act_buffer_inst_act_buffer_inst_U5 ( .A(rst), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n2) );
  INV_X8 wrap_act_buffer_inst_act_buffer_inst_U4 ( .A(rst), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n1) );
  NOR3_X1 wrap_act_buffer_inst_act_buffer_inst_U3 ( .A1(ps_int_L0_ptr[1]), 
        .A2(ps_int_L0_ptr[2]), .A3(ps_int_L0_ptr[0]), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n15) );
  NOR3_X1 wrap_act_buffer_inst_act_buffer_inst_U2 ( .A1(ps_int_L0_ptr[1]), 
        .A2(ps_int_L0_ptr[2]), .A3(wrap_act_buffer_inst_act_buffer_inst_n192), 
        .ZN(wrap_act_buffer_inst_act_buffer_inst_n17) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_4__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4624), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[8]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_4__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4624), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[9]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_4__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4624), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[10]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_4__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4624), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[11]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_4__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4624), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[12]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_4__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4624), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[13]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_4__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4624), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[14]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_4__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4624), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[15]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_5__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4629), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[0]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_5__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4629), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[1]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_5__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4629), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[2]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_5__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4629), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[3]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_5__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4629), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[4]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_5__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4629), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[5]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_5__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4629), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[6]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_5__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4629), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[7]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_0__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4634), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[40]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_0__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4634), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[41]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_0__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4634), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[42]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_0__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4634), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[43]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_0__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4634), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[44]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_0__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4634), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[45]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_0__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4634), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[46]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_0__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4634), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[47]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_1__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4639), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[32]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_1__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4639), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[33]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_1__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4639), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[34]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_1__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4639), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[35]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_1__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4639), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[36]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_1__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4639), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[37]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_1__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4639), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[38]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_1__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4639), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[39]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_2__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4644), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[24]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_2__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4644), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[25]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_2__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4644), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[26]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_2__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4644), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[27]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_2__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4644), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[28]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_2__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4644), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[29]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_2__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4644), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[30]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_2__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4644), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[31]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_3__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4649), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[16]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_3__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4649), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[17]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_3__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4649), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[18]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_3__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4649), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[19]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_3__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4649), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[20]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_3__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4649), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[21]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_3__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4649), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[22]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_3__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4649), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[23]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_4__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4654), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[8]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_4__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4654), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[9]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_4__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4654), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[10]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_4__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4654), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[11]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_4__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4654), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[12]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_4__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4654), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[13]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_4__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4654), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[14]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_4__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4654), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[15]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_5__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4659), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[0]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_5__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4659), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[1]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_5__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4659), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[2]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_5__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4659), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[3]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_5__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4659), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[4]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_5__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4659), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[5]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_5__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4659), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[6]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_5__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4659), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[7]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_0__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4664), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[40]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_0__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4664), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[41]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_0__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4664), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[42]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_0__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4664), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[43]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_0__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4664), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[44]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_0__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4664), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[45]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_0__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4664), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[46]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_0__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4664), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[47]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_1__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4669), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[32]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_1__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4669), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[33]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_1__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4669), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[34]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_1__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4669), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[35]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_1__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4669), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[36]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_1__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4669), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[37]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_1__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4669), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[38]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_1__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4669), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[39]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_2__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4674), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[24]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_2__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4674), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[25]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_2__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4674), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[26]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_2__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4674), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[27]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_2__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4674), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[28]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_2__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4674), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[29]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_2__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4674), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[30]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_2__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4674), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[31]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_3__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4679), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[16]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_3__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4679), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[17]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_3__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4679), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[18]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_3__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4679), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[19]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_3__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4679), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[20]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_3__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4679), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[21]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_3__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4679), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[22]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_3__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4679), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[23]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_4__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4684), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[8]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_4__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4684), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[9]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_4__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4684), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[10]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_4__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4684), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[11]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_4__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4684), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[12]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_4__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4684), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[13]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_4__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4684), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[14]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_4__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4684), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[15]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_5__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4689), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[0]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_5__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4689), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[1]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_5__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4689), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[2]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_5__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4689), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[3]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_5__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4689), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[4]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_5__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4689), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[5]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_5__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4689), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[6]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_5__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4689), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[7]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_0__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4694), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[40]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_0__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4694), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[41]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_0__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4694), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[42]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_0__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4694), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[43]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_0__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4694), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[44]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_0__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4694), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[45]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_0__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4694), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[46]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_0__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4694), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[47]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_1__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4699), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[32]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_1__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4699), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[33]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_1__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4699), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[34]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_1__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4699), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[35]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_1__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4699), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[36]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_1__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4699), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[37]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_1__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4699), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[38]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_1__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4699), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[39]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_2__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4704), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[24]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_2__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4704), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[25]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_2__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4704), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[26]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_2__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4704), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[27]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_2__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4704), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[28]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_2__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4704), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[29]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_2__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4704), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[30]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_2__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4704), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[31]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_3__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4709), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[16]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_3__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4709), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[17]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_3__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4709), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[18]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_3__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4709), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[19]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_3__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4709), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[20]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_3__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4709), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[21]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_3__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4709), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[22]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_3__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4709), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[23]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_4__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4714), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[8]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_4__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4714), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[9]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_4__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4714), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[10]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_4__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4714), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[11]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_4__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4714), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[12]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_4__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4714), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[13]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_4__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4714), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[14]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_4__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4714), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[15]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_5__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4719), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[0]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_5__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4719), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[1]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_5__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4719), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[2]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_5__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4719), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[3]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_5__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4719), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[4]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_5__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4719), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[5]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_5__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4719), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[6]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_5__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4719), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[7]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_0__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4724), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[40]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_0__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4724), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[41]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_0__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4724), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[42]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_0__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4724), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[43]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_0__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4724), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[44]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_0__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4724), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[45]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_0__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4724), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[46]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_0__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4724), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[47]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_1__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4729), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[32]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_1__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4729), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[33]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_1__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4729), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[34]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_1__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4729), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[35]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_1__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4729), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[36]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_1__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4729), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[37]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_1__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4729), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[38]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_1__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4729), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[39]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_2__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4734), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[24]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_2__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4734), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[25]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_2__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4734), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[26]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_2__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4734), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[27]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_2__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4734), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[28]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_2__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4734), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[29]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_2__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4734), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[30]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_2__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4734), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[31]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_3__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4739), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[16]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_3__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4739), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[17]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_3__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4739), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[18]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_3__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4739), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[19]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_3__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4739), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[20]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_3__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4739), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[21]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_3__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4739), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[22]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_3__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4739), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[23]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_4__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4744), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[8]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_4__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4744), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[9]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_4__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4744), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[10]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_4__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4744), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[11]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_4__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4744), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[12]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_4__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4744), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[13]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_4__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4744), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[14]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_4__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4744), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[15]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_5__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4749), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[0]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_5__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4749), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[1]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_5__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4749), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[2]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_5__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4749), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[3]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_5__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4749), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[4]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_5__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4749), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[5]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_5__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4749), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[6]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_5__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4749), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[7]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_0__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4754), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[40]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_0__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4754), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[41]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_0__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4754), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[42]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_0__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4754), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[43]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_0__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4754), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[44]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_0__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4754), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[45]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_0__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4754), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[46]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_0__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4754), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[47]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_1__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4759), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[32]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_1__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4759), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[33]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_1__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4759), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[34]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_1__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4759), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[35]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_1__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4759), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[36]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_1__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4759), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[37]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_1__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4759), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[38]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_1__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4759), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[39]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_2__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4764), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[24]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_2__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4764), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[25]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_2__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4764), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[26]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_2__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4764), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[27]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_2__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4764), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[28]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_2__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4764), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[29]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_2__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4764), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[30]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_2__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4764), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[31]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_3__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4769), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[16]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_3__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4769), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[17]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_3__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4769), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[18]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_3__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4769), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[19]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_3__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4769), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[20]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_3__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4769), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[21]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_3__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4769), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[22]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_3__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4769), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[23]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_4__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4774), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[8]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_4__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4774), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[9]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_4__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4774), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[10]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_4__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4774), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[11]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_4__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4774), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[12]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_4__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4774), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[13]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_4__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4774), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[14]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_4__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4774), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[15]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_5__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4779), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[0]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_5__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4779), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[1]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_5__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4779), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[2]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_5__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4779), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[3]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_5__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4779), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[4]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_5__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4779), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[5]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_5__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4779), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[6]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_5__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4779), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[7]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_0__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4784), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[40]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_0__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4784), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[41]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_0__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4784), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[42]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_0__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4784), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[43]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_0__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4784), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[44]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_0__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4784), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[45]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_0__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4784), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[46]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_0__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4784), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[47]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_1__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4789), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[32]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_1__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4789), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[33]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_1__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4789), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[34]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_1__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4789), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[35]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_1__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4789), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[36]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_1__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4789), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[37]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_1__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4789), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[38]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_1__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4789), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[39]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_2__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4794), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[24]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_2__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4794), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[25]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_2__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4794), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[26]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_2__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4794), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[27]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_2__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4794), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[28]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_2__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4794), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[29]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_2__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4794), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[30]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_2__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4794), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[31]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_3__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4799), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[16]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_3__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4799), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[17]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_3__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4799), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[18]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_3__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4799), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[19]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_3__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4799), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[20]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_3__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4799), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[21]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_3__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4799), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[22]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_3__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4799), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[23]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_4__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4804), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[8]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_4__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4804), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[9]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_4__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4804), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[10]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_4__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4804), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[11]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_4__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4804), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[12]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_4__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4804), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[13]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_4__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4804), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[14]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_4__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4804), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[15]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_5__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4809), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[0]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_5__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4809), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[1]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_5__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4809), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[2]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_5__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4809), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[3]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_5__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4809), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[4]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_5__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4809), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[5]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_5__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4809), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[6]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_5__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4809), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[7]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_0__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4814), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[40]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_0__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4814), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[41]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_0__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4814), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[42]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_0__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4814), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[43]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_0__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4814), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[44]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_0__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4814), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[45]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_0__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4814), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[46]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_0__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4814), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[47]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_1__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4819), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[32]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_1__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4819), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[33]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_1__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4819), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[34]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_1__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4819), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[35]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_1__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4819), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[36]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_1__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4819), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[37]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_1__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4819), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[38]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_1__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4819), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[39]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_2__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4824), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[24]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_2__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4824), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[25]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_2__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4824), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[26]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_2__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4824), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[27]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_2__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4824), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[28]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_2__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4824), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[29]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_2__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4824), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[30]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_2__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4824), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[31]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_3__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4829), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[16]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_3__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4829), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[17]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_3__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4829), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[18]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_3__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4829), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[19]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_3__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4829), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[20]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_3__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4829), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[21]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_3__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4829), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[22]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_3__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4829), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[23]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_4__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4834), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[8]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_4__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4834), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[9]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_4__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4834), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[10]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_4__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4834), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[11]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_4__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4834), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[12]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_4__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4834), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[13]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_4__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4834), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[14]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_4__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4834), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[15]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_5__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4839), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[0]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_5__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4839), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[1]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_5__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4839), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[2]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_5__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4839), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[3]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_5__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4839), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[4]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_5__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4839), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[5]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_5__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4839), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[6]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_5__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4839), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[7]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_0__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4603), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[40]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_0__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4603), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[41]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_0__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4603), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[42]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_0__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4603), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[43]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_0__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4603), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[44]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_0__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4603), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[45]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_0__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4603), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[46]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_0__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4603), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[47]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_1__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4609), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[32]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_1__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4609), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[33]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_1__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4609), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[34]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_1__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4609), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[35]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_1__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4609), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[36]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_1__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4609), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[37]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_1__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4609), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[38]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_1__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4609), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[39]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_2__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4614), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[24]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_2__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4614), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[25]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_2__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4614), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[26]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_2__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4614), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[27]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_2__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4614), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[28]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_2__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4614), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[29]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_2__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4614), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[30]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_2__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4614), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[31]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_3__0_ ( .D(
        i_acth[8]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4619), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[16]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_3__1_ ( .D(
        i_acth[9]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4619), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[17]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_3__2_ ( .D(
        i_acth[10]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4619), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[18]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_3__3_ ( .D(
        i_acth[11]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4619), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[19]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_3__4_ ( .D(
        i_acth[12]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4619), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[20]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_3__5_ ( .D(
        i_acth[13]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4619), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n1), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[21]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_3__6_ ( .D(
        i_acth[14]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4619), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n2), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[22]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_3__7_ ( .D(
        i_acth[15]), .CK(wrap_act_buffer_inst_act_buffer_inst_net4619), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n3), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[23]) );
  NAND3_X1 wrap_act_buffer_inst_act_buffer_inst_U271 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n189), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n191), .A3(int_L1_ptr[1]), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n155) );
  NAND3_X1 wrap_act_buffer_inst_act_buffer_inst_U270 ( .A1(int_L1_ptr[0]), 
        .A2(wrap_act_buffer_inst_act_buffer_inst_n191), .A3(int_L1_ptr[1]), 
        .ZN(wrap_act_buffer_inst_act_buffer_inst_n154) );
  NAND3_X1 wrap_act_buffer_inst_act_buffer_inst_U269 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n190), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n191), .A3(int_L1_ptr[0]), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n156) );
  NAND3_X1 wrap_act_buffer_inst_act_buffer_inst_U268 ( .A1(int_L1_ptr[1]), 
        .A2(int_L1_ptr[0]), .A3(int_L1_ptr[2]), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n144) );
  NAND3_X1 wrap_act_buffer_inst_act_buffer_inst_U267 ( .A1(int_L1_ptr[1]), 
        .A2(wrap_act_buffer_inst_act_buffer_inst_n189), .A3(int_L1_ptr[2]), 
        .ZN(wrap_act_buffer_inst_act_buffer_inst_n151) );
  NAND3_X1 wrap_act_buffer_inst_act_buffer_inst_U266 ( .A1(int_L1_ptr[0]), 
        .A2(wrap_act_buffer_inst_act_buffer_inst_n190), .A3(int_L1_ptr[2]), 
        .ZN(wrap_act_buffer_inst_act_buffer_inst_n152) );
  NAND3_X1 wrap_act_buffer_inst_act_buffer_inst_U265 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n189), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n190), .A3(int_L1_ptr[2]), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n153) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data1_reg_0__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N120), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4603) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data1_reg_1__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N119), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4609) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data1_reg_2__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N118), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4614) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data1_reg_3__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N117), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4619) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data1_reg_4__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N116), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4624) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data1_reg_5__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N115), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4629) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data2_reg_0__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N126), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4634) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data2_reg_1__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N125), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4639) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data2_reg_2__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N124), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4644) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data2_reg_3__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N123), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4649) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data2_reg_4__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N122), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4654) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data2_reg_5__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N121), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4659) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data3_reg_0__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N132), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4664) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data3_reg_1__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N131), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4669) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data3_reg_2__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N130), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4674) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data3_reg_3__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N129), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4679) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data3_reg_4__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N128), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4684) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data3_reg_5__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N127), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4689) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data4_reg_0__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N138), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4694) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data4_reg_1__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N137), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4699) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data4_reg_2__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N136), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4704) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data4_reg_3__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N135), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4709) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data4_reg_4__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N134), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4714) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data4_reg_5__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N133), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4719) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data5_reg_0__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N144), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4724) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data5_reg_1__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N143), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4729) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data5_reg_2__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N142), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4734) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data5_reg_3__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N141), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4739) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data5_reg_4__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N140), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4744) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data5_reg_5__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N139), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4749) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data6_reg_0__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N150), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4754) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data6_reg_1__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N149), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4759) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data6_reg_2__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N148), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4764) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data6_reg_3__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N147), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4769) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data6_reg_4__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N146), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4774) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data6_reg_5__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N145), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4779) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data7_reg_0__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N156), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4784) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data7_reg_1__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N155), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4789) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data7_reg_2__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N154), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4794) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data7_reg_3__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N153), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4799) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data7_reg_4__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N152), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4804) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data7_reg_5__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N151), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4809) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data8_reg_0__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N162), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4814) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data8_reg_1__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N161), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4819) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data8_reg_2__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N160), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4824) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data8_reg_3__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N159), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4829) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data8_reg_4__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N158), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4834) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data8_reg_5__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N157), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4839) );
  NOR3_X4 wrap_act_buffer_inst_act_if_inst_U392 ( .A1(ps_int_hmode_cnt[0]), 
        .A2(1'b0), .A3(wrap_act_buffer_inst_act_if_inst_n312), .ZN(
        wrap_act_buffer_inst_act_if_inst_n7) );
  CLKBUF_X1 wrap_act_buffer_inst_act_if_inst_U391 ( .A(int_L1_ptr[0]), .Z(
        wrap_act_buffer_inst_act_if_inst_n305) );
  CLKBUF_X1 wrap_act_buffer_inst_act_if_inst_U390 ( .A(int_L1_ptr[1]), .Z(
        wrap_act_buffer_inst_act_if_inst_n299) );
  CLKBUF_X1 wrap_act_buffer_inst_act_if_inst_U389 ( .A(int_L1_ptr[2]), .Z(
        wrap_act_buffer_inst_act_if_inst_n293) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U388 ( .A(
        wrap_act_buffer_inst_act_if_inst_n130), .B(
        wrap_act_buffer_inst_act_if_inst_n131), .S(
        wrap_act_buffer_inst_act_if_inst_n298), .Z(
        wrap_act_buffer_inst_act_if_inst_n164) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U387 ( .A(
        wrap_act_buffer_inst_act_if_inst_n124), .B(
        wrap_act_buffer_inst_act_if_inst_n125), .S(
        wrap_act_buffer_inst_act_if_inst_n298), .Z(
        wrap_act_buffer_inst_act_if_inst_n163) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U386 ( .A(
        wrap_act_buffer_inst_act_if_inst_n118), .B(
        wrap_act_buffer_inst_act_if_inst_n119), .S(
        wrap_act_buffer_inst_act_if_inst_n298), .Z(
        wrap_act_buffer_inst_act_if_inst_n162) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U385 ( .A(
        wrap_act_buffer_inst_act_if_inst_n112), .B(
        wrap_act_buffer_inst_act_if_inst_n113), .S(
        wrap_act_buffer_inst_act_if_inst_n298), .Z(
        wrap_act_buffer_inst_act_if_inst_n161) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U384 ( .A(
        wrap_act_buffer_inst_act_if_inst_n106), .B(
        wrap_act_buffer_inst_act_if_inst_n107), .S(
        wrap_act_buffer_inst_act_if_inst_n298), .Z(
        wrap_act_buffer_inst_act_if_inst_n160) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U383 ( .A(
        wrap_act_buffer_inst_act_if_inst_n100), .B(
        wrap_act_buffer_inst_act_if_inst_n101), .S(
        wrap_act_buffer_inst_act_if_inst_n298), .Z(
        wrap_act_buffer_inst_act_if_inst_n159) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U382 ( .A(
        wrap_act_buffer_inst_act_if_inst_n94), .B(
        wrap_act_buffer_inst_act_if_inst_n95), .S(
        wrap_act_buffer_inst_act_if_inst_n298), .Z(
        wrap_act_buffer_inst_act_if_inst_n158) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U381 ( .A(
        wrap_act_buffer_inst_act_if_inst_n88), .B(
        wrap_act_buffer_inst_act_if_inst_n89), .S(
        wrap_act_buffer_inst_act_if_inst_n298), .Z(
        wrap_act_buffer_inst_act_if_inst_n157) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U380 ( .A(
        wrap_act_buffer_inst_act_if_inst_n82), .B(
        wrap_act_buffer_inst_act_if_inst_n83), .S(
        wrap_act_buffer_inst_act_if_inst_n298), .Z(
        wrap_act_buffer_inst_act_if_inst_n156) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U379 ( .A(
        wrap_act_buffer_inst_act_if_inst_n76), .B(
        wrap_act_buffer_inst_act_if_inst_n77), .S(
        wrap_act_buffer_inst_act_if_inst_n298), .Z(
        wrap_act_buffer_inst_act_if_inst_n155) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U378 ( .A(
        wrap_act_buffer_inst_act_if_inst_n70), .B(
        wrap_act_buffer_inst_act_if_inst_n71), .S(
        wrap_act_buffer_inst_act_if_inst_n298), .Z(
        wrap_act_buffer_inst_act_if_inst_n154) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U377 ( .A(
        wrap_act_buffer_inst_act_if_inst_n64), .B(
        wrap_act_buffer_inst_act_if_inst_n65), .S(
        wrap_act_buffer_inst_act_if_inst_n298), .Z(
        wrap_act_buffer_inst_act_if_inst_n153) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U376 ( .A(
        wrap_act_buffer_inst_act_if_inst_n58), .B(
        wrap_act_buffer_inst_act_if_inst_n59), .S(
        wrap_act_buffer_inst_act_if_inst_n297), .Z(
        wrap_act_buffer_inst_act_if_inst_n152) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U375 ( .A(
        wrap_act_buffer_inst_act_if_inst_n52), .B(
        wrap_act_buffer_inst_act_if_inst_n53), .S(
        wrap_act_buffer_inst_act_if_inst_n297), .Z(
        wrap_act_buffer_inst_act_if_inst_n151) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U374 ( .A(
        wrap_act_buffer_inst_act_if_inst_n46), .B(
        wrap_act_buffer_inst_act_if_inst_n47), .S(
        wrap_act_buffer_inst_act_if_inst_n297), .Z(
        wrap_act_buffer_inst_act_if_inst_n150) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U373 ( .A(
        wrap_act_buffer_inst_act_if_inst_n40), .B(
        wrap_act_buffer_inst_act_if_inst_n41), .S(
        wrap_act_buffer_inst_act_if_inst_n297), .Z(
        wrap_act_buffer_inst_act_if_inst_n149) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U372 ( .A(
        wrap_act_buffer_inst_act_if_inst_n127), .B(
        wrap_act_buffer_inst_act_if_inst_n128), .S(
        wrap_act_buffer_inst_act_if_inst_n297), .Z(
        wrap_act_buffer_inst_act_if_inst_n148) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U371 ( .A(
        wrap_act_buffer_inst_act_if_inst_n121), .B(
        wrap_act_buffer_inst_act_if_inst_n122), .S(
        wrap_act_buffer_inst_act_if_inst_n297), .Z(
        wrap_act_buffer_inst_act_if_inst_n147) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U370 ( .A(
        wrap_act_buffer_inst_act_if_inst_n115), .B(
        wrap_act_buffer_inst_act_if_inst_n116), .S(
        wrap_act_buffer_inst_act_if_inst_n297), .Z(
        wrap_act_buffer_inst_act_if_inst_n146) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U369 ( .A(
        wrap_act_buffer_inst_act_if_inst_n109), .B(
        wrap_act_buffer_inst_act_if_inst_n110), .S(
        wrap_act_buffer_inst_act_if_inst_n297), .Z(
        wrap_act_buffer_inst_act_if_inst_n145) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U368 ( .A(
        wrap_act_buffer_inst_act_if_inst_n103), .B(
        wrap_act_buffer_inst_act_if_inst_n104), .S(
        wrap_act_buffer_inst_act_if_inst_n297), .Z(
        wrap_act_buffer_inst_act_if_inst_n144) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U367 ( .A(
        wrap_act_buffer_inst_act_if_inst_n97), .B(
        wrap_act_buffer_inst_act_if_inst_n98), .S(
        wrap_act_buffer_inst_act_if_inst_n297), .Z(
        wrap_act_buffer_inst_act_if_inst_n143) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U366 ( .A(
        wrap_act_buffer_inst_act_if_inst_n91), .B(
        wrap_act_buffer_inst_act_if_inst_n92), .S(
        wrap_act_buffer_inst_act_if_inst_n297), .Z(
        wrap_act_buffer_inst_act_if_inst_n142) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U365 ( .A(
        wrap_act_buffer_inst_act_if_inst_n85), .B(
        wrap_act_buffer_inst_act_if_inst_n86), .S(
        wrap_act_buffer_inst_act_if_inst_n297), .Z(
        wrap_act_buffer_inst_act_if_inst_n141) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U364 ( .A(
        wrap_act_buffer_inst_act_if_inst_n79), .B(
        wrap_act_buffer_inst_act_if_inst_n80), .S(
        wrap_act_buffer_inst_act_if_inst_n296), .Z(
        wrap_act_buffer_inst_act_if_inst_n140) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U363 ( .A(
        wrap_act_buffer_inst_act_if_inst_n73), .B(
        wrap_act_buffer_inst_act_if_inst_n74), .S(
        wrap_act_buffer_inst_act_if_inst_n296), .Z(
        wrap_act_buffer_inst_act_if_inst_n139) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U362 ( .A(
        wrap_act_buffer_inst_act_if_inst_n67), .B(
        wrap_act_buffer_inst_act_if_inst_n68), .S(
        wrap_act_buffer_inst_act_if_inst_n296), .Z(
        wrap_act_buffer_inst_act_if_inst_n138) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U361 ( .A(
        wrap_act_buffer_inst_act_if_inst_n61), .B(
        wrap_act_buffer_inst_act_if_inst_n62), .S(
        wrap_act_buffer_inst_act_if_inst_n296), .Z(
        wrap_act_buffer_inst_act_if_inst_n137) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U360 ( .A(
        wrap_act_buffer_inst_act_if_inst_n55), .B(
        wrap_act_buffer_inst_act_if_inst_n56), .S(
        wrap_act_buffer_inst_act_if_inst_n296), .Z(
        wrap_act_buffer_inst_act_if_inst_n136) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U359 ( .A(
        wrap_act_buffer_inst_act_if_inst_n49), .B(
        wrap_act_buffer_inst_act_if_inst_n50), .S(
        wrap_act_buffer_inst_act_if_inst_n296), .Z(
        wrap_act_buffer_inst_act_if_inst_n135) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U358 ( .A(
        wrap_act_buffer_inst_act_if_inst_n43), .B(
        wrap_act_buffer_inst_act_if_inst_n44), .S(
        wrap_act_buffer_inst_act_if_inst_n296), .Z(
        wrap_act_buffer_inst_act_if_inst_n134) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U357 ( .A(
        wrap_act_buffer_inst_act_if_inst_n1), .B(
        wrap_act_buffer_inst_act_if_inst_n2), .S(
        wrap_act_buffer_inst_act_if_inst_n296), .Z(
        wrap_act_buffer_inst_act_if_inst_n133) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U356 ( .A(
        wrap_act_buffer_inst_act_if_inst_n131), .B(
        wrap_act_buffer_inst_act_if_inst_n130), .S(
        wrap_act_buffer_inst_act_if_inst_n296), .Z(
        wrap_act_buffer_inst_act_if_inst_n132) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U355 ( .A(
        wrap_act_buffer_inst_act_if_inst_n180), .B(
        wrap_act_buffer_inst_act_if_inst_n172), .S(
        wrap_act_buffer_inst_act_if_inst_n310), .Z(
        wrap_act_buffer_inst_act_if_inst_n131) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U354 ( .A(
        wrap_act_buffer_inst_act_if_inst_n226), .B(
        wrap_act_buffer_inst_act_if_inst_n204), .S(
        wrap_act_buffer_inst_act_if_inst_n310), .Z(
        wrap_act_buffer_inst_act_if_inst_n130) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U353 ( .A(
        wrap_act_buffer_inst_act_if_inst_n128), .B(
        wrap_act_buffer_inst_act_if_inst_n127), .S(
        wrap_act_buffer_inst_act_if_inst_n296), .Z(
        wrap_act_buffer_inst_act_if_inst_n129) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U352 ( .A(
        wrap_act_buffer_inst_act_if_inst_n288), .B(
        wrap_act_buffer_inst_act_if_inst_n250), .S(
        wrap_act_buffer_inst_act_if_inst_n310), .Z(
        wrap_act_buffer_inst_act_if_inst_n128) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U351 ( .A(
        wrap_act_buffer_inst_act_if_inst_n196), .B(
        wrap_act_buffer_inst_act_if_inst_n188), .S(
        wrap_act_buffer_inst_act_if_inst_n310), .Z(
        wrap_act_buffer_inst_act_if_inst_n127) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U350 ( .A(
        wrap_act_buffer_inst_act_if_inst_n125), .B(
        wrap_act_buffer_inst_act_if_inst_n124), .S(
        wrap_act_buffer_inst_act_if_inst_n296), .Z(
        wrap_act_buffer_inst_act_if_inst_n126) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U349 ( .A(
        wrap_act_buffer_inst_act_if_inst_n179), .B(
        wrap_act_buffer_inst_act_if_inst_n171), .S(
        wrap_act_buffer_inst_act_if_inst_n310), .Z(
        wrap_act_buffer_inst_act_if_inst_n125) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U348 ( .A(
        wrap_act_buffer_inst_act_if_inst_n223), .B(
        wrap_act_buffer_inst_act_if_inst_n203), .S(
        wrap_act_buffer_inst_act_if_inst_n310), .Z(
        wrap_act_buffer_inst_act_if_inst_n124) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U347 ( .A(
        wrap_act_buffer_inst_act_if_inst_n122), .B(
        wrap_act_buffer_inst_act_if_inst_n121), .S(
        wrap_act_buffer_inst_act_if_inst_n296), .Z(
        wrap_act_buffer_inst_act_if_inst_n123) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U346 ( .A(
        wrap_act_buffer_inst_act_if_inst_n283), .B(
        wrap_act_buffer_inst_act_if_inst_n247), .S(
        wrap_act_buffer_inst_act_if_inst_n310), .Z(
        wrap_act_buffer_inst_act_if_inst_n122) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U345 ( .A(
        wrap_act_buffer_inst_act_if_inst_n195), .B(
        wrap_act_buffer_inst_act_if_inst_n187), .S(
        wrap_act_buffer_inst_act_if_inst_n310), .Z(
        wrap_act_buffer_inst_act_if_inst_n121) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U344 ( .A(
        wrap_act_buffer_inst_act_if_inst_n119), .B(
        wrap_act_buffer_inst_act_if_inst_n118), .S(
        wrap_act_buffer_inst_act_if_inst_n295), .Z(
        wrap_act_buffer_inst_act_if_inst_n120) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U343 ( .A(
        wrap_act_buffer_inst_act_if_inst_n178), .B(
        wrap_act_buffer_inst_act_if_inst_n170), .S(
        wrap_act_buffer_inst_act_if_inst_n310), .Z(
        wrap_act_buffer_inst_act_if_inst_n119) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U342 ( .A(
        wrap_act_buffer_inst_act_if_inst_n220), .B(
        wrap_act_buffer_inst_act_if_inst_n202), .S(
        wrap_act_buffer_inst_act_if_inst_n310), .Z(
        wrap_act_buffer_inst_act_if_inst_n118) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U341 ( .A(
        wrap_act_buffer_inst_act_if_inst_n116), .B(
        wrap_act_buffer_inst_act_if_inst_n115), .S(
        wrap_act_buffer_inst_act_if_inst_n295), .Z(
        wrap_act_buffer_inst_act_if_inst_n117) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U340 ( .A(
        wrap_act_buffer_inst_act_if_inst_n278), .B(
        wrap_act_buffer_inst_act_if_inst_n244), .S(
        wrap_act_buffer_inst_act_if_inst_n310), .Z(
        wrap_act_buffer_inst_act_if_inst_n116) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U339 ( .A(
        wrap_act_buffer_inst_act_if_inst_n194), .B(
        wrap_act_buffer_inst_act_if_inst_n186), .S(
        wrap_act_buffer_inst_act_if_inst_n310), .Z(
        wrap_act_buffer_inst_act_if_inst_n115) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U338 ( .A(
        wrap_act_buffer_inst_act_if_inst_n113), .B(
        wrap_act_buffer_inst_act_if_inst_n112), .S(
        wrap_act_buffer_inst_act_if_inst_n295), .Z(
        wrap_act_buffer_inst_act_if_inst_n114) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U337 ( .A(
        wrap_act_buffer_inst_act_if_inst_n177), .B(
        wrap_act_buffer_inst_act_if_inst_n169), .S(
        wrap_act_buffer_inst_act_if_inst_n309), .Z(
        wrap_act_buffer_inst_act_if_inst_n113) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U336 ( .A(
        wrap_act_buffer_inst_act_if_inst_n217), .B(
        wrap_act_buffer_inst_act_if_inst_n201), .S(
        wrap_act_buffer_inst_act_if_inst_n309), .Z(
        wrap_act_buffer_inst_act_if_inst_n112) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U335 ( .A(
        wrap_act_buffer_inst_act_if_inst_n110), .B(
        wrap_act_buffer_inst_act_if_inst_n109), .S(
        wrap_act_buffer_inst_act_if_inst_n295), .Z(
        wrap_act_buffer_inst_act_if_inst_n111) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U334 ( .A(
        wrap_act_buffer_inst_act_if_inst_n273), .B(
        wrap_act_buffer_inst_act_if_inst_n241), .S(
        wrap_act_buffer_inst_act_if_inst_n309), .Z(
        wrap_act_buffer_inst_act_if_inst_n110) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U333 ( .A(
        wrap_act_buffer_inst_act_if_inst_n193), .B(
        wrap_act_buffer_inst_act_if_inst_n185), .S(
        wrap_act_buffer_inst_act_if_inst_n309), .Z(
        wrap_act_buffer_inst_act_if_inst_n109) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U332 ( .A(
        wrap_act_buffer_inst_act_if_inst_n107), .B(
        wrap_act_buffer_inst_act_if_inst_n106), .S(
        wrap_act_buffer_inst_act_if_inst_n295), .Z(
        wrap_act_buffer_inst_act_if_inst_n108) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U331 ( .A(
        wrap_act_buffer_inst_act_if_inst_n176), .B(
        wrap_act_buffer_inst_act_if_inst_n168), .S(
        wrap_act_buffer_inst_act_if_inst_n309), .Z(
        wrap_act_buffer_inst_act_if_inst_n107) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U330 ( .A(
        wrap_act_buffer_inst_act_if_inst_n214), .B(
        wrap_act_buffer_inst_act_if_inst_n200), .S(
        wrap_act_buffer_inst_act_if_inst_n309), .Z(
        wrap_act_buffer_inst_act_if_inst_n106) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U329 ( .A(
        wrap_act_buffer_inst_act_if_inst_n104), .B(
        wrap_act_buffer_inst_act_if_inst_n103), .S(
        wrap_act_buffer_inst_act_if_inst_n295), .Z(
        wrap_act_buffer_inst_act_if_inst_n105) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U328 ( .A(
        wrap_act_buffer_inst_act_if_inst_n268), .B(
        wrap_act_buffer_inst_act_if_inst_n238), .S(
        wrap_act_buffer_inst_act_if_inst_n309), .Z(
        wrap_act_buffer_inst_act_if_inst_n104) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U327 ( .A(
        wrap_act_buffer_inst_act_if_inst_n192), .B(
        wrap_act_buffer_inst_act_if_inst_n184), .S(
        wrap_act_buffer_inst_act_if_inst_n309), .Z(
        wrap_act_buffer_inst_act_if_inst_n103) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U326 ( .A(
        wrap_act_buffer_inst_act_if_inst_n101), .B(
        wrap_act_buffer_inst_act_if_inst_n100), .S(
        wrap_act_buffer_inst_act_if_inst_n295), .Z(
        wrap_act_buffer_inst_act_if_inst_n102) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U325 ( .A(
        wrap_act_buffer_inst_act_if_inst_n175), .B(
        wrap_act_buffer_inst_act_if_inst_n167), .S(
        wrap_act_buffer_inst_act_if_inst_n309), .Z(
        wrap_act_buffer_inst_act_if_inst_n101) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U324 ( .A(
        wrap_act_buffer_inst_act_if_inst_n211), .B(
        wrap_act_buffer_inst_act_if_inst_n199), .S(
        wrap_act_buffer_inst_act_if_inst_n309), .Z(
        wrap_act_buffer_inst_act_if_inst_n100) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U323 ( .A(
        wrap_act_buffer_inst_act_if_inst_n98), .B(
        wrap_act_buffer_inst_act_if_inst_n97), .S(
        wrap_act_buffer_inst_act_if_inst_n295), .Z(
        wrap_act_buffer_inst_act_if_inst_n99) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U322 ( .A(
        wrap_act_buffer_inst_act_if_inst_n263), .B(
        wrap_act_buffer_inst_act_if_inst_n235), .S(
        wrap_act_buffer_inst_act_if_inst_n309), .Z(
        wrap_act_buffer_inst_act_if_inst_n98) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U321 ( .A(
        wrap_act_buffer_inst_act_if_inst_n191), .B(
        wrap_act_buffer_inst_act_if_inst_n183), .S(
        wrap_act_buffer_inst_act_if_inst_n309), .Z(
        wrap_act_buffer_inst_act_if_inst_n97) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U320 ( .A(
        wrap_act_buffer_inst_act_if_inst_n95), .B(
        wrap_act_buffer_inst_act_if_inst_n94), .S(
        wrap_act_buffer_inst_act_if_inst_n295), .Z(
        wrap_act_buffer_inst_act_if_inst_n96) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U319 ( .A(
        wrap_act_buffer_inst_act_if_inst_n174), .B(
        wrap_act_buffer_inst_act_if_inst_n166), .S(
        wrap_act_buffer_inst_act_if_inst_n308), .Z(
        wrap_act_buffer_inst_act_if_inst_n95) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U318 ( .A(
        wrap_act_buffer_inst_act_if_inst_n208), .B(
        wrap_act_buffer_inst_act_if_inst_n198), .S(
        wrap_act_buffer_inst_act_if_inst_n308), .Z(
        wrap_act_buffer_inst_act_if_inst_n94) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U317 ( .A(
        wrap_act_buffer_inst_act_if_inst_n92), .B(
        wrap_act_buffer_inst_act_if_inst_n91), .S(
        wrap_act_buffer_inst_act_if_inst_n295), .Z(
        wrap_act_buffer_inst_act_if_inst_n93) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U316 ( .A(
        wrap_act_buffer_inst_act_if_inst_n258), .B(
        wrap_act_buffer_inst_act_if_inst_n232), .S(
        wrap_act_buffer_inst_act_if_inst_n308), .Z(
        wrap_act_buffer_inst_act_if_inst_n92) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U315 ( .A(
        wrap_act_buffer_inst_act_if_inst_n190), .B(
        wrap_act_buffer_inst_act_if_inst_n182), .S(
        wrap_act_buffer_inst_act_if_inst_n308), .Z(
        wrap_act_buffer_inst_act_if_inst_n91) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U314 ( .A(
        wrap_act_buffer_inst_act_if_inst_n89), .B(
        wrap_act_buffer_inst_act_if_inst_n88), .S(
        wrap_act_buffer_inst_act_if_inst_n295), .Z(
        wrap_act_buffer_inst_act_if_inst_n90) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U313 ( .A(
        wrap_act_buffer_inst_act_if_inst_n173), .B(
        wrap_act_buffer_inst_act_if_inst_n165), .S(
        wrap_act_buffer_inst_act_if_inst_n308), .Z(
        wrap_act_buffer_inst_act_if_inst_n89) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U312 ( .A(
        wrap_act_buffer_inst_act_if_inst_n205), .B(
        wrap_act_buffer_inst_act_if_inst_n197), .S(
        wrap_act_buffer_inst_act_if_inst_n308), .Z(
        wrap_act_buffer_inst_act_if_inst_n88) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U311 ( .A(
        wrap_act_buffer_inst_act_if_inst_n86), .B(
        wrap_act_buffer_inst_act_if_inst_n85), .S(
        wrap_act_buffer_inst_act_if_inst_n295), .Z(
        wrap_act_buffer_inst_act_if_inst_n87) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U310 ( .A(
        wrap_act_buffer_inst_act_if_inst_n253), .B(
        wrap_act_buffer_inst_act_if_inst_n229), .S(
        wrap_act_buffer_inst_act_if_inst_n308), .Z(
        wrap_act_buffer_inst_act_if_inst_n86) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U309 ( .A(
        wrap_act_buffer_inst_act_if_inst_n189), .B(
        wrap_act_buffer_inst_act_if_inst_n181), .S(
        wrap_act_buffer_inst_act_if_inst_n308), .Z(
        wrap_act_buffer_inst_act_if_inst_n85) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U308 ( .A(
        wrap_act_buffer_inst_act_if_inst_n83), .B(
        wrap_act_buffer_inst_act_if_inst_n82), .S(
        wrap_act_buffer_inst_act_if_inst_n294), .Z(
        wrap_act_buffer_inst_act_if_inst_n84) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U307 ( .A(
        wrap_act_buffer_inst_act_if_inst_n172), .B(
        wrap_act_buffer_inst_act_if_inst_n288), .S(
        wrap_act_buffer_inst_act_if_inst_n308), .Z(
        wrap_act_buffer_inst_act_if_inst_n83) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U306 ( .A(
        wrap_act_buffer_inst_act_if_inst_n204), .B(
        wrap_act_buffer_inst_act_if_inst_n196), .S(
        wrap_act_buffer_inst_act_if_inst_n308), .Z(
        wrap_act_buffer_inst_act_if_inst_n82) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U305 ( .A(
        wrap_act_buffer_inst_act_if_inst_n80), .B(
        wrap_act_buffer_inst_act_if_inst_n79), .S(
        wrap_act_buffer_inst_act_if_inst_n294), .Z(
        wrap_act_buffer_inst_act_if_inst_n81) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U304 ( .A(
        wrap_act_buffer_inst_act_if_inst_n250), .B(
        wrap_act_buffer_inst_act_if_inst_n226), .S(
        wrap_act_buffer_inst_act_if_inst_n308), .Z(
        wrap_act_buffer_inst_act_if_inst_n80) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U303 ( .A(
        wrap_act_buffer_inst_act_if_inst_n188), .B(
        wrap_act_buffer_inst_act_if_inst_n180), .S(
        wrap_act_buffer_inst_act_if_inst_n308), .Z(
        wrap_act_buffer_inst_act_if_inst_n79) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U302 ( .A(
        wrap_act_buffer_inst_act_if_inst_n77), .B(
        wrap_act_buffer_inst_act_if_inst_n76), .S(
        wrap_act_buffer_inst_act_if_inst_n294), .Z(
        wrap_act_buffer_inst_act_if_inst_n78) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U301 ( .A(
        wrap_act_buffer_inst_act_if_inst_n171), .B(
        wrap_act_buffer_inst_act_if_inst_n283), .S(
        wrap_act_buffer_inst_act_if_inst_n307), .Z(
        wrap_act_buffer_inst_act_if_inst_n77) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U300 ( .A(
        wrap_act_buffer_inst_act_if_inst_n203), .B(
        wrap_act_buffer_inst_act_if_inst_n195), .S(
        wrap_act_buffer_inst_act_if_inst_n307), .Z(
        wrap_act_buffer_inst_act_if_inst_n76) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U299 ( .A(
        wrap_act_buffer_inst_act_if_inst_n74), .B(
        wrap_act_buffer_inst_act_if_inst_n73), .S(
        wrap_act_buffer_inst_act_if_inst_n294), .Z(
        wrap_act_buffer_inst_act_if_inst_n75) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U298 ( .A(
        wrap_act_buffer_inst_act_if_inst_n247), .B(
        wrap_act_buffer_inst_act_if_inst_n223), .S(
        wrap_act_buffer_inst_act_if_inst_n307), .Z(
        wrap_act_buffer_inst_act_if_inst_n74) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U297 ( .A(
        wrap_act_buffer_inst_act_if_inst_n187), .B(
        wrap_act_buffer_inst_act_if_inst_n179), .S(
        wrap_act_buffer_inst_act_if_inst_n307), .Z(
        wrap_act_buffer_inst_act_if_inst_n73) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U296 ( .A(
        wrap_act_buffer_inst_act_if_inst_n71), .B(
        wrap_act_buffer_inst_act_if_inst_n70), .S(
        wrap_act_buffer_inst_act_if_inst_n294), .Z(
        wrap_act_buffer_inst_act_if_inst_n72) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U295 ( .A(
        wrap_act_buffer_inst_act_if_inst_n170), .B(
        wrap_act_buffer_inst_act_if_inst_n278), .S(
        wrap_act_buffer_inst_act_if_inst_n307), .Z(
        wrap_act_buffer_inst_act_if_inst_n71) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U294 ( .A(
        wrap_act_buffer_inst_act_if_inst_n202), .B(
        wrap_act_buffer_inst_act_if_inst_n194), .S(
        wrap_act_buffer_inst_act_if_inst_n307), .Z(
        wrap_act_buffer_inst_act_if_inst_n70) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U293 ( .A(
        wrap_act_buffer_inst_act_if_inst_n68), .B(
        wrap_act_buffer_inst_act_if_inst_n67), .S(
        wrap_act_buffer_inst_act_if_inst_n294), .Z(
        wrap_act_buffer_inst_act_if_inst_n69) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U292 ( .A(
        wrap_act_buffer_inst_act_if_inst_n244), .B(
        wrap_act_buffer_inst_act_if_inst_n220), .S(
        wrap_act_buffer_inst_act_if_inst_n307), .Z(
        wrap_act_buffer_inst_act_if_inst_n68) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U291 ( .A(
        wrap_act_buffer_inst_act_if_inst_n186), .B(
        wrap_act_buffer_inst_act_if_inst_n178), .S(
        wrap_act_buffer_inst_act_if_inst_n307), .Z(
        wrap_act_buffer_inst_act_if_inst_n67) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U290 ( .A(
        wrap_act_buffer_inst_act_if_inst_n65), .B(
        wrap_act_buffer_inst_act_if_inst_n64), .S(
        wrap_act_buffer_inst_act_if_inst_n294), .Z(
        wrap_act_buffer_inst_act_if_inst_n66) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U289 ( .A(
        wrap_act_buffer_inst_act_if_inst_n169), .B(
        wrap_act_buffer_inst_act_if_inst_n273), .S(
        wrap_act_buffer_inst_act_if_inst_n307), .Z(
        wrap_act_buffer_inst_act_if_inst_n65) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U288 ( .A(
        wrap_act_buffer_inst_act_if_inst_n201), .B(
        wrap_act_buffer_inst_act_if_inst_n193), .S(
        wrap_act_buffer_inst_act_if_inst_n307), .Z(
        wrap_act_buffer_inst_act_if_inst_n64) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U287 ( .A(
        wrap_act_buffer_inst_act_if_inst_n62), .B(
        wrap_act_buffer_inst_act_if_inst_n61), .S(
        wrap_act_buffer_inst_act_if_inst_n294), .Z(
        wrap_act_buffer_inst_act_if_inst_n63) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U286 ( .A(
        wrap_act_buffer_inst_act_if_inst_n241), .B(
        wrap_act_buffer_inst_act_if_inst_n217), .S(
        wrap_act_buffer_inst_act_if_inst_n307), .Z(
        wrap_act_buffer_inst_act_if_inst_n62) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U285 ( .A(
        wrap_act_buffer_inst_act_if_inst_n185), .B(
        wrap_act_buffer_inst_act_if_inst_n177), .S(
        wrap_act_buffer_inst_act_if_inst_n307), .Z(
        wrap_act_buffer_inst_act_if_inst_n61) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U284 ( .A(
        wrap_act_buffer_inst_act_if_inst_n59), .B(
        wrap_act_buffer_inst_act_if_inst_n58), .S(
        wrap_act_buffer_inst_act_if_inst_n294), .Z(
        wrap_act_buffer_inst_act_if_inst_n60) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U283 ( .A(
        wrap_act_buffer_inst_act_if_inst_n168), .B(
        wrap_act_buffer_inst_act_if_inst_n268), .S(
        wrap_act_buffer_inst_act_if_inst_n306), .Z(
        wrap_act_buffer_inst_act_if_inst_n59) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U282 ( .A(
        wrap_act_buffer_inst_act_if_inst_n200), .B(
        wrap_act_buffer_inst_act_if_inst_n192), .S(
        wrap_act_buffer_inst_act_if_inst_n306), .Z(
        wrap_act_buffer_inst_act_if_inst_n58) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U281 ( .A(
        wrap_act_buffer_inst_act_if_inst_n56), .B(
        wrap_act_buffer_inst_act_if_inst_n55), .S(
        wrap_act_buffer_inst_act_if_inst_n294), .Z(
        wrap_act_buffer_inst_act_if_inst_n57) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U280 ( .A(
        wrap_act_buffer_inst_act_if_inst_n238), .B(
        wrap_act_buffer_inst_act_if_inst_n214), .S(
        wrap_act_buffer_inst_act_if_inst_n306), .Z(
        wrap_act_buffer_inst_act_if_inst_n56) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U279 ( .A(
        wrap_act_buffer_inst_act_if_inst_n184), .B(
        wrap_act_buffer_inst_act_if_inst_n176), .S(
        wrap_act_buffer_inst_act_if_inst_n306), .Z(
        wrap_act_buffer_inst_act_if_inst_n55) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U278 ( .A(
        wrap_act_buffer_inst_act_if_inst_n53), .B(
        wrap_act_buffer_inst_act_if_inst_n52), .S(
        wrap_act_buffer_inst_act_if_inst_n294), .Z(
        wrap_act_buffer_inst_act_if_inst_n54) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U277 ( .A(
        wrap_act_buffer_inst_act_if_inst_n167), .B(
        wrap_act_buffer_inst_act_if_inst_n263), .S(
        wrap_act_buffer_inst_act_if_inst_n306), .Z(
        wrap_act_buffer_inst_act_if_inst_n53) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U276 ( .A(
        wrap_act_buffer_inst_act_if_inst_n199), .B(
        wrap_act_buffer_inst_act_if_inst_n191), .S(
        wrap_act_buffer_inst_act_if_inst_n306), .Z(
        wrap_act_buffer_inst_act_if_inst_n52) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U275 ( .A(
        wrap_act_buffer_inst_act_if_inst_n50), .B(
        wrap_act_buffer_inst_act_if_inst_n49), .S(
        wrap_act_buffer_inst_act_if_inst_n294), .Z(
        wrap_act_buffer_inst_act_if_inst_n51) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U274 ( .A(
        wrap_act_buffer_inst_act_if_inst_n235), .B(
        wrap_act_buffer_inst_act_if_inst_n211), .S(
        wrap_act_buffer_inst_act_if_inst_n306), .Z(
        wrap_act_buffer_inst_act_if_inst_n50) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U273 ( .A(
        wrap_act_buffer_inst_act_if_inst_n183), .B(
        wrap_act_buffer_inst_act_if_inst_n175), .S(
        wrap_act_buffer_inst_act_if_inst_n306), .Z(
        wrap_act_buffer_inst_act_if_inst_n49) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U272 ( .A(
        wrap_act_buffer_inst_act_if_inst_n47), .B(
        wrap_act_buffer_inst_act_if_inst_n46), .S(
        wrap_act_buffer_inst_act_if_inst_n293), .Z(
        wrap_act_buffer_inst_act_if_inst_n48) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U271 ( .A(
        wrap_act_buffer_inst_act_if_inst_n166), .B(
        wrap_act_buffer_inst_act_if_inst_n258), .S(
        wrap_act_buffer_inst_act_if_inst_n306), .Z(
        wrap_act_buffer_inst_act_if_inst_n47) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U270 ( .A(
        wrap_act_buffer_inst_act_if_inst_n198), .B(
        wrap_act_buffer_inst_act_if_inst_n190), .S(
        wrap_act_buffer_inst_act_if_inst_n306), .Z(
        wrap_act_buffer_inst_act_if_inst_n46) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U269 ( .A(
        wrap_act_buffer_inst_act_if_inst_n44), .B(
        wrap_act_buffer_inst_act_if_inst_n43), .S(
        wrap_act_buffer_inst_act_if_inst_n293), .Z(
        wrap_act_buffer_inst_act_if_inst_n45) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U268 ( .A(
        wrap_act_buffer_inst_act_if_inst_n232), .B(
        wrap_act_buffer_inst_act_if_inst_n208), .S(
        wrap_act_buffer_inst_act_if_inst_n306), .Z(
        wrap_act_buffer_inst_act_if_inst_n44) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U267 ( .A(
        wrap_act_buffer_inst_act_if_inst_n182), .B(
        wrap_act_buffer_inst_act_if_inst_n174), .S(
        wrap_act_buffer_inst_act_if_inst_n306), .Z(
        wrap_act_buffer_inst_act_if_inst_n43) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U266 ( .A(
        wrap_act_buffer_inst_act_if_inst_n41), .B(
        wrap_act_buffer_inst_act_if_inst_n40), .S(
        wrap_act_buffer_inst_act_if_inst_n293), .Z(
        wrap_act_buffer_inst_act_if_inst_n42) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U265 ( .A(
        wrap_act_buffer_inst_act_if_inst_n165), .B(
        wrap_act_buffer_inst_act_if_inst_n253), .S(
        wrap_act_buffer_inst_act_if_inst_n305), .Z(
        wrap_act_buffer_inst_act_if_inst_n41) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U264 ( .A(
        wrap_act_buffer_inst_act_if_inst_n197), .B(
        wrap_act_buffer_inst_act_if_inst_n189), .S(
        wrap_act_buffer_inst_act_if_inst_n305), .Z(
        wrap_act_buffer_inst_act_if_inst_n40) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U263 ( .A(
        wrap_act_buffer_inst_act_if_inst_n2), .B(
        wrap_act_buffer_inst_act_if_inst_n1), .S(
        wrap_act_buffer_inst_act_if_inst_n293), .Z(
        wrap_act_buffer_inst_act_if_inst_n39) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U262 ( .A(
        wrap_act_buffer_inst_act_if_inst_n229), .B(
        wrap_act_buffer_inst_act_if_inst_n205), .S(
        wrap_act_buffer_inst_act_if_inst_n305), .Z(
        wrap_act_buffer_inst_act_if_inst_n2) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U261 ( .A(
        wrap_act_buffer_inst_act_if_inst_n181), .B(
        wrap_act_buffer_inst_act_if_inst_n173), .S(
        wrap_act_buffer_inst_act_if_inst_n305), .Z(
        wrap_act_buffer_inst_act_if_inst_n1) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U260 ( .A(
        wrap_act_buffer_inst_act_if_inst_n289), .B(
        wrap_act_buffer_inst_act_if_inst_n228), .S(
        wrap_act_buffer_inst_act_if_inst_n304), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data1[7]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U259 ( .A(
        wrap_act_buffer_inst_act_if_inst_n284), .B(
        wrap_act_buffer_inst_act_if_inst_n225), .S(
        wrap_act_buffer_inst_act_if_inst_n304), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data1[6]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U258 ( .A(
        wrap_act_buffer_inst_act_if_inst_n279), .B(
        wrap_act_buffer_inst_act_if_inst_n222), .S(
        wrap_act_buffer_inst_act_if_inst_n304), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data1[5]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U257 ( .A(
        wrap_act_buffer_inst_act_if_inst_n274), .B(
        wrap_act_buffer_inst_act_if_inst_n219), .S(
        wrap_act_buffer_inst_act_if_inst_n304), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data1[4]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U256 ( .A(
        wrap_act_buffer_inst_act_if_inst_n269), .B(
        wrap_act_buffer_inst_act_if_inst_n216), .S(
        wrap_act_buffer_inst_act_if_inst_n304), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data1[3]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U255 ( .A(
        wrap_act_buffer_inst_act_if_inst_n264), .B(
        wrap_act_buffer_inst_act_if_inst_n213), .S(
        wrap_act_buffer_inst_act_if_inst_n304), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data1[2]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U254 ( .A(
        wrap_act_buffer_inst_act_if_inst_n259), .B(
        wrap_act_buffer_inst_act_if_inst_n210), .S(
        wrap_act_buffer_inst_act_if_inst_n304), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data1[1]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U253 ( .A(
        wrap_act_buffer_inst_act_if_inst_n254), .B(
        wrap_act_buffer_inst_act_if_inst_n207), .S(
        wrap_act_buffer_inst_act_if_inst_n304), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data1[0]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U252 ( .A(
        wrap_act_buffer_inst_act_if_inst_n251), .B(
        wrap_act_buffer_inst_act_if_inst_n292), .S(
        wrap_act_buffer_inst_act_if_inst_n304), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data2[7]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U251 ( .A(
        wrap_act_buffer_inst_act_if_inst_n248), .B(
        wrap_act_buffer_inst_act_if_inst_n287), .S(
        wrap_act_buffer_inst_act_if_inst_n304), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data2[6]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U250 ( .A(
        wrap_act_buffer_inst_act_if_inst_n245), .B(
        wrap_act_buffer_inst_act_if_inst_n282), .S(
        wrap_act_buffer_inst_act_if_inst_n304), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data2[5]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U249 ( .A(
        wrap_act_buffer_inst_act_if_inst_n242), .B(
        wrap_act_buffer_inst_act_if_inst_n277), .S(
        wrap_act_buffer_inst_act_if_inst_n304), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data2[4]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U248 ( .A(
        wrap_act_buffer_inst_act_if_inst_n239), .B(
        wrap_act_buffer_inst_act_if_inst_n272), .S(
        wrap_act_buffer_inst_act_if_inst_n303), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data2[3]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U247 ( .A(
        wrap_act_buffer_inst_act_if_inst_n236), .B(
        wrap_act_buffer_inst_act_if_inst_n267), .S(
        wrap_act_buffer_inst_act_if_inst_n303), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data2[2]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U246 ( .A(
        wrap_act_buffer_inst_act_if_inst_n233), .B(
        wrap_act_buffer_inst_act_if_inst_n262), .S(
        wrap_act_buffer_inst_act_if_inst_n303), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data2[1]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U245 ( .A(
        wrap_act_buffer_inst_act_if_inst_n230), .B(
        wrap_act_buffer_inst_act_if_inst_n257), .S(
        wrap_act_buffer_inst_act_if_inst_n303), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data2[0]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U244 ( .A(
        wrap_act_buffer_inst_act_if_inst_n228), .B(
        wrap_act_buffer_inst_act_if_inst_n290), .S(
        wrap_act_buffer_inst_act_if_inst_n303), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data3[7]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U243 ( .A(
        wrap_act_buffer_inst_act_if_inst_n225), .B(
        wrap_act_buffer_inst_act_if_inst_n285), .S(
        wrap_act_buffer_inst_act_if_inst_n303), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data3[6]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U242 ( .A(
        wrap_act_buffer_inst_act_if_inst_n222), .B(
        wrap_act_buffer_inst_act_if_inst_n280), .S(
        wrap_act_buffer_inst_act_if_inst_n303), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data3[5]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U241 ( .A(
        wrap_act_buffer_inst_act_if_inst_n219), .B(
        wrap_act_buffer_inst_act_if_inst_n275), .S(
        wrap_act_buffer_inst_act_if_inst_n303), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data3[4]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U240 ( .A(
        wrap_act_buffer_inst_act_if_inst_n216), .B(
        wrap_act_buffer_inst_act_if_inst_n270), .S(
        wrap_act_buffer_inst_act_if_inst_n303), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data3[3]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U239 ( .A(
        wrap_act_buffer_inst_act_if_inst_n213), .B(
        wrap_act_buffer_inst_act_if_inst_n265), .S(
        wrap_act_buffer_inst_act_if_inst_n303), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data3[2]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U238 ( .A(
        wrap_act_buffer_inst_act_if_inst_n210), .B(
        wrap_act_buffer_inst_act_if_inst_n260), .S(
        wrap_act_buffer_inst_act_if_inst_n303), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data3[1]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U237 ( .A(
        wrap_act_buffer_inst_act_if_inst_n207), .B(
        wrap_act_buffer_inst_act_if_inst_n255), .S(
        wrap_act_buffer_inst_act_if_inst_n303), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data3[0]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U236 ( .A(
        wrap_act_buffer_inst_act_if_inst_n292), .B(
        wrap_act_buffer_inst_act_if_inst_n252), .S(
        wrap_act_buffer_inst_act_if_inst_n302), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data4[7]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U235 ( .A(
        wrap_act_buffer_inst_act_if_inst_n287), .B(
        wrap_act_buffer_inst_act_if_inst_n249), .S(
        wrap_act_buffer_inst_act_if_inst_n302), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data4[6]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U234 ( .A(
        wrap_act_buffer_inst_act_if_inst_n282), .B(
        wrap_act_buffer_inst_act_if_inst_n246), .S(
        wrap_act_buffer_inst_act_if_inst_n302), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data4[5]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U233 ( .A(
        wrap_act_buffer_inst_act_if_inst_n277), .B(
        wrap_act_buffer_inst_act_if_inst_n243), .S(
        wrap_act_buffer_inst_act_if_inst_n302), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data4[4]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U232 ( .A(
        wrap_act_buffer_inst_act_if_inst_n272), .B(
        wrap_act_buffer_inst_act_if_inst_n240), .S(
        wrap_act_buffer_inst_act_if_inst_n302), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data4[3]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U231 ( .A(
        wrap_act_buffer_inst_act_if_inst_n267), .B(
        wrap_act_buffer_inst_act_if_inst_n237), .S(
        wrap_act_buffer_inst_act_if_inst_n302), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data4[2]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U230 ( .A(
        wrap_act_buffer_inst_act_if_inst_n262), .B(
        wrap_act_buffer_inst_act_if_inst_n234), .S(
        wrap_act_buffer_inst_act_if_inst_n302), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data4[1]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U229 ( .A(
        wrap_act_buffer_inst_act_if_inst_n257), .B(
        wrap_act_buffer_inst_act_if_inst_n231), .S(
        wrap_act_buffer_inst_act_if_inst_n302), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data4[0]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U228 ( .A(
        wrap_act_buffer_inst_act_if_inst_n290), .B(
        wrap_act_buffer_inst_act_if_inst_n227), .S(
        wrap_act_buffer_inst_act_if_inst_n302), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data5[7]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U227 ( .A(
        wrap_act_buffer_inst_act_if_inst_n285), .B(
        wrap_act_buffer_inst_act_if_inst_n224), .S(
        wrap_act_buffer_inst_act_if_inst_n302), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data5[6]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U226 ( .A(
        wrap_act_buffer_inst_act_if_inst_n280), .B(
        wrap_act_buffer_inst_act_if_inst_n221), .S(
        wrap_act_buffer_inst_act_if_inst_n302), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data5[5]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U225 ( .A(
        wrap_act_buffer_inst_act_if_inst_n275), .B(
        wrap_act_buffer_inst_act_if_inst_n218), .S(
        wrap_act_buffer_inst_act_if_inst_n302), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data5[4]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U224 ( .A(
        wrap_act_buffer_inst_act_if_inst_n270), .B(
        wrap_act_buffer_inst_act_if_inst_n215), .S(
        wrap_act_buffer_inst_act_if_inst_n301), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data5[3]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U223 ( .A(
        wrap_act_buffer_inst_act_if_inst_n265), .B(
        wrap_act_buffer_inst_act_if_inst_n212), .S(
        wrap_act_buffer_inst_act_if_inst_n301), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data5[2]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U222 ( .A(
        wrap_act_buffer_inst_act_if_inst_n260), .B(
        wrap_act_buffer_inst_act_if_inst_n209), .S(
        wrap_act_buffer_inst_act_if_inst_n301), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data5[1]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U221 ( .A(
        wrap_act_buffer_inst_act_if_inst_n255), .B(
        wrap_act_buffer_inst_act_if_inst_n206), .S(
        wrap_act_buffer_inst_act_if_inst_n301), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data5[0]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U220 ( .A(
        wrap_act_buffer_inst_act_if_inst_n252), .B(
        wrap_act_buffer_inst_act_if_inst_n291), .S(
        wrap_act_buffer_inst_act_if_inst_n301), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data6[7]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U219 ( .A(
        wrap_act_buffer_inst_act_if_inst_n249), .B(
        wrap_act_buffer_inst_act_if_inst_n286), .S(
        wrap_act_buffer_inst_act_if_inst_n301), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data6[6]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U218 ( .A(
        wrap_act_buffer_inst_act_if_inst_n246), .B(
        wrap_act_buffer_inst_act_if_inst_n281), .S(
        wrap_act_buffer_inst_act_if_inst_n301), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data6[5]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U217 ( .A(
        wrap_act_buffer_inst_act_if_inst_n243), .B(
        wrap_act_buffer_inst_act_if_inst_n276), .S(
        wrap_act_buffer_inst_act_if_inst_n301), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data6[4]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U216 ( .A(
        wrap_act_buffer_inst_act_if_inst_n240), .B(
        wrap_act_buffer_inst_act_if_inst_n271), .S(
        wrap_act_buffer_inst_act_if_inst_n301), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data6[3]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U215 ( .A(
        wrap_act_buffer_inst_act_if_inst_n237), .B(
        wrap_act_buffer_inst_act_if_inst_n266), .S(
        wrap_act_buffer_inst_act_if_inst_n301), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data6[2]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U214 ( .A(
        wrap_act_buffer_inst_act_if_inst_n234), .B(
        wrap_act_buffer_inst_act_if_inst_n261), .S(
        wrap_act_buffer_inst_act_if_inst_n301), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data6[1]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U213 ( .A(
        wrap_act_buffer_inst_act_if_inst_n231), .B(
        wrap_act_buffer_inst_act_if_inst_n256), .S(
        wrap_act_buffer_inst_act_if_inst_n301), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data6[0]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U212 ( .A(
        wrap_act_buffer_inst_act_if_inst_n227), .B(
        wrap_act_buffer_inst_act_if_inst_n289), .S(
        wrap_act_buffer_inst_act_if_inst_n300), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data7[7]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U211 ( .A(
        wrap_act_buffer_inst_act_if_inst_n224), .B(
        wrap_act_buffer_inst_act_if_inst_n284), .S(
        wrap_act_buffer_inst_act_if_inst_n300), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data7[6]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U210 ( .A(
        wrap_act_buffer_inst_act_if_inst_n221), .B(
        wrap_act_buffer_inst_act_if_inst_n279), .S(
        wrap_act_buffer_inst_act_if_inst_n300), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data7[5]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U209 ( .A(
        wrap_act_buffer_inst_act_if_inst_n218), .B(
        wrap_act_buffer_inst_act_if_inst_n274), .S(
        wrap_act_buffer_inst_act_if_inst_n300), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data7[4]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U208 ( .A(
        wrap_act_buffer_inst_act_if_inst_n215), .B(
        wrap_act_buffer_inst_act_if_inst_n269), .S(
        wrap_act_buffer_inst_act_if_inst_n300), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data7[3]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U207 ( .A(
        wrap_act_buffer_inst_act_if_inst_n212), .B(
        wrap_act_buffer_inst_act_if_inst_n264), .S(
        wrap_act_buffer_inst_act_if_inst_n300), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data7[2]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U206 ( .A(
        wrap_act_buffer_inst_act_if_inst_n209), .B(
        wrap_act_buffer_inst_act_if_inst_n259), .S(
        wrap_act_buffer_inst_act_if_inst_n300), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data7[1]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U205 ( .A(
        wrap_act_buffer_inst_act_if_inst_n206), .B(
        wrap_act_buffer_inst_act_if_inst_n254), .S(
        wrap_act_buffer_inst_act_if_inst_n300), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data7[0]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U204 ( .A(
        wrap_act_buffer_inst_act_if_inst_n291), .B(
        wrap_act_buffer_inst_act_if_inst_n251), .S(
        wrap_act_buffer_inst_act_if_inst_n300), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data8[7]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U203 ( .A(
        wrap_act_buffer_inst_act_if_inst_n286), .B(
        wrap_act_buffer_inst_act_if_inst_n248), .S(
        wrap_act_buffer_inst_act_if_inst_n300), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data8[6]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U202 ( .A(
        wrap_act_buffer_inst_act_if_inst_n281), .B(
        wrap_act_buffer_inst_act_if_inst_n245), .S(
        wrap_act_buffer_inst_act_if_inst_n300), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data8[5]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U201 ( .A(
        wrap_act_buffer_inst_act_if_inst_n276), .B(
        wrap_act_buffer_inst_act_if_inst_n242), .S(
        wrap_act_buffer_inst_act_if_inst_n300), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data8[4]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U200 ( .A(
        wrap_act_buffer_inst_act_if_inst_n271), .B(
        wrap_act_buffer_inst_act_if_inst_n239), .S(
        wrap_act_buffer_inst_act_if_inst_n299), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data8[3]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U199 ( .A(
        wrap_act_buffer_inst_act_if_inst_n266), .B(
        wrap_act_buffer_inst_act_if_inst_n236), .S(
        wrap_act_buffer_inst_act_if_inst_n299), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data8[2]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U198 ( .A(
        wrap_act_buffer_inst_act_if_inst_n261), .B(
        wrap_act_buffer_inst_act_if_inst_n233), .S(
        wrap_act_buffer_inst_act_if_inst_n299), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data8[1]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U197 ( .A(
        wrap_act_buffer_inst_act_if_inst_n256), .B(
        wrap_act_buffer_inst_act_if_inst_n230), .S(
        wrap_act_buffer_inst_act_if_inst_n299), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data8[0]) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U196 ( .A(1'b0), .ZN(
        wrap_act_buffer_inst_act_if_inst_n311) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U195 ( .A(ps_int_hmode_cnt[1]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n312) );
  BUF_X1 wrap_act_buffer_inst_act_if_inst_U194 ( .A(int_L1_ptr[1]), .Z(
        wrap_act_buffer_inst_act_if_inst_n304) );
  BUF_X1 wrap_act_buffer_inst_act_if_inst_U193 ( .A(int_L1_ptr[1]), .Z(
        wrap_act_buffer_inst_act_if_inst_n303) );
  BUF_X1 wrap_act_buffer_inst_act_if_inst_U192 ( .A(int_L1_ptr[1]), .Z(
        wrap_act_buffer_inst_act_if_inst_n302) );
  BUF_X1 wrap_act_buffer_inst_act_if_inst_U191 ( .A(int_L1_ptr[1]), .Z(
        wrap_act_buffer_inst_act_if_inst_n301) );
  BUF_X1 wrap_act_buffer_inst_act_if_inst_U190 ( .A(int_L1_ptr[1]), .Z(
        wrap_act_buffer_inst_act_if_inst_n300) );
  BUF_X1 wrap_act_buffer_inst_act_if_inst_U189 ( .A(int_L1_ptr[2]), .Z(
        wrap_act_buffer_inst_act_if_inst_n295) );
  BUF_X1 wrap_act_buffer_inst_act_if_inst_U188 ( .A(int_L1_ptr[2]), .Z(
        wrap_act_buffer_inst_act_if_inst_n298) );
  BUF_X1 wrap_act_buffer_inst_act_if_inst_U187 ( .A(int_L1_ptr[2]), .Z(
        wrap_act_buffer_inst_act_if_inst_n296) );
  BUF_X1 wrap_act_buffer_inst_act_if_inst_U186 ( .A(int_L1_ptr[2]), .Z(
        wrap_act_buffer_inst_act_if_inst_n294) );
  BUF_X1 wrap_act_buffer_inst_act_if_inst_U185 ( .A(int_L1_ptr[2]), .Z(
        wrap_act_buffer_inst_act_if_inst_n297) );
  BUF_X1 wrap_act_buffer_inst_act_if_inst_U184 ( .A(int_L1_ptr[0]), .Z(
        wrap_act_buffer_inst_act_if_inst_n309) );
  BUF_X1 wrap_act_buffer_inst_act_if_inst_U183 ( .A(int_L1_ptr[0]), .Z(
        wrap_act_buffer_inst_act_if_inst_n310) );
  BUF_X1 wrap_act_buffer_inst_act_if_inst_U182 ( .A(int_L1_ptr[0]), .Z(
        wrap_act_buffer_inst_act_if_inst_n308) );
  BUF_X1 wrap_act_buffer_inst_act_if_inst_U181 ( .A(int_L1_ptr[0]), .Z(
        wrap_act_buffer_inst_act_if_inst_n306) );
  BUF_X1 wrap_act_buffer_inst_act_if_inst_U180 ( .A(int_L1_ptr[0]), .Z(
        wrap_act_buffer_inst_act_if_inst_n307) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U179 ( .A(
        wrap_act_buffer_inst_int_i_data_if1[3]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n268) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U178 ( .A(
        wrap_act_buffer_inst_int_i_data_if2[3]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n238) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U177 ( .A(
        wrap_act_buffer_inst_int_i_data_if5[3]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n192) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U176 ( .A(
        wrap_act_buffer_inst_int_i_data_if3[3]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n214) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U175 ( .A(
        wrap_act_buffer_inst_int_i_data_if4[3]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n200) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U174 ( .A(
        wrap_act_buffer_inst_int_i_data_if1[5]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n278) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U173 ( .A(
        wrap_act_buffer_inst_int_i_data_if2[5]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n244) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U172 ( .A(
        wrap_act_buffer_inst_int_i_data_if3[5]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n220) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U171 ( .A(
        wrap_act_buffer_inst_int_i_data_if4[5]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n202) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U170 ( .A(
        wrap_act_buffer_inst_int_i_data_if1[7]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n288) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U169 ( .A(
        wrap_act_buffer_inst_int_i_data_if2[7]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n250) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U168 ( .A(
        wrap_act_buffer_inst_int_i_data_if3[7]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n226) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U167 ( .A(
        wrap_act_buffer_inst_int_i_data_if4[7]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n204) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U166 ( .A(
        wrap_act_buffer_inst_int_i_data_if1[1]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n258) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U165 ( .A(
        wrap_act_buffer_inst_int_i_data_if2[1]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n232) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U164 ( .A(
        wrap_act_buffer_inst_int_i_data_if5[1]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n190) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U163 ( .A(
        wrap_act_buffer_inst_int_i_data_if3[1]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n208) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U162 ( .A(
        wrap_act_buffer_inst_int_i_data_if4[1]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n198) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U161 ( .A(
        wrap_act_buffer_inst_int_i_data_if1[2]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n263) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U160 ( .A(
        wrap_act_buffer_inst_int_i_data_if2[2]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n235) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U159 ( .A(
        wrap_act_buffer_inst_int_i_data_if5[2]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n191) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U158 ( .A(
        wrap_act_buffer_inst_int_i_data_if3[2]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n211) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U157 ( .A(
        wrap_act_buffer_inst_int_i_data_if4[2]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n199) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U156 ( .A(
        wrap_act_buffer_inst_int_i_data_if1[4]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n273) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U155 ( .A(
        wrap_act_buffer_inst_int_i_data_if2[4]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n241) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U154 ( .A(
        wrap_act_buffer_inst_int_i_data_if3[4]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n217) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U153 ( .A(
        wrap_act_buffer_inst_int_i_data_if4[4]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n201) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U152 ( .A(
        wrap_act_buffer_inst_int_i_data_if1[6]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n283) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U151 ( .A(
        wrap_act_buffer_inst_int_i_data_if2[6]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n247) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U150 ( .A(
        wrap_act_buffer_inst_int_i_data_if3[6]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n223) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U149 ( .A(
        wrap_act_buffer_inst_int_i_data_if4[6]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n203) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U148 ( .A(
        wrap_act_buffer_inst_int_i_data_if1[0]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n253) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U147 ( .A(
        wrap_act_buffer_inst_int_i_data_if2[0]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n229) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U146 ( .A(
        wrap_act_buffer_inst_int_i_data_if5[0]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n189) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U145 ( .A(
        wrap_act_buffer_inst_int_i_data_if4[0]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n197) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U144 ( .A(
        wrap_act_buffer_inst_int_i_data_if3[0]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n205) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U143 ( .A(
        wrap_act_buffer_inst_int_i_data_if6[3]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n184) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U142 ( .A(
        wrap_act_buffer_inst_int_i_data_if7[3]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n176) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U141 ( .A(
        wrap_act_buffer_inst_int_i_data_if8[3]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n168) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U140 ( .A(
        wrap_act_buffer_inst_int_i_data_if5[5]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n194) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U139 ( .A(
        wrap_act_buffer_inst_int_i_data_if6[5]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n186) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U138 ( .A(
        wrap_act_buffer_inst_int_i_data_if8[5]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n170) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U137 ( .A(
        wrap_act_buffer_inst_int_i_data_if7[5]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n178) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U136 ( .A(
        wrap_act_buffer_inst_int_i_data_if5[7]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n196) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U135 ( .A(
        wrap_act_buffer_inst_int_i_data_if6[7]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n188) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U134 ( .A(
        wrap_act_buffer_inst_int_i_data_if8[7]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n172) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U133 ( .A(
        wrap_act_buffer_inst_int_i_data_if7[7]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n180) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U132 ( .A(
        wrap_act_buffer_inst_int_i_data_if6[1]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n182) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U131 ( .A(
        wrap_act_buffer_inst_int_i_data_if8[1]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n166) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U130 ( .A(
        wrap_act_buffer_inst_int_i_data_if7[1]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n174) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U129 ( .A(
        wrap_act_buffer_inst_int_i_data_if6[2]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n183) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U128 ( .A(
        wrap_act_buffer_inst_int_i_data_if7[2]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n175) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U127 ( .A(
        wrap_act_buffer_inst_int_i_data_if8[2]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n167) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U126 ( .A(
        wrap_act_buffer_inst_int_i_data_if5[4]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n193) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U125 ( .A(
        wrap_act_buffer_inst_int_i_data_if6[4]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n185) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U124 ( .A(
        wrap_act_buffer_inst_int_i_data_if8[4]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n169) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U123 ( .A(
        wrap_act_buffer_inst_int_i_data_if7[4]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n177) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U122 ( .A(
        wrap_act_buffer_inst_int_i_data_if5[6]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n195) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U121 ( .A(
        wrap_act_buffer_inst_int_i_data_if6[6]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n187) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U120 ( .A(
        wrap_act_buffer_inst_int_i_data_if8[6]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n171) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U119 ( .A(
        wrap_act_buffer_inst_int_i_data_if7[6]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n179) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U118 ( .A(
        wrap_act_buffer_inst_int_i_data_if6[0]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n181) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U117 ( .A(
        wrap_act_buffer_inst_int_i_data_if8[0]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n165) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U116 ( .A(
        wrap_act_buffer_inst_int_i_data_if7[0]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n173) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U115 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data8[6]), .A2(
        wrap_act_buffer_inst_act_if_inst_n5), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data8[0]), .B2(
        wrap_act_buffer_inst_act_if_inst_n6), .ZN(
        wrap_act_buffer_inst_act_if_inst_n10) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U114 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data8[2]), .A2(
        wrap_act_buffer_inst_act_if_inst_n7), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data8[4]), .B2(
        wrap_act_buffer_inst_act_if_inst_n8), .ZN(
        wrap_act_buffer_inst_act_if_inst_n9) );
  NAND2_X1 wrap_act_buffer_inst_act_if_inst_U113 ( .A1(
        wrap_act_buffer_inst_act_if_inst_n9), .A2(
        wrap_act_buffer_inst_act_if_inst_n10), .ZN(int_i_data_h_npu[0]) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U112 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data8[7]), .A2(
        wrap_act_buffer_inst_act_if_inst_n5), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data8[1]), .B2(
        wrap_act_buffer_inst_act_if_inst_n6), .ZN(
        wrap_act_buffer_inst_act_if_inst_n4) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U111 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data8[3]), .A2(
        wrap_act_buffer_inst_act_if_inst_n7), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data8[5]), .B2(
        wrap_act_buffer_inst_act_if_inst_n8), .ZN(
        wrap_act_buffer_inst_act_if_inst_n3) );
  NAND2_X1 wrap_act_buffer_inst_act_if_inst_U110 ( .A1(
        wrap_act_buffer_inst_act_if_inst_n3), .A2(
        wrap_act_buffer_inst_act_if_inst_n4), .ZN(int_i_data_h_npu[1]) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U109 ( .A(
        wrap_act_buffer_inst_act_if_inst_n105), .ZN(
        wrap_act_buffer_inst_act_if_inst_n269) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U108 ( .A(
        wrap_act_buffer_inst_act_if_inst_n160), .ZN(
        wrap_act_buffer_inst_act_if_inst_n216) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U107 ( .A(
        wrap_act_buffer_inst_act_if_inst_n117), .ZN(
        wrap_act_buffer_inst_act_if_inst_n279) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U106 ( .A(
        wrap_act_buffer_inst_act_if_inst_n162), .ZN(
        wrap_act_buffer_inst_act_if_inst_n222) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U105 ( .A(
        wrap_act_buffer_inst_act_if_inst_n129), .ZN(
        wrap_act_buffer_inst_act_if_inst_n289) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U104 ( .A(
        wrap_act_buffer_inst_act_if_inst_n164), .ZN(
        wrap_act_buffer_inst_act_if_inst_n228) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U103 ( .A(
        wrap_act_buffer_inst_act_if_inst_n93), .ZN(
        wrap_act_buffer_inst_act_if_inst_n259) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U102 ( .A(
        wrap_act_buffer_inst_act_if_inst_n158), .ZN(
        wrap_act_buffer_inst_act_if_inst_n210) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U101 ( .A(
        wrap_act_buffer_inst_act_if_inst_n99), .ZN(
        wrap_act_buffer_inst_act_if_inst_n264) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U100 ( .A(
        wrap_act_buffer_inst_act_if_inst_n159), .ZN(
        wrap_act_buffer_inst_act_if_inst_n213) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U99 ( .A(
        wrap_act_buffer_inst_act_if_inst_n111), .ZN(
        wrap_act_buffer_inst_act_if_inst_n274) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U98 ( .A(
        wrap_act_buffer_inst_act_if_inst_n161), .ZN(
        wrap_act_buffer_inst_act_if_inst_n219) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U97 ( .A(
        wrap_act_buffer_inst_act_if_inst_n123), .ZN(
        wrap_act_buffer_inst_act_if_inst_n284) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U96 ( .A(
        wrap_act_buffer_inst_act_if_inst_n163), .ZN(
        wrap_act_buffer_inst_act_if_inst_n225) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U95 ( .A(
        wrap_act_buffer_inst_act_if_inst_n87), .ZN(
        wrap_act_buffer_inst_act_if_inst_n254) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U94 ( .A(
        wrap_act_buffer_inst_act_if_inst_n157), .ZN(
        wrap_act_buffer_inst_act_if_inst_n207) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U93 ( .A(
        wrap_act_buffer_inst_act_if_inst_n57), .ZN(
        wrap_act_buffer_inst_act_if_inst_n239) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U92 ( .A(
        wrap_act_buffer_inst_act_if_inst_n152), .ZN(
        wrap_act_buffer_inst_act_if_inst_n272) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U91 ( .A(
        wrap_act_buffer_inst_act_if_inst_n69), .ZN(
        wrap_act_buffer_inst_act_if_inst_n245) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U90 ( .A(
        wrap_act_buffer_inst_act_if_inst_n154), .ZN(
        wrap_act_buffer_inst_act_if_inst_n282) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U89 ( .A(
        wrap_act_buffer_inst_act_if_inst_n81), .ZN(
        wrap_act_buffer_inst_act_if_inst_n251) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U88 ( .A(
        wrap_act_buffer_inst_act_if_inst_n156), .ZN(
        wrap_act_buffer_inst_act_if_inst_n292) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U87 ( .A(
        wrap_act_buffer_inst_act_if_inst_n45), .ZN(
        wrap_act_buffer_inst_act_if_inst_n233) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U86 ( .A(
        wrap_act_buffer_inst_act_if_inst_n150), .ZN(
        wrap_act_buffer_inst_act_if_inst_n262) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U85 ( .A(
        wrap_act_buffer_inst_act_if_inst_n51), .ZN(
        wrap_act_buffer_inst_act_if_inst_n236) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U84 ( .A(
        wrap_act_buffer_inst_act_if_inst_n151), .ZN(
        wrap_act_buffer_inst_act_if_inst_n267) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U83 ( .A(
        wrap_act_buffer_inst_act_if_inst_n63), .ZN(
        wrap_act_buffer_inst_act_if_inst_n242) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U82 ( .A(
        wrap_act_buffer_inst_act_if_inst_n153), .ZN(
        wrap_act_buffer_inst_act_if_inst_n277) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U81 ( .A(
        wrap_act_buffer_inst_act_if_inst_n75), .ZN(
        wrap_act_buffer_inst_act_if_inst_n248) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U80 ( .A(
        wrap_act_buffer_inst_act_if_inst_n155), .ZN(
        wrap_act_buffer_inst_act_if_inst_n287) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U79 ( .A(
        wrap_act_buffer_inst_act_if_inst_n39), .ZN(
        wrap_act_buffer_inst_act_if_inst_n230) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U78 ( .A(
        wrap_act_buffer_inst_act_if_inst_n149), .ZN(
        wrap_act_buffer_inst_act_if_inst_n257) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U77 ( .A(
        wrap_act_buffer_inst_act_if_inst_n144), .ZN(
        wrap_act_buffer_inst_act_if_inst_n270) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U76 ( .A(
        wrap_act_buffer_inst_act_if_inst_n146), .ZN(
        wrap_act_buffer_inst_act_if_inst_n280) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U75 ( .A(
        wrap_act_buffer_inst_act_if_inst_n148), .ZN(
        wrap_act_buffer_inst_act_if_inst_n290) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U74 ( .A(
        wrap_act_buffer_inst_act_if_inst_n142), .ZN(
        wrap_act_buffer_inst_act_if_inst_n260) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U73 ( .A(
        wrap_act_buffer_inst_act_if_inst_n143), .ZN(
        wrap_act_buffer_inst_act_if_inst_n265) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U72 ( .A(
        wrap_act_buffer_inst_act_if_inst_n145), .ZN(
        wrap_act_buffer_inst_act_if_inst_n275) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U71 ( .A(
        wrap_act_buffer_inst_act_if_inst_n147), .ZN(
        wrap_act_buffer_inst_act_if_inst_n285) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U70 ( .A(
        wrap_act_buffer_inst_act_if_inst_n141), .ZN(
        wrap_act_buffer_inst_act_if_inst_n255) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U69 ( .A(
        wrap_act_buffer_inst_act_if_inst_n136), .ZN(
        wrap_act_buffer_inst_act_if_inst_n240) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U68 ( .A(
        wrap_act_buffer_inst_act_if_inst_n138), .ZN(
        wrap_act_buffer_inst_act_if_inst_n246) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U67 ( .A(
        wrap_act_buffer_inst_act_if_inst_n140), .ZN(
        wrap_act_buffer_inst_act_if_inst_n252) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U66 ( .A(
        wrap_act_buffer_inst_act_if_inst_n134), .ZN(
        wrap_act_buffer_inst_act_if_inst_n234) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U65 ( .A(
        wrap_act_buffer_inst_act_if_inst_n135), .ZN(
        wrap_act_buffer_inst_act_if_inst_n237) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U64 ( .A(
        wrap_act_buffer_inst_act_if_inst_n137), .ZN(
        wrap_act_buffer_inst_act_if_inst_n243) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U63 ( .A(
        wrap_act_buffer_inst_act_if_inst_n139), .ZN(
        wrap_act_buffer_inst_act_if_inst_n249) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U62 ( .A(
        wrap_act_buffer_inst_act_if_inst_n133), .ZN(
        wrap_act_buffer_inst_act_if_inst_n231) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U61 ( .A(
        wrap_act_buffer_inst_act_if_inst_n108), .ZN(
        wrap_act_buffer_inst_act_if_inst_n215) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U60 ( .A(
        wrap_act_buffer_inst_act_if_inst_n120), .ZN(
        wrap_act_buffer_inst_act_if_inst_n221) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U59 ( .A(
        wrap_act_buffer_inst_act_if_inst_n132), .ZN(
        wrap_act_buffer_inst_act_if_inst_n227) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U58 ( .A(
        wrap_act_buffer_inst_act_if_inst_n96), .ZN(
        wrap_act_buffer_inst_act_if_inst_n209) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U57 ( .A(
        wrap_act_buffer_inst_act_if_inst_n102), .ZN(
        wrap_act_buffer_inst_act_if_inst_n212) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U56 ( .A(
        wrap_act_buffer_inst_act_if_inst_n114), .ZN(
        wrap_act_buffer_inst_act_if_inst_n218) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U55 ( .A(
        wrap_act_buffer_inst_act_if_inst_n126), .ZN(
        wrap_act_buffer_inst_act_if_inst_n224) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U54 ( .A(
        wrap_act_buffer_inst_act_if_inst_n90), .ZN(
        wrap_act_buffer_inst_act_if_inst_n206) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U53 ( .A(
        wrap_act_buffer_inst_act_if_inst_n60), .ZN(
        wrap_act_buffer_inst_act_if_inst_n271) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U52 ( .A(
        wrap_act_buffer_inst_act_if_inst_n72), .ZN(
        wrap_act_buffer_inst_act_if_inst_n281) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U51 ( .A(
        wrap_act_buffer_inst_act_if_inst_n84), .ZN(
        wrap_act_buffer_inst_act_if_inst_n291) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U50 ( .A(
        wrap_act_buffer_inst_act_if_inst_n48), .ZN(
        wrap_act_buffer_inst_act_if_inst_n261) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U49 ( .A(
        wrap_act_buffer_inst_act_if_inst_n54), .ZN(
        wrap_act_buffer_inst_act_if_inst_n266) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U48 ( .A(
        wrap_act_buffer_inst_act_if_inst_n66), .ZN(
        wrap_act_buffer_inst_act_if_inst_n276) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U47 ( .A(
        wrap_act_buffer_inst_act_if_inst_n78), .ZN(
        wrap_act_buffer_inst_act_if_inst_n286) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U46 ( .A(
        wrap_act_buffer_inst_act_if_inst_n42), .ZN(
        wrap_act_buffer_inst_act_if_inst_n256) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U45 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data1[7]), .A2(
        wrap_act_buffer_inst_act_if_inst_n5), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data1[1]), .B2(
        wrap_act_buffer_inst_act_if_inst_n6), .ZN(
        wrap_act_buffer_inst_act_if_inst_n36) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U44 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data1[3]), .A2(
        wrap_act_buffer_inst_act_if_inst_n7), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data1[5]), .B2(
        wrap_act_buffer_inst_act_if_inst_n8), .ZN(
        wrap_act_buffer_inst_act_if_inst_n35) );
  NAND2_X1 wrap_act_buffer_inst_act_if_inst_U43 ( .A1(
        wrap_act_buffer_inst_act_if_inst_n35), .A2(
        wrap_act_buffer_inst_act_if_inst_n36), .ZN(int_i_data_h_npu[15]) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U42 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data1[6]), .A2(
        wrap_act_buffer_inst_act_if_inst_n5), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data1[0]), .B2(
        wrap_act_buffer_inst_act_if_inst_n6), .ZN(
        wrap_act_buffer_inst_act_if_inst_n38) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U41 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data1[2]), .A2(
        wrap_act_buffer_inst_act_if_inst_n7), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data1[4]), .B2(
        wrap_act_buffer_inst_act_if_inst_n8), .ZN(
        wrap_act_buffer_inst_act_if_inst_n37) );
  NAND2_X1 wrap_act_buffer_inst_act_if_inst_U40 ( .A1(
        wrap_act_buffer_inst_act_if_inst_n37), .A2(
        wrap_act_buffer_inst_act_if_inst_n38), .ZN(int_i_data_h_npu[14]) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U39 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data2[7]), .A2(
        wrap_act_buffer_inst_act_if_inst_n5), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data2[1]), .B2(
        wrap_act_buffer_inst_act_if_inst_n6), .ZN(
        wrap_act_buffer_inst_act_if_inst_n32) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U38 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data2[3]), .A2(
        wrap_act_buffer_inst_act_if_inst_n7), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data2[5]), .B2(
        wrap_act_buffer_inst_act_if_inst_n8), .ZN(
        wrap_act_buffer_inst_act_if_inst_n31) );
  NAND2_X1 wrap_act_buffer_inst_act_if_inst_U37 ( .A1(
        wrap_act_buffer_inst_act_if_inst_n31), .A2(
        wrap_act_buffer_inst_act_if_inst_n32), .ZN(int_i_data_h_npu[13]) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U36 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data2[6]), .A2(
        wrap_act_buffer_inst_act_if_inst_n5), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data2[0]), .B2(
        wrap_act_buffer_inst_act_if_inst_n6), .ZN(
        wrap_act_buffer_inst_act_if_inst_n34) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U35 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data2[2]), .A2(
        wrap_act_buffer_inst_act_if_inst_n7), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data2[4]), .B2(
        wrap_act_buffer_inst_act_if_inst_n8), .ZN(
        wrap_act_buffer_inst_act_if_inst_n33) );
  NAND2_X1 wrap_act_buffer_inst_act_if_inst_U34 ( .A1(
        wrap_act_buffer_inst_act_if_inst_n33), .A2(
        wrap_act_buffer_inst_act_if_inst_n34), .ZN(int_i_data_h_npu[12]) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U33 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data3[7]), .A2(
        wrap_act_buffer_inst_act_if_inst_n5), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data3[1]), .B2(
        wrap_act_buffer_inst_act_if_inst_n6), .ZN(
        wrap_act_buffer_inst_act_if_inst_n28) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U32 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data3[3]), .A2(
        wrap_act_buffer_inst_act_if_inst_n7), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data3[5]), .B2(
        wrap_act_buffer_inst_act_if_inst_n8), .ZN(
        wrap_act_buffer_inst_act_if_inst_n27) );
  NAND2_X1 wrap_act_buffer_inst_act_if_inst_U31 ( .A1(
        wrap_act_buffer_inst_act_if_inst_n27), .A2(
        wrap_act_buffer_inst_act_if_inst_n28), .ZN(int_i_data_h_npu[11]) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U30 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data3[6]), .A2(
        wrap_act_buffer_inst_act_if_inst_n5), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data3[0]), .B2(
        wrap_act_buffer_inst_act_if_inst_n6), .ZN(
        wrap_act_buffer_inst_act_if_inst_n30) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U29 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data3[2]), .A2(
        wrap_act_buffer_inst_act_if_inst_n7), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data3[4]), .B2(
        wrap_act_buffer_inst_act_if_inst_n8), .ZN(
        wrap_act_buffer_inst_act_if_inst_n29) );
  NAND2_X1 wrap_act_buffer_inst_act_if_inst_U28 ( .A1(
        wrap_act_buffer_inst_act_if_inst_n29), .A2(
        wrap_act_buffer_inst_act_if_inst_n30), .ZN(int_i_data_h_npu[10]) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U27 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data4[7]), .A2(
        wrap_act_buffer_inst_act_if_inst_n5), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data4[1]), .B2(
        wrap_act_buffer_inst_act_if_inst_n6), .ZN(
        wrap_act_buffer_inst_act_if_inst_n24) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U26 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data4[3]), .A2(
        wrap_act_buffer_inst_act_if_inst_n7), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data4[5]), .B2(
        wrap_act_buffer_inst_act_if_inst_n8), .ZN(
        wrap_act_buffer_inst_act_if_inst_n23) );
  NAND2_X1 wrap_act_buffer_inst_act_if_inst_U25 ( .A1(
        wrap_act_buffer_inst_act_if_inst_n23), .A2(
        wrap_act_buffer_inst_act_if_inst_n24), .ZN(int_i_data_h_npu[9]) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U24 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data4[6]), .A2(
        wrap_act_buffer_inst_act_if_inst_n5), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data4[0]), .B2(
        wrap_act_buffer_inst_act_if_inst_n6), .ZN(
        wrap_act_buffer_inst_act_if_inst_n26) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U23 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data4[2]), .A2(
        wrap_act_buffer_inst_act_if_inst_n7), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data4[4]), .B2(
        wrap_act_buffer_inst_act_if_inst_n8), .ZN(
        wrap_act_buffer_inst_act_if_inst_n25) );
  NAND2_X1 wrap_act_buffer_inst_act_if_inst_U22 ( .A1(
        wrap_act_buffer_inst_act_if_inst_n25), .A2(
        wrap_act_buffer_inst_act_if_inst_n26), .ZN(int_i_data_h_npu[8]) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U21 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data5[7]), .A2(
        wrap_act_buffer_inst_act_if_inst_n5), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data5[1]), .B2(
        wrap_act_buffer_inst_act_if_inst_n6), .ZN(
        wrap_act_buffer_inst_act_if_inst_n20) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U20 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data5[3]), .A2(
        wrap_act_buffer_inst_act_if_inst_n7), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data5[5]), .B2(
        wrap_act_buffer_inst_act_if_inst_n8), .ZN(
        wrap_act_buffer_inst_act_if_inst_n19) );
  NAND2_X1 wrap_act_buffer_inst_act_if_inst_U19 ( .A1(
        wrap_act_buffer_inst_act_if_inst_n19), .A2(
        wrap_act_buffer_inst_act_if_inst_n20), .ZN(int_i_data_h_npu[7]) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U18 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data5[6]), .A2(
        wrap_act_buffer_inst_act_if_inst_n5), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data5[0]), .B2(
        wrap_act_buffer_inst_act_if_inst_n6), .ZN(
        wrap_act_buffer_inst_act_if_inst_n22) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U17 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data5[2]), .A2(
        wrap_act_buffer_inst_act_if_inst_n7), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data5[4]), .B2(
        wrap_act_buffer_inst_act_if_inst_n8), .ZN(
        wrap_act_buffer_inst_act_if_inst_n21) );
  NAND2_X1 wrap_act_buffer_inst_act_if_inst_U16 ( .A1(
        wrap_act_buffer_inst_act_if_inst_n21), .A2(
        wrap_act_buffer_inst_act_if_inst_n22), .ZN(int_i_data_h_npu[6]) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U15 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data6[7]), .A2(
        wrap_act_buffer_inst_act_if_inst_n5), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data6[1]), .B2(
        wrap_act_buffer_inst_act_if_inst_n6), .ZN(
        wrap_act_buffer_inst_act_if_inst_n16) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U14 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data6[3]), .A2(
        wrap_act_buffer_inst_act_if_inst_n7), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data6[5]), .B2(
        wrap_act_buffer_inst_act_if_inst_n8), .ZN(
        wrap_act_buffer_inst_act_if_inst_n15) );
  NAND2_X1 wrap_act_buffer_inst_act_if_inst_U13 ( .A1(
        wrap_act_buffer_inst_act_if_inst_n15), .A2(
        wrap_act_buffer_inst_act_if_inst_n16), .ZN(int_i_data_h_npu[5]) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U12 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data6[6]), .A2(
        wrap_act_buffer_inst_act_if_inst_n5), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data6[0]), .B2(
        wrap_act_buffer_inst_act_if_inst_n6), .ZN(
        wrap_act_buffer_inst_act_if_inst_n18) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U11 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data6[2]), .A2(
        wrap_act_buffer_inst_act_if_inst_n7), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data6[4]), .B2(
        wrap_act_buffer_inst_act_if_inst_n8), .ZN(
        wrap_act_buffer_inst_act_if_inst_n17) );
  NAND2_X1 wrap_act_buffer_inst_act_if_inst_U10 ( .A1(
        wrap_act_buffer_inst_act_if_inst_n17), .A2(
        wrap_act_buffer_inst_act_if_inst_n18), .ZN(int_i_data_h_npu[4]) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U9 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data7[7]), .A2(
        wrap_act_buffer_inst_act_if_inst_n5), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data7[1]), .B2(
        wrap_act_buffer_inst_act_if_inst_n6), .ZN(
        wrap_act_buffer_inst_act_if_inst_n12) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U8 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data7[3]), .A2(
        wrap_act_buffer_inst_act_if_inst_n7), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data7[5]), .B2(
        wrap_act_buffer_inst_act_if_inst_n8), .ZN(
        wrap_act_buffer_inst_act_if_inst_n11) );
  NAND2_X1 wrap_act_buffer_inst_act_if_inst_U7 ( .A1(
        wrap_act_buffer_inst_act_if_inst_n11), .A2(
        wrap_act_buffer_inst_act_if_inst_n12), .ZN(int_i_data_h_npu[3]) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U6 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data7[6]), .A2(
        wrap_act_buffer_inst_act_if_inst_n5), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data7[0]), .B2(
        wrap_act_buffer_inst_act_if_inst_n6), .ZN(
        wrap_act_buffer_inst_act_if_inst_n14) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U5 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data7[2]), .A2(
        wrap_act_buffer_inst_act_if_inst_n7), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data7[4]), .B2(
        wrap_act_buffer_inst_act_if_inst_n8), .ZN(
        wrap_act_buffer_inst_act_if_inst_n13) );
  NAND2_X1 wrap_act_buffer_inst_act_if_inst_U4 ( .A1(
        wrap_act_buffer_inst_act_if_inst_n13), .A2(
        wrap_act_buffer_inst_act_if_inst_n14), .ZN(int_i_data_h_npu[2]) );
  AND3_X1 wrap_act_buffer_inst_act_if_inst_U3 ( .A1(
        wrap_act_buffer_inst_act_if_inst_n312), .A2(
        wrap_act_buffer_inst_act_if_inst_n311), .A3(ps_int_hmode_cnt[0]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n8) );
  AND3_X1 wrap_act_buffer_inst_act_if_inst_U2 ( .A1(ps_int_hmode_cnt[0]), .A2(
        wrap_act_buffer_inst_act_if_inst_n311), .A3(ps_int_hmode_cnt[1]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n6) );
  NOR3_X4 wrap_act_buffer_inst_act_if_inst_U1 ( .A1(
        wrap_act_buffer_inst_act_if_inst_n7), .A2(
        wrap_act_buffer_inst_act_if_inst_n8), .A3(
        wrap_act_buffer_inst_act_if_inst_n6), .ZN(
        wrap_act_buffer_inst_act_if_inst_n5) );
  CLKGATETST_X1 wrap_act_buffer_inst_clk_gate_int_i_data_v_npu_reg_latch ( 
        .CK(ck), .E(ctrl_ldh_v_n), .SE(1'b0), .GCK(
        wrap_act_buffer_inst_net4585) );
  CLKBUF_X1 npu_inst_U207 ( .A(i_weight[1]), .Z(npu_inst_n119) );
  CLKBUF_X1 npu_inst_U206 ( .A(i_weight[0]), .Z(npu_inst_n113) );
  CLKBUF_X1 npu_inst_U205 ( .A(ps_int_L0_ptr[0]), .Z(npu_inst_n72) );
  INV_X1 npu_inst_U204 ( .A(1'b0), .ZN(npu_inst_n129) );
  INV_X1 npu_inst_U203 ( .A(1'b0), .ZN(npu_inst_n128) );
  NAND2_X1 npu_inst_U202 ( .A1(npu_inst_n129), .A2(npu_inst_n128), .ZN(
        npu_inst_int_ckg[63]) );
  NAND2_X1 npu_inst_U201 ( .A1(npu_inst_n129), .A2(npu_inst_n136), .ZN(
        npu_inst_int_ckg[59]) );
  NAND2_X1 npu_inst_U200 ( .A1(npu_inst_n143), .A2(npu_inst_n128), .ZN(
        npu_inst_int_ckg[31]) );
  NAND2_X1 npu_inst_U199 ( .A1(npu_inst_n143), .A2(npu_inst_n136), .ZN(
        npu_inst_int_ckg[27]) );
  BUF_X1 npu_inst_U198 ( .A(ps_ctrl_wr_pipe), .Z(npu_inst_n5) );
  BUF_X1 npu_inst_U197 ( .A(ps_ctrl_ldh_v_n), .Z(npu_inst_n51) );
  BUF_X1 npu_inst_U196 ( .A(ps_ctrl_ldh_v_n), .Z(npu_inst_n50) );
  BUF_X1 npu_inst_U195 ( .A(ps_ctrl_en_npu), .Z(npu_inst_n66) );
  BUF_X1 npu_inst_U194 ( .A(ps_ctrl_en_npu), .Z(npu_inst_n61) );
  BUF_X1 npu_inst_U193 ( .A(ps_ctrl_en_npu), .Z(npu_inst_n62) );
  BUF_X1 npu_inst_U192 ( .A(ps_ctrl_en_npu), .Z(npu_inst_n63) );
  BUF_X1 npu_inst_U191 ( .A(ps_ctrl_en_npu), .Z(npu_inst_n64) );
  BUF_X1 npu_inst_U190 ( .A(ps_ctrl_en_npu), .Z(npu_inst_n65) );
  BUF_X1 npu_inst_U189 ( .A(i_weight[1]), .Z(npu_inst_n118) );
  BUF_X1 npu_inst_U188 ( .A(i_weight[0]), .Z(npu_inst_n112) );
  BUF_X1 npu_inst_U187 ( .A(i_weight[1]), .Z(npu_inst_n117) );
  BUF_X1 npu_inst_U186 ( .A(i_weight[0]), .Z(npu_inst_n111) );
  BUF_X1 npu_inst_U185 ( .A(i_weight[1]), .Z(npu_inst_n116) );
  BUF_X1 npu_inst_U184 ( .A(i_weight[0]), .Z(npu_inst_n110) );
  BUF_X1 npu_inst_U183 ( .A(i_weight[1]), .Z(npu_inst_n115) );
  BUF_X1 npu_inst_U182 ( .A(i_weight[0]), .Z(npu_inst_n109) );
  BUF_X1 npu_inst_U181 ( .A(i_weight[1]), .Z(npu_inst_n114) );
  BUF_X1 npu_inst_U180 ( .A(i_weight[0]), .Z(npu_inst_n108) );
  INV_X1 npu_inst_U179 ( .A(int_ckg_rmask[4]), .ZN(npu_inst_n143) );
  INV_X1 npu_inst_U178 ( .A(int_ckg_cmask[4]), .ZN(npu_inst_n136) );
  NAND2_X1 npu_inst_U177 ( .A1(npu_inst_n129), .A2(npu_inst_n130), .ZN(
        npu_inst_int_ckg[62]) );
  NAND2_X1 npu_inst_U176 ( .A1(npu_inst_n129), .A2(npu_inst_n135), .ZN(
        npu_inst_int_ckg[61]) );
  NAND2_X1 npu_inst_U175 ( .A1(npu_inst_n129), .A2(npu_inst_n132), .ZN(
        npu_inst_int_ckg[60]) );
  NAND2_X1 npu_inst_U174 ( .A1(npu_inst_n129), .A2(npu_inst_n137), .ZN(
        npu_inst_int_ckg[58]) );
  NAND2_X1 npu_inst_U173 ( .A1(npu_inst_n129), .A2(npu_inst_n138), .ZN(
        npu_inst_int_ckg[57]) );
  NAND2_X1 npu_inst_U172 ( .A1(npu_inst_n129), .A2(npu_inst_n139), .ZN(
        npu_inst_int_ckg[56]) );
  NAND2_X1 npu_inst_U171 ( .A1(npu_inst_n131), .A2(npu_inst_n128), .ZN(
        npu_inst_int_ckg[55]) );
  NAND2_X1 npu_inst_U170 ( .A1(npu_inst_n131), .A2(npu_inst_n130), .ZN(
        npu_inst_int_ckg[54]) );
  NAND2_X1 npu_inst_U169 ( .A1(npu_inst_n131), .A2(npu_inst_n135), .ZN(
        npu_inst_int_ckg[53]) );
  NAND2_X1 npu_inst_U168 ( .A1(npu_inst_n131), .A2(npu_inst_n132), .ZN(
        npu_inst_int_ckg[52]) );
  NAND2_X1 npu_inst_U167 ( .A1(npu_inst_n131), .A2(npu_inst_n136), .ZN(
        npu_inst_int_ckg[51]) );
  NAND2_X1 npu_inst_U166 ( .A1(npu_inst_n131), .A2(npu_inst_n137), .ZN(
        npu_inst_int_ckg[50]) );
  NAND2_X1 npu_inst_U165 ( .A1(npu_inst_n131), .A2(npu_inst_n138), .ZN(
        npu_inst_int_ckg[49]) );
  NAND2_X1 npu_inst_U164 ( .A1(npu_inst_n131), .A2(npu_inst_n139), .ZN(
        npu_inst_int_ckg[48]) );
  NAND2_X1 npu_inst_U163 ( .A1(npu_inst_n134), .A2(npu_inst_n128), .ZN(
        npu_inst_int_ckg[47]) );
  NAND2_X1 npu_inst_U162 ( .A1(npu_inst_n134), .A2(npu_inst_n130), .ZN(
        npu_inst_int_ckg[46]) );
  NAND2_X1 npu_inst_U161 ( .A1(npu_inst_n134), .A2(npu_inst_n135), .ZN(
        npu_inst_int_ckg[45]) );
  NAND2_X1 npu_inst_U160 ( .A1(npu_inst_n134), .A2(npu_inst_n132), .ZN(
        npu_inst_int_ckg[44]) );
  NAND2_X1 npu_inst_U159 ( .A1(npu_inst_n134), .A2(npu_inst_n136), .ZN(
        npu_inst_int_ckg[43]) );
  NAND2_X1 npu_inst_U158 ( .A1(npu_inst_n134), .A2(npu_inst_n137), .ZN(
        npu_inst_int_ckg[42]) );
  NAND2_X1 npu_inst_U157 ( .A1(npu_inst_n134), .A2(npu_inst_n138), .ZN(
        npu_inst_int_ckg[41]) );
  NAND2_X1 npu_inst_U156 ( .A1(npu_inst_n134), .A2(npu_inst_n139), .ZN(
        npu_inst_int_ckg[40]) );
  NAND2_X1 npu_inst_U155 ( .A1(npu_inst_n133), .A2(npu_inst_n128), .ZN(
        npu_inst_int_ckg[39]) );
  NAND2_X1 npu_inst_U154 ( .A1(npu_inst_n133), .A2(npu_inst_n130), .ZN(
        npu_inst_int_ckg[38]) );
  NAND2_X1 npu_inst_U153 ( .A1(npu_inst_n133), .A2(npu_inst_n135), .ZN(
        npu_inst_int_ckg[37]) );
  NAND2_X1 npu_inst_U152 ( .A1(npu_inst_n133), .A2(npu_inst_n132), .ZN(
        npu_inst_int_ckg[36]) );
  NAND2_X1 npu_inst_U151 ( .A1(npu_inst_n133), .A2(npu_inst_n136), .ZN(
        npu_inst_int_ckg[35]) );
  NAND2_X1 npu_inst_U150 ( .A1(npu_inst_n133), .A2(npu_inst_n137), .ZN(
        npu_inst_int_ckg[34]) );
  NAND2_X1 npu_inst_U149 ( .A1(npu_inst_n133), .A2(npu_inst_n138), .ZN(
        npu_inst_int_ckg[33]) );
  NAND2_X1 npu_inst_U148 ( .A1(npu_inst_n133), .A2(npu_inst_n139), .ZN(
        npu_inst_int_ckg[32]) );
  NAND2_X1 npu_inst_U147 ( .A1(npu_inst_n143), .A2(npu_inst_n130), .ZN(
        npu_inst_int_ckg[30]) );
  NAND2_X1 npu_inst_U146 ( .A1(npu_inst_n143), .A2(npu_inst_n135), .ZN(
        npu_inst_int_ckg[29]) );
  NAND2_X1 npu_inst_U145 ( .A1(npu_inst_n143), .A2(npu_inst_n132), .ZN(
        npu_inst_int_ckg[28]) );
  NAND2_X1 npu_inst_U144 ( .A1(npu_inst_n143), .A2(npu_inst_n137), .ZN(
        npu_inst_int_ckg[26]) );
  NAND2_X1 npu_inst_U143 ( .A1(npu_inst_n143), .A2(npu_inst_n138), .ZN(
        npu_inst_int_ckg[25]) );
  NAND2_X1 npu_inst_U142 ( .A1(npu_inst_n143), .A2(npu_inst_n139), .ZN(
        npu_inst_int_ckg[24]) );
  NAND2_X1 npu_inst_U141 ( .A1(npu_inst_n141), .A2(npu_inst_n128), .ZN(
        npu_inst_int_ckg[23]) );
  NAND2_X1 npu_inst_U140 ( .A1(npu_inst_n141), .A2(npu_inst_n130), .ZN(
        npu_inst_int_ckg[22]) );
  NAND2_X1 npu_inst_U139 ( .A1(npu_inst_n141), .A2(npu_inst_n135), .ZN(
        npu_inst_int_ckg[21]) );
  NAND2_X1 npu_inst_U138 ( .A1(npu_inst_n141), .A2(npu_inst_n132), .ZN(
        npu_inst_int_ckg[20]) );
  NAND2_X1 npu_inst_U137 ( .A1(npu_inst_n141), .A2(npu_inst_n136), .ZN(
        npu_inst_int_ckg[19]) );
  NAND2_X1 npu_inst_U136 ( .A1(npu_inst_n141), .A2(npu_inst_n137), .ZN(
        npu_inst_int_ckg[18]) );
  NAND2_X1 npu_inst_U135 ( .A1(npu_inst_n141), .A2(npu_inst_n138), .ZN(
        npu_inst_int_ckg[17]) );
  NAND2_X1 npu_inst_U134 ( .A1(npu_inst_n141), .A2(npu_inst_n139), .ZN(
        npu_inst_int_ckg[16]) );
  NAND2_X1 npu_inst_U133 ( .A1(npu_inst_n142), .A2(npu_inst_n128), .ZN(
        npu_inst_int_ckg[15]) );
  NAND2_X1 npu_inst_U132 ( .A1(npu_inst_n142), .A2(npu_inst_n130), .ZN(
        npu_inst_int_ckg[14]) );
  NAND2_X1 npu_inst_U131 ( .A1(npu_inst_n142), .A2(npu_inst_n135), .ZN(
        npu_inst_int_ckg[13]) );
  NAND2_X1 npu_inst_U130 ( .A1(npu_inst_n142), .A2(npu_inst_n132), .ZN(
        npu_inst_int_ckg[12]) );
  NAND2_X1 npu_inst_U129 ( .A1(npu_inst_n142), .A2(npu_inst_n136), .ZN(
        npu_inst_int_ckg[11]) );
  NAND2_X1 npu_inst_U128 ( .A1(npu_inst_n142), .A2(npu_inst_n137), .ZN(
        npu_inst_int_ckg[10]) );
  NAND2_X1 npu_inst_U127 ( .A1(npu_inst_n142), .A2(npu_inst_n138), .ZN(
        npu_inst_int_ckg[9]) );
  NAND2_X1 npu_inst_U126 ( .A1(npu_inst_n142), .A2(npu_inst_n139), .ZN(
        npu_inst_int_ckg[8]) );
  NAND2_X1 npu_inst_U125 ( .A1(npu_inst_n140), .A2(npu_inst_n139), .ZN(
        npu_inst_int_ckg[0]) );
  BUF_X1 npu_inst_U124 ( .A(ps_ctrl_wr_pipe), .Z(npu_inst_n6) );
  BUF_X1 npu_inst_U123 ( .A(ps_int_L0_ptr[2]), .Z(npu_inst_n91) );
  BUF_X1 npu_inst_U122 ( .A(ps_int_L0_ptr[2]), .Z(npu_inst_n89) );
  BUF_X1 npu_inst_U121 ( .A(ps_int_L0_ptr[2]), .Z(npu_inst_n90) );
  BUF_X1 npu_inst_U120 ( .A(ps_int_L0_ptr[1]), .Z(npu_inst_n74) );
  NAND2_X1 npu_inst_U119 ( .A1(npu_inst_n140), .A2(npu_inst_n128), .ZN(
        npu_inst_int_ckg[7]) );
  NAND2_X1 npu_inst_U118 ( .A1(npu_inst_n140), .A2(npu_inst_n130), .ZN(
        npu_inst_int_ckg[6]) );
  NAND2_X1 npu_inst_U117 ( .A1(npu_inst_n140), .A2(npu_inst_n135), .ZN(
        npu_inst_int_ckg[5]) );
  NAND2_X1 npu_inst_U116 ( .A1(npu_inst_n140), .A2(npu_inst_n132), .ZN(
        npu_inst_int_ckg[4]) );
  NAND2_X1 npu_inst_U115 ( .A1(npu_inst_n140), .A2(npu_inst_n136), .ZN(
        npu_inst_int_ckg[3]) );
  NAND2_X1 npu_inst_U114 ( .A1(npu_inst_n140), .A2(npu_inst_n137), .ZN(
        npu_inst_int_ckg[2]) );
  NAND2_X1 npu_inst_U113 ( .A1(npu_inst_n140), .A2(npu_inst_n138), .ZN(
        npu_inst_int_ckg[1]) );
  BUF_X1 npu_inst_U112 ( .A(ps_int_L0_ptr[1]), .Z(npu_inst_n73) );
  BUF_X1 npu_inst_U111 ( .A(ps_int_L0_ptr[0]), .Z(npu_inst_n71) );
  BUF_X1 npu_inst_U110 ( .A(ps_int_L0_ptr[0]), .Z(npu_inst_n70) );
  BUF_X1 npu_inst_U109 ( .A(ps_int_L0_ptr[0]), .Z(npu_inst_n69) );
  BUF_X1 npu_inst_U108 ( .A(ps_int_L0_ptr[0]), .Z(npu_inst_n68) );
  BUF_X1 npu_inst_U107 ( .A(ps_int_L0_ptr[0]), .Z(npu_inst_n67) );
  INV_X1 npu_inst_U106 ( .A(int_ckg_rmask[1]), .ZN(npu_inst_n131) );
  INV_X1 npu_inst_U105 ( .A(int_ckg_rmask[2]), .ZN(npu_inst_n134) );
  INV_X1 npu_inst_U104 ( .A(int_ckg_rmask[3]), .ZN(npu_inst_n133) );
  INV_X1 npu_inst_U103 ( .A(int_ckg_rmask[7]), .ZN(npu_inst_n140) );
  INV_X1 npu_inst_U102 ( .A(int_ckg_cmask[1]), .ZN(npu_inst_n130) );
  INV_X1 npu_inst_U101 ( .A(int_ckg_cmask[2]), .ZN(npu_inst_n135) );
  INV_X1 npu_inst_U100 ( .A(int_ckg_cmask[3]), .ZN(npu_inst_n132) );
  INV_X1 npu_inst_U99 ( .A(int_ckg_cmask[7]), .ZN(npu_inst_n139) );
  INV_X1 npu_inst_U98 ( .A(int_ckg_cmask[6]), .ZN(npu_inst_n138) );
  BUF_X1 npu_inst_U97 ( .A(npu_inst_n5), .Z(npu_inst_n4) );
  BUF_X1 npu_inst_U96 ( .A(npu_inst_n6), .Z(npu_inst_n2) );
  BUF_X1 npu_inst_U95 ( .A(npu_inst_n5), .Z(npu_inst_n3) );
  BUF_X2 npu_inst_U94 ( .A(npu_inst_n51), .Z(npu_inst_n60) );
  BUF_X2 npu_inst_U93 ( .A(npu_inst_n51), .Z(npu_inst_n59) );
  BUF_X2 npu_inst_U92 ( .A(npu_inst_n51), .Z(npu_inst_n58) );
  BUF_X2 npu_inst_U91 ( .A(npu_inst_n51), .Z(npu_inst_n57) );
  BUF_X2 npu_inst_U90 ( .A(npu_inst_n50), .Z(npu_inst_n56) );
  BUF_X2 npu_inst_U89 ( .A(npu_inst_n50), .Z(npu_inst_n55) );
  BUF_X2 npu_inst_U88 ( .A(npu_inst_n50), .Z(npu_inst_n54) );
  BUF_X2 npu_inst_U87 ( .A(npu_inst_n50), .Z(npu_inst_n53) );
  BUF_X2 npu_inst_U86 ( .A(npu_inst_n50), .Z(npu_inst_n52) );
  BUF_X1 npu_inst_U85 ( .A(npu_inst_n91), .Z(npu_inst_n82) );
  BUF_X1 npu_inst_U84 ( .A(npu_inst_n91), .Z(npu_inst_n81) );
  BUF_X1 npu_inst_U83 ( .A(npu_inst_n89), .Z(npu_inst_n88) );
  BUF_X1 npu_inst_U82 ( .A(npu_inst_n89), .Z(npu_inst_n87) );
  BUF_X1 npu_inst_U81 ( .A(npu_inst_n89), .Z(npu_inst_n86) );
  BUF_X1 npu_inst_U80 ( .A(npu_inst_n90), .Z(npu_inst_n85) );
  BUF_X1 npu_inst_U79 ( .A(npu_inst_n90), .Z(npu_inst_n84) );
  BUF_X1 npu_inst_U78 ( .A(npu_inst_n90), .Z(npu_inst_n83) );
  BUF_X1 npu_inst_U77 ( .A(npu_inst_n6), .Z(npu_inst_n1) );
  BUF_X1 npu_inst_U76 ( .A(npu_inst_n74), .Z(npu_inst_n80) );
  INV_X1 npu_inst_U75 ( .A(n40), .ZN(npu_inst_n141) );
  INV_X1 npu_inst_U74 ( .A(int_ckg_rmask[6]), .ZN(npu_inst_n142) );
  BUF_X1 npu_inst_U73 ( .A(npu_inst_n74), .Z(npu_inst_n79) );
  BUF_X1 npu_inst_U72 ( .A(npu_inst_n74), .Z(npu_inst_n78) );
  BUF_X1 npu_inst_U71 ( .A(npu_inst_n73), .Z(npu_inst_n77) );
  BUF_X1 npu_inst_U70 ( .A(npu_inst_n73), .Z(npu_inst_n76) );
  BUF_X1 npu_inst_U69 ( .A(npu_inst_n73), .Z(npu_inst_n75) );
  INV_X1 npu_inst_U68 ( .A(n39), .ZN(npu_inst_n137) );
  BUF_X1 npu_inst_U67 ( .A(rst), .Z(npu_inst_n121) );
  BUF_X1 npu_inst_U66 ( .A(rst), .Z(npu_inst_n120) );
  BUF_X1 npu_inst_U65 ( .A(npu_inst_n4), .Z(npu_inst_n49) );
  BUF_X1 npu_inst_U64 ( .A(npu_inst_n4), .Z(npu_inst_n48) );
  BUF_X1 npu_inst_U63 ( .A(npu_inst_n1), .Z(npu_inst_n41) );
  BUF_X1 npu_inst_U62 ( .A(npu_inst_n2), .Z(npu_inst_n42) );
  BUF_X1 npu_inst_U61 ( .A(npu_inst_n2), .Z(npu_inst_n43) );
  BUF_X1 npu_inst_U60 ( .A(npu_inst_n2), .Z(npu_inst_n44) );
  BUF_X1 npu_inst_U59 ( .A(npu_inst_n3), .Z(npu_inst_n45) );
  BUF_X1 npu_inst_U58 ( .A(npu_inst_n3), .Z(npu_inst_n46) );
  BUF_X1 npu_inst_U57 ( .A(npu_inst_n3), .Z(npu_inst_n47) );
  BUF_X1 npu_inst_U56 ( .A(npu_inst_n1), .Z(npu_inst_n39) );
  BUF_X1 npu_inst_U55 ( .A(npu_inst_n1), .Z(npu_inst_n40) );
  BUF_X1 npu_inst_U54 ( .A(npu_inst_n88), .Z(npu_inst_n107) );
  BUF_X1 npu_inst_U53 ( .A(npu_inst_n88), .Z(npu_inst_n106) );
  BUF_X1 npu_inst_U52 ( .A(npu_inst_n87), .Z(npu_inst_n105) );
  BUF_X1 npu_inst_U51 ( .A(npu_inst_n87), .Z(npu_inst_n104) );
  BUF_X1 npu_inst_U50 ( .A(npu_inst_n86), .Z(npu_inst_n103) );
  BUF_X1 npu_inst_U49 ( .A(npu_inst_n86), .Z(npu_inst_n102) );
  BUF_X1 npu_inst_U48 ( .A(npu_inst_n85), .Z(npu_inst_n101) );
  BUF_X1 npu_inst_U47 ( .A(npu_inst_n85), .Z(npu_inst_n100) );
  BUF_X1 npu_inst_U46 ( .A(npu_inst_n84), .Z(npu_inst_n99) );
  BUF_X1 npu_inst_U45 ( .A(npu_inst_n84), .Z(npu_inst_n98) );
  BUF_X1 npu_inst_U44 ( .A(npu_inst_n83), .Z(npu_inst_n97) );
  BUF_X1 npu_inst_U43 ( .A(npu_inst_n83), .Z(npu_inst_n96) );
  BUF_X1 npu_inst_U42 ( .A(npu_inst_n82), .Z(npu_inst_n95) );
  BUF_X1 npu_inst_U41 ( .A(npu_inst_n82), .Z(npu_inst_n94) );
  BUF_X1 npu_inst_U40 ( .A(npu_inst_n81), .Z(npu_inst_n93) );
  BUF_X1 npu_inst_U39 ( .A(npu_inst_n81), .Z(npu_inst_n92) );
  BUF_X1 npu_inst_U38 ( .A(npu_inst_n121), .Z(npu_inst_n127) );
  BUF_X1 npu_inst_U37 ( .A(npu_inst_n49), .Z(npu_inst_n8) );
  BUF_X1 npu_inst_U36 ( .A(npu_inst_n49), .Z(npu_inst_n7) );
  BUF_X1 npu_inst_U35 ( .A(npu_inst_n40), .Z(npu_inst_n34) );
  BUF_X1 npu_inst_U34 ( .A(npu_inst_n40), .Z(npu_inst_n33) );
  BUF_X1 npu_inst_U33 ( .A(npu_inst_n41), .Z(npu_inst_n32) );
  BUF_X1 npu_inst_U32 ( .A(npu_inst_n41), .Z(npu_inst_n31) );
  BUF_X1 npu_inst_U31 ( .A(npu_inst_n41), .Z(npu_inst_n30) );
  BUF_X1 npu_inst_U30 ( .A(npu_inst_n42), .Z(npu_inst_n29) );
  BUF_X1 npu_inst_U29 ( .A(npu_inst_n42), .Z(npu_inst_n28) );
  BUF_X1 npu_inst_U28 ( .A(npu_inst_n42), .Z(npu_inst_n27) );
  BUF_X1 npu_inst_U27 ( .A(npu_inst_n43), .Z(npu_inst_n26) );
  BUF_X1 npu_inst_U26 ( .A(npu_inst_n43), .Z(npu_inst_n25) );
  BUF_X1 npu_inst_U25 ( .A(npu_inst_n43), .Z(npu_inst_n24) );
  BUF_X1 npu_inst_U24 ( .A(npu_inst_n44), .Z(npu_inst_n23) );
  BUF_X1 npu_inst_U23 ( .A(npu_inst_n44), .Z(npu_inst_n22) );
  BUF_X1 npu_inst_U22 ( .A(npu_inst_n44), .Z(npu_inst_n21) );
  BUF_X1 npu_inst_U21 ( .A(npu_inst_n45), .Z(npu_inst_n20) );
  BUF_X1 npu_inst_U20 ( .A(npu_inst_n45), .Z(npu_inst_n19) );
  BUF_X1 npu_inst_U19 ( .A(npu_inst_n45), .Z(npu_inst_n18) );
  BUF_X1 npu_inst_U18 ( .A(npu_inst_n46), .Z(npu_inst_n17) );
  BUF_X1 npu_inst_U17 ( .A(npu_inst_n46), .Z(npu_inst_n16) );
  BUF_X1 npu_inst_U16 ( .A(npu_inst_n46), .Z(npu_inst_n15) );
  BUF_X1 npu_inst_U15 ( .A(npu_inst_n47), .Z(npu_inst_n14) );
  BUF_X1 npu_inst_U14 ( .A(npu_inst_n47), .Z(npu_inst_n13) );
  BUF_X1 npu_inst_U13 ( .A(npu_inst_n47), .Z(npu_inst_n12) );
  BUF_X1 npu_inst_U12 ( .A(npu_inst_n48), .Z(npu_inst_n11) );
  BUF_X1 npu_inst_U11 ( .A(npu_inst_n48), .Z(npu_inst_n10) );
  BUF_X1 npu_inst_U10 ( .A(npu_inst_n48), .Z(npu_inst_n9) );
  BUF_X1 npu_inst_U9 ( .A(npu_inst_n39), .Z(npu_inst_n38) );
  BUF_X1 npu_inst_U8 ( .A(npu_inst_n39), .Z(npu_inst_n37) );
  BUF_X1 npu_inst_U7 ( .A(npu_inst_n39), .Z(npu_inst_n36) );
  BUF_X1 npu_inst_U6 ( .A(npu_inst_n40), .Z(npu_inst_n35) );
  BUF_X1 npu_inst_U5 ( .A(npu_inst_n121), .Z(npu_inst_n126) );
  BUF_X1 npu_inst_U4 ( .A(npu_inst_n121), .Z(npu_inst_n125) );
  BUF_X1 npu_inst_U3 ( .A(npu_inst_n120), .Z(npu_inst_n124) );
  BUF_X1 npu_inst_U2 ( .A(npu_inst_n120), .Z(npu_inst_n123) );
  BUF_X1 npu_inst_U1 ( .A(npu_inst_n120), .Z(npu_inst_n122) );
  MUX2_X1 npu_inst_pe_1_0_0_U161 ( .A(npu_inst_pe_1_0_0_n31), .B(
        npu_inst_pe_1_0_0_n28), .S(npu_inst_pe_1_0_0_n7), .Z(
        npu_inst_pe_1_0_0_N93) );
  MUX2_X1 npu_inst_pe_1_0_0_U160 ( .A(npu_inst_pe_1_0_0_n30), .B(
        npu_inst_pe_1_0_0_n29), .S(npu_inst_n80), .Z(npu_inst_pe_1_0_0_n31) );
  MUX2_X1 npu_inst_pe_1_0_0_U159 ( .A(npu_inst_pe_1_0_0_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_0_0_int_q_reg_v_1__0_), .S(npu_inst_pe_1_0_0_n4), .Z(
        npu_inst_pe_1_0_0_n30) );
  MUX2_X1 npu_inst_pe_1_0_0_U158 ( .A(npu_inst_pe_1_0_0_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_0_0_int_q_reg_v_3__0_), .S(npu_inst_pe_1_0_0_n4), .Z(
        npu_inst_pe_1_0_0_n29) );
  MUX2_X1 npu_inst_pe_1_0_0_U157 ( .A(npu_inst_pe_1_0_0_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_0_0_int_q_reg_v_5__0_), .S(npu_inst_pe_1_0_0_n4), .Z(
        npu_inst_pe_1_0_0_n28) );
  MUX2_X1 npu_inst_pe_1_0_0_U156 ( .A(npu_inst_pe_1_0_0_n25), .B(
        npu_inst_pe_1_0_0_n22), .S(npu_inst_pe_1_0_0_n7), .Z(
        npu_inst_pe_1_0_0_N94) );
  MUX2_X1 npu_inst_pe_1_0_0_U155 ( .A(npu_inst_pe_1_0_0_n24), .B(
        npu_inst_pe_1_0_0_n23), .S(npu_inst_n80), .Z(npu_inst_pe_1_0_0_n25) );
  MUX2_X1 npu_inst_pe_1_0_0_U154 ( .A(npu_inst_pe_1_0_0_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_0_0_int_q_reg_v_1__1_), .S(npu_inst_pe_1_0_0_n4), .Z(
        npu_inst_pe_1_0_0_n24) );
  MUX2_X1 npu_inst_pe_1_0_0_U153 ( .A(npu_inst_pe_1_0_0_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_0_0_int_q_reg_v_3__1_), .S(npu_inst_pe_1_0_0_n4), .Z(
        npu_inst_pe_1_0_0_n23) );
  MUX2_X1 npu_inst_pe_1_0_0_U152 ( .A(npu_inst_pe_1_0_0_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_0_0_int_q_reg_v_5__1_), .S(npu_inst_pe_1_0_0_n4), .Z(
        npu_inst_pe_1_0_0_n22) );
  MUX2_X1 npu_inst_pe_1_0_0_U151 ( .A(npu_inst_pe_1_0_0_n21), .B(
        npu_inst_pe_1_0_0_n18), .S(npu_inst_pe_1_0_0_n7), .Z(
        npu_inst_pe_1_0_0_o_data_h_1_) );
  MUX2_X1 npu_inst_pe_1_0_0_U150 ( .A(npu_inst_pe_1_0_0_n20), .B(
        npu_inst_pe_1_0_0_n19), .S(npu_inst_n80), .Z(npu_inst_pe_1_0_0_n21) );
  MUX2_X1 npu_inst_pe_1_0_0_U149 ( .A(npu_inst_pe_1_0_0_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_0_0_int_q_reg_h_1__1_), .S(npu_inst_pe_1_0_0_n4), .Z(
        npu_inst_pe_1_0_0_n20) );
  MUX2_X1 npu_inst_pe_1_0_0_U148 ( .A(npu_inst_pe_1_0_0_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_0_0_int_q_reg_h_3__1_), .S(npu_inst_pe_1_0_0_n4), .Z(
        npu_inst_pe_1_0_0_n19) );
  MUX2_X1 npu_inst_pe_1_0_0_U147 ( .A(npu_inst_pe_1_0_0_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_0_0_int_q_reg_h_5__1_), .S(npu_inst_pe_1_0_0_n4), .Z(
        npu_inst_pe_1_0_0_n18) );
  MUX2_X1 npu_inst_pe_1_0_0_U146 ( .A(npu_inst_pe_1_0_0_n17), .B(
        npu_inst_pe_1_0_0_n14), .S(npu_inst_pe_1_0_0_n7), .Z(
        npu_inst_pe_1_0_0_o_data_h_0_) );
  MUX2_X1 npu_inst_pe_1_0_0_U145 ( .A(npu_inst_pe_1_0_0_n16), .B(
        npu_inst_pe_1_0_0_n15), .S(npu_inst_n80), .Z(npu_inst_pe_1_0_0_n17) );
  MUX2_X1 npu_inst_pe_1_0_0_U144 ( .A(npu_inst_pe_1_0_0_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_0_0_int_q_reg_h_1__0_), .S(npu_inst_pe_1_0_0_n4), .Z(
        npu_inst_pe_1_0_0_n16) );
  MUX2_X1 npu_inst_pe_1_0_0_U143 ( .A(npu_inst_pe_1_0_0_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_0_0_int_q_reg_h_3__0_), .S(npu_inst_pe_1_0_0_n4), .Z(
        npu_inst_pe_1_0_0_n15) );
  MUX2_X1 npu_inst_pe_1_0_0_U142 ( .A(npu_inst_pe_1_0_0_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_0_0_int_q_reg_h_5__0_), .S(npu_inst_pe_1_0_0_n4), .Z(
        npu_inst_pe_1_0_0_n14) );
  XOR2_X1 npu_inst_pe_1_0_0_U141 ( .A(npu_inst_pe_1_0_0_int_data_0_), .B(
        npu_inst_pe_1_0_0_int_q_acc_0_), .Z(npu_inst_pe_1_0_0_N73) );
  AND2_X1 npu_inst_pe_1_0_0_U140 ( .A1(npu_inst_pe_1_0_0_int_q_acc_0_), .A2(
        npu_inst_pe_1_0_0_int_data_0_), .ZN(npu_inst_pe_1_0_0_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_0_0_U139 ( .A(npu_inst_pe_1_0_0_int_q_acc_0_), .B(
        npu_inst_pe_1_0_0_n12), .ZN(npu_inst_pe_1_0_0_N65) );
  OR2_X1 npu_inst_pe_1_0_0_U138 ( .A1(npu_inst_pe_1_0_0_n12), .A2(
        npu_inst_pe_1_0_0_int_q_acc_0_), .ZN(npu_inst_pe_1_0_0_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_0_0_U137 ( .A(npu_inst_pe_1_0_0_int_q_acc_2_), .B(
        npu_inst_pe_1_0_0_add_69_carry_2_), .Z(npu_inst_pe_1_0_0_N75) );
  AND2_X1 npu_inst_pe_1_0_0_U136 ( .A1(npu_inst_pe_1_0_0_add_69_carry_2_), 
        .A2(npu_inst_pe_1_0_0_int_q_acc_2_), .ZN(
        npu_inst_pe_1_0_0_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_0_0_U135 ( .A(npu_inst_pe_1_0_0_int_q_acc_3_), .B(
        npu_inst_pe_1_0_0_add_69_carry_3_), .Z(npu_inst_pe_1_0_0_N76) );
  AND2_X1 npu_inst_pe_1_0_0_U134 ( .A1(npu_inst_pe_1_0_0_add_69_carry_3_), 
        .A2(npu_inst_pe_1_0_0_int_q_acc_3_), .ZN(
        npu_inst_pe_1_0_0_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_0_0_U133 ( .A(npu_inst_pe_1_0_0_int_q_acc_4_), .B(
        npu_inst_pe_1_0_0_add_69_carry_4_), .Z(npu_inst_pe_1_0_0_N77) );
  AND2_X1 npu_inst_pe_1_0_0_U132 ( .A1(npu_inst_pe_1_0_0_add_69_carry_4_), 
        .A2(npu_inst_pe_1_0_0_int_q_acc_4_), .ZN(
        npu_inst_pe_1_0_0_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_0_0_U131 ( .A(npu_inst_pe_1_0_0_int_q_acc_5_), .B(
        npu_inst_pe_1_0_0_add_69_carry_5_), .Z(npu_inst_pe_1_0_0_N78) );
  AND2_X1 npu_inst_pe_1_0_0_U130 ( .A1(npu_inst_pe_1_0_0_add_69_carry_5_), 
        .A2(npu_inst_pe_1_0_0_int_q_acc_5_), .ZN(
        npu_inst_pe_1_0_0_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_0_0_U129 ( .A(npu_inst_pe_1_0_0_int_q_acc_6_), .B(
        npu_inst_pe_1_0_0_add_69_carry_6_), .Z(npu_inst_pe_1_0_0_N79) );
  AND2_X1 npu_inst_pe_1_0_0_U128 ( .A1(npu_inst_pe_1_0_0_add_69_carry_6_), 
        .A2(npu_inst_pe_1_0_0_int_q_acc_6_), .ZN(
        npu_inst_pe_1_0_0_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_0_0_U127 ( .A(npu_inst_pe_1_0_0_int_q_acc_7_), .B(
        npu_inst_pe_1_0_0_add_69_carry_7_), .Z(npu_inst_pe_1_0_0_N80) );
  XNOR2_X1 npu_inst_pe_1_0_0_U126 ( .A(npu_inst_pe_1_0_0_sub_67_carry_2_), .B(
        npu_inst_pe_1_0_0_int_q_acc_2_), .ZN(npu_inst_pe_1_0_0_N67) );
  OR2_X1 npu_inst_pe_1_0_0_U125 ( .A1(npu_inst_pe_1_0_0_int_q_acc_2_), .A2(
        npu_inst_pe_1_0_0_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_0_0_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_0_0_U124 ( .A(npu_inst_pe_1_0_0_sub_67_carry_3_), .B(
        npu_inst_pe_1_0_0_int_q_acc_3_), .ZN(npu_inst_pe_1_0_0_N68) );
  OR2_X1 npu_inst_pe_1_0_0_U123 ( .A1(npu_inst_pe_1_0_0_int_q_acc_3_), .A2(
        npu_inst_pe_1_0_0_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_0_0_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_0_0_U122 ( .A(npu_inst_pe_1_0_0_sub_67_carry_4_), .B(
        npu_inst_pe_1_0_0_int_q_acc_4_), .ZN(npu_inst_pe_1_0_0_N69) );
  OR2_X1 npu_inst_pe_1_0_0_U121 ( .A1(npu_inst_pe_1_0_0_int_q_acc_4_), .A2(
        npu_inst_pe_1_0_0_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_0_0_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_0_0_U120 ( .A(npu_inst_pe_1_0_0_sub_67_carry_5_), .B(
        npu_inst_pe_1_0_0_int_q_acc_5_), .ZN(npu_inst_pe_1_0_0_N70) );
  OR2_X1 npu_inst_pe_1_0_0_U119 ( .A1(npu_inst_pe_1_0_0_int_q_acc_5_), .A2(
        npu_inst_pe_1_0_0_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_0_0_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_0_0_U118 ( .A(npu_inst_pe_1_0_0_sub_67_carry_6_), .B(
        npu_inst_pe_1_0_0_int_q_acc_6_), .ZN(npu_inst_pe_1_0_0_N71) );
  OR2_X1 npu_inst_pe_1_0_0_U117 ( .A1(npu_inst_pe_1_0_0_int_q_acc_6_), .A2(
        npu_inst_pe_1_0_0_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_0_0_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_0_0_U116 ( .A(npu_inst_pe_1_0_0_int_q_acc_7_), .B(
        npu_inst_pe_1_0_0_sub_67_carry_7_), .ZN(npu_inst_pe_1_0_0_N72) );
  INV_X1 npu_inst_pe_1_0_0_U115 ( .A(npu_inst_n80), .ZN(npu_inst_pe_1_0_0_n6)
         );
  INV_X1 npu_inst_pe_1_0_0_U114 ( .A(npu_inst_n57), .ZN(npu_inst_pe_1_0_0_n3)
         );
  AOI22_X1 npu_inst_pe_1_0_0_U113 ( .A1(npu_inst_int_data_y_1__0__0_), .A2(
        npu_inst_pe_1_0_0_n58), .B1(npu_inst_pe_1_0_0_n118), .B2(
        npu_inst_pe_1_0_0_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_0_0_n57) );
  INV_X1 npu_inst_pe_1_0_0_U112 ( .A(npu_inst_pe_1_0_0_n57), .ZN(
        npu_inst_pe_1_0_0_n107) );
  AOI22_X1 npu_inst_pe_1_0_0_U111 ( .A1(npu_inst_int_data_y_1__0__0_), .A2(
        npu_inst_pe_1_0_0_n54), .B1(npu_inst_pe_1_0_0_n117), .B2(
        npu_inst_pe_1_0_0_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_0_0_n53) );
  INV_X1 npu_inst_pe_1_0_0_U110 ( .A(npu_inst_pe_1_0_0_n53), .ZN(
        npu_inst_pe_1_0_0_n108) );
  AOI22_X1 npu_inst_pe_1_0_0_U107 ( .A1(npu_inst_int_data_y_1__0__0_), .A2(
        npu_inst_pe_1_0_0_n50), .B1(npu_inst_pe_1_0_0_n116), .B2(
        npu_inst_pe_1_0_0_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_0_0_n49) );
  INV_X1 npu_inst_pe_1_0_0_U106 ( .A(npu_inst_pe_1_0_0_n49), .ZN(
        npu_inst_pe_1_0_0_n109) );
  AOI22_X1 npu_inst_pe_1_0_0_U105 ( .A1(npu_inst_int_data_y_1__0__0_), .A2(
        npu_inst_pe_1_0_0_n46), .B1(npu_inst_pe_1_0_0_n115), .B2(
        npu_inst_pe_1_0_0_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_0_0_n45) );
  INV_X1 npu_inst_pe_1_0_0_U104 ( .A(npu_inst_pe_1_0_0_n45), .ZN(
        npu_inst_pe_1_0_0_n110) );
  AOI22_X1 npu_inst_pe_1_0_0_U103 ( .A1(npu_inst_int_data_y_1__0__0_), .A2(
        npu_inst_pe_1_0_0_n42), .B1(npu_inst_pe_1_0_0_n114), .B2(
        npu_inst_pe_1_0_0_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_0_0_n41) );
  INV_X1 npu_inst_pe_1_0_0_U102 ( .A(npu_inst_pe_1_0_0_n41), .ZN(
        npu_inst_pe_1_0_0_n111) );
  AOI22_X1 npu_inst_pe_1_0_0_U101 ( .A1(npu_inst_int_data_y_1__0__1_), .A2(
        npu_inst_pe_1_0_0_n58), .B1(npu_inst_pe_1_0_0_n118), .B2(
        npu_inst_pe_1_0_0_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_0_0_n59) );
  INV_X1 npu_inst_pe_1_0_0_U100 ( .A(npu_inst_pe_1_0_0_n59), .ZN(
        npu_inst_pe_1_0_0_n101) );
  AOI22_X1 npu_inst_pe_1_0_0_U99 ( .A1(npu_inst_int_data_y_1__0__1_), .A2(
        npu_inst_pe_1_0_0_n54), .B1(npu_inst_pe_1_0_0_n117), .B2(
        npu_inst_pe_1_0_0_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_0_0_n55) );
  INV_X1 npu_inst_pe_1_0_0_U98 ( .A(npu_inst_pe_1_0_0_n55), .ZN(
        npu_inst_pe_1_0_0_n102) );
  AOI22_X1 npu_inst_pe_1_0_0_U97 ( .A1(npu_inst_int_data_y_1__0__1_), .A2(
        npu_inst_pe_1_0_0_n50), .B1(npu_inst_pe_1_0_0_n116), .B2(
        npu_inst_pe_1_0_0_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_0_0_n51) );
  INV_X1 npu_inst_pe_1_0_0_U96 ( .A(npu_inst_pe_1_0_0_n51), .ZN(
        npu_inst_pe_1_0_0_n103) );
  AOI22_X1 npu_inst_pe_1_0_0_U95 ( .A1(npu_inst_int_data_y_1__0__1_), .A2(
        npu_inst_pe_1_0_0_n46), .B1(npu_inst_pe_1_0_0_n115), .B2(
        npu_inst_pe_1_0_0_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_0_0_n47) );
  INV_X1 npu_inst_pe_1_0_0_U94 ( .A(npu_inst_pe_1_0_0_n47), .ZN(
        npu_inst_pe_1_0_0_n104) );
  AOI22_X1 npu_inst_pe_1_0_0_U93 ( .A1(npu_inst_int_data_y_1__0__1_), .A2(
        npu_inst_pe_1_0_0_n42), .B1(npu_inst_pe_1_0_0_n114), .B2(
        npu_inst_pe_1_0_0_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_0_0_n43) );
  INV_X1 npu_inst_pe_1_0_0_U92 ( .A(npu_inst_pe_1_0_0_n43), .ZN(
        npu_inst_pe_1_0_0_n105) );
  AOI22_X1 npu_inst_pe_1_0_0_U91 ( .A1(npu_inst_pe_1_0_0_n38), .A2(
        npu_inst_int_data_y_1__0__1_), .B1(npu_inst_pe_1_0_0_n113), .B2(
        npu_inst_pe_1_0_0_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_0_0_n39) );
  INV_X1 npu_inst_pe_1_0_0_U90 ( .A(npu_inst_pe_1_0_0_n39), .ZN(
        npu_inst_pe_1_0_0_n106) );
  AOI22_X1 npu_inst_pe_1_0_0_U89 ( .A1(npu_inst_pe_1_0_0_n38), .A2(
        npu_inst_int_data_y_1__0__0_), .B1(npu_inst_pe_1_0_0_n113), .B2(
        npu_inst_pe_1_0_0_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_0_0_n37) );
  INV_X1 npu_inst_pe_1_0_0_U88 ( .A(npu_inst_pe_1_0_0_n37), .ZN(
        npu_inst_pe_1_0_0_n112) );
  NOR3_X1 npu_inst_pe_1_0_0_U87 ( .A1(npu_inst_pe_1_0_0_n26), .A2(npu_inst_n57), .A3(npu_inst_int_ckg[63]), .ZN(npu_inst_pe_1_0_0_n85) );
  OR2_X1 npu_inst_pe_1_0_0_U86 ( .A1(npu_inst_pe_1_0_0_n85), .A2(
        npu_inst_pe_1_0_0_n2), .ZN(npu_inst_pe_1_0_0_N84) );
  NAND2_X1 npu_inst_pe_1_0_0_U85 ( .A1(npu_inst_pe_1_0_0_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_0_0_n60), .ZN(npu_inst_pe_1_0_0_n74) );
  OAI21_X1 npu_inst_pe_1_0_0_U84 ( .B1(npu_inst_pe_1_0_0_n63), .B2(
        npu_inst_pe_1_0_0_n60), .A(npu_inst_pe_1_0_0_n74), .ZN(
        npu_inst_pe_1_0_0_n97) );
  NAND2_X1 npu_inst_pe_1_0_0_U83 ( .A1(npu_inst_pe_1_0_0_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_0_0_n60), .ZN(npu_inst_pe_1_0_0_n73) );
  OAI21_X1 npu_inst_pe_1_0_0_U82 ( .B1(npu_inst_pe_1_0_0_n61), .B2(
        npu_inst_pe_1_0_0_n60), .A(npu_inst_pe_1_0_0_n73), .ZN(
        npu_inst_pe_1_0_0_n96) );
  NAND2_X1 npu_inst_pe_1_0_0_U81 ( .A1(npu_inst_pe_1_0_0_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_0_0_n56), .ZN(npu_inst_pe_1_0_0_n72) );
  OAI21_X1 npu_inst_pe_1_0_0_U80 ( .B1(npu_inst_pe_1_0_0_n63), .B2(
        npu_inst_pe_1_0_0_n56), .A(npu_inst_pe_1_0_0_n72), .ZN(
        npu_inst_pe_1_0_0_n95) );
  NAND2_X1 npu_inst_pe_1_0_0_U79 ( .A1(npu_inst_pe_1_0_0_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_0_0_n56), .ZN(npu_inst_pe_1_0_0_n71) );
  OAI21_X1 npu_inst_pe_1_0_0_U78 ( .B1(npu_inst_pe_1_0_0_n61), .B2(
        npu_inst_pe_1_0_0_n56), .A(npu_inst_pe_1_0_0_n71), .ZN(
        npu_inst_pe_1_0_0_n94) );
  NAND2_X1 npu_inst_pe_1_0_0_U77 ( .A1(npu_inst_pe_1_0_0_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_0_0_n52), .ZN(npu_inst_pe_1_0_0_n70) );
  OAI21_X1 npu_inst_pe_1_0_0_U76 ( .B1(npu_inst_pe_1_0_0_n63), .B2(
        npu_inst_pe_1_0_0_n52), .A(npu_inst_pe_1_0_0_n70), .ZN(
        npu_inst_pe_1_0_0_n93) );
  NAND2_X1 npu_inst_pe_1_0_0_U75 ( .A1(npu_inst_pe_1_0_0_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_0_0_n52), .ZN(npu_inst_pe_1_0_0_n69) );
  OAI21_X1 npu_inst_pe_1_0_0_U74 ( .B1(npu_inst_pe_1_0_0_n61), .B2(
        npu_inst_pe_1_0_0_n52), .A(npu_inst_pe_1_0_0_n69), .ZN(
        npu_inst_pe_1_0_0_n92) );
  NAND2_X1 npu_inst_pe_1_0_0_U73 ( .A1(npu_inst_pe_1_0_0_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_0_0_n48), .ZN(npu_inst_pe_1_0_0_n68) );
  OAI21_X1 npu_inst_pe_1_0_0_U72 ( .B1(npu_inst_pe_1_0_0_n63), .B2(
        npu_inst_pe_1_0_0_n48), .A(npu_inst_pe_1_0_0_n68), .ZN(
        npu_inst_pe_1_0_0_n91) );
  NAND2_X1 npu_inst_pe_1_0_0_U71 ( .A1(npu_inst_pe_1_0_0_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_0_0_n48), .ZN(npu_inst_pe_1_0_0_n67) );
  OAI21_X1 npu_inst_pe_1_0_0_U70 ( .B1(npu_inst_pe_1_0_0_n61), .B2(
        npu_inst_pe_1_0_0_n48), .A(npu_inst_pe_1_0_0_n67), .ZN(
        npu_inst_pe_1_0_0_n90) );
  NAND2_X1 npu_inst_pe_1_0_0_U69 ( .A1(npu_inst_pe_1_0_0_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_0_0_n44), .ZN(npu_inst_pe_1_0_0_n66) );
  OAI21_X1 npu_inst_pe_1_0_0_U68 ( .B1(npu_inst_pe_1_0_0_n63), .B2(
        npu_inst_pe_1_0_0_n44), .A(npu_inst_pe_1_0_0_n66), .ZN(
        npu_inst_pe_1_0_0_n89) );
  NAND2_X1 npu_inst_pe_1_0_0_U67 ( .A1(npu_inst_pe_1_0_0_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_0_0_n44), .ZN(npu_inst_pe_1_0_0_n65) );
  OAI21_X1 npu_inst_pe_1_0_0_U66 ( .B1(npu_inst_pe_1_0_0_n61), .B2(
        npu_inst_pe_1_0_0_n44), .A(npu_inst_pe_1_0_0_n65), .ZN(
        npu_inst_pe_1_0_0_n88) );
  NAND2_X1 npu_inst_pe_1_0_0_U65 ( .A1(npu_inst_pe_1_0_0_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_0_0_n40), .ZN(npu_inst_pe_1_0_0_n64) );
  OAI21_X1 npu_inst_pe_1_0_0_U64 ( .B1(npu_inst_pe_1_0_0_n63), .B2(
        npu_inst_pe_1_0_0_n40), .A(npu_inst_pe_1_0_0_n64), .ZN(
        npu_inst_pe_1_0_0_n87) );
  NAND2_X1 npu_inst_pe_1_0_0_U63 ( .A1(npu_inst_pe_1_0_0_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_0_0_n40), .ZN(npu_inst_pe_1_0_0_n62) );
  OAI21_X1 npu_inst_pe_1_0_0_U62 ( .B1(npu_inst_pe_1_0_0_n61), .B2(
        npu_inst_pe_1_0_0_n40), .A(npu_inst_pe_1_0_0_n62), .ZN(
        npu_inst_pe_1_0_0_n86) );
  AND2_X1 npu_inst_pe_1_0_0_U61 ( .A1(npu_inst_pe_1_0_0_int_q_acc_2_), .A2(
        npu_inst_pe_1_0_0_n1), .ZN(int_o_data_npu[58]) );
  AND2_X1 npu_inst_pe_1_0_0_U60 ( .A1(npu_inst_pe_1_0_0_int_q_acc_3_), .A2(
        npu_inst_pe_1_0_0_n2), .ZN(int_o_data_npu[59]) );
  AND2_X1 npu_inst_pe_1_0_0_U59 ( .A1(npu_inst_pe_1_0_0_int_q_acc_6_), .A2(
        npu_inst_pe_1_0_0_n2), .ZN(int_o_data_npu[62]) );
  AND2_X1 npu_inst_pe_1_0_0_U58 ( .A1(npu_inst_pe_1_0_0_int_q_acc_5_), .A2(
        npu_inst_pe_1_0_0_n2), .ZN(int_o_data_npu[61]) );
  AND2_X1 npu_inst_pe_1_0_0_U57 ( .A1(npu_inst_pe_1_0_0_int_q_acc_4_), .A2(
        npu_inst_pe_1_0_0_n2), .ZN(int_o_data_npu[60]) );
  AOI222_X1 npu_inst_pe_1_0_0_U56 ( .A1(npu_inst_int_data_res_1__0__0_), .A2(
        npu_inst_pe_1_0_0_n1), .B1(npu_inst_pe_1_0_0_N73), .B2(
        npu_inst_pe_1_0_0_n76), .C1(npu_inst_pe_1_0_0_N65), .C2(
        npu_inst_pe_1_0_0_n77), .ZN(npu_inst_pe_1_0_0_n84) );
  INV_X1 npu_inst_pe_1_0_0_U55 ( .A(npu_inst_pe_1_0_0_n84), .ZN(
        npu_inst_pe_1_0_0_n100) );
  AOI222_X1 npu_inst_pe_1_0_0_U54 ( .A1(npu_inst_int_data_res_1__0__7_), .A2(
        npu_inst_pe_1_0_0_n1), .B1(npu_inst_pe_1_0_0_N80), .B2(
        npu_inst_pe_1_0_0_n76), .C1(npu_inst_pe_1_0_0_N72), .C2(
        npu_inst_pe_1_0_0_n77), .ZN(npu_inst_pe_1_0_0_n75) );
  INV_X1 npu_inst_pe_1_0_0_U53 ( .A(npu_inst_pe_1_0_0_n75), .ZN(
        npu_inst_pe_1_0_0_n32) );
  AOI222_X1 npu_inst_pe_1_0_0_U52 ( .A1(npu_inst_int_data_res_1__0__1_), .A2(
        npu_inst_pe_1_0_0_n1), .B1(npu_inst_pe_1_0_0_N74), .B2(
        npu_inst_pe_1_0_0_n76), .C1(npu_inst_pe_1_0_0_N66), .C2(
        npu_inst_pe_1_0_0_n77), .ZN(npu_inst_pe_1_0_0_n83) );
  INV_X1 npu_inst_pe_1_0_0_U51 ( .A(npu_inst_pe_1_0_0_n83), .ZN(
        npu_inst_pe_1_0_0_n99) );
  AOI222_X1 npu_inst_pe_1_0_0_U50 ( .A1(npu_inst_int_data_res_1__0__2_), .A2(
        npu_inst_pe_1_0_0_n1), .B1(npu_inst_pe_1_0_0_N75), .B2(
        npu_inst_pe_1_0_0_n76), .C1(npu_inst_pe_1_0_0_N67), .C2(
        npu_inst_pe_1_0_0_n77), .ZN(npu_inst_pe_1_0_0_n82) );
  INV_X1 npu_inst_pe_1_0_0_U49 ( .A(npu_inst_pe_1_0_0_n82), .ZN(
        npu_inst_pe_1_0_0_n98) );
  AOI222_X1 npu_inst_pe_1_0_0_U48 ( .A1(npu_inst_int_data_res_1__0__3_), .A2(
        npu_inst_pe_1_0_0_n1), .B1(npu_inst_pe_1_0_0_N76), .B2(
        npu_inst_pe_1_0_0_n76), .C1(npu_inst_pe_1_0_0_N68), .C2(
        npu_inst_pe_1_0_0_n77), .ZN(npu_inst_pe_1_0_0_n81) );
  INV_X1 npu_inst_pe_1_0_0_U47 ( .A(npu_inst_pe_1_0_0_n81), .ZN(
        npu_inst_pe_1_0_0_n36) );
  AOI222_X1 npu_inst_pe_1_0_0_U46 ( .A1(npu_inst_int_data_res_1__0__4_), .A2(
        npu_inst_pe_1_0_0_n1), .B1(npu_inst_pe_1_0_0_N77), .B2(
        npu_inst_pe_1_0_0_n76), .C1(npu_inst_pe_1_0_0_N69), .C2(
        npu_inst_pe_1_0_0_n77), .ZN(npu_inst_pe_1_0_0_n80) );
  INV_X1 npu_inst_pe_1_0_0_U45 ( .A(npu_inst_pe_1_0_0_n80), .ZN(
        npu_inst_pe_1_0_0_n35) );
  AOI222_X1 npu_inst_pe_1_0_0_U44 ( .A1(npu_inst_int_data_res_1__0__5_), .A2(
        npu_inst_pe_1_0_0_n1), .B1(npu_inst_pe_1_0_0_N78), .B2(
        npu_inst_pe_1_0_0_n76), .C1(npu_inst_pe_1_0_0_N70), .C2(
        npu_inst_pe_1_0_0_n77), .ZN(npu_inst_pe_1_0_0_n79) );
  INV_X1 npu_inst_pe_1_0_0_U43 ( .A(npu_inst_pe_1_0_0_n79), .ZN(
        npu_inst_pe_1_0_0_n34) );
  AOI222_X1 npu_inst_pe_1_0_0_U42 ( .A1(npu_inst_int_data_res_1__0__6_), .A2(
        npu_inst_pe_1_0_0_n1), .B1(npu_inst_pe_1_0_0_N79), .B2(
        npu_inst_pe_1_0_0_n76), .C1(npu_inst_pe_1_0_0_N71), .C2(
        npu_inst_pe_1_0_0_n77), .ZN(npu_inst_pe_1_0_0_n78) );
  INV_X1 npu_inst_pe_1_0_0_U41 ( .A(npu_inst_pe_1_0_0_n78), .ZN(
        npu_inst_pe_1_0_0_n33) );
  AND2_X1 npu_inst_pe_1_0_0_U40 ( .A1(npu_inst_pe_1_0_0_o_data_h_1_), .A2(
        npu_inst_pe_1_0_0_int_q_weight_1_), .ZN(npu_inst_pe_1_0_0_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_0_0_U39 ( .A1(npu_inst_pe_1_0_0_o_data_h_0_), .A2(
        npu_inst_pe_1_0_0_int_q_weight_1_), .ZN(npu_inst_pe_1_0_0_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_0_0_U38 ( .A(npu_inst_pe_1_0_0_int_data_1_), .ZN(
        npu_inst_pe_1_0_0_n13) );
  AND2_X1 npu_inst_pe_1_0_0_U37 ( .A1(npu_inst_pe_1_0_0_n2), .A2(
        npu_inst_pe_1_0_0_int_q_acc_7_), .ZN(int_o_data_npu[63]) );
  AND2_X1 npu_inst_pe_1_0_0_U36 ( .A1(npu_inst_pe_1_0_0_int_q_acc_1_), .A2(
        npu_inst_pe_1_0_0_n1), .ZN(int_o_data_npu[57]) );
  AND2_X1 npu_inst_pe_1_0_0_U35 ( .A1(npu_inst_pe_1_0_0_int_q_acc_0_), .A2(
        npu_inst_pe_1_0_0_n1), .ZN(int_o_data_npu[56]) );
  AND2_X1 npu_inst_pe_1_0_0_U34 ( .A1(npu_inst_pe_1_0_0_N93), .A2(npu_inst_n57), .ZN(npu_inst_pe_1_0_0_o_data_v_0_) );
  AND2_X1 npu_inst_pe_1_0_0_U33 ( .A1(npu_inst_n57), .A2(npu_inst_pe_1_0_0_N94), .ZN(npu_inst_pe_1_0_0_o_data_v_1_) );
  AOI22_X1 npu_inst_pe_1_0_0_U32 ( .A1(npu_inst_n57), .A2(
        npu_inst_int_data_y_1__0__1_), .B1(npu_inst_pe_1_0_0_n3), .B2(
        npu_inst_int_data_x_0__1__1_), .ZN(npu_inst_pe_1_0_0_n63) );
  AOI22_X1 npu_inst_pe_1_0_0_U31 ( .A1(npu_inst_n57), .A2(
        npu_inst_int_data_y_1__0__0_), .B1(npu_inst_pe_1_0_0_n3), .B2(
        npu_inst_int_data_x_0__1__0_), .ZN(npu_inst_pe_1_0_0_n61) );
  INV_X1 npu_inst_pe_1_0_0_U30 ( .A(npu_inst_pe_1_0_0_int_data_0_), .ZN(
        npu_inst_pe_1_0_0_n12) );
  INV_X1 npu_inst_pe_1_0_0_U29 ( .A(npu_inst_n72), .ZN(npu_inst_pe_1_0_0_n5)
         );
  OR3_X1 npu_inst_pe_1_0_0_U28 ( .A1(npu_inst_n80), .A2(npu_inst_pe_1_0_0_n7), 
        .A3(npu_inst_pe_1_0_0_n5), .ZN(npu_inst_pe_1_0_0_n56) );
  OR3_X1 npu_inst_pe_1_0_0_U27 ( .A1(npu_inst_pe_1_0_0_n5), .A2(
        npu_inst_pe_1_0_0_n7), .A3(npu_inst_pe_1_0_0_n6), .ZN(
        npu_inst_pe_1_0_0_n48) );
  INV_X1 npu_inst_pe_1_0_0_U26 ( .A(npu_inst_pe_1_0_0_n5), .ZN(
        npu_inst_pe_1_0_0_n4) );
  OR3_X1 npu_inst_pe_1_0_0_U25 ( .A1(npu_inst_pe_1_0_0_n4), .A2(
        npu_inst_pe_1_0_0_n7), .A3(npu_inst_pe_1_0_0_n6), .ZN(
        npu_inst_pe_1_0_0_n52) );
  OR3_X1 npu_inst_pe_1_0_0_U24 ( .A1(npu_inst_n80), .A2(npu_inst_pe_1_0_0_n7), 
        .A3(npu_inst_pe_1_0_0_n4), .ZN(npu_inst_pe_1_0_0_n60) );
  NOR2_X1 npu_inst_pe_1_0_0_U23 ( .A1(npu_inst_pe_1_0_0_n60), .A2(
        npu_inst_pe_1_0_0_n3), .ZN(npu_inst_pe_1_0_0_n58) );
  NOR2_X1 npu_inst_pe_1_0_0_U22 ( .A1(npu_inst_pe_1_0_0_n56), .A2(
        npu_inst_pe_1_0_0_n3), .ZN(npu_inst_pe_1_0_0_n54) );
  NOR2_X1 npu_inst_pe_1_0_0_U21 ( .A1(npu_inst_pe_1_0_0_n52), .A2(
        npu_inst_pe_1_0_0_n3), .ZN(npu_inst_pe_1_0_0_n50) );
  NOR2_X1 npu_inst_pe_1_0_0_U20 ( .A1(npu_inst_pe_1_0_0_n48), .A2(
        npu_inst_pe_1_0_0_n3), .ZN(npu_inst_pe_1_0_0_n46) );
  NOR2_X1 npu_inst_pe_1_0_0_U19 ( .A1(npu_inst_pe_1_0_0_n40), .A2(
        npu_inst_pe_1_0_0_n3), .ZN(npu_inst_pe_1_0_0_n38) );
  NOR2_X1 npu_inst_pe_1_0_0_U18 ( .A1(npu_inst_pe_1_0_0_n44), .A2(
        npu_inst_pe_1_0_0_n3), .ZN(npu_inst_pe_1_0_0_n42) );
  BUF_X1 npu_inst_pe_1_0_0_U17 ( .A(npu_inst_n107), .Z(npu_inst_pe_1_0_0_n7)
         );
  INV_X1 npu_inst_pe_1_0_0_U16 ( .A(npu_inst_n127), .ZN(npu_inst_pe_1_0_0_n11)
         );
  INV_X1 npu_inst_pe_1_0_0_U15 ( .A(npu_inst_pe_1_0_0_n38), .ZN(
        npu_inst_pe_1_0_0_n113) );
  INV_X1 npu_inst_pe_1_0_0_U14 ( .A(npu_inst_pe_1_0_0_n58), .ZN(
        npu_inst_pe_1_0_0_n118) );
  INV_X1 npu_inst_pe_1_0_0_U13 ( .A(npu_inst_pe_1_0_0_n54), .ZN(
        npu_inst_pe_1_0_0_n117) );
  INV_X1 npu_inst_pe_1_0_0_U12 ( .A(npu_inst_pe_1_0_0_n50), .ZN(
        npu_inst_pe_1_0_0_n116) );
  INV_X1 npu_inst_pe_1_0_0_U11 ( .A(npu_inst_pe_1_0_0_n46), .ZN(
        npu_inst_pe_1_0_0_n115) );
  INV_X1 npu_inst_pe_1_0_0_U10 ( .A(npu_inst_pe_1_0_0_n42), .ZN(
        npu_inst_pe_1_0_0_n114) );
  BUF_X1 npu_inst_pe_1_0_0_U9 ( .A(npu_inst_n38), .Z(npu_inst_pe_1_0_0_n2) );
  BUF_X1 npu_inst_pe_1_0_0_U8 ( .A(npu_inst_n38), .Z(npu_inst_pe_1_0_0_n1) );
  BUF_X1 npu_inst_pe_1_0_0_U7 ( .A(npu_inst_pe_1_0_0_n11), .Z(
        npu_inst_pe_1_0_0_n10) );
  BUF_X1 npu_inst_pe_1_0_0_U6 ( .A(npu_inst_pe_1_0_0_n11), .Z(
        npu_inst_pe_1_0_0_n9) );
  BUF_X1 npu_inst_pe_1_0_0_U5 ( .A(npu_inst_pe_1_0_0_n11), .Z(
        npu_inst_pe_1_0_0_n8) );
  NOR2_X1 npu_inst_pe_1_0_0_U4 ( .A1(npu_inst_pe_1_0_0_int_q_weight_0_), .A2(
        npu_inst_pe_1_0_0_n1), .ZN(npu_inst_pe_1_0_0_n76) );
  NOR2_X1 npu_inst_pe_1_0_0_U3 ( .A1(npu_inst_pe_1_0_0_n27), .A2(
        npu_inst_pe_1_0_0_n1), .ZN(npu_inst_pe_1_0_0_n77) );
  FA_X1 npu_inst_pe_1_0_0_sub_67_U2_1 ( .A(npu_inst_pe_1_0_0_int_q_acc_1_), 
        .B(npu_inst_pe_1_0_0_n13), .CI(npu_inst_pe_1_0_0_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_0_0_sub_67_carry_2_), .S(npu_inst_pe_1_0_0_N66) );
  FA_X1 npu_inst_pe_1_0_0_add_69_U1_1 ( .A(npu_inst_pe_1_0_0_int_q_acc_1_), 
        .B(npu_inst_pe_1_0_0_int_data_1_), .CI(
        npu_inst_pe_1_0_0_add_69_carry_1_), .CO(
        npu_inst_pe_1_0_0_add_69_carry_2_), .S(npu_inst_pe_1_0_0_N74) );
  NAND3_X1 npu_inst_pe_1_0_0_U109 ( .A1(npu_inst_pe_1_0_0_n5), .A2(
        npu_inst_pe_1_0_0_n6), .A3(npu_inst_pe_1_0_0_n7), .ZN(
        npu_inst_pe_1_0_0_n44) );
  NAND3_X1 npu_inst_pe_1_0_0_U108 ( .A1(npu_inst_pe_1_0_0_n4), .A2(
        npu_inst_pe_1_0_0_n6), .A3(npu_inst_pe_1_0_0_n7), .ZN(
        npu_inst_pe_1_0_0_n40) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_0_0_n33), .CK(
        npu_inst_pe_1_0_0_net4562), .RN(npu_inst_pe_1_0_0_n8), .Q(
        npu_inst_pe_1_0_0_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_0_0_n34), .CK(
        npu_inst_pe_1_0_0_net4562), .RN(npu_inst_pe_1_0_0_n8), .Q(
        npu_inst_pe_1_0_0_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_0_0_n35), .CK(
        npu_inst_pe_1_0_0_net4562), .RN(npu_inst_pe_1_0_0_n8), .Q(
        npu_inst_pe_1_0_0_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_0_0_n36), .CK(
        npu_inst_pe_1_0_0_net4562), .RN(npu_inst_pe_1_0_0_n8), .Q(
        npu_inst_pe_1_0_0_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_0_0_n98), .CK(
        npu_inst_pe_1_0_0_net4562), .RN(npu_inst_pe_1_0_0_n8), .Q(
        npu_inst_pe_1_0_0_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_0_0_n99), .CK(
        npu_inst_pe_1_0_0_net4562), .RN(npu_inst_pe_1_0_0_n8), .Q(
        npu_inst_pe_1_0_0_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_0_0_n32), .CK(
        npu_inst_pe_1_0_0_net4562), .RN(npu_inst_pe_1_0_0_n8), .Q(
        npu_inst_pe_1_0_0_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_0_0_n100), 
        .CK(npu_inst_pe_1_0_0_net4562), .RN(npu_inst_pe_1_0_0_n8), .Q(
        npu_inst_pe_1_0_0_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_weight_reg_0_ ( .D(npu_inst_n113), .CK(
        npu_inst_pe_1_0_0_net4568), .RN(npu_inst_pe_1_0_0_n8), .Q(
        npu_inst_pe_1_0_0_int_q_weight_0_), .QN(npu_inst_pe_1_0_0_n27) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_weight_reg_1_ ( .D(npu_inst_n119), .CK(
        npu_inst_pe_1_0_0_net4568), .RN(npu_inst_pe_1_0_0_n8), .Q(
        npu_inst_pe_1_0_0_int_q_weight_1_), .QN(npu_inst_pe_1_0_0_n26) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_0_0_n112), 
        .CK(npu_inst_pe_1_0_0_net4568), .RN(npu_inst_pe_1_0_0_n8), .Q(
        npu_inst_pe_1_0_0_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_0_0_n106), 
        .CK(npu_inst_pe_1_0_0_net4568), .RN(npu_inst_pe_1_0_0_n8), .Q(
        npu_inst_pe_1_0_0_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_0_0_n111), 
        .CK(npu_inst_pe_1_0_0_net4568), .RN(npu_inst_pe_1_0_0_n9), .Q(
        npu_inst_pe_1_0_0_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_0_0_n105), 
        .CK(npu_inst_pe_1_0_0_net4568), .RN(npu_inst_pe_1_0_0_n9), .Q(
        npu_inst_pe_1_0_0_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_0_0_n110), 
        .CK(npu_inst_pe_1_0_0_net4568), .RN(npu_inst_pe_1_0_0_n9), .Q(
        npu_inst_pe_1_0_0_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_0_0_n104), 
        .CK(npu_inst_pe_1_0_0_net4568), .RN(npu_inst_pe_1_0_0_n9), .Q(
        npu_inst_pe_1_0_0_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_0_0_n109), 
        .CK(npu_inst_pe_1_0_0_net4568), .RN(npu_inst_pe_1_0_0_n9), .Q(
        npu_inst_pe_1_0_0_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_0_0_n103), 
        .CK(npu_inst_pe_1_0_0_net4568), .RN(npu_inst_pe_1_0_0_n9), .Q(
        npu_inst_pe_1_0_0_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_0_0_n108), 
        .CK(npu_inst_pe_1_0_0_net4568), .RN(npu_inst_pe_1_0_0_n9), .Q(
        npu_inst_pe_1_0_0_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_0_0_n102), 
        .CK(npu_inst_pe_1_0_0_net4568), .RN(npu_inst_pe_1_0_0_n9), .Q(
        npu_inst_pe_1_0_0_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_0_0_n107), 
        .CK(npu_inst_pe_1_0_0_net4568), .RN(npu_inst_pe_1_0_0_n9), .Q(
        npu_inst_pe_1_0_0_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_0_0_n101), 
        .CK(npu_inst_pe_1_0_0_net4568), .RN(npu_inst_pe_1_0_0_n9), .Q(
        npu_inst_pe_1_0_0_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_0_0_n86), 
        .CK(npu_inst_pe_1_0_0_net4568), .RN(npu_inst_pe_1_0_0_n9), .Q(
        npu_inst_pe_1_0_0_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_0_0_n87), 
        .CK(npu_inst_pe_1_0_0_net4568), .RN(npu_inst_pe_1_0_0_n9), .Q(
        npu_inst_pe_1_0_0_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_0_0_n88), 
        .CK(npu_inst_pe_1_0_0_net4568), .RN(npu_inst_pe_1_0_0_n10), .Q(
        npu_inst_pe_1_0_0_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_0_0_n89), 
        .CK(npu_inst_pe_1_0_0_net4568), .RN(npu_inst_pe_1_0_0_n10), .Q(
        npu_inst_pe_1_0_0_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_0_0_n90), 
        .CK(npu_inst_pe_1_0_0_net4568), .RN(npu_inst_pe_1_0_0_n10), .Q(
        npu_inst_pe_1_0_0_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_0_0_n91), 
        .CK(npu_inst_pe_1_0_0_net4568), .RN(npu_inst_pe_1_0_0_n10), .Q(
        npu_inst_pe_1_0_0_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_0_0_n92), 
        .CK(npu_inst_pe_1_0_0_net4568), .RN(npu_inst_pe_1_0_0_n10), .Q(
        npu_inst_pe_1_0_0_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_0_0_n93), 
        .CK(npu_inst_pe_1_0_0_net4568), .RN(npu_inst_pe_1_0_0_n10), .Q(
        npu_inst_pe_1_0_0_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_0_0_n94), 
        .CK(npu_inst_pe_1_0_0_net4568), .RN(npu_inst_pe_1_0_0_n10), .Q(
        npu_inst_pe_1_0_0_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_0_0_n95), 
        .CK(npu_inst_pe_1_0_0_net4568), .RN(npu_inst_pe_1_0_0_n10), .Q(
        npu_inst_pe_1_0_0_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_0_0_n96), 
        .CK(npu_inst_pe_1_0_0_net4568), .RN(npu_inst_pe_1_0_0_n10), .Q(
        npu_inst_pe_1_0_0_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_0_0_n97), 
        .CK(npu_inst_pe_1_0_0_net4568), .RN(npu_inst_pe_1_0_0_n10), .Q(
        npu_inst_pe_1_0_0_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_0_0_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_0_0_N84), .SE(1'b0), .GCK(npu_inst_pe_1_0_0_net4562) );
  CLKGATETST_X1 npu_inst_pe_1_0_0_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n66), .SE(1'b0), .GCK(npu_inst_pe_1_0_0_net4568) );
  MUX2_X1 npu_inst_pe_1_0_1_U160 ( .A(npu_inst_pe_1_0_1_n30), .B(
        npu_inst_pe_1_0_1_n25), .S(npu_inst_pe_1_0_1_n6), .Z(
        npu_inst_pe_1_0_1_N93) );
  MUX2_X1 npu_inst_pe_1_0_1_U159 ( .A(npu_inst_pe_1_0_1_n29), .B(
        npu_inst_pe_1_0_1_n28), .S(npu_inst_n80), .Z(npu_inst_pe_1_0_1_n30) );
  MUX2_X1 npu_inst_pe_1_0_1_U158 ( .A(npu_inst_pe_1_0_1_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_0_1_int_q_reg_v_1__0_), .S(npu_inst_n72), .Z(
        npu_inst_pe_1_0_1_n29) );
  MUX2_X1 npu_inst_pe_1_0_1_U157 ( .A(npu_inst_pe_1_0_1_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_0_1_int_q_reg_v_3__0_), .S(npu_inst_n72), .Z(
        npu_inst_pe_1_0_1_n28) );
  MUX2_X1 npu_inst_pe_1_0_1_U156 ( .A(npu_inst_pe_1_0_1_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_0_1_int_q_reg_v_5__0_), .S(npu_inst_n72), .Z(
        npu_inst_pe_1_0_1_n25) );
  MUX2_X1 npu_inst_pe_1_0_1_U155 ( .A(npu_inst_pe_1_0_1_n24), .B(
        npu_inst_pe_1_0_1_n21), .S(npu_inst_pe_1_0_1_n6), .Z(
        npu_inst_pe_1_0_1_N94) );
  MUX2_X1 npu_inst_pe_1_0_1_U154 ( .A(npu_inst_pe_1_0_1_n23), .B(
        npu_inst_pe_1_0_1_n22), .S(npu_inst_n80), .Z(npu_inst_pe_1_0_1_n24) );
  MUX2_X1 npu_inst_pe_1_0_1_U153 ( .A(npu_inst_pe_1_0_1_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_0_1_int_q_reg_v_1__1_), .S(npu_inst_n72), .Z(
        npu_inst_pe_1_0_1_n23) );
  MUX2_X1 npu_inst_pe_1_0_1_U152 ( .A(npu_inst_pe_1_0_1_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_0_1_int_q_reg_v_3__1_), .S(npu_inst_n72), .Z(
        npu_inst_pe_1_0_1_n22) );
  MUX2_X1 npu_inst_pe_1_0_1_U151 ( .A(npu_inst_pe_1_0_1_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_0_1_int_q_reg_v_5__1_), .S(npu_inst_n72), .Z(
        npu_inst_pe_1_0_1_n21) );
  MUX2_X1 npu_inst_pe_1_0_1_U150 ( .A(npu_inst_pe_1_0_1_n20), .B(
        npu_inst_pe_1_0_1_n17), .S(npu_inst_pe_1_0_1_n6), .Z(
        npu_inst_int_data_x_0__1__1_) );
  MUX2_X1 npu_inst_pe_1_0_1_U149 ( .A(npu_inst_pe_1_0_1_n19), .B(
        npu_inst_pe_1_0_1_n18), .S(npu_inst_n80), .Z(npu_inst_pe_1_0_1_n20) );
  MUX2_X1 npu_inst_pe_1_0_1_U148 ( .A(npu_inst_pe_1_0_1_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_0_1_int_q_reg_h_1__1_), .S(npu_inst_n72), .Z(
        npu_inst_pe_1_0_1_n19) );
  MUX2_X1 npu_inst_pe_1_0_1_U147 ( .A(npu_inst_pe_1_0_1_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_0_1_int_q_reg_h_3__1_), .S(npu_inst_n72), .Z(
        npu_inst_pe_1_0_1_n18) );
  MUX2_X1 npu_inst_pe_1_0_1_U146 ( .A(npu_inst_pe_1_0_1_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_0_1_int_q_reg_h_5__1_), .S(npu_inst_n72), .Z(
        npu_inst_pe_1_0_1_n17) );
  MUX2_X1 npu_inst_pe_1_0_1_U145 ( .A(npu_inst_pe_1_0_1_n16), .B(
        npu_inst_pe_1_0_1_n13), .S(npu_inst_pe_1_0_1_n6), .Z(
        npu_inst_int_data_x_0__1__0_) );
  MUX2_X1 npu_inst_pe_1_0_1_U144 ( .A(npu_inst_pe_1_0_1_n15), .B(
        npu_inst_pe_1_0_1_n14), .S(npu_inst_n80), .Z(npu_inst_pe_1_0_1_n16) );
  MUX2_X1 npu_inst_pe_1_0_1_U143 ( .A(npu_inst_pe_1_0_1_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_0_1_int_q_reg_h_1__0_), .S(npu_inst_n72), .Z(
        npu_inst_pe_1_0_1_n15) );
  MUX2_X1 npu_inst_pe_1_0_1_U142 ( .A(npu_inst_pe_1_0_1_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_0_1_int_q_reg_h_3__0_), .S(npu_inst_n72), .Z(
        npu_inst_pe_1_0_1_n14) );
  MUX2_X1 npu_inst_pe_1_0_1_U141 ( .A(npu_inst_pe_1_0_1_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_0_1_int_q_reg_h_5__0_), .S(npu_inst_n72), .Z(
        npu_inst_pe_1_0_1_n13) );
  XOR2_X1 npu_inst_pe_1_0_1_U140 ( .A(npu_inst_pe_1_0_1_int_data_0_), .B(
        npu_inst_pe_1_0_1_int_q_acc_0_), .Z(npu_inst_pe_1_0_1_N73) );
  AND2_X1 npu_inst_pe_1_0_1_U139 ( .A1(npu_inst_pe_1_0_1_int_q_acc_0_), .A2(
        npu_inst_pe_1_0_1_int_data_0_), .ZN(npu_inst_pe_1_0_1_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_0_1_U138 ( .A(npu_inst_pe_1_0_1_int_q_acc_0_), .B(
        npu_inst_pe_1_0_1_n11), .ZN(npu_inst_pe_1_0_1_N65) );
  OR2_X1 npu_inst_pe_1_0_1_U137 ( .A1(npu_inst_pe_1_0_1_n11), .A2(
        npu_inst_pe_1_0_1_int_q_acc_0_), .ZN(npu_inst_pe_1_0_1_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_0_1_U136 ( .A(npu_inst_pe_1_0_1_int_q_acc_2_), .B(
        npu_inst_pe_1_0_1_add_69_carry_2_), .Z(npu_inst_pe_1_0_1_N75) );
  AND2_X1 npu_inst_pe_1_0_1_U135 ( .A1(npu_inst_pe_1_0_1_add_69_carry_2_), 
        .A2(npu_inst_pe_1_0_1_int_q_acc_2_), .ZN(
        npu_inst_pe_1_0_1_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_0_1_U134 ( .A(npu_inst_pe_1_0_1_int_q_acc_3_), .B(
        npu_inst_pe_1_0_1_add_69_carry_3_), .Z(npu_inst_pe_1_0_1_N76) );
  AND2_X1 npu_inst_pe_1_0_1_U133 ( .A1(npu_inst_pe_1_0_1_add_69_carry_3_), 
        .A2(npu_inst_pe_1_0_1_int_q_acc_3_), .ZN(
        npu_inst_pe_1_0_1_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_0_1_U132 ( .A(npu_inst_pe_1_0_1_int_q_acc_4_), .B(
        npu_inst_pe_1_0_1_add_69_carry_4_), .Z(npu_inst_pe_1_0_1_N77) );
  AND2_X1 npu_inst_pe_1_0_1_U131 ( .A1(npu_inst_pe_1_0_1_add_69_carry_4_), 
        .A2(npu_inst_pe_1_0_1_int_q_acc_4_), .ZN(
        npu_inst_pe_1_0_1_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_0_1_U130 ( .A(npu_inst_pe_1_0_1_int_q_acc_5_), .B(
        npu_inst_pe_1_0_1_add_69_carry_5_), .Z(npu_inst_pe_1_0_1_N78) );
  AND2_X1 npu_inst_pe_1_0_1_U129 ( .A1(npu_inst_pe_1_0_1_add_69_carry_5_), 
        .A2(npu_inst_pe_1_0_1_int_q_acc_5_), .ZN(
        npu_inst_pe_1_0_1_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_0_1_U128 ( .A(npu_inst_pe_1_0_1_int_q_acc_6_), .B(
        npu_inst_pe_1_0_1_add_69_carry_6_), .Z(npu_inst_pe_1_0_1_N79) );
  AND2_X1 npu_inst_pe_1_0_1_U127 ( .A1(npu_inst_pe_1_0_1_add_69_carry_6_), 
        .A2(npu_inst_pe_1_0_1_int_q_acc_6_), .ZN(
        npu_inst_pe_1_0_1_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_0_1_U126 ( .A(npu_inst_pe_1_0_1_int_q_acc_7_), .B(
        npu_inst_pe_1_0_1_add_69_carry_7_), .Z(npu_inst_pe_1_0_1_N80) );
  XNOR2_X1 npu_inst_pe_1_0_1_U125 ( .A(npu_inst_pe_1_0_1_sub_67_carry_2_), .B(
        npu_inst_pe_1_0_1_int_q_acc_2_), .ZN(npu_inst_pe_1_0_1_N67) );
  OR2_X1 npu_inst_pe_1_0_1_U124 ( .A1(npu_inst_pe_1_0_1_int_q_acc_2_), .A2(
        npu_inst_pe_1_0_1_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_0_1_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_0_1_U123 ( .A(npu_inst_pe_1_0_1_sub_67_carry_3_), .B(
        npu_inst_pe_1_0_1_int_q_acc_3_), .ZN(npu_inst_pe_1_0_1_N68) );
  OR2_X1 npu_inst_pe_1_0_1_U122 ( .A1(npu_inst_pe_1_0_1_int_q_acc_3_), .A2(
        npu_inst_pe_1_0_1_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_0_1_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_0_1_U121 ( .A(npu_inst_pe_1_0_1_sub_67_carry_4_), .B(
        npu_inst_pe_1_0_1_int_q_acc_4_), .ZN(npu_inst_pe_1_0_1_N69) );
  OR2_X1 npu_inst_pe_1_0_1_U120 ( .A1(npu_inst_pe_1_0_1_int_q_acc_4_), .A2(
        npu_inst_pe_1_0_1_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_0_1_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_0_1_U119 ( .A(npu_inst_pe_1_0_1_sub_67_carry_5_), .B(
        npu_inst_pe_1_0_1_int_q_acc_5_), .ZN(npu_inst_pe_1_0_1_N70) );
  OR2_X1 npu_inst_pe_1_0_1_U118 ( .A1(npu_inst_pe_1_0_1_int_q_acc_5_), .A2(
        npu_inst_pe_1_0_1_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_0_1_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_0_1_U117 ( .A(npu_inst_pe_1_0_1_sub_67_carry_6_), .B(
        npu_inst_pe_1_0_1_int_q_acc_6_), .ZN(npu_inst_pe_1_0_1_N71) );
  OR2_X1 npu_inst_pe_1_0_1_U116 ( .A1(npu_inst_pe_1_0_1_int_q_acc_6_), .A2(
        npu_inst_pe_1_0_1_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_0_1_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_0_1_U115 ( .A(npu_inst_pe_1_0_1_int_q_acc_7_), .B(
        npu_inst_pe_1_0_1_sub_67_carry_7_), .ZN(npu_inst_pe_1_0_1_N72) );
  INV_X1 npu_inst_pe_1_0_1_U114 ( .A(npu_inst_n80), .ZN(npu_inst_pe_1_0_1_n5)
         );
  INV_X1 npu_inst_pe_1_0_1_U113 ( .A(npu_inst_n60), .ZN(npu_inst_pe_1_0_1_n3)
         );
  AOI22_X1 npu_inst_pe_1_0_1_U112 ( .A1(npu_inst_int_data_y_1__1__0_), .A2(
        npu_inst_pe_1_0_1_n58), .B1(npu_inst_pe_1_0_1_n117), .B2(
        npu_inst_pe_1_0_1_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_0_1_n57) );
  INV_X1 npu_inst_pe_1_0_1_U111 ( .A(npu_inst_pe_1_0_1_n57), .ZN(
        npu_inst_pe_1_0_1_n106) );
  AOI22_X1 npu_inst_pe_1_0_1_U110 ( .A1(npu_inst_int_data_y_1__1__0_), .A2(
        npu_inst_pe_1_0_1_n54), .B1(npu_inst_pe_1_0_1_n116), .B2(
        npu_inst_pe_1_0_1_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_0_1_n53) );
  INV_X1 npu_inst_pe_1_0_1_U107 ( .A(npu_inst_pe_1_0_1_n53), .ZN(
        npu_inst_pe_1_0_1_n107) );
  AOI22_X1 npu_inst_pe_1_0_1_U106 ( .A1(npu_inst_int_data_y_1__1__0_), .A2(
        npu_inst_pe_1_0_1_n50), .B1(npu_inst_pe_1_0_1_n115), .B2(
        npu_inst_pe_1_0_1_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_0_1_n49) );
  INV_X1 npu_inst_pe_1_0_1_U105 ( .A(npu_inst_pe_1_0_1_n49), .ZN(
        npu_inst_pe_1_0_1_n108) );
  AOI22_X1 npu_inst_pe_1_0_1_U104 ( .A1(npu_inst_int_data_y_1__1__0_), .A2(
        npu_inst_pe_1_0_1_n46), .B1(npu_inst_pe_1_0_1_n114), .B2(
        npu_inst_pe_1_0_1_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_0_1_n45) );
  INV_X1 npu_inst_pe_1_0_1_U103 ( .A(npu_inst_pe_1_0_1_n45), .ZN(
        npu_inst_pe_1_0_1_n109) );
  AOI22_X1 npu_inst_pe_1_0_1_U102 ( .A1(npu_inst_int_data_y_1__1__0_), .A2(
        npu_inst_pe_1_0_1_n42), .B1(npu_inst_pe_1_0_1_n113), .B2(
        npu_inst_pe_1_0_1_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_0_1_n41) );
  INV_X1 npu_inst_pe_1_0_1_U101 ( .A(npu_inst_pe_1_0_1_n41), .ZN(
        npu_inst_pe_1_0_1_n110) );
  AOI22_X1 npu_inst_pe_1_0_1_U100 ( .A1(npu_inst_int_data_y_1__1__1_), .A2(
        npu_inst_pe_1_0_1_n58), .B1(npu_inst_pe_1_0_1_n117), .B2(
        npu_inst_pe_1_0_1_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_0_1_n59) );
  INV_X1 npu_inst_pe_1_0_1_U99 ( .A(npu_inst_pe_1_0_1_n59), .ZN(
        npu_inst_pe_1_0_1_n100) );
  AOI22_X1 npu_inst_pe_1_0_1_U98 ( .A1(npu_inst_int_data_y_1__1__1_), .A2(
        npu_inst_pe_1_0_1_n54), .B1(npu_inst_pe_1_0_1_n116), .B2(
        npu_inst_pe_1_0_1_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_0_1_n55) );
  INV_X1 npu_inst_pe_1_0_1_U97 ( .A(npu_inst_pe_1_0_1_n55), .ZN(
        npu_inst_pe_1_0_1_n101) );
  AOI22_X1 npu_inst_pe_1_0_1_U96 ( .A1(npu_inst_int_data_y_1__1__1_), .A2(
        npu_inst_pe_1_0_1_n50), .B1(npu_inst_pe_1_0_1_n115), .B2(
        npu_inst_pe_1_0_1_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_0_1_n51) );
  INV_X1 npu_inst_pe_1_0_1_U95 ( .A(npu_inst_pe_1_0_1_n51), .ZN(
        npu_inst_pe_1_0_1_n102) );
  AOI22_X1 npu_inst_pe_1_0_1_U94 ( .A1(npu_inst_int_data_y_1__1__1_), .A2(
        npu_inst_pe_1_0_1_n46), .B1(npu_inst_pe_1_0_1_n114), .B2(
        npu_inst_pe_1_0_1_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_0_1_n47) );
  INV_X1 npu_inst_pe_1_0_1_U93 ( .A(npu_inst_pe_1_0_1_n47), .ZN(
        npu_inst_pe_1_0_1_n103) );
  AOI22_X1 npu_inst_pe_1_0_1_U92 ( .A1(npu_inst_int_data_y_1__1__1_), .A2(
        npu_inst_pe_1_0_1_n42), .B1(npu_inst_pe_1_0_1_n113), .B2(
        npu_inst_pe_1_0_1_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_0_1_n43) );
  INV_X1 npu_inst_pe_1_0_1_U91 ( .A(npu_inst_pe_1_0_1_n43), .ZN(
        npu_inst_pe_1_0_1_n104) );
  AOI22_X1 npu_inst_pe_1_0_1_U90 ( .A1(npu_inst_pe_1_0_1_n38), .A2(
        npu_inst_int_data_y_1__1__1_), .B1(npu_inst_pe_1_0_1_n112), .B2(
        npu_inst_pe_1_0_1_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_0_1_n39) );
  INV_X1 npu_inst_pe_1_0_1_U89 ( .A(npu_inst_pe_1_0_1_n39), .ZN(
        npu_inst_pe_1_0_1_n105) );
  AOI22_X1 npu_inst_pe_1_0_1_U88 ( .A1(npu_inst_pe_1_0_1_n38), .A2(
        npu_inst_int_data_y_1__1__0_), .B1(npu_inst_pe_1_0_1_n112), .B2(
        npu_inst_pe_1_0_1_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_0_1_n37) );
  INV_X1 npu_inst_pe_1_0_1_U87 ( .A(npu_inst_pe_1_0_1_n37), .ZN(
        npu_inst_pe_1_0_1_n111) );
  NAND2_X1 npu_inst_pe_1_0_1_U86 ( .A1(npu_inst_pe_1_0_1_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_0_1_n60), .ZN(npu_inst_pe_1_0_1_n74) );
  OAI21_X1 npu_inst_pe_1_0_1_U85 ( .B1(npu_inst_pe_1_0_1_n63), .B2(
        npu_inst_pe_1_0_1_n60), .A(npu_inst_pe_1_0_1_n74), .ZN(
        npu_inst_pe_1_0_1_n97) );
  NAND2_X1 npu_inst_pe_1_0_1_U84 ( .A1(npu_inst_pe_1_0_1_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_0_1_n60), .ZN(npu_inst_pe_1_0_1_n73) );
  OAI21_X1 npu_inst_pe_1_0_1_U83 ( .B1(npu_inst_pe_1_0_1_n61), .B2(
        npu_inst_pe_1_0_1_n60), .A(npu_inst_pe_1_0_1_n73), .ZN(
        npu_inst_pe_1_0_1_n96) );
  NAND2_X1 npu_inst_pe_1_0_1_U82 ( .A1(npu_inst_pe_1_0_1_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_0_1_n56), .ZN(npu_inst_pe_1_0_1_n72) );
  OAI21_X1 npu_inst_pe_1_0_1_U81 ( .B1(npu_inst_pe_1_0_1_n63), .B2(
        npu_inst_pe_1_0_1_n56), .A(npu_inst_pe_1_0_1_n72), .ZN(
        npu_inst_pe_1_0_1_n95) );
  NAND2_X1 npu_inst_pe_1_0_1_U80 ( .A1(npu_inst_pe_1_0_1_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_0_1_n56), .ZN(npu_inst_pe_1_0_1_n71) );
  OAI21_X1 npu_inst_pe_1_0_1_U79 ( .B1(npu_inst_pe_1_0_1_n61), .B2(
        npu_inst_pe_1_0_1_n56), .A(npu_inst_pe_1_0_1_n71), .ZN(
        npu_inst_pe_1_0_1_n94) );
  NAND2_X1 npu_inst_pe_1_0_1_U78 ( .A1(npu_inst_pe_1_0_1_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_0_1_n52), .ZN(npu_inst_pe_1_0_1_n70) );
  OAI21_X1 npu_inst_pe_1_0_1_U77 ( .B1(npu_inst_pe_1_0_1_n63), .B2(
        npu_inst_pe_1_0_1_n52), .A(npu_inst_pe_1_0_1_n70), .ZN(
        npu_inst_pe_1_0_1_n93) );
  NAND2_X1 npu_inst_pe_1_0_1_U76 ( .A1(npu_inst_pe_1_0_1_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_0_1_n52), .ZN(npu_inst_pe_1_0_1_n69) );
  OAI21_X1 npu_inst_pe_1_0_1_U75 ( .B1(npu_inst_pe_1_0_1_n61), .B2(
        npu_inst_pe_1_0_1_n52), .A(npu_inst_pe_1_0_1_n69), .ZN(
        npu_inst_pe_1_0_1_n92) );
  NAND2_X1 npu_inst_pe_1_0_1_U74 ( .A1(npu_inst_pe_1_0_1_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_0_1_n48), .ZN(npu_inst_pe_1_0_1_n68) );
  OAI21_X1 npu_inst_pe_1_0_1_U73 ( .B1(npu_inst_pe_1_0_1_n63), .B2(
        npu_inst_pe_1_0_1_n48), .A(npu_inst_pe_1_0_1_n68), .ZN(
        npu_inst_pe_1_0_1_n91) );
  NAND2_X1 npu_inst_pe_1_0_1_U72 ( .A1(npu_inst_pe_1_0_1_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_0_1_n48), .ZN(npu_inst_pe_1_0_1_n67) );
  OAI21_X1 npu_inst_pe_1_0_1_U71 ( .B1(npu_inst_pe_1_0_1_n61), .B2(
        npu_inst_pe_1_0_1_n48), .A(npu_inst_pe_1_0_1_n67), .ZN(
        npu_inst_pe_1_0_1_n90) );
  NAND2_X1 npu_inst_pe_1_0_1_U70 ( .A1(npu_inst_pe_1_0_1_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_0_1_n44), .ZN(npu_inst_pe_1_0_1_n66) );
  OAI21_X1 npu_inst_pe_1_0_1_U69 ( .B1(npu_inst_pe_1_0_1_n63), .B2(
        npu_inst_pe_1_0_1_n44), .A(npu_inst_pe_1_0_1_n66), .ZN(
        npu_inst_pe_1_0_1_n89) );
  NAND2_X1 npu_inst_pe_1_0_1_U68 ( .A1(npu_inst_pe_1_0_1_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_0_1_n44), .ZN(npu_inst_pe_1_0_1_n65) );
  OAI21_X1 npu_inst_pe_1_0_1_U67 ( .B1(npu_inst_pe_1_0_1_n61), .B2(
        npu_inst_pe_1_0_1_n44), .A(npu_inst_pe_1_0_1_n65), .ZN(
        npu_inst_pe_1_0_1_n88) );
  NAND2_X1 npu_inst_pe_1_0_1_U66 ( .A1(npu_inst_pe_1_0_1_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_0_1_n40), .ZN(npu_inst_pe_1_0_1_n64) );
  OAI21_X1 npu_inst_pe_1_0_1_U65 ( .B1(npu_inst_pe_1_0_1_n63), .B2(
        npu_inst_pe_1_0_1_n40), .A(npu_inst_pe_1_0_1_n64), .ZN(
        npu_inst_pe_1_0_1_n87) );
  NAND2_X1 npu_inst_pe_1_0_1_U64 ( .A1(npu_inst_pe_1_0_1_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_0_1_n40), .ZN(npu_inst_pe_1_0_1_n62) );
  OAI21_X1 npu_inst_pe_1_0_1_U63 ( .B1(npu_inst_pe_1_0_1_n61), .B2(
        npu_inst_pe_1_0_1_n40), .A(npu_inst_pe_1_0_1_n62), .ZN(
        npu_inst_pe_1_0_1_n86) );
  AND2_X1 npu_inst_pe_1_0_1_U62 ( .A1(npu_inst_pe_1_0_1_int_q_acc_2_), .A2(
        npu_inst_pe_1_0_1_n1), .ZN(int_o_data_npu[50]) );
  AND2_X1 npu_inst_pe_1_0_1_U61 ( .A1(npu_inst_pe_1_0_1_int_q_acc_3_), .A2(
        npu_inst_pe_1_0_1_n2), .ZN(int_o_data_npu[51]) );
  NOR3_X1 npu_inst_pe_1_0_1_U60 ( .A1(npu_inst_pe_1_0_1_n26), .A2(npu_inst_n60), .A3(npu_inst_int_ckg[62]), .ZN(npu_inst_pe_1_0_1_n85) );
  OR2_X1 npu_inst_pe_1_0_1_U59 ( .A1(npu_inst_pe_1_0_1_n85), .A2(
        npu_inst_pe_1_0_1_n2), .ZN(npu_inst_pe_1_0_1_N84) );
  AND2_X1 npu_inst_pe_1_0_1_U58 ( .A1(npu_inst_pe_1_0_1_int_q_acc_6_), .A2(
        npu_inst_pe_1_0_1_n2), .ZN(int_o_data_npu[54]) );
  AND2_X1 npu_inst_pe_1_0_1_U57 ( .A1(npu_inst_pe_1_0_1_int_q_acc_5_), .A2(
        npu_inst_pe_1_0_1_n2), .ZN(int_o_data_npu[53]) );
  AND2_X1 npu_inst_pe_1_0_1_U56 ( .A1(npu_inst_pe_1_0_1_int_q_acc_4_), .A2(
        npu_inst_pe_1_0_1_n2), .ZN(int_o_data_npu[52]) );
  AOI222_X1 npu_inst_pe_1_0_1_U55 ( .A1(npu_inst_int_data_res_1__1__0_), .A2(
        npu_inst_pe_1_0_1_n1), .B1(npu_inst_pe_1_0_1_N73), .B2(
        npu_inst_pe_1_0_1_n76), .C1(npu_inst_pe_1_0_1_N65), .C2(
        npu_inst_pe_1_0_1_n77), .ZN(npu_inst_pe_1_0_1_n84) );
  INV_X1 npu_inst_pe_1_0_1_U54 ( .A(npu_inst_pe_1_0_1_n84), .ZN(
        npu_inst_pe_1_0_1_n99) );
  AOI222_X1 npu_inst_pe_1_0_1_U53 ( .A1(npu_inst_int_data_res_1__1__7_), .A2(
        npu_inst_pe_1_0_1_n1), .B1(npu_inst_pe_1_0_1_N80), .B2(
        npu_inst_pe_1_0_1_n76), .C1(npu_inst_pe_1_0_1_N72), .C2(
        npu_inst_pe_1_0_1_n77), .ZN(npu_inst_pe_1_0_1_n75) );
  INV_X1 npu_inst_pe_1_0_1_U52 ( .A(npu_inst_pe_1_0_1_n75), .ZN(
        npu_inst_pe_1_0_1_n31) );
  AOI222_X1 npu_inst_pe_1_0_1_U51 ( .A1(npu_inst_int_data_res_1__1__1_), .A2(
        npu_inst_pe_1_0_1_n1), .B1(npu_inst_pe_1_0_1_N74), .B2(
        npu_inst_pe_1_0_1_n76), .C1(npu_inst_pe_1_0_1_N66), .C2(
        npu_inst_pe_1_0_1_n77), .ZN(npu_inst_pe_1_0_1_n83) );
  INV_X1 npu_inst_pe_1_0_1_U50 ( .A(npu_inst_pe_1_0_1_n83), .ZN(
        npu_inst_pe_1_0_1_n98) );
  AOI222_X1 npu_inst_pe_1_0_1_U49 ( .A1(npu_inst_int_data_res_1__1__2_), .A2(
        npu_inst_pe_1_0_1_n1), .B1(npu_inst_pe_1_0_1_N75), .B2(
        npu_inst_pe_1_0_1_n76), .C1(npu_inst_pe_1_0_1_N67), .C2(
        npu_inst_pe_1_0_1_n77), .ZN(npu_inst_pe_1_0_1_n82) );
  INV_X1 npu_inst_pe_1_0_1_U48 ( .A(npu_inst_pe_1_0_1_n82), .ZN(
        npu_inst_pe_1_0_1_n36) );
  AOI222_X1 npu_inst_pe_1_0_1_U47 ( .A1(npu_inst_int_data_res_1__1__3_), .A2(
        npu_inst_pe_1_0_1_n1), .B1(npu_inst_pe_1_0_1_N76), .B2(
        npu_inst_pe_1_0_1_n76), .C1(npu_inst_pe_1_0_1_N68), .C2(
        npu_inst_pe_1_0_1_n77), .ZN(npu_inst_pe_1_0_1_n81) );
  INV_X1 npu_inst_pe_1_0_1_U46 ( .A(npu_inst_pe_1_0_1_n81), .ZN(
        npu_inst_pe_1_0_1_n35) );
  AOI222_X1 npu_inst_pe_1_0_1_U45 ( .A1(npu_inst_int_data_res_1__1__4_), .A2(
        npu_inst_pe_1_0_1_n1), .B1(npu_inst_pe_1_0_1_N77), .B2(
        npu_inst_pe_1_0_1_n76), .C1(npu_inst_pe_1_0_1_N69), .C2(
        npu_inst_pe_1_0_1_n77), .ZN(npu_inst_pe_1_0_1_n80) );
  INV_X1 npu_inst_pe_1_0_1_U44 ( .A(npu_inst_pe_1_0_1_n80), .ZN(
        npu_inst_pe_1_0_1_n34) );
  AOI222_X1 npu_inst_pe_1_0_1_U43 ( .A1(npu_inst_int_data_res_1__1__5_), .A2(
        npu_inst_pe_1_0_1_n1), .B1(npu_inst_pe_1_0_1_N78), .B2(
        npu_inst_pe_1_0_1_n76), .C1(npu_inst_pe_1_0_1_N70), .C2(
        npu_inst_pe_1_0_1_n77), .ZN(npu_inst_pe_1_0_1_n79) );
  INV_X1 npu_inst_pe_1_0_1_U42 ( .A(npu_inst_pe_1_0_1_n79), .ZN(
        npu_inst_pe_1_0_1_n33) );
  AOI222_X1 npu_inst_pe_1_0_1_U41 ( .A1(npu_inst_int_data_res_1__1__6_), .A2(
        npu_inst_pe_1_0_1_n1), .B1(npu_inst_pe_1_0_1_N79), .B2(
        npu_inst_pe_1_0_1_n76), .C1(npu_inst_pe_1_0_1_N71), .C2(
        npu_inst_pe_1_0_1_n77), .ZN(npu_inst_pe_1_0_1_n78) );
  INV_X1 npu_inst_pe_1_0_1_U40 ( .A(npu_inst_pe_1_0_1_n78), .ZN(
        npu_inst_pe_1_0_1_n32) );
  INV_X1 npu_inst_pe_1_0_1_U39 ( .A(npu_inst_pe_1_0_1_int_data_1_), .ZN(
        npu_inst_pe_1_0_1_n12) );
  AND2_X1 npu_inst_pe_1_0_1_U38 ( .A1(npu_inst_int_data_x_0__1__1_), .A2(
        npu_inst_pe_1_0_1_int_q_weight_1_), .ZN(npu_inst_pe_1_0_1_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_0_1_U37 ( .A1(npu_inst_int_data_x_0__1__0_), .A2(
        npu_inst_pe_1_0_1_int_q_weight_1_), .ZN(npu_inst_pe_1_0_1_int_data_0_)
         );
  AND2_X1 npu_inst_pe_1_0_1_U36 ( .A1(npu_inst_pe_1_0_1_n2), .A2(
        npu_inst_pe_1_0_1_int_q_acc_7_), .ZN(int_o_data_npu[55]) );
  AND2_X1 npu_inst_pe_1_0_1_U35 ( .A1(npu_inst_pe_1_0_1_int_q_acc_1_), .A2(
        npu_inst_pe_1_0_1_n1), .ZN(int_o_data_npu[49]) );
  AND2_X1 npu_inst_pe_1_0_1_U34 ( .A1(npu_inst_pe_1_0_1_int_q_acc_0_), .A2(
        npu_inst_pe_1_0_1_n1), .ZN(int_o_data_npu[48]) );
  AND2_X1 npu_inst_pe_1_0_1_U33 ( .A1(npu_inst_pe_1_0_1_N93), .A2(npu_inst_n60), .ZN(npu_inst_pe_1_0_1_o_data_v_0_) );
  AND2_X1 npu_inst_pe_1_0_1_U32 ( .A1(npu_inst_n60), .A2(npu_inst_pe_1_0_1_N94), .ZN(npu_inst_pe_1_0_1_o_data_v_1_) );
  AOI22_X1 npu_inst_pe_1_0_1_U31 ( .A1(npu_inst_n60), .A2(
        npu_inst_int_data_y_1__1__1_), .B1(npu_inst_pe_1_0_1_n3), .B2(
        npu_inst_int_data_x_0__2__1_), .ZN(npu_inst_pe_1_0_1_n63) );
  AOI22_X1 npu_inst_pe_1_0_1_U30 ( .A1(npu_inst_n60), .A2(
        npu_inst_int_data_y_1__1__0_), .B1(npu_inst_pe_1_0_1_n3), .B2(
        npu_inst_int_data_x_0__2__0_), .ZN(npu_inst_pe_1_0_1_n61) );
  INV_X1 npu_inst_pe_1_0_1_U29 ( .A(npu_inst_pe_1_0_1_int_data_0_), .ZN(
        npu_inst_pe_1_0_1_n11) );
  INV_X1 npu_inst_pe_1_0_1_U28 ( .A(npu_inst_n72), .ZN(npu_inst_pe_1_0_1_n4)
         );
  OR3_X1 npu_inst_pe_1_0_1_U27 ( .A1(npu_inst_n80), .A2(npu_inst_pe_1_0_1_n6), 
        .A3(npu_inst_pe_1_0_1_n4), .ZN(npu_inst_pe_1_0_1_n56) );
  OR3_X1 npu_inst_pe_1_0_1_U26 ( .A1(npu_inst_pe_1_0_1_n4), .A2(
        npu_inst_pe_1_0_1_n6), .A3(npu_inst_pe_1_0_1_n5), .ZN(
        npu_inst_pe_1_0_1_n48) );
  OR3_X1 npu_inst_pe_1_0_1_U25 ( .A1(npu_inst_n72), .A2(npu_inst_pe_1_0_1_n6), 
        .A3(npu_inst_pe_1_0_1_n5), .ZN(npu_inst_pe_1_0_1_n52) );
  OR3_X1 npu_inst_pe_1_0_1_U24 ( .A1(npu_inst_n80), .A2(npu_inst_pe_1_0_1_n6), 
        .A3(npu_inst_n72), .ZN(npu_inst_pe_1_0_1_n60) );
  NOR2_X1 npu_inst_pe_1_0_1_U23 ( .A1(npu_inst_pe_1_0_1_n60), .A2(
        npu_inst_pe_1_0_1_n3), .ZN(npu_inst_pe_1_0_1_n58) );
  NOR2_X1 npu_inst_pe_1_0_1_U22 ( .A1(npu_inst_pe_1_0_1_n56), .A2(
        npu_inst_pe_1_0_1_n3), .ZN(npu_inst_pe_1_0_1_n54) );
  NOR2_X1 npu_inst_pe_1_0_1_U21 ( .A1(npu_inst_pe_1_0_1_n52), .A2(
        npu_inst_pe_1_0_1_n3), .ZN(npu_inst_pe_1_0_1_n50) );
  NOR2_X1 npu_inst_pe_1_0_1_U20 ( .A1(npu_inst_pe_1_0_1_n48), .A2(
        npu_inst_pe_1_0_1_n3), .ZN(npu_inst_pe_1_0_1_n46) );
  NOR2_X1 npu_inst_pe_1_0_1_U19 ( .A1(npu_inst_pe_1_0_1_n40), .A2(
        npu_inst_pe_1_0_1_n3), .ZN(npu_inst_pe_1_0_1_n38) );
  NOR2_X1 npu_inst_pe_1_0_1_U18 ( .A1(npu_inst_pe_1_0_1_n44), .A2(
        npu_inst_pe_1_0_1_n3), .ZN(npu_inst_pe_1_0_1_n42) );
  BUF_X1 npu_inst_pe_1_0_1_U17 ( .A(npu_inst_n107), .Z(npu_inst_pe_1_0_1_n6)
         );
  INV_X1 npu_inst_pe_1_0_1_U16 ( .A(npu_inst_n127), .ZN(npu_inst_pe_1_0_1_n10)
         );
  INV_X1 npu_inst_pe_1_0_1_U15 ( .A(npu_inst_pe_1_0_1_n38), .ZN(
        npu_inst_pe_1_0_1_n112) );
  INV_X1 npu_inst_pe_1_0_1_U14 ( .A(npu_inst_pe_1_0_1_n58), .ZN(
        npu_inst_pe_1_0_1_n117) );
  INV_X1 npu_inst_pe_1_0_1_U13 ( .A(npu_inst_pe_1_0_1_n54), .ZN(
        npu_inst_pe_1_0_1_n116) );
  INV_X1 npu_inst_pe_1_0_1_U12 ( .A(npu_inst_pe_1_0_1_n50), .ZN(
        npu_inst_pe_1_0_1_n115) );
  INV_X1 npu_inst_pe_1_0_1_U11 ( .A(npu_inst_pe_1_0_1_n46), .ZN(
        npu_inst_pe_1_0_1_n114) );
  INV_X1 npu_inst_pe_1_0_1_U10 ( .A(npu_inst_pe_1_0_1_n42), .ZN(
        npu_inst_pe_1_0_1_n113) );
  BUF_X1 npu_inst_pe_1_0_1_U9 ( .A(npu_inst_n38), .Z(npu_inst_pe_1_0_1_n2) );
  BUF_X1 npu_inst_pe_1_0_1_U8 ( .A(npu_inst_n38), .Z(npu_inst_pe_1_0_1_n1) );
  BUF_X1 npu_inst_pe_1_0_1_U7 ( .A(npu_inst_pe_1_0_1_n10), .Z(
        npu_inst_pe_1_0_1_n9) );
  BUF_X1 npu_inst_pe_1_0_1_U6 ( .A(npu_inst_pe_1_0_1_n10), .Z(
        npu_inst_pe_1_0_1_n8) );
  BUF_X1 npu_inst_pe_1_0_1_U5 ( .A(npu_inst_pe_1_0_1_n10), .Z(
        npu_inst_pe_1_0_1_n7) );
  NOR2_X1 npu_inst_pe_1_0_1_U4 ( .A1(npu_inst_pe_1_0_1_int_q_weight_0_), .A2(
        npu_inst_pe_1_0_1_n1), .ZN(npu_inst_pe_1_0_1_n76) );
  NOR2_X1 npu_inst_pe_1_0_1_U3 ( .A1(npu_inst_pe_1_0_1_n27), .A2(
        npu_inst_pe_1_0_1_n1), .ZN(npu_inst_pe_1_0_1_n77) );
  FA_X1 npu_inst_pe_1_0_1_sub_67_U2_1 ( .A(npu_inst_pe_1_0_1_int_q_acc_1_), 
        .B(npu_inst_pe_1_0_1_n12), .CI(npu_inst_pe_1_0_1_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_0_1_sub_67_carry_2_), .S(npu_inst_pe_1_0_1_N66) );
  FA_X1 npu_inst_pe_1_0_1_add_69_U1_1 ( .A(npu_inst_pe_1_0_1_int_q_acc_1_), 
        .B(npu_inst_pe_1_0_1_int_data_1_), .CI(
        npu_inst_pe_1_0_1_add_69_carry_1_), .CO(
        npu_inst_pe_1_0_1_add_69_carry_2_), .S(npu_inst_pe_1_0_1_N74) );
  NAND3_X1 npu_inst_pe_1_0_1_U109 ( .A1(npu_inst_pe_1_0_1_n4), .A2(
        npu_inst_pe_1_0_1_n5), .A3(npu_inst_pe_1_0_1_n6), .ZN(
        npu_inst_pe_1_0_1_n44) );
  NAND3_X1 npu_inst_pe_1_0_1_U108 ( .A1(npu_inst_n72), .A2(
        npu_inst_pe_1_0_1_n5), .A3(npu_inst_pe_1_0_1_n6), .ZN(
        npu_inst_pe_1_0_1_n40) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_0_1_n32), .CK(
        npu_inst_pe_1_0_1_net4539), .RN(npu_inst_pe_1_0_1_n7), .Q(
        npu_inst_pe_1_0_1_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_0_1_n33), .CK(
        npu_inst_pe_1_0_1_net4539), .RN(npu_inst_pe_1_0_1_n7), .Q(
        npu_inst_pe_1_0_1_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_0_1_n34), .CK(
        npu_inst_pe_1_0_1_net4539), .RN(npu_inst_pe_1_0_1_n7), .Q(
        npu_inst_pe_1_0_1_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_0_1_n35), .CK(
        npu_inst_pe_1_0_1_net4539), .RN(npu_inst_pe_1_0_1_n7), .Q(
        npu_inst_pe_1_0_1_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_0_1_n36), .CK(
        npu_inst_pe_1_0_1_net4539), .RN(npu_inst_pe_1_0_1_n7), .Q(
        npu_inst_pe_1_0_1_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_0_1_n98), .CK(
        npu_inst_pe_1_0_1_net4539), .RN(npu_inst_pe_1_0_1_n7), .Q(
        npu_inst_pe_1_0_1_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_0_1_n31), .CK(
        npu_inst_pe_1_0_1_net4539), .RN(npu_inst_pe_1_0_1_n7), .Q(
        npu_inst_pe_1_0_1_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_0_1_n99), .CK(
        npu_inst_pe_1_0_1_net4539), .RN(npu_inst_pe_1_0_1_n7), .Q(
        npu_inst_pe_1_0_1_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_weight_reg_0_ ( .D(npu_inst_n113), .CK(
        npu_inst_pe_1_0_1_net4545), .RN(npu_inst_pe_1_0_1_n7), .Q(
        npu_inst_pe_1_0_1_int_q_weight_0_), .QN(npu_inst_pe_1_0_1_n27) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_weight_reg_1_ ( .D(npu_inst_n119), .CK(
        npu_inst_pe_1_0_1_net4545), .RN(npu_inst_pe_1_0_1_n7), .Q(
        npu_inst_pe_1_0_1_int_q_weight_1_), .QN(npu_inst_pe_1_0_1_n26) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_0_1_n111), 
        .CK(npu_inst_pe_1_0_1_net4545), .RN(npu_inst_pe_1_0_1_n7), .Q(
        npu_inst_pe_1_0_1_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_0_1_n105), 
        .CK(npu_inst_pe_1_0_1_net4545), .RN(npu_inst_pe_1_0_1_n7), .Q(
        npu_inst_pe_1_0_1_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_0_1_n110), 
        .CK(npu_inst_pe_1_0_1_net4545), .RN(npu_inst_pe_1_0_1_n8), .Q(
        npu_inst_pe_1_0_1_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_0_1_n104), 
        .CK(npu_inst_pe_1_0_1_net4545), .RN(npu_inst_pe_1_0_1_n8), .Q(
        npu_inst_pe_1_0_1_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_0_1_n109), 
        .CK(npu_inst_pe_1_0_1_net4545), .RN(npu_inst_pe_1_0_1_n8), .Q(
        npu_inst_pe_1_0_1_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_0_1_n103), 
        .CK(npu_inst_pe_1_0_1_net4545), .RN(npu_inst_pe_1_0_1_n8), .Q(
        npu_inst_pe_1_0_1_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_0_1_n108), 
        .CK(npu_inst_pe_1_0_1_net4545), .RN(npu_inst_pe_1_0_1_n8), .Q(
        npu_inst_pe_1_0_1_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_0_1_n102), 
        .CK(npu_inst_pe_1_0_1_net4545), .RN(npu_inst_pe_1_0_1_n8), .Q(
        npu_inst_pe_1_0_1_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_0_1_n107), 
        .CK(npu_inst_pe_1_0_1_net4545), .RN(npu_inst_pe_1_0_1_n8), .Q(
        npu_inst_pe_1_0_1_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_0_1_n101), 
        .CK(npu_inst_pe_1_0_1_net4545), .RN(npu_inst_pe_1_0_1_n8), .Q(
        npu_inst_pe_1_0_1_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_0_1_n106), 
        .CK(npu_inst_pe_1_0_1_net4545), .RN(npu_inst_pe_1_0_1_n8), .Q(
        npu_inst_pe_1_0_1_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_0_1_n100), 
        .CK(npu_inst_pe_1_0_1_net4545), .RN(npu_inst_pe_1_0_1_n8), .Q(
        npu_inst_pe_1_0_1_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_0_1_n86), 
        .CK(npu_inst_pe_1_0_1_net4545), .RN(npu_inst_pe_1_0_1_n8), .Q(
        npu_inst_pe_1_0_1_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_0_1_n87), 
        .CK(npu_inst_pe_1_0_1_net4545), .RN(npu_inst_pe_1_0_1_n8), .Q(
        npu_inst_pe_1_0_1_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_0_1_n88), 
        .CK(npu_inst_pe_1_0_1_net4545), .RN(npu_inst_pe_1_0_1_n9), .Q(
        npu_inst_pe_1_0_1_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_0_1_n89), 
        .CK(npu_inst_pe_1_0_1_net4545), .RN(npu_inst_pe_1_0_1_n9), .Q(
        npu_inst_pe_1_0_1_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_0_1_n90), 
        .CK(npu_inst_pe_1_0_1_net4545), .RN(npu_inst_pe_1_0_1_n9), .Q(
        npu_inst_pe_1_0_1_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_0_1_n91), 
        .CK(npu_inst_pe_1_0_1_net4545), .RN(npu_inst_pe_1_0_1_n9), .Q(
        npu_inst_pe_1_0_1_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_0_1_n92), 
        .CK(npu_inst_pe_1_0_1_net4545), .RN(npu_inst_pe_1_0_1_n9), .Q(
        npu_inst_pe_1_0_1_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_0_1_n93), 
        .CK(npu_inst_pe_1_0_1_net4545), .RN(npu_inst_pe_1_0_1_n9), .Q(
        npu_inst_pe_1_0_1_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_0_1_n94), 
        .CK(npu_inst_pe_1_0_1_net4545), .RN(npu_inst_pe_1_0_1_n9), .Q(
        npu_inst_pe_1_0_1_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_0_1_n95), 
        .CK(npu_inst_pe_1_0_1_net4545), .RN(npu_inst_pe_1_0_1_n9), .Q(
        npu_inst_pe_1_0_1_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_0_1_n96), 
        .CK(npu_inst_pe_1_0_1_net4545), .RN(npu_inst_pe_1_0_1_n9), .Q(
        npu_inst_pe_1_0_1_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_0_1_n97), 
        .CK(npu_inst_pe_1_0_1_net4545), .RN(npu_inst_pe_1_0_1_n9), .Q(
        npu_inst_pe_1_0_1_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_0_1_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_0_1_N84), .SE(1'b0), .GCK(npu_inst_pe_1_0_1_net4539) );
  CLKGATETST_X1 npu_inst_pe_1_0_1_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n66), .SE(1'b0), .GCK(npu_inst_pe_1_0_1_net4545) );
  MUX2_X1 npu_inst_pe_1_0_2_U161 ( .A(npu_inst_pe_1_0_2_n31), .B(
        npu_inst_pe_1_0_2_n28), .S(npu_inst_pe_1_0_2_n7), .Z(
        npu_inst_pe_1_0_2_N93) );
  MUX2_X1 npu_inst_pe_1_0_2_U160 ( .A(npu_inst_pe_1_0_2_n30), .B(
        npu_inst_pe_1_0_2_n29), .S(npu_inst_n80), .Z(npu_inst_pe_1_0_2_n31) );
  MUX2_X1 npu_inst_pe_1_0_2_U159 ( .A(npu_inst_pe_1_0_2_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_0_2_int_q_reg_v_1__0_), .S(npu_inst_pe_1_0_2_n4), .Z(
        npu_inst_pe_1_0_2_n30) );
  MUX2_X1 npu_inst_pe_1_0_2_U158 ( .A(npu_inst_pe_1_0_2_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_0_2_int_q_reg_v_3__0_), .S(npu_inst_pe_1_0_2_n4), .Z(
        npu_inst_pe_1_0_2_n29) );
  MUX2_X1 npu_inst_pe_1_0_2_U157 ( .A(npu_inst_pe_1_0_2_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_0_2_int_q_reg_v_5__0_), .S(npu_inst_pe_1_0_2_n4), .Z(
        npu_inst_pe_1_0_2_n28) );
  MUX2_X1 npu_inst_pe_1_0_2_U156 ( .A(npu_inst_pe_1_0_2_n25), .B(
        npu_inst_pe_1_0_2_n22), .S(npu_inst_pe_1_0_2_n7), .Z(
        npu_inst_pe_1_0_2_N94) );
  MUX2_X1 npu_inst_pe_1_0_2_U155 ( .A(npu_inst_pe_1_0_2_n24), .B(
        npu_inst_pe_1_0_2_n23), .S(npu_inst_n80), .Z(npu_inst_pe_1_0_2_n25) );
  MUX2_X1 npu_inst_pe_1_0_2_U154 ( .A(npu_inst_pe_1_0_2_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_0_2_int_q_reg_v_1__1_), .S(npu_inst_pe_1_0_2_n4), .Z(
        npu_inst_pe_1_0_2_n24) );
  MUX2_X1 npu_inst_pe_1_0_2_U153 ( .A(npu_inst_pe_1_0_2_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_0_2_int_q_reg_v_3__1_), .S(npu_inst_pe_1_0_2_n4), .Z(
        npu_inst_pe_1_0_2_n23) );
  MUX2_X1 npu_inst_pe_1_0_2_U152 ( .A(npu_inst_pe_1_0_2_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_0_2_int_q_reg_v_5__1_), .S(npu_inst_pe_1_0_2_n4), .Z(
        npu_inst_pe_1_0_2_n22) );
  MUX2_X1 npu_inst_pe_1_0_2_U151 ( .A(npu_inst_pe_1_0_2_n21), .B(
        npu_inst_pe_1_0_2_n18), .S(npu_inst_pe_1_0_2_n7), .Z(
        npu_inst_int_data_x_0__2__1_) );
  MUX2_X1 npu_inst_pe_1_0_2_U150 ( .A(npu_inst_pe_1_0_2_n20), .B(
        npu_inst_pe_1_0_2_n19), .S(npu_inst_n80), .Z(npu_inst_pe_1_0_2_n21) );
  MUX2_X1 npu_inst_pe_1_0_2_U149 ( .A(npu_inst_pe_1_0_2_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_0_2_int_q_reg_h_1__1_), .S(npu_inst_pe_1_0_2_n4), .Z(
        npu_inst_pe_1_0_2_n20) );
  MUX2_X1 npu_inst_pe_1_0_2_U148 ( .A(npu_inst_pe_1_0_2_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_0_2_int_q_reg_h_3__1_), .S(npu_inst_pe_1_0_2_n4), .Z(
        npu_inst_pe_1_0_2_n19) );
  MUX2_X1 npu_inst_pe_1_0_2_U147 ( .A(npu_inst_pe_1_0_2_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_0_2_int_q_reg_h_5__1_), .S(npu_inst_pe_1_0_2_n4), .Z(
        npu_inst_pe_1_0_2_n18) );
  MUX2_X1 npu_inst_pe_1_0_2_U146 ( .A(npu_inst_pe_1_0_2_n17), .B(
        npu_inst_pe_1_0_2_n14), .S(npu_inst_pe_1_0_2_n7), .Z(
        npu_inst_int_data_x_0__2__0_) );
  MUX2_X1 npu_inst_pe_1_0_2_U145 ( .A(npu_inst_pe_1_0_2_n16), .B(
        npu_inst_pe_1_0_2_n15), .S(npu_inst_n80), .Z(npu_inst_pe_1_0_2_n17) );
  MUX2_X1 npu_inst_pe_1_0_2_U144 ( .A(npu_inst_pe_1_0_2_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_0_2_int_q_reg_h_1__0_), .S(npu_inst_pe_1_0_2_n4), .Z(
        npu_inst_pe_1_0_2_n16) );
  MUX2_X1 npu_inst_pe_1_0_2_U143 ( .A(npu_inst_pe_1_0_2_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_0_2_int_q_reg_h_3__0_), .S(npu_inst_pe_1_0_2_n4), .Z(
        npu_inst_pe_1_0_2_n15) );
  MUX2_X1 npu_inst_pe_1_0_2_U142 ( .A(npu_inst_pe_1_0_2_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_0_2_int_q_reg_h_5__0_), .S(npu_inst_pe_1_0_2_n4), .Z(
        npu_inst_pe_1_0_2_n14) );
  XOR2_X1 npu_inst_pe_1_0_2_U141 ( .A(npu_inst_pe_1_0_2_int_data_0_), .B(
        npu_inst_pe_1_0_2_int_q_acc_0_), .Z(npu_inst_pe_1_0_2_N73) );
  AND2_X1 npu_inst_pe_1_0_2_U140 ( .A1(npu_inst_pe_1_0_2_int_q_acc_0_), .A2(
        npu_inst_pe_1_0_2_int_data_0_), .ZN(npu_inst_pe_1_0_2_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_0_2_U139 ( .A(npu_inst_pe_1_0_2_int_q_acc_0_), .B(
        npu_inst_pe_1_0_2_n12), .ZN(npu_inst_pe_1_0_2_N65) );
  OR2_X1 npu_inst_pe_1_0_2_U138 ( .A1(npu_inst_pe_1_0_2_n12), .A2(
        npu_inst_pe_1_0_2_int_q_acc_0_), .ZN(npu_inst_pe_1_0_2_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_0_2_U137 ( .A(npu_inst_pe_1_0_2_int_q_acc_2_), .B(
        npu_inst_pe_1_0_2_add_69_carry_2_), .Z(npu_inst_pe_1_0_2_N75) );
  AND2_X1 npu_inst_pe_1_0_2_U136 ( .A1(npu_inst_pe_1_0_2_add_69_carry_2_), 
        .A2(npu_inst_pe_1_0_2_int_q_acc_2_), .ZN(
        npu_inst_pe_1_0_2_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_0_2_U135 ( .A(npu_inst_pe_1_0_2_int_q_acc_3_), .B(
        npu_inst_pe_1_0_2_add_69_carry_3_), .Z(npu_inst_pe_1_0_2_N76) );
  AND2_X1 npu_inst_pe_1_0_2_U134 ( .A1(npu_inst_pe_1_0_2_add_69_carry_3_), 
        .A2(npu_inst_pe_1_0_2_int_q_acc_3_), .ZN(
        npu_inst_pe_1_0_2_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_0_2_U133 ( .A(npu_inst_pe_1_0_2_int_q_acc_4_), .B(
        npu_inst_pe_1_0_2_add_69_carry_4_), .Z(npu_inst_pe_1_0_2_N77) );
  AND2_X1 npu_inst_pe_1_0_2_U132 ( .A1(npu_inst_pe_1_0_2_add_69_carry_4_), 
        .A2(npu_inst_pe_1_0_2_int_q_acc_4_), .ZN(
        npu_inst_pe_1_0_2_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_0_2_U131 ( .A(npu_inst_pe_1_0_2_int_q_acc_5_), .B(
        npu_inst_pe_1_0_2_add_69_carry_5_), .Z(npu_inst_pe_1_0_2_N78) );
  AND2_X1 npu_inst_pe_1_0_2_U130 ( .A1(npu_inst_pe_1_0_2_add_69_carry_5_), 
        .A2(npu_inst_pe_1_0_2_int_q_acc_5_), .ZN(
        npu_inst_pe_1_0_2_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_0_2_U129 ( .A(npu_inst_pe_1_0_2_int_q_acc_6_), .B(
        npu_inst_pe_1_0_2_add_69_carry_6_), .Z(npu_inst_pe_1_0_2_N79) );
  AND2_X1 npu_inst_pe_1_0_2_U128 ( .A1(npu_inst_pe_1_0_2_add_69_carry_6_), 
        .A2(npu_inst_pe_1_0_2_int_q_acc_6_), .ZN(
        npu_inst_pe_1_0_2_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_0_2_U127 ( .A(npu_inst_pe_1_0_2_int_q_acc_7_), .B(
        npu_inst_pe_1_0_2_add_69_carry_7_), .Z(npu_inst_pe_1_0_2_N80) );
  XNOR2_X1 npu_inst_pe_1_0_2_U126 ( .A(npu_inst_pe_1_0_2_sub_67_carry_2_), .B(
        npu_inst_pe_1_0_2_int_q_acc_2_), .ZN(npu_inst_pe_1_0_2_N67) );
  OR2_X1 npu_inst_pe_1_0_2_U125 ( .A1(npu_inst_pe_1_0_2_int_q_acc_2_), .A2(
        npu_inst_pe_1_0_2_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_0_2_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_0_2_U124 ( .A(npu_inst_pe_1_0_2_sub_67_carry_3_), .B(
        npu_inst_pe_1_0_2_int_q_acc_3_), .ZN(npu_inst_pe_1_0_2_N68) );
  OR2_X1 npu_inst_pe_1_0_2_U123 ( .A1(npu_inst_pe_1_0_2_int_q_acc_3_), .A2(
        npu_inst_pe_1_0_2_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_0_2_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_0_2_U122 ( .A(npu_inst_pe_1_0_2_sub_67_carry_4_), .B(
        npu_inst_pe_1_0_2_int_q_acc_4_), .ZN(npu_inst_pe_1_0_2_N69) );
  OR2_X1 npu_inst_pe_1_0_2_U121 ( .A1(npu_inst_pe_1_0_2_int_q_acc_4_), .A2(
        npu_inst_pe_1_0_2_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_0_2_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_0_2_U120 ( .A(npu_inst_pe_1_0_2_sub_67_carry_5_), .B(
        npu_inst_pe_1_0_2_int_q_acc_5_), .ZN(npu_inst_pe_1_0_2_N70) );
  OR2_X1 npu_inst_pe_1_0_2_U119 ( .A1(npu_inst_pe_1_0_2_int_q_acc_5_), .A2(
        npu_inst_pe_1_0_2_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_0_2_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_0_2_U118 ( .A(npu_inst_pe_1_0_2_sub_67_carry_6_), .B(
        npu_inst_pe_1_0_2_int_q_acc_6_), .ZN(npu_inst_pe_1_0_2_N71) );
  OR2_X1 npu_inst_pe_1_0_2_U117 ( .A1(npu_inst_pe_1_0_2_int_q_acc_6_), .A2(
        npu_inst_pe_1_0_2_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_0_2_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_0_2_U116 ( .A(npu_inst_pe_1_0_2_int_q_acc_7_), .B(
        npu_inst_pe_1_0_2_sub_67_carry_7_), .ZN(npu_inst_pe_1_0_2_N72) );
  INV_X1 npu_inst_pe_1_0_2_U115 ( .A(npu_inst_n80), .ZN(npu_inst_pe_1_0_2_n6)
         );
  INV_X1 npu_inst_pe_1_0_2_U114 ( .A(npu_inst_n60), .ZN(npu_inst_pe_1_0_2_n3)
         );
  AOI22_X1 npu_inst_pe_1_0_2_U113 ( .A1(npu_inst_int_data_y_1__2__0_), .A2(
        npu_inst_pe_1_0_2_n58), .B1(npu_inst_pe_1_0_2_n118), .B2(
        npu_inst_pe_1_0_2_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_0_2_n57) );
  INV_X1 npu_inst_pe_1_0_2_U112 ( .A(npu_inst_pe_1_0_2_n57), .ZN(
        npu_inst_pe_1_0_2_n107) );
  AOI22_X1 npu_inst_pe_1_0_2_U111 ( .A1(npu_inst_int_data_y_1__2__0_), .A2(
        npu_inst_pe_1_0_2_n54), .B1(npu_inst_pe_1_0_2_n117), .B2(
        npu_inst_pe_1_0_2_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_0_2_n53) );
  INV_X1 npu_inst_pe_1_0_2_U110 ( .A(npu_inst_pe_1_0_2_n53), .ZN(
        npu_inst_pe_1_0_2_n108) );
  AOI22_X1 npu_inst_pe_1_0_2_U107 ( .A1(npu_inst_int_data_y_1__2__0_), .A2(
        npu_inst_pe_1_0_2_n50), .B1(npu_inst_pe_1_0_2_n116), .B2(
        npu_inst_pe_1_0_2_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_0_2_n49) );
  INV_X1 npu_inst_pe_1_0_2_U106 ( .A(npu_inst_pe_1_0_2_n49), .ZN(
        npu_inst_pe_1_0_2_n109) );
  AOI22_X1 npu_inst_pe_1_0_2_U105 ( .A1(npu_inst_int_data_y_1__2__0_), .A2(
        npu_inst_pe_1_0_2_n46), .B1(npu_inst_pe_1_0_2_n115), .B2(
        npu_inst_pe_1_0_2_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_0_2_n45) );
  INV_X1 npu_inst_pe_1_0_2_U104 ( .A(npu_inst_pe_1_0_2_n45), .ZN(
        npu_inst_pe_1_0_2_n110) );
  AOI22_X1 npu_inst_pe_1_0_2_U103 ( .A1(npu_inst_int_data_y_1__2__0_), .A2(
        npu_inst_pe_1_0_2_n42), .B1(npu_inst_pe_1_0_2_n114), .B2(
        npu_inst_pe_1_0_2_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_0_2_n41) );
  INV_X1 npu_inst_pe_1_0_2_U102 ( .A(npu_inst_pe_1_0_2_n41), .ZN(
        npu_inst_pe_1_0_2_n111) );
  AOI22_X1 npu_inst_pe_1_0_2_U101 ( .A1(npu_inst_int_data_y_1__2__1_), .A2(
        npu_inst_pe_1_0_2_n58), .B1(npu_inst_pe_1_0_2_n118), .B2(
        npu_inst_pe_1_0_2_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_0_2_n59) );
  INV_X1 npu_inst_pe_1_0_2_U100 ( .A(npu_inst_pe_1_0_2_n59), .ZN(
        npu_inst_pe_1_0_2_n101) );
  AOI22_X1 npu_inst_pe_1_0_2_U99 ( .A1(npu_inst_int_data_y_1__2__1_), .A2(
        npu_inst_pe_1_0_2_n54), .B1(npu_inst_pe_1_0_2_n117), .B2(
        npu_inst_pe_1_0_2_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_0_2_n55) );
  INV_X1 npu_inst_pe_1_0_2_U98 ( .A(npu_inst_pe_1_0_2_n55), .ZN(
        npu_inst_pe_1_0_2_n102) );
  AOI22_X1 npu_inst_pe_1_0_2_U97 ( .A1(npu_inst_int_data_y_1__2__1_), .A2(
        npu_inst_pe_1_0_2_n50), .B1(npu_inst_pe_1_0_2_n116), .B2(
        npu_inst_pe_1_0_2_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_0_2_n51) );
  INV_X1 npu_inst_pe_1_0_2_U96 ( .A(npu_inst_pe_1_0_2_n51), .ZN(
        npu_inst_pe_1_0_2_n103) );
  AOI22_X1 npu_inst_pe_1_0_2_U95 ( .A1(npu_inst_int_data_y_1__2__1_), .A2(
        npu_inst_pe_1_0_2_n46), .B1(npu_inst_pe_1_0_2_n115), .B2(
        npu_inst_pe_1_0_2_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_0_2_n47) );
  INV_X1 npu_inst_pe_1_0_2_U94 ( .A(npu_inst_pe_1_0_2_n47), .ZN(
        npu_inst_pe_1_0_2_n104) );
  AOI22_X1 npu_inst_pe_1_0_2_U93 ( .A1(npu_inst_int_data_y_1__2__1_), .A2(
        npu_inst_pe_1_0_2_n42), .B1(npu_inst_pe_1_0_2_n114), .B2(
        npu_inst_pe_1_0_2_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_0_2_n43) );
  INV_X1 npu_inst_pe_1_0_2_U92 ( .A(npu_inst_pe_1_0_2_n43), .ZN(
        npu_inst_pe_1_0_2_n105) );
  AOI22_X1 npu_inst_pe_1_0_2_U91 ( .A1(npu_inst_pe_1_0_2_n38), .A2(
        npu_inst_int_data_y_1__2__1_), .B1(npu_inst_pe_1_0_2_n113), .B2(
        npu_inst_pe_1_0_2_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_0_2_n39) );
  INV_X1 npu_inst_pe_1_0_2_U90 ( .A(npu_inst_pe_1_0_2_n39), .ZN(
        npu_inst_pe_1_0_2_n106) );
  AOI22_X1 npu_inst_pe_1_0_2_U89 ( .A1(npu_inst_pe_1_0_2_n38), .A2(
        npu_inst_int_data_y_1__2__0_), .B1(npu_inst_pe_1_0_2_n113), .B2(
        npu_inst_pe_1_0_2_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_0_2_n37) );
  INV_X1 npu_inst_pe_1_0_2_U88 ( .A(npu_inst_pe_1_0_2_n37), .ZN(
        npu_inst_pe_1_0_2_n112) );
  NAND2_X1 npu_inst_pe_1_0_2_U87 ( .A1(npu_inst_pe_1_0_2_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_0_2_n60), .ZN(npu_inst_pe_1_0_2_n74) );
  OAI21_X1 npu_inst_pe_1_0_2_U86 ( .B1(npu_inst_pe_1_0_2_n63), .B2(
        npu_inst_pe_1_0_2_n60), .A(npu_inst_pe_1_0_2_n74), .ZN(
        npu_inst_pe_1_0_2_n97) );
  NAND2_X1 npu_inst_pe_1_0_2_U85 ( .A1(npu_inst_pe_1_0_2_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_0_2_n60), .ZN(npu_inst_pe_1_0_2_n73) );
  OAI21_X1 npu_inst_pe_1_0_2_U84 ( .B1(npu_inst_pe_1_0_2_n61), .B2(
        npu_inst_pe_1_0_2_n60), .A(npu_inst_pe_1_0_2_n73), .ZN(
        npu_inst_pe_1_0_2_n96) );
  NAND2_X1 npu_inst_pe_1_0_2_U83 ( .A1(npu_inst_pe_1_0_2_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_0_2_n56), .ZN(npu_inst_pe_1_0_2_n72) );
  OAI21_X1 npu_inst_pe_1_0_2_U82 ( .B1(npu_inst_pe_1_0_2_n63), .B2(
        npu_inst_pe_1_0_2_n56), .A(npu_inst_pe_1_0_2_n72), .ZN(
        npu_inst_pe_1_0_2_n95) );
  NAND2_X1 npu_inst_pe_1_0_2_U81 ( .A1(npu_inst_pe_1_0_2_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_0_2_n56), .ZN(npu_inst_pe_1_0_2_n71) );
  OAI21_X1 npu_inst_pe_1_0_2_U80 ( .B1(npu_inst_pe_1_0_2_n61), .B2(
        npu_inst_pe_1_0_2_n56), .A(npu_inst_pe_1_0_2_n71), .ZN(
        npu_inst_pe_1_0_2_n94) );
  NAND2_X1 npu_inst_pe_1_0_2_U79 ( .A1(npu_inst_pe_1_0_2_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_0_2_n52), .ZN(npu_inst_pe_1_0_2_n70) );
  OAI21_X1 npu_inst_pe_1_0_2_U78 ( .B1(npu_inst_pe_1_0_2_n63), .B2(
        npu_inst_pe_1_0_2_n52), .A(npu_inst_pe_1_0_2_n70), .ZN(
        npu_inst_pe_1_0_2_n93) );
  NAND2_X1 npu_inst_pe_1_0_2_U77 ( .A1(npu_inst_pe_1_0_2_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_0_2_n52), .ZN(npu_inst_pe_1_0_2_n69) );
  OAI21_X1 npu_inst_pe_1_0_2_U76 ( .B1(npu_inst_pe_1_0_2_n61), .B2(
        npu_inst_pe_1_0_2_n52), .A(npu_inst_pe_1_0_2_n69), .ZN(
        npu_inst_pe_1_0_2_n92) );
  NAND2_X1 npu_inst_pe_1_0_2_U75 ( .A1(npu_inst_pe_1_0_2_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_0_2_n48), .ZN(npu_inst_pe_1_0_2_n68) );
  OAI21_X1 npu_inst_pe_1_0_2_U74 ( .B1(npu_inst_pe_1_0_2_n63), .B2(
        npu_inst_pe_1_0_2_n48), .A(npu_inst_pe_1_0_2_n68), .ZN(
        npu_inst_pe_1_0_2_n91) );
  NAND2_X1 npu_inst_pe_1_0_2_U73 ( .A1(npu_inst_pe_1_0_2_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_0_2_n48), .ZN(npu_inst_pe_1_0_2_n67) );
  OAI21_X1 npu_inst_pe_1_0_2_U72 ( .B1(npu_inst_pe_1_0_2_n61), .B2(
        npu_inst_pe_1_0_2_n48), .A(npu_inst_pe_1_0_2_n67), .ZN(
        npu_inst_pe_1_0_2_n90) );
  NAND2_X1 npu_inst_pe_1_0_2_U71 ( .A1(npu_inst_pe_1_0_2_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_0_2_n44), .ZN(npu_inst_pe_1_0_2_n66) );
  OAI21_X1 npu_inst_pe_1_0_2_U70 ( .B1(npu_inst_pe_1_0_2_n63), .B2(
        npu_inst_pe_1_0_2_n44), .A(npu_inst_pe_1_0_2_n66), .ZN(
        npu_inst_pe_1_0_2_n89) );
  NAND2_X1 npu_inst_pe_1_0_2_U69 ( .A1(npu_inst_pe_1_0_2_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_0_2_n44), .ZN(npu_inst_pe_1_0_2_n65) );
  OAI21_X1 npu_inst_pe_1_0_2_U68 ( .B1(npu_inst_pe_1_0_2_n61), .B2(
        npu_inst_pe_1_0_2_n44), .A(npu_inst_pe_1_0_2_n65), .ZN(
        npu_inst_pe_1_0_2_n88) );
  NAND2_X1 npu_inst_pe_1_0_2_U67 ( .A1(npu_inst_pe_1_0_2_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_0_2_n40), .ZN(npu_inst_pe_1_0_2_n64) );
  OAI21_X1 npu_inst_pe_1_0_2_U66 ( .B1(npu_inst_pe_1_0_2_n63), .B2(
        npu_inst_pe_1_0_2_n40), .A(npu_inst_pe_1_0_2_n64), .ZN(
        npu_inst_pe_1_0_2_n87) );
  NAND2_X1 npu_inst_pe_1_0_2_U65 ( .A1(npu_inst_pe_1_0_2_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_0_2_n40), .ZN(npu_inst_pe_1_0_2_n62) );
  OAI21_X1 npu_inst_pe_1_0_2_U64 ( .B1(npu_inst_pe_1_0_2_n61), .B2(
        npu_inst_pe_1_0_2_n40), .A(npu_inst_pe_1_0_2_n62), .ZN(
        npu_inst_pe_1_0_2_n86) );
  AND2_X1 npu_inst_pe_1_0_2_U63 ( .A1(npu_inst_pe_1_0_2_int_q_acc_2_), .A2(
        npu_inst_pe_1_0_2_n1), .ZN(int_o_data_npu[42]) );
  AND2_X1 npu_inst_pe_1_0_2_U62 ( .A1(npu_inst_pe_1_0_2_int_q_acc_3_), .A2(
        npu_inst_pe_1_0_2_n2), .ZN(int_o_data_npu[43]) );
  NOR3_X1 npu_inst_pe_1_0_2_U61 ( .A1(npu_inst_pe_1_0_2_n26), .A2(npu_inst_n60), .A3(npu_inst_int_ckg[61]), .ZN(npu_inst_pe_1_0_2_n85) );
  OR2_X1 npu_inst_pe_1_0_2_U60 ( .A1(npu_inst_pe_1_0_2_n85), .A2(
        npu_inst_pe_1_0_2_n2), .ZN(npu_inst_pe_1_0_2_N84) );
  AND2_X1 npu_inst_pe_1_0_2_U59 ( .A1(npu_inst_pe_1_0_2_int_q_acc_6_), .A2(
        npu_inst_pe_1_0_2_n2), .ZN(int_o_data_npu[46]) );
  AND2_X1 npu_inst_pe_1_0_2_U58 ( .A1(npu_inst_pe_1_0_2_int_q_acc_5_), .A2(
        npu_inst_pe_1_0_2_n2), .ZN(int_o_data_npu[45]) );
  AND2_X1 npu_inst_pe_1_0_2_U57 ( .A1(npu_inst_pe_1_0_2_int_q_acc_4_), .A2(
        npu_inst_pe_1_0_2_n2), .ZN(int_o_data_npu[44]) );
  AOI222_X1 npu_inst_pe_1_0_2_U56 ( .A1(npu_inst_int_data_res_1__2__0_), .A2(
        npu_inst_pe_1_0_2_n1), .B1(npu_inst_pe_1_0_2_N73), .B2(
        npu_inst_pe_1_0_2_n76), .C1(npu_inst_pe_1_0_2_N65), .C2(
        npu_inst_pe_1_0_2_n77), .ZN(npu_inst_pe_1_0_2_n84) );
  INV_X1 npu_inst_pe_1_0_2_U55 ( .A(npu_inst_pe_1_0_2_n84), .ZN(
        npu_inst_pe_1_0_2_n100) );
  AOI222_X1 npu_inst_pe_1_0_2_U54 ( .A1(npu_inst_int_data_res_1__2__7_), .A2(
        npu_inst_pe_1_0_2_n1), .B1(npu_inst_pe_1_0_2_N80), .B2(
        npu_inst_pe_1_0_2_n76), .C1(npu_inst_pe_1_0_2_N72), .C2(
        npu_inst_pe_1_0_2_n77), .ZN(npu_inst_pe_1_0_2_n75) );
  INV_X1 npu_inst_pe_1_0_2_U53 ( .A(npu_inst_pe_1_0_2_n75), .ZN(
        npu_inst_pe_1_0_2_n32) );
  AOI222_X1 npu_inst_pe_1_0_2_U52 ( .A1(npu_inst_int_data_res_1__2__1_), .A2(
        npu_inst_pe_1_0_2_n1), .B1(npu_inst_pe_1_0_2_N74), .B2(
        npu_inst_pe_1_0_2_n76), .C1(npu_inst_pe_1_0_2_N66), .C2(
        npu_inst_pe_1_0_2_n77), .ZN(npu_inst_pe_1_0_2_n83) );
  INV_X1 npu_inst_pe_1_0_2_U51 ( .A(npu_inst_pe_1_0_2_n83), .ZN(
        npu_inst_pe_1_0_2_n99) );
  AOI222_X1 npu_inst_pe_1_0_2_U50 ( .A1(npu_inst_int_data_res_1__2__2_), .A2(
        npu_inst_pe_1_0_2_n1), .B1(npu_inst_pe_1_0_2_N75), .B2(
        npu_inst_pe_1_0_2_n76), .C1(npu_inst_pe_1_0_2_N67), .C2(
        npu_inst_pe_1_0_2_n77), .ZN(npu_inst_pe_1_0_2_n82) );
  INV_X1 npu_inst_pe_1_0_2_U49 ( .A(npu_inst_pe_1_0_2_n82), .ZN(
        npu_inst_pe_1_0_2_n98) );
  AOI222_X1 npu_inst_pe_1_0_2_U48 ( .A1(npu_inst_int_data_res_1__2__3_), .A2(
        npu_inst_pe_1_0_2_n1), .B1(npu_inst_pe_1_0_2_N76), .B2(
        npu_inst_pe_1_0_2_n76), .C1(npu_inst_pe_1_0_2_N68), .C2(
        npu_inst_pe_1_0_2_n77), .ZN(npu_inst_pe_1_0_2_n81) );
  INV_X1 npu_inst_pe_1_0_2_U47 ( .A(npu_inst_pe_1_0_2_n81), .ZN(
        npu_inst_pe_1_0_2_n36) );
  AOI222_X1 npu_inst_pe_1_0_2_U46 ( .A1(npu_inst_int_data_res_1__2__4_), .A2(
        npu_inst_pe_1_0_2_n1), .B1(npu_inst_pe_1_0_2_N77), .B2(
        npu_inst_pe_1_0_2_n76), .C1(npu_inst_pe_1_0_2_N69), .C2(
        npu_inst_pe_1_0_2_n77), .ZN(npu_inst_pe_1_0_2_n80) );
  INV_X1 npu_inst_pe_1_0_2_U45 ( .A(npu_inst_pe_1_0_2_n80), .ZN(
        npu_inst_pe_1_0_2_n35) );
  AOI222_X1 npu_inst_pe_1_0_2_U44 ( .A1(npu_inst_int_data_res_1__2__5_), .A2(
        npu_inst_pe_1_0_2_n1), .B1(npu_inst_pe_1_0_2_N78), .B2(
        npu_inst_pe_1_0_2_n76), .C1(npu_inst_pe_1_0_2_N70), .C2(
        npu_inst_pe_1_0_2_n77), .ZN(npu_inst_pe_1_0_2_n79) );
  INV_X1 npu_inst_pe_1_0_2_U43 ( .A(npu_inst_pe_1_0_2_n79), .ZN(
        npu_inst_pe_1_0_2_n34) );
  AOI222_X1 npu_inst_pe_1_0_2_U42 ( .A1(npu_inst_int_data_res_1__2__6_), .A2(
        npu_inst_pe_1_0_2_n1), .B1(npu_inst_pe_1_0_2_N79), .B2(
        npu_inst_pe_1_0_2_n76), .C1(npu_inst_pe_1_0_2_N71), .C2(
        npu_inst_pe_1_0_2_n77), .ZN(npu_inst_pe_1_0_2_n78) );
  INV_X1 npu_inst_pe_1_0_2_U41 ( .A(npu_inst_pe_1_0_2_n78), .ZN(
        npu_inst_pe_1_0_2_n33) );
  INV_X1 npu_inst_pe_1_0_2_U40 ( .A(npu_inst_pe_1_0_2_int_data_1_), .ZN(
        npu_inst_pe_1_0_2_n13) );
  AND2_X1 npu_inst_pe_1_0_2_U39 ( .A1(npu_inst_int_data_x_0__2__1_), .A2(
        npu_inst_pe_1_0_2_int_q_weight_1_), .ZN(npu_inst_pe_1_0_2_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_0_2_U38 ( .A1(npu_inst_int_data_x_0__2__0_), .A2(
        npu_inst_pe_1_0_2_int_q_weight_1_), .ZN(npu_inst_pe_1_0_2_int_data_0_)
         );
  AND2_X1 npu_inst_pe_1_0_2_U37 ( .A1(npu_inst_pe_1_0_2_n2), .A2(
        npu_inst_pe_1_0_2_int_q_acc_7_), .ZN(int_o_data_npu[47]) );
  AND2_X1 npu_inst_pe_1_0_2_U36 ( .A1(npu_inst_pe_1_0_2_int_q_acc_1_), .A2(
        npu_inst_pe_1_0_2_n1), .ZN(int_o_data_npu[41]) );
  AND2_X1 npu_inst_pe_1_0_2_U35 ( .A1(npu_inst_pe_1_0_2_int_q_acc_0_), .A2(
        npu_inst_pe_1_0_2_n1), .ZN(int_o_data_npu[40]) );
  AND2_X1 npu_inst_pe_1_0_2_U34 ( .A1(npu_inst_pe_1_0_2_N93), .A2(npu_inst_n60), .ZN(npu_inst_pe_1_0_2_o_data_v_0_) );
  AND2_X1 npu_inst_pe_1_0_2_U33 ( .A1(npu_inst_n60), .A2(npu_inst_pe_1_0_2_N94), .ZN(npu_inst_pe_1_0_2_o_data_v_1_) );
  AOI22_X1 npu_inst_pe_1_0_2_U32 ( .A1(npu_inst_n60), .A2(
        npu_inst_int_data_y_1__2__1_), .B1(npu_inst_pe_1_0_2_n3), .B2(
        npu_inst_int_data_x_0__3__1_), .ZN(npu_inst_pe_1_0_2_n63) );
  AOI22_X1 npu_inst_pe_1_0_2_U31 ( .A1(npu_inst_n60), .A2(
        npu_inst_int_data_y_1__2__0_), .B1(npu_inst_pe_1_0_2_n3), .B2(
        npu_inst_int_data_x_0__3__0_), .ZN(npu_inst_pe_1_0_2_n61) );
  INV_X1 npu_inst_pe_1_0_2_U30 ( .A(npu_inst_pe_1_0_2_int_data_0_), .ZN(
        npu_inst_pe_1_0_2_n12) );
  INV_X1 npu_inst_pe_1_0_2_U29 ( .A(npu_inst_n72), .ZN(npu_inst_pe_1_0_2_n5)
         );
  OR3_X1 npu_inst_pe_1_0_2_U28 ( .A1(npu_inst_n80), .A2(npu_inst_pe_1_0_2_n7), 
        .A3(npu_inst_pe_1_0_2_n5), .ZN(npu_inst_pe_1_0_2_n56) );
  OR3_X1 npu_inst_pe_1_0_2_U27 ( .A1(npu_inst_pe_1_0_2_n5), .A2(
        npu_inst_pe_1_0_2_n7), .A3(npu_inst_pe_1_0_2_n6), .ZN(
        npu_inst_pe_1_0_2_n48) );
  INV_X1 npu_inst_pe_1_0_2_U26 ( .A(npu_inst_pe_1_0_2_n5), .ZN(
        npu_inst_pe_1_0_2_n4) );
  OR3_X1 npu_inst_pe_1_0_2_U25 ( .A1(npu_inst_pe_1_0_2_n4), .A2(
        npu_inst_pe_1_0_2_n7), .A3(npu_inst_pe_1_0_2_n6), .ZN(
        npu_inst_pe_1_0_2_n52) );
  OR3_X1 npu_inst_pe_1_0_2_U24 ( .A1(npu_inst_n80), .A2(npu_inst_pe_1_0_2_n7), 
        .A3(npu_inst_pe_1_0_2_n4), .ZN(npu_inst_pe_1_0_2_n60) );
  NOR2_X1 npu_inst_pe_1_0_2_U23 ( .A1(npu_inst_pe_1_0_2_n60), .A2(
        npu_inst_pe_1_0_2_n3), .ZN(npu_inst_pe_1_0_2_n58) );
  NOR2_X1 npu_inst_pe_1_0_2_U22 ( .A1(npu_inst_pe_1_0_2_n56), .A2(
        npu_inst_pe_1_0_2_n3), .ZN(npu_inst_pe_1_0_2_n54) );
  NOR2_X1 npu_inst_pe_1_0_2_U21 ( .A1(npu_inst_pe_1_0_2_n52), .A2(
        npu_inst_pe_1_0_2_n3), .ZN(npu_inst_pe_1_0_2_n50) );
  NOR2_X1 npu_inst_pe_1_0_2_U20 ( .A1(npu_inst_pe_1_0_2_n48), .A2(
        npu_inst_pe_1_0_2_n3), .ZN(npu_inst_pe_1_0_2_n46) );
  NOR2_X1 npu_inst_pe_1_0_2_U19 ( .A1(npu_inst_pe_1_0_2_n40), .A2(
        npu_inst_pe_1_0_2_n3), .ZN(npu_inst_pe_1_0_2_n38) );
  NOR2_X1 npu_inst_pe_1_0_2_U18 ( .A1(npu_inst_pe_1_0_2_n44), .A2(
        npu_inst_pe_1_0_2_n3), .ZN(npu_inst_pe_1_0_2_n42) );
  BUF_X1 npu_inst_pe_1_0_2_U17 ( .A(npu_inst_n107), .Z(npu_inst_pe_1_0_2_n7)
         );
  INV_X1 npu_inst_pe_1_0_2_U16 ( .A(npu_inst_n127), .ZN(npu_inst_pe_1_0_2_n11)
         );
  INV_X1 npu_inst_pe_1_0_2_U15 ( .A(npu_inst_pe_1_0_2_n38), .ZN(
        npu_inst_pe_1_0_2_n113) );
  INV_X1 npu_inst_pe_1_0_2_U14 ( .A(npu_inst_pe_1_0_2_n58), .ZN(
        npu_inst_pe_1_0_2_n118) );
  INV_X1 npu_inst_pe_1_0_2_U13 ( .A(npu_inst_pe_1_0_2_n54), .ZN(
        npu_inst_pe_1_0_2_n117) );
  INV_X1 npu_inst_pe_1_0_2_U12 ( .A(npu_inst_pe_1_0_2_n50), .ZN(
        npu_inst_pe_1_0_2_n116) );
  INV_X1 npu_inst_pe_1_0_2_U11 ( .A(npu_inst_pe_1_0_2_n46), .ZN(
        npu_inst_pe_1_0_2_n115) );
  INV_X1 npu_inst_pe_1_0_2_U10 ( .A(npu_inst_pe_1_0_2_n42), .ZN(
        npu_inst_pe_1_0_2_n114) );
  BUF_X1 npu_inst_pe_1_0_2_U9 ( .A(npu_inst_n37), .Z(npu_inst_pe_1_0_2_n2) );
  BUF_X1 npu_inst_pe_1_0_2_U8 ( .A(npu_inst_n37), .Z(npu_inst_pe_1_0_2_n1) );
  BUF_X1 npu_inst_pe_1_0_2_U7 ( .A(npu_inst_pe_1_0_2_n11), .Z(
        npu_inst_pe_1_0_2_n10) );
  BUF_X1 npu_inst_pe_1_0_2_U6 ( .A(npu_inst_pe_1_0_2_n11), .Z(
        npu_inst_pe_1_0_2_n9) );
  BUF_X1 npu_inst_pe_1_0_2_U5 ( .A(npu_inst_pe_1_0_2_n11), .Z(
        npu_inst_pe_1_0_2_n8) );
  NOR2_X1 npu_inst_pe_1_0_2_U4 ( .A1(npu_inst_pe_1_0_2_int_q_weight_0_), .A2(
        npu_inst_pe_1_0_2_n1), .ZN(npu_inst_pe_1_0_2_n76) );
  NOR2_X1 npu_inst_pe_1_0_2_U3 ( .A1(npu_inst_pe_1_0_2_n27), .A2(
        npu_inst_pe_1_0_2_n1), .ZN(npu_inst_pe_1_0_2_n77) );
  FA_X1 npu_inst_pe_1_0_2_sub_67_U2_1 ( .A(npu_inst_pe_1_0_2_int_q_acc_1_), 
        .B(npu_inst_pe_1_0_2_n13), .CI(npu_inst_pe_1_0_2_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_0_2_sub_67_carry_2_), .S(npu_inst_pe_1_0_2_N66) );
  FA_X1 npu_inst_pe_1_0_2_add_69_U1_1 ( .A(npu_inst_pe_1_0_2_int_q_acc_1_), 
        .B(npu_inst_pe_1_0_2_int_data_1_), .CI(
        npu_inst_pe_1_0_2_add_69_carry_1_), .CO(
        npu_inst_pe_1_0_2_add_69_carry_2_), .S(npu_inst_pe_1_0_2_N74) );
  NAND3_X1 npu_inst_pe_1_0_2_U109 ( .A1(npu_inst_pe_1_0_2_n5), .A2(
        npu_inst_pe_1_0_2_n6), .A3(npu_inst_pe_1_0_2_n7), .ZN(
        npu_inst_pe_1_0_2_n44) );
  NAND3_X1 npu_inst_pe_1_0_2_U108 ( .A1(npu_inst_pe_1_0_2_n4), .A2(
        npu_inst_pe_1_0_2_n6), .A3(npu_inst_pe_1_0_2_n7), .ZN(
        npu_inst_pe_1_0_2_n40) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_0_2_n33), .CK(
        npu_inst_pe_1_0_2_net4516), .RN(npu_inst_pe_1_0_2_n8), .Q(
        npu_inst_pe_1_0_2_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_0_2_n34), .CK(
        npu_inst_pe_1_0_2_net4516), .RN(npu_inst_pe_1_0_2_n8), .Q(
        npu_inst_pe_1_0_2_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_0_2_n35), .CK(
        npu_inst_pe_1_0_2_net4516), .RN(npu_inst_pe_1_0_2_n8), .Q(
        npu_inst_pe_1_0_2_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_0_2_n36), .CK(
        npu_inst_pe_1_0_2_net4516), .RN(npu_inst_pe_1_0_2_n8), .Q(
        npu_inst_pe_1_0_2_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_0_2_n98), .CK(
        npu_inst_pe_1_0_2_net4516), .RN(npu_inst_pe_1_0_2_n8), .Q(
        npu_inst_pe_1_0_2_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_0_2_n99), .CK(
        npu_inst_pe_1_0_2_net4516), .RN(npu_inst_pe_1_0_2_n8), .Q(
        npu_inst_pe_1_0_2_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_0_2_n32), .CK(
        npu_inst_pe_1_0_2_net4516), .RN(npu_inst_pe_1_0_2_n8), .Q(
        npu_inst_pe_1_0_2_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_0_2_n100), 
        .CK(npu_inst_pe_1_0_2_net4516), .RN(npu_inst_pe_1_0_2_n8), .Q(
        npu_inst_pe_1_0_2_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_weight_reg_0_ ( .D(npu_inst_n113), .CK(
        npu_inst_pe_1_0_2_net4522), .RN(npu_inst_pe_1_0_2_n8), .Q(
        npu_inst_pe_1_0_2_int_q_weight_0_), .QN(npu_inst_pe_1_0_2_n27) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_weight_reg_1_ ( .D(npu_inst_n119), .CK(
        npu_inst_pe_1_0_2_net4522), .RN(npu_inst_pe_1_0_2_n8), .Q(
        npu_inst_pe_1_0_2_int_q_weight_1_), .QN(npu_inst_pe_1_0_2_n26) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_0_2_n112), 
        .CK(npu_inst_pe_1_0_2_net4522), .RN(npu_inst_pe_1_0_2_n8), .Q(
        npu_inst_pe_1_0_2_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_0_2_n106), 
        .CK(npu_inst_pe_1_0_2_net4522), .RN(npu_inst_pe_1_0_2_n8), .Q(
        npu_inst_pe_1_0_2_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_0_2_n111), 
        .CK(npu_inst_pe_1_0_2_net4522), .RN(npu_inst_pe_1_0_2_n9), .Q(
        npu_inst_pe_1_0_2_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_0_2_n105), 
        .CK(npu_inst_pe_1_0_2_net4522), .RN(npu_inst_pe_1_0_2_n9), .Q(
        npu_inst_pe_1_0_2_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_0_2_n110), 
        .CK(npu_inst_pe_1_0_2_net4522), .RN(npu_inst_pe_1_0_2_n9), .Q(
        npu_inst_pe_1_0_2_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_0_2_n104), 
        .CK(npu_inst_pe_1_0_2_net4522), .RN(npu_inst_pe_1_0_2_n9), .Q(
        npu_inst_pe_1_0_2_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_0_2_n109), 
        .CK(npu_inst_pe_1_0_2_net4522), .RN(npu_inst_pe_1_0_2_n9), .Q(
        npu_inst_pe_1_0_2_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_0_2_n103), 
        .CK(npu_inst_pe_1_0_2_net4522), .RN(npu_inst_pe_1_0_2_n9), .Q(
        npu_inst_pe_1_0_2_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_0_2_n108), 
        .CK(npu_inst_pe_1_0_2_net4522), .RN(npu_inst_pe_1_0_2_n9), .Q(
        npu_inst_pe_1_0_2_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_0_2_n102), 
        .CK(npu_inst_pe_1_0_2_net4522), .RN(npu_inst_pe_1_0_2_n9), .Q(
        npu_inst_pe_1_0_2_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_0_2_n107), 
        .CK(npu_inst_pe_1_0_2_net4522), .RN(npu_inst_pe_1_0_2_n9), .Q(
        npu_inst_pe_1_0_2_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_0_2_n101), 
        .CK(npu_inst_pe_1_0_2_net4522), .RN(npu_inst_pe_1_0_2_n9), .Q(
        npu_inst_pe_1_0_2_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_0_2_n86), 
        .CK(npu_inst_pe_1_0_2_net4522), .RN(npu_inst_pe_1_0_2_n9), .Q(
        npu_inst_pe_1_0_2_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_0_2_n87), 
        .CK(npu_inst_pe_1_0_2_net4522), .RN(npu_inst_pe_1_0_2_n9), .Q(
        npu_inst_pe_1_0_2_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_0_2_n88), 
        .CK(npu_inst_pe_1_0_2_net4522), .RN(npu_inst_pe_1_0_2_n10), .Q(
        npu_inst_pe_1_0_2_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_0_2_n89), 
        .CK(npu_inst_pe_1_0_2_net4522), .RN(npu_inst_pe_1_0_2_n10), .Q(
        npu_inst_pe_1_0_2_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_0_2_n90), 
        .CK(npu_inst_pe_1_0_2_net4522), .RN(npu_inst_pe_1_0_2_n10), .Q(
        npu_inst_pe_1_0_2_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_0_2_n91), 
        .CK(npu_inst_pe_1_0_2_net4522), .RN(npu_inst_pe_1_0_2_n10), .Q(
        npu_inst_pe_1_0_2_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_0_2_n92), 
        .CK(npu_inst_pe_1_0_2_net4522), .RN(npu_inst_pe_1_0_2_n10), .Q(
        npu_inst_pe_1_0_2_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_0_2_n93), 
        .CK(npu_inst_pe_1_0_2_net4522), .RN(npu_inst_pe_1_0_2_n10), .Q(
        npu_inst_pe_1_0_2_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_0_2_n94), 
        .CK(npu_inst_pe_1_0_2_net4522), .RN(npu_inst_pe_1_0_2_n10), .Q(
        npu_inst_pe_1_0_2_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_0_2_n95), 
        .CK(npu_inst_pe_1_0_2_net4522), .RN(npu_inst_pe_1_0_2_n10), .Q(
        npu_inst_pe_1_0_2_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_0_2_n96), 
        .CK(npu_inst_pe_1_0_2_net4522), .RN(npu_inst_pe_1_0_2_n10), .Q(
        npu_inst_pe_1_0_2_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_0_2_n97), 
        .CK(npu_inst_pe_1_0_2_net4522), .RN(npu_inst_pe_1_0_2_n10), .Q(
        npu_inst_pe_1_0_2_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_0_2_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_0_2_N84), .SE(1'b0), .GCK(npu_inst_pe_1_0_2_net4516) );
  CLKGATETST_X1 npu_inst_pe_1_0_2_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n66), .SE(1'b0), .GCK(npu_inst_pe_1_0_2_net4522) );
  MUX2_X1 npu_inst_pe_1_0_3_U162 ( .A(npu_inst_pe_1_0_3_n32), .B(
        npu_inst_pe_1_0_3_n29), .S(npu_inst_pe_1_0_3_n8), .Z(
        npu_inst_pe_1_0_3_N93) );
  MUX2_X1 npu_inst_pe_1_0_3_U161 ( .A(npu_inst_pe_1_0_3_n31), .B(
        npu_inst_pe_1_0_3_n30), .S(npu_inst_pe_1_0_3_n6), .Z(
        npu_inst_pe_1_0_3_n32) );
  MUX2_X1 npu_inst_pe_1_0_3_U160 ( .A(npu_inst_pe_1_0_3_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_0_3_int_q_reg_v_1__0_), .S(npu_inst_pe_1_0_3_n4), .Z(
        npu_inst_pe_1_0_3_n31) );
  MUX2_X1 npu_inst_pe_1_0_3_U159 ( .A(npu_inst_pe_1_0_3_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_0_3_int_q_reg_v_3__0_), .S(npu_inst_pe_1_0_3_n4), .Z(
        npu_inst_pe_1_0_3_n30) );
  MUX2_X1 npu_inst_pe_1_0_3_U158 ( .A(npu_inst_pe_1_0_3_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_0_3_int_q_reg_v_5__0_), .S(npu_inst_pe_1_0_3_n4), .Z(
        npu_inst_pe_1_0_3_n29) );
  MUX2_X1 npu_inst_pe_1_0_3_U157 ( .A(npu_inst_pe_1_0_3_n28), .B(
        npu_inst_pe_1_0_3_n23), .S(npu_inst_pe_1_0_3_n8), .Z(
        npu_inst_pe_1_0_3_N94) );
  MUX2_X1 npu_inst_pe_1_0_3_U156 ( .A(npu_inst_pe_1_0_3_n25), .B(
        npu_inst_pe_1_0_3_n24), .S(npu_inst_pe_1_0_3_n6), .Z(
        npu_inst_pe_1_0_3_n28) );
  MUX2_X1 npu_inst_pe_1_0_3_U155 ( .A(npu_inst_pe_1_0_3_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_0_3_int_q_reg_v_1__1_), .S(npu_inst_pe_1_0_3_n4), .Z(
        npu_inst_pe_1_0_3_n25) );
  MUX2_X1 npu_inst_pe_1_0_3_U154 ( .A(npu_inst_pe_1_0_3_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_0_3_int_q_reg_v_3__1_), .S(npu_inst_pe_1_0_3_n4), .Z(
        npu_inst_pe_1_0_3_n24) );
  MUX2_X1 npu_inst_pe_1_0_3_U153 ( .A(npu_inst_pe_1_0_3_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_0_3_int_q_reg_v_5__1_), .S(npu_inst_pe_1_0_3_n4), .Z(
        npu_inst_pe_1_0_3_n23) );
  MUX2_X1 npu_inst_pe_1_0_3_U152 ( .A(npu_inst_pe_1_0_3_n22), .B(
        npu_inst_pe_1_0_3_n19), .S(npu_inst_pe_1_0_3_n8), .Z(
        npu_inst_int_data_x_0__3__1_) );
  MUX2_X1 npu_inst_pe_1_0_3_U151 ( .A(npu_inst_pe_1_0_3_n21), .B(
        npu_inst_pe_1_0_3_n20), .S(npu_inst_pe_1_0_3_n6), .Z(
        npu_inst_pe_1_0_3_n22) );
  MUX2_X1 npu_inst_pe_1_0_3_U150 ( .A(npu_inst_pe_1_0_3_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_0_3_int_q_reg_h_1__1_), .S(npu_inst_pe_1_0_3_n4), .Z(
        npu_inst_pe_1_0_3_n21) );
  MUX2_X1 npu_inst_pe_1_0_3_U149 ( .A(npu_inst_pe_1_0_3_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_0_3_int_q_reg_h_3__1_), .S(npu_inst_pe_1_0_3_n4), .Z(
        npu_inst_pe_1_0_3_n20) );
  MUX2_X1 npu_inst_pe_1_0_3_U148 ( .A(npu_inst_pe_1_0_3_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_0_3_int_q_reg_h_5__1_), .S(npu_inst_pe_1_0_3_n4), .Z(
        npu_inst_pe_1_0_3_n19) );
  MUX2_X1 npu_inst_pe_1_0_3_U147 ( .A(npu_inst_pe_1_0_3_n18), .B(
        npu_inst_pe_1_0_3_n15), .S(npu_inst_pe_1_0_3_n8), .Z(
        npu_inst_int_data_x_0__3__0_) );
  MUX2_X1 npu_inst_pe_1_0_3_U146 ( .A(npu_inst_pe_1_0_3_n17), .B(
        npu_inst_pe_1_0_3_n16), .S(npu_inst_pe_1_0_3_n6), .Z(
        npu_inst_pe_1_0_3_n18) );
  MUX2_X1 npu_inst_pe_1_0_3_U145 ( .A(npu_inst_pe_1_0_3_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_0_3_int_q_reg_h_1__0_), .S(npu_inst_pe_1_0_3_n4), .Z(
        npu_inst_pe_1_0_3_n17) );
  MUX2_X1 npu_inst_pe_1_0_3_U144 ( .A(npu_inst_pe_1_0_3_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_0_3_int_q_reg_h_3__0_), .S(npu_inst_pe_1_0_3_n4), .Z(
        npu_inst_pe_1_0_3_n16) );
  MUX2_X1 npu_inst_pe_1_0_3_U143 ( .A(npu_inst_pe_1_0_3_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_0_3_int_q_reg_h_5__0_), .S(npu_inst_pe_1_0_3_n4), .Z(
        npu_inst_pe_1_0_3_n15) );
  XOR2_X1 npu_inst_pe_1_0_3_U142 ( .A(npu_inst_pe_1_0_3_int_data_0_), .B(
        npu_inst_pe_1_0_3_int_q_acc_0_), .Z(npu_inst_pe_1_0_3_N73) );
  AND2_X1 npu_inst_pe_1_0_3_U141 ( .A1(npu_inst_pe_1_0_3_int_q_acc_0_), .A2(
        npu_inst_pe_1_0_3_int_data_0_), .ZN(npu_inst_pe_1_0_3_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_0_3_U140 ( .A(npu_inst_pe_1_0_3_int_q_acc_0_), .B(
        npu_inst_pe_1_0_3_n13), .ZN(npu_inst_pe_1_0_3_N65) );
  OR2_X1 npu_inst_pe_1_0_3_U139 ( .A1(npu_inst_pe_1_0_3_n13), .A2(
        npu_inst_pe_1_0_3_int_q_acc_0_), .ZN(npu_inst_pe_1_0_3_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_0_3_U138 ( .A(npu_inst_pe_1_0_3_int_q_acc_2_), .B(
        npu_inst_pe_1_0_3_add_69_carry_2_), .Z(npu_inst_pe_1_0_3_N75) );
  AND2_X1 npu_inst_pe_1_0_3_U137 ( .A1(npu_inst_pe_1_0_3_add_69_carry_2_), 
        .A2(npu_inst_pe_1_0_3_int_q_acc_2_), .ZN(
        npu_inst_pe_1_0_3_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_0_3_U136 ( .A(npu_inst_pe_1_0_3_int_q_acc_3_), .B(
        npu_inst_pe_1_0_3_add_69_carry_3_), .Z(npu_inst_pe_1_0_3_N76) );
  AND2_X1 npu_inst_pe_1_0_3_U135 ( .A1(npu_inst_pe_1_0_3_add_69_carry_3_), 
        .A2(npu_inst_pe_1_0_3_int_q_acc_3_), .ZN(
        npu_inst_pe_1_0_3_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_0_3_U134 ( .A(npu_inst_pe_1_0_3_int_q_acc_4_), .B(
        npu_inst_pe_1_0_3_add_69_carry_4_), .Z(npu_inst_pe_1_0_3_N77) );
  AND2_X1 npu_inst_pe_1_0_3_U133 ( .A1(npu_inst_pe_1_0_3_add_69_carry_4_), 
        .A2(npu_inst_pe_1_0_3_int_q_acc_4_), .ZN(
        npu_inst_pe_1_0_3_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_0_3_U132 ( .A(npu_inst_pe_1_0_3_int_q_acc_5_), .B(
        npu_inst_pe_1_0_3_add_69_carry_5_), .Z(npu_inst_pe_1_0_3_N78) );
  AND2_X1 npu_inst_pe_1_0_3_U131 ( .A1(npu_inst_pe_1_0_3_add_69_carry_5_), 
        .A2(npu_inst_pe_1_0_3_int_q_acc_5_), .ZN(
        npu_inst_pe_1_0_3_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_0_3_U130 ( .A(npu_inst_pe_1_0_3_int_q_acc_6_), .B(
        npu_inst_pe_1_0_3_add_69_carry_6_), .Z(npu_inst_pe_1_0_3_N79) );
  AND2_X1 npu_inst_pe_1_0_3_U129 ( .A1(npu_inst_pe_1_0_3_add_69_carry_6_), 
        .A2(npu_inst_pe_1_0_3_int_q_acc_6_), .ZN(
        npu_inst_pe_1_0_3_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_0_3_U128 ( .A(npu_inst_pe_1_0_3_int_q_acc_7_), .B(
        npu_inst_pe_1_0_3_add_69_carry_7_), .Z(npu_inst_pe_1_0_3_N80) );
  XNOR2_X1 npu_inst_pe_1_0_3_U127 ( .A(npu_inst_pe_1_0_3_sub_67_carry_2_), .B(
        npu_inst_pe_1_0_3_int_q_acc_2_), .ZN(npu_inst_pe_1_0_3_N67) );
  OR2_X1 npu_inst_pe_1_0_3_U126 ( .A1(npu_inst_pe_1_0_3_int_q_acc_2_), .A2(
        npu_inst_pe_1_0_3_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_0_3_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_0_3_U125 ( .A(npu_inst_pe_1_0_3_sub_67_carry_3_), .B(
        npu_inst_pe_1_0_3_int_q_acc_3_), .ZN(npu_inst_pe_1_0_3_N68) );
  OR2_X1 npu_inst_pe_1_0_3_U124 ( .A1(npu_inst_pe_1_0_3_int_q_acc_3_), .A2(
        npu_inst_pe_1_0_3_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_0_3_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_0_3_U123 ( .A(npu_inst_pe_1_0_3_sub_67_carry_4_), .B(
        npu_inst_pe_1_0_3_int_q_acc_4_), .ZN(npu_inst_pe_1_0_3_N69) );
  OR2_X1 npu_inst_pe_1_0_3_U122 ( .A1(npu_inst_pe_1_0_3_int_q_acc_4_), .A2(
        npu_inst_pe_1_0_3_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_0_3_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_0_3_U121 ( .A(npu_inst_pe_1_0_3_sub_67_carry_5_), .B(
        npu_inst_pe_1_0_3_int_q_acc_5_), .ZN(npu_inst_pe_1_0_3_N70) );
  OR2_X1 npu_inst_pe_1_0_3_U120 ( .A1(npu_inst_pe_1_0_3_int_q_acc_5_), .A2(
        npu_inst_pe_1_0_3_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_0_3_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_0_3_U119 ( .A(npu_inst_pe_1_0_3_sub_67_carry_6_), .B(
        npu_inst_pe_1_0_3_int_q_acc_6_), .ZN(npu_inst_pe_1_0_3_N71) );
  OR2_X1 npu_inst_pe_1_0_3_U118 ( .A1(npu_inst_pe_1_0_3_int_q_acc_6_), .A2(
        npu_inst_pe_1_0_3_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_0_3_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_0_3_U117 ( .A(npu_inst_pe_1_0_3_int_q_acc_7_), .B(
        npu_inst_pe_1_0_3_sub_67_carry_7_), .ZN(npu_inst_pe_1_0_3_N72) );
  INV_X1 npu_inst_pe_1_0_3_U116 ( .A(npu_inst_n80), .ZN(npu_inst_pe_1_0_3_n7)
         );
  INV_X1 npu_inst_pe_1_0_3_U115 ( .A(npu_inst_pe_1_0_3_n7), .ZN(
        npu_inst_pe_1_0_3_n6) );
  INV_X1 npu_inst_pe_1_0_3_U114 ( .A(npu_inst_n60), .ZN(npu_inst_pe_1_0_3_n3)
         );
  AOI22_X1 npu_inst_pe_1_0_3_U113 ( .A1(npu_inst_int_data_y_1__3__0_), .A2(
        npu_inst_pe_1_0_3_n58), .B1(npu_inst_pe_1_0_3_n119), .B2(
        npu_inst_pe_1_0_3_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_0_3_n57) );
  INV_X1 npu_inst_pe_1_0_3_U112 ( .A(npu_inst_pe_1_0_3_n57), .ZN(
        npu_inst_pe_1_0_3_n108) );
  AOI22_X1 npu_inst_pe_1_0_3_U111 ( .A1(npu_inst_int_data_y_1__3__0_), .A2(
        npu_inst_pe_1_0_3_n54), .B1(npu_inst_pe_1_0_3_n118), .B2(
        npu_inst_pe_1_0_3_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_0_3_n53) );
  INV_X1 npu_inst_pe_1_0_3_U110 ( .A(npu_inst_pe_1_0_3_n53), .ZN(
        npu_inst_pe_1_0_3_n109) );
  AOI22_X1 npu_inst_pe_1_0_3_U107 ( .A1(npu_inst_int_data_y_1__3__0_), .A2(
        npu_inst_pe_1_0_3_n50), .B1(npu_inst_pe_1_0_3_n117), .B2(
        npu_inst_pe_1_0_3_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_0_3_n49) );
  INV_X1 npu_inst_pe_1_0_3_U106 ( .A(npu_inst_pe_1_0_3_n49), .ZN(
        npu_inst_pe_1_0_3_n110) );
  AOI22_X1 npu_inst_pe_1_0_3_U105 ( .A1(npu_inst_int_data_y_1__3__0_), .A2(
        npu_inst_pe_1_0_3_n46), .B1(npu_inst_pe_1_0_3_n116), .B2(
        npu_inst_pe_1_0_3_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_0_3_n45) );
  INV_X1 npu_inst_pe_1_0_3_U104 ( .A(npu_inst_pe_1_0_3_n45), .ZN(
        npu_inst_pe_1_0_3_n111) );
  AOI22_X1 npu_inst_pe_1_0_3_U103 ( .A1(npu_inst_int_data_y_1__3__0_), .A2(
        npu_inst_pe_1_0_3_n42), .B1(npu_inst_pe_1_0_3_n115), .B2(
        npu_inst_pe_1_0_3_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_0_3_n41) );
  INV_X1 npu_inst_pe_1_0_3_U102 ( .A(npu_inst_pe_1_0_3_n41), .ZN(
        npu_inst_pe_1_0_3_n112) );
  AOI22_X1 npu_inst_pe_1_0_3_U101 ( .A1(npu_inst_int_data_y_1__3__1_), .A2(
        npu_inst_pe_1_0_3_n58), .B1(npu_inst_pe_1_0_3_n119), .B2(
        npu_inst_pe_1_0_3_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_0_3_n59) );
  INV_X1 npu_inst_pe_1_0_3_U100 ( .A(npu_inst_pe_1_0_3_n59), .ZN(
        npu_inst_pe_1_0_3_n102) );
  AOI22_X1 npu_inst_pe_1_0_3_U99 ( .A1(npu_inst_int_data_y_1__3__1_), .A2(
        npu_inst_pe_1_0_3_n54), .B1(npu_inst_pe_1_0_3_n118), .B2(
        npu_inst_pe_1_0_3_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_0_3_n55) );
  INV_X1 npu_inst_pe_1_0_3_U98 ( .A(npu_inst_pe_1_0_3_n55), .ZN(
        npu_inst_pe_1_0_3_n103) );
  AOI22_X1 npu_inst_pe_1_0_3_U97 ( .A1(npu_inst_int_data_y_1__3__1_), .A2(
        npu_inst_pe_1_0_3_n50), .B1(npu_inst_pe_1_0_3_n117), .B2(
        npu_inst_pe_1_0_3_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_0_3_n51) );
  INV_X1 npu_inst_pe_1_0_3_U96 ( .A(npu_inst_pe_1_0_3_n51), .ZN(
        npu_inst_pe_1_0_3_n104) );
  AOI22_X1 npu_inst_pe_1_0_3_U95 ( .A1(npu_inst_int_data_y_1__3__1_), .A2(
        npu_inst_pe_1_0_3_n46), .B1(npu_inst_pe_1_0_3_n116), .B2(
        npu_inst_pe_1_0_3_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_0_3_n47) );
  INV_X1 npu_inst_pe_1_0_3_U94 ( .A(npu_inst_pe_1_0_3_n47), .ZN(
        npu_inst_pe_1_0_3_n105) );
  AOI22_X1 npu_inst_pe_1_0_3_U93 ( .A1(npu_inst_int_data_y_1__3__1_), .A2(
        npu_inst_pe_1_0_3_n42), .B1(npu_inst_pe_1_0_3_n115), .B2(
        npu_inst_pe_1_0_3_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_0_3_n43) );
  INV_X1 npu_inst_pe_1_0_3_U92 ( .A(npu_inst_pe_1_0_3_n43), .ZN(
        npu_inst_pe_1_0_3_n106) );
  AOI22_X1 npu_inst_pe_1_0_3_U91 ( .A1(npu_inst_pe_1_0_3_n38), .A2(
        npu_inst_int_data_y_1__3__1_), .B1(npu_inst_pe_1_0_3_n114), .B2(
        npu_inst_pe_1_0_3_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_0_3_n39) );
  INV_X1 npu_inst_pe_1_0_3_U90 ( .A(npu_inst_pe_1_0_3_n39), .ZN(
        npu_inst_pe_1_0_3_n107) );
  AOI22_X1 npu_inst_pe_1_0_3_U89 ( .A1(npu_inst_pe_1_0_3_n38), .A2(
        npu_inst_int_data_y_1__3__0_), .B1(npu_inst_pe_1_0_3_n114), .B2(
        npu_inst_pe_1_0_3_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_0_3_n37) );
  INV_X1 npu_inst_pe_1_0_3_U88 ( .A(npu_inst_pe_1_0_3_n37), .ZN(
        npu_inst_pe_1_0_3_n113) );
  NAND2_X1 npu_inst_pe_1_0_3_U87 ( .A1(npu_inst_pe_1_0_3_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_0_3_n60), .ZN(npu_inst_pe_1_0_3_n74) );
  OAI21_X1 npu_inst_pe_1_0_3_U86 ( .B1(npu_inst_pe_1_0_3_n63), .B2(
        npu_inst_pe_1_0_3_n60), .A(npu_inst_pe_1_0_3_n74), .ZN(
        npu_inst_pe_1_0_3_n97) );
  NAND2_X1 npu_inst_pe_1_0_3_U85 ( .A1(npu_inst_pe_1_0_3_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_0_3_n60), .ZN(npu_inst_pe_1_0_3_n73) );
  OAI21_X1 npu_inst_pe_1_0_3_U84 ( .B1(npu_inst_pe_1_0_3_n61), .B2(
        npu_inst_pe_1_0_3_n60), .A(npu_inst_pe_1_0_3_n73), .ZN(
        npu_inst_pe_1_0_3_n96) );
  NAND2_X1 npu_inst_pe_1_0_3_U83 ( .A1(npu_inst_pe_1_0_3_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_0_3_n56), .ZN(npu_inst_pe_1_0_3_n72) );
  OAI21_X1 npu_inst_pe_1_0_3_U82 ( .B1(npu_inst_pe_1_0_3_n63), .B2(
        npu_inst_pe_1_0_3_n56), .A(npu_inst_pe_1_0_3_n72), .ZN(
        npu_inst_pe_1_0_3_n95) );
  NAND2_X1 npu_inst_pe_1_0_3_U81 ( .A1(npu_inst_pe_1_0_3_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_0_3_n56), .ZN(npu_inst_pe_1_0_3_n71) );
  OAI21_X1 npu_inst_pe_1_0_3_U80 ( .B1(npu_inst_pe_1_0_3_n61), .B2(
        npu_inst_pe_1_0_3_n56), .A(npu_inst_pe_1_0_3_n71), .ZN(
        npu_inst_pe_1_0_3_n94) );
  NAND2_X1 npu_inst_pe_1_0_3_U79 ( .A1(npu_inst_pe_1_0_3_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_0_3_n52), .ZN(npu_inst_pe_1_0_3_n70) );
  OAI21_X1 npu_inst_pe_1_0_3_U78 ( .B1(npu_inst_pe_1_0_3_n63), .B2(
        npu_inst_pe_1_0_3_n52), .A(npu_inst_pe_1_0_3_n70), .ZN(
        npu_inst_pe_1_0_3_n93) );
  NAND2_X1 npu_inst_pe_1_0_3_U77 ( .A1(npu_inst_pe_1_0_3_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_0_3_n52), .ZN(npu_inst_pe_1_0_3_n69) );
  OAI21_X1 npu_inst_pe_1_0_3_U76 ( .B1(npu_inst_pe_1_0_3_n61), .B2(
        npu_inst_pe_1_0_3_n52), .A(npu_inst_pe_1_0_3_n69), .ZN(
        npu_inst_pe_1_0_3_n92) );
  NAND2_X1 npu_inst_pe_1_0_3_U75 ( .A1(npu_inst_pe_1_0_3_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_0_3_n48), .ZN(npu_inst_pe_1_0_3_n68) );
  OAI21_X1 npu_inst_pe_1_0_3_U74 ( .B1(npu_inst_pe_1_0_3_n63), .B2(
        npu_inst_pe_1_0_3_n48), .A(npu_inst_pe_1_0_3_n68), .ZN(
        npu_inst_pe_1_0_3_n91) );
  NAND2_X1 npu_inst_pe_1_0_3_U73 ( .A1(npu_inst_pe_1_0_3_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_0_3_n48), .ZN(npu_inst_pe_1_0_3_n67) );
  OAI21_X1 npu_inst_pe_1_0_3_U72 ( .B1(npu_inst_pe_1_0_3_n61), .B2(
        npu_inst_pe_1_0_3_n48), .A(npu_inst_pe_1_0_3_n67), .ZN(
        npu_inst_pe_1_0_3_n90) );
  NAND2_X1 npu_inst_pe_1_0_3_U71 ( .A1(npu_inst_pe_1_0_3_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_0_3_n44), .ZN(npu_inst_pe_1_0_3_n66) );
  OAI21_X1 npu_inst_pe_1_0_3_U70 ( .B1(npu_inst_pe_1_0_3_n63), .B2(
        npu_inst_pe_1_0_3_n44), .A(npu_inst_pe_1_0_3_n66), .ZN(
        npu_inst_pe_1_0_3_n89) );
  NAND2_X1 npu_inst_pe_1_0_3_U69 ( .A1(npu_inst_pe_1_0_3_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_0_3_n44), .ZN(npu_inst_pe_1_0_3_n65) );
  OAI21_X1 npu_inst_pe_1_0_3_U68 ( .B1(npu_inst_pe_1_0_3_n61), .B2(
        npu_inst_pe_1_0_3_n44), .A(npu_inst_pe_1_0_3_n65), .ZN(
        npu_inst_pe_1_0_3_n88) );
  NAND2_X1 npu_inst_pe_1_0_3_U67 ( .A1(npu_inst_pe_1_0_3_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_0_3_n40), .ZN(npu_inst_pe_1_0_3_n64) );
  OAI21_X1 npu_inst_pe_1_0_3_U66 ( .B1(npu_inst_pe_1_0_3_n63), .B2(
        npu_inst_pe_1_0_3_n40), .A(npu_inst_pe_1_0_3_n64), .ZN(
        npu_inst_pe_1_0_3_n87) );
  NAND2_X1 npu_inst_pe_1_0_3_U65 ( .A1(npu_inst_pe_1_0_3_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_0_3_n40), .ZN(npu_inst_pe_1_0_3_n62) );
  OAI21_X1 npu_inst_pe_1_0_3_U64 ( .B1(npu_inst_pe_1_0_3_n61), .B2(
        npu_inst_pe_1_0_3_n40), .A(npu_inst_pe_1_0_3_n62), .ZN(
        npu_inst_pe_1_0_3_n86) );
  AND2_X1 npu_inst_pe_1_0_3_U63 ( .A1(npu_inst_pe_1_0_3_int_q_acc_2_), .A2(
        npu_inst_pe_1_0_3_n1), .ZN(int_o_data_npu[34]) );
  AND2_X1 npu_inst_pe_1_0_3_U62 ( .A1(npu_inst_pe_1_0_3_int_q_acc_3_), .A2(
        npu_inst_pe_1_0_3_n2), .ZN(int_o_data_npu[35]) );
  NOR3_X1 npu_inst_pe_1_0_3_U61 ( .A1(npu_inst_pe_1_0_3_n26), .A2(npu_inst_n60), .A3(npu_inst_int_ckg[60]), .ZN(npu_inst_pe_1_0_3_n85) );
  OR2_X1 npu_inst_pe_1_0_3_U60 ( .A1(npu_inst_pe_1_0_3_n85), .A2(
        npu_inst_pe_1_0_3_n2), .ZN(npu_inst_pe_1_0_3_N84) );
  AND2_X1 npu_inst_pe_1_0_3_U59 ( .A1(npu_inst_pe_1_0_3_int_q_acc_6_), .A2(
        npu_inst_pe_1_0_3_n2), .ZN(int_o_data_npu[38]) );
  AND2_X1 npu_inst_pe_1_0_3_U58 ( .A1(npu_inst_pe_1_0_3_int_q_acc_5_), .A2(
        npu_inst_pe_1_0_3_n2), .ZN(int_o_data_npu[37]) );
  AND2_X1 npu_inst_pe_1_0_3_U57 ( .A1(npu_inst_pe_1_0_3_int_q_acc_4_), .A2(
        npu_inst_pe_1_0_3_n2), .ZN(int_o_data_npu[36]) );
  AOI222_X1 npu_inst_pe_1_0_3_U56 ( .A1(npu_inst_int_data_res_1__3__0_), .A2(
        npu_inst_pe_1_0_3_n1), .B1(npu_inst_pe_1_0_3_N73), .B2(
        npu_inst_pe_1_0_3_n76), .C1(npu_inst_pe_1_0_3_N65), .C2(
        npu_inst_pe_1_0_3_n77), .ZN(npu_inst_pe_1_0_3_n84) );
  INV_X1 npu_inst_pe_1_0_3_U55 ( .A(npu_inst_pe_1_0_3_n84), .ZN(
        npu_inst_pe_1_0_3_n101) );
  AOI222_X1 npu_inst_pe_1_0_3_U54 ( .A1(npu_inst_int_data_res_1__3__7_), .A2(
        npu_inst_pe_1_0_3_n1), .B1(npu_inst_pe_1_0_3_N80), .B2(
        npu_inst_pe_1_0_3_n76), .C1(npu_inst_pe_1_0_3_N72), .C2(
        npu_inst_pe_1_0_3_n77), .ZN(npu_inst_pe_1_0_3_n75) );
  INV_X1 npu_inst_pe_1_0_3_U53 ( .A(npu_inst_pe_1_0_3_n75), .ZN(
        npu_inst_pe_1_0_3_n33) );
  AOI222_X1 npu_inst_pe_1_0_3_U52 ( .A1(npu_inst_int_data_res_1__3__1_), .A2(
        npu_inst_pe_1_0_3_n1), .B1(npu_inst_pe_1_0_3_N74), .B2(
        npu_inst_pe_1_0_3_n76), .C1(npu_inst_pe_1_0_3_N66), .C2(
        npu_inst_pe_1_0_3_n77), .ZN(npu_inst_pe_1_0_3_n83) );
  INV_X1 npu_inst_pe_1_0_3_U51 ( .A(npu_inst_pe_1_0_3_n83), .ZN(
        npu_inst_pe_1_0_3_n100) );
  AOI222_X1 npu_inst_pe_1_0_3_U50 ( .A1(npu_inst_int_data_res_1__3__2_), .A2(
        npu_inst_pe_1_0_3_n1), .B1(npu_inst_pe_1_0_3_N75), .B2(
        npu_inst_pe_1_0_3_n76), .C1(npu_inst_pe_1_0_3_N67), .C2(
        npu_inst_pe_1_0_3_n77), .ZN(npu_inst_pe_1_0_3_n82) );
  INV_X1 npu_inst_pe_1_0_3_U49 ( .A(npu_inst_pe_1_0_3_n82), .ZN(
        npu_inst_pe_1_0_3_n99) );
  AOI222_X1 npu_inst_pe_1_0_3_U48 ( .A1(npu_inst_int_data_res_1__3__3_), .A2(
        npu_inst_pe_1_0_3_n1), .B1(npu_inst_pe_1_0_3_N76), .B2(
        npu_inst_pe_1_0_3_n76), .C1(npu_inst_pe_1_0_3_N68), .C2(
        npu_inst_pe_1_0_3_n77), .ZN(npu_inst_pe_1_0_3_n81) );
  INV_X1 npu_inst_pe_1_0_3_U47 ( .A(npu_inst_pe_1_0_3_n81), .ZN(
        npu_inst_pe_1_0_3_n98) );
  AOI222_X1 npu_inst_pe_1_0_3_U46 ( .A1(npu_inst_int_data_res_1__3__4_), .A2(
        npu_inst_pe_1_0_3_n1), .B1(npu_inst_pe_1_0_3_N77), .B2(
        npu_inst_pe_1_0_3_n76), .C1(npu_inst_pe_1_0_3_N69), .C2(
        npu_inst_pe_1_0_3_n77), .ZN(npu_inst_pe_1_0_3_n80) );
  INV_X1 npu_inst_pe_1_0_3_U45 ( .A(npu_inst_pe_1_0_3_n80), .ZN(
        npu_inst_pe_1_0_3_n36) );
  AOI222_X1 npu_inst_pe_1_0_3_U44 ( .A1(npu_inst_int_data_res_1__3__5_), .A2(
        npu_inst_pe_1_0_3_n1), .B1(npu_inst_pe_1_0_3_N78), .B2(
        npu_inst_pe_1_0_3_n76), .C1(npu_inst_pe_1_0_3_N70), .C2(
        npu_inst_pe_1_0_3_n77), .ZN(npu_inst_pe_1_0_3_n79) );
  INV_X1 npu_inst_pe_1_0_3_U43 ( .A(npu_inst_pe_1_0_3_n79), .ZN(
        npu_inst_pe_1_0_3_n35) );
  AOI222_X1 npu_inst_pe_1_0_3_U42 ( .A1(npu_inst_int_data_res_1__3__6_), .A2(
        npu_inst_pe_1_0_3_n1), .B1(npu_inst_pe_1_0_3_N79), .B2(
        npu_inst_pe_1_0_3_n76), .C1(npu_inst_pe_1_0_3_N71), .C2(
        npu_inst_pe_1_0_3_n77), .ZN(npu_inst_pe_1_0_3_n78) );
  INV_X1 npu_inst_pe_1_0_3_U41 ( .A(npu_inst_pe_1_0_3_n78), .ZN(
        npu_inst_pe_1_0_3_n34) );
  INV_X1 npu_inst_pe_1_0_3_U40 ( .A(npu_inst_pe_1_0_3_int_data_1_), .ZN(
        npu_inst_pe_1_0_3_n14) );
  AND2_X1 npu_inst_pe_1_0_3_U39 ( .A1(npu_inst_int_data_x_0__3__1_), .A2(
        npu_inst_pe_1_0_3_int_q_weight_1_), .ZN(npu_inst_pe_1_0_3_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_0_3_U38 ( .A1(npu_inst_int_data_x_0__3__0_), .A2(
        npu_inst_pe_1_0_3_int_q_weight_1_), .ZN(npu_inst_pe_1_0_3_int_data_0_)
         );
  AND2_X1 npu_inst_pe_1_0_3_U37 ( .A1(npu_inst_pe_1_0_3_n2), .A2(
        npu_inst_pe_1_0_3_int_q_acc_7_), .ZN(int_o_data_npu[39]) );
  AND2_X1 npu_inst_pe_1_0_3_U36 ( .A1(npu_inst_pe_1_0_3_int_q_acc_1_), .A2(
        npu_inst_pe_1_0_3_n1), .ZN(int_o_data_npu[33]) );
  AND2_X1 npu_inst_pe_1_0_3_U35 ( .A1(npu_inst_pe_1_0_3_int_q_acc_0_), .A2(
        npu_inst_pe_1_0_3_n1), .ZN(int_o_data_npu[32]) );
  AND2_X1 npu_inst_pe_1_0_3_U34 ( .A1(npu_inst_pe_1_0_3_N93), .A2(npu_inst_n60), .ZN(npu_inst_pe_1_0_3_o_data_v_0_) );
  AND2_X1 npu_inst_pe_1_0_3_U33 ( .A1(npu_inst_n60), .A2(npu_inst_pe_1_0_3_N94), .ZN(npu_inst_pe_1_0_3_o_data_v_1_) );
  AOI22_X1 npu_inst_pe_1_0_3_U32 ( .A1(npu_inst_n60), .A2(
        npu_inst_int_data_y_1__3__1_), .B1(npu_inst_pe_1_0_3_n3), .B2(
        npu_inst_int_data_x_0__4__1_), .ZN(npu_inst_pe_1_0_3_n63) );
  AOI22_X1 npu_inst_pe_1_0_3_U31 ( .A1(npu_inst_n60), .A2(
        npu_inst_int_data_y_1__3__0_), .B1(npu_inst_pe_1_0_3_n3), .B2(
        npu_inst_int_data_x_0__4__0_), .ZN(npu_inst_pe_1_0_3_n61) );
  INV_X1 npu_inst_pe_1_0_3_U30 ( .A(npu_inst_pe_1_0_3_int_data_0_), .ZN(
        npu_inst_pe_1_0_3_n13) );
  INV_X1 npu_inst_pe_1_0_3_U29 ( .A(npu_inst_n72), .ZN(npu_inst_pe_1_0_3_n5)
         );
  OR3_X1 npu_inst_pe_1_0_3_U28 ( .A1(npu_inst_pe_1_0_3_n6), .A2(
        npu_inst_pe_1_0_3_n8), .A3(npu_inst_pe_1_0_3_n5), .ZN(
        npu_inst_pe_1_0_3_n56) );
  OR3_X1 npu_inst_pe_1_0_3_U27 ( .A1(npu_inst_pe_1_0_3_n5), .A2(
        npu_inst_pe_1_0_3_n8), .A3(npu_inst_pe_1_0_3_n7), .ZN(
        npu_inst_pe_1_0_3_n48) );
  INV_X1 npu_inst_pe_1_0_3_U26 ( .A(npu_inst_pe_1_0_3_n5), .ZN(
        npu_inst_pe_1_0_3_n4) );
  OR3_X1 npu_inst_pe_1_0_3_U25 ( .A1(npu_inst_pe_1_0_3_n4), .A2(
        npu_inst_pe_1_0_3_n8), .A3(npu_inst_pe_1_0_3_n7), .ZN(
        npu_inst_pe_1_0_3_n52) );
  OR3_X1 npu_inst_pe_1_0_3_U24 ( .A1(npu_inst_pe_1_0_3_n6), .A2(
        npu_inst_pe_1_0_3_n8), .A3(npu_inst_pe_1_0_3_n4), .ZN(
        npu_inst_pe_1_0_3_n60) );
  NOR2_X1 npu_inst_pe_1_0_3_U23 ( .A1(npu_inst_pe_1_0_3_n60), .A2(
        npu_inst_pe_1_0_3_n3), .ZN(npu_inst_pe_1_0_3_n58) );
  NOR2_X1 npu_inst_pe_1_0_3_U22 ( .A1(npu_inst_pe_1_0_3_n56), .A2(
        npu_inst_pe_1_0_3_n3), .ZN(npu_inst_pe_1_0_3_n54) );
  NOR2_X1 npu_inst_pe_1_0_3_U21 ( .A1(npu_inst_pe_1_0_3_n52), .A2(
        npu_inst_pe_1_0_3_n3), .ZN(npu_inst_pe_1_0_3_n50) );
  NOR2_X1 npu_inst_pe_1_0_3_U20 ( .A1(npu_inst_pe_1_0_3_n48), .A2(
        npu_inst_pe_1_0_3_n3), .ZN(npu_inst_pe_1_0_3_n46) );
  NOR2_X1 npu_inst_pe_1_0_3_U19 ( .A1(npu_inst_pe_1_0_3_n40), .A2(
        npu_inst_pe_1_0_3_n3), .ZN(npu_inst_pe_1_0_3_n38) );
  NOR2_X1 npu_inst_pe_1_0_3_U18 ( .A1(npu_inst_pe_1_0_3_n44), .A2(
        npu_inst_pe_1_0_3_n3), .ZN(npu_inst_pe_1_0_3_n42) );
  BUF_X1 npu_inst_pe_1_0_3_U17 ( .A(npu_inst_n107), .Z(npu_inst_pe_1_0_3_n8)
         );
  INV_X1 npu_inst_pe_1_0_3_U16 ( .A(npu_inst_n127), .ZN(npu_inst_pe_1_0_3_n12)
         );
  INV_X1 npu_inst_pe_1_0_3_U15 ( .A(npu_inst_pe_1_0_3_n38), .ZN(
        npu_inst_pe_1_0_3_n114) );
  INV_X1 npu_inst_pe_1_0_3_U14 ( .A(npu_inst_pe_1_0_3_n58), .ZN(
        npu_inst_pe_1_0_3_n119) );
  INV_X1 npu_inst_pe_1_0_3_U13 ( .A(npu_inst_pe_1_0_3_n54), .ZN(
        npu_inst_pe_1_0_3_n118) );
  INV_X1 npu_inst_pe_1_0_3_U12 ( .A(npu_inst_pe_1_0_3_n50), .ZN(
        npu_inst_pe_1_0_3_n117) );
  INV_X1 npu_inst_pe_1_0_3_U11 ( .A(npu_inst_pe_1_0_3_n46), .ZN(
        npu_inst_pe_1_0_3_n116) );
  INV_X1 npu_inst_pe_1_0_3_U10 ( .A(npu_inst_pe_1_0_3_n42), .ZN(
        npu_inst_pe_1_0_3_n115) );
  BUF_X1 npu_inst_pe_1_0_3_U9 ( .A(npu_inst_n37), .Z(npu_inst_pe_1_0_3_n2) );
  BUF_X1 npu_inst_pe_1_0_3_U8 ( .A(npu_inst_n37), .Z(npu_inst_pe_1_0_3_n1) );
  BUF_X1 npu_inst_pe_1_0_3_U7 ( .A(npu_inst_pe_1_0_3_n12), .Z(
        npu_inst_pe_1_0_3_n11) );
  BUF_X1 npu_inst_pe_1_0_3_U6 ( .A(npu_inst_pe_1_0_3_n12), .Z(
        npu_inst_pe_1_0_3_n10) );
  BUF_X1 npu_inst_pe_1_0_3_U5 ( .A(npu_inst_pe_1_0_3_n12), .Z(
        npu_inst_pe_1_0_3_n9) );
  NOR2_X1 npu_inst_pe_1_0_3_U4 ( .A1(npu_inst_pe_1_0_3_int_q_weight_0_), .A2(
        npu_inst_pe_1_0_3_n1), .ZN(npu_inst_pe_1_0_3_n76) );
  NOR2_X1 npu_inst_pe_1_0_3_U3 ( .A1(npu_inst_pe_1_0_3_n27), .A2(
        npu_inst_pe_1_0_3_n1), .ZN(npu_inst_pe_1_0_3_n77) );
  FA_X1 npu_inst_pe_1_0_3_sub_67_U2_1 ( .A(npu_inst_pe_1_0_3_int_q_acc_1_), 
        .B(npu_inst_pe_1_0_3_n14), .CI(npu_inst_pe_1_0_3_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_0_3_sub_67_carry_2_), .S(npu_inst_pe_1_0_3_N66) );
  FA_X1 npu_inst_pe_1_0_3_add_69_U1_1 ( .A(npu_inst_pe_1_0_3_int_q_acc_1_), 
        .B(npu_inst_pe_1_0_3_int_data_1_), .CI(
        npu_inst_pe_1_0_3_add_69_carry_1_), .CO(
        npu_inst_pe_1_0_3_add_69_carry_2_), .S(npu_inst_pe_1_0_3_N74) );
  NAND3_X1 npu_inst_pe_1_0_3_U109 ( .A1(npu_inst_pe_1_0_3_n5), .A2(
        npu_inst_pe_1_0_3_n7), .A3(npu_inst_pe_1_0_3_n8), .ZN(
        npu_inst_pe_1_0_3_n44) );
  NAND3_X1 npu_inst_pe_1_0_3_U108 ( .A1(npu_inst_pe_1_0_3_n4), .A2(
        npu_inst_pe_1_0_3_n7), .A3(npu_inst_pe_1_0_3_n8), .ZN(
        npu_inst_pe_1_0_3_n40) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_0_3_n34), .CK(
        npu_inst_pe_1_0_3_net4493), .RN(npu_inst_pe_1_0_3_n9), .Q(
        npu_inst_pe_1_0_3_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_0_3_n35), .CK(
        npu_inst_pe_1_0_3_net4493), .RN(npu_inst_pe_1_0_3_n9), .Q(
        npu_inst_pe_1_0_3_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_0_3_n36), .CK(
        npu_inst_pe_1_0_3_net4493), .RN(npu_inst_pe_1_0_3_n9), .Q(
        npu_inst_pe_1_0_3_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_0_3_n98), .CK(
        npu_inst_pe_1_0_3_net4493), .RN(npu_inst_pe_1_0_3_n9), .Q(
        npu_inst_pe_1_0_3_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_0_3_n99), .CK(
        npu_inst_pe_1_0_3_net4493), .RN(npu_inst_pe_1_0_3_n9), .Q(
        npu_inst_pe_1_0_3_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_0_3_n100), 
        .CK(npu_inst_pe_1_0_3_net4493), .RN(npu_inst_pe_1_0_3_n9), .Q(
        npu_inst_pe_1_0_3_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_0_3_n33), .CK(
        npu_inst_pe_1_0_3_net4493), .RN(npu_inst_pe_1_0_3_n9), .Q(
        npu_inst_pe_1_0_3_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_0_3_n101), 
        .CK(npu_inst_pe_1_0_3_net4493), .RN(npu_inst_pe_1_0_3_n9), .Q(
        npu_inst_pe_1_0_3_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_weight_reg_0_ ( .D(npu_inst_n113), .CK(
        npu_inst_pe_1_0_3_net4499), .RN(npu_inst_pe_1_0_3_n9), .Q(
        npu_inst_pe_1_0_3_int_q_weight_0_), .QN(npu_inst_pe_1_0_3_n27) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_weight_reg_1_ ( .D(npu_inst_n119), .CK(
        npu_inst_pe_1_0_3_net4499), .RN(npu_inst_pe_1_0_3_n9), .Q(
        npu_inst_pe_1_0_3_int_q_weight_1_), .QN(npu_inst_pe_1_0_3_n26) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_0_3_n113), 
        .CK(npu_inst_pe_1_0_3_net4499), .RN(npu_inst_pe_1_0_3_n9), .Q(
        npu_inst_pe_1_0_3_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_0_3_n107), 
        .CK(npu_inst_pe_1_0_3_net4499), .RN(npu_inst_pe_1_0_3_n9), .Q(
        npu_inst_pe_1_0_3_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_0_3_n112), 
        .CK(npu_inst_pe_1_0_3_net4499), .RN(npu_inst_pe_1_0_3_n10), .Q(
        npu_inst_pe_1_0_3_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_0_3_n106), 
        .CK(npu_inst_pe_1_0_3_net4499), .RN(npu_inst_pe_1_0_3_n10), .Q(
        npu_inst_pe_1_0_3_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_0_3_n111), 
        .CK(npu_inst_pe_1_0_3_net4499), .RN(npu_inst_pe_1_0_3_n10), .Q(
        npu_inst_pe_1_0_3_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_0_3_n105), 
        .CK(npu_inst_pe_1_0_3_net4499), .RN(npu_inst_pe_1_0_3_n10), .Q(
        npu_inst_pe_1_0_3_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_0_3_n110), 
        .CK(npu_inst_pe_1_0_3_net4499), .RN(npu_inst_pe_1_0_3_n10), .Q(
        npu_inst_pe_1_0_3_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_0_3_n104), 
        .CK(npu_inst_pe_1_0_3_net4499), .RN(npu_inst_pe_1_0_3_n10), .Q(
        npu_inst_pe_1_0_3_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_0_3_n109), 
        .CK(npu_inst_pe_1_0_3_net4499), .RN(npu_inst_pe_1_0_3_n10), .Q(
        npu_inst_pe_1_0_3_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_0_3_n103), 
        .CK(npu_inst_pe_1_0_3_net4499), .RN(npu_inst_pe_1_0_3_n10), .Q(
        npu_inst_pe_1_0_3_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_0_3_n108), 
        .CK(npu_inst_pe_1_0_3_net4499), .RN(npu_inst_pe_1_0_3_n10), .Q(
        npu_inst_pe_1_0_3_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_0_3_n102), 
        .CK(npu_inst_pe_1_0_3_net4499), .RN(npu_inst_pe_1_0_3_n10), .Q(
        npu_inst_pe_1_0_3_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_0_3_n86), 
        .CK(npu_inst_pe_1_0_3_net4499), .RN(npu_inst_pe_1_0_3_n10), .Q(
        npu_inst_pe_1_0_3_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_0_3_n87), 
        .CK(npu_inst_pe_1_0_3_net4499), .RN(npu_inst_pe_1_0_3_n10), .Q(
        npu_inst_pe_1_0_3_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_0_3_n88), 
        .CK(npu_inst_pe_1_0_3_net4499), .RN(npu_inst_pe_1_0_3_n11), .Q(
        npu_inst_pe_1_0_3_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_0_3_n89), 
        .CK(npu_inst_pe_1_0_3_net4499), .RN(npu_inst_pe_1_0_3_n11), .Q(
        npu_inst_pe_1_0_3_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_0_3_n90), 
        .CK(npu_inst_pe_1_0_3_net4499), .RN(npu_inst_pe_1_0_3_n11), .Q(
        npu_inst_pe_1_0_3_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_0_3_n91), 
        .CK(npu_inst_pe_1_0_3_net4499), .RN(npu_inst_pe_1_0_3_n11), .Q(
        npu_inst_pe_1_0_3_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_0_3_n92), 
        .CK(npu_inst_pe_1_0_3_net4499), .RN(npu_inst_pe_1_0_3_n11), .Q(
        npu_inst_pe_1_0_3_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_0_3_n93), 
        .CK(npu_inst_pe_1_0_3_net4499), .RN(npu_inst_pe_1_0_3_n11), .Q(
        npu_inst_pe_1_0_3_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_0_3_n94), 
        .CK(npu_inst_pe_1_0_3_net4499), .RN(npu_inst_pe_1_0_3_n11), .Q(
        npu_inst_pe_1_0_3_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_0_3_n95), 
        .CK(npu_inst_pe_1_0_3_net4499), .RN(npu_inst_pe_1_0_3_n11), .Q(
        npu_inst_pe_1_0_3_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_0_3_n96), 
        .CK(npu_inst_pe_1_0_3_net4499), .RN(npu_inst_pe_1_0_3_n11), .Q(
        npu_inst_pe_1_0_3_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_0_3_n97), 
        .CK(npu_inst_pe_1_0_3_net4499), .RN(npu_inst_pe_1_0_3_n11), .Q(
        npu_inst_pe_1_0_3_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_0_3_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_0_3_N84), .SE(1'b0), .GCK(npu_inst_pe_1_0_3_net4493) );
  CLKGATETST_X1 npu_inst_pe_1_0_3_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n66), .SE(1'b0), .GCK(npu_inst_pe_1_0_3_net4499) );
  MUX2_X1 npu_inst_pe_1_0_4_U161 ( .A(npu_inst_pe_1_0_4_n31), .B(
        npu_inst_pe_1_0_4_n28), .S(npu_inst_pe_1_0_4_n7), .Z(
        npu_inst_pe_1_0_4_N93) );
  MUX2_X1 npu_inst_pe_1_0_4_U160 ( .A(npu_inst_pe_1_0_4_n30), .B(
        npu_inst_pe_1_0_4_n29), .S(npu_inst_n79), .Z(npu_inst_pe_1_0_4_n31) );
  MUX2_X1 npu_inst_pe_1_0_4_U159 ( .A(npu_inst_pe_1_0_4_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_0_4_int_q_reg_v_1__0_), .S(npu_inst_pe_1_0_4_n4), .Z(
        npu_inst_pe_1_0_4_n30) );
  MUX2_X1 npu_inst_pe_1_0_4_U158 ( .A(npu_inst_pe_1_0_4_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_0_4_int_q_reg_v_3__0_), .S(npu_inst_pe_1_0_4_n4), .Z(
        npu_inst_pe_1_0_4_n29) );
  MUX2_X1 npu_inst_pe_1_0_4_U157 ( .A(npu_inst_pe_1_0_4_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_0_4_int_q_reg_v_5__0_), .S(npu_inst_pe_1_0_4_n4), .Z(
        npu_inst_pe_1_0_4_n28) );
  MUX2_X1 npu_inst_pe_1_0_4_U156 ( .A(npu_inst_pe_1_0_4_n25), .B(
        npu_inst_pe_1_0_4_n22), .S(npu_inst_pe_1_0_4_n7), .Z(
        npu_inst_pe_1_0_4_N94) );
  MUX2_X1 npu_inst_pe_1_0_4_U155 ( .A(npu_inst_pe_1_0_4_n24), .B(
        npu_inst_pe_1_0_4_n23), .S(npu_inst_n79), .Z(npu_inst_pe_1_0_4_n25) );
  MUX2_X1 npu_inst_pe_1_0_4_U154 ( .A(npu_inst_pe_1_0_4_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_0_4_int_q_reg_v_1__1_), .S(npu_inst_pe_1_0_4_n4), .Z(
        npu_inst_pe_1_0_4_n24) );
  MUX2_X1 npu_inst_pe_1_0_4_U153 ( .A(npu_inst_pe_1_0_4_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_0_4_int_q_reg_v_3__1_), .S(npu_inst_pe_1_0_4_n4), .Z(
        npu_inst_pe_1_0_4_n23) );
  MUX2_X1 npu_inst_pe_1_0_4_U152 ( .A(npu_inst_pe_1_0_4_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_0_4_int_q_reg_v_5__1_), .S(npu_inst_pe_1_0_4_n4), .Z(
        npu_inst_pe_1_0_4_n22) );
  MUX2_X1 npu_inst_pe_1_0_4_U151 ( .A(npu_inst_pe_1_0_4_n21), .B(
        npu_inst_pe_1_0_4_n18), .S(npu_inst_pe_1_0_4_n7), .Z(
        npu_inst_int_data_x_0__4__1_) );
  MUX2_X1 npu_inst_pe_1_0_4_U150 ( .A(npu_inst_pe_1_0_4_n20), .B(
        npu_inst_pe_1_0_4_n19), .S(npu_inst_n79), .Z(npu_inst_pe_1_0_4_n21) );
  MUX2_X1 npu_inst_pe_1_0_4_U149 ( .A(npu_inst_pe_1_0_4_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_0_4_int_q_reg_h_1__1_), .S(npu_inst_pe_1_0_4_n4), .Z(
        npu_inst_pe_1_0_4_n20) );
  MUX2_X1 npu_inst_pe_1_0_4_U148 ( .A(npu_inst_pe_1_0_4_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_0_4_int_q_reg_h_3__1_), .S(npu_inst_pe_1_0_4_n4), .Z(
        npu_inst_pe_1_0_4_n19) );
  MUX2_X1 npu_inst_pe_1_0_4_U147 ( .A(npu_inst_pe_1_0_4_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_0_4_int_q_reg_h_5__1_), .S(npu_inst_pe_1_0_4_n4), .Z(
        npu_inst_pe_1_0_4_n18) );
  MUX2_X1 npu_inst_pe_1_0_4_U146 ( .A(npu_inst_pe_1_0_4_n17), .B(
        npu_inst_pe_1_0_4_n14), .S(npu_inst_pe_1_0_4_n7), .Z(
        npu_inst_int_data_x_0__4__0_) );
  MUX2_X1 npu_inst_pe_1_0_4_U145 ( .A(npu_inst_pe_1_0_4_n16), .B(
        npu_inst_pe_1_0_4_n15), .S(npu_inst_n79), .Z(npu_inst_pe_1_0_4_n17) );
  MUX2_X1 npu_inst_pe_1_0_4_U144 ( .A(npu_inst_pe_1_0_4_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_0_4_int_q_reg_h_1__0_), .S(npu_inst_pe_1_0_4_n4), .Z(
        npu_inst_pe_1_0_4_n16) );
  MUX2_X1 npu_inst_pe_1_0_4_U143 ( .A(npu_inst_pe_1_0_4_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_0_4_int_q_reg_h_3__0_), .S(npu_inst_pe_1_0_4_n4), .Z(
        npu_inst_pe_1_0_4_n15) );
  MUX2_X1 npu_inst_pe_1_0_4_U142 ( .A(npu_inst_pe_1_0_4_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_0_4_int_q_reg_h_5__0_), .S(npu_inst_pe_1_0_4_n4), .Z(
        npu_inst_pe_1_0_4_n14) );
  XOR2_X1 npu_inst_pe_1_0_4_U141 ( .A(npu_inst_pe_1_0_4_int_data_0_), .B(
        npu_inst_pe_1_0_4_int_q_acc_0_), .Z(npu_inst_pe_1_0_4_N73) );
  AND2_X1 npu_inst_pe_1_0_4_U140 ( .A1(npu_inst_pe_1_0_4_int_q_acc_0_), .A2(
        npu_inst_pe_1_0_4_int_data_0_), .ZN(npu_inst_pe_1_0_4_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_0_4_U139 ( .A(npu_inst_pe_1_0_4_int_q_acc_0_), .B(
        npu_inst_pe_1_0_4_n12), .ZN(npu_inst_pe_1_0_4_N65) );
  OR2_X1 npu_inst_pe_1_0_4_U138 ( .A1(npu_inst_pe_1_0_4_n12), .A2(
        npu_inst_pe_1_0_4_int_q_acc_0_), .ZN(npu_inst_pe_1_0_4_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_0_4_U137 ( .A(npu_inst_pe_1_0_4_int_q_acc_2_), .B(
        npu_inst_pe_1_0_4_add_69_carry_2_), .Z(npu_inst_pe_1_0_4_N75) );
  AND2_X1 npu_inst_pe_1_0_4_U136 ( .A1(npu_inst_pe_1_0_4_add_69_carry_2_), 
        .A2(npu_inst_pe_1_0_4_int_q_acc_2_), .ZN(
        npu_inst_pe_1_0_4_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_0_4_U135 ( .A(npu_inst_pe_1_0_4_int_q_acc_3_), .B(
        npu_inst_pe_1_0_4_add_69_carry_3_), .Z(npu_inst_pe_1_0_4_N76) );
  AND2_X1 npu_inst_pe_1_0_4_U134 ( .A1(npu_inst_pe_1_0_4_add_69_carry_3_), 
        .A2(npu_inst_pe_1_0_4_int_q_acc_3_), .ZN(
        npu_inst_pe_1_0_4_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_0_4_U133 ( .A(npu_inst_pe_1_0_4_int_q_acc_4_), .B(
        npu_inst_pe_1_0_4_add_69_carry_4_), .Z(npu_inst_pe_1_0_4_N77) );
  AND2_X1 npu_inst_pe_1_0_4_U132 ( .A1(npu_inst_pe_1_0_4_add_69_carry_4_), 
        .A2(npu_inst_pe_1_0_4_int_q_acc_4_), .ZN(
        npu_inst_pe_1_0_4_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_0_4_U131 ( .A(npu_inst_pe_1_0_4_int_q_acc_5_), .B(
        npu_inst_pe_1_0_4_add_69_carry_5_), .Z(npu_inst_pe_1_0_4_N78) );
  AND2_X1 npu_inst_pe_1_0_4_U130 ( .A1(npu_inst_pe_1_0_4_add_69_carry_5_), 
        .A2(npu_inst_pe_1_0_4_int_q_acc_5_), .ZN(
        npu_inst_pe_1_0_4_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_0_4_U129 ( .A(npu_inst_pe_1_0_4_int_q_acc_6_), .B(
        npu_inst_pe_1_0_4_add_69_carry_6_), .Z(npu_inst_pe_1_0_4_N79) );
  AND2_X1 npu_inst_pe_1_0_4_U128 ( .A1(npu_inst_pe_1_0_4_add_69_carry_6_), 
        .A2(npu_inst_pe_1_0_4_int_q_acc_6_), .ZN(
        npu_inst_pe_1_0_4_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_0_4_U127 ( .A(npu_inst_pe_1_0_4_int_q_acc_7_), .B(
        npu_inst_pe_1_0_4_add_69_carry_7_), .Z(npu_inst_pe_1_0_4_N80) );
  XNOR2_X1 npu_inst_pe_1_0_4_U126 ( .A(npu_inst_pe_1_0_4_sub_67_carry_2_), .B(
        npu_inst_pe_1_0_4_int_q_acc_2_), .ZN(npu_inst_pe_1_0_4_N67) );
  OR2_X1 npu_inst_pe_1_0_4_U125 ( .A1(npu_inst_pe_1_0_4_int_q_acc_2_), .A2(
        npu_inst_pe_1_0_4_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_0_4_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_0_4_U124 ( .A(npu_inst_pe_1_0_4_sub_67_carry_3_), .B(
        npu_inst_pe_1_0_4_int_q_acc_3_), .ZN(npu_inst_pe_1_0_4_N68) );
  OR2_X1 npu_inst_pe_1_0_4_U123 ( .A1(npu_inst_pe_1_0_4_int_q_acc_3_), .A2(
        npu_inst_pe_1_0_4_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_0_4_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_0_4_U122 ( .A(npu_inst_pe_1_0_4_sub_67_carry_4_), .B(
        npu_inst_pe_1_0_4_int_q_acc_4_), .ZN(npu_inst_pe_1_0_4_N69) );
  OR2_X1 npu_inst_pe_1_0_4_U121 ( .A1(npu_inst_pe_1_0_4_int_q_acc_4_), .A2(
        npu_inst_pe_1_0_4_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_0_4_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_0_4_U120 ( .A(npu_inst_pe_1_0_4_sub_67_carry_5_), .B(
        npu_inst_pe_1_0_4_int_q_acc_5_), .ZN(npu_inst_pe_1_0_4_N70) );
  OR2_X1 npu_inst_pe_1_0_4_U119 ( .A1(npu_inst_pe_1_0_4_int_q_acc_5_), .A2(
        npu_inst_pe_1_0_4_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_0_4_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_0_4_U118 ( .A(npu_inst_pe_1_0_4_sub_67_carry_6_), .B(
        npu_inst_pe_1_0_4_int_q_acc_6_), .ZN(npu_inst_pe_1_0_4_N71) );
  OR2_X1 npu_inst_pe_1_0_4_U117 ( .A1(npu_inst_pe_1_0_4_int_q_acc_6_), .A2(
        npu_inst_pe_1_0_4_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_0_4_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_0_4_U116 ( .A(npu_inst_pe_1_0_4_int_q_acc_7_), .B(
        npu_inst_pe_1_0_4_sub_67_carry_7_), .ZN(npu_inst_pe_1_0_4_N72) );
  INV_X1 npu_inst_pe_1_0_4_U115 ( .A(npu_inst_n79), .ZN(npu_inst_pe_1_0_4_n6)
         );
  INV_X1 npu_inst_pe_1_0_4_U114 ( .A(npu_inst_n60), .ZN(npu_inst_pe_1_0_4_n3)
         );
  AOI22_X1 npu_inst_pe_1_0_4_U113 ( .A1(npu_inst_int_data_y_1__4__0_), .A2(
        npu_inst_pe_1_0_4_n58), .B1(npu_inst_pe_1_0_4_n118), .B2(
        npu_inst_pe_1_0_4_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_0_4_n57) );
  INV_X1 npu_inst_pe_1_0_4_U112 ( .A(npu_inst_pe_1_0_4_n57), .ZN(
        npu_inst_pe_1_0_4_n107) );
  AOI22_X1 npu_inst_pe_1_0_4_U111 ( .A1(npu_inst_int_data_y_1__4__0_), .A2(
        npu_inst_pe_1_0_4_n54), .B1(npu_inst_pe_1_0_4_n117), .B2(
        npu_inst_pe_1_0_4_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_0_4_n53) );
  INV_X1 npu_inst_pe_1_0_4_U110 ( .A(npu_inst_pe_1_0_4_n53), .ZN(
        npu_inst_pe_1_0_4_n108) );
  AOI22_X1 npu_inst_pe_1_0_4_U107 ( .A1(npu_inst_int_data_y_1__4__0_), .A2(
        npu_inst_pe_1_0_4_n50), .B1(npu_inst_pe_1_0_4_n116), .B2(
        npu_inst_pe_1_0_4_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_0_4_n49) );
  INV_X1 npu_inst_pe_1_0_4_U106 ( .A(npu_inst_pe_1_0_4_n49), .ZN(
        npu_inst_pe_1_0_4_n109) );
  AOI22_X1 npu_inst_pe_1_0_4_U105 ( .A1(npu_inst_int_data_y_1__4__0_), .A2(
        npu_inst_pe_1_0_4_n46), .B1(npu_inst_pe_1_0_4_n115), .B2(
        npu_inst_pe_1_0_4_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_0_4_n45) );
  INV_X1 npu_inst_pe_1_0_4_U104 ( .A(npu_inst_pe_1_0_4_n45), .ZN(
        npu_inst_pe_1_0_4_n110) );
  AOI22_X1 npu_inst_pe_1_0_4_U103 ( .A1(npu_inst_int_data_y_1__4__0_), .A2(
        npu_inst_pe_1_0_4_n42), .B1(npu_inst_pe_1_0_4_n114), .B2(
        npu_inst_pe_1_0_4_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_0_4_n41) );
  INV_X1 npu_inst_pe_1_0_4_U102 ( .A(npu_inst_pe_1_0_4_n41), .ZN(
        npu_inst_pe_1_0_4_n111) );
  AOI22_X1 npu_inst_pe_1_0_4_U101 ( .A1(npu_inst_int_data_y_1__4__1_), .A2(
        npu_inst_pe_1_0_4_n58), .B1(npu_inst_pe_1_0_4_n118), .B2(
        npu_inst_pe_1_0_4_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_0_4_n59) );
  INV_X1 npu_inst_pe_1_0_4_U100 ( .A(npu_inst_pe_1_0_4_n59), .ZN(
        npu_inst_pe_1_0_4_n101) );
  AOI22_X1 npu_inst_pe_1_0_4_U99 ( .A1(npu_inst_int_data_y_1__4__1_), .A2(
        npu_inst_pe_1_0_4_n54), .B1(npu_inst_pe_1_0_4_n117), .B2(
        npu_inst_pe_1_0_4_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_0_4_n55) );
  INV_X1 npu_inst_pe_1_0_4_U98 ( .A(npu_inst_pe_1_0_4_n55), .ZN(
        npu_inst_pe_1_0_4_n102) );
  AOI22_X1 npu_inst_pe_1_0_4_U97 ( .A1(npu_inst_int_data_y_1__4__1_), .A2(
        npu_inst_pe_1_0_4_n50), .B1(npu_inst_pe_1_0_4_n116), .B2(
        npu_inst_pe_1_0_4_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_0_4_n51) );
  INV_X1 npu_inst_pe_1_0_4_U96 ( .A(npu_inst_pe_1_0_4_n51), .ZN(
        npu_inst_pe_1_0_4_n103) );
  AOI22_X1 npu_inst_pe_1_0_4_U95 ( .A1(npu_inst_int_data_y_1__4__1_), .A2(
        npu_inst_pe_1_0_4_n46), .B1(npu_inst_pe_1_0_4_n115), .B2(
        npu_inst_pe_1_0_4_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_0_4_n47) );
  INV_X1 npu_inst_pe_1_0_4_U94 ( .A(npu_inst_pe_1_0_4_n47), .ZN(
        npu_inst_pe_1_0_4_n104) );
  AOI22_X1 npu_inst_pe_1_0_4_U93 ( .A1(npu_inst_int_data_y_1__4__1_), .A2(
        npu_inst_pe_1_0_4_n42), .B1(npu_inst_pe_1_0_4_n114), .B2(
        npu_inst_pe_1_0_4_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_0_4_n43) );
  INV_X1 npu_inst_pe_1_0_4_U92 ( .A(npu_inst_pe_1_0_4_n43), .ZN(
        npu_inst_pe_1_0_4_n105) );
  AOI22_X1 npu_inst_pe_1_0_4_U91 ( .A1(npu_inst_pe_1_0_4_n38), .A2(
        npu_inst_int_data_y_1__4__1_), .B1(npu_inst_pe_1_0_4_n113), .B2(
        npu_inst_pe_1_0_4_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_0_4_n39) );
  INV_X1 npu_inst_pe_1_0_4_U90 ( .A(npu_inst_pe_1_0_4_n39), .ZN(
        npu_inst_pe_1_0_4_n106) );
  AOI22_X1 npu_inst_pe_1_0_4_U89 ( .A1(npu_inst_pe_1_0_4_n38), .A2(
        npu_inst_int_data_y_1__4__0_), .B1(npu_inst_pe_1_0_4_n113), .B2(
        npu_inst_pe_1_0_4_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_0_4_n37) );
  INV_X1 npu_inst_pe_1_0_4_U88 ( .A(npu_inst_pe_1_0_4_n37), .ZN(
        npu_inst_pe_1_0_4_n112) );
  NOR3_X1 npu_inst_pe_1_0_4_U87 ( .A1(npu_inst_pe_1_0_4_n26), .A2(npu_inst_n60), .A3(npu_inst_int_ckg[59]), .ZN(npu_inst_pe_1_0_4_n85) );
  OR2_X1 npu_inst_pe_1_0_4_U86 ( .A1(npu_inst_pe_1_0_4_n85), .A2(
        npu_inst_pe_1_0_4_n2), .ZN(npu_inst_pe_1_0_4_N84) );
  NAND2_X1 npu_inst_pe_1_0_4_U85 ( .A1(npu_inst_pe_1_0_4_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_0_4_n60), .ZN(npu_inst_pe_1_0_4_n74) );
  OAI21_X1 npu_inst_pe_1_0_4_U84 ( .B1(npu_inst_pe_1_0_4_n63), .B2(
        npu_inst_pe_1_0_4_n60), .A(npu_inst_pe_1_0_4_n74), .ZN(
        npu_inst_pe_1_0_4_n97) );
  NAND2_X1 npu_inst_pe_1_0_4_U83 ( .A1(npu_inst_pe_1_0_4_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_0_4_n60), .ZN(npu_inst_pe_1_0_4_n73) );
  OAI21_X1 npu_inst_pe_1_0_4_U82 ( .B1(npu_inst_pe_1_0_4_n61), .B2(
        npu_inst_pe_1_0_4_n60), .A(npu_inst_pe_1_0_4_n73), .ZN(
        npu_inst_pe_1_0_4_n96) );
  NAND2_X1 npu_inst_pe_1_0_4_U81 ( .A1(npu_inst_pe_1_0_4_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_0_4_n56), .ZN(npu_inst_pe_1_0_4_n72) );
  OAI21_X1 npu_inst_pe_1_0_4_U80 ( .B1(npu_inst_pe_1_0_4_n63), .B2(
        npu_inst_pe_1_0_4_n56), .A(npu_inst_pe_1_0_4_n72), .ZN(
        npu_inst_pe_1_0_4_n95) );
  NAND2_X1 npu_inst_pe_1_0_4_U79 ( .A1(npu_inst_pe_1_0_4_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_0_4_n56), .ZN(npu_inst_pe_1_0_4_n71) );
  OAI21_X1 npu_inst_pe_1_0_4_U78 ( .B1(npu_inst_pe_1_0_4_n61), .B2(
        npu_inst_pe_1_0_4_n56), .A(npu_inst_pe_1_0_4_n71), .ZN(
        npu_inst_pe_1_0_4_n94) );
  NAND2_X1 npu_inst_pe_1_0_4_U77 ( .A1(npu_inst_pe_1_0_4_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_0_4_n52), .ZN(npu_inst_pe_1_0_4_n70) );
  OAI21_X1 npu_inst_pe_1_0_4_U76 ( .B1(npu_inst_pe_1_0_4_n63), .B2(
        npu_inst_pe_1_0_4_n52), .A(npu_inst_pe_1_0_4_n70), .ZN(
        npu_inst_pe_1_0_4_n93) );
  NAND2_X1 npu_inst_pe_1_0_4_U75 ( .A1(npu_inst_pe_1_0_4_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_0_4_n52), .ZN(npu_inst_pe_1_0_4_n69) );
  OAI21_X1 npu_inst_pe_1_0_4_U74 ( .B1(npu_inst_pe_1_0_4_n61), .B2(
        npu_inst_pe_1_0_4_n52), .A(npu_inst_pe_1_0_4_n69), .ZN(
        npu_inst_pe_1_0_4_n92) );
  NAND2_X1 npu_inst_pe_1_0_4_U73 ( .A1(npu_inst_pe_1_0_4_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_0_4_n48), .ZN(npu_inst_pe_1_0_4_n68) );
  OAI21_X1 npu_inst_pe_1_0_4_U72 ( .B1(npu_inst_pe_1_0_4_n63), .B2(
        npu_inst_pe_1_0_4_n48), .A(npu_inst_pe_1_0_4_n68), .ZN(
        npu_inst_pe_1_0_4_n91) );
  NAND2_X1 npu_inst_pe_1_0_4_U71 ( .A1(npu_inst_pe_1_0_4_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_0_4_n48), .ZN(npu_inst_pe_1_0_4_n67) );
  OAI21_X1 npu_inst_pe_1_0_4_U70 ( .B1(npu_inst_pe_1_0_4_n61), .B2(
        npu_inst_pe_1_0_4_n48), .A(npu_inst_pe_1_0_4_n67), .ZN(
        npu_inst_pe_1_0_4_n90) );
  NAND2_X1 npu_inst_pe_1_0_4_U69 ( .A1(npu_inst_pe_1_0_4_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_0_4_n44), .ZN(npu_inst_pe_1_0_4_n66) );
  OAI21_X1 npu_inst_pe_1_0_4_U68 ( .B1(npu_inst_pe_1_0_4_n63), .B2(
        npu_inst_pe_1_0_4_n44), .A(npu_inst_pe_1_0_4_n66), .ZN(
        npu_inst_pe_1_0_4_n89) );
  NAND2_X1 npu_inst_pe_1_0_4_U67 ( .A1(npu_inst_pe_1_0_4_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_0_4_n44), .ZN(npu_inst_pe_1_0_4_n65) );
  OAI21_X1 npu_inst_pe_1_0_4_U66 ( .B1(npu_inst_pe_1_0_4_n61), .B2(
        npu_inst_pe_1_0_4_n44), .A(npu_inst_pe_1_0_4_n65), .ZN(
        npu_inst_pe_1_0_4_n88) );
  NAND2_X1 npu_inst_pe_1_0_4_U65 ( .A1(npu_inst_pe_1_0_4_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_0_4_n40), .ZN(npu_inst_pe_1_0_4_n64) );
  OAI21_X1 npu_inst_pe_1_0_4_U64 ( .B1(npu_inst_pe_1_0_4_n63), .B2(
        npu_inst_pe_1_0_4_n40), .A(npu_inst_pe_1_0_4_n64), .ZN(
        npu_inst_pe_1_0_4_n87) );
  NAND2_X1 npu_inst_pe_1_0_4_U63 ( .A1(npu_inst_pe_1_0_4_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_0_4_n40), .ZN(npu_inst_pe_1_0_4_n62) );
  OAI21_X1 npu_inst_pe_1_0_4_U62 ( .B1(npu_inst_pe_1_0_4_n61), .B2(
        npu_inst_pe_1_0_4_n40), .A(npu_inst_pe_1_0_4_n62), .ZN(
        npu_inst_pe_1_0_4_n86) );
  AND2_X1 npu_inst_pe_1_0_4_U61 ( .A1(npu_inst_pe_1_0_4_int_q_acc_2_), .A2(
        npu_inst_pe_1_0_4_n1), .ZN(int_o_data_npu[26]) );
  AND2_X1 npu_inst_pe_1_0_4_U60 ( .A1(npu_inst_pe_1_0_4_int_q_acc_3_), .A2(
        npu_inst_pe_1_0_4_n2), .ZN(int_o_data_npu[27]) );
  AND2_X1 npu_inst_pe_1_0_4_U59 ( .A1(npu_inst_pe_1_0_4_int_q_acc_6_), .A2(
        npu_inst_pe_1_0_4_n2), .ZN(int_o_data_npu[30]) );
  AND2_X1 npu_inst_pe_1_0_4_U58 ( .A1(npu_inst_pe_1_0_4_int_q_acc_5_), .A2(
        npu_inst_pe_1_0_4_n2), .ZN(int_o_data_npu[29]) );
  AND2_X1 npu_inst_pe_1_0_4_U57 ( .A1(npu_inst_pe_1_0_4_int_q_acc_4_), .A2(
        npu_inst_pe_1_0_4_n2), .ZN(int_o_data_npu[28]) );
  AOI222_X1 npu_inst_pe_1_0_4_U56 ( .A1(npu_inst_int_data_res_1__4__0_), .A2(
        npu_inst_pe_1_0_4_n1), .B1(npu_inst_pe_1_0_4_N73), .B2(
        npu_inst_pe_1_0_4_n76), .C1(npu_inst_pe_1_0_4_N65), .C2(
        npu_inst_pe_1_0_4_n77), .ZN(npu_inst_pe_1_0_4_n84) );
  INV_X1 npu_inst_pe_1_0_4_U55 ( .A(npu_inst_pe_1_0_4_n84), .ZN(
        npu_inst_pe_1_0_4_n100) );
  AOI222_X1 npu_inst_pe_1_0_4_U54 ( .A1(npu_inst_int_data_res_1__4__7_), .A2(
        npu_inst_pe_1_0_4_n1), .B1(npu_inst_pe_1_0_4_N80), .B2(
        npu_inst_pe_1_0_4_n76), .C1(npu_inst_pe_1_0_4_N72), .C2(
        npu_inst_pe_1_0_4_n77), .ZN(npu_inst_pe_1_0_4_n75) );
  INV_X1 npu_inst_pe_1_0_4_U53 ( .A(npu_inst_pe_1_0_4_n75), .ZN(
        npu_inst_pe_1_0_4_n32) );
  AOI222_X1 npu_inst_pe_1_0_4_U52 ( .A1(npu_inst_int_data_res_1__4__1_), .A2(
        npu_inst_pe_1_0_4_n1), .B1(npu_inst_pe_1_0_4_N74), .B2(
        npu_inst_pe_1_0_4_n76), .C1(npu_inst_pe_1_0_4_N66), .C2(
        npu_inst_pe_1_0_4_n77), .ZN(npu_inst_pe_1_0_4_n83) );
  INV_X1 npu_inst_pe_1_0_4_U51 ( .A(npu_inst_pe_1_0_4_n83), .ZN(
        npu_inst_pe_1_0_4_n99) );
  AOI222_X1 npu_inst_pe_1_0_4_U50 ( .A1(npu_inst_int_data_res_1__4__2_), .A2(
        npu_inst_pe_1_0_4_n1), .B1(npu_inst_pe_1_0_4_N75), .B2(
        npu_inst_pe_1_0_4_n76), .C1(npu_inst_pe_1_0_4_N67), .C2(
        npu_inst_pe_1_0_4_n77), .ZN(npu_inst_pe_1_0_4_n82) );
  INV_X1 npu_inst_pe_1_0_4_U49 ( .A(npu_inst_pe_1_0_4_n82), .ZN(
        npu_inst_pe_1_0_4_n98) );
  AOI222_X1 npu_inst_pe_1_0_4_U48 ( .A1(npu_inst_int_data_res_1__4__3_), .A2(
        npu_inst_pe_1_0_4_n1), .B1(npu_inst_pe_1_0_4_N76), .B2(
        npu_inst_pe_1_0_4_n76), .C1(npu_inst_pe_1_0_4_N68), .C2(
        npu_inst_pe_1_0_4_n77), .ZN(npu_inst_pe_1_0_4_n81) );
  INV_X1 npu_inst_pe_1_0_4_U47 ( .A(npu_inst_pe_1_0_4_n81), .ZN(
        npu_inst_pe_1_0_4_n36) );
  AOI222_X1 npu_inst_pe_1_0_4_U46 ( .A1(npu_inst_int_data_res_1__4__4_), .A2(
        npu_inst_pe_1_0_4_n1), .B1(npu_inst_pe_1_0_4_N77), .B2(
        npu_inst_pe_1_0_4_n76), .C1(npu_inst_pe_1_0_4_N69), .C2(
        npu_inst_pe_1_0_4_n77), .ZN(npu_inst_pe_1_0_4_n80) );
  INV_X1 npu_inst_pe_1_0_4_U45 ( .A(npu_inst_pe_1_0_4_n80), .ZN(
        npu_inst_pe_1_0_4_n35) );
  AOI222_X1 npu_inst_pe_1_0_4_U44 ( .A1(npu_inst_int_data_res_1__4__5_), .A2(
        npu_inst_pe_1_0_4_n1), .B1(npu_inst_pe_1_0_4_N78), .B2(
        npu_inst_pe_1_0_4_n76), .C1(npu_inst_pe_1_0_4_N70), .C2(
        npu_inst_pe_1_0_4_n77), .ZN(npu_inst_pe_1_0_4_n79) );
  INV_X1 npu_inst_pe_1_0_4_U43 ( .A(npu_inst_pe_1_0_4_n79), .ZN(
        npu_inst_pe_1_0_4_n34) );
  AOI222_X1 npu_inst_pe_1_0_4_U42 ( .A1(npu_inst_int_data_res_1__4__6_), .A2(
        npu_inst_pe_1_0_4_n1), .B1(npu_inst_pe_1_0_4_N79), .B2(
        npu_inst_pe_1_0_4_n76), .C1(npu_inst_pe_1_0_4_N71), .C2(
        npu_inst_pe_1_0_4_n77), .ZN(npu_inst_pe_1_0_4_n78) );
  INV_X1 npu_inst_pe_1_0_4_U41 ( .A(npu_inst_pe_1_0_4_n78), .ZN(
        npu_inst_pe_1_0_4_n33) );
  INV_X1 npu_inst_pe_1_0_4_U40 ( .A(npu_inst_pe_1_0_4_int_data_1_), .ZN(
        npu_inst_pe_1_0_4_n13) );
  AND2_X1 npu_inst_pe_1_0_4_U39 ( .A1(npu_inst_int_data_x_0__4__1_), .A2(
        npu_inst_pe_1_0_4_int_q_weight_1_), .ZN(npu_inst_pe_1_0_4_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_0_4_U38 ( .A1(npu_inst_int_data_x_0__4__0_), .A2(
        npu_inst_pe_1_0_4_int_q_weight_1_), .ZN(npu_inst_pe_1_0_4_int_data_0_)
         );
  AND2_X1 npu_inst_pe_1_0_4_U37 ( .A1(npu_inst_pe_1_0_4_n2), .A2(
        npu_inst_pe_1_0_4_int_q_acc_7_), .ZN(int_o_data_npu[31]) );
  AND2_X1 npu_inst_pe_1_0_4_U36 ( .A1(npu_inst_pe_1_0_4_int_q_acc_1_), .A2(
        npu_inst_pe_1_0_4_n1), .ZN(int_o_data_npu[25]) );
  AND2_X1 npu_inst_pe_1_0_4_U35 ( .A1(npu_inst_pe_1_0_4_int_q_acc_0_), .A2(
        npu_inst_pe_1_0_4_n1), .ZN(int_o_data_npu[24]) );
  AND2_X1 npu_inst_pe_1_0_4_U34 ( .A1(npu_inst_pe_1_0_4_N93), .A2(npu_inst_n60), .ZN(npu_inst_pe_1_0_4_o_data_v_0_) );
  AND2_X1 npu_inst_pe_1_0_4_U33 ( .A1(npu_inst_n60), .A2(npu_inst_pe_1_0_4_N94), .ZN(npu_inst_pe_1_0_4_o_data_v_1_) );
  AOI22_X1 npu_inst_pe_1_0_4_U32 ( .A1(npu_inst_n60), .A2(
        npu_inst_int_data_y_1__4__1_), .B1(npu_inst_pe_1_0_4_n3), .B2(
        npu_inst_int_data_x_0__5__1_), .ZN(npu_inst_pe_1_0_4_n63) );
  AOI22_X1 npu_inst_pe_1_0_4_U31 ( .A1(npu_inst_n60), .A2(
        npu_inst_int_data_y_1__4__0_), .B1(npu_inst_pe_1_0_4_n3), .B2(
        npu_inst_int_data_x_0__5__0_), .ZN(npu_inst_pe_1_0_4_n61) );
  INV_X1 npu_inst_pe_1_0_4_U30 ( .A(npu_inst_pe_1_0_4_int_data_0_), .ZN(
        npu_inst_pe_1_0_4_n12) );
  INV_X1 npu_inst_pe_1_0_4_U29 ( .A(npu_inst_n71), .ZN(npu_inst_pe_1_0_4_n5)
         );
  OR3_X1 npu_inst_pe_1_0_4_U28 ( .A1(npu_inst_n79), .A2(npu_inst_pe_1_0_4_n7), 
        .A3(npu_inst_pe_1_0_4_n5), .ZN(npu_inst_pe_1_0_4_n56) );
  OR3_X1 npu_inst_pe_1_0_4_U27 ( .A1(npu_inst_pe_1_0_4_n5), .A2(
        npu_inst_pe_1_0_4_n7), .A3(npu_inst_pe_1_0_4_n6), .ZN(
        npu_inst_pe_1_0_4_n48) );
  INV_X1 npu_inst_pe_1_0_4_U26 ( .A(npu_inst_pe_1_0_4_n5), .ZN(
        npu_inst_pe_1_0_4_n4) );
  OR3_X1 npu_inst_pe_1_0_4_U25 ( .A1(npu_inst_pe_1_0_4_n4), .A2(
        npu_inst_pe_1_0_4_n7), .A3(npu_inst_pe_1_0_4_n6), .ZN(
        npu_inst_pe_1_0_4_n52) );
  OR3_X1 npu_inst_pe_1_0_4_U24 ( .A1(npu_inst_n79), .A2(npu_inst_pe_1_0_4_n7), 
        .A3(npu_inst_pe_1_0_4_n4), .ZN(npu_inst_pe_1_0_4_n60) );
  NOR2_X1 npu_inst_pe_1_0_4_U23 ( .A1(npu_inst_pe_1_0_4_n60), .A2(
        npu_inst_pe_1_0_4_n3), .ZN(npu_inst_pe_1_0_4_n58) );
  NOR2_X1 npu_inst_pe_1_0_4_U22 ( .A1(npu_inst_pe_1_0_4_n56), .A2(
        npu_inst_pe_1_0_4_n3), .ZN(npu_inst_pe_1_0_4_n54) );
  NOR2_X1 npu_inst_pe_1_0_4_U21 ( .A1(npu_inst_pe_1_0_4_n52), .A2(
        npu_inst_pe_1_0_4_n3), .ZN(npu_inst_pe_1_0_4_n50) );
  NOR2_X1 npu_inst_pe_1_0_4_U20 ( .A1(npu_inst_pe_1_0_4_n48), .A2(
        npu_inst_pe_1_0_4_n3), .ZN(npu_inst_pe_1_0_4_n46) );
  NOR2_X1 npu_inst_pe_1_0_4_U19 ( .A1(npu_inst_pe_1_0_4_n40), .A2(
        npu_inst_pe_1_0_4_n3), .ZN(npu_inst_pe_1_0_4_n38) );
  NOR2_X1 npu_inst_pe_1_0_4_U18 ( .A1(npu_inst_pe_1_0_4_n44), .A2(
        npu_inst_pe_1_0_4_n3), .ZN(npu_inst_pe_1_0_4_n42) );
  BUF_X1 npu_inst_pe_1_0_4_U17 ( .A(npu_inst_n106), .Z(npu_inst_pe_1_0_4_n7)
         );
  INV_X1 npu_inst_pe_1_0_4_U16 ( .A(npu_inst_n126), .ZN(npu_inst_pe_1_0_4_n11)
         );
  INV_X1 npu_inst_pe_1_0_4_U15 ( .A(npu_inst_pe_1_0_4_n38), .ZN(
        npu_inst_pe_1_0_4_n113) );
  INV_X1 npu_inst_pe_1_0_4_U14 ( .A(npu_inst_pe_1_0_4_n58), .ZN(
        npu_inst_pe_1_0_4_n118) );
  INV_X1 npu_inst_pe_1_0_4_U13 ( .A(npu_inst_pe_1_0_4_n54), .ZN(
        npu_inst_pe_1_0_4_n117) );
  INV_X1 npu_inst_pe_1_0_4_U12 ( .A(npu_inst_pe_1_0_4_n50), .ZN(
        npu_inst_pe_1_0_4_n116) );
  INV_X1 npu_inst_pe_1_0_4_U11 ( .A(npu_inst_pe_1_0_4_n46), .ZN(
        npu_inst_pe_1_0_4_n115) );
  INV_X1 npu_inst_pe_1_0_4_U10 ( .A(npu_inst_pe_1_0_4_n42), .ZN(
        npu_inst_pe_1_0_4_n114) );
  BUF_X1 npu_inst_pe_1_0_4_U9 ( .A(npu_inst_n36), .Z(npu_inst_pe_1_0_4_n2) );
  BUF_X1 npu_inst_pe_1_0_4_U8 ( .A(npu_inst_n36), .Z(npu_inst_pe_1_0_4_n1) );
  BUF_X1 npu_inst_pe_1_0_4_U7 ( .A(npu_inst_pe_1_0_4_n11), .Z(
        npu_inst_pe_1_0_4_n10) );
  BUF_X1 npu_inst_pe_1_0_4_U6 ( .A(npu_inst_pe_1_0_4_n11), .Z(
        npu_inst_pe_1_0_4_n9) );
  BUF_X1 npu_inst_pe_1_0_4_U5 ( .A(npu_inst_pe_1_0_4_n11), .Z(
        npu_inst_pe_1_0_4_n8) );
  NOR2_X1 npu_inst_pe_1_0_4_U4 ( .A1(npu_inst_pe_1_0_4_int_q_weight_0_), .A2(
        npu_inst_pe_1_0_4_n1), .ZN(npu_inst_pe_1_0_4_n76) );
  NOR2_X1 npu_inst_pe_1_0_4_U3 ( .A1(npu_inst_pe_1_0_4_n27), .A2(
        npu_inst_pe_1_0_4_n1), .ZN(npu_inst_pe_1_0_4_n77) );
  FA_X1 npu_inst_pe_1_0_4_sub_67_U2_1 ( .A(npu_inst_pe_1_0_4_int_q_acc_1_), 
        .B(npu_inst_pe_1_0_4_n13), .CI(npu_inst_pe_1_0_4_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_0_4_sub_67_carry_2_), .S(npu_inst_pe_1_0_4_N66) );
  FA_X1 npu_inst_pe_1_0_4_add_69_U1_1 ( .A(npu_inst_pe_1_0_4_int_q_acc_1_), 
        .B(npu_inst_pe_1_0_4_int_data_1_), .CI(
        npu_inst_pe_1_0_4_add_69_carry_1_), .CO(
        npu_inst_pe_1_0_4_add_69_carry_2_), .S(npu_inst_pe_1_0_4_N74) );
  NAND3_X1 npu_inst_pe_1_0_4_U109 ( .A1(npu_inst_pe_1_0_4_n5), .A2(
        npu_inst_pe_1_0_4_n6), .A3(npu_inst_pe_1_0_4_n7), .ZN(
        npu_inst_pe_1_0_4_n44) );
  NAND3_X1 npu_inst_pe_1_0_4_U108 ( .A1(npu_inst_pe_1_0_4_n4), .A2(
        npu_inst_pe_1_0_4_n6), .A3(npu_inst_pe_1_0_4_n7), .ZN(
        npu_inst_pe_1_0_4_n40) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_0_4_n33), .CK(
        npu_inst_pe_1_0_4_net4470), .RN(npu_inst_pe_1_0_4_n8), .Q(
        npu_inst_pe_1_0_4_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_0_4_n34), .CK(
        npu_inst_pe_1_0_4_net4470), .RN(npu_inst_pe_1_0_4_n8), .Q(
        npu_inst_pe_1_0_4_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_0_4_n35), .CK(
        npu_inst_pe_1_0_4_net4470), .RN(npu_inst_pe_1_0_4_n8), .Q(
        npu_inst_pe_1_0_4_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_0_4_n36), .CK(
        npu_inst_pe_1_0_4_net4470), .RN(npu_inst_pe_1_0_4_n8), .Q(
        npu_inst_pe_1_0_4_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_0_4_n98), .CK(
        npu_inst_pe_1_0_4_net4470), .RN(npu_inst_pe_1_0_4_n8), .Q(
        npu_inst_pe_1_0_4_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_0_4_n99), .CK(
        npu_inst_pe_1_0_4_net4470), .RN(npu_inst_pe_1_0_4_n8), .Q(
        npu_inst_pe_1_0_4_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_0_4_n32), .CK(
        npu_inst_pe_1_0_4_net4470), .RN(npu_inst_pe_1_0_4_n8), .Q(
        npu_inst_pe_1_0_4_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_0_4_n100), 
        .CK(npu_inst_pe_1_0_4_net4470), .RN(npu_inst_pe_1_0_4_n8), .Q(
        npu_inst_pe_1_0_4_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_weight_reg_0_ ( .D(npu_inst_n112), .CK(
        npu_inst_pe_1_0_4_net4476), .RN(npu_inst_pe_1_0_4_n8), .Q(
        npu_inst_pe_1_0_4_int_q_weight_0_), .QN(npu_inst_pe_1_0_4_n27) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_weight_reg_1_ ( .D(npu_inst_n118), .CK(
        npu_inst_pe_1_0_4_net4476), .RN(npu_inst_pe_1_0_4_n8), .Q(
        npu_inst_pe_1_0_4_int_q_weight_1_), .QN(npu_inst_pe_1_0_4_n26) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_0_4_n112), 
        .CK(npu_inst_pe_1_0_4_net4476), .RN(npu_inst_pe_1_0_4_n8), .Q(
        npu_inst_pe_1_0_4_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_0_4_n106), 
        .CK(npu_inst_pe_1_0_4_net4476), .RN(npu_inst_pe_1_0_4_n8), .Q(
        npu_inst_pe_1_0_4_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_0_4_n111), 
        .CK(npu_inst_pe_1_0_4_net4476), .RN(npu_inst_pe_1_0_4_n9), .Q(
        npu_inst_pe_1_0_4_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_0_4_n105), 
        .CK(npu_inst_pe_1_0_4_net4476), .RN(npu_inst_pe_1_0_4_n9), .Q(
        npu_inst_pe_1_0_4_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_0_4_n110), 
        .CK(npu_inst_pe_1_0_4_net4476), .RN(npu_inst_pe_1_0_4_n9), .Q(
        npu_inst_pe_1_0_4_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_0_4_n104), 
        .CK(npu_inst_pe_1_0_4_net4476), .RN(npu_inst_pe_1_0_4_n9), .Q(
        npu_inst_pe_1_0_4_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_0_4_n109), 
        .CK(npu_inst_pe_1_0_4_net4476), .RN(npu_inst_pe_1_0_4_n9), .Q(
        npu_inst_pe_1_0_4_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_0_4_n103), 
        .CK(npu_inst_pe_1_0_4_net4476), .RN(npu_inst_pe_1_0_4_n9), .Q(
        npu_inst_pe_1_0_4_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_0_4_n108), 
        .CK(npu_inst_pe_1_0_4_net4476), .RN(npu_inst_pe_1_0_4_n9), .Q(
        npu_inst_pe_1_0_4_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_0_4_n102), 
        .CK(npu_inst_pe_1_0_4_net4476), .RN(npu_inst_pe_1_0_4_n9), .Q(
        npu_inst_pe_1_0_4_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_0_4_n107), 
        .CK(npu_inst_pe_1_0_4_net4476), .RN(npu_inst_pe_1_0_4_n9), .Q(
        npu_inst_pe_1_0_4_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_0_4_n101), 
        .CK(npu_inst_pe_1_0_4_net4476), .RN(npu_inst_pe_1_0_4_n9), .Q(
        npu_inst_pe_1_0_4_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_0_4_n86), 
        .CK(npu_inst_pe_1_0_4_net4476), .RN(npu_inst_pe_1_0_4_n9), .Q(
        npu_inst_pe_1_0_4_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_0_4_n87), 
        .CK(npu_inst_pe_1_0_4_net4476), .RN(npu_inst_pe_1_0_4_n9), .Q(
        npu_inst_pe_1_0_4_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_0_4_n88), 
        .CK(npu_inst_pe_1_0_4_net4476), .RN(npu_inst_pe_1_0_4_n10), .Q(
        npu_inst_pe_1_0_4_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_0_4_n89), 
        .CK(npu_inst_pe_1_0_4_net4476), .RN(npu_inst_pe_1_0_4_n10), .Q(
        npu_inst_pe_1_0_4_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_0_4_n90), 
        .CK(npu_inst_pe_1_0_4_net4476), .RN(npu_inst_pe_1_0_4_n10), .Q(
        npu_inst_pe_1_0_4_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_0_4_n91), 
        .CK(npu_inst_pe_1_0_4_net4476), .RN(npu_inst_pe_1_0_4_n10), .Q(
        npu_inst_pe_1_0_4_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_0_4_n92), 
        .CK(npu_inst_pe_1_0_4_net4476), .RN(npu_inst_pe_1_0_4_n10), .Q(
        npu_inst_pe_1_0_4_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_0_4_n93), 
        .CK(npu_inst_pe_1_0_4_net4476), .RN(npu_inst_pe_1_0_4_n10), .Q(
        npu_inst_pe_1_0_4_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_0_4_n94), 
        .CK(npu_inst_pe_1_0_4_net4476), .RN(npu_inst_pe_1_0_4_n10), .Q(
        npu_inst_pe_1_0_4_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_0_4_n95), 
        .CK(npu_inst_pe_1_0_4_net4476), .RN(npu_inst_pe_1_0_4_n10), .Q(
        npu_inst_pe_1_0_4_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_0_4_n96), 
        .CK(npu_inst_pe_1_0_4_net4476), .RN(npu_inst_pe_1_0_4_n10), .Q(
        npu_inst_pe_1_0_4_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_0_4_n97), 
        .CK(npu_inst_pe_1_0_4_net4476), .RN(npu_inst_pe_1_0_4_n10), .Q(
        npu_inst_pe_1_0_4_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_0_4_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_0_4_N84), .SE(1'b0), .GCK(npu_inst_pe_1_0_4_net4470) );
  CLKGATETST_X1 npu_inst_pe_1_0_4_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n66), .SE(1'b0), .GCK(npu_inst_pe_1_0_4_net4476) );
  MUX2_X1 npu_inst_pe_1_0_5_U162 ( .A(npu_inst_pe_1_0_5_n32), .B(
        npu_inst_pe_1_0_5_n29), .S(npu_inst_pe_1_0_5_n8), .Z(
        npu_inst_pe_1_0_5_N93) );
  MUX2_X1 npu_inst_pe_1_0_5_U161 ( .A(npu_inst_pe_1_0_5_n31), .B(
        npu_inst_pe_1_0_5_n30), .S(npu_inst_pe_1_0_5_n6), .Z(
        npu_inst_pe_1_0_5_n32) );
  MUX2_X1 npu_inst_pe_1_0_5_U160 ( .A(npu_inst_pe_1_0_5_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_0_5_int_q_reg_v_1__0_), .S(npu_inst_pe_1_0_5_n4), .Z(
        npu_inst_pe_1_0_5_n31) );
  MUX2_X1 npu_inst_pe_1_0_5_U159 ( .A(npu_inst_pe_1_0_5_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_0_5_int_q_reg_v_3__0_), .S(npu_inst_pe_1_0_5_n4), .Z(
        npu_inst_pe_1_0_5_n30) );
  MUX2_X1 npu_inst_pe_1_0_5_U158 ( .A(npu_inst_pe_1_0_5_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_0_5_int_q_reg_v_5__0_), .S(npu_inst_pe_1_0_5_n4), .Z(
        npu_inst_pe_1_0_5_n29) );
  MUX2_X1 npu_inst_pe_1_0_5_U157 ( .A(npu_inst_pe_1_0_5_n28), .B(
        npu_inst_pe_1_0_5_n23), .S(npu_inst_pe_1_0_5_n8), .Z(
        npu_inst_pe_1_0_5_N94) );
  MUX2_X1 npu_inst_pe_1_0_5_U156 ( .A(npu_inst_pe_1_0_5_n25), .B(
        npu_inst_pe_1_0_5_n24), .S(npu_inst_pe_1_0_5_n6), .Z(
        npu_inst_pe_1_0_5_n28) );
  MUX2_X1 npu_inst_pe_1_0_5_U155 ( .A(npu_inst_pe_1_0_5_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_0_5_int_q_reg_v_1__1_), .S(npu_inst_pe_1_0_5_n4), .Z(
        npu_inst_pe_1_0_5_n25) );
  MUX2_X1 npu_inst_pe_1_0_5_U154 ( .A(npu_inst_pe_1_0_5_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_0_5_int_q_reg_v_3__1_), .S(npu_inst_pe_1_0_5_n4), .Z(
        npu_inst_pe_1_0_5_n24) );
  MUX2_X1 npu_inst_pe_1_0_5_U153 ( .A(npu_inst_pe_1_0_5_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_0_5_int_q_reg_v_5__1_), .S(npu_inst_pe_1_0_5_n4), .Z(
        npu_inst_pe_1_0_5_n23) );
  MUX2_X1 npu_inst_pe_1_0_5_U152 ( .A(npu_inst_pe_1_0_5_n22), .B(
        npu_inst_pe_1_0_5_n19), .S(npu_inst_pe_1_0_5_n8), .Z(
        npu_inst_int_data_x_0__5__1_) );
  MUX2_X1 npu_inst_pe_1_0_5_U151 ( .A(npu_inst_pe_1_0_5_n21), .B(
        npu_inst_pe_1_0_5_n20), .S(npu_inst_pe_1_0_5_n6), .Z(
        npu_inst_pe_1_0_5_n22) );
  MUX2_X1 npu_inst_pe_1_0_5_U150 ( .A(npu_inst_pe_1_0_5_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_0_5_int_q_reg_h_1__1_), .S(npu_inst_pe_1_0_5_n4), .Z(
        npu_inst_pe_1_0_5_n21) );
  MUX2_X1 npu_inst_pe_1_0_5_U149 ( .A(npu_inst_pe_1_0_5_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_0_5_int_q_reg_h_3__1_), .S(npu_inst_pe_1_0_5_n4), .Z(
        npu_inst_pe_1_0_5_n20) );
  MUX2_X1 npu_inst_pe_1_0_5_U148 ( .A(npu_inst_pe_1_0_5_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_0_5_int_q_reg_h_5__1_), .S(npu_inst_pe_1_0_5_n4), .Z(
        npu_inst_pe_1_0_5_n19) );
  MUX2_X1 npu_inst_pe_1_0_5_U147 ( .A(npu_inst_pe_1_0_5_n18), .B(
        npu_inst_pe_1_0_5_n15), .S(npu_inst_pe_1_0_5_n8), .Z(
        npu_inst_int_data_x_0__5__0_) );
  MUX2_X1 npu_inst_pe_1_0_5_U146 ( .A(npu_inst_pe_1_0_5_n17), .B(
        npu_inst_pe_1_0_5_n16), .S(npu_inst_pe_1_0_5_n6), .Z(
        npu_inst_pe_1_0_5_n18) );
  MUX2_X1 npu_inst_pe_1_0_5_U145 ( .A(npu_inst_pe_1_0_5_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_0_5_int_q_reg_h_1__0_), .S(npu_inst_pe_1_0_5_n4), .Z(
        npu_inst_pe_1_0_5_n17) );
  MUX2_X1 npu_inst_pe_1_0_5_U144 ( .A(npu_inst_pe_1_0_5_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_0_5_int_q_reg_h_3__0_), .S(npu_inst_pe_1_0_5_n4), .Z(
        npu_inst_pe_1_0_5_n16) );
  MUX2_X1 npu_inst_pe_1_0_5_U143 ( .A(npu_inst_pe_1_0_5_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_0_5_int_q_reg_h_5__0_), .S(npu_inst_pe_1_0_5_n4), .Z(
        npu_inst_pe_1_0_5_n15) );
  XOR2_X1 npu_inst_pe_1_0_5_U142 ( .A(npu_inst_pe_1_0_5_int_data_0_), .B(
        npu_inst_pe_1_0_5_int_q_acc_0_), .Z(npu_inst_pe_1_0_5_N73) );
  AND2_X1 npu_inst_pe_1_0_5_U141 ( .A1(npu_inst_pe_1_0_5_int_q_acc_0_), .A2(
        npu_inst_pe_1_0_5_int_data_0_), .ZN(npu_inst_pe_1_0_5_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_0_5_U140 ( .A(npu_inst_pe_1_0_5_int_q_acc_0_), .B(
        npu_inst_pe_1_0_5_n13), .ZN(npu_inst_pe_1_0_5_N65) );
  OR2_X1 npu_inst_pe_1_0_5_U139 ( .A1(npu_inst_pe_1_0_5_n13), .A2(
        npu_inst_pe_1_0_5_int_q_acc_0_), .ZN(npu_inst_pe_1_0_5_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_0_5_U138 ( .A(npu_inst_pe_1_0_5_int_q_acc_2_), .B(
        npu_inst_pe_1_0_5_add_69_carry_2_), .Z(npu_inst_pe_1_0_5_N75) );
  AND2_X1 npu_inst_pe_1_0_5_U137 ( .A1(npu_inst_pe_1_0_5_add_69_carry_2_), 
        .A2(npu_inst_pe_1_0_5_int_q_acc_2_), .ZN(
        npu_inst_pe_1_0_5_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_0_5_U136 ( .A(npu_inst_pe_1_0_5_int_q_acc_3_), .B(
        npu_inst_pe_1_0_5_add_69_carry_3_), .Z(npu_inst_pe_1_0_5_N76) );
  AND2_X1 npu_inst_pe_1_0_5_U135 ( .A1(npu_inst_pe_1_0_5_add_69_carry_3_), 
        .A2(npu_inst_pe_1_0_5_int_q_acc_3_), .ZN(
        npu_inst_pe_1_0_5_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_0_5_U134 ( .A(npu_inst_pe_1_0_5_int_q_acc_4_), .B(
        npu_inst_pe_1_0_5_add_69_carry_4_), .Z(npu_inst_pe_1_0_5_N77) );
  AND2_X1 npu_inst_pe_1_0_5_U133 ( .A1(npu_inst_pe_1_0_5_add_69_carry_4_), 
        .A2(npu_inst_pe_1_0_5_int_q_acc_4_), .ZN(
        npu_inst_pe_1_0_5_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_0_5_U132 ( .A(npu_inst_pe_1_0_5_int_q_acc_5_), .B(
        npu_inst_pe_1_0_5_add_69_carry_5_), .Z(npu_inst_pe_1_0_5_N78) );
  AND2_X1 npu_inst_pe_1_0_5_U131 ( .A1(npu_inst_pe_1_0_5_add_69_carry_5_), 
        .A2(npu_inst_pe_1_0_5_int_q_acc_5_), .ZN(
        npu_inst_pe_1_0_5_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_0_5_U130 ( .A(npu_inst_pe_1_0_5_int_q_acc_6_), .B(
        npu_inst_pe_1_0_5_add_69_carry_6_), .Z(npu_inst_pe_1_0_5_N79) );
  AND2_X1 npu_inst_pe_1_0_5_U129 ( .A1(npu_inst_pe_1_0_5_add_69_carry_6_), 
        .A2(npu_inst_pe_1_0_5_int_q_acc_6_), .ZN(
        npu_inst_pe_1_0_5_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_0_5_U128 ( .A(npu_inst_pe_1_0_5_int_q_acc_7_), .B(
        npu_inst_pe_1_0_5_add_69_carry_7_), .Z(npu_inst_pe_1_0_5_N80) );
  XNOR2_X1 npu_inst_pe_1_0_5_U127 ( .A(npu_inst_pe_1_0_5_sub_67_carry_2_), .B(
        npu_inst_pe_1_0_5_int_q_acc_2_), .ZN(npu_inst_pe_1_0_5_N67) );
  OR2_X1 npu_inst_pe_1_0_5_U126 ( .A1(npu_inst_pe_1_0_5_int_q_acc_2_), .A2(
        npu_inst_pe_1_0_5_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_0_5_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_0_5_U125 ( .A(npu_inst_pe_1_0_5_sub_67_carry_3_), .B(
        npu_inst_pe_1_0_5_int_q_acc_3_), .ZN(npu_inst_pe_1_0_5_N68) );
  OR2_X1 npu_inst_pe_1_0_5_U124 ( .A1(npu_inst_pe_1_0_5_int_q_acc_3_), .A2(
        npu_inst_pe_1_0_5_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_0_5_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_0_5_U123 ( .A(npu_inst_pe_1_0_5_sub_67_carry_4_), .B(
        npu_inst_pe_1_0_5_int_q_acc_4_), .ZN(npu_inst_pe_1_0_5_N69) );
  OR2_X1 npu_inst_pe_1_0_5_U122 ( .A1(npu_inst_pe_1_0_5_int_q_acc_4_), .A2(
        npu_inst_pe_1_0_5_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_0_5_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_0_5_U121 ( .A(npu_inst_pe_1_0_5_sub_67_carry_5_), .B(
        npu_inst_pe_1_0_5_int_q_acc_5_), .ZN(npu_inst_pe_1_0_5_N70) );
  OR2_X1 npu_inst_pe_1_0_5_U120 ( .A1(npu_inst_pe_1_0_5_int_q_acc_5_), .A2(
        npu_inst_pe_1_0_5_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_0_5_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_0_5_U119 ( .A(npu_inst_pe_1_0_5_sub_67_carry_6_), .B(
        npu_inst_pe_1_0_5_int_q_acc_6_), .ZN(npu_inst_pe_1_0_5_N71) );
  OR2_X1 npu_inst_pe_1_0_5_U118 ( .A1(npu_inst_pe_1_0_5_int_q_acc_6_), .A2(
        npu_inst_pe_1_0_5_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_0_5_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_0_5_U117 ( .A(npu_inst_pe_1_0_5_int_q_acc_7_), .B(
        npu_inst_pe_1_0_5_sub_67_carry_7_), .ZN(npu_inst_pe_1_0_5_N72) );
  INV_X1 npu_inst_pe_1_0_5_U116 ( .A(npu_inst_n79), .ZN(npu_inst_pe_1_0_5_n7)
         );
  INV_X1 npu_inst_pe_1_0_5_U115 ( .A(npu_inst_pe_1_0_5_n7), .ZN(
        npu_inst_pe_1_0_5_n6) );
  INV_X1 npu_inst_pe_1_0_5_U114 ( .A(npu_inst_n60), .ZN(npu_inst_pe_1_0_5_n3)
         );
  AOI22_X1 npu_inst_pe_1_0_5_U113 ( .A1(npu_inst_int_data_y_1__5__0_), .A2(
        npu_inst_pe_1_0_5_n58), .B1(npu_inst_pe_1_0_5_n119), .B2(
        npu_inst_pe_1_0_5_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_0_5_n57) );
  INV_X1 npu_inst_pe_1_0_5_U112 ( .A(npu_inst_pe_1_0_5_n57), .ZN(
        npu_inst_pe_1_0_5_n108) );
  AOI22_X1 npu_inst_pe_1_0_5_U111 ( .A1(npu_inst_int_data_y_1__5__0_), .A2(
        npu_inst_pe_1_0_5_n54), .B1(npu_inst_pe_1_0_5_n118), .B2(
        npu_inst_pe_1_0_5_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_0_5_n53) );
  INV_X1 npu_inst_pe_1_0_5_U110 ( .A(npu_inst_pe_1_0_5_n53), .ZN(
        npu_inst_pe_1_0_5_n109) );
  AOI22_X1 npu_inst_pe_1_0_5_U107 ( .A1(npu_inst_int_data_y_1__5__0_), .A2(
        npu_inst_pe_1_0_5_n50), .B1(npu_inst_pe_1_0_5_n117), .B2(
        npu_inst_pe_1_0_5_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_0_5_n49) );
  INV_X1 npu_inst_pe_1_0_5_U106 ( .A(npu_inst_pe_1_0_5_n49), .ZN(
        npu_inst_pe_1_0_5_n110) );
  AOI22_X1 npu_inst_pe_1_0_5_U105 ( .A1(npu_inst_int_data_y_1__5__0_), .A2(
        npu_inst_pe_1_0_5_n46), .B1(npu_inst_pe_1_0_5_n116), .B2(
        npu_inst_pe_1_0_5_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_0_5_n45) );
  INV_X1 npu_inst_pe_1_0_5_U104 ( .A(npu_inst_pe_1_0_5_n45), .ZN(
        npu_inst_pe_1_0_5_n111) );
  AOI22_X1 npu_inst_pe_1_0_5_U103 ( .A1(npu_inst_int_data_y_1__5__0_), .A2(
        npu_inst_pe_1_0_5_n42), .B1(npu_inst_pe_1_0_5_n115), .B2(
        npu_inst_pe_1_0_5_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_0_5_n41) );
  INV_X1 npu_inst_pe_1_0_5_U102 ( .A(npu_inst_pe_1_0_5_n41), .ZN(
        npu_inst_pe_1_0_5_n112) );
  AOI22_X1 npu_inst_pe_1_0_5_U101 ( .A1(npu_inst_int_data_y_1__5__1_), .A2(
        npu_inst_pe_1_0_5_n58), .B1(npu_inst_pe_1_0_5_n119), .B2(
        npu_inst_pe_1_0_5_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_0_5_n59) );
  INV_X1 npu_inst_pe_1_0_5_U100 ( .A(npu_inst_pe_1_0_5_n59), .ZN(
        npu_inst_pe_1_0_5_n102) );
  AOI22_X1 npu_inst_pe_1_0_5_U99 ( .A1(npu_inst_int_data_y_1__5__1_), .A2(
        npu_inst_pe_1_0_5_n54), .B1(npu_inst_pe_1_0_5_n118), .B2(
        npu_inst_pe_1_0_5_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_0_5_n55) );
  INV_X1 npu_inst_pe_1_0_5_U98 ( .A(npu_inst_pe_1_0_5_n55), .ZN(
        npu_inst_pe_1_0_5_n103) );
  AOI22_X1 npu_inst_pe_1_0_5_U97 ( .A1(npu_inst_int_data_y_1__5__1_), .A2(
        npu_inst_pe_1_0_5_n50), .B1(npu_inst_pe_1_0_5_n117), .B2(
        npu_inst_pe_1_0_5_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_0_5_n51) );
  INV_X1 npu_inst_pe_1_0_5_U96 ( .A(npu_inst_pe_1_0_5_n51), .ZN(
        npu_inst_pe_1_0_5_n104) );
  AOI22_X1 npu_inst_pe_1_0_5_U95 ( .A1(npu_inst_int_data_y_1__5__1_), .A2(
        npu_inst_pe_1_0_5_n46), .B1(npu_inst_pe_1_0_5_n116), .B2(
        npu_inst_pe_1_0_5_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_0_5_n47) );
  INV_X1 npu_inst_pe_1_0_5_U94 ( .A(npu_inst_pe_1_0_5_n47), .ZN(
        npu_inst_pe_1_0_5_n105) );
  AOI22_X1 npu_inst_pe_1_0_5_U93 ( .A1(npu_inst_int_data_y_1__5__1_), .A2(
        npu_inst_pe_1_0_5_n42), .B1(npu_inst_pe_1_0_5_n115), .B2(
        npu_inst_pe_1_0_5_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_0_5_n43) );
  INV_X1 npu_inst_pe_1_0_5_U92 ( .A(npu_inst_pe_1_0_5_n43), .ZN(
        npu_inst_pe_1_0_5_n106) );
  AOI22_X1 npu_inst_pe_1_0_5_U91 ( .A1(npu_inst_pe_1_0_5_n38), .A2(
        npu_inst_int_data_y_1__5__1_), .B1(npu_inst_pe_1_0_5_n114), .B2(
        npu_inst_pe_1_0_5_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_0_5_n39) );
  INV_X1 npu_inst_pe_1_0_5_U90 ( .A(npu_inst_pe_1_0_5_n39), .ZN(
        npu_inst_pe_1_0_5_n107) );
  AOI22_X1 npu_inst_pe_1_0_5_U89 ( .A1(npu_inst_pe_1_0_5_n38), .A2(
        npu_inst_int_data_y_1__5__0_), .B1(npu_inst_pe_1_0_5_n114), .B2(
        npu_inst_pe_1_0_5_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_0_5_n37) );
  INV_X1 npu_inst_pe_1_0_5_U88 ( .A(npu_inst_pe_1_0_5_n37), .ZN(
        npu_inst_pe_1_0_5_n113) );
  NAND2_X1 npu_inst_pe_1_0_5_U87 ( .A1(npu_inst_pe_1_0_5_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_0_5_n60), .ZN(npu_inst_pe_1_0_5_n74) );
  OAI21_X1 npu_inst_pe_1_0_5_U86 ( .B1(npu_inst_pe_1_0_5_n63), .B2(
        npu_inst_pe_1_0_5_n60), .A(npu_inst_pe_1_0_5_n74), .ZN(
        npu_inst_pe_1_0_5_n97) );
  NAND2_X1 npu_inst_pe_1_0_5_U85 ( .A1(npu_inst_pe_1_0_5_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_0_5_n60), .ZN(npu_inst_pe_1_0_5_n73) );
  OAI21_X1 npu_inst_pe_1_0_5_U84 ( .B1(npu_inst_pe_1_0_5_n61), .B2(
        npu_inst_pe_1_0_5_n60), .A(npu_inst_pe_1_0_5_n73), .ZN(
        npu_inst_pe_1_0_5_n96) );
  NAND2_X1 npu_inst_pe_1_0_5_U83 ( .A1(npu_inst_pe_1_0_5_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_0_5_n56), .ZN(npu_inst_pe_1_0_5_n72) );
  OAI21_X1 npu_inst_pe_1_0_5_U82 ( .B1(npu_inst_pe_1_0_5_n63), .B2(
        npu_inst_pe_1_0_5_n56), .A(npu_inst_pe_1_0_5_n72), .ZN(
        npu_inst_pe_1_0_5_n95) );
  NAND2_X1 npu_inst_pe_1_0_5_U81 ( .A1(npu_inst_pe_1_0_5_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_0_5_n56), .ZN(npu_inst_pe_1_0_5_n71) );
  OAI21_X1 npu_inst_pe_1_0_5_U80 ( .B1(npu_inst_pe_1_0_5_n61), .B2(
        npu_inst_pe_1_0_5_n56), .A(npu_inst_pe_1_0_5_n71), .ZN(
        npu_inst_pe_1_0_5_n94) );
  NAND2_X1 npu_inst_pe_1_0_5_U79 ( .A1(npu_inst_pe_1_0_5_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_0_5_n52), .ZN(npu_inst_pe_1_0_5_n70) );
  OAI21_X1 npu_inst_pe_1_0_5_U78 ( .B1(npu_inst_pe_1_0_5_n63), .B2(
        npu_inst_pe_1_0_5_n52), .A(npu_inst_pe_1_0_5_n70), .ZN(
        npu_inst_pe_1_0_5_n93) );
  NAND2_X1 npu_inst_pe_1_0_5_U77 ( .A1(npu_inst_pe_1_0_5_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_0_5_n52), .ZN(npu_inst_pe_1_0_5_n69) );
  OAI21_X1 npu_inst_pe_1_0_5_U76 ( .B1(npu_inst_pe_1_0_5_n61), .B2(
        npu_inst_pe_1_0_5_n52), .A(npu_inst_pe_1_0_5_n69), .ZN(
        npu_inst_pe_1_0_5_n92) );
  NAND2_X1 npu_inst_pe_1_0_5_U75 ( .A1(npu_inst_pe_1_0_5_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_0_5_n48), .ZN(npu_inst_pe_1_0_5_n68) );
  OAI21_X1 npu_inst_pe_1_0_5_U74 ( .B1(npu_inst_pe_1_0_5_n63), .B2(
        npu_inst_pe_1_0_5_n48), .A(npu_inst_pe_1_0_5_n68), .ZN(
        npu_inst_pe_1_0_5_n91) );
  NAND2_X1 npu_inst_pe_1_0_5_U73 ( .A1(npu_inst_pe_1_0_5_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_0_5_n48), .ZN(npu_inst_pe_1_0_5_n67) );
  OAI21_X1 npu_inst_pe_1_0_5_U72 ( .B1(npu_inst_pe_1_0_5_n61), .B2(
        npu_inst_pe_1_0_5_n48), .A(npu_inst_pe_1_0_5_n67), .ZN(
        npu_inst_pe_1_0_5_n90) );
  NAND2_X1 npu_inst_pe_1_0_5_U71 ( .A1(npu_inst_pe_1_0_5_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_0_5_n44), .ZN(npu_inst_pe_1_0_5_n66) );
  OAI21_X1 npu_inst_pe_1_0_5_U70 ( .B1(npu_inst_pe_1_0_5_n63), .B2(
        npu_inst_pe_1_0_5_n44), .A(npu_inst_pe_1_0_5_n66), .ZN(
        npu_inst_pe_1_0_5_n89) );
  NAND2_X1 npu_inst_pe_1_0_5_U69 ( .A1(npu_inst_pe_1_0_5_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_0_5_n44), .ZN(npu_inst_pe_1_0_5_n65) );
  OAI21_X1 npu_inst_pe_1_0_5_U68 ( .B1(npu_inst_pe_1_0_5_n61), .B2(
        npu_inst_pe_1_0_5_n44), .A(npu_inst_pe_1_0_5_n65), .ZN(
        npu_inst_pe_1_0_5_n88) );
  NAND2_X1 npu_inst_pe_1_0_5_U67 ( .A1(npu_inst_pe_1_0_5_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_0_5_n40), .ZN(npu_inst_pe_1_0_5_n64) );
  OAI21_X1 npu_inst_pe_1_0_5_U66 ( .B1(npu_inst_pe_1_0_5_n63), .B2(
        npu_inst_pe_1_0_5_n40), .A(npu_inst_pe_1_0_5_n64), .ZN(
        npu_inst_pe_1_0_5_n87) );
  NAND2_X1 npu_inst_pe_1_0_5_U65 ( .A1(npu_inst_pe_1_0_5_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_0_5_n40), .ZN(npu_inst_pe_1_0_5_n62) );
  OAI21_X1 npu_inst_pe_1_0_5_U64 ( .B1(npu_inst_pe_1_0_5_n61), .B2(
        npu_inst_pe_1_0_5_n40), .A(npu_inst_pe_1_0_5_n62), .ZN(
        npu_inst_pe_1_0_5_n86) );
  AND2_X1 npu_inst_pe_1_0_5_U63 ( .A1(npu_inst_pe_1_0_5_int_q_acc_2_), .A2(
        npu_inst_pe_1_0_5_n1), .ZN(int_o_data_npu[18]) );
  AND2_X1 npu_inst_pe_1_0_5_U62 ( .A1(npu_inst_pe_1_0_5_int_q_acc_3_), .A2(
        npu_inst_pe_1_0_5_n2), .ZN(int_o_data_npu[19]) );
  NOR3_X1 npu_inst_pe_1_0_5_U61 ( .A1(npu_inst_pe_1_0_5_n26), .A2(npu_inst_n60), .A3(npu_inst_int_ckg[58]), .ZN(npu_inst_pe_1_0_5_n85) );
  OR2_X1 npu_inst_pe_1_0_5_U60 ( .A1(npu_inst_pe_1_0_5_n85), .A2(
        npu_inst_pe_1_0_5_n2), .ZN(npu_inst_pe_1_0_5_N84) );
  AND2_X1 npu_inst_pe_1_0_5_U59 ( .A1(npu_inst_pe_1_0_5_int_q_acc_6_), .A2(
        npu_inst_pe_1_0_5_n2), .ZN(int_o_data_npu[22]) );
  AND2_X1 npu_inst_pe_1_0_5_U58 ( .A1(npu_inst_pe_1_0_5_int_q_acc_5_), .A2(
        npu_inst_pe_1_0_5_n2), .ZN(int_o_data_npu[21]) );
  AND2_X1 npu_inst_pe_1_0_5_U57 ( .A1(npu_inst_pe_1_0_5_int_q_acc_4_), .A2(
        npu_inst_pe_1_0_5_n2), .ZN(int_o_data_npu[20]) );
  AOI222_X1 npu_inst_pe_1_0_5_U56 ( .A1(npu_inst_int_data_res_1__5__0_), .A2(
        npu_inst_pe_1_0_5_n1), .B1(npu_inst_pe_1_0_5_N73), .B2(
        npu_inst_pe_1_0_5_n76), .C1(npu_inst_pe_1_0_5_N65), .C2(
        npu_inst_pe_1_0_5_n77), .ZN(npu_inst_pe_1_0_5_n84) );
  INV_X1 npu_inst_pe_1_0_5_U55 ( .A(npu_inst_pe_1_0_5_n84), .ZN(
        npu_inst_pe_1_0_5_n101) );
  AOI222_X1 npu_inst_pe_1_0_5_U54 ( .A1(npu_inst_int_data_res_1__5__7_), .A2(
        npu_inst_pe_1_0_5_n1), .B1(npu_inst_pe_1_0_5_N80), .B2(
        npu_inst_pe_1_0_5_n76), .C1(npu_inst_pe_1_0_5_N72), .C2(
        npu_inst_pe_1_0_5_n77), .ZN(npu_inst_pe_1_0_5_n75) );
  INV_X1 npu_inst_pe_1_0_5_U53 ( .A(npu_inst_pe_1_0_5_n75), .ZN(
        npu_inst_pe_1_0_5_n33) );
  AOI222_X1 npu_inst_pe_1_0_5_U52 ( .A1(npu_inst_int_data_res_1__5__1_), .A2(
        npu_inst_pe_1_0_5_n1), .B1(npu_inst_pe_1_0_5_N74), .B2(
        npu_inst_pe_1_0_5_n76), .C1(npu_inst_pe_1_0_5_N66), .C2(
        npu_inst_pe_1_0_5_n77), .ZN(npu_inst_pe_1_0_5_n83) );
  INV_X1 npu_inst_pe_1_0_5_U51 ( .A(npu_inst_pe_1_0_5_n83), .ZN(
        npu_inst_pe_1_0_5_n100) );
  AOI222_X1 npu_inst_pe_1_0_5_U50 ( .A1(npu_inst_int_data_res_1__5__2_), .A2(
        npu_inst_pe_1_0_5_n1), .B1(npu_inst_pe_1_0_5_N75), .B2(
        npu_inst_pe_1_0_5_n76), .C1(npu_inst_pe_1_0_5_N67), .C2(
        npu_inst_pe_1_0_5_n77), .ZN(npu_inst_pe_1_0_5_n82) );
  INV_X1 npu_inst_pe_1_0_5_U49 ( .A(npu_inst_pe_1_0_5_n82), .ZN(
        npu_inst_pe_1_0_5_n99) );
  AOI222_X1 npu_inst_pe_1_0_5_U48 ( .A1(npu_inst_int_data_res_1__5__3_), .A2(
        npu_inst_pe_1_0_5_n1), .B1(npu_inst_pe_1_0_5_N76), .B2(
        npu_inst_pe_1_0_5_n76), .C1(npu_inst_pe_1_0_5_N68), .C2(
        npu_inst_pe_1_0_5_n77), .ZN(npu_inst_pe_1_0_5_n81) );
  INV_X1 npu_inst_pe_1_0_5_U47 ( .A(npu_inst_pe_1_0_5_n81), .ZN(
        npu_inst_pe_1_0_5_n98) );
  AOI222_X1 npu_inst_pe_1_0_5_U46 ( .A1(npu_inst_int_data_res_1__5__4_), .A2(
        npu_inst_pe_1_0_5_n1), .B1(npu_inst_pe_1_0_5_N77), .B2(
        npu_inst_pe_1_0_5_n76), .C1(npu_inst_pe_1_0_5_N69), .C2(
        npu_inst_pe_1_0_5_n77), .ZN(npu_inst_pe_1_0_5_n80) );
  INV_X1 npu_inst_pe_1_0_5_U45 ( .A(npu_inst_pe_1_0_5_n80), .ZN(
        npu_inst_pe_1_0_5_n36) );
  AOI222_X1 npu_inst_pe_1_0_5_U44 ( .A1(npu_inst_int_data_res_1__5__5_), .A2(
        npu_inst_pe_1_0_5_n1), .B1(npu_inst_pe_1_0_5_N78), .B2(
        npu_inst_pe_1_0_5_n76), .C1(npu_inst_pe_1_0_5_N70), .C2(
        npu_inst_pe_1_0_5_n77), .ZN(npu_inst_pe_1_0_5_n79) );
  INV_X1 npu_inst_pe_1_0_5_U43 ( .A(npu_inst_pe_1_0_5_n79), .ZN(
        npu_inst_pe_1_0_5_n35) );
  AOI222_X1 npu_inst_pe_1_0_5_U42 ( .A1(npu_inst_int_data_res_1__5__6_), .A2(
        npu_inst_pe_1_0_5_n1), .B1(npu_inst_pe_1_0_5_N79), .B2(
        npu_inst_pe_1_0_5_n76), .C1(npu_inst_pe_1_0_5_N71), .C2(
        npu_inst_pe_1_0_5_n77), .ZN(npu_inst_pe_1_0_5_n78) );
  INV_X1 npu_inst_pe_1_0_5_U41 ( .A(npu_inst_pe_1_0_5_n78), .ZN(
        npu_inst_pe_1_0_5_n34) );
  INV_X1 npu_inst_pe_1_0_5_U40 ( .A(npu_inst_pe_1_0_5_int_data_1_), .ZN(
        npu_inst_pe_1_0_5_n14) );
  AND2_X1 npu_inst_pe_1_0_5_U39 ( .A1(npu_inst_int_data_x_0__5__1_), .A2(
        npu_inst_pe_1_0_5_int_q_weight_1_), .ZN(npu_inst_pe_1_0_5_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_0_5_U38 ( .A1(npu_inst_int_data_x_0__5__0_), .A2(
        npu_inst_pe_1_0_5_int_q_weight_1_), .ZN(npu_inst_pe_1_0_5_int_data_0_)
         );
  AND2_X1 npu_inst_pe_1_0_5_U37 ( .A1(npu_inst_pe_1_0_5_n2), .A2(
        npu_inst_pe_1_0_5_int_q_acc_7_), .ZN(int_o_data_npu[23]) );
  AND2_X1 npu_inst_pe_1_0_5_U36 ( .A1(npu_inst_pe_1_0_5_int_q_acc_1_), .A2(
        npu_inst_pe_1_0_5_n1), .ZN(int_o_data_npu[17]) );
  AND2_X1 npu_inst_pe_1_0_5_U35 ( .A1(npu_inst_pe_1_0_5_int_q_acc_0_), .A2(
        npu_inst_pe_1_0_5_n1), .ZN(int_o_data_npu[16]) );
  AND2_X1 npu_inst_pe_1_0_5_U34 ( .A1(npu_inst_pe_1_0_5_N93), .A2(npu_inst_n60), .ZN(npu_inst_pe_1_0_5_o_data_v_0_) );
  AND2_X1 npu_inst_pe_1_0_5_U33 ( .A1(npu_inst_n60), .A2(npu_inst_pe_1_0_5_N94), .ZN(npu_inst_pe_1_0_5_o_data_v_1_) );
  AOI22_X1 npu_inst_pe_1_0_5_U32 ( .A1(npu_inst_n60), .A2(
        npu_inst_int_data_y_1__5__1_), .B1(npu_inst_pe_1_0_5_n3), .B2(
        npu_inst_int_data_x_0__6__1_), .ZN(npu_inst_pe_1_0_5_n63) );
  AOI22_X1 npu_inst_pe_1_0_5_U31 ( .A1(npu_inst_n60), .A2(
        npu_inst_int_data_y_1__5__0_), .B1(npu_inst_pe_1_0_5_n3), .B2(
        npu_inst_int_data_x_0__6__0_), .ZN(npu_inst_pe_1_0_5_n61) );
  INV_X1 npu_inst_pe_1_0_5_U30 ( .A(npu_inst_pe_1_0_5_int_data_0_), .ZN(
        npu_inst_pe_1_0_5_n13) );
  INV_X1 npu_inst_pe_1_0_5_U29 ( .A(npu_inst_n71), .ZN(npu_inst_pe_1_0_5_n5)
         );
  OR3_X1 npu_inst_pe_1_0_5_U28 ( .A1(npu_inst_pe_1_0_5_n6), .A2(
        npu_inst_pe_1_0_5_n8), .A3(npu_inst_pe_1_0_5_n5), .ZN(
        npu_inst_pe_1_0_5_n56) );
  OR3_X1 npu_inst_pe_1_0_5_U27 ( .A1(npu_inst_pe_1_0_5_n5), .A2(
        npu_inst_pe_1_0_5_n8), .A3(npu_inst_pe_1_0_5_n7), .ZN(
        npu_inst_pe_1_0_5_n48) );
  INV_X1 npu_inst_pe_1_0_5_U26 ( .A(npu_inst_pe_1_0_5_n5), .ZN(
        npu_inst_pe_1_0_5_n4) );
  OR3_X1 npu_inst_pe_1_0_5_U25 ( .A1(npu_inst_pe_1_0_5_n4), .A2(
        npu_inst_pe_1_0_5_n8), .A3(npu_inst_pe_1_0_5_n7), .ZN(
        npu_inst_pe_1_0_5_n52) );
  OR3_X1 npu_inst_pe_1_0_5_U24 ( .A1(npu_inst_pe_1_0_5_n6), .A2(
        npu_inst_pe_1_0_5_n8), .A3(npu_inst_pe_1_0_5_n4), .ZN(
        npu_inst_pe_1_0_5_n60) );
  NOR2_X1 npu_inst_pe_1_0_5_U23 ( .A1(npu_inst_pe_1_0_5_n60), .A2(
        npu_inst_pe_1_0_5_n3), .ZN(npu_inst_pe_1_0_5_n58) );
  NOR2_X1 npu_inst_pe_1_0_5_U22 ( .A1(npu_inst_pe_1_0_5_n56), .A2(
        npu_inst_pe_1_0_5_n3), .ZN(npu_inst_pe_1_0_5_n54) );
  NOR2_X1 npu_inst_pe_1_0_5_U21 ( .A1(npu_inst_pe_1_0_5_n52), .A2(
        npu_inst_pe_1_0_5_n3), .ZN(npu_inst_pe_1_0_5_n50) );
  NOR2_X1 npu_inst_pe_1_0_5_U20 ( .A1(npu_inst_pe_1_0_5_n48), .A2(
        npu_inst_pe_1_0_5_n3), .ZN(npu_inst_pe_1_0_5_n46) );
  NOR2_X1 npu_inst_pe_1_0_5_U19 ( .A1(npu_inst_pe_1_0_5_n40), .A2(
        npu_inst_pe_1_0_5_n3), .ZN(npu_inst_pe_1_0_5_n38) );
  NOR2_X1 npu_inst_pe_1_0_5_U18 ( .A1(npu_inst_pe_1_0_5_n44), .A2(
        npu_inst_pe_1_0_5_n3), .ZN(npu_inst_pe_1_0_5_n42) );
  BUF_X1 npu_inst_pe_1_0_5_U17 ( .A(npu_inst_n106), .Z(npu_inst_pe_1_0_5_n8)
         );
  INV_X1 npu_inst_pe_1_0_5_U16 ( .A(npu_inst_n126), .ZN(npu_inst_pe_1_0_5_n12)
         );
  INV_X1 npu_inst_pe_1_0_5_U15 ( .A(npu_inst_pe_1_0_5_n38), .ZN(
        npu_inst_pe_1_0_5_n114) );
  INV_X1 npu_inst_pe_1_0_5_U14 ( .A(npu_inst_pe_1_0_5_n58), .ZN(
        npu_inst_pe_1_0_5_n119) );
  INV_X1 npu_inst_pe_1_0_5_U13 ( .A(npu_inst_pe_1_0_5_n54), .ZN(
        npu_inst_pe_1_0_5_n118) );
  INV_X1 npu_inst_pe_1_0_5_U12 ( .A(npu_inst_pe_1_0_5_n50), .ZN(
        npu_inst_pe_1_0_5_n117) );
  INV_X1 npu_inst_pe_1_0_5_U11 ( .A(npu_inst_pe_1_0_5_n46), .ZN(
        npu_inst_pe_1_0_5_n116) );
  INV_X1 npu_inst_pe_1_0_5_U10 ( .A(npu_inst_pe_1_0_5_n42), .ZN(
        npu_inst_pe_1_0_5_n115) );
  BUF_X1 npu_inst_pe_1_0_5_U9 ( .A(npu_inst_n36), .Z(npu_inst_pe_1_0_5_n2) );
  BUF_X1 npu_inst_pe_1_0_5_U8 ( .A(npu_inst_n36), .Z(npu_inst_pe_1_0_5_n1) );
  BUF_X1 npu_inst_pe_1_0_5_U7 ( .A(npu_inst_pe_1_0_5_n12), .Z(
        npu_inst_pe_1_0_5_n11) );
  BUF_X1 npu_inst_pe_1_0_5_U6 ( .A(npu_inst_pe_1_0_5_n12), .Z(
        npu_inst_pe_1_0_5_n10) );
  BUF_X1 npu_inst_pe_1_0_5_U5 ( .A(npu_inst_pe_1_0_5_n12), .Z(
        npu_inst_pe_1_0_5_n9) );
  NOR2_X1 npu_inst_pe_1_0_5_U4 ( .A1(npu_inst_pe_1_0_5_int_q_weight_0_), .A2(
        npu_inst_pe_1_0_5_n1), .ZN(npu_inst_pe_1_0_5_n76) );
  NOR2_X1 npu_inst_pe_1_0_5_U3 ( .A1(npu_inst_pe_1_0_5_n27), .A2(
        npu_inst_pe_1_0_5_n1), .ZN(npu_inst_pe_1_0_5_n77) );
  FA_X1 npu_inst_pe_1_0_5_sub_67_U2_1 ( .A(npu_inst_pe_1_0_5_int_q_acc_1_), 
        .B(npu_inst_pe_1_0_5_n14), .CI(npu_inst_pe_1_0_5_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_0_5_sub_67_carry_2_), .S(npu_inst_pe_1_0_5_N66) );
  FA_X1 npu_inst_pe_1_0_5_add_69_U1_1 ( .A(npu_inst_pe_1_0_5_int_q_acc_1_), 
        .B(npu_inst_pe_1_0_5_int_data_1_), .CI(
        npu_inst_pe_1_0_5_add_69_carry_1_), .CO(
        npu_inst_pe_1_0_5_add_69_carry_2_), .S(npu_inst_pe_1_0_5_N74) );
  NAND3_X1 npu_inst_pe_1_0_5_U109 ( .A1(npu_inst_pe_1_0_5_n5), .A2(
        npu_inst_pe_1_0_5_n7), .A3(npu_inst_pe_1_0_5_n8), .ZN(
        npu_inst_pe_1_0_5_n44) );
  NAND3_X1 npu_inst_pe_1_0_5_U108 ( .A1(npu_inst_pe_1_0_5_n4), .A2(
        npu_inst_pe_1_0_5_n7), .A3(npu_inst_pe_1_0_5_n8), .ZN(
        npu_inst_pe_1_0_5_n40) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_0_5_n34), .CK(
        npu_inst_pe_1_0_5_net4447), .RN(npu_inst_pe_1_0_5_n9), .Q(
        npu_inst_pe_1_0_5_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_0_5_n35), .CK(
        npu_inst_pe_1_0_5_net4447), .RN(npu_inst_pe_1_0_5_n9), .Q(
        npu_inst_pe_1_0_5_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_0_5_n36), .CK(
        npu_inst_pe_1_0_5_net4447), .RN(npu_inst_pe_1_0_5_n9), .Q(
        npu_inst_pe_1_0_5_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_0_5_n98), .CK(
        npu_inst_pe_1_0_5_net4447), .RN(npu_inst_pe_1_0_5_n9), .Q(
        npu_inst_pe_1_0_5_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_0_5_n99), .CK(
        npu_inst_pe_1_0_5_net4447), .RN(npu_inst_pe_1_0_5_n9), .Q(
        npu_inst_pe_1_0_5_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_0_5_n100), 
        .CK(npu_inst_pe_1_0_5_net4447), .RN(npu_inst_pe_1_0_5_n9), .Q(
        npu_inst_pe_1_0_5_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_0_5_n33), .CK(
        npu_inst_pe_1_0_5_net4447), .RN(npu_inst_pe_1_0_5_n9), .Q(
        npu_inst_pe_1_0_5_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_0_5_n101), 
        .CK(npu_inst_pe_1_0_5_net4447), .RN(npu_inst_pe_1_0_5_n9), .Q(
        npu_inst_pe_1_0_5_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_weight_reg_0_ ( .D(npu_inst_n112), .CK(
        npu_inst_pe_1_0_5_net4453), .RN(npu_inst_pe_1_0_5_n9), .Q(
        npu_inst_pe_1_0_5_int_q_weight_0_), .QN(npu_inst_pe_1_0_5_n27) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_weight_reg_1_ ( .D(npu_inst_n118), .CK(
        npu_inst_pe_1_0_5_net4453), .RN(npu_inst_pe_1_0_5_n9), .Q(
        npu_inst_pe_1_0_5_int_q_weight_1_), .QN(npu_inst_pe_1_0_5_n26) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_0_5_n113), 
        .CK(npu_inst_pe_1_0_5_net4453), .RN(npu_inst_pe_1_0_5_n9), .Q(
        npu_inst_pe_1_0_5_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_0_5_n107), 
        .CK(npu_inst_pe_1_0_5_net4453), .RN(npu_inst_pe_1_0_5_n9), .Q(
        npu_inst_pe_1_0_5_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_0_5_n112), 
        .CK(npu_inst_pe_1_0_5_net4453), .RN(npu_inst_pe_1_0_5_n10), .Q(
        npu_inst_pe_1_0_5_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_0_5_n106), 
        .CK(npu_inst_pe_1_0_5_net4453), .RN(npu_inst_pe_1_0_5_n10), .Q(
        npu_inst_pe_1_0_5_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_0_5_n111), 
        .CK(npu_inst_pe_1_0_5_net4453), .RN(npu_inst_pe_1_0_5_n10), .Q(
        npu_inst_pe_1_0_5_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_0_5_n105), 
        .CK(npu_inst_pe_1_0_5_net4453), .RN(npu_inst_pe_1_0_5_n10), .Q(
        npu_inst_pe_1_0_5_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_0_5_n110), 
        .CK(npu_inst_pe_1_0_5_net4453), .RN(npu_inst_pe_1_0_5_n10), .Q(
        npu_inst_pe_1_0_5_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_0_5_n104), 
        .CK(npu_inst_pe_1_0_5_net4453), .RN(npu_inst_pe_1_0_5_n10), .Q(
        npu_inst_pe_1_0_5_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_0_5_n109), 
        .CK(npu_inst_pe_1_0_5_net4453), .RN(npu_inst_pe_1_0_5_n10), .Q(
        npu_inst_pe_1_0_5_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_0_5_n103), 
        .CK(npu_inst_pe_1_0_5_net4453), .RN(npu_inst_pe_1_0_5_n10), .Q(
        npu_inst_pe_1_0_5_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_0_5_n108), 
        .CK(npu_inst_pe_1_0_5_net4453), .RN(npu_inst_pe_1_0_5_n10), .Q(
        npu_inst_pe_1_0_5_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_0_5_n102), 
        .CK(npu_inst_pe_1_0_5_net4453), .RN(npu_inst_pe_1_0_5_n10), .Q(
        npu_inst_pe_1_0_5_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_0_5_n86), 
        .CK(npu_inst_pe_1_0_5_net4453), .RN(npu_inst_pe_1_0_5_n10), .Q(
        npu_inst_pe_1_0_5_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_0_5_n87), 
        .CK(npu_inst_pe_1_0_5_net4453), .RN(npu_inst_pe_1_0_5_n10), .Q(
        npu_inst_pe_1_0_5_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_0_5_n88), 
        .CK(npu_inst_pe_1_0_5_net4453), .RN(npu_inst_pe_1_0_5_n11), .Q(
        npu_inst_pe_1_0_5_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_0_5_n89), 
        .CK(npu_inst_pe_1_0_5_net4453), .RN(npu_inst_pe_1_0_5_n11), .Q(
        npu_inst_pe_1_0_5_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_0_5_n90), 
        .CK(npu_inst_pe_1_0_5_net4453), .RN(npu_inst_pe_1_0_5_n11), .Q(
        npu_inst_pe_1_0_5_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_0_5_n91), 
        .CK(npu_inst_pe_1_0_5_net4453), .RN(npu_inst_pe_1_0_5_n11), .Q(
        npu_inst_pe_1_0_5_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_0_5_n92), 
        .CK(npu_inst_pe_1_0_5_net4453), .RN(npu_inst_pe_1_0_5_n11), .Q(
        npu_inst_pe_1_0_5_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_0_5_n93), 
        .CK(npu_inst_pe_1_0_5_net4453), .RN(npu_inst_pe_1_0_5_n11), .Q(
        npu_inst_pe_1_0_5_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_0_5_n94), 
        .CK(npu_inst_pe_1_0_5_net4453), .RN(npu_inst_pe_1_0_5_n11), .Q(
        npu_inst_pe_1_0_5_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_0_5_n95), 
        .CK(npu_inst_pe_1_0_5_net4453), .RN(npu_inst_pe_1_0_5_n11), .Q(
        npu_inst_pe_1_0_5_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_0_5_n96), 
        .CK(npu_inst_pe_1_0_5_net4453), .RN(npu_inst_pe_1_0_5_n11), .Q(
        npu_inst_pe_1_0_5_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_0_5_n97), 
        .CK(npu_inst_pe_1_0_5_net4453), .RN(npu_inst_pe_1_0_5_n11), .Q(
        npu_inst_pe_1_0_5_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_0_5_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_0_5_N84), .SE(1'b0), .GCK(npu_inst_pe_1_0_5_net4447) );
  CLKGATETST_X1 npu_inst_pe_1_0_5_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n66), .SE(1'b0), .GCK(npu_inst_pe_1_0_5_net4453) );
  MUX2_X1 npu_inst_pe_1_0_6_U162 ( .A(npu_inst_pe_1_0_6_n32), .B(
        npu_inst_pe_1_0_6_n29), .S(npu_inst_pe_1_0_6_n8), .Z(
        npu_inst_pe_1_0_6_N93) );
  MUX2_X1 npu_inst_pe_1_0_6_U161 ( .A(npu_inst_pe_1_0_6_n31), .B(
        npu_inst_pe_1_0_6_n30), .S(npu_inst_pe_1_0_6_n6), .Z(
        npu_inst_pe_1_0_6_n32) );
  MUX2_X1 npu_inst_pe_1_0_6_U160 ( .A(npu_inst_pe_1_0_6_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_0_6_int_q_reg_v_1__0_), .S(npu_inst_pe_1_0_6_n4), .Z(
        npu_inst_pe_1_0_6_n31) );
  MUX2_X1 npu_inst_pe_1_0_6_U159 ( .A(npu_inst_pe_1_0_6_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_0_6_int_q_reg_v_3__0_), .S(npu_inst_pe_1_0_6_n4), .Z(
        npu_inst_pe_1_0_6_n30) );
  MUX2_X1 npu_inst_pe_1_0_6_U158 ( .A(npu_inst_pe_1_0_6_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_0_6_int_q_reg_v_5__0_), .S(npu_inst_pe_1_0_6_n4), .Z(
        npu_inst_pe_1_0_6_n29) );
  MUX2_X1 npu_inst_pe_1_0_6_U157 ( .A(npu_inst_pe_1_0_6_n28), .B(
        npu_inst_pe_1_0_6_n23), .S(npu_inst_pe_1_0_6_n8), .Z(
        npu_inst_pe_1_0_6_N94) );
  MUX2_X1 npu_inst_pe_1_0_6_U156 ( .A(npu_inst_pe_1_0_6_n25), .B(
        npu_inst_pe_1_0_6_n24), .S(npu_inst_pe_1_0_6_n6), .Z(
        npu_inst_pe_1_0_6_n28) );
  MUX2_X1 npu_inst_pe_1_0_6_U155 ( .A(npu_inst_pe_1_0_6_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_0_6_int_q_reg_v_1__1_), .S(npu_inst_pe_1_0_6_n4), .Z(
        npu_inst_pe_1_0_6_n25) );
  MUX2_X1 npu_inst_pe_1_0_6_U154 ( .A(npu_inst_pe_1_0_6_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_0_6_int_q_reg_v_3__1_), .S(npu_inst_pe_1_0_6_n4), .Z(
        npu_inst_pe_1_0_6_n24) );
  MUX2_X1 npu_inst_pe_1_0_6_U153 ( .A(npu_inst_pe_1_0_6_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_0_6_int_q_reg_v_5__1_), .S(npu_inst_pe_1_0_6_n4), .Z(
        npu_inst_pe_1_0_6_n23) );
  MUX2_X1 npu_inst_pe_1_0_6_U152 ( .A(npu_inst_pe_1_0_6_n22), .B(
        npu_inst_pe_1_0_6_n19), .S(npu_inst_pe_1_0_6_n8), .Z(
        npu_inst_int_data_x_0__6__1_) );
  MUX2_X1 npu_inst_pe_1_0_6_U151 ( .A(npu_inst_pe_1_0_6_n21), .B(
        npu_inst_pe_1_0_6_n20), .S(npu_inst_pe_1_0_6_n6), .Z(
        npu_inst_pe_1_0_6_n22) );
  MUX2_X1 npu_inst_pe_1_0_6_U150 ( .A(npu_inst_pe_1_0_6_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_0_6_int_q_reg_h_1__1_), .S(npu_inst_pe_1_0_6_n4), .Z(
        npu_inst_pe_1_0_6_n21) );
  MUX2_X1 npu_inst_pe_1_0_6_U149 ( .A(npu_inst_pe_1_0_6_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_0_6_int_q_reg_h_3__1_), .S(npu_inst_pe_1_0_6_n4), .Z(
        npu_inst_pe_1_0_6_n20) );
  MUX2_X1 npu_inst_pe_1_0_6_U148 ( .A(npu_inst_pe_1_0_6_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_0_6_int_q_reg_h_5__1_), .S(npu_inst_pe_1_0_6_n4), .Z(
        npu_inst_pe_1_0_6_n19) );
  MUX2_X1 npu_inst_pe_1_0_6_U147 ( .A(npu_inst_pe_1_0_6_n18), .B(
        npu_inst_pe_1_0_6_n15), .S(npu_inst_pe_1_0_6_n8), .Z(
        npu_inst_int_data_x_0__6__0_) );
  MUX2_X1 npu_inst_pe_1_0_6_U146 ( .A(npu_inst_pe_1_0_6_n17), .B(
        npu_inst_pe_1_0_6_n16), .S(npu_inst_pe_1_0_6_n6), .Z(
        npu_inst_pe_1_0_6_n18) );
  MUX2_X1 npu_inst_pe_1_0_6_U145 ( .A(npu_inst_pe_1_0_6_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_0_6_int_q_reg_h_1__0_), .S(npu_inst_pe_1_0_6_n4), .Z(
        npu_inst_pe_1_0_6_n17) );
  MUX2_X1 npu_inst_pe_1_0_6_U144 ( .A(npu_inst_pe_1_0_6_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_0_6_int_q_reg_h_3__0_), .S(npu_inst_pe_1_0_6_n4), .Z(
        npu_inst_pe_1_0_6_n16) );
  MUX2_X1 npu_inst_pe_1_0_6_U143 ( .A(npu_inst_pe_1_0_6_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_0_6_int_q_reg_h_5__0_), .S(npu_inst_pe_1_0_6_n4), .Z(
        npu_inst_pe_1_0_6_n15) );
  XOR2_X1 npu_inst_pe_1_0_6_U142 ( .A(npu_inst_pe_1_0_6_int_data_0_), .B(
        npu_inst_pe_1_0_6_int_q_acc_0_), .Z(npu_inst_pe_1_0_6_N73) );
  AND2_X1 npu_inst_pe_1_0_6_U141 ( .A1(npu_inst_pe_1_0_6_int_q_acc_0_), .A2(
        npu_inst_pe_1_0_6_int_data_0_), .ZN(npu_inst_pe_1_0_6_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_0_6_U140 ( .A(npu_inst_pe_1_0_6_int_q_acc_0_), .B(
        npu_inst_pe_1_0_6_n13), .ZN(npu_inst_pe_1_0_6_N65) );
  OR2_X1 npu_inst_pe_1_0_6_U139 ( .A1(npu_inst_pe_1_0_6_n13), .A2(
        npu_inst_pe_1_0_6_int_q_acc_0_), .ZN(npu_inst_pe_1_0_6_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_0_6_U138 ( .A(npu_inst_pe_1_0_6_int_q_acc_2_), .B(
        npu_inst_pe_1_0_6_add_69_carry_2_), .Z(npu_inst_pe_1_0_6_N75) );
  AND2_X1 npu_inst_pe_1_0_6_U137 ( .A1(npu_inst_pe_1_0_6_add_69_carry_2_), 
        .A2(npu_inst_pe_1_0_6_int_q_acc_2_), .ZN(
        npu_inst_pe_1_0_6_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_0_6_U136 ( .A(npu_inst_pe_1_0_6_int_q_acc_3_), .B(
        npu_inst_pe_1_0_6_add_69_carry_3_), .Z(npu_inst_pe_1_0_6_N76) );
  AND2_X1 npu_inst_pe_1_0_6_U135 ( .A1(npu_inst_pe_1_0_6_add_69_carry_3_), 
        .A2(npu_inst_pe_1_0_6_int_q_acc_3_), .ZN(
        npu_inst_pe_1_0_6_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_0_6_U134 ( .A(npu_inst_pe_1_0_6_int_q_acc_4_), .B(
        npu_inst_pe_1_0_6_add_69_carry_4_), .Z(npu_inst_pe_1_0_6_N77) );
  AND2_X1 npu_inst_pe_1_0_6_U133 ( .A1(npu_inst_pe_1_0_6_add_69_carry_4_), 
        .A2(npu_inst_pe_1_0_6_int_q_acc_4_), .ZN(
        npu_inst_pe_1_0_6_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_0_6_U132 ( .A(npu_inst_pe_1_0_6_int_q_acc_5_), .B(
        npu_inst_pe_1_0_6_add_69_carry_5_), .Z(npu_inst_pe_1_0_6_N78) );
  AND2_X1 npu_inst_pe_1_0_6_U131 ( .A1(npu_inst_pe_1_0_6_add_69_carry_5_), 
        .A2(npu_inst_pe_1_0_6_int_q_acc_5_), .ZN(
        npu_inst_pe_1_0_6_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_0_6_U130 ( .A(npu_inst_pe_1_0_6_int_q_acc_6_), .B(
        npu_inst_pe_1_0_6_add_69_carry_6_), .Z(npu_inst_pe_1_0_6_N79) );
  AND2_X1 npu_inst_pe_1_0_6_U129 ( .A1(npu_inst_pe_1_0_6_add_69_carry_6_), 
        .A2(npu_inst_pe_1_0_6_int_q_acc_6_), .ZN(
        npu_inst_pe_1_0_6_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_0_6_U128 ( .A(npu_inst_pe_1_0_6_int_q_acc_7_), .B(
        npu_inst_pe_1_0_6_add_69_carry_7_), .Z(npu_inst_pe_1_0_6_N80) );
  XNOR2_X1 npu_inst_pe_1_0_6_U127 ( .A(npu_inst_pe_1_0_6_sub_67_carry_2_), .B(
        npu_inst_pe_1_0_6_int_q_acc_2_), .ZN(npu_inst_pe_1_0_6_N67) );
  OR2_X1 npu_inst_pe_1_0_6_U126 ( .A1(npu_inst_pe_1_0_6_int_q_acc_2_), .A2(
        npu_inst_pe_1_0_6_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_0_6_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_0_6_U125 ( .A(npu_inst_pe_1_0_6_sub_67_carry_3_), .B(
        npu_inst_pe_1_0_6_int_q_acc_3_), .ZN(npu_inst_pe_1_0_6_N68) );
  OR2_X1 npu_inst_pe_1_0_6_U124 ( .A1(npu_inst_pe_1_0_6_int_q_acc_3_), .A2(
        npu_inst_pe_1_0_6_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_0_6_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_0_6_U123 ( .A(npu_inst_pe_1_0_6_sub_67_carry_4_), .B(
        npu_inst_pe_1_0_6_int_q_acc_4_), .ZN(npu_inst_pe_1_0_6_N69) );
  OR2_X1 npu_inst_pe_1_0_6_U122 ( .A1(npu_inst_pe_1_0_6_int_q_acc_4_), .A2(
        npu_inst_pe_1_0_6_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_0_6_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_0_6_U121 ( .A(npu_inst_pe_1_0_6_sub_67_carry_5_), .B(
        npu_inst_pe_1_0_6_int_q_acc_5_), .ZN(npu_inst_pe_1_0_6_N70) );
  OR2_X1 npu_inst_pe_1_0_6_U120 ( .A1(npu_inst_pe_1_0_6_int_q_acc_5_), .A2(
        npu_inst_pe_1_0_6_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_0_6_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_0_6_U119 ( .A(npu_inst_pe_1_0_6_sub_67_carry_6_), .B(
        npu_inst_pe_1_0_6_int_q_acc_6_), .ZN(npu_inst_pe_1_0_6_N71) );
  OR2_X1 npu_inst_pe_1_0_6_U118 ( .A1(npu_inst_pe_1_0_6_int_q_acc_6_), .A2(
        npu_inst_pe_1_0_6_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_0_6_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_0_6_U117 ( .A(npu_inst_pe_1_0_6_int_q_acc_7_), .B(
        npu_inst_pe_1_0_6_sub_67_carry_7_), .ZN(npu_inst_pe_1_0_6_N72) );
  INV_X1 npu_inst_pe_1_0_6_U116 ( .A(npu_inst_n79), .ZN(npu_inst_pe_1_0_6_n7)
         );
  INV_X1 npu_inst_pe_1_0_6_U115 ( .A(npu_inst_pe_1_0_6_n7), .ZN(
        npu_inst_pe_1_0_6_n6) );
  INV_X1 npu_inst_pe_1_0_6_U114 ( .A(npu_inst_n60), .ZN(npu_inst_pe_1_0_6_n3)
         );
  AOI22_X1 npu_inst_pe_1_0_6_U113 ( .A1(npu_inst_int_data_y_1__6__0_), .A2(
        npu_inst_pe_1_0_6_n58), .B1(npu_inst_pe_1_0_6_n119), .B2(
        npu_inst_pe_1_0_6_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_0_6_n57) );
  INV_X1 npu_inst_pe_1_0_6_U112 ( .A(npu_inst_pe_1_0_6_n57), .ZN(
        npu_inst_pe_1_0_6_n108) );
  AOI22_X1 npu_inst_pe_1_0_6_U111 ( .A1(npu_inst_int_data_y_1__6__0_), .A2(
        npu_inst_pe_1_0_6_n54), .B1(npu_inst_pe_1_0_6_n118), .B2(
        npu_inst_pe_1_0_6_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_0_6_n53) );
  INV_X1 npu_inst_pe_1_0_6_U110 ( .A(npu_inst_pe_1_0_6_n53), .ZN(
        npu_inst_pe_1_0_6_n109) );
  AOI22_X1 npu_inst_pe_1_0_6_U107 ( .A1(npu_inst_int_data_y_1__6__0_), .A2(
        npu_inst_pe_1_0_6_n50), .B1(npu_inst_pe_1_0_6_n117), .B2(
        npu_inst_pe_1_0_6_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_0_6_n49) );
  INV_X1 npu_inst_pe_1_0_6_U106 ( .A(npu_inst_pe_1_0_6_n49), .ZN(
        npu_inst_pe_1_0_6_n110) );
  AOI22_X1 npu_inst_pe_1_0_6_U105 ( .A1(npu_inst_int_data_y_1__6__0_), .A2(
        npu_inst_pe_1_0_6_n46), .B1(npu_inst_pe_1_0_6_n116), .B2(
        npu_inst_pe_1_0_6_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_0_6_n45) );
  INV_X1 npu_inst_pe_1_0_6_U104 ( .A(npu_inst_pe_1_0_6_n45), .ZN(
        npu_inst_pe_1_0_6_n111) );
  AOI22_X1 npu_inst_pe_1_0_6_U103 ( .A1(npu_inst_int_data_y_1__6__0_), .A2(
        npu_inst_pe_1_0_6_n42), .B1(npu_inst_pe_1_0_6_n115), .B2(
        npu_inst_pe_1_0_6_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_0_6_n41) );
  INV_X1 npu_inst_pe_1_0_6_U102 ( .A(npu_inst_pe_1_0_6_n41), .ZN(
        npu_inst_pe_1_0_6_n112) );
  AOI22_X1 npu_inst_pe_1_0_6_U101 ( .A1(npu_inst_int_data_y_1__6__1_), .A2(
        npu_inst_pe_1_0_6_n58), .B1(npu_inst_pe_1_0_6_n119), .B2(
        npu_inst_pe_1_0_6_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_0_6_n59) );
  INV_X1 npu_inst_pe_1_0_6_U100 ( .A(npu_inst_pe_1_0_6_n59), .ZN(
        npu_inst_pe_1_0_6_n102) );
  AOI22_X1 npu_inst_pe_1_0_6_U99 ( .A1(npu_inst_int_data_y_1__6__1_), .A2(
        npu_inst_pe_1_0_6_n54), .B1(npu_inst_pe_1_0_6_n118), .B2(
        npu_inst_pe_1_0_6_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_0_6_n55) );
  INV_X1 npu_inst_pe_1_0_6_U98 ( .A(npu_inst_pe_1_0_6_n55), .ZN(
        npu_inst_pe_1_0_6_n103) );
  AOI22_X1 npu_inst_pe_1_0_6_U97 ( .A1(npu_inst_int_data_y_1__6__1_), .A2(
        npu_inst_pe_1_0_6_n50), .B1(npu_inst_pe_1_0_6_n117), .B2(
        npu_inst_pe_1_0_6_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_0_6_n51) );
  INV_X1 npu_inst_pe_1_0_6_U96 ( .A(npu_inst_pe_1_0_6_n51), .ZN(
        npu_inst_pe_1_0_6_n104) );
  AOI22_X1 npu_inst_pe_1_0_6_U95 ( .A1(npu_inst_int_data_y_1__6__1_), .A2(
        npu_inst_pe_1_0_6_n46), .B1(npu_inst_pe_1_0_6_n116), .B2(
        npu_inst_pe_1_0_6_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_0_6_n47) );
  INV_X1 npu_inst_pe_1_0_6_U94 ( .A(npu_inst_pe_1_0_6_n47), .ZN(
        npu_inst_pe_1_0_6_n105) );
  AOI22_X1 npu_inst_pe_1_0_6_U93 ( .A1(npu_inst_int_data_y_1__6__1_), .A2(
        npu_inst_pe_1_0_6_n42), .B1(npu_inst_pe_1_0_6_n115), .B2(
        npu_inst_pe_1_0_6_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_0_6_n43) );
  INV_X1 npu_inst_pe_1_0_6_U92 ( .A(npu_inst_pe_1_0_6_n43), .ZN(
        npu_inst_pe_1_0_6_n106) );
  AOI22_X1 npu_inst_pe_1_0_6_U91 ( .A1(npu_inst_pe_1_0_6_n38), .A2(
        npu_inst_int_data_y_1__6__1_), .B1(npu_inst_pe_1_0_6_n114), .B2(
        npu_inst_pe_1_0_6_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_0_6_n39) );
  INV_X1 npu_inst_pe_1_0_6_U90 ( .A(npu_inst_pe_1_0_6_n39), .ZN(
        npu_inst_pe_1_0_6_n107) );
  AOI22_X1 npu_inst_pe_1_0_6_U89 ( .A1(npu_inst_pe_1_0_6_n38), .A2(
        npu_inst_int_data_y_1__6__0_), .B1(npu_inst_pe_1_0_6_n114), .B2(
        npu_inst_pe_1_0_6_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_0_6_n37) );
  INV_X1 npu_inst_pe_1_0_6_U88 ( .A(npu_inst_pe_1_0_6_n37), .ZN(
        npu_inst_pe_1_0_6_n113) );
  NAND2_X1 npu_inst_pe_1_0_6_U87 ( .A1(npu_inst_pe_1_0_6_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_0_6_n60), .ZN(npu_inst_pe_1_0_6_n74) );
  OAI21_X1 npu_inst_pe_1_0_6_U86 ( .B1(npu_inst_pe_1_0_6_n63), .B2(
        npu_inst_pe_1_0_6_n60), .A(npu_inst_pe_1_0_6_n74), .ZN(
        npu_inst_pe_1_0_6_n97) );
  NAND2_X1 npu_inst_pe_1_0_6_U85 ( .A1(npu_inst_pe_1_0_6_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_0_6_n60), .ZN(npu_inst_pe_1_0_6_n73) );
  OAI21_X1 npu_inst_pe_1_0_6_U84 ( .B1(npu_inst_pe_1_0_6_n61), .B2(
        npu_inst_pe_1_0_6_n60), .A(npu_inst_pe_1_0_6_n73), .ZN(
        npu_inst_pe_1_0_6_n96) );
  NAND2_X1 npu_inst_pe_1_0_6_U83 ( .A1(npu_inst_pe_1_0_6_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_0_6_n56), .ZN(npu_inst_pe_1_0_6_n72) );
  OAI21_X1 npu_inst_pe_1_0_6_U82 ( .B1(npu_inst_pe_1_0_6_n63), .B2(
        npu_inst_pe_1_0_6_n56), .A(npu_inst_pe_1_0_6_n72), .ZN(
        npu_inst_pe_1_0_6_n95) );
  NAND2_X1 npu_inst_pe_1_0_6_U81 ( .A1(npu_inst_pe_1_0_6_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_0_6_n56), .ZN(npu_inst_pe_1_0_6_n71) );
  OAI21_X1 npu_inst_pe_1_0_6_U80 ( .B1(npu_inst_pe_1_0_6_n61), .B2(
        npu_inst_pe_1_0_6_n56), .A(npu_inst_pe_1_0_6_n71), .ZN(
        npu_inst_pe_1_0_6_n94) );
  NAND2_X1 npu_inst_pe_1_0_6_U79 ( .A1(npu_inst_pe_1_0_6_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_0_6_n52), .ZN(npu_inst_pe_1_0_6_n70) );
  OAI21_X1 npu_inst_pe_1_0_6_U78 ( .B1(npu_inst_pe_1_0_6_n63), .B2(
        npu_inst_pe_1_0_6_n52), .A(npu_inst_pe_1_0_6_n70), .ZN(
        npu_inst_pe_1_0_6_n93) );
  NAND2_X1 npu_inst_pe_1_0_6_U77 ( .A1(npu_inst_pe_1_0_6_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_0_6_n52), .ZN(npu_inst_pe_1_0_6_n69) );
  OAI21_X1 npu_inst_pe_1_0_6_U76 ( .B1(npu_inst_pe_1_0_6_n61), .B2(
        npu_inst_pe_1_0_6_n52), .A(npu_inst_pe_1_0_6_n69), .ZN(
        npu_inst_pe_1_0_6_n92) );
  NAND2_X1 npu_inst_pe_1_0_6_U75 ( .A1(npu_inst_pe_1_0_6_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_0_6_n48), .ZN(npu_inst_pe_1_0_6_n68) );
  OAI21_X1 npu_inst_pe_1_0_6_U74 ( .B1(npu_inst_pe_1_0_6_n63), .B2(
        npu_inst_pe_1_0_6_n48), .A(npu_inst_pe_1_0_6_n68), .ZN(
        npu_inst_pe_1_0_6_n91) );
  NAND2_X1 npu_inst_pe_1_0_6_U73 ( .A1(npu_inst_pe_1_0_6_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_0_6_n48), .ZN(npu_inst_pe_1_0_6_n67) );
  OAI21_X1 npu_inst_pe_1_0_6_U72 ( .B1(npu_inst_pe_1_0_6_n61), .B2(
        npu_inst_pe_1_0_6_n48), .A(npu_inst_pe_1_0_6_n67), .ZN(
        npu_inst_pe_1_0_6_n90) );
  NAND2_X1 npu_inst_pe_1_0_6_U71 ( .A1(npu_inst_pe_1_0_6_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_0_6_n44), .ZN(npu_inst_pe_1_0_6_n66) );
  OAI21_X1 npu_inst_pe_1_0_6_U70 ( .B1(npu_inst_pe_1_0_6_n63), .B2(
        npu_inst_pe_1_0_6_n44), .A(npu_inst_pe_1_0_6_n66), .ZN(
        npu_inst_pe_1_0_6_n89) );
  NAND2_X1 npu_inst_pe_1_0_6_U69 ( .A1(npu_inst_pe_1_0_6_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_0_6_n44), .ZN(npu_inst_pe_1_0_6_n65) );
  OAI21_X1 npu_inst_pe_1_0_6_U68 ( .B1(npu_inst_pe_1_0_6_n61), .B2(
        npu_inst_pe_1_0_6_n44), .A(npu_inst_pe_1_0_6_n65), .ZN(
        npu_inst_pe_1_0_6_n88) );
  NAND2_X1 npu_inst_pe_1_0_6_U67 ( .A1(npu_inst_pe_1_0_6_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_0_6_n40), .ZN(npu_inst_pe_1_0_6_n64) );
  OAI21_X1 npu_inst_pe_1_0_6_U66 ( .B1(npu_inst_pe_1_0_6_n63), .B2(
        npu_inst_pe_1_0_6_n40), .A(npu_inst_pe_1_0_6_n64), .ZN(
        npu_inst_pe_1_0_6_n87) );
  NAND2_X1 npu_inst_pe_1_0_6_U65 ( .A1(npu_inst_pe_1_0_6_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_0_6_n40), .ZN(npu_inst_pe_1_0_6_n62) );
  OAI21_X1 npu_inst_pe_1_0_6_U64 ( .B1(npu_inst_pe_1_0_6_n61), .B2(
        npu_inst_pe_1_0_6_n40), .A(npu_inst_pe_1_0_6_n62), .ZN(
        npu_inst_pe_1_0_6_n86) );
  AND2_X1 npu_inst_pe_1_0_6_U63 ( .A1(npu_inst_pe_1_0_6_int_q_acc_2_), .A2(
        npu_inst_pe_1_0_6_n1), .ZN(int_o_data_npu[10]) );
  AND2_X1 npu_inst_pe_1_0_6_U62 ( .A1(npu_inst_pe_1_0_6_int_q_acc_3_), .A2(
        npu_inst_pe_1_0_6_n2), .ZN(int_o_data_npu[11]) );
  NOR3_X1 npu_inst_pe_1_0_6_U61 ( .A1(npu_inst_pe_1_0_6_n26), .A2(npu_inst_n60), .A3(npu_inst_int_ckg[57]), .ZN(npu_inst_pe_1_0_6_n85) );
  OR2_X1 npu_inst_pe_1_0_6_U60 ( .A1(npu_inst_pe_1_0_6_n85), .A2(
        npu_inst_pe_1_0_6_n2), .ZN(npu_inst_pe_1_0_6_N84) );
  AND2_X1 npu_inst_pe_1_0_6_U59 ( .A1(npu_inst_pe_1_0_6_int_q_acc_6_), .A2(
        npu_inst_pe_1_0_6_n2), .ZN(int_o_data_npu[14]) );
  AND2_X1 npu_inst_pe_1_0_6_U58 ( .A1(npu_inst_pe_1_0_6_int_q_acc_5_), .A2(
        npu_inst_pe_1_0_6_n2), .ZN(int_o_data_npu[13]) );
  AND2_X1 npu_inst_pe_1_0_6_U57 ( .A1(npu_inst_pe_1_0_6_int_q_acc_4_), .A2(
        npu_inst_pe_1_0_6_n2), .ZN(int_o_data_npu[12]) );
  AOI222_X1 npu_inst_pe_1_0_6_U56 ( .A1(npu_inst_int_data_res_1__6__0_), .A2(
        npu_inst_pe_1_0_6_n1), .B1(npu_inst_pe_1_0_6_N73), .B2(
        npu_inst_pe_1_0_6_n76), .C1(npu_inst_pe_1_0_6_N65), .C2(
        npu_inst_pe_1_0_6_n77), .ZN(npu_inst_pe_1_0_6_n84) );
  INV_X1 npu_inst_pe_1_0_6_U55 ( .A(npu_inst_pe_1_0_6_n84), .ZN(
        npu_inst_pe_1_0_6_n101) );
  AOI222_X1 npu_inst_pe_1_0_6_U54 ( .A1(npu_inst_int_data_res_1__6__7_), .A2(
        npu_inst_pe_1_0_6_n1), .B1(npu_inst_pe_1_0_6_N80), .B2(
        npu_inst_pe_1_0_6_n76), .C1(npu_inst_pe_1_0_6_N72), .C2(
        npu_inst_pe_1_0_6_n77), .ZN(npu_inst_pe_1_0_6_n75) );
  INV_X1 npu_inst_pe_1_0_6_U53 ( .A(npu_inst_pe_1_0_6_n75), .ZN(
        npu_inst_pe_1_0_6_n33) );
  AOI222_X1 npu_inst_pe_1_0_6_U52 ( .A1(npu_inst_int_data_res_1__6__1_), .A2(
        npu_inst_pe_1_0_6_n1), .B1(npu_inst_pe_1_0_6_N74), .B2(
        npu_inst_pe_1_0_6_n76), .C1(npu_inst_pe_1_0_6_N66), .C2(
        npu_inst_pe_1_0_6_n77), .ZN(npu_inst_pe_1_0_6_n83) );
  INV_X1 npu_inst_pe_1_0_6_U51 ( .A(npu_inst_pe_1_0_6_n83), .ZN(
        npu_inst_pe_1_0_6_n100) );
  AOI222_X1 npu_inst_pe_1_0_6_U50 ( .A1(npu_inst_int_data_res_1__6__2_), .A2(
        npu_inst_pe_1_0_6_n1), .B1(npu_inst_pe_1_0_6_N75), .B2(
        npu_inst_pe_1_0_6_n76), .C1(npu_inst_pe_1_0_6_N67), .C2(
        npu_inst_pe_1_0_6_n77), .ZN(npu_inst_pe_1_0_6_n82) );
  INV_X1 npu_inst_pe_1_0_6_U49 ( .A(npu_inst_pe_1_0_6_n82), .ZN(
        npu_inst_pe_1_0_6_n99) );
  AOI222_X1 npu_inst_pe_1_0_6_U48 ( .A1(npu_inst_int_data_res_1__6__3_), .A2(
        npu_inst_pe_1_0_6_n1), .B1(npu_inst_pe_1_0_6_N76), .B2(
        npu_inst_pe_1_0_6_n76), .C1(npu_inst_pe_1_0_6_N68), .C2(
        npu_inst_pe_1_0_6_n77), .ZN(npu_inst_pe_1_0_6_n81) );
  INV_X1 npu_inst_pe_1_0_6_U47 ( .A(npu_inst_pe_1_0_6_n81), .ZN(
        npu_inst_pe_1_0_6_n98) );
  AOI222_X1 npu_inst_pe_1_0_6_U46 ( .A1(npu_inst_int_data_res_1__6__4_), .A2(
        npu_inst_pe_1_0_6_n1), .B1(npu_inst_pe_1_0_6_N77), .B2(
        npu_inst_pe_1_0_6_n76), .C1(npu_inst_pe_1_0_6_N69), .C2(
        npu_inst_pe_1_0_6_n77), .ZN(npu_inst_pe_1_0_6_n80) );
  INV_X1 npu_inst_pe_1_0_6_U45 ( .A(npu_inst_pe_1_0_6_n80), .ZN(
        npu_inst_pe_1_0_6_n36) );
  AOI222_X1 npu_inst_pe_1_0_6_U44 ( .A1(npu_inst_int_data_res_1__6__5_), .A2(
        npu_inst_pe_1_0_6_n1), .B1(npu_inst_pe_1_0_6_N78), .B2(
        npu_inst_pe_1_0_6_n76), .C1(npu_inst_pe_1_0_6_N70), .C2(
        npu_inst_pe_1_0_6_n77), .ZN(npu_inst_pe_1_0_6_n79) );
  INV_X1 npu_inst_pe_1_0_6_U43 ( .A(npu_inst_pe_1_0_6_n79), .ZN(
        npu_inst_pe_1_0_6_n35) );
  AOI222_X1 npu_inst_pe_1_0_6_U42 ( .A1(npu_inst_int_data_res_1__6__6_), .A2(
        npu_inst_pe_1_0_6_n1), .B1(npu_inst_pe_1_0_6_N79), .B2(
        npu_inst_pe_1_0_6_n76), .C1(npu_inst_pe_1_0_6_N71), .C2(
        npu_inst_pe_1_0_6_n77), .ZN(npu_inst_pe_1_0_6_n78) );
  INV_X1 npu_inst_pe_1_0_6_U41 ( .A(npu_inst_pe_1_0_6_n78), .ZN(
        npu_inst_pe_1_0_6_n34) );
  INV_X1 npu_inst_pe_1_0_6_U40 ( .A(npu_inst_pe_1_0_6_int_data_1_), .ZN(
        npu_inst_pe_1_0_6_n14) );
  AND2_X1 npu_inst_pe_1_0_6_U39 ( .A1(npu_inst_int_data_x_0__6__1_), .A2(
        npu_inst_pe_1_0_6_int_q_weight_1_), .ZN(npu_inst_pe_1_0_6_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_0_6_U38 ( .A1(npu_inst_int_data_x_0__6__0_), .A2(
        npu_inst_pe_1_0_6_int_q_weight_1_), .ZN(npu_inst_pe_1_0_6_int_data_0_)
         );
  AND2_X1 npu_inst_pe_1_0_6_U37 ( .A1(npu_inst_pe_1_0_6_n2), .A2(
        npu_inst_pe_1_0_6_int_q_acc_7_), .ZN(int_o_data_npu[15]) );
  AND2_X1 npu_inst_pe_1_0_6_U36 ( .A1(npu_inst_pe_1_0_6_int_q_acc_1_), .A2(
        npu_inst_pe_1_0_6_n1), .ZN(int_o_data_npu[9]) );
  AND2_X1 npu_inst_pe_1_0_6_U35 ( .A1(npu_inst_pe_1_0_6_int_q_acc_0_), .A2(
        npu_inst_pe_1_0_6_n1), .ZN(int_o_data_npu[8]) );
  AND2_X1 npu_inst_pe_1_0_6_U34 ( .A1(npu_inst_pe_1_0_6_N93), .A2(npu_inst_n60), .ZN(npu_inst_pe_1_0_6_o_data_v_0_) );
  AND2_X1 npu_inst_pe_1_0_6_U33 ( .A1(npu_inst_n60), .A2(npu_inst_pe_1_0_6_N94), .ZN(npu_inst_pe_1_0_6_o_data_v_1_) );
  AOI22_X1 npu_inst_pe_1_0_6_U32 ( .A1(npu_inst_n60), .A2(
        npu_inst_int_data_y_1__6__1_), .B1(npu_inst_pe_1_0_6_n3), .B2(
        npu_inst_int_data_x_0__7__1_), .ZN(npu_inst_pe_1_0_6_n63) );
  AOI22_X1 npu_inst_pe_1_0_6_U31 ( .A1(npu_inst_n60), .A2(
        npu_inst_int_data_y_1__6__0_), .B1(npu_inst_pe_1_0_6_n3), .B2(
        npu_inst_int_data_x_0__7__0_), .ZN(npu_inst_pe_1_0_6_n61) );
  INV_X1 npu_inst_pe_1_0_6_U30 ( .A(npu_inst_pe_1_0_6_int_data_0_), .ZN(
        npu_inst_pe_1_0_6_n13) );
  INV_X1 npu_inst_pe_1_0_6_U29 ( .A(npu_inst_n71), .ZN(npu_inst_pe_1_0_6_n5)
         );
  OR3_X1 npu_inst_pe_1_0_6_U28 ( .A1(npu_inst_pe_1_0_6_n6), .A2(
        npu_inst_pe_1_0_6_n8), .A3(npu_inst_pe_1_0_6_n5), .ZN(
        npu_inst_pe_1_0_6_n56) );
  OR3_X1 npu_inst_pe_1_0_6_U27 ( .A1(npu_inst_pe_1_0_6_n5), .A2(
        npu_inst_pe_1_0_6_n8), .A3(npu_inst_pe_1_0_6_n7), .ZN(
        npu_inst_pe_1_0_6_n48) );
  INV_X1 npu_inst_pe_1_0_6_U26 ( .A(npu_inst_pe_1_0_6_n5), .ZN(
        npu_inst_pe_1_0_6_n4) );
  OR3_X1 npu_inst_pe_1_0_6_U25 ( .A1(npu_inst_pe_1_0_6_n4), .A2(
        npu_inst_pe_1_0_6_n8), .A3(npu_inst_pe_1_0_6_n7), .ZN(
        npu_inst_pe_1_0_6_n52) );
  OR3_X1 npu_inst_pe_1_0_6_U24 ( .A1(npu_inst_pe_1_0_6_n6), .A2(
        npu_inst_pe_1_0_6_n8), .A3(npu_inst_pe_1_0_6_n4), .ZN(
        npu_inst_pe_1_0_6_n60) );
  NOR2_X1 npu_inst_pe_1_0_6_U23 ( .A1(npu_inst_pe_1_0_6_n60), .A2(
        npu_inst_pe_1_0_6_n3), .ZN(npu_inst_pe_1_0_6_n58) );
  NOR2_X1 npu_inst_pe_1_0_6_U22 ( .A1(npu_inst_pe_1_0_6_n56), .A2(
        npu_inst_pe_1_0_6_n3), .ZN(npu_inst_pe_1_0_6_n54) );
  NOR2_X1 npu_inst_pe_1_0_6_U21 ( .A1(npu_inst_pe_1_0_6_n52), .A2(
        npu_inst_pe_1_0_6_n3), .ZN(npu_inst_pe_1_0_6_n50) );
  NOR2_X1 npu_inst_pe_1_0_6_U20 ( .A1(npu_inst_pe_1_0_6_n48), .A2(
        npu_inst_pe_1_0_6_n3), .ZN(npu_inst_pe_1_0_6_n46) );
  NOR2_X1 npu_inst_pe_1_0_6_U19 ( .A1(npu_inst_pe_1_0_6_n40), .A2(
        npu_inst_pe_1_0_6_n3), .ZN(npu_inst_pe_1_0_6_n38) );
  NOR2_X1 npu_inst_pe_1_0_6_U18 ( .A1(npu_inst_pe_1_0_6_n44), .A2(
        npu_inst_pe_1_0_6_n3), .ZN(npu_inst_pe_1_0_6_n42) );
  BUF_X1 npu_inst_pe_1_0_6_U17 ( .A(npu_inst_n106), .Z(npu_inst_pe_1_0_6_n8)
         );
  INV_X1 npu_inst_pe_1_0_6_U16 ( .A(npu_inst_n126), .ZN(npu_inst_pe_1_0_6_n12)
         );
  INV_X1 npu_inst_pe_1_0_6_U15 ( .A(npu_inst_pe_1_0_6_n38), .ZN(
        npu_inst_pe_1_0_6_n114) );
  INV_X1 npu_inst_pe_1_0_6_U14 ( .A(npu_inst_pe_1_0_6_n58), .ZN(
        npu_inst_pe_1_0_6_n119) );
  INV_X1 npu_inst_pe_1_0_6_U13 ( .A(npu_inst_pe_1_0_6_n54), .ZN(
        npu_inst_pe_1_0_6_n118) );
  INV_X1 npu_inst_pe_1_0_6_U12 ( .A(npu_inst_pe_1_0_6_n50), .ZN(
        npu_inst_pe_1_0_6_n117) );
  INV_X1 npu_inst_pe_1_0_6_U11 ( .A(npu_inst_pe_1_0_6_n46), .ZN(
        npu_inst_pe_1_0_6_n116) );
  INV_X1 npu_inst_pe_1_0_6_U10 ( .A(npu_inst_pe_1_0_6_n42), .ZN(
        npu_inst_pe_1_0_6_n115) );
  BUF_X1 npu_inst_pe_1_0_6_U9 ( .A(npu_inst_n35), .Z(npu_inst_pe_1_0_6_n2) );
  BUF_X1 npu_inst_pe_1_0_6_U8 ( .A(npu_inst_n35), .Z(npu_inst_pe_1_0_6_n1) );
  BUF_X1 npu_inst_pe_1_0_6_U7 ( .A(npu_inst_pe_1_0_6_n12), .Z(
        npu_inst_pe_1_0_6_n11) );
  BUF_X1 npu_inst_pe_1_0_6_U6 ( .A(npu_inst_pe_1_0_6_n12), .Z(
        npu_inst_pe_1_0_6_n10) );
  BUF_X1 npu_inst_pe_1_0_6_U5 ( .A(npu_inst_pe_1_0_6_n12), .Z(
        npu_inst_pe_1_0_6_n9) );
  NOR2_X1 npu_inst_pe_1_0_6_U4 ( .A1(npu_inst_pe_1_0_6_int_q_weight_0_), .A2(
        npu_inst_pe_1_0_6_n1), .ZN(npu_inst_pe_1_0_6_n76) );
  NOR2_X1 npu_inst_pe_1_0_6_U3 ( .A1(npu_inst_pe_1_0_6_n27), .A2(
        npu_inst_pe_1_0_6_n1), .ZN(npu_inst_pe_1_0_6_n77) );
  FA_X1 npu_inst_pe_1_0_6_sub_67_U2_1 ( .A(npu_inst_pe_1_0_6_int_q_acc_1_), 
        .B(npu_inst_pe_1_0_6_n14), .CI(npu_inst_pe_1_0_6_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_0_6_sub_67_carry_2_), .S(npu_inst_pe_1_0_6_N66) );
  FA_X1 npu_inst_pe_1_0_6_add_69_U1_1 ( .A(npu_inst_pe_1_0_6_int_q_acc_1_), 
        .B(npu_inst_pe_1_0_6_int_data_1_), .CI(
        npu_inst_pe_1_0_6_add_69_carry_1_), .CO(
        npu_inst_pe_1_0_6_add_69_carry_2_), .S(npu_inst_pe_1_0_6_N74) );
  NAND3_X1 npu_inst_pe_1_0_6_U109 ( .A1(npu_inst_pe_1_0_6_n5), .A2(
        npu_inst_pe_1_0_6_n7), .A3(npu_inst_pe_1_0_6_n8), .ZN(
        npu_inst_pe_1_0_6_n44) );
  NAND3_X1 npu_inst_pe_1_0_6_U108 ( .A1(npu_inst_pe_1_0_6_n4), .A2(
        npu_inst_pe_1_0_6_n7), .A3(npu_inst_pe_1_0_6_n8), .ZN(
        npu_inst_pe_1_0_6_n40) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_0_6_n34), .CK(
        npu_inst_pe_1_0_6_net4424), .RN(npu_inst_pe_1_0_6_n9), .Q(
        npu_inst_pe_1_0_6_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_0_6_n35), .CK(
        npu_inst_pe_1_0_6_net4424), .RN(npu_inst_pe_1_0_6_n9), .Q(
        npu_inst_pe_1_0_6_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_0_6_n36), .CK(
        npu_inst_pe_1_0_6_net4424), .RN(npu_inst_pe_1_0_6_n9), .Q(
        npu_inst_pe_1_0_6_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_0_6_n98), .CK(
        npu_inst_pe_1_0_6_net4424), .RN(npu_inst_pe_1_0_6_n9), .Q(
        npu_inst_pe_1_0_6_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_0_6_n99), .CK(
        npu_inst_pe_1_0_6_net4424), .RN(npu_inst_pe_1_0_6_n9), .Q(
        npu_inst_pe_1_0_6_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_0_6_n100), 
        .CK(npu_inst_pe_1_0_6_net4424), .RN(npu_inst_pe_1_0_6_n9), .Q(
        npu_inst_pe_1_0_6_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_0_6_n33), .CK(
        npu_inst_pe_1_0_6_net4424), .RN(npu_inst_pe_1_0_6_n9), .Q(
        npu_inst_pe_1_0_6_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_0_6_n101), 
        .CK(npu_inst_pe_1_0_6_net4424), .RN(npu_inst_pe_1_0_6_n9), .Q(
        npu_inst_pe_1_0_6_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_weight_reg_0_ ( .D(npu_inst_n112), .CK(
        npu_inst_pe_1_0_6_net4430), .RN(npu_inst_pe_1_0_6_n9), .Q(
        npu_inst_pe_1_0_6_int_q_weight_0_), .QN(npu_inst_pe_1_0_6_n27) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_weight_reg_1_ ( .D(npu_inst_n118), .CK(
        npu_inst_pe_1_0_6_net4430), .RN(npu_inst_pe_1_0_6_n9), .Q(
        npu_inst_pe_1_0_6_int_q_weight_1_), .QN(npu_inst_pe_1_0_6_n26) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_0_6_n113), 
        .CK(npu_inst_pe_1_0_6_net4430), .RN(npu_inst_pe_1_0_6_n9), .Q(
        npu_inst_pe_1_0_6_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_0_6_n107), 
        .CK(npu_inst_pe_1_0_6_net4430), .RN(npu_inst_pe_1_0_6_n9), .Q(
        npu_inst_pe_1_0_6_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_0_6_n112), 
        .CK(npu_inst_pe_1_0_6_net4430), .RN(npu_inst_pe_1_0_6_n10), .Q(
        npu_inst_pe_1_0_6_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_0_6_n106), 
        .CK(npu_inst_pe_1_0_6_net4430), .RN(npu_inst_pe_1_0_6_n10), .Q(
        npu_inst_pe_1_0_6_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_0_6_n111), 
        .CK(npu_inst_pe_1_0_6_net4430), .RN(npu_inst_pe_1_0_6_n10), .Q(
        npu_inst_pe_1_0_6_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_0_6_n105), 
        .CK(npu_inst_pe_1_0_6_net4430), .RN(npu_inst_pe_1_0_6_n10), .Q(
        npu_inst_pe_1_0_6_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_0_6_n110), 
        .CK(npu_inst_pe_1_0_6_net4430), .RN(npu_inst_pe_1_0_6_n10), .Q(
        npu_inst_pe_1_0_6_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_0_6_n104), 
        .CK(npu_inst_pe_1_0_6_net4430), .RN(npu_inst_pe_1_0_6_n10), .Q(
        npu_inst_pe_1_0_6_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_0_6_n109), 
        .CK(npu_inst_pe_1_0_6_net4430), .RN(npu_inst_pe_1_0_6_n10), .Q(
        npu_inst_pe_1_0_6_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_0_6_n103), 
        .CK(npu_inst_pe_1_0_6_net4430), .RN(npu_inst_pe_1_0_6_n10), .Q(
        npu_inst_pe_1_0_6_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_0_6_n108), 
        .CK(npu_inst_pe_1_0_6_net4430), .RN(npu_inst_pe_1_0_6_n10), .Q(
        npu_inst_pe_1_0_6_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_0_6_n102), 
        .CK(npu_inst_pe_1_0_6_net4430), .RN(npu_inst_pe_1_0_6_n10), .Q(
        npu_inst_pe_1_0_6_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_0_6_n86), 
        .CK(npu_inst_pe_1_0_6_net4430), .RN(npu_inst_pe_1_0_6_n10), .Q(
        npu_inst_pe_1_0_6_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_0_6_n87), 
        .CK(npu_inst_pe_1_0_6_net4430), .RN(npu_inst_pe_1_0_6_n10), .Q(
        npu_inst_pe_1_0_6_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_0_6_n88), 
        .CK(npu_inst_pe_1_0_6_net4430), .RN(npu_inst_pe_1_0_6_n11), .Q(
        npu_inst_pe_1_0_6_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_0_6_n89), 
        .CK(npu_inst_pe_1_0_6_net4430), .RN(npu_inst_pe_1_0_6_n11), .Q(
        npu_inst_pe_1_0_6_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_0_6_n90), 
        .CK(npu_inst_pe_1_0_6_net4430), .RN(npu_inst_pe_1_0_6_n11), .Q(
        npu_inst_pe_1_0_6_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_0_6_n91), 
        .CK(npu_inst_pe_1_0_6_net4430), .RN(npu_inst_pe_1_0_6_n11), .Q(
        npu_inst_pe_1_0_6_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_0_6_n92), 
        .CK(npu_inst_pe_1_0_6_net4430), .RN(npu_inst_pe_1_0_6_n11), .Q(
        npu_inst_pe_1_0_6_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_0_6_n93), 
        .CK(npu_inst_pe_1_0_6_net4430), .RN(npu_inst_pe_1_0_6_n11), .Q(
        npu_inst_pe_1_0_6_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_0_6_n94), 
        .CK(npu_inst_pe_1_0_6_net4430), .RN(npu_inst_pe_1_0_6_n11), .Q(
        npu_inst_pe_1_0_6_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_0_6_n95), 
        .CK(npu_inst_pe_1_0_6_net4430), .RN(npu_inst_pe_1_0_6_n11), .Q(
        npu_inst_pe_1_0_6_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_0_6_n96), 
        .CK(npu_inst_pe_1_0_6_net4430), .RN(npu_inst_pe_1_0_6_n11), .Q(
        npu_inst_pe_1_0_6_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_0_6_n97), 
        .CK(npu_inst_pe_1_0_6_net4430), .RN(npu_inst_pe_1_0_6_n11), .Q(
        npu_inst_pe_1_0_6_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_0_6_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_0_6_N84), .SE(1'b0), .GCK(npu_inst_pe_1_0_6_net4424) );
  CLKGATETST_X1 npu_inst_pe_1_0_6_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n66), .SE(1'b0), .GCK(npu_inst_pe_1_0_6_net4430) );
  MUX2_X1 npu_inst_pe_1_0_7_U162 ( .A(npu_inst_pe_1_0_7_n32), .B(
        npu_inst_pe_1_0_7_n29), .S(npu_inst_pe_1_0_7_n8), .Z(
        npu_inst_pe_1_0_7_N93) );
  MUX2_X1 npu_inst_pe_1_0_7_U161 ( .A(npu_inst_pe_1_0_7_n31), .B(
        npu_inst_pe_1_0_7_n30), .S(npu_inst_pe_1_0_7_n6), .Z(
        npu_inst_pe_1_0_7_n32) );
  MUX2_X1 npu_inst_pe_1_0_7_U160 ( .A(npu_inst_pe_1_0_7_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_0_7_int_q_reg_v_1__0_), .S(npu_inst_pe_1_0_7_n4), .Z(
        npu_inst_pe_1_0_7_n31) );
  MUX2_X1 npu_inst_pe_1_0_7_U159 ( .A(npu_inst_pe_1_0_7_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_0_7_int_q_reg_v_3__0_), .S(npu_inst_pe_1_0_7_n4), .Z(
        npu_inst_pe_1_0_7_n30) );
  MUX2_X1 npu_inst_pe_1_0_7_U158 ( .A(npu_inst_pe_1_0_7_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_0_7_int_q_reg_v_5__0_), .S(npu_inst_pe_1_0_7_n4), .Z(
        npu_inst_pe_1_0_7_n29) );
  MUX2_X1 npu_inst_pe_1_0_7_U157 ( .A(npu_inst_pe_1_0_7_n28), .B(
        npu_inst_pe_1_0_7_n23), .S(npu_inst_pe_1_0_7_n8), .Z(
        npu_inst_pe_1_0_7_N94) );
  MUX2_X1 npu_inst_pe_1_0_7_U156 ( .A(npu_inst_pe_1_0_7_n25), .B(
        npu_inst_pe_1_0_7_n24), .S(npu_inst_pe_1_0_7_n6), .Z(
        npu_inst_pe_1_0_7_n28) );
  MUX2_X1 npu_inst_pe_1_0_7_U155 ( .A(npu_inst_pe_1_0_7_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_0_7_int_q_reg_v_1__1_), .S(npu_inst_pe_1_0_7_n4), .Z(
        npu_inst_pe_1_0_7_n25) );
  MUX2_X1 npu_inst_pe_1_0_7_U154 ( .A(npu_inst_pe_1_0_7_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_0_7_int_q_reg_v_3__1_), .S(npu_inst_pe_1_0_7_n4), .Z(
        npu_inst_pe_1_0_7_n24) );
  MUX2_X1 npu_inst_pe_1_0_7_U153 ( .A(npu_inst_pe_1_0_7_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_0_7_int_q_reg_v_5__1_), .S(npu_inst_pe_1_0_7_n4), .Z(
        npu_inst_pe_1_0_7_n23) );
  MUX2_X1 npu_inst_pe_1_0_7_U152 ( .A(npu_inst_pe_1_0_7_n22), .B(
        npu_inst_pe_1_0_7_n19), .S(npu_inst_pe_1_0_7_n8), .Z(
        npu_inst_int_data_x_0__7__1_) );
  MUX2_X1 npu_inst_pe_1_0_7_U151 ( .A(npu_inst_pe_1_0_7_n21), .B(
        npu_inst_pe_1_0_7_n20), .S(npu_inst_pe_1_0_7_n6), .Z(
        npu_inst_pe_1_0_7_n22) );
  MUX2_X1 npu_inst_pe_1_0_7_U150 ( .A(npu_inst_pe_1_0_7_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_0_7_int_q_reg_h_1__1_), .S(npu_inst_pe_1_0_7_n4), .Z(
        npu_inst_pe_1_0_7_n21) );
  MUX2_X1 npu_inst_pe_1_0_7_U149 ( .A(npu_inst_pe_1_0_7_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_0_7_int_q_reg_h_3__1_), .S(npu_inst_pe_1_0_7_n4), .Z(
        npu_inst_pe_1_0_7_n20) );
  MUX2_X1 npu_inst_pe_1_0_7_U148 ( .A(npu_inst_pe_1_0_7_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_0_7_int_q_reg_h_5__1_), .S(npu_inst_pe_1_0_7_n4), .Z(
        npu_inst_pe_1_0_7_n19) );
  MUX2_X1 npu_inst_pe_1_0_7_U147 ( .A(npu_inst_pe_1_0_7_n18), .B(
        npu_inst_pe_1_0_7_n15), .S(npu_inst_pe_1_0_7_n8), .Z(
        npu_inst_int_data_x_0__7__0_) );
  MUX2_X1 npu_inst_pe_1_0_7_U146 ( .A(npu_inst_pe_1_0_7_n17), .B(
        npu_inst_pe_1_0_7_n16), .S(npu_inst_pe_1_0_7_n6), .Z(
        npu_inst_pe_1_0_7_n18) );
  MUX2_X1 npu_inst_pe_1_0_7_U145 ( .A(npu_inst_pe_1_0_7_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_0_7_int_q_reg_h_1__0_), .S(npu_inst_pe_1_0_7_n4), .Z(
        npu_inst_pe_1_0_7_n17) );
  MUX2_X1 npu_inst_pe_1_0_7_U144 ( .A(npu_inst_pe_1_0_7_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_0_7_int_q_reg_h_3__0_), .S(npu_inst_pe_1_0_7_n4), .Z(
        npu_inst_pe_1_0_7_n16) );
  MUX2_X1 npu_inst_pe_1_0_7_U143 ( .A(npu_inst_pe_1_0_7_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_0_7_int_q_reg_h_5__0_), .S(npu_inst_pe_1_0_7_n4), .Z(
        npu_inst_pe_1_0_7_n15) );
  XOR2_X1 npu_inst_pe_1_0_7_U142 ( .A(npu_inst_pe_1_0_7_int_data_0_), .B(
        npu_inst_pe_1_0_7_int_q_acc_0_), .Z(npu_inst_pe_1_0_7_N73) );
  AND2_X1 npu_inst_pe_1_0_7_U141 ( .A1(npu_inst_pe_1_0_7_int_q_acc_0_), .A2(
        npu_inst_pe_1_0_7_int_data_0_), .ZN(npu_inst_pe_1_0_7_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_0_7_U140 ( .A(npu_inst_pe_1_0_7_int_q_acc_0_), .B(
        npu_inst_pe_1_0_7_n13), .ZN(npu_inst_pe_1_0_7_N65) );
  OR2_X1 npu_inst_pe_1_0_7_U139 ( .A1(npu_inst_pe_1_0_7_n13), .A2(
        npu_inst_pe_1_0_7_int_q_acc_0_), .ZN(npu_inst_pe_1_0_7_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_0_7_U138 ( .A(npu_inst_pe_1_0_7_int_q_acc_2_), .B(
        npu_inst_pe_1_0_7_add_69_carry_2_), .Z(npu_inst_pe_1_0_7_N75) );
  AND2_X1 npu_inst_pe_1_0_7_U137 ( .A1(npu_inst_pe_1_0_7_add_69_carry_2_), 
        .A2(npu_inst_pe_1_0_7_int_q_acc_2_), .ZN(
        npu_inst_pe_1_0_7_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_0_7_U136 ( .A(npu_inst_pe_1_0_7_int_q_acc_3_), .B(
        npu_inst_pe_1_0_7_add_69_carry_3_), .Z(npu_inst_pe_1_0_7_N76) );
  AND2_X1 npu_inst_pe_1_0_7_U135 ( .A1(npu_inst_pe_1_0_7_add_69_carry_3_), 
        .A2(npu_inst_pe_1_0_7_int_q_acc_3_), .ZN(
        npu_inst_pe_1_0_7_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_0_7_U134 ( .A(npu_inst_pe_1_0_7_int_q_acc_4_), .B(
        npu_inst_pe_1_0_7_add_69_carry_4_), .Z(npu_inst_pe_1_0_7_N77) );
  AND2_X1 npu_inst_pe_1_0_7_U133 ( .A1(npu_inst_pe_1_0_7_add_69_carry_4_), 
        .A2(npu_inst_pe_1_0_7_int_q_acc_4_), .ZN(
        npu_inst_pe_1_0_7_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_0_7_U132 ( .A(npu_inst_pe_1_0_7_int_q_acc_5_), .B(
        npu_inst_pe_1_0_7_add_69_carry_5_), .Z(npu_inst_pe_1_0_7_N78) );
  AND2_X1 npu_inst_pe_1_0_7_U131 ( .A1(npu_inst_pe_1_0_7_add_69_carry_5_), 
        .A2(npu_inst_pe_1_0_7_int_q_acc_5_), .ZN(
        npu_inst_pe_1_0_7_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_0_7_U130 ( .A(npu_inst_pe_1_0_7_int_q_acc_6_), .B(
        npu_inst_pe_1_0_7_add_69_carry_6_), .Z(npu_inst_pe_1_0_7_N79) );
  AND2_X1 npu_inst_pe_1_0_7_U129 ( .A1(npu_inst_pe_1_0_7_add_69_carry_6_), 
        .A2(npu_inst_pe_1_0_7_int_q_acc_6_), .ZN(
        npu_inst_pe_1_0_7_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_0_7_U128 ( .A(npu_inst_pe_1_0_7_int_q_acc_7_), .B(
        npu_inst_pe_1_0_7_add_69_carry_7_), .Z(npu_inst_pe_1_0_7_N80) );
  XNOR2_X1 npu_inst_pe_1_0_7_U127 ( .A(npu_inst_pe_1_0_7_sub_67_carry_2_), .B(
        npu_inst_pe_1_0_7_int_q_acc_2_), .ZN(npu_inst_pe_1_0_7_N67) );
  OR2_X1 npu_inst_pe_1_0_7_U126 ( .A1(npu_inst_pe_1_0_7_int_q_acc_2_), .A2(
        npu_inst_pe_1_0_7_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_0_7_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_0_7_U125 ( .A(npu_inst_pe_1_0_7_sub_67_carry_3_), .B(
        npu_inst_pe_1_0_7_int_q_acc_3_), .ZN(npu_inst_pe_1_0_7_N68) );
  OR2_X1 npu_inst_pe_1_0_7_U124 ( .A1(npu_inst_pe_1_0_7_int_q_acc_3_), .A2(
        npu_inst_pe_1_0_7_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_0_7_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_0_7_U123 ( .A(npu_inst_pe_1_0_7_sub_67_carry_4_), .B(
        npu_inst_pe_1_0_7_int_q_acc_4_), .ZN(npu_inst_pe_1_0_7_N69) );
  OR2_X1 npu_inst_pe_1_0_7_U122 ( .A1(npu_inst_pe_1_0_7_int_q_acc_4_), .A2(
        npu_inst_pe_1_0_7_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_0_7_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_0_7_U121 ( .A(npu_inst_pe_1_0_7_sub_67_carry_5_), .B(
        npu_inst_pe_1_0_7_int_q_acc_5_), .ZN(npu_inst_pe_1_0_7_N70) );
  OR2_X1 npu_inst_pe_1_0_7_U120 ( .A1(npu_inst_pe_1_0_7_int_q_acc_5_), .A2(
        npu_inst_pe_1_0_7_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_0_7_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_0_7_U119 ( .A(npu_inst_pe_1_0_7_sub_67_carry_6_), .B(
        npu_inst_pe_1_0_7_int_q_acc_6_), .ZN(npu_inst_pe_1_0_7_N71) );
  OR2_X1 npu_inst_pe_1_0_7_U118 ( .A1(npu_inst_pe_1_0_7_int_q_acc_6_), .A2(
        npu_inst_pe_1_0_7_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_0_7_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_0_7_U117 ( .A(npu_inst_pe_1_0_7_int_q_acc_7_), .B(
        npu_inst_pe_1_0_7_sub_67_carry_7_), .ZN(npu_inst_pe_1_0_7_N72) );
  INV_X1 npu_inst_pe_1_0_7_U116 ( .A(npu_inst_n79), .ZN(npu_inst_pe_1_0_7_n7)
         );
  INV_X1 npu_inst_pe_1_0_7_U115 ( .A(npu_inst_pe_1_0_7_n7), .ZN(
        npu_inst_pe_1_0_7_n6) );
  INV_X1 npu_inst_pe_1_0_7_U114 ( .A(npu_inst_n60), .ZN(npu_inst_pe_1_0_7_n3)
         );
  AOI22_X1 npu_inst_pe_1_0_7_U113 ( .A1(npu_inst_int_data_y_1__7__0_), .A2(
        npu_inst_pe_1_0_7_n58), .B1(npu_inst_pe_1_0_7_n119), .B2(
        npu_inst_pe_1_0_7_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_0_7_n57) );
  INV_X1 npu_inst_pe_1_0_7_U112 ( .A(npu_inst_pe_1_0_7_n57), .ZN(
        npu_inst_pe_1_0_7_n108) );
  AOI22_X1 npu_inst_pe_1_0_7_U111 ( .A1(npu_inst_int_data_y_1__7__0_), .A2(
        npu_inst_pe_1_0_7_n54), .B1(npu_inst_pe_1_0_7_n118), .B2(
        npu_inst_pe_1_0_7_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_0_7_n53) );
  INV_X1 npu_inst_pe_1_0_7_U110 ( .A(npu_inst_pe_1_0_7_n53), .ZN(
        npu_inst_pe_1_0_7_n109) );
  AOI22_X1 npu_inst_pe_1_0_7_U107 ( .A1(npu_inst_int_data_y_1__7__0_), .A2(
        npu_inst_pe_1_0_7_n50), .B1(npu_inst_pe_1_0_7_n117), .B2(
        npu_inst_pe_1_0_7_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_0_7_n49) );
  INV_X1 npu_inst_pe_1_0_7_U106 ( .A(npu_inst_pe_1_0_7_n49), .ZN(
        npu_inst_pe_1_0_7_n110) );
  AOI22_X1 npu_inst_pe_1_0_7_U105 ( .A1(npu_inst_int_data_y_1__7__0_), .A2(
        npu_inst_pe_1_0_7_n46), .B1(npu_inst_pe_1_0_7_n116), .B2(
        npu_inst_pe_1_0_7_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_0_7_n45) );
  INV_X1 npu_inst_pe_1_0_7_U104 ( .A(npu_inst_pe_1_0_7_n45), .ZN(
        npu_inst_pe_1_0_7_n111) );
  AOI22_X1 npu_inst_pe_1_0_7_U103 ( .A1(npu_inst_int_data_y_1__7__0_), .A2(
        npu_inst_pe_1_0_7_n42), .B1(npu_inst_pe_1_0_7_n115), .B2(
        npu_inst_pe_1_0_7_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_0_7_n41) );
  INV_X1 npu_inst_pe_1_0_7_U102 ( .A(npu_inst_pe_1_0_7_n41), .ZN(
        npu_inst_pe_1_0_7_n112) );
  AOI22_X1 npu_inst_pe_1_0_7_U101 ( .A1(npu_inst_int_data_y_1__7__1_), .A2(
        npu_inst_pe_1_0_7_n58), .B1(npu_inst_pe_1_0_7_n119), .B2(
        npu_inst_pe_1_0_7_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_0_7_n59) );
  INV_X1 npu_inst_pe_1_0_7_U100 ( .A(npu_inst_pe_1_0_7_n59), .ZN(
        npu_inst_pe_1_0_7_n102) );
  AOI22_X1 npu_inst_pe_1_0_7_U99 ( .A1(npu_inst_int_data_y_1__7__1_), .A2(
        npu_inst_pe_1_0_7_n54), .B1(npu_inst_pe_1_0_7_n118), .B2(
        npu_inst_pe_1_0_7_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_0_7_n55) );
  INV_X1 npu_inst_pe_1_0_7_U98 ( .A(npu_inst_pe_1_0_7_n55), .ZN(
        npu_inst_pe_1_0_7_n103) );
  AOI22_X1 npu_inst_pe_1_0_7_U97 ( .A1(npu_inst_int_data_y_1__7__1_), .A2(
        npu_inst_pe_1_0_7_n50), .B1(npu_inst_pe_1_0_7_n117), .B2(
        npu_inst_pe_1_0_7_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_0_7_n51) );
  INV_X1 npu_inst_pe_1_0_7_U96 ( .A(npu_inst_pe_1_0_7_n51), .ZN(
        npu_inst_pe_1_0_7_n104) );
  AOI22_X1 npu_inst_pe_1_0_7_U95 ( .A1(npu_inst_int_data_y_1__7__1_), .A2(
        npu_inst_pe_1_0_7_n46), .B1(npu_inst_pe_1_0_7_n116), .B2(
        npu_inst_pe_1_0_7_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_0_7_n47) );
  INV_X1 npu_inst_pe_1_0_7_U94 ( .A(npu_inst_pe_1_0_7_n47), .ZN(
        npu_inst_pe_1_0_7_n105) );
  AOI22_X1 npu_inst_pe_1_0_7_U93 ( .A1(npu_inst_int_data_y_1__7__1_), .A2(
        npu_inst_pe_1_0_7_n42), .B1(npu_inst_pe_1_0_7_n115), .B2(
        npu_inst_pe_1_0_7_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_0_7_n43) );
  INV_X1 npu_inst_pe_1_0_7_U92 ( .A(npu_inst_pe_1_0_7_n43), .ZN(
        npu_inst_pe_1_0_7_n106) );
  AOI22_X1 npu_inst_pe_1_0_7_U91 ( .A1(npu_inst_pe_1_0_7_n38), .A2(
        npu_inst_int_data_y_1__7__1_), .B1(npu_inst_pe_1_0_7_n114), .B2(
        npu_inst_pe_1_0_7_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_0_7_n39) );
  INV_X1 npu_inst_pe_1_0_7_U90 ( .A(npu_inst_pe_1_0_7_n39), .ZN(
        npu_inst_pe_1_0_7_n107) );
  AOI22_X1 npu_inst_pe_1_0_7_U89 ( .A1(npu_inst_pe_1_0_7_n38), .A2(
        npu_inst_int_data_y_1__7__0_), .B1(npu_inst_pe_1_0_7_n114), .B2(
        npu_inst_pe_1_0_7_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_0_7_n37) );
  INV_X1 npu_inst_pe_1_0_7_U88 ( .A(npu_inst_pe_1_0_7_n37), .ZN(
        npu_inst_pe_1_0_7_n113) );
  AND2_X1 npu_inst_pe_1_0_7_U87 ( .A1(npu_inst_pe_1_0_7_int_q_acc_2_), .A2(
        npu_inst_pe_1_0_7_n1), .ZN(int_o_data_npu[2]) );
  AND2_X1 npu_inst_pe_1_0_7_U86 ( .A1(npu_inst_pe_1_0_7_int_q_acc_3_), .A2(
        npu_inst_pe_1_0_7_n2), .ZN(int_o_data_npu[3]) );
  NOR3_X1 npu_inst_pe_1_0_7_U85 ( .A1(npu_inst_pe_1_0_7_n26), .A2(npu_inst_n60), .A3(npu_inst_int_ckg[56]), .ZN(npu_inst_pe_1_0_7_n85) );
  OR2_X1 npu_inst_pe_1_0_7_U84 ( .A1(npu_inst_pe_1_0_7_n85), .A2(
        npu_inst_pe_1_0_7_n2), .ZN(npu_inst_pe_1_0_7_N84) );
  AND2_X1 npu_inst_pe_1_0_7_U83 ( .A1(npu_inst_pe_1_0_7_int_q_acc_6_), .A2(
        npu_inst_pe_1_0_7_n2), .ZN(int_o_data_npu[6]) );
  AND2_X1 npu_inst_pe_1_0_7_U82 ( .A1(npu_inst_pe_1_0_7_int_q_acc_5_), .A2(
        npu_inst_pe_1_0_7_n2), .ZN(int_o_data_npu[5]) );
  AND2_X1 npu_inst_pe_1_0_7_U81 ( .A1(npu_inst_pe_1_0_7_int_q_acc_4_), .A2(
        npu_inst_pe_1_0_7_n2), .ZN(int_o_data_npu[4]) );
  AOI222_X1 npu_inst_pe_1_0_7_U80 ( .A1(npu_inst_int_data_res_1__7__0_), .A2(
        npu_inst_pe_1_0_7_n1), .B1(npu_inst_pe_1_0_7_N73), .B2(
        npu_inst_pe_1_0_7_n76), .C1(npu_inst_pe_1_0_7_N65), .C2(
        npu_inst_pe_1_0_7_n77), .ZN(npu_inst_pe_1_0_7_n84) );
  INV_X1 npu_inst_pe_1_0_7_U79 ( .A(npu_inst_pe_1_0_7_n84), .ZN(
        npu_inst_pe_1_0_7_n101) );
  AOI222_X1 npu_inst_pe_1_0_7_U78 ( .A1(npu_inst_int_data_res_1__7__7_), .A2(
        npu_inst_pe_1_0_7_n1), .B1(npu_inst_pe_1_0_7_N80), .B2(
        npu_inst_pe_1_0_7_n76), .C1(npu_inst_pe_1_0_7_N72), .C2(
        npu_inst_pe_1_0_7_n77), .ZN(npu_inst_pe_1_0_7_n75) );
  INV_X1 npu_inst_pe_1_0_7_U77 ( .A(npu_inst_pe_1_0_7_n75), .ZN(
        npu_inst_pe_1_0_7_n33) );
  AOI222_X1 npu_inst_pe_1_0_7_U76 ( .A1(npu_inst_int_data_res_1__7__1_), .A2(
        npu_inst_pe_1_0_7_n1), .B1(npu_inst_pe_1_0_7_N74), .B2(
        npu_inst_pe_1_0_7_n76), .C1(npu_inst_pe_1_0_7_N66), .C2(
        npu_inst_pe_1_0_7_n77), .ZN(npu_inst_pe_1_0_7_n83) );
  INV_X1 npu_inst_pe_1_0_7_U75 ( .A(npu_inst_pe_1_0_7_n83), .ZN(
        npu_inst_pe_1_0_7_n100) );
  AOI222_X1 npu_inst_pe_1_0_7_U74 ( .A1(npu_inst_int_data_res_1__7__2_), .A2(
        npu_inst_pe_1_0_7_n1), .B1(npu_inst_pe_1_0_7_N75), .B2(
        npu_inst_pe_1_0_7_n76), .C1(npu_inst_pe_1_0_7_N67), .C2(
        npu_inst_pe_1_0_7_n77), .ZN(npu_inst_pe_1_0_7_n82) );
  INV_X1 npu_inst_pe_1_0_7_U73 ( .A(npu_inst_pe_1_0_7_n82), .ZN(
        npu_inst_pe_1_0_7_n99) );
  AOI222_X1 npu_inst_pe_1_0_7_U72 ( .A1(npu_inst_int_data_res_1__7__3_), .A2(
        npu_inst_pe_1_0_7_n1), .B1(npu_inst_pe_1_0_7_N76), .B2(
        npu_inst_pe_1_0_7_n76), .C1(npu_inst_pe_1_0_7_N68), .C2(
        npu_inst_pe_1_0_7_n77), .ZN(npu_inst_pe_1_0_7_n81) );
  INV_X1 npu_inst_pe_1_0_7_U71 ( .A(npu_inst_pe_1_0_7_n81), .ZN(
        npu_inst_pe_1_0_7_n98) );
  AOI222_X1 npu_inst_pe_1_0_7_U70 ( .A1(npu_inst_int_data_res_1__7__4_), .A2(
        npu_inst_pe_1_0_7_n1), .B1(npu_inst_pe_1_0_7_N77), .B2(
        npu_inst_pe_1_0_7_n76), .C1(npu_inst_pe_1_0_7_N69), .C2(
        npu_inst_pe_1_0_7_n77), .ZN(npu_inst_pe_1_0_7_n80) );
  INV_X1 npu_inst_pe_1_0_7_U69 ( .A(npu_inst_pe_1_0_7_n80), .ZN(
        npu_inst_pe_1_0_7_n36) );
  AOI222_X1 npu_inst_pe_1_0_7_U68 ( .A1(npu_inst_int_data_res_1__7__5_), .A2(
        npu_inst_pe_1_0_7_n1), .B1(npu_inst_pe_1_0_7_N78), .B2(
        npu_inst_pe_1_0_7_n76), .C1(npu_inst_pe_1_0_7_N70), .C2(
        npu_inst_pe_1_0_7_n77), .ZN(npu_inst_pe_1_0_7_n79) );
  INV_X1 npu_inst_pe_1_0_7_U67 ( .A(npu_inst_pe_1_0_7_n79), .ZN(
        npu_inst_pe_1_0_7_n35) );
  AOI222_X1 npu_inst_pe_1_0_7_U66 ( .A1(npu_inst_int_data_res_1__7__6_), .A2(
        npu_inst_pe_1_0_7_n1), .B1(npu_inst_pe_1_0_7_N79), .B2(
        npu_inst_pe_1_0_7_n76), .C1(npu_inst_pe_1_0_7_N71), .C2(
        npu_inst_pe_1_0_7_n77), .ZN(npu_inst_pe_1_0_7_n78) );
  INV_X1 npu_inst_pe_1_0_7_U65 ( .A(npu_inst_pe_1_0_7_n78), .ZN(
        npu_inst_pe_1_0_7_n34) );
  INV_X1 npu_inst_pe_1_0_7_U64 ( .A(npu_inst_pe_1_0_7_int_data_1_), .ZN(
        npu_inst_pe_1_0_7_n14) );
  AND2_X1 npu_inst_pe_1_0_7_U63 ( .A1(npu_inst_int_data_x_0__7__1_), .A2(
        npu_inst_pe_1_0_7_int_q_weight_1_), .ZN(npu_inst_pe_1_0_7_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_0_7_U62 ( .A1(npu_inst_int_data_x_0__7__0_), .A2(
        npu_inst_pe_1_0_7_int_q_weight_1_), .ZN(npu_inst_pe_1_0_7_int_data_0_)
         );
  AND2_X1 npu_inst_pe_1_0_7_U61 ( .A1(npu_inst_pe_1_0_7_n2), .A2(
        npu_inst_pe_1_0_7_int_q_acc_7_), .ZN(int_o_data_npu[7]) );
  NAND2_X1 npu_inst_pe_1_0_7_U60 ( .A1(npu_inst_pe_1_0_7_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_0_7_n60), .ZN(npu_inst_pe_1_0_7_n74) );
  OAI21_X1 npu_inst_pe_1_0_7_U59 ( .B1(npu_inst_pe_1_0_7_n63), .B2(
        npu_inst_pe_1_0_7_n60), .A(npu_inst_pe_1_0_7_n74), .ZN(
        npu_inst_pe_1_0_7_n97) );
  NAND2_X1 npu_inst_pe_1_0_7_U58 ( .A1(npu_inst_pe_1_0_7_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_0_7_n60), .ZN(npu_inst_pe_1_0_7_n73) );
  OAI21_X1 npu_inst_pe_1_0_7_U57 ( .B1(npu_inst_pe_1_0_7_n61), .B2(
        npu_inst_pe_1_0_7_n60), .A(npu_inst_pe_1_0_7_n73), .ZN(
        npu_inst_pe_1_0_7_n96) );
  NAND2_X1 npu_inst_pe_1_0_7_U56 ( .A1(npu_inst_pe_1_0_7_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_0_7_n56), .ZN(npu_inst_pe_1_0_7_n72) );
  OAI21_X1 npu_inst_pe_1_0_7_U55 ( .B1(npu_inst_pe_1_0_7_n63), .B2(
        npu_inst_pe_1_0_7_n56), .A(npu_inst_pe_1_0_7_n72), .ZN(
        npu_inst_pe_1_0_7_n95) );
  NAND2_X1 npu_inst_pe_1_0_7_U54 ( .A1(npu_inst_pe_1_0_7_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_0_7_n56), .ZN(npu_inst_pe_1_0_7_n71) );
  OAI21_X1 npu_inst_pe_1_0_7_U53 ( .B1(npu_inst_pe_1_0_7_n61), .B2(
        npu_inst_pe_1_0_7_n56), .A(npu_inst_pe_1_0_7_n71), .ZN(
        npu_inst_pe_1_0_7_n94) );
  NAND2_X1 npu_inst_pe_1_0_7_U52 ( .A1(npu_inst_pe_1_0_7_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_0_7_n52), .ZN(npu_inst_pe_1_0_7_n70) );
  OAI21_X1 npu_inst_pe_1_0_7_U51 ( .B1(npu_inst_pe_1_0_7_n63), .B2(
        npu_inst_pe_1_0_7_n52), .A(npu_inst_pe_1_0_7_n70), .ZN(
        npu_inst_pe_1_0_7_n93) );
  NAND2_X1 npu_inst_pe_1_0_7_U50 ( .A1(npu_inst_pe_1_0_7_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_0_7_n52), .ZN(npu_inst_pe_1_0_7_n69) );
  OAI21_X1 npu_inst_pe_1_0_7_U49 ( .B1(npu_inst_pe_1_0_7_n61), .B2(
        npu_inst_pe_1_0_7_n52), .A(npu_inst_pe_1_0_7_n69), .ZN(
        npu_inst_pe_1_0_7_n92) );
  NAND2_X1 npu_inst_pe_1_0_7_U48 ( .A1(npu_inst_pe_1_0_7_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_0_7_n48), .ZN(npu_inst_pe_1_0_7_n68) );
  OAI21_X1 npu_inst_pe_1_0_7_U47 ( .B1(npu_inst_pe_1_0_7_n63), .B2(
        npu_inst_pe_1_0_7_n48), .A(npu_inst_pe_1_0_7_n68), .ZN(
        npu_inst_pe_1_0_7_n91) );
  NAND2_X1 npu_inst_pe_1_0_7_U46 ( .A1(npu_inst_pe_1_0_7_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_0_7_n48), .ZN(npu_inst_pe_1_0_7_n67) );
  OAI21_X1 npu_inst_pe_1_0_7_U45 ( .B1(npu_inst_pe_1_0_7_n61), .B2(
        npu_inst_pe_1_0_7_n48), .A(npu_inst_pe_1_0_7_n67), .ZN(
        npu_inst_pe_1_0_7_n90) );
  NAND2_X1 npu_inst_pe_1_0_7_U44 ( .A1(npu_inst_pe_1_0_7_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_0_7_n44), .ZN(npu_inst_pe_1_0_7_n66) );
  OAI21_X1 npu_inst_pe_1_0_7_U43 ( .B1(npu_inst_pe_1_0_7_n63), .B2(
        npu_inst_pe_1_0_7_n44), .A(npu_inst_pe_1_0_7_n66), .ZN(
        npu_inst_pe_1_0_7_n89) );
  NAND2_X1 npu_inst_pe_1_0_7_U42 ( .A1(npu_inst_pe_1_0_7_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_0_7_n44), .ZN(npu_inst_pe_1_0_7_n65) );
  OAI21_X1 npu_inst_pe_1_0_7_U41 ( .B1(npu_inst_pe_1_0_7_n61), .B2(
        npu_inst_pe_1_0_7_n44), .A(npu_inst_pe_1_0_7_n65), .ZN(
        npu_inst_pe_1_0_7_n88) );
  NAND2_X1 npu_inst_pe_1_0_7_U40 ( .A1(npu_inst_pe_1_0_7_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_0_7_n40), .ZN(npu_inst_pe_1_0_7_n64) );
  OAI21_X1 npu_inst_pe_1_0_7_U39 ( .B1(npu_inst_pe_1_0_7_n63), .B2(
        npu_inst_pe_1_0_7_n40), .A(npu_inst_pe_1_0_7_n64), .ZN(
        npu_inst_pe_1_0_7_n87) );
  NAND2_X1 npu_inst_pe_1_0_7_U38 ( .A1(npu_inst_pe_1_0_7_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_0_7_n40), .ZN(npu_inst_pe_1_0_7_n62) );
  OAI21_X1 npu_inst_pe_1_0_7_U37 ( .B1(npu_inst_pe_1_0_7_n61), .B2(
        npu_inst_pe_1_0_7_n40), .A(npu_inst_pe_1_0_7_n62), .ZN(
        npu_inst_pe_1_0_7_n86) );
  AND2_X1 npu_inst_pe_1_0_7_U36 ( .A1(npu_inst_pe_1_0_7_int_q_acc_1_), .A2(
        npu_inst_pe_1_0_7_n1), .ZN(int_o_data_npu[1]) );
  AND2_X1 npu_inst_pe_1_0_7_U35 ( .A1(npu_inst_pe_1_0_7_int_q_acc_0_), .A2(
        npu_inst_pe_1_0_7_n1), .ZN(int_o_data_npu[0]) );
  AND2_X1 npu_inst_pe_1_0_7_U34 ( .A1(npu_inst_pe_1_0_7_N93), .A2(npu_inst_n60), .ZN(npu_inst_pe_1_0_7_o_data_v_0_) );
  AND2_X1 npu_inst_pe_1_0_7_U33 ( .A1(npu_inst_n60), .A2(npu_inst_pe_1_0_7_N94), .ZN(npu_inst_pe_1_0_7_o_data_v_1_) );
  INV_X1 npu_inst_pe_1_0_7_U32 ( .A(npu_inst_pe_1_0_7_int_data_0_), .ZN(
        npu_inst_pe_1_0_7_n13) );
  INV_X1 npu_inst_pe_1_0_7_U31 ( .A(npu_inst_n71), .ZN(npu_inst_pe_1_0_7_n5)
         );
  AOI22_X1 npu_inst_pe_1_0_7_U30 ( .A1(npu_inst_n60), .A2(
        npu_inst_int_data_y_1__7__1_), .B1(npu_inst_pe_1_0_7_n3), .B2(
        int_i_data_h_npu[15]), .ZN(npu_inst_pe_1_0_7_n63) );
  AOI22_X1 npu_inst_pe_1_0_7_U29 ( .A1(npu_inst_n60), .A2(
        npu_inst_int_data_y_1__7__0_), .B1(npu_inst_pe_1_0_7_n3), .B2(
        int_i_data_h_npu[14]), .ZN(npu_inst_pe_1_0_7_n61) );
  OR3_X1 npu_inst_pe_1_0_7_U28 ( .A1(npu_inst_pe_1_0_7_n6), .A2(
        npu_inst_pe_1_0_7_n8), .A3(npu_inst_pe_1_0_7_n5), .ZN(
        npu_inst_pe_1_0_7_n56) );
  OR3_X1 npu_inst_pe_1_0_7_U27 ( .A1(npu_inst_pe_1_0_7_n5), .A2(
        npu_inst_pe_1_0_7_n8), .A3(npu_inst_pe_1_0_7_n7), .ZN(
        npu_inst_pe_1_0_7_n48) );
  INV_X1 npu_inst_pe_1_0_7_U26 ( .A(npu_inst_pe_1_0_7_n5), .ZN(
        npu_inst_pe_1_0_7_n4) );
  OR3_X1 npu_inst_pe_1_0_7_U25 ( .A1(npu_inst_pe_1_0_7_n4), .A2(
        npu_inst_pe_1_0_7_n8), .A3(npu_inst_pe_1_0_7_n7), .ZN(
        npu_inst_pe_1_0_7_n52) );
  OR3_X1 npu_inst_pe_1_0_7_U24 ( .A1(npu_inst_pe_1_0_7_n6), .A2(
        npu_inst_pe_1_0_7_n8), .A3(npu_inst_pe_1_0_7_n4), .ZN(
        npu_inst_pe_1_0_7_n60) );
  NOR2_X1 npu_inst_pe_1_0_7_U23 ( .A1(npu_inst_pe_1_0_7_n60), .A2(
        npu_inst_pe_1_0_7_n3), .ZN(npu_inst_pe_1_0_7_n58) );
  NOR2_X1 npu_inst_pe_1_0_7_U22 ( .A1(npu_inst_pe_1_0_7_n56), .A2(
        npu_inst_pe_1_0_7_n3), .ZN(npu_inst_pe_1_0_7_n54) );
  NOR2_X1 npu_inst_pe_1_0_7_U21 ( .A1(npu_inst_pe_1_0_7_n52), .A2(
        npu_inst_pe_1_0_7_n3), .ZN(npu_inst_pe_1_0_7_n50) );
  NOR2_X1 npu_inst_pe_1_0_7_U20 ( .A1(npu_inst_pe_1_0_7_n48), .A2(
        npu_inst_pe_1_0_7_n3), .ZN(npu_inst_pe_1_0_7_n46) );
  NOR2_X1 npu_inst_pe_1_0_7_U19 ( .A1(npu_inst_pe_1_0_7_n40), .A2(
        npu_inst_pe_1_0_7_n3), .ZN(npu_inst_pe_1_0_7_n38) );
  NOR2_X1 npu_inst_pe_1_0_7_U18 ( .A1(npu_inst_pe_1_0_7_n44), .A2(
        npu_inst_pe_1_0_7_n3), .ZN(npu_inst_pe_1_0_7_n42) );
  BUF_X1 npu_inst_pe_1_0_7_U17 ( .A(npu_inst_n106), .Z(npu_inst_pe_1_0_7_n8)
         );
  INV_X1 npu_inst_pe_1_0_7_U16 ( .A(npu_inst_n126), .ZN(npu_inst_pe_1_0_7_n12)
         );
  INV_X1 npu_inst_pe_1_0_7_U15 ( .A(npu_inst_pe_1_0_7_n38), .ZN(
        npu_inst_pe_1_0_7_n114) );
  INV_X1 npu_inst_pe_1_0_7_U14 ( .A(npu_inst_pe_1_0_7_n58), .ZN(
        npu_inst_pe_1_0_7_n119) );
  INV_X1 npu_inst_pe_1_0_7_U13 ( .A(npu_inst_pe_1_0_7_n54), .ZN(
        npu_inst_pe_1_0_7_n118) );
  INV_X1 npu_inst_pe_1_0_7_U12 ( .A(npu_inst_pe_1_0_7_n50), .ZN(
        npu_inst_pe_1_0_7_n117) );
  INV_X1 npu_inst_pe_1_0_7_U11 ( .A(npu_inst_pe_1_0_7_n46), .ZN(
        npu_inst_pe_1_0_7_n116) );
  INV_X1 npu_inst_pe_1_0_7_U10 ( .A(npu_inst_pe_1_0_7_n42), .ZN(
        npu_inst_pe_1_0_7_n115) );
  BUF_X1 npu_inst_pe_1_0_7_U9 ( .A(npu_inst_n35), .Z(npu_inst_pe_1_0_7_n2) );
  BUF_X1 npu_inst_pe_1_0_7_U8 ( .A(npu_inst_n35), .Z(npu_inst_pe_1_0_7_n1) );
  BUF_X1 npu_inst_pe_1_0_7_U7 ( .A(npu_inst_pe_1_0_7_n12), .Z(
        npu_inst_pe_1_0_7_n11) );
  BUF_X1 npu_inst_pe_1_0_7_U6 ( .A(npu_inst_pe_1_0_7_n12), .Z(
        npu_inst_pe_1_0_7_n10) );
  BUF_X1 npu_inst_pe_1_0_7_U5 ( .A(npu_inst_pe_1_0_7_n12), .Z(
        npu_inst_pe_1_0_7_n9) );
  NOR2_X1 npu_inst_pe_1_0_7_U4 ( .A1(npu_inst_pe_1_0_7_int_q_weight_0_), .A2(
        npu_inst_pe_1_0_7_n1), .ZN(npu_inst_pe_1_0_7_n76) );
  NOR2_X1 npu_inst_pe_1_0_7_U3 ( .A1(npu_inst_pe_1_0_7_n27), .A2(
        npu_inst_pe_1_0_7_n1), .ZN(npu_inst_pe_1_0_7_n77) );
  FA_X1 npu_inst_pe_1_0_7_sub_67_U2_1 ( .A(npu_inst_pe_1_0_7_int_q_acc_1_), 
        .B(npu_inst_pe_1_0_7_n14), .CI(npu_inst_pe_1_0_7_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_0_7_sub_67_carry_2_), .S(npu_inst_pe_1_0_7_N66) );
  FA_X1 npu_inst_pe_1_0_7_add_69_U1_1 ( .A(npu_inst_pe_1_0_7_int_q_acc_1_), 
        .B(npu_inst_pe_1_0_7_int_data_1_), .CI(
        npu_inst_pe_1_0_7_add_69_carry_1_), .CO(
        npu_inst_pe_1_0_7_add_69_carry_2_), .S(npu_inst_pe_1_0_7_N74) );
  NAND3_X1 npu_inst_pe_1_0_7_U109 ( .A1(npu_inst_pe_1_0_7_n5), .A2(
        npu_inst_pe_1_0_7_n7), .A3(npu_inst_pe_1_0_7_n8), .ZN(
        npu_inst_pe_1_0_7_n44) );
  NAND3_X1 npu_inst_pe_1_0_7_U108 ( .A1(npu_inst_pe_1_0_7_n4), .A2(
        npu_inst_pe_1_0_7_n7), .A3(npu_inst_pe_1_0_7_n8), .ZN(
        npu_inst_pe_1_0_7_n40) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_0_7_n34), .CK(
        npu_inst_pe_1_0_7_net4401), .RN(npu_inst_pe_1_0_7_n9), .Q(
        npu_inst_pe_1_0_7_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_0_7_n35), .CK(
        npu_inst_pe_1_0_7_net4401), .RN(npu_inst_pe_1_0_7_n9), .Q(
        npu_inst_pe_1_0_7_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_0_7_n36), .CK(
        npu_inst_pe_1_0_7_net4401), .RN(npu_inst_pe_1_0_7_n9), .Q(
        npu_inst_pe_1_0_7_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_0_7_n98), .CK(
        npu_inst_pe_1_0_7_net4401), .RN(npu_inst_pe_1_0_7_n9), .Q(
        npu_inst_pe_1_0_7_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_0_7_n99), .CK(
        npu_inst_pe_1_0_7_net4401), .RN(npu_inst_pe_1_0_7_n9), .Q(
        npu_inst_pe_1_0_7_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_0_7_n100), 
        .CK(npu_inst_pe_1_0_7_net4401), .RN(npu_inst_pe_1_0_7_n9), .Q(
        npu_inst_pe_1_0_7_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_0_7_n33), .CK(
        npu_inst_pe_1_0_7_net4401), .RN(npu_inst_pe_1_0_7_n9), .Q(
        npu_inst_pe_1_0_7_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_0_7_n101), 
        .CK(npu_inst_pe_1_0_7_net4401), .RN(npu_inst_pe_1_0_7_n9), .Q(
        npu_inst_pe_1_0_7_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_weight_reg_0_ ( .D(npu_inst_n112), .CK(
        npu_inst_pe_1_0_7_net4407), .RN(npu_inst_pe_1_0_7_n9), .Q(
        npu_inst_pe_1_0_7_int_q_weight_0_), .QN(npu_inst_pe_1_0_7_n27) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_weight_reg_1_ ( .D(npu_inst_n118), .CK(
        npu_inst_pe_1_0_7_net4407), .RN(npu_inst_pe_1_0_7_n9), .Q(
        npu_inst_pe_1_0_7_int_q_weight_1_), .QN(npu_inst_pe_1_0_7_n26) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_0_7_n113), 
        .CK(npu_inst_pe_1_0_7_net4407), .RN(npu_inst_pe_1_0_7_n9), .Q(
        npu_inst_pe_1_0_7_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_0_7_n107), 
        .CK(npu_inst_pe_1_0_7_net4407), .RN(npu_inst_pe_1_0_7_n9), .Q(
        npu_inst_pe_1_0_7_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_0_7_n112), 
        .CK(npu_inst_pe_1_0_7_net4407), .RN(npu_inst_pe_1_0_7_n10), .Q(
        npu_inst_pe_1_0_7_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_0_7_n106), 
        .CK(npu_inst_pe_1_0_7_net4407), .RN(npu_inst_pe_1_0_7_n10), .Q(
        npu_inst_pe_1_0_7_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_0_7_n111), 
        .CK(npu_inst_pe_1_0_7_net4407), .RN(npu_inst_pe_1_0_7_n10), .Q(
        npu_inst_pe_1_0_7_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_0_7_n105), 
        .CK(npu_inst_pe_1_0_7_net4407), .RN(npu_inst_pe_1_0_7_n10), .Q(
        npu_inst_pe_1_0_7_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_0_7_n110), 
        .CK(npu_inst_pe_1_0_7_net4407), .RN(npu_inst_pe_1_0_7_n10), .Q(
        npu_inst_pe_1_0_7_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_0_7_n104), 
        .CK(npu_inst_pe_1_0_7_net4407), .RN(npu_inst_pe_1_0_7_n10), .Q(
        npu_inst_pe_1_0_7_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_0_7_n109), 
        .CK(npu_inst_pe_1_0_7_net4407), .RN(npu_inst_pe_1_0_7_n10), .Q(
        npu_inst_pe_1_0_7_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_0_7_n103), 
        .CK(npu_inst_pe_1_0_7_net4407), .RN(npu_inst_pe_1_0_7_n10), .Q(
        npu_inst_pe_1_0_7_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_0_7_n108), 
        .CK(npu_inst_pe_1_0_7_net4407), .RN(npu_inst_pe_1_0_7_n10), .Q(
        npu_inst_pe_1_0_7_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_0_7_n102), 
        .CK(npu_inst_pe_1_0_7_net4407), .RN(npu_inst_pe_1_0_7_n10), .Q(
        npu_inst_pe_1_0_7_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_0_7_n86), 
        .CK(npu_inst_pe_1_0_7_net4407), .RN(npu_inst_pe_1_0_7_n10), .Q(
        npu_inst_pe_1_0_7_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_0_7_n87), 
        .CK(npu_inst_pe_1_0_7_net4407), .RN(npu_inst_pe_1_0_7_n10), .Q(
        npu_inst_pe_1_0_7_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_0_7_n88), 
        .CK(npu_inst_pe_1_0_7_net4407), .RN(npu_inst_pe_1_0_7_n11), .Q(
        npu_inst_pe_1_0_7_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_0_7_n89), 
        .CK(npu_inst_pe_1_0_7_net4407), .RN(npu_inst_pe_1_0_7_n11), .Q(
        npu_inst_pe_1_0_7_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_0_7_n90), 
        .CK(npu_inst_pe_1_0_7_net4407), .RN(npu_inst_pe_1_0_7_n11), .Q(
        npu_inst_pe_1_0_7_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_0_7_n91), 
        .CK(npu_inst_pe_1_0_7_net4407), .RN(npu_inst_pe_1_0_7_n11), .Q(
        npu_inst_pe_1_0_7_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_0_7_n92), 
        .CK(npu_inst_pe_1_0_7_net4407), .RN(npu_inst_pe_1_0_7_n11), .Q(
        npu_inst_pe_1_0_7_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_0_7_n93), 
        .CK(npu_inst_pe_1_0_7_net4407), .RN(npu_inst_pe_1_0_7_n11), .Q(
        npu_inst_pe_1_0_7_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_0_7_n94), 
        .CK(npu_inst_pe_1_0_7_net4407), .RN(npu_inst_pe_1_0_7_n11), .Q(
        npu_inst_pe_1_0_7_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_0_7_n95), 
        .CK(npu_inst_pe_1_0_7_net4407), .RN(npu_inst_pe_1_0_7_n11), .Q(
        npu_inst_pe_1_0_7_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_0_7_n96), 
        .CK(npu_inst_pe_1_0_7_net4407), .RN(npu_inst_pe_1_0_7_n11), .Q(
        npu_inst_pe_1_0_7_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_0_7_n97), 
        .CK(npu_inst_pe_1_0_7_net4407), .RN(npu_inst_pe_1_0_7_n11), .Q(
        npu_inst_pe_1_0_7_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_0_7_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_0_7_N84), .SE(1'b0), .GCK(npu_inst_pe_1_0_7_net4401) );
  CLKGATETST_X1 npu_inst_pe_1_0_7_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n66), .SE(1'b0), .GCK(npu_inst_pe_1_0_7_net4407) );
  MUX2_X1 npu_inst_pe_1_1_0_U162 ( .A(npu_inst_pe_1_1_0_n32), .B(
        npu_inst_pe_1_1_0_n29), .S(npu_inst_pe_1_1_0_n8), .Z(
        npu_inst_pe_1_1_0_N93) );
  MUX2_X1 npu_inst_pe_1_1_0_U161 ( .A(npu_inst_pe_1_1_0_n31), .B(
        npu_inst_pe_1_1_0_n30), .S(npu_inst_pe_1_1_0_n6), .Z(
        npu_inst_pe_1_1_0_n32) );
  MUX2_X1 npu_inst_pe_1_1_0_U160 ( .A(npu_inst_pe_1_1_0_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_1_0_int_q_reg_v_1__0_), .S(npu_inst_pe_1_1_0_n4), .Z(
        npu_inst_pe_1_1_0_n31) );
  MUX2_X1 npu_inst_pe_1_1_0_U159 ( .A(npu_inst_pe_1_1_0_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_1_0_int_q_reg_v_3__0_), .S(npu_inst_pe_1_1_0_n4), .Z(
        npu_inst_pe_1_1_0_n30) );
  MUX2_X1 npu_inst_pe_1_1_0_U158 ( .A(npu_inst_pe_1_1_0_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_1_0_int_q_reg_v_5__0_), .S(npu_inst_pe_1_1_0_n4), .Z(
        npu_inst_pe_1_1_0_n29) );
  MUX2_X1 npu_inst_pe_1_1_0_U157 ( .A(npu_inst_pe_1_1_0_n28), .B(
        npu_inst_pe_1_1_0_n23), .S(npu_inst_pe_1_1_0_n8), .Z(
        npu_inst_pe_1_1_0_N94) );
  MUX2_X1 npu_inst_pe_1_1_0_U156 ( .A(npu_inst_pe_1_1_0_n25), .B(
        npu_inst_pe_1_1_0_n24), .S(npu_inst_pe_1_1_0_n6), .Z(
        npu_inst_pe_1_1_0_n28) );
  MUX2_X1 npu_inst_pe_1_1_0_U155 ( .A(npu_inst_pe_1_1_0_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_1_0_int_q_reg_v_1__1_), .S(npu_inst_pe_1_1_0_n4), .Z(
        npu_inst_pe_1_1_0_n25) );
  MUX2_X1 npu_inst_pe_1_1_0_U154 ( .A(npu_inst_pe_1_1_0_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_1_0_int_q_reg_v_3__1_), .S(npu_inst_pe_1_1_0_n4), .Z(
        npu_inst_pe_1_1_0_n24) );
  MUX2_X1 npu_inst_pe_1_1_0_U153 ( .A(npu_inst_pe_1_1_0_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_1_0_int_q_reg_v_5__1_), .S(npu_inst_pe_1_1_0_n4), .Z(
        npu_inst_pe_1_1_0_n23) );
  MUX2_X1 npu_inst_pe_1_1_0_U152 ( .A(npu_inst_pe_1_1_0_n22), .B(
        npu_inst_pe_1_1_0_n19), .S(npu_inst_pe_1_1_0_n8), .Z(
        npu_inst_pe_1_1_0_o_data_h_1_) );
  MUX2_X1 npu_inst_pe_1_1_0_U151 ( .A(npu_inst_pe_1_1_0_n21), .B(
        npu_inst_pe_1_1_0_n20), .S(npu_inst_pe_1_1_0_n6), .Z(
        npu_inst_pe_1_1_0_n22) );
  MUX2_X1 npu_inst_pe_1_1_0_U150 ( .A(npu_inst_pe_1_1_0_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_1_0_int_q_reg_h_1__1_), .S(npu_inst_pe_1_1_0_n4), .Z(
        npu_inst_pe_1_1_0_n21) );
  MUX2_X1 npu_inst_pe_1_1_0_U149 ( .A(npu_inst_pe_1_1_0_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_1_0_int_q_reg_h_3__1_), .S(npu_inst_pe_1_1_0_n4), .Z(
        npu_inst_pe_1_1_0_n20) );
  MUX2_X1 npu_inst_pe_1_1_0_U148 ( .A(npu_inst_pe_1_1_0_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_1_0_int_q_reg_h_5__1_), .S(npu_inst_pe_1_1_0_n4), .Z(
        npu_inst_pe_1_1_0_n19) );
  MUX2_X1 npu_inst_pe_1_1_0_U147 ( .A(npu_inst_pe_1_1_0_n18), .B(
        npu_inst_pe_1_1_0_n15), .S(npu_inst_pe_1_1_0_n8), .Z(
        npu_inst_pe_1_1_0_o_data_h_0_) );
  MUX2_X1 npu_inst_pe_1_1_0_U146 ( .A(npu_inst_pe_1_1_0_n17), .B(
        npu_inst_pe_1_1_0_n16), .S(npu_inst_pe_1_1_0_n6), .Z(
        npu_inst_pe_1_1_0_n18) );
  MUX2_X1 npu_inst_pe_1_1_0_U145 ( .A(npu_inst_pe_1_1_0_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_1_0_int_q_reg_h_1__0_), .S(npu_inst_pe_1_1_0_n4), .Z(
        npu_inst_pe_1_1_0_n17) );
  MUX2_X1 npu_inst_pe_1_1_0_U144 ( .A(npu_inst_pe_1_1_0_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_1_0_int_q_reg_h_3__0_), .S(npu_inst_pe_1_1_0_n4), .Z(
        npu_inst_pe_1_1_0_n16) );
  MUX2_X1 npu_inst_pe_1_1_0_U143 ( .A(npu_inst_pe_1_1_0_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_1_0_int_q_reg_h_5__0_), .S(npu_inst_pe_1_1_0_n4), .Z(
        npu_inst_pe_1_1_0_n15) );
  XOR2_X1 npu_inst_pe_1_1_0_U142 ( .A(npu_inst_pe_1_1_0_int_data_0_), .B(
        npu_inst_pe_1_1_0_int_q_acc_0_), .Z(npu_inst_pe_1_1_0_N73) );
  AND2_X1 npu_inst_pe_1_1_0_U141 ( .A1(npu_inst_pe_1_1_0_int_q_acc_0_), .A2(
        npu_inst_pe_1_1_0_int_data_0_), .ZN(npu_inst_pe_1_1_0_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_1_0_U140 ( .A(npu_inst_pe_1_1_0_int_q_acc_0_), .B(
        npu_inst_pe_1_1_0_n13), .ZN(npu_inst_pe_1_1_0_N65) );
  OR2_X1 npu_inst_pe_1_1_0_U139 ( .A1(npu_inst_pe_1_1_0_n13), .A2(
        npu_inst_pe_1_1_0_int_q_acc_0_), .ZN(npu_inst_pe_1_1_0_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_1_0_U138 ( .A(npu_inst_pe_1_1_0_int_q_acc_2_), .B(
        npu_inst_pe_1_1_0_add_69_carry_2_), .Z(npu_inst_pe_1_1_0_N75) );
  AND2_X1 npu_inst_pe_1_1_0_U137 ( .A1(npu_inst_pe_1_1_0_add_69_carry_2_), 
        .A2(npu_inst_pe_1_1_0_int_q_acc_2_), .ZN(
        npu_inst_pe_1_1_0_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_1_0_U136 ( .A(npu_inst_pe_1_1_0_int_q_acc_3_), .B(
        npu_inst_pe_1_1_0_add_69_carry_3_), .Z(npu_inst_pe_1_1_0_N76) );
  AND2_X1 npu_inst_pe_1_1_0_U135 ( .A1(npu_inst_pe_1_1_0_add_69_carry_3_), 
        .A2(npu_inst_pe_1_1_0_int_q_acc_3_), .ZN(
        npu_inst_pe_1_1_0_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_1_0_U134 ( .A(npu_inst_pe_1_1_0_int_q_acc_4_), .B(
        npu_inst_pe_1_1_0_add_69_carry_4_), .Z(npu_inst_pe_1_1_0_N77) );
  AND2_X1 npu_inst_pe_1_1_0_U133 ( .A1(npu_inst_pe_1_1_0_add_69_carry_4_), 
        .A2(npu_inst_pe_1_1_0_int_q_acc_4_), .ZN(
        npu_inst_pe_1_1_0_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_1_0_U132 ( .A(npu_inst_pe_1_1_0_int_q_acc_5_), .B(
        npu_inst_pe_1_1_0_add_69_carry_5_), .Z(npu_inst_pe_1_1_0_N78) );
  AND2_X1 npu_inst_pe_1_1_0_U131 ( .A1(npu_inst_pe_1_1_0_add_69_carry_5_), 
        .A2(npu_inst_pe_1_1_0_int_q_acc_5_), .ZN(
        npu_inst_pe_1_1_0_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_1_0_U130 ( .A(npu_inst_pe_1_1_0_int_q_acc_6_), .B(
        npu_inst_pe_1_1_0_add_69_carry_6_), .Z(npu_inst_pe_1_1_0_N79) );
  AND2_X1 npu_inst_pe_1_1_0_U129 ( .A1(npu_inst_pe_1_1_0_add_69_carry_6_), 
        .A2(npu_inst_pe_1_1_0_int_q_acc_6_), .ZN(
        npu_inst_pe_1_1_0_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_1_0_U128 ( .A(npu_inst_pe_1_1_0_int_q_acc_7_), .B(
        npu_inst_pe_1_1_0_add_69_carry_7_), .Z(npu_inst_pe_1_1_0_N80) );
  XNOR2_X1 npu_inst_pe_1_1_0_U127 ( .A(npu_inst_pe_1_1_0_sub_67_carry_2_), .B(
        npu_inst_pe_1_1_0_int_q_acc_2_), .ZN(npu_inst_pe_1_1_0_N67) );
  OR2_X1 npu_inst_pe_1_1_0_U126 ( .A1(npu_inst_pe_1_1_0_int_q_acc_2_), .A2(
        npu_inst_pe_1_1_0_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_1_0_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_1_0_U125 ( .A(npu_inst_pe_1_1_0_sub_67_carry_3_), .B(
        npu_inst_pe_1_1_0_int_q_acc_3_), .ZN(npu_inst_pe_1_1_0_N68) );
  OR2_X1 npu_inst_pe_1_1_0_U124 ( .A1(npu_inst_pe_1_1_0_int_q_acc_3_), .A2(
        npu_inst_pe_1_1_0_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_1_0_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_1_0_U123 ( .A(npu_inst_pe_1_1_0_sub_67_carry_4_), .B(
        npu_inst_pe_1_1_0_int_q_acc_4_), .ZN(npu_inst_pe_1_1_0_N69) );
  OR2_X1 npu_inst_pe_1_1_0_U122 ( .A1(npu_inst_pe_1_1_0_int_q_acc_4_), .A2(
        npu_inst_pe_1_1_0_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_1_0_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_1_0_U121 ( .A(npu_inst_pe_1_1_0_sub_67_carry_5_), .B(
        npu_inst_pe_1_1_0_int_q_acc_5_), .ZN(npu_inst_pe_1_1_0_N70) );
  OR2_X1 npu_inst_pe_1_1_0_U120 ( .A1(npu_inst_pe_1_1_0_int_q_acc_5_), .A2(
        npu_inst_pe_1_1_0_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_1_0_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_1_0_U119 ( .A(npu_inst_pe_1_1_0_sub_67_carry_6_), .B(
        npu_inst_pe_1_1_0_int_q_acc_6_), .ZN(npu_inst_pe_1_1_0_N71) );
  OR2_X1 npu_inst_pe_1_1_0_U118 ( .A1(npu_inst_pe_1_1_0_int_q_acc_6_), .A2(
        npu_inst_pe_1_1_0_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_1_0_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_1_0_U117 ( .A(npu_inst_pe_1_1_0_int_q_acc_7_), .B(
        npu_inst_pe_1_1_0_sub_67_carry_7_), .ZN(npu_inst_pe_1_1_0_N72) );
  INV_X1 npu_inst_pe_1_1_0_U116 ( .A(npu_inst_n79), .ZN(npu_inst_pe_1_1_0_n7)
         );
  INV_X1 npu_inst_pe_1_1_0_U115 ( .A(npu_inst_pe_1_1_0_n7), .ZN(
        npu_inst_pe_1_1_0_n6) );
  INV_X1 npu_inst_pe_1_1_0_U114 ( .A(npu_inst_n59), .ZN(npu_inst_pe_1_1_0_n3)
         );
  AOI22_X1 npu_inst_pe_1_1_0_U113 ( .A1(npu_inst_int_data_y_2__0__0_), .A2(
        npu_inst_pe_1_1_0_n58), .B1(npu_inst_pe_1_1_0_n119), .B2(
        npu_inst_pe_1_1_0_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_1_0_n57) );
  INV_X1 npu_inst_pe_1_1_0_U112 ( .A(npu_inst_pe_1_1_0_n57), .ZN(
        npu_inst_pe_1_1_0_n108) );
  AOI22_X1 npu_inst_pe_1_1_0_U111 ( .A1(npu_inst_int_data_y_2__0__0_), .A2(
        npu_inst_pe_1_1_0_n54), .B1(npu_inst_pe_1_1_0_n118), .B2(
        npu_inst_pe_1_1_0_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_1_0_n53) );
  INV_X1 npu_inst_pe_1_1_0_U110 ( .A(npu_inst_pe_1_1_0_n53), .ZN(
        npu_inst_pe_1_1_0_n109) );
  AOI22_X1 npu_inst_pe_1_1_0_U107 ( .A1(npu_inst_int_data_y_2__0__0_), .A2(
        npu_inst_pe_1_1_0_n50), .B1(npu_inst_pe_1_1_0_n117), .B2(
        npu_inst_pe_1_1_0_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_1_0_n49) );
  INV_X1 npu_inst_pe_1_1_0_U106 ( .A(npu_inst_pe_1_1_0_n49), .ZN(
        npu_inst_pe_1_1_0_n110) );
  AOI22_X1 npu_inst_pe_1_1_0_U105 ( .A1(npu_inst_int_data_y_2__0__0_), .A2(
        npu_inst_pe_1_1_0_n46), .B1(npu_inst_pe_1_1_0_n116), .B2(
        npu_inst_pe_1_1_0_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_1_0_n45) );
  INV_X1 npu_inst_pe_1_1_0_U104 ( .A(npu_inst_pe_1_1_0_n45), .ZN(
        npu_inst_pe_1_1_0_n111) );
  AOI22_X1 npu_inst_pe_1_1_0_U103 ( .A1(npu_inst_int_data_y_2__0__0_), .A2(
        npu_inst_pe_1_1_0_n42), .B1(npu_inst_pe_1_1_0_n115), .B2(
        npu_inst_pe_1_1_0_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_1_0_n41) );
  INV_X1 npu_inst_pe_1_1_0_U102 ( .A(npu_inst_pe_1_1_0_n41), .ZN(
        npu_inst_pe_1_1_0_n112) );
  AOI22_X1 npu_inst_pe_1_1_0_U101 ( .A1(npu_inst_int_data_y_2__0__1_), .A2(
        npu_inst_pe_1_1_0_n58), .B1(npu_inst_pe_1_1_0_n119), .B2(
        npu_inst_pe_1_1_0_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_1_0_n59) );
  INV_X1 npu_inst_pe_1_1_0_U100 ( .A(npu_inst_pe_1_1_0_n59), .ZN(
        npu_inst_pe_1_1_0_n102) );
  AOI22_X1 npu_inst_pe_1_1_0_U99 ( .A1(npu_inst_int_data_y_2__0__1_), .A2(
        npu_inst_pe_1_1_0_n54), .B1(npu_inst_pe_1_1_0_n118), .B2(
        npu_inst_pe_1_1_0_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_1_0_n55) );
  INV_X1 npu_inst_pe_1_1_0_U98 ( .A(npu_inst_pe_1_1_0_n55), .ZN(
        npu_inst_pe_1_1_0_n103) );
  AOI22_X1 npu_inst_pe_1_1_0_U97 ( .A1(npu_inst_int_data_y_2__0__1_), .A2(
        npu_inst_pe_1_1_0_n50), .B1(npu_inst_pe_1_1_0_n117), .B2(
        npu_inst_pe_1_1_0_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_1_0_n51) );
  INV_X1 npu_inst_pe_1_1_0_U96 ( .A(npu_inst_pe_1_1_0_n51), .ZN(
        npu_inst_pe_1_1_0_n104) );
  AOI22_X1 npu_inst_pe_1_1_0_U95 ( .A1(npu_inst_int_data_y_2__0__1_), .A2(
        npu_inst_pe_1_1_0_n46), .B1(npu_inst_pe_1_1_0_n116), .B2(
        npu_inst_pe_1_1_0_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_1_0_n47) );
  INV_X1 npu_inst_pe_1_1_0_U94 ( .A(npu_inst_pe_1_1_0_n47), .ZN(
        npu_inst_pe_1_1_0_n105) );
  AOI22_X1 npu_inst_pe_1_1_0_U93 ( .A1(npu_inst_int_data_y_2__0__1_), .A2(
        npu_inst_pe_1_1_0_n42), .B1(npu_inst_pe_1_1_0_n115), .B2(
        npu_inst_pe_1_1_0_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_1_0_n43) );
  INV_X1 npu_inst_pe_1_1_0_U92 ( .A(npu_inst_pe_1_1_0_n43), .ZN(
        npu_inst_pe_1_1_0_n106) );
  AOI22_X1 npu_inst_pe_1_1_0_U91 ( .A1(npu_inst_pe_1_1_0_n38), .A2(
        npu_inst_int_data_y_2__0__1_), .B1(npu_inst_pe_1_1_0_n114), .B2(
        npu_inst_pe_1_1_0_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_1_0_n39) );
  INV_X1 npu_inst_pe_1_1_0_U90 ( .A(npu_inst_pe_1_1_0_n39), .ZN(
        npu_inst_pe_1_1_0_n107) );
  AOI22_X1 npu_inst_pe_1_1_0_U89 ( .A1(npu_inst_pe_1_1_0_n38), .A2(
        npu_inst_int_data_y_2__0__0_), .B1(npu_inst_pe_1_1_0_n114), .B2(
        npu_inst_pe_1_1_0_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_1_0_n37) );
  INV_X1 npu_inst_pe_1_1_0_U88 ( .A(npu_inst_pe_1_1_0_n37), .ZN(
        npu_inst_pe_1_1_0_n113) );
  NAND2_X1 npu_inst_pe_1_1_0_U87 ( .A1(npu_inst_pe_1_1_0_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_1_0_n60), .ZN(npu_inst_pe_1_1_0_n74) );
  OAI21_X1 npu_inst_pe_1_1_0_U86 ( .B1(npu_inst_pe_1_1_0_n63), .B2(
        npu_inst_pe_1_1_0_n60), .A(npu_inst_pe_1_1_0_n74), .ZN(
        npu_inst_pe_1_1_0_n97) );
  NAND2_X1 npu_inst_pe_1_1_0_U85 ( .A1(npu_inst_pe_1_1_0_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_1_0_n60), .ZN(npu_inst_pe_1_1_0_n73) );
  OAI21_X1 npu_inst_pe_1_1_0_U84 ( .B1(npu_inst_pe_1_1_0_n61), .B2(
        npu_inst_pe_1_1_0_n60), .A(npu_inst_pe_1_1_0_n73), .ZN(
        npu_inst_pe_1_1_0_n96) );
  NAND2_X1 npu_inst_pe_1_1_0_U83 ( .A1(npu_inst_pe_1_1_0_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_1_0_n56), .ZN(npu_inst_pe_1_1_0_n72) );
  OAI21_X1 npu_inst_pe_1_1_0_U82 ( .B1(npu_inst_pe_1_1_0_n63), .B2(
        npu_inst_pe_1_1_0_n56), .A(npu_inst_pe_1_1_0_n72), .ZN(
        npu_inst_pe_1_1_0_n95) );
  NAND2_X1 npu_inst_pe_1_1_0_U81 ( .A1(npu_inst_pe_1_1_0_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_1_0_n56), .ZN(npu_inst_pe_1_1_0_n71) );
  OAI21_X1 npu_inst_pe_1_1_0_U80 ( .B1(npu_inst_pe_1_1_0_n61), .B2(
        npu_inst_pe_1_1_0_n56), .A(npu_inst_pe_1_1_0_n71), .ZN(
        npu_inst_pe_1_1_0_n94) );
  NAND2_X1 npu_inst_pe_1_1_0_U79 ( .A1(npu_inst_pe_1_1_0_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_1_0_n52), .ZN(npu_inst_pe_1_1_0_n70) );
  OAI21_X1 npu_inst_pe_1_1_0_U78 ( .B1(npu_inst_pe_1_1_0_n63), .B2(
        npu_inst_pe_1_1_0_n52), .A(npu_inst_pe_1_1_0_n70), .ZN(
        npu_inst_pe_1_1_0_n93) );
  NAND2_X1 npu_inst_pe_1_1_0_U77 ( .A1(npu_inst_pe_1_1_0_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_1_0_n52), .ZN(npu_inst_pe_1_1_0_n69) );
  OAI21_X1 npu_inst_pe_1_1_0_U76 ( .B1(npu_inst_pe_1_1_0_n61), .B2(
        npu_inst_pe_1_1_0_n52), .A(npu_inst_pe_1_1_0_n69), .ZN(
        npu_inst_pe_1_1_0_n92) );
  NAND2_X1 npu_inst_pe_1_1_0_U75 ( .A1(npu_inst_pe_1_1_0_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_1_0_n48), .ZN(npu_inst_pe_1_1_0_n68) );
  OAI21_X1 npu_inst_pe_1_1_0_U74 ( .B1(npu_inst_pe_1_1_0_n63), .B2(
        npu_inst_pe_1_1_0_n48), .A(npu_inst_pe_1_1_0_n68), .ZN(
        npu_inst_pe_1_1_0_n91) );
  NAND2_X1 npu_inst_pe_1_1_0_U73 ( .A1(npu_inst_pe_1_1_0_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_1_0_n48), .ZN(npu_inst_pe_1_1_0_n67) );
  OAI21_X1 npu_inst_pe_1_1_0_U72 ( .B1(npu_inst_pe_1_1_0_n61), .B2(
        npu_inst_pe_1_1_0_n48), .A(npu_inst_pe_1_1_0_n67), .ZN(
        npu_inst_pe_1_1_0_n90) );
  NAND2_X1 npu_inst_pe_1_1_0_U71 ( .A1(npu_inst_pe_1_1_0_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_1_0_n44), .ZN(npu_inst_pe_1_1_0_n66) );
  OAI21_X1 npu_inst_pe_1_1_0_U70 ( .B1(npu_inst_pe_1_1_0_n63), .B2(
        npu_inst_pe_1_1_0_n44), .A(npu_inst_pe_1_1_0_n66), .ZN(
        npu_inst_pe_1_1_0_n89) );
  NAND2_X1 npu_inst_pe_1_1_0_U69 ( .A1(npu_inst_pe_1_1_0_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_1_0_n44), .ZN(npu_inst_pe_1_1_0_n65) );
  OAI21_X1 npu_inst_pe_1_1_0_U68 ( .B1(npu_inst_pe_1_1_0_n61), .B2(
        npu_inst_pe_1_1_0_n44), .A(npu_inst_pe_1_1_0_n65), .ZN(
        npu_inst_pe_1_1_0_n88) );
  NAND2_X1 npu_inst_pe_1_1_0_U67 ( .A1(npu_inst_pe_1_1_0_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_1_0_n40), .ZN(npu_inst_pe_1_1_0_n64) );
  OAI21_X1 npu_inst_pe_1_1_0_U66 ( .B1(npu_inst_pe_1_1_0_n63), .B2(
        npu_inst_pe_1_1_0_n40), .A(npu_inst_pe_1_1_0_n64), .ZN(
        npu_inst_pe_1_1_0_n87) );
  NAND2_X1 npu_inst_pe_1_1_0_U65 ( .A1(npu_inst_pe_1_1_0_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_1_0_n40), .ZN(npu_inst_pe_1_1_0_n62) );
  OAI21_X1 npu_inst_pe_1_1_0_U64 ( .B1(npu_inst_pe_1_1_0_n61), .B2(
        npu_inst_pe_1_1_0_n40), .A(npu_inst_pe_1_1_0_n62), .ZN(
        npu_inst_pe_1_1_0_n86) );
  AND2_X1 npu_inst_pe_1_1_0_U63 ( .A1(npu_inst_pe_1_1_0_N93), .A2(npu_inst_n59), .ZN(npu_inst_int_data_y_1__0__0_) );
  AND2_X1 npu_inst_pe_1_1_0_U62 ( .A1(npu_inst_n59), .A2(npu_inst_pe_1_1_0_N94), .ZN(npu_inst_int_data_y_1__0__1_) );
  NOR3_X1 npu_inst_pe_1_1_0_U61 ( .A1(npu_inst_pe_1_1_0_n26), .A2(npu_inst_n59), .A3(npu_inst_int_ckg[55]), .ZN(npu_inst_pe_1_1_0_n85) );
  OR2_X1 npu_inst_pe_1_1_0_U60 ( .A1(npu_inst_pe_1_1_0_n85), .A2(
        npu_inst_pe_1_1_0_n2), .ZN(npu_inst_pe_1_1_0_N84) );
  AND2_X1 npu_inst_pe_1_1_0_U59 ( .A1(npu_inst_pe_1_1_0_int_q_acc_0_), .A2(
        npu_inst_pe_1_1_0_n1), .ZN(npu_inst_int_data_res_1__0__0_) );
  AND2_X1 npu_inst_pe_1_1_0_U58 ( .A1(npu_inst_pe_1_1_0_n2), .A2(
        npu_inst_pe_1_1_0_int_q_acc_7_), .ZN(npu_inst_int_data_res_1__0__7_)
         );
  AND2_X1 npu_inst_pe_1_1_0_U57 ( .A1(npu_inst_pe_1_1_0_int_q_acc_1_), .A2(
        npu_inst_pe_1_1_0_n1), .ZN(npu_inst_int_data_res_1__0__1_) );
  AND2_X1 npu_inst_pe_1_1_0_U56 ( .A1(npu_inst_pe_1_1_0_int_q_acc_2_), .A2(
        npu_inst_pe_1_1_0_n1), .ZN(npu_inst_int_data_res_1__0__2_) );
  AND2_X1 npu_inst_pe_1_1_0_U55 ( .A1(npu_inst_pe_1_1_0_int_q_acc_3_), .A2(
        npu_inst_pe_1_1_0_n2), .ZN(npu_inst_int_data_res_1__0__3_) );
  AND2_X1 npu_inst_pe_1_1_0_U54 ( .A1(npu_inst_pe_1_1_0_int_q_acc_4_), .A2(
        npu_inst_pe_1_1_0_n2), .ZN(npu_inst_int_data_res_1__0__4_) );
  AND2_X1 npu_inst_pe_1_1_0_U53 ( .A1(npu_inst_pe_1_1_0_int_q_acc_5_), .A2(
        npu_inst_pe_1_1_0_n2), .ZN(npu_inst_int_data_res_1__0__5_) );
  AND2_X1 npu_inst_pe_1_1_0_U52 ( .A1(npu_inst_pe_1_1_0_int_q_acc_6_), .A2(
        npu_inst_pe_1_1_0_n2), .ZN(npu_inst_int_data_res_1__0__6_) );
  AOI222_X1 npu_inst_pe_1_1_0_U51 ( .A1(npu_inst_int_data_res_2__0__0_), .A2(
        npu_inst_pe_1_1_0_n1), .B1(npu_inst_pe_1_1_0_N73), .B2(
        npu_inst_pe_1_1_0_n76), .C1(npu_inst_pe_1_1_0_N65), .C2(
        npu_inst_pe_1_1_0_n77), .ZN(npu_inst_pe_1_1_0_n84) );
  INV_X1 npu_inst_pe_1_1_0_U50 ( .A(npu_inst_pe_1_1_0_n84), .ZN(
        npu_inst_pe_1_1_0_n101) );
  AOI222_X1 npu_inst_pe_1_1_0_U49 ( .A1(npu_inst_int_data_res_2__0__7_), .A2(
        npu_inst_pe_1_1_0_n1), .B1(npu_inst_pe_1_1_0_N80), .B2(
        npu_inst_pe_1_1_0_n76), .C1(npu_inst_pe_1_1_0_N72), .C2(
        npu_inst_pe_1_1_0_n77), .ZN(npu_inst_pe_1_1_0_n75) );
  INV_X1 npu_inst_pe_1_1_0_U48 ( .A(npu_inst_pe_1_1_0_n75), .ZN(
        npu_inst_pe_1_1_0_n33) );
  AOI222_X1 npu_inst_pe_1_1_0_U47 ( .A1(npu_inst_int_data_res_2__0__1_), .A2(
        npu_inst_pe_1_1_0_n1), .B1(npu_inst_pe_1_1_0_N74), .B2(
        npu_inst_pe_1_1_0_n76), .C1(npu_inst_pe_1_1_0_N66), .C2(
        npu_inst_pe_1_1_0_n77), .ZN(npu_inst_pe_1_1_0_n83) );
  INV_X1 npu_inst_pe_1_1_0_U46 ( .A(npu_inst_pe_1_1_0_n83), .ZN(
        npu_inst_pe_1_1_0_n100) );
  AOI222_X1 npu_inst_pe_1_1_0_U45 ( .A1(npu_inst_int_data_res_2__0__2_), .A2(
        npu_inst_pe_1_1_0_n1), .B1(npu_inst_pe_1_1_0_N75), .B2(
        npu_inst_pe_1_1_0_n76), .C1(npu_inst_pe_1_1_0_N67), .C2(
        npu_inst_pe_1_1_0_n77), .ZN(npu_inst_pe_1_1_0_n82) );
  INV_X1 npu_inst_pe_1_1_0_U44 ( .A(npu_inst_pe_1_1_0_n82), .ZN(
        npu_inst_pe_1_1_0_n99) );
  AOI222_X1 npu_inst_pe_1_1_0_U43 ( .A1(npu_inst_int_data_res_2__0__3_), .A2(
        npu_inst_pe_1_1_0_n1), .B1(npu_inst_pe_1_1_0_N76), .B2(
        npu_inst_pe_1_1_0_n76), .C1(npu_inst_pe_1_1_0_N68), .C2(
        npu_inst_pe_1_1_0_n77), .ZN(npu_inst_pe_1_1_0_n81) );
  INV_X1 npu_inst_pe_1_1_0_U42 ( .A(npu_inst_pe_1_1_0_n81), .ZN(
        npu_inst_pe_1_1_0_n98) );
  AOI222_X1 npu_inst_pe_1_1_0_U41 ( .A1(npu_inst_int_data_res_2__0__4_), .A2(
        npu_inst_pe_1_1_0_n1), .B1(npu_inst_pe_1_1_0_N77), .B2(
        npu_inst_pe_1_1_0_n76), .C1(npu_inst_pe_1_1_0_N69), .C2(
        npu_inst_pe_1_1_0_n77), .ZN(npu_inst_pe_1_1_0_n80) );
  INV_X1 npu_inst_pe_1_1_0_U40 ( .A(npu_inst_pe_1_1_0_n80), .ZN(
        npu_inst_pe_1_1_0_n36) );
  AOI222_X1 npu_inst_pe_1_1_0_U39 ( .A1(npu_inst_int_data_res_2__0__5_), .A2(
        npu_inst_pe_1_1_0_n1), .B1(npu_inst_pe_1_1_0_N78), .B2(
        npu_inst_pe_1_1_0_n76), .C1(npu_inst_pe_1_1_0_N70), .C2(
        npu_inst_pe_1_1_0_n77), .ZN(npu_inst_pe_1_1_0_n79) );
  INV_X1 npu_inst_pe_1_1_0_U38 ( .A(npu_inst_pe_1_1_0_n79), .ZN(
        npu_inst_pe_1_1_0_n35) );
  AOI222_X1 npu_inst_pe_1_1_0_U37 ( .A1(npu_inst_int_data_res_2__0__6_), .A2(
        npu_inst_pe_1_1_0_n1), .B1(npu_inst_pe_1_1_0_N79), .B2(
        npu_inst_pe_1_1_0_n76), .C1(npu_inst_pe_1_1_0_N71), .C2(
        npu_inst_pe_1_1_0_n77), .ZN(npu_inst_pe_1_1_0_n78) );
  INV_X1 npu_inst_pe_1_1_0_U36 ( .A(npu_inst_pe_1_1_0_n78), .ZN(
        npu_inst_pe_1_1_0_n34) );
  AND2_X1 npu_inst_pe_1_1_0_U35 ( .A1(npu_inst_pe_1_1_0_o_data_h_1_), .A2(
        npu_inst_pe_1_1_0_int_q_weight_1_), .ZN(npu_inst_pe_1_1_0_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_1_0_U34 ( .A1(npu_inst_pe_1_1_0_o_data_h_0_), .A2(
        npu_inst_pe_1_1_0_int_q_weight_1_), .ZN(npu_inst_pe_1_1_0_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_1_0_U33 ( .A(npu_inst_pe_1_1_0_int_data_1_), .ZN(
        npu_inst_pe_1_1_0_n14) );
  AOI22_X1 npu_inst_pe_1_1_0_U32 ( .A1(npu_inst_n59), .A2(
        npu_inst_int_data_y_2__0__1_), .B1(npu_inst_pe_1_1_0_n3), .B2(
        npu_inst_int_data_x_1__1__1_), .ZN(npu_inst_pe_1_1_0_n63) );
  AOI22_X1 npu_inst_pe_1_1_0_U31 ( .A1(npu_inst_n59), .A2(
        npu_inst_int_data_y_2__0__0_), .B1(npu_inst_pe_1_1_0_n3), .B2(
        npu_inst_int_data_x_1__1__0_), .ZN(npu_inst_pe_1_1_0_n61) );
  INV_X1 npu_inst_pe_1_1_0_U30 ( .A(npu_inst_pe_1_1_0_int_data_0_), .ZN(
        npu_inst_pe_1_1_0_n13) );
  INV_X1 npu_inst_pe_1_1_0_U29 ( .A(npu_inst_n71), .ZN(npu_inst_pe_1_1_0_n5)
         );
  OR3_X1 npu_inst_pe_1_1_0_U28 ( .A1(npu_inst_pe_1_1_0_n6), .A2(
        npu_inst_pe_1_1_0_n8), .A3(npu_inst_pe_1_1_0_n5), .ZN(
        npu_inst_pe_1_1_0_n56) );
  OR3_X1 npu_inst_pe_1_1_0_U27 ( .A1(npu_inst_pe_1_1_0_n5), .A2(
        npu_inst_pe_1_1_0_n8), .A3(npu_inst_pe_1_1_0_n7), .ZN(
        npu_inst_pe_1_1_0_n48) );
  INV_X1 npu_inst_pe_1_1_0_U26 ( .A(npu_inst_pe_1_1_0_n5), .ZN(
        npu_inst_pe_1_1_0_n4) );
  OR3_X1 npu_inst_pe_1_1_0_U25 ( .A1(npu_inst_pe_1_1_0_n4), .A2(
        npu_inst_pe_1_1_0_n8), .A3(npu_inst_pe_1_1_0_n7), .ZN(
        npu_inst_pe_1_1_0_n52) );
  OR3_X1 npu_inst_pe_1_1_0_U24 ( .A1(npu_inst_pe_1_1_0_n6), .A2(
        npu_inst_pe_1_1_0_n8), .A3(npu_inst_pe_1_1_0_n4), .ZN(
        npu_inst_pe_1_1_0_n60) );
  NOR2_X1 npu_inst_pe_1_1_0_U23 ( .A1(npu_inst_pe_1_1_0_n60), .A2(
        npu_inst_pe_1_1_0_n3), .ZN(npu_inst_pe_1_1_0_n58) );
  NOR2_X1 npu_inst_pe_1_1_0_U22 ( .A1(npu_inst_pe_1_1_0_n56), .A2(
        npu_inst_pe_1_1_0_n3), .ZN(npu_inst_pe_1_1_0_n54) );
  NOR2_X1 npu_inst_pe_1_1_0_U21 ( .A1(npu_inst_pe_1_1_0_n52), .A2(
        npu_inst_pe_1_1_0_n3), .ZN(npu_inst_pe_1_1_0_n50) );
  NOR2_X1 npu_inst_pe_1_1_0_U20 ( .A1(npu_inst_pe_1_1_0_n48), .A2(
        npu_inst_pe_1_1_0_n3), .ZN(npu_inst_pe_1_1_0_n46) );
  NOR2_X1 npu_inst_pe_1_1_0_U19 ( .A1(npu_inst_pe_1_1_0_n40), .A2(
        npu_inst_pe_1_1_0_n3), .ZN(npu_inst_pe_1_1_0_n38) );
  NOR2_X1 npu_inst_pe_1_1_0_U18 ( .A1(npu_inst_pe_1_1_0_n44), .A2(
        npu_inst_pe_1_1_0_n3), .ZN(npu_inst_pe_1_1_0_n42) );
  BUF_X1 npu_inst_pe_1_1_0_U17 ( .A(npu_inst_n105), .Z(npu_inst_pe_1_1_0_n8)
         );
  INV_X1 npu_inst_pe_1_1_0_U16 ( .A(npu_inst_n126), .ZN(npu_inst_pe_1_1_0_n12)
         );
  INV_X1 npu_inst_pe_1_1_0_U15 ( .A(npu_inst_pe_1_1_0_n38), .ZN(
        npu_inst_pe_1_1_0_n114) );
  INV_X1 npu_inst_pe_1_1_0_U14 ( .A(npu_inst_pe_1_1_0_n58), .ZN(
        npu_inst_pe_1_1_0_n119) );
  INV_X1 npu_inst_pe_1_1_0_U13 ( .A(npu_inst_pe_1_1_0_n54), .ZN(
        npu_inst_pe_1_1_0_n118) );
  INV_X1 npu_inst_pe_1_1_0_U12 ( .A(npu_inst_pe_1_1_0_n50), .ZN(
        npu_inst_pe_1_1_0_n117) );
  INV_X1 npu_inst_pe_1_1_0_U11 ( .A(npu_inst_pe_1_1_0_n46), .ZN(
        npu_inst_pe_1_1_0_n116) );
  INV_X1 npu_inst_pe_1_1_0_U10 ( .A(npu_inst_pe_1_1_0_n42), .ZN(
        npu_inst_pe_1_1_0_n115) );
  BUF_X1 npu_inst_pe_1_1_0_U9 ( .A(npu_inst_n34), .Z(npu_inst_pe_1_1_0_n2) );
  BUF_X1 npu_inst_pe_1_1_0_U8 ( .A(npu_inst_n34), .Z(npu_inst_pe_1_1_0_n1) );
  BUF_X1 npu_inst_pe_1_1_0_U7 ( .A(npu_inst_pe_1_1_0_n12), .Z(
        npu_inst_pe_1_1_0_n11) );
  BUF_X1 npu_inst_pe_1_1_0_U6 ( .A(npu_inst_pe_1_1_0_n12), .Z(
        npu_inst_pe_1_1_0_n10) );
  BUF_X1 npu_inst_pe_1_1_0_U5 ( .A(npu_inst_pe_1_1_0_n12), .Z(
        npu_inst_pe_1_1_0_n9) );
  NOR2_X1 npu_inst_pe_1_1_0_U4 ( .A1(npu_inst_pe_1_1_0_int_q_weight_0_), .A2(
        npu_inst_pe_1_1_0_n1), .ZN(npu_inst_pe_1_1_0_n76) );
  NOR2_X1 npu_inst_pe_1_1_0_U3 ( .A1(npu_inst_pe_1_1_0_n27), .A2(
        npu_inst_pe_1_1_0_n1), .ZN(npu_inst_pe_1_1_0_n77) );
  FA_X1 npu_inst_pe_1_1_0_sub_67_U2_1 ( .A(npu_inst_pe_1_1_0_int_q_acc_1_), 
        .B(npu_inst_pe_1_1_0_n14), .CI(npu_inst_pe_1_1_0_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_1_0_sub_67_carry_2_), .S(npu_inst_pe_1_1_0_N66) );
  FA_X1 npu_inst_pe_1_1_0_add_69_U1_1 ( .A(npu_inst_pe_1_1_0_int_q_acc_1_), 
        .B(npu_inst_pe_1_1_0_int_data_1_), .CI(
        npu_inst_pe_1_1_0_add_69_carry_1_), .CO(
        npu_inst_pe_1_1_0_add_69_carry_2_), .S(npu_inst_pe_1_1_0_N74) );
  NAND3_X1 npu_inst_pe_1_1_0_U109 ( .A1(npu_inst_pe_1_1_0_n5), .A2(
        npu_inst_pe_1_1_0_n7), .A3(npu_inst_pe_1_1_0_n8), .ZN(
        npu_inst_pe_1_1_0_n44) );
  NAND3_X1 npu_inst_pe_1_1_0_U108 ( .A1(npu_inst_pe_1_1_0_n4), .A2(
        npu_inst_pe_1_1_0_n7), .A3(npu_inst_pe_1_1_0_n8), .ZN(
        npu_inst_pe_1_1_0_n40) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_1_0_n34), .CK(
        npu_inst_pe_1_1_0_net4378), .RN(npu_inst_pe_1_1_0_n9), .Q(
        npu_inst_pe_1_1_0_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_1_0_n35), .CK(
        npu_inst_pe_1_1_0_net4378), .RN(npu_inst_pe_1_1_0_n9), .Q(
        npu_inst_pe_1_1_0_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_1_0_n36), .CK(
        npu_inst_pe_1_1_0_net4378), .RN(npu_inst_pe_1_1_0_n9), .Q(
        npu_inst_pe_1_1_0_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_1_0_n98), .CK(
        npu_inst_pe_1_1_0_net4378), .RN(npu_inst_pe_1_1_0_n9), .Q(
        npu_inst_pe_1_1_0_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_1_0_n99), .CK(
        npu_inst_pe_1_1_0_net4378), .RN(npu_inst_pe_1_1_0_n9), .Q(
        npu_inst_pe_1_1_0_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_1_0_n100), 
        .CK(npu_inst_pe_1_1_0_net4378), .RN(npu_inst_pe_1_1_0_n9), .Q(
        npu_inst_pe_1_1_0_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_1_0_n33), .CK(
        npu_inst_pe_1_1_0_net4378), .RN(npu_inst_pe_1_1_0_n9), .Q(
        npu_inst_pe_1_1_0_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_1_0_n101), 
        .CK(npu_inst_pe_1_1_0_net4378), .RN(npu_inst_pe_1_1_0_n9), .Q(
        npu_inst_pe_1_1_0_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_weight_reg_0_ ( .D(npu_inst_n112), .CK(
        npu_inst_pe_1_1_0_net4384), .RN(npu_inst_pe_1_1_0_n9), .Q(
        npu_inst_pe_1_1_0_int_q_weight_0_), .QN(npu_inst_pe_1_1_0_n27) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_weight_reg_1_ ( .D(npu_inst_n118), .CK(
        npu_inst_pe_1_1_0_net4384), .RN(npu_inst_pe_1_1_0_n9), .Q(
        npu_inst_pe_1_1_0_int_q_weight_1_), .QN(npu_inst_pe_1_1_0_n26) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_1_0_n113), 
        .CK(npu_inst_pe_1_1_0_net4384), .RN(npu_inst_pe_1_1_0_n9), .Q(
        npu_inst_pe_1_1_0_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_1_0_n107), 
        .CK(npu_inst_pe_1_1_0_net4384), .RN(npu_inst_pe_1_1_0_n9), .Q(
        npu_inst_pe_1_1_0_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_1_0_n112), 
        .CK(npu_inst_pe_1_1_0_net4384), .RN(npu_inst_pe_1_1_0_n10), .Q(
        npu_inst_pe_1_1_0_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_1_0_n106), 
        .CK(npu_inst_pe_1_1_0_net4384), .RN(npu_inst_pe_1_1_0_n10), .Q(
        npu_inst_pe_1_1_0_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_1_0_n111), 
        .CK(npu_inst_pe_1_1_0_net4384), .RN(npu_inst_pe_1_1_0_n10), .Q(
        npu_inst_pe_1_1_0_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_1_0_n105), 
        .CK(npu_inst_pe_1_1_0_net4384), .RN(npu_inst_pe_1_1_0_n10), .Q(
        npu_inst_pe_1_1_0_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_1_0_n110), 
        .CK(npu_inst_pe_1_1_0_net4384), .RN(npu_inst_pe_1_1_0_n10), .Q(
        npu_inst_pe_1_1_0_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_1_0_n104), 
        .CK(npu_inst_pe_1_1_0_net4384), .RN(npu_inst_pe_1_1_0_n10), .Q(
        npu_inst_pe_1_1_0_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_1_0_n109), 
        .CK(npu_inst_pe_1_1_0_net4384), .RN(npu_inst_pe_1_1_0_n10), .Q(
        npu_inst_pe_1_1_0_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_1_0_n103), 
        .CK(npu_inst_pe_1_1_0_net4384), .RN(npu_inst_pe_1_1_0_n10), .Q(
        npu_inst_pe_1_1_0_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_1_0_n108), 
        .CK(npu_inst_pe_1_1_0_net4384), .RN(npu_inst_pe_1_1_0_n10), .Q(
        npu_inst_pe_1_1_0_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_1_0_n102), 
        .CK(npu_inst_pe_1_1_0_net4384), .RN(npu_inst_pe_1_1_0_n10), .Q(
        npu_inst_pe_1_1_0_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_1_0_n86), 
        .CK(npu_inst_pe_1_1_0_net4384), .RN(npu_inst_pe_1_1_0_n10), .Q(
        npu_inst_pe_1_1_0_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_1_0_n87), 
        .CK(npu_inst_pe_1_1_0_net4384), .RN(npu_inst_pe_1_1_0_n10), .Q(
        npu_inst_pe_1_1_0_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_1_0_n88), 
        .CK(npu_inst_pe_1_1_0_net4384), .RN(npu_inst_pe_1_1_0_n11), .Q(
        npu_inst_pe_1_1_0_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_1_0_n89), 
        .CK(npu_inst_pe_1_1_0_net4384), .RN(npu_inst_pe_1_1_0_n11), .Q(
        npu_inst_pe_1_1_0_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_1_0_n90), 
        .CK(npu_inst_pe_1_1_0_net4384), .RN(npu_inst_pe_1_1_0_n11), .Q(
        npu_inst_pe_1_1_0_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_1_0_n91), 
        .CK(npu_inst_pe_1_1_0_net4384), .RN(npu_inst_pe_1_1_0_n11), .Q(
        npu_inst_pe_1_1_0_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_1_0_n92), 
        .CK(npu_inst_pe_1_1_0_net4384), .RN(npu_inst_pe_1_1_0_n11), .Q(
        npu_inst_pe_1_1_0_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_1_0_n93), 
        .CK(npu_inst_pe_1_1_0_net4384), .RN(npu_inst_pe_1_1_0_n11), .Q(
        npu_inst_pe_1_1_0_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_1_0_n94), 
        .CK(npu_inst_pe_1_1_0_net4384), .RN(npu_inst_pe_1_1_0_n11), .Q(
        npu_inst_pe_1_1_0_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_1_0_n95), 
        .CK(npu_inst_pe_1_1_0_net4384), .RN(npu_inst_pe_1_1_0_n11), .Q(
        npu_inst_pe_1_1_0_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_1_0_n96), 
        .CK(npu_inst_pe_1_1_0_net4384), .RN(npu_inst_pe_1_1_0_n11), .Q(
        npu_inst_pe_1_1_0_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_1_0_n97), 
        .CK(npu_inst_pe_1_1_0_net4384), .RN(npu_inst_pe_1_1_0_n11), .Q(
        npu_inst_pe_1_1_0_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_1_0_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_1_0_N84), .SE(1'b0), .GCK(npu_inst_pe_1_1_0_net4378) );
  CLKGATETST_X1 npu_inst_pe_1_1_0_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n66), .SE(1'b0), .GCK(npu_inst_pe_1_1_0_net4384) );
  MUX2_X1 npu_inst_pe_1_1_1_U162 ( .A(npu_inst_pe_1_1_1_n32), .B(
        npu_inst_pe_1_1_1_n29), .S(npu_inst_pe_1_1_1_n8), .Z(
        npu_inst_pe_1_1_1_N93) );
  MUX2_X1 npu_inst_pe_1_1_1_U161 ( .A(npu_inst_pe_1_1_1_n31), .B(
        npu_inst_pe_1_1_1_n30), .S(npu_inst_pe_1_1_1_n6), .Z(
        npu_inst_pe_1_1_1_n32) );
  MUX2_X1 npu_inst_pe_1_1_1_U160 ( .A(npu_inst_pe_1_1_1_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_1_1_int_q_reg_v_1__0_), .S(npu_inst_pe_1_1_1_n4), .Z(
        npu_inst_pe_1_1_1_n31) );
  MUX2_X1 npu_inst_pe_1_1_1_U159 ( .A(npu_inst_pe_1_1_1_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_1_1_int_q_reg_v_3__0_), .S(npu_inst_pe_1_1_1_n4), .Z(
        npu_inst_pe_1_1_1_n30) );
  MUX2_X1 npu_inst_pe_1_1_1_U158 ( .A(npu_inst_pe_1_1_1_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_1_1_int_q_reg_v_5__0_), .S(npu_inst_pe_1_1_1_n4), .Z(
        npu_inst_pe_1_1_1_n29) );
  MUX2_X1 npu_inst_pe_1_1_1_U157 ( .A(npu_inst_pe_1_1_1_n28), .B(
        npu_inst_pe_1_1_1_n23), .S(npu_inst_pe_1_1_1_n8), .Z(
        npu_inst_pe_1_1_1_N94) );
  MUX2_X1 npu_inst_pe_1_1_1_U156 ( .A(npu_inst_pe_1_1_1_n25), .B(
        npu_inst_pe_1_1_1_n24), .S(npu_inst_pe_1_1_1_n6), .Z(
        npu_inst_pe_1_1_1_n28) );
  MUX2_X1 npu_inst_pe_1_1_1_U155 ( .A(npu_inst_pe_1_1_1_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_1_1_int_q_reg_v_1__1_), .S(npu_inst_pe_1_1_1_n4), .Z(
        npu_inst_pe_1_1_1_n25) );
  MUX2_X1 npu_inst_pe_1_1_1_U154 ( .A(npu_inst_pe_1_1_1_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_1_1_int_q_reg_v_3__1_), .S(npu_inst_pe_1_1_1_n4), .Z(
        npu_inst_pe_1_1_1_n24) );
  MUX2_X1 npu_inst_pe_1_1_1_U153 ( .A(npu_inst_pe_1_1_1_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_1_1_int_q_reg_v_5__1_), .S(npu_inst_pe_1_1_1_n4), .Z(
        npu_inst_pe_1_1_1_n23) );
  MUX2_X1 npu_inst_pe_1_1_1_U152 ( .A(npu_inst_pe_1_1_1_n22), .B(
        npu_inst_pe_1_1_1_n19), .S(npu_inst_pe_1_1_1_n8), .Z(
        npu_inst_int_data_x_1__1__1_) );
  MUX2_X1 npu_inst_pe_1_1_1_U151 ( .A(npu_inst_pe_1_1_1_n21), .B(
        npu_inst_pe_1_1_1_n20), .S(npu_inst_pe_1_1_1_n6), .Z(
        npu_inst_pe_1_1_1_n22) );
  MUX2_X1 npu_inst_pe_1_1_1_U150 ( .A(npu_inst_pe_1_1_1_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_1_1_int_q_reg_h_1__1_), .S(npu_inst_pe_1_1_1_n4), .Z(
        npu_inst_pe_1_1_1_n21) );
  MUX2_X1 npu_inst_pe_1_1_1_U149 ( .A(npu_inst_pe_1_1_1_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_1_1_int_q_reg_h_3__1_), .S(npu_inst_pe_1_1_1_n4), .Z(
        npu_inst_pe_1_1_1_n20) );
  MUX2_X1 npu_inst_pe_1_1_1_U148 ( .A(npu_inst_pe_1_1_1_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_1_1_int_q_reg_h_5__1_), .S(npu_inst_pe_1_1_1_n4), .Z(
        npu_inst_pe_1_1_1_n19) );
  MUX2_X1 npu_inst_pe_1_1_1_U147 ( .A(npu_inst_pe_1_1_1_n18), .B(
        npu_inst_pe_1_1_1_n15), .S(npu_inst_pe_1_1_1_n8), .Z(
        npu_inst_int_data_x_1__1__0_) );
  MUX2_X1 npu_inst_pe_1_1_1_U146 ( .A(npu_inst_pe_1_1_1_n17), .B(
        npu_inst_pe_1_1_1_n16), .S(npu_inst_pe_1_1_1_n6), .Z(
        npu_inst_pe_1_1_1_n18) );
  MUX2_X1 npu_inst_pe_1_1_1_U145 ( .A(npu_inst_pe_1_1_1_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_1_1_int_q_reg_h_1__0_), .S(npu_inst_pe_1_1_1_n4), .Z(
        npu_inst_pe_1_1_1_n17) );
  MUX2_X1 npu_inst_pe_1_1_1_U144 ( .A(npu_inst_pe_1_1_1_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_1_1_int_q_reg_h_3__0_), .S(npu_inst_pe_1_1_1_n4), .Z(
        npu_inst_pe_1_1_1_n16) );
  MUX2_X1 npu_inst_pe_1_1_1_U143 ( .A(npu_inst_pe_1_1_1_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_1_1_int_q_reg_h_5__0_), .S(npu_inst_pe_1_1_1_n4), .Z(
        npu_inst_pe_1_1_1_n15) );
  XOR2_X1 npu_inst_pe_1_1_1_U142 ( .A(npu_inst_pe_1_1_1_int_data_0_), .B(
        npu_inst_pe_1_1_1_int_q_acc_0_), .Z(npu_inst_pe_1_1_1_N73) );
  AND2_X1 npu_inst_pe_1_1_1_U141 ( .A1(npu_inst_pe_1_1_1_int_q_acc_0_), .A2(
        npu_inst_pe_1_1_1_int_data_0_), .ZN(npu_inst_pe_1_1_1_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_1_1_U140 ( .A(npu_inst_pe_1_1_1_int_q_acc_0_), .B(
        npu_inst_pe_1_1_1_n13), .ZN(npu_inst_pe_1_1_1_N65) );
  OR2_X1 npu_inst_pe_1_1_1_U139 ( .A1(npu_inst_pe_1_1_1_n13), .A2(
        npu_inst_pe_1_1_1_int_q_acc_0_), .ZN(npu_inst_pe_1_1_1_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_1_1_U138 ( .A(npu_inst_pe_1_1_1_int_q_acc_2_), .B(
        npu_inst_pe_1_1_1_add_69_carry_2_), .Z(npu_inst_pe_1_1_1_N75) );
  AND2_X1 npu_inst_pe_1_1_1_U137 ( .A1(npu_inst_pe_1_1_1_add_69_carry_2_), 
        .A2(npu_inst_pe_1_1_1_int_q_acc_2_), .ZN(
        npu_inst_pe_1_1_1_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_1_1_U136 ( .A(npu_inst_pe_1_1_1_int_q_acc_3_), .B(
        npu_inst_pe_1_1_1_add_69_carry_3_), .Z(npu_inst_pe_1_1_1_N76) );
  AND2_X1 npu_inst_pe_1_1_1_U135 ( .A1(npu_inst_pe_1_1_1_add_69_carry_3_), 
        .A2(npu_inst_pe_1_1_1_int_q_acc_3_), .ZN(
        npu_inst_pe_1_1_1_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_1_1_U134 ( .A(npu_inst_pe_1_1_1_int_q_acc_4_), .B(
        npu_inst_pe_1_1_1_add_69_carry_4_), .Z(npu_inst_pe_1_1_1_N77) );
  AND2_X1 npu_inst_pe_1_1_1_U133 ( .A1(npu_inst_pe_1_1_1_add_69_carry_4_), 
        .A2(npu_inst_pe_1_1_1_int_q_acc_4_), .ZN(
        npu_inst_pe_1_1_1_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_1_1_U132 ( .A(npu_inst_pe_1_1_1_int_q_acc_5_), .B(
        npu_inst_pe_1_1_1_add_69_carry_5_), .Z(npu_inst_pe_1_1_1_N78) );
  AND2_X1 npu_inst_pe_1_1_1_U131 ( .A1(npu_inst_pe_1_1_1_add_69_carry_5_), 
        .A2(npu_inst_pe_1_1_1_int_q_acc_5_), .ZN(
        npu_inst_pe_1_1_1_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_1_1_U130 ( .A(npu_inst_pe_1_1_1_int_q_acc_6_), .B(
        npu_inst_pe_1_1_1_add_69_carry_6_), .Z(npu_inst_pe_1_1_1_N79) );
  AND2_X1 npu_inst_pe_1_1_1_U129 ( .A1(npu_inst_pe_1_1_1_add_69_carry_6_), 
        .A2(npu_inst_pe_1_1_1_int_q_acc_6_), .ZN(
        npu_inst_pe_1_1_1_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_1_1_U128 ( .A(npu_inst_pe_1_1_1_int_q_acc_7_), .B(
        npu_inst_pe_1_1_1_add_69_carry_7_), .Z(npu_inst_pe_1_1_1_N80) );
  XNOR2_X1 npu_inst_pe_1_1_1_U127 ( .A(npu_inst_pe_1_1_1_sub_67_carry_2_), .B(
        npu_inst_pe_1_1_1_int_q_acc_2_), .ZN(npu_inst_pe_1_1_1_N67) );
  OR2_X1 npu_inst_pe_1_1_1_U126 ( .A1(npu_inst_pe_1_1_1_int_q_acc_2_), .A2(
        npu_inst_pe_1_1_1_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_1_1_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_1_1_U125 ( .A(npu_inst_pe_1_1_1_sub_67_carry_3_), .B(
        npu_inst_pe_1_1_1_int_q_acc_3_), .ZN(npu_inst_pe_1_1_1_N68) );
  OR2_X1 npu_inst_pe_1_1_1_U124 ( .A1(npu_inst_pe_1_1_1_int_q_acc_3_), .A2(
        npu_inst_pe_1_1_1_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_1_1_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_1_1_U123 ( .A(npu_inst_pe_1_1_1_sub_67_carry_4_), .B(
        npu_inst_pe_1_1_1_int_q_acc_4_), .ZN(npu_inst_pe_1_1_1_N69) );
  OR2_X1 npu_inst_pe_1_1_1_U122 ( .A1(npu_inst_pe_1_1_1_int_q_acc_4_), .A2(
        npu_inst_pe_1_1_1_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_1_1_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_1_1_U121 ( .A(npu_inst_pe_1_1_1_sub_67_carry_5_), .B(
        npu_inst_pe_1_1_1_int_q_acc_5_), .ZN(npu_inst_pe_1_1_1_N70) );
  OR2_X1 npu_inst_pe_1_1_1_U120 ( .A1(npu_inst_pe_1_1_1_int_q_acc_5_), .A2(
        npu_inst_pe_1_1_1_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_1_1_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_1_1_U119 ( .A(npu_inst_pe_1_1_1_sub_67_carry_6_), .B(
        npu_inst_pe_1_1_1_int_q_acc_6_), .ZN(npu_inst_pe_1_1_1_N71) );
  OR2_X1 npu_inst_pe_1_1_1_U118 ( .A1(npu_inst_pe_1_1_1_int_q_acc_6_), .A2(
        npu_inst_pe_1_1_1_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_1_1_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_1_1_U117 ( .A(npu_inst_pe_1_1_1_int_q_acc_7_), .B(
        npu_inst_pe_1_1_1_sub_67_carry_7_), .ZN(npu_inst_pe_1_1_1_N72) );
  INV_X1 npu_inst_pe_1_1_1_U116 ( .A(npu_inst_n79), .ZN(npu_inst_pe_1_1_1_n7)
         );
  INV_X1 npu_inst_pe_1_1_1_U115 ( .A(npu_inst_pe_1_1_1_n7), .ZN(
        npu_inst_pe_1_1_1_n6) );
  INV_X1 npu_inst_pe_1_1_1_U114 ( .A(npu_inst_n59), .ZN(npu_inst_pe_1_1_1_n3)
         );
  AOI22_X1 npu_inst_pe_1_1_1_U113 ( .A1(npu_inst_int_data_y_2__1__0_), .A2(
        npu_inst_pe_1_1_1_n58), .B1(npu_inst_pe_1_1_1_n119), .B2(
        npu_inst_pe_1_1_1_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_1_1_n57) );
  INV_X1 npu_inst_pe_1_1_1_U112 ( .A(npu_inst_pe_1_1_1_n57), .ZN(
        npu_inst_pe_1_1_1_n108) );
  AOI22_X1 npu_inst_pe_1_1_1_U111 ( .A1(npu_inst_int_data_y_2__1__0_), .A2(
        npu_inst_pe_1_1_1_n54), .B1(npu_inst_pe_1_1_1_n118), .B2(
        npu_inst_pe_1_1_1_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_1_1_n53) );
  INV_X1 npu_inst_pe_1_1_1_U110 ( .A(npu_inst_pe_1_1_1_n53), .ZN(
        npu_inst_pe_1_1_1_n109) );
  AOI22_X1 npu_inst_pe_1_1_1_U107 ( .A1(npu_inst_int_data_y_2__1__0_), .A2(
        npu_inst_pe_1_1_1_n50), .B1(npu_inst_pe_1_1_1_n117), .B2(
        npu_inst_pe_1_1_1_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_1_1_n49) );
  INV_X1 npu_inst_pe_1_1_1_U106 ( .A(npu_inst_pe_1_1_1_n49), .ZN(
        npu_inst_pe_1_1_1_n110) );
  AOI22_X1 npu_inst_pe_1_1_1_U105 ( .A1(npu_inst_int_data_y_2__1__0_), .A2(
        npu_inst_pe_1_1_1_n46), .B1(npu_inst_pe_1_1_1_n116), .B2(
        npu_inst_pe_1_1_1_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_1_1_n45) );
  INV_X1 npu_inst_pe_1_1_1_U104 ( .A(npu_inst_pe_1_1_1_n45), .ZN(
        npu_inst_pe_1_1_1_n111) );
  AOI22_X1 npu_inst_pe_1_1_1_U103 ( .A1(npu_inst_int_data_y_2__1__0_), .A2(
        npu_inst_pe_1_1_1_n42), .B1(npu_inst_pe_1_1_1_n115), .B2(
        npu_inst_pe_1_1_1_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_1_1_n41) );
  INV_X1 npu_inst_pe_1_1_1_U102 ( .A(npu_inst_pe_1_1_1_n41), .ZN(
        npu_inst_pe_1_1_1_n112) );
  AOI22_X1 npu_inst_pe_1_1_1_U101 ( .A1(npu_inst_int_data_y_2__1__1_), .A2(
        npu_inst_pe_1_1_1_n58), .B1(npu_inst_pe_1_1_1_n119), .B2(
        npu_inst_pe_1_1_1_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_1_1_n59) );
  INV_X1 npu_inst_pe_1_1_1_U100 ( .A(npu_inst_pe_1_1_1_n59), .ZN(
        npu_inst_pe_1_1_1_n102) );
  AOI22_X1 npu_inst_pe_1_1_1_U99 ( .A1(npu_inst_int_data_y_2__1__1_), .A2(
        npu_inst_pe_1_1_1_n54), .B1(npu_inst_pe_1_1_1_n118), .B2(
        npu_inst_pe_1_1_1_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_1_1_n55) );
  INV_X1 npu_inst_pe_1_1_1_U98 ( .A(npu_inst_pe_1_1_1_n55), .ZN(
        npu_inst_pe_1_1_1_n103) );
  AOI22_X1 npu_inst_pe_1_1_1_U97 ( .A1(npu_inst_int_data_y_2__1__1_), .A2(
        npu_inst_pe_1_1_1_n50), .B1(npu_inst_pe_1_1_1_n117), .B2(
        npu_inst_pe_1_1_1_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_1_1_n51) );
  INV_X1 npu_inst_pe_1_1_1_U96 ( .A(npu_inst_pe_1_1_1_n51), .ZN(
        npu_inst_pe_1_1_1_n104) );
  AOI22_X1 npu_inst_pe_1_1_1_U95 ( .A1(npu_inst_int_data_y_2__1__1_), .A2(
        npu_inst_pe_1_1_1_n46), .B1(npu_inst_pe_1_1_1_n116), .B2(
        npu_inst_pe_1_1_1_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_1_1_n47) );
  INV_X1 npu_inst_pe_1_1_1_U94 ( .A(npu_inst_pe_1_1_1_n47), .ZN(
        npu_inst_pe_1_1_1_n105) );
  AOI22_X1 npu_inst_pe_1_1_1_U93 ( .A1(npu_inst_int_data_y_2__1__1_), .A2(
        npu_inst_pe_1_1_1_n42), .B1(npu_inst_pe_1_1_1_n115), .B2(
        npu_inst_pe_1_1_1_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_1_1_n43) );
  INV_X1 npu_inst_pe_1_1_1_U92 ( .A(npu_inst_pe_1_1_1_n43), .ZN(
        npu_inst_pe_1_1_1_n106) );
  AOI22_X1 npu_inst_pe_1_1_1_U91 ( .A1(npu_inst_pe_1_1_1_n38), .A2(
        npu_inst_int_data_y_2__1__1_), .B1(npu_inst_pe_1_1_1_n114), .B2(
        npu_inst_pe_1_1_1_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_1_1_n39) );
  INV_X1 npu_inst_pe_1_1_1_U90 ( .A(npu_inst_pe_1_1_1_n39), .ZN(
        npu_inst_pe_1_1_1_n107) );
  AOI22_X1 npu_inst_pe_1_1_1_U89 ( .A1(npu_inst_pe_1_1_1_n38), .A2(
        npu_inst_int_data_y_2__1__0_), .B1(npu_inst_pe_1_1_1_n114), .B2(
        npu_inst_pe_1_1_1_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_1_1_n37) );
  INV_X1 npu_inst_pe_1_1_1_U88 ( .A(npu_inst_pe_1_1_1_n37), .ZN(
        npu_inst_pe_1_1_1_n113) );
  NAND2_X1 npu_inst_pe_1_1_1_U87 ( .A1(npu_inst_pe_1_1_1_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_1_1_n60), .ZN(npu_inst_pe_1_1_1_n74) );
  OAI21_X1 npu_inst_pe_1_1_1_U86 ( .B1(npu_inst_pe_1_1_1_n63), .B2(
        npu_inst_pe_1_1_1_n60), .A(npu_inst_pe_1_1_1_n74), .ZN(
        npu_inst_pe_1_1_1_n97) );
  NAND2_X1 npu_inst_pe_1_1_1_U85 ( .A1(npu_inst_pe_1_1_1_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_1_1_n60), .ZN(npu_inst_pe_1_1_1_n73) );
  OAI21_X1 npu_inst_pe_1_1_1_U84 ( .B1(npu_inst_pe_1_1_1_n61), .B2(
        npu_inst_pe_1_1_1_n60), .A(npu_inst_pe_1_1_1_n73), .ZN(
        npu_inst_pe_1_1_1_n96) );
  NAND2_X1 npu_inst_pe_1_1_1_U83 ( .A1(npu_inst_pe_1_1_1_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_1_1_n56), .ZN(npu_inst_pe_1_1_1_n72) );
  OAI21_X1 npu_inst_pe_1_1_1_U82 ( .B1(npu_inst_pe_1_1_1_n63), .B2(
        npu_inst_pe_1_1_1_n56), .A(npu_inst_pe_1_1_1_n72), .ZN(
        npu_inst_pe_1_1_1_n95) );
  NAND2_X1 npu_inst_pe_1_1_1_U81 ( .A1(npu_inst_pe_1_1_1_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_1_1_n56), .ZN(npu_inst_pe_1_1_1_n71) );
  OAI21_X1 npu_inst_pe_1_1_1_U80 ( .B1(npu_inst_pe_1_1_1_n61), .B2(
        npu_inst_pe_1_1_1_n56), .A(npu_inst_pe_1_1_1_n71), .ZN(
        npu_inst_pe_1_1_1_n94) );
  NAND2_X1 npu_inst_pe_1_1_1_U79 ( .A1(npu_inst_pe_1_1_1_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_1_1_n52), .ZN(npu_inst_pe_1_1_1_n70) );
  OAI21_X1 npu_inst_pe_1_1_1_U78 ( .B1(npu_inst_pe_1_1_1_n63), .B2(
        npu_inst_pe_1_1_1_n52), .A(npu_inst_pe_1_1_1_n70), .ZN(
        npu_inst_pe_1_1_1_n93) );
  NAND2_X1 npu_inst_pe_1_1_1_U77 ( .A1(npu_inst_pe_1_1_1_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_1_1_n52), .ZN(npu_inst_pe_1_1_1_n69) );
  OAI21_X1 npu_inst_pe_1_1_1_U76 ( .B1(npu_inst_pe_1_1_1_n61), .B2(
        npu_inst_pe_1_1_1_n52), .A(npu_inst_pe_1_1_1_n69), .ZN(
        npu_inst_pe_1_1_1_n92) );
  NAND2_X1 npu_inst_pe_1_1_1_U75 ( .A1(npu_inst_pe_1_1_1_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_1_1_n48), .ZN(npu_inst_pe_1_1_1_n68) );
  OAI21_X1 npu_inst_pe_1_1_1_U74 ( .B1(npu_inst_pe_1_1_1_n63), .B2(
        npu_inst_pe_1_1_1_n48), .A(npu_inst_pe_1_1_1_n68), .ZN(
        npu_inst_pe_1_1_1_n91) );
  NAND2_X1 npu_inst_pe_1_1_1_U73 ( .A1(npu_inst_pe_1_1_1_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_1_1_n48), .ZN(npu_inst_pe_1_1_1_n67) );
  OAI21_X1 npu_inst_pe_1_1_1_U72 ( .B1(npu_inst_pe_1_1_1_n61), .B2(
        npu_inst_pe_1_1_1_n48), .A(npu_inst_pe_1_1_1_n67), .ZN(
        npu_inst_pe_1_1_1_n90) );
  NAND2_X1 npu_inst_pe_1_1_1_U71 ( .A1(npu_inst_pe_1_1_1_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_1_1_n44), .ZN(npu_inst_pe_1_1_1_n66) );
  OAI21_X1 npu_inst_pe_1_1_1_U70 ( .B1(npu_inst_pe_1_1_1_n63), .B2(
        npu_inst_pe_1_1_1_n44), .A(npu_inst_pe_1_1_1_n66), .ZN(
        npu_inst_pe_1_1_1_n89) );
  NAND2_X1 npu_inst_pe_1_1_1_U69 ( .A1(npu_inst_pe_1_1_1_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_1_1_n44), .ZN(npu_inst_pe_1_1_1_n65) );
  OAI21_X1 npu_inst_pe_1_1_1_U68 ( .B1(npu_inst_pe_1_1_1_n61), .B2(
        npu_inst_pe_1_1_1_n44), .A(npu_inst_pe_1_1_1_n65), .ZN(
        npu_inst_pe_1_1_1_n88) );
  NAND2_X1 npu_inst_pe_1_1_1_U67 ( .A1(npu_inst_pe_1_1_1_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_1_1_n40), .ZN(npu_inst_pe_1_1_1_n64) );
  OAI21_X1 npu_inst_pe_1_1_1_U66 ( .B1(npu_inst_pe_1_1_1_n63), .B2(
        npu_inst_pe_1_1_1_n40), .A(npu_inst_pe_1_1_1_n64), .ZN(
        npu_inst_pe_1_1_1_n87) );
  NAND2_X1 npu_inst_pe_1_1_1_U65 ( .A1(npu_inst_pe_1_1_1_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_1_1_n40), .ZN(npu_inst_pe_1_1_1_n62) );
  OAI21_X1 npu_inst_pe_1_1_1_U64 ( .B1(npu_inst_pe_1_1_1_n61), .B2(
        npu_inst_pe_1_1_1_n40), .A(npu_inst_pe_1_1_1_n62), .ZN(
        npu_inst_pe_1_1_1_n86) );
  AND2_X1 npu_inst_pe_1_1_1_U63 ( .A1(npu_inst_pe_1_1_1_N93), .A2(npu_inst_n59), .ZN(npu_inst_int_data_y_1__1__0_) );
  AND2_X1 npu_inst_pe_1_1_1_U62 ( .A1(npu_inst_n59), .A2(npu_inst_pe_1_1_1_N94), .ZN(npu_inst_int_data_y_1__1__1_) );
  NOR3_X1 npu_inst_pe_1_1_1_U61 ( .A1(npu_inst_pe_1_1_1_n26), .A2(npu_inst_n59), .A3(npu_inst_int_ckg[54]), .ZN(npu_inst_pe_1_1_1_n85) );
  OR2_X1 npu_inst_pe_1_1_1_U60 ( .A1(npu_inst_pe_1_1_1_n85), .A2(
        npu_inst_pe_1_1_1_n2), .ZN(npu_inst_pe_1_1_1_N84) );
  AND2_X1 npu_inst_pe_1_1_1_U59 ( .A1(npu_inst_pe_1_1_1_int_q_acc_0_), .A2(
        npu_inst_pe_1_1_1_n1), .ZN(npu_inst_int_data_res_1__1__0_) );
  AND2_X1 npu_inst_pe_1_1_1_U58 ( .A1(npu_inst_pe_1_1_1_n2), .A2(
        npu_inst_pe_1_1_1_int_q_acc_7_), .ZN(npu_inst_int_data_res_1__1__7_)
         );
  AND2_X1 npu_inst_pe_1_1_1_U57 ( .A1(npu_inst_pe_1_1_1_int_q_acc_1_), .A2(
        npu_inst_pe_1_1_1_n1), .ZN(npu_inst_int_data_res_1__1__1_) );
  AND2_X1 npu_inst_pe_1_1_1_U56 ( .A1(npu_inst_pe_1_1_1_int_q_acc_2_), .A2(
        npu_inst_pe_1_1_1_n1), .ZN(npu_inst_int_data_res_1__1__2_) );
  AND2_X1 npu_inst_pe_1_1_1_U55 ( .A1(npu_inst_pe_1_1_1_int_q_acc_3_), .A2(
        npu_inst_pe_1_1_1_n2), .ZN(npu_inst_int_data_res_1__1__3_) );
  AND2_X1 npu_inst_pe_1_1_1_U54 ( .A1(npu_inst_pe_1_1_1_int_q_acc_4_), .A2(
        npu_inst_pe_1_1_1_n2), .ZN(npu_inst_int_data_res_1__1__4_) );
  AND2_X1 npu_inst_pe_1_1_1_U53 ( .A1(npu_inst_pe_1_1_1_int_q_acc_5_), .A2(
        npu_inst_pe_1_1_1_n2), .ZN(npu_inst_int_data_res_1__1__5_) );
  AND2_X1 npu_inst_pe_1_1_1_U52 ( .A1(npu_inst_pe_1_1_1_int_q_acc_6_), .A2(
        npu_inst_pe_1_1_1_n2), .ZN(npu_inst_int_data_res_1__1__6_) );
  AOI222_X1 npu_inst_pe_1_1_1_U51 ( .A1(npu_inst_int_data_res_2__1__0_), .A2(
        npu_inst_pe_1_1_1_n1), .B1(npu_inst_pe_1_1_1_N73), .B2(
        npu_inst_pe_1_1_1_n76), .C1(npu_inst_pe_1_1_1_N65), .C2(
        npu_inst_pe_1_1_1_n77), .ZN(npu_inst_pe_1_1_1_n84) );
  INV_X1 npu_inst_pe_1_1_1_U50 ( .A(npu_inst_pe_1_1_1_n84), .ZN(
        npu_inst_pe_1_1_1_n101) );
  AOI222_X1 npu_inst_pe_1_1_1_U49 ( .A1(npu_inst_int_data_res_2__1__7_), .A2(
        npu_inst_pe_1_1_1_n1), .B1(npu_inst_pe_1_1_1_N80), .B2(
        npu_inst_pe_1_1_1_n76), .C1(npu_inst_pe_1_1_1_N72), .C2(
        npu_inst_pe_1_1_1_n77), .ZN(npu_inst_pe_1_1_1_n75) );
  INV_X1 npu_inst_pe_1_1_1_U48 ( .A(npu_inst_pe_1_1_1_n75), .ZN(
        npu_inst_pe_1_1_1_n33) );
  AOI222_X1 npu_inst_pe_1_1_1_U47 ( .A1(npu_inst_int_data_res_2__1__1_), .A2(
        npu_inst_pe_1_1_1_n1), .B1(npu_inst_pe_1_1_1_N74), .B2(
        npu_inst_pe_1_1_1_n76), .C1(npu_inst_pe_1_1_1_N66), .C2(
        npu_inst_pe_1_1_1_n77), .ZN(npu_inst_pe_1_1_1_n83) );
  INV_X1 npu_inst_pe_1_1_1_U46 ( .A(npu_inst_pe_1_1_1_n83), .ZN(
        npu_inst_pe_1_1_1_n100) );
  AOI222_X1 npu_inst_pe_1_1_1_U45 ( .A1(npu_inst_int_data_res_2__1__2_), .A2(
        npu_inst_pe_1_1_1_n1), .B1(npu_inst_pe_1_1_1_N75), .B2(
        npu_inst_pe_1_1_1_n76), .C1(npu_inst_pe_1_1_1_N67), .C2(
        npu_inst_pe_1_1_1_n77), .ZN(npu_inst_pe_1_1_1_n82) );
  INV_X1 npu_inst_pe_1_1_1_U44 ( .A(npu_inst_pe_1_1_1_n82), .ZN(
        npu_inst_pe_1_1_1_n99) );
  AOI222_X1 npu_inst_pe_1_1_1_U43 ( .A1(npu_inst_int_data_res_2__1__3_), .A2(
        npu_inst_pe_1_1_1_n1), .B1(npu_inst_pe_1_1_1_N76), .B2(
        npu_inst_pe_1_1_1_n76), .C1(npu_inst_pe_1_1_1_N68), .C2(
        npu_inst_pe_1_1_1_n77), .ZN(npu_inst_pe_1_1_1_n81) );
  INV_X1 npu_inst_pe_1_1_1_U42 ( .A(npu_inst_pe_1_1_1_n81), .ZN(
        npu_inst_pe_1_1_1_n98) );
  AOI222_X1 npu_inst_pe_1_1_1_U41 ( .A1(npu_inst_int_data_res_2__1__4_), .A2(
        npu_inst_pe_1_1_1_n1), .B1(npu_inst_pe_1_1_1_N77), .B2(
        npu_inst_pe_1_1_1_n76), .C1(npu_inst_pe_1_1_1_N69), .C2(
        npu_inst_pe_1_1_1_n77), .ZN(npu_inst_pe_1_1_1_n80) );
  INV_X1 npu_inst_pe_1_1_1_U40 ( .A(npu_inst_pe_1_1_1_n80), .ZN(
        npu_inst_pe_1_1_1_n36) );
  AOI222_X1 npu_inst_pe_1_1_1_U39 ( .A1(npu_inst_int_data_res_2__1__5_), .A2(
        npu_inst_pe_1_1_1_n1), .B1(npu_inst_pe_1_1_1_N78), .B2(
        npu_inst_pe_1_1_1_n76), .C1(npu_inst_pe_1_1_1_N70), .C2(
        npu_inst_pe_1_1_1_n77), .ZN(npu_inst_pe_1_1_1_n79) );
  INV_X1 npu_inst_pe_1_1_1_U38 ( .A(npu_inst_pe_1_1_1_n79), .ZN(
        npu_inst_pe_1_1_1_n35) );
  AOI222_X1 npu_inst_pe_1_1_1_U37 ( .A1(npu_inst_int_data_res_2__1__6_), .A2(
        npu_inst_pe_1_1_1_n1), .B1(npu_inst_pe_1_1_1_N79), .B2(
        npu_inst_pe_1_1_1_n76), .C1(npu_inst_pe_1_1_1_N71), .C2(
        npu_inst_pe_1_1_1_n77), .ZN(npu_inst_pe_1_1_1_n78) );
  INV_X1 npu_inst_pe_1_1_1_U36 ( .A(npu_inst_pe_1_1_1_n78), .ZN(
        npu_inst_pe_1_1_1_n34) );
  INV_X1 npu_inst_pe_1_1_1_U35 ( .A(npu_inst_pe_1_1_1_int_data_1_), .ZN(
        npu_inst_pe_1_1_1_n14) );
  AND2_X1 npu_inst_pe_1_1_1_U34 ( .A1(npu_inst_int_data_x_1__1__1_), .A2(
        npu_inst_pe_1_1_1_int_q_weight_1_), .ZN(npu_inst_pe_1_1_1_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_1_1_U33 ( .A1(npu_inst_int_data_x_1__1__0_), .A2(
        npu_inst_pe_1_1_1_int_q_weight_1_), .ZN(npu_inst_pe_1_1_1_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_1_1_U32 ( .A1(npu_inst_n59), .A2(
        npu_inst_int_data_y_2__1__1_), .B1(npu_inst_pe_1_1_1_n3), .B2(
        npu_inst_int_data_x_1__2__1_), .ZN(npu_inst_pe_1_1_1_n63) );
  AOI22_X1 npu_inst_pe_1_1_1_U31 ( .A1(npu_inst_n59), .A2(
        npu_inst_int_data_y_2__1__0_), .B1(npu_inst_pe_1_1_1_n3), .B2(
        npu_inst_int_data_x_1__2__0_), .ZN(npu_inst_pe_1_1_1_n61) );
  INV_X1 npu_inst_pe_1_1_1_U30 ( .A(npu_inst_pe_1_1_1_int_data_0_), .ZN(
        npu_inst_pe_1_1_1_n13) );
  INV_X1 npu_inst_pe_1_1_1_U29 ( .A(npu_inst_n71), .ZN(npu_inst_pe_1_1_1_n5)
         );
  OR3_X1 npu_inst_pe_1_1_1_U28 ( .A1(npu_inst_pe_1_1_1_n6), .A2(
        npu_inst_pe_1_1_1_n8), .A3(npu_inst_pe_1_1_1_n5), .ZN(
        npu_inst_pe_1_1_1_n56) );
  OR3_X1 npu_inst_pe_1_1_1_U27 ( .A1(npu_inst_pe_1_1_1_n5), .A2(
        npu_inst_pe_1_1_1_n8), .A3(npu_inst_pe_1_1_1_n7), .ZN(
        npu_inst_pe_1_1_1_n48) );
  INV_X1 npu_inst_pe_1_1_1_U26 ( .A(npu_inst_pe_1_1_1_n5), .ZN(
        npu_inst_pe_1_1_1_n4) );
  OR3_X1 npu_inst_pe_1_1_1_U25 ( .A1(npu_inst_pe_1_1_1_n4), .A2(
        npu_inst_pe_1_1_1_n8), .A3(npu_inst_pe_1_1_1_n7), .ZN(
        npu_inst_pe_1_1_1_n52) );
  OR3_X1 npu_inst_pe_1_1_1_U24 ( .A1(npu_inst_pe_1_1_1_n6), .A2(
        npu_inst_pe_1_1_1_n8), .A3(npu_inst_pe_1_1_1_n4), .ZN(
        npu_inst_pe_1_1_1_n60) );
  NOR2_X1 npu_inst_pe_1_1_1_U23 ( .A1(npu_inst_pe_1_1_1_n60), .A2(
        npu_inst_pe_1_1_1_n3), .ZN(npu_inst_pe_1_1_1_n58) );
  NOR2_X1 npu_inst_pe_1_1_1_U22 ( .A1(npu_inst_pe_1_1_1_n56), .A2(
        npu_inst_pe_1_1_1_n3), .ZN(npu_inst_pe_1_1_1_n54) );
  NOR2_X1 npu_inst_pe_1_1_1_U21 ( .A1(npu_inst_pe_1_1_1_n52), .A2(
        npu_inst_pe_1_1_1_n3), .ZN(npu_inst_pe_1_1_1_n50) );
  NOR2_X1 npu_inst_pe_1_1_1_U20 ( .A1(npu_inst_pe_1_1_1_n48), .A2(
        npu_inst_pe_1_1_1_n3), .ZN(npu_inst_pe_1_1_1_n46) );
  NOR2_X1 npu_inst_pe_1_1_1_U19 ( .A1(npu_inst_pe_1_1_1_n40), .A2(
        npu_inst_pe_1_1_1_n3), .ZN(npu_inst_pe_1_1_1_n38) );
  NOR2_X1 npu_inst_pe_1_1_1_U18 ( .A1(npu_inst_pe_1_1_1_n44), .A2(
        npu_inst_pe_1_1_1_n3), .ZN(npu_inst_pe_1_1_1_n42) );
  BUF_X1 npu_inst_pe_1_1_1_U17 ( .A(npu_inst_n105), .Z(npu_inst_pe_1_1_1_n8)
         );
  INV_X1 npu_inst_pe_1_1_1_U16 ( .A(npu_inst_n126), .ZN(npu_inst_pe_1_1_1_n12)
         );
  INV_X1 npu_inst_pe_1_1_1_U15 ( .A(npu_inst_pe_1_1_1_n38), .ZN(
        npu_inst_pe_1_1_1_n114) );
  INV_X1 npu_inst_pe_1_1_1_U14 ( .A(npu_inst_pe_1_1_1_n58), .ZN(
        npu_inst_pe_1_1_1_n119) );
  INV_X1 npu_inst_pe_1_1_1_U13 ( .A(npu_inst_pe_1_1_1_n54), .ZN(
        npu_inst_pe_1_1_1_n118) );
  INV_X1 npu_inst_pe_1_1_1_U12 ( .A(npu_inst_pe_1_1_1_n50), .ZN(
        npu_inst_pe_1_1_1_n117) );
  INV_X1 npu_inst_pe_1_1_1_U11 ( .A(npu_inst_pe_1_1_1_n46), .ZN(
        npu_inst_pe_1_1_1_n116) );
  INV_X1 npu_inst_pe_1_1_1_U10 ( .A(npu_inst_pe_1_1_1_n42), .ZN(
        npu_inst_pe_1_1_1_n115) );
  BUF_X1 npu_inst_pe_1_1_1_U9 ( .A(npu_inst_n34), .Z(npu_inst_pe_1_1_1_n2) );
  BUF_X1 npu_inst_pe_1_1_1_U8 ( .A(npu_inst_n34), .Z(npu_inst_pe_1_1_1_n1) );
  BUF_X1 npu_inst_pe_1_1_1_U7 ( .A(npu_inst_pe_1_1_1_n12), .Z(
        npu_inst_pe_1_1_1_n11) );
  BUF_X1 npu_inst_pe_1_1_1_U6 ( .A(npu_inst_pe_1_1_1_n12), .Z(
        npu_inst_pe_1_1_1_n10) );
  BUF_X1 npu_inst_pe_1_1_1_U5 ( .A(npu_inst_pe_1_1_1_n12), .Z(
        npu_inst_pe_1_1_1_n9) );
  NOR2_X1 npu_inst_pe_1_1_1_U4 ( .A1(npu_inst_pe_1_1_1_int_q_weight_0_), .A2(
        npu_inst_pe_1_1_1_n1), .ZN(npu_inst_pe_1_1_1_n76) );
  NOR2_X1 npu_inst_pe_1_1_1_U3 ( .A1(npu_inst_pe_1_1_1_n27), .A2(
        npu_inst_pe_1_1_1_n1), .ZN(npu_inst_pe_1_1_1_n77) );
  FA_X1 npu_inst_pe_1_1_1_sub_67_U2_1 ( .A(npu_inst_pe_1_1_1_int_q_acc_1_), 
        .B(npu_inst_pe_1_1_1_n14), .CI(npu_inst_pe_1_1_1_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_1_1_sub_67_carry_2_), .S(npu_inst_pe_1_1_1_N66) );
  FA_X1 npu_inst_pe_1_1_1_add_69_U1_1 ( .A(npu_inst_pe_1_1_1_int_q_acc_1_), 
        .B(npu_inst_pe_1_1_1_int_data_1_), .CI(
        npu_inst_pe_1_1_1_add_69_carry_1_), .CO(
        npu_inst_pe_1_1_1_add_69_carry_2_), .S(npu_inst_pe_1_1_1_N74) );
  NAND3_X1 npu_inst_pe_1_1_1_U109 ( .A1(npu_inst_pe_1_1_1_n5), .A2(
        npu_inst_pe_1_1_1_n7), .A3(npu_inst_pe_1_1_1_n8), .ZN(
        npu_inst_pe_1_1_1_n44) );
  NAND3_X1 npu_inst_pe_1_1_1_U108 ( .A1(npu_inst_pe_1_1_1_n4), .A2(
        npu_inst_pe_1_1_1_n7), .A3(npu_inst_pe_1_1_1_n8), .ZN(
        npu_inst_pe_1_1_1_n40) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_1_1_n34), .CK(
        npu_inst_pe_1_1_1_net4355), .RN(npu_inst_pe_1_1_1_n9), .Q(
        npu_inst_pe_1_1_1_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_1_1_n35), .CK(
        npu_inst_pe_1_1_1_net4355), .RN(npu_inst_pe_1_1_1_n9), .Q(
        npu_inst_pe_1_1_1_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_1_1_n36), .CK(
        npu_inst_pe_1_1_1_net4355), .RN(npu_inst_pe_1_1_1_n9), .Q(
        npu_inst_pe_1_1_1_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_1_1_n98), .CK(
        npu_inst_pe_1_1_1_net4355), .RN(npu_inst_pe_1_1_1_n9), .Q(
        npu_inst_pe_1_1_1_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_1_1_n99), .CK(
        npu_inst_pe_1_1_1_net4355), .RN(npu_inst_pe_1_1_1_n9), .Q(
        npu_inst_pe_1_1_1_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_1_1_n100), 
        .CK(npu_inst_pe_1_1_1_net4355), .RN(npu_inst_pe_1_1_1_n9), .Q(
        npu_inst_pe_1_1_1_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_1_1_n33), .CK(
        npu_inst_pe_1_1_1_net4355), .RN(npu_inst_pe_1_1_1_n9), .Q(
        npu_inst_pe_1_1_1_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_1_1_n101), 
        .CK(npu_inst_pe_1_1_1_net4355), .RN(npu_inst_pe_1_1_1_n9), .Q(
        npu_inst_pe_1_1_1_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_weight_reg_0_ ( .D(npu_inst_n112), .CK(
        npu_inst_pe_1_1_1_net4361), .RN(npu_inst_pe_1_1_1_n9), .Q(
        npu_inst_pe_1_1_1_int_q_weight_0_), .QN(npu_inst_pe_1_1_1_n27) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_weight_reg_1_ ( .D(npu_inst_n118), .CK(
        npu_inst_pe_1_1_1_net4361), .RN(npu_inst_pe_1_1_1_n9), .Q(
        npu_inst_pe_1_1_1_int_q_weight_1_), .QN(npu_inst_pe_1_1_1_n26) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_1_1_n113), 
        .CK(npu_inst_pe_1_1_1_net4361), .RN(npu_inst_pe_1_1_1_n9), .Q(
        npu_inst_pe_1_1_1_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_1_1_n107), 
        .CK(npu_inst_pe_1_1_1_net4361), .RN(npu_inst_pe_1_1_1_n9), .Q(
        npu_inst_pe_1_1_1_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_1_1_n112), 
        .CK(npu_inst_pe_1_1_1_net4361), .RN(npu_inst_pe_1_1_1_n10), .Q(
        npu_inst_pe_1_1_1_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_1_1_n106), 
        .CK(npu_inst_pe_1_1_1_net4361), .RN(npu_inst_pe_1_1_1_n10), .Q(
        npu_inst_pe_1_1_1_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_1_1_n111), 
        .CK(npu_inst_pe_1_1_1_net4361), .RN(npu_inst_pe_1_1_1_n10), .Q(
        npu_inst_pe_1_1_1_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_1_1_n105), 
        .CK(npu_inst_pe_1_1_1_net4361), .RN(npu_inst_pe_1_1_1_n10), .Q(
        npu_inst_pe_1_1_1_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_1_1_n110), 
        .CK(npu_inst_pe_1_1_1_net4361), .RN(npu_inst_pe_1_1_1_n10), .Q(
        npu_inst_pe_1_1_1_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_1_1_n104), 
        .CK(npu_inst_pe_1_1_1_net4361), .RN(npu_inst_pe_1_1_1_n10), .Q(
        npu_inst_pe_1_1_1_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_1_1_n109), 
        .CK(npu_inst_pe_1_1_1_net4361), .RN(npu_inst_pe_1_1_1_n10), .Q(
        npu_inst_pe_1_1_1_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_1_1_n103), 
        .CK(npu_inst_pe_1_1_1_net4361), .RN(npu_inst_pe_1_1_1_n10), .Q(
        npu_inst_pe_1_1_1_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_1_1_n108), 
        .CK(npu_inst_pe_1_1_1_net4361), .RN(npu_inst_pe_1_1_1_n10), .Q(
        npu_inst_pe_1_1_1_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_1_1_n102), 
        .CK(npu_inst_pe_1_1_1_net4361), .RN(npu_inst_pe_1_1_1_n10), .Q(
        npu_inst_pe_1_1_1_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_1_1_n86), 
        .CK(npu_inst_pe_1_1_1_net4361), .RN(npu_inst_pe_1_1_1_n10), .Q(
        npu_inst_pe_1_1_1_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_1_1_n87), 
        .CK(npu_inst_pe_1_1_1_net4361), .RN(npu_inst_pe_1_1_1_n10), .Q(
        npu_inst_pe_1_1_1_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_1_1_n88), 
        .CK(npu_inst_pe_1_1_1_net4361), .RN(npu_inst_pe_1_1_1_n11), .Q(
        npu_inst_pe_1_1_1_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_1_1_n89), 
        .CK(npu_inst_pe_1_1_1_net4361), .RN(npu_inst_pe_1_1_1_n11), .Q(
        npu_inst_pe_1_1_1_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_1_1_n90), 
        .CK(npu_inst_pe_1_1_1_net4361), .RN(npu_inst_pe_1_1_1_n11), .Q(
        npu_inst_pe_1_1_1_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_1_1_n91), 
        .CK(npu_inst_pe_1_1_1_net4361), .RN(npu_inst_pe_1_1_1_n11), .Q(
        npu_inst_pe_1_1_1_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_1_1_n92), 
        .CK(npu_inst_pe_1_1_1_net4361), .RN(npu_inst_pe_1_1_1_n11), .Q(
        npu_inst_pe_1_1_1_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_1_1_n93), 
        .CK(npu_inst_pe_1_1_1_net4361), .RN(npu_inst_pe_1_1_1_n11), .Q(
        npu_inst_pe_1_1_1_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_1_1_n94), 
        .CK(npu_inst_pe_1_1_1_net4361), .RN(npu_inst_pe_1_1_1_n11), .Q(
        npu_inst_pe_1_1_1_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_1_1_n95), 
        .CK(npu_inst_pe_1_1_1_net4361), .RN(npu_inst_pe_1_1_1_n11), .Q(
        npu_inst_pe_1_1_1_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_1_1_n96), 
        .CK(npu_inst_pe_1_1_1_net4361), .RN(npu_inst_pe_1_1_1_n11), .Q(
        npu_inst_pe_1_1_1_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_1_1_n97), 
        .CK(npu_inst_pe_1_1_1_net4361), .RN(npu_inst_pe_1_1_1_n11), .Q(
        npu_inst_pe_1_1_1_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_1_1_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_1_1_N84), .SE(1'b0), .GCK(npu_inst_pe_1_1_1_net4355) );
  CLKGATETST_X1 npu_inst_pe_1_1_1_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n65), .SE(1'b0), .GCK(npu_inst_pe_1_1_1_net4361) );
  MUX2_X1 npu_inst_pe_1_1_2_U162 ( .A(npu_inst_pe_1_1_2_n32), .B(
        npu_inst_pe_1_1_2_n29), .S(npu_inst_pe_1_1_2_n8), .Z(
        npu_inst_pe_1_1_2_N93) );
  MUX2_X1 npu_inst_pe_1_1_2_U161 ( .A(npu_inst_pe_1_1_2_n31), .B(
        npu_inst_pe_1_1_2_n30), .S(npu_inst_pe_1_1_2_n6), .Z(
        npu_inst_pe_1_1_2_n32) );
  MUX2_X1 npu_inst_pe_1_1_2_U160 ( .A(npu_inst_pe_1_1_2_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_1_2_int_q_reg_v_1__0_), .S(npu_inst_pe_1_1_2_n4), .Z(
        npu_inst_pe_1_1_2_n31) );
  MUX2_X1 npu_inst_pe_1_1_2_U159 ( .A(npu_inst_pe_1_1_2_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_1_2_int_q_reg_v_3__0_), .S(npu_inst_pe_1_1_2_n4), .Z(
        npu_inst_pe_1_1_2_n30) );
  MUX2_X1 npu_inst_pe_1_1_2_U158 ( .A(npu_inst_pe_1_1_2_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_1_2_int_q_reg_v_5__0_), .S(npu_inst_pe_1_1_2_n4), .Z(
        npu_inst_pe_1_1_2_n29) );
  MUX2_X1 npu_inst_pe_1_1_2_U157 ( .A(npu_inst_pe_1_1_2_n28), .B(
        npu_inst_pe_1_1_2_n23), .S(npu_inst_pe_1_1_2_n8), .Z(
        npu_inst_pe_1_1_2_N94) );
  MUX2_X1 npu_inst_pe_1_1_2_U156 ( .A(npu_inst_pe_1_1_2_n25), .B(
        npu_inst_pe_1_1_2_n24), .S(npu_inst_pe_1_1_2_n6), .Z(
        npu_inst_pe_1_1_2_n28) );
  MUX2_X1 npu_inst_pe_1_1_2_U155 ( .A(npu_inst_pe_1_1_2_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_1_2_int_q_reg_v_1__1_), .S(npu_inst_pe_1_1_2_n4), .Z(
        npu_inst_pe_1_1_2_n25) );
  MUX2_X1 npu_inst_pe_1_1_2_U154 ( .A(npu_inst_pe_1_1_2_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_1_2_int_q_reg_v_3__1_), .S(npu_inst_pe_1_1_2_n4), .Z(
        npu_inst_pe_1_1_2_n24) );
  MUX2_X1 npu_inst_pe_1_1_2_U153 ( .A(npu_inst_pe_1_1_2_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_1_2_int_q_reg_v_5__1_), .S(npu_inst_pe_1_1_2_n4), .Z(
        npu_inst_pe_1_1_2_n23) );
  MUX2_X1 npu_inst_pe_1_1_2_U152 ( .A(npu_inst_pe_1_1_2_n22), .B(
        npu_inst_pe_1_1_2_n19), .S(npu_inst_pe_1_1_2_n8), .Z(
        npu_inst_int_data_x_1__2__1_) );
  MUX2_X1 npu_inst_pe_1_1_2_U151 ( .A(npu_inst_pe_1_1_2_n21), .B(
        npu_inst_pe_1_1_2_n20), .S(npu_inst_pe_1_1_2_n6), .Z(
        npu_inst_pe_1_1_2_n22) );
  MUX2_X1 npu_inst_pe_1_1_2_U150 ( .A(npu_inst_pe_1_1_2_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_1_2_int_q_reg_h_1__1_), .S(npu_inst_pe_1_1_2_n4), .Z(
        npu_inst_pe_1_1_2_n21) );
  MUX2_X1 npu_inst_pe_1_1_2_U149 ( .A(npu_inst_pe_1_1_2_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_1_2_int_q_reg_h_3__1_), .S(npu_inst_pe_1_1_2_n4), .Z(
        npu_inst_pe_1_1_2_n20) );
  MUX2_X1 npu_inst_pe_1_1_2_U148 ( .A(npu_inst_pe_1_1_2_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_1_2_int_q_reg_h_5__1_), .S(npu_inst_pe_1_1_2_n4), .Z(
        npu_inst_pe_1_1_2_n19) );
  MUX2_X1 npu_inst_pe_1_1_2_U147 ( .A(npu_inst_pe_1_1_2_n18), .B(
        npu_inst_pe_1_1_2_n15), .S(npu_inst_pe_1_1_2_n8), .Z(
        npu_inst_int_data_x_1__2__0_) );
  MUX2_X1 npu_inst_pe_1_1_2_U146 ( .A(npu_inst_pe_1_1_2_n17), .B(
        npu_inst_pe_1_1_2_n16), .S(npu_inst_pe_1_1_2_n6), .Z(
        npu_inst_pe_1_1_2_n18) );
  MUX2_X1 npu_inst_pe_1_1_2_U145 ( .A(npu_inst_pe_1_1_2_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_1_2_int_q_reg_h_1__0_), .S(npu_inst_pe_1_1_2_n4), .Z(
        npu_inst_pe_1_1_2_n17) );
  MUX2_X1 npu_inst_pe_1_1_2_U144 ( .A(npu_inst_pe_1_1_2_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_1_2_int_q_reg_h_3__0_), .S(npu_inst_pe_1_1_2_n4), .Z(
        npu_inst_pe_1_1_2_n16) );
  MUX2_X1 npu_inst_pe_1_1_2_U143 ( .A(npu_inst_pe_1_1_2_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_1_2_int_q_reg_h_5__0_), .S(npu_inst_pe_1_1_2_n4), .Z(
        npu_inst_pe_1_1_2_n15) );
  XOR2_X1 npu_inst_pe_1_1_2_U142 ( .A(npu_inst_pe_1_1_2_int_data_0_), .B(
        npu_inst_pe_1_1_2_int_q_acc_0_), .Z(npu_inst_pe_1_1_2_N73) );
  AND2_X1 npu_inst_pe_1_1_2_U141 ( .A1(npu_inst_pe_1_1_2_int_q_acc_0_), .A2(
        npu_inst_pe_1_1_2_int_data_0_), .ZN(npu_inst_pe_1_1_2_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_1_2_U140 ( .A(npu_inst_pe_1_1_2_int_q_acc_0_), .B(
        npu_inst_pe_1_1_2_n13), .ZN(npu_inst_pe_1_1_2_N65) );
  OR2_X1 npu_inst_pe_1_1_2_U139 ( .A1(npu_inst_pe_1_1_2_n13), .A2(
        npu_inst_pe_1_1_2_int_q_acc_0_), .ZN(npu_inst_pe_1_1_2_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_1_2_U138 ( .A(npu_inst_pe_1_1_2_int_q_acc_2_), .B(
        npu_inst_pe_1_1_2_add_69_carry_2_), .Z(npu_inst_pe_1_1_2_N75) );
  AND2_X1 npu_inst_pe_1_1_2_U137 ( .A1(npu_inst_pe_1_1_2_add_69_carry_2_), 
        .A2(npu_inst_pe_1_1_2_int_q_acc_2_), .ZN(
        npu_inst_pe_1_1_2_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_1_2_U136 ( .A(npu_inst_pe_1_1_2_int_q_acc_3_), .B(
        npu_inst_pe_1_1_2_add_69_carry_3_), .Z(npu_inst_pe_1_1_2_N76) );
  AND2_X1 npu_inst_pe_1_1_2_U135 ( .A1(npu_inst_pe_1_1_2_add_69_carry_3_), 
        .A2(npu_inst_pe_1_1_2_int_q_acc_3_), .ZN(
        npu_inst_pe_1_1_2_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_1_2_U134 ( .A(npu_inst_pe_1_1_2_int_q_acc_4_), .B(
        npu_inst_pe_1_1_2_add_69_carry_4_), .Z(npu_inst_pe_1_1_2_N77) );
  AND2_X1 npu_inst_pe_1_1_2_U133 ( .A1(npu_inst_pe_1_1_2_add_69_carry_4_), 
        .A2(npu_inst_pe_1_1_2_int_q_acc_4_), .ZN(
        npu_inst_pe_1_1_2_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_1_2_U132 ( .A(npu_inst_pe_1_1_2_int_q_acc_5_), .B(
        npu_inst_pe_1_1_2_add_69_carry_5_), .Z(npu_inst_pe_1_1_2_N78) );
  AND2_X1 npu_inst_pe_1_1_2_U131 ( .A1(npu_inst_pe_1_1_2_add_69_carry_5_), 
        .A2(npu_inst_pe_1_1_2_int_q_acc_5_), .ZN(
        npu_inst_pe_1_1_2_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_1_2_U130 ( .A(npu_inst_pe_1_1_2_int_q_acc_6_), .B(
        npu_inst_pe_1_1_2_add_69_carry_6_), .Z(npu_inst_pe_1_1_2_N79) );
  AND2_X1 npu_inst_pe_1_1_2_U129 ( .A1(npu_inst_pe_1_1_2_add_69_carry_6_), 
        .A2(npu_inst_pe_1_1_2_int_q_acc_6_), .ZN(
        npu_inst_pe_1_1_2_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_1_2_U128 ( .A(npu_inst_pe_1_1_2_int_q_acc_7_), .B(
        npu_inst_pe_1_1_2_add_69_carry_7_), .Z(npu_inst_pe_1_1_2_N80) );
  XNOR2_X1 npu_inst_pe_1_1_2_U127 ( .A(npu_inst_pe_1_1_2_sub_67_carry_2_), .B(
        npu_inst_pe_1_1_2_int_q_acc_2_), .ZN(npu_inst_pe_1_1_2_N67) );
  OR2_X1 npu_inst_pe_1_1_2_U126 ( .A1(npu_inst_pe_1_1_2_int_q_acc_2_), .A2(
        npu_inst_pe_1_1_2_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_1_2_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_1_2_U125 ( .A(npu_inst_pe_1_1_2_sub_67_carry_3_), .B(
        npu_inst_pe_1_1_2_int_q_acc_3_), .ZN(npu_inst_pe_1_1_2_N68) );
  OR2_X1 npu_inst_pe_1_1_2_U124 ( .A1(npu_inst_pe_1_1_2_int_q_acc_3_), .A2(
        npu_inst_pe_1_1_2_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_1_2_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_1_2_U123 ( .A(npu_inst_pe_1_1_2_sub_67_carry_4_), .B(
        npu_inst_pe_1_1_2_int_q_acc_4_), .ZN(npu_inst_pe_1_1_2_N69) );
  OR2_X1 npu_inst_pe_1_1_2_U122 ( .A1(npu_inst_pe_1_1_2_int_q_acc_4_), .A2(
        npu_inst_pe_1_1_2_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_1_2_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_1_2_U121 ( .A(npu_inst_pe_1_1_2_sub_67_carry_5_), .B(
        npu_inst_pe_1_1_2_int_q_acc_5_), .ZN(npu_inst_pe_1_1_2_N70) );
  OR2_X1 npu_inst_pe_1_1_2_U120 ( .A1(npu_inst_pe_1_1_2_int_q_acc_5_), .A2(
        npu_inst_pe_1_1_2_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_1_2_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_1_2_U119 ( .A(npu_inst_pe_1_1_2_sub_67_carry_6_), .B(
        npu_inst_pe_1_1_2_int_q_acc_6_), .ZN(npu_inst_pe_1_1_2_N71) );
  OR2_X1 npu_inst_pe_1_1_2_U118 ( .A1(npu_inst_pe_1_1_2_int_q_acc_6_), .A2(
        npu_inst_pe_1_1_2_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_1_2_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_1_2_U117 ( .A(npu_inst_pe_1_1_2_int_q_acc_7_), .B(
        npu_inst_pe_1_1_2_sub_67_carry_7_), .ZN(npu_inst_pe_1_1_2_N72) );
  INV_X1 npu_inst_pe_1_1_2_U116 ( .A(npu_inst_n79), .ZN(npu_inst_pe_1_1_2_n7)
         );
  INV_X1 npu_inst_pe_1_1_2_U115 ( .A(npu_inst_pe_1_1_2_n7), .ZN(
        npu_inst_pe_1_1_2_n6) );
  INV_X1 npu_inst_pe_1_1_2_U114 ( .A(npu_inst_n59), .ZN(npu_inst_pe_1_1_2_n3)
         );
  AOI22_X1 npu_inst_pe_1_1_2_U113 ( .A1(npu_inst_int_data_y_2__2__0_), .A2(
        npu_inst_pe_1_1_2_n58), .B1(npu_inst_pe_1_1_2_n119), .B2(
        npu_inst_pe_1_1_2_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_1_2_n57) );
  INV_X1 npu_inst_pe_1_1_2_U112 ( .A(npu_inst_pe_1_1_2_n57), .ZN(
        npu_inst_pe_1_1_2_n108) );
  AOI22_X1 npu_inst_pe_1_1_2_U111 ( .A1(npu_inst_int_data_y_2__2__0_), .A2(
        npu_inst_pe_1_1_2_n54), .B1(npu_inst_pe_1_1_2_n118), .B2(
        npu_inst_pe_1_1_2_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_1_2_n53) );
  INV_X1 npu_inst_pe_1_1_2_U110 ( .A(npu_inst_pe_1_1_2_n53), .ZN(
        npu_inst_pe_1_1_2_n109) );
  AOI22_X1 npu_inst_pe_1_1_2_U107 ( .A1(npu_inst_int_data_y_2__2__0_), .A2(
        npu_inst_pe_1_1_2_n50), .B1(npu_inst_pe_1_1_2_n117), .B2(
        npu_inst_pe_1_1_2_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_1_2_n49) );
  INV_X1 npu_inst_pe_1_1_2_U106 ( .A(npu_inst_pe_1_1_2_n49), .ZN(
        npu_inst_pe_1_1_2_n110) );
  AOI22_X1 npu_inst_pe_1_1_2_U105 ( .A1(npu_inst_int_data_y_2__2__0_), .A2(
        npu_inst_pe_1_1_2_n46), .B1(npu_inst_pe_1_1_2_n116), .B2(
        npu_inst_pe_1_1_2_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_1_2_n45) );
  INV_X1 npu_inst_pe_1_1_2_U104 ( .A(npu_inst_pe_1_1_2_n45), .ZN(
        npu_inst_pe_1_1_2_n111) );
  AOI22_X1 npu_inst_pe_1_1_2_U103 ( .A1(npu_inst_int_data_y_2__2__0_), .A2(
        npu_inst_pe_1_1_2_n42), .B1(npu_inst_pe_1_1_2_n115), .B2(
        npu_inst_pe_1_1_2_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_1_2_n41) );
  INV_X1 npu_inst_pe_1_1_2_U102 ( .A(npu_inst_pe_1_1_2_n41), .ZN(
        npu_inst_pe_1_1_2_n112) );
  AOI22_X1 npu_inst_pe_1_1_2_U101 ( .A1(npu_inst_int_data_y_2__2__1_), .A2(
        npu_inst_pe_1_1_2_n58), .B1(npu_inst_pe_1_1_2_n119), .B2(
        npu_inst_pe_1_1_2_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_1_2_n59) );
  INV_X1 npu_inst_pe_1_1_2_U100 ( .A(npu_inst_pe_1_1_2_n59), .ZN(
        npu_inst_pe_1_1_2_n102) );
  AOI22_X1 npu_inst_pe_1_1_2_U99 ( .A1(npu_inst_int_data_y_2__2__1_), .A2(
        npu_inst_pe_1_1_2_n54), .B1(npu_inst_pe_1_1_2_n118), .B2(
        npu_inst_pe_1_1_2_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_1_2_n55) );
  INV_X1 npu_inst_pe_1_1_2_U98 ( .A(npu_inst_pe_1_1_2_n55), .ZN(
        npu_inst_pe_1_1_2_n103) );
  AOI22_X1 npu_inst_pe_1_1_2_U97 ( .A1(npu_inst_int_data_y_2__2__1_), .A2(
        npu_inst_pe_1_1_2_n50), .B1(npu_inst_pe_1_1_2_n117), .B2(
        npu_inst_pe_1_1_2_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_1_2_n51) );
  INV_X1 npu_inst_pe_1_1_2_U96 ( .A(npu_inst_pe_1_1_2_n51), .ZN(
        npu_inst_pe_1_1_2_n104) );
  AOI22_X1 npu_inst_pe_1_1_2_U95 ( .A1(npu_inst_int_data_y_2__2__1_), .A2(
        npu_inst_pe_1_1_2_n46), .B1(npu_inst_pe_1_1_2_n116), .B2(
        npu_inst_pe_1_1_2_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_1_2_n47) );
  INV_X1 npu_inst_pe_1_1_2_U94 ( .A(npu_inst_pe_1_1_2_n47), .ZN(
        npu_inst_pe_1_1_2_n105) );
  AOI22_X1 npu_inst_pe_1_1_2_U93 ( .A1(npu_inst_int_data_y_2__2__1_), .A2(
        npu_inst_pe_1_1_2_n42), .B1(npu_inst_pe_1_1_2_n115), .B2(
        npu_inst_pe_1_1_2_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_1_2_n43) );
  INV_X1 npu_inst_pe_1_1_2_U92 ( .A(npu_inst_pe_1_1_2_n43), .ZN(
        npu_inst_pe_1_1_2_n106) );
  AOI22_X1 npu_inst_pe_1_1_2_U91 ( .A1(npu_inst_pe_1_1_2_n38), .A2(
        npu_inst_int_data_y_2__2__1_), .B1(npu_inst_pe_1_1_2_n114), .B2(
        npu_inst_pe_1_1_2_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_1_2_n39) );
  INV_X1 npu_inst_pe_1_1_2_U90 ( .A(npu_inst_pe_1_1_2_n39), .ZN(
        npu_inst_pe_1_1_2_n107) );
  AOI22_X1 npu_inst_pe_1_1_2_U89 ( .A1(npu_inst_pe_1_1_2_n38), .A2(
        npu_inst_int_data_y_2__2__0_), .B1(npu_inst_pe_1_1_2_n114), .B2(
        npu_inst_pe_1_1_2_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_1_2_n37) );
  INV_X1 npu_inst_pe_1_1_2_U88 ( .A(npu_inst_pe_1_1_2_n37), .ZN(
        npu_inst_pe_1_1_2_n113) );
  NAND2_X1 npu_inst_pe_1_1_2_U87 ( .A1(npu_inst_pe_1_1_2_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_1_2_n60), .ZN(npu_inst_pe_1_1_2_n74) );
  OAI21_X1 npu_inst_pe_1_1_2_U86 ( .B1(npu_inst_pe_1_1_2_n63), .B2(
        npu_inst_pe_1_1_2_n60), .A(npu_inst_pe_1_1_2_n74), .ZN(
        npu_inst_pe_1_1_2_n97) );
  NAND2_X1 npu_inst_pe_1_1_2_U85 ( .A1(npu_inst_pe_1_1_2_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_1_2_n60), .ZN(npu_inst_pe_1_1_2_n73) );
  OAI21_X1 npu_inst_pe_1_1_2_U84 ( .B1(npu_inst_pe_1_1_2_n61), .B2(
        npu_inst_pe_1_1_2_n60), .A(npu_inst_pe_1_1_2_n73), .ZN(
        npu_inst_pe_1_1_2_n96) );
  NAND2_X1 npu_inst_pe_1_1_2_U83 ( .A1(npu_inst_pe_1_1_2_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_1_2_n56), .ZN(npu_inst_pe_1_1_2_n72) );
  OAI21_X1 npu_inst_pe_1_1_2_U82 ( .B1(npu_inst_pe_1_1_2_n63), .B2(
        npu_inst_pe_1_1_2_n56), .A(npu_inst_pe_1_1_2_n72), .ZN(
        npu_inst_pe_1_1_2_n95) );
  NAND2_X1 npu_inst_pe_1_1_2_U81 ( .A1(npu_inst_pe_1_1_2_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_1_2_n56), .ZN(npu_inst_pe_1_1_2_n71) );
  OAI21_X1 npu_inst_pe_1_1_2_U80 ( .B1(npu_inst_pe_1_1_2_n61), .B2(
        npu_inst_pe_1_1_2_n56), .A(npu_inst_pe_1_1_2_n71), .ZN(
        npu_inst_pe_1_1_2_n94) );
  NAND2_X1 npu_inst_pe_1_1_2_U79 ( .A1(npu_inst_pe_1_1_2_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_1_2_n52), .ZN(npu_inst_pe_1_1_2_n70) );
  OAI21_X1 npu_inst_pe_1_1_2_U78 ( .B1(npu_inst_pe_1_1_2_n63), .B2(
        npu_inst_pe_1_1_2_n52), .A(npu_inst_pe_1_1_2_n70), .ZN(
        npu_inst_pe_1_1_2_n93) );
  NAND2_X1 npu_inst_pe_1_1_2_U77 ( .A1(npu_inst_pe_1_1_2_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_1_2_n52), .ZN(npu_inst_pe_1_1_2_n69) );
  OAI21_X1 npu_inst_pe_1_1_2_U76 ( .B1(npu_inst_pe_1_1_2_n61), .B2(
        npu_inst_pe_1_1_2_n52), .A(npu_inst_pe_1_1_2_n69), .ZN(
        npu_inst_pe_1_1_2_n92) );
  NAND2_X1 npu_inst_pe_1_1_2_U75 ( .A1(npu_inst_pe_1_1_2_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_1_2_n48), .ZN(npu_inst_pe_1_1_2_n68) );
  OAI21_X1 npu_inst_pe_1_1_2_U74 ( .B1(npu_inst_pe_1_1_2_n63), .B2(
        npu_inst_pe_1_1_2_n48), .A(npu_inst_pe_1_1_2_n68), .ZN(
        npu_inst_pe_1_1_2_n91) );
  NAND2_X1 npu_inst_pe_1_1_2_U73 ( .A1(npu_inst_pe_1_1_2_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_1_2_n48), .ZN(npu_inst_pe_1_1_2_n67) );
  OAI21_X1 npu_inst_pe_1_1_2_U72 ( .B1(npu_inst_pe_1_1_2_n61), .B2(
        npu_inst_pe_1_1_2_n48), .A(npu_inst_pe_1_1_2_n67), .ZN(
        npu_inst_pe_1_1_2_n90) );
  NAND2_X1 npu_inst_pe_1_1_2_U71 ( .A1(npu_inst_pe_1_1_2_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_1_2_n44), .ZN(npu_inst_pe_1_1_2_n66) );
  OAI21_X1 npu_inst_pe_1_1_2_U70 ( .B1(npu_inst_pe_1_1_2_n63), .B2(
        npu_inst_pe_1_1_2_n44), .A(npu_inst_pe_1_1_2_n66), .ZN(
        npu_inst_pe_1_1_2_n89) );
  NAND2_X1 npu_inst_pe_1_1_2_U69 ( .A1(npu_inst_pe_1_1_2_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_1_2_n44), .ZN(npu_inst_pe_1_1_2_n65) );
  OAI21_X1 npu_inst_pe_1_1_2_U68 ( .B1(npu_inst_pe_1_1_2_n61), .B2(
        npu_inst_pe_1_1_2_n44), .A(npu_inst_pe_1_1_2_n65), .ZN(
        npu_inst_pe_1_1_2_n88) );
  NAND2_X1 npu_inst_pe_1_1_2_U67 ( .A1(npu_inst_pe_1_1_2_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_1_2_n40), .ZN(npu_inst_pe_1_1_2_n64) );
  OAI21_X1 npu_inst_pe_1_1_2_U66 ( .B1(npu_inst_pe_1_1_2_n63), .B2(
        npu_inst_pe_1_1_2_n40), .A(npu_inst_pe_1_1_2_n64), .ZN(
        npu_inst_pe_1_1_2_n87) );
  NAND2_X1 npu_inst_pe_1_1_2_U65 ( .A1(npu_inst_pe_1_1_2_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_1_2_n40), .ZN(npu_inst_pe_1_1_2_n62) );
  OAI21_X1 npu_inst_pe_1_1_2_U64 ( .B1(npu_inst_pe_1_1_2_n61), .B2(
        npu_inst_pe_1_1_2_n40), .A(npu_inst_pe_1_1_2_n62), .ZN(
        npu_inst_pe_1_1_2_n86) );
  AND2_X1 npu_inst_pe_1_1_2_U63 ( .A1(npu_inst_pe_1_1_2_N93), .A2(npu_inst_n59), .ZN(npu_inst_int_data_y_1__2__0_) );
  AND2_X1 npu_inst_pe_1_1_2_U62 ( .A1(npu_inst_n59), .A2(npu_inst_pe_1_1_2_N94), .ZN(npu_inst_int_data_y_1__2__1_) );
  NOR3_X1 npu_inst_pe_1_1_2_U61 ( .A1(npu_inst_pe_1_1_2_n26), .A2(npu_inst_n59), .A3(npu_inst_int_ckg[53]), .ZN(npu_inst_pe_1_1_2_n85) );
  OR2_X1 npu_inst_pe_1_1_2_U60 ( .A1(npu_inst_pe_1_1_2_n85), .A2(
        npu_inst_pe_1_1_2_n2), .ZN(npu_inst_pe_1_1_2_N84) );
  AND2_X1 npu_inst_pe_1_1_2_U59 ( .A1(npu_inst_pe_1_1_2_int_q_acc_0_), .A2(
        npu_inst_pe_1_1_2_n1), .ZN(npu_inst_int_data_res_1__2__0_) );
  AND2_X1 npu_inst_pe_1_1_2_U58 ( .A1(npu_inst_pe_1_1_2_n2), .A2(
        npu_inst_pe_1_1_2_int_q_acc_7_), .ZN(npu_inst_int_data_res_1__2__7_)
         );
  AND2_X1 npu_inst_pe_1_1_2_U57 ( .A1(npu_inst_pe_1_1_2_int_q_acc_1_), .A2(
        npu_inst_pe_1_1_2_n1), .ZN(npu_inst_int_data_res_1__2__1_) );
  AND2_X1 npu_inst_pe_1_1_2_U56 ( .A1(npu_inst_pe_1_1_2_int_q_acc_2_), .A2(
        npu_inst_pe_1_1_2_n1), .ZN(npu_inst_int_data_res_1__2__2_) );
  AND2_X1 npu_inst_pe_1_1_2_U55 ( .A1(npu_inst_pe_1_1_2_int_q_acc_3_), .A2(
        npu_inst_pe_1_1_2_n2), .ZN(npu_inst_int_data_res_1__2__3_) );
  AND2_X1 npu_inst_pe_1_1_2_U54 ( .A1(npu_inst_pe_1_1_2_int_q_acc_4_), .A2(
        npu_inst_pe_1_1_2_n2), .ZN(npu_inst_int_data_res_1__2__4_) );
  AND2_X1 npu_inst_pe_1_1_2_U53 ( .A1(npu_inst_pe_1_1_2_int_q_acc_5_), .A2(
        npu_inst_pe_1_1_2_n2), .ZN(npu_inst_int_data_res_1__2__5_) );
  AND2_X1 npu_inst_pe_1_1_2_U52 ( .A1(npu_inst_pe_1_1_2_int_q_acc_6_), .A2(
        npu_inst_pe_1_1_2_n2), .ZN(npu_inst_int_data_res_1__2__6_) );
  AOI222_X1 npu_inst_pe_1_1_2_U51 ( .A1(npu_inst_int_data_res_2__2__0_), .A2(
        npu_inst_pe_1_1_2_n1), .B1(npu_inst_pe_1_1_2_N73), .B2(
        npu_inst_pe_1_1_2_n76), .C1(npu_inst_pe_1_1_2_N65), .C2(
        npu_inst_pe_1_1_2_n77), .ZN(npu_inst_pe_1_1_2_n84) );
  INV_X1 npu_inst_pe_1_1_2_U50 ( .A(npu_inst_pe_1_1_2_n84), .ZN(
        npu_inst_pe_1_1_2_n101) );
  AOI222_X1 npu_inst_pe_1_1_2_U49 ( .A1(npu_inst_int_data_res_2__2__7_), .A2(
        npu_inst_pe_1_1_2_n1), .B1(npu_inst_pe_1_1_2_N80), .B2(
        npu_inst_pe_1_1_2_n76), .C1(npu_inst_pe_1_1_2_N72), .C2(
        npu_inst_pe_1_1_2_n77), .ZN(npu_inst_pe_1_1_2_n75) );
  INV_X1 npu_inst_pe_1_1_2_U48 ( .A(npu_inst_pe_1_1_2_n75), .ZN(
        npu_inst_pe_1_1_2_n33) );
  AOI222_X1 npu_inst_pe_1_1_2_U47 ( .A1(npu_inst_int_data_res_2__2__1_), .A2(
        npu_inst_pe_1_1_2_n1), .B1(npu_inst_pe_1_1_2_N74), .B2(
        npu_inst_pe_1_1_2_n76), .C1(npu_inst_pe_1_1_2_N66), .C2(
        npu_inst_pe_1_1_2_n77), .ZN(npu_inst_pe_1_1_2_n83) );
  INV_X1 npu_inst_pe_1_1_2_U46 ( .A(npu_inst_pe_1_1_2_n83), .ZN(
        npu_inst_pe_1_1_2_n100) );
  AOI222_X1 npu_inst_pe_1_1_2_U45 ( .A1(npu_inst_int_data_res_2__2__2_), .A2(
        npu_inst_pe_1_1_2_n1), .B1(npu_inst_pe_1_1_2_N75), .B2(
        npu_inst_pe_1_1_2_n76), .C1(npu_inst_pe_1_1_2_N67), .C2(
        npu_inst_pe_1_1_2_n77), .ZN(npu_inst_pe_1_1_2_n82) );
  INV_X1 npu_inst_pe_1_1_2_U44 ( .A(npu_inst_pe_1_1_2_n82), .ZN(
        npu_inst_pe_1_1_2_n99) );
  AOI222_X1 npu_inst_pe_1_1_2_U43 ( .A1(npu_inst_int_data_res_2__2__3_), .A2(
        npu_inst_pe_1_1_2_n1), .B1(npu_inst_pe_1_1_2_N76), .B2(
        npu_inst_pe_1_1_2_n76), .C1(npu_inst_pe_1_1_2_N68), .C2(
        npu_inst_pe_1_1_2_n77), .ZN(npu_inst_pe_1_1_2_n81) );
  INV_X1 npu_inst_pe_1_1_2_U42 ( .A(npu_inst_pe_1_1_2_n81), .ZN(
        npu_inst_pe_1_1_2_n98) );
  AOI222_X1 npu_inst_pe_1_1_2_U41 ( .A1(npu_inst_int_data_res_2__2__4_), .A2(
        npu_inst_pe_1_1_2_n1), .B1(npu_inst_pe_1_1_2_N77), .B2(
        npu_inst_pe_1_1_2_n76), .C1(npu_inst_pe_1_1_2_N69), .C2(
        npu_inst_pe_1_1_2_n77), .ZN(npu_inst_pe_1_1_2_n80) );
  INV_X1 npu_inst_pe_1_1_2_U40 ( .A(npu_inst_pe_1_1_2_n80), .ZN(
        npu_inst_pe_1_1_2_n36) );
  AOI222_X1 npu_inst_pe_1_1_2_U39 ( .A1(npu_inst_int_data_res_2__2__5_), .A2(
        npu_inst_pe_1_1_2_n1), .B1(npu_inst_pe_1_1_2_N78), .B2(
        npu_inst_pe_1_1_2_n76), .C1(npu_inst_pe_1_1_2_N70), .C2(
        npu_inst_pe_1_1_2_n77), .ZN(npu_inst_pe_1_1_2_n79) );
  INV_X1 npu_inst_pe_1_1_2_U38 ( .A(npu_inst_pe_1_1_2_n79), .ZN(
        npu_inst_pe_1_1_2_n35) );
  AOI222_X1 npu_inst_pe_1_1_2_U37 ( .A1(npu_inst_int_data_res_2__2__6_), .A2(
        npu_inst_pe_1_1_2_n1), .B1(npu_inst_pe_1_1_2_N79), .B2(
        npu_inst_pe_1_1_2_n76), .C1(npu_inst_pe_1_1_2_N71), .C2(
        npu_inst_pe_1_1_2_n77), .ZN(npu_inst_pe_1_1_2_n78) );
  INV_X1 npu_inst_pe_1_1_2_U36 ( .A(npu_inst_pe_1_1_2_n78), .ZN(
        npu_inst_pe_1_1_2_n34) );
  INV_X1 npu_inst_pe_1_1_2_U35 ( .A(npu_inst_pe_1_1_2_int_data_1_), .ZN(
        npu_inst_pe_1_1_2_n14) );
  AND2_X1 npu_inst_pe_1_1_2_U34 ( .A1(npu_inst_int_data_x_1__2__1_), .A2(
        npu_inst_pe_1_1_2_int_q_weight_1_), .ZN(npu_inst_pe_1_1_2_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_1_2_U33 ( .A1(npu_inst_int_data_x_1__2__0_), .A2(
        npu_inst_pe_1_1_2_int_q_weight_1_), .ZN(npu_inst_pe_1_1_2_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_1_2_U32 ( .A1(npu_inst_n59), .A2(
        npu_inst_int_data_y_2__2__1_), .B1(npu_inst_pe_1_1_2_n3), .B2(
        npu_inst_int_data_x_1__3__1_), .ZN(npu_inst_pe_1_1_2_n63) );
  AOI22_X1 npu_inst_pe_1_1_2_U31 ( .A1(npu_inst_n59), .A2(
        npu_inst_int_data_y_2__2__0_), .B1(npu_inst_pe_1_1_2_n3), .B2(
        npu_inst_int_data_x_1__3__0_), .ZN(npu_inst_pe_1_1_2_n61) );
  INV_X1 npu_inst_pe_1_1_2_U30 ( .A(npu_inst_pe_1_1_2_int_data_0_), .ZN(
        npu_inst_pe_1_1_2_n13) );
  INV_X1 npu_inst_pe_1_1_2_U29 ( .A(npu_inst_n71), .ZN(npu_inst_pe_1_1_2_n5)
         );
  OR3_X1 npu_inst_pe_1_1_2_U28 ( .A1(npu_inst_pe_1_1_2_n6), .A2(
        npu_inst_pe_1_1_2_n8), .A3(npu_inst_pe_1_1_2_n5), .ZN(
        npu_inst_pe_1_1_2_n56) );
  OR3_X1 npu_inst_pe_1_1_2_U27 ( .A1(npu_inst_pe_1_1_2_n5), .A2(
        npu_inst_pe_1_1_2_n8), .A3(npu_inst_pe_1_1_2_n7), .ZN(
        npu_inst_pe_1_1_2_n48) );
  INV_X1 npu_inst_pe_1_1_2_U26 ( .A(npu_inst_pe_1_1_2_n5), .ZN(
        npu_inst_pe_1_1_2_n4) );
  OR3_X1 npu_inst_pe_1_1_2_U25 ( .A1(npu_inst_pe_1_1_2_n4), .A2(
        npu_inst_pe_1_1_2_n8), .A3(npu_inst_pe_1_1_2_n7), .ZN(
        npu_inst_pe_1_1_2_n52) );
  OR3_X1 npu_inst_pe_1_1_2_U24 ( .A1(npu_inst_pe_1_1_2_n6), .A2(
        npu_inst_pe_1_1_2_n8), .A3(npu_inst_pe_1_1_2_n4), .ZN(
        npu_inst_pe_1_1_2_n60) );
  NOR2_X1 npu_inst_pe_1_1_2_U23 ( .A1(npu_inst_pe_1_1_2_n60), .A2(
        npu_inst_pe_1_1_2_n3), .ZN(npu_inst_pe_1_1_2_n58) );
  NOR2_X1 npu_inst_pe_1_1_2_U22 ( .A1(npu_inst_pe_1_1_2_n56), .A2(
        npu_inst_pe_1_1_2_n3), .ZN(npu_inst_pe_1_1_2_n54) );
  NOR2_X1 npu_inst_pe_1_1_2_U21 ( .A1(npu_inst_pe_1_1_2_n52), .A2(
        npu_inst_pe_1_1_2_n3), .ZN(npu_inst_pe_1_1_2_n50) );
  NOR2_X1 npu_inst_pe_1_1_2_U20 ( .A1(npu_inst_pe_1_1_2_n48), .A2(
        npu_inst_pe_1_1_2_n3), .ZN(npu_inst_pe_1_1_2_n46) );
  NOR2_X1 npu_inst_pe_1_1_2_U19 ( .A1(npu_inst_pe_1_1_2_n40), .A2(
        npu_inst_pe_1_1_2_n3), .ZN(npu_inst_pe_1_1_2_n38) );
  NOR2_X1 npu_inst_pe_1_1_2_U18 ( .A1(npu_inst_pe_1_1_2_n44), .A2(
        npu_inst_pe_1_1_2_n3), .ZN(npu_inst_pe_1_1_2_n42) );
  BUF_X1 npu_inst_pe_1_1_2_U17 ( .A(npu_inst_n105), .Z(npu_inst_pe_1_1_2_n8)
         );
  INV_X1 npu_inst_pe_1_1_2_U16 ( .A(npu_inst_n126), .ZN(npu_inst_pe_1_1_2_n12)
         );
  INV_X1 npu_inst_pe_1_1_2_U15 ( .A(npu_inst_pe_1_1_2_n38), .ZN(
        npu_inst_pe_1_1_2_n114) );
  INV_X1 npu_inst_pe_1_1_2_U14 ( .A(npu_inst_pe_1_1_2_n58), .ZN(
        npu_inst_pe_1_1_2_n119) );
  INV_X1 npu_inst_pe_1_1_2_U13 ( .A(npu_inst_pe_1_1_2_n54), .ZN(
        npu_inst_pe_1_1_2_n118) );
  INV_X1 npu_inst_pe_1_1_2_U12 ( .A(npu_inst_pe_1_1_2_n50), .ZN(
        npu_inst_pe_1_1_2_n117) );
  INV_X1 npu_inst_pe_1_1_2_U11 ( .A(npu_inst_pe_1_1_2_n46), .ZN(
        npu_inst_pe_1_1_2_n116) );
  INV_X1 npu_inst_pe_1_1_2_U10 ( .A(npu_inst_pe_1_1_2_n42), .ZN(
        npu_inst_pe_1_1_2_n115) );
  BUF_X1 npu_inst_pe_1_1_2_U9 ( .A(npu_inst_n33), .Z(npu_inst_pe_1_1_2_n2) );
  BUF_X1 npu_inst_pe_1_1_2_U8 ( .A(npu_inst_n33), .Z(npu_inst_pe_1_1_2_n1) );
  BUF_X1 npu_inst_pe_1_1_2_U7 ( .A(npu_inst_pe_1_1_2_n12), .Z(
        npu_inst_pe_1_1_2_n11) );
  BUF_X1 npu_inst_pe_1_1_2_U6 ( .A(npu_inst_pe_1_1_2_n12), .Z(
        npu_inst_pe_1_1_2_n10) );
  BUF_X1 npu_inst_pe_1_1_2_U5 ( .A(npu_inst_pe_1_1_2_n12), .Z(
        npu_inst_pe_1_1_2_n9) );
  NOR2_X1 npu_inst_pe_1_1_2_U4 ( .A1(npu_inst_pe_1_1_2_int_q_weight_0_), .A2(
        npu_inst_pe_1_1_2_n1), .ZN(npu_inst_pe_1_1_2_n76) );
  NOR2_X1 npu_inst_pe_1_1_2_U3 ( .A1(npu_inst_pe_1_1_2_n27), .A2(
        npu_inst_pe_1_1_2_n1), .ZN(npu_inst_pe_1_1_2_n77) );
  FA_X1 npu_inst_pe_1_1_2_sub_67_U2_1 ( .A(npu_inst_pe_1_1_2_int_q_acc_1_), 
        .B(npu_inst_pe_1_1_2_n14), .CI(npu_inst_pe_1_1_2_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_1_2_sub_67_carry_2_), .S(npu_inst_pe_1_1_2_N66) );
  FA_X1 npu_inst_pe_1_1_2_add_69_U1_1 ( .A(npu_inst_pe_1_1_2_int_q_acc_1_), 
        .B(npu_inst_pe_1_1_2_int_data_1_), .CI(
        npu_inst_pe_1_1_2_add_69_carry_1_), .CO(
        npu_inst_pe_1_1_2_add_69_carry_2_), .S(npu_inst_pe_1_1_2_N74) );
  NAND3_X1 npu_inst_pe_1_1_2_U109 ( .A1(npu_inst_pe_1_1_2_n5), .A2(
        npu_inst_pe_1_1_2_n7), .A3(npu_inst_pe_1_1_2_n8), .ZN(
        npu_inst_pe_1_1_2_n44) );
  NAND3_X1 npu_inst_pe_1_1_2_U108 ( .A1(npu_inst_pe_1_1_2_n4), .A2(
        npu_inst_pe_1_1_2_n7), .A3(npu_inst_pe_1_1_2_n8), .ZN(
        npu_inst_pe_1_1_2_n40) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_1_2_n34), .CK(
        npu_inst_pe_1_1_2_net4332), .RN(npu_inst_pe_1_1_2_n9), .Q(
        npu_inst_pe_1_1_2_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_1_2_n35), .CK(
        npu_inst_pe_1_1_2_net4332), .RN(npu_inst_pe_1_1_2_n9), .Q(
        npu_inst_pe_1_1_2_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_1_2_n36), .CK(
        npu_inst_pe_1_1_2_net4332), .RN(npu_inst_pe_1_1_2_n9), .Q(
        npu_inst_pe_1_1_2_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_1_2_n98), .CK(
        npu_inst_pe_1_1_2_net4332), .RN(npu_inst_pe_1_1_2_n9), .Q(
        npu_inst_pe_1_1_2_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_1_2_n99), .CK(
        npu_inst_pe_1_1_2_net4332), .RN(npu_inst_pe_1_1_2_n9), .Q(
        npu_inst_pe_1_1_2_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_1_2_n100), 
        .CK(npu_inst_pe_1_1_2_net4332), .RN(npu_inst_pe_1_1_2_n9), .Q(
        npu_inst_pe_1_1_2_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_1_2_n33), .CK(
        npu_inst_pe_1_1_2_net4332), .RN(npu_inst_pe_1_1_2_n9), .Q(
        npu_inst_pe_1_1_2_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_1_2_n101), 
        .CK(npu_inst_pe_1_1_2_net4332), .RN(npu_inst_pe_1_1_2_n9), .Q(
        npu_inst_pe_1_1_2_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_weight_reg_0_ ( .D(npu_inst_n112), .CK(
        npu_inst_pe_1_1_2_net4338), .RN(npu_inst_pe_1_1_2_n9), .Q(
        npu_inst_pe_1_1_2_int_q_weight_0_), .QN(npu_inst_pe_1_1_2_n27) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_weight_reg_1_ ( .D(npu_inst_n118), .CK(
        npu_inst_pe_1_1_2_net4338), .RN(npu_inst_pe_1_1_2_n9), .Q(
        npu_inst_pe_1_1_2_int_q_weight_1_), .QN(npu_inst_pe_1_1_2_n26) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_1_2_n113), 
        .CK(npu_inst_pe_1_1_2_net4338), .RN(npu_inst_pe_1_1_2_n9), .Q(
        npu_inst_pe_1_1_2_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_1_2_n107), 
        .CK(npu_inst_pe_1_1_2_net4338), .RN(npu_inst_pe_1_1_2_n9), .Q(
        npu_inst_pe_1_1_2_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_1_2_n112), 
        .CK(npu_inst_pe_1_1_2_net4338), .RN(npu_inst_pe_1_1_2_n10), .Q(
        npu_inst_pe_1_1_2_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_1_2_n106), 
        .CK(npu_inst_pe_1_1_2_net4338), .RN(npu_inst_pe_1_1_2_n10), .Q(
        npu_inst_pe_1_1_2_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_1_2_n111), 
        .CK(npu_inst_pe_1_1_2_net4338), .RN(npu_inst_pe_1_1_2_n10), .Q(
        npu_inst_pe_1_1_2_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_1_2_n105), 
        .CK(npu_inst_pe_1_1_2_net4338), .RN(npu_inst_pe_1_1_2_n10), .Q(
        npu_inst_pe_1_1_2_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_1_2_n110), 
        .CK(npu_inst_pe_1_1_2_net4338), .RN(npu_inst_pe_1_1_2_n10), .Q(
        npu_inst_pe_1_1_2_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_1_2_n104), 
        .CK(npu_inst_pe_1_1_2_net4338), .RN(npu_inst_pe_1_1_2_n10), .Q(
        npu_inst_pe_1_1_2_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_1_2_n109), 
        .CK(npu_inst_pe_1_1_2_net4338), .RN(npu_inst_pe_1_1_2_n10), .Q(
        npu_inst_pe_1_1_2_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_1_2_n103), 
        .CK(npu_inst_pe_1_1_2_net4338), .RN(npu_inst_pe_1_1_2_n10), .Q(
        npu_inst_pe_1_1_2_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_1_2_n108), 
        .CK(npu_inst_pe_1_1_2_net4338), .RN(npu_inst_pe_1_1_2_n10), .Q(
        npu_inst_pe_1_1_2_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_1_2_n102), 
        .CK(npu_inst_pe_1_1_2_net4338), .RN(npu_inst_pe_1_1_2_n10), .Q(
        npu_inst_pe_1_1_2_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_1_2_n86), 
        .CK(npu_inst_pe_1_1_2_net4338), .RN(npu_inst_pe_1_1_2_n10), .Q(
        npu_inst_pe_1_1_2_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_1_2_n87), 
        .CK(npu_inst_pe_1_1_2_net4338), .RN(npu_inst_pe_1_1_2_n10), .Q(
        npu_inst_pe_1_1_2_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_1_2_n88), 
        .CK(npu_inst_pe_1_1_2_net4338), .RN(npu_inst_pe_1_1_2_n11), .Q(
        npu_inst_pe_1_1_2_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_1_2_n89), 
        .CK(npu_inst_pe_1_1_2_net4338), .RN(npu_inst_pe_1_1_2_n11), .Q(
        npu_inst_pe_1_1_2_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_1_2_n90), 
        .CK(npu_inst_pe_1_1_2_net4338), .RN(npu_inst_pe_1_1_2_n11), .Q(
        npu_inst_pe_1_1_2_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_1_2_n91), 
        .CK(npu_inst_pe_1_1_2_net4338), .RN(npu_inst_pe_1_1_2_n11), .Q(
        npu_inst_pe_1_1_2_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_1_2_n92), 
        .CK(npu_inst_pe_1_1_2_net4338), .RN(npu_inst_pe_1_1_2_n11), .Q(
        npu_inst_pe_1_1_2_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_1_2_n93), 
        .CK(npu_inst_pe_1_1_2_net4338), .RN(npu_inst_pe_1_1_2_n11), .Q(
        npu_inst_pe_1_1_2_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_1_2_n94), 
        .CK(npu_inst_pe_1_1_2_net4338), .RN(npu_inst_pe_1_1_2_n11), .Q(
        npu_inst_pe_1_1_2_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_1_2_n95), 
        .CK(npu_inst_pe_1_1_2_net4338), .RN(npu_inst_pe_1_1_2_n11), .Q(
        npu_inst_pe_1_1_2_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_1_2_n96), 
        .CK(npu_inst_pe_1_1_2_net4338), .RN(npu_inst_pe_1_1_2_n11), .Q(
        npu_inst_pe_1_1_2_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_1_2_n97), 
        .CK(npu_inst_pe_1_1_2_net4338), .RN(npu_inst_pe_1_1_2_n11), .Q(
        npu_inst_pe_1_1_2_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_1_2_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_1_2_N84), .SE(1'b0), .GCK(npu_inst_pe_1_1_2_net4332) );
  CLKGATETST_X1 npu_inst_pe_1_1_2_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n65), .SE(1'b0), .GCK(npu_inst_pe_1_1_2_net4338) );
  MUX2_X1 npu_inst_pe_1_1_3_U162 ( .A(npu_inst_pe_1_1_3_n32), .B(
        npu_inst_pe_1_1_3_n29), .S(npu_inst_pe_1_1_3_n8), .Z(
        npu_inst_pe_1_1_3_N93) );
  MUX2_X1 npu_inst_pe_1_1_3_U161 ( .A(npu_inst_pe_1_1_3_n31), .B(
        npu_inst_pe_1_1_3_n30), .S(npu_inst_pe_1_1_3_n6), .Z(
        npu_inst_pe_1_1_3_n32) );
  MUX2_X1 npu_inst_pe_1_1_3_U160 ( .A(npu_inst_pe_1_1_3_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_1_3_int_q_reg_v_1__0_), .S(npu_inst_pe_1_1_3_n4), .Z(
        npu_inst_pe_1_1_3_n31) );
  MUX2_X1 npu_inst_pe_1_1_3_U159 ( .A(npu_inst_pe_1_1_3_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_1_3_int_q_reg_v_3__0_), .S(npu_inst_pe_1_1_3_n4), .Z(
        npu_inst_pe_1_1_3_n30) );
  MUX2_X1 npu_inst_pe_1_1_3_U158 ( .A(npu_inst_pe_1_1_3_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_1_3_int_q_reg_v_5__0_), .S(npu_inst_pe_1_1_3_n4), .Z(
        npu_inst_pe_1_1_3_n29) );
  MUX2_X1 npu_inst_pe_1_1_3_U157 ( .A(npu_inst_pe_1_1_3_n28), .B(
        npu_inst_pe_1_1_3_n23), .S(npu_inst_pe_1_1_3_n8), .Z(
        npu_inst_pe_1_1_3_N94) );
  MUX2_X1 npu_inst_pe_1_1_3_U156 ( .A(npu_inst_pe_1_1_3_n25), .B(
        npu_inst_pe_1_1_3_n24), .S(npu_inst_pe_1_1_3_n6), .Z(
        npu_inst_pe_1_1_3_n28) );
  MUX2_X1 npu_inst_pe_1_1_3_U155 ( .A(npu_inst_pe_1_1_3_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_1_3_int_q_reg_v_1__1_), .S(npu_inst_pe_1_1_3_n4), .Z(
        npu_inst_pe_1_1_3_n25) );
  MUX2_X1 npu_inst_pe_1_1_3_U154 ( .A(npu_inst_pe_1_1_3_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_1_3_int_q_reg_v_3__1_), .S(npu_inst_pe_1_1_3_n4), .Z(
        npu_inst_pe_1_1_3_n24) );
  MUX2_X1 npu_inst_pe_1_1_3_U153 ( .A(npu_inst_pe_1_1_3_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_1_3_int_q_reg_v_5__1_), .S(npu_inst_pe_1_1_3_n4), .Z(
        npu_inst_pe_1_1_3_n23) );
  MUX2_X1 npu_inst_pe_1_1_3_U152 ( .A(npu_inst_pe_1_1_3_n22), .B(
        npu_inst_pe_1_1_3_n19), .S(npu_inst_pe_1_1_3_n8), .Z(
        npu_inst_int_data_x_1__3__1_) );
  MUX2_X1 npu_inst_pe_1_1_3_U151 ( .A(npu_inst_pe_1_1_3_n21), .B(
        npu_inst_pe_1_1_3_n20), .S(npu_inst_pe_1_1_3_n6), .Z(
        npu_inst_pe_1_1_3_n22) );
  MUX2_X1 npu_inst_pe_1_1_3_U150 ( .A(npu_inst_pe_1_1_3_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_1_3_int_q_reg_h_1__1_), .S(npu_inst_pe_1_1_3_n4), .Z(
        npu_inst_pe_1_1_3_n21) );
  MUX2_X1 npu_inst_pe_1_1_3_U149 ( .A(npu_inst_pe_1_1_3_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_1_3_int_q_reg_h_3__1_), .S(npu_inst_pe_1_1_3_n4), .Z(
        npu_inst_pe_1_1_3_n20) );
  MUX2_X1 npu_inst_pe_1_1_3_U148 ( .A(npu_inst_pe_1_1_3_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_1_3_int_q_reg_h_5__1_), .S(npu_inst_pe_1_1_3_n4), .Z(
        npu_inst_pe_1_1_3_n19) );
  MUX2_X1 npu_inst_pe_1_1_3_U147 ( .A(npu_inst_pe_1_1_3_n18), .B(
        npu_inst_pe_1_1_3_n15), .S(npu_inst_pe_1_1_3_n8), .Z(
        npu_inst_int_data_x_1__3__0_) );
  MUX2_X1 npu_inst_pe_1_1_3_U146 ( .A(npu_inst_pe_1_1_3_n17), .B(
        npu_inst_pe_1_1_3_n16), .S(npu_inst_pe_1_1_3_n6), .Z(
        npu_inst_pe_1_1_3_n18) );
  MUX2_X1 npu_inst_pe_1_1_3_U145 ( .A(npu_inst_pe_1_1_3_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_1_3_int_q_reg_h_1__0_), .S(npu_inst_pe_1_1_3_n4), .Z(
        npu_inst_pe_1_1_3_n17) );
  MUX2_X1 npu_inst_pe_1_1_3_U144 ( .A(npu_inst_pe_1_1_3_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_1_3_int_q_reg_h_3__0_), .S(npu_inst_pe_1_1_3_n4), .Z(
        npu_inst_pe_1_1_3_n16) );
  MUX2_X1 npu_inst_pe_1_1_3_U143 ( .A(npu_inst_pe_1_1_3_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_1_3_int_q_reg_h_5__0_), .S(npu_inst_pe_1_1_3_n4), .Z(
        npu_inst_pe_1_1_3_n15) );
  XOR2_X1 npu_inst_pe_1_1_3_U142 ( .A(npu_inst_pe_1_1_3_int_data_0_), .B(
        npu_inst_pe_1_1_3_int_q_acc_0_), .Z(npu_inst_pe_1_1_3_N73) );
  AND2_X1 npu_inst_pe_1_1_3_U141 ( .A1(npu_inst_pe_1_1_3_int_q_acc_0_), .A2(
        npu_inst_pe_1_1_3_int_data_0_), .ZN(npu_inst_pe_1_1_3_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_1_3_U140 ( .A(npu_inst_pe_1_1_3_int_q_acc_0_), .B(
        npu_inst_pe_1_1_3_n13), .ZN(npu_inst_pe_1_1_3_N65) );
  OR2_X1 npu_inst_pe_1_1_3_U139 ( .A1(npu_inst_pe_1_1_3_n13), .A2(
        npu_inst_pe_1_1_3_int_q_acc_0_), .ZN(npu_inst_pe_1_1_3_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_1_3_U138 ( .A(npu_inst_pe_1_1_3_int_q_acc_2_), .B(
        npu_inst_pe_1_1_3_add_69_carry_2_), .Z(npu_inst_pe_1_1_3_N75) );
  AND2_X1 npu_inst_pe_1_1_3_U137 ( .A1(npu_inst_pe_1_1_3_add_69_carry_2_), 
        .A2(npu_inst_pe_1_1_3_int_q_acc_2_), .ZN(
        npu_inst_pe_1_1_3_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_1_3_U136 ( .A(npu_inst_pe_1_1_3_int_q_acc_3_), .B(
        npu_inst_pe_1_1_3_add_69_carry_3_), .Z(npu_inst_pe_1_1_3_N76) );
  AND2_X1 npu_inst_pe_1_1_3_U135 ( .A1(npu_inst_pe_1_1_3_add_69_carry_3_), 
        .A2(npu_inst_pe_1_1_3_int_q_acc_3_), .ZN(
        npu_inst_pe_1_1_3_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_1_3_U134 ( .A(npu_inst_pe_1_1_3_int_q_acc_4_), .B(
        npu_inst_pe_1_1_3_add_69_carry_4_), .Z(npu_inst_pe_1_1_3_N77) );
  AND2_X1 npu_inst_pe_1_1_3_U133 ( .A1(npu_inst_pe_1_1_3_add_69_carry_4_), 
        .A2(npu_inst_pe_1_1_3_int_q_acc_4_), .ZN(
        npu_inst_pe_1_1_3_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_1_3_U132 ( .A(npu_inst_pe_1_1_3_int_q_acc_5_), .B(
        npu_inst_pe_1_1_3_add_69_carry_5_), .Z(npu_inst_pe_1_1_3_N78) );
  AND2_X1 npu_inst_pe_1_1_3_U131 ( .A1(npu_inst_pe_1_1_3_add_69_carry_5_), 
        .A2(npu_inst_pe_1_1_3_int_q_acc_5_), .ZN(
        npu_inst_pe_1_1_3_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_1_3_U130 ( .A(npu_inst_pe_1_1_3_int_q_acc_6_), .B(
        npu_inst_pe_1_1_3_add_69_carry_6_), .Z(npu_inst_pe_1_1_3_N79) );
  AND2_X1 npu_inst_pe_1_1_3_U129 ( .A1(npu_inst_pe_1_1_3_add_69_carry_6_), 
        .A2(npu_inst_pe_1_1_3_int_q_acc_6_), .ZN(
        npu_inst_pe_1_1_3_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_1_3_U128 ( .A(npu_inst_pe_1_1_3_int_q_acc_7_), .B(
        npu_inst_pe_1_1_3_add_69_carry_7_), .Z(npu_inst_pe_1_1_3_N80) );
  XNOR2_X1 npu_inst_pe_1_1_3_U127 ( .A(npu_inst_pe_1_1_3_sub_67_carry_2_), .B(
        npu_inst_pe_1_1_3_int_q_acc_2_), .ZN(npu_inst_pe_1_1_3_N67) );
  OR2_X1 npu_inst_pe_1_1_3_U126 ( .A1(npu_inst_pe_1_1_3_int_q_acc_2_), .A2(
        npu_inst_pe_1_1_3_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_1_3_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_1_3_U125 ( .A(npu_inst_pe_1_1_3_sub_67_carry_3_), .B(
        npu_inst_pe_1_1_3_int_q_acc_3_), .ZN(npu_inst_pe_1_1_3_N68) );
  OR2_X1 npu_inst_pe_1_1_3_U124 ( .A1(npu_inst_pe_1_1_3_int_q_acc_3_), .A2(
        npu_inst_pe_1_1_3_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_1_3_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_1_3_U123 ( .A(npu_inst_pe_1_1_3_sub_67_carry_4_), .B(
        npu_inst_pe_1_1_3_int_q_acc_4_), .ZN(npu_inst_pe_1_1_3_N69) );
  OR2_X1 npu_inst_pe_1_1_3_U122 ( .A1(npu_inst_pe_1_1_3_int_q_acc_4_), .A2(
        npu_inst_pe_1_1_3_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_1_3_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_1_3_U121 ( .A(npu_inst_pe_1_1_3_sub_67_carry_5_), .B(
        npu_inst_pe_1_1_3_int_q_acc_5_), .ZN(npu_inst_pe_1_1_3_N70) );
  OR2_X1 npu_inst_pe_1_1_3_U120 ( .A1(npu_inst_pe_1_1_3_int_q_acc_5_), .A2(
        npu_inst_pe_1_1_3_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_1_3_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_1_3_U119 ( .A(npu_inst_pe_1_1_3_sub_67_carry_6_), .B(
        npu_inst_pe_1_1_3_int_q_acc_6_), .ZN(npu_inst_pe_1_1_3_N71) );
  OR2_X1 npu_inst_pe_1_1_3_U118 ( .A1(npu_inst_pe_1_1_3_int_q_acc_6_), .A2(
        npu_inst_pe_1_1_3_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_1_3_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_1_3_U117 ( .A(npu_inst_pe_1_1_3_int_q_acc_7_), .B(
        npu_inst_pe_1_1_3_sub_67_carry_7_), .ZN(npu_inst_pe_1_1_3_N72) );
  INV_X1 npu_inst_pe_1_1_3_U116 ( .A(npu_inst_n79), .ZN(npu_inst_pe_1_1_3_n7)
         );
  INV_X1 npu_inst_pe_1_1_3_U115 ( .A(npu_inst_pe_1_1_3_n7), .ZN(
        npu_inst_pe_1_1_3_n6) );
  INV_X1 npu_inst_pe_1_1_3_U114 ( .A(npu_inst_n59), .ZN(npu_inst_pe_1_1_3_n3)
         );
  AOI22_X1 npu_inst_pe_1_1_3_U113 ( .A1(npu_inst_int_data_y_2__3__0_), .A2(
        npu_inst_pe_1_1_3_n58), .B1(npu_inst_pe_1_1_3_n119), .B2(
        npu_inst_pe_1_1_3_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_1_3_n57) );
  INV_X1 npu_inst_pe_1_1_3_U112 ( .A(npu_inst_pe_1_1_3_n57), .ZN(
        npu_inst_pe_1_1_3_n108) );
  AOI22_X1 npu_inst_pe_1_1_3_U111 ( .A1(npu_inst_int_data_y_2__3__0_), .A2(
        npu_inst_pe_1_1_3_n54), .B1(npu_inst_pe_1_1_3_n118), .B2(
        npu_inst_pe_1_1_3_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_1_3_n53) );
  INV_X1 npu_inst_pe_1_1_3_U110 ( .A(npu_inst_pe_1_1_3_n53), .ZN(
        npu_inst_pe_1_1_3_n109) );
  AOI22_X1 npu_inst_pe_1_1_3_U107 ( .A1(npu_inst_int_data_y_2__3__0_), .A2(
        npu_inst_pe_1_1_3_n50), .B1(npu_inst_pe_1_1_3_n117), .B2(
        npu_inst_pe_1_1_3_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_1_3_n49) );
  INV_X1 npu_inst_pe_1_1_3_U106 ( .A(npu_inst_pe_1_1_3_n49), .ZN(
        npu_inst_pe_1_1_3_n110) );
  AOI22_X1 npu_inst_pe_1_1_3_U105 ( .A1(npu_inst_int_data_y_2__3__0_), .A2(
        npu_inst_pe_1_1_3_n46), .B1(npu_inst_pe_1_1_3_n116), .B2(
        npu_inst_pe_1_1_3_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_1_3_n45) );
  INV_X1 npu_inst_pe_1_1_3_U104 ( .A(npu_inst_pe_1_1_3_n45), .ZN(
        npu_inst_pe_1_1_3_n111) );
  AOI22_X1 npu_inst_pe_1_1_3_U103 ( .A1(npu_inst_int_data_y_2__3__0_), .A2(
        npu_inst_pe_1_1_3_n42), .B1(npu_inst_pe_1_1_3_n115), .B2(
        npu_inst_pe_1_1_3_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_1_3_n41) );
  INV_X1 npu_inst_pe_1_1_3_U102 ( .A(npu_inst_pe_1_1_3_n41), .ZN(
        npu_inst_pe_1_1_3_n112) );
  AOI22_X1 npu_inst_pe_1_1_3_U101 ( .A1(npu_inst_int_data_y_2__3__1_), .A2(
        npu_inst_pe_1_1_3_n58), .B1(npu_inst_pe_1_1_3_n119), .B2(
        npu_inst_pe_1_1_3_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_1_3_n59) );
  INV_X1 npu_inst_pe_1_1_3_U100 ( .A(npu_inst_pe_1_1_3_n59), .ZN(
        npu_inst_pe_1_1_3_n102) );
  AOI22_X1 npu_inst_pe_1_1_3_U99 ( .A1(npu_inst_int_data_y_2__3__1_), .A2(
        npu_inst_pe_1_1_3_n54), .B1(npu_inst_pe_1_1_3_n118), .B2(
        npu_inst_pe_1_1_3_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_1_3_n55) );
  INV_X1 npu_inst_pe_1_1_3_U98 ( .A(npu_inst_pe_1_1_3_n55), .ZN(
        npu_inst_pe_1_1_3_n103) );
  AOI22_X1 npu_inst_pe_1_1_3_U97 ( .A1(npu_inst_int_data_y_2__3__1_), .A2(
        npu_inst_pe_1_1_3_n50), .B1(npu_inst_pe_1_1_3_n117), .B2(
        npu_inst_pe_1_1_3_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_1_3_n51) );
  INV_X1 npu_inst_pe_1_1_3_U96 ( .A(npu_inst_pe_1_1_3_n51), .ZN(
        npu_inst_pe_1_1_3_n104) );
  AOI22_X1 npu_inst_pe_1_1_3_U95 ( .A1(npu_inst_int_data_y_2__3__1_), .A2(
        npu_inst_pe_1_1_3_n46), .B1(npu_inst_pe_1_1_3_n116), .B2(
        npu_inst_pe_1_1_3_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_1_3_n47) );
  INV_X1 npu_inst_pe_1_1_3_U94 ( .A(npu_inst_pe_1_1_3_n47), .ZN(
        npu_inst_pe_1_1_3_n105) );
  AOI22_X1 npu_inst_pe_1_1_3_U93 ( .A1(npu_inst_int_data_y_2__3__1_), .A2(
        npu_inst_pe_1_1_3_n42), .B1(npu_inst_pe_1_1_3_n115), .B2(
        npu_inst_pe_1_1_3_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_1_3_n43) );
  INV_X1 npu_inst_pe_1_1_3_U92 ( .A(npu_inst_pe_1_1_3_n43), .ZN(
        npu_inst_pe_1_1_3_n106) );
  AOI22_X1 npu_inst_pe_1_1_3_U91 ( .A1(npu_inst_pe_1_1_3_n38), .A2(
        npu_inst_int_data_y_2__3__1_), .B1(npu_inst_pe_1_1_3_n114), .B2(
        npu_inst_pe_1_1_3_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_1_3_n39) );
  INV_X1 npu_inst_pe_1_1_3_U90 ( .A(npu_inst_pe_1_1_3_n39), .ZN(
        npu_inst_pe_1_1_3_n107) );
  AOI22_X1 npu_inst_pe_1_1_3_U89 ( .A1(npu_inst_pe_1_1_3_n38), .A2(
        npu_inst_int_data_y_2__3__0_), .B1(npu_inst_pe_1_1_3_n114), .B2(
        npu_inst_pe_1_1_3_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_1_3_n37) );
  INV_X1 npu_inst_pe_1_1_3_U88 ( .A(npu_inst_pe_1_1_3_n37), .ZN(
        npu_inst_pe_1_1_3_n113) );
  NAND2_X1 npu_inst_pe_1_1_3_U87 ( .A1(npu_inst_pe_1_1_3_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_1_3_n60), .ZN(npu_inst_pe_1_1_3_n74) );
  OAI21_X1 npu_inst_pe_1_1_3_U86 ( .B1(npu_inst_pe_1_1_3_n63), .B2(
        npu_inst_pe_1_1_3_n60), .A(npu_inst_pe_1_1_3_n74), .ZN(
        npu_inst_pe_1_1_3_n97) );
  NAND2_X1 npu_inst_pe_1_1_3_U85 ( .A1(npu_inst_pe_1_1_3_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_1_3_n60), .ZN(npu_inst_pe_1_1_3_n73) );
  OAI21_X1 npu_inst_pe_1_1_3_U84 ( .B1(npu_inst_pe_1_1_3_n61), .B2(
        npu_inst_pe_1_1_3_n60), .A(npu_inst_pe_1_1_3_n73), .ZN(
        npu_inst_pe_1_1_3_n96) );
  NAND2_X1 npu_inst_pe_1_1_3_U83 ( .A1(npu_inst_pe_1_1_3_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_1_3_n56), .ZN(npu_inst_pe_1_1_3_n72) );
  OAI21_X1 npu_inst_pe_1_1_3_U82 ( .B1(npu_inst_pe_1_1_3_n63), .B2(
        npu_inst_pe_1_1_3_n56), .A(npu_inst_pe_1_1_3_n72), .ZN(
        npu_inst_pe_1_1_3_n95) );
  NAND2_X1 npu_inst_pe_1_1_3_U81 ( .A1(npu_inst_pe_1_1_3_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_1_3_n56), .ZN(npu_inst_pe_1_1_3_n71) );
  OAI21_X1 npu_inst_pe_1_1_3_U80 ( .B1(npu_inst_pe_1_1_3_n61), .B2(
        npu_inst_pe_1_1_3_n56), .A(npu_inst_pe_1_1_3_n71), .ZN(
        npu_inst_pe_1_1_3_n94) );
  NAND2_X1 npu_inst_pe_1_1_3_U79 ( .A1(npu_inst_pe_1_1_3_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_1_3_n52), .ZN(npu_inst_pe_1_1_3_n70) );
  OAI21_X1 npu_inst_pe_1_1_3_U78 ( .B1(npu_inst_pe_1_1_3_n63), .B2(
        npu_inst_pe_1_1_3_n52), .A(npu_inst_pe_1_1_3_n70), .ZN(
        npu_inst_pe_1_1_3_n93) );
  NAND2_X1 npu_inst_pe_1_1_3_U77 ( .A1(npu_inst_pe_1_1_3_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_1_3_n52), .ZN(npu_inst_pe_1_1_3_n69) );
  OAI21_X1 npu_inst_pe_1_1_3_U76 ( .B1(npu_inst_pe_1_1_3_n61), .B2(
        npu_inst_pe_1_1_3_n52), .A(npu_inst_pe_1_1_3_n69), .ZN(
        npu_inst_pe_1_1_3_n92) );
  NAND2_X1 npu_inst_pe_1_1_3_U75 ( .A1(npu_inst_pe_1_1_3_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_1_3_n48), .ZN(npu_inst_pe_1_1_3_n68) );
  OAI21_X1 npu_inst_pe_1_1_3_U74 ( .B1(npu_inst_pe_1_1_3_n63), .B2(
        npu_inst_pe_1_1_3_n48), .A(npu_inst_pe_1_1_3_n68), .ZN(
        npu_inst_pe_1_1_3_n91) );
  NAND2_X1 npu_inst_pe_1_1_3_U73 ( .A1(npu_inst_pe_1_1_3_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_1_3_n48), .ZN(npu_inst_pe_1_1_3_n67) );
  OAI21_X1 npu_inst_pe_1_1_3_U72 ( .B1(npu_inst_pe_1_1_3_n61), .B2(
        npu_inst_pe_1_1_3_n48), .A(npu_inst_pe_1_1_3_n67), .ZN(
        npu_inst_pe_1_1_3_n90) );
  NAND2_X1 npu_inst_pe_1_1_3_U71 ( .A1(npu_inst_pe_1_1_3_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_1_3_n44), .ZN(npu_inst_pe_1_1_3_n66) );
  OAI21_X1 npu_inst_pe_1_1_3_U70 ( .B1(npu_inst_pe_1_1_3_n63), .B2(
        npu_inst_pe_1_1_3_n44), .A(npu_inst_pe_1_1_3_n66), .ZN(
        npu_inst_pe_1_1_3_n89) );
  NAND2_X1 npu_inst_pe_1_1_3_U69 ( .A1(npu_inst_pe_1_1_3_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_1_3_n44), .ZN(npu_inst_pe_1_1_3_n65) );
  OAI21_X1 npu_inst_pe_1_1_3_U68 ( .B1(npu_inst_pe_1_1_3_n61), .B2(
        npu_inst_pe_1_1_3_n44), .A(npu_inst_pe_1_1_3_n65), .ZN(
        npu_inst_pe_1_1_3_n88) );
  NAND2_X1 npu_inst_pe_1_1_3_U67 ( .A1(npu_inst_pe_1_1_3_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_1_3_n40), .ZN(npu_inst_pe_1_1_3_n64) );
  OAI21_X1 npu_inst_pe_1_1_3_U66 ( .B1(npu_inst_pe_1_1_3_n63), .B2(
        npu_inst_pe_1_1_3_n40), .A(npu_inst_pe_1_1_3_n64), .ZN(
        npu_inst_pe_1_1_3_n87) );
  NAND2_X1 npu_inst_pe_1_1_3_U65 ( .A1(npu_inst_pe_1_1_3_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_1_3_n40), .ZN(npu_inst_pe_1_1_3_n62) );
  OAI21_X1 npu_inst_pe_1_1_3_U64 ( .B1(npu_inst_pe_1_1_3_n61), .B2(
        npu_inst_pe_1_1_3_n40), .A(npu_inst_pe_1_1_3_n62), .ZN(
        npu_inst_pe_1_1_3_n86) );
  AND2_X1 npu_inst_pe_1_1_3_U63 ( .A1(npu_inst_pe_1_1_3_N93), .A2(npu_inst_n59), .ZN(npu_inst_int_data_y_1__3__0_) );
  AND2_X1 npu_inst_pe_1_1_3_U62 ( .A1(npu_inst_n59), .A2(npu_inst_pe_1_1_3_N94), .ZN(npu_inst_int_data_y_1__3__1_) );
  NOR3_X1 npu_inst_pe_1_1_3_U61 ( .A1(npu_inst_pe_1_1_3_n26), .A2(npu_inst_n59), .A3(npu_inst_int_ckg[52]), .ZN(npu_inst_pe_1_1_3_n85) );
  OR2_X1 npu_inst_pe_1_1_3_U60 ( .A1(npu_inst_pe_1_1_3_n85), .A2(
        npu_inst_pe_1_1_3_n2), .ZN(npu_inst_pe_1_1_3_N84) );
  AND2_X1 npu_inst_pe_1_1_3_U59 ( .A1(npu_inst_pe_1_1_3_int_q_acc_0_), .A2(
        npu_inst_pe_1_1_3_n1), .ZN(npu_inst_int_data_res_1__3__0_) );
  AND2_X1 npu_inst_pe_1_1_3_U58 ( .A1(npu_inst_pe_1_1_3_n2), .A2(
        npu_inst_pe_1_1_3_int_q_acc_7_), .ZN(npu_inst_int_data_res_1__3__7_)
         );
  AND2_X1 npu_inst_pe_1_1_3_U57 ( .A1(npu_inst_pe_1_1_3_int_q_acc_1_), .A2(
        npu_inst_pe_1_1_3_n1), .ZN(npu_inst_int_data_res_1__3__1_) );
  AND2_X1 npu_inst_pe_1_1_3_U56 ( .A1(npu_inst_pe_1_1_3_int_q_acc_2_), .A2(
        npu_inst_pe_1_1_3_n1), .ZN(npu_inst_int_data_res_1__3__2_) );
  AND2_X1 npu_inst_pe_1_1_3_U55 ( .A1(npu_inst_pe_1_1_3_int_q_acc_3_), .A2(
        npu_inst_pe_1_1_3_n2), .ZN(npu_inst_int_data_res_1__3__3_) );
  AND2_X1 npu_inst_pe_1_1_3_U54 ( .A1(npu_inst_pe_1_1_3_int_q_acc_4_), .A2(
        npu_inst_pe_1_1_3_n2), .ZN(npu_inst_int_data_res_1__3__4_) );
  AND2_X1 npu_inst_pe_1_1_3_U53 ( .A1(npu_inst_pe_1_1_3_int_q_acc_5_), .A2(
        npu_inst_pe_1_1_3_n2), .ZN(npu_inst_int_data_res_1__3__5_) );
  AND2_X1 npu_inst_pe_1_1_3_U52 ( .A1(npu_inst_pe_1_1_3_int_q_acc_6_), .A2(
        npu_inst_pe_1_1_3_n2), .ZN(npu_inst_int_data_res_1__3__6_) );
  AOI222_X1 npu_inst_pe_1_1_3_U51 ( .A1(npu_inst_int_data_res_2__3__0_), .A2(
        npu_inst_pe_1_1_3_n1), .B1(npu_inst_pe_1_1_3_N73), .B2(
        npu_inst_pe_1_1_3_n76), .C1(npu_inst_pe_1_1_3_N65), .C2(
        npu_inst_pe_1_1_3_n77), .ZN(npu_inst_pe_1_1_3_n84) );
  INV_X1 npu_inst_pe_1_1_3_U50 ( .A(npu_inst_pe_1_1_3_n84), .ZN(
        npu_inst_pe_1_1_3_n101) );
  AOI222_X1 npu_inst_pe_1_1_3_U49 ( .A1(npu_inst_int_data_res_2__3__7_), .A2(
        npu_inst_pe_1_1_3_n1), .B1(npu_inst_pe_1_1_3_N80), .B2(
        npu_inst_pe_1_1_3_n76), .C1(npu_inst_pe_1_1_3_N72), .C2(
        npu_inst_pe_1_1_3_n77), .ZN(npu_inst_pe_1_1_3_n75) );
  INV_X1 npu_inst_pe_1_1_3_U48 ( .A(npu_inst_pe_1_1_3_n75), .ZN(
        npu_inst_pe_1_1_3_n33) );
  AOI222_X1 npu_inst_pe_1_1_3_U47 ( .A1(npu_inst_int_data_res_2__3__1_), .A2(
        npu_inst_pe_1_1_3_n1), .B1(npu_inst_pe_1_1_3_N74), .B2(
        npu_inst_pe_1_1_3_n76), .C1(npu_inst_pe_1_1_3_N66), .C2(
        npu_inst_pe_1_1_3_n77), .ZN(npu_inst_pe_1_1_3_n83) );
  INV_X1 npu_inst_pe_1_1_3_U46 ( .A(npu_inst_pe_1_1_3_n83), .ZN(
        npu_inst_pe_1_1_3_n100) );
  AOI222_X1 npu_inst_pe_1_1_3_U45 ( .A1(npu_inst_int_data_res_2__3__2_), .A2(
        npu_inst_pe_1_1_3_n1), .B1(npu_inst_pe_1_1_3_N75), .B2(
        npu_inst_pe_1_1_3_n76), .C1(npu_inst_pe_1_1_3_N67), .C2(
        npu_inst_pe_1_1_3_n77), .ZN(npu_inst_pe_1_1_3_n82) );
  INV_X1 npu_inst_pe_1_1_3_U44 ( .A(npu_inst_pe_1_1_3_n82), .ZN(
        npu_inst_pe_1_1_3_n99) );
  AOI222_X1 npu_inst_pe_1_1_3_U43 ( .A1(npu_inst_int_data_res_2__3__3_), .A2(
        npu_inst_pe_1_1_3_n1), .B1(npu_inst_pe_1_1_3_N76), .B2(
        npu_inst_pe_1_1_3_n76), .C1(npu_inst_pe_1_1_3_N68), .C2(
        npu_inst_pe_1_1_3_n77), .ZN(npu_inst_pe_1_1_3_n81) );
  INV_X1 npu_inst_pe_1_1_3_U42 ( .A(npu_inst_pe_1_1_3_n81), .ZN(
        npu_inst_pe_1_1_3_n98) );
  AOI222_X1 npu_inst_pe_1_1_3_U41 ( .A1(npu_inst_int_data_res_2__3__4_), .A2(
        npu_inst_pe_1_1_3_n1), .B1(npu_inst_pe_1_1_3_N77), .B2(
        npu_inst_pe_1_1_3_n76), .C1(npu_inst_pe_1_1_3_N69), .C2(
        npu_inst_pe_1_1_3_n77), .ZN(npu_inst_pe_1_1_3_n80) );
  INV_X1 npu_inst_pe_1_1_3_U40 ( .A(npu_inst_pe_1_1_3_n80), .ZN(
        npu_inst_pe_1_1_3_n36) );
  AOI222_X1 npu_inst_pe_1_1_3_U39 ( .A1(npu_inst_int_data_res_2__3__5_), .A2(
        npu_inst_pe_1_1_3_n1), .B1(npu_inst_pe_1_1_3_N78), .B2(
        npu_inst_pe_1_1_3_n76), .C1(npu_inst_pe_1_1_3_N70), .C2(
        npu_inst_pe_1_1_3_n77), .ZN(npu_inst_pe_1_1_3_n79) );
  INV_X1 npu_inst_pe_1_1_3_U38 ( .A(npu_inst_pe_1_1_3_n79), .ZN(
        npu_inst_pe_1_1_3_n35) );
  AOI222_X1 npu_inst_pe_1_1_3_U37 ( .A1(npu_inst_int_data_res_2__3__6_), .A2(
        npu_inst_pe_1_1_3_n1), .B1(npu_inst_pe_1_1_3_N79), .B2(
        npu_inst_pe_1_1_3_n76), .C1(npu_inst_pe_1_1_3_N71), .C2(
        npu_inst_pe_1_1_3_n77), .ZN(npu_inst_pe_1_1_3_n78) );
  INV_X1 npu_inst_pe_1_1_3_U36 ( .A(npu_inst_pe_1_1_3_n78), .ZN(
        npu_inst_pe_1_1_3_n34) );
  INV_X1 npu_inst_pe_1_1_3_U35 ( .A(npu_inst_pe_1_1_3_int_data_1_), .ZN(
        npu_inst_pe_1_1_3_n14) );
  AND2_X1 npu_inst_pe_1_1_3_U34 ( .A1(npu_inst_int_data_x_1__3__1_), .A2(
        npu_inst_pe_1_1_3_int_q_weight_1_), .ZN(npu_inst_pe_1_1_3_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_1_3_U33 ( .A1(npu_inst_int_data_x_1__3__0_), .A2(
        npu_inst_pe_1_1_3_int_q_weight_1_), .ZN(npu_inst_pe_1_1_3_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_1_3_U32 ( .A1(npu_inst_n59), .A2(
        npu_inst_int_data_y_2__3__1_), .B1(npu_inst_pe_1_1_3_n3), .B2(
        npu_inst_int_data_x_1__4__1_), .ZN(npu_inst_pe_1_1_3_n63) );
  AOI22_X1 npu_inst_pe_1_1_3_U31 ( .A1(npu_inst_n59), .A2(
        npu_inst_int_data_y_2__3__0_), .B1(npu_inst_pe_1_1_3_n3), .B2(
        npu_inst_int_data_x_1__4__0_), .ZN(npu_inst_pe_1_1_3_n61) );
  INV_X1 npu_inst_pe_1_1_3_U30 ( .A(npu_inst_pe_1_1_3_int_data_0_), .ZN(
        npu_inst_pe_1_1_3_n13) );
  INV_X1 npu_inst_pe_1_1_3_U29 ( .A(npu_inst_n71), .ZN(npu_inst_pe_1_1_3_n5)
         );
  OR3_X1 npu_inst_pe_1_1_3_U28 ( .A1(npu_inst_pe_1_1_3_n6), .A2(
        npu_inst_pe_1_1_3_n8), .A3(npu_inst_pe_1_1_3_n5), .ZN(
        npu_inst_pe_1_1_3_n56) );
  OR3_X1 npu_inst_pe_1_1_3_U27 ( .A1(npu_inst_pe_1_1_3_n5), .A2(
        npu_inst_pe_1_1_3_n8), .A3(npu_inst_pe_1_1_3_n7), .ZN(
        npu_inst_pe_1_1_3_n48) );
  INV_X1 npu_inst_pe_1_1_3_U26 ( .A(npu_inst_pe_1_1_3_n5), .ZN(
        npu_inst_pe_1_1_3_n4) );
  OR3_X1 npu_inst_pe_1_1_3_U25 ( .A1(npu_inst_pe_1_1_3_n4), .A2(
        npu_inst_pe_1_1_3_n8), .A3(npu_inst_pe_1_1_3_n7), .ZN(
        npu_inst_pe_1_1_3_n52) );
  OR3_X1 npu_inst_pe_1_1_3_U24 ( .A1(npu_inst_pe_1_1_3_n6), .A2(
        npu_inst_pe_1_1_3_n8), .A3(npu_inst_pe_1_1_3_n4), .ZN(
        npu_inst_pe_1_1_3_n60) );
  NOR2_X1 npu_inst_pe_1_1_3_U23 ( .A1(npu_inst_pe_1_1_3_n60), .A2(
        npu_inst_pe_1_1_3_n3), .ZN(npu_inst_pe_1_1_3_n58) );
  NOR2_X1 npu_inst_pe_1_1_3_U22 ( .A1(npu_inst_pe_1_1_3_n56), .A2(
        npu_inst_pe_1_1_3_n3), .ZN(npu_inst_pe_1_1_3_n54) );
  NOR2_X1 npu_inst_pe_1_1_3_U21 ( .A1(npu_inst_pe_1_1_3_n52), .A2(
        npu_inst_pe_1_1_3_n3), .ZN(npu_inst_pe_1_1_3_n50) );
  NOR2_X1 npu_inst_pe_1_1_3_U20 ( .A1(npu_inst_pe_1_1_3_n48), .A2(
        npu_inst_pe_1_1_3_n3), .ZN(npu_inst_pe_1_1_3_n46) );
  NOR2_X1 npu_inst_pe_1_1_3_U19 ( .A1(npu_inst_pe_1_1_3_n40), .A2(
        npu_inst_pe_1_1_3_n3), .ZN(npu_inst_pe_1_1_3_n38) );
  NOR2_X1 npu_inst_pe_1_1_3_U18 ( .A1(npu_inst_pe_1_1_3_n44), .A2(
        npu_inst_pe_1_1_3_n3), .ZN(npu_inst_pe_1_1_3_n42) );
  BUF_X1 npu_inst_pe_1_1_3_U17 ( .A(npu_inst_n105), .Z(npu_inst_pe_1_1_3_n8)
         );
  INV_X1 npu_inst_pe_1_1_3_U16 ( .A(npu_inst_n126), .ZN(npu_inst_pe_1_1_3_n12)
         );
  INV_X1 npu_inst_pe_1_1_3_U15 ( .A(npu_inst_pe_1_1_3_n38), .ZN(
        npu_inst_pe_1_1_3_n114) );
  INV_X1 npu_inst_pe_1_1_3_U14 ( .A(npu_inst_pe_1_1_3_n58), .ZN(
        npu_inst_pe_1_1_3_n119) );
  INV_X1 npu_inst_pe_1_1_3_U13 ( .A(npu_inst_pe_1_1_3_n54), .ZN(
        npu_inst_pe_1_1_3_n118) );
  INV_X1 npu_inst_pe_1_1_3_U12 ( .A(npu_inst_pe_1_1_3_n50), .ZN(
        npu_inst_pe_1_1_3_n117) );
  INV_X1 npu_inst_pe_1_1_3_U11 ( .A(npu_inst_pe_1_1_3_n46), .ZN(
        npu_inst_pe_1_1_3_n116) );
  INV_X1 npu_inst_pe_1_1_3_U10 ( .A(npu_inst_pe_1_1_3_n42), .ZN(
        npu_inst_pe_1_1_3_n115) );
  BUF_X1 npu_inst_pe_1_1_3_U9 ( .A(npu_inst_n33), .Z(npu_inst_pe_1_1_3_n2) );
  BUF_X1 npu_inst_pe_1_1_3_U8 ( .A(npu_inst_n33), .Z(npu_inst_pe_1_1_3_n1) );
  BUF_X1 npu_inst_pe_1_1_3_U7 ( .A(npu_inst_pe_1_1_3_n12), .Z(
        npu_inst_pe_1_1_3_n11) );
  BUF_X1 npu_inst_pe_1_1_3_U6 ( .A(npu_inst_pe_1_1_3_n12), .Z(
        npu_inst_pe_1_1_3_n10) );
  BUF_X1 npu_inst_pe_1_1_3_U5 ( .A(npu_inst_pe_1_1_3_n12), .Z(
        npu_inst_pe_1_1_3_n9) );
  NOR2_X1 npu_inst_pe_1_1_3_U4 ( .A1(npu_inst_pe_1_1_3_int_q_weight_0_), .A2(
        npu_inst_pe_1_1_3_n1), .ZN(npu_inst_pe_1_1_3_n76) );
  NOR2_X1 npu_inst_pe_1_1_3_U3 ( .A1(npu_inst_pe_1_1_3_n27), .A2(
        npu_inst_pe_1_1_3_n1), .ZN(npu_inst_pe_1_1_3_n77) );
  FA_X1 npu_inst_pe_1_1_3_sub_67_U2_1 ( .A(npu_inst_pe_1_1_3_int_q_acc_1_), 
        .B(npu_inst_pe_1_1_3_n14), .CI(npu_inst_pe_1_1_3_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_1_3_sub_67_carry_2_), .S(npu_inst_pe_1_1_3_N66) );
  FA_X1 npu_inst_pe_1_1_3_add_69_U1_1 ( .A(npu_inst_pe_1_1_3_int_q_acc_1_), 
        .B(npu_inst_pe_1_1_3_int_data_1_), .CI(
        npu_inst_pe_1_1_3_add_69_carry_1_), .CO(
        npu_inst_pe_1_1_3_add_69_carry_2_), .S(npu_inst_pe_1_1_3_N74) );
  NAND3_X1 npu_inst_pe_1_1_3_U109 ( .A1(npu_inst_pe_1_1_3_n5), .A2(
        npu_inst_pe_1_1_3_n7), .A3(npu_inst_pe_1_1_3_n8), .ZN(
        npu_inst_pe_1_1_3_n44) );
  NAND3_X1 npu_inst_pe_1_1_3_U108 ( .A1(npu_inst_pe_1_1_3_n4), .A2(
        npu_inst_pe_1_1_3_n7), .A3(npu_inst_pe_1_1_3_n8), .ZN(
        npu_inst_pe_1_1_3_n40) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_1_3_n34), .CK(
        npu_inst_pe_1_1_3_net4309), .RN(npu_inst_pe_1_1_3_n9), .Q(
        npu_inst_pe_1_1_3_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_1_3_n35), .CK(
        npu_inst_pe_1_1_3_net4309), .RN(npu_inst_pe_1_1_3_n9), .Q(
        npu_inst_pe_1_1_3_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_1_3_n36), .CK(
        npu_inst_pe_1_1_3_net4309), .RN(npu_inst_pe_1_1_3_n9), .Q(
        npu_inst_pe_1_1_3_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_1_3_n98), .CK(
        npu_inst_pe_1_1_3_net4309), .RN(npu_inst_pe_1_1_3_n9), .Q(
        npu_inst_pe_1_1_3_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_1_3_n99), .CK(
        npu_inst_pe_1_1_3_net4309), .RN(npu_inst_pe_1_1_3_n9), .Q(
        npu_inst_pe_1_1_3_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_1_3_n100), 
        .CK(npu_inst_pe_1_1_3_net4309), .RN(npu_inst_pe_1_1_3_n9), .Q(
        npu_inst_pe_1_1_3_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_1_3_n33), .CK(
        npu_inst_pe_1_1_3_net4309), .RN(npu_inst_pe_1_1_3_n9), .Q(
        npu_inst_pe_1_1_3_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_1_3_n101), 
        .CK(npu_inst_pe_1_1_3_net4309), .RN(npu_inst_pe_1_1_3_n9), .Q(
        npu_inst_pe_1_1_3_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_weight_reg_0_ ( .D(npu_inst_n112), .CK(
        npu_inst_pe_1_1_3_net4315), .RN(npu_inst_pe_1_1_3_n9), .Q(
        npu_inst_pe_1_1_3_int_q_weight_0_), .QN(npu_inst_pe_1_1_3_n27) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_weight_reg_1_ ( .D(npu_inst_n118), .CK(
        npu_inst_pe_1_1_3_net4315), .RN(npu_inst_pe_1_1_3_n9), .Q(
        npu_inst_pe_1_1_3_int_q_weight_1_), .QN(npu_inst_pe_1_1_3_n26) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_1_3_n113), 
        .CK(npu_inst_pe_1_1_3_net4315), .RN(npu_inst_pe_1_1_3_n9), .Q(
        npu_inst_pe_1_1_3_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_1_3_n107), 
        .CK(npu_inst_pe_1_1_3_net4315), .RN(npu_inst_pe_1_1_3_n9), .Q(
        npu_inst_pe_1_1_3_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_1_3_n112), 
        .CK(npu_inst_pe_1_1_3_net4315), .RN(npu_inst_pe_1_1_3_n10), .Q(
        npu_inst_pe_1_1_3_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_1_3_n106), 
        .CK(npu_inst_pe_1_1_3_net4315), .RN(npu_inst_pe_1_1_3_n10), .Q(
        npu_inst_pe_1_1_3_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_1_3_n111), 
        .CK(npu_inst_pe_1_1_3_net4315), .RN(npu_inst_pe_1_1_3_n10), .Q(
        npu_inst_pe_1_1_3_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_1_3_n105), 
        .CK(npu_inst_pe_1_1_3_net4315), .RN(npu_inst_pe_1_1_3_n10), .Q(
        npu_inst_pe_1_1_3_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_1_3_n110), 
        .CK(npu_inst_pe_1_1_3_net4315), .RN(npu_inst_pe_1_1_3_n10), .Q(
        npu_inst_pe_1_1_3_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_1_3_n104), 
        .CK(npu_inst_pe_1_1_3_net4315), .RN(npu_inst_pe_1_1_3_n10), .Q(
        npu_inst_pe_1_1_3_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_1_3_n109), 
        .CK(npu_inst_pe_1_1_3_net4315), .RN(npu_inst_pe_1_1_3_n10), .Q(
        npu_inst_pe_1_1_3_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_1_3_n103), 
        .CK(npu_inst_pe_1_1_3_net4315), .RN(npu_inst_pe_1_1_3_n10), .Q(
        npu_inst_pe_1_1_3_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_1_3_n108), 
        .CK(npu_inst_pe_1_1_3_net4315), .RN(npu_inst_pe_1_1_3_n10), .Q(
        npu_inst_pe_1_1_3_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_1_3_n102), 
        .CK(npu_inst_pe_1_1_3_net4315), .RN(npu_inst_pe_1_1_3_n10), .Q(
        npu_inst_pe_1_1_3_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_1_3_n86), 
        .CK(npu_inst_pe_1_1_3_net4315), .RN(npu_inst_pe_1_1_3_n10), .Q(
        npu_inst_pe_1_1_3_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_1_3_n87), 
        .CK(npu_inst_pe_1_1_3_net4315), .RN(npu_inst_pe_1_1_3_n10), .Q(
        npu_inst_pe_1_1_3_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_1_3_n88), 
        .CK(npu_inst_pe_1_1_3_net4315), .RN(npu_inst_pe_1_1_3_n11), .Q(
        npu_inst_pe_1_1_3_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_1_3_n89), 
        .CK(npu_inst_pe_1_1_3_net4315), .RN(npu_inst_pe_1_1_3_n11), .Q(
        npu_inst_pe_1_1_3_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_1_3_n90), 
        .CK(npu_inst_pe_1_1_3_net4315), .RN(npu_inst_pe_1_1_3_n11), .Q(
        npu_inst_pe_1_1_3_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_1_3_n91), 
        .CK(npu_inst_pe_1_1_3_net4315), .RN(npu_inst_pe_1_1_3_n11), .Q(
        npu_inst_pe_1_1_3_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_1_3_n92), 
        .CK(npu_inst_pe_1_1_3_net4315), .RN(npu_inst_pe_1_1_3_n11), .Q(
        npu_inst_pe_1_1_3_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_1_3_n93), 
        .CK(npu_inst_pe_1_1_3_net4315), .RN(npu_inst_pe_1_1_3_n11), .Q(
        npu_inst_pe_1_1_3_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_1_3_n94), 
        .CK(npu_inst_pe_1_1_3_net4315), .RN(npu_inst_pe_1_1_3_n11), .Q(
        npu_inst_pe_1_1_3_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_1_3_n95), 
        .CK(npu_inst_pe_1_1_3_net4315), .RN(npu_inst_pe_1_1_3_n11), .Q(
        npu_inst_pe_1_1_3_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_1_3_n96), 
        .CK(npu_inst_pe_1_1_3_net4315), .RN(npu_inst_pe_1_1_3_n11), .Q(
        npu_inst_pe_1_1_3_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_1_3_n97), 
        .CK(npu_inst_pe_1_1_3_net4315), .RN(npu_inst_pe_1_1_3_n11), .Q(
        npu_inst_pe_1_1_3_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_1_3_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_1_3_N84), .SE(1'b0), .GCK(npu_inst_pe_1_1_3_net4309) );
  CLKGATETST_X1 npu_inst_pe_1_1_3_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n65), .SE(1'b0), .GCK(npu_inst_pe_1_1_3_net4315) );
  MUX2_X1 npu_inst_pe_1_1_4_U162 ( .A(npu_inst_pe_1_1_4_n32), .B(
        npu_inst_pe_1_1_4_n29), .S(npu_inst_pe_1_1_4_n8), .Z(
        npu_inst_pe_1_1_4_N93) );
  MUX2_X1 npu_inst_pe_1_1_4_U161 ( .A(npu_inst_pe_1_1_4_n31), .B(
        npu_inst_pe_1_1_4_n30), .S(npu_inst_pe_1_1_4_n6), .Z(
        npu_inst_pe_1_1_4_n32) );
  MUX2_X1 npu_inst_pe_1_1_4_U160 ( .A(npu_inst_pe_1_1_4_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_1_4_int_q_reg_v_1__0_), .S(npu_inst_pe_1_1_4_n4), .Z(
        npu_inst_pe_1_1_4_n31) );
  MUX2_X1 npu_inst_pe_1_1_4_U159 ( .A(npu_inst_pe_1_1_4_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_1_4_int_q_reg_v_3__0_), .S(npu_inst_pe_1_1_4_n4), .Z(
        npu_inst_pe_1_1_4_n30) );
  MUX2_X1 npu_inst_pe_1_1_4_U158 ( .A(npu_inst_pe_1_1_4_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_1_4_int_q_reg_v_5__0_), .S(npu_inst_pe_1_1_4_n4), .Z(
        npu_inst_pe_1_1_4_n29) );
  MUX2_X1 npu_inst_pe_1_1_4_U157 ( .A(npu_inst_pe_1_1_4_n28), .B(
        npu_inst_pe_1_1_4_n23), .S(npu_inst_pe_1_1_4_n8), .Z(
        npu_inst_pe_1_1_4_N94) );
  MUX2_X1 npu_inst_pe_1_1_4_U156 ( .A(npu_inst_pe_1_1_4_n25), .B(
        npu_inst_pe_1_1_4_n24), .S(npu_inst_pe_1_1_4_n6), .Z(
        npu_inst_pe_1_1_4_n28) );
  MUX2_X1 npu_inst_pe_1_1_4_U155 ( .A(npu_inst_pe_1_1_4_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_1_4_int_q_reg_v_1__1_), .S(npu_inst_pe_1_1_4_n4), .Z(
        npu_inst_pe_1_1_4_n25) );
  MUX2_X1 npu_inst_pe_1_1_4_U154 ( .A(npu_inst_pe_1_1_4_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_1_4_int_q_reg_v_3__1_), .S(npu_inst_pe_1_1_4_n4), .Z(
        npu_inst_pe_1_1_4_n24) );
  MUX2_X1 npu_inst_pe_1_1_4_U153 ( .A(npu_inst_pe_1_1_4_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_1_4_int_q_reg_v_5__1_), .S(npu_inst_pe_1_1_4_n4), .Z(
        npu_inst_pe_1_1_4_n23) );
  MUX2_X1 npu_inst_pe_1_1_4_U152 ( .A(npu_inst_pe_1_1_4_n22), .B(
        npu_inst_pe_1_1_4_n19), .S(npu_inst_pe_1_1_4_n8), .Z(
        npu_inst_int_data_x_1__4__1_) );
  MUX2_X1 npu_inst_pe_1_1_4_U151 ( .A(npu_inst_pe_1_1_4_n21), .B(
        npu_inst_pe_1_1_4_n20), .S(npu_inst_pe_1_1_4_n6), .Z(
        npu_inst_pe_1_1_4_n22) );
  MUX2_X1 npu_inst_pe_1_1_4_U150 ( .A(npu_inst_pe_1_1_4_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_1_4_int_q_reg_h_1__1_), .S(npu_inst_pe_1_1_4_n4), .Z(
        npu_inst_pe_1_1_4_n21) );
  MUX2_X1 npu_inst_pe_1_1_4_U149 ( .A(npu_inst_pe_1_1_4_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_1_4_int_q_reg_h_3__1_), .S(npu_inst_pe_1_1_4_n4), .Z(
        npu_inst_pe_1_1_4_n20) );
  MUX2_X1 npu_inst_pe_1_1_4_U148 ( .A(npu_inst_pe_1_1_4_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_1_4_int_q_reg_h_5__1_), .S(npu_inst_pe_1_1_4_n4), .Z(
        npu_inst_pe_1_1_4_n19) );
  MUX2_X1 npu_inst_pe_1_1_4_U147 ( .A(npu_inst_pe_1_1_4_n18), .B(
        npu_inst_pe_1_1_4_n15), .S(npu_inst_pe_1_1_4_n8), .Z(
        npu_inst_int_data_x_1__4__0_) );
  MUX2_X1 npu_inst_pe_1_1_4_U146 ( .A(npu_inst_pe_1_1_4_n17), .B(
        npu_inst_pe_1_1_4_n16), .S(npu_inst_pe_1_1_4_n6), .Z(
        npu_inst_pe_1_1_4_n18) );
  MUX2_X1 npu_inst_pe_1_1_4_U145 ( .A(npu_inst_pe_1_1_4_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_1_4_int_q_reg_h_1__0_), .S(npu_inst_pe_1_1_4_n4), .Z(
        npu_inst_pe_1_1_4_n17) );
  MUX2_X1 npu_inst_pe_1_1_4_U144 ( .A(npu_inst_pe_1_1_4_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_1_4_int_q_reg_h_3__0_), .S(npu_inst_pe_1_1_4_n4), .Z(
        npu_inst_pe_1_1_4_n16) );
  MUX2_X1 npu_inst_pe_1_1_4_U143 ( .A(npu_inst_pe_1_1_4_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_1_4_int_q_reg_h_5__0_), .S(npu_inst_pe_1_1_4_n4), .Z(
        npu_inst_pe_1_1_4_n15) );
  XOR2_X1 npu_inst_pe_1_1_4_U142 ( .A(npu_inst_pe_1_1_4_int_data_0_), .B(
        npu_inst_pe_1_1_4_int_q_acc_0_), .Z(npu_inst_pe_1_1_4_N73) );
  AND2_X1 npu_inst_pe_1_1_4_U141 ( .A1(npu_inst_pe_1_1_4_int_q_acc_0_), .A2(
        npu_inst_pe_1_1_4_int_data_0_), .ZN(npu_inst_pe_1_1_4_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_1_4_U140 ( .A(npu_inst_pe_1_1_4_int_q_acc_0_), .B(
        npu_inst_pe_1_1_4_n13), .ZN(npu_inst_pe_1_1_4_N65) );
  OR2_X1 npu_inst_pe_1_1_4_U139 ( .A1(npu_inst_pe_1_1_4_n13), .A2(
        npu_inst_pe_1_1_4_int_q_acc_0_), .ZN(npu_inst_pe_1_1_4_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_1_4_U138 ( .A(npu_inst_pe_1_1_4_int_q_acc_2_), .B(
        npu_inst_pe_1_1_4_add_69_carry_2_), .Z(npu_inst_pe_1_1_4_N75) );
  AND2_X1 npu_inst_pe_1_1_4_U137 ( .A1(npu_inst_pe_1_1_4_add_69_carry_2_), 
        .A2(npu_inst_pe_1_1_4_int_q_acc_2_), .ZN(
        npu_inst_pe_1_1_4_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_1_4_U136 ( .A(npu_inst_pe_1_1_4_int_q_acc_3_), .B(
        npu_inst_pe_1_1_4_add_69_carry_3_), .Z(npu_inst_pe_1_1_4_N76) );
  AND2_X1 npu_inst_pe_1_1_4_U135 ( .A1(npu_inst_pe_1_1_4_add_69_carry_3_), 
        .A2(npu_inst_pe_1_1_4_int_q_acc_3_), .ZN(
        npu_inst_pe_1_1_4_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_1_4_U134 ( .A(npu_inst_pe_1_1_4_int_q_acc_4_), .B(
        npu_inst_pe_1_1_4_add_69_carry_4_), .Z(npu_inst_pe_1_1_4_N77) );
  AND2_X1 npu_inst_pe_1_1_4_U133 ( .A1(npu_inst_pe_1_1_4_add_69_carry_4_), 
        .A2(npu_inst_pe_1_1_4_int_q_acc_4_), .ZN(
        npu_inst_pe_1_1_4_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_1_4_U132 ( .A(npu_inst_pe_1_1_4_int_q_acc_5_), .B(
        npu_inst_pe_1_1_4_add_69_carry_5_), .Z(npu_inst_pe_1_1_4_N78) );
  AND2_X1 npu_inst_pe_1_1_4_U131 ( .A1(npu_inst_pe_1_1_4_add_69_carry_5_), 
        .A2(npu_inst_pe_1_1_4_int_q_acc_5_), .ZN(
        npu_inst_pe_1_1_4_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_1_4_U130 ( .A(npu_inst_pe_1_1_4_int_q_acc_6_), .B(
        npu_inst_pe_1_1_4_add_69_carry_6_), .Z(npu_inst_pe_1_1_4_N79) );
  AND2_X1 npu_inst_pe_1_1_4_U129 ( .A1(npu_inst_pe_1_1_4_add_69_carry_6_), 
        .A2(npu_inst_pe_1_1_4_int_q_acc_6_), .ZN(
        npu_inst_pe_1_1_4_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_1_4_U128 ( .A(npu_inst_pe_1_1_4_int_q_acc_7_), .B(
        npu_inst_pe_1_1_4_add_69_carry_7_), .Z(npu_inst_pe_1_1_4_N80) );
  XNOR2_X1 npu_inst_pe_1_1_4_U127 ( .A(npu_inst_pe_1_1_4_sub_67_carry_2_), .B(
        npu_inst_pe_1_1_4_int_q_acc_2_), .ZN(npu_inst_pe_1_1_4_N67) );
  OR2_X1 npu_inst_pe_1_1_4_U126 ( .A1(npu_inst_pe_1_1_4_int_q_acc_2_), .A2(
        npu_inst_pe_1_1_4_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_1_4_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_1_4_U125 ( .A(npu_inst_pe_1_1_4_sub_67_carry_3_), .B(
        npu_inst_pe_1_1_4_int_q_acc_3_), .ZN(npu_inst_pe_1_1_4_N68) );
  OR2_X1 npu_inst_pe_1_1_4_U124 ( .A1(npu_inst_pe_1_1_4_int_q_acc_3_), .A2(
        npu_inst_pe_1_1_4_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_1_4_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_1_4_U123 ( .A(npu_inst_pe_1_1_4_sub_67_carry_4_), .B(
        npu_inst_pe_1_1_4_int_q_acc_4_), .ZN(npu_inst_pe_1_1_4_N69) );
  OR2_X1 npu_inst_pe_1_1_4_U122 ( .A1(npu_inst_pe_1_1_4_int_q_acc_4_), .A2(
        npu_inst_pe_1_1_4_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_1_4_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_1_4_U121 ( .A(npu_inst_pe_1_1_4_sub_67_carry_5_), .B(
        npu_inst_pe_1_1_4_int_q_acc_5_), .ZN(npu_inst_pe_1_1_4_N70) );
  OR2_X1 npu_inst_pe_1_1_4_U120 ( .A1(npu_inst_pe_1_1_4_int_q_acc_5_), .A2(
        npu_inst_pe_1_1_4_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_1_4_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_1_4_U119 ( .A(npu_inst_pe_1_1_4_sub_67_carry_6_), .B(
        npu_inst_pe_1_1_4_int_q_acc_6_), .ZN(npu_inst_pe_1_1_4_N71) );
  OR2_X1 npu_inst_pe_1_1_4_U118 ( .A1(npu_inst_pe_1_1_4_int_q_acc_6_), .A2(
        npu_inst_pe_1_1_4_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_1_4_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_1_4_U117 ( .A(npu_inst_pe_1_1_4_int_q_acc_7_), .B(
        npu_inst_pe_1_1_4_sub_67_carry_7_), .ZN(npu_inst_pe_1_1_4_N72) );
  INV_X1 npu_inst_pe_1_1_4_U116 ( .A(npu_inst_n79), .ZN(npu_inst_pe_1_1_4_n7)
         );
  INV_X1 npu_inst_pe_1_1_4_U115 ( .A(npu_inst_pe_1_1_4_n7), .ZN(
        npu_inst_pe_1_1_4_n6) );
  INV_X1 npu_inst_pe_1_1_4_U114 ( .A(npu_inst_n59), .ZN(npu_inst_pe_1_1_4_n3)
         );
  AOI22_X1 npu_inst_pe_1_1_4_U113 ( .A1(npu_inst_int_data_y_2__4__0_), .A2(
        npu_inst_pe_1_1_4_n58), .B1(npu_inst_pe_1_1_4_n119), .B2(
        npu_inst_pe_1_1_4_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_1_4_n57) );
  INV_X1 npu_inst_pe_1_1_4_U112 ( .A(npu_inst_pe_1_1_4_n57), .ZN(
        npu_inst_pe_1_1_4_n108) );
  AOI22_X1 npu_inst_pe_1_1_4_U111 ( .A1(npu_inst_int_data_y_2__4__0_), .A2(
        npu_inst_pe_1_1_4_n54), .B1(npu_inst_pe_1_1_4_n118), .B2(
        npu_inst_pe_1_1_4_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_1_4_n53) );
  INV_X1 npu_inst_pe_1_1_4_U110 ( .A(npu_inst_pe_1_1_4_n53), .ZN(
        npu_inst_pe_1_1_4_n109) );
  AOI22_X1 npu_inst_pe_1_1_4_U107 ( .A1(npu_inst_int_data_y_2__4__0_), .A2(
        npu_inst_pe_1_1_4_n50), .B1(npu_inst_pe_1_1_4_n117), .B2(
        npu_inst_pe_1_1_4_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_1_4_n49) );
  INV_X1 npu_inst_pe_1_1_4_U106 ( .A(npu_inst_pe_1_1_4_n49), .ZN(
        npu_inst_pe_1_1_4_n110) );
  AOI22_X1 npu_inst_pe_1_1_4_U105 ( .A1(npu_inst_int_data_y_2__4__0_), .A2(
        npu_inst_pe_1_1_4_n46), .B1(npu_inst_pe_1_1_4_n116), .B2(
        npu_inst_pe_1_1_4_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_1_4_n45) );
  INV_X1 npu_inst_pe_1_1_4_U104 ( .A(npu_inst_pe_1_1_4_n45), .ZN(
        npu_inst_pe_1_1_4_n111) );
  AOI22_X1 npu_inst_pe_1_1_4_U103 ( .A1(npu_inst_int_data_y_2__4__0_), .A2(
        npu_inst_pe_1_1_4_n42), .B1(npu_inst_pe_1_1_4_n115), .B2(
        npu_inst_pe_1_1_4_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_1_4_n41) );
  INV_X1 npu_inst_pe_1_1_4_U102 ( .A(npu_inst_pe_1_1_4_n41), .ZN(
        npu_inst_pe_1_1_4_n112) );
  AOI22_X1 npu_inst_pe_1_1_4_U101 ( .A1(npu_inst_int_data_y_2__4__1_), .A2(
        npu_inst_pe_1_1_4_n58), .B1(npu_inst_pe_1_1_4_n119), .B2(
        npu_inst_pe_1_1_4_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_1_4_n59) );
  INV_X1 npu_inst_pe_1_1_4_U100 ( .A(npu_inst_pe_1_1_4_n59), .ZN(
        npu_inst_pe_1_1_4_n102) );
  AOI22_X1 npu_inst_pe_1_1_4_U99 ( .A1(npu_inst_int_data_y_2__4__1_), .A2(
        npu_inst_pe_1_1_4_n54), .B1(npu_inst_pe_1_1_4_n118), .B2(
        npu_inst_pe_1_1_4_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_1_4_n55) );
  INV_X1 npu_inst_pe_1_1_4_U98 ( .A(npu_inst_pe_1_1_4_n55), .ZN(
        npu_inst_pe_1_1_4_n103) );
  AOI22_X1 npu_inst_pe_1_1_4_U97 ( .A1(npu_inst_int_data_y_2__4__1_), .A2(
        npu_inst_pe_1_1_4_n50), .B1(npu_inst_pe_1_1_4_n117), .B2(
        npu_inst_pe_1_1_4_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_1_4_n51) );
  INV_X1 npu_inst_pe_1_1_4_U96 ( .A(npu_inst_pe_1_1_4_n51), .ZN(
        npu_inst_pe_1_1_4_n104) );
  AOI22_X1 npu_inst_pe_1_1_4_U95 ( .A1(npu_inst_int_data_y_2__4__1_), .A2(
        npu_inst_pe_1_1_4_n46), .B1(npu_inst_pe_1_1_4_n116), .B2(
        npu_inst_pe_1_1_4_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_1_4_n47) );
  INV_X1 npu_inst_pe_1_1_4_U94 ( .A(npu_inst_pe_1_1_4_n47), .ZN(
        npu_inst_pe_1_1_4_n105) );
  AOI22_X1 npu_inst_pe_1_1_4_U93 ( .A1(npu_inst_int_data_y_2__4__1_), .A2(
        npu_inst_pe_1_1_4_n42), .B1(npu_inst_pe_1_1_4_n115), .B2(
        npu_inst_pe_1_1_4_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_1_4_n43) );
  INV_X1 npu_inst_pe_1_1_4_U92 ( .A(npu_inst_pe_1_1_4_n43), .ZN(
        npu_inst_pe_1_1_4_n106) );
  AOI22_X1 npu_inst_pe_1_1_4_U91 ( .A1(npu_inst_pe_1_1_4_n38), .A2(
        npu_inst_int_data_y_2__4__1_), .B1(npu_inst_pe_1_1_4_n114), .B2(
        npu_inst_pe_1_1_4_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_1_4_n39) );
  INV_X1 npu_inst_pe_1_1_4_U90 ( .A(npu_inst_pe_1_1_4_n39), .ZN(
        npu_inst_pe_1_1_4_n107) );
  AOI22_X1 npu_inst_pe_1_1_4_U89 ( .A1(npu_inst_pe_1_1_4_n38), .A2(
        npu_inst_int_data_y_2__4__0_), .B1(npu_inst_pe_1_1_4_n114), .B2(
        npu_inst_pe_1_1_4_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_1_4_n37) );
  INV_X1 npu_inst_pe_1_1_4_U88 ( .A(npu_inst_pe_1_1_4_n37), .ZN(
        npu_inst_pe_1_1_4_n113) );
  NAND2_X1 npu_inst_pe_1_1_4_U87 ( .A1(npu_inst_pe_1_1_4_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_1_4_n60), .ZN(npu_inst_pe_1_1_4_n74) );
  OAI21_X1 npu_inst_pe_1_1_4_U86 ( .B1(npu_inst_pe_1_1_4_n63), .B2(
        npu_inst_pe_1_1_4_n60), .A(npu_inst_pe_1_1_4_n74), .ZN(
        npu_inst_pe_1_1_4_n97) );
  NAND2_X1 npu_inst_pe_1_1_4_U85 ( .A1(npu_inst_pe_1_1_4_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_1_4_n60), .ZN(npu_inst_pe_1_1_4_n73) );
  OAI21_X1 npu_inst_pe_1_1_4_U84 ( .B1(npu_inst_pe_1_1_4_n61), .B2(
        npu_inst_pe_1_1_4_n60), .A(npu_inst_pe_1_1_4_n73), .ZN(
        npu_inst_pe_1_1_4_n96) );
  NAND2_X1 npu_inst_pe_1_1_4_U83 ( .A1(npu_inst_pe_1_1_4_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_1_4_n56), .ZN(npu_inst_pe_1_1_4_n72) );
  OAI21_X1 npu_inst_pe_1_1_4_U82 ( .B1(npu_inst_pe_1_1_4_n63), .B2(
        npu_inst_pe_1_1_4_n56), .A(npu_inst_pe_1_1_4_n72), .ZN(
        npu_inst_pe_1_1_4_n95) );
  NAND2_X1 npu_inst_pe_1_1_4_U81 ( .A1(npu_inst_pe_1_1_4_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_1_4_n56), .ZN(npu_inst_pe_1_1_4_n71) );
  OAI21_X1 npu_inst_pe_1_1_4_U80 ( .B1(npu_inst_pe_1_1_4_n61), .B2(
        npu_inst_pe_1_1_4_n56), .A(npu_inst_pe_1_1_4_n71), .ZN(
        npu_inst_pe_1_1_4_n94) );
  NAND2_X1 npu_inst_pe_1_1_4_U79 ( .A1(npu_inst_pe_1_1_4_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_1_4_n52), .ZN(npu_inst_pe_1_1_4_n70) );
  OAI21_X1 npu_inst_pe_1_1_4_U78 ( .B1(npu_inst_pe_1_1_4_n63), .B2(
        npu_inst_pe_1_1_4_n52), .A(npu_inst_pe_1_1_4_n70), .ZN(
        npu_inst_pe_1_1_4_n93) );
  NAND2_X1 npu_inst_pe_1_1_4_U77 ( .A1(npu_inst_pe_1_1_4_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_1_4_n52), .ZN(npu_inst_pe_1_1_4_n69) );
  OAI21_X1 npu_inst_pe_1_1_4_U76 ( .B1(npu_inst_pe_1_1_4_n61), .B2(
        npu_inst_pe_1_1_4_n52), .A(npu_inst_pe_1_1_4_n69), .ZN(
        npu_inst_pe_1_1_4_n92) );
  NAND2_X1 npu_inst_pe_1_1_4_U75 ( .A1(npu_inst_pe_1_1_4_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_1_4_n48), .ZN(npu_inst_pe_1_1_4_n68) );
  OAI21_X1 npu_inst_pe_1_1_4_U74 ( .B1(npu_inst_pe_1_1_4_n63), .B2(
        npu_inst_pe_1_1_4_n48), .A(npu_inst_pe_1_1_4_n68), .ZN(
        npu_inst_pe_1_1_4_n91) );
  NAND2_X1 npu_inst_pe_1_1_4_U73 ( .A1(npu_inst_pe_1_1_4_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_1_4_n48), .ZN(npu_inst_pe_1_1_4_n67) );
  OAI21_X1 npu_inst_pe_1_1_4_U72 ( .B1(npu_inst_pe_1_1_4_n61), .B2(
        npu_inst_pe_1_1_4_n48), .A(npu_inst_pe_1_1_4_n67), .ZN(
        npu_inst_pe_1_1_4_n90) );
  NAND2_X1 npu_inst_pe_1_1_4_U71 ( .A1(npu_inst_pe_1_1_4_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_1_4_n44), .ZN(npu_inst_pe_1_1_4_n66) );
  OAI21_X1 npu_inst_pe_1_1_4_U70 ( .B1(npu_inst_pe_1_1_4_n63), .B2(
        npu_inst_pe_1_1_4_n44), .A(npu_inst_pe_1_1_4_n66), .ZN(
        npu_inst_pe_1_1_4_n89) );
  NAND2_X1 npu_inst_pe_1_1_4_U69 ( .A1(npu_inst_pe_1_1_4_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_1_4_n44), .ZN(npu_inst_pe_1_1_4_n65) );
  OAI21_X1 npu_inst_pe_1_1_4_U68 ( .B1(npu_inst_pe_1_1_4_n61), .B2(
        npu_inst_pe_1_1_4_n44), .A(npu_inst_pe_1_1_4_n65), .ZN(
        npu_inst_pe_1_1_4_n88) );
  NAND2_X1 npu_inst_pe_1_1_4_U67 ( .A1(npu_inst_pe_1_1_4_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_1_4_n40), .ZN(npu_inst_pe_1_1_4_n64) );
  OAI21_X1 npu_inst_pe_1_1_4_U66 ( .B1(npu_inst_pe_1_1_4_n63), .B2(
        npu_inst_pe_1_1_4_n40), .A(npu_inst_pe_1_1_4_n64), .ZN(
        npu_inst_pe_1_1_4_n87) );
  NAND2_X1 npu_inst_pe_1_1_4_U65 ( .A1(npu_inst_pe_1_1_4_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_1_4_n40), .ZN(npu_inst_pe_1_1_4_n62) );
  OAI21_X1 npu_inst_pe_1_1_4_U64 ( .B1(npu_inst_pe_1_1_4_n61), .B2(
        npu_inst_pe_1_1_4_n40), .A(npu_inst_pe_1_1_4_n62), .ZN(
        npu_inst_pe_1_1_4_n86) );
  AND2_X1 npu_inst_pe_1_1_4_U63 ( .A1(npu_inst_pe_1_1_4_N93), .A2(npu_inst_n59), .ZN(npu_inst_int_data_y_1__4__0_) );
  AND2_X1 npu_inst_pe_1_1_4_U62 ( .A1(npu_inst_n59), .A2(npu_inst_pe_1_1_4_N94), .ZN(npu_inst_int_data_y_1__4__1_) );
  NOR3_X1 npu_inst_pe_1_1_4_U61 ( .A1(npu_inst_pe_1_1_4_n26), .A2(npu_inst_n59), .A3(npu_inst_int_ckg[51]), .ZN(npu_inst_pe_1_1_4_n85) );
  OR2_X1 npu_inst_pe_1_1_4_U60 ( .A1(npu_inst_pe_1_1_4_n85), .A2(
        npu_inst_pe_1_1_4_n2), .ZN(npu_inst_pe_1_1_4_N84) );
  AND2_X1 npu_inst_pe_1_1_4_U59 ( .A1(npu_inst_pe_1_1_4_int_q_acc_0_), .A2(
        npu_inst_pe_1_1_4_n1), .ZN(npu_inst_int_data_res_1__4__0_) );
  AND2_X1 npu_inst_pe_1_1_4_U58 ( .A1(npu_inst_pe_1_1_4_n2), .A2(
        npu_inst_pe_1_1_4_int_q_acc_7_), .ZN(npu_inst_int_data_res_1__4__7_)
         );
  AND2_X1 npu_inst_pe_1_1_4_U57 ( .A1(npu_inst_pe_1_1_4_int_q_acc_1_), .A2(
        npu_inst_pe_1_1_4_n1), .ZN(npu_inst_int_data_res_1__4__1_) );
  AND2_X1 npu_inst_pe_1_1_4_U56 ( .A1(npu_inst_pe_1_1_4_int_q_acc_2_), .A2(
        npu_inst_pe_1_1_4_n1), .ZN(npu_inst_int_data_res_1__4__2_) );
  AND2_X1 npu_inst_pe_1_1_4_U55 ( .A1(npu_inst_pe_1_1_4_int_q_acc_3_), .A2(
        npu_inst_pe_1_1_4_n2), .ZN(npu_inst_int_data_res_1__4__3_) );
  AND2_X1 npu_inst_pe_1_1_4_U54 ( .A1(npu_inst_pe_1_1_4_int_q_acc_4_), .A2(
        npu_inst_pe_1_1_4_n2), .ZN(npu_inst_int_data_res_1__4__4_) );
  AND2_X1 npu_inst_pe_1_1_4_U53 ( .A1(npu_inst_pe_1_1_4_int_q_acc_5_), .A2(
        npu_inst_pe_1_1_4_n2), .ZN(npu_inst_int_data_res_1__4__5_) );
  AND2_X1 npu_inst_pe_1_1_4_U52 ( .A1(npu_inst_pe_1_1_4_int_q_acc_6_), .A2(
        npu_inst_pe_1_1_4_n2), .ZN(npu_inst_int_data_res_1__4__6_) );
  AOI222_X1 npu_inst_pe_1_1_4_U51 ( .A1(npu_inst_int_data_res_2__4__0_), .A2(
        npu_inst_pe_1_1_4_n1), .B1(npu_inst_pe_1_1_4_N73), .B2(
        npu_inst_pe_1_1_4_n76), .C1(npu_inst_pe_1_1_4_N65), .C2(
        npu_inst_pe_1_1_4_n77), .ZN(npu_inst_pe_1_1_4_n84) );
  INV_X1 npu_inst_pe_1_1_4_U50 ( .A(npu_inst_pe_1_1_4_n84), .ZN(
        npu_inst_pe_1_1_4_n101) );
  AOI222_X1 npu_inst_pe_1_1_4_U49 ( .A1(npu_inst_int_data_res_2__4__7_), .A2(
        npu_inst_pe_1_1_4_n1), .B1(npu_inst_pe_1_1_4_N80), .B2(
        npu_inst_pe_1_1_4_n76), .C1(npu_inst_pe_1_1_4_N72), .C2(
        npu_inst_pe_1_1_4_n77), .ZN(npu_inst_pe_1_1_4_n75) );
  INV_X1 npu_inst_pe_1_1_4_U48 ( .A(npu_inst_pe_1_1_4_n75), .ZN(
        npu_inst_pe_1_1_4_n33) );
  AOI222_X1 npu_inst_pe_1_1_4_U47 ( .A1(npu_inst_int_data_res_2__4__1_), .A2(
        npu_inst_pe_1_1_4_n1), .B1(npu_inst_pe_1_1_4_N74), .B2(
        npu_inst_pe_1_1_4_n76), .C1(npu_inst_pe_1_1_4_N66), .C2(
        npu_inst_pe_1_1_4_n77), .ZN(npu_inst_pe_1_1_4_n83) );
  INV_X1 npu_inst_pe_1_1_4_U46 ( .A(npu_inst_pe_1_1_4_n83), .ZN(
        npu_inst_pe_1_1_4_n100) );
  AOI222_X1 npu_inst_pe_1_1_4_U45 ( .A1(npu_inst_int_data_res_2__4__2_), .A2(
        npu_inst_pe_1_1_4_n1), .B1(npu_inst_pe_1_1_4_N75), .B2(
        npu_inst_pe_1_1_4_n76), .C1(npu_inst_pe_1_1_4_N67), .C2(
        npu_inst_pe_1_1_4_n77), .ZN(npu_inst_pe_1_1_4_n82) );
  INV_X1 npu_inst_pe_1_1_4_U44 ( .A(npu_inst_pe_1_1_4_n82), .ZN(
        npu_inst_pe_1_1_4_n99) );
  AOI222_X1 npu_inst_pe_1_1_4_U43 ( .A1(npu_inst_int_data_res_2__4__3_), .A2(
        npu_inst_pe_1_1_4_n1), .B1(npu_inst_pe_1_1_4_N76), .B2(
        npu_inst_pe_1_1_4_n76), .C1(npu_inst_pe_1_1_4_N68), .C2(
        npu_inst_pe_1_1_4_n77), .ZN(npu_inst_pe_1_1_4_n81) );
  INV_X1 npu_inst_pe_1_1_4_U42 ( .A(npu_inst_pe_1_1_4_n81), .ZN(
        npu_inst_pe_1_1_4_n98) );
  AOI222_X1 npu_inst_pe_1_1_4_U41 ( .A1(npu_inst_int_data_res_2__4__4_), .A2(
        npu_inst_pe_1_1_4_n1), .B1(npu_inst_pe_1_1_4_N77), .B2(
        npu_inst_pe_1_1_4_n76), .C1(npu_inst_pe_1_1_4_N69), .C2(
        npu_inst_pe_1_1_4_n77), .ZN(npu_inst_pe_1_1_4_n80) );
  INV_X1 npu_inst_pe_1_1_4_U40 ( .A(npu_inst_pe_1_1_4_n80), .ZN(
        npu_inst_pe_1_1_4_n36) );
  AOI222_X1 npu_inst_pe_1_1_4_U39 ( .A1(npu_inst_int_data_res_2__4__5_), .A2(
        npu_inst_pe_1_1_4_n1), .B1(npu_inst_pe_1_1_4_N78), .B2(
        npu_inst_pe_1_1_4_n76), .C1(npu_inst_pe_1_1_4_N70), .C2(
        npu_inst_pe_1_1_4_n77), .ZN(npu_inst_pe_1_1_4_n79) );
  INV_X1 npu_inst_pe_1_1_4_U38 ( .A(npu_inst_pe_1_1_4_n79), .ZN(
        npu_inst_pe_1_1_4_n35) );
  AOI222_X1 npu_inst_pe_1_1_4_U37 ( .A1(npu_inst_int_data_res_2__4__6_), .A2(
        npu_inst_pe_1_1_4_n1), .B1(npu_inst_pe_1_1_4_N79), .B2(
        npu_inst_pe_1_1_4_n76), .C1(npu_inst_pe_1_1_4_N71), .C2(
        npu_inst_pe_1_1_4_n77), .ZN(npu_inst_pe_1_1_4_n78) );
  INV_X1 npu_inst_pe_1_1_4_U36 ( .A(npu_inst_pe_1_1_4_n78), .ZN(
        npu_inst_pe_1_1_4_n34) );
  INV_X1 npu_inst_pe_1_1_4_U35 ( .A(npu_inst_pe_1_1_4_int_data_1_), .ZN(
        npu_inst_pe_1_1_4_n14) );
  AND2_X1 npu_inst_pe_1_1_4_U34 ( .A1(npu_inst_int_data_x_1__4__1_), .A2(
        npu_inst_pe_1_1_4_int_q_weight_1_), .ZN(npu_inst_pe_1_1_4_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_1_4_U33 ( .A1(npu_inst_int_data_x_1__4__0_), .A2(
        npu_inst_pe_1_1_4_int_q_weight_1_), .ZN(npu_inst_pe_1_1_4_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_1_4_U32 ( .A1(npu_inst_n59), .A2(
        npu_inst_int_data_y_2__4__1_), .B1(npu_inst_pe_1_1_4_n3), .B2(
        npu_inst_int_data_x_1__5__1_), .ZN(npu_inst_pe_1_1_4_n63) );
  AOI22_X1 npu_inst_pe_1_1_4_U31 ( .A1(npu_inst_n59), .A2(
        npu_inst_int_data_y_2__4__0_), .B1(npu_inst_pe_1_1_4_n3), .B2(
        npu_inst_int_data_x_1__5__0_), .ZN(npu_inst_pe_1_1_4_n61) );
  INV_X1 npu_inst_pe_1_1_4_U30 ( .A(npu_inst_pe_1_1_4_int_data_0_), .ZN(
        npu_inst_pe_1_1_4_n13) );
  INV_X1 npu_inst_pe_1_1_4_U29 ( .A(npu_inst_n71), .ZN(npu_inst_pe_1_1_4_n5)
         );
  OR3_X1 npu_inst_pe_1_1_4_U28 ( .A1(npu_inst_pe_1_1_4_n6), .A2(
        npu_inst_pe_1_1_4_n8), .A3(npu_inst_pe_1_1_4_n5), .ZN(
        npu_inst_pe_1_1_4_n56) );
  OR3_X1 npu_inst_pe_1_1_4_U27 ( .A1(npu_inst_pe_1_1_4_n5), .A2(
        npu_inst_pe_1_1_4_n8), .A3(npu_inst_pe_1_1_4_n7), .ZN(
        npu_inst_pe_1_1_4_n48) );
  INV_X1 npu_inst_pe_1_1_4_U26 ( .A(npu_inst_pe_1_1_4_n5), .ZN(
        npu_inst_pe_1_1_4_n4) );
  OR3_X1 npu_inst_pe_1_1_4_U25 ( .A1(npu_inst_pe_1_1_4_n4), .A2(
        npu_inst_pe_1_1_4_n8), .A3(npu_inst_pe_1_1_4_n7), .ZN(
        npu_inst_pe_1_1_4_n52) );
  OR3_X1 npu_inst_pe_1_1_4_U24 ( .A1(npu_inst_pe_1_1_4_n6), .A2(
        npu_inst_pe_1_1_4_n8), .A3(npu_inst_pe_1_1_4_n4), .ZN(
        npu_inst_pe_1_1_4_n60) );
  NOR2_X1 npu_inst_pe_1_1_4_U23 ( .A1(npu_inst_pe_1_1_4_n60), .A2(
        npu_inst_pe_1_1_4_n3), .ZN(npu_inst_pe_1_1_4_n58) );
  NOR2_X1 npu_inst_pe_1_1_4_U22 ( .A1(npu_inst_pe_1_1_4_n56), .A2(
        npu_inst_pe_1_1_4_n3), .ZN(npu_inst_pe_1_1_4_n54) );
  NOR2_X1 npu_inst_pe_1_1_4_U21 ( .A1(npu_inst_pe_1_1_4_n52), .A2(
        npu_inst_pe_1_1_4_n3), .ZN(npu_inst_pe_1_1_4_n50) );
  NOR2_X1 npu_inst_pe_1_1_4_U20 ( .A1(npu_inst_pe_1_1_4_n48), .A2(
        npu_inst_pe_1_1_4_n3), .ZN(npu_inst_pe_1_1_4_n46) );
  NOR2_X1 npu_inst_pe_1_1_4_U19 ( .A1(npu_inst_pe_1_1_4_n40), .A2(
        npu_inst_pe_1_1_4_n3), .ZN(npu_inst_pe_1_1_4_n38) );
  NOR2_X1 npu_inst_pe_1_1_4_U18 ( .A1(npu_inst_pe_1_1_4_n44), .A2(
        npu_inst_pe_1_1_4_n3), .ZN(npu_inst_pe_1_1_4_n42) );
  BUF_X1 npu_inst_pe_1_1_4_U17 ( .A(npu_inst_n104), .Z(npu_inst_pe_1_1_4_n8)
         );
  INV_X1 npu_inst_pe_1_1_4_U16 ( .A(npu_inst_n126), .ZN(npu_inst_pe_1_1_4_n12)
         );
  INV_X1 npu_inst_pe_1_1_4_U15 ( .A(npu_inst_pe_1_1_4_n38), .ZN(
        npu_inst_pe_1_1_4_n114) );
  INV_X1 npu_inst_pe_1_1_4_U14 ( .A(npu_inst_pe_1_1_4_n58), .ZN(
        npu_inst_pe_1_1_4_n119) );
  INV_X1 npu_inst_pe_1_1_4_U13 ( .A(npu_inst_pe_1_1_4_n54), .ZN(
        npu_inst_pe_1_1_4_n118) );
  INV_X1 npu_inst_pe_1_1_4_U12 ( .A(npu_inst_pe_1_1_4_n50), .ZN(
        npu_inst_pe_1_1_4_n117) );
  INV_X1 npu_inst_pe_1_1_4_U11 ( .A(npu_inst_pe_1_1_4_n46), .ZN(
        npu_inst_pe_1_1_4_n116) );
  INV_X1 npu_inst_pe_1_1_4_U10 ( .A(npu_inst_pe_1_1_4_n42), .ZN(
        npu_inst_pe_1_1_4_n115) );
  BUF_X1 npu_inst_pe_1_1_4_U9 ( .A(npu_inst_n32), .Z(npu_inst_pe_1_1_4_n2) );
  BUF_X1 npu_inst_pe_1_1_4_U8 ( .A(npu_inst_n32), .Z(npu_inst_pe_1_1_4_n1) );
  BUF_X1 npu_inst_pe_1_1_4_U7 ( .A(npu_inst_pe_1_1_4_n12), .Z(
        npu_inst_pe_1_1_4_n11) );
  BUF_X1 npu_inst_pe_1_1_4_U6 ( .A(npu_inst_pe_1_1_4_n12), .Z(
        npu_inst_pe_1_1_4_n10) );
  BUF_X1 npu_inst_pe_1_1_4_U5 ( .A(npu_inst_pe_1_1_4_n12), .Z(
        npu_inst_pe_1_1_4_n9) );
  NOR2_X1 npu_inst_pe_1_1_4_U4 ( .A1(npu_inst_pe_1_1_4_int_q_weight_0_), .A2(
        npu_inst_pe_1_1_4_n1), .ZN(npu_inst_pe_1_1_4_n76) );
  NOR2_X1 npu_inst_pe_1_1_4_U3 ( .A1(npu_inst_pe_1_1_4_n27), .A2(
        npu_inst_pe_1_1_4_n1), .ZN(npu_inst_pe_1_1_4_n77) );
  FA_X1 npu_inst_pe_1_1_4_sub_67_U2_1 ( .A(npu_inst_pe_1_1_4_int_q_acc_1_), 
        .B(npu_inst_pe_1_1_4_n14), .CI(npu_inst_pe_1_1_4_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_1_4_sub_67_carry_2_), .S(npu_inst_pe_1_1_4_N66) );
  FA_X1 npu_inst_pe_1_1_4_add_69_U1_1 ( .A(npu_inst_pe_1_1_4_int_q_acc_1_), 
        .B(npu_inst_pe_1_1_4_int_data_1_), .CI(
        npu_inst_pe_1_1_4_add_69_carry_1_), .CO(
        npu_inst_pe_1_1_4_add_69_carry_2_), .S(npu_inst_pe_1_1_4_N74) );
  NAND3_X1 npu_inst_pe_1_1_4_U109 ( .A1(npu_inst_pe_1_1_4_n5), .A2(
        npu_inst_pe_1_1_4_n7), .A3(npu_inst_pe_1_1_4_n8), .ZN(
        npu_inst_pe_1_1_4_n44) );
  NAND3_X1 npu_inst_pe_1_1_4_U108 ( .A1(npu_inst_pe_1_1_4_n4), .A2(
        npu_inst_pe_1_1_4_n7), .A3(npu_inst_pe_1_1_4_n8), .ZN(
        npu_inst_pe_1_1_4_n40) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_1_4_n34), .CK(
        npu_inst_pe_1_1_4_net4286), .RN(npu_inst_pe_1_1_4_n9), .Q(
        npu_inst_pe_1_1_4_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_1_4_n35), .CK(
        npu_inst_pe_1_1_4_net4286), .RN(npu_inst_pe_1_1_4_n9), .Q(
        npu_inst_pe_1_1_4_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_1_4_n36), .CK(
        npu_inst_pe_1_1_4_net4286), .RN(npu_inst_pe_1_1_4_n9), .Q(
        npu_inst_pe_1_1_4_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_1_4_n98), .CK(
        npu_inst_pe_1_1_4_net4286), .RN(npu_inst_pe_1_1_4_n9), .Q(
        npu_inst_pe_1_1_4_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_1_4_n99), .CK(
        npu_inst_pe_1_1_4_net4286), .RN(npu_inst_pe_1_1_4_n9), .Q(
        npu_inst_pe_1_1_4_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_1_4_n100), 
        .CK(npu_inst_pe_1_1_4_net4286), .RN(npu_inst_pe_1_1_4_n9), .Q(
        npu_inst_pe_1_1_4_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_1_4_n33), .CK(
        npu_inst_pe_1_1_4_net4286), .RN(npu_inst_pe_1_1_4_n9), .Q(
        npu_inst_pe_1_1_4_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_1_4_n101), 
        .CK(npu_inst_pe_1_1_4_net4286), .RN(npu_inst_pe_1_1_4_n9), .Q(
        npu_inst_pe_1_1_4_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_weight_reg_0_ ( .D(npu_inst_n112), .CK(
        npu_inst_pe_1_1_4_net4292), .RN(npu_inst_pe_1_1_4_n9), .Q(
        npu_inst_pe_1_1_4_int_q_weight_0_), .QN(npu_inst_pe_1_1_4_n27) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_weight_reg_1_ ( .D(npu_inst_n118), .CK(
        npu_inst_pe_1_1_4_net4292), .RN(npu_inst_pe_1_1_4_n9), .Q(
        npu_inst_pe_1_1_4_int_q_weight_1_), .QN(npu_inst_pe_1_1_4_n26) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_1_4_n113), 
        .CK(npu_inst_pe_1_1_4_net4292), .RN(npu_inst_pe_1_1_4_n9), .Q(
        npu_inst_pe_1_1_4_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_1_4_n107), 
        .CK(npu_inst_pe_1_1_4_net4292), .RN(npu_inst_pe_1_1_4_n9), .Q(
        npu_inst_pe_1_1_4_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_1_4_n112), 
        .CK(npu_inst_pe_1_1_4_net4292), .RN(npu_inst_pe_1_1_4_n10), .Q(
        npu_inst_pe_1_1_4_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_1_4_n106), 
        .CK(npu_inst_pe_1_1_4_net4292), .RN(npu_inst_pe_1_1_4_n10), .Q(
        npu_inst_pe_1_1_4_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_1_4_n111), 
        .CK(npu_inst_pe_1_1_4_net4292), .RN(npu_inst_pe_1_1_4_n10), .Q(
        npu_inst_pe_1_1_4_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_1_4_n105), 
        .CK(npu_inst_pe_1_1_4_net4292), .RN(npu_inst_pe_1_1_4_n10), .Q(
        npu_inst_pe_1_1_4_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_1_4_n110), 
        .CK(npu_inst_pe_1_1_4_net4292), .RN(npu_inst_pe_1_1_4_n10), .Q(
        npu_inst_pe_1_1_4_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_1_4_n104), 
        .CK(npu_inst_pe_1_1_4_net4292), .RN(npu_inst_pe_1_1_4_n10), .Q(
        npu_inst_pe_1_1_4_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_1_4_n109), 
        .CK(npu_inst_pe_1_1_4_net4292), .RN(npu_inst_pe_1_1_4_n10), .Q(
        npu_inst_pe_1_1_4_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_1_4_n103), 
        .CK(npu_inst_pe_1_1_4_net4292), .RN(npu_inst_pe_1_1_4_n10), .Q(
        npu_inst_pe_1_1_4_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_1_4_n108), 
        .CK(npu_inst_pe_1_1_4_net4292), .RN(npu_inst_pe_1_1_4_n10), .Q(
        npu_inst_pe_1_1_4_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_1_4_n102), 
        .CK(npu_inst_pe_1_1_4_net4292), .RN(npu_inst_pe_1_1_4_n10), .Q(
        npu_inst_pe_1_1_4_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_1_4_n86), 
        .CK(npu_inst_pe_1_1_4_net4292), .RN(npu_inst_pe_1_1_4_n10), .Q(
        npu_inst_pe_1_1_4_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_1_4_n87), 
        .CK(npu_inst_pe_1_1_4_net4292), .RN(npu_inst_pe_1_1_4_n10), .Q(
        npu_inst_pe_1_1_4_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_1_4_n88), 
        .CK(npu_inst_pe_1_1_4_net4292), .RN(npu_inst_pe_1_1_4_n11), .Q(
        npu_inst_pe_1_1_4_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_1_4_n89), 
        .CK(npu_inst_pe_1_1_4_net4292), .RN(npu_inst_pe_1_1_4_n11), .Q(
        npu_inst_pe_1_1_4_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_1_4_n90), 
        .CK(npu_inst_pe_1_1_4_net4292), .RN(npu_inst_pe_1_1_4_n11), .Q(
        npu_inst_pe_1_1_4_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_1_4_n91), 
        .CK(npu_inst_pe_1_1_4_net4292), .RN(npu_inst_pe_1_1_4_n11), .Q(
        npu_inst_pe_1_1_4_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_1_4_n92), 
        .CK(npu_inst_pe_1_1_4_net4292), .RN(npu_inst_pe_1_1_4_n11), .Q(
        npu_inst_pe_1_1_4_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_1_4_n93), 
        .CK(npu_inst_pe_1_1_4_net4292), .RN(npu_inst_pe_1_1_4_n11), .Q(
        npu_inst_pe_1_1_4_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_1_4_n94), 
        .CK(npu_inst_pe_1_1_4_net4292), .RN(npu_inst_pe_1_1_4_n11), .Q(
        npu_inst_pe_1_1_4_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_1_4_n95), 
        .CK(npu_inst_pe_1_1_4_net4292), .RN(npu_inst_pe_1_1_4_n11), .Q(
        npu_inst_pe_1_1_4_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_1_4_n96), 
        .CK(npu_inst_pe_1_1_4_net4292), .RN(npu_inst_pe_1_1_4_n11), .Q(
        npu_inst_pe_1_1_4_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_1_4_n97), 
        .CK(npu_inst_pe_1_1_4_net4292), .RN(npu_inst_pe_1_1_4_n11), .Q(
        npu_inst_pe_1_1_4_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_1_4_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_1_4_N84), .SE(1'b0), .GCK(npu_inst_pe_1_1_4_net4286) );
  CLKGATETST_X1 npu_inst_pe_1_1_4_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n65), .SE(1'b0), .GCK(npu_inst_pe_1_1_4_net4292) );
  MUX2_X1 npu_inst_pe_1_1_5_U162 ( .A(npu_inst_pe_1_1_5_n32), .B(
        npu_inst_pe_1_1_5_n29), .S(npu_inst_pe_1_1_5_n8), .Z(
        npu_inst_pe_1_1_5_N93) );
  MUX2_X1 npu_inst_pe_1_1_5_U161 ( .A(npu_inst_pe_1_1_5_n31), .B(
        npu_inst_pe_1_1_5_n30), .S(npu_inst_pe_1_1_5_n6), .Z(
        npu_inst_pe_1_1_5_n32) );
  MUX2_X1 npu_inst_pe_1_1_5_U160 ( .A(npu_inst_pe_1_1_5_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_1_5_int_q_reg_v_1__0_), .S(npu_inst_pe_1_1_5_n4), .Z(
        npu_inst_pe_1_1_5_n31) );
  MUX2_X1 npu_inst_pe_1_1_5_U159 ( .A(npu_inst_pe_1_1_5_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_1_5_int_q_reg_v_3__0_), .S(npu_inst_pe_1_1_5_n4), .Z(
        npu_inst_pe_1_1_5_n30) );
  MUX2_X1 npu_inst_pe_1_1_5_U158 ( .A(npu_inst_pe_1_1_5_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_1_5_int_q_reg_v_5__0_), .S(npu_inst_pe_1_1_5_n4), .Z(
        npu_inst_pe_1_1_5_n29) );
  MUX2_X1 npu_inst_pe_1_1_5_U157 ( .A(npu_inst_pe_1_1_5_n28), .B(
        npu_inst_pe_1_1_5_n23), .S(npu_inst_pe_1_1_5_n8), .Z(
        npu_inst_pe_1_1_5_N94) );
  MUX2_X1 npu_inst_pe_1_1_5_U156 ( .A(npu_inst_pe_1_1_5_n25), .B(
        npu_inst_pe_1_1_5_n24), .S(npu_inst_pe_1_1_5_n6), .Z(
        npu_inst_pe_1_1_5_n28) );
  MUX2_X1 npu_inst_pe_1_1_5_U155 ( .A(npu_inst_pe_1_1_5_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_1_5_int_q_reg_v_1__1_), .S(npu_inst_pe_1_1_5_n4), .Z(
        npu_inst_pe_1_1_5_n25) );
  MUX2_X1 npu_inst_pe_1_1_5_U154 ( .A(npu_inst_pe_1_1_5_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_1_5_int_q_reg_v_3__1_), .S(npu_inst_pe_1_1_5_n4), .Z(
        npu_inst_pe_1_1_5_n24) );
  MUX2_X1 npu_inst_pe_1_1_5_U153 ( .A(npu_inst_pe_1_1_5_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_1_5_int_q_reg_v_5__1_), .S(npu_inst_pe_1_1_5_n4), .Z(
        npu_inst_pe_1_1_5_n23) );
  MUX2_X1 npu_inst_pe_1_1_5_U152 ( .A(npu_inst_pe_1_1_5_n22), .B(
        npu_inst_pe_1_1_5_n19), .S(npu_inst_pe_1_1_5_n8), .Z(
        npu_inst_int_data_x_1__5__1_) );
  MUX2_X1 npu_inst_pe_1_1_5_U151 ( .A(npu_inst_pe_1_1_5_n21), .B(
        npu_inst_pe_1_1_5_n20), .S(npu_inst_pe_1_1_5_n6), .Z(
        npu_inst_pe_1_1_5_n22) );
  MUX2_X1 npu_inst_pe_1_1_5_U150 ( .A(npu_inst_pe_1_1_5_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_1_5_int_q_reg_h_1__1_), .S(npu_inst_pe_1_1_5_n4), .Z(
        npu_inst_pe_1_1_5_n21) );
  MUX2_X1 npu_inst_pe_1_1_5_U149 ( .A(npu_inst_pe_1_1_5_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_1_5_int_q_reg_h_3__1_), .S(npu_inst_pe_1_1_5_n4), .Z(
        npu_inst_pe_1_1_5_n20) );
  MUX2_X1 npu_inst_pe_1_1_5_U148 ( .A(npu_inst_pe_1_1_5_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_1_5_int_q_reg_h_5__1_), .S(npu_inst_pe_1_1_5_n4), .Z(
        npu_inst_pe_1_1_5_n19) );
  MUX2_X1 npu_inst_pe_1_1_5_U147 ( .A(npu_inst_pe_1_1_5_n18), .B(
        npu_inst_pe_1_1_5_n15), .S(npu_inst_pe_1_1_5_n8), .Z(
        npu_inst_int_data_x_1__5__0_) );
  MUX2_X1 npu_inst_pe_1_1_5_U146 ( .A(npu_inst_pe_1_1_5_n17), .B(
        npu_inst_pe_1_1_5_n16), .S(npu_inst_pe_1_1_5_n6), .Z(
        npu_inst_pe_1_1_5_n18) );
  MUX2_X1 npu_inst_pe_1_1_5_U145 ( .A(npu_inst_pe_1_1_5_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_1_5_int_q_reg_h_1__0_), .S(npu_inst_pe_1_1_5_n4), .Z(
        npu_inst_pe_1_1_5_n17) );
  MUX2_X1 npu_inst_pe_1_1_5_U144 ( .A(npu_inst_pe_1_1_5_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_1_5_int_q_reg_h_3__0_), .S(npu_inst_pe_1_1_5_n4), .Z(
        npu_inst_pe_1_1_5_n16) );
  MUX2_X1 npu_inst_pe_1_1_5_U143 ( .A(npu_inst_pe_1_1_5_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_1_5_int_q_reg_h_5__0_), .S(npu_inst_pe_1_1_5_n4), .Z(
        npu_inst_pe_1_1_5_n15) );
  XOR2_X1 npu_inst_pe_1_1_5_U142 ( .A(npu_inst_pe_1_1_5_int_data_0_), .B(
        npu_inst_pe_1_1_5_int_q_acc_0_), .Z(npu_inst_pe_1_1_5_N73) );
  AND2_X1 npu_inst_pe_1_1_5_U141 ( .A1(npu_inst_pe_1_1_5_int_q_acc_0_), .A2(
        npu_inst_pe_1_1_5_int_data_0_), .ZN(npu_inst_pe_1_1_5_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_1_5_U140 ( .A(npu_inst_pe_1_1_5_int_q_acc_0_), .B(
        npu_inst_pe_1_1_5_n13), .ZN(npu_inst_pe_1_1_5_N65) );
  OR2_X1 npu_inst_pe_1_1_5_U139 ( .A1(npu_inst_pe_1_1_5_n13), .A2(
        npu_inst_pe_1_1_5_int_q_acc_0_), .ZN(npu_inst_pe_1_1_5_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_1_5_U138 ( .A(npu_inst_pe_1_1_5_int_q_acc_2_), .B(
        npu_inst_pe_1_1_5_add_69_carry_2_), .Z(npu_inst_pe_1_1_5_N75) );
  AND2_X1 npu_inst_pe_1_1_5_U137 ( .A1(npu_inst_pe_1_1_5_add_69_carry_2_), 
        .A2(npu_inst_pe_1_1_5_int_q_acc_2_), .ZN(
        npu_inst_pe_1_1_5_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_1_5_U136 ( .A(npu_inst_pe_1_1_5_int_q_acc_3_), .B(
        npu_inst_pe_1_1_5_add_69_carry_3_), .Z(npu_inst_pe_1_1_5_N76) );
  AND2_X1 npu_inst_pe_1_1_5_U135 ( .A1(npu_inst_pe_1_1_5_add_69_carry_3_), 
        .A2(npu_inst_pe_1_1_5_int_q_acc_3_), .ZN(
        npu_inst_pe_1_1_5_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_1_5_U134 ( .A(npu_inst_pe_1_1_5_int_q_acc_4_), .B(
        npu_inst_pe_1_1_5_add_69_carry_4_), .Z(npu_inst_pe_1_1_5_N77) );
  AND2_X1 npu_inst_pe_1_1_5_U133 ( .A1(npu_inst_pe_1_1_5_add_69_carry_4_), 
        .A2(npu_inst_pe_1_1_5_int_q_acc_4_), .ZN(
        npu_inst_pe_1_1_5_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_1_5_U132 ( .A(npu_inst_pe_1_1_5_int_q_acc_5_), .B(
        npu_inst_pe_1_1_5_add_69_carry_5_), .Z(npu_inst_pe_1_1_5_N78) );
  AND2_X1 npu_inst_pe_1_1_5_U131 ( .A1(npu_inst_pe_1_1_5_add_69_carry_5_), 
        .A2(npu_inst_pe_1_1_5_int_q_acc_5_), .ZN(
        npu_inst_pe_1_1_5_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_1_5_U130 ( .A(npu_inst_pe_1_1_5_int_q_acc_6_), .B(
        npu_inst_pe_1_1_5_add_69_carry_6_), .Z(npu_inst_pe_1_1_5_N79) );
  AND2_X1 npu_inst_pe_1_1_5_U129 ( .A1(npu_inst_pe_1_1_5_add_69_carry_6_), 
        .A2(npu_inst_pe_1_1_5_int_q_acc_6_), .ZN(
        npu_inst_pe_1_1_5_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_1_5_U128 ( .A(npu_inst_pe_1_1_5_int_q_acc_7_), .B(
        npu_inst_pe_1_1_5_add_69_carry_7_), .Z(npu_inst_pe_1_1_5_N80) );
  XNOR2_X1 npu_inst_pe_1_1_5_U127 ( .A(npu_inst_pe_1_1_5_sub_67_carry_2_), .B(
        npu_inst_pe_1_1_5_int_q_acc_2_), .ZN(npu_inst_pe_1_1_5_N67) );
  OR2_X1 npu_inst_pe_1_1_5_U126 ( .A1(npu_inst_pe_1_1_5_int_q_acc_2_), .A2(
        npu_inst_pe_1_1_5_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_1_5_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_1_5_U125 ( .A(npu_inst_pe_1_1_5_sub_67_carry_3_), .B(
        npu_inst_pe_1_1_5_int_q_acc_3_), .ZN(npu_inst_pe_1_1_5_N68) );
  OR2_X1 npu_inst_pe_1_1_5_U124 ( .A1(npu_inst_pe_1_1_5_int_q_acc_3_), .A2(
        npu_inst_pe_1_1_5_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_1_5_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_1_5_U123 ( .A(npu_inst_pe_1_1_5_sub_67_carry_4_), .B(
        npu_inst_pe_1_1_5_int_q_acc_4_), .ZN(npu_inst_pe_1_1_5_N69) );
  OR2_X1 npu_inst_pe_1_1_5_U122 ( .A1(npu_inst_pe_1_1_5_int_q_acc_4_), .A2(
        npu_inst_pe_1_1_5_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_1_5_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_1_5_U121 ( .A(npu_inst_pe_1_1_5_sub_67_carry_5_), .B(
        npu_inst_pe_1_1_5_int_q_acc_5_), .ZN(npu_inst_pe_1_1_5_N70) );
  OR2_X1 npu_inst_pe_1_1_5_U120 ( .A1(npu_inst_pe_1_1_5_int_q_acc_5_), .A2(
        npu_inst_pe_1_1_5_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_1_5_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_1_5_U119 ( .A(npu_inst_pe_1_1_5_sub_67_carry_6_), .B(
        npu_inst_pe_1_1_5_int_q_acc_6_), .ZN(npu_inst_pe_1_1_5_N71) );
  OR2_X1 npu_inst_pe_1_1_5_U118 ( .A1(npu_inst_pe_1_1_5_int_q_acc_6_), .A2(
        npu_inst_pe_1_1_5_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_1_5_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_1_5_U117 ( .A(npu_inst_pe_1_1_5_int_q_acc_7_), .B(
        npu_inst_pe_1_1_5_sub_67_carry_7_), .ZN(npu_inst_pe_1_1_5_N72) );
  INV_X1 npu_inst_pe_1_1_5_U116 ( .A(npu_inst_n79), .ZN(npu_inst_pe_1_1_5_n7)
         );
  INV_X1 npu_inst_pe_1_1_5_U115 ( .A(npu_inst_pe_1_1_5_n7), .ZN(
        npu_inst_pe_1_1_5_n6) );
  INV_X1 npu_inst_pe_1_1_5_U114 ( .A(npu_inst_n59), .ZN(npu_inst_pe_1_1_5_n3)
         );
  AOI22_X1 npu_inst_pe_1_1_5_U113 ( .A1(npu_inst_int_data_y_2__5__0_), .A2(
        npu_inst_pe_1_1_5_n58), .B1(npu_inst_pe_1_1_5_n119), .B2(
        npu_inst_pe_1_1_5_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_1_5_n57) );
  INV_X1 npu_inst_pe_1_1_5_U112 ( .A(npu_inst_pe_1_1_5_n57), .ZN(
        npu_inst_pe_1_1_5_n108) );
  AOI22_X1 npu_inst_pe_1_1_5_U111 ( .A1(npu_inst_int_data_y_2__5__0_), .A2(
        npu_inst_pe_1_1_5_n54), .B1(npu_inst_pe_1_1_5_n118), .B2(
        npu_inst_pe_1_1_5_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_1_5_n53) );
  INV_X1 npu_inst_pe_1_1_5_U110 ( .A(npu_inst_pe_1_1_5_n53), .ZN(
        npu_inst_pe_1_1_5_n109) );
  AOI22_X1 npu_inst_pe_1_1_5_U107 ( .A1(npu_inst_int_data_y_2__5__0_), .A2(
        npu_inst_pe_1_1_5_n50), .B1(npu_inst_pe_1_1_5_n117), .B2(
        npu_inst_pe_1_1_5_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_1_5_n49) );
  INV_X1 npu_inst_pe_1_1_5_U106 ( .A(npu_inst_pe_1_1_5_n49), .ZN(
        npu_inst_pe_1_1_5_n110) );
  AOI22_X1 npu_inst_pe_1_1_5_U105 ( .A1(npu_inst_int_data_y_2__5__0_), .A2(
        npu_inst_pe_1_1_5_n46), .B1(npu_inst_pe_1_1_5_n116), .B2(
        npu_inst_pe_1_1_5_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_1_5_n45) );
  INV_X1 npu_inst_pe_1_1_5_U104 ( .A(npu_inst_pe_1_1_5_n45), .ZN(
        npu_inst_pe_1_1_5_n111) );
  AOI22_X1 npu_inst_pe_1_1_5_U103 ( .A1(npu_inst_int_data_y_2__5__0_), .A2(
        npu_inst_pe_1_1_5_n42), .B1(npu_inst_pe_1_1_5_n115), .B2(
        npu_inst_pe_1_1_5_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_1_5_n41) );
  INV_X1 npu_inst_pe_1_1_5_U102 ( .A(npu_inst_pe_1_1_5_n41), .ZN(
        npu_inst_pe_1_1_5_n112) );
  AOI22_X1 npu_inst_pe_1_1_5_U101 ( .A1(npu_inst_int_data_y_2__5__1_), .A2(
        npu_inst_pe_1_1_5_n58), .B1(npu_inst_pe_1_1_5_n119), .B2(
        npu_inst_pe_1_1_5_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_1_5_n59) );
  INV_X1 npu_inst_pe_1_1_5_U100 ( .A(npu_inst_pe_1_1_5_n59), .ZN(
        npu_inst_pe_1_1_5_n102) );
  AOI22_X1 npu_inst_pe_1_1_5_U99 ( .A1(npu_inst_int_data_y_2__5__1_), .A2(
        npu_inst_pe_1_1_5_n54), .B1(npu_inst_pe_1_1_5_n118), .B2(
        npu_inst_pe_1_1_5_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_1_5_n55) );
  INV_X1 npu_inst_pe_1_1_5_U98 ( .A(npu_inst_pe_1_1_5_n55), .ZN(
        npu_inst_pe_1_1_5_n103) );
  AOI22_X1 npu_inst_pe_1_1_5_U97 ( .A1(npu_inst_int_data_y_2__5__1_), .A2(
        npu_inst_pe_1_1_5_n50), .B1(npu_inst_pe_1_1_5_n117), .B2(
        npu_inst_pe_1_1_5_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_1_5_n51) );
  INV_X1 npu_inst_pe_1_1_5_U96 ( .A(npu_inst_pe_1_1_5_n51), .ZN(
        npu_inst_pe_1_1_5_n104) );
  AOI22_X1 npu_inst_pe_1_1_5_U95 ( .A1(npu_inst_int_data_y_2__5__1_), .A2(
        npu_inst_pe_1_1_5_n46), .B1(npu_inst_pe_1_1_5_n116), .B2(
        npu_inst_pe_1_1_5_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_1_5_n47) );
  INV_X1 npu_inst_pe_1_1_5_U94 ( .A(npu_inst_pe_1_1_5_n47), .ZN(
        npu_inst_pe_1_1_5_n105) );
  AOI22_X1 npu_inst_pe_1_1_5_U93 ( .A1(npu_inst_int_data_y_2__5__1_), .A2(
        npu_inst_pe_1_1_5_n42), .B1(npu_inst_pe_1_1_5_n115), .B2(
        npu_inst_pe_1_1_5_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_1_5_n43) );
  INV_X1 npu_inst_pe_1_1_5_U92 ( .A(npu_inst_pe_1_1_5_n43), .ZN(
        npu_inst_pe_1_1_5_n106) );
  AOI22_X1 npu_inst_pe_1_1_5_U91 ( .A1(npu_inst_pe_1_1_5_n38), .A2(
        npu_inst_int_data_y_2__5__1_), .B1(npu_inst_pe_1_1_5_n114), .B2(
        npu_inst_pe_1_1_5_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_1_5_n39) );
  INV_X1 npu_inst_pe_1_1_5_U90 ( .A(npu_inst_pe_1_1_5_n39), .ZN(
        npu_inst_pe_1_1_5_n107) );
  AOI22_X1 npu_inst_pe_1_1_5_U89 ( .A1(npu_inst_pe_1_1_5_n38), .A2(
        npu_inst_int_data_y_2__5__0_), .B1(npu_inst_pe_1_1_5_n114), .B2(
        npu_inst_pe_1_1_5_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_1_5_n37) );
  INV_X1 npu_inst_pe_1_1_5_U88 ( .A(npu_inst_pe_1_1_5_n37), .ZN(
        npu_inst_pe_1_1_5_n113) );
  NAND2_X1 npu_inst_pe_1_1_5_U87 ( .A1(npu_inst_pe_1_1_5_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_1_5_n60), .ZN(npu_inst_pe_1_1_5_n74) );
  OAI21_X1 npu_inst_pe_1_1_5_U86 ( .B1(npu_inst_pe_1_1_5_n63), .B2(
        npu_inst_pe_1_1_5_n60), .A(npu_inst_pe_1_1_5_n74), .ZN(
        npu_inst_pe_1_1_5_n97) );
  NAND2_X1 npu_inst_pe_1_1_5_U85 ( .A1(npu_inst_pe_1_1_5_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_1_5_n60), .ZN(npu_inst_pe_1_1_5_n73) );
  OAI21_X1 npu_inst_pe_1_1_5_U84 ( .B1(npu_inst_pe_1_1_5_n61), .B2(
        npu_inst_pe_1_1_5_n60), .A(npu_inst_pe_1_1_5_n73), .ZN(
        npu_inst_pe_1_1_5_n96) );
  NAND2_X1 npu_inst_pe_1_1_5_U83 ( .A1(npu_inst_pe_1_1_5_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_1_5_n56), .ZN(npu_inst_pe_1_1_5_n72) );
  OAI21_X1 npu_inst_pe_1_1_5_U82 ( .B1(npu_inst_pe_1_1_5_n63), .B2(
        npu_inst_pe_1_1_5_n56), .A(npu_inst_pe_1_1_5_n72), .ZN(
        npu_inst_pe_1_1_5_n95) );
  NAND2_X1 npu_inst_pe_1_1_5_U81 ( .A1(npu_inst_pe_1_1_5_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_1_5_n56), .ZN(npu_inst_pe_1_1_5_n71) );
  OAI21_X1 npu_inst_pe_1_1_5_U80 ( .B1(npu_inst_pe_1_1_5_n61), .B2(
        npu_inst_pe_1_1_5_n56), .A(npu_inst_pe_1_1_5_n71), .ZN(
        npu_inst_pe_1_1_5_n94) );
  NAND2_X1 npu_inst_pe_1_1_5_U79 ( .A1(npu_inst_pe_1_1_5_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_1_5_n52), .ZN(npu_inst_pe_1_1_5_n70) );
  OAI21_X1 npu_inst_pe_1_1_5_U78 ( .B1(npu_inst_pe_1_1_5_n63), .B2(
        npu_inst_pe_1_1_5_n52), .A(npu_inst_pe_1_1_5_n70), .ZN(
        npu_inst_pe_1_1_5_n93) );
  NAND2_X1 npu_inst_pe_1_1_5_U77 ( .A1(npu_inst_pe_1_1_5_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_1_5_n52), .ZN(npu_inst_pe_1_1_5_n69) );
  OAI21_X1 npu_inst_pe_1_1_5_U76 ( .B1(npu_inst_pe_1_1_5_n61), .B2(
        npu_inst_pe_1_1_5_n52), .A(npu_inst_pe_1_1_5_n69), .ZN(
        npu_inst_pe_1_1_5_n92) );
  NAND2_X1 npu_inst_pe_1_1_5_U75 ( .A1(npu_inst_pe_1_1_5_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_1_5_n48), .ZN(npu_inst_pe_1_1_5_n68) );
  OAI21_X1 npu_inst_pe_1_1_5_U74 ( .B1(npu_inst_pe_1_1_5_n63), .B2(
        npu_inst_pe_1_1_5_n48), .A(npu_inst_pe_1_1_5_n68), .ZN(
        npu_inst_pe_1_1_5_n91) );
  NAND2_X1 npu_inst_pe_1_1_5_U73 ( .A1(npu_inst_pe_1_1_5_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_1_5_n48), .ZN(npu_inst_pe_1_1_5_n67) );
  OAI21_X1 npu_inst_pe_1_1_5_U72 ( .B1(npu_inst_pe_1_1_5_n61), .B2(
        npu_inst_pe_1_1_5_n48), .A(npu_inst_pe_1_1_5_n67), .ZN(
        npu_inst_pe_1_1_5_n90) );
  NAND2_X1 npu_inst_pe_1_1_5_U71 ( .A1(npu_inst_pe_1_1_5_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_1_5_n44), .ZN(npu_inst_pe_1_1_5_n66) );
  OAI21_X1 npu_inst_pe_1_1_5_U70 ( .B1(npu_inst_pe_1_1_5_n63), .B2(
        npu_inst_pe_1_1_5_n44), .A(npu_inst_pe_1_1_5_n66), .ZN(
        npu_inst_pe_1_1_5_n89) );
  NAND2_X1 npu_inst_pe_1_1_5_U69 ( .A1(npu_inst_pe_1_1_5_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_1_5_n44), .ZN(npu_inst_pe_1_1_5_n65) );
  OAI21_X1 npu_inst_pe_1_1_5_U68 ( .B1(npu_inst_pe_1_1_5_n61), .B2(
        npu_inst_pe_1_1_5_n44), .A(npu_inst_pe_1_1_5_n65), .ZN(
        npu_inst_pe_1_1_5_n88) );
  NAND2_X1 npu_inst_pe_1_1_5_U67 ( .A1(npu_inst_pe_1_1_5_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_1_5_n40), .ZN(npu_inst_pe_1_1_5_n64) );
  OAI21_X1 npu_inst_pe_1_1_5_U66 ( .B1(npu_inst_pe_1_1_5_n63), .B2(
        npu_inst_pe_1_1_5_n40), .A(npu_inst_pe_1_1_5_n64), .ZN(
        npu_inst_pe_1_1_5_n87) );
  NAND2_X1 npu_inst_pe_1_1_5_U65 ( .A1(npu_inst_pe_1_1_5_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_1_5_n40), .ZN(npu_inst_pe_1_1_5_n62) );
  OAI21_X1 npu_inst_pe_1_1_5_U64 ( .B1(npu_inst_pe_1_1_5_n61), .B2(
        npu_inst_pe_1_1_5_n40), .A(npu_inst_pe_1_1_5_n62), .ZN(
        npu_inst_pe_1_1_5_n86) );
  AND2_X1 npu_inst_pe_1_1_5_U63 ( .A1(npu_inst_pe_1_1_5_N93), .A2(npu_inst_n59), .ZN(npu_inst_int_data_y_1__5__0_) );
  AND2_X1 npu_inst_pe_1_1_5_U62 ( .A1(npu_inst_n59), .A2(npu_inst_pe_1_1_5_N94), .ZN(npu_inst_int_data_y_1__5__1_) );
  NOR3_X1 npu_inst_pe_1_1_5_U61 ( .A1(npu_inst_pe_1_1_5_n26), .A2(npu_inst_n59), .A3(npu_inst_int_ckg[50]), .ZN(npu_inst_pe_1_1_5_n85) );
  OR2_X1 npu_inst_pe_1_1_5_U60 ( .A1(npu_inst_pe_1_1_5_n85), .A2(
        npu_inst_pe_1_1_5_n2), .ZN(npu_inst_pe_1_1_5_N84) );
  AND2_X1 npu_inst_pe_1_1_5_U59 ( .A1(npu_inst_pe_1_1_5_int_q_acc_0_), .A2(
        npu_inst_pe_1_1_5_n1), .ZN(npu_inst_int_data_res_1__5__0_) );
  AND2_X1 npu_inst_pe_1_1_5_U58 ( .A1(npu_inst_pe_1_1_5_n2), .A2(
        npu_inst_pe_1_1_5_int_q_acc_7_), .ZN(npu_inst_int_data_res_1__5__7_)
         );
  AND2_X1 npu_inst_pe_1_1_5_U57 ( .A1(npu_inst_pe_1_1_5_int_q_acc_1_), .A2(
        npu_inst_pe_1_1_5_n1), .ZN(npu_inst_int_data_res_1__5__1_) );
  AND2_X1 npu_inst_pe_1_1_5_U56 ( .A1(npu_inst_pe_1_1_5_int_q_acc_2_), .A2(
        npu_inst_pe_1_1_5_n1), .ZN(npu_inst_int_data_res_1__5__2_) );
  AND2_X1 npu_inst_pe_1_1_5_U55 ( .A1(npu_inst_pe_1_1_5_int_q_acc_3_), .A2(
        npu_inst_pe_1_1_5_n2), .ZN(npu_inst_int_data_res_1__5__3_) );
  AND2_X1 npu_inst_pe_1_1_5_U54 ( .A1(npu_inst_pe_1_1_5_int_q_acc_4_), .A2(
        npu_inst_pe_1_1_5_n2), .ZN(npu_inst_int_data_res_1__5__4_) );
  AND2_X1 npu_inst_pe_1_1_5_U53 ( .A1(npu_inst_pe_1_1_5_int_q_acc_5_), .A2(
        npu_inst_pe_1_1_5_n2), .ZN(npu_inst_int_data_res_1__5__5_) );
  AND2_X1 npu_inst_pe_1_1_5_U52 ( .A1(npu_inst_pe_1_1_5_int_q_acc_6_), .A2(
        npu_inst_pe_1_1_5_n2), .ZN(npu_inst_int_data_res_1__5__6_) );
  AOI222_X1 npu_inst_pe_1_1_5_U51 ( .A1(npu_inst_int_data_res_2__5__0_), .A2(
        npu_inst_pe_1_1_5_n1), .B1(npu_inst_pe_1_1_5_N73), .B2(
        npu_inst_pe_1_1_5_n76), .C1(npu_inst_pe_1_1_5_N65), .C2(
        npu_inst_pe_1_1_5_n77), .ZN(npu_inst_pe_1_1_5_n84) );
  INV_X1 npu_inst_pe_1_1_5_U50 ( .A(npu_inst_pe_1_1_5_n84), .ZN(
        npu_inst_pe_1_1_5_n101) );
  AOI222_X1 npu_inst_pe_1_1_5_U49 ( .A1(npu_inst_int_data_res_2__5__7_), .A2(
        npu_inst_pe_1_1_5_n1), .B1(npu_inst_pe_1_1_5_N80), .B2(
        npu_inst_pe_1_1_5_n76), .C1(npu_inst_pe_1_1_5_N72), .C2(
        npu_inst_pe_1_1_5_n77), .ZN(npu_inst_pe_1_1_5_n75) );
  INV_X1 npu_inst_pe_1_1_5_U48 ( .A(npu_inst_pe_1_1_5_n75), .ZN(
        npu_inst_pe_1_1_5_n33) );
  AOI222_X1 npu_inst_pe_1_1_5_U47 ( .A1(npu_inst_int_data_res_2__5__1_), .A2(
        npu_inst_pe_1_1_5_n1), .B1(npu_inst_pe_1_1_5_N74), .B2(
        npu_inst_pe_1_1_5_n76), .C1(npu_inst_pe_1_1_5_N66), .C2(
        npu_inst_pe_1_1_5_n77), .ZN(npu_inst_pe_1_1_5_n83) );
  INV_X1 npu_inst_pe_1_1_5_U46 ( .A(npu_inst_pe_1_1_5_n83), .ZN(
        npu_inst_pe_1_1_5_n100) );
  AOI222_X1 npu_inst_pe_1_1_5_U45 ( .A1(npu_inst_int_data_res_2__5__2_), .A2(
        npu_inst_pe_1_1_5_n1), .B1(npu_inst_pe_1_1_5_N75), .B2(
        npu_inst_pe_1_1_5_n76), .C1(npu_inst_pe_1_1_5_N67), .C2(
        npu_inst_pe_1_1_5_n77), .ZN(npu_inst_pe_1_1_5_n82) );
  INV_X1 npu_inst_pe_1_1_5_U44 ( .A(npu_inst_pe_1_1_5_n82), .ZN(
        npu_inst_pe_1_1_5_n99) );
  AOI222_X1 npu_inst_pe_1_1_5_U43 ( .A1(npu_inst_int_data_res_2__5__3_), .A2(
        npu_inst_pe_1_1_5_n1), .B1(npu_inst_pe_1_1_5_N76), .B2(
        npu_inst_pe_1_1_5_n76), .C1(npu_inst_pe_1_1_5_N68), .C2(
        npu_inst_pe_1_1_5_n77), .ZN(npu_inst_pe_1_1_5_n81) );
  INV_X1 npu_inst_pe_1_1_5_U42 ( .A(npu_inst_pe_1_1_5_n81), .ZN(
        npu_inst_pe_1_1_5_n98) );
  AOI222_X1 npu_inst_pe_1_1_5_U41 ( .A1(npu_inst_int_data_res_2__5__4_), .A2(
        npu_inst_pe_1_1_5_n1), .B1(npu_inst_pe_1_1_5_N77), .B2(
        npu_inst_pe_1_1_5_n76), .C1(npu_inst_pe_1_1_5_N69), .C2(
        npu_inst_pe_1_1_5_n77), .ZN(npu_inst_pe_1_1_5_n80) );
  INV_X1 npu_inst_pe_1_1_5_U40 ( .A(npu_inst_pe_1_1_5_n80), .ZN(
        npu_inst_pe_1_1_5_n36) );
  AOI222_X1 npu_inst_pe_1_1_5_U39 ( .A1(npu_inst_int_data_res_2__5__5_), .A2(
        npu_inst_pe_1_1_5_n1), .B1(npu_inst_pe_1_1_5_N78), .B2(
        npu_inst_pe_1_1_5_n76), .C1(npu_inst_pe_1_1_5_N70), .C2(
        npu_inst_pe_1_1_5_n77), .ZN(npu_inst_pe_1_1_5_n79) );
  INV_X1 npu_inst_pe_1_1_5_U38 ( .A(npu_inst_pe_1_1_5_n79), .ZN(
        npu_inst_pe_1_1_5_n35) );
  AOI222_X1 npu_inst_pe_1_1_5_U37 ( .A1(npu_inst_int_data_res_2__5__6_), .A2(
        npu_inst_pe_1_1_5_n1), .B1(npu_inst_pe_1_1_5_N79), .B2(
        npu_inst_pe_1_1_5_n76), .C1(npu_inst_pe_1_1_5_N71), .C2(
        npu_inst_pe_1_1_5_n77), .ZN(npu_inst_pe_1_1_5_n78) );
  INV_X1 npu_inst_pe_1_1_5_U36 ( .A(npu_inst_pe_1_1_5_n78), .ZN(
        npu_inst_pe_1_1_5_n34) );
  INV_X1 npu_inst_pe_1_1_5_U35 ( .A(npu_inst_pe_1_1_5_int_data_1_), .ZN(
        npu_inst_pe_1_1_5_n14) );
  AND2_X1 npu_inst_pe_1_1_5_U34 ( .A1(npu_inst_int_data_x_1__5__1_), .A2(
        npu_inst_pe_1_1_5_int_q_weight_1_), .ZN(npu_inst_pe_1_1_5_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_1_5_U33 ( .A1(npu_inst_int_data_x_1__5__0_), .A2(
        npu_inst_pe_1_1_5_int_q_weight_1_), .ZN(npu_inst_pe_1_1_5_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_1_5_U32 ( .A1(npu_inst_n59), .A2(
        npu_inst_int_data_y_2__5__1_), .B1(npu_inst_pe_1_1_5_n3), .B2(
        npu_inst_int_data_x_1__6__1_), .ZN(npu_inst_pe_1_1_5_n63) );
  AOI22_X1 npu_inst_pe_1_1_5_U31 ( .A1(npu_inst_n59), .A2(
        npu_inst_int_data_y_2__5__0_), .B1(npu_inst_pe_1_1_5_n3), .B2(
        npu_inst_int_data_x_1__6__0_), .ZN(npu_inst_pe_1_1_5_n61) );
  INV_X1 npu_inst_pe_1_1_5_U30 ( .A(npu_inst_pe_1_1_5_int_data_0_), .ZN(
        npu_inst_pe_1_1_5_n13) );
  INV_X1 npu_inst_pe_1_1_5_U29 ( .A(npu_inst_n71), .ZN(npu_inst_pe_1_1_5_n5)
         );
  OR3_X1 npu_inst_pe_1_1_5_U28 ( .A1(npu_inst_pe_1_1_5_n6), .A2(
        npu_inst_pe_1_1_5_n8), .A3(npu_inst_pe_1_1_5_n5), .ZN(
        npu_inst_pe_1_1_5_n56) );
  OR3_X1 npu_inst_pe_1_1_5_U27 ( .A1(npu_inst_pe_1_1_5_n5), .A2(
        npu_inst_pe_1_1_5_n8), .A3(npu_inst_pe_1_1_5_n7), .ZN(
        npu_inst_pe_1_1_5_n48) );
  INV_X1 npu_inst_pe_1_1_5_U26 ( .A(npu_inst_pe_1_1_5_n5), .ZN(
        npu_inst_pe_1_1_5_n4) );
  OR3_X1 npu_inst_pe_1_1_5_U25 ( .A1(npu_inst_pe_1_1_5_n4), .A2(
        npu_inst_pe_1_1_5_n8), .A3(npu_inst_pe_1_1_5_n7), .ZN(
        npu_inst_pe_1_1_5_n52) );
  OR3_X1 npu_inst_pe_1_1_5_U24 ( .A1(npu_inst_pe_1_1_5_n6), .A2(
        npu_inst_pe_1_1_5_n8), .A3(npu_inst_pe_1_1_5_n4), .ZN(
        npu_inst_pe_1_1_5_n60) );
  NOR2_X1 npu_inst_pe_1_1_5_U23 ( .A1(npu_inst_pe_1_1_5_n60), .A2(
        npu_inst_pe_1_1_5_n3), .ZN(npu_inst_pe_1_1_5_n58) );
  NOR2_X1 npu_inst_pe_1_1_5_U22 ( .A1(npu_inst_pe_1_1_5_n56), .A2(
        npu_inst_pe_1_1_5_n3), .ZN(npu_inst_pe_1_1_5_n54) );
  NOR2_X1 npu_inst_pe_1_1_5_U21 ( .A1(npu_inst_pe_1_1_5_n52), .A2(
        npu_inst_pe_1_1_5_n3), .ZN(npu_inst_pe_1_1_5_n50) );
  NOR2_X1 npu_inst_pe_1_1_5_U20 ( .A1(npu_inst_pe_1_1_5_n48), .A2(
        npu_inst_pe_1_1_5_n3), .ZN(npu_inst_pe_1_1_5_n46) );
  NOR2_X1 npu_inst_pe_1_1_5_U19 ( .A1(npu_inst_pe_1_1_5_n40), .A2(
        npu_inst_pe_1_1_5_n3), .ZN(npu_inst_pe_1_1_5_n38) );
  NOR2_X1 npu_inst_pe_1_1_5_U18 ( .A1(npu_inst_pe_1_1_5_n44), .A2(
        npu_inst_pe_1_1_5_n3), .ZN(npu_inst_pe_1_1_5_n42) );
  BUF_X1 npu_inst_pe_1_1_5_U17 ( .A(npu_inst_n104), .Z(npu_inst_pe_1_1_5_n8)
         );
  INV_X1 npu_inst_pe_1_1_5_U16 ( .A(npu_inst_n126), .ZN(npu_inst_pe_1_1_5_n12)
         );
  INV_X1 npu_inst_pe_1_1_5_U15 ( .A(npu_inst_pe_1_1_5_n38), .ZN(
        npu_inst_pe_1_1_5_n114) );
  INV_X1 npu_inst_pe_1_1_5_U14 ( .A(npu_inst_pe_1_1_5_n58), .ZN(
        npu_inst_pe_1_1_5_n119) );
  INV_X1 npu_inst_pe_1_1_5_U13 ( .A(npu_inst_pe_1_1_5_n54), .ZN(
        npu_inst_pe_1_1_5_n118) );
  INV_X1 npu_inst_pe_1_1_5_U12 ( .A(npu_inst_pe_1_1_5_n50), .ZN(
        npu_inst_pe_1_1_5_n117) );
  INV_X1 npu_inst_pe_1_1_5_U11 ( .A(npu_inst_pe_1_1_5_n46), .ZN(
        npu_inst_pe_1_1_5_n116) );
  INV_X1 npu_inst_pe_1_1_5_U10 ( .A(npu_inst_pe_1_1_5_n42), .ZN(
        npu_inst_pe_1_1_5_n115) );
  BUF_X1 npu_inst_pe_1_1_5_U9 ( .A(npu_inst_n32), .Z(npu_inst_pe_1_1_5_n2) );
  BUF_X1 npu_inst_pe_1_1_5_U8 ( .A(npu_inst_n32), .Z(npu_inst_pe_1_1_5_n1) );
  BUF_X1 npu_inst_pe_1_1_5_U7 ( .A(npu_inst_pe_1_1_5_n12), .Z(
        npu_inst_pe_1_1_5_n11) );
  BUF_X1 npu_inst_pe_1_1_5_U6 ( .A(npu_inst_pe_1_1_5_n12), .Z(
        npu_inst_pe_1_1_5_n10) );
  BUF_X1 npu_inst_pe_1_1_5_U5 ( .A(npu_inst_pe_1_1_5_n12), .Z(
        npu_inst_pe_1_1_5_n9) );
  NOR2_X1 npu_inst_pe_1_1_5_U4 ( .A1(npu_inst_pe_1_1_5_int_q_weight_0_), .A2(
        npu_inst_pe_1_1_5_n1), .ZN(npu_inst_pe_1_1_5_n76) );
  NOR2_X1 npu_inst_pe_1_1_5_U3 ( .A1(npu_inst_pe_1_1_5_n27), .A2(
        npu_inst_pe_1_1_5_n1), .ZN(npu_inst_pe_1_1_5_n77) );
  FA_X1 npu_inst_pe_1_1_5_sub_67_U2_1 ( .A(npu_inst_pe_1_1_5_int_q_acc_1_), 
        .B(npu_inst_pe_1_1_5_n14), .CI(npu_inst_pe_1_1_5_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_1_5_sub_67_carry_2_), .S(npu_inst_pe_1_1_5_N66) );
  FA_X1 npu_inst_pe_1_1_5_add_69_U1_1 ( .A(npu_inst_pe_1_1_5_int_q_acc_1_), 
        .B(npu_inst_pe_1_1_5_int_data_1_), .CI(
        npu_inst_pe_1_1_5_add_69_carry_1_), .CO(
        npu_inst_pe_1_1_5_add_69_carry_2_), .S(npu_inst_pe_1_1_5_N74) );
  NAND3_X1 npu_inst_pe_1_1_5_U109 ( .A1(npu_inst_pe_1_1_5_n5), .A2(
        npu_inst_pe_1_1_5_n7), .A3(npu_inst_pe_1_1_5_n8), .ZN(
        npu_inst_pe_1_1_5_n44) );
  NAND3_X1 npu_inst_pe_1_1_5_U108 ( .A1(npu_inst_pe_1_1_5_n4), .A2(
        npu_inst_pe_1_1_5_n7), .A3(npu_inst_pe_1_1_5_n8), .ZN(
        npu_inst_pe_1_1_5_n40) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_1_5_n34), .CK(
        npu_inst_pe_1_1_5_net4263), .RN(npu_inst_pe_1_1_5_n9), .Q(
        npu_inst_pe_1_1_5_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_1_5_n35), .CK(
        npu_inst_pe_1_1_5_net4263), .RN(npu_inst_pe_1_1_5_n9), .Q(
        npu_inst_pe_1_1_5_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_1_5_n36), .CK(
        npu_inst_pe_1_1_5_net4263), .RN(npu_inst_pe_1_1_5_n9), .Q(
        npu_inst_pe_1_1_5_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_1_5_n98), .CK(
        npu_inst_pe_1_1_5_net4263), .RN(npu_inst_pe_1_1_5_n9), .Q(
        npu_inst_pe_1_1_5_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_1_5_n99), .CK(
        npu_inst_pe_1_1_5_net4263), .RN(npu_inst_pe_1_1_5_n9), .Q(
        npu_inst_pe_1_1_5_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_1_5_n100), 
        .CK(npu_inst_pe_1_1_5_net4263), .RN(npu_inst_pe_1_1_5_n9), .Q(
        npu_inst_pe_1_1_5_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_1_5_n33), .CK(
        npu_inst_pe_1_1_5_net4263), .RN(npu_inst_pe_1_1_5_n9), .Q(
        npu_inst_pe_1_1_5_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_1_5_n101), 
        .CK(npu_inst_pe_1_1_5_net4263), .RN(npu_inst_pe_1_1_5_n9), .Q(
        npu_inst_pe_1_1_5_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_weight_reg_0_ ( .D(npu_inst_n112), .CK(
        npu_inst_pe_1_1_5_net4269), .RN(npu_inst_pe_1_1_5_n9), .Q(
        npu_inst_pe_1_1_5_int_q_weight_0_), .QN(npu_inst_pe_1_1_5_n27) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_weight_reg_1_ ( .D(npu_inst_n118), .CK(
        npu_inst_pe_1_1_5_net4269), .RN(npu_inst_pe_1_1_5_n9), .Q(
        npu_inst_pe_1_1_5_int_q_weight_1_), .QN(npu_inst_pe_1_1_5_n26) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_1_5_n113), 
        .CK(npu_inst_pe_1_1_5_net4269), .RN(npu_inst_pe_1_1_5_n9), .Q(
        npu_inst_pe_1_1_5_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_1_5_n107), 
        .CK(npu_inst_pe_1_1_5_net4269), .RN(npu_inst_pe_1_1_5_n9), .Q(
        npu_inst_pe_1_1_5_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_1_5_n112), 
        .CK(npu_inst_pe_1_1_5_net4269), .RN(npu_inst_pe_1_1_5_n10), .Q(
        npu_inst_pe_1_1_5_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_1_5_n106), 
        .CK(npu_inst_pe_1_1_5_net4269), .RN(npu_inst_pe_1_1_5_n10), .Q(
        npu_inst_pe_1_1_5_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_1_5_n111), 
        .CK(npu_inst_pe_1_1_5_net4269), .RN(npu_inst_pe_1_1_5_n10), .Q(
        npu_inst_pe_1_1_5_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_1_5_n105), 
        .CK(npu_inst_pe_1_1_5_net4269), .RN(npu_inst_pe_1_1_5_n10), .Q(
        npu_inst_pe_1_1_5_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_1_5_n110), 
        .CK(npu_inst_pe_1_1_5_net4269), .RN(npu_inst_pe_1_1_5_n10), .Q(
        npu_inst_pe_1_1_5_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_1_5_n104), 
        .CK(npu_inst_pe_1_1_5_net4269), .RN(npu_inst_pe_1_1_5_n10), .Q(
        npu_inst_pe_1_1_5_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_1_5_n109), 
        .CK(npu_inst_pe_1_1_5_net4269), .RN(npu_inst_pe_1_1_5_n10), .Q(
        npu_inst_pe_1_1_5_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_1_5_n103), 
        .CK(npu_inst_pe_1_1_5_net4269), .RN(npu_inst_pe_1_1_5_n10), .Q(
        npu_inst_pe_1_1_5_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_1_5_n108), 
        .CK(npu_inst_pe_1_1_5_net4269), .RN(npu_inst_pe_1_1_5_n10), .Q(
        npu_inst_pe_1_1_5_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_1_5_n102), 
        .CK(npu_inst_pe_1_1_5_net4269), .RN(npu_inst_pe_1_1_5_n10), .Q(
        npu_inst_pe_1_1_5_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_1_5_n86), 
        .CK(npu_inst_pe_1_1_5_net4269), .RN(npu_inst_pe_1_1_5_n10), .Q(
        npu_inst_pe_1_1_5_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_1_5_n87), 
        .CK(npu_inst_pe_1_1_5_net4269), .RN(npu_inst_pe_1_1_5_n10), .Q(
        npu_inst_pe_1_1_5_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_1_5_n88), 
        .CK(npu_inst_pe_1_1_5_net4269), .RN(npu_inst_pe_1_1_5_n11), .Q(
        npu_inst_pe_1_1_5_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_1_5_n89), 
        .CK(npu_inst_pe_1_1_5_net4269), .RN(npu_inst_pe_1_1_5_n11), .Q(
        npu_inst_pe_1_1_5_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_1_5_n90), 
        .CK(npu_inst_pe_1_1_5_net4269), .RN(npu_inst_pe_1_1_5_n11), .Q(
        npu_inst_pe_1_1_5_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_1_5_n91), 
        .CK(npu_inst_pe_1_1_5_net4269), .RN(npu_inst_pe_1_1_5_n11), .Q(
        npu_inst_pe_1_1_5_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_1_5_n92), 
        .CK(npu_inst_pe_1_1_5_net4269), .RN(npu_inst_pe_1_1_5_n11), .Q(
        npu_inst_pe_1_1_5_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_1_5_n93), 
        .CK(npu_inst_pe_1_1_5_net4269), .RN(npu_inst_pe_1_1_5_n11), .Q(
        npu_inst_pe_1_1_5_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_1_5_n94), 
        .CK(npu_inst_pe_1_1_5_net4269), .RN(npu_inst_pe_1_1_5_n11), .Q(
        npu_inst_pe_1_1_5_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_1_5_n95), 
        .CK(npu_inst_pe_1_1_5_net4269), .RN(npu_inst_pe_1_1_5_n11), .Q(
        npu_inst_pe_1_1_5_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_1_5_n96), 
        .CK(npu_inst_pe_1_1_5_net4269), .RN(npu_inst_pe_1_1_5_n11), .Q(
        npu_inst_pe_1_1_5_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_1_5_n97), 
        .CK(npu_inst_pe_1_1_5_net4269), .RN(npu_inst_pe_1_1_5_n11), .Q(
        npu_inst_pe_1_1_5_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_1_5_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_1_5_N84), .SE(1'b0), .GCK(npu_inst_pe_1_1_5_net4263) );
  CLKGATETST_X1 npu_inst_pe_1_1_5_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n65), .SE(1'b0), .GCK(npu_inst_pe_1_1_5_net4269) );
  MUX2_X1 npu_inst_pe_1_1_6_U162 ( .A(npu_inst_pe_1_1_6_n32), .B(
        npu_inst_pe_1_1_6_n29), .S(npu_inst_pe_1_1_6_n8), .Z(
        npu_inst_pe_1_1_6_N93) );
  MUX2_X1 npu_inst_pe_1_1_6_U161 ( .A(npu_inst_pe_1_1_6_n31), .B(
        npu_inst_pe_1_1_6_n30), .S(npu_inst_pe_1_1_6_n6), .Z(
        npu_inst_pe_1_1_6_n32) );
  MUX2_X1 npu_inst_pe_1_1_6_U160 ( .A(npu_inst_pe_1_1_6_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_1_6_int_q_reg_v_1__0_), .S(npu_inst_pe_1_1_6_n4), .Z(
        npu_inst_pe_1_1_6_n31) );
  MUX2_X1 npu_inst_pe_1_1_6_U159 ( .A(npu_inst_pe_1_1_6_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_1_6_int_q_reg_v_3__0_), .S(npu_inst_pe_1_1_6_n4), .Z(
        npu_inst_pe_1_1_6_n30) );
  MUX2_X1 npu_inst_pe_1_1_6_U158 ( .A(npu_inst_pe_1_1_6_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_1_6_int_q_reg_v_5__0_), .S(npu_inst_pe_1_1_6_n4), .Z(
        npu_inst_pe_1_1_6_n29) );
  MUX2_X1 npu_inst_pe_1_1_6_U157 ( .A(npu_inst_pe_1_1_6_n28), .B(
        npu_inst_pe_1_1_6_n23), .S(npu_inst_pe_1_1_6_n8), .Z(
        npu_inst_pe_1_1_6_N94) );
  MUX2_X1 npu_inst_pe_1_1_6_U156 ( .A(npu_inst_pe_1_1_6_n25), .B(
        npu_inst_pe_1_1_6_n24), .S(npu_inst_pe_1_1_6_n6), .Z(
        npu_inst_pe_1_1_6_n28) );
  MUX2_X1 npu_inst_pe_1_1_6_U155 ( .A(npu_inst_pe_1_1_6_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_1_6_int_q_reg_v_1__1_), .S(npu_inst_pe_1_1_6_n4), .Z(
        npu_inst_pe_1_1_6_n25) );
  MUX2_X1 npu_inst_pe_1_1_6_U154 ( .A(npu_inst_pe_1_1_6_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_1_6_int_q_reg_v_3__1_), .S(npu_inst_pe_1_1_6_n4), .Z(
        npu_inst_pe_1_1_6_n24) );
  MUX2_X1 npu_inst_pe_1_1_6_U153 ( .A(npu_inst_pe_1_1_6_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_1_6_int_q_reg_v_5__1_), .S(npu_inst_pe_1_1_6_n4), .Z(
        npu_inst_pe_1_1_6_n23) );
  MUX2_X1 npu_inst_pe_1_1_6_U152 ( .A(npu_inst_pe_1_1_6_n22), .B(
        npu_inst_pe_1_1_6_n19), .S(npu_inst_pe_1_1_6_n8), .Z(
        npu_inst_int_data_x_1__6__1_) );
  MUX2_X1 npu_inst_pe_1_1_6_U151 ( .A(npu_inst_pe_1_1_6_n21), .B(
        npu_inst_pe_1_1_6_n20), .S(npu_inst_pe_1_1_6_n6), .Z(
        npu_inst_pe_1_1_6_n22) );
  MUX2_X1 npu_inst_pe_1_1_6_U150 ( .A(npu_inst_pe_1_1_6_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_1_6_int_q_reg_h_1__1_), .S(npu_inst_pe_1_1_6_n4), .Z(
        npu_inst_pe_1_1_6_n21) );
  MUX2_X1 npu_inst_pe_1_1_6_U149 ( .A(npu_inst_pe_1_1_6_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_1_6_int_q_reg_h_3__1_), .S(npu_inst_pe_1_1_6_n4), .Z(
        npu_inst_pe_1_1_6_n20) );
  MUX2_X1 npu_inst_pe_1_1_6_U148 ( .A(npu_inst_pe_1_1_6_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_1_6_int_q_reg_h_5__1_), .S(npu_inst_pe_1_1_6_n4), .Z(
        npu_inst_pe_1_1_6_n19) );
  MUX2_X1 npu_inst_pe_1_1_6_U147 ( .A(npu_inst_pe_1_1_6_n18), .B(
        npu_inst_pe_1_1_6_n15), .S(npu_inst_pe_1_1_6_n8), .Z(
        npu_inst_int_data_x_1__6__0_) );
  MUX2_X1 npu_inst_pe_1_1_6_U146 ( .A(npu_inst_pe_1_1_6_n17), .B(
        npu_inst_pe_1_1_6_n16), .S(npu_inst_pe_1_1_6_n6), .Z(
        npu_inst_pe_1_1_6_n18) );
  MUX2_X1 npu_inst_pe_1_1_6_U145 ( .A(npu_inst_pe_1_1_6_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_1_6_int_q_reg_h_1__0_), .S(npu_inst_pe_1_1_6_n4), .Z(
        npu_inst_pe_1_1_6_n17) );
  MUX2_X1 npu_inst_pe_1_1_6_U144 ( .A(npu_inst_pe_1_1_6_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_1_6_int_q_reg_h_3__0_), .S(npu_inst_pe_1_1_6_n4), .Z(
        npu_inst_pe_1_1_6_n16) );
  MUX2_X1 npu_inst_pe_1_1_6_U143 ( .A(npu_inst_pe_1_1_6_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_1_6_int_q_reg_h_5__0_), .S(npu_inst_pe_1_1_6_n4), .Z(
        npu_inst_pe_1_1_6_n15) );
  XOR2_X1 npu_inst_pe_1_1_6_U142 ( .A(npu_inst_pe_1_1_6_int_data_0_), .B(
        npu_inst_pe_1_1_6_int_q_acc_0_), .Z(npu_inst_pe_1_1_6_N73) );
  AND2_X1 npu_inst_pe_1_1_6_U141 ( .A1(npu_inst_pe_1_1_6_int_q_acc_0_), .A2(
        npu_inst_pe_1_1_6_int_data_0_), .ZN(npu_inst_pe_1_1_6_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_1_6_U140 ( .A(npu_inst_pe_1_1_6_int_q_acc_0_), .B(
        npu_inst_pe_1_1_6_n13), .ZN(npu_inst_pe_1_1_6_N65) );
  OR2_X1 npu_inst_pe_1_1_6_U139 ( .A1(npu_inst_pe_1_1_6_n13), .A2(
        npu_inst_pe_1_1_6_int_q_acc_0_), .ZN(npu_inst_pe_1_1_6_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_1_6_U138 ( .A(npu_inst_pe_1_1_6_int_q_acc_2_), .B(
        npu_inst_pe_1_1_6_add_69_carry_2_), .Z(npu_inst_pe_1_1_6_N75) );
  AND2_X1 npu_inst_pe_1_1_6_U137 ( .A1(npu_inst_pe_1_1_6_add_69_carry_2_), 
        .A2(npu_inst_pe_1_1_6_int_q_acc_2_), .ZN(
        npu_inst_pe_1_1_6_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_1_6_U136 ( .A(npu_inst_pe_1_1_6_int_q_acc_3_), .B(
        npu_inst_pe_1_1_6_add_69_carry_3_), .Z(npu_inst_pe_1_1_6_N76) );
  AND2_X1 npu_inst_pe_1_1_6_U135 ( .A1(npu_inst_pe_1_1_6_add_69_carry_3_), 
        .A2(npu_inst_pe_1_1_6_int_q_acc_3_), .ZN(
        npu_inst_pe_1_1_6_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_1_6_U134 ( .A(npu_inst_pe_1_1_6_int_q_acc_4_), .B(
        npu_inst_pe_1_1_6_add_69_carry_4_), .Z(npu_inst_pe_1_1_6_N77) );
  AND2_X1 npu_inst_pe_1_1_6_U133 ( .A1(npu_inst_pe_1_1_6_add_69_carry_4_), 
        .A2(npu_inst_pe_1_1_6_int_q_acc_4_), .ZN(
        npu_inst_pe_1_1_6_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_1_6_U132 ( .A(npu_inst_pe_1_1_6_int_q_acc_5_), .B(
        npu_inst_pe_1_1_6_add_69_carry_5_), .Z(npu_inst_pe_1_1_6_N78) );
  AND2_X1 npu_inst_pe_1_1_6_U131 ( .A1(npu_inst_pe_1_1_6_add_69_carry_5_), 
        .A2(npu_inst_pe_1_1_6_int_q_acc_5_), .ZN(
        npu_inst_pe_1_1_6_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_1_6_U130 ( .A(npu_inst_pe_1_1_6_int_q_acc_6_), .B(
        npu_inst_pe_1_1_6_add_69_carry_6_), .Z(npu_inst_pe_1_1_6_N79) );
  AND2_X1 npu_inst_pe_1_1_6_U129 ( .A1(npu_inst_pe_1_1_6_add_69_carry_6_), 
        .A2(npu_inst_pe_1_1_6_int_q_acc_6_), .ZN(
        npu_inst_pe_1_1_6_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_1_6_U128 ( .A(npu_inst_pe_1_1_6_int_q_acc_7_), .B(
        npu_inst_pe_1_1_6_add_69_carry_7_), .Z(npu_inst_pe_1_1_6_N80) );
  XNOR2_X1 npu_inst_pe_1_1_6_U127 ( .A(npu_inst_pe_1_1_6_sub_67_carry_2_), .B(
        npu_inst_pe_1_1_6_int_q_acc_2_), .ZN(npu_inst_pe_1_1_6_N67) );
  OR2_X1 npu_inst_pe_1_1_6_U126 ( .A1(npu_inst_pe_1_1_6_int_q_acc_2_), .A2(
        npu_inst_pe_1_1_6_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_1_6_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_1_6_U125 ( .A(npu_inst_pe_1_1_6_sub_67_carry_3_), .B(
        npu_inst_pe_1_1_6_int_q_acc_3_), .ZN(npu_inst_pe_1_1_6_N68) );
  OR2_X1 npu_inst_pe_1_1_6_U124 ( .A1(npu_inst_pe_1_1_6_int_q_acc_3_), .A2(
        npu_inst_pe_1_1_6_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_1_6_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_1_6_U123 ( .A(npu_inst_pe_1_1_6_sub_67_carry_4_), .B(
        npu_inst_pe_1_1_6_int_q_acc_4_), .ZN(npu_inst_pe_1_1_6_N69) );
  OR2_X1 npu_inst_pe_1_1_6_U122 ( .A1(npu_inst_pe_1_1_6_int_q_acc_4_), .A2(
        npu_inst_pe_1_1_6_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_1_6_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_1_6_U121 ( .A(npu_inst_pe_1_1_6_sub_67_carry_5_), .B(
        npu_inst_pe_1_1_6_int_q_acc_5_), .ZN(npu_inst_pe_1_1_6_N70) );
  OR2_X1 npu_inst_pe_1_1_6_U120 ( .A1(npu_inst_pe_1_1_6_int_q_acc_5_), .A2(
        npu_inst_pe_1_1_6_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_1_6_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_1_6_U119 ( .A(npu_inst_pe_1_1_6_sub_67_carry_6_), .B(
        npu_inst_pe_1_1_6_int_q_acc_6_), .ZN(npu_inst_pe_1_1_6_N71) );
  OR2_X1 npu_inst_pe_1_1_6_U118 ( .A1(npu_inst_pe_1_1_6_int_q_acc_6_), .A2(
        npu_inst_pe_1_1_6_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_1_6_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_1_6_U117 ( .A(npu_inst_pe_1_1_6_int_q_acc_7_), .B(
        npu_inst_pe_1_1_6_sub_67_carry_7_), .ZN(npu_inst_pe_1_1_6_N72) );
  INV_X1 npu_inst_pe_1_1_6_U116 ( .A(npu_inst_n79), .ZN(npu_inst_pe_1_1_6_n7)
         );
  INV_X1 npu_inst_pe_1_1_6_U115 ( .A(npu_inst_pe_1_1_6_n7), .ZN(
        npu_inst_pe_1_1_6_n6) );
  INV_X1 npu_inst_pe_1_1_6_U114 ( .A(npu_inst_n59), .ZN(npu_inst_pe_1_1_6_n3)
         );
  AOI22_X1 npu_inst_pe_1_1_6_U113 ( .A1(npu_inst_int_data_y_2__6__0_), .A2(
        npu_inst_pe_1_1_6_n58), .B1(npu_inst_pe_1_1_6_n119), .B2(
        npu_inst_pe_1_1_6_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_1_6_n57) );
  INV_X1 npu_inst_pe_1_1_6_U112 ( .A(npu_inst_pe_1_1_6_n57), .ZN(
        npu_inst_pe_1_1_6_n108) );
  AOI22_X1 npu_inst_pe_1_1_6_U111 ( .A1(npu_inst_int_data_y_2__6__0_), .A2(
        npu_inst_pe_1_1_6_n54), .B1(npu_inst_pe_1_1_6_n118), .B2(
        npu_inst_pe_1_1_6_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_1_6_n53) );
  INV_X1 npu_inst_pe_1_1_6_U110 ( .A(npu_inst_pe_1_1_6_n53), .ZN(
        npu_inst_pe_1_1_6_n109) );
  AOI22_X1 npu_inst_pe_1_1_6_U107 ( .A1(npu_inst_int_data_y_2__6__0_), .A2(
        npu_inst_pe_1_1_6_n50), .B1(npu_inst_pe_1_1_6_n117), .B2(
        npu_inst_pe_1_1_6_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_1_6_n49) );
  INV_X1 npu_inst_pe_1_1_6_U106 ( .A(npu_inst_pe_1_1_6_n49), .ZN(
        npu_inst_pe_1_1_6_n110) );
  AOI22_X1 npu_inst_pe_1_1_6_U105 ( .A1(npu_inst_int_data_y_2__6__0_), .A2(
        npu_inst_pe_1_1_6_n46), .B1(npu_inst_pe_1_1_6_n116), .B2(
        npu_inst_pe_1_1_6_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_1_6_n45) );
  INV_X1 npu_inst_pe_1_1_6_U104 ( .A(npu_inst_pe_1_1_6_n45), .ZN(
        npu_inst_pe_1_1_6_n111) );
  AOI22_X1 npu_inst_pe_1_1_6_U103 ( .A1(npu_inst_int_data_y_2__6__0_), .A2(
        npu_inst_pe_1_1_6_n42), .B1(npu_inst_pe_1_1_6_n115), .B2(
        npu_inst_pe_1_1_6_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_1_6_n41) );
  INV_X1 npu_inst_pe_1_1_6_U102 ( .A(npu_inst_pe_1_1_6_n41), .ZN(
        npu_inst_pe_1_1_6_n112) );
  AOI22_X1 npu_inst_pe_1_1_6_U101 ( .A1(npu_inst_int_data_y_2__6__1_), .A2(
        npu_inst_pe_1_1_6_n58), .B1(npu_inst_pe_1_1_6_n119), .B2(
        npu_inst_pe_1_1_6_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_1_6_n59) );
  INV_X1 npu_inst_pe_1_1_6_U100 ( .A(npu_inst_pe_1_1_6_n59), .ZN(
        npu_inst_pe_1_1_6_n102) );
  AOI22_X1 npu_inst_pe_1_1_6_U99 ( .A1(npu_inst_int_data_y_2__6__1_), .A2(
        npu_inst_pe_1_1_6_n54), .B1(npu_inst_pe_1_1_6_n118), .B2(
        npu_inst_pe_1_1_6_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_1_6_n55) );
  INV_X1 npu_inst_pe_1_1_6_U98 ( .A(npu_inst_pe_1_1_6_n55), .ZN(
        npu_inst_pe_1_1_6_n103) );
  AOI22_X1 npu_inst_pe_1_1_6_U97 ( .A1(npu_inst_int_data_y_2__6__1_), .A2(
        npu_inst_pe_1_1_6_n50), .B1(npu_inst_pe_1_1_6_n117), .B2(
        npu_inst_pe_1_1_6_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_1_6_n51) );
  INV_X1 npu_inst_pe_1_1_6_U96 ( .A(npu_inst_pe_1_1_6_n51), .ZN(
        npu_inst_pe_1_1_6_n104) );
  AOI22_X1 npu_inst_pe_1_1_6_U95 ( .A1(npu_inst_int_data_y_2__6__1_), .A2(
        npu_inst_pe_1_1_6_n46), .B1(npu_inst_pe_1_1_6_n116), .B2(
        npu_inst_pe_1_1_6_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_1_6_n47) );
  INV_X1 npu_inst_pe_1_1_6_U94 ( .A(npu_inst_pe_1_1_6_n47), .ZN(
        npu_inst_pe_1_1_6_n105) );
  AOI22_X1 npu_inst_pe_1_1_6_U93 ( .A1(npu_inst_int_data_y_2__6__1_), .A2(
        npu_inst_pe_1_1_6_n42), .B1(npu_inst_pe_1_1_6_n115), .B2(
        npu_inst_pe_1_1_6_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_1_6_n43) );
  INV_X1 npu_inst_pe_1_1_6_U92 ( .A(npu_inst_pe_1_1_6_n43), .ZN(
        npu_inst_pe_1_1_6_n106) );
  AOI22_X1 npu_inst_pe_1_1_6_U91 ( .A1(npu_inst_pe_1_1_6_n38), .A2(
        npu_inst_int_data_y_2__6__1_), .B1(npu_inst_pe_1_1_6_n114), .B2(
        npu_inst_pe_1_1_6_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_1_6_n39) );
  INV_X1 npu_inst_pe_1_1_6_U90 ( .A(npu_inst_pe_1_1_6_n39), .ZN(
        npu_inst_pe_1_1_6_n107) );
  AOI22_X1 npu_inst_pe_1_1_6_U89 ( .A1(npu_inst_pe_1_1_6_n38), .A2(
        npu_inst_int_data_y_2__6__0_), .B1(npu_inst_pe_1_1_6_n114), .B2(
        npu_inst_pe_1_1_6_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_1_6_n37) );
  INV_X1 npu_inst_pe_1_1_6_U88 ( .A(npu_inst_pe_1_1_6_n37), .ZN(
        npu_inst_pe_1_1_6_n113) );
  NAND2_X1 npu_inst_pe_1_1_6_U87 ( .A1(npu_inst_pe_1_1_6_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_1_6_n60), .ZN(npu_inst_pe_1_1_6_n74) );
  OAI21_X1 npu_inst_pe_1_1_6_U86 ( .B1(npu_inst_pe_1_1_6_n63), .B2(
        npu_inst_pe_1_1_6_n60), .A(npu_inst_pe_1_1_6_n74), .ZN(
        npu_inst_pe_1_1_6_n97) );
  NAND2_X1 npu_inst_pe_1_1_6_U85 ( .A1(npu_inst_pe_1_1_6_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_1_6_n60), .ZN(npu_inst_pe_1_1_6_n73) );
  OAI21_X1 npu_inst_pe_1_1_6_U84 ( .B1(npu_inst_pe_1_1_6_n61), .B2(
        npu_inst_pe_1_1_6_n60), .A(npu_inst_pe_1_1_6_n73), .ZN(
        npu_inst_pe_1_1_6_n96) );
  NAND2_X1 npu_inst_pe_1_1_6_U83 ( .A1(npu_inst_pe_1_1_6_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_1_6_n56), .ZN(npu_inst_pe_1_1_6_n72) );
  OAI21_X1 npu_inst_pe_1_1_6_U82 ( .B1(npu_inst_pe_1_1_6_n63), .B2(
        npu_inst_pe_1_1_6_n56), .A(npu_inst_pe_1_1_6_n72), .ZN(
        npu_inst_pe_1_1_6_n95) );
  NAND2_X1 npu_inst_pe_1_1_6_U81 ( .A1(npu_inst_pe_1_1_6_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_1_6_n56), .ZN(npu_inst_pe_1_1_6_n71) );
  OAI21_X1 npu_inst_pe_1_1_6_U80 ( .B1(npu_inst_pe_1_1_6_n61), .B2(
        npu_inst_pe_1_1_6_n56), .A(npu_inst_pe_1_1_6_n71), .ZN(
        npu_inst_pe_1_1_6_n94) );
  NAND2_X1 npu_inst_pe_1_1_6_U79 ( .A1(npu_inst_pe_1_1_6_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_1_6_n52), .ZN(npu_inst_pe_1_1_6_n70) );
  OAI21_X1 npu_inst_pe_1_1_6_U78 ( .B1(npu_inst_pe_1_1_6_n63), .B2(
        npu_inst_pe_1_1_6_n52), .A(npu_inst_pe_1_1_6_n70), .ZN(
        npu_inst_pe_1_1_6_n93) );
  NAND2_X1 npu_inst_pe_1_1_6_U77 ( .A1(npu_inst_pe_1_1_6_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_1_6_n52), .ZN(npu_inst_pe_1_1_6_n69) );
  OAI21_X1 npu_inst_pe_1_1_6_U76 ( .B1(npu_inst_pe_1_1_6_n61), .B2(
        npu_inst_pe_1_1_6_n52), .A(npu_inst_pe_1_1_6_n69), .ZN(
        npu_inst_pe_1_1_6_n92) );
  NAND2_X1 npu_inst_pe_1_1_6_U75 ( .A1(npu_inst_pe_1_1_6_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_1_6_n48), .ZN(npu_inst_pe_1_1_6_n68) );
  OAI21_X1 npu_inst_pe_1_1_6_U74 ( .B1(npu_inst_pe_1_1_6_n63), .B2(
        npu_inst_pe_1_1_6_n48), .A(npu_inst_pe_1_1_6_n68), .ZN(
        npu_inst_pe_1_1_6_n91) );
  NAND2_X1 npu_inst_pe_1_1_6_U73 ( .A1(npu_inst_pe_1_1_6_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_1_6_n48), .ZN(npu_inst_pe_1_1_6_n67) );
  OAI21_X1 npu_inst_pe_1_1_6_U72 ( .B1(npu_inst_pe_1_1_6_n61), .B2(
        npu_inst_pe_1_1_6_n48), .A(npu_inst_pe_1_1_6_n67), .ZN(
        npu_inst_pe_1_1_6_n90) );
  NAND2_X1 npu_inst_pe_1_1_6_U71 ( .A1(npu_inst_pe_1_1_6_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_1_6_n44), .ZN(npu_inst_pe_1_1_6_n66) );
  OAI21_X1 npu_inst_pe_1_1_6_U70 ( .B1(npu_inst_pe_1_1_6_n63), .B2(
        npu_inst_pe_1_1_6_n44), .A(npu_inst_pe_1_1_6_n66), .ZN(
        npu_inst_pe_1_1_6_n89) );
  NAND2_X1 npu_inst_pe_1_1_6_U69 ( .A1(npu_inst_pe_1_1_6_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_1_6_n44), .ZN(npu_inst_pe_1_1_6_n65) );
  OAI21_X1 npu_inst_pe_1_1_6_U68 ( .B1(npu_inst_pe_1_1_6_n61), .B2(
        npu_inst_pe_1_1_6_n44), .A(npu_inst_pe_1_1_6_n65), .ZN(
        npu_inst_pe_1_1_6_n88) );
  NAND2_X1 npu_inst_pe_1_1_6_U67 ( .A1(npu_inst_pe_1_1_6_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_1_6_n40), .ZN(npu_inst_pe_1_1_6_n64) );
  OAI21_X1 npu_inst_pe_1_1_6_U66 ( .B1(npu_inst_pe_1_1_6_n63), .B2(
        npu_inst_pe_1_1_6_n40), .A(npu_inst_pe_1_1_6_n64), .ZN(
        npu_inst_pe_1_1_6_n87) );
  NAND2_X1 npu_inst_pe_1_1_6_U65 ( .A1(npu_inst_pe_1_1_6_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_1_6_n40), .ZN(npu_inst_pe_1_1_6_n62) );
  OAI21_X1 npu_inst_pe_1_1_6_U64 ( .B1(npu_inst_pe_1_1_6_n61), .B2(
        npu_inst_pe_1_1_6_n40), .A(npu_inst_pe_1_1_6_n62), .ZN(
        npu_inst_pe_1_1_6_n86) );
  AND2_X1 npu_inst_pe_1_1_6_U63 ( .A1(npu_inst_pe_1_1_6_N93), .A2(npu_inst_n59), .ZN(npu_inst_int_data_y_1__6__0_) );
  AND2_X1 npu_inst_pe_1_1_6_U62 ( .A1(npu_inst_n59), .A2(npu_inst_pe_1_1_6_N94), .ZN(npu_inst_int_data_y_1__6__1_) );
  NOR3_X1 npu_inst_pe_1_1_6_U61 ( .A1(npu_inst_pe_1_1_6_n26), .A2(npu_inst_n59), .A3(npu_inst_int_ckg[49]), .ZN(npu_inst_pe_1_1_6_n85) );
  OR2_X1 npu_inst_pe_1_1_6_U60 ( .A1(npu_inst_pe_1_1_6_n85), .A2(
        npu_inst_pe_1_1_6_n2), .ZN(npu_inst_pe_1_1_6_N84) );
  AND2_X1 npu_inst_pe_1_1_6_U59 ( .A1(npu_inst_pe_1_1_6_int_q_acc_0_), .A2(
        npu_inst_pe_1_1_6_n1), .ZN(npu_inst_int_data_res_1__6__0_) );
  AND2_X1 npu_inst_pe_1_1_6_U58 ( .A1(npu_inst_pe_1_1_6_n2), .A2(
        npu_inst_pe_1_1_6_int_q_acc_7_), .ZN(npu_inst_int_data_res_1__6__7_)
         );
  AND2_X1 npu_inst_pe_1_1_6_U57 ( .A1(npu_inst_pe_1_1_6_int_q_acc_1_), .A2(
        npu_inst_pe_1_1_6_n1), .ZN(npu_inst_int_data_res_1__6__1_) );
  AND2_X1 npu_inst_pe_1_1_6_U56 ( .A1(npu_inst_pe_1_1_6_int_q_acc_2_), .A2(
        npu_inst_pe_1_1_6_n1), .ZN(npu_inst_int_data_res_1__6__2_) );
  AND2_X1 npu_inst_pe_1_1_6_U55 ( .A1(npu_inst_pe_1_1_6_int_q_acc_3_), .A2(
        npu_inst_pe_1_1_6_n2), .ZN(npu_inst_int_data_res_1__6__3_) );
  AND2_X1 npu_inst_pe_1_1_6_U54 ( .A1(npu_inst_pe_1_1_6_int_q_acc_4_), .A2(
        npu_inst_pe_1_1_6_n2), .ZN(npu_inst_int_data_res_1__6__4_) );
  AND2_X1 npu_inst_pe_1_1_6_U53 ( .A1(npu_inst_pe_1_1_6_int_q_acc_5_), .A2(
        npu_inst_pe_1_1_6_n2), .ZN(npu_inst_int_data_res_1__6__5_) );
  AND2_X1 npu_inst_pe_1_1_6_U52 ( .A1(npu_inst_pe_1_1_6_int_q_acc_6_), .A2(
        npu_inst_pe_1_1_6_n2), .ZN(npu_inst_int_data_res_1__6__6_) );
  AOI222_X1 npu_inst_pe_1_1_6_U51 ( .A1(npu_inst_int_data_res_2__6__0_), .A2(
        npu_inst_pe_1_1_6_n1), .B1(npu_inst_pe_1_1_6_N73), .B2(
        npu_inst_pe_1_1_6_n76), .C1(npu_inst_pe_1_1_6_N65), .C2(
        npu_inst_pe_1_1_6_n77), .ZN(npu_inst_pe_1_1_6_n84) );
  INV_X1 npu_inst_pe_1_1_6_U50 ( .A(npu_inst_pe_1_1_6_n84), .ZN(
        npu_inst_pe_1_1_6_n101) );
  AOI222_X1 npu_inst_pe_1_1_6_U49 ( .A1(npu_inst_int_data_res_2__6__7_), .A2(
        npu_inst_pe_1_1_6_n1), .B1(npu_inst_pe_1_1_6_N80), .B2(
        npu_inst_pe_1_1_6_n76), .C1(npu_inst_pe_1_1_6_N72), .C2(
        npu_inst_pe_1_1_6_n77), .ZN(npu_inst_pe_1_1_6_n75) );
  INV_X1 npu_inst_pe_1_1_6_U48 ( .A(npu_inst_pe_1_1_6_n75), .ZN(
        npu_inst_pe_1_1_6_n33) );
  AOI222_X1 npu_inst_pe_1_1_6_U47 ( .A1(npu_inst_int_data_res_2__6__1_), .A2(
        npu_inst_pe_1_1_6_n1), .B1(npu_inst_pe_1_1_6_N74), .B2(
        npu_inst_pe_1_1_6_n76), .C1(npu_inst_pe_1_1_6_N66), .C2(
        npu_inst_pe_1_1_6_n77), .ZN(npu_inst_pe_1_1_6_n83) );
  INV_X1 npu_inst_pe_1_1_6_U46 ( .A(npu_inst_pe_1_1_6_n83), .ZN(
        npu_inst_pe_1_1_6_n100) );
  AOI222_X1 npu_inst_pe_1_1_6_U45 ( .A1(npu_inst_int_data_res_2__6__2_), .A2(
        npu_inst_pe_1_1_6_n1), .B1(npu_inst_pe_1_1_6_N75), .B2(
        npu_inst_pe_1_1_6_n76), .C1(npu_inst_pe_1_1_6_N67), .C2(
        npu_inst_pe_1_1_6_n77), .ZN(npu_inst_pe_1_1_6_n82) );
  INV_X1 npu_inst_pe_1_1_6_U44 ( .A(npu_inst_pe_1_1_6_n82), .ZN(
        npu_inst_pe_1_1_6_n99) );
  AOI222_X1 npu_inst_pe_1_1_6_U43 ( .A1(npu_inst_int_data_res_2__6__3_), .A2(
        npu_inst_pe_1_1_6_n1), .B1(npu_inst_pe_1_1_6_N76), .B2(
        npu_inst_pe_1_1_6_n76), .C1(npu_inst_pe_1_1_6_N68), .C2(
        npu_inst_pe_1_1_6_n77), .ZN(npu_inst_pe_1_1_6_n81) );
  INV_X1 npu_inst_pe_1_1_6_U42 ( .A(npu_inst_pe_1_1_6_n81), .ZN(
        npu_inst_pe_1_1_6_n98) );
  AOI222_X1 npu_inst_pe_1_1_6_U41 ( .A1(npu_inst_int_data_res_2__6__4_), .A2(
        npu_inst_pe_1_1_6_n1), .B1(npu_inst_pe_1_1_6_N77), .B2(
        npu_inst_pe_1_1_6_n76), .C1(npu_inst_pe_1_1_6_N69), .C2(
        npu_inst_pe_1_1_6_n77), .ZN(npu_inst_pe_1_1_6_n80) );
  INV_X1 npu_inst_pe_1_1_6_U40 ( .A(npu_inst_pe_1_1_6_n80), .ZN(
        npu_inst_pe_1_1_6_n36) );
  AOI222_X1 npu_inst_pe_1_1_6_U39 ( .A1(npu_inst_int_data_res_2__6__5_), .A2(
        npu_inst_pe_1_1_6_n1), .B1(npu_inst_pe_1_1_6_N78), .B2(
        npu_inst_pe_1_1_6_n76), .C1(npu_inst_pe_1_1_6_N70), .C2(
        npu_inst_pe_1_1_6_n77), .ZN(npu_inst_pe_1_1_6_n79) );
  INV_X1 npu_inst_pe_1_1_6_U38 ( .A(npu_inst_pe_1_1_6_n79), .ZN(
        npu_inst_pe_1_1_6_n35) );
  AOI222_X1 npu_inst_pe_1_1_6_U37 ( .A1(npu_inst_int_data_res_2__6__6_), .A2(
        npu_inst_pe_1_1_6_n1), .B1(npu_inst_pe_1_1_6_N79), .B2(
        npu_inst_pe_1_1_6_n76), .C1(npu_inst_pe_1_1_6_N71), .C2(
        npu_inst_pe_1_1_6_n77), .ZN(npu_inst_pe_1_1_6_n78) );
  INV_X1 npu_inst_pe_1_1_6_U36 ( .A(npu_inst_pe_1_1_6_n78), .ZN(
        npu_inst_pe_1_1_6_n34) );
  INV_X1 npu_inst_pe_1_1_6_U35 ( .A(npu_inst_pe_1_1_6_int_data_1_), .ZN(
        npu_inst_pe_1_1_6_n14) );
  AND2_X1 npu_inst_pe_1_1_6_U34 ( .A1(npu_inst_int_data_x_1__6__1_), .A2(
        npu_inst_pe_1_1_6_int_q_weight_1_), .ZN(npu_inst_pe_1_1_6_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_1_6_U33 ( .A1(npu_inst_int_data_x_1__6__0_), .A2(
        npu_inst_pe_1_1_6_int_q_weight_1_), .ZN(npu_inst_pe_1_1_6_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_1_6_U32 ( .A1(npu_inst_n59), .A2(
        npu_inst_int_data_y_2__6__1_), .B1(npu_inst_pe_1_1_6_n3), .B2(
        npu_inst_int_data_x_1__7__1_), .ZN(npu_inst_pe_1_1_6_n63) );
  AOI22_X1 npu_inst_pe_1_1_6_U31 ( .A1(npu_inst_n59), .A2(
        npu_inst_int_data_y_2__6__0_), .B1(npu_inst_pe_1_1_6_n3), .B2(
        npu_inst_int_data_x_1__7__0_), .ZN(npu_inst_pe_1_1_6_n61) );
  INV_X1 npu_inst_pe_1_1_6_U30 ( .A(npu_inst_pe_1_1_6_int_data_0_), .ZN(
        npu_inst_pe_1_1_6_n13) );
  INV_X1 npu_inst_pe_1_1_6_U29 ( .A(npu_inst_n71), .ZN(npu_inst_pe_1_1_6_n5)
         );
  OR3_X1 npu_inst_pe_1_1_6_U28 ( .A1(npu_inst_pe_1_1_6_n6), .A2(
        npu_inst_pe_1_1_6_n8), .A3(npu_inst_pe_1_1_6_n5), .ZN(
        npu_inst_pe_1_1_6_n56) );
  OR3_X1 npu_inst_pe_1_1_6_U27 ( .A1(npu_inst_pe_1_1_6_n5), .A2(
        npu_inst_pe_1_1_6_n8), .A3(npu_inst_pe_1_1_6_n7), .ZN(
        npu_inst_pe_1_1_6_n48) );
  INV_X1 npu_inst_pe_1_1_6_U26 ( .A(npu_inst_pe_1_1_6_n5), .ZN(
        npu_inst_pe_1_1_6_n4) );
  OR3_X1 npu_inst_pe_1_1_6_U25 ( .A1(npu_inst_pe_1_1_6_n4), .A2(
        npu_inst_pe_1_1_6_n8), .A3(npu_inst_pe_1_1_6_n7), .ZN(
        npu_inst_pe_1_1_6_n52) );
  OR3_X1 npu_inst_pe_1_1_6_U24 ( .A1(npu_inst_pe_1_1_6_n6), .A2(
        npu_inst_pe_1_1_6_n8), .A3(npu_inst_pe_1_1_6_n4), .ZN(
        npu_inst_pe_1_1_6_n60) );
  NOR2_X1 npu_inst_pe_1_1_6_U23 ( .A1(npu_inst_pe_1_1_6_n60), .A2(
        npu_inst_pe_1_1_6_n3), .ZN(npu_inst_pe_1_1_6_n58) );
  NOR2_X1 npu_inst_pe_1_1_6_U22 ( .A1(npu_inst_pe_1_1_6_n56), .A2(
        npu_inst_pe_1_1_6_n3), .ZN(npu_inst_pe_1_1_6_n54) );
  NOR2_X1 npu_inst_pe_1_1_6_U21 ( .A1(npu_inst_pe_1_1_6_n52), .A2(
        npu_inst_pe_1_1_6_n3), .ZN(npu_inst_pe_1_1_6_n50) );
  NOR2_X1 npu_inst_pe_1_1_6_U20 ( .A1(npu_inst_pe_1_1_6_n48), .A2(
        npu_inst_pe_1_1_6_n3), .ZN(npu_inst_pe_1_1_6_n46) );
  NOR2_X1 npu_inst_pe_1_1_6_U19 ( .A1(npu_inst_pe_1_1_6_n40), .A2(
        npu_inst_pe_1_1_6_n3), .ZN(npu_inst_pe_1_1_6_n38) );
  NOR2_X1 npu_inst_pe_1_1_6_U18 ( .A1(npu_inst_pe_1_1_6_n44), .A2(
        npu_inst_pe_1_1_6_n3), .ZN(npu_inst_pe_1_1_6_n42) );
  BUF_X1 npu_inst_pe_1_1_6_U17 ( .A(npu_inst_n104), .Z(npu_inst_pe_1_1_6_n8)
         );
  INV_X1 npu_inst_pe_1_1_6_U16 ( .A(npu_inst_n126), .ZN(npu_inst_pe_1_1_6_n12)
         );
  INV_X1 npu_inst_pe_1_1_6_U15 ( .A(npu_inst_pe_1_1_6_n38), .ZN(
        npu_inst_pe_1_1_6_n114) );
  INV_X1 npu_inst_pe_1_1_6_U14 ( .A(npu_inst_pe_1_1_6_n58), .ZN(
        npu_inst_pe_1_1_6_n119) );
  INV_X1 npu_inst_pe_1_1_6_U13 ( .A(npu_inst_pe_1_1_6_n54), .ZN(
        npu_inst_pe_1_1_6_n118) );
  INV_X1 npu_inst_pe_1_1_6_U12 ( .A(npu_inst_pe_1_1_6_n50), .ZN(
        npu_inst_pe_1_1_6_n117) );
  INV_X1 npu_inst_pe_1_1_6_U11 ( .A(npu_inst_pe_1_1_6_n46), .ZN(
        npu_inst_pe_1_1_6_n116) );
  INV_X1 npu_inst_pe_1_1_6_U10 ( .A(npu_inst_pe_1_1_6_n42), .ZN(
        npu_inst_pe_1_1_6_n115) );
  BUF_X1 npu_inst_pe_1_1_6_U9 ( .A(npu_inst_n31), .Z(npu_inst_pe_1_1_6_n2) );
  BUF_X1 npu_inst_pe_1_1_6_U8 ( .A(npu_inst_n31), .Z(npu_inst_pe_1_1_6_n1) );
  BUF_X1 npu_inst_pe_1_1_6_U7 ( .A(npu_inst_pe_1_1_6_n12), .Z(
        npu_inst_pe_1_1_6_n11) );
  BUF_X1 npu_inst_pe_1_1_6_U6 ( .A(npu_inst_pe_1_1_6_n12), .Z(
        npu_inst_pe_1_1_6_n10) );
  BUF_X1 npu_inst_pe_1_1_6_U5 ( .A(npu_inst_pe_1_1_6_n12), .Z(
        npu_inst_pe_1_1_6_n9) );
  NOR2_X1 npu_inst_pe_1_1_6_U4 ( .A1(npu_inst_pe_1_1_6_int_q_weight_0_), .A2(
        npu_inst_pe_1_1_6_n1), .ZN(npu_inst_pe_1_1_6_n76) );
  NOR2_X1 npu_inst_pe_1_1_6_U3 ( .A1(npu_inst_pe_1_1_6_n27), .A2(
        npu_inst_pe_1_1_6_n1), .ZN(npu_inst_pe_1_1_6_n77) );
  FA_X1 npu_inst_pe_1_1_6_sub_67_U2_1 ( .A(npu_inst_pe_1_1_6_int_q_acc_1_), 
        .B(npu_inst_pe_1_1_6_n14), .CI(npu_inst_pe_1_1_6_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_1_6_sub_67_carry_2_), .S(npu_inst_pe_1_1_6_N66) );
  FA_X1 npu_inst_pe_1_1_6_add_69_U1_1 ( .A(npu_inst_pe_1_1_6_int_q_acc_1_), 
        .B(npu_inst_pe_1_1_6_int_data_1_), .CI(
        npu_inst_pe_1_1_6_add_69_carry_1_), .CO(
        npu_inst_pe_1_1_6_add_69_carry_2_), .S(npu_inst_pe_1_1_6_N74) );
  NAND3_X1 npu_inst_pe_1_1_6_U109 ( .A1(npu_inst_pe_1_1_6_n5), .A2(
        npu_inst_pe_1_1_6_n7), .A3(npu_inst_pe_1_1_6_n8), .ZN(
        npu_inst_pe_1_1_6_n44) );
  NAND3_X1 npu_inst_pe_1_1_6_U108 ( .A1(npu_inst_pe_1_1_6_n4), .A2(
        npu_inst_pe_1_1_6_n7), .A3(npu_inst_pe_1_1_6_n8), .ZN(
        npu_inst_pe_1_1_6_n40) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_1_6_n34), .CK(
        npu_inst_pe_1_1_6_net4240), .RN(npu_inst_pe_1_1_6_n9), .Q(
        npu_inst_pe_1_1_6_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_1_6_n35), .CK(
        npu_inst_pe_1_1_6_net4240), .RN(npu_inst_pe_1_1_6_n9), .Q(
        npu_inst_pe_1_1_6_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_1_6_n36), .CK(
        npu_inst_pe_1_1_6_net4240), .RN(npu_inst_pe_1_1_6_n9), .Q(
        npu_inst_pe_1_1_6_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_1_6_n98), .CK(
        npu_inst_pe_1_1_6_net4240), .RN(npu_inst_pe_1_1_6_n9), .Q(
        npu_inst_pe_1_1_6_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_1_6_n99), .CK(
        npu_inst_pe_1_1_6_net4240), .RN(npu_inst_pe_1_1_6_n9), .Q(
        npu_inst_pe_1_1_6_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_1_6_n100), 
        .CK(npu_inst_pe_1_1_6_net4240), .RN(npu_inst_pe_1_1_6_n9), .Q(
        npu_inst_pe_1_1_6_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_1_6_n33), .CK(
        npu_inst_pe_1_1_6_net4240), .RN(npu_inst_pe_1_1_6_n9), .Q(
        npu_inst_pe_1_1_6_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_1_6_n101), 
        .CK(npu_inst_pe_1_1_6_net4240), .RN(npu_inst_pe_1_1_6_n9), .Q(
        npu_inst_pe_1_1_6_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_weight_reg_0_ ( .D(npu_inst_n112), .CK(
        npu_inst_pe_1_1_6_net4246), .RN(npu_inst_pe_1_1_6_n9), .Q(
        npu_inst_pe_1_1_6_int_q_weight_0_), .QN(npu_inst_pe_1_1_6_n27) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_weight_reg_1_ ( .D(npu_inst_n118), .CK(
        npu_inst_pe_1_1_6_net4246), .RN(npu_inst_pe_1_1_6_n9), .Q(
        npu_inst_pe_1_1_6_int_q_weight_1_), .QN(npu_inst_pe_1_1_6_n26) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_1_6_n113), 
        .CK(npu_inst_pe_1_1_6_net4246), .RN(npu_inst_pe_1_1_6_n9), .Q(
        npu_inst_pe_1_1_6_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_1_6_n107), 
        .CK(npu_inst_pe_1_1_6_net4246), .RN(npu_inst_pe_1_1_6_n9), .Q(
        npu_inst_pe_1_1_6_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_1_6_n112), 
        .CK(npu_inst_pe_1_1_6_net4246), .RN(npu_inst_pe_1_1_6_n10), .Q(
        npu_inst_pe_1_1_6_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_1_6_n106), 
        .CK(npu_inst_pe_1_1_6_net4246), .RN(npu_inst_pe_1_1_6_n10), .Q(
        npu_inst_pe_1_1_6_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_1_6_n111), 
        .CK(npu_inst_pe_1_1_6_net4246), .RN(npu_inst_pe_1_1_6_n10), .Q(
        npu_inst_pe_1_1_6_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_1_6_n105), 
        .CK(npu_inst_pe_1_1_6_net4246), .RN(npu_inst_pe_1_1_6_n10), .Q(
        npu_inst_pe_1_1_6_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_1_6_n110), 
        .CK(npu_inst_pe_1_1_6_net4246), .RN(npu_inst_pe_1_1_6_n10), .Q(
        npu_inst_pe_1_1_6_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_1_6_n104), 
        .CK(npu_inst_pe_1_1_6_net4246), .RN(npu_inst_pe_1_1_6_n10), .Q(
        npu_inst_pe_1_1_6_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_1_6_n109), 
        .CK(npu_inst_pe_1_1_6_net4246), .RN(npu_inst_pe_1_1_6_n10), .Q(
        npu_inst_pe_1_1_6_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_1_6_n103), 
        .CK(npu_inst_pe_1_1_6_net4246), .RN(npu_inst_pe_1_1_6_n10), .Q(
        npu_inst_pe_1_1_6_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_1_6_n108), 
        .CK(npu_inst_pe_1_1_6_net4246), .RN(npu_inst_pe_1_1_6_n10), .Q(
        npu_inst_pe_1_1_6_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_1_6_n102), 
        .CK(npu_inst_pe_1_1_6_net4246), .RN(npu_inst_pe_1_1_6_n10), .Q(
        npu_inst_pe_1_1_6_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_1_6_n86), 
        .CK(npu_inst_pe_1_1_6_net4246), .RN(npu_inst_pe_1_1_6_n10), .Q(
        npu_inst_pe_1_1_6_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_1_6_n87), 
        .CK(npu_inst_pe_1_1_6_net4246), .RN(npu_inst_pe_1_1_6_n10), .Q(
        npu_inst_pe_1_1_6_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_1_6_n88), 
        .CK(npu_inst_pe_1_1_6_net4246), .RN(npu_inst_pe_1_1_6_n11), .Q(
        npu_inst_pe_1_1_6_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_1_6_n89), 
        .CK(npu_inst_pe_1_1_6_net4246), .RN(npu_inst_pe_1_1_6_n11), .Q(
        npu_inst_pe_1_1_6_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_1_6_n90), 
        .CK(npu_inst_pe_1_1_6_net4246), .RN(npu_inst_pe_1_1_6_n11), .Q(
        npu_inst_pe_1_1_6_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_1_6_n91), 
        .CK(npu_inst_pe_1_1_6_net4246), .RN(npu_inst_pe_1_1_6_n11), .Q(
        npu_inst_pe_1_1_6_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_1_6_n92), 
        .CK(npu_inst_pe_1_1_6_net4246), .RN(npu_inst_pe_1_1_6_n11), .Q(
        npu_inst_pe_1_1_6_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_1_6_n93), 
        .CK(npu_inst_pe_1_1_6_net4246), .RN(npu_inst_pe_1_1_6_n11), .Q(
        npu_inst_pe_1_1_6_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_1_6_n94), 
        .CK(npu_inst_pe_1_1_6_net4246), .RN(npu_inst_pe_1_1_6_n11), .Q(
        npu_inst_pe_1_1_6_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_1_6_n95), 
        .CK(npu_inst_pe_1_1_6_net4246), .RN(npu_inst_pe_1_1_6_n11), .Q(
        npu_inst_pe_1_1_6_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_1_6_n96), 
        .CK(npu_inst_pe_1_1_6_net4246), .RN(npu_inst_pe_1_1_6_n11), .Q(
        npu_inst_pe_1_1_6_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_1_6_n97), 
        .CK(npu_inst_pe_1_1_6_net4246), .RN(npu_inst_pe_1_1_6_n11), .Q(
        npu_inst_pe_1_1_6_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_1_6_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_1_6_N84), .SE(1'b0), .GCK(npu_inst_pe_1_1_6_net4240) );
  CLKGATETST_X1 npu_inst_pe_1_1_6_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n65), .SE(1'b0), .GCK(npu_inst_pe_1_1_6_net4246) );
  MUX2_X1 npu_inst_pe_1_1_7_U162 ( .A(npu_inst_pe_1_1_7_n32), .B(
        npu_inst_pe_1_1_7_n29), .S(npu_inst_pe_1_1_7_n8), .Z(
        npu_inst_pe_1_1_7_N93) );
  MUX2_X1 npu_inst_pe_1_1_7_U161 ( .A(npu_inst_pe_1_1_7_n31), .B(
        npu_inst_pe_1_1_7_n30), .S(npu_inst_pe_1_1_7_n6), .Z(
        npu_inst_pe_1_1_7_n32) );
  MUX2_X1 npu_inst_pe_1_1_7_U160 ( .A(npu_inst_pe_1_1_7_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_1_7_int_q_reg_v_1__0_), .S(npu_inst_pe_1_1_7_n4), .Z(
        npu_inst_pe_1_1_7_n31) );
  MUX2_X1 npu_inst_pe_1_1_7_U159 ( .A(npu_inst_pe_1_1_7_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_1_7_int_q_reg_v_3__0_), .S(npu_inst_pe_1_1_7_n4), .Z(
        npu_inst_pe_1_1_7_n30) );
  MUX2_X1 npu_inst_pe_1_1_7_U158 ( .A(npu_inst_pe_1_1_7_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_1_7_int_q_reg_v_5__0_), .S(npu_inst_pe_1_1_7_n4), .Z(
        npu_inst_pe_1_1_7_n29) );
  MUX2_X1 npu_inst_pe_1_1_7_U157 ( .A(npu_inst_pe_1_1_7_n28), .B(
        npu_inst_pe_1_1_7_n23), .S(npu_inst_pe_1_1_7_n8), .Z(
        npu_inst_pe_1_1_7_N94) );
  MUX2_X1 npu_inst_pe_1_1_7_U156 ( .A(npu_inst_pe_1_1_7_n25), .B(
        npu_inst_pe_1_1_7_n24), .S(npu_inst_pe_1_1_7_n6), .Z(
        npu_inst_pe_1_1_7_n28) );
  MUX2_X1 npu_inst_pe_1_1_7_U155 ( .A(npu_inst_pe_1_1_7_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_1_7_int_q_reg_v_1__1_), .S(npu_inst_pe_1_1_7_n4), .Z(
        npu_inst_pe_1_1_7_n25) );
  MUX2_X1 npu_inst_pe_1_1_7_U154 ( .A(npu_inst_pe_1_1_7_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_1_7_int_q_reg_v_3__1_), .S(npu_inst_pe_1_1_7_n4), .Z(
        npu_inst_pe_1_1_7_n24) );
  MUX2_X1 npu_inst_pe_1_1_7_U153 ( .A(npu_inst_pe_1_1_7_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_1_7_int_q_reg_v_5__1_), .S(npu_inst_pe_1_1_7_n4), .Z(
        npu_inst_pe_1_1_7_n23) );
  MUX2_X1 npu_inst_pe_1_1_7_U152 ( .A(npu_inst_pe_1_1_7_n22), .B(
        npu_inst_pe_1_1_7_n19), .S(npu_inst_pe_1_1_7_n8), .Z(
        npu_inst_int_data_x_1__7__1_) );
  MUX2_X1 npu_inst_pe_1_1_7_U151 ( .A(npu_inst_pe_1_1_7_n21), .B(
        npu_inst_pe_1_1_7_n20), .S(npu_inst_pe_1_1_7_n6), .Z(
        npu_inst_pe_1_1_7_n22) );
  MUX2_X1 npu_inst_pe_1_1_7_U150 ( .A(npu_inst_pe_1_1_7_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_1_7_int_q_reg_h_1__1_), .S(npu_inst_pe_1_1_7_n4), .Z(
        npu_inst_pe_1_1_7_n21) );
  MUX2_X1 npu_inst_pe_1_1_7_U149 ( .A(npu_inst_pe_1_1_7_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_1_7_int_q_reg_h_3__1_), .S(npu_inst_pe_1_1_7_n4), .Z(
        npu_inst_pe_1_1_7_n20) );
  MUX2_X1 npu_inst_pe_1_1_7_U148 ( .A(npu_inst_pe_1_1_7_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_1_7_int_q_reg_h_5__1_), .S(npu_inst_pe_1_1_7_n4), .Z(
        npu_inst_pe_1_1_7_n19) );
  MUX2_X1 npu_inst_pe_1_1_7_U147 ( .A(npu_inst_pe_1_1_7_n18), .B(
        npu_inst_pe_1_1_7_n15), .S(npu_inst_pe_1_1_7_n8), .Z(
        npu_inst_int_data_x_1__7__0_) );
  MUX2_X1 npu_inst_pe_1_1_7_U146 ( .A(npu_inst_pe_1_1_7_n17), .B(
        npu_inst_pe_1_1_7_n16), .S(npu_inst_pe_1_1_7_n6), .Z(
        npu_inst_pe_1_1_7_n18) );
  MUX2_X1 npu_inst_pe_1_1_7_U145 ( .A(npu_inst_pe_1_1_7_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_1_7_int_q_reg_h_1__0_), .S(npu_inst_pe_1_1_7_n4), .Z(
        npu_inst_pe_1_1_7_n17) );
  MUX2_X1 npu_inst_pe_1_1_7_U144 ( .A(npu_inst_pe_1_1_7_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_1_7_int_q_reg_h_3__0_), .S(npu_inst_pe_1_1_7_n4), .Z(
        npu_inst_pe_1_1_7_n16) );
  MUX2_X1 npu_inst_pe_1_1_7_U143 ( .A(npu_inst_pe_1_1_7_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_1_7_int_q_reg_h_5__0_), .S(npu_inst_pe_1_1_7_n4), .Z(
        npu_inst_pe_1_1_7_n15) );
  XOR2_X1 npu_inst_pe_1_1_7_U142 ( .A(npu_inst_pe_1_1_7_int_data_0_), .B(
        npu_inst_pe_1_1_7_int_q_acc_0_), .Z(npu_inst_pe_1_1_7_N73) );
  AND2_X1 npu_inst_pe_1_1_7_U141 ( .A1(npu_inst_pe_1_1_7_int_q_acc_0_), .A2(
        npu_inst_pe_1_1_7_int_data_0_), .ZN(npu_inst_pe_1_1_7_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_1_7_U140 ( .A(npu_inst_pe_1_1_7_int_q_acc_0_), .B(
        npu_inst_pe_1_1_7_n13), .ZN(npu_inst_pe_1_1_7_N65) );
  OR2_X1 npu_inst_pe_1_1_7_U139 ( .A1(npu_inst_pe_1_1_7_n13), .A2(
        npu_inst_pe_1_1_7_int_q_acc_0_), .ZN(npu_inst_pe_1_1_7_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_1_7_U138 ( .A(npu_inst_pe_1_1_7_int_q_acc_2_), .B(
        npu_inst_pe_1_1_7_add_69_carry_2_), .Z(npu_inst_pe_1_1_7_N75) );
  AND2_X1 npu_inst_pe_1_1_7_U137 ( .A1(npu_inst_pe_1_1_7_add_69_carry_2_), 
        .A2(npu_inst_pe_1_1_7_int_q_acc_2_), .ZN(
        npu_inst_pe_1_1_7_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_1_7_U136 ( .A(npu_inst_pe_1_1_7_int_q_acc_3_), .B(
        npu_inst_pe_1_1_7_add_69_carry_3_), .Z(npu_inst_pe_1_1_7_N76) );
  AND2_X1 npu_inst_pe_1_1_7_U135 ( .A1(npu_inst_pe_1_1_7_add_69_carry_3_), 
        .A2(npu_inst_pe_1_1_7_int_q_acc_3_), .ZN(
        npu_inst_pe_1_1_7_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_1_7_U134 ( .A(npu_inst_pe_1_1_7_int_q_acc_4_), .B(
        npu_inst_pe_1_1_7_add_69_carry_4_), .Z(npu_inst_pe_1_1_7_N77) );
  AND2_X1 npu_inst_pe_1_1_7_U133 ( .A1(npu_inst_pe_1_1_7_add_69_carry_4_), 
        .A2(npu_inst_pe_1_1_7_int_q_acc_4_), .ZN(
        npu_inst_pe_1_1_7_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_1_7_U132 ( .A(npu_inst_pe_1_1_7_int_q_acc_5_), .B(
        npu_inst_pe_1_1_7_add_69_carry_5_), .Z(npu_inst_pe_1_1_7_N78) );
  AND2_X1 npu_inst_pe_1_1_7_U131 ( .A1(npu_inst_pe_1_1_7_add_69_carry_5_), 
        .A2(npu_inst_pe_1_1_7_int_q_acc_5_), .ZN(
        npu_inst_pe_1_1_7_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_1_7_U130 ( .A(npu_inst_pe_1_1_7_int_q_acc_6_), .B(
        npu_inst_pe_1_1_7_add_69_carry_6_), .Z(npu_inst_pe_1_1_7_N79) );
  AND2_X1 npu_inst_pe_1_1_7_U129 ( .A1(npu_inst_pe_1_1_7_add_69_carry_6_), 
        .A2(npu_inst_pe_1_1_7_int_q_acc_6_), .ZN(
        npu_inst_pe_1_1_7_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_1_7_U128 ( .A(npu_inst_pe_1_1_7_int_q_acc_7_), .B(
        npu_inst_pe_1_1_7_add_69_carry_7_), .Z(npu_inst_pe_1_1_7_N80) );
  XNOR2_X1 npu_inst_pe_1_1_7_U127 ( .A(npu_inst_pe_1_1_7_sub_67_carry_2_), .B(
        npu_inst_pe_1_1_7_int_q_acc_2_), .ZN(npu_inst_pe_1_1_7_N67) );
  OR2_X1 npu_inst_pe_1_1_7_U126 ( .A1(npu_inst_pe_1_1_7_int_q_acc_2_), .A2(
        npu_inst_pe_1_1_7_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_1_7_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_1_7_U125 ( .A(npu_inst_pe_1_1_7_sub_67_carry_3_), .B(
        npu_inst_pe_1_1_7_int_q_acc_3_), .ZN(npu_inst_pe_1_1_7_N68) );
  OR2_X1 npu_inst_pe_1_1_7_U124 ( .A1(npu_inst_pe_1_1_7_int_q_acc_3_), .A2(
        npu_inst_pe_1_1_7_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_1_7_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_1_7_U123 ( .A(npu_inst_pe_1_1_7_sub_67_carry_4_), .B(
        npu_inst_pe_1_1_7_int_q_acc_4_), .ZN(npu_inst_pe_1_1_7_N69) );
  OR2_X1 npu_inst_pe_1_1_7_U122 ( .A1(npu_inst_pe_1_1_7_int_q_acc_4_), .A2(
        npu_inst_pe_1_1_7_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_1_7_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_1_7_U121 ( .A(npu_inst_pe_1_1_7_sub_67_carry_5_), .B(
        npu_inst_pe_1_1_7_int_q_acc_5_), .ZN(npu_inst_pe_1_1_7_N70) );
  OR2_X1 npu_inst_pe_1_1_7_U120 ( .A1(npu_inst_pe_1_1_7_int_q_acc_5_), .A2(
        npu_inst_pe_1_1_7_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_1_7_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_1_7_U119 ( .A(npu_inst_pe_1_1_7_sub_67_carry_6_), .B(
        npu_inst_pe_1_1_7_int_q_acc_6_), .ZN(npu_inst_pe_1_1_7_N71) );
  OR2_X1 npu_inst_pe_1_1_7_U118 ( .A1(npu_inst_pe_1_1_7_int_q_acc_6_), .A2(
        npu_inst_pe_1_1_7_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_1_7_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_1_7_U117 ( .A(npu_inst_pe_1_1_7_int_q_acc_7_), .B(
        npu_inst_pe_1_1_7_sub_67_carry_7_), .ZN(npu_inst_pe_1_1_7_N72) );
  INV_X1 npu_inst_pe_1_1_7_U116 ( .A(npu_inst_n79), .ZN(npu_inst_pe_1_1_7_n7)
         );
  INV_X1 npu_inst_pe_1_1_7_U115 ( .A(npu_inst_pe_1_1_7_n7), .ZN(
        npu_inst_pe_1_1_7_n6) );
  INV_X1 npu_inst_pe_1_1_7_U114 ( .A(npu_inst_n58), .ZN(npu_inst_pe_1_1_7_n3)
         );
  AOI22_X1 npu_inst_pe_1_1_7_U113 ( .A1(npu_inst_int_data_y_2__7__0_), .A2(
        npu_inst_pe_1_1_7_n58), .B1(npu_inst_pe_1_1_7_n119), .B2(
        npu_inst_pe_1_1_7_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_1_7_n57) );
  INV_X1 npu_inst_pe_1_1_7_U112 ( .A(npu_inst_pe_1_1_7_n57), .ZN(
        npu_inst_pe_1_1_7_n108) );
  AOI22_X1 npu_inst_pe_1_1_7_U111 ( .A1(npu_inst_int_data_y_2__7__0_), .A2(
        npu_inst_pe_1_1_7_n54), .B1(npu_inst_pe_1_1_7_n118), .B2(
        npu_inst_pe_1_1_7_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_1_7_n53) );
  INV_X1 npu_inst_pe_1_1_7_U110 ( .A(npu_inst_pe_1_1_7_n53), .ZN(
        npu_inst_pe_1_1_7_n109) );
  AOI22_X1 npu_inst_pe_1_1_7_U107 ( .A1(npu_inst_int_data_y_2__7__0_), .A2(
        npu_inst_pe_1_1_7_n50), .B1(npu_inst_pe_1_1_7_n117), .B2(
        npu_inst_pe_1_1_7_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_1_7_n49) );
  INV_X1 npu_inst_pe_1_1_7_U106 ( .A(npu_inst_pe_1_1_7_n49), .ZN(
        npu_inst_pe_1_1_7_n110) );
  AOI22_X1 npu_inst_pe_1_1_7_U105 ( .A1(npu_inst_int_data_y_2__7__0_), .A2(
        npu_inst_pe_1_1_7_n46), .B1(npu_inst_pe_1_1_7_n116), .B2(
        npu_inst_pe_1_1_7_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_1_7_n45) );
  INV_X1 npu_inst_pe_1_1_7_U104 ( .A(npu_inst_pe_1_1_7_n45), .ZN(
        npu_inst_pe_1_1_7_n111) );
  AOI22_X1 npu_inst_pe_1_1_7_U103 ( .A1(npu_inst_int_data_y_2__7__0_), .A2(
        npu_inst_pe_1_1_7_n42), .B1(npu_inst_pe_1_1_7_n115), .B2(
        npu_inst_pe_1_1_7_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_1_7_n41) );
  INV_X1 npu_inst_pe_1_1_7_U102 ( .A(npu_inst_pe_1_1_7_n41), .ZN(
        npu_inst_pe_1_1_7_n112) );
  AOI22_X1 npu_inst_pe_1_1_7_U101 ( .A1(npu_inst_int_data_y_2__7__1_), .A2(
        npu_inst_pe_1_1_7_n58), .B1(npu_inst_pe_1_1_7_n119), .B2(
        npu_inst_pe_1_1_7_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_1_7_n59) );
  INV_X1 npu_inst_pe_1_1_7_U100 ( .A(npu_inst_pe_1_1_7_n59), .ZN(
        npu_inst_pe_1_1_7_n102) );
  AOI22_X1 npu_inst_pe_1_1_7_U99 ( .A1(npu_inst_int_data_y_2__7__1_), .A2(
        npu_inst_pe_1_1_7_n54), .B1(npu_inst_pe_1_1_7_n118), .B2(
        npu_inst_pe_1_1_7_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_1_7_n55) );
  INV_X1 npu_inst_pe_1_1_7_U98 ( .A(npu_inst_pe_1_1_7_n55), .ZN(
        npu_inst_pe_1_1_7_n103) );
  AOI22_X1 npu_inst_pe_1_1_7_U97 ( .A1(npu_inst_int_data_y_2__7__1_), .A2(
        npu_inst_pe_1_1_7_n50), .B1(npu_inst_pe_1_1_7_n117), .B2(
        npu_inst_pe_1_1_7_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_1_7_n51) );
  INV_X1 npu_inst_pe_1_1_7_U96 ( .A(npu_inst_pe_1_1_7_n51), .ZN(
        npu_inst_pe_1_1_7_n104) );
  AOI22_X1 npu_inst_pe_1_1_7_U95 ( .A1(npu_inst_int_data_y_2__7__1_), .A2(
        npu_inst_pe_1_1_7_n46), .B1(npu_inst_pe_1_1_7_n116), .B2(
        npu_inst_pe_1_1_7_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_1_7_n47) );
  INV_X1 npu_inst_pe_1_1_7_U94 ( .A(npu_inst_pe_1_1_7_n47), .ZN(
        npu_inst_pe_1_1_7_n105) );
  AOI22_X1 npu_inst_pe_1_1_7_U93 ( .A1(npu_inst_int_data_y_2__7__1_), .A2(
        npu_inst_pe_1_1_7_n42), .B1(npu_inst_pe_1_1_7_n115), .B2(
        npu_inst_pe_1_1_7_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_1_7_n43) );
  INV_X1 npu_inst_pe_1_1_7_U92 ( .A(npu_inst_pe_1_1_7_n43), .ZN(
        npu_inst_pe_1_1_7_n106) );
  AOI22_X1 npu_inst_pe_1_1_7_U91 ( .A1(npu_inst_pe_1_1_7_n38), .A2(
        npu_inst_int_data_y_2__7__1_), .B1(npu_inst_pe_1_1_7_n114), .B2(
        npu_inst_pe_1_1_7_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_1_7_n39) );
  INV_X1 npu_inst_pe_1_1_7_U90 ( .A(npu_inst_pe_1_1_7_n39), .ZN(
        npu_inst_pe_1_1_7_n107) );
  AOI22_X1 npu_inst_pe_1_1_7_U89 ( .A1(npu_inst_pe_1_1_7_n38), .A2(
        npu_inst_int_data_y_2__7__0_), .B1(npu_inst_pe_1_1_7_n114), .B2(
        npu_inst_pe_1_1_7_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_1_7_n37) );
  INV_X1 npu_inst_pe_1_1_7_U88 ( .A(npu_inst_pe_1_1_7_n37), .ZN(
        npu_inst_pe_1_1_7_n113) );
  AND2_X1 npu_inst_pe_1_1_7_U87 ( .A1(npu_inst_pe_1_1_7_N93), .A2(npu_inst_n58), .ZN(npu_inst_int_data_y_1__7__0_) );
  AND2_X1 npu_inst_pe_1_1_7_U86 ( .A1(npu_inst_n58), .A2(npu_inst_pe_1_1_7_N94), .ZN(npu_inst_int_data_y_1__7__1_) );
  NOR3_X1 npu_inst_pe_1_1_7_U85 ( .A1(npu_inst_pe_1_1_7_n26), .A2(npu_inst_n58), .A3(npu_inst_int_ckg[48]), .ZN(npu_inst_pe_1_1_7_n85) );
  OR2_X1 npu_inst_pe_1_1_7_U84 ( .A1(npu_inst_pe_1_1_7_n85), .A2(
        npu_inst_pe_1_1_7_n2), .ZN(npu_inst_pe_1_1_7_N84) );
  AND2_X1 npu_inst_pe_1_1_7_U83 ( .A1(npu_inst_pe_1_1_7_int_q_acc_0_), .A2(
        npu_inst_pe_1_1_7_n1), .ZN(npu_inst_int_data_res_1__7__0_) );
  AND2_X1 npu_inst_pe_1_1_7_U82 ( .A1(npu_inst_pe_1_1_7_n2), .A2(
        npu_inst_pe_1_1_7_int_q_acc_7_), .ZN(npu_inst_int_data_res_1__7__7_)
         );
  AND2_X1 npu_inst_pe_1_1_7_U81 ( .A1(npu_inst_pe_1_1_7_int_q_acc_1_), .A2(
        npu_inst_pe_1_1_7_n1), .ZN(npu_inst_int_data_res_1__7__1_) );
  AND2_X1 npu_inst_pe_1_1_7_U80 ( .A1(npu_inst_pe_1_1_7_int_q_acc_2_), .A2(
        npu_inst_pe_1_1_7_n1), .ZN(npu_inst_int_data_res_1__7__2_) );
  AND2_X1 npu_inst_pe_1_1_7_U79 ( .A1(npu_inst_pe_1_1_7_int_q_acc_3_), .A2(
        npu_inst_pe_1_1_7_n2), .ZN(npu_inst_int_data_res_1__7__3_) );
  AND2_X1 npu_inst_pe_1_1_7_U78 ( .A1(npu_inst_pe_1_1_7_int_q_acc_4_), .A2(
        npu_inst_pe_1_1_7_n2), .ZN(npu_inst_int_data_res_1__7__4_) );
  AND2_X1 npu_inst_pe_1_1_7_U77 ( .A1(npu_inst_pe_1_1_7_int_q_acc_5_), .A2(
        npu_inst_pe_1_1_7_n2), .ZN(npu_inst_int_data_res_1__7__5_) );
  AND2_X1 npu_inst_pe_1_1_7_U76 ( .A1(npu_inst_pe_1_1_7_int_q_acc_6_), .A2(
        npu_inst_pe_1_1_7_n2), .ZN(npu_inst_int_data_res_1__7__6_) );
  AOI222_X1 npu_inst_pe_1_1_7_U75 ( .A1(npu_inst_int_data_res_2__7__0_), .A2(
        npu_inst_pe_1_1_7_n1), .B1(npu_inst_pe_1_1_7_N73), .B2(
        npu_inst_pe_1_1_7_n76), .C1(npu_inst_pe_1_1_7_N65), .C2(
        npu_inst_pe_1_1_7_n77), .ZN(npu_inst_pe_1_1_7_n84) );
  INV_X1 npu_inst_pe_1_1_7_U74 ( .A(npu_inst_pe_1_1_7_n84), .ZN(
        npu_inst_pe_1_1_7_n101) );
  AOI222_X1 npu_inst_pe_1_1_7_U73 ( .A1(npu_inst_int_data_res_2__7__7_), .A2(
        npu_inst_pe_1_1_7_n1), .B1(npu_inst_pe_1_1_7_N80), .B2(
        npu_inst_pe_1_1_7_n76), .C1(npu_inst_pe_1_1_7_N72), .C2(
        npu_inst_pe_1_1_7_n77), .ZN(npu_inst_pe_1_1_7_n75) );
  INV_X1 npu_inst_pe_1_1_7_U72 ( .A(npu_inst_pe_1_1_7_n75), .ZN(
        npu_inst_pe_1_1_7_n33) );
  AOI222_X1 npu_inst_pe_1_1_7_U71 ( .A1(npu_inst_int_data_res_2__7__1_), .A2(
        npu_inst_pe_1_1_7_n1), .B1(npu_inst_pe_1_1_7_N74), .B2(
        npu_inst_pe_1_1_7_n76), .C1(npu_inst_pe_1_1_7_N66), .C2(
        npu_inst_pe_1_1_7_n77), .ZN(npu_inst_pe_1_1_7_n83) );
  INV_X1 npu_inst_pe_1_1_7_U70 ( .A(npu_inst_pe_1_1_7_n83), .ZN(
        npu_inst_pe_1_1_7_n100) );
  AOI222_X1 npu_inst_pe_1_1_7_U69 ( .A1(npu_inst_int_data_res_2__7__2_), .A2(
        npu_inst_pe_1_1_7_n1), .B1(npu_inst_pe_1_1_7_N75), .B2(
        npu_inst_pe_1_1_7_n76), .C1(npu_inst_pe_1_1_7_N67), .C2(
        npu_inst_pe_1_1_7_n77), .ZN(npu_inst_pe_1_1_7_n82) );
  INV_X1 npu_inst_pe_1_1_7_U68 ( .A(npu_inst_pe_1_1_7_n82), .ZN(
        npu_inst_pe_1_1_7_n99) );
  AOI222_X1 npu_inst_pe_1_1_7_U67 ( .A1(npu_inst_int_data_res_2__7__3_), .A2(
        npu_inst_pe_1_1_7_n1), .B1(npu_inst_pe_1_1_7_N76), .B2(
        npu_inst_pe_1_1_7_n76), .C1(npu_inst_pe_1_1_7_N68), .C2(
        npu_inst_pe_1_1_7_n77), .ZN(npu_inst_pe_1_1_7_n81) );
  INV_X1 npu_inst_pe_1_1_7_U66 ( .A(npu_inst_pe_1_1_7_n81), .ZN(
        npu_inst_pe_1_1_7_n98) );
  AOI222_X1 npu_inst_pe_1_1_7_U65 ( .A1(npu_inst_int_data_res_2__7__4_), .A2(
        npu_inst_pe_1_1_7_n1), .B1(npu_inst_pe_1_1_7_N77), .B2(
        npu_inst_pe_1_1_7_n76), .C1(npu_inst_pe_1_1_7_N69), .C2(
        npu_inst_pe_1_1_7_n77), .ZN(npu_inst_pe_1_1_7_n80) );
  INV_X1 npu_inst_pe_1_1_7_U64 ( .A(npu_inst_pe_1_1_7_n80), .ZN(
        npu_inst_pe_1_1_7_n36) );
  AOI222_X1 npu_inst_pe_1_1_7_U63 ( .A1(npu_inst_int_data_res_2__7__5_), .A2(
        npu_inst_pe_1_1_7_n1), .B1(npu_inst_pe_1_1_7_N78), .B2(
        npu_inst_pe_1_1_7_n76), .C1(npu_inst_pe_1_1_7_N70), .C2(
        npu_inst_pe_1_1_7_n77), .ZN(npu_inst_pe_1_1_7_n79) );
  INV_X1 npu_inst_pe_1_1_7_U62 ( .A(npu_inst_pe_1_1_7_n79), .ZN(
        npu_inst_pe_1_1_7_n35) );
  AOI222_X1 npu_inst_pe_1_1_7_U61 ( .A1(npu_inst_int_data_res_2__7__6_), .A2(
        npu_inst_pe_1_1_7_n1), .B1(npu_inst_pe_1_1_7_N79), .B2(
        npu_inst_pe_1_1_7_n76), .C1(npu_inst_pe_1_1_7_N71), .C2(
        npu_inst_pe_1_1_7_n77), .ZN(npu_inst_pe_1_1_7_n78) );
  INV_X1 npu_inst_pe_1_1_7_U60 ( .A(npu_inst_pe_1_1_7_n78), .ZN(
        npu_inst_pe_1_1_7_n34) );
  INV_X1 npu_inst_pe_1_1_7_U59 ( .A(npu_inst_pe_1_1_7_int_data_1_), .ZN(
        npu_inst_pe_1_1_7_n14) );
  AND2_X1 npu_inst_pe_1_1_7_U58 ( .A1(npu_inst_int_data_x_1__7__1_), .A2(
        npu_inst_pe_1_1_7_int_q_weight_1_), .ZN(npu_inst_pe_1_1_7_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_1_7_U57 ( .A1(npu_inst_int_data_x_1__7__0_), .A2(
        npu_inst_pe_1_1_7_int_q_weight_1_), .ZN(npu_inst_pe_1_1_7_int_data_0_)
         );
  NAND2_X1 npu_inst_pe_1_1_7_U56 ( .A1(npu_inst_pe_1_1_7_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_1_7_n60), .ZN(npu_inst_pe_1_1_7_n74) );
  OAI21_X1 npu_inst_pe_1_1_7_U55 ( .B1(npu_inst_pe_1_1_7_n63), .B2(
        npu_inst_pe_1_1_7_n60), .A(npu_inst_pe_1_1_7_n74), .ZN(
        npu_inst_pe_1_1_7_n97) );
  NAND2_X1 npu_inst_pe_1_1_7_U54 ( .A1(npu_inst_pe_1_1_7_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_1_7_n60), .ZN(npu_inst_pe_1_1_7_n73) );
  OAI21_X1 npu_inst_pe_1_1_7_U53 ( .B1(npu_inst_pe_1_1_7_n61), .B2(
        npu_inst_pe_1_1_7_n60), .A(npu_inst_pe_1_1_7_n73), .ZN(
        npu_inst_pe_1_1_7_n96) );
  NAND2_X1 npu_inst_pe_1_1_7_U52 ( .A1(npu_inst_pe_1_1_7_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_1_7_n56), .ZN(npu_inst_pe_1_1_7_n72) );
  OAI21_X1 npu_inst_pe_1_1_7_U51 ( .B1(npu_inst_pe_1_1_7_n63), .B2(
        npu_inst_pe_1_1_7_n56), .A(npu_inst_pe_1_1_7_n72), .ZN(
        npu_inst_pe_1_1_7_n95) );
  NAND2_X1 npu_inst_pe_1_1_7_U50 ( .A1(npu_inst_pe_1_1_7_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_1_7_n56), .ZN(npu_inst_pe_1_1_7_n71) );
  OAI21_X1 npu_inst_pe_1_1_7_U49 ( .B1(npu_inst_pe_1_1_7_n61), .B2(
        npu_inst_pe_1_1_7_n56), .A(npu_inst_pe_1_1_7_n71), .ZN(
        npu_inst_pe_1_1_7_n94) );
  NAND2_X1 npu_inst_pe_1_1_7_U48 ( .A1(npu_inst_pe_1_1_7_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_1_7_n52), .ZN(npu_inst_pe_1_1_7_n70) );
  OAI21_X1 npu_inst_pe_1_1_7_U47 ( .B1(npu_inst_pe_1_1_7_n63), .B2(
        npu_inst_pe_1_1_7_n52), .A(npu_inst_pe_1_1_7_n70), .ZN(
        npu_inst_pe_1_1_7_n93) );
  NAND2_X1 npu_inst_pe_1_1_7_U46 ( .A1(npu_inst_pe_1_1_7_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_1_7_n52), .ZN(npu_inst_pe_1_1_7_n69) );
  OAI21_X1 npu_inst_pe_1_1_7_U45 ( .B1(npu_inst_pe_1_1_7_n61), .B2(
        npu_inst_pe_1_1_7_n52), .A(npu_inst_pe_1_1_7_n69), .ZN(
        npu_inst_pe_1_1_7_n92) );
  NAND2_X1 npu_inst_pe_1_1_7_U44 ( .A1(npu_inst_pe_1_1_7_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_1_7_n48), .ZN(npu_inst_pe_1_1_7_n68) );
  OAI21_X1 npu_inst_pe_1_1_7_U43 ( .B1(npu_inst_pe_1_1_7_n63), .B2(
        npu_inst_pe_1_1_7_n48), .A(npu_inst_pe_1_1_7_n68), .ZN(
        npu_inst_pe_1_1_7_n91) );
  NAND2_X1 npu_inst_pe_1_1_7_U42 ( .A1(npu_inst_pe_1_1_7_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_1_7_n48), .ZN(npu_inst_pe_1_1_7_n67) );
  OAI21_X1 npu_inst_pe_1_1_7_U41 ( .B1(npu_inst_pe_1_1_7_n61), .B2(
        npu_inst_pe_1_1_7_n48), .A(npu_inst_pe_1_1_7_n67), .ZN(
        npu_inst_pe_1_1_7_n90) );
  NAND2_X1 npu_inst_pe_1_1_7_U40 ( .A1(npu_inst_pe_1_1_7_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_1_7_n44), .ZN(npu_inst_pe_1_1_7_n66) );
  OAI21_X1 npu_inst_pe_1_1_7_U39 ( .B1(npu_inst_pe_1_1_7_n63), .B2(
        npu_inst_pe_1_1_7_n44), .A(npu_inst_pe_1_1_7_n66), .ZN(
        npu_inst_pe_1_1_7_n89) );
  NAND2_X1 npu_inst_pe_1_1_7_U38 ( .A1(npu_inst_pe_1_1_7_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_1_7_n44), .ZN(npu_inst_pe_1_1_7_n65) );
  OAI21_X1 npu_inst_pe_1_1_7_U37 ( .B1(npu_inst_pe_1_1_7_n61), .B2(
        npu_inst_pe_1_1_7_n44), .A(npu_inst_pe_1_1_7_n65), .ZN(
        npu_inst_pe_1_1_7_n88) );
  NAND2_X1 npu_inst_pe_1_1_7_U36 ( .A1(npu_inst_pe_1_1_7_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_1_7_n40), .ZN(npu_inst_pe_1_1_7_n64) );
  OAI21_X1 npu_inst_pe_1_1_7_U35 ( .B1(npu_inst_pe_1_1_7_n63), .B2(
        npu_inst_pe_1_1_7_n40), .A(npu_inst_pe_1_1_7_n64), .ZN(
        npu_inst_pe_1_1_7_n87) );
  NAND2_X1 npu_inst_pe_1_1_7_U34 ( .A1(npu_inst_pe_1_1_7_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_1_7_n40), .ZN(npu_inst_pe_1_1_7_n62) );
  OAI21_X1 npu_inst_pe_1_1_7_U33 ( .B1(npu_inst_pe_1_1_7_n61), .B2(
        npu_inst_pe_1_1_7_n40), .A(npu_inst_pe_1_1_7_n62), .ZN(
        npu_inst_pe_1_1_7_n86) );
  INV_X1 npu_inst_pe_1_1_7_U32 ( .A(npu_inst_pe_1_1_7_int_data_0_), .ZN(
        npu_inst_pe_1_1_7_n13) );
  INV_X1 npu_inst_pe_1_1_7_U31 ( .A(npu_inst_n71), .ZN(npu_inst_pe_1_1_7_n5)
         );
  AOI22_X1 npu_inst_pe_1_1_7_U30 ( .A1(npu_inst_n58), .A2(
        npu_inst_int_data_y_2__7__1_), .B1(npu_inst_pe_1_1_7_n3), .B2(
        int_i_data_h_npu[13]), .ZN(npu_inst_pe_1_1_7_n63) );
  AOI22_X1 npu_inst_pe_1_1_7_U29 ( .A1(npu_inst_n58), .A2(
        npu_inst_int_data_y_2__7__0_), .B1(npu_inst_pe_1_1_7_n3), .B2(
        int_i_data_h_npu[12]), .ZN(npu_inst_pe_1_1_7_n61) );
  OR3_X1 npu_inst_pe_1_1_7_U28 ( .A1(npu_inst_pe_1_1_7_n6), .A2(
        npu_inst_pe_1_1_7_n8), .A3(npu_inst_pe_1_1_7_n5), .ZN(
        npu_inst_pe_1_1_7_n56) );
  OR3_X1 npu_inst_pe_1_1_7_U27 ( .A1(npu_inst_pe_1_1_7_n5), .A2(
        npu_inst_pe_1_1_7_n8), .A3(npu_inst_pe_1_1_7_n7), .ZN(
        npu_inst_pe_1_1_7_n48) );
  INV_X1 npu_inst_pe_1_1_7_U26 ( .A(npu_inst_pe_1_1_7_n5), .ZN(
        npu_inst_pe_1_1_7_n4) );
  OR3_X1 npu_inst_pe_1_1_7_U25 ( .A1(npu_inst_pe_1_1_7_n4), .A2(
        npu_inst_pe_1_1_7_n8), .A3(npu_inst_pe_1_1_7_n7), .ZN(
        npu_inst_pe_1_1_7_n52) );
  OR3_X1 npu_inst_pe_1_1_7_U24 ( .A1(npu_inst_pe_1_1_7_n6), .A2(
        npu_inst_pe_1_1_7_n8), .A3(npu_inst_pe_1_1_7_n4), .ZN(
        npu_inst_pe_1_1_7_n60) );
  NOR2_X1 npu_inst_pe_1_1_7_U23 ( .A1(npu_inst_pe_1_1_7_n60), .A2(
        npu_inst_pe_1_1_7_n3), .ZN(npu_inst_pe_1_1_7_n58) );
  NOR2_X1 npu_inst_pe_1_1_7_U22 ( .A1(npu_inst_pe_1_1_7_n56), .A2(
        npu_inst_pe_1_1_7_n3), .ZN(npu_inst_pe_1_1_7_n54) );
  NOR2_X1 npu_inst_pe_1_1_7_U21 ( .A1(npu_inst_pe_1_1_7_n52), .A2(
        npu_inst_pe_1_1_7_n3), .ZN(npu_inst_pe_1_1_7_n50) );
  NOR2_X1 npu_inst_pe_1_1_7_U20 ( .A1(npu_inst_pe_1_1_7_n48), .A2(
        npu_inst_pe_1_1_7_n3), .ZN(npu_inst_pe_1_1_7_n46) );
  NOR2_X1 npu_inst_pe_1_1_7_U19 ( .A1(npu_inst_pe_1_1_7_n40), .A2(
        npu_inst_pe_1_1_7_n3), .ZN(npu_inst_pe_1_1_7_n38) );
  NOR2_X1 npu_inst_pe_1_1_7_U18 ( .A1(npu_inst_pe_1_1_7_n44), .A2(
        npu_inst_pe_1_1_7_n3), .ZN(npu_inst_pe_1_1_7_n42) );
  BUF_X1 npu_inst_pe_1_1_7_U17 ( .A(npu_inst_n104), .Z(npu_inst_pe_1_1_7_n8)
         );
  INV_X1 npu_inst_pe_1_1_7_U16 ( .A(npu_inst_n126), .ZN(npu_inst_pe_1_1_7_n12)
         );
  INV_X1 npu_inst_pe_1_1_7_U15 ( .A(npu_inst_pe_1_1_7_n38), .ZN(
        npu_inst_pe_1_1_7_n114) );
  INV_X1 npu_inst_pe_1_1_7_U14 ( .A(npu_inst_pe_1_1_7_n58), .ZN(
        npu_inst_pe_1_1_7_n119) );
  INV_X1 npu_inst_pe_1_1_7_U13 ( .A(npu_inst_pe_1_1_7_n54), .ZN(
        npu_inst_pe_1_1_7_n118) );
  INV_X1 npu_inst_pe_1_1_7_U12 ( .A(npu_inst_pe_1_1_7_n50), .ZN(
        npu_inst_pe_1_1_7_n117) );
  INV_X1 npu_inst_pe_1_1_7_U11 ( .A(npu_inst_pe_1_1_7_n46), .ZN(
        npu_inst_pe_1_1_7_n116) );
  INV_X1 npu_inst_pe_1_1_7_U10 ( .A(npu_inst_pe_1_1_7_n42), .ZN(
        npu_inst_pe_1_1_7_n115) );
  BUF_X1 npu_inst_pe_1_1_7_U9 ( .A(npu_inst_n31), .Z(npu_inst_pe_1_1_7_n2) );
  BUF_X1 npu_inst_pe_1_1_7_U8 ( .A(npu_inst_n31), .Z(npu_inst_pe_1_1_7_n1) );
  BUF_X1 npu_inst_pe_1_1_7_U7 ( .A(npu_inst_pe_1_1_7_n12), .Z(
        npu_inst_pe_1_1_7_n11) );
  BUF_X1 npu_inst_pe_1_1_7_U6 ( .A(npu_inst_pe_1_1_7_n12), .Z(
        npu_inst_pe_1_1_7_n10) );
  BUF_X1 npu_inst_pe_1_1_7_U5 ( .A(npu_inst_pe_1_1_7_n12), .Z(
        npu_inst_pe_1_1_7_n9) );
  NOR2_X1 npu_inst_pe_1_1_7_U4 ( .A1(npu_inst_pe_1_1_7_int_q_weight_0_), .A2(
        npu_inst_pe_1_1_7_n1), .ZN(npu_inst_pe_1_1_7_n76) );
  NOR2_X1 npu_inst_pe_1_1_7_U3 ( .A1(npu_inst_pe_1_1_7_n27), .A2(
        npu_inst_pe_1_1_7_n1), .ZN(npu_inst_pe_1_1_7_n77) );
  FA_X1 npu_inst_pe_1_1_7_sub_67_U2_1 ( .A(npu_inst_pe_1_1_7_int_q_acc_1_), 
        .B(npu_inst_pe_1_1_7_n14), .CI(npu_inst_pe_1_1_7_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_1_7_sub_67_carry_2_), .S(npu_inst_pe_1_1_7_N66) );
  FA_X1 npu_inst_pe_1_1_7_add_69_U1_1 ( .A(npu_inst_pe_1_1_7_int_q_acc_1_), 
        .B(npu_inst_pe_1_1_7_int_data_1_), .CI(
        npu_inst_pe_1_1_7_add_69_carry_1_), .CO(
        npu_inst_pe_1_1_7_add_69_carry_2_), .S(npu_inst_pe_1_1_7_N74) );
  NAND3_X1 npu_inst_pe_1_1_7_U109 ( .A1(npu_inst_pe_1_1_7_n5), .A2(
        npu_inst_pe_1_1_7_n7), .A3(npu_inst_pe_1_1_7_n8), .ZN(
        npu_inst_pe_1_1_7_n44) );
  NAND3_X1 npu_inst_pe_1_1_7_U108 ( .A1(npu_inst_pe_1_1_7_n4), .A2(
        npu_inst_pe_1_1_7_n7), .A3(npu_inst_pe_1_1_7_n8), .ZN(
        npu_inst_pe_1_1_7_n40) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_1_7_n34), .CK(
        npu_inst_pe_1_1_7_net4217), .RN(npu_inst_pe_1_1_7_n9), .Q(
        npu_inst_pe_1_1_7_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_1_7_n35), .CK(
        npu_inst_pe_1_1_7_net4217), .RN(npu_inst_pe_1_1_7_n9), .Q(
        npu_inst_pe_1_1_7_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_1_7_n36), .CK(
        npu_inst_pe_1_1_7_net4217), .RN(npu_inst_pe_1_1_7_n9), .Q(
        npu_inst_pe_1_1_7_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_1_7_n98), .CK(
        npu_inst_pe_1_1_7_net4217), .RN(npu_inst_pe_1_1_7_n9), .Q(
        npu_inst_pe_1_1_7_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_1_7_n99), .CK(
        npu_inst_pe_1_1_7_net4217), .RN(npu_inst_pe_1_1_7_n9), .Q(
        npu_inst_pe_1_1_7_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_1_7_n100), 
        .CK(npu_inst_pe_1_1_7_net4217), .RN(npu_inst_pe_1_1_7_n9), .Q(
        npu_inst_pe_1_1_7_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_1_7_n33), .CK(
        npu_inst_pe_1_1_7_net4217), .RN(npu_inst_pe_1_1_7_n9), .Q(
        npu_inst_pe_1_1_7_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_1_7_n101), 
        .CK(npu_inst_pe_1_1_7_net4217), .RN(npu_inst_pe_1_1_7_n9), .Q(
        npu_inst_pe_1_1_7_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_weight_reg_0_ ( .D(npu_inst_n112), .CK(
        npu_inst_pe_1_1_7_net4223), .RN(npu_inst_pe_1_1_7_n9), .Q(
        npu_inst_pe_1_1_7_int_q_weight_0_), .QN(npu_inst_pe_1_1_7_n27) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_weight_reg_1_ ( .D(npu_inst_n118), .CK(
        npu_inst_pe_1_1_7_net4223), .RN(npu_inst_pe_1_1_7_n9), .Q(
        npu_inst_pe_1_1_7_int_q_weight_1_), .QN(npu_inst_pe_1_1_7_n26) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_1_7_n113), 
        .CK(npu_inst_pe_1_1_7_net4223), .RN(npu_inst_pe_1_1_7_n9), .Q(
        npu_inst_pe_1_1_7_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_1_7_n107), 
        .CK(npu_inst_pe_1_1_7_net4223), .RN(npu_inst_pe_1_1_7_n9), .Q(
        npu_inst_pe_1_1_7_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_1_7_n112), 
        .CK(npu_inst_pe_1_1_7_net4223), .RN(npu_inst_pe_1_1_7_n10), .Q(
        npu_inst_pe_1_1_7_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_1_7_n106), 
        .CK(npu_inst_pe_1_1_7_net4223), .RN(npu_inst_pe_1_1_7_n10), .Q(
        npu_inst_pe_1_1_7_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_1_7_n111), 
        .CK(npu_inst_pe_1_1_7_net4223), .RN(npu_inst_pe_1_1_7_n10), .Q(
        npu_inst_pe_1_1_7_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_1_7_n105), 
        .CK(npu_inst_pe_1_1_7_net4223), .RN(npu_inst_pe_1_1_7_n10), .Q(
        npu_inst_pe_1_1_7_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_1_7_n110), 
        .CK(npu_inst_pe_1_1_7_net4223), .RN(npu_inst_pe_1_1_7_n10), .Q(
        npu_inst_pe_1_1_7_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_1_7_n104), 
        .CK(npu_inst_pe_1_1_7_net4223), .RN(npu_inst_pe_1_1_7_n10), .Q(
        npu_inst_pe_1_1_7_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_1_7_n109), 
        .CK(npu_inst_pe_1_1_7_net4223), .RN(npu_inst_pe_1_1_7_n10), .Q(
        npu_inst_pe_1_1_7_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_1_7_n103), 
        .CK(npu_inst_pe_1_1_7_net4223), .RN(npu_inst_pe_1_1_7_n10), .Q(
        npu_inst_pe_1_1_7_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_1_7_n108), 
        .CK(npu_inst_pe_1_1_7_net4223), .RN(npu_inst_pe_1_1_7_n10), .Q(
        npu_inst_pe_1_1_7_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_1_7_n102), 
        .CK(npu_inst_pe_1_1_7_net4223), .RN(npu_inst_pe_1_1_7_n10), .Q(
        npu_inst_pe_1_1_7_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_1_7_n86), 
        .CK(npu_inst_pe_1_1_7_net4223), .RN(npu_inst_pe_1_1_7_n10), .Q(
        npu_inst_pe_1_1_7_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_1_7_n87), 
        .CK(npu_inst_pe_1_1_7_net4223), .RN(npu_inst_pe_1_1_7_n10), .Q(
        npu_inst_pe_1_1_7_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_1_7_n88), 
        .CK(npu_inst_pe_1_1_7_net4223), .RN(npu_inst_pe_1_1_7_n11), .Q(
        npu_inst_pe_1_1_7_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_1_7_n89), 
        .CK(npu_inst_pe_1_1_7_net4223), .RN(npu_inst_pe_1_1_7_n11), .Q(
        npu_inst_pe_1_1_7_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_1_7_n90), 
        .CK(npu_inst_pe_1_1_7_net4223), .RN(npu_inst_pe_1_1_7_n11), .Q(
        npu_inst_pe_1_1_7_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_1_7_n91), 
        .CK(npu_inst_pe_1_1_7_net4223), .RN(npu_inst_pe_1_1_7_n11), .Q(
        npu_inst_pe_1_1_7_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_1_7_n92), 
        .CK(npu_inst_pe_1_1_7_net4223), .RN(npu_inst_pe_1_1_7_n11), .Q(
        npu_inst_pe_1_1_7_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_1_7_n93), 
        .CK(npu_inst_pe_1_1_7_net4223), .RN(npu_inst_pe_1_1_7_n11), .Q(
        npu_inst_pe_1_1_7_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_1_7_n94), 
        .CK(npu_inst_pe_1_1_7_net4223), .RN(npu_inst_pe_1_1_7_n11), .Q(
        npu_inst_pe_1_1_7_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_1_7_n95), 
        .CK(npu_inst_pe_1_1_7_net4223), .RN(npu_inst_pe_1_1_7_n11), .Q(
        npu_inst_pe_1_1_7_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_1_7_n96), 
        .CK(npu_inst_pe_1_1_7_net4223), .RN(npu_inst_pe_1_1_7_n11), .Q(
        npu_inst_pe_1_1_7_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_1_7_n97), 
        .CK(npu_inst_pe_1_1_7_net4223), .RN(npu_inst_pe_1_1_7_n11), .Q(
        npu_inst_pe_1_1_7_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_1_7_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_1_7_N84), .SE(1'b0), .GCK(npu_inst_pe_1_1_7_net4217) );
  CLKGATETST_X1 npu_inst_pe_1_1_7_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n65), .SE(1'b0), .GCK(npu_inst_pe_1_1_7_net4223) );
  MUX2_X1 npu_inst_pe_1_2_0_U161 ( .A(npu_inst_pe_1_2_0_n31), .B(
        npu_inst_pe_1_2_0_n28), .S(npu_inst_pe_1_2_0_n7), .Z(
        npu_inst_pe_1_2_0_N93) );
  MUX2_X1 npu_inst_pe_1_2_0_U160 ( .A(npu_inst_pe_1_2_0_n30), .B(
        npu_inst_pe_1_2_0_n29), .S(npu_inst_n78), .Z(npu_inst_pe_1_2_0_n31) );
  MUX2_X1 npu_inst_pe_1_2_0_U159 ( .A(npu_inst_pe_1_2_0_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_2_0_int_q_reg_v_1__0_), .S(npu_inst_pe_1_2_0_n4), .Z(
        npu_inst_pe_1_2_0_n30) );
  MUX2_X1 npu_inst_pe_1_2_0_U158 ( .A(npu_inst_pe_1_2_0_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_2_0_int_q_reg_v_3__0_), .S(npu_inst_pe_1_2_0_n4), .Z(
        npu_inst_pe_1_2_0_n29) );
  MUX2_X1 npu_inst_pe_1_2_0_U157 ( .A(npu_inst_pe_1_2_0_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_2_0_int_q_reg_v_5__0_), .S(npu_inst_pe_1_2_0_n4), .Z(
        npu_inst_pe_1_2_0_n28) );
  MUX2_X1 npu_inst_pe_1_2_0_U156 ( .A(npu_inst_pe_1_2_0_n25), .B(
        npu_inst_pe_1_2_0_n22), .S(npu_inst_pe_1_2_0_n7), .Z(
        npu_inst_pe_1_2_0_N94) );
  MUX2_X1 npu_inst_pe_1_2_0_U155 ( .A(npu_inst_pe_1_2_0_n24), .B(
        npu_inst_pe_1_2_0_n23), .S(npu_inst_n78), .Z(npu_inst_pe_1_2_0_n25) );
  MUX2_X1 npu_inst_pe_1_2_0_U154 ( .A(npu_inst_pe_1_2_0_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_2_0_int_q_reg_v_1__1_), .S(npu_inst_pe_1_2_0_n4), .Z(
        npu_inst_pe_1_2_0_n24) );
  MUX2_X1 npu_inst_pe_1_2_0_U153 ( .A(npu_inst_pe_1_2_0_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_2_0_int_q_reg_v_3__1_), .S(npu_inst_pe_1_2_0_n4), .Z(
        npu_inst_pe_1_2_0_n23) );
  MUX2_X1 npu_inst_pe_1_2_0_U152 ( .A(npu_inst_pe_1_2_0_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_2_0_int_q_reg_v_5__1_), .S(npu_inst_pe_1_2_0_n4), .Z(
        npu_inst_pe_1_2_0_n22) );
  MUX2_X1 npu_inst_pe_1_2_0_U151 ( .A(npu_inst_pe_1_2_0_n21), .B(
        npu_inst_pe_1_2_0_n18), .S(npu_inst_pe_1_2_0_n7), .Z(
        npu_inst_pe_1_2_0_o_data_h_1_) );
  MUX2_X1 npu_inst_pe_1_2_0_U150 ( .A(npu_inst_pe_1_2_0_n20), .B(
        npu_inst_pe_1_2_0_n19), .S(npu_inst_n78), .Z(npu_inst_pe_1_2_0_n21) );
  MUX2_X1 npu_inst_pe_1_2_0_U149 ( .A(npu_inst_pe_1_2_0_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_2_0_int_q_reg_h_1__1_), .S(npu_inst_pe_1_2_0_n4), .Z(
        npu_inst_pe_1_2_0_n20) );
  MUX2_X1 npu_inst_pe_1_2_0_U148 ( .A(npu_inst_pe_1_2_0_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_2_0_int_q_reg_h_3__1_), .S(npu_inst_pe_1_2_0_n4), .Z(
        npu_inst_pe_1_2_0_n19) );
  MUX2_X1 npu_inst_pe_1_2_0_U147 ( .A(npu_inst_pe_1_2_0_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_2_0_int_q_reg_h_5__1_), .S(npu_inst_pe_1_2_0_n4), .Z(
        npu_inst_pe_1_2_0_n18) );
  MUX2_X1 npu_inst_pe_1_2_0_U146 ( .A(npu_inst_pe_1_2_0_n17), .B(
        npu_inst_pe_1_2_0_n14), .S(npu_inst_pe_1_2_0_n7), .Z(
        npu_inst_pe_1_2_0_o_data_h_0_) );
  MUX2_X1 npu_inst_pe_1_2_0_U145 ( .A(npu_inst_pe_1_2_0_n16), .B(
        npu_inst_pe_1_2_0_n15), .S(npu_inst_n78), .Z(npu_inst_pe_1_2_0_n17) );
  MUX2_X1 npu_inst_pe_1_2_0_U144 ( .A(npu_inst_pe_1_2_0_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_2_0_int_q_reg_h_1__0_), .S(npu_inst_pe_1_2_0_n4), .Z(
        npu_inst_pe_1_2_0_n16) );
  MUX2_X1 npu_inst_pe_1_2_0_U143 ( .A(npu_inst_pe_1_2_0_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_2_0_int_q_reg_h_3__0_), .S(npu_inst_pe_1_2_0_n4), .Z(
        npu_inst_pe_1_2_0_n15) );
  MUX2_X1 npu_inst_pe_1_2_0_U142 ( .A(npu_inst_pe_1_2_0_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_2_0_int_q_reg_h_5__0_), .S(npu_inst_pe_1_2_0_n4), .Z(
        npu_inst_pe_1_2_0_n14) );
  XOR2_X1 npu_inst_pe_1_2_0_U141 ( .A(npu_inst_pe_1_2_0_int_data_0_), .B(
        npu_inst_pe_1_2_0_int_q_acc_0_), .Z(npu_inst_pe_1_2_0_N73) );
  AND2_X1 npu_inst_pe_1_2_0_U140 ( .A1(npu_inst_pe_1_2_0_int_q_acc_0_), .A2(
        npu_inst_pe_1_2_0_int_data_0_), .ZN(npu_inst_pe_1_2_0_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_2_0_U139 ( .A(npu_inst_pe_1_2_0_int_q_acc_0_), .B(
        npu_inst_pe_1_2_0_n12), .ZN(npu_inst_pe_1_2_0_N65) );
  OR2_X1 npu_inst_pe_1_2_0_U138 ( .A1(npu_inst_pe_1_2_0_n12), .A2(
        npu_inst_pe_1_2_0_int_q_acc_0_), .ZN(npu_inst_pe_1_2_0_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_2_0_U137 ( .A(npu_inst_pe_1_2_0_int_q_acc_2_), .B(
        npu_inst_pe_1_2_0_add_69_carry_2_), .Z(npu_inst_pe_1_2_0_N75) );
  AND2_X1 npu_inst_pe_1_2_0_U136 ( .A1(npu_inst_pe_1_2_0_add_69_carry_2_), 
        .A2(npu_inst_pe_1_2_0_int_q_acc_2_), .ZN(
        npu_inst_pe_1_2_0_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_2_0_U135 ( .A(npu_inst_pe_1_2_0_int_q_acc_3_), .B(
        npu_inst_pe_1_2_0_add_69_carry_3_), .Z(npu_inst_pe_1_2_0_N76) );
  AND2_X1 npu_inst_pe_1_2_0_U134 ( .A1(npu_inst_pe_1_2_0_add_69_carry_3_), 
        .A2(npu_inst_pe_1_2_0_int_q_acc_3_), .ZN(
        npu_inst_pe_1_2_0_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_2_0_U133 ( .A(npu_inst_pe_1_2_0_int_q_acc_4_), .B(
        npu_inst_pe_1_2_0_add_69_carry_4_), .Z(npu_inst_pe_1_2_0_N77) );
  AND2_X1 npu_inst_pe_1_2_0_U132 ( .A1(npu_inst_pe_1_2_0_add_69_carry_4_), 
        .A2(npu_inst_pe_1_2_0_int_q_acc_4_), .ZN(
        npu_inst_pe_1_2_0_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_2_0_U131 ( .A(npu_inst_pe_1_2_0_int_q_acc_5_), .B(
        npu_inst_pe_1_2_0_add_69_carry_5_), .Z(npu_inst_pe_1_2_0_N78) );
  AND2_X1 npu_inst_pe_1_2_0_U130 ( .A1(npu_inst_pe_1_2_0_add_69_carry_5_), 
        .A2(npu_inst_pe_1_2_0_int_q_acc_5_), .ZN(
        npu_inst_pe_1_2_0_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_2_0_U129 ( .A(npu_inst_pe_1_2_0_int_q_acc_6_), .B(
        npu_inst_pe_1_2_0_add_69_carry_6_), .Z(npu_inst_pe_1_2_0_N79) );
  AND2_X1 npu_inst_pe_1_2_0_U128 ( .A1(npu_inst_pe_1_2_0_add_69_carry_6_), 
        .A2(npu_inst_pe_1_2_0_int_q_acc_6_), .ZN(
        npu_inst_pe_1_2_0_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_2_0_U127 ( .A(npu_inst_pe_1_2_0_int_q_acc_7_), .B(
        npu_inst_pe_1_2_0_add_69_carry_7_), .Z(npu_inst_pe_1_2_0_N80) );
  XNOR2_X1 npu_inst_pe_1_2_0_U126 ( .A(npu_inst_pe_1_2_0_sub_67_carry_2_), .B(
        npu_inst_pe_1_2_0_int_q_acc_2_), .ZN(npu_inst_pe_1_2_0_N67) );
  OR2_X1 npu_inst_pe_1_2_0_U125 ( .A1(npu_inst_pe_1_2_0_int_q_acc_2_), .A2(
        npu_inst_pe_1_2_0_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_2_0_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_2_0_U124 ( .A(npu_inst_pe_1_2_0_sub_67_carry_3_), .B(
        npu_inst_pe_1_2_0_int_q_acc_3_), .ZN(npu_inst_pe_1_2_0_N68) );
  OR2_X1 npu_inst_pe_1_2_0_U123 ( .A1(npu_inst_pe_1_2_0_int_q_acc_3_), .A2(
        npu_inst_pe_1_2_0_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_2_0_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_2_0_U122 ( .A(npu_inst_pe_1_2_0_sub_67_carry_4_), .B(
        npu_inst_pe_1_2_0_int_q_acc_4_), .ZN(npu_inst_pe_1_2_0_N69) );
  OR2_X1 npu_inst_pe_1_2_0_U121 ( .A1(npu_inst_pe_1_2_0_int_q_acc_4_), .A2(
        npu_inst_pe_1_2_0_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_2_0_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_2_0_U120 ( .A(npu_inst_pe_1_2_0_sub_67_carry_5_), .B(
        npu_inst_pe_1_2_0_int_q_acc_5_), .ZN(npu_inst_pe_1_2_0_N70) );
  OR2_X1 npu_inst_pe_1_2_0_U119 ( .A1(npu_inst_pe_1_2_0_int_q_acc_5_), .A2(
        npu_inst_pe_1_2_0_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_2_0_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_2_0_U118 ( .A(npu_inst_pe_1_2_0_sub_67_carry_6_), .B(
        npu_inst_pe_1_2_0_int_q_acc_6_), .ZN(npu_inst_pe_1_2_0_N71) );
  OR2_X1 npu_inst_pe_1_2_0_U117 ( .A1(npu_inst_pe_1_2_0_int_q_acc_6_), .A2(
        npu_inst_pe_1_2_0_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_2_0_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_2_0_U116 ( .A(npu_inst_pe_1_2_0_int_q_acc_7_), .B(
        npu_inst_pe_1_2_0_sub_67_carry_7_), .ZN(npu_inst_pe_1_2_0_N72) );
  INV_X1 npu_inst_pe_1_2_0_U115 ( .A(npu_inst_n78), .ZN(npu_inst_pe_1_2_0_n6)
         );
  INV_X1 npu_inst_pe_1_2_0_U114 ( .A(npu_inst_n58), .ZN(npu_inst_pe_1_2_0_n3)
         );
  AOI22_X1 npu_inst_pe_1_2_0_U113 ( .A1(npu_inst_int_data_y_3__0__0_), .A2(
        npu_inst_pe_1_2_0_n58), .B1(npu_inst_pe_1_2_0_n118), .B2(
        npu_inst_pe_1_2_0_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_2_0_n57) );
  INV_X1 npu_inst_pe_1_2_0_U112 ( .A(npu_inst_pe_1_2_0_n57), .ZN(
        npu_inst_pe_1_2_0_n107) );
  AOI22_X1 npu_inst_pe_1_2_0_U111 ( .A1(npu_inst_int_data_y_3__0__0_), .A2(
        npu_inst_pe_1_2_0_n54), .B1(npu_inst_pe_1_2_0_n117), .B2(
        npu_inst_pe_1_2_0_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_2_0_n53) );
  INV_X1 npu_inst_pe_1_2_0_U110 ( .A(npu_inst_pe_1_2_0_n53), .ZN(
        npu_inst_pe_1_2_0_n108) );
  AOI22_X1 npu_inst_pe_1_2_0_U107 ( .A1(npu_inst_int_data_y_3__0__0_), .A2(
        npu_inst_pe_1_2_0_n50), .B1(npu_inst_pe_1_2_0_n116), .B2(
        npu_inst_pe_1_2_0_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_2_0_n49) );
  INV_X1 npu_inst_pe_1_2_0_U106 ( .A(npu_inst_pe_1_2_0_n49), .ZN(
        npu_inst_pe_1_2_0_n109) );
  AOI22_X1 npu_inst_pe_1_2_0_U105 ( .A1(npu_inst_int_data_y_3__0__0_), .A2(
        npu_inst_pe_1_2_0_n46), .B1(npu_inst_pe_1_2_0_n115), .B2(
        npu_inst_pe_1_2_0_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_2_0_n45) );
  INV_X1 npu_inst_pe_1_2_0_U104 ( .A(npu_inst_pe_1_2_0_n45), .ZN(
        npu_inst_pe_1_2_0_n110) );
  AOI22_X1 npu_inst_pe_1_2_0_U103 ( .A1(npu_inst_int_data_y_3__0__0_), .A2(
        npu_inst_pe_1_2_0_n42), .B1(npu_inst_pe_1_2_0_n114), .B2(
        npu_inst_pe_1_2_0_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_2_0_n41) );
  INV_X1 npu_inst_pe_1_2_0_U102 ( .A(npu_inst_pe_1_2_0_n41), .ZN(
        npu_inst_pe_1_2_0_n111) );
  AOI22_X1 npu_inst_pe_1_2_0_U101 ( .A1(npu_inst_int_data_y_3__0__1_), .A2(
        npu_inst_pe_1_2_0_n58), .B1(npu_inst_pe_1_2_0_n118), .B2(
        npu_inst_pe_1_2_0_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_2_0_n59) );
  INV_X1 npu_inst_pe_1_2_0_U100 ( .A(npu_inst_pe_1_2_0_n59), .ZN(
        npu_inst_pe_1_2_0_n101) );
  AOI22_X1 npu_inst_pe_1_2_0_U99 ( .A1(npu_inst_int_data_y_3__0__1_), .A2(
        npu_inst_pe_1_2_0_n54), .B1(npu_inst_pe_1_2_0_n117), .B2(
        npu_inst_pe_1_2_0_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_2_0_n55) );
  INV_X1 npu_inst_pe_1_2_0_U98 ( .A(npu_inst_pe_1_2_0_n55), .ZN(
        npu_inst_pe_1_2_0_n102) );
  AOI22_X1 npu_inst_pe_1_2_0_U97 ( .A1(npu_inst_int_data_y_3__0__1_), .A2(
        npu_inst_pe_1_2_0_n50), .B1(npu_inst_pe_1_2_0_n116), .B2(
        npu_inst_pe_1_2_0_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_2_0_n51) );
  INV_X1 npu_inst_pe_1_2_0_U96 ( .A(npu_inst_pe_1_2_0_n51), .ZN(
        npu_inst_pe_1_2_0_n103) );
  AOI22_X1 npu_inst_pe_1_2_0_U95 ( .A1(npu_inst_int_data_y_3__0__1_), .A2(
        npu_inst_pe_1_2_0_n46), .B1(npu_inst_pe_1_2_0_n115), .B2(
        npu_inst_pe_1_2_0_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_2_0_n47) );
  INV_X1 npu_inst_pe_1_2_0_U94 ( .A(npu_inst_pe_1_2_0_n47), .ZN(
        npu_inst_pe_1_2_0_n104) );
  AOI22_X1 npu_inst_pe_1_2_0_U93 ( .A1(npu_inst_int_data_y_3__0__1_), .A2(
        npu_inst_pe_1_2_0_n42), .B1(npu_inst_pe_1_2_0_n114), .B2(
        npu_inst_pe_1_2_0_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_2_0_n43) );
  INV_X1 npu_inst_pe_1_2_0_U92 ( .A(npu_inst_pe_1_2_0_n43), .ZN(
        npu_inst_pe_1_2_0_n105) );
  AOI22_X1 npu_inst_pe_1_2_0_U91 ( .A1(npu_inst_pe_1_2_0_n38), .A2(
        npu_inst_int_data_y_3__0__1_), .B1(npu_inst_pe_1_2_0_n113), .B2(
        npu_inst_pe_1_2_0_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_2_0_n39) );
  INV_X1 npu_inst_pe_1_2_0_U90 ( .A(npu_inst_pe_1_2_0_n39), .ZN(
        npu_inst_pe_1_2_0_n106) );
  AOI22_X1 npu_inst_pe_1_2_0_U89 ( .A1(npu_inst_pe_1_2_0_n38), .A2(
        npu_inst_int_data_y_3__0__0_), .B1(npu_inst_pe_1_2_0_n113), .B2(
        npu_inst_pe_1_2_0_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_2_0_n37) );
  INV_X1 npu_inst_pe_1_2_0_U88 ( .A(npu_inst_pe_1_2_0_n37), .ZN(
        npu_inst_pe_1_2_0_n112) );
  NAND2_X1 npu_inst_pe_1_2_0_U87 ( .A1(npu_inst_pe_1_2_0_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_2_0_n60), .ZN(npu_inst_pe_1_2_0_n74) );
  OAI21_X1 npu_inst_pe_1_2_0_U86 ( .B1(npu_inst_pe_1_2_0_n63), .B2(
        npu_inst_pe_1_2_0_n60), .A(npu_inst_pe_1_2_0_n74), .ZN(
        npu_inst_pe_1_2_0_n97) );
  NAND2_X1 npu_inst_pe_1_2_0_U85 ( .A1(npu_inst_pe_1_2_0_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_2_0_n60), .ZN(npu_inst_pe_1_2_0_n73) );
  OAI21_X1 npu_inst_pe_1_2_0_U84 ( .B1(npu_inst_pe_1_2_0_n61), .B2(
        npu_inst_pe_1_2_0_n60), .A(npu_inst_pe_1_2_0_n73), .ZN(
        npu_inst_pe_1_2_0_n96) );
  NAND2_X1 npu_inst_pe_1_2_0_U83 ( .A1(npu_inst_pe_1_2_0_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_2_0_n56), .ZN(npu_inst_pe_1_2_0_n72) );
  OAI21_X1 npu_inst_pe_1_2_0_U82 ( .B1(npu_inst_pe_1_2_0_n63), .B2(
        npu_inst_pe_1_2_0_n56), .A(npu_inst_pe_1_2_0_n72), .ZN(
        npu_inst_pe_1_2_0_n95) );
  NAND2_X1 npu_inst_pe_1_2_0_U81 ( .A1(npu_inst_pe_1_2_0_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_2_0_n56), .ZN(npu_inst_pe_1_2_0_n71) );
  OAI21_X1 npu_inst_pe_1_2_0_U80 ( .B1(npu_inst_pe_1_2_0_n61), .B2(
        npu_inst_pe_1_2_0_n56), .A(npu_inst_pe_1_2_0_n71), .ZN(
        npu_inst_pe_1_2_0_n94) );
  NAND2_X1 npu_inst_pe_1_2_0_U79 ( .A1(npu_inst_pe_1_2_0_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_2_0_n52), .ZN(npu_inst_pe_1_2_0_n70) );
  OAI21_X1 npu_inst_pe_1_2_0_U78 ( .B1(npu_inst_pe_1_2_0_n63), .B2(
        npu_inst_pe_1_2_0_n52), .A(npu_inst_pe_1_2_0_n70), .ZN(
        npu_inst_pe_1_2_0_n93) );
  NAND2_X1 npu_inst_pe_1_2_0_U77 ( .A1(npu_inst_pe_1_2_0_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_2_0_n52), .ZN(npu_inst_pe_1_2_0_n69) );
  OAI21_X1 npu_inst_pe_1_2_0_U76 ( .B1(npu_inst_pe_1_2_0_n61), .B2(
        npu_inst_pe_1_2_0_n52), .A(npu_inst_pe_1_2_0_n69), .ZN(
        npu_inst_pe_1_2_0_n92) );
  NAND2_X1 npu_inst_pe_1_2_0_U75 ( .A1(npu_inst_pe_1_2_0_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_2_0_n48), .ZN(npu_inst_pe_1_2_0_n68) );
  OAI21_X1 npu_inst_pe_1_2_0_U74 ( .B1(npu_inst_pe_1_2_0_n63), .B2(
        npu_inst_pe_1_2_0_n48), .A(npu_inst_pe_1_2_0_n68), .ZN(
        npu_inst_pe_1_2_0_n91) );
  NAND2_X1 npu_inst_pe_1_2_0_U73 ( .A1(npu_inst_pe_1_2_0_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_2_0_n48), .ZN(npu_inst_pe_1_2_0_n67) );
  OAI21_X1 npu_inst_pe_1_2_0_U72 ( .B1(npu_inst_pe_1_2_0_n61), .B2(
        npu_inst_pe_1_2_0_n48), .A(npu_inst_pe_1_2_0_n67), .ZN(
        npu_inst_pe_1_2_0_n90) );
  NAND2_X1 npu_inst_pe_1_2_0_U71 ( .A1(npu_inst_pe_1_2_0_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_2_0_n44), .ZN(npu_inst_pe_1_2_0_n66) );
  OAI21_X1 npu_inst_pe_1_2_0_U70 ( .B1(npu_inst_pe_1_2_0_n63), .B2(
        npu_inst_pe_1_2_0_n44), .A(npu_inst_pe_1_2_0_n66), .ZN(
        npu_inst_pe_1_2_0_n89) );
  NAND2_X1 npu_inst_pe_1_2_0_U69 ( .A1(npu_inst_pe_1_2_0_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_2_0_n44), .ZN(npu_inst_pe_1_2_0_n65) );
  OAI21_X1 npu_inst_pe_1_2_0_U68 ( .B1(npu_inst_pe_1_2_0_n61), .B2(
        npu_inst_pe_1_2_0_n44), .A(npu_inst_pe_1_2_0_n65), .ZN(
        npu_inst_pe_1_2_0_n88) );
  NAND2_X1 npu_inst_pe_1_2_0_U67 ( .A1(npu_inst_pe_1_2_0_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_2_0_n40), .ZN(npu_inst_pe_1_2_0_n64) );
  OAI21_X1 npu_inst_pe_1_2_0_U66 ( .B1(npu_inst_pe_1_2_0_n63), .B2(
        npu_inst_pe_1_2_0_n40), .A(npu_inst_pe_1_2_0_n64), .ZN(
        npu_inst_pe_1_2_0_n87) );
  NAND2_X1 npu_inst_pe_1_2_0_U65 ( .A1(npu_inst_pe_1_2_0_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_2_0_n40), .ZN(npu_inst_pe_1_2_0_n62) );
  OAI21_X1 npu_inst_pe_1_2_0_U64 ( .B1(npu_inst_pe_1_2_0_n61), .B2(
        npu_inst_pe_1_2_0_n40), .A(npu_inst_pe_1_2_0_n62), .ZN(
        npu_inst_pe_1_2_0_n86) );
  AND2_X1 npu_inst_pe_1_2_0_U63 ( .A1(npu_inst_pe_1_2_0_N93), .A2(npu_inst_n58), .ZN(npu_inst_int_data_y_2__0__0_) );
  AND2_X1 npu_inst_pe_1_2_0_U62 ( .A1(npu_inst_n58), .A2(npu_inst_pe_1_2_0_N94), .ZN(npu_inst_int_data_y_2__0__1_) );
  NOR3_X1 npu_inst_pe_1_2_0_U61 ( .A1(npu_inst_pe_1_2_0_n26), .A2(npu_inst_n58), .A3(npu_inst_int_ckg[47]), .ZN(npu_inst_pe_1_2_0_n85) );
  OR2_X1 npu_inst_pe_1_2_0_U60 ( .A1(npu_inst_pe_1_2_0_n85), .A2(
        npu_inst_pe_1_2_0_n2), .ZN(npu_inst_pe_1_2_0_N84) );
  AND2_X1 npu_inst_pe_1_2_0_U59 ( .A1(npu_inst_pe_1_2_0_int_q_acc_0_), .A2(
        npu_inst_pe_1_2_0_n1), .ZN(npu_inst_int_data_res_2__0__0_) );
  AND2_X1 npu_inst_pe_1_2_0_U58 ( .A1(npu_inst_pe_1_2_0_n2), .A2(
        npu_inst_pe_1_2_0_int_q_acc_7_), .ZN(npu_inst_int_data_res_2__0__7_)
         );
  AND2_X1 npu_inst_pe_1_2_0_U57 ( .A1(npu_inst_pe_1_2_0_int_q_acc_1_), .A2(
        npu_inst_pe_1_2_0_n1), .ZN(npu_inst_int_data_res_2__0__1_) );
  AND2_X1 npu_inst_pe_1_2_0_U56 ( .A1(npu_inst_pe_1_2_0_int_q_acc_2_), .A2(
        npu_inst_pe_1_2_0_n1), .ZN(npu_inst_int_data_res_2__0__2_) );
  AND2_X1 npu_inst_pe_1_2_0_U55 ( .A1(npu_inst_pe_1_2_0_int_q_acc_3_), .A2(
        npu_inst_pe_1_2_0_n2), .ZN(npu_inst_int_data_res_2__0__3_) );
  AND2_X1 npu_inst_pe_1_2_0_U54 ( .A1(npu_inst_pe_1_2_0_int_q_acc_4_), .A2(
        npu_inst_pe_1_2_0_n2), .ZN(npu_inst_int_data_res_2__0__4_) );
  AND2_X1 npu_inst_pe_1_2_0_U53 ( .A1(npu_inst_pe_1_2_0_int_q_acc_5_), .A2(
        npu_inst_pe_1_2_0_n2), .ZN(npu_inst_int_data_res_2__0__5_) );
  AND2_X1 npu_inst_pe_1_2_0_U52 ( .A1(npu_inst_pe_1_2_0_int_q_acc_6_), .A2(
        npu_inst_pe_1_2_0_n2), .ZN(npu_inst_int_data_res_2__0__6_) );
  AOI222_X1 npu_inst_pe_1_2_0_U51 ( .A1(npu_inst_int_data_res_3__0__0_), .A2(
        npu_inst_pe_1_2_0_n1), .B1(npu_inst_pe_1_2_0_N73), .B2(
        npu_inst_pe_1_2_0_n76), .C1(npu_inst_pe_1_2_0_N65), .C2(
        npu_inst_pe_1_2_0_n77), .ZN(npu_inst_pe_1_2_0_n84) );
  INV_X1 npu_inst_pe_1_2_0_U50 ( .A(npu_inst_pe_1_2_0_n84), .ZN(
        npu_inst_pe_1_2_0_n100) );
  AOI222_X1 npu_inst_pe_1_2_0_U49 ( .A1(npu_inst_int_data_res_3__0__7_), .A2(
        npu_inst_pe_1_2_0_n1), .B1(npu_inst_pe_1_2_0_N80), .B2(
        npu_inst_pe_1_2_0_n76), .C1(npu_inst_pe_1_2_0_N72), .C2(
        npu_inst_pe_1_2_0_n77), .ZN(npu_inst_pe_1_2_0_n75) );
  INV_X1 npu_inst_pe_1_2_0_U48 ( .A(npu_inst_pe_1_2_0_n75), .ZN(
        npu_inst_pe_1_2_0_n32) );
  AOI222_X1 npu_inst_pe_1_2_0_U47 ( .A1(npu_inst_int_data_res_3__0__1_), .A2(
        npu_inst_pe_1_2_0_n1), .B1(npu_inst_pe_1_2_0_N74), .B2(
        npu_inst_pe_1_2_0_n76), .C1(npu_inst_pe_1_2_0_N66), .C2(
        npu_inst_pe_1_2_0_n77), .ZN(npu_inst_pe_1_2_0_n83) );
  INV_X1 npu_inst_pe_1_2_0_U46 ( .A(npu_inst_pe_1_2_0_n83), .ZN(
        npu_inst_pe_1_2_0_n99) );
  AOI222_X1 npu_inst_pe_1_2_0_U45 ( .A1(npu_inst_int_data_res_3__0__2_), .A2(
        npu_inst_pe_1_2_0_n1), .B1(npu_inst_pe_1_2_0_N75), .B2(
        npu_inst_pe_1_2_0_n76), .C1(npu_inst_pe_1_2_0_N67), .C2(
        npu_inst_pe_1_2_0_n77), .ZN(npu_inst_pe_1_2_0_n82) );
  INV_X1 npu_inst_pe_1_2_0_U44 ( .A(npu_inst_pe_1_2_0_n82), .ZN(
        npu_inst_pe_1_2_0_n98) );
  AOI222_X1 npu_inst_pe_1_2_0_U43 ( .A1(npu_inst_int_data_res_3__0__3_), .A2(
        npu_inst_pe_1_2_0_n1), .B1(npu_inst_pe_1_2_0_N76), .B2(
        npu_inst_pe_1_2_0_n76), .C1(npu_inst_pe_1_2_0_N68), .C2(
        npu_inst_pe_1_2_0_n77), .ZN(npu_inst_pe_1_2_0_n81) );
  INV_X1 npu_inst_pe_1_2_0_U42 ( .A(npu_inst_pe_1_2_0_n81), .ZN(
        npu_inst_pe_1_2_0_n36) );
  AOI222_X1 npu_inst_pe_1_2_0_U41 ( .A1(npu_inst_int_data_res_3__0__4_), .A2(
        npu_inst_pe_1_2_0_n1), .B1(npu_inst_pe_1_2_0_N77), .B2(
        npu_inst_pe_1_2_0_n76), .C1(npu_inst_pe_1_2_0_N69), .C2(
        npu_inst_pe_1_2_0_n77), .ZN(npu_inst_pe_1_2_0_n80) );
  INV_X1 npu_inst_pe_1_2_0_U40 ( .A(npu_inst_pe_1_2_0_n80), .ZN(
        npu_inst_pe_1_2_0_n35) );
  AOI222_X1 npu_inst_pe_1_2_0_U39 ( .A1(npu_inst_int_data_res_3__0__5_), .A2(
        npu_inst_pe_1_2_0_n1), .B1(npu_inst_pe_1_2_0_N78), .B2(
        npu_inst_pe_1_2_0_n76), .C1(npu_inst_pe_1_2_0_N70), .C2(
        npu_inst_pe_1_2_0_n77), .ZN(npu_inst_pe_1_2_0_n79) );
  INV_X1 npu_inst_pe_1_2_0_U38 ( .A(npu_inst_pe_1_2_0_n79), .ZN(
        npu_inst_pe_1_2_0_n34) );
  AOI222_X1 npu_inst_pe_1_2_0_U37 ( .A1(npu_inst_int_data_res_3__0__6_), .A2(
        npu_inst_pe_1_2_0_n1), .B1(npu_inst_pe_1_2_0_N79), .B2(
        npu_inst_pe_1_2_0_n76), .C1(npu_inst_pe_1_2_0_N71), .C2(
        npu_inst_pe_1_2_0_n77), .ZN(npu_inst_pe_1_2_0_n78) );
  INV_X1 npu_inst_pe_1_2_0_U36 ( .A(npu_inst_pe_1_2_0_n78), .ZN(
        npu_inst_pe_1_2_0_n33) );
  AND2_X1 npu_inst_pe_1_2_0_U35 ( .A1(npu_inst_pe_1_2_0_o_data_h_1_), .A2(
        npu_inst_pe_1_2_0_int_q_weight_1_), .ZN(npu_inst_pe_1_2_0_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_2_0_U34 ( .A1(npu_inst_pe_1_2_0_o_data_h_0_), .A2(
        npu_inst_pe_1_2_0_int_q_weight_1_), .ZN(npu_inst_pe_1_2_0_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_2_0_U33 ( .A(npu_inst_pe_1_2_0_int_data_1_), .ZN(
        npu_inst_pe_1_2_0_n13) );
  AOI22_X1 npu_inst_pe_1_2_0_U32 ( .A1(npu_inst_n58), .A2(
        npu_inst_int_data_y_3__0__1_), .B1(npu_inst_pe_1_2_0_n3), .B2(
        npu_inst_int_data_x_2__1__1_), .ZN(npu_inst_pe_1_2_0_n63) );
  AOI22_X1 npu_inst_pe_1_2_0_U31 ( .A1(npu_inst_n58), .A2(
        npu_inst_int_data_y_3__0__0_), .B1(npu_inst_pe_1_2_0_n3), .B2(
        npu_inst_int_data_x_2__1__0_), .ZN(npu_inst_pe_1_2_0_n61) );
  INV_X1 npu_inst_pe_1_2_0_U30 ( .A(npu_inst_pe_1_2_0_int_data_0_), .ZN(
        npu_inst_pe_1_2_0_n12) );
  INV_X1 npu_inst_pe_1_2_0_U29 ( .A(npu_inst_n70), .ZN(npu_inst_pe_1_2_0_n5)
         );
  OR3_X1 npu_inst_pe_1_2_0_U28 ( .A1(npu_inst_n78), .A2(npu_inst_pe_1_2_0_n7), 
        .A3(npu_inst_pe_1_2_0_n5), .ZN(npu_inst_pe_1_2_0_n56) );
  OR3_X1 npu_inst_pe_1_2_0_U27 ( .A1(npu_inst_pe_1_2_0_n5), .A2(
        npu_inst_pe_1_2_0_n7), .A3(npu_inst_pe_1_2_0_n6), .ZN(
        npu_inst_pe_1_2_0_n48) );
  INV_X1 npu_inst_pe_1_2_0_U26 ( .A(npu_inst_pe_1_2_0_n5), .ZN(
        npu_inst_pe_1_2_0_n4) );
  OR3_X1 npu_inst_pe_1_2_0_U25 ( .A1(npu_inst_pe_1_2_0_n4), .A2(
        npu_inst_pe_1_2_0_n7), .A3(npu_inst_pe_1_2_0_n6), .ZN(
        npu_inst_pe_1_2_0_n52) );
  OR3_X1 npu_inst_pe_1_2_0_U24 ( .A1(npu_inst_n78), .A2(npu_inst_pe_1_2_0_n7), 
        .A3(npu_inst_pe_1_2_0_n4), .ZN(npu_inst_pe_1_2_0_n60) );
  NOR2_X1 npu_inst_pe_1_2_0_U23 ( .A1(npu_inst_pe_1_2_0_n60), .A2(
        npu_inst_pe_1_2_0_n3), .ZN(npu_inst_pe_1_2_0_n58) );
  NOR2_X1 npu_inst_pe_1_2_0_U22 ( .A1(npu_inst_pe_1_2_0_n56), .A2(
        npu_inst_pe_1_2_0_n3), .ZN(npu_inst_pe_1_2_0_n54) );
  NOR2_X1 npu_inst_pe_1_2_0_U21 ( .A1(npu_inst_pe_1_2_0_n52), .A2(
        npu_inst_pe_1_2_0_n3), .ZN(npu_inst_pe_1_2_0_n50) );
  NOR2_X1 npu_inst_pe_1_2_0_U20 ( .A1(npu_inst_pe_1_2_0_n48), .A2(
        npu_inst_pe_1_2_0_n3), .ZN(npu_inst_pe_1_2_0_n46) );
  NOR2_X1 npu_inst_pe_1_2_0_U19 ( .A1(npu_inst_pe_1_2_0_n40), .A2(
        npu_inst_pe_1_2_0_n3), .ZN(npu_inst_pe_1_2_0_n38) );
  NOR2_X1 npu_inst_pe_1_2_0_U18 ( .A1(npu_inst_pe_1_2_0_n44), .A2(
        npu_inst_pe_1_2_0_n3), .ZN(npu_inst_pe_1_2_0_n42) );
  BUF_X1 npu_inst_pe_1_2_0_U17 ( .A(npu_inst_n103), .Z(npu_inst_pe_1_2_0_n7)
         );
  INV_X1 npu_inst_pe_1_2_0_U16 ( .A(npu_inst_n125), .ZN(npu_inst_pe_1_2_0_n11)
         );
  INV_X1 npu_inst_pe_1_2_0_U15 ( .A(npu_inst_pe_1_2_0_n38), .ZN(
        npu_inst_pe_1_2_0_n113) );
  INV_X1 npu_inst_pe_1_2_0_U14 ( .A(npu_inst_pe_1_2_0_n58), .ZN(
        npu_inst_pe_1_2_0_n118) );
  INV_X1 npu_inst_pe_1_2_0_U13 ( .A(npu_inst_pe_1_2_0_n54), .ZN(
        npu_inst_pe_1_2_0_n117) );
  INV_X1 npu_inst_pe_1_2_0_U12 ( .A(npu_inst_pe_1_2_0_n50), .ZN(
        npu_inst_pe_1_2_0_n116) );
  INV_X1 npu_inst_pe_1_2_0_U11 ( .A(npu_inst_pe_1_2_0_n46), .ZN(
        npu_inst_pe_1_2_0_n115) );
  INV_X1 npu_inst_pe_1_2_0_U10 ( .A(npu_inst_pe_1_2_0_n42), .ZN(
        npu_inst_pe_1_2_0_n114) );
  BUF_X1 npu_inst_pe_1_2_0_U9 ( .A(npu_inst_n30), .Z(npu_inst_pe_1_2_0_n2) );
  BUF_X1 npu_inst_pe_1_2_0_U8 ( .A(npu_inst_n30), .Z(npu_inst_pe_1_2_0_n1) );
  BUF_X1 npu_inst_pe_1_2_0_U7 ( .A(npu_inst_pe_1_2_0_n11), .Z(
        npu_inst_pe_1_2_0_n10) );
  BUF_X1 npu_inst_pe_1_2_0_U6 ( .A(npu_inst_pe_1_2_0_n11), .Z(
        npu_inst_pe_1_2_0_n9) );
  BUF_X1 npu_inst_pe_1_2_0_U5 ( .A(npu_inst_pe_1_2_0_n11), .Z(
        npu_inst_pe_1_2_0_n8) );
  NOR2_X1 npu_inst_pe_1_2_0_U4 ( .A1(npu_inst_pe_1_2_0_int_q_weight_0_), .A2(
        npu_inst_pe_1_2_0_n1), .ZN(npu_inst_pe_1_2_0_n76) );
  NOR2_X1 npu_inst_pe_1_2_0_U3 ( .A1(npu_inst_pe_1_2_0_n27), .A2(
        npu_inst_pe_1_2_0_n1), .ZN(npu_inst_pe_1_2_0_n77) );
  FA_X1 npu_inst_pe_1_2_0_sub_67_U2_1 ( .A(npu_inst_pe_1_2_0_int_q_acc_1_), 
        .B(npu_inst_pe_1_2_0_n13), .CI(npu_inst_pe_1_2_0_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_2_0_sub_67_carry_2_), .S(npu_inst_pe_1_2_0_N66) );
  FA_X1 npu_inst_pe_1_2_0_add_69_U1_1 ( .A(npu_inst_pe_1_2_0_int_q_acc_1_), 
        .B(npu_inst_pe_1_2_0_int_data_1_), .CI(
        npu_inst_pe_1_2_0_add_69_carry_1_), .CO(
        npu_inst_pe_1_2_0_add_69_carry_2_), .S(npu_inst_pe_1_2_0_N74) );
  NAND3_X1 npu_inst_pe_1_2_0_U109 ( .A1(npu_inst_pe_1_2_0_n5), .A2(
        npu_inst_pe_1_2_0_n6), .A3(npu_inst_pe_1_2_0_n7), .ZN(
        npu_inst_pe_1_2_0_n44) );
  NAND3_X1 npu_inst_pe_1_2_0_U108 ( .A1(npu_inst_pe_1_2_0_n4), .A2(
        npu_inst_pe_1_2_0_n6), .A3(npu_inst_pe_1_2_0_n7), .ZN(
        npu_inst_pe_1_2_0_n40) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_2_0_n33), .CK(
        npu_inst_pe_1_2_0_net4194), .RN(npu_inst_pe_1_2_0_n8), .Q(
        npu_inst_pe_1_2_0_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_2_0_n34), .CK(
        npu_inst_pe_1_2_0_net4194), .RN(npu_inst_pe_1_2_0_n8), .Q(
        npu_inst_pe_1_2_0_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_2_0_n35), .CK(
        npu_inst_pe_1_2_0_net4194), .RN(npu_inst_pe_1_2_0_n8), .Q(
        npu_inst_pe_1_2_0_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_2_0_n36), .CK(
        npu_inst_pe_1_2_0_net4194), .RN(npu_inst_pe_1_2_0_n8), .Q(
        npu_inst_pe_1_2_0_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_2_0_n98), .CK(
        npu_inst_pe_1_2_0_net4194), .RN(npu_inst_pe_1_2_0_n8), .Q(
        npu_inst_pe_1_2_0_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_2_0_n99), .CK(
        npu_inst_pe_1_2_0_net4194), .RN(npu_inst_pe_1_2_0_n8), .Q(
        npu_inst_pe_1_2_0_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_2_0_n32), .CK(
        npu_inst_pe_1_2_0_net4194), .RN(npu_inst_pe_1_2_0_n8), .Q(
        npu_inst_pe_1_2_0_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_2_0_n100), 
        .CK(npu_inst_pe_1_2_0_net4194), .RN(npu_inst_pe_1_2_0_n8), .Q(
        npu_inst_pe_1_2_0_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_weight_reg_0_ ( .D(npu_inst_n111), .CK(
        npu_inst_pe_1_2_0_net4200), .RN(npu_inst_pe_1_2_0_n8), .Q(
        npu_inst_pe_1_2_0_int_q_weight_0_), .QN(npu_inst_pe_1_2_0_n27) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_weight_reg_1_ ( .D(npu_inst_n117), .CK(
        npu_inst_pe_1_2_0_net4200), .RN(npu_inst_pe_1_2_0_n8), .Q(
        npu_inst_pe_1_2_0_int_q_weight_1_), .QN(npu_inst_pe_1_2_0_n26) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_2_0_n112), 
        .CK(npu_inst_pe_1_2_0_net4200), .RN(npu_inst_pe_1_2_0_n8), .Q(
        npu_inst_pe_1_2_0_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_2_0_n106), 
        .CK(npu_inst_pe_1_2_0_net4200), .RN(npu_inst_pe_1_2_0_n8), .Q(
        npu_inst_pe_1_2_0_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_2_0_n111), 
        .CK(npu_inst_pe_1_2_0_net4200), .RN(npu_inst_pe_1_2_0_n9), .Q(
        npu_inst_pe_1_2_0_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_2_0_n105), 
        .CK(npu_inst_pe_1_2_0_net4200), .RN(npu_inst_pe_1_2_0_n9), .Q(
        npu_inst_pe_1_2_0_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_2_0_n110), 
        .CK(npu_inst_pe_1_2_0_net4200), .RN(npu_inst_pe_1_2_0_n9), .Q(
        npu_inst_pe_1_2_0_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_2_0_n104), 
        .CK(npu_inst_pe_1_2_0_net4200), .RN(npu_inst_pe_1_2_0_n9), .Q(
        npu_inst_pe_1_2_0_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_2_0_n109), 
        .CK(npu_inst_pe_1_2_0_net4200), .RN(npu_inst_pe_1_2_0_n9), .Q(
        npu_inst_pe_1_2_0_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_2_0_n103), 
        .CK(npu_inst_pe_1_2_0_net4200), .RN(npu_inst_pe_1_2_0_n9), .Q(
        npu_inst_pe_1_2_0_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_2_0_n108), 
        .CK(npu_inst_pe_1_2_0_net4200), .RN(npu_inst_pe_1_2_0_n9), .Q(
        npu_inst_pe_1_2_0_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_2_0_n102), 
        .CK(npu_inst_pe_1_2_0_net4200), .RN(npu_inst_pe_1_2_0_n9), .Q(
        npu_inst_pe_1_2_0_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_2_0_n107), 
        .CK(npu_inst_pe_1_2_0_net4200), .RN(npu_inst_pe_1_2_0_n9), .Q(
        npu_inst_pe_1_2_0_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_2_0_n101), 
        .CK(npu_inst_pe_1_2_0_net4200), .RN(npu_inst_pe_1_2_0_n9), .Q(
        npu_inst_pe_1_2_0_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_2_0_n86), 
        .CK(npu_inst_pe_1_2_0_net4200), .RN(npu_inst_pe_1_2_0_n9), .Q(
        npu_inst_pe_1_2_0_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_2_0_n87), 
        .CK(npu_inst_pe_1_2_0_net4200), .RN(npu_inst_pe_1_2_0_n9), .Q(
        npu_inst_pe_1_2_0_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_2_0_n88), 
        .CK(npu_inst_pe_1_2_0_net4200), .RN(npu_inst_pe_1_2_0_n10), .Q(
        npu_inst_pe_1_2_0_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_2_0_n89), 
        .CK(npu_inst_pe_1_2_0_net4200), .RN(npu_inst_pe_1_2_0_n10), .Q(
        npu_inst_pe_1_2_0_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_2_0_n90), 
        .CK(npu_inst_pe_1_2_0_net4200), .RN(npu_inst_pe_1_2_0_n10), .Q(
        npu_inst_pe_1_2_0_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_2_0_n91), 
        .CK(npu_inst_pe_1_2_0_net4200), .RN(npu_inst_pe_1_2_0_n10), .Q(
        npu_inst_pe_1_2_0_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_2_0_n92), 
        .CK(npu_inst_pe_1_2_0_net4200), .RN(npu_inst_pe_1_2_0_n10), .Q(
        npu_inst_pe_1_2_0_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_2_0_n93), 
        .CK(npu_inst_pe_1_2_0_net4200), .RN(npu_inst_pe_1_2_0_n10), .Q(
        npu_inst_pe_1_2_0_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_2_0_n94), 
        .CK(npu_inst_pe_1_2_0_net4200), .RN(npu_inst_pe_1_2_0_n10), .Q(
        npu_inst_pe_1_2_0_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_2_0_n95), 
        .CK(npu_inst_pe_1_2_0_net4200), .RN(npu_inst_pe_1_2_0_n10), .Q(
        npu_inst_pe_1_2_0_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_2_0_n96), 
        .CK(npu_inst_pe_1_2_0_net4200), .RN(npu_inst_pe_1_2_0_n10), .Q(
        npu_inst_pe_1_2_0_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_2_0_n97), 
        .CK(npu_inst_pe_1_2_0_net4200), .RN(npu_inst_pe_1_2_0_n10), .Q(
        npu_inst_pe_1_2_0_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_2_0_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_2_0_N84), .SE(1'b0), .GCK(npu_inst_pe_1_2_0_net4194) );
  CLKGATETST_X1 npu_inst_pe_1_2_0_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n65), .SE(1'b0), .GCK(npu_inst_pe_1_2_0_net4200) );
  MUX2_X1 npu_inst_pe_1_2_1_U162 ( .A(npu_inst_pe_1_2_1_n32), .B(
        npu_inst_pe_1_2_1_n29), .S(npu_inst_pe_1_2_1_n8), .Z(
        npu_inst_pe_1_2_1_N93) );
  MUX2_X1 npu_inst_pe_1_2_1_U161 ( .A(npu_inst_pe_1_2_1_n31), .B(
        npu_inst_pe_1_2_1_n30), .S(npu_inst_pe_1_2_1_n6), .Z(
        npu_inst_pe_1_2_1_n32) );
  MUX2_X1 npu_inst_pe_1_2_1_U160 ( .A(npu_inst_pe_1_2_1_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_2_1_int_q_reg_v_1__0_), .S(npu_inst_pe_1_2_1_n4), .Z(
        npu_inst_pe_1_2_1_n31) );
  MUX2_X1 npu_inst_pe_1_2_1_U159 ( .A(npu_inst_pe_1_2_1_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_2_1_int_q_reg_v_3__0_), .S(npu_inst_pe_1_2_1_n4), .Z(
        npu_inst_pe_1_2_1_n30) );
  MUX2_X1 npu_inst_pe_1_2_1_U158 ( .A(npu_inst_pe_1_2_1_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_2_1_int_q_reg_v_5__0_), .S(npu_inst_pe_1_2_1_n4), .Z(
        npu_inst_pe_1_2_1_n29) );
  MUX2_X1 npu_inst_pe_1_2_1_U157 ( .A(npu_inst_pe_1_2_1_n28), .B(
        npu_inst_pe_1_2_1_n23), .S(npu_inst_pe_1_2_1_n8), .Z(
        npu_inst_pe_1_2_1_N94) );
  MUX2_X1 npu_inst_pe_1_2_1_U156 ( .A(npu_inst_pe_1_2_1_n25), .B(
        npu_inst_pe_1_2_1_n24), .S(npu_inst_pe_1_2_1_n6), .Z(
        npu_inst_pe_1_2_1_n28) );
  MUX2_X1 npu_inst_pe_1_2_1_U155 ( .A(npu_inst_pe_1_2_1_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_2_1_int_q_reg_v_1__1_), .S(npu_inst_pe_1_2_1_n4), .Z(
        npu_inst_pe_1_2_1_n25) );
  MUX2_X1 npu_inst_pe_1_2_1_U154 ( .A(npu_inst_pe_1_2_1_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_2_1_int_q_reg_v_3__1_), .S(npu_inst_pe_1_2_1_n4), .Z(
        npu_inst_pe_1_2_1_n24) );
  MUX2_X1 npu_inst_pe_1_2_1_U153 ( .A(npu_inst_pe_1_2_1_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_2_1_int_q_reg_v_5__1_), .S(npu_inst_pe_1_2_1_n4), .Z(
        npu_inst_pe_1_2_1_n23) );
  MUX2_X1 npu_inst_pe_1_2_1_U152 ( .A(npu_inst_pe_1_2_1_n22), .B(
        npu_inst_pe_1_2_1_n19), .S(npu_inst_pe_1_2_1_n8), .Z(
        npu_inst_int_data_x_2__1__1_) );
  MUX2_X1 npu_inst_pe_1_2_1_U151 ( .A(npu_inst_pe_1_2_1_n21), .B(
        npu_inst_pe_1_2_1_n20), .S(npu_inst_pe_1_2_1_n6), .Z(
        npu_inst_pe_1_2_1_n22) );
  MUX2_X1 npu_inst_pe_1_2_1_U150 ( .A(npu_inst_pe_1_2_1_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_2_1_int_q_reg_h_1__1_), .S(npu_inst_pe_1_2_1_n4), .Z(
        npu_inst_pe_1_2_1_n21) );
  MUX2_X1 npu_inst_pe_1_2_1_U149 ( .A(npu_inst_pe_1_2_1_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_2_1_int_q_reg_h_3__1_), .S(npu_inst_pe_1_2_1_n4), .Z(
        npu_inst_pe_1_2_1_n20) );
  MUX2_X1 npu_inst_pe_1_2_1_U148 ( .A(npu_inst_pe_1_2_1_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_2_1_int_q_reg_h_5__1_), .S(npu_inst_pe_1_2_1_n4), .Z(
        npu_inst_pe_1_2_1_n19) );
  MUX2_X1 npu_inst_pe_1_2_1_U147 ( .A(npu_inst_pe_1_2_1_n18), .B(
        npu_inst_pe_1_2_1_n15), .S(npu_inst_pe_1_2_1_n8), .Z(
        npu_inst_int_data_x_2__1__0_) );
  MUX2_X1 npu_inst_pe_1_2_1_U146 ( .A(npu_inst_pe_1_2_1_n17), .B(
        npu_inst_pe_1_2_1_n16), .S(npu_inst_pe_1_2_1_n6), .Z(
        npu_inst_pe_1_2_1_n18) );
  MUX2_X1 npu_inst_pe_1_2_1_U145 ( .A(npu_inst_pe_1_2_1_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_2_1_int_q_reg_h_1__0_), .S(npu_inst_pe_1_2_1_n4), .Z(
        npu_inst_pe_1_2_1_n17) );
  MUX2_X1 npu_inst_pe_1_2_1_U144 ( .A(npu_inst_pe_1_2_1_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_2_1_int_q_reg_h_3__0_), .S(npu_inst_pe_1_2_1_n4), .Z(
        npu_inst_pe_1_2_1_n16) );
  MUX2_X1 npu_inst_pe_1_2_1_U143 ( .A(npu_inst_pe_1_2_1_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_2_1_int_q_reg_h_5__0_), .S(npu_inst_pe_1_2_1_n4), .Z(
        npu_inst_pe_1_2_1_n15) );
  XOR2_X1 npu_inst_pe_1_2_1_U142 ( .A(npu_inst_pe_1_2_1_int_data_0_), .B(
        npu_inst_pe_1_2_1_int_q_acc_0_), .Z(npu_inst_pe_1_2_1_N73) );
  AND2_X1 npu_inst_pe_1_2_1_U141 ( .A1(npu_inst_pe_1_2_1_int_q_acc_0_), .A2(
        npu_inst_pe_1_2_1_int_data_0_), .ZN(npu_inst_pe_1_2_1_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_2_1_U140 ( .A(npu_inst_pe_1_2_1_int_q_acc_0_), .B(
        npu_inst_pe_1_2_1_n13), .ZN(npu_inst_pe_1_2_1_N65) );
  OR2_X1 npu_inst_pe_1_2_1_U139 ( .A1(npu_inst_pe_1_2_1_n13), .A2(
        npu_inst_pe_1_2_1_int_q_acc_0_), .ZN(npu_inst_pe_1_2_1_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_2_1_U138 ( .A(npu_inst_pe_1_2_1_int_q_acc_2_), .B(
        npu_inst_pe_1_2_1_add_69_carry_2_), .Z(npu_inst_pe_1_2_1_N75) );
  AND2_X1 npu_inst_pe_1_2_1_U137 ( .A1(npu_inst_pe_1_2_1_add_69_carry_2_), 
        .A2(npu_inst_pe_1_2_1_int_q_acc_2_), .ZN(
        npu_inst_pe_1_2_1_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_2_1_U136 ( .A(npu_inst_pe_1_2_1_int_q_acc_3_), .B(
        npu_inst_pe_1_2_1_add_69_carry_3_), .Z(npu_inst_pe_1_2_1_N76) );
  AND2_X1 npu_inst_pe_1_2_1_U135 ( .A1(npu_inst_pe_1_2_1_add_69_carry_3_), 
        .A2(npu_inst_pe_1_2_1_int_q_acc_3_), .ZN(
        npu_inst_pe_1_2_1_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_2_1_U134 ( .A(npu_inst_pe_1_2_1_int_q_acc_4_), .B(
        npu_inst_pe_1_2_1_add_69_carry_4_), .Z(npu_inst_pe_1_2_1_N77) );
  AND2_X1 npu_inst_pe_1_2_1_U133 ( .A1(npu_inst_pe_1_2_1_add_69_carry_4_), 
        .A2(npu_inst_pe_1_2_1_int_q_acc_4_), .ZN(
        npu_inst_pe_1_2_1_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_2_1_U132 ( .A(npu_inst_pe_1_2_1_int_q_acc_5_), .B(
        npu_inst_pe_1_2_1_add_69_carry_5_), .Z(npu_inst_pe_1_2_1_N78) );
  AND2_X1 npu_inst_pe_1_2_1_U131 ( .A1(npu_inst_pe_1_2_1_add_69_carry_5_), 
        .A2(npu_inst_pe_1_2_1_int_q_acc_5_), .ZN(
        npu_inst_pe_1_2_1_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_2_1_U130 ( .A(npu_inst_pe_1_2_1_int_q_acc_6_), .B(
        npu_inst_pe_1_2_1_add_69_carry_6_), .Z(npu_inst_pe_1_2_1_N79) );
  AND2_X1 npu_inst_pe_1_2_1_U129 ( .A1(npu_inst_pe_1_2_1_add_69_carry_6_), 
        .A2(npu_inst_pe_1_2_1_int_q_acc_6_), .ZN(
        npu_inst_pe_1_2_1_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_2_1_U128 ( .A(npu_inst_pe_1_2_1_int_q_acc_7_), .B(
        npu_inst_pe_1_2_1_add_69_carry_7_), .Z(npu_inst_pe_1_2_1_N80) );
  XNOR2_X1 npu_inst_pe_1_2_1_U127 ( .A(npu_inst_pe_1_2_1_sub_67_carry_2_), .B(
        npu_inst_pe_1_2_1_int_q_acc_2_), .ZN(npu_inst_pe_1_2_1_N67) );
  OR2_X1 npu_inst_pe_1_2_1_U126 ( .A1(npu_inst_pe_1_2_1_int_q_acc_2_), .A2(
        npu_inst_pe_1_2_1_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_2_1_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_2_1_U125 ( .A(npu_inst_pe_1_2_1_sub_67_carry_3_), .B(
        npu_inst_pe_1_2_1_int_q_acc_3_), .ZN(npu_inst_pe_1_2_1_N68) );
  OR2_X1 npu_inst_pe_1_2_1_U124 ( .A1(npu_inst_pe_1_2_1_int_q_acc_3_), .A2(
        npu_inst_pe_1_2_1_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_2_1_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_2_1_U123 ( .A(npu_inst_pe_1_2_1_sub_67_carry_4_), .B(
        npu_inst_pe_1_2_1_int_q_acc_4_), .ZN(npu_inst_pe_1_2_1_N69) );
  OR2_X1 npu_inst_pe_1_2_1_U122 ( .A1(npu_inst_pe_1_2_1_int_q_acc_4_), .A2(
        npu_inst_pe_1_2_1_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_2_1_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_2_1_U121 ( .A(npu_inst_pe_1_2_1_sub_67_carry_5_), .B(
        npu_inst_pe_1_2_1_int_q_acc_5_), .ZN(npu_inst_pe_1_2_1_N70) );
  OR2_X1 npu_inst_pe_1_2_1_U120 ( .A1(npu_inst_pe_1_2_1_int_q_acc_5_), .A2(
        npu_inst_pe_1_2_1_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_2_1_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_2_1_U119 ( .A(npu_inst_pe_1_2_1_sub_67_carry_6_), .B(
        npu_inst_pe_1_2_1_int_q_acc_6_), .ZN(npu_inst_pe_1_2_1_N71) );
  OR2_X1 npu_inst_pe_1_2_1_U118 ( .A1(npu_inst_pe_1_2_1_int_q_acc_6_), .A2(
        npu_inst_pe_1_2_1_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_2_1_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_2_1_U117 ( .A(npu_inst_pe_1_2_1_int_q_acc_7_), .B(
        npu_inst_pe_1_2_1_sub_67_carry_7_), .ZN(npu_inst_pe_1_2_1_N72) );
  INV_X1 npu_inst_pe_1_2_1_U116 ( .A(npu_inst_n78), .ZN(npu_inst_pe_1_2_1_n7)
         );
  INV_X1 npu_inst_pe_1_2_1_U115 ( .A(npu_inst_pe_1_2_1_n7), .ZN(
        npu_inst_pe_1_2_1_n6) );
  INV_X1 npu_inst_pe_1_2_1_U114 ( .A(npu_inst_n58), .ZN(npu_inst_pe_1_2_1_n3)
         );
  AOI22_X1 npu_inst_pe_1_2_1_U113 ( .A1(npu_inst_int_data_y_3__1__0_), .A2(
        npu_inst_pe_1_2_1_n58), .B1(npu_inst_pe_1_2_1_n119), .B2(
        npu_inst_pe_1_2_1_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_2_1_n57) );
  INV_X1 npu_inst_pe_1_2_1_U112 ( .A(npu_inst_pe_1_2_1_n57), .ZN(
        npu_inst_pe_1_2_1_n108) );
  AOI22_X1 npu_inst_pe_1_2_1_U111 ( .A1(npu_inst_int_data_y_3__1__0_), .A2(
        npu_inst_pe_1_2_1_n54), .B1(npu_inst_pe_1_2_1_n118), .B2(
        npu_inst_pe_1_2_1_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_2_1_n53) );
  INV_X1 npu_inst_pe_1_2_1_U110 ( .A(npu_inst_pe_1_2_1_n53), .ZN(
        npu_inst_pe_1_2_1_n109) );
  AOI22_X1 npu_inst_pe_1_2_1_U107 ( .A1(npu_inst_int_data_y_3__1__0_), .A2(
        npu_inst_pe_1_2_1_n50), .B1(npu_inst_pe_1_2_1_n117), .B2(
        npu_inst_pe_1_2_1_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_2_1_n49) );
  INV_X1 npu_inst_pe_1_2_1_U106 ( .A(npu_inst_pe_1_2_1_n49), .ZN(
        npu_inst_pe_1_2_1_n110) );
  AOI22_X1 npu_inst_pe_1_2_1_U105 ( .A1(npu_inst_int_data_y_3__1__0_), .A2(
        npu_inst_pe_1_2_1_n46), .B1(npu_inst_pe_1_2_1_n116), .B2(
        npu_inst_pe_1_2_1_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_2_1_n45) );
  INV_X1 npu_inst_pe_1_2_1_U104 ( .A(npu_inst_pe_1_2_1_n45), .ZN(
        npu_inst_pe_1_2_1_n111) );
  AOI22_X1 npu_inst_pe_1_2_1_U103 ( .A1(npu_inst_int_data_y_3__1__0_), .A2(
        npu_inst_pe_1_2_1_n42), .B1(npu_inst_pe_1_2_1_n115), .B2(
        npu_inst_pe_1_2_1_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_2_1_n41) );
  INV_X1 npu_inst_pe_1_2_1_U102 ( .A(npu_inst_pe_1_2_1_n41), .ZN(
        npu_inst_pe_1_2_1_n112) );
  AOI22_X1 npu_inst_pe_1_2_1_U101 ( .A1(npu_inst_int_data_y_3__1__1_), .A2(
        npu_inst_pe_1_2_1_n58), .B1(npu_inst_pe_1_2_1_n119), .B2(
        npu_inst_pe_1_2_1_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_2_1_n59) );
  INV_X1 npu_inst_pe_1_2_1_U100 ( .A(npu_inst_pe_1_2_1_n59), .ZN(
        npu_inst_pe_1_2_1_n102) );
  AOI22_X1 npu_inst_pe_1_2_1_U99 ( .A1(npu_inst_int_data_y_3__1__1_), .A2(
        npu_inst_pe_1_2_1_n54), .B1(npu_inst_pe_1_2_1_n118), .B2(
        npu_inst_pe_1_2_1_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_2_1_n55) );
  INV_X1 npu_inst_pe_1_2_1_U98 ( .A(npu_inst_pe_1_2_1_n55), .ZN(
        npu_inst_pe_1_2_1_n103) );
  AOI22_X1 npu_inst_pe_1_2_1_U97 ( .A1(npu_inst_int_data_y_3__1__1_), .A2(
        npu_inst_pe_1_2_1_n50), .B1(npu_inst_pe_1_2_1_n117), .B2(
        npu_inst_pe_1_2_1_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_2_1_n51) );
  INV_X1 npu_inst_pe_1_2_1_U96 ( .A(npu_inst_pe_1_2_1_n51), .ZN(
        npu_inst_pe_1_2_1_n104) );
  AOI22_X1 npu_inst_pe_1_2_1_U95 ( .A1(npu_inst_int_data_y_3__1__1_), .A2(
        npu_inst_pe_1_2_1_n46), .B1(npu_inst_pe_1_2_1_n116), .B2(
        npu_inst_pe_1_2_1_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_2_1_n47) );
  INV_X1 npu_inst_pe_1_2_1_U94 ( .A(npu_inst_pe_1_2_1_n47), .ZN(
        npu_inst_pe_1_2_1_n105) );
  AOI22_X1 npu_inst_pe_1_2_1_U93 ( .A1(npu_inst_int_data_y_3__1__1_), .A2(
        npu_inst_pe_1_2_1_n42), .B1(npu_inst_pe_1_2_1_n115), .B2(
        npu_inst_pe_1_2_1_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_2_1_n43) );
  INV_X1 npu_inst_pe_1_2_1_U92 ( .A(npu_inst_pe_1_2_1_n43), .ZN(
        npu_inst_pe_1_2_1_n106) );
  AOI22_X1 npu_inst_pe_1_2_1_U91 ( .A1(npu_inst_pe_1_2_1_n38), .A2(
        npu_inst_int_data_y_3__1__1_), .B1(npu_inst_pe_1_2_1_n114), .B2(
        npu_inst_pe_1_2_1_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_2_1_n39) );
  INV_X1 npu_inst_pe_1_2_1_U90 ( .A(npu_inst_pe_1_2_1_n39), .ZN(
        npu_inst_pe_1_2_1_n107) );
  AOI22_X1 npu_inst_pe_1_2_1_U89 ( .A1(npu_inst_pe_1_2_1_n38), .A2(
        npu_inst_int_data_y_3__1__0_), .B1(npu_inst_pe_1_2_1_n114), .B2(
        npu_inst_pe_1_2_1_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_2_1_n37) );
  INV_X1 npu_inst_pe_1_2_1_U88 ( .A(npu_inst_pe_1_2_1_n37), .ZN(
        npu_inst_pe_1_2_1_n113) );
  NAND2_X1 npu_inst_pe_1_2_1_U87 ( .A1(npu_inst_pe_1_2_1_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_2_1_n60), .ZN(npu_inst_pe_1_2_1_n74) );
  OAI21_X1 npu_inst_pe_1_2_1_U86 ( .B1(npu_inst_pe_1_2_1_n63), .B2(
        npu_inst_pe_1_2_1_n60), .A(npu_inst_pe_1_2_1_n74), .ZN(
        npu_inst_pe_1_2_1_n97) );
  NAND2_X1 npu_inst_pe_1_2_1_U85 ( .A1(npu_inst_pe_1_2_1_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_2_1_n60), .ZN(npu_inst_pe_1_2_1_n73) );
  OAI21_X1 npu_inst_pe_1_2_1_U84 ( .B1(npu_inst_pe_1_2_1_n61), .B2(
        npu_inst_pe_1_2_1_n60), .A(npu_inst_pe_1_2_1_n73), .ZN(
        npu_inst_pe_1_2_1_n96) );
  NAND2_X1 npu_inst_pe_1_2_1_U83 ( .A1(npu_inst_pe_1_2_1_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_2_1_n56), .ZN(npu_inst_pe_1_2_1_n72) );
  OAI21_X1 npu_inst_pe_1_2_1_U82 ( .B1(npu_inst_pe_1_2_1_n63), .B2(
        npu_inst_pe_1_2_1_n56), .A(npu_inst_pe_1_2_1_n72), .ZN(
        npu_inst_pe_1_2_1_n95) );
  NAND2_X1 npu_inst_pe_1_2_1_U81 ( .A1(npu_inst_pe_1_2_1_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_2_1_n56), .ZN(npu_inst_pe_1_2_1_n71) );
  OAI21_X1 npu_inst_pe_1_2_1_U80 ( .B1(npu_inst_pe_1_2_1_n61), .B2(
        npu_inst_pe_1_2_1_n56), .A(npu_inst_pe_1_2_1_n71), .ZN(
        npu_inst_pe_1_2_1_n94) );
  NAND2_X1 npu_inst_pe_1_2_1_U79 ( .A1(npu_inst_pe_1_2_1_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_2_1_n52), .ZN(npu_inst_pe_1_2_1_n70) );
  OAI21_X1 npu_inst_pe_1_2_1_U78 ( .B1(npu_inst_pe_1_2_1_n63), .B2(
        npu_inst_pe_1_2_1_n52), .A(npu_inst_pe_1_2_1_n70), .ZN(
        npu_inst_pe_1_2_1_n93) );
  NAND2_X1 npu_inst_pe_1_2_1_U77 ( .A1(npu_inst_pe_1_2_1_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_2_1_n52), .ZN(npu_inst_pe_1_2_1_n69) );
  OAI21_X1 npu_inst_pe_1_2_1_U76 ( .B1(npu_inst_pe_1_2_1_n61), .B2(
        npu_inst_pe_1_2_1_n52), .A(npu_inst_pe_1_2_1_n69), .ZN(
        npu_inst_pe_1_2_1_n92) );
  NAND2_X1 npu_inst_pe_1_2_1_U75 ( .A1(npu_inst_pe_1_2_1_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_2_1_n48), .ZN(npu_inst_pe_1_2_1_n68) );
  OAI21_X1 npu_inst_pe_1_2_1_U74 ( .B1(npu_inst_pe_1_2_1_n63), .B2(
        npu_inst_pe_1_2_1_n48), .A(npu_inst_pe_1_2_1_n68), .ZN(
        npu_inst_pe_1_2_1_n91) );
  NAND2_X1 npu_inst_pe_1_2_1_U73 ( .A1(npu_inst_pe_1_2_1_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_2_1_n48), .ZN(npu_inst_pe_1_2_1_n67) );
  OAI21_X1 npu_inst_pe_1_2_1_U72 ( .B1(npu_inst_pe_1_2_1_n61), .B2(
        npu_inst_pe_1_2_1_n48), .A(npu_inst_pe_1_2_1_n67), .ZN(
        npu_inst_pe_1_2_1_n90) );
  NAND2_X1 npu_inst_pe_1_2_1_U71 ( .A1(npu_inst_pe_1_2_1_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_2_1_n44), .ZN(npu_inst_pe_1_2_1_n66) );
  OAI21_X1 npu_inst_pe_1_2_1_U70 ( .B1(npu_inst_pe_1_2_1_n63), .B2(
        npu_inst_pe_1_2_1_n44), .A(npu_inst_pe_1_2_1_n66), .ZN(
        npu_inst_pe_1_2_1_n89) );
  NAND2_X1 npu_inst_pe_1_2_1_U69 ( .A1(npu_inst_pe_1_2_1_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_2_1_n44), .ZN(npu_inst_pe_1_2_1_n65) );
  OAI21_X1 npu_inst_pe_1_2_1_U68 ( .B1(npu_inst_pe_1_2_1_n61), .B2(
        npu_inst_pe_1_2_1_n44), .A(npu_inst_pe_1_2_1_n65), .ZN(
        npu_inst_pe_1_2_1_n88) );
  NAND2_X1 npu_inst_pe_1_2_1_U67 ( .A1(npu_inst_pe_1_2_1_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_2_1_n40), .ZN(npu_inst_pe_1_2_1_n64) );
  OAI21_X1 npu_inst_pe_1_2_1_U66 ( .B1(npu_inst_pe_1_2_1_n63), .B2(
        npu_inst_pe_1_2_1_n40), .A(npu_inst_pe_1_2_1_n64), .ZN(
        npu_inst_pe_1_2_1_n87) );
  NAND2_X1 npu_inst_pe_1_2_1_U65 ( .A1(npu_inst_pe_1_2_1_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_2_1_n40), .ZN(npu_inst_pe_1_2_1_n62) );
  OAI21_X1 npu_inst_pe_1_2_1_U64 ( .B1(npu_inst_pe_1_2_1_n61), .B2(
        npu_inst_pe_1_2_1_n40), .A(npu_inst_pe_1_2_1_n62), .ZN(
        npu_inst_pe_1_2_1_n86) );
  AND2_X1 npu_inst_pe_1_2_1_U63 ( .A1(npu_inst_pe_1_2_1_N93), .A2(npu_inst_n58), .ZN(npu_inst_int_data_y_2__1__0_) );
  AND2_X1 npu_inst_pe_1_2_1_U62 ( .A1(npu_inst_n58), .A2(npu_inst_pe_1_2_1_N94), .ZN(npu_inst_int_data_y_2__1__1_) );
  NOR3_X1 npu_inst_pe_1_2_1_U61 ( .A1(npu_inst_pe_1_2_1_n26), .A2(npu_inst_n58), .A3(npu_inst_int_ckg[46]), .ZN(npu_inst_pe_1_2_1_n85) );
  OR2_X1 npu_inst_pe_1_2_1_U60 ( .A1(npu_inst_pe_1_2_1_n85), .A2(
        npu_inst_pe_1_2_1_n2), .ZN(npu_inst_pe_1_2_1_N84) );
  AND2_X1 npu_inst_pe_1_2_1_U59 ( .A1(npu_inst_pe_1_2_1_int_q_acc_0_), .A2(
        npu_inst_pe_1_2_1_n1), .ZN(npu_inst_int_data_res_2__1__0_) );
  AND2_X1 npu_inst_pe_1_2_1_U58 ( .A1(npu_inst_pe_1_2_1_n2), .A2(
        npu_inst_pe_1_2_1_int_q_acc_7_), .ZN(npu_inst_int_data_res_2__1__7_)
         );
  AND2_X1 npu_inst_pe_1_2_1_U57 ( .A1(npu_inst_pe_1_2_1_int_q_acc_1_), .A2(
        npu_inst_pe_1_2_1_n1), .ZN(npu_inst_int_data_res_2__1__1_) );
  AND2_X1 npu_inst_pe_1_2_1_U56 ( .A1(npu_inst_pe_1_2_1_int_q_acc_2_), .A2(
        npu_inst_pe_1_2_1_n1), .ZN(npu_inst_int_data_res_2__1__2_) );
  AND2_X1 npu_inst_pe_1_2_1_U55 ( .A1(npu_inst_pe_1_2_1_int_q_acc_3_), .A2(
        npu_inst_pe_1_2_1_n2), .ZN(npu_inst_int_data_res_2__1__3_) );
  AND2_X1 npu_inst_pe_1_2_1_U54 ( .A1(npu_inst_pe_1_2_1_int_q_acc_4_), .A2(
        npu_inst_pe_1_2_1_n2), .ZN(npu_inst_int_data_res_2__1__4_) );
  AND2_X1 npu_inst_pe_1_2_1_U53 ( .A1(npu_inst_pe_1_2_1_int_q_acc_5_), .A2(
        npu_inst_pe_1_2_1_n2), .ZN(npu_inst_int_data_res_2__1__5_) );
  AND2_X1 npu_inst_pe_1_2_1_U52 ( .A1(npu_inst_pe_1_2_1_int_q_acc_6_), .A2(
        npu_inst_pe_1_2_1_n2), .ZN(npu_inst_int_data_res_2__1__6_) );
  AOI222_X1 npu_inst_pe_1_2_1_U51 ( .A1(npu_inst_int_data_res_3__1__0_), .A2(
        npu_inst_pe_1_2_1_n1), .B1(npu_inst_pe_1_2_1_N73), .B2(
        npu_inst_pe_1_2_1_n76), .C1(npu_inst_pe_1_2_1_N65), .C2(
        npu_inst_pe_1_2_1_n77), .ZN(npu_inst_pe_1_2_1_n84) );
  INV_X1 npu_inst_pe_1_2_1_U50 ( .A(npu_inst_pe_1_2_1_n84), .ZN(
        npu_inst_pe_1_2_1_n101) );
  AOI222_X1 npu_inst_pe_1_2_1_U49 ( .A1(npu_inst_int_data_res_3__1__7_), .A2(
        npu_inst_pe_1_2_1_n1), .B1(npu_inst_pe_1_2_1_N80), .B2(
        npu_inst_pe_1_2_1_n76), .C1(npu_inst_pe_1_2_1_N72), .C2(
        npu_inst_pe_1_2_1_n77), .ZN(npu_inst_pe_1_2_1_n75) );
  INV_X1 npu_inst_pe_1_2_1_U48 ( .A(npu_inst_pe_1_2_1_n75), .ZN(
        npu_inst_pe_1_2_1_n33) );
  AOI222_X1 npu_inst_pe_1_2_1_U47 ( .A1(npu_inst_int_data_res_3__1__1_), .A2(
        npu_inst_pe_1_2_1_n1), .B1(npu_inst_pe_1_2_1_N74), .B2(
        npu_inst_pe_1_2_1_n76), .C1(npu_inst_pe_1_2_1_N66), .C2(
        npu_inst_pe_1_2_1_n77), .ZN(npu_inst_pe_1_2_1_n83) );
  INV_X1 npu_inst_pe_1_2_1_U46 ( .A(npu_inst_pe_1_2_1_n83), .ZN(
        npu_inst_pe_1_2_1_n100) );
  AOI222_X1 npu_inst_pe_1_2_1_U45 ( .A1(npu_inst_int_data_res_3__1__2_), .A2(
        npu_inst_pe_1_2_1_n1), .B1(npu_inst_pe_1_2_1_N75), .B2(
        npu_inst_pe_1_2_1_n76), .C1(npu_inst_pe_1_2_1_N67), .C2(
        npu_inst_pe_1_2_1_n77), .ZN(npu_inst_pe_1_2_1_n82) );
  INV_X1 npu_inst_pe_1_2_1_U44 ( .A(npu_inst_pe_1_2_1_n82), .ZN(
        npu_inst_pe_1_2_1_n99) );
  AOI222_X1 npu_inst_pe_1_2_1_U43 ( .A1(npu_inst_int_data_res_3__1__3_), .A2(
        npu_inst_pe_1_2_1_n1), .B1(npu_inst_pe_1_2_1_N76), .B2(
        npu_inst_pe_1_2_1_n76), .C1(npu_inst_pe_1_2_1_N68), .C2(
        npu_inst_pe_1_2_1_n77), .ZN(npu_inst_pe_1_2_1_n81) );
  INV_X1 npu_inst_pe_1_2_1_U42 ( .A(npu_inst_pe_1_2_1_n81), .ZN(
        npu_inst_pe_1_2_1_n98) );
  AOI222_X1 npu_inst_pe_1_2_1_U41 ( .A1(npu_inst_int_data_res_3__1__4_), .A2(
        npu_inst_pe_1_2_1_n1), .B1(npu_inst_pe_1_2_1_N77), .B2(
        npu_inst_pe_1_2_1_n76), .C1(npu_inst_pe_1_2_1_N69), .C2(
        npu_inst_pe_1_2_1_n77), .ZN(npu_inst_pe_1_2_1_n80) );
  INV_X1 npu_inst_pe_1_2_1_U40 ( .A(npu_inst_pe_1_2_1_n80), .ZN(
        npu_inst_pe_1_2_1_n36) );
  AOI222_X1 npu_inst_pe_1_2_1_U39 ( .A1(npu_inst_int_data_res_3__1__5_), .A2(
        npu_inst_pe_1_2_1_n1), .B1(npu_inst_pe_1_2_1_N78), .B2(
        npu_inst_pe_1_2_1_n76), .C1(npu_inst_pe_1_2_1_N70), .C2(
        npu_inst_pe_1_2_1_n77), .ZN(npu_inst_pe_1_2_1_n79) );
  INV_X1 npu_inst_pe_1_2_1_U38 ( .A(npu_inst_pe_1_2_1_n79), .ZN(
        npu_inst_pe_1_2_1_n35) );
  AOI222_X1 npu_inst_pe_1_2_1_U37 ( .A1(npu_inst_int_data_res_3__1__6_), .A2(
        npu_inst_pe_1_2_1_n1), .B1(npu_inst_pe_1_2_1_N79), .B2(
        npu_inst_pe_1_2_1_n76), .C1(npu_inst_pe_1_2_1_N71), .C2(
        npu_inst_pe_1_2_1_n77), .ZN(npu_inst_pe_1_2_1_n78) );
  INV_X1 npu_inst_pe_1_2_1_U36 ( .A(npu_inst_pe_1_2_1_n78), .ZN(
        npu_inst_pe_1_2_1_n34) );
  INV_X1 npu_inst_pe_1_2_1_U35 ( .A(npu_inst_pe_1_2_1_int_data_1_), .ZN(
        npu_inst_pe_1_2_1_n14) );
  AND2_X1 npu_inst_pe_1_2_1_U34 ( .A1(npu_inst_int_data_x_2__1__1_), .A2(
        npu_inst_pe_1_2_1_int_q_weight_1_), .ZN(npu_inst_pe_1_2_1_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_2_1_U33 ( .A1(npu_inst_int_data_x_2__1__0_), .A2(
        npu_inst_pe_1_2_1_int_q_weight_1_), .ZN(npu_inst_pe_1_2_1_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_2_1_U32 ( .A1(npu_inst_n58), .A2(
        npu_inst_int_data_y_3__1__1_), .B1(npu_inst_pe_1_2_1_n3), .B2(
        npu_inst_int_data_x_2__2__1_), .ZN(npu_inst_pe_1_2_1_n63) );
  AOI22_X1 npu_inst_pe_1_2_1_U31 ( .A1(npu_inst_n58), .A2(
        npu_inst_int_data_y_3__1__0_), .B1(npu_inst_pe_1_2_1_n3), .B2(
        npu_inst_int_data_x_2__2__0_), .ZN(npu_inst_pe_1_2_1_n61) );
  INV_X1 npu_inst_pe_1_2_1_U30 ( .A(npu_inst_pe_1_2_1_int_data_0_), .ZN(
        npu_inst_pe_1_2_1_n13) );
  INV_X1 npu_inst_pe_1_2_1_U29 ( .A(npu_inst_n70), .ZN(npu_inst_pe_1_2_1_n5)
         );
  OR3_X1 npu_inst_pe_1_2_1_U28 ( .A1(npu_inst_pe_1_2_1_n6), .A2(
        npu_inst_pe_1_2_1_n8), .A3(npu_inst_pe_1_2_1_n5), .ZN(
        npu_inst_pe_1_2_1_n56) );
  OR3_X1 npu_inst_pe_1_2_1_U27 ( .A1(npu_inst_pe_1_2_1_n5), .A2(
        npu_inst_pe_1_2_1_n8), .A3(npu_inst_pe_1_2_1_n7), .ZN(
        npu_inst_pe_1_2_1_n48) );
  INV_X1 npu_inst_pe_1_2_1_U26 ( .A(npu_inst_pe_1_2_1_n5), .ZN(
        npu_inst_pe_1_2_1_n4) );
  OR3_X1 npu_inst_pe_1_2_1_U25 ( .A1(npu_inst_pe_1_2_1_n4), .A2(
        npu_inst_pe_1_2_1_n8), .A3(npu_inst_pe_1_2_1_n7), .ZN(
        npu_inst_pe_1_2_1_n52) );
  OR3_X1 npu_inst_pe_1_2_1_U24 ( .A1(npu_inst_pe_1_2_1_n6), .A2(
        npu_inst_pe_1_2_1_n8), .A3(npu_inst_pe_1_2_1_n4), .ZN(
        npu_inst_pe_1_2_1_n60) );
  NOR2_X1 npu_inst_pe_1_2_1_U23 ( .A1(npu_inst_pe_1_2_1_n60), .A2(
        npu_inst_pe_1_2_1_n3), .ZN(npu_inst_pe_1_2_1_n58) );
  NOR2_X1 npu_inst_pe_1_2_1_U22 ( .A1(npu_inst_pe_1_2_1_n56), .A2(
        npu_inst_pe_1_2_1_n3), .ZN(npu_inst_pe_1_2_1_n54) );
  NOR2_X1 npu_inst_pe_1_2_1_U21 ( .A1(npu_inst_pe_1_2_1_n52), .A2(
        npu_inst_pe_1_2_1_n3), .ZN(npu_inst_pe_1_2_1_n50) );
  NOR2_X1 npu_inst_pe_1_2_1_U20 ( .A1(npu_inst_pe_1_2_1_n48), .A2(
        npu_inst_pe_1_2_1_n3), .ZN(npu_inst_pe_1_2_1_n46) );
  NOR2_X1 npu_inst_pe_1_2_1_U19 ( .A1(npu_inst_pe_1_2_1_n40), .A2(
        npu_inst_pe_1_2_1_n3), .ZN(npu_inst_pe_1_2_1_n38) );
  NOR2_X1 npu_inst_pe_1_2_1_U18 ( .A1(npu_inst_pe_1_2_1_n44), .A2(
        npu_inst_pe_1_2_1_n3), .ZN(npu_inst_pe_1_2_1_n42) );
  BUF_X1 npu_inst_pe_1_2_1_U17 ( .A(npu_inst_n103), .Z(npu_inst_pe_1_2_1_n8)
         );
  INV_X1 npu_inst_pe_1_2_1_U16 ( .A(npu_inst_n125), .ZN(npu_inst_pe_1_2_1_n12)
         );
  INV_X1 npu_inst_pe_1_2_1_U15 ( .A(npu_inst_pe_1_2_1_n38), .ZN(
        npu_inst_pe_1_2_1_n114) );
  INV_X1 npu_inst_pe_1_2_1_U14 ( .A(npu_inst_pe_1_2_1_n58), .ZN(
        npu_inst_pe_1_2_1_n119) );
  INV_X1 npu_inst_pe_1_2_1_U13 ( .A(npu_inst_pe_1_2_1_n54), .ZN(
        npu_inst_pe_1_2_1_n118) );
  INV_X1 npu_inst_pe_1_2_1_U12 ( .A(npu_inst_pe_1_2_1_n50), .ZN(
        npu_inst_pe_1_2_1_n117) );
  INV_X1 npu_inst_pe_1_2_1_U11 ( .A(npu_inst_pe_1_2_1_n46), .ZN(
        npu_inst_pe_1_2_1_n116) );
  INV_X1 npu_inst_pe_1_2_1_U10 ( .A(npu_inst_pe_1_2_1_n42), .ZN(
        npu_inst_pe_1_2_1_n115) );
  BUF_X1 npu_inst_pe_1_2_1_U9 ( .A(npu_inst_n30), .Z(npu_inst_pe_1_2_1_n2) );
  BUF_X1 npu_inst_pe_1_2_1_U8 ( .A(npu_inst_n30), .Z(npu_inst_pe_1_2_1_n1) );
  BUF_X1 npu_inst_pe_1_2_1_U7 ( .A(npu_inst_pe_1_2_1_n12), .Z(
        npu_inst_pe_1_2_1_n11) );
  BUF_X1 npu_inst_pe_1_2_1_U6 ( .A(npu_inst_pe_1_2_1_n12), .Z(
        npu_inst_pe_1_2_1_n10) );
  BUF_X1 npu_inst_pe_1_2_1_U5 ( .A(npu_inst_pe_1_2_1_n12), .Z(
        npu_inst_pe_1_2_1_n9) );
  NOR2_X1 npu_inst_pe_1_2_1_U4 ( .A1(npu_inst_pe_1_2_1_int_q_weight_0_), .A2(
        npu_inst_pe_1_2_1_n1), .ZN(npu_inst_pe_1_2_1_n76) );
  NOR2_X1 npu_inst_pe_1_2_1_U3 ( .A1(npu_inst_pe_1_2_1_n27), .A2(
        npu_inst_pe_1_2_1_n1), .ZN(npu_inst_pe_1_2_1_n77) );
  FA_X1 npu_inst_pe_1_2_1_sub_67_U2_1 ( .A(npu_inst_pe_1_2_1_int_q_acc_1_), 
        .B(npu_inst_pe_1_2_1_n14), .CI(npu_inst_pe_1_2_1_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_2_1_sub_67_carry_2_), .S(npu_inst_pe_1_2_1_N66) );
  FA_X1 npu_inst_pe_1_2_1_add_69_U1_1 ( .A(npu_inst_pe_1_2_1_int_q_acc_1_), 
        .B(npu_inst_pe_1_2_1_int_data_1_), .CI(
        npu_inst_pe_1_2_1_add_69_carry_1_), .CO(
        npu_inst_pe_1_2_1_add_69_carry_2_), .S(npu_inst_pe_1_2_1_N74) );
  NAND3_X1 npu_inst_pe_1_2_1_U109 ( .A1(npu_inst_pe_1_2_1_n5), .A2(
        npu_inst_pe_1_2_1_n7), .A3(npu_inst_pe_1_2_1_n8), .ZN(
        npu_inst_pe_1_2_1_n44) );
  NAND3_X1 npu_inst_pe_1_2_1_U108 ( .A1(npu_inst_pe_1_2_1_n4), .A2(
        npu_inst_pe_1_2_1_n7), .A3(npu_inst_pe_1_2_1_n8), .ZN(
        npu_inst_pe_1_2_1_n40) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_2_1_n34), .CK(
        npu_inst_pe_1_2_1_net4171), .RN(npu_inst_pe_1_2_1_n9), .Q(
        npu_inst_pe_1_2_1_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_2_1_n35), .CK(
        npu_inst_pe_1_2_1_net4171), .RN(npu_inst_pe_1_2_1_n9), .Q(
        npu_inst_pe_1_2_1_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_2_1_n36), .CK(
        npu_inst_pe_1_2_1_net4171), .RN(npu_inst_pe_1_2_1_n9), .Q(
        npu_inst_pe_1_2_1_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_2_1_n98), .CK(
        npu_inst_pe_1_2_1_net4171), .RN(npu_inst_pe_1_2_1_n9), .Q(
        npu_inst_pe_1_2_1_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_2_1_n99), .CK(
        npu_inst_pe_1_2_1_net4171), .RN(npu_inst_pe_1_2_1_n9), .Q(
        npu_inst_pe_1_2_1_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_2_1_n100), 
        .CK(npu_inst_pe_1_2_1_net4171), .RN(npu_inst_pe_1_2_1_n9), .Q(
        npu_inst_pe_1_2_1_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_2_1_n33), .CK(
        npu_inst_pe_1_2_1_net4171), .RN(npu_inst_pe_1_2_1_n9), .Q(
        npu_inst_pe_1_2_1_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_2_1_n101), 
        .CK(npu_inst_pe_1_2_1_net4171), .RN(npu_inst_pe_1_2_1_n9), .Q(
        npu_inst_pe_1_2_1_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_weight_reg_0_ ( .D(npu_inst_n111), .CK(
        npu_inst_pe_1_2_1_net4177), .RN(npu_inst_pe_1_2_1_n9), .Q(
        npu_inst_pe_1_2_1_int_q_weight_0_), .QN(npu_inst_pe_1_2_1_n27) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_weight_reg_1_ ( .D(npu_inst_n117), .CK(
        npu_inst_pe_1_2_1_net4177), .RN(npu_inst_pe_1_2_1_n9), .Q(
        npu_inst_pe_1_2_1_int_q_weight_1_), .QN(npu_inst_pe_1_2_1_n26) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_2_1_n113), 
        .CK(npu_inst_pe_1_2_1_net4177), .RN(npu_inst_pe_1_2_1_n9), .Q(
        npu_inst_pe_1_2_1_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_2_1_n107), 
        .CK(npu_inst_pe_1_2_1_net4177), .RN(npu_inst_pe_1_2_1_n9), .Q(
        npu_inst_pe_1_2_1_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_2_1_n112), 
        .CK(npu_inst_pe_1_2_1_net4177), .RN(npu_inst_pe_1_2_1_n10), .Q(
        npu_inst_pe_1_2_1_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_2_1_n106), 
        .CK(npu_inst_pe_1_2_1_net4177), .RN(npu_inst_pe_1_2_1_n10), .Q(
        npu_inst_pe_1_2_1_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_2_1_n111), 
        .CK(npu_inst_pe_1_2_1_net4177), .RN(npu_inst_pe_1_2_1_n10), .Q(
        npu_inst_pe_1_2_1_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_2_1_n105), 
        .CK(npu_inst_pe_1_2_1_net4177), .RN(npu_inst_pe_1_2_1_n10), .Q(
        npu_inst_pe_1_2_1_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_2_1_n110), 
        .CK(npu_inst_pe_1_2_1_net4177), .RN(npu_inst_pe_1_2_1_n10), .Q(
        npu_inst_pe_1_2_1_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_2_1_n104), 
        .CK(npu_inst_pe_1_2_1_net4177), .RN(npu_inst_pe_1_2_1_n10), .Q(
        npu_inst_pe_1_2_1_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_2_1_n109), 
        .CK(npu_inst_pe_1_2_1_net4177), .RN(npu_inst_pe_1_2_1_n10), .Q(
        npu_inst_pe_1_2_1_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_2_1_n103), 
        .CK(npu_inst_pe_1_2_1_net4177), .RN(npu_inst_pe_1_2_1_n10), .Q(
        npu_inst_pe_1_2_1_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_2_1_n108), 
        .CK(npu_inst_pe_1_2_1_net4177), .RN(npu_inst_pe_1_2_1_n10), .Q(
        npu_inst_pe_1_2_1_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_2_1_n102), 
        .CK(npu_inst_pe_1_2_1_net4177), .RN(npu_inst_pe_1_2_1_n10), .Q(
        npu_inst_pe_1_2_1_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_2_1_n86), 
        .CK(npu_inst_pe_1_2_1_net4177), .RN(npu_inst_pe_1_2_1_n10), .Q(
        npu_inst_pe_1_2_1_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_2_1_n87), 
        .CK(npu_inst_pe_1_2_1_net4177), .RN(npu_inst_pe_1_2_1_n10), .Q(
        npu_inst_pe_1_2_1_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_2_1_n88), 
        .CK(npu_inst_pe_1_2_1_net4177), .RN(npu_inst_pe_1_2_1_n11), .Q(
        npu_inst_pe_1_2_1_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_2_1_n89), 
        .CK(npu_inst_pe_1_2_1_net4177), .RN(npu_inst_pe_1_2_1_n11), .Q(
        npu_inst_pe_1_2_1_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_2_1_n90), 
        .CK(npu_inst_pe_1_2_1_net4177), .RN(npu_inst_pe_1_2_1_n11), .Q(
        npu_inst_pe_1_2_1_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_2_1_n91), 
        .CK(npu_inst_pe_1_2_1_net4177), .RN(npu_inst_pe_1_2_1_n11), .Q(
        npu_inst_pe_1_2_1_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_2_1_n92), 
        .CK(npu_inst_pe_1_2_1_net4177), .RN(npu_inst_pe_1_2_1_n11), .Q(
        npu_inst_pe_1_2_1_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_2_1_n93), 
        .CK(npu_inst_pe_1_2_1_net4177), .RN(npu_inst_pe_1_2_1_n11), .Q(
        npu_inst_pe_1_2_1_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_2_1_n94), 
        .CK(npu_inst_pe_1_2_1_net4177), .RN(npu_inst_pe_1_2_1_n11), .Q(
        npu_inst_pe_1_2_1_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_2_1_n95), 
        .CK(npu_inst_pe_1_2_1_net4177), .RN(npu_inst_pe_1_2_1_n11), .Q(
        npu_inst_pe_1_2_1_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_2_1_n96), 
        .CK(npu_inst_pe_1_2_1_net4177), .RN(npu_inst_pe_1_2_1_n11), .Q(
        npu_inst_pe_1_2_1_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_2_1_n97), 
        .CK(npu_inst_pe_1_2_1_net4177), .RN(npu_inst_pe_1_2_1_n11), .Q(
        npu_inst_pe_1_2_1_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_2_1_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_2_1_N84), .SE(1'b0), .GCK(npu_inst_pe_1_2_1_net4171) );
  CLKGATETST_X1 npu_inst_pe_1_2_1_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n65), .SE(1'b0), .GCK(npu_inst_pe_1_2_1_net4177) );
  MUX2_X1 npu_inst_pe_1_2_2_U162 ( .A(npu_inst_pe_1_2_2_n32), .B(
        npu_inst_pe_1_2_2_n29), .S(npu_inst_pe_1_2_2_n8), .Z(
        npu_inst_pe_1_2_2_N93) );
  MUX2_X1 npu_inst_pe_1_2_2_U161 ( .A(npu_inst_pe_1_2_2_n31), .B(
        npu_inst_pe_1_2_2_n30), .S(npu_inst_pe_1_2_2_n6), .Z(
        npu_inst_pe_1_2_2_n32) );
  MUX2_X1 npu_inst_pe_1_2_2_U160 ( .A(npu_inst_pe_1_2_2_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_2_2_int_q_reg_v_1__0_), .S(npu_inst_pe_1_2_2_n4), .Z(
        npu_inst_pe_1_2_2_n31) );
  MUX2_X1 npu_inst_pe_1_2_2_U159 ( .A(npu_inst_pe_1_2_2_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_2_2_int_q_reg_v_3__0_), .S(npu_inst_pe_1_2_2_n4), .Z(
        npu_inst_pe_1_2_2_n30) );
  MUX2_X1 npu_inst_pe_1_2_2_U158 ( .A(npu_inst_pe_1_2_2_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_2_2_int_q_reg_v_5__0_), .S(npu_inst_pe_1_2_2_n4), .Z(
        npu_inst_pe_1_2_2_n29) );
  MUX2_X1 npu_inst_pe_1_2_2_U157 ( .A(npu_inst_pe_1_2_2_n28), .B(
        npu_inst_pe_1_2_2_n23), .S(npu_inst_pe_1_2_2_n8), .Z(
        npu_inst_pe_1_2_2_N94) );
  MUX2_X1 npu_inst_pe_1_2_2_U156 ( .A(npu_inst_pe_1_2_2_n25), .B(
        npu_inst_pe_1_2_2_n24), .S(npu_inst_pe_1_2_2_n6), .Z(
        npu_inst_pe_1_2_2_n28) );
  MUX2_X1 npu_inst_pe_1_2_2_U155 ( .A(npu_inst_pe_1_2_2_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_2_2_int_q_reg_v_1__1_), .S(npu_inst_pe_1_2_2_n4), .Z(
        npu_inst_pe_1_2_2_n25) );
  MUX2_X1 npu_inst_pe_1_2_2_U154 ( .A(npu_inst_pe_1_2_2_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_2_2_int_q_reg_v_3__1_), .S(npu_inst_pe_1_2_2_n4), .Z(
        npu_inst_pe_1_2_2_n24) );
  MUX2_X1 npu_inst_pe_1_2_2_U153 ( .A(npu_inst_pe_1_2_2_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_2_2_int_q_reg_v_5__1_), .S(npu_inst_pe_1_2_2_n4), .Z(
        npu_inst_pe_1_2_2_n23) );
  MUX2_X1 npu_inst_pe_1_2_2_U152 ( .A(npu_inst_pe_1_2_2_n22), .B(
        npu_inst_pe_1_2_2_n19), .S(npu_inst_pe_1_2_2_n8), .Z(
        npu_inst_int_data_x_2__2__1_) );
  MUX2_X1 npu_inst_pe_1_2_2_U151 ( .A(npu_inst_pe_1_2_2_n21), .B(
        npu_inst_pe_1_2_2_n20), .S(npu_inst_pe_1_2_2_n6), .Z(
        npu_inst_pe_1_2_2_n22) );
  MUX2_X1 npu_inst_pe_1_2_2_U150 ( .A(npu_inst_pe_1_2_2_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_2_2_int_q_reg_h_1__1_), .S(npu_inst_pe_1_2_2_n4), .Z(
        npu_inst_pe_1_2_2_n21) );
  MUX2_X1 npu_inst_pe_1_2_2_U149 ( .A(npu_inst_pe_1_2_2_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_2_2_int_q_reg_h_3__1_), .S(npu_inst_pe_1_2_2_n4), .Z(
        npu_inst_pe_1_2_2_n20) );
  MUX2_X1 npu_inst_pe_1_2_2_U148 ( .A(npu_inst_pe_1_2_2_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_2_2_int_q_reg_h_5__1_), .S(npu_inst_pe_1_2_2_n4), .Z(
        npu_inst_pe_1_2_2_n19) );
  MUX2_X1 npu_inst_pe_1_2_2_U147 ( .A(npu_inst_pe_1_2_2_n18), .B(
        npu_inst_pe_1_2_2_n15), .S(npu_inst_pe_1_2_2_n8), .Z(
        npu_inst_int_data_x_2__2__0_) );
  MUX2_X1 npu_inst_pe_1_2_2_U146 ( .A(npu_inst_pe_1_2_2_n17), .B(
        npu_inst_pe_1_2_2_n16), .S(npu_inst_pe_1_2_2_n6), .Z(
        npu_inst_pe_1_2_2_n18) );
  MUX2_X1 npu_inst_pe_1_2_2_U145 ( .A(npu_inst_pe_1_2_2_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_2_2_int_q_reg_h_1__0_), .S(npu_inst_pe_1_2_2_n4), .Z(
        npu_inst_pe_1_2_2_n17) );
  MUX2_X1 npu_inst_pe_1_2_2_U144 ( .A(npu_inst_pe_1_2_2_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_2_2_int_q_reg_h_3__0_), .S(npu_inst_pe_1_2_2_n4), .Z(
        npu_inst_pe_1_2_2_n16) );
  MUX2_X1 npu_inst_pe_1_2_2_U143 ( .A(npu_inst_pe_1_2_2_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_2_2_int_q_reg_h_5__0_), .S(npu_inst_pe_1_2_2_n4), .Z(
        npu_inst_pe_1_2_2_n15) );
  XOR2_X1 npu_inst_pe_1_2_2_U142 ( .A(npu_inst_pe_1_2_2_int_data_0_), .B(
        npu_inst_pe_1_2_2_int_q_acc_0_), .Z(npu_inst_pe_1_2_2_N73) );
  AND2_X1 npu_inst_pe_1_2_2_U141 ( .A1(npu_inst_pe_1_2_2_int_q_acc_0_), .A2(
        npu_inst_pe_1_2_2_int_data_0_), .ZN(npu_inst_pe_1_2_2_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_2_2_U140 ( .A(npu_inst_pe_1_2_2_int_q_acc_0_), .B(
        npu_inst_pe_1_2_2_n13), .ZN(npu_inst_pe_1_2_2_N65) );
  OR2_X1 npu_inst_pe_1_2_2_U139 ( .A1(npu_inst_pe_1_2_2_n13), .A2(
        npu_inst_pe_1_2_2_int_q_acc_0_), .ZN(npu_inst_pe_1_2_2_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_2_2_U138 ( .A(npu_inst_pe_1_2_2_int_q_acc_2_), .B(
        npu_inst_pe_1_2_2_add_69_carry_2_), .Z(npu_inst_pe_1_2_2_N75) );
  AND2_X1 npu_inst_pe_1_2_2_U137 ( .A1(npu_inst_pe_1_2_2_add_69_carry_2_), 
        .A2(npu_inst_pe_1_2_2_int_q_acc_2_), .ZN(
        npu_inst_pe_1_2_2_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_2_2_U136 ( .A(npu_inst_pe_1_2_2_int_q_acc_3_), .B(
        npu_inst_pe_1_2_2_add_69_carry_3_), .Z(npu_inst_pe_1_2_2_N76) );
  AND2_X1 npu_inst_pe_1_2_2_U135 ( .A1(npu_inst_pe_1_2_2_add_69_carry_3_), 
        .A2(npu_inst_pe_1_2_2_int_q_acc_3_), .ZN(
        npu_inst_pe_1_2_2_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_2_2_U134 ( .A(npu_inst_pe_1_2_2_int_q_acc_4_), .B(
        npu_inst_pe_1_2_2_add_69_carry_4_), .Z(npu_inst_pe_1_2_2_N77) );
  AND2_X1 npu_inst_pe_1_2_2_U133 ( .A1(npu_inst_pe_1_2_2_add_69_carry_4_), 
        .A2(npu_inst_pe_1_2_2_int_q_acc_4_), .ZN(
        npu_inst_pe_1_2_2_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_2_2_U132 ( .A(npu_inst_pe_1_2_2_int_q_acc_5_), .B(
        npu_inst_pe_1_2_2_add_69_carry_5_), .Z(npu_inst_pe_1_2_2_N78) );
  AND2_X1 npu_inst_pe_1_2_2_U131 ( .A1(npu_inst_pe_1_2_2_add_69_carry_5_), 
        .A2(npu_inst_pe_1_2_2_int_q_acc_5_), .ZN(
        npu_inst_pe_1_2_2_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_2_2_U130 ( .A(npu_inst_pe_1_2_2_int_q_acc_6_), .B(
        npu_inst_pe_1_2_2_add_69_carry_6_), .Z(npu_inst_pe_1_2_2_N79) );
  AND2_X1 npu_inst_pe_1_2_2_U129 ( .A1(npu_inst_pe_1_2_2_add_69_carry_6_), 
        .A2(npu_inst_pe_1_2_2_int_q_acc_6_), .ZN(
        npu_inst_pe_1_2_2_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_2_2_U128 ( .A(npu_inst_pe_1_2_2_int_q_acc_7_), .B(
        npu_inst_pe_1_2_2_add_69_carry_7_), .Z(npu_inst_pe_1_2_2_N80) );
  XNOR2_X1 npu_inst_pe_1_2_2_U127 ( .A(npu_inst_pe_1_2_2_sub_67_carry_2_), .B(
        npu_inst_pe_1_2_2_int_q_acc_2_), .ZN(npu_inst_pe_1_2_2_N67) );
  OR2_X1 npu_inst_pe_1_2_2_U126 ( .A1(npu_inst_pe_1_2_2_int_q_acc_2_), .A2(
        npu_inst_pe_1_2_2_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_2_2_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_2_2_U125 ( .A(npu_inst_pe_1_2_2_sub_67_carry_3_), .B(
        npu_inst_pe_1_2_2_int_q_acc_3_), .ZN(npu_inst_pe_1_2_2_N68) );
  OR2_X1 npu_inst_pe_1_2_2_U124 ( .A1(npu_inst_pe_1_2_2_int_q_acc_3_), .A2(
        npu_inst_pe_1_2_2_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_2_2_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_2_2_U123 ( .A(npu_inst_pe_1_2_2_sub_67_carry_4_), .B(
        npu_inst_pe_1_2_2_int_q_acc_4_), .ZN(npu_inst_pe_1_2_2_N69) );
  OR2_X1 npu_inst_pe_1_2_2_U122 ( .A1(npu_inst_pe_1_2_2_int_q_acc_4_), .A2(
        npu_inst_pe_1_2_2_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_2_2_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_2_2_U121 ( .A(npu_inst_pe_1_2_2_sub_67_carry_5_), .B(
        npu_inst_pe_1_2_2_int_q_acc_5_), .ZN(npu_inst_pe_1_2_2_N70) );
  OR2_X1 npu_inst_pe_1_2_2_U120 ( .A1(npu_inst_pe_1_2_2_int_q_acc_5_), .A2(
        npu_inst_pe_1_2_2_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_2_2_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_2_2_U119 ( .A(npu_inst_pe_1_2_2_sub_67_carry_6_), .B(
        npu_inst_pe_1_2_2_int_q_acc_6_), .ZN(npu_inst_pe_1_2_2_N71) );
  OR2_X1 npu_inst_pe_1_2_2_U118 ( .A1(npu_inst_pe_1_2_2_int_q_acc_6_), .A2(
        npu_inst_pe_1_2_2_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_2_2_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_2_2_U117 ( .A(npu_inst_pe_1_2_2_int_q_acc_7_), .B(
        npu_inst_pe_1_2_2_sub_67_carry_7_), .ZN(npu_inst_pe_1_2_2_N72) );
  INV_X1 npu_inst_pe_1_2_2_U116 ( .A(npu_inst_n78), .ZN(npu_inst_pe_1_2_2_n7)
         );
  INV_X1 npu_inst_pe_1_2_2_U115 ( .A(npu_inst_pe_1_2_2_n7), .ZN(
        npu_inst_pe_1_2_2_n6) );
  INV_X1 npu_inst_pe_1_2_2_U114 ( .A(npu_inst_n58), .ZN(npu_inst_pe_1_2_2_n3)
         );
  AOI22_X1 npu_inst_pe_1_2_2_U113 ( .A1(npu_inst_int_data_y_3__2__0_), .A2(
        npu_inst_pe_1_2_2_n58), .B1(npu_inst_pe_1_2_2_n119), .B2(
        npu_inst_pe_1_2_2_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_2_2_n57) );
  INV_X1 npu_inst_pe_1_2_2_U112 ( .A(npu_inst_pe_1_2_2_n57), .ZN(
        npu_inst_pe_1_2_2_n108) );
  AOI22_X1 npu_inst_pe_1_2_2_U111 ( .A1(npu_inst_int_data_y_3__2__0_), .A2(
        npu_inst_pe_1_2_2_n54), .B1(npu_inst_pe_1_2_2_n118), .B2(
        npu_inst_pe_1_2_2_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_2_2_n53) );
  INV_X1 npu_inst_pe_1_2_2_U110 ( .A(npu_inst_pe_1_2_2_n53), .ZN(
        npu_inst_pe_1_2_2_n109) );
  AOI22_X1 npu_inst_pe_1_2_2_U107 ( .A1(npu_inst_int_data_y_3__2__0_), .A2(
        npu_inst_pe_1_2_2_n50), .B1(npu_inst_pe_1_2_2_n117), .B2(
        npu_inst_pe_1_2_2_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_2_2_n49) );
  INV_X1 npu_inst_pe_1_2_2_U106 ( .A(npu_inst_pe_1_2_2_n49), .ZN(
        npu_inst_pe_1_2_2_n110) );
  AOI22_X1 npu_inst_pe_1_2_2_U105 ( .A1(npu_inst_int_data_y_3__2__0_), .A2(
        npu_inst_pe_1_2_2_n46), .B1(npu_inst_pe_1_2_2_n116), .B2(
        npu_inst_pe_1_2_2_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_2_2_n45) );
  INV_X1 npu_inst_pe_1_2_2_U104 ( .A(npu_inst_pe_1_2_2_n45), .ZN(
        npu_inst_pe_1_2_2_n111) );
  AOI22_X1 npu_inst_pe_1_2_2_U103 ( .A1(npu_inst_int_data_y_3__2__0_), .A2(
        npu_inst_pe_1_2_2_n42), .B1(npu_inst_pe_1_2_2_n115), .B2(
        npu_inst_pe_1_2_2_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_2_2_n41) );
  INV_X1 npu_inst_pe_1_2_2_U102 ( .A(npu_inst_pe_1_2_2_n41), .ZN(
        npu_inst_pe_1_2_2_n112) );
  AOI22_X1 npu_inst_pe_1_2_2_U101 ( .A1(npu_inst_int_data_y_3__2__1_), .A2(
        npu_inst_pe_1_2_2_n58), .B1(npu_inst_pe_1_2_2_n119), .B2(
        npu_inst_pe_1_2_2_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_2_2_n59) );
  INV_X1 npu_inst_pe_1_2_2_U100 ( .A(npu_inst_pe_1_2_2_n59), .ZN(
        npu_inst_pe_1_2_2_n102) );
  AOI22_X1 npu_inst_pe_1_2_2_U99 ( .A1(npu_inst_int_data_y_3__2__1_), .A2(
        npu_inst_pe_1_2_2_n54), .B1(npu_inst_pe_1_2_2_n118), .B2(
        npu_inst_pe_1_2_2_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_2_2_n55) );
  INV_X1 npu_inst_pe_1_2_2_U98 ( .A(npu_inst_pe_1_2_2_n55), .ZN(
        npu_inst_pe_1_2_2_n103) );
  AOI22_X1 npu_inst_pe_1_2_2_U97 ( .A1(npu_inst_int_data_y_3__2__1_), .A2(
        npu_inst_pe_1_2_2_n50), .B1(npu_inst_pe_1_2_2_n117), .B2(
        npu_inst_pe_1_2_2_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_2_2_n51) );
  INV_X1 npu_inst_pe_1_2_2_U96 ( .A(npu_inst_pe_1_2_2_n51), .ZN(
        npu_inst_pe_1_2_2_n104) );
  AOI22_X1 npu_inst_pe_1_2_2_U95 ( .A1(npu_inst_int_data_y_3__2__1_), .A2(
        npu_inst_pe_1_2_2_n46), .B1(npu_inst_pe_1_2_2_n116), .B2(
        npu_inst_pe_1_2_2_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_2_2_n47) );
  INV_X1 npu_inst_pe_1_2_2_U94 ( .A(npu_inst_pe_1_2_2_n47), .ZN(
        npu_inst_pe_1_2_2_n105) );
  AOI22_X1 npu_inst_pe_1_2_2_U93 ( .A1(npu_inst_int_data_y_3__2__1_), .A2(
        npu_inst_pe_1_2_2_n42), .B1(npu_inst_pe_1_2_2_n115), .B2(
        npu_inst_pe_1_2_2_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_2_2_n43) );
  INV_X1 npu_inst_pe_1_2_2_U92 ( .A(npu_inst_pe_1_2_2_n43), .ZN(
        npu_inst_pe_1_2_2_n106) );
  AOI22_X1 npu_inst_pe_1_2_2_U91 ( .A1(npu_inst_pe_1_2_2_n38), .A2(
        npu_inst_int_data_y_3__2__1_), .B1(npu_inst_pe_1_2_2_n114), .B2(
        npu_inst_pe_1_2_2_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_2_2_n39) );
  INV_X1 npu_inst_pe_1_2_2_U90 ( .A(npu_inst_pe_1_2_2_n39), .ZN(
        npu_inst_pe_1_2_2_n107) );
  AOI22_X1 npu_inst_pe_1_2_2_U89 ( .A1(npu_inst_pe_1_2_2_n38), .A2(
        npu_inst_int_data_y_3__2__0_), .B1(npu_inst_pe_1_2_2_n114), .B2(
        npu_inst_pe_1_2_2_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_2_2_n37) );
  INV_X1 npu_inst_pe_1_2_2_U88 ( .A(npu_inst_pe_1_2_2_n37), .ZN(
        npu_inst_pe_1_2_2_n113) );
  NAND2_X1 npu_inst_pe_1_2_2_U87 ( .A1(npu_inst_pe_1_2_2_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_2_2_n60), .ZN(npu_inst_pe_1_2_2_n74) );
  OAI21_X1 npu_inst_pe_1_2_2_U86 ( .B1(npu_inst_pe_1_2_2_n63), .B2(
        npu_inst_pe_1_2_2_n60), .A(npu_inst_pe_1_2_2_n74), .ZN(
        npu_inst_pe_1_2_2_n97) );
  NAND2_X1 npu_inst_pe_1_2_2_U85 ( .A1(npu_inst_pe_1_2_2_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_2_2_n60), .ZN(npu_inst_pe_1_2_2_n73) );
  OAI21_X1 npu_inst_pe_1_2_2_U84 ( .B1(npu_inst_pe_1_2_2_n61), .B2(
        npu_inst_pe_1_2_2_n60), .A(npu_inst_pe_1_2_2_n73), .ZN(
        npu_inst_pe_1_2_2_n96) );
  NAND2_X1 npu_inst_pe_1_2_2_U83 ( .A1(npu_inst_pe_1_2_2_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_2_2_n56), .ZN(npu_inst_pe_1_2_2_n72) );
  OAI21_X1 npu_inst_pe_1_2_2_U82 ( .B1(npu_inst_pe_1_2_2_n63), .B2(
        npu_inst_pe_1_2_2_n56), .A(npu_inst_pe_1_2_2_n72), .ZN(
        npu_inst_pe_1_2_2_n95) );
  NAND2_X1 npu_inst_pe_1_2_2_U81 ( .A1(npu_inst_pe_1_2_2_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_2_2_n56), .ZN(npu_inst_pe_1_2_2_n71) );
  OAI21_X1 npu_inst_pe_1_2_2_U80 ( .B1(npu_inst_pe_1_2_2_n61), .B2(
        npu_inst_pe_1_2_2_n56), .A(npu_inst_pe_1_2_2_n71), .ZN(
        npu_inst_pe_1_2_2_n94) );
  NAND2_X1 npu_inst_pe_1_2_2_U79 ( .A1(npu_inst_pe_1_2_2_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_2_2_n52), .ZN(npu_inst_pe_1_2_2_n70) );
  OAI21_X1 npu_inst_pe_1_2_2_U78 ( .B1(npu_inst_pe_1_2_2_n63), .B2(
        npu_inst_pe_1_2_2_n52), .A(npu_inst_pe_1_2_2_n70), .ZN(
        npu_inst_pe_1_2_2_n93) );
  NAND2_X1 npu_inst_pe_1_2_2_U77 ( .A1(npu_inst_pe_1_2_2_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_2_2_n52), .ZN(npu_inst_pe_1_2_2_n69) );
  OAI21_X1 npu_inst_pe_1_2_2_U76 ( .B1(npu_inst_pe_1_2_2_n61), .B2(
        npu_inst_pe_1_2_2_n52), .A(npu_inst_pe_1_2_2_n69), .ZN(
        npu_inst_pe_1_2_2_n92) );
  NAND2_X1 npu_inst_pe_1_2_2_U75 ( .A1(npu_inst_pe_1_2_2_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_2_2_n48), .ZN(npu_inst_pe_1_2_2_n68) );
  OAI21_X1 npu_inst_pe_1_2_2_U74 ( .B1(npu_inst_pe_1_2_2_n63), .B2(
        npu_inst_pe_1_2_2_n48), .A(npu_inst_pe_1_2_2_n68), .ZN(
        npu_inst_pe_1_2_2_n91) );
  NAND2_X1 npu_inst_pe_1_2_2_U73 ( .A1(npu_inst_pe_1_2_2_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_2_2_n48), .ZN(npu_inst_pe_1_2_2_n67) );
  OAI21_X1 npu_inst_pe_1_2_2_U72 ( .B1(npu_inst_pe_1_2_2_n61), .B2(
        npu_inst_pe_1_2_2_n48), .A(npu_inst_pe_1_2_2_n67), .ZN(
        npu_inst_pe_1_2_2_n90) );
  NAND2_X1 npu_inst_pe_1_2_2_U71 ( .A1(npu_inst_pe_1_2_2_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_2_2_n44), .ZN(npu_inst_pe_1_2_2_n66) );
  OAI21_X1 npu_inst_pe_1_2_2_U70 ( .B1(npu_inst_pe_1_2_2_n63), .B2(
        npu_inst_pe_1_2_2_n44), .A(npu_inst_pe_1_2_2_n66), .ZN(
        npu_inst_pe_1_2_2_n89) );
  NAND2_X1 npu_inst_pe_1_2_2_U69 ( .A1(npu_inst_pe_1_2_2_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_2_2_n44), .ZN(npu_inst_pe_1_2_2_n65) );
  OAI21_X1 npu_inst_pe_1_2_2_U68 ( .B1(npu_inst_pe_1_2_2_n61), .B2(
        npu_inst_pe_1_2_2_n44), .A(npu_inst_pe_1_2_2_n65), .ZN(
        npu_inst_pe_1_2_2_n88) );
  NAND2_X1 npu_inst_pe_1_2_2_U67 ( .A1(npu_inst_pe_1_2_2_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_2_2_n40), .ZN(npu_inst_pe_1_2_2_n64) );
  OAI21_X1 npu_inst_pe_1_2_2_U66 ( .B1(npu_inst_pe_1_2_2_n63), .B2(
        npu_inst_pe_1_2_2_n40), .A(npu_inst_pe_1_2_2_n64), .ZN(
        npu_inst_pe_1_2_2_n87) );
  NAND2_X1 npu_inst_pe_1_2_2_U65 ( .A1(npu_inst_pe_1_2_2_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_2_2_n40), .ZN(npu_inst_pe_1_2_2_n62) );
  OAI21_X1 npu_inst_pe_1_2_2_U64 ( .B1(npu_inst_pe_1_2_2_n61), .B2(
        npu_inst_pe_1_2_2_n40), .A(npu_inst_pe_1_2_2_n62), .ZN(
        npu_inst_pe_1_2_2_n86) );
  AND2_X1 npu_inst_pe_1_2_2_U63 ( .A1(npu_inst_pe_1_2_2_N93), .A2(npu_inst_n58), .ZN(npu_inst_int_data_y_2__2__0_) );
  AND2_X1 npu_inst_pe_1_2_2_U62 ( .A1(npu_inst_n58), .A2(npu_inst_pe_1_2_2_N94), .ZN(npu_inst_int_data_y_2__2__1_) );
  NOR3_X1 npu_inst_pe_1_2_2_U61 ( .A1(npu_inst_pe_1_2_2_n26), .A2(npu_inst_n58), .A3(npu_inst_int_ckg[45]), .ZN(npu_inst_pe_1_2_2_n85) );
  OR2_X1 npu_inst_pe_1_2_2_U60 ( .A1(npu_inst_pe_1_2_2_n85), .A2(
        npu_inst_pe_1_2_2_n2), .ZN(npu_inst_pe_1_2_2_N84) );
  AND2_X1 npu_inst_pe_1_2_2_U59 ( .A1(npu_inst_pe_1_2_2_int_q_acc_0_), .A2(
        npu_inst_pe_1_2_2_n1), .ZN(npu_inst_int_data_res_2__2__0_) );
  AND2_X1 npu_inst_pe_1_2_2_U58 ( .A1(npu_inst_pe_1_2_2_n2), .A2(
        npu_inst_pe_1_2_2_int_q_acc_7_), .ZN(npu_inst_int_data_res_2__2__7_)
         );
  AND2_X1 npu_inst_pe_1_2_2_U57 ( .A1(npu_inst_pe_1_2_2_int_q_acc_1_), .A2(
        npu_inst_pe_1_2_2_n1), .ZN(npu_inst_int_data_res_2__2__1_) );
  AND2_X1 npu_inst_pe_1_2_2_U56 ( .A1(npu_inst_pe_1_2_2_int_q_acc_2_), .A2(
        npu_inst_pe_1_2_2_n1), .ZN(npu_inst_int_data_res_2__2__2_) );
  AND2_X1 npu_inst_pe_1_2_2_U55 ( .A1(npu_inst_pe_1_2_2_int_q_acc_3_), .A2(
        npu_inst_pe_1_2_2_n2), .ZN(npu_inst_int_data_res_2__2__3_) );
  AND2_X1 npu_inst_pe_1_2_2_U54 ( .A1(npu_inst_pe_1_2_2_int_q_acc_4_), .A2(
        npu_inst_pe_1_2_2_n2), .ZN(npu_inst_int_data_res_2__2__4_) );
  AND2_X1 npu_inst_pe_1_2_2_U53 ( .A1(npu_inst_pe_1_2_2_int_q_acc_5_), .A2(
        npu_inst_pe_1_2_2_n2), .ZN(npu_inst_int_data_res_2__2__5_) );
  AND2_X1 npu_inst_pe_1_2_2_U52 ( .A1(npu_inst_pe_1_2_2_int_q_acc_6_), .A2(
        npu_inst_pe_1_2_2_n2), .ZN(npu_inst_int_data_res_2__2__6_) );
  AOI222_X1 npu_inst_pe_1_2_2_U51 ( .A1(npu_inst_int_data_res_3__2__0_), .A2(
        npu_inst_pe_1_2_2_n1), .B1(npu_inst_pe_1_2_2_N73), .B2(
        npu_inst_pe_1_2_2_n76), .C1(npu_inst_pe_1_2_2_N65), .C2(
        npu_inst_pe_1_2_2_n77), .ZN(npu_inst_pe_1_2_2_n84) );
  INV_X1 npu_inst_pe_1_2_2_U50 ( .A(npu_inst_pe_1_2_2_n84), .ZN(
        npu_inst_pe_1_2_2_n101) );
  AOI222_X1 npu_inst_pe_1_2_2_U49 ( .A1(npu_inst_int_data_res_3__2__7_), .A2(
        npu_inst_pe_1_2_2_n1), .B1(npu_inst_pe_1_2_2_N80), .B2(
        npu_inst_pe_1_2_2_n76), .C1(npu_inst_pe_1_2_2_N72), .C2(
        npu_inst_pe_1_2_2_n77), .ZN(npu_inst_pe_1_2_2_n75) );
  INV_X1 npu_inst_pe_1_2_2_U48 ( .A(npu_inst_pe_1_2_2_n75), .ZN(
        npu_inst_pe_1_2_2_n33) );
  AOI222_X1 npu_inst_pe_1_2_2_U47 ( .A1(npu_inst_int_data_res_3__2__1_), .A2(
        npu_inst_pe_1_2_2_n1), .B1(npu_inst_pe_1_2_2_N74), .B2(
        npu_inst_pe_1_2_2_n76), .C1(npu_inst_pe_1_2_2_N66), .C2(
        npu_inst_pe_1_2_2_n77), .ZN(npu_inst_pe_1_2_2_n83) );
  INV_X1 npu_inst_pe_1_2_2_U46 ( .A(npu_inst_pe_1_2_2_n83), .ZN(
        npu_inst_pe_1_2_2_n100) );
  AOI222_X1 npu_inst_pe_1_2_2_U45 ( .A1(npu_inst_int_data_res_3__2__2_), .A2(
        npu_inst_pe_1_2_2_n1), .B1(npu_inst_pe_1_2_2_N75), .B2(
        npu_inst_pe_1_2_2_n76), .C1(npu_inst_pe_1_2_2_N67), .C2(
        npu_inst_pe_1_2_2_n77), .ZN(npu_inst_pe_1_2_2_n82) );
  INV_X1 npu_inst_pe_1_2_2_U44 ( .A(npu_inst_pe_1_2_2_n82), .ZN(
        npu_inst_pe_1_2_2_n99) );
  AOI222_X1 npu_inst_pe_1_2_2_U43 ( .A1(npu_inst_int_data_res_3__2__3_), .A2(
        npu_inst_pe_1_2_2_n1), .B1(npu_inst_pe_1_2_2_N76), .B2(
        npu_inst_pe_1_2_2_n76), .C1(npu_inst_pe_1_2_2_N68), .C2(
        npu_inst_pe_1_2_2_n77), .ZN(npu_inst_pe_1_2_2_n81) );
  INV_X1 npu_inst_pe_1_2_2_U42 ( .A(npu_inst_pe_1_2_2_n81), .ZN(
        npu_inst_pe_1_2_2_n98) );
  AOI222_X1 npu_inst_pe_1_2_2_U41 ( .A1(npu_inst_int_data_res_3__2__4_), .A2(
        npu_inst_pe_1_2_2_n1), .B1(npu_inst_pe_1_2_2_N77), .B2(
        npu_inst_pe_1_2_2_n76), .C1(npu_inst_pe_1_2_2_N69), .C2(
        npu_inst_pe_1_2_2_n77), .ZN(npu_inst_pe_1_2_2_n80) );
  INV_X1 npu_inst_pe_1_2_2_U40 ( .A(npu_inst_pe_1_2_2_n80), .ZN(
        npu_inst_pe_1_2_2_n36) );
  AOI222_X1 npu_inst_pe_1_2_2_U39 ( .A1(npu_inst_int_data_res_3__2__5_), .A2(
        npu_inst_pe_1_2_2_n1), .B1(npu_inst_pe_1_2_2_N78), .B2(
        npu_inst_pe_1_2_2_n76), .C1(npu_inst_pe_1_2_2_N70), .C2(
        npu_inst_pe_1_2_2_n77), .ZN(npu_inst_pe_1_2_2_n79) );
  INV_X1 npu_inst_pe_1_2_2_U38 ( .A(npu_inst_pe_1_2_2_n79), .ZN(
        npu_inst_pe_1_2_2_n35) );
  AOI222_X1 npu_inst_pe_1_2_2_U37 ( .A1(npu_inst_int_data_res_3__2__6_), .A2(
        npu_inst_pe_1_2_2_n1), .B1(npu_inst_pe_1_2_2_N79), .B2(
        npu_inst_pe_1_2_2_n76), .C1(npu_inst_pe_1_2_2_N71), .C2(
        npu_inst_pe_1_2_2_n77), .ZN(npu_inst_pe_1_2_2_n78) );
  INV_X1 npu_inst_pe_1_2_2_U36 ( .A(npu_inst_pe_1_2_2_n78), .ZN(
        npu_inst_pe_1_2_2_n34) );
  INV_X1 npu_inst_pe_1_2_2_U35 ( .A(npu_inst_pe_1_2_2_int_data_1_), .ZN(
        npu_inst_pe_1_2_2_n14) );
  AND2_X1 npu_inst_pe_1_2_2_U34 ( .A1(npu_inst_int_data_x_2__2__1_), .A2(
        npu_inst_pe_1_2_2_int_q_weight_1_), .ZN(npu_inst_pe_1_2_2_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_2_2_U33 ( .A1(npu_inst_int_data_x_2__2__0_), .A2(
        npu_inst_pe_1_2_2_int_q_weight_1_), .ZN(npu_inst_pe_1_2_2_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_2_2_U32 ( .A1(npu_inst_n58), .A2(
        npu_inst_int_data_y_3__2__1_), .B1(npu_inst_pe_1_2_2_n3), .B2(
        npu_inst_int_data_x_2__3__1_), .ZN(npu_inst_pe_1_2_2_n63) );
  AOI22_X1 npu_inst_pe_1_2_2_U31 ( .A1(npu_inst_n58), .A2(
        npu_inst_int_data_y_3__2__0_), .B1(npu_inst_pe_1_2_2_n3), .B2(
        npu_inst_int_data_x_2__3__0_), .ZN(npu_inst_pe_1_2_2_n61) );
  INV_X1 npu_inst_pe_1_2_2_U30 ( .A(npu_inst_pe_1_2_2_int_data_0_), .ZN(
        npu_inst_pe_1_2_2_n13) );
  INV_X1 npu_inst_pe_1_2_2_U29 ( .A(npu_inst_n70), .ZN(npu_inst_pe_1_2_2_n5)
         );
  OR3_X1 npu_inst_pe_1_2_2_U28 ( .A1(npu_inst_pe_1_2_2_n6), .A2(
        npu_inst_pe_1_2_2_n8), .A3(npu_inst_pe_1_2_2_n5), .ZN(
        npu_inst_pe_1_2_2_n56) );
  OR3_X1 npu_inst_pe_1_2_2_U27 ( .A1(npu_inst_pe_1_2_2_n5), .A2(
        npu_inst_pe_1_2_2_n8), .A3(npu_inst_pe_1_2_2_n7), .ZN(
        npu_inst_pe_1_2_2_n48) );
  INV_X1 npu_inst_pe_1_2_2_U26 ( .A(npu_inst_pe_1_2_2_n5), .ZN(
        npu_inst_pe_1_2_2_n4) );
  OR3_X1 npu_inst_pe_1_2_2_U25 ( .A1(npu_inst_pe_1_2_2_n4), .A2(
        npu_inst_pe_1_2_2_n8), .A3(npu_inst_pe_1_2_2_n7), .ZN(
        npu_inst_pe_1_2_2_n52) );
  OR3_X1 npu_inst_pe_1_2_2_U24 ( .A1(npu_inst_pe_1_2_2_n6), .A2(
        npu_inst_pe_1_2_2_n8), .A3(npu_inst_pe_1_2_2_n4), .ZN(
        npu_inst_pe_1_2_2_n60) );
  NOR2_X1 npu_inst_pe_1_2_2_U23 ( .A1(npu_inst_pe_1_2_2_n60), .A2(
        npu_inst_pe_1_2_2_n3), .ZN(npu_inst_pe_1_2_2_n58) );
  NOR2_X1 npu_inst_pe_1_2_2_U22 ( .A1(npu_inst_pe_1_2_2_n56), .A2(
        npu_inst_pe_1_2_2_n3), .ZN(npu_inst_pe_1_2_2_n54) );
  NOR2_X1 npu_inst_pe_1_2_2_U21 ( .A1(npu_inst_pe_1_2_2_n52), .A2(
        npu_inst_pe_1_2_2_n3), .ZN(npu_inst_pe_1_2_2_n50) );
  NOR2_X1 npu_inst_pe_1_2_2_U20 ( .A1(npu_inst_pe_1_2_2_n48), .A2(
        npu_inst_pe_1_2_2_n3), .ZN(npu_inst_pe_1_2_2_n46) );
  NOR2_X1 npu_inst_pe_1_2_2_U19 ( .A1(npu_inst_pe_1_2_2_n40), .A2(
        npu_inst_pe_1_2_2_n3), .ZN(npu_inst_pe_1_2_2_n38) );
  NOR2_X1 npu_inst_pe_1_2_2_U18 ( .A1(npu_inst_pe_1_2_2_n44), .A2(
        npu_inst_pe_1_2_2_n3), .ZN(npu_inst_pe_1_2_2_n42) );
  BUF_X1 npu_inst_pe_1_2_2_U17 ( .A(npu_inst_n103), .Z(npu_inst_pe_1_2_2_n8)
         );
  INV_X1 npu_inst_pe_1_2_2_U16 ( .A(npu_inst_n125), .ZN(npu_inst_pe_1_2_2_n12)
         );
  INV_X1 npu_inst_pe_1_2_2_U15 ( .A(npu_inst_pe_1_2_2_n38), .ZN(
        npu_inst_pe_1_2_2_n114) );
  INV_X1 npu_inst_pe_1_2_2_U14 ( .A(npu_inst_pe_1_2_2_n58), .ZN(
        npu_inst_pe_1_2_2_n119) );
  INV_X1 npu_inst_pe_1_2_2_U13 ( .A(npu_inst_pe_1_2_2_n54), .ZN(
        npu_inst_pe_1_2_2_n118) );
  INV_X1 npu_inst_pe_1_2_2_U12 ( .A(npu_inst_pe_1_2_2_n50), .ZN(
        npu_inst_pe_1_2_2_n117) );
  INV_X1 npu_inst_pe_1_2_2_U11 ( .A(npu_inst_pe_1_2_2_n46), .ZN(
        npu_inst_pe_1_2_2_n116) );
  INV_X1 npu_inst_pe_1_2_2_U10 ( .A(npu_inst_pe_1_2_2_n42), .ZN(
        npu_inst_pe_1_2_2_n115) );
  BUF_X1 npu_inst_pe_1_2_2_U9 ( .A(npu_inst_n29), .Z(npu_inst_pe_1_2_2_n2) );
  BUF_X1 npu_inst_pe_1_2_2_U8 ( .A(npu_inst_n29), .Z(npu_inst_pe_1_2_2_n1) );
  BUF_X1 npu_inst_pe_1_2_2_U7 ( .A(npu_inst_pe_1_2_2_n12), .Z(
        npu_inst_pe_1_2_2_n11) );
  BUF_X1 npu_inst_pe_1_2_2_U6 ( .A(npu_inst_pe_1_2_2_n12), .Z(
        npu_inst_pe_1_2_2_n10) );
  BUF_X1 npu_inst_pe_1_2_2_U5 ( .A(npu_inst_pe_1_2_2_n12), .Z(
        npu_inst_pe_1_2_2_n9) );
  NOR2_X1 npu_inst_pe_1_2_2_U4 ( .A1(npu_inst_pe_1_2_2_int_q_weight_0_), .A2(
        npu_inst_pe_1_2_2_n1), .ZN(npu_inst_pe_1_2_2_n76) );
  NOR2_X1 npu_inst_pe_1_2_2_U3 ( .A1(npu_inst_pe_1_2_2_n27), .A2(
        npu_inst_pe_1_2_2_n1), .ZN(npu_inst_pe_1_2_2_n77) );
  FA_X1 npu_inst_pe_1_2_2_sub_67_U2_1 ( .A(npu_inst_pe_1_2_2_int_q_acc_1_), 
        .B(npu_inst_pe_1_2_2_n14), .CI(npu_inst_pe_1_2_2_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_2_2_sub_67_carry_2_), .S(npu_inst_pe_1_2_2_N66) );
  FA_X1 npu_inst_pe_1_2_2_add_69_U1_1 ( .A(npu_inst_pe_1_2_2_int_q_acc_1_), 
        .B(npu_inst_pe_1_2_2_int_data_1_), .CI(
        npu_inst_pe_1_2_2_add_69_carry_1_), .CO(
        npu_inst_pe_1_2_2_add_69_carry_2_), .S(npu_inst_pe_1_2_2_N74) );
  NAND3_X1 npu_inst_pe_1_2_2_U109 ( .A1(npu_inst_pe_1_2_2_n5), .A2(
        npu_inst_pe_1_2_2_n7), .A3(npu_inst_pe_1_2_2_n8), .ZN(
        npu_inst_pe_1_2_2_n44) );
  NAND3_X1 npu_inst_pe_1_2_2_U108 ( .A1(npu_inst_pe_1_2_2_n4), .A2(
        npu_inst_pe_1_2_2_n7), .A3(npu_inst_pe_1_2_2_n8), .ZN(
        npu_inst_pe_1_2_2_n40) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_2_2_n34), .CK(
        npu_inst_pe_1_2_2_net4148), .RN(npu_inst_pe_1_2_2_n9), .Q(
        npu_inst_pe_1_2_2_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_2_2_n35), .CK(
        npu_inst_pe_1_2_2_net4148), .RN(npu_inst_pe_1_2_2_n9), .Q(
        npu_inst_pe_1_2_2_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_2_2_n36), .CK(
        npu_inst_pe_1_2_2_net4148), .RN(npu_inst_pe_1_2_2_n9), .Q(
        npu_inst_pe_1_2_2_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_2_2_n98), .CK(
        npu_inst_pe_1_2_2_net4148), .RN(npu_inst_pe_1_2_2_n9), .Q(
        npu_inst_pe_1_2_2_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_2_2_n99), .CK(
        npu_inst_pe_1_2_2_net4148), .RN(npu_inst_pe_1_2_2_n9), .Q(
        npu_inst_pe_1_2_2_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_2_2_n100), 
        .CK(npu_inst_pe_1_2_2_net4148), .RN(npu_inst_pe_1_2_2_n9), .Q(
        npu_inst_pe_1_2_2_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_2_2_n33), .CK(
        npu_inst_pe_1_2_2_net4148), .RN(npu_inst_pe_1_2_2_n9), .Q(
        npu_inst_pe_1_2_2_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_2_2_n101), 
        .CK(npu_inst_pe_1_2_2_net4148), .RN(npu_inst_pe_1_2_2_n9), .Q(
        npu_inst_pe_1_2_2_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_weight_reg_0_ ( .D(npu_inst_n111), .CK(
        npu_inst_pe_1_2_2_net4154), .RN(npu_inst_pe_1_2_2_n9), .Q(
        npu_inst_pe_1_2_2_int_q_weight_0_), .QN(npu_inst_pe_1_2_2_n27) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_weight_reg_1_ ( .D(npu_inst_n117), .CK(
        npu_inst_pe_1_2_2_net4154), .RN(npu_inst_pe_1_2_2_n9), .Q(
        npu_inst_pe_1_2_2_int_q_weight_1_), .QN(npu_inst_pe_1_2_2_n26) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_2_2_n113), 
        .CK(npu_inst_pe_1_2_2_net4154), .RN(npu_inst_pe_1_2_2_n9), .Q(
        npu_inst_pe_1_2_2_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_2_2_n107), 
        .CK(npu_inst_pe_1_2_2_net4154), .RN(npu_inst_pe_1_2_2_n9), .Q(
        npu_inst_pe_1_2_2_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_2_2_n112), 
        .CK(npu_inst_pe_1_2_2_net4154), .RN(npu_inst_pe_1_2_2_n10), .Q(
        npu_inst_pe_1_2_2_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_2_2_n106), 
        .CK(npu_inst_pe_1_2_2_net4154), .RN(npu_inst_pe_1_2_2_n10), .Q(
        npu_inst_pe_1_2_2_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_2_2_n111), 
        .CK(npu_inst_pe_1_2_2_net4154), .RN(npu_inst_pe_1_2_2_n10), .Q(
        npu_inst_pe_1_2_2_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_2_2_n105), 
        .CK(npu_inst_pe_1_2_2_net4154), .RN(npu_inst_pe_1_2_2_n10), .Q(
        npu_inst_pe_1_2_2_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_2_2_n110), 
        .CK(npu_inst_pe_1_2_2_net4154), .RN(npu_inst_pe_1_2_2_n10), .Q(
        npu_inst_pe_1_2_2_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_2_2_n104), 
        .CK(npu_inst_pe_1_2_2_net4154), .RN(npu_inst_pe_1_2_2_n10), .Q(
        npu_inst_pe_1_2_2_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_2_2_n109), 
        .CK(npu_inst_pe_1_2_2_net4154), .RN(npu_inst_pe_1_2_2_n10), .Q(
        npu_inst_pe_1_2_2_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_2_2_n103), 
        .CK(npu_inst_pe_1_2_2_net4154), .RN(npu_inst_pe_1_2_2_n10), .Q(
        npu_inst_pe_1_2_2_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_2_2_n108), 
        .CK(npu_inst_pe_1_2_2_net4154), .RN(npu_inst_pe_1_2_2_n10), .Q(
        npu_inst_pe_1_2_2_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_2_2_n102), 
        .CK(npu_inst_pe_1_2_2_net4154), .RN(npu_inst_pe_1_2_2_n10), .Q(
        npu_inst_pe_1_2_2_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_2_2_n86), 
        .CK(npu_inst_pe_1_2_2_net4154), .RN(npu_inst_pe_1_2_2_n10), .Q(
        npu_inst_pe_1_2_2_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_2_2_n87), 
        .CK(npu_inst_pe_1_2_2_net4154), .RN(npu_inst_pe_1_2_2_n10), .Q(
        npu_inst_pe_1_2_2_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_2_2_n88), 
        .CK(npu_inst_pe_1_2_2_net4154), .RN(npu_inst_pe_1_2_2_n11), .Q(
        npu_inst_pe_1_2_2_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_2_2_n89), 
        .CK(npu_inst_pe_1_2_2_net4154), .RN(npu_inst_pe_1_2_2_n11), .Q(
        npu_inst_pe_1_2_2_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_2_2_n90), 
        .CK(npu_inst_pe_1_2_2_net4154), .RN(npu_inst_pe_1_2_2_n11), .Q(
        npu_inst_pe_1_2_2_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_2_2_n91), 
        .CK(npu_inst_pe_1_2_2_net4154), .RN(npu_inst_pe_1_2_2_n11), .Q(
        npu_inst_pe_1_2_2_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_2_2_n92), 
        .CK(npu_inst_pe_1_2_2_net4154), .RN(npu_inst_pe_1_2_2_n11), .Q(
        npu_inst_pe_1_2_2_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_2_2_n93), 
        .CK(npu_inst_pe_1_2_2_net4154), .RN(npu_inst_pe_1_2_2_n11), .Q(
        npu_inst_pe_1_2_2_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_2_2_n94), 
        .CK(npu_inst_pe_1_2_2_net4154), .RN(npu_inst_pe_1_2_2_n11), .Q(
        npu_inst_pe_1_2_2_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_2_2_n95), 
        .CK(npu_inst_pe_1_2_2_net4154), .RN(npu_inst_pe_1_2_2_n11), .Q(
        npu_inst_pe_1_2_2_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_2_2_n96), 
        .CK(npu_inst_pe_1_2_2_net4154), .RN(npu_inst_pe_1_2_2_n11), .Q(
        npu_inst_pe_1_2_2_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_2_2_n97), 
        .CK(npu_inst_pe_1_2_2_net4154), .RN(npu_inst_pe_1_2_2_n11), .Q(
        npu_inst_pe_1_2_2_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_2_2_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_2_2_N84), .SE(1'b0), .GCK(npu_inst_pe_1_2_2_net4148) );
  CLKGATETST_X1 npu_inst_pe_1_2_2_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n65), .SE(1'b0), .GCK(npu_inst_pe_1_2_2_net4154) );
  MUX2_X1 npu_inst_pe_1_2_3_U162 ( .A(npu_inst_pe_1_2_3_n32), .B(
        npu_inst_pe_1_2_3_n29), .S(npu_inst_pe_1_2_3_n8), .Z(
        npu_inst_pe_1_2_3_N93) );
  MUX2_X1 npu_inst_pe_1_2_3_U161 ( .A(npu_inst_pe_1_2_3_n31), .B(
        npu_inst_pe_1_2_3_n30), .S(npu_inst_pe_1_2_3_n6), .Z(
        npu_inst_pe_1_2_3_n32) );
  MUX2_X1 npu_inst_pe_1_2_3_U160 ( .A(npu_inst_pe_1_2_3_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_2_3_int_q_reg_v_1__0_), .S(npu_inst_pe_1_2_3_n4), .Z(
        npu_inst_pe_1_2_3_n31) );
  MUX2_X1 npu_inst_pe_1_2_3_U159 ( .A(npu_inst_pe_1_2_3_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_2_3_int_q_reg_v_3__0_), .S(npu_inst_pe_1_2_3_n4), .Z(
        npu_inst_pe_1_2_3_n30) );
  MUX2_X1 npu_inst_pe_1_2_3_U158 ( .A(npu_inst_pe_1_2_3_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_2_3_int_q_reg_v_5__0_), .S(npu_inst_pe_1_2_3_n4), .Z(
        npu_inst_pe_1_2_3_n29) );
  MUX2_X1 npu_inst_pe_1_2_3_U157 ( .A(npu_inst_pe_1_2_3_n28), .B(
        npu_inst_pe_1_2_3_n23), .S(npu_inst_pe_1_2_3_n8), .Z(
        npu_inst_pe_1_2_3_N94) );
  MUX2_X1 npu_inst_pe_1_2_3_U156 ( .A(npu_inst_pe_1_2_3_n25), .B(
        npu_inst_pe_1_2_3_n24), .S(npu_inst_pe_1_2_3_n6), .Z(
        npu_inst_pe_1_2_3_n28) );
  MUX2_X1 npu_inst_pe_1_2_3_U155 ( .A(npu_inst_pe_1_2_3_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_2_3_int_q_reg_v_1__1_), .S(npu_inst_pe_1_2_3_n4), .Z(
        npu_inst_pe_1_2_3_n25) );
  MUX2_X1 npu_inst_pe_1_2_3_U154 ( .A(npu_inst_pe_1_2_3_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_2_3_int_q_reg_v_3__1_), .S(npu_inst_pe_1_2_3_n4), .Z(
        npu_inst_pe_1_2_3_n24) );
  MUX2_X1 npu_inst_pe_1_2_3_U153 ( .A(npu_inst_pe_1_2_3_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_2_3_int_q_reg_v_5__1_), .S(npu_inst_pe_1_2_3_n4), .Z(
        npu_inst_pe_1_2_3_n23) );
  MUX2_X1 npu_inst_pe_1_2_3_U152 ( .A(npu_inst_pe_1_2_3_n22), .B(
        npu_inst_pe_1_2_3_n19), .S(npu_inst_pe_1_2_3_n8), .Z(
        npu_inst_int_data_x_2__3__1_) );
  MUX2_X1 npu_inst_pe_1_2_3_U151 ( .A(npu_inst_pe_1_2_3_n21), .B(
        npu_inst_pe_1_2_3_n20), .S(npu_inst_pe_1_2_3_n6), .Z(
        npu_inst_pe_1_2_3_n22) );
  MUX2_X1 npu_inst_pe_1_2_3_U150 ( .A(npu_inst_pe_1_2_3_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_2_3_int_q_reg_h_1__1_), .S(npu_inst_pe_1_2_3_n4), .Z(
        npu_inst_pe_1_2_3_n21) );
  MUX2_X1 npu_inst_pe_1_2_3_U149 ( .A(npu_inst_pe_1_2_3_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_2_3_int_q_reg_h_3__1_), .S(npu_inst_pe_1_2_3_n4), .Z(
        npu_inst_pe_1_2_3_n20) );
  MUX2_X1 npu_inst_pe_1_2_3_U148 ( .A(npu_inst_pe_1_2_3_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_2_3_int_q_reg_h_5__1_), .S(npu_inst_pe_1_2_3_n4), .Z(
        npu_inst_pe_1_2_3_n19) );
  MUX2_X1 npu_inst_pe_1_2_3_U147 ( .A(npu_inst_pe_1_2_3_n18), .B(
        npu_inst_pe_1_2_3_n15), .S(npu_inst_pe_1_2_3_n8), .Z(
        npu_inst_int_data_x_2__3__0_) );
  MUX2_X1 npu_inst_pe_1_2_3_U146 ( .A(npu_inst_pe_1_2_3_n17), .B(
        npu_inst_pe_1_2_3_n16), .S(npu_inst_pe_1_2_3_n6), .Z(
        npu_inst_pe_1_2_3_n18) );
  MUX2_X1 npu_inst_pe_1_2_3_U145 ( .A(npu_inst_pe_1_2_3_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_2_3_int_q_reg_h_1__0_), .S(npu_inst_pe_1_2_3_n4), .Z(
        npu_inst_pe_1_2_3_n17) );
  MUX2_X1 npu_inst_pe_1_2_3_U144 ( .A(npu_inst_pe_1_2_3_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_2_3_int_q_reg_h_3__0_), .S(npu_inst_pe_1_2_3_n4), .Z(
        npu_inst_pe_1_2_3_n16) );
  MUX2_X1 npu_inst_pe_1_2_3_U143 ( .A(npu_inst_pe_1_2_3_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_2_3_int_q_reg_h_5__0_), .S(npu_inst_pe_1_2_3_n4), .Z(
        npu_inst_pe_1_2_3_n15) );
  XOR2_X1 npu_inst_pe_1_2_3_U142 ( .A(npu_inst_pe_1_2_3_int_data_0_), .B(
        npu_inst_pe_1_2_3_int_q_acc_0_), .Z(npu_inst_pe_1_2_3_N73) );
  AND2_X1 npu_inst_pe_1_2_3_U141 ( .A1(npu_inst_pe_1_2_3_int_q_acc_0_), .A2(
        npu_inst_pe_1_2_3_int_data_0_), .ZN(npu_inst_pe_1_2_3_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_2_3_U140 ( .A(npu_inst_pe_1_2_3_int_q_acc_0_), .B(
        npu_inst_pe_1_2_3_n13), .ZN(npu_inst_pe_1_2_3_N65) );
  OR2_X1 npu_inst_pe_1_2_3_U139 ( .A1(npu_inst_pe_1_2_3_n13), .A2(
        npu_inst_pe_1_2_3_int_q_acc_0_), .ZN(npu_inst_pe_1_2_3_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_2_3_U138 ( .A(npu_inst_pe_1_2_3_int_q_acc_2_), .B(
        npu_inst_pe_1_2_3_add_69_carry_2_), .Z(npu_inst_pe_1_2_3_N75) );
  AND2_X1 npu_inst_pe_1_2_3_U137 ( .A1(npu_inst_pe_1_2_3_add_69_carry_2_), 
        .A2(npu_inst_pe_1_2_3_int_q_acc_2_), .ZN(
        npu_inst_pe_1_2_3_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_2_3_U136 ( .A(npu_inst_pe_1_2_3_int_q_acc_3_), .B(
        npu_inst_pe_1_2_3_add_69_carry_3_), .Z(npu_inst_pe_1_2_3_N76) );
  AND2_X1 npu_inst_pe_1_2_3_U135 ( .A1(npu_inst_pe_1_2_3_add_69_carry_3_), 
        .A2(npu_inst_pe_1_2_3_int_q_acc_3_), .ZN(
        npu_inst_pe_1_2_3_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_2_3_U134 ( .A(npu_inst_pe_1_2_3_int_q_acc_4_), .B(
        npu_inst_pe_1_2_3_add_69_carry_4_), .Z(npu_inst_pe_1_2_3_N77) );
  AND2_X1 npu_inst_pe_1_2_3_U133 ( .A1(npu_inst_pe_1_2_3_add_69_carry_4_), 
        .A2(npu_inst_pe_1_2_3_int_q_acc_4_), .ZN(
        npu_inst_pe_1_2_3_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_2_3_U132 ( .A(npu_inst_pe_1_2_3_int_q_acc_5_), .B(
        npu_inst_pe_1_2_3_add_69_carry_5_), .Z(npu_inst_pe_1_2_3_N78) );
  AND2_X1 npu_inst_pe_1_2_3_U131 ( .A1(npu_inst_pe_1_2_3_add_69_carry_5_), 
        .A2(npu_inst_pe_1_2_3_int_q_acc_5_), .ZN(
        npu_inst_pe_1_2_3_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_2_3_U130 ( .A(npu_inst_pe_1_2_3_int_q_acc_6_), .B(
        npu_inst_pe_1_2_3_add_69_carry_6_), .Z(npu_inst_pe_1_2_3_N79) );
  AND2_X1 npu_inst_pe_1_2_3_U129 ( .A1(npu_inst_pe_1_2_3_add_69_carry_6_), 
        .A2(npu_inst_pe_1_2_3_int_q_acc_6_), .ZN(
        npu_inst_pe_1_2_3_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_2_3_U128 ( .A(npu_inst_pe_1_2_3_int_q_acc_7_), .B(
        npu_inst_pe_1_2_3_add_69_carry_7_), .Z(npu_inst_pe_1_2_3_N80) );
  XNOR2_X1 npu_inst_pe_1_2_3_U127 ( .A(npu_inst_pe_1_2_3_sub_67_carry_2_), .B(
        npu_inst_pe_1_2_3_int_q_acc_2_), .ZN(npu_inst_pe_1_2_3_N67) );
  OR2_X1 npu_inst_pe_1_2_3_U126 ( .A1(npu_inst_pe_1_2_3_int_q_acc_2_), .A2(
        npu_inst_pe_1_2_3_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_2_3_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_2_3_U125 ( .A(npu_inst_pe_1_2_3_sub_67_carry_3_), .B(
        npu_inst_pe_1_2_3_int_q_acc_3_), .ZN(npu_inst_pe_1_2_3_N68) );
  OR2_X1 npu_inst_pe_1_2_3_U124 ( .A1(npu_inst_pe_1_2_3_int_q_acc_3_), .A2(
        npu_inst_pe_1_2_3_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_2_3_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_2_3_U123 ( .A(npu_inst_pe_1_2_3_sub_67_carry_4_), .B(
        npu_inst_pe_1_2_3_int_q_acc_4_), .ZN(npu_inst_pe_1_2_3_N69) );
  OR2_X1 npu_inst_pe_1_2_3_U122 ( .A1(npu_inst_pe_1_2_3_int_q_acc_4_), .A2(
        npu_inst_pe_1_2_3_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_2_3_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_2_3_U121 ( .A(npu_inst_pe_1_2_3_sub_67_carry_5_), .B(
        npu_inst_pe_1_2_3_int_q_acc_5_), .ZN(npu_inst_pe_1_2_3_N70) );
  OR2_X1 npu_inst_pe_1_2_3_U120 ( .A1(npu_inst_pe_1_2_3_int_q_acc_5_), .A2(
        npu_inst_pe_1_2_3_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_2_3_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_2_3_U119 ( .A(npu_inst_pe_1_2_3_sub_67_carry_6_), .B(
        npu_inst_pe_1_2_3_int_q_acc_6_), .ZN(npu_inst_pe_1_2_3_N71) );
  OR2_X1 npu_inst_pe_1_2_3_U118 ( .A1(npu_inst_pe_1_2_3_int_q_acc_6_), .A2(
        npu_inst_pe_1_2_3_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_2_3_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_2_3_U117 ( .A(npu_inst_pe_1_2_3_int_q_acc_7_), .B(
        npu_inst_pe_1_2_3_sub_67_carry_7_), .ZN(npu_inst_pe_1_2_3_N72) );
  INV_X1 npu_inst_pe_1_2_3_U116 ( .A(npu_inst_n78), .ZN(npu_inst_pe_1_2_3_n7)
         );
  INV_X1 npu_inst_pe_1_2_3_U115 ( .A(npu_inst_pe_1_2_3_n7), .ZN(
        npu_inst_pe_1_2_3_n6) );
  INV_X1 npu_inst_pe_1_2_3_U114 ( .A(npu_inst_n58), .ZN(npu_inst_pe_1_2_3_n3)
         );
  AOI22_X1 npu_inst_pe_1_2_3_U113 ( .A1(npu_inst_int_data_y_3__3__0_), .A2(
        npu_inst_pe_1_2_3_n58), .B1(npu_inst_pe_1_2_3_n119), .B2(
        npu_inst_pe_1_2_3_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_2_3_n57) );
  INV_X1 npu_inst_pe_1_2_3_U112 ( .A(npu_inst_pe_1_2_3_n57), .ZN(
        npu_inst_pe_1_2_3_n108) );
  AOI22_X1 npu_inst_pe_1_2_3_U111 ( .A1(npu_inst_int_data_y_3__3__0_), .A2(
        npu_inst_pe_1_2_3_n54), .B1(npu_inst_pe_1_2_3_n118), .B2(
        npu_inst_pe_1_2_3_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_2_3_n53) );
  INV_X1 npu_inst_pe_1_2_3_U110 ( .A(npu_inst_pe_1_2_3_n53), .ZN(
        npu_inst_pe_1_2_3_n109) );
  AOI22_X1 npu_inst_pe_1_2_3_U107 ( .A1(npu_inst_int_data_y_3__3__0_), .A2(
        npu_inst_pe_1_2_3_n50), .B1(npu_inst_pe_1_2_3_n117), .B2(
        npu_inst_pe_1_2_3_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_2_3_n49) );
  INV_X1 npu_inst_pe_1_2_3_U106 ( .A(npu_inst_pe_1_2_3_n49), .ZN(
        npu_inst_pe_1_2_3_n110) );
  AOI22_X1 npu_inst_pe_1_2_3_U105 ( .A1(npu_inst_int_data_y_3__3__0_), .A2(
        npu_inst_pe_1_2_3_n46), .B1(npu_inst_pe_1_2_3_n116), .B2(
        npu_inst_pe_1_2_3_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_2_3_n45) );
  INV_X1 npu_inst_pe_1_2_3_U104 ( .A(npu_inst_pe_1_2_3_n45), .ZN(
        npu_inst_pe_1_2_3_n111) );
  AOI22_X1 npu_inst_pe_1_2_3_U103 ( .A1(npu_inst_int_data_y_3__3__0_), .A2(
        npu_inst_pe_1_2_3_n42), .B1(npu_inst_pe_1_2_3_n115), .B2(
        npu_inst_pe_1_2_3_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_2_3_n41) );
  INV_X1 npu_inst_pe_1_2_3_U102 ( .A(npu_inst_pe_1_2_3_n41), .ZN(
        npu_inst_pe_1_2_3_n112) );
  AOI22_X1 npu_inst_pe_1_2_3_U101 ( .A1(npu_inst_int_data_y_3__3__1_), .A2(
        npu_inst_pe_1_2_3_n58), .B1(npu_inst_pe_1_2_3_n119), .B2(
        npu_inst_pe_1_2_3_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_2_3_n59) );
  INV_X1 npu_inst_pe_1_2_3_U100 ( .A(npu_inst_pe_1_2_3_n59), .ZN(
        npu_inst_pe_1_2_3_n102) );
  AOI22_X1 npu_inst_pe_1_2_3_U99 ( .A1(npu_inst_int_data_y_3__3__1_), .A2(
        npu_inst_pe_1_2_3_n54), .B1(npu_inst_pe_1_2_3_n118), .B2(
        npu_inst_pe_1_2_3_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_2_3_n55) );
  INV_X1 npu_inst_pe_1_2_3_U98 ( .A(npu_inst_pe_1_2_3_n55), .ZN(
        npu_inst_pe_1_2_3_n103) );
  AOI22_X1 npu_inst_pe_1_2_3_U97 ( .A1(npu_inst_int_data_y_3__3__1_), .A2(
        npu_inst_pe_1_2_3_n50), .B1(npu_inst_pe_1_2_3_n117), .B2(
        npu_inst_pe_1_2_3_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_2_3_n51) );
  INV_X1 npu_inst_pe_1_2_3_U96 ( .A(npu_inst_pe_1_2_3_n51), .ZN(
        npu_inst_pe_1_2_3_n104) );
  AOI22_X1 npu_inst_pe_1_2_3_U95 ( .A1(npu_inst_int_data_y_3__3__1_), .A2(
        npu_inst_pe_1_2_3_n46), .B1(npu_inst_pe_1_2_3_n116), .B2(
        npu_inst_pe_1_2_3_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_2_3_n47) );
  INV_X1 npu_inst_pe_1_2_3_U94 ( .A(npu_inst_pe_1_2_3_n47), .ZN(
        npu_inst_pe_1_2_3_n105) );
  AOI22_X1 npu_inst_pe_1_2_3_U93 ( .A1(npu_inst_int_data_y_3__3__1_), .A2(
        npu_inst_pe_1_2_3_n42), .B1(npu_inst_pe_1_2_3_n115), .B2(
        npu_inst_pe_1_2_3_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_2_3_n43) );
  INV_X1 npu_inst_pe_1_2_3_U92 ( .A(npu_inst_pe_1_2_3_n43), .ZN(
        npu_inst_pe_1_2_3_n106) );
  AOI22_X1 npu_inst_pe_1_2_3_U91 ( .A1(npu_inst_pe_1_2_3_n38), .A2(
        npu_inst_int_data_y_3__3__1_), .B1(npu_inst_pe_1_2_3_n114), .B2(
        npu_inst_pe_1_2_3_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_2_3_n39) );
  INV_X1 npu_inst_pe_1_2_3_U90 ( .A(npu_inst_pe_1_2_3_n39), .ZN(
        npu_inst_pe_1_2_3_n107) );
  AOI22_X1 npu_inst_pe_1_2_3_U89 ( .A1(npu_inst_pe_1_2_3_n38), .A2(
        npu_inst_int_data_y_3__3__0_), .B1(npu_inst_pe_1_2_3_n114), .B2(
        npu_inst_pe_1_2_3_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_2_3_n37) );
  INV_X1 npu_inst_pe_1_2_3_U88 ( .A(npu_inst_pe_1_2_3_n37), .ZN(
        npu_inst_pe_1_2_3_n113) );
  NAND2_X1 npu_inst_pe_1_2_3_U87 ( .A1(npu_inst_pe_1_2_3_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_2_3_n60), .ZN(npu_inst_pe_1_2_3_n74) );
  OAI21_X1 npu_inst_pe_1_2_3_U86 ( .B1(npu_inst_pe_1_2_3_n63), .B2(
        npu_inst_pe_1_2_3_n60), .A(npu_inst_pe_1_2_3_n74), .ZN(
        npu_inst_pe_1_2_3_n97) );
  NAND2_X1 npu_inst_pe_1_2_3_U85 ( .A1(npu_inst_pe_1_2_3_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_2_3_n60), .ZN(npu_inst_pe_1_2_3_n73) );
  OAI21_X1 npu_inst_pe_1_2_3_U84 ( .B1(npu_inst_pe_1_2_3_n61), .B2(
        npu_inst_pe_1_2_3_n60), .A(npu_inst_pe_1_2_3_n73), .ZN(
        npu_inst_pe_1_2_3_n96) );
  NAND2_X1 npu_inst_pe_1_2_3_U83 ( .A1(npu_inst_pe_1_2_3_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_2_3_n56), .ZN(npu_inst_pe_1_2_3_n72) );
  OAI21_X1 npu_inst_pe_1_2_3_U82 ( .B1(npu_inst_pe_1_2_3_n63), .B2(
        npu_inst_pe_1_2_3_n56), .A(npu_inst_pe_1_2_3_n72), .ZN(
        npu_inst_pe_1_2_3_n95) );
  NAND2_X1 npu_inst_pe_1_2_3_U81 ( .A1(npu_inst_pe_1_2_3_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_2_3_n56), .ZN(npu_inst_pe_1_2_3_n71) );
  OAI21_X1 npu_inst_pe_1_2_3_U80 ( .B1(npu_inst_pe_1_2_3_n61), .B2(
        npu_inst_pe_1_2_3_n56), .A(npu_inst_pe_1_2_3_n71), .ZN(
        npu_inst_pe_1_2_3_n94) );
  NAND2_X1 npu_inst_pe_1_2_3_U79 ( .A1(npu_inst_pe_1_2_3_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_2_3_n52), .ZN(npu_inst_pe_1_2_3_n70) );
  OAI21_X1 npu_inst_pe_1_2_3_U78 ( .B1(npu_inst_pe_1_2_3_n63), .B2(
        npu_inst_pe_1_2_3_n52), .A(npu_inst_pe_1_2_3_n70), .ZN(
        npu_inst_pe_1_2_3_n93) );
  NAND2_X1 npu_inst_pe_1_2_3_U77 ( .A1(npu_inst_pe_1_2_3_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_2_3_n52), .ZN(npu_inst_pe_1_2_3_n69) );
  OAI21_X1 npu_inst_pe_1_2_3_U76 ( .B1(npu_inst_pe_1_2_3_n61), .B2(
        npu_inst_pe_1_2_3_n52), .A(npu_inst_pe_1_2_3_n69), .ZN(
        npu_inst_pe_1_2_3_n92) );
  NAND2_X1 npu_inst_pe_1_2_3_U75 ( .A1(npu_inst_pe_1_2_3_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_2_3_n48), .ZN(npu_inst_pe_1_2_3_n68) );
  OAI21_X1 npu_inst_pe_1_2_3_U74 ( .B1(npu_inst_pe_1_2_3_n63), .B2(
        npu_inst_pe_1_2_3_n48), .A(npu_inst_pe_1_2_3_n68), .ZN(
        npu_inst_pe_1_2_3_n91) );
  NAND2_X1 npu_inst_pe_1_2_3_U73 ( .A1(npu_inst_pe_1_2_3_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_2_3_n48), .ZN(npu_inst_pe_1_2_3_n67) );
  OAI21_X1 npu_inst_pe_1_2_3_U72 ( .B1(npu_inst_pe_1_2_3_n61), .B2(
        npu_inst_pe_1_2_3_n48), .A(npu_inst_pe_1_2_3_n67), .ZN(
        npu_inst_pe_1_2_3_n90) );
  NAND2_X1 npu_inst_pe_1_2_3_U71 ( .A1(npu_inst_pe_1_2_3_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_2_3_n44), .ZN(npu_inst_pe_1_2_3_n66) );
  OAI21_X1 npu_inst_pe_1_2_3_U70 ( .B1(npu_inst_pe_1_2_3_n63), .B2(
        npu_inst_pe_1_2_3_n44), .A(npu_inst_pe_1_2_3_n66), .ZN(
        npu_inst_pe_1_2_3_n89) );
  NAND2_X1 npu_inst_pe_1_2_3_U69 ( .A1(npu_inst_pe_1_2_3_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_2_3_n44), .ZN(npu_inst_pe_1_2_3_n65) );
  OAI21_X1 npu_inst_pe_1_2_3_U68 ( .B1(npu_inst_pe_1_2_3_n61), .B2(
        npu_inst_pe_1_2_3_n44), .A(npu_inst_pe_1_2_3_n65), .ZN(
        npu_inst_pe_1_2_3_n88) );
  NAND2_X1 npu_inst_pe_1_2_3_U67 ( .A1(npu_inst_pe_1_2_3_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_2_3_n40), .ZN(npu_inst_pe_1_2_3_n64) );
  OAI21_X1 npu_inst_pe_1_2_3_U66 ( .B1(npu_inst_pe_1_2_3_n63), .B2(
        npu_inst_pe_1_2_3_n40), .A(npu_inst_pe_1_2_3_n64), .ZN(
        npu_inst_pe_1_2_3_n87) );
  NAND2_X1 npu_inst_pe_1_2_3_U65 ( .A1(npu_inst_pe_1_2_3_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_2_3_n40), .ZN(npu_inst_pe_1_2_3_n62) );
  OAI21_X1 npu_inst_pe_1_2_3_U64 ( .B1(npu_inst_pe_1_2_3_n61), .B2(
        npu_inst_pe_1_2_3_n40), .A(npu_inst_pe_1_2_3_n62), .ZN(
        npu_inst_pe_1_2_3_n86) );
  AND2_X1 npu_inst_pe_1_2_3_U63 ( .A1(npu_inst_pe_1_2_3_N93), .A2(npu_inst_n58), .ZN(npu_inst_int_data_y_2__3__0_) );
  AND2_X1 npu_inst_pe_1_2_3_U62 ( .A1(npu_inst_n58), .A2(npu_inst_pe_1_2_3_N94), .ZN(npu_inst_int_data_y_2__3__1_) );
  NOR3_X1 npu_inst_pe_1_2_3_U61 ( .A1(npu_inst_pe_1_2_3_n26), .A2(npu_inst_n58), .A3(npu_inst_int_ckg[44]), .ZN(npu_inst_pe_1_2_3_n85) );
  OR2_X1 npu_inst_pe_1_2_3_U60 ( .A1(npu_inst_pe_1_2_3_n85), .A2(
        npu_inst_pe_1_2_3_n2), .ZN(npu_inst_pe_1_2_3_N84) );
  AND2_X1 npu_inst_pe_1_2_3_U59 ( .A1(npu_inst_pe_1_2_3_int_q_acc_0_), .A2(
        npu_inst_pe_1_2_3_n1), .ZN(npu_inst_int_data_res_2__3__0_) );
  AND2_X1 npu_inst_pe_1_2_3_U58 ( .A1(npu_inst_pe_1_2_3_n2), .A2(
        npu_inst_pe_1_2_3_int_q_acc_7_), .ZN(npu_inst_int_data_res_2__3__7_)
         );
  AND2_X1 npu_inst_pe_1_2_3_U57 ( .A1(npu_inst_pe_1_2_3_int_q_acc_1_), .A2(
        npu_inst_pe_1_2_3_n1), .ZN(npu_inst_int_data_res_2__3__1_) );
  AND2_X1 npu_inst_pe_1_2_3_U56 ( .A1(npu_inst_pe_1_2_3_int_q_acc_2_), .A2(
        npu_inst_pe_1_2_3_n1), .ZN(npu_inst_int_data_res_2__3__2_) );
  AND2_X1 npu_inst_pe_1_2_3_U55 ( .A1(npu_inst_pe_1_2_3_int_q_acc_3_), .A2(
        npu_inst_pe_1_2_3_n2), .ZN(npu_inst_int_data_res_2__3__3_) );
  AND2_X1 npu_inst_pe_1_2_3_U54 ( .A1(npu_inst_pe_1_2_3_int_q_acc_4_), .A2(
        npu_inst_pe_1_2_3_n2), .ZN(npu_inst_int_data_res_2__3__4_) );
  AND2_X1 npu_inst_pe_1_2_3_U53 ( .A1(npu_inst_pe_1_2_3_int_q_acc_5_), .A2(
        npu_inst_pe_1_2_3_n2), .ZN(npu_inst_int_data_res_2__3__5_) );
  AND2_X1 npu_inst_pe_1_2_3_U52 ( .A1(npu_inst_pe_1_2_3_int_q_acc_6_), .A2(
        npu_inst_pe_1_2_3_n2), .ZN(npu_inst_int_data_res_2__3__6_) );
  AOI222_X1 npu_inst_pe_1_2_3_U51 ( .A1(npu_inst_int_data_res_3__3__0_), .A2(
        npu_inst_pe_1_2_3_n1), .B1(npu_inst_pe_1_2_3_N73), .B2(
        npu_inst_pe_1_2_3_n76), .C1(npu_inst_pe_1_2_3_N65), .C2(
        npu_inst_pe_1_2_3_n77), .ZN(npu_inst_pe_1_2_3_n84) );
  INV_X1 npu_inst_pe_1_2_3_U50 ( .A(npu_inst_pe_1_2_3_n84), .ZN(
        npu_inst_pe_1_2_3_n101) );
  AOI222_X1 npu_inst_pe_1_2_3_U49 ( .A1(npu_inst_int_data_res_3__3__7_), .A2(
        npu_inst_pe_1_2_3_n1), .B1(npu_inst_pe_1_2_3_N80), .B2(
        npu_inst_pe_1_2_3_n76), .C1(npu_inst_pe_1_2_3_N72), .C2(
        npu_inst_pe_1_2_3_n77), .ZN(npu_inst_pe_1_2_3_n75) );
  INV_X1 npu_inst_pe_1_2_3_U48 ( .A(npu_inst_pe_1_2_3_n75), .ZN(
        npu_inst_pe_1_2_3_n33) );
  AOI222_X1 npu_inst_pe_1_2_3_U47 ( .A1(npu_inst_int_data_res_3__3__1_), .A2(
        npu_inst_pe_1_2_3_n1), .B1(npu_inst_pe_1_2_3_N74), .B2(
        npu_inst_pe_1_2_3_n76), .C1(npu_inst_pe_1_2_3_N66), .C2(
        npu_inst_pe_1_2_3_n77), .ZN(npu_inst_pe_1_2_3_n83) );
  INV_X1 npu_inst_pe_1_2_3_U46 ( .A(npu_inst_pe_1_2_3_n83), .ZN(
        npu_inst_pe_1_2_3_n100) );
  AOI222_X1 npu_inst_pe_1_2_3_U45 ( .A1(npu_inst_int_data_res_3__3__2_), .A2(
        npu_inst_pe_1_2_3_n1), .B1(npu_inst_pe_1_2_3_N75), .B2(
        npu_inst_pe_1_2_3_n76), .C1(npu_inst_pe_1_2_3_N67), .C2(
        npu_inst_pe_1_2_3_n77), .ZN(npu_inst_pe_1_2_3_n82) );
  INV_X1 npu_inst_pe_1_2_3_U44 ( .A(npu_inst_pe_1_2_3_n82), .ZN(
        npu_inst_pe_1_2_3_n99) );
  AOI222_X1 npu_inst_pe_1_2_3_U43 ( .A1(npu_inst_int_data_res_3__3__3_), .A2(
        npu_inst_pe_1_2_3_n1), .B1(npu_inst_pe_1_2_3_N76), .B2(
        npu_inst_pe_1_2_3_n76), .C1(npu_inst_pe_1_2_3_N68), .C2(
        npu_inst_pe_1_2_3_n77), .ZN(npu_inst_pe_1_2_3_n81) );
  INV_X1 npu_inst_pe_1_2_3_U42 ( .A(npu_inst_pe_1_2_3_n81), .ZN(
        npu_inst_pe_1_2_3_n98) );
  AOI222_X1 npu_inst_pe_1_2_3_U41 ( .A1(npu_inst_int_data_res_3__3__4_), .A2(
        npu_inst_pe_1_2_3_n1), .B1(npu_inst_pe_1_2_3_N77), .B2(
        npu_inst_pe_1_2_3_n76), .C1(npu_inst_pe_1_2_3_N69), .C2(
        npu_inst_pe_1_2_3_n77), .ZN(npu_inst_pe_1_2_3_n80) );
  INV_X1 npu_inst_pe_1_2_3_U40 ( .A(npu_inst_pe_1_2_3_n80), .ZN(
        npu_inst_pe_1_2_3_n36) );
  AOI222_X1 npu_inst_pe_1_2_3_U39 ( .A1(npu_inst_int_data_res_3__3__5_), .A2(
        npu_inst_pe_1_2_3_n1), .B1(npu_inst_pe_1_2_3_N78), .B2(
        npu_inst_pe_1_2_3_n76), .C1(npu_inst_pe_1_2_3_N70), .C2(
        npu_inst_pe_1_2_3_n77), .ZN(npu_inst_pe_1_2_3_n79) );
  INV_X1 npu_inst_pe_1_2_3_U38 ( .A(npu_inst_pe_1_2_3_n79), .ZN(
        npu_inst_pe_1_2_3_n35) );
  AOI222_X1 npu_inst_pe_1_2_3_U37 ( .A1(npu_inst_int_data_res_3__3__6_), .A2(
        npu_inst_pe_1_2_3_n1), .B1(npu_inst_pe_1_2_3_N79), .B2(
        npu_inst_pe_1_2_3_n76), .C1(npu_inst_pe_1_2_3_N71), .C2(
        npu_inst_pe_1_2_3_n77), .ZN(npu_inst_pe_1_2_3_n78) );
  INV_X1 npu_inst_pe_1_2_3_U36 ( .A(npu_inst_pe_1_2_3_n78), .ZN(
        npu_inst_pe_1_2_3_n34) );
  INV_X1 npu_inst_pe_1_2_3_U35 ( .A(npu_inst_pe_1_2_3_int_data_1_), .ZN(
        npu_inst_pe_1_2_3_n14) );
  AND2_X1 npu_inst_pe_1_2_3_U34 ( .A1(npu_inst_int_data_x_2__3__1_), .A2(
        npu_inst_pe_1_2_3_int_q_weight_1_), .ZN(npu_inst_pe_1_2_3_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_2_3_U33 ( .A1(npu_inst_int_data_x_2__3__0_), .A2(
        npu_inst_pe_1_2_3_int_q_weight_1_), .ZN(npu_inst_pe_1_2_3_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_2_3_U32 ( .A1(npu_inst_n58), .A2(
        npu_inst_int_data_y_3__3__1_), .B1(npu_inst_pe_1_2_3_n3), .B2(
        npu_inst_int_data_x_2__4__1_), .ZN(npu_inst_pe_1_2_3_n63) );
  AOI22_X1 npu_inst_pe_1_2_3_U31 ( .A1(npu_inst_n58), .A2(
        npu_inst_int_data_y_3__3__0_), .B1(npu_inst_pe_1_2_3_n3), .B2(
        npu_inst_int_data_x_2__4__0_), .ZN(npu_inst_pe_1_2_3_n61) );
  INV_X1 npu_inst_pe_1_2_3_U30 ( .A(npu_inst_pe_1_2_3_int_data_0_), .ZN(
        npu_inst_pe_1_2_3_n13) );
  INV_X1 npu_inst_pe_1_2_3_U29 ( .A(npu_inst_n70), .ZN(npu_inst_pe_1_2_3_n5)
         );
  OR3_X1 npu_inst_pe_1_2_3_U28 ( .A1(npu_inst_pe_1_2_3_n6), .A2(
        npu_inst_pe_1_2_3_n8), .A3(npu_inst_pe_1_2_3_n5), .ZN(
        npu_inst_pe_1_2_3_n56) );
  OR3_X1 npu_inst_pe_1_2_3_U27 ( .A1(npu_inst_pe_1_2_3_n5), .A2(
        npu_inst_pe_1_2_3_n8), .A3(npu_inst_pe_1_2_3_n7), .ZN(
        npu_inst_pe_1_2_3_n48) );
  INV_X1 npu_inst_pe_1_2_3_U26 ( .A(npu_inst_pe_1_2_3_n5), .ZN(
        npu_inst_pe_1_2_3_n4) );
  OR3_X1 npu_inst_pe_1_2_3_U25 ( .A1(npu_inst_pe_1_2_3_n4), .A2(
        npu_inst_pe_1_2_3_n8), .A3(npu_inst_pe_1_2_3_n7), .ZN(
        npu_inst_pe_1_2_3_n52) );
  OR3_X1 npu_inst_pe_1_2_3_U24 ( .A1(npu_inst_pe_1_2_3_n6), .A2(
        npu_inst_pe_1_2_3_n8), .A3(npu_inst_pe_1_2_3_n4), .ZN(
        npu_inst_pe_1_2_3_n60) );
  NOR2_X1 npu_inst_pe_1_2_3_U23 ( .A1(npu_inst_pe_1_2_3_n60), .A2(
        npu_inst_pe_1_2_3_n3), .ZN(npu_inst_pe_1_2_3_n58) );
  NOR2_X1 npu_inst_pe_1_2_3_U22 ( .A1(npu_inst_pe_1_2_3_n56), .A2(
        npu_inst_pe_1_2_3_n3), .ZN(npu_inst_pe_1_2_3_n54) );
  NOR2_X1 npu_inst_pe_1_2_3_U21 ( .A1(npu_inst_pe_1_2_3_n52), .A2(
        npu_inst_pe_1_2_3_n3), .ZN(npu_inst_pe_1_2_3_n50) );
  NOR2_X1 npu_inst_pe_1_2_3_U20 ( .A1(npu_inst_pe_1_2_3_n48), .A2(
        npu_inst_pe_1_2_3_n3), .ZN(npu_inst_pe_1_2_3_n46) );
  NOR2_X1 npu_inst_pe_1_2_3_U19 ( .A1(npu_inst_pe_1_2_3_n40), .A2(
        npu_inst_pe_1_2_3_n3), .ZN(npu_inst_pe_1_2_3_n38) );
  NOR2_X1 npu_inst_pe_1_2_3_U18 ( .A1(npu_inst_pe_1_2_3_n44), .A2(
        npu_inst_pe_1_2_3_n3), .ZN(npu_inst_pe_1_2_3_n42) );
  BUF_X1 npu_inst_pe_1_2_3_U17 ( .A(npu_inst_n103), .Z(npu_inst_pe_1_2_3_n8)
         );
  INV_X1 npu_inst_pe_1_2_3_U16 ( .A(npu_inst_n125), .ZN(npu_inst_pe_1_2_3_n12)
         );
  INV_X1 npu_inst_pe_1_2_3_U15 ( .A(npu_inst_pe_1_2_3_n38), .ZN(
        npu_inst_pe_1_2_3_n114) );
  INV_X1 npu_inst_pe_1_2_3_U14 ( .A(npu_inst_pe_1_2_3_n58), .ZN(
        npu_inst_pe_1_2_3_n119) );
  INV_X1 npu_inst_pe_1_2_3_U13 ( .A(npu_inst_pe_1_2_3_n54), .ZN(
        npu_inst_pe_1_2_3_n118) );
  INV_X1 npu_inst_pe_1_2_3_U12 ( .A(npu_inst_pe_1_2_3_n50), .ZN(
        npu_inst_pe_1_2_3_n117) );
  INV_X1 npu_inst_pe_1_2_3_U11 ( .A(npu_inst_pe_1_2_3_n46), .ZN(
        npu_inst_pe_1_2_3_n116) );
  INV_X1 npu_inst_pe_1_2_3_U10 ( .A(npu_inst_pe_1_2_3_n42), .ZN(
        npu_inst_pe_1_2_3_n115) );
  BUF_X1 npu_inst_pe_1_2_3_U9 ( .A(npu_inst_n29), .Z(npu_inst_pe_1_2_3_n2) );
  BUF_X1 npu_inst_pe_1_2_3_U8 ( .A(npu_inst_n29), .Z(npu_inst_pe_1_2_3_n1) );
  BUF_X1 npu_inst_pe_1_2_3_U7 ( .A(npu_inst_pe_1_2_3_n12), .Z(
        npu_inst_pe_1_2_3_n11) );
  BUF_X1 npu_inst_pe_1_2_3_U6 ( .A(npu_inst_pe_1_2_3_n12), .Z(
        npu_inst_pe_1_2_3_n10) );
  BUF_X1 npu_inst_pe_1_2_3_U5 ( .A(npu_inst_pe_1_2_3_n12), .Z(
        npu_inst_pe_1_2_3_n9) );
  NOR2_X1 npu_inst_pe_1_2_3_U4 ( .A1(npu_inst_pe_1_2_3_int_q_weight_0_), .A2(
        npu_inst_pe_1_2_3_n1), .ZN(npu_inst_pe_1_2_3_n76) );
  NOR2_X1 npu_inst_pe_1_2_3_U3 ( .A1(npu_inst_pe_1_2_3_n27), .A2(
        npu_inst_pe_1_2_3_n1), .ZN(npu_inst_pe_1_2_3_n77) );
  FA_X1 npu_inst_pe_1_2_3_sub_67_U2_1 ( .A(npu_inst_pe_1_2_3_int_q_acc_1_), 
        .B(npu_inst_pe_1_2_3_n14), .CI(npu_inst_pe_1_2_3_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_2_3_sub_67_carry_2_), .S(npu_inst_pe_1_2_3_N66) );
  FA_X1 npu_inst_pe_1_2_3_add_69_U1_1 ( .A(npu_inst_pe_1_2_3_int_q_acc_1_), 
        .B(npu_inst_pe_1_2_3_int_data_1_), .CI(
        npu_inst_pe_1_2_3_add_69_carry_1_), .CO(
        npu_inst_pe_1_2_3_add_69_carry_2_), .S(npu_inst_pe_1_2_3_N74) );
  NAND3_X1 npu_inst_pe_1_2_3_U109 ( .A1(npu_inst_pe_1_2_3_n5), .A2(
        npu_inst_pe_1_2_3_n7), .A3(npu_inst_pe_1_2_3_n8), .ZN(
        npu_inst_pe_1_2_3_n44) );
  NAND3_X1 npu_inst_pe_1_2_3_U108 ( .A1(npu_inst_pe_1_2_3_n4), .A2(
        npu_inst_pe_1_2_3_n7), .A3(npu_inst_pe_1_2_3_n8), .ZN(
        npu_inst_pe_1_2_3_n40) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_2_3_n34), .CK(
        npu_inst_pe_1_2_3_net4125), .RN(npu_inst_pe_1_2_3_n9), .Q(
        npu_inst_pe_1_2_3_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_2_3_n35), .CK(
        npu_inst_pe_1_2_3_net4125), .RN(npu_inst_pe_1_2_3_n9), .Q(
        npu_inst_pe_1_2_3_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_2_3_n36), .CK(
        npu_inst_pe_1_2_3_net4125), .RN(npu_inst_pe_1_2_3_n9), .Q(
        npu_inst_pe_1_2_3_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_2_3_n98), .CK(
        npu_inst_pe_1_2_3_net4125), .RN(npu_inst_pe_1_2_3_n9), .Q(
        npu_inst_pe_1_2_3_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_2_3_n99), .CK(
        npu_inst_pe_1_2_3_net4125), .RN(npu_inst_pe_1_2_3_n9), .Q(
        npu_inst_pe_1_2_3_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_2_3_n100), 
        .CK(npu_inst_pe_1_2_3_net4125), .RN(npu_inst_pe_1_2_3_n9), .Q(
        npu_inst_pe_1_2_3_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_2_3_n33), .CK(
        npu_inst_pe_1_2_3_net4125), .RN(npu_inst_pe_1_2_3_n9), .Q(
        npu_inst_pe_1_2_3_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_2_3_n101), 
        .CK(npu_inst_pe_1_2_3_net4125), .RN(npu_inst_pe_1_2_3_n9), .Q(
        npu_inst_pe_1_2_3_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_weight_reg_0_ ( .D(npu_inst_n111), .CK(
        npu_inst_pe_1_2_3_net4131), .RN(npu_inst_pe_1_2_3_n9), .Q(
        npu_inst_pe_1_2_3_int_q_weight_0_), .QN(npu_inst_pe_1_2_3_n27) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_weight_reg_1_ ( .D(npu_inst_n117), .CK(
        npu_inst_pe_1_2_3_net4131), .RN(npu_inst_pe_1_2_3_n9), .Q(
        npu_inst_pe_1_2_3_int_q_weight_1_), .QN(npu_inst_pe_1_2_3_n26) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_2_3_n113), 
        .CK(npu_inst_pe_1_2_3_net4131), .RN(npu_inst_pe_1_2_3_n9), .Q(
        npu_inst_pe_1_2_3_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_2_3_n107), 
        .CK(npu_inst_pe_1_2_3_net4131), .RN(npu_inst_pe_1_2_3_n9), .Q(
        npu_inst_pe_1_2_3_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_2_3_n112), 
        .CK(npu_inst_pe_1_2_3_net4131), .RN(npu_inst_pe_1_2_3_n10), .Q(
        npu_inst_pe_1_2_3_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_2_3_n106), 
        .CK(npu_inst_pe_1_2_3_net4131), .RN(npu_inst_pe_1_2_3_n10), .Q(
        npu_inst_pe_1_2_3_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_2_3_n111), 
        .CK(npu_inst_pe_1_2_3_net4131), .RN(npu_inst_pe_1_2_3_n10), .Q(
        npu_inst_pe_1_2_3_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_2_3_n105), 
        .CK(npu_inst_pe_1_2_3_net4131), .RN(npu_inst_pe_1_2_3_n10), .Q(
        npu_inst_pe_1_2_3_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_2_3_n110), 
        .CK(npu_inst_pe_1_2_3_net4131), .RN(npu_inst_pe_1_2_3_n10), .Q(
        npu_inst_pe_1_2_3_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_2_3_n104), 
        .CK(npu_inst_pe_1_2_3_net4131), .RN(npu_inst_pe_1_2_3_n10), .Q(
        npu_inst_pe_1_2_3_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_2_3_n109), 
        .CK(npu_inst_pe_1_2_3_net4131), .RN(npu_inst_pe_1_2_3_n10), .Q(
        npu_inst_pe_1_2_3_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_2_3_n103), 
        .CK(npu_inst_pe_1_2_3_net4131), .RN(npu_inst_pe_1_2_3_n10), .Q(
        npu_inst_pe_1_2_3_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_2_3_n108), 
        .CK(npu_inst_pe_1_2_3_net4131), .RN(npu_inst_pe_1_2_3_n10), .Q(
        npu_inst_pe_1_2_3_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_2_3_n102), 
        .CK(npu_inst_pe_1_2_3_net4131), .RN(npu_inst_pe_1_2_3_n10), .Q(
        npu_inst_pe_1_2_3_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_2_3_n86), 
        .CK(npu_inst_pe_1_2_3_net4131), .RN(npu_inst_pe_1_2_3_n10), .Q(
        npu_inst_pe_1_2_3_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_2_3_n87), 
        .CK(npu_inst_pe_1_2_3_net4131), .RN(npu_inst_pe_1_2_3_n10), .Q(
        npu_inst_pe_1_2_3_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_2_3_n88), 
        .CK(npu_inst_pe_1_2_3_net4131), .RN(npu_inst_pe_1_2_3_n11), .Q(
        npu_inst_pe_1_2_3_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_2_3_n89), 
        .CK(npu_inst_pe_1_2_3_net4131), .RN(npu_inst_pe_1_2_3_n11), .Q(
        npu_inst_pe_1_2_3_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_2_3_n90), 
        .CK(npu_inst_pe_1_2_3_net4131), .RN(npu_inst_pe_1_2_3_n11), .Q(
        npu_inst_pe_1_2_3_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_2_3_n91), 
        .CK(npu_inst_pe_1_2_3_net4131), .RN(npu_inst_pe_1_2_3_n11), .Q(
        npu_inst_pe_1_2_3_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_2_3_n92), 
        .CK(npu_inst_pe_1_2_3_net4131), .RN(npu_inst_pe_1_2_3_n11), .Q(
        npu_inst_pe_1_2_3_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_2_3_n93), 
        .CK(npu_inst_pe_1_2_3_net4131), .RN(npu_inst_pe_1_2_3_n11), .Q(
        npu_inst_pe_1_2_3_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_2_3_n94), 
        .CK(npu_inst_pe_1_2_3_net4131), .RN(npu_inst_pe_1_2_3_n11), .Q(
        npu_inst_pe_1_2_3_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_2_3_n95), 
        .CK(npu_inst_pe_1_2_3_net4131), .RN(npu_inst_pe_1_2_3_n11), .Q(
        npu_inst_pe_1_2_3_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_2_3_n96), 
        .CK(npu_inst_pe_1_2_3_net4131), .RN(npu_inst_pe_1_2_3_n11), .Q(
        npu_inst_pe_1_2_3_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_2_3_n97), 
        .CK(npu_inst_pe_1_2_3_net4131), .RN(npu_inst_pe_1_2_3_n11), .Q(
        npu_inst_pe_1_2_3_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_2_3_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_2_3_N84), .SE(1'b0), .GCK(npu_inst_pe_1_2_3_net4125) );
  CLKGATETST_X1 npu_inst_pe_1_2_3_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n65), .SE(1'b0), .GCK(npu_inst_pe_1_2_3_net4131) );
  MUX2_X1 npu_inst_pe_1_2_4_U162 ( .A(npu_inst_pe_1_2_4_n32), .B(
        npu_inst_pe_1_2_4_n29), .S(npu_inst_pe_1_2_4_n8), .Z(
        npu_inst_pe_1_2_4_N93) );
  MUX2_X1 npu_inst_pe_1_2_4_U161 ( .A(npu_inst_pe_1_2_4_n31), .B(
        npu_inst_pe_1_2_4_n30), .S(npu_inst_pe_1_2_4_n6), .Z(
        npu_inst_pe_1_2_4_n32) );
  MUX2_X1 npu_inst_pe_1_2_4_U160 ( .A(npu_inst_pe_1_2_4_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_2_4_int_q_reg_v_1__0_), .S(npu_inst_pe_1_2_4_n4), .Z(
        npu_inst_pe_1_2_4_n31) );
  MUX2_X1 npu_inst_pe_1_2_4_U159 ( .A(npu_inst_pe_1_2_4_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_2_4_int_q_reg_v_3__0_), .S(npu_inst_pe_1_2_4_n4), .Z(
        npu_inst_pe_1_2_4_n30) );
  MUX2_X1 npu_inst_pe_1_2_4_U158 ( .A(npu_inst_pe_1_2_4_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_2_4_int_q_reg_v_5__0_), .S(npu_inst_pe_1_2_4_n4), .Z(
        npu_inst_pe_1_2_4_n29) );
  MUX2_X1 npu_inst_pe_1_2_4_U157 ( .A(npu_inst_pe_1_2_4_n28), .B(
        npu_inst_pe_1_2_4_n23), .S(npu_inst_pe_1_2_4_n8), .Z(
        npu_inst_pe_1_2_4_N94) );
  MUX2_X1 npu_inst_pe_1_2_4_U156 ( .A(npu_inst_pe_1_2_4_n25), .B(
        npu_inst_pe_1_2_4_n24), .S(npu_inst_pe_1_2_4_n6), .Z(
        npu_inst_pe_1_2_4_n28) );
  MUX2_X1 npu_inst_pe_1_2_4_U155 ( .A(npu_inst_pe_1_2_4_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_2_4_int_q_reg_v_1__1_), .S(npu_inst_pe_1_2_4_n4), .Z(
        npu_inst_pe_1_2_4_n25) );
  MUX2_X1 npu_inst_pe_1_2_4_U154 ( .A(npu_inst_pe_1_2_4_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_2_4_int_q_reg_v_3__1_), .S(npu_inst_pe_1_2_4_n4), .Z(
        npu_inst_pe_1_2_4_n24) );
  MUX2_X1 npu_inst_pe_1_2_4_U153 ( .A(npu_inst_pe_1_2_4_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_2_4_int_q_reg_v_5__1_), .S(npu_inst_pe_1_2_4_n4), .Z(
        npu_inst_pe_1_2_4_n23) );
  MUX2_X1 npu_inst_pe_1_2_4_U152 ( .A(npu_inst_pe_1_2_4_n22), .B(
        npu_inst_pe_1_2_4_n19), .S(npu_inst_pe_1_2_4_n8), .Z(
        npu_inst_int_data_x_2__4__1_) );
  MUX2_X1 npu_inst_pe_1_2_4_U151 ( .A(npu_inst_pe_1_2_4_n21), .B(
        npu_inst_pe_1_2_4_n20), .S(npu_inst_pe_1_2_4_n6), .Z(
        npu_inst_pe_1_2_4_n22) );
  MUX2_X1 npu_inst_pe_1_2_4_U150 ( .A(npu_inst_pe_1_2_4_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_2_4_int_q_reg_h_1__1_), .S(npu_inst_pe_1_2_4_n4), .Z(
        npu_inst_pe_1_2_4_n21) );
  MUX2_X1 npu_inst_pe_1_2_4_U149 ( .A(npu_inst_pe_1_2_4_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_2_4_int_q_reg_h_3__1_), .S(npu_inst_pe_1_2_4_n4), .Z(
        npu_inst_pe_1_2_4_n20) );
  MUX2_X1 npu_inst_pe_1_2_4_U148 ( .A(npu_inst_pe_1_2_4_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_2_4_int_q_reg_h_5__1_), .S(npu_inst_pe_1_2_4_n4), .Z(
        npu_inst_pe_1_2_4_n19) );
  MUX2_X1 npu_inst_pe_1_2_4_U147 ( .A(npu_inst_pe_1_2_4_n18), .B(
        npu_inst_pe_1_2_4_n15), .S(npu_inst_pe_1_2_4_n8), .Z(
        npu_inst_int_data_x_2__4__0_) );
  MUX2_X1 npu_inst_pe_1_2_4_U146 ( .A(npu_inst_pe_1_2_4_n17), .B(
        npu_inst_pe_1_2_4_n16), .S(npu_inst_pe_1_2_4_n6), .Z(
        npu_inst_pe_1_2_4_n18) );
  MUX2_X1 npu_inst_pe_1_2_4_U145 ( .A(npu_inst_pe_1_2_4_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_2_4_int_q_reg_h_1__0_), .S(npu_inst_pe_1_2_4_n4), .Z(
        npu_inst_pe_1_2_4_n17) );
  MUX2_X1 npu_inst_pe_1_2_4_U144 ( .A(npu_inst_pe_1_2_4_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_2_4_int_q_reg_h_3__0_), .S(npu_inst_pe_1_2_4_n4), .Z(
        npu_inst_pe_1_2_4_n16) );
  MUX2_X1 npu_inst_pe_1_2_4_U143 ( .A(npu_inst_pe_1_2_4_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_2_4_int_q_reg_h_5__0_), .S(npu_inst_pe_1_2_4_n4), .Z(
        npu_inst_pe_1_2_4_n15) );
  XOR2_X1 npu_inst_pe_1_2_4_U142 ( .A(npu_inst_pe_1_2_4_int_data_0_), .B(
        npu_inst_pe_1_2_4_int_q_acc_0_), .Z(npu_inst_pe_1_2_4_N73) );
  AND2_X1 npu_inst_pe_1_2_4_U141 ( .A1(npu_inst_pe_1_2_4_int_q_acc_0_), .A2(
        npu_inst_pe_1_2_4_int_data_0_), .ZN(npu_inst_pe_1_2_4_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_2_4_U140 ( .A(npu_inst_pe_1_2_4_int_q_acc_0_), .B(
        npu_inst_pe_1_2_4_n13), .ZN(npu_inst_pe_1_2_4_N65) );
  OR2_X1 npu_inst_pe_1_2_4_U139 ( .A1(npu_inst_pe_1_2_4_n13), .A2(
        npu_inst_pe_1_2_4_int_q_acc_0_), .ZN(npu_inst_pe_1_2_4_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_2_4_U138 ( .A(npu_inst_pe_1_2_4_int_q_acc_2_), .B(
        npu_inst_pe_1_2_4_add_69_carry_2_), .Z(npu_inst_pe_1_2_4_N75) );
  AND2_X1 npu_inst_pe_1_2_4_U137 ( .A1(npu_inst_pe_1_2_4_add_69_carry_2_), 
        .A2(npu_inst_pe_1_2_4_int_q_acc_2_), .ZN(
        npu_inst_pe_1_2_4_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_2_4_U136 ( .A(npu_inst_pe_1_2_4_int_q_acc_3_), .B(
        npu_inst_pe_1_2_4_add_69_carry_3_), .Z(npu_inst_pe_1_2_4_N76) );
  AND2_X1 npu_inst_pe_1_2_4_U135 ( .A1(npu_inst_pe_1_2_4_add_69_carry_3_), 
        .A2(npu_inst_pe_1_2_4_int_q_acc_3_), .ZN(
        npu_inst_pe_1_2_4_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_2_4_U134 ( .A(npu_inst_pe_1_2_4_int_q_acc_4_), .B(
        npu_inst_pe_1_2_4_add_69_carry_4_), .Z(npu_inst_pe_1_2_4_N77) );
  AND2_X1 npu_inst_pe_1_2_4_U133 ( .A1(npu_inst_pe_1_2_4_add_69_carry_4_), 
        .A2(npu_inst_pe_1_2_4_int_q_acc_4_), .ZN(
        npu_inst_pe_1_2_4_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_2_4_U132 ( .A(npu_inst_pe_1_2_4_int_q_acc_5_), .B(
        npu_inst_pe_1_2_4_add_69_carry_5_), .Z(npu_inst_pe_1_2_4_N78) );
  AND2_X1 npu_inst_pe_1_2_4_U131 ( .A1(npu_inst_pe_1_2_4_add_69_carry_5_), 
        .A2(npu_inst_pe_1_2_4_int_q_acc_5_), .ZN(
        npu_inst_pe_1_2_4_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_2_4_U130 ( .A(npu_inst_pe_1_2_4_int_q_acc_6_), .B(
        npu_inst_pe_1_2_4_add_69_carry_6_), .Z(npu_inst_pe_1_2_4_N79) );
  AND2_X1 npu_inst_pe_1_2_4_U129 ( .A1(npu_inst_pe_1_2_4_add_69_carry_6_), 
        .A2(npu_inst_pe_1_2_4_int_q_acc_6_), .ZN(
        npu_inst_pe_1_2_4_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_2_4_U128 ( .A(npu_inst_pe_1_2_4_int_q_acc_7_), .B(
        npu_inst_pe_1_2_4_add_69_carry_7_), .Z(npu_inst_pe_1_2_4_N80) );
  XNOR2_X1 npu_inst_pe_1_2_4_U127 ( .A(npu_inst_pe_1_2_4_sub_67_carry_2_), .B(
        npu_inst_pe_1_2_4_int_q_acc_2_), .ZN(npu_inst_pe_1_2_4_N67) );
  OR2_X1 npu_inst_pe_1_2_4_U126 ( .A1(npu_inst_pe_1_2_4_int_q_acc_2_), .A2(
        npu_inst_pe_1_2_4_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_2_4_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_2_4_U125 ( .A(npu_inst_pe_1_2_4_sub_67_carry_3_), .B(
        npu_inst_pe_1_2_4_int_q_acc_3_), .ZN(npu_inst_pe_1_2_4_N68) );
  OR2_X1 npu_inst_pe_1_2_4_U124 ( .A1(npu_inst_pe_1_2_4_int_q_acc_3_), .A2(
        npu_inst_pe_1_2_4_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_2_4_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_2_4_U123 ( .A(npu_inst_pe_1_2_4_sub_67_carry_4_), .B(
        npu_inst_pe_1_2_4_int_q_acc_4_), .ZN(npu_inst_pe_1_2_4_N69) );
  OR2_X1 npu_inst_pe_1_2_4_U122 ( .A1(npu_inst_pe_1_2_4_int_q_acc_4_), .A2(
        npu_inst_pe_1_2_4_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_2_4_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_2_4_U121 ( .A(npu_inst_pe_1_2_4_sub_67_carry_5_), .B(
        npu_inst_pe_1_2_4_int_q_acc_5_), .ZN(npu_inst_pe_1_2_4_N70) );
  OR2_X1 npu_inst_pe_1_2_4_U120 ( .A1(npu_inst_pe_1_2_4_int_q_acc_5_), .A2(
        npu_inst_pe_1_2_4_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_2_4_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_2_4_U119 ( .A(npu_inst_pe_1_2_4_sub_67_carry_6_), .B(
        npu_inst_pe_1_2_4_int_q_acc_6_), .ZN(npu_inst_pe_1_2_4_N71) );
  OR2_X1 npu_inst_pe_1_2_4_U118 ( .A1(npu_inst_pe_1_2_4_int_q_acc_6_), .A2(
        npu_inst_pe_1_2_4_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_2_4_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_2_4_U117 ( .A(npu_inst_pe_1_2_4_int_q_acc_7_), .B(
        npu_inst_pe_1_2_4_sub_67_carry_7_), .ZN(npu_inst_pe_1_2_4_N72) );
  INV_X1 npu_inst_pe_1_2_4_U116 ( .A(npu_inst_n78), .ZN(npu_inst_pe_1_2_4_n7)
         );
  INV_X1 npu_inst_pe_1_2_4_U115 ( .A(npu_inst_pe_1_2_4_n7), .ZN(
        npu_inst_pe_1_2_4_n6) );
  INV_X1 npu_inst_pe_1_2_4_U114 ( .A(npu_inst_n58), .ZN(npu_inst_pe_1_2_4_n3)
         );
  AOI22_X1 npu_inst_pe_1_2_4_U113 ( .A1(npu_inst_int_data_y_3__4__0_), .A2(
        npu_inst_pe_1_2_4_n58), .B1(npu_inst_pe_1_2_4_n119), .B2(
        npu_inst_pe_1_2_4_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_2_4_n57) );
  INV_X1 npu_inst_pe_1_2_4_U112 ( .A(npu_inst_pe_1_2_4_n57), .ZN(
        npu_inst_pe_1_2_4_n108) );
  AOI22_X1 npu_inst_pe_1_2_4_U111 ( .A1(npu_inst_int_data_y_3__4__0_), .A2(
        npu_inst_pe_1_2_4_n54), .B1(npu_inst_pe_1_2_4_n118), .B2(
        npu_inst_pe_1_2_4_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_2_4_n53) );
  INV_X1 npu_inst_pe_1_2_4_U110 ( .A(npu_inst_pe_1_2_4_n53), .ZN(
        npu_inst_pe_1_2_4_n109) );
  AOI22_X1 npu_inst_pe_1_2_4_U107 ( .A1(npu_inst_int_data_y_3__4__0_), .A2(
        npu_inst_pe_1_2_4_n50), .B1(npu_inst_pe_1_2_4_n117), .B2(
        npu_inst_pe_1_2_4_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_2_4_n49) );
  INV_X1 npu_inst_pe_1_2_4_U106 ( .A(npu_inst_pe_1_2_4_n49), .ZN(
        npu_inst_pe_1_2_4_n110) );
  AOI22_X1 npu_inst_pe_1_2_4_U105 ( .A1(npu_inst_int_data_y_3__4__0_), .A2(
        npu_inst_pe_1_2_4_n46), .B1(npu_inst_pe_1_2_4_n116), .B2(
        npu_inst_pe_1_2_4_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_2_4_n45) );
  INV_X1 npu_inst_pe_1_2_4_U104 ( .A(npu_inst_pe_1_2_4_n45), .ZN(
        npu_inst_pe_1_2_4_n111) );
  AOI22_X1 npu_inst_pe_1_2_4_U103 ( .A1(npu_inst_int_data_y_3__4__0_), .A2(
        npu_inst_pe_1_2_4_n42), .B1(npu_inst_pe_1_2_4_n115), .B2(
        npu_inst_pe_1_2_4_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_2_4_n41) );
  INV_X1 npu_inst_pe_1_2_4_U102 ( .A(npu_inst_pe_1_2_4_n41), .ZN(
        npu_inst_pe_1_2_4_n112) );
  AOI22_X1 npu_inst_pe_1_2_4_U101 ( .A1(npu_inst_int_data_y_3__4__1_), .A2(
        npu_inst_pe_1_2_4_n58), .B1(npu_inst_pe_1_2_4_n119), .B2(
        npu_inst_pe_1_2_4_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_2_4_n59) );
  INV_X1 npu_inst_pe_1_2_4_U100 ( .A(npu_inst_pe_1_2_4_n59), .ZN(
        npu_inst_pe_1_2_4_n102) );
  AOI22_X1 npu_inst_pe_1_2_4_U99 ( .A1(npu_inst_int_data_y_3__4__1_), .A2(
        npu_inst_pe_1_2_4_n54), .B1(npu_inst_pe_1_2_4_n118), .B2(
        npu_inst_pe_1_2_4_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_2_4_n55) );
  INV_X1 npu_inst_pe_1_2_4_U98 ( .A(npu_inst_pe_1_2_4_n55), .ZN(
        npu_inst_pe_1_2_4_n103) );
  AOI22_X1 npu_inst_pe_1_2_4_U97 ( .A1(npu_inst_int_data_y_3__4__1_), .A2(
        npu_inst_pe_1_2_4_n50), .B1(npu_inst_pe_1_2_4_n117), .B2(
        npu_inst_pe_1_2_4_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_2_4_n51) );
  INV_X1 npu_inst_pe_1_2_4_U96 ( .A(npu_inst_pe_1_2_4_n51), .ZN(
        npu_inst_pe_1_2_4_n104) );
  AOI22_X1 npu_inst_pe_1_2_4_U95 ( .A1(npu_inst_int_data_y_3__4__1_), .A2(
        npu_inst_pe_1_2_4_n46), .B1(npu_inst_pe_1_2_4_n116), .B2(
        npu_inst_pe_1_2_4_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_2_4_n47) );
  INV_X1 npu_inst_pe_1_2_4_U94 ( .A(npu_inst_pe_1_2_4_n47), .ZN(
        npu_inst_pe_1_2_4_n105) );
  AOI22_X1 npu_inst_pe_1_2_4_U93 ( .A1(npu_inst_int_data_y_3__4__1_), .A2(
        npu_inst_pe_1_2_4_n42), .B1(npu_inst_pe_1_2_4_n115), .B2(
        npu_inst_pe_1_2_4_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_2_4_n43) );
  INV_X1 npu_inst_pe_1_2_4_U92 ( .A(npu_inst_pe_1_2_4_n43), .ZN(
        npu_inst_pe_1_2_4_n106) );
  AOI22_X1 npu_inst_pe_1_2_4_U91 ( .A1(npu_inst_pe_1_2_4_n38), .A2(
        npu_inst_int_data_y_3__4__1_), .B1(npu_inst_pe_1_2_4_n114), .B2(
        npu_inst_pe_1_2_4_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_2_4_n39) );
  INV_X1 npu_inst_pe_1_2_4_U90 ( .A(npu_inst_pe_1_2_4_n39), .ZN(
        npu_inst_pe_1_2_4_n107) );
  AOI22_X1 npu_inst_pe_1_2_4_U89 ( .A1(npu_inst_pe_1_2_4_n38), .A2(
        npu_inst_int_data_y_3__4__0_), .B1(npu_inst_pe_1_2_4_n114), .B2(
        npu_inst_pe_1_2_4_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_2_4_n37) );
  INV_X1 npu_inst_pe_1_2_4_U88 ( .A(npu_inst_pe_1_2_4_n37), .ZN(
        npu_inst_pe_1_2_4_n113) );
  NAND2_X1 npu_inst_pe_1_2_4_U87 ( .A1(npu_inst_pe_1_2_4_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_2_4_n60), .ZN(npu_inst_pe_1_2_4_n74) );
  OAI21_X1 npu_inst_pe_1_2_4_U86 ( .B1(npu_inst_pe_1_2_4_n63), .B2(
        npu_inst_pe_1_2_4_n60), .A(npu_inst_pe_1_2_4_n74), .ZN(
        npu_inst_pe_1_2_4_n97) );
  NAND2_X1 npu_inst_pe_1_2_4_U85 ( .A1(npu_inst_pe_1_2_4_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_2_4_n60), .ZN(npu_inst_pe_1_2_4_n73) );
  OAI21_X1 npu_inst_pe_1_2_4_U84 ( .B1(npu_inst_pe_1_2_4_n61), .B2(
        npu_inst_pe_1_2_4_n60), .A(npu_inst_pe_1_2_4_n73), .ZN(
        npu_inst_pe_1_2_4_n96) );
  NAND2_X1 npu_inst_pe_1_2_4_U83 ( .A1(npu_inst_pe_1_2_4_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_2_4_n56), .ZN(npu_inst_pe_1_2_4_n72) );
  OAI21_X1 npu_inst_pe_1_2_4_U82 ( .B1(npu_inst_pe_1_2_4_n63), .B2(
        npu_inst_pe_1_2_4_n56), .A(npu_inst_pe_1_2_4_n72), .ZN(
        npu_inst_pe_1_2_4_n95) );
  NAND2_X1 npu_inst_pe_1_2_4_U81 ( .A1(npu_inst_pe_1_2_4_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_2_4_n56), .ZN(npu_inst_pe_1_2_4_n71) );
  OAI21_X1 npu_inst_pe_1_2_4_U80 ( .B1(npu_inst_pe_1_2_4_n61), .B2(
        npu_inst_pe_1_2_4_n56), .A(npu_inst_pe_1_2_4_n71), .ZN(
        npu_inst_pe_1_2_4_n94) );
  NAND2_X1 npu_inst_pe_1_2_4_U79 ( .A1(npu_inst_pe_1_2_4_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_2_4_n52), .ZN(npu_inst_pe_1_2_4_n70) );
  OAI21_X1 npu_inst_pe_1_2_4_U78 ( .B1(npu_inst_pe_1_2_4_n63), .B2(
        npu_inst_pe_1_2_4_n52), .A(npu_inst_pe_1_2_4_n70), .ZN(
        npu_inst_pe_1_2_4_n93) );
  NAND2_X1 npu_inst_pe_1_2_4_U77 ( .A1(npu_inst_pe_1_2_4_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_2_4_n52), .ZN(npu_inst_pe_1_2_4_n69) );
  OAI21_X1 npu_inst_pe_1_2_4_U76 ( .B1(npu_inst_pe_1_2_4_n61), .B2(
        npu_inst_pe_1_2_4_n52), .A(npu_inst_pe_1_2_4_n69), .ZN(
        npu_inst_pe_1_2_4_n92) );
  NAND2_X1 npu_inst_pe_1_2_4_U75 ( .A1(npu_inst_pe_1_2_4_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_2_4_n48), .ZN(npu_inst_pe_1_2_4_n68) );
  OAI21_X1 npu_inst_pe_1_2_4_U74 ( .B1(npu_inst_pe_1_2_4_n63), .B2(
        npu_inst_pe_1_2_4_n48), .A(npu_inst_pe_1_2_4_n68), .ZN(
        npu_inst_pe_1_2_4_n91) );
  NAND2_X1 npu_inst_pe_1_2_4_U73 ( .A1(npu_inst_pe_1_2_4_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_2_4_n48), .ZN(npu_inst_pe_1_2_4_n67) );
  OAI21_X1 npu_inst_pe_1_2_4_U72 ( .B1(npu_inst_pe_1_2_4_n61), .B2(
        npu_inst_pe_1_2_4_n48), .A(npu_inst_pe_1_2_4_n67), .ZN(
        npu_inst_pe_1_2_4_n90) );
  NAND2_X1 npu_inst_pe_1_2_4_U71 ( .A1(npu_inst_pe_1_2_4_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_2_4_n44), .ZN(npu_inst_pe_1_2_4_n66) );
  OAI21_X1 npu_inst_pe_1_2_4_U70 ( .B1(npu_inst_pe_1_2_4_n63), .B2(
        npu_inst_pe_1_2_4_n44), .A(npu_inst_pe_1_2_4_n66), .ZN(
        npu_inst_pe_1_2_4_n89) );
  NAND2_X1 npu_inst_pe_1_2_4_U69 ( .A1(npu_inst_pe_1_2_4_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_2_4_n44), .ZN(npu_inst_pe_1_2_4_n65) );
  OAI21_X1 npu_inst_pe_1_2_4_U68 ( .B1(npu_inst_pe_1_2_4_n61), .B2(
        npu_inst_pe_1_2_4_n44), .A(npu_inst_pe_1_2_4_n65), .ZN(
        npu_inst_pe_1_2_4_n88) );
  NAND2_X1 npu_inst_pe_1_2_4_U67 ( .A1(npu_inst_pe_1_2_4_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_2_4_n40), .ZN(npu_inst_pe_1_2_4_n64) );
  OAI21_X1 npu_inst_pe_1_2_4_U66 ( .B1(npu_inst_pe_1_2_4_n63), .B2(
        npu_inst_pe_1_2_4_n40), .A(npu_inst_pe_1_2_4_n64), .ZN(
        npu_inst_pe_1_2_4_n87) );
  NAND2_X1 npu_inst_pe_1_2_4_U65 ( .A1(npu_inst_pe_1_2_4_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_2_4_n40), .ZN(npu_inst_pe_1_2_4_n62) );
  OAI21_X1 npu_inst_pe_1_2_4_U64 ( .B1(npu_inst_pe_1_2_4_n61), .B2(
        npu_inst_pe_1_2_4_n40), .A(npu_inst_pe_1_2_4_n62), .ZN(
        npu_inst_pe_1_2_4_n86) );
  AND2_X1 npu_inst_pe_1_2_4_U63 ( .A1(npu_inst_pe_1_2_4_N93), .A2(npu_inst_n58), .ZN(npu_inst_int_data_y_2__4__0_) );
  AND2_X1 npu_inst_pe_1_2_4_U62 ( .A1(npu_inst_n58), .A2(npu_inst_pe_1_2_4_N94), .ZN(npu_inst_int_data_y_2__4__1_) );
  NOR3_X1 npu_inst_pe_1_2_4_U61 ( .A1(npu_inst_pe_1_2_4_n26), .A2(npu_inst_n58), .A3(npu_inst_int_ckg[43]), .ZN(npu_inst_pe_1_2_4_n85) );
  OR2_X1 npu_inst_pe_1_2_4_U60 ( .A1(npu_inst_pe_1_2_4_n85), .A2(
        npu_inst_pe_1_2_4_n2), .ZN(npu_inst_pe_1_2_4_N84) );
  AND2_X1 npu_inst_pe_1_2_4_U59 ( .A1(npu_inst_pe_1_2_4_int_q_acc_0_), .A2(
        npu_inst_pe_1_2_4_n1), .ZN(npu_inst_int_data_res_2__4__0_) );
  AND2_X1 npu_inst_pe_1_2_4_U58 ( .A1(npu_inst_pe_1_2_4_n2), .A2(
        npu_inst_pe_1_2_4_int_q_acc_7_), .ZN(npu_inst_int_data_res_2__4__7_)
         );
  AND2_X1 npu_inst_pe_1_2_4_U57 ( .A1(npu_inst_pe_1_2_4_int_q_acc_1_), .A2(
        npu_inst_pe_1_2_4_n1), .ZN(npu_inst_int_data_res_2__4__1_) );
  AND2_X1 npu_inst_pe_1_2_4_U56 ( .A1(npu_inst_pe_1_2_4_int_q_acc_2_), .A2(
        npu_inst_pe_1_2_4_n1), .ZN(npu_inst_int_data_res_2__4__2_) );
  AND2_X1 npu_inst_pe_1_2_4_U55 ( .A1(npu_inst_pe_1_2_4_int_q_acc_3_), .A2(
        npu_inst_pe_1_2_4_n2), .ZN(npu_inst_int_data_res_2__4__3_) );
  AND2_X1 npu_inst_pe_1_2_4_U54 ( .A1(npu_inst_pe_1_2_4_int_q_acc_4_), .A2(
        npu_inst_pe_1_2_4_n2), .ZN(npu_inst_int_data_res_2__4__4_) );
  AND2_X1 npu_inst_pe_1_2_4_U53 ( .A1(npu_inst_pe_1_2_4_int_q_acc_5_), .A2(
        npu_inst_pe_1_2_4_n2), .ZN(npu_inst_int_data_res_2__4__5_) );
  AND2_X1 npu_inst_pe_1_2_4_U52 ( .A1(npu_inst_pe_1_2_4_int_q_acc_6_), .A2(
        npu_inst_pe_1_2_4_n2), .ZN(npu_inst_int_data_res_2__4__6_) );
  AOI222_X1 npu_inst_pe_1_2_4_U51 ( .A1(npu_inst_int_data_res_3__4__0_), .A2(
        npu_inst_pe_1_2_4_n1), .B1(npu_inst_pe_1_2_4_N73), .B2(
        npu_inst_pe_1_2_4_n76), .C1(npu_inst_pe_1_2_4_N65), .C2(
        npu_inst_pe_1_2_4_n77), .ZN(npu_inst_pe_1_2_4_n84) );
  INV_X1 npu_inst_pe_1_2_4_U50 ( .A(npu_inst_pe_1_2_4_n84), .ZN(
        npu_inst_pe_1_2_4_n101) );
  AOI222_X1 npu_inst_pe_1_2_4_U49 ( .A1(npu_inst_int_data_res_3__4__7_), .A2(
        npu_inst_pe_1_2_4_n1), .B1(npu_inst_pe_1_2_4_N80), .B2(
        npu_inst_pe_1_2_4_n76), .C1(npu_inst_pe_1_2_4_N72), .C2(
        npu_inst_pe_1_2_4_n77), .ZN(npu_inst_pe_1_2_4_n75) );
  INV_X1 npu_inst_pe_1_2_4_U48 ( .A(npu_inst_pe_1_2_4_n75), .ZN(
        npu_inst_pe_1_2_4_n33) );
  AOI222_X1 npu_inst_pe_1_2_4_U47 ( .A1(npu_inst_int_data_res_3__4__1_), .A2(
        npu_inst_pe_1_2_4_n1), .B1(npu_inst_pe_1_2_4_N74), .B2(
        npu_inst_pe_1_2_4_n76), .C1(npu_inst_pe_1_2_4_N66), .C2(
        npu_inst_pe_1_2_4_n77), .ZN(npu_inst_pe_1_2_4_n83) );
  INV_X1 npu_inst_pe_1_2_4_U46 ( .A(npu_inst_pe_1_2_4_n83), .ZN(
        npu_inst_pe_1_2_4_n100) );
  AOI222_X1 npu_inst_pe_1_2_4_U45 ( .A1(npu_inst_int_data_res_3__4__2_), .A2(
        npu_inst_pe_1_2_4_n1), .B1(npu_inst_pe_1_2_4_N75), .B2(
        npu_inst_pe_1_2_4_n76), .C1(npu_inst_pe_1_2_4_N67), .C2(
        npu_inst_pe_1_2_4_n77), .ZN(npu_inst_pe_1_2_4_n82) );
  INV_X1 npu_inst_pe_1_2_4_U44 ( .A(npu_inst_pe_1_2_4_n82), .ZN(
        npu_inst_pe_1_2_4_n99) );
  AOI222_X1 npu_inst_pe_1_2_4_U43 ( .A1(npu_inst_int_data_res_3__4__3_), .A2(
        npu_inst_pe_1_2_4_n1), .B1(npu_inst_pe_1_2_4_N76), .B2(
        npu_inst_pe_1_2_4_n76), .C1(npu_inst_pe_1_2_4_N68), .C2(
        npu_inst_pe_1_2_4_n77), .ZN(npu_inst_pe_1_2_4_n81) );
  INV_X1 npu_inst_pe_1_2_4_U42 ( .A(npu_inst_pe_1_2_4_n81), .ZN(
        npu_inst_pe_1_2_4_n98) );
  AOI222_X1 npu_inst_pe_1_2_4_U41 ( .A1(npu_inst_int_data_res_3__4__4_), .A2(
        npu_inst_pe_1_2_4_n1), .B1(npu_inst_pe_1_2_4_N77), .B2(
        npu_inst_pe_1_2_4_n76), .C1(npu_inst_pe_1_2_4_N69), .C2(
        npu_inst_pe_1_2_4_n77), .ZN(npu_inst_pe_1_2_4_n80) );
  INV_X1 npu_inst_pe_1_2_4_U40 ( .A(npu_inst_pe_1_2_4_n80), .ZN(
        npu_inst_pe_1_2_4_n36) );
  AOI222_X1 npu_inst_pe_1_2_4_U39 ( .A1(npu_inst_int_data_res_3__4__5_), .A2(
        npu_inst_pe_1_2_4_n1), .B1(npu_inst_pe_1_2_4_N78), .B2(
        npu_inst_pe_1_2_4_n76), .C1(npu_inst_pe_1_2_4_N70), .C2(
        npu_inst_pe_1_2_4_n77), .ZN(npu_inst_pe_1_2_4_n79) );
  INV_X1 npu_inst_pe_1_2_4_U38 ( .A(npu_inst_pe_1_2_4_n79), .ZN(
        npu_inst_pe_1_2_4_n35) );
  AOI222_X1 npu_inst_pe_1_2_4_U37 ( .A1(npu_inst_int_data_res_3__4__6_), .A2(
        npu_inst_pe_1_2_4_n1), .B1(npu_inst_pe_1_2_4_N79), .B2(
        npu_inst_pe_1_2_4_n76), .C1(npu_inst_pe_1_2_4_N71), .C2(
        npu_inst_pe_1_2_4_n77), .ZN(npu_inst_pe_1_2_4_n78) );
  INV_X1 npu_inst_pe_1_2_4_U36 ( .A(npu_inst_pe_1_2_4_n78), .ZN(
        npu_inst_pe_1_2_4_n34) );
  INV_X1 npu_inst_pe_1_2_4_U35 ( .A(npu_inst_pe_1_2_4_int_data_1_), .ZN(
        npu_inst_pe_1_2_4_n14) );
  AND2_X1 npu_inst_pe_1_2_4_U34 ( .A1(npu_inst_int_data_x_2__4__1_), .A2(
        npu_inst_pe_1_2_4_int_q_weight_1_), .ZN(npu_inst_pe_1_2_4_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_2_4_U33 ( .A1(npu_inst_int_data_x_2__4__0_), .A2(
        npu_inst_pe_1_2_4_int_q_weight_1_), .ZN(npu_inst_pe_1_2_4_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_2_4_U32 ( .A1(npu_inst_n58), .A2(
        npu_inst_int_data_y_3__4__1_), .B1(npu_inst_pe_1_2_4_n3), .B2(
        npu_inst_int_data_x_2__5__1_), .ZN(npu_inst_pe_1_2_4_n63) );
  AOI22_X1 npu_inst_pe_1_2_4_U31 ( .A1(npu_inst_n58), .A2(
        npu_inst_int_data_y_3__4__0_), .B1(npu_inst_pe_1_2_4_n3), .B2(
        npu_inst_int_data_x_2__5__0_), .ZN(npu_inst_pe_1_2_4_n61) );
  INV_X1 npu_inst_pe_1_2_4_U30 ( .A(npu_inst_pe_1_2_4_int_data_0_), .ZN(
        npu_inst_pe_1_2_4_n13) );
  INV_X1 npu_inst_pe_1_2_4_U29 ( .A(npu_inst_n70), .ZN(npu_inst_pe_1_2_4_n5)
         );
  OR3_X1 npu_inst_pe_1_2_4_U28 ( .A1(npu_inst_pe_1_2_4_n6), .A2(
        npu_inst_pe_1_2_4_n8), .A3(npu_inst_pe_1_2_4_n5), .ZN(
        npu_inst_pe_1_2_4_n56) );
  OR3_X1 npu_inst_pe_1_2_4_U27 ( .A1(npu_inst_pe_1_2_4_n5), .A2(
        npu_inst_pe_1_2_4_n8), .A3(npu_inst_pe_1_2_4_n7), .ZN(
        npu_inst_pe_1_2_4_n48) );
  INV_X1 npu_inst_pe_1_2_4_U26 ( .A(npu_inst_pe_1_2_4_n5), .ZN(
        npu_inst_pe_1_2_4_n4) );
  OR3_X1 npu_inst_pe_1_2_4_U25 ( .A1(npu_inst_pe_1_2_4_n4), .A2(
        npu_inst_pe_1_2_4_n8), .A3(npu_inst_pe_1_2_4_n7), .ZN(
        npu_inst_pe_1_2_4_n52) );
  OR3_X1 npu_inst_pe_1_2_4_U24 ( .A1(npu_inst_pe_1_2_4_n6), .A2(
        npu_inst_pe_1_2_4_n8), .A3(npu_inst_pe_1_2_4_n4), .ZN(
        npu_inst_pe_1_2_4_n60) );
  NOR2_X1 npu_inst_pe_1_2_4_U23 ( .A1(npu_inst_pe_1_2_4_n60), .A2(
        npu_inst_pe_1_2_4_n3), .ZN(npu_inst_pe_1_2_4_n58) );
  NOR2_X1 npu_inst_pe_1_2_4_U22 ( .A1(npu_inst_pe_1_2_4_n56), .A2(
        npu_inst_pe_1_2_4_n3), .ZN(npu_inst_pe_1_2_4_n54) );
  NOR2_X1 npu_inst_pe_1_2_4_U21 ( .A1(npu_inst_pe_1_2_4_n52), .A2(
        npu_inst_pe_1_2_4_n3), .ZN(npu_inst_pe_1_2_4_n50) );
  NOR2_X1 npu_inst_pe_1_2_4_U20 ( .A1(npu_inst_pe_1_2_4_n48), .A2(
        npu_inst_pe_1_2_4_n3), .ZN(npu_inst_pe_1_2_4_n46) );
  NOR2_X1 npu_inst_pe_1_2_4_U19 ( .A1(npu_inst_pe_1_2_4_n40), .A2(
        npu_inst_pe_1_2_4_n3), .ZN(npu_inst_pe_1_2_4_n38) );
  NOR2_X1 npu_inst_pe_1_2_4_U18 ( .A1(npu_inst_pe_1_2_4_n44), .A2(
        npu_inst_pe_1_2_4_n3), .ZN(npu_inst_pe_1_2_4_n42) );
  BUF_X1 npu_inst_pe_1_2_4_U17 ( .A(npu_inst_n102), .Z(npu_inst_pe_1_2_4_n8)
         );
  INV_X1 npu_inst_pe_1_2_4_U16 ( .A(npu_inst_n125), .ZN(npu_inst_pe_1_2_4_n12)
         );
  INV_X1 npu_inst_pe_1_2_4_U15 ( .A(npu_inst_pe_1_2_4_n38), .ZN(
        npu_inst_pe_1_2_4_n114) );
  INV_X1 npu_inst_pe_1_2_4_U14 ( .A(npu_inst_pe_1_2_4_n58), .ZN(
        npu_inst_pe_1_2_4_n119) );
  INV_X1 npu_inst_pe_1_2_4_U13 ( .A(npu_inst_pe_1_2_4_n54), .ZN(
        npu_inst_pe_1_2_4_n118) );
  INV_X1 npu_inst_pe_1_2_4_U12 ( .A(npu_inst_pe_1_2_4_n50), .ZN(
        npu_inst_pe_1_2_4_n117) );
  INV_X1 npu_inst_pe_1_2_4_U11 ( .A(npu_inst_pe_1_2_4_n46), .ZN(
        npu_inst_pe_1_2_4_n116) );
  INV_X1 npu_inst_pe_1_2_4_U10 ( .A(npu_inst_pe_1_2_4_n42), .ZN(
        npu_inst_pe_1_2_4_n115) );
  BUF_X1 npu_inst_pe_1_2_4_U9 ( .A(npu_inst_n28), .Z(npu_inst_pe_1_2_4_n2) );
  BUF_X1 npu_inst_pe_1_2_4_U8 ( .A(npu_inst_n28), .Z(npu_inst_pe_1_2_4_n1) );
  BUF_X1 npu_inst_pe_1_2_4_U7 ( .A(npu_inst_pe_1_2_4_n12), .Z(
        npu_inst_pe_1_2_4_n11) );
  BUF_X1 npu_inst_pe_1_2_4_U6 ( .A(npu_inst_pe_1_2_4_n12), .Z(
        npu_inst_pe_1_2_4_n10) );
  BUF_X1 npu_inst_pe_1_2_4_U5 ( .A(npu_inst_pe_1_2_4_n12), .Z(
        npu_inst_pe_1_2_4_n9) );
  NOR2_X1 npu_inst_pe_1_2_4_U4 ( .A1(npu_inst_pe_1_2_4_int_q_weight_0_), .A2(
        npu_inst_pe_1_2_4_n1), .ZN(npu_inst_pe_1_2_4_n76) );
  NOR2_X1 npu_inst_pe_1_2_4_U3 ( .A1(npu_inst_pe_1_2_4_n27), .A2(
        npu_inst_pe_1_2_4_n1), .ZN(npu_inst_pe_1_2_4_n77) );
  FA_X1 npu_inst_pe_1_2_4_sub_67_U2_1 ( .A(npu_inst_pe_1_2_4_int_q_acc_1_), 
        .B(npu_inst_pe_1_2_4_n14), .CI(npu_inst_pe_1_2_4_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_2_4_sub_67_carry_2_), .S(npu_inst_pe_1_2_4_N66) );
  FA_X1 npu_inst_pe_1_2_4_add_69_U1_1 ( .A(npu_inst_pe_1_2_4_int_q_acc_1_), 
        .B(npu_inst_pe_1_2_4_int_data_1_), .CI(
        npu_inst_pe_1_2_4_add_69_carry_1_), .CO(
        npu_inst_pe_1_2_4_add_69_carry_2_), .S(npu_inst_pe_1_2_4_N74) );
  NAND3_X1 npu_inst_pe_1_2_4_U109 ( .A1(npu_inst_pe_1_2_4_n5), .A2(
        npu_inst_pe_1_2_4_n7), .A3(npu_inst_pe_1_2_4_n8), .ZN(
        npu_inst_pe_1_2_4_n44) );
  NAND3_X1 npu_inst_pe_1_2_4_U108 ( .A1(npu_inst_pe_1_2_4_n4), .A2(
        npu_inst_pe_1_2_4_n7), .A3(npu_inst_pe_1_2_4_n8), .ZN(
        npu_inst_pe_1_2_4_n40) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_2_4_n34), .CK(
        npu_inst_pe_1_2_4_net4102), .RN(npu_inst_pe_1_2_4_n9), .Q(
        npu_inst_pe_1_2_4_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_2_4_n35), .CK(
        npu_inst_pe_1_2_4_net4102), .RN(npu_inst_pe_1_2_4_n9), .Q(
        npu_inst_pe_1_2_4_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_2_4_n36), .CK(
        npu_inst_pe_1_2_4_net4102), .RN(npu_inst_pe_1_2_4_n9), .Q(
        npu_inst_pe_1_2_4_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_2_4_n98), .CK(
        npu_inst_pe_1_2_4_net4102), .RN(npu_inst_pe_1_2_4_n9), .Q(
        npu_inst_pe_1_2_4_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_2_4_n99), .CK(
        npu_inst_pe_1_2_4_net4102), .RN(npu_inst_pe_1_2_4_n9), .Q(
        npu_inst_pe_1_2_4_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_2_4_n100), 
        .CK(npu_inst_pe_1_2_4_net4102), .RN(npu_inst_pe_1_2_4_n9), .Q(
        npu_inst_pe_1_2_4_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_2_4_n33), .CK(
        npu_inst_pe_1_2_4_net4102), .RN(npu_inst_pe_1_2_4_n9), .Q(
        npu_inst_pe_1_2_4_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_2_4_n101), 
        .CK(npu_inst_pe_1_2_4_net4102), .RN(npu_inst_pe_1_2_4_n9), .Q(
        npu_inst_pe_1_2_4_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_weight_reg_0_ ( .D(npu_inst_n111), .CK(
        npu_inst_pe_1_2_4_net4108), .RN(npu_inst_pe_1_2_4_n9), .Q(
        npu_inst_pe_1_2_4_int_q_weight_0_), .QN(npu_inst_pe_1_2_4_n27) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_weight_reg_1_ ( .D(npu_inst_n117), .CK(
        npu_inst_pe_1_2_4_net4108), .RN(npu_inst_pe_1_2_4_n9), .Q(
        npu_inst_pe_1_2_4_int_q_weight_1_), .QN(npu_inst_pe_1_2_4_n26) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_2_4_n113), 
        .CK(npu_inst_pe_1_2_4_net4108), .RN(npu_inst_pe_1_2_4_n9), .Q(
        npu_inst_pe_1_2_4_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_2_4_n107), 
        .CK(npu_inst_pe_1_2_4_net4108), .RN(npu_inst_pe_1_2_4_n9), .Q(
        npu_inst_pe_1_2_4_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_2_4_n112), 
        .CK(npu_inst_pe_1_2_4_net4108), .RN(npu_inst_pe_1_2_4_n10), .Q(
        npu_inst_pe_1_2_4_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_2_4_n106), 
        .CK(npu_inst_pe_1_2_4_net4108), .RN(npu_inst_pe_1_2_4_n10), .Q(
        npu_inst_pe_1_2_4_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_2_4_n111), 
        .CK(npu_inst_pe_1_2_4_net4108), .RN(npu_inst_pe_1_2_4_n10), .Q(
        npu_inst_pe_1_2_4_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_2_4_n105), 
        .CK(npu_inst_pe_1_2_4_net4108), .RN(npu_inst_pe_1_2_4_n10), .Q(
        npu_inst_pe_1_2_4_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_2_4_n110), 
        .CK(npu_inst_pe_1_2_4_net4108), .RN(npu_inst_pe_1_2_4_n10), .Q(
        npu_inst_pe_1_2_4_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_2_4_n104), 
        .CK(npu_inst_pe_1_2_4_net4108), .RN(npu_inst_pe_1_2_4_n10), .Q(
        npu_inst_pe_1_2_4_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_2_4_n109), 
        .CK(npu_inst_pe_1_2_4_net4108), .RN(npu_inst_pe_1_2_4_n10), .Q(
        npu_inst_pe_1_2_4_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_2_4_n103), 
        .CK(npu_inst_pe_1_2_4_net4108), .RN(npu_inst_pe_1_2_4_n10), .Q(
        npu_inst_pe_1_2_4_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_2_4_n108), 
        .CK(npu_inst_pe_1_2_4_net4108), .RN(npu_inst_pe_1_2_4_n10), .Q(
        npu_inst_pe_1_2_4_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_2_4_n102), 
        .CK(npu_inst_pe_1_2_4_net4108), .RN(npu_inst_pe_1_2_4_n10), .Q(
        npu_inst_pe_1_2_4_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_2_4_n86), 
        .CK(npu_inst_pe_1_2_4_net4108), .RN(npu_inst_pe_1_2_4_n10), .Q(
        npu_inst_pe_1_2_4_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_2_4_n87), 
        .CK(npu_inst_pe_1_2_4_net4108), .RN(npu_inst_pe_1_2_4_n10), .Q(
        npu_inst_pe_1_2_4_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_2_4_n88), 
        .CK(npu_inst_pe_1_2_4_net4108), .RN(npu_inst_pe_1_2_4_n11), .Q(
        npu_inst_pe_1_2_4_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_2_4_n89), 
        .CK(npu_inst_pe_1_2_4_net4108), .RN(npu_inst_pe_1_2_4_n11), .Q(
        npu_inst_pe_1_2_4_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_2_4_n90), 
        .CK(npu_inst_pe_1_2_4_net4108), .RN(npu_inst_pe_1_2_4_n11), .Q(
        npu_inst_pe_1_2_4_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_2_4_n91), 
        .CK(npu_inst_pe_1_2_4_net4108), .RN(npu_inst_pe_1_2_4_n11), .Q(
        npu_inst_pe_1_2_4_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_2_4_n92), 
        .CK(npu_inst_pe_1_2_4_net4108), .RN(npu_inst_pe_1_2_4_n11), .Q(
        npu_inst_pe_1_2_4_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_2_4_n93), 
        .CK(npu_inst_pe_1_2_4_net4108), .RN(npu_inst_pe_1_2_4_n11), .Q(
        npu_inst_pe_1_2_4_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_2_4_n94), 
        .CK(npu_inst_pe_1_2_4_net4108), .RN(npu_inst_pe_1_2_4_n11), .Q(
        npu_inst_pe_1_2_4_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_2_4_n95), 
        .CK(npu_inst_pe_1_2_4_net4108), .RN(npu_inst_pe_1_2_4_n11), .Q(
        npu_inst_pe_1_2_4_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_2_4_n96), 
        .CK(npu_inst_pe_1_2_4_net4108), .RN(npu_inst_pe_1_2_4_n11), .Q(
        npu_inst_pe_1_2_4_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_2_4_n97), 
        .CK(npu_inst_pe_1_2_4_net4108), .RN(npu_inst_pe_1_2_4_n11), .Q(
        npu_inst_pe_1_2_4_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_2_4_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_2_4_N84), .SE(1'b0), .GCK(npu_inst_pe_1_2_4_net4102) );
  CLKGATETST_X1 npu_inst_pe_1_2_4_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n64), .SE(1'b0), .GCK(npu_inst_pe_1_2_4_net4108) );
  MUX2_X1 npu_inst_pe_1_2_5_U162 ( .A(npu_inst_pe_1_2_5_n32), .B(
        npu_inst_pe_1_2_5_n29), .S(npu_inst_pe_1_2_5_n8), .Z(
        npu_inst_pe_1_2_5_N93) );
  MUX2_X1 npu_inst_pe_1_2_5_U161 ( .A(npu_inst_pe_1_2_5_n31), .B(
        npu_inst_pe_1_2_5_n30), .S(npu_inst_pe_1_2_5_n6), .Z(
        npu_inst_pe_1_2_5_n32) );
  MUX2_X1 npu_inst_pe_1_2_5_U160 ( .A(npu_inst_pe_1_2_5_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_2_5_int_q_reg_v_1__0_), .S(npu_inst_pe_1_2_5_n4), .Z(
        npu_inst_pe_1_2_5_n31) );
  MUX2_X1 npu_inst_pe_1_2_5_U159 ( .A(npu_inst_pe_1_2_5_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_2_5_int_q_reg_v_3__0_), .S(npu_inst_pe_1_2_5_n4), .Z(
        npu_inst_pe_1_2_5_n30) );
  MUX2_X1 npu_inst_pe_1_2_5_U158 ( .A(npu_inst_pe_1_2_5_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_2_5_int_q_reg_v_5__0_), .S(npu_inst_pe_1_2_5_n4), .Z(
        npu_inst_pe_1_2_5_n29) );
  MUX2_X1 npu_inst_pe_1_2_5_U157 ( .A(npu_inst_pe_1_2_5_n28), .B(
        npu_inst_pe_1_2_5_n23), .S(npu_inst_pe_1_2_5_n8), .Z(
        npu_inst_pe_1_2_5_N94) );
  MUX2_X1 npu_inst_pe_1_2_5_U156 ( .A(npu_inst_pe_1_2_5_n25), .B(
        npu_inst_pe_1_2_5_n24), .S(npu_inst_pe_1_2_5_n6), .Z(
        npu_inst_pe_1_2_5_n28) );
  MUX2_X1 npu_inst_pe_1_2_5_U155 ( .A(npu_inst_pe_1_2_5_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_2_5_int_q_reg_v_1__1_), .S(npu_inst_pe_1_2_5_n4), .Z(
        npu_inst_pe_1_2_5_n25) );
  MUX2_X1 npu_inst_pe_1_2_5_U154 ( .A(npu_inst_pe_1_2_5_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_2_5_int_q_reg_v_3__1_), .S(npu_inst_pe_1_2_5_n4), .Z(
        npu_inst_pe_1_2_5_n24) );
  MUX2_X1 npu_inst_pe_1_2_5_U153 ( .A(npu_inst_pe_1_2_5_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_2_5_int_q_reg_v_5__1_), .S(npu_inst_pe_1_2_5_n4), .Z(
        npu_inst_pe_1_2_5_n23) );
  MUX2_X1 npu_inst_pe_1_2_5_U152 ( .A(npu_inst_pe_1_2_5_n22), .B(
        npu_inst_pe_1_2_5_n19), .S(npu_inst_pe_1_2_5_n8), .Z(
        npu_inst_int_data_x_2__5__1_) );
  MUX2_X1 npu_inst_pe_1_2_5_U151 ( .A(npu_inst_pe_1_2_5_n21), .B(
        npu_inst_pe_1_2_5_n20), .S(npu_inst_pe_1_2_5_n6), .Z(
        npu_inst_pe_1_2_5_n22) );
  MUX2_X1 npu_inst_pe_1_2_5_U150 ( .A(npu_inst_pe_1_2_5_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_2_5_int_q_reg_h_1__1_), .S(npu_inst_pe_1_2_5_n4), .Z(
        npu_inst_pe_1_2_5_n21) );
  MUX2_X1 npu_inst_pe_1_2_5_U149 ( .A(npu_inst_pe_1_2_5_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_2_5_int_q_reg_h_3__1_), .S(npu_inst_pe_1_2_5_n4), .Z(
        npu_inst_pe_1_2_5_n20) );
  MUX2_X1 npu_inst_pe_1_2_5_U148 ( .A(npu_inst_pe_1_2_5_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_2_5_int_q_reg_h_5__1_), .S(npu_inst_pe_1_2_5_n4), .Z(
        npu_inst_pe_1_2_5_n19) );
  MUX2_X1 npu_inst_pe_1_2_5_U147 ( .A(npu_inst_pe_1_2_5_n18), .B(
        npu_inst_pe_1_2_5_n15), .S(npu_inst_pe_1_2_5_n8), .Z(
        npu_inst_int_data_x_2__5__0_) );
  MUX2_X1 npu_inst_pe_1_2_5_U146 ( .A(npu_inst_pe_1_2_5_n17), .B(
        npu_inst_pe_1_2_5_n16), .S(npu_inst_pe_1_2_5_n6), .Z(
        npu_inst_pe_1_2_5_n18) );
  MUX2_X1 npu_inst_pe_1_2_5_U145 ( .A(npu_inst_pe_1_2_5_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_2_5_int_q_reg_h_1__0_), .S(npu_inst_pe_1_2_5_n4), .Z(
        npu_inst_pe_1_2_5_n17) );
  MUX2_X1 npu_inst_pe_1_2_5_U144 ( .A(npu_inst_pe_1_2_5_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_2_5_int_q_reg_h_3__0_), .S(npu_inst_pe_1_2_5_n4), .Z(
        npu_inst_pe_1_2_5_n16) );
  MUX2_X1 npu_inst_pe_1_2_5_U143 ( .A(npu_inst_pe_1_2_5_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_2_5_int_q_reg_h_5__0_), .S(npu_inst_pe_1_2_5_n4), .Z(
        npu_inst_pe_1_2_5_n15) );
  XOR2_X1 npu_inst_pe_1_2_5_U142 ( .A(npu_inst_pe_1_2_5_int_data_0_), .B(
        npu_inst_pe_1_2_5_int_q_acc_0_), .Z(npu_inst_pe_1_2_5_N73) );
  AND2_X1 npu_inst_pe_1_2_5_U141 ( .A1(npu_inst_pe_1_2_5_int_q_acc_0_), .A2(
        npu_inst_pe_1_2_5_int_data_0_), .ZN(npu_inst_pe_1_2_5_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_2_5_U140 ( .A(npu_inst_pe_1_2_5_int_q_acc_0_), .B(
        npu_inst_pe_1_2_5_n13), .ZN(npu_inst_pe_1_2_5_N65) );
  OR2_X1 npu_inst_pe_1_2_5_U139 ( .A1(npu_inst_pe_1_2_5_n13), .A2(
        npu_inst_pe_1_2_5_int_q_acc_0_), .ZN(npu_inst_pe_1_2_5_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_2_5_U138 ( .A(npu_inst_pe_1_2_5_int_q_acc_2_), .B(
        npu_inst_pe_1_2_5_add_69_carry_2_), .Z(npu_inst_pe_1_2_5_N75) );
  AND2_X1 npu_inst_pe_1_2_5_U137 ( .A1(npu_inst_pe_1_2_5_add_69_carry_2_), 
        .A2(npu_inst_pe_1_2_5_int_q_acc_2_), .ZN(
        npu_inst_pe_1_2_5_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_2_5_U136 ( .A(npu_inst_pe_1_2_5_int_q_acc_3_), .B(
        npu_inst_pe_1_2_5_add_69_carry_3_), .Z(npu_inst_pe_1_2_5_N76) );
  AND2_X1 npu_inst_pe_1_2_5_U135 ( .A1(npu_inst_pe_1_2_5_add_69_carry_3_), 
        .A2(npu_inst_pe_1_2_5_int_q_acc_3_), .ZN(
        npu_inst_pe_1_2_5_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_2_5_U134 ( .A(npu_inst_pe_1_2_5_int_q_acc_4_), .B(
        npu_inst_pe_1_2_5_add_69_carry_4_), .Z(npu_inst_pe_1_2_5_N77) );
  AND2_X1 npu_inst_pe_1_2_5_U133 ( .A1(npu_inst_pe_1_2_5_add_69_carry_4_), 
        .A2(npu_inst_pe_1_2_5_int_q_acc_4_), .ZN(
        npu_inst_pe_1_2_5_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_2_5_U132 ( .A(npu_inst_pe_1_2_5_int_q_acc_5_), .B(
        npu_inst_pe_1_2_5_add_69_carry_5_), .Z(npu_inst_pe_1_2_5_N78) );
  AND2_X1 npu_inst_pe_1_2_5_U131 ( .A1(npu_inst_pe_1_2_5_add_69_carry_5_), 
        .A2(npu_inst_pe_1_2_5_int_q_acc_5_), .ZN(
        npu_inst_pe_1_2_5_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_2_5_U130 ( .A(npu_inst_pe_1_2_5_int_q_acc_6_), .B(
        npu_inst_pe_1_2_5_add_69_carry_6_), .Z(npu_inst_pe_1_2_5_N79) );
  AND2_X1 npu_inst_pe_1_2_5_U129 ( .A1(npu_inst_pe_1_2_5_add_69_carry_6_), 
        .A2(npu_inst_pe_1_2_5_int_q_acc_6_), .ZN(
        npu_inst_pe_1_2_5_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_2_5_U128 ( .A(npu_inst_pe_1_2_5_int_q_acc_7_), .B(
        npu_inst_pe_1_2_5_add_69_carry_7_), .Z(npu_inst_pe_1_2_5_N80) );
  XNOR2_X1 npu_inst_pe_1_2_5_U127 ( .A(npu_inst_pe_1_2_5_sub_67_carry_2_), .B(
        npu_inst_pe_1_2_5_int_q_acc_2_), .ZN(npu_inst_pe_1_2_5_N67) );
  OR2_X1 npu_inst_pe_1_2_5_U126 ( .A1(npu_inst_pe_1_2_5_int_q_acc_2_), .A2(
        npu_inst_pe_1_2_5_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_2_5_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_2_5_U125 ( .A(npu_inst_pe_1_2_5_sub_67_carry_3_), .B(
        npu_inst_pe_1_2_5_int_q_acc_3_), .ZN(npu_inst_pe_1_2_5_N68) );
  OR2_X1 npu_inst_pe_1_2_5_U124 ( .A1(npu_inst_pe_1_2_5_int_q_acc_3_), .A2(
        npu_inst_pe_1_2_5_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_2_5_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_2_5_U123 ( .A(npu_inst_pe_1_2_5_sub_67_carry_4_), .B(
        npu_inst_pe_1_2_5_int_q_acc_4_), .ZN(npu_inst_pe_1_2_5_N69) );
  OR2_X1 npu_inst_pe_1_2_5_U122 ( .A1(npu_inst_pe_1_2_5_int_q_acc_4_), .A2(
        npu_inst_pe_1_2_5_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_2_5_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_2_5_U121 ( .A(npu_inst_pe_1_2_5_sub_67_carry_5_), .B(
        npu_inst_pe_1_2_5_int_q_acc_5_), .ZN(npu_inst_pe_1_2_5_N70) );
  OR2_X1 npu_inst_pe_1_2_5_U120 ( .A1(npu_inst_pe_1_2_5_int_q_acc_5_), .A2(
        npu_inst_pe_1_2_5_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_2_5_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_2_5_U119 ( .A(npu_inst_pe_1_2_5_sub_67_carry_6_), .B(
        npu_inst_pe_1_2_5_int_q_acc_6_), .ZN(npu_inst_pe_1_2_5_N71) );
  OR2_X1 npu_inst_pe_1_2_5_U118 ( .A1(npu_inst_pe_1_2_5_int_q_acc_6_), .A2(
        npu_inst_pe_1_2_5_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_2_5_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_2_5_U117 ( .A(npu_inst_pe_1_2_5_int_q_acc_7_), .B(
        npu_inst_pe_1_2_5_sub_67_carry_7_), .ZN(npu_inst_pe_1_2_5_N72) );
  INV_X1 npu_inst_pe_1_2_5_U116 ( .A(npu_inst_n78), .ZN(npu_inst_pe_1_2_5_n7)
         );
  INV_X1 npu_inst_pe_1_2_5_U115 ( .A(npu_inst_pe_1_2_5_n7), .ZN(
        npu_inst_pe_1_2_5_n6) );
  INV_X1 npu_inst_pe_1_2_5_U114 ( .A(npu_inst_n58), .ZN(npu_inst_pe_1_2_5_n3)
         );
  AOI22_X1 npu_inst_pe_1_2_5_U113 ( .A1(npu_inst_int_data_y_3__5__0_), .A2(
        npu_inst_pe_1_2_5_n58), .B1(npu_inst_pe_1_2_5_n119), .B2(
        npu_inst_pe_1_2_5_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_2_5_n57) );
  INV_X1 npu_inst_pe_1_2_5_U112 ( .A(npu_inst_pe_1_2_5_n57), .ZN(
        npu_inst_pe_1_2_5_n108) );
  AOI22_X1 npu_inst_pe_1_2_5_U111 ( .A1(npu_inst_int_data_y_3__5__0_), .A2(
        npu_inst_pe_1_2_5_n54), .B1(npu_inst_pe_1_2_5_n118), .B2(
        npu_inst_pe_1_2_5_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_2_5_n53) );
  INV_X1 npu_inst_pe_1_2_5_U110 ( .A(npu_inst_pe_1_2_5_n53), .ZN(
        npu_inst_pe_1_2_5_n109) );
  AOI22_X1 npu_inst_pe_1_2_5_U107 ( .A1(npu_inst_int_data_y_3__5__0_), .A2(
        npu_inst_pe_1_2_5_n50), .B1(npu_inst_pe_1_2_5_n117), .B2(
        npu_inst_pe_1_2_5_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_2_5_n49) );
  INV_X1 npu_inst_pe_1_2_5_U106 ( .A(npu_inst_pe_1_2_5_n49), .ZN(
        npu_inst_pe_1_2_5_n110) );
  AOI22_X1 npu_inst_pe_1_2_5_U105 ( .A1(npu_inst_int_data_y_3__5__0_), .A2(
        npu_inst_pe_1_2_5_n46), .B1(npu_inst_pe_1_2_5_n116), .B2(
        npu_inst_pe_1_2_5_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_2_5_n45) );
  INV_X1 npu_inst_pe_1_2_5_U104 ( .A(npu_inst_pe_1_2_5_n45), .ZN(
        npu_inst_pe_1_2_5_n111) );
  AOI22_X1 npu_inst_pe_1_2_5_U103 ( .A1(npu_inst_int_data_y_3__5__0_), .A2(
        npu_inst_pe_1_2_5_n42), .B1(npu_inst_pe_1_2_5_n115), .B2(
        npu_inst_pe_1_2_5_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_2_5_n41) );
  INV_X1 npu_inst_pe_1_2_5_U102 ( .A(npu_inst_pe_1_2_5_n41), .ZN(
        npu_inst_pe_1_2_5_n112) );
  AOI22_X1 npu_inst_pe_1_2_5_U101 ( .A1(npu_inst_int_data_y_3__5__1_), .A2(
        npu_inst_pe_1_2_5_n58), .B1(npu_inst_pe_1_2_5_n119), .B2(
        npu_inst_pe_1_2_5_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_2_5_n59) );
  INV_X1 npu_inst_pe_1_2_5_U100 ( .A(npu_inst_pe_1_2_5_n59), .ZN(
        npu_inst_pe_1_2_5_n102) );
  AOI22_X1 npu_inst_pe_1_2_5_U99 ( .A1(npu_inst_int_data_y_3__5__1_), .A2(
        npu_inst_pe_1_2_5_n54), .B1(npu_inst_pe_1_2_5_n118), .B2(
        npu_inst_pe_1_2_5_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_2_5_n55) );
  INV_X1 npu_inst_pe_1_2_5_U98 ( .A(npu_inst_pe_1_2_5_n55), .ZN(
        npu_inst_pe_1_2_5_n103) );
  AOI22_X1 npu_inst_pe_1_2_5_U97 ( .A1(npu_inst_int_data_y_3__5__1_), .A2(
        npu_inst_pe_1_2_5_n50), .B1(npu_inst_pe_1_2_5_n117), .B2(
        npu_inst_pe_1_2_5_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_2_5_n51) );
  INV_X1 npu_inst_pe_1_2_5_U96 ( .A(npu_inst_pe_1_2_5_n51), .ZN(
        npu_inst_pe_1_2_5_n104) );
  AOI22_X1 npu_inst_pe_1_2_5_U95 ( .A1(npu_inst_int_data_y_3__5__1_), .A2(
        npu_inst_pe_1_2_5_n46), .B1(npu_inst_pe_1_2_5_n116), .B2(
        npu_inst_pe_1_2_5_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_2_5_n47) );
  INV_X1 npu_inst_pe_1_2_5_U94 ( .A(npu_inst_pe_1_2_5_n47), .ZN(
        npu_inst_pe_1_2_5_n105) );
  AOI22_X1 npu_inst_pe_1_2_5_U93 ( .A1(npu_inst_int_data_y_3__5__1_), .A2(
        npu_inst_pe_1_2_5_n42), .B1(npu_inst_pe_1_2_5_n115), .B2(
        npu_inst_pe_1_2_5_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_2_5_n43) );
  INV_X1 npu_inst_pe_1_2_5_U92 ( .A(npu_inst_pe_1_2_5_n43), .ZN(
        npu_inst_pe_1_2_5_n106) );
  AOI22_X1 npu_inst_pe_1_2_5_U91 ( .A1(npu_inst_pe_1_2_5_n38), .A2(
        npu_inst_int_data_y_3__5__1_), .B1(npu_inst_pe_1_2_5_n114), .B2(
        npu_inst_pe_1_2_5_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_2_5_n39) );
  INV_X1 npu_inst_pe_1_2_5_U90 ( .A(npu_inst_pe_1_2_5_n39), .ZN(
        npu_inst_pe_1_2_5_n107) );
  AOI22_X1 npu_inst_pe_1_2_5_U89 ( .A1(npu_inst_pe_1_2_5_n38), .A2(
        npu_inst_int_data_y_3__5__0_), .B1(npu_inst_pe_1_2_5_n114), .B2(
        npu_inst_pe_1_2_5_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_2_5_n37) );
  INV_X1 npu_inst_pe_1_2_5_U88 ( .A(npu_inst_pe_1_2_5_n37), .ZN(
        npu_inst_pe_1_2_5_n113) );
  NAND2_X1 npu_inst_pe_1_2_5_U87 ( .A1(npu_inst_pe_1_2_5_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_2_5_n60), .ZN(npu_inst_pe_1_2_5_n74) );
  OAI21_X1 npu_inst_pe_1_2_5_U86 ( .B1(npu_inst_pe_1_2_5_n63), .B2(
        npu_inst_pe_1_2_5_n60), .A(npu_inst_pe_1_2_5_n74), .ZN(
        npu_inst_pe_1_2_5_n97) );
  NAND2_X1 npu_inst_pe_1_2_5_U85 ( .A1(npu_inst_pe_1_2_5_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_2_5_n60), .ZN(npu_inst_pe_1_2_5_n73) );
  OAI21_X1 npu_inst_pe_1_2_5_U84 ( .B1(npu_inst_pe_1_2_5_n61), .B2(
        npu_inst_pe_1_2_5_n60), .A(npu_inst_pe_1_2_5_n73), .ZN(
        npu_inst_pe_1_2_5_n96) );
  NAND2_X1 npu_inst_pe_1_2_5_U83 ( .A1(npu_inst_pe_1_2_5_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_2_5_n56), .ZN(npu_inst_pe_1_2_5_n72) );
  OAI21_X1 npu_inst_pe_1_2_5_U82 ( .B1(npu_inst_pe_1_2_5_n63), .B2(
        npu_inst_pe_1_2_5_n56), .A(npu_inst_pe_1_2_5_n72), .ZN(
        npu_inst_pe_1_2_5_n95) );
  NAND2_X1 npu_inst_pe_1_2_5_U81 ( .A1(npu_inst_pe_1_2_5_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_2_5_n56), .ZN(npu_inst_pe_1_2_5_n71) );
  OAI21_X1 npu_inst_pe_1_2_5_U80 ( .B1(npu_inst_pe_1_2_5_n61), .B2(
        npu_inst_pe_1_2_5_n56), .A(npu_inst_pe_1_2_5_n71), .ZN(
        npu_inst_pe_1_2_5_n94) );
  NAND2_X1 npu_inst_pe_1_2_5_U79 ( .A1(npu_inst_pe_1_2_5_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_2_5_n52), .ZN(npu_inst_pe_1_2_5_n70) );
  OAI21_X1 npu_inst_pe_1_2_5_U78 ( .B1(npu_inst_pe_1_2_5_n63), .B2(
        npu_inst_pe_1_2_5_n52), .A(npu_inst_pe_1_2_5_n70), .ZN(
        npu_inst_pe_1_2_5_n93) );
  NAND2_X1 npu_inst_pe_1_2_5_U77 ( .A1(npu_inst_pe_1_2_5_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_2_5_n52), .ZN(npu_inst_pe_1_2_5_n69) );
  OAI21_X1 npu_inst_pe_1_2_5_U76 ( .B1(npu_inst_pe_1_2_5_n61), .B2(
        npu_inst_pe_1_2_5_n52), .A(npu_inst_pe_1_2_5_n69), .ZN(
        npu_inst_pe_1_2_5_n92) );
  NAND2_X1 npu_inst_pe_1_2_5_U75 ( .A1(npu_inst_pe_1_2_5_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_2_5_n48), .ZN(npu_inst_pe_1_2_5_n68) );
  OAI21_X1 npu_inst_pe_1_2_5_U74 ( .B1(npu_inst_pe_1_2_5_n63), .B2(
        npu_inst_pe_1_2_5_n48), .A(npu_inst_pe_1_2_5_n68), .ZN(
        npu_inst_pe_1_2_5_n91) );
  NAND2_X1 npu_inst_pe_1_2_5_U73 ( .A1(npu_inst_pe_1_2_5_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_2_5_n48), .ZN(npu_inst_pe_1_2_5_n67) );
  OAI21_X1 npu_inst_pe_1_2_5_U72 ( .B1(npu_inst_pe_1_2_5_n61), .B2(
        npu_inst_pe_1_2_5_n48), .A(npu_inst_pe_1_2_5_n67), .ZN(
        npu_inst_pe_1_2_5_n90) );
  NAND2_X1 npu_inst_pe_1_2_5_U71 ( .A1(npu_inst_pe_1_2_5_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_2_5_n44), .ZN(npu_inst_pe_1_2_5_n66) );
  OAI21_X1 npu_inst_pe_1_2_5_U70 ( .B1(npu_inst_pe_1_2_5_n63), .B2(
        npu_inst_pe_1_2_5_n44), .A(npu_inst_pe_1_2_5_n66), .ZN(
        npu_inst_pe_1_2_5_n89) );
  NAND2_X1 npu_inst_pe_1_2_5_U69 ( .A1(npu_inst_pe_1_2_5_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_2_5_n44), .ZN(npu_inst_pe_1_2_5_n65) );
  OAI21_X1 npu_inst_pe_1_2_5_U68 ( .B1(npu_inst_pe_1_2_5_n61), .B2(
        npu_inst_pe_1_2_5_n44), .A(npu_inst_pe_1_2_5_n65), .ZN(
        npu_inst_pe_1_2_5_n88) );
  NAND2_X1 npu_inst_pe_1_2_5_U67 ( .A1(npu_inst_pe_1_2_5_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_2_5_n40), .ZN(npu_inst_pe_1_2_5_n64) );
  OAI21_X1 npu_inst_pe_1_2_5_U66 ( .B1(npu_inst_pe_1_2_5_n63), .B2(
        npu_inst_pe_1_2_5_n40), .A(npu_inst_pe_1_2_5_n64), .ZN(
        npu_inst_pe_1_2_5_n87) );
  NAND2_X1 npu_inst_pe_1_2_5_U65 ( .A1(npu_inst_pe_1_2_5_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_2_5_n40), .ZN(npu_inst_pe_1_2_5_n62) );
  OAI21_X1 npu_inst_pe_1_2_5_U64 ( .B1(npu_inst_pe_1_2_5_n61), .B2(
        npu_inst_pe_1_2_5_n40), .A(npu_inst_pe_1_2_5_n62), .ZN(
        npu_inst_pe_1_2_5_n86) );
  AND2_X1 npu_inst_pe_1_2_5_U63 ( .A1(npu_inst_pe_1_2_5_N93), .A2(npu_inst_n58), .ZN(npu_inst_int_data_y_2__5__0_) );
  AND2_X1 npu_inst_pe_1_2_5_U62 ( .A1(npu_inst_n58), .A2(npu_inst_pe_1_2_5_N94), .ZN(npu_inst_int_data_y_2__5__1_) );
  NOR3_X1 npu_inst_pe_1_2_5_U61 ( .A1(npu_inst_pe_1_2_5_n26), .A2(npu_inst_n58), .A3(npu_inst_int_ckg[42]), .ZN(npu_inst_pe_1_2_5_n85) );
  OR2_X1 npu_inst_pe_1_2_5_U60 ( .A1(npu_inst_pe_1_2_5_n85), .A2(
        npu_inst_pe_1_2_5_n2), .ZN(npu_inst_pe_1_2_5_N84) );
  AND2_X1 npu_inst_pe_1_2_5_U59 ( .A1(npu_inst_pe_1_2_5_int_q_acc_0_), .A2(
        npu_inst_pe_1_2_5_n1), .ZN(npu_inst_int_data_res_2__5__0_) );
  AND2_X1 npu_inst_pe_1_2_5_U58 ( .A1(npu_inst_pe_1_2_5_n2), .A2(
        npu_inst_pe_1_2_5_int_q_acc_7_), .ZN(npu_inst_int_data_res_2__5__7_)
         );
  AND2_X1 npu_inst_pe_1_2_5_U57 ( .A1(npu_inst_pe_1_2_5_int_q_acc_1_), .A2(
        npu_inst_pe_1_2_5_n1), .ZN(npu_inst_int_data_res_2__5__1_) );
  AND2_X1 npu_inst_pe_1_2_5_U56 ( .A1(npu_inst_pe_1_2_5_int_q_acc_2_), .A2(
        npu_inst_pe_1_2_5_n1), .ZN(npu_inst_int_data_res_2__5__2_) );
  AND2_X1 npu_inst_pe_1_2_5_U55 ( .A1(npu_inst_pe_1_2_5_int_q_acc_3_), .A2(
        npu_inst_pe_1_2_5_n2), .ZN(npu_inst_int_data_res_2__5__3_) );
  AND2_X1 npu_inst_pe_1_2_5_U54 ( .A1(npu_inst_pe_1_2_5_int_q_acc_4_), .A2(
        npu_inst_pe_1_2_5_n2), .ZN(npu_inst_int_data_res_2__5__4_) );
  AND2_X1 npu_inst_pe_1_2_5_U53 ( .A1(npu_inst_pe_1_2_5_int_q_acc_5_), .A2(
        npu_inst_pe_1_2_5_n2), .ZN(npu_inst_int_data_res_2__5__5_) );
  AND2_X1 npu_inst_pe_1_2_5_U52 ( .A1(npu_inst_pe_1_2_5_int_q_acc_6_), .A2(
        npu_inst_pe_1_2_5_n2), .ZN(npu_inst_int_data_res_2__5__6_) );
  AOI222_X1 npu_inst_pe_1_2_5_U51 ( .A1(npu_inst_int_data_res_3__5__0_), .A2(
        npu_inst_pe_1_2_5_n1), .B1(npu_inst_pe_1_2_5_N73), .B2(
        npu_inst_pe_1_2_5_n76), .C1(npu_inst_pe_1_2_5_N65), .C2(
        npu_inst_pe_1_2_5_n77), .ZN(npu_inst_pe_1_2_5_n84) );
  INV_X1 npu_inst_pe_1_2_5_U50 ( .A(npu_inst_pe_1_2_5_n84), .ZN(
        npu_inst_pe_1_2_5_n101) );
  AOI222_X1 npu_inst_pe_1_2_5_U49 ( .A1(npu_inst_int_data_res_3__5__7_), .A2(
        npu_inst_pe_1_2_5_n1), .B1(npu_inst_pe_1_2_5_N80), .B2(
        npu_inst_pe_1_2_5_n76), .C1(npu_inst_pe_1_2_5_N72), .C2(
        npu_inst_pe_1_2_5_n77), .ZN(npu_inst_pe_1_2_5_n75) );
  INV_X1 npu_inst_pe_1_2_5_U48 ( .A(npu_inst_pe_1_2_5_n75), .ZN(
        npu_inst_pe_1_2_5_n33) );
  AOI222_X1 npu_inst_pe_1_2_5_U47 ( .A1(npu_inst_int_data_res_3__5__1_), .A2(
        npu_inst_pe_1_2_5_n1), .B1(npu_inst_pe_1_2_5_N74), .B2(
        npu_inst_pe_1_2_5_n76), .C1(npu_inst_pe_1_2_5_N66), .C2(
        npu_inst_pe_1_2_5_n77), .ZN(npu_inst_pe_1_2_5_n83) );
  INV_X1 npu_inst_pe_1_2_5_U46 ( .A(npu_inst_pe_1_2_5_n83), .ZN(
        npu_inst_pe_1_2_5_n100) );
  AOI222_X1 npu_inst_pe_1_2_5_U45 ( .A1(npu_inst_int_data_res_3__5__2_), .A2(
        npu_inst_pe_1_2_5_n1), .B1(npu_inst_pe_1_2_5_N75), .B2(
        npu_inst_pe_1_2_5_n76), .C1(npu_inst_pe_1_2_5_N67), .C2(
        npu_inst_pe_1_2_5_n77), .ZN(npu_inst_pe_1_2_5_n82) );
  INV_X1 npu_inst_pe_1_2_5_U44 ( .A(npu_inst_pe_1_2_5_n82), .ZN(
        npu_inst_pe_1_2_5_n99) );
  AOI222_X1 npu_inst_pe_1_2_5_U43 ( .A1(npu_inst_int_data_res_3__5__3_), .A2(
        npu_inst_pe_1_2_5_n1), .B1(npu_inst_pe_1_2_5_N76), .B2(
        npu_inst_pe_1_2_5_n76), .C1(npu_inst_pe_1_2_5_N68), .C2(
        npu_inst_pe_1_2_5_n77), .ZN(npu_inst_pe_1_2_5_n81) );
  INV_X1 npu_inst_pe_1_2_5_U42 ( .A(npu_inst_pe_1_2_5_n81), .ZN(
        npu_inst_pe_1_2_5_n98) );
  AOI222_X1 npu_inst_pe_1_2_5_U41 ( .A1(npu_inst_int_data_res_3__5__4_), .A2(
        npu_inst_pe_1_2_5_n1), .B1(npu_inst_pe_1_2_5_N77), .B2(
        npu_inst_pe_1_2_5_n76), .C1(npu_inst_pe_1_2_5_N69), .C2(
        npu_inst_pe_1_2_5_n77), .ZN(npu_inst_pe_1_2_5_n80) );
  INV_X1 npu_inst_pe_1_2_5_U40 ( .A(npu_inst_pe_1_2_5_n80), .ZN(
        npu_inst_pe_1_2_5_n36) );
  AOI222_X1 npu_inst_pe_1_2_5_U39 ( .A1(npu_inst_int_data_res_3__5__5_), .A2(
        npu_inst_pe_1_2_5_n1), .B1(npu_inst_pe_1_2_5_N78), .B2(
        npu_inst_pe_1_2_5_n76), .C1(npu_inst_pe_1_2_5_N70), .C2(
        npu_inst_pe_1_2_5_n77), .ZN(npu_inst_pe_1_2_5_n79) );
  INV_X1 npu_inst_pe_1_2_5_U38 ( .A(npu_inst_pe_1_2_5_n79), .ZN(
        npu_inst_pe_1_2_5_n35) );
  AOI222_X1 npu_inst_pe_1_2_5_U37 ( .A1(npu_inst_int_data_res_3__5__6_), .A2(
        npu_inst_pe_1_2_5_n1), .B1(npu_inst_pe_1_2_5_N79), .B2(
        npu_inst_pe_1_2_5_n76), .C1(npu_inst_pe_1_2_5_N71), .C2(
        npu_inst_pe_1_2_5_n77), .ZN(npu_inst_pe_1_2_5_n78) );
  INV_X1 npu_inst_pe_1_2_5_U36 ( .A(npu_inst_pe_1_2_5_n78), .ZN(
        npu_inst_pe_1_2_5_n34) );
  INV_X1 npu_inst_pe_1_2_5_U35 ( .A(npu_inst_pe_1_2_5_int_data_1_), .ZN(
        npu_inst_pe_1_2_5_n14) );
  AND2_X1 npu_inst_pe_1_2_5_U34 ( .A1(npu_inst_int_data_x_2__5__1_), .A2(
        npu_inst_pe_1_2_5_int_q_weight_1_), .ZN(npu_inst_pe_1_2_5_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_2_5_U33 ( .A1(npu_inst_int_data_x_2__5__0_), .A2(
        npu_inst_pe_1_2_5_int_q_weight_1_), .ZN(npu_inst_pe_1_2_5_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_2_5_U32 ( .A1(npu_inst_n58), .A2(
        npu_inst_int_data_y_3__5__1_), .B1(npu_inst_pe_1_2_5_n3), .B2(
        npu_inst_int_data_x_2__6__1_), .ZN(npu_inst_pe_1_2_5_n63) );
  AOI22_X1 npu_inst_pe_1_2_5_U31 ( .A1(npu_inst_n58), .A2(
        npu_inst_int_data_y_3__5__0_), .B1(npu_inst_pe_1_2_5_n3), .B2(
        npu_inst_int_data_x_2__6__0_), .ZN(npu_inst_pe_1_2_5_n61) );
  INV_X1 npu_inst_pe_1_2_5_U30 ( .A(npu_inst_pe_1_2_5_int_data_0_), .ZN(
        npu_inst_pe_1_2_5_n13) );
  INV_X1 npu_inst_pe_1_2_5_U29 ( .A(npu_inst_n70), .ZN(npu_inst_pe_1_2_5_n5)
         );
  OR3_X1 npu_inst_pe_1_2_5_U28 ( .A1(npu_inst_pe_1_2_5_n6), .A2(
        npu_inst_pe_1_2_5_n8), .A3(npu_inst_pe_1_2_5_n5), .ZN(
        npu_inst_pe_1_2_5_n56) );
  OR3_X1 npu_inst_pe_1_2_5_U27 ( .A1(npu_inst_pe_1_2_5_n5), .A2(
        npu_inst_pe_1_2_5_n8), .A3(npu_inst_pe_1_2_5_n7), .ZN(
        npu_inst_pe_1_2_5_n48) );
  INV_X1 npu_inst_pe_1_2_5_U26 ( .A(npu_inst_pe_1_2_5_n5), .ZN(
        npu_inst_pe_1_2_5_n4) );
  OR3_X1 npu_inst_pe_1_2_5_U25 ( .A1(npu_inst_pe_1_2_5_n4), .A2(
        npu_inst_pe_1_2_5_n8), .A3(npu_inst_pe_1_2_5_n7), .ZN(
        npu_inst_pe_1_2_5_n52) );
  OR3_X1 npu_inst_pe_1_2_5_U24 ( .A1(npu_inst_pe_1_2_5_n6), .A2(
        npu_inst_pe_1_2_5_n8), .A3(npu_inst_pe_1_2_5_n4), .ZN(
        npu_inst_pe_1_2_5_n60) );
  NOR2_X1 npu_inst_pe_1_2_5_U23 ( .A1(npu_inst_pe_1_2_5_n60), .A2(
        npu_inst_pe_1_2_5_n3), .ZN(npu_inst_pe_1_2_5_n58) );
  NOR2_X1 npu_inst_pe_1_2_5_U22 ( .A1(npu_inst_pe_1_2_5_n56), .A2(
        npu_inst_pe_1_2_5_n3), .ZN(npu_inst_pe_1_2_5_n54) );
  NOR2_X1 npu_inst_pe_1_2_5_U21 ( .A1(npu_inst_pe_1_2_5_n52), .A2(
        npu_inst_pe_1_2_5_n3), .ZN(npu_inst_pe_1_2_5_n50) );
  NOR2_X1 npu_inst_pe_1_2_5_U20 ( .A1(npu_inst_pe_1_2_5_n48), .A2(
        npu_inst_pe_1_2_5_n3), .ZN(npu_inst_pe_1_2_5_n46) );
  NOR2_X1 npu_inst_pe_1_2_5_U19 ( .A1(npu_inst_pe_1_2_5_n40), .A2(
        npu_inst_pe_1_2_5_n3), .ZN(npu_inst_pe_1_2_5_n38) );
  NOR2_X1 npu_inst_pe_1_2_5_U18 ( .A1(npu_inst_pe_1_2_5_n44), .A2(
        npu_inst_pe_1_2_5_n3), .ZN(npu_inst_pe_1_2_5_n42) );
  BUF_X1 npu_inst_pe_1_2_5_U17 ( .A(npu_inst_n102), .Z(npu_inst_pe_1_2_5_n8)
         );
  INV_X1 npu_inst_pe_1_2_5_U16 ( .A(npu_inst_n125), .ZN(npu_inst_pe_1_2_5_n12)
         );
  INV_X1 npu_inst_pe_1_2_5_U15 ( .A(npu_inst_pe_1_2_5_n38), .ZN(
        npu_inst_pe_1_2_5_n114) );
  INV_X1 npu_inst_pe_1_2_5_U14 ( .A(npu_inst_pe_1_2_5_n58), .ZN(
        npu_inst_pe_1_2_5_n119) );
  INV_X1 npu_inst_pe_1_2_5_U13 ( .A(npu_inst_pe_1_2_5_n54), .ZN(
        npu_inst_pe_1_2_5_n118) );
  INV_X1 npu_inst_pe_1_2_5_U12 ( .A(npu_inst_pe_1_2_5_n50), .ZN(
        npu_inst_pe_1_2_5_n117) );
  INV_X1 npu_inst_pe_1_2_5_U11 ( .A(npu_inst_pe_1_2_5_n46), .ZN(
        npu_inst_pe_1_2_5_n116) );
  INV_X1 npu_inst_pe_1_2_5_U10 ( .A(npu_inst_pe_1_2_5_n42), .ZN(
        npu_inst_pe_1_2_5_n115) );
  BUF_X1 npu_inst_pe_1_2_5_U9 ( .A(npu_inst_n28), .Z(npu_inst_pe_1_2_5_n2) );
  BUF_X1 npu_inst_pe_1_2_5_U8 ( .A(npu_inst_n28), .Z(npu_inst_pe_1_2_5_n1) );
  BUF_X1 npu_inst_pe_1_2_5_U7 ( .A(npu_inst_pe_1_2_5_n12), .Z(
        npu_inst_pe_1_2_5_n11) );
  BUF_X1 npu_inst_pe_1_2_5_U6 ( .A(npu_inst_pe_1_2_5_n12), .Z(
        npu_inst_pe_1_2_5_n10) );
  BUF_X1 npu_inst_pe_1_2_5_U5 ( .A(npu_inst_pe_1_2_5_n12), .Z(
        npu_inst_pe_1_2_5_n9) );
  NOR2_X1 npu_inst_pe_1_2_5_U4 ( .A1(npu_inst_pe_1_2_5_int_q_weight_0_), .A2(
        npu_inst_pe_1_2_5_n1), .ZN(npu_inst_pe_1_2_5_n76) );
  NOR2_X1 npu_inst_pe_1_2_5_U3 ( .A1(npu_inst_pe_1_2_5_n27), .A2(
        npu_inst_pe_1_2_5_n1), .ZN(npu_inst_pe_1_2_5_n77) );
  FA_X1 npu_inst_pe_1_2_5_sub_67_U2_1 ( .A(npu_inst_pe_1_2_5_int_q_acc_1_), 
        .B(npu_inst_pe_1_2_5_n14), .CI(npu_inst_pe_1_2_5_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_2_5_sub_67_carry_2_), .S(npu_inst_pe_1_2_5_N66) );
  FA_X1 npu_inst_pe_1_2_5_add_69_U1_1 ( .A(npu_inst_pe_1_2_5_int_q_acc_1_), 
        .B(npu_inst_pe_1_2_5_int_data_1_), .CI(
        npu_inst_pe_1_2_5_add_69_carry_1_), .CO(
        npu_inst_pe_1_2_5_add_69_carry_2_), .S(npu_inst_pe_1_2_5_N74) );
  NAND3_X1 npu_inst_pe_1_2_5_U109 ( .A1(npu_inst_pe_1_2_5_n5), .A2(
        npu_inst_pe_1_2_5_n7), .A3(npu_inst_pe_1_2_5_n8), .ZN(
        npu_inst_pe_1_2_5_n44) );
  NAND3_X1 npu_inst_pe_1_2_5_U108 ( .A1(npu_inst_pe_1_2_5_n4), .A2(
        npu_inst_pe_1_2_5_n7), .A3(npu_inst_pe_1_2_5_n8), .ZN(
        npu_inst_pe_1_2_5_n40) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_2_5_n34), .CK(
        npu_inst_pe_1_2_5_net4079), .RN(npu_inst_pe_1_2_5_n9), .Q(
        npu_inst_pe_1_2_5_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_2_5_n35), .CK(
        npu_inst_pe_1_2_5_net4079), .RN(npu_inst_pe_1_2_5_n9), .Q(
        npu_inst_pe_1_2_5_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_2_5_n36), .CK(
        npu_inst_pe_1_2_5_net4079), .RN(npu_inst_pe_1_2_5_n9), .Q(
        npu_inst_pe_1_2_5_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_2_5_n98), .CK(
        npu_inst_pe_1_2_5_net4079), .RN(npu_inst_pe_1_2_5_n9), .Q(
        npu_inst_pe_1_2_5_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_2_5_n99), .CK(
        npu_inst_pe_1_2_5_net4079), .RN(npu_inst_pe_1_2_5_n9), .Q(
        npu_inst_pe_1_2_5_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_2_5_n100), 
        .CK(npu_inst_pe_1_2_5_net4079), .RN(npu_inst_pe_1_2_5_n9), .Q(
        npu_inst_pe_1_2_5_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_2_5_n33), .CK(
        npu_inst_pe_1_2_5_net4079), .RN(npu_inst_pe_1_2_5_n9), .Q(
        npu_inst_pe_1_2_5_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_2_5_n101), 
        .CK(npu_inst_pe_1_2_5_net4079), .RN(npu_inst_pe_1_2_5_n9), .Q(
        npu_inst_pe_1_2_5_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_weight_reg_0_ ( .D(npu_inst_n111), .CK(
        npu_inst_pe_1_2_5_net4085), .RN(npu_inst_pe_1_2_5_n9), .Q(
        npu_inst_pe_1_2_5_int_q_weight_0_), .QN(npu_inst_pe_1_2_5_n27) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_weight_reg_1_ ( .D(npu_inst_n117), .CK(
        npu_inst_pe_1_2_5_net4085), .RN(npu_inst_pe_1_2_5_n9), .Q(
        npu_inst_pe_1_2_5_int_q_weight_1_), .QN(npu_inst_pe_1_2_5_n26) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_2_5_n113), 
        .CK(npu_inst_pe_1_2_5_net4085), .RN(npu_inst_pe_1_2_5_n9), .Q(
        npu_inst_pe_1_2_5_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_2_5_n107), 
        .CK(npu_inst_pe_1_2_5_net4085), .RN(npu_inst_pe_1_2_5_n9), .Q(
        npu_inst_pe_1_2_5_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_2_5_n112), 
        .CK(npu_inst_pe_1_2_5_net4085), .RN(npu_inst_pe_1_2_5_n10), .Q(
        npu_inst_pe_1_2_5_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_2_5_n106), 
        .CK(npu_inst_pe_1_2_5_net4085), .RN(npu_inst_pe_1_2_5_n10), .Q(
        npu_inst_pe_1_2_5_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_2_5_n111), 
        .CK(npu_inst_pe_1_2_5_net4085), .RN(npu_inst_pe_1_2_5_n10), .Q(
        npu_inst_pe_1_2_5_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_2_5_n105), 
        .CK(npu_inst_pe_1_2_5_net4085), .RN(npu_inst_pe_1_2_5_n10), .Q(
        npu_inst_pe_1_2_5_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_2_5_n110), 
        .CK(npu_inst_pe_1_2_5_net4085), .RN(npu_inst_pe_1_2_5_n10), .Q(
        npu_inst_pe_1_2_5_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_2_5_n104), 
        .CK(npu_inst_pe_1_2_5_net4085), .RN(npu_inst_pe_1_2_5_n10), .Q(
        npu_inst_pe_1_2_5_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_2_5_n109), 
        .CK(npu_inst_pe_1_2_5_net4085), .RN(npu_inst_pe_1_2_5_n10), .Q(
        npu_inst_pe_1_2_5_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_2_5_n103), 
        .CK(npu_inst_pe_1_2_5_net4085), .RN(npu_inst_pe_1_2_5_n10), .Q(
        npu_inst_pe_1_2_5_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_2_5_n108), 
        .CK(npu_inst_pe_1_2_5_net4085), .RN(npu_inst_pe_1_2_5_n10), .Q(
        npu_inst_pe_1_2_5_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_2_5_n102), 
        .CK(npu_inst_pe_1_2_5_net4085), .RN(npu_inst_pe_1_2_5_n10), .Q(
        npu_inst_pe_1_2_5_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_2_5_n86), 
        .CK(npu_inst_pe_1_2_5_net4085), .RN(npu_inst_pe_1_2_5_n10), .Q(
        npu_inst_pe_1_2_5_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_2_5_n87), 
        .CK(npu_inst_pe_1_2_5_net4085), .RN(npu_inst_pe_1_2_5_n10), .Q(
        npu_inst_pe_1_2_5_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_2_5_n88), 
        .CK(npu_inst_pe_1_2_5_net4085), .RN(npu_inst_pe_1_2_5_n11), .Q(
        npu_inst_pe_1_2_5_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_2_5_n89), 
        .CK(npu_inst_pe_1_2_5_net4085), .RN(npu_inst_pe_1_2_5_n11), .Q(
        npu_inst_pe_1_2_5_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_2_5_n90), 
        .CK(npu_inst_pe_1_2_5_net4085), .RN(npu_inst_pe_1_2_5_n11), .Q(
        npu_inst_pe_1_2_5_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_2_5_n91), 
        .CK(npu_inst_pe_1_2_5_net4085), .RN(npu_inst_pe_1_2_5_n11), .Q(
        npu_inst_pe_1_2_5_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_2_5_n92), 
        .CK(npu_inst_pe_1_2_5_net4085), .RN(npu_inst_pe_1_2_5_n11), .Q(
        npu_inst_pe_1_2_5_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_2_5_n93), 
        .CK(npu_inst_pe_1_2_5_net4085), .RN(npu_inst_pe_1_2_5_n11), .Q(
        npu_inst_pe_1_2_5_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_2_5_n94), 
        .CK(npu_inst_pe_1_2_5_net4085), .RN(npu_inst_pe_1_2_5_n11), .Q(
        npu_inst_pe_1_2_5_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_2_5_n95), 
        .CK(npu_inst_pe_1_2_5_net4085), .RN(npu_inst_pe_1_2_5_n11), .Q(
        npu_inst_pe_1_2_5_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_2_5_n96), 
        .CK(npu_inst_pe_1_2_5_net4085), .RN(npu_inst_pe_1_2_5_n11), .Q(
        npu_inst_pe_1_2_5_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_2_5_n97), 
        .CK(npu_inst_pe_1_2_5_net4085), .RN(npu_inst_pe_1_2_5_n11), .Q(
        npu_inst_pe_1_2_5_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_2_5_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_2_5_N84), .SE(1'b0), .GCK(npu_inst_pe_1_2_5_net4079) );
  CLKGATETST_X1 npu_inst_pe_1_2_5_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n64), .SE(1'b0), .GCK(npu_inst_pe_1_2_5_net4085) );
  MUX2_X1 npu_inst_pe_1_2_6_U162 ( .A(npu_inst_pe_1_2_6_n32), .B(
        npu_inst_pe_1_2_6_n29), .S(npu_inst_pe_1_2_6_n8), .Z(
        npu_inst_pe_1_2_6_N93) );
  MUX2_X1 npu_inst_pe_1_2_6_U161 ( .A(npu_inst_pe_1_2_6_n31), .B(
        npu_inst_pe_1_2_6_n30), .S(npu_inst_pe_1_2_6_n6), .Z(
        npu_inst_pe_1_2_6_n32) );
  MUX2_X1 npu_inst_pe_1_2_6_U160 ( .A(npu_inst_pe_1_2_6_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_2_6_int_q_reg_v_1__0_), .S(npu_inst_pe_1_2_6_n4), .Z(
        npu_inst_pe_1_2_6_n31) );
  MUX2_X1 npu_inst_pe_1_2_6_U159 ( .A(npu_inst_pe_1_2_6_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_2_6_int_q_reg_v_3__0_), .S(npu_inst_pe_1_2_6_n4), .Z(
        npu_inst_pe_1_2_6_n30) );
  MUX2_X1 npu_inst_pe_1_2_6_U158 ( .A(npu_inst_pe_1_2_6_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_2_6_int_q_reg_v_5__0_), .S(npu_inst_pe_1_2_6_n4), .Z(
        npu_inst_pe_1_2_6_n29) );
  MUX2_X1 npu_inst_pe_1_2_6_U157 ( .A(npu_inst_pe_1_2_6_n28), .B(
        npu_inst_pe_1_2_6_n23), .S(npu_inst_pe_1_2_6_n8), .Z(
        npu_inst_pe_1_2_6_N94) );
  MUX2_X1 npu_inst_pe_1_2_6_U156 ( .A(npu_inst_pe_1_2_6_n25), .B(
        npu_inst_pe_1_2_6_n24), .S(npu_inst_pe_1_2_6_n6), .Z(
        npu_inst_pe_1_2_6_n28) );
  MUX2_X1 npu_inst_pe_1_2_6_U155 ( .A(npu_inst_pe_1_2_6_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_2_6_int_q_reg_v_1__1_), .S(npu_inst_pe_1_2_6_n4), .Z(
        npu_inst_pe_1_2_6_n25) );
  MUX2_X1 npu_inst_pe_1_2_6_U154 ( .A(npu_inst_pe_1_2_6_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_2_6_int_q_reg_v_3__1_), .S(npu_inst_pe_1_2_6_n4), .Z(
        npu_inst_pe_1_2_6_n24) );
  MUX2_X1 npu_inst_pe_1_2_6_U153 ( .A(npu_inst_pe_1_2_6_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_2_6_int_q_reg_v_5__1_), .S(npu_inst_pe_1_2_6_n4), .Z(
        npu_inst_pe_1_2_6_n23) );
  MUX2_X1 npu_inst_pe_1_2_6_U152 ( .A(npu_inst_pe_1_2_6_n22), .B(
        npu_inst_pe_1_2_6_n19), .S(npu_inst_pe_1_2_6_n8), .Z(
        npu_inst_int_data_x_2__6__1_) );
  MUX2_X1 npu_inst_pe_1_2_6_U151 ( .A(npu_inst_pe_1_2_6_n21), .B(
        npu_inst_pe_1_2_6_n20), .S(npu_inst_pe_1_2_6_n6), .Z(
        npu_inst_pe_1_2_6_n22) );
  MUX2_X1 npu_inst_pe_1_2_6_U150 ( .A(npu_inst_pe_1_2_6_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_2_6_int_q_reg_h_1__1_), .S(npu_inst_pe_1_2_6_n4), .Z(
        npu_inst_pe_1_2_6_n21) );
  MUX2_X1 npu_inst_pe_1_2_6_U149 ( .A(npu_inst_pe_1_2_6_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_2_6_int_q_reg_h_3__1_), .S(npu_inst_pe_1_2_6_n4), .Z(
        npu_inst_pe_1_2_6_n20) );
  MUX2_X1 npu_inst_pe_1_2_6_U148 ( .A(npu_inst_pe_1_2_6_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_2_6_int_q_reg_h_5__1_), .S(npu_inst_pe_1_2_6_n4), .Z(
        npu_inst_pe_1_2_6_n19) );
  MUX2_X1 npu_inst_pe_1_2_6_U147 ( .A(npu_inst_pe_1_2_6_n18), .B(
        npu_inst_pe_1_2_6_n15), .S(npu_inst_pe_1_2_6_n8), .Z(
        npu_inst_int_data_x_2__6__0_) );
  MUX2_X1 npu_inst_pe_1_2_6_U146 ( .A(npu_inst_pe_1_2_6_n17), .B(
        npu_inst_pe_1_2_6_n16), .S(npu_inst_pe_1_2_6_n6), .Z(
        npu_inst_pe_1_2_6_n18) );
  MUX2_X1 npu_inst_pe_1_2_6_U145 ( .A(npu_inst_pe_1_2_6_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_2_6_int_q_reg_h_1__0_), .S(npu_inst_pe_1_2_6_n4), .Z(
        npu_inst_pe_1_2_6_n17) );
  MUX2_X1 npu_inst_pe_1_2_6_U144 ( .A(npu_inst_pe_1_2_6_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_2_6_int_q_reg_h_3__0_), .S(npu_inst_pe_1_2_6_n4), .Z(
        npu_inst_pe_1_2_6_n16) );
  MUX2_X1 npu_inst_pe_1_2_6_U143 ( .A(npu_inst_pe_1_2_6_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_2_6_int_q_reg_h_5__0_), .S(npu_inst_pe_1_2_6_n4), .Z(
        npu_inst_pe_1_2_6_n15) );
  XOR2_X1 npu_inst_pe_1_2_6_U142 ( .A(npu_inst_pe_1_2_6_int_data_0_), .B(
        npu_inst_pe_1_2_6_int_q_acc_0_), .Z(npu_inst_pe_1_2_6_N73) );
  AND2_X1 npu_inst_pe_1_2_6_U141 ( .A1(npu_inst_pe_1_2_6_int_q_acc_0_), .A2(
        npu_inst_pe_1_2_6_int_data_0_), .ZN(npu_inst_pe_1_2_6_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_2_6_U140 ( .A(npu_inst_pe_1_2_6_int_q_acc_0_), .B(
        npu_inst_pe_1_2_6_n13), .ZN(npu_inst_pe_1_2_6_N65) );
  OR2_X1 npu_inst_pe_1_2_6_U139 ( .A1(npu_inst_pe_1_2_6_n13), .A2(
        npu_inst_pe_1_2_6_int_q_acc_0_), .ZN(npu_inst_pe_1_2_6_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_2_6_U138 ( .A(npu_inst_pe_1_2_6_int_q_acc_2_), .B(
        npu_inst_pe_1_2_6_add_69_carry_2_), .Z(npu_inst_pe_1_2_6_N75) );
  AND2_X1 npu_inst_pe_1_2_6_U137 ( .A1(npu_inst_pe_1_2_6_add_69_carry_2_), 
        .A2(npu_inst_pe_1_2_6_int_q_acc_2_), .ZN(
        npu_inst_pe_1_2_6_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_2_6_U136 ( .A(npu_inst_pe_1_2_6_int_q_acc_3_), .B(
        npu_inst_pe_1_2_6_add_69_carry_3_), .Z(npu_inst_pe_1_2_6_N76) );
  AND2_X1 npu_inst_pe_1_2_6_U135 ( .A1(npu_inst_pe_1_2_6_add_69_carry_3_), 
        .A2(npu_inst_pe_1_2_6_int_q_acc_3_), .ZN(
        npu_inst_pe_1_2_6_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_2_6_U134 ( .A(npu_inst_pe_1_2_6_int_q_acc_4_), .B(
        npu_inst_pe_1_2_6_add_69_carry_4_), .Z(npu_inst_pe_1_2_6_N77) );
  AND2_X1 npu_inst_pe_1_2_6_U133 ( .A1(npu_inst_pe_1_2_6_add_69_carry_4_), 
        .A2(npu_inst_pe_1_2_6_int_q_acc_4_), .ZN(
        npu_inst_pe_1_2_6_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_2_6_U132 ( .A(npu_inst_pe_1_2_6_int_q_acc_5_), .B(
        npu_inst_pe_1_2_6_add_69_carry_5_), .Z(npu_inst_pe_1_2_6_N78) );
  AND2_X1 npu_inst_pe_1_2_6_U131 ( .A1(npu_inst_pe_1_2_6_add_69_carry_5_), 
        .A2(npu_inst_pe_1_2_6_int_q_acc_5_), .ZN(
        npu_inst_pe_1_2_6_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_2_6_U130 ( .A(npu_inst_pe_1_2_6_int_q_acc_6_), .B(
        npu_inst_pe_1_2_6_add_69_carry_6_), .Z(npu_inst_pe_1_2_6_N79) );
  AND2_X1 npu_inst_pe_1_2_6_U129 ( .A1(npu_inst_pe_1_2_6_add_69_carry_6_), 
        .A2(npu_inst_pe_1_2_6_int_q_acc_6_), .ZN(
        npu_inst_pe_1_2_6_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_2_6_U128 ( .A(npu_inst_pe_1_2_6_int_q_acc_7_), .B(
        npu_inst_pe_1_2_6_add_69_carry_7_), .Z(npu_inst_pe_1_2_6_N80) );
  XNOR2_X1 npu_inst_pe_1_2_6_U127 ( .A(npu_inst_pe_1_2_6_sub_67_carry_2_), .B(
        npu_inst_pe_1_2_6_int_q_acc_2_), .ZN(npu_inst_pe_1_2_6_N67) );
  OR2_X1 npu_inst_pe_1_2_6_U126 ( .A1(npu_inst_pe_1_2_6_int_q_acc_2_), .A2(
        npu_inst_pe_1_2_6_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_2_6_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_2_6_U125 ( .A(npu_inst_pe_1_2_6_sub_67_carry_3_), .B(
        npu_inst_pe_1_2_6_int_q_acc_3_), .ZN(npu_inst_pe_1_2_6_N68) );
  OR2_X1 npu_inst_pe_1_2_6_U124 ( .A1(npu_inst_pe_1_2_6_int_q_acc_3_), .A2(
        npu_inst_pe_1_2_6_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_2_6_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_2_6_U123 ( .A(npu_inst_pe_1_2_6_sub_67_carry_4_), .B(
        npu_inst_pe_1_2_6_int_q_acc_4_), .ZN(npu_inst_pe_1_2_6_N69) );
  OR2_X1 npu_inst_pe_1_2_6_U122 ( .A1(npu_inst_pe_1_2_6_int_q_acc_4_), .A2(
        npu_inst_pe_1_2_6_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_2_6_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_2_6_U121 ( .A(npu_inst_pe_1_2_6_sub_67_carry_5_), .B(
        npu_inst_pe_1_2_6_int_q_acc_5_), .ZN(npu_inst_pe_1_2_6_N70) );
  OR2_X1 npu_inst_pe_1_2_6_U120 ( .A1(npu_inst_pe_1_2_6_int_q_acc_5_), .A2(
        npu_inst_pe_1_2_6_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_2_6_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_2_6_U119 ( .A(npu_inst_pe_1_2_6_sub_67_carry_6_), .B(
        npu_inst_pe_1_2_6_int_q_acc_6_), .ZN(npu_inst_pe_1_2_6_N71) );
  OR2_X1 npu_inst_pe_1_2_6_U118 ( .A1(npu_inst_pe_1_2_6_int_q_acc_6_), .A2(
        npu_inst_pe_1_2_6_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_2_6_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_2_6_U117 ( .A(npu_inst_pe_1_2_6_int_q_acc_7_), .B(
        npu_inst_pe_1_2_6_sub_67_carry_7_), .ZN(npu_inst_pe_1_2_6_N72) );
  INV_X1 npu_inst_pe_1_2_6_U116 ( .A(npu_inst_n78), .ZN(npu_inst_pe_1_2_6_n7)
         );
  INV_X1 npu_inst_pe_1_2_6_U115 ( .A(npu_inst_pe_1_2_6_n7), .ZN(
        npu_inst_pe_1_2_6_n6) );
  INV_X1 npu_inst_pe_1_2_6_U114 ( .A(npu_inst_n57), .ZN(npu_inst_pe_1_2_6_n3)
         );
  AOI22_X1 npu_inst_pe_1_2_6_U113 ( .A1(npu_inst_int_data_y_3__6__0_), .A2(
        npu_inst_pe_1_2_6_n58), .B1(npu_inst_pe_1_2_6_n119), .B2(
        npu_inst_pe_1_2_6_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_2_6_n57) );
  INV_X1 npu_inst_pe_1_2_6_U112 ( .A(npu_inst_pe_1_2_6_n57), .ZN(
        npu_inst_pe_1_2_6_n108) );
  AOI22_X1 npu_inst_pe_1_2_6_U111 ( .A1(npu_inst_int_data_y_3__6__0_), .A2(
        npu_inst_pe_1_2_6_n54), .B1(npu_inst_pe_1_2_6_n118), .B2(
        npu_inst_pe_1_2_6_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_2_6_n53) );
  INV_X1 npu_inst_pe_1_2_6_U110 ( .A(npu_inst_pe_1_2_6_n53), .ZN(
        npu_inst_pe_1_2_6_n109) );
  AOI22_X1 npu_inst_pe_1_2_6_U107 ( .A1(npu_inst_int_data_y_3__6__0_), .A2(
        npu_inst_pe_1_2_6_n50), .B1(npu_inst_pe_1_2_6_n117), .B2(
        npu_inst_pe_1_2_6_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_2_6_n49) );
  INV_X1 npu_inst_pe_1_2_6_U106 ( .A(npu_inst_pe_1_2_6_n49), .ZN(
        npu_inst_pe_1_2_6_n110) );
  AOI22_X1 npu_inst_pe_1_2_6_U105 ( .A1(npu_inst_int_data_y_3__6__0_), .A2(
        npu_inst_pe_1_2_6_n46), .B1(npu_inst_pe_1_2_6_n116), .B2(
        npu_inst_pe_1_2_6_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_2_6_n45) );
  INV_X1 npu_inst_pe_1_2_6_U104 ( .A(npu_inst_pe_1_2_6_n45), .ZN(
        npu_inst_pe_1_2_6_n111) );
  AOI22_X1 npu_inst_pe_1_2_6_U103 ( .A1(npu_inst_int_data_y_3__6__0_), .A2(
        npu_inst_pe_1_2_6_n42), .B1(npu_inst_pe_1_2_6_n115), .B2(
        npu_inst_pe_1_2_6_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_2_6_n41) );
  INV_X1 npu_inst_pe_1_2_6_U102 ( .A(npu_inst_pe_1_2_6_n41), .ZN(
        npu_inst_pe_1_2_6_n112) );
  AOI22_X1 npu_inst_pe_1_2_6_U101 ( .A1(npu_inst_int_data_y_3__6__1_), .A2(
        npu_inst_pe_1_2_6_n58), .B1(npu_inst_pe_1_2_6_n119), .B2(
        npu_inst_pe_1_2_6_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_2_6_n59) );
  INV_X1 npu_inst_pe_1_2_6_U100 ( .A(npu_inst_pe_1_2_6_n59), .ZN(
        npu_inst_pe_1_2_6_n102) );
  AOI22_X1 npu_inst_pe_1_2_6_U99 ( .A1(npu_inst_int_data_y_3__6__1_), .A2(
        npu_inst_pe_1_2_6_n54), .B1(npu_inst_pe_1_2_6_n118), .B2(
        npu_inst_pe_1_2_6_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_2_6_n55) );
  INV_X1 npu_inst_pe_1_2_6_U98 ( .A(npu_inst_pe_1_2_6_n55), .ZN(
        npu_inst_pe_1_2_6_n103) );
  AOI22_X1 npu_inst_pe_1_2_6_U97 ( .A1(npu_inst_int_data_y_3__6__1_), .A2(
        npu_inst_pe_1_2_6_n50), .B1(npu_inst_pe_1_2_6_n117), .B2(
        npu_inst_pe_1_2_6_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_2_6_n51) );
  INV_X1 npu_inst_pe_1_2_6_U96 ( .A(npu_inst_pe_1_2_6_n51), .ZN(
        npu_inst_pe_1_2_6_n104) );
  AOI22_X1 npu_inst_pe_1_2_6_U95 ( .A1(npu_inst_int_data_y_3__6__1_), .A2(
        npu_inst_pe_1_2_6_n46), .B1(npu_inst_pe_1_2_6_n116), .B2(
        npu_inst_pe_1_2_6_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_2_6_n47) );
  INV_X1 npu_inst_pe_1_2_6_U94 ( .A(npu_inst_pe_1_2_6_n47), .ZN(
        npu_inst_pe_1_2_6_n105) );
  AOI22_X1 npu_inst_pe_1_2_6_U93 ( .A1(npu_inst_int_data_y_3__6__1_), .A2(
        npu_inst_pe_1_2_6_n42), .B1(npu_inst_pe_1_2_6_n115), .B2(
        npu_inst_pe_1_2_6_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_2_6_n43) );
  INV_X1 npu_inst_pe_1_2_6_U92 ( .A(npu_inst_pe_1_2_6_n43), .ZN(
        npu_inst_pe_1_2_6_n106) );
  AOI22_X1 npu_inst_pe_1_2_6_U91 ( .A1(npu_inst_pe_1_2_6_n38), .A2(
        npu_inst_int_data_y_3__6__1_), .B1(npu_inst_pe_1_2_6_n114), .B2(
        npu_inst_pe_1_2_6_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_2_6_n39) );
  INV_X1 npu_inst_pe_1_2_6_U90 ( .A(npu_inst_pe_1_2_6_n39), .ZN(
        npu_inst_pe_1_2_6_n107) );
  AOI22_X1 npu_inst_pe_1_2_6_U89 ( .A1(npu_inst_pe_1_2_6_n38), .A2(
        npu_inst_int_data_y_3__6__0_), .B1(npu_inst_pe_1_2_6_n114), .B2(
        npu_inst_pe_1_2_6_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_2_6_n37) );
  INV_X1 npu_inst_pe_1_2_6_U88 ( .A(npu_inst_pe_1_2_6_n37), .ZN(
        npu_inst_pe_1_2_6_n113) );
  NAND2_X1 npu_inst_pe_1_2_6_U87 ( .A1(npu_inst_pe_1_2_6_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_2_6_n60), .ZN(npu_inst_pe_1_2_6_n74) );
  OAI21_X1 npu_inst_pe_1_2_6_U86 ( .B1(npu_inst_pe_1_2_6_n63), .B2(
        npu_inst_pe_1_2_6_n60), .A(npu_inst_pe_1_2_6_n74), .ZN(
        npu_inst_pe_1_2_6_n97) );
  NAND2_X1 npu_inst_pe_1_2_6_U85 ( .A1(npu_inst_pe_1_2_6_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_2_6_n60), .ZN(npu_inst_pe_1_2_6_n73) );
  OAI21_X1 npu_inst_pe_1_2_6_U84 ( .B1(npu_inst_pe_1_2_6_n61), .B2(
        npu_inst_pe_1_2_6_n60), .A(npu_inst_pe_1_2_6_n73), .ZN(
        npu_inst_pe_1_2_6_n96) );
  NAND2_X1 npu_inst_pe_1_2_6_U83 ( .A1(npu_inst_pe_1_2_6_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_2_6_n56), .ZN(npu_inst_pe_1_2_6_n72) );
  OAI21_X1 npu_inst_pe_1_2_6_U82 ( .B1(npu_inst_pe_1_2_6_n63), .B2(
        npu_inst_pe_1_2_6_n56), .A(npu_inst_pe_1_2_6_n72), .ZN(
        npu_inst_pe_1_2_6_n95) );
  NAND2_X1 npu_inst_pe_1_2_6_U81 ( .A1(npu_inst_pe_1_2_6_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_2_6_n56), .ZN(npu_inst_pe_1_2_6_n71) );
  OAI21_X1 npu_inst_pe_1_2_6_U80 ( .B1(npu_inst_pe_1_2_6_n61), .B2(
        npu_inst_pe_1_2_6_n56), .A(npu_inst_pe_1_2_6_n71), .ZN(
        npu_inst_pe_1_2_6_n94) );
  NAND2_X1 npu_inst_pe_1_2_6_U79 ( .A1(npu_inst_pe_1_2_6_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_2_6_n52), .ZN(npu_inst_pe_1_2_6_n70) );
  OAI21_X1 npu_inst_pe_1_2_6_U78 ( .B1(npu_inst_pe_1_2_6_n63), .B2(
        npu_inst_pe_1_2_6_n52), .A(npu_inst_pe_1_2_6_n70), .ZN(
        npu_inst_pe_1_2_6_n93) );
  NAND2_X1 npu_inst_pe_1_2_6_U77 ( .A1(npu_inst_pe_1_2_6_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_2_6_n52), .ZN(npu_inst_pe_1_2_6_n69) );
  OAI21_X1 npu_inst_pe_1_2_6_U76 ( .B1(npu_inst_pe_1_2_6_n61), .B2(
        npu_inst_pe_1_2_6_n52), .A(npu_inst_pe_1_2_6_n69), .ZN(
        npu_inst_pe_1_2_6_n92) );
  NAND2_X1 npu_inst_pe_1_2_6_U75 ( .A1(npu_inst_pe_1_2_6_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_2_6_n48), .ZN(npu_inst_pe_1_2_6_n68) );
  OAI21_X1 npu_inst_pe_1_2_6_U74 ( .B1(npu_inst_pe_1_2_6_n63), .B2(
        npu_inst_pe_1_2_6_n48), .A(npu_inst_pe_1_2_6_n68), .ZN(
        npu_inst_pe_1_2_6_n91) );
  NAND2_X1 npu_inst_pe_1_2_6_U73 ( .A1(npu_inst_pe_1_2_6_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_2_6_n48), .ZN(npu_inst_pe_1_2_6_n67) );
  OAI21_X1 npu_inst_pe_1_2_6_U72 ( .B1(npu_inst_pe_1_2_6_n61), .B2(
        npu_inst_pe_1_2_6_n48), .A(npu_inst_pe_1_2_6_n67), .ZN(
        npu_inst_pe_1_2_6_n90) );
  NAND2_X1 npu_inst_pe_1_2_6_U71 ( .A1(npu_inst_pe_1_2_6_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_2_6_n44), .ZN(npu_inst_pe_1_2_6_n66) );
  OAI21_X1 npu_inst_pe_1_2_6_U70 ( .B1(npu_inst_pe_1_2_6_n63), .B2(
        npu_inst_pe_1_2_6_n44), .A(npu_inst_pe_1_2_6_n66), .ZN(
        npu_inst_pe_1_2_6_n89) );
  NAND2_X1 npu_inst_pe_1_2_6_U69 ( .A1(npu_inst_pe_1_2_6_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_2_6_n44), .ZN(npu_inst_pe_1_2_6_n65) );
  OAI21_X1 npu_inst_pe_1_2_6_U68 ( .B1(npu_inst_pe_1_2_6_n61), .B2(
        npu_inst_pe_1_2_6_n44), .A(npu_inst_pe_1_2_6_n65), .ZN(
        npu_inst_pe_1_2_6_n88) );
  NAND2_X1 npu_inst_pe_1_2_6_U67 ( .A1(npu_inst_pe_1_2_6_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_2_6_n40), .ZN(npu_inst_pe_1_2_6_n64) );
  OAI21_X1 npu_inst_pe_1_2_6_U66 ( .B1(npu_inst_pe_1_2_6_n63), .B2(
        npu_inst_pe_1_2_6_n40), .A(npu_inst_pe_1_2_6_n64), .ZN(
        npu_inst_pe_1_2_6_n87) );
  NAND2_X1 npu_inst_pe_1_2_6_U65 ( .A1(npu_inst_pe_1_2_6_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_2_6_n40), .ZN(npu_inst_pe_1_2_6_n62) );
  OAI21_X1 npu_inst_pe_1_2_6_U64 ( .B1(npu_inst_pe_1_2_6_n61), .B2(
        npu_inst_pe_1_2_6_n40), .A(npu_inst_pe_1_2_6_n62), .ZN(
        npu_inst_pe_1_2_6_n86) );
  AND2_X1 npu_inst_pe_1_2_6_U63 ( .A1(npu_inst_pe_1_2_6_N93), .A2(npu_inst_n57), .ZN(npu_inst_int_data_y_2__6__0_) );
  AND2_X1 npu_inst_pe_1_2_6_U62 ( .A1(npu_inst_n57), .A2(npu_inst_pe_1_2_6_N94), .ZN(npu_inst_int_data_y_2__6__1_) );
  NOR3_X1 npu_inst_pe_1_2_6_U61 ( .A1(npu_inst_pe_1_2_6_n26), .A2(npu_inst_n57), .A3(npu_inst_int_ckg[41]), .ZN(npu_inst_pe_1_2_6_n85) );
  OR2_X1 npu_inst_pe_1_2_6_U60 ( .A1(npu_inst_pe_1_2_6_n85), .A2(
        npu_inst_pe_1_2_6_n2), .ZN(npu_inst_pe_1_2_6_N84) );
  AND2_X1 npu_inst_pe_1_2_6_U59 ( .A1(npu_inst_pe_1_2_6_int_q_acc_0_), .A2(
        npu_inst_pe_1_2_6_n1), .ZN(npu_inst_int_data_res_2__6__0_) );
  AND2_X1 npu_inst_pe_1_2_6_U58 ( .A1(npu_inst_pe_1_2_6_n2), .A2(
        npu_inst_pe_1_2_6_int_q_acc_7_), .ZN(npu_inst_int_data_res_2__6__7_)
         );
  AND2_X1 npu_inst_pe_1_2_6_U57 ( .A1(npu_inst_pe_1_2_6_int_q_acc_1_), .A2(
        npu_inst_pe_1_2_6_n1), .ZN(npu_inst_int_data_res_2__6__1_) );
  AND2_X1 npu_inst_pe_1_2_6_U56 ( .A1(npu_inst_pe_1_2_6_int_q_acc_2_), .A2(
        npu_inst_pe_1_2_6_n1), .ZN(npu_inst_int_data_res_2__6__2_) );
  AND2_X1 npu_inst_pe_1_2_6_U55 ( .A1(npu_inst_pe_1_2_6_int_q_acc_3_), .A2(
        npu_inst_pe_1_2_6_n2), .ZN(npu_inst_int_data_res_2__6__3_) );
  AND2_X1 npu_inst_pe_1_2_6_U54 ( .A1(npu_inst_pe_1_2_6_int_q_acc_4_), .A2(
        npu_inst_pe_1_2_6_n2), .ZN(npu_inst_int_data_res_2__6__4_) );
  AND2_X1 npu_inst_pe_1_2_6_U53 ( .A1(npu_inst_pe_1_2_6_int_q_acc_5_), .A2(
        npu_inst_pe_1_2_6_n2), .ZN(npu_inst_int_data_res_2__6__5_) );
  AND2_X1 npu_inst_pe_1_2_6_U52 ( .A1(npu_inst_pe_1_2_6_int_q_acc_6_), .A2(
        npu_inst_pe_1_2_6_n2), .ZN(npu_inst_int_data_res_2__6__6_) );
  AOI222_X1 npu_inst_pe_1_2_6_U51 ( .A1(npu_inst_int_data_res_3__6__0_), .A2(
        npu_inst_pe_1_2_6_n1), .B1(npu_inst_pe_1_2_6_N73), .B2(
        npu_inst_pe_1_2_6_n76), .C1(npu_inst_pe_1_2_6_N65), .C2(
        npu_inst_pe_1_2_6_n77), .ZN(npu_inst_pe_1_2_6_n84) );
  INV_X1 npu_inst_pe_1_2_6_U50 ( .A(npu_inst_pe_1_2_6_n84), .ZN(
        npu_inst_pe_1_2_6_n101) );
  AOI222_X1 npu_inst_pe_1_2_6_U49 ( .A1(npu_inst_int_data_res_3__6__7_), .A2(
        npu_inst_pe_1_2_6_n1), .B1(npu_inst_pe_1_2_6_N80), .B2(
        npu_inst_pe_1_2_6_n76), .C1(npu_inst_pe_1_2_6_N72), .C2(
        npu_inst_pe_1_2_6_n77), .ZN(npu_inst_pe_1_2_6_n75) );
  INV_X1 npu_inst_pe_1_2_6_U48 ( .A(npu_inst_pe_1_2_6_n75), .ZN(
        npu_inst_pe_1_2_6_n33) );
  AOI222_X1 npu_inst_pe_1_2_6_U47 ( .A1(npu_inst_int_data_res_3__6__1_), .A2(
        npu_inst_pe_1_2_6_n1), .B1(npu_inst_pe_1_2_6_N74), .B2(
        npu_inst_pe_1_2_6_n76), .C1(npu_inst_pe_1_2_6_N66), .C2(
        npu_inst_pe_1_2_6_n77), .ZN(npu_inst_pe_1_2_6_n83) );
  INV_X1 npu_inst_pe_1_2_6_U46 ( .A(npu_inst_pe_1_2_6_n83), .ZN(
        npu_inst_pe_1_2_6_n100) );
  AOI222_X1 npu_inst_pe_1_2_6_U45 ( .A1(npu_inst_int_data_res_3__6__2_), .A2(
        npu_inst_pe_1_2_6_n1), .B1(npu_inst_pe_1_2_6_N75), .B2(
        npu_inst_pe_1_2_6_n76), .C1(npu_inst_pe_1_2_6_N67), .C2(
        npu_inst_pe_1_2_6_n77), .ZN(npu_inst_pe_1_2_6_n82) );
  INV_X1 npu_inst_pe_1_2_6_U44 ( .A(npu_inst_pe_1_2_6_n82), .ZN(
        npu_inst_pe_1_2_6_n99) );
  AOI222_X1 npu_inst_pe_1_2_6_U43 ( .A1(npu_inst_int_data_res_3__6__3_), .A2(
        npu_inst_pe_1_2_6_n1), .B1(npu_inst_pe_1_2_6_N76), .B2(
        npu_inst_pe_1_2_6_n76), .C1(npu_inst_pe_1_2_6_N68), .C2(
        npu_inst_pe_1_2_6_n77), .ZN(npu_inst_pe_1_2_6_n81) );
  INV_X1 npu_inst_pe_1_2_6_U42 ( .A(npu_inst_pe_1_2_6_n81), .ZN(
        npu_inst_pe_1_2_6_n98) );
  AOI222_X1 npu_inst_pe_1_2_6_U41 ( .A1(npu_inst_int_data_res_3__6__4_), .A2(
        npu_inst_pe_1_2_6_n1), .B1(npu_inst_pe_1_2_6_N77), .B2(
        npu_inst_pe_1_2_6_n76), .C1(npu_inst_pe_1_2_6_N69), .C2(
        npu_inst_pe_1_2_6_n77), .ZN(npu_inst_pe_1_2_6_n80) );
  INV_X1 npu_inst_pe_1_2_6_U40 ( .A(npu_inst_pe_1_2_6_n80), .ZN(
        npu_inst_pe_1_2_6_n36) );
  AOI222_X1 npu_inst_pe_1_2_6_U39 ( .A1(npu_inst_int_data_res_3__6__5_), .A2(
        npu_inst_pe_1_2_6_n1), .B1(npu_inst_pe_1_2_6_N78), .B2(
        npu_inst_pe_1_2_6_n76), .C1(npu_inst_pe_1_2_6_N70), .C2(
        npu_inst_pe_1_2_6_n77), .ZN(npu_inst_pe_1_2_6_n79) );
  INV_X1 npu_inst_pe_1_2_6_U38 ( .A(npu_inst_pe_1_2_6_n79), .ZN(
        npu_inst_pe_1_2_6_n35) );
  AOI222_X1 npu_inst_pe_1_2_6_U37 ( .A1(npu_inst_int_data_res_3__6__6_), .A2(
        npu_inst_pe_1_2_6_n1), .B1(npu_inst_pe_1_2_6_N79), .B2(
        npu_inst_pe_1_2_6_n76), .C1(npu_inst_pe_1_2_6_N71), .C2(
        npu_inst_pe_1_2_6_n77), .ZN(npu_inst_pe_1_2_6_n78) );
  INV_X1 npu_inst_pe_1_2_6_U36 ( .A(npu_inst_pe_1_2_6_n78), .ZN(
        npu_inst_pe_1_2_6_n34) );
  INV_X1 npu_inst_pe_1_2_6_U35 ( .A(npu_inst_pe_1_2_6_int_data_1_), .ZN(
        npu_inst_pe_1_2_6_n14) );
  AND2_X1 npu_inst_pe_1_2_6_U34 ( .A1(npu_inst_int_data_x_2__6__1_), .A2(
        npu_inst_pe_1_2_6_int_q_weight_1_), .ZN(npu_inst_pe_1_2_6_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_2_6_U33 ( .A1(npu_inst_int_data_x_2__6__0_), .A2(
        npu_inst_pe_1_2_6_int_q_weight_1_), .ZN(npu_inst_pe_1_2_6_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_2_6_U32 ( .A1(npu_inst_n57), .A2(
        npu_inst_int_data_y_3__6__1_), .B1(npu_inst_pe_1_2_6_n3), .B2(
        npu_inst_int_data_x_2__7__1_), .ZN(npu_inst_pe_1_2_6_n63) );
  AOI22_X1 npu_inst_pe_1_2_6_U31 ( .A1(npu_inst_n57), .A2(
        npu_inst_int_data_y_3__6__0_), .B1(npu_inst_pe_1_2_6_n3), .B2(
        npu_inst_int_data_x_2__7__0_), .ZN(npu_inst_pe_1_2_6_n61) );
  INV_X1 npu_inst_pe_1_2_6_U30 ( .A(npu_inst_pe_1_2_6_int_data_0_), .ZN(
        npu_inst_pe_1_2_6_n13) );
  INV_X1 npu_inst_pe_1_2_6_U29 ( .A(npu_inst_n70), .ZN(npu_inst_pe_1_2_6_n5)
         );
  OR3_X1 npu_inst_pe_1_2_6_U28 ( .A1(npu_inst_pe_1_2_6_n6), .A2(
        npu_inst_pe_1_2_6_n8), .A3(npu_inst_pe_1_2_6_n5), .ZN(
        npu_inst_pe_1_2_6_n56) );
  OR3_X1 npu_inst_pe_1_2_6_U27 ( .A1(npu_inst_pe_1_2_6_n5), .A2(
        npu_inst_pe_1_2_6_n8), .A3(npu_inst_pe_1_2_6_n7), .ZN(
        npu_inst_pe_1_2_6_n48) );
  INV_X1 npu_inst_pe_1_2_6_U26 ( .A(npu_inst_pe_1_2_6_n5), .ZN(
        npu_inst_pe_1_2_6_n4) );
  OR3_X1 npu_inst_pe_1_2_6_U25 ( .A1(npu_inst_pe_1_2_6_n4), .A2(
        npu_inst_pe_1_2_6_n8), .A3(npu_inst_pe_1_2_6_n7), .ZN(
        npu_inst_pe_1_2_6_n52) );
  OR3_X1 npu_inst_pe_1_2_6_U24 ( .A1(npu_inst_pe_1_2_6_n6), .A2(
        npu_inst_pe_1_2_6_n8), .A3(npu_inst_pe_1_2_6_n4), .ZN(
        npu_inst_pe_1_2_6_n60) );
  NOR2_X1 npu_inst_pe_1_2_6_U23 ( .A1(npu_inst_pe_1_2_6_n60), .A2(
        npu_inst_pe_1_2_6_n3), .ZN(npu_inst_pe_1_2_6_n58) );
  NOR2_X1 npu_inst_pe_1_2_6_U22 ( .A1(npu_inst_pe_1_2_6_n56), .A2(
        npu_inst_pe_1_2_6_n3), .ZN(npu_inst_pe_1_2_6_n54) );
  NOR2_X1 npu_inst_pe_1_2_6_U21 ( .A1(npu_inst_pe_1_2_6_n52), .A2(
        npu_inst_pe_1_2_6_n3), .ZN(npu_inst_pe_1_2_6_n50) );
  NOR2_X1 npu_inst_pe_1_2_6_U20 ( .A1(npu_inst_pe_1_2_6_n48), .A2(
        npu_inst_pe_1_2_6_n3), .ZN(npu_inst_pe_1_2_6_n46) );
  NOR2_X1 npu_inst_pe_1_2_6_U19 ( .A1(npu_inst_pe_1_2_6_n40), .A2(
        npu_inst_pe_1_2_6_n3), .ZN(npu_inst_pe_1_2_6_n38) );
  NOR2_X1 npu_inst_pe_1_2_6_U18 ( .A1(npu_inst_pe_1_2_6_n44), .A2(
        npu_inst_pe_1_2_6_n3), .ZN(npu_inst_pe_1_2_6_n42) );
  BUF_X1 npu_inst_pe_1_2_6_U17 ( .A(npu_inst_n102), .Z(npu_inst_pe_1_2_6_n8)
         );
  INV_X1 npu_inst_pe_1_2_6_U16 ( .A(npu_inst_n125), .ZN(npu_inst_pe_1_2_6_n12)
         );
  INV_X1 npu_inst_pe_1_2_6_U15 ( .A(npu_inst_pe_1_2_6_n38), .ZN(
        npu_inst_pe_1_2_6_n114) );
  INV_X1 npu_inst_pe_1_2_6_U14 ( .A(npu_inst_pe_1_2_6_n58), .ZN(
        npu_inst_pe_1_2_6_n119) );
  INV_X1 npu_inst_pe_1_2_6_U13 ( .A(npu_inst_pe_1_2_6_n54), .ZN(
        npu_inst_pe_1_2_6_n118) );
  INV_X1 npu_inst_pe_1_2_6_U12 ( .A(npu_inst_pe_1_2_6_n50), .ZN(
        npu_inst_pe_1_2_6_n117) );
  INV_X1 npu_inst_pe_1_2_6_U11 ( .A(npu_inst_pe_1_2_6_n46), .ZN(
        npu_inst_pe_1_2_6_n116) );
  INV_X1 npu_inst_pe_1_2_6_U10 ( .A(npu_inst_pe_1_2_6_n42), .ZN(
        npu_inst_pe_1_2_6_n115) );
  BUF_X1 npu_inst_pe_1_2_6_U9 ( .A(npu_inst_n27), .Z(npu_inst_pe_1_2_6_n2) );
  BUF_X1 npu_inst_pe_1_2_6_U8 ( .A(npu_inst_n27), .Z(npu_inst_pe_1_2_6_n1) );
  BUF_X1 npu_inst_pe_1_2_6_U7 ( .A(npu_inst_pe_1_2_6_n12), .Z(
        npu_inst_pe_1_2_6_n11) );
  BUF_X1 npu_inst_pe_1_2_6_U6 ( .A(npu_inst_pe_1_2_6_n12), .Z(
        npu_inst_pe_1_2_6_n10) );
  BUF_X1 npu_inst_pe_1_2_6_U5 ( .A(npu_inst_pe_1_2_6_n12), .Z(
        npu_inst_pe_1_2_6_n9) );
  NOR2_X1 npu_inst_pe_1_2_6_U4 ( .A1(npu_inst_pe_1_2_6_int_q_weight_0_), .A2(
        npu_inst_pe_1_2_6_n1), .ZN(npu_inst_pe_1_2_6_n76) );
  NOR2_X1 npu_inst_pe_1_2_6_U3 ( .A1(npu_inst_pe_1_2_6_n27), .A2(
        npu_inst_pe_1_2_6_n1), .ZN(npu_inst_pe_1_2_6_n77) );
  FA_X1 npu_inst_pe_1_2_6_sub_67_U2_1 ( .A(npu_inst_pe_1_2_6_int_q_acc_1_), 
        .B(npu_inst_pe_1_2_6_n14), .CI(npu_inst_pe_1_2_6_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_2_6_sub_67_carry_2_), .S(npu_inst_pe_1_2_6_N66) );
  FA_X1 npu_inst_pe_1_2_6_add_69_U1_1 ( .A(npu_inst_pe_1_2_6_int_q_acc_1_), 
        .B(npu_inst_pe_1_2_6_int_data_1_), .CI(
        npu_inst_pe_1_2_6_add_69_carry_1_), .CO(
        npu_inst_pe_1_2_6_add_69_carry_2_), .S(npu_inst_pe_1_2_6_N74) );
  NAND3_X1 npu_inst_pe_1_2_6_U109 ( .A1(npu_inst_pe_1_2_6_n5), .A2(
        npu_inst_pe_1_2_6_n7), .A3(npu_inst_pe_1_2_6_n8), .ZN(
        npu_inst_pe_1_2_6_n44) );
  NAND3_X1 npu_inst_pe_1_2_6_U108 ( .A1(npu_inst_pe_1_2_6_n4), .A2(
        npu_inst_pe_1_2_6_n7), .A3(npu_inst_pe_1_2_6_n8), .ZN(
        npu_inst_pe_1_2_6_n40) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_2_6_n34), .CK(
        npu_inst_pe_1_2_6_net4056), .RN(npu_inst_pe_1_2_6_n9), .Q(
        npu_inst_pe_1_2_6_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_2_6_n35), .CK(
        npu_inst_pe_1_2_6_net4056), .RN(npu_inst_pe_1_2_6_n9), .Q(
        npu_inst_pe_1_2_6_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_2_6_n36), .CK(
        npu_inst_pe_1_2_6_net4056), .RN(npu_inst_pe_1_2_6_n9), .Q(
        npu_inst_pe_1_2_6_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_2_6_n98), .CK(
        npu_inst_pe_1_2_6_net4056), .RN(npu_inst_pe_1_2_6_n9), .Q(
        npu_inst_pe_1_2_6_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_2_6_n99), .CK(
        npu_inst_pe_1_2_6_net4056), .RN(npu_inst_pe_1_2_6_n9), .Q(
        npu_inst_pe_1_2_6_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_2_6_n100), 
        .CK(npu_inst_pe_1_2_6_net4056), .RN(npu_inst_pe_1_2_6_n9), .Q(
        npu_inst_pe_1_2_6_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_2_6_n33), .CK(
        npu_inst_pe_1_2_6_net4056), .RN(npu_inst_pe_1_2_6_n9), .Q(
        npu_inst_pe_1_2_6_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_2_6_n101), 
        .CK(npu_inst_pe_1_2_6_net4056), .RN(npu_inst_pe_1_2_6_n9), .Q(
        npu_inst_pe_1_2_6_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_weight_reg_0_ ( .D(npu_inst_n111), .CK(
        npu_inst_pe_1_2_6_net4062), .RN(npu_inst_pe_1_2_6_n9), .Q(
        npu_inst_pe_1_2_6_int_q_weight_0_), .QN(npu_inst_pe_1_2_6_n27) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_weight_reg_1_ ( .D(npu_inst_n117), .CK(
        npu_inst_pe_1_2_6_net4062), .RN(npu_inst_pe_1_2_6_n9), .Q(
        npu_inst_pe_1_2_6_int_q_weight_1_), .QN(npu_inst_pe_1_2_6_n26) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_2_6_n113), 
        .CK(npu_inst_pe_1_2_6_net4062), .RN(npu_inst_pe_1_2_6_n9), .Q(
        npu_inst_pe_1_2_6_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_2_6_n107), 
        .CK(npu_inst_pe_1_2_6_net4062), .RN(npu_inst_pe_1_2_6_n9), .Q(
        npu_inst_pe_1_2_6_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_2_6_n112), 
        .CK(npu_inst_pe_1_2_6_net4062), .RN(npu_inst_pe_1_2_6_n10), .Q(
        npu_inst_pe_1_2_6_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_2_6_n106), 
        .CK(npu_inst_pe_1_2_6_net4062), .RN(npu_inst_pe_1_2_6_n10), .Q(
        npu_inst_pe_1_2_6_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_2_6_n111), 
        .CK(npu_inst_pe_1_2_6_net4062), .RN(npu_inst_pe_1_2_6_n10), .Q(
        npu_inst_pe_1_2_6_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_2_6_n105), 
        .CK(npu_inst_pe_1_2_6_net4062), .RN(npu_inst_pe_1_2_6_n10), .Q(
        npu_inst_pe_1_2_6_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_2_6_n110), 
        .CK(npu_inst_pe_1_2_6_net4062), .RN(npu_inst_pe_1_2_6_n10), .Q(
        npu_inst_pe_1_2_6_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_2_6_n104), 
        .CK(npu_inst_pe_1_2_6_net4062), .RN(npu_inst_pe_1_2_6_n10), .Q(
        npu_inst_pe_1_2_6_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_2_6_n109), 
        .CK(npu_inst_pe_1_2_6_net4062), .RN(npu_inst_pe_1_2_6_n10), .Q(
        npu_inst_pe_1_2_6_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_2_6_n103), 
        .CK(npu_inst_pe_1_2_6_net4062), .RN(npu_inst_pe_1_2_6_n10), .Q(
        npu_inst_pe_1_2_6_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_2_6_n108), 
        .CK(npu_inst_pe_1_2_6_net4062), .RN(npu_inst_pe_1_2_6_n10), .Q(
        npu_inst_pe_1_2_6_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_2_6_n102), 
        .CK(npu_inst_pe_1_2_6_net4062), .RN(npu_inst_pe_1_2_6_n10), .Q(
        npu_inst_pe_1_2_6_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_2_6_n86), 
        .CK(npu_inst_pe_1_2_6_net4062), .RN(npu_inst_pe_1_2_6_n10), .Q(
        npu_inst_pe_1_2_6_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_2_6_n87), 
        .CK(npu_inst_pe_1_2_6_net4062), .RN(npu_inst_pe_1_2_6_n10), .Q(
        npu_inst_pe_1_2_6_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_2_6_n88), 
        .CK(npu_inst_pe_1_2_6_net4062), .RN(npu_inst_pe_1_2_6_n11), .Q(
        npu_inst_pe_1_2_6_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_2_6_n89), 
        .CK(npu_inst_pe_1_2_6_net4062), .RN(npu_inst_pe_1_2_6_n11), .Q(
        npu_inst_pe_1_2_6_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_2_6_n90), 
        .CK(npu_inst_pe_1_2_6_net4062), .RN(npu_inst_pe_1_2_6_n11), .Q(
        npu_inst_pe_1_2_6_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_2_6_n91), 
        .CK(npu_inst_pe_1_2_6_net4062), .RN(npu_inst_pe_1_2_6_n11), .Q(
        npu_inst_pe_1_2_6_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_2_6_n92), 
        .CK(npu_inst_pe_1_2_6_net4062), .RN(npu_inst_pe_1_2_6_n11), .Q(
        npu_inst_pe_1_2_6_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_2_6_n93), 
        .CK(npu_inst_pe_1_2_6_net4062), .RN(npu_inst_pe_1_2_6_n11), .Q(
        npu_inst_pe_1_2_6_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_2_6_n94), 
        .CK(npu_inst_pe_1_2_6_net4062), .RN(npu_inst_pe_1_2_6_n11), .Q(
        npu_inst_pe_1_2_6_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_2_6_n95), 
        .CK(npu_inst_pe_1_2_6_net4062), .RN(npu_inst_pe_1_2_6_n11), .Q(
        npu_inst_pe_1_2_6_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_2_6_n96), 
        .CK(npu_inst_pe_1_2_6_net4062), .RN(npu_inst_pe_1_2_6_n11), .Q(
        npu_inst_pe_1_2_6_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_2_6_n97), 
        .CK(npu_inst_pe_1_2_6_net4062), .RN(npu_inst_pe_1_2_6_n11), .Q(
        npu_inst_pe_1_2_6_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_2_6_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_2_6_N84), .SE(1'b0), .GCK(npu_inst_pe_1_2_6_net4056) );
  CLKGATETST_X1 npu_inst_pe_1_2_6_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n64), .SE(1'b0), .GCK(npu_inst_pe_1_2_6_net4062) );
  MUX2_X1 npu_inst_pe_1_2_7_U162 ( .A(npu_inst_pe_1_2_7_n32), .B(
        npu_inst_pe_1_2_7_n29), .S(npu_inst_pe_1_2_7_n8), .Z(
        npu_inst_pe_1_2_7_N93) );
  MUX2_X1 npu_inst_pe_1_2_7_U161 ( .A(npu_inst_pe_1_2_7_n31), .B(
        npu_inst_pe_1_2_7_n30), .S(npu_inst_pe_1_2_7_n6), .Z(
        npu_inst_pe_1_2_7_n32) );
  MUX2_X1 npu_inst_pe_1_2_7_U160 ( .A(npu_inst_pe_1_2_7_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_2_7_int_q_reg_v_1__0_), .S(npu_inst_pe_1_2_7_n4), .Z(
        npu_inst_pe_1_2_7_n31) );
  MUX2_X1 npu_inst_pe_1_2_7_U159 ( .A(npu_inst_pe_1_2_7_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_2_7_int_q_reg_v_3__0_), .S(npu_inst_pe_1_2_7_n4), .Z(
        npu_inst_pe_1_2_7_n30) );
  MUX2_X1 npu_inst_pe_1_2_7_U158 ( .A(npu_inst_pe_1_2_7_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_2_7_int_q_reg_v_5__0_), .S(npu_inst_pe_1_2_7_n4), .Z(
        npu_inst_pe_1_2_7_n29) );
  MUX2_X1 npu_inst_pe_1_2_7_U157 ( .A(npu_inst_pe_1_2_7_n28), .B(
        npu_inst_pe_1_2_7_n23), .S(npu_inst_pe_1_2_7_n8), .Z(
        npu_inst_pe_1_2_7_N94) );
  MUX2_X1 npu_inst_pe_1_2_7_U156 ( .A(npu_inst_pe_1_2_7_n25), .B(
        npu_inst_pe_1_2_7_n24), .S(npu_inst_pe_1_2_7_n6), .Z(
        npu_inst_pe_1_2_7_n28) );
  MUX2_X1 npu_inst_pe_1_2_7_U155 ( .A(npu_inst_pe_1_2_7_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_2_7_int_q_reg_v_1__1_), .S(npu_inst_pe_1_2_7_n4), .Z(
        npu_inst_pe_1_2_7_n25) );
  MUX2_X1 npu_inst_pe_1_2_7_U154 ( .A(npu_inst_pe_1_2_7_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_2_7_int_q_reg_v_3__1_), .S(npu_inst_pe_1_2_7_n4), .Z(
        npu_inst_pe_1_2_7_n24) );
  MUX2_X1 npu_inst_pe_1_2_7_U153 ( .A(npu_inst_pe_1_2_7_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_2_7_int_q_reg_v_5__1_), .S(npu_inst_pe_1_2_7_n4), .Z(
        npu_inst_pe_1_2_7_n23) );
  MUX2_X1 npu_inst_pe_1_2_7_U152 ( .A(npu_inst_pe_1_2_7_n22), .B(
        npu_inst_pe_1_2_7_n19), .S(npu_inst_pe_1_2_7_n8), .Z(
        npu_inst_int_data_x_2__7__1_) );
  MUX2_X1 npu_inst_pe_1_2_7_U151 ( .A(npu_inst_pe_1_2_7_n21), .B(
        npu_inst_pe_1_2_7_n20), .S(npu_inst_pe_1_2_7_n6), .Z(
        npu_inst_pe_1_2_7_n22) );
  MUX2_X1 npu_inst_pe_1_2_7_U150 ( .A(npu_inst_pe_1_2_7_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_2_7_int_q_reg_h_1__1_), .S(npu_inst_pe_1_2_7_n4), .Z(
        npu_inst_pe_1_2_7_n21) );
  MUX2_X1 npu_inst_pe_1_2_7_U149 ( .A(npu_inst_pe_1_2_7_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_2_7_int_q_reg_h_3__1_), .S(npu_inst_pe_1_2_7_n4), .Z(
        npu_inst_pe_1_2_7_n20) );
  MUX2_X1 npu_inst_pe_1_2_7_U148 ( .A(npu_inst_pe_1_2_7_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_2_7_int_q_reg_h_5__1_), .S(npu_inst_pe_1_2_7_n4), .Z(
        npu_inst_pe_1_2_7_n19) );
  MUX2_X1 npu_inst_pe_1_2_7_U147 ( .A(npu_inst_pe_1_2_7_n18), .B(
        npu_inst_pe_1_2_7_n15), .S(npu_inst_pe_1_2_7_n8), .Z(
        npu_inst_int_data_x_2__7__0_) );
  MUX2_X1 npu_inst_pe_1_2_7_U146 ( .A(npu_inst_pe_1_2_7_n17), .B(
        npu_inst_pe_1_2_7_n16), .S(npu_inst_pe_1_2_7_n6), .Z(
        npu_inst_pe_1_2_7_n18) );
  MUX2_X1 npu_inst_pe_1_2_7_U145 ( .A(npu_inst_pe_1_2_7_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_2_7_int_q_reg_h_1__0_), .S(npu_inst_pe_1_2_7_n4), .Z(
        npu_inst_pe_1_2_7_n17) );
  MUX2_X1 npu_inst_pe_1_2_7_U144 ( .A(npu_inst_pe_1_2_7_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_2_7_int_q_reg_h_3__0_), .S(npu_inst_pe_1_2_7_n4), .Z(
        npu_inst_pe_1_2_7_n16) );
  MUX2_X1 npu_inst_pe_1_2_7_U143 ( .A(npu_inst_pe_1_2_7_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_2_7_int_q_reg_h_5__0_), .S(npu_inst_pe_1_2_7_n4), .Z(
        npu_inst_pe_1_2_7_n15) );
  XOR2_X1 npu_inst_pe_1_2_7_U142 ( .A(npu_inst_pe_1_2_7_int_data_0_), .B(
        npu_inst_pe_1_2_7_int_q_acc_0_), .Z(npu_inst_pe_1_2_7_N73) );
  AND2_X1 npu_inst_pe_1_2_7_U141 ( .A1(npu_inst_pe_1_2_7_int_q_acc_0_), .A2(
        npu_inst_pe_1_2_7_int_data_0_), .ZN(npu_inst_pe_1_2_7_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_2_7_U140 ( .A(npu_inst_pe_1_2_7_int_q_acc_0_), .B(
        npu_inst_pe_1_2_7_n13), .ZN(npu_inst_pe_1_2_7_N65) );
  OR2_X1 npu_inst_pe_1_2_7_U139 ( .A1(npu_inst_pe_1_2_7_n13), .A2(
        npu_inst_pe_1_2_7_int_q_acc_0_), .ZN(npu_inst_pe_1_2_7_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_2_7_U138 ( .A(npu_inst_pe_1_2_7_int_q_acc_2_), .B(
        npu_inst_pe_1_2_7_add_69_carry_2_), .Z(npu_inst_pe_1_2_7_N75) );
  AND2_X1 npu_inst_pe_1_2_7_U137 ( .A1(npu_inst_pe_1_2_7_add_69_carry_2_), 
        .A2(npu_inst_pe_1_2_7_int_q_acc_2_), .ZN(
        npu_inst_pe_1_2_7_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_2_7_U136 ( .A(npu_inst_pe_1_2_7_int_q_acc_3_), .B(
        npu_inst_pe_1_2_7_add_69_carry_3_), .Z(npu_inst_pe_1_2_7_N76) );
  AND2_X1 npu_inst_pe_1_2_7_U135 ( .A1(npu_inst_pe_1_2_7_add_69_carry_3_), 
        .A2(npu_inst_pe_1_2_7_int_q_acc_3_), .ZN(
        npu_inst_pe_1_2_7_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_2_7_U134 ( .A(npu_inst_pe_1_2_7_int_q_acc_4_), .B(
        npu_inst_pe_1_2_7_add_69_carry_4_), .Z(npu_inst_pe_1_2_7_N77) );
  AND2_X1 npu_inst_pe_1_2_7_U133 ( .A1(npu_inst_pe_1_2_7_add_69_carry_4_), 
        .A2(npu_inst_pe_1_2_7_int_q_acc_4_), .ZN(
        npu_inst_pe_1_2_7_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_2_7_U132 ( .A(npu_inst_pe_1_2_7_int_q_acc_5_), .B(
        npu_inst_pe_1_2_7_add_69_carry_5_), .Z(npu_inst_pe_1_2_7_N78) );
  AND2_X1 npu_inst_pe_1_2_7_U131 ( .A1(npu_inst_pe_1_2_7_add_69_carry_5_), 
        .A2(npu_inst_pe_1_2_7_int_q_acc_5_), .ZN(
        npu_inst_pe_1_2_7_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_2_7_U130 ( .A(npu_inst_pe_1_2_7_int_q_acc_6_), .B(
        npu_inst_pe_1_2_7_add_69_carry_6_), .Z(npu_inst_pe_1_2_7_N79) );
  AND2_X1 npu_inst_pe_1_2_7_U129 ( .A1(npu_inst_pe_1_2_7_add_69_carry_6_), 
        .A2(npu_inst_pe_1_2_7_int_q_acc_6_), .ZN(
        npu_inst_pe_1_2_7_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_2_7_U128 ( .A(npu_inst_pe_1_2_7_int_q_acc_7_), .B(
        npu_inst_pe_1_2_7_add_69_carry_7_), .Z(npu_inst_pe_1_2_7_N80) );
  XNOR2_X1 npu_inst_pe_1_2_7_U127 ( .A(npu_inst_pe_1_2_7_sub_67_carry_2_), .B(
        npu_inst_pe_1_2_7_int_q_acc_2_), .ZN(npu_inst_pe_1_2_7_N67) );
  OR2_X1 npu_inst_pe_1_2_7_U126 ( .A1(npu_inst_pe_1_2_7_int_q_acc_2_), .A2(
        npu_inst_pe_1_2_7_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_2_7_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_2_7_U125 ( .A(npu_inst_pe_1_2_7_sub_67_carry_3_), .B(
        npu_inst_pe_1_2_7_int_q_acc_3_), .ZN(npu_inst_pe_1_2_7_N68) );
  OR2_X1 npu_inst_pe_1_2_7_U124 ( .A1(npu_inst_pe_1_2_7_int_q_acc_3_), .A2(
        npu_inst_pe_1_2_7_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_2_7_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_2_7_U123 ( .A(npu_inst_pe_1_2_7_sub_67_carry_4_), .B(
        npu_inst_pe_1_2_7_int_q_acc_4_), .ZN(npu_inst_pe_1_2_7_N69) );
  OR2_X1 npu_inst_pe_1_2_7_U122 ( .A1(npu_inst_pe_1_2_7_int_q_acc_4_), .A2(
        npu_inst_pe_1_2_7_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_2_7_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_2_7_U121 ( .A(npu_inst_pe_1_2_7_sub_67_carry_5_), .B(
        npu_inst_pe_1_2_7_int_q_acc_5_), .ZN(npu_inst_pe_1_2_7_N70) );
  OR2_X1 npu_inst_pe_1_2_7_U120 ( .A1(npu_inst_pe_1_2_7_int_q_acc_5_), .A2(
        npu_inst_pe_1_2_7_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_2_7_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_2_7_U119 ( .A(npu_inst_pe_1_2_7_sub_67_carry_6_), .B(
        npu_inst_pe_1_2_7_int_q_acc_6_), .ZN(npu_inst_pe_1_2_7_N71) );
  OR2_X1 npu_inst_pe_1_2_7_U118 ( .A1(npu_inst_pe_1_2_7_int_q_acc_6_), .A2(
        npu_inst_pe_1_2_7_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_2_7_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_2_7_U117 ( .A(npu_inst_pe_1_2_7_int_q_acc_7_), .B(
        npu_inst_pe_1_2_7_sub_67_carry_7_), .ZN(npu_inst_pe_1_2_7_N72) );
  INV_X1 npu_inst_pe_1_2_7_U116 ( .A(npu_inst_n78), .ZN(npu_inst_pe_1_2_7_n7)
         );
  INV_X1 npu_inst_pe_1_2_7_U115 ( .A(npu_inst_pe_1_2_7_n7), .ZN(
        npu_inst_pe_1_2_7_n6) );
  INV_X1 npu_inst_pe_1_2_7_U114 ( .A(npu_inst_n57), .ZN(npu_inst_pe_1_2_7_n3)
         );
  AOI22_X1 npu_inst_pe_1_2_7_U113 ( .A1(npu_inst_int_data_y_3__7__0_), .A2(
        npu_inst_pe_1_2_7_n58), .B1(npu_inst_pe_1_2_7_n119), .B2(
        npu_inst_pe_1_2_7_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_2_7_n57) );
  INV_X1 npu_inst_pe_1_2_7_U112 ( .A(npu_inst_pe_1_2_7_n57), .ZN(
        npu_inst_pe_1_2_7_n108) );
  AOI22_X1 npu_inst_pe_1_2_7_U111 ( .A1(npu_inst_int_data_y_3__7__0_), .A2(
        npu_inst_pe_1_2_7_n54), .B1(npu_inst_pe_1_2_7_n118), .B2(
        npu_inst_pe_1_2_7_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_2_7_n53) );
  INV_X1 npu_inst_pe_1_2_7_U110 ( .A(npu_inst_pe_1_2_7_n53), .ZN(
        npu_inst_pe_1_2_7_n109) );
  AOI22_X1 npu_inst_pe_1_2_7_U107 ( .A1(npu_inst_int_data_y_3__7__0_), .A2(
        npu_inst_pe_1_2_7_n50), .B1(npu_inst_pe_1_2_7_n117), .B2(
        npu_inst_pe_1_2_7_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_2_7_n49) );
  INV_X1 npu_inst_pe_1_2_7_U106 ( .A(npu_inst_pe_1_2_7_n49), .ZN(
        npu_inst_pe_1_2_7_n110) );
  AOI22_X1 npu_inst_pe_1_2_7_U105 ( .A1(npu_inst_int_data_y_3__7__0_), .A2(
        npu_inst_pe_1_2_7_n46), .B1(npu_inst_pe_1_2_7_n116), .B2(
        npu_inst_pe_1_2_7_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_2_7_n45) );
  INV_X1 npu_inst_pe_1_2_7_U104 ( .A(npu_inst_pe_1_2_7_n45), .ZN(
        npu_inst_pe_1_2_7_n111) );
  AOI22_X1 npu_inst_pe_1_2_7_U103 ( .A1(npu_inst_int_data_y_3__7__0_), .A2(
        npu_inst_pe_1_2_7_n42), .B1(npu_inst_pe_1_2_7_n115), .B2(
        npu_inst_pe_1_2_7_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_2_7_n41) );
  INV_X1 npu_inst_pe_1_2_7_U102 ( .A(npu_inst_pe_1_2_7_n41), .ZN(
        npu_inst_pe_1_2_7_n112) );
  AOI22_X1 npu_inst_pe_1_2_7_U101 ( .A1(npu_inst_int_data_y_3__7__1_), .A2(
        npu_inst_pe_1_2_7_n58), .B1(npu_inst_pe_1_2_7_n119), .B2(
        npu_inst_pe_1_2_7_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_2_7_n59) );
  INV_X1 npu_inst_pe_1_2_7_U100 ( .A(npu_inst_pe_1_2_7_n59), .ZN(
        npu_inst_pe_1_2_7_n102) );
  AOI22_X1 npu_inst_pe_1_2_7_U99 ( .A1(npu_inst_int_data_y_3__7__1_), .A2(
        npu_inst_pe_1_2_7_n54), .B1(npu_inst_pe_1_2_7_n118), .B2(
        npu_inst_pe_1_2_7_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_2_7_n55) );
  INV_X1 npu_inst_pe_1_2_7_U98 ( .A(npu_inst_pe_1_2_7_n55), .ZN(
        npu_inst_pe_1_2_7_n103) );
  AOI22_X1 npu_inst_pe_1_2_7_U97 ( .A1(npu_inst_int_data_y_3__7__1_), .A2(
        npu_inst_pe_1_2_7_n50), .B1(npu_inst_pe_1_2_7_n117), .B2(
        npu_inst_pe_1_2_7_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_2_7_n51) );
  INV_X1 npu_inst_pe_1_2_7_U96 ( .A(npu_inst_pe_1_2_7_n51), .ZN(
        npu_inst_pe_1_2_7_n104) );
  AOI22_X1 npu_inst_pe_1_2_7_U95 ( .A1(npu_inst_int_data_y_3__7__1_), .A2(
        npu_inst_pe_1_2_7_n46), .B1(npu_inst_pe_1_2_7_n116), .B2(
        npu_inst_pe_1_2_7_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_2_7_n47) );
  INV_X1 npu_inst_pe_1_2_7_U94 ( .A(npu_inst_pe_1_2_7_n47), .ZN(
        npu_inst_pe_1_2_7_n105) );
  AOI22_X1 npu_inst_pe_1_2_7_U93 ( .A1(npu_inst_int_data_y_3__7__1_), .A2(
        npu_inst_pe_1_2_7_n42), .B1(npu_inst_pe_1_2_7_n115), .B2(
        npu_inst_pe_1_2_7_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_2_7_n43) );
  INV_X1 npu_inst_pe_1_2_7_U92 ( .A(npu_inst_pe_1_2_7_n43), .ZN(
        npu_inst_pe_1_2_7_n106) );
  AOI22_X1 npu_inst_pe_1_2_7_U91 ( .A1(npu_inst_pe_1_2_7_n38), .A2(
        npu_inst_int_data_y_3__7__1_), .B1(npu_inst_pe_1_2_7_n114), .B2(
        npu_inst_pe_1_2_7_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_2_7_n39) );
  INV_X1 npu_inst_pe_1_2_7_U90 ( .A(npu_inst_pe_1_2_7_n39), .ZN(
        npu_inst_pe_1_2_7_n107) );
  AOI22_X1 npu_inst_pe_1_2_7_U89 ( .A1(npu_inst_pe_1_2_7_n38), .A2(
        npu_inst_int_data_y_3__7__0_), .B1(npu_inst_pe_1_2_7_n114), .B2(
        npu_inst_pe_1_2_7_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_2_7_n37) );
  INV_X1 npu_inst_pe_1_2_7_U88 ( .A(npu_inst_pe_1_2_7_n37), .ZN(
        npu_inst_pe_1_2_7_n113) );
  AND2_X1 npu_inst_pe_1_2_7_U87 ( .A1(npu_inst_pe_1_2_7_N93), .A2(npu_inst_n57), .ZN(npu_inst_int_data_y_2__7__0_) );
  AND2_X1 npu_inst_pe_1_2_7_U86 ( .A1(npu_inst_n57), .A2(npu_inst_pe_1_2_7_N94), .ZN(npu_inst_int_data_y_2__7__1_) );
  NOR3_X1 npu_inst_pe_1_2_7_U85 ( .A1(npu_inst_pe_1_2_7_n26), .A2(npu_inst_n57), .A3(npu_inst_int_ckg[40]), .ZN(npu_inst_pe_1_2_7_n85) );
  OR2_X1 npu_inst_pe_1_2_7_U84 ( .A1(npu_inst_pe_1_2_7_n85), .A2(
        npu_inst_pe_1_2_7_n2), .ZN(npu_inst_pe_1_2_7_N84) );
  AND2_X1 npu_inst_pe_1_2_7_U83 ( .A1(npu_inst_pe_1_2_7_int_q_acc_0_), .A2(
        npu_inst_pe_1_2_7_n1), .ZN(npu_inst_int_data_res_2__7__0_) );
  AND2_X1 npu_inst_pe_1_2_7_U82 ( .A1(npu_inst_pe_1_2_7_n2), .A2(
        npu_inst_pe_1_2_7_int_q_acc_7_), .ZN(npu_inst_int_data_res_2__7__7_)
         );
  AND2_X1 npu_inst_pe_1_2_7_U81 ( .A1(npu_inst_pe_1_2_7_int_q_acc_1_), .A2(
        npu_inst_pe_1_2_7_n1), .ZN(npu_inst_int_data_res_2__7__1_) );
  AND2_X1 npu_inst_pe_1_2_7_U80 ( .A1(npu_inst_pe_1_2_7_int_q_acc_2_), .A2(
        npu_inst_pe_1_2_7_n1), .ZN(npu_inst_int_data_res_2__7__2_) );
  AND2_X1 npu_inst_pe_1_2_7_U79 ( .A1(npu_inst_pe_1_2_7_int_q_acc_3_), .A2(
        npu_inst_pe_1_2_7_n2), .ZN(npu_inst_int_data_res_2__7__3_) );
  AND2_X1 npu_inst_pe_1_2_7_U78 ( .A1(npu_inst_pe_1_2_7_int_q_acc_4_), .A2(
        npu_inst_pe_1_2_7_n2), .ZN(npu_inst_int_data_res_2__7__4_) );
  AND2_X1 npu_inst_pe_1_2_7_U77 ( .A1(npu_inst_pe_1_2_7_int_q_acc_5_), .A2(
        npu_inst_pe_1_2_7_n2), .ZN(npu_inst_int_data_res_2__7__5_) );
  AND2_X1 npu_inst_pe_1_2_7_U76 ( .A1(npu_inst_pe_1_2_7_int_q_acc_6_), .A2(
        npu_inst_pe_1_2_7_n2), .ZN(npu_inst_int_data_res_2__7__6_) );
  AOI222_X1 npu_inst_pe_1_2_7_U75 ( .A1(npu_inst_int_data_res_3__7__0_), .A2(
        npu_inst_pe_1_2_7_n1), .B1(npu_inst_pe_1_2_7_N73), .B2(
        npu_inst_pe_1_2_7_n76), .C1(npu_inst_pe_1_2_7_N65), .C2(
        npu_inst_pe_1_2_7_n77), .ZN(npu_inst_pe_1_2_7_n84) );
  INV_X1 npu_inst_pe_1_2_7_U74 ( .A(npu_inst_pe_1_2_7_n84), .ZN(
        npu_inst_pe_1_2_7_n101) );
  AOI222_X1 npu_inst_pe_1_2_7_U73 ( .A1(npu_inst_int_data_res_3__7__7_), .A2(
        npu_inst_pe_1_2_7_n1), .B1(npu_inst_pe_1_2_7_N80), .B2(
        npu_inst_pe_1_2_7_n76), .C1(npu_inst_pe_1_2_7_N72), .C2(
        npu_inst_pe_1_2_7_n77), .ZN(npu_inst_pe_1_2_7_n75) );
  INV_X1 npu_inst_pe_1_2_7_U72 ( .A(npu_inst_pe_1_2_7_n75), .ZN(
        npu_inst_pe_1_2_7_n33) );
  AOI222_X1 npu_inst_pe_1_2_7_U71 ( .A1(npu_inst_int_data_res_3__7__1_), .A2(
        npu_inst_pe_1_2_7_n1), .B1(npu_inst_pe_1_2_7_N74), .B2(
        npu_inst_pe_1_2_7_n76), .C1(npu_inst_pe_1_2_7_N66), .C2(
        npu_inst_pe_1_2_7_n77), .ZN(npu_inst_pe_1_2_7_n83) );
  INV_X1 npu_inst_pe_1_2_7_U70 ( .A(npu_inst_pe_1_2_7_n83), .ZN(
        npu_inst_pe_1_2_7_n100) );
  AOI222_X1 npu_inst_pe_1_2_7_U69 ( .A1(npu_inst_int_data_res_3__7__2_), .A2(
        npu_inst_pe_1_2_7_n1), .B1(npu_inst_pe_1_2_7_N75), .B2(
        npu_inst_pe_1_2_7_n76), .C1(npu_inst_pe_1_2_7_N67), .C2(
        npu_inst_pe_1_2_7_n77), .ZN(npu_inst_pe_1_2_7_n82) );
  INV_X1 npu_inst_pe_1_2_7_U68 ( .A(npu_inst_pe_1_2_7_n82), .ZN(
        npu_inst_pe_1_2_7_n99) );
  AOI222_X1 npu_inst_pe_1_2_7_U67 ( .A1(npu_inst_int_data_res_3__7__3_), .A2(
        npu_inst_pe_1_2_7_n1), .B1(npu_inst_pe_1_2_7_N76), .B2(
        npu_inst_pe_1_2_7_n76), .C1(npu_inst_pe_1_2_7_N68), .C2(
        npu_inst_pe_1_2_7_n77), .ZN(npu_inst_pe_1_2_7_n81) );
  INV_X1 npu_inst_pe_1_2_7_U66 ( .A(npu_inst_pe_1_2_7_n81), .ZN(
        npu_inst_pe_1_2_7_n98) );
  AOI222_X1 npu_inst_pe_1_2_7_U65 ( .A1(npu_inst_int_data_res_3__7__4_), .A2(
        npu_inst_pe_1_2_7_n1), .B1(npu_inst_pe_1_2_7_N77), .B2(
        npu_inst_pe_1_2_7_n76), .C1(npu_inst_pe_1_2_7_N69), .C2(
        npu_inst_pe_1_2_7_n77), .ZN(npu_inst_pe_1_2_7_n80) );
  INV_X1 npu_inst_pe_1_2_7_U64 ( .A(npu_inst_pe_1_2_7_n80), .ZN(
        npu_inst_pe_1_2_7_n36) );
  AOI222_X1 npu_inst_pe_1_2_7_U63 ( .A1(npu_inst_int_data_res_3__7__5_), .A2(
        npu_inst_pe_1_2_7_n1), .B1(npu_inst_pe_1_2_7_N78), .B2(
        npu_inst_pe_1_2_7_n76), .C1(npu_inst_pe_1_2_7_N70), .C2(
        npu_inst_pe_1_2_7_n77), .ZN(npu_inst_pe_1_2_7_n79) );
  INV_X1 npu_inst_pe_1_2_7_U62 ( .A(npu_inst_pe_1_2_7_n79), .ZN(
        npu_inst_pe_1_2_7_n35) );
  AOI222_X1 npu_inst_pe_1_2_7_U61 ( .A1(npu_inst_int_data_res_3__7__6_), .A2(
        npu_inst_pe_1_2_7_n1), .B1(npu_inst_pe_1_2_7_N79), .B2(
        npu_inst_pe_1_2_7_n76), .C1(npu_inst_pe_1_2_7_N71), .C2(
        npu_inst_pe_1_2_7_n77), .ZN(npu_inst_pe_1_2_7_n78) );
  INV_X1 npu_inst_pe_1_2_7_U60 ( .A(npu_inst_pe_1_2_7_n78), .ZN(
        npu_inst_pe_1_2_7_n34) );
  INV_X1 npu_inst_pe_1_2_7_U59 ( .A(npu_inst_pe_1_2_7_int_data_1_), .ZN(
        npu_inst_pe_1_2_7_n14) );
  AND2_X1 npu_inst_pe_1_2_7_U58 ( .A1(npu_inst_int_data_x_2__7__1_), .A2(
        npu_inst_pe_1_2_7_int_q_weight_1_), .ZN(npu_inst_pe_1_2_7_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_2_7_U57 ( .A1(npu_inst_int_data_x_2__7__0_), .A2(
        npu_inst_pe_1_2_7_int_q_weight_1_), .ZN(npu_inst_pe_1_2_7_int_data_0_)
         );
  NAND2_X1 npu_inst_pe_1_2_7_U56 ( .A1(npu_inst_pe_1_2_7_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_2_7_n60), .ZN(npu_inst_pe_1_2_7_n74) );
  OAI21_X1 npu_inst_pe_1_2_7_U55 ( .B1(npu_inst_pe_1_2_7_n63), .B2(
        npu_inst_pe_1_2_7_n60), .A(npu_inst_pe_1_2_7_n74), .ZN(
        npu_inst_pe_1_2_7_n97) );
  NAND2_X1 npu_inst_pe_1_2_7_U54 ( .A1(npu_inst_pe_1_2_7_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_2_7_n60), .ZN(npu_inst_pe_1_2_7_n73) );
  OAI21_X1 npu_inst_pe_1_2_7_U53 ( .B1(npu_inst_pe_1_2_7_n61), .B2(
        npu_inst_pe_1_2_7_n60), .A(npu_inst_pe_1_2_7_n73), .ZN(
        npu_inst_pe_1_2_7_n96) );
  NAND2_X1 npu_inst_pe_1_2_7_U52 ( .A1(npu_inst_pe_1_2_7_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_2_7_n56), .ZN(npu_inst_pe_1_2_7_n72) );
  OAI21_X1 npu_inst_pe_1_2_7_U51 ( .B1(npu_inst_pe_1_2_7_n63), .B2(
        npu_inst_pe_1_2_7_n56), .A(npu_inst_pe_1_2_7_n72), .ZN(
        npu_inst_pe_1_2_7_n95) );
  NAND2_X1 npu_inst_pe_1_2_7_U50 ( .A1(npu_inst_pe_1_2_7_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_2_7_n56), .ZN(npu_inst_pe_1_2_7_n71) );
  OAI21_X1 npu_inst_pe_1_2_7_U49 ( .B1(npu_inst_pe_1_2_7_n61), .B2(
        npu_inst_pe_1_2_7_n56), .A(npu_inst_pe_1_2_7_n71), .ZN(
        npu_inst_pe_1_2_7_n94) );
  NAND2_X1 npu_inst_pe_1_2_7_U48 ( .A1(npu_inst_pe_1_2_7_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_2_7_n52), .ZN(npu_inst_pe_1_2_7_n70) );
  OAI21_X1 npu_inst_pe_1_2_7_U47 ( .B1(npu_inst_pe_1_2_7_n63), .B2(
        npu_inst_pe_1_2_7_n52), .A(npu_inst_pe_1_2_7_n70), .ZN(
        npu_inst_pe_1_2_7_n93) );
  NAND2_X1 npu_inst_pe_1_2_7_U46 ( .A1(npu_inst_pe_1_2_7_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_2_7_n52), .ZN(npu_inst_pe_1_2_7_n69) );
  OAI21_X1 npu_inst_pe_1_2_7_U45 ( .B1(npu_inst_pe_1_2_7_n61), .B2(
        npu_inst_pe_1_2_7_n52), .A(npu_inst_pe_1_2_7_n69), .ZN(
        npu_inst_pe_1_2_7_n92) );
  NAND2_X1 npu_inst_pe_1_2_7_U44 ( .A1(npu_inst_pe_1_2_7_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_2_7_n48), .ZN(npu_inst_pe_1_2_7_n68) );
  OAI21_X1 npu_inst_pe_1_2_7_U43 ( .B1(npu_inst_pe_1_2_7_n63), .B2(
        npu_inst_pe_1_2_7_n48), .A(npu_inst_pe_1_2_7_n68), .ZN(
        npu_inst_pe_1_2_7_n91) );
  NAND2_X1 npu_inst_pe_1_2_7_U42 ( .A1(npu_inst_pe_1_2_7_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_2_7_n48), .ZN(npu_inst_pe_1_2_7_n67) );
  OAI21_X1 npu_inst_pe_1_2_7_U41 ( .B1(npu_inst_pe_1_2_7_n61), .B2(
        npu_inst_pe_1_2_7_n48), .A(npu_inst_pe_1_2_7_n67), .ZN(
        npu_inst_pe_1_2_7_n90) );
  NAND2_X1 npu_inst_pe_1_2_7_U40 ( .A1(npu_inst_pe_1_2_7_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_2_7_n44), .ZN(npu_inst_pe_1_2_7_n66) );
  OAI21_X1 npu_inst_pe_1_2_7_U39 ( .B1(npu_inst_pe_1_2_7_n63), .B2(
        npu_inst_pe_1_2_7_n44), .A(npu_inst_pe_1_2_7_n66), .ZN(
        npu_inst_pe_1_2_7_n89) );
  NAND2_X1 npu_inst_pe_1_2_7_U38 ( .A1(npu_inst_pe_1_2_7_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_2_7_n44), .ZN(npu_inst_pe_1_2_7_n65) );
  OAI21_X1 npu_inst_pe_1_2_7_U37 ( .B1(npu_inst_pe_1_2_7_n61), .B2(
        npu_inst_pe_1_2_7_n44), .A(npu_inst_pe_1_2_7_n65), .ZN(
        npu_inst_pe_1_2_7_n88) );
  NAND2_X1 npu_inst_pe_1_2_7_U36 ( .A1(npu_inst_pe_1_2_7_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_2_7_n40), .ZN(npu_inst_pe_1_2_7_n64) );
  OAI21_X1 npu_inst_pe_1_2_7_U35 ( .B1(npu_inst_pe_1_2_7_n63), .B2(
        npu_inst_pe_1_2_7_n40), .A(npu_inst_pe_1_2_7_n64), .ZN(
        npu_inst_pe_1_2_7_n87) );
  NAND2_X1 npu_inst_pe_1_2_7_U34 ( .A1(npu_inst_pe_1_2_7_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_2_7_n40), .ZN(npu_inst_pe_1_2_7_n62) );
  OAI21_X1 npu_inst_pe_1_2_7_U33 ( .B1(npu_inst_pe_1_2_7_n61), .B2(
        npu_inst_pe_1_2_7_n40), .A(npu_inst_pe_1_2_7_n62), .ZN(
        npu_inst_pe_1_2_7_n86) );
  INV_X1 npu_inst_pe_1_2_7_U32 ( .A(npu_inst_pe_1_2_7_int_data_0_), .ZN(
        npu_inst_pe_1_2_7_n13) );
  INV_X1 npu_inst_pe_1_2_7_U31 ( .A(npu_inst_n70), .ZN(npu_inst_pe_1_2_7_n5)
         );
  AOI22_X1 npu_inst_pe_1_2_7_U30 ( .A1(npu_inst_n57), .A2(
        npu_inst_int_data_y_3__7__1_), .B1(npu_inst_pe_1_2_7_n3), .B2(
        int_i_data_h_npu[11]), .ZN(npu_inst_pe_1_2_7_n63) );
  AOI22_X1 npu_inst_pe_1_2_7_U29 ( .A1(npu_inst_n57), .A2(
        npu_inst_int_data_y_3__7__0_), .B1(npu_inst_pe_1_2_7_n3), .B2(
        int_i_data_h_npu[10]), .ZN(npu_inst_pe_1_2_7_n61) );
  OR3_X1 npu_inst_pe_1_2_7_U28 ( .A1(npu_inst_pe_1_2_7_n6), .A2(
        npu_inst_pe_1_2_7_n8), .A3(npu_inst_pe_1_2_7_n5), .ZN(
        npu_inst_pe_1_2_7_n56) );
  OR3_X1 npu_inst_pe_1_2_7_U27 ( .A1(npu_inst_pe_1_2_7_n5), .A2(
        npu_inst_pe_1_2_7_n8), .A3(npu_inst_pe_1_2_7_n7), .ZN(
        npu_inst_pe_1_2_7_n48) );
  INV_X1 npu_inst_pe_1_2_7_U26 ( .A(npu_inst_pe_1_2_7_n5), .ZN(
        npu_inst_pe_1_2_7_n4) );
  OR3_X1 npu_inst_pe_1_2_7_U25 ( .A1(npu_inst_pe_1_2_7_n4), .A2(
        npu_inst_pe_1_2_7_n8), .A3(npu_inst_pe_1_2_7_n7), .ZN(
        npu_inst_pe_1_2_7_n52) );
  OR3_X1 npu_inst_pe_1_2_7_U24 ( .A1(npu_inst_pe_1_2_7_n6), .A2(
        npu_inst_pe_1_2_7_n8), .A3(npu_inst_pe_1_2_7_n4), .ZN(
        npu_inst_pe_1_2_7_n60) );
  NOR2_X1 npu_inst_pe_1_2_7_U23 ( .A1(npu_inst_pe_1_2_7_n60), .A2(
        npu_inst_pe_1_2_7_n3), .ZN(npu_inst_pe_1_2_7_n58) );
  NOR2_X1 npu_inst_pe_1_2_7_U22 ( .A1(npu_inst_pe_1_2_7_n56), .A2(
        npu_inst_pe_1_2_7_n3), .ZN(npu_inst_pe_1_2_7_n54) );
  NOR2_X1 npu_inst_pe_1_2_7_U21 ( .A1(npu_inst_pe_1_2_7_n52), .A2(
        npu_inst_pe_1_2_7_n3), .ZN(npu_inst_pe_1_2_7_n50) );
  NOR2_X1 npu_inst_pe_1_2_7_U20 ( .A1(npu_inst_pe_1_2_7_n48), .A2(
        npu_inst_pe_1_2_7_n3), .ZN(npu_inst_pe_1_2_7_n46) );
  NOR2_X1 npu_inst_pe_1_2_7_U19 ( .A1(npu_inst_pe_1_2_7_n40), .A2(
        npu_inst_pe_1_2_7_n3), .ZN(npu_inst_pe_1_2_7_n38) );
  NOR2_X1 npu_inst_pe_1_2_7_U18 ( .A1(npu_inst_pe_1_2_7_n44), .A2(
        npu_inst_pe_1_2_7_n3), .ZN(npu_inst_pe_1_2_7_n42) );
  BUF_X1 npu_inst_pe_1_2_7_U17 ( .A(npu_inst_n102), .Z(npu_inst_pe_1_2_7_n8)
         );
  INV_X1 npu_inst_pe_1_2_7_U16 ( .A(npu_inst_n125), .ZN(npu_inst_pe_1_2_7_n12)
         );
  INV_X1 npu_inst_pe_1_2_7_U15 ( .A(npu_inst_pe_1_2_7_n38), .ZN(
        npu_inst_pe_1_2_7_n114) );
  INV_X1 npu_inst_pe_1_2_7_U14 ( .A(npu_inst_pe_1_2_7_n58), .ZN(
        npu_inst_pe_1_2_7_n119) );
  INV_X1 npu_inst_pe_1_2_7_U13 ( .A(npu_inst_pe_1_2_7_n54), .ZN(
        npu_inst_pe_1_2_7_n118) );
  INV_X1 npu_inst_pe_1_2_7_U12 ( .A(npu_inst_pe_1_2_7_n50), .ZN(
        npu_inst_pe_1_2_7_n117) );
  INV_X1 npu_inst_pe_1_2_7_U11 ( .A(npu_inst_pe_1_2_7_n46), .ZN(
        npu_inst_pe_1_2_7_n116) );
  INV_X1 npu_inst_pe_1_2_7_U10 ( .A(npu_inst_pe_1_2_7_n42), .ZN(
        npu_inst_pe_1_2_7_n115) );
  BUF_X1 npu_inst_pe_1_2_7_U9 ( .A(npu_inst_n27), .Z(npu_inst_pe_1_2_7_n2) );
  BUF_X1 npu_inst_pe_1_2_7_U8 ( .A(npu_inst_n27), .Z(npu_inst_pe_1_2_7_n1) );
  BUF_X1 npu_inst_pe_1_2_7_U7 ( .A(npu_inst_pe_1_2_7_n12), .Z(
        npu_inst_pe_1_2_7_n11) );
  BUF_X1 npu_inst_pe_1_2_7_U6 ( .A(npu_inst_pe_1_2_7_n12), .Z(
        npu_inst_pe_1_2_7_n10) );
  BUF_X1 npu_inst_pe_1_2_7_U5 ( .A(npu_inst_pe_1_2_7_n12), .Z(
        npu_inst_pe_1_2_7_n9) );
  NOR2_X1 npu_inst_pe_1_2_7_U4 ( .A1(npu_inst_pe_1_2_7_int_q_weight_0_), .A2(
        npu_inst_pe_1_2_7_n1), .ZN(npu_inst_pe_1_2_7_n76) );
  NOR2_X1 npu_inst_pe_1_2_7_U3 ( .A1(npu_inst_pe_1_2_7_n27), .A2(
        npu_inst_pe_1_2_7_n1), .ZN(npu_inst_pe_1_2_7_n77) );
  FA_X1 npu_inst_pe_1_2_7_sub_67_U2_1 ( .A(npu_inst_pe_1_2_7_int_q_acc_1_), 
        .B(npu_inst_pe_1_2_7_n14), .CI(npu_inst_pe_1_2_7_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_2_7_sub_67_carry_2_), .S(npu_inst_pe_1_2_7_N66) );
  FA_X1 npu_inst_pe_1_2_7_add_69_U1_1 ( .A(npu_inst_pe_1_2_7_int_q_acc_1_), 
        .B(npu_inst_pe_1_2_7_int_data_1_), .CI(
        npu_inst_pe_1_2_7_add_69_carry_1_), .CO(
        npu_inst_pe_1_2_7_add_69_carry_2_), .S(npu_inst_pe_1_2_7_N74) );
  NAND3_X1 npu_inst_pe_1_2_7_U109 ( .A1(npu_inst_pe_1_2_7_n5), .A2(
        npu_inst_pe_1_2_7_n7), .A3(npu_inst_pe_1_2_7_n8), .ZN(
        npu_inst_pe_1_2_7_n44) );
  NAND3_X1 npu_inst_pe_1_2_7_U108 ( .A1(npu_inst_pe_1_2_7_n4), .A2(
        npu_inst_pe_1_2_7_n7), .A3(npu_inst_pe_1_2_7_n8), .ZN(
        npu_inst_pe_1_2_7_n40) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_2_7_n34), .CK(
        npu_inst_pe_1_2_7_net4033), .RN(npu_inst_pe_1_2_7_n9), .Q(
        npu_inst_pe_1_2_7_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_2_7_n35), .CK(
        npu_inst_pe_1_2_7_net4033), .RN(npu_inst_pe_1_2_7_n9), .Q(
        npu_inst_pe_1_2_7_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_2_7_n36), .CK(
        npu_inst_pe_1_2_7_net4033), .RN(npu_inst_pe_1_2_7_n9), .Q(
        npu_inst_pe_1_2_7_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_2_7_n98), .CK(
        npu_inst_pe_1_2_7_net4033), .RN(npu_inst_pe_1_2_7_n9), .Q(
        npu_inst_pe_1_2_7_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_2_7_n99), .CK(
        npu_inst_pe_1_2_7_net4033), .RN(npu_inst_pe_1_2_7_n9), .Q(
        npu_inst_pe_1_2_7_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_2_7_n100), 
        .CK(npu_inst_pe_1_2_7_net4033), .RN(npu_inst_pe_1_2_7_n9), .Q(
        npu_inst_pe_1_2_7_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_2_7_n33), .CK(
        npu_inst_pe_1_2_7_net4033), .RN(npu_inst_pe_1_2_7_n9), .Q(
        npu_inst_pe_1_2_7_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_2_7_n101), 
        .CK(npu_inst_pe_1_2_7_net4033), .RN(npu_inst_pe_1_2_7_n9), .Q(
        npu_inst_pe_1_2_7_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_weight_reg_0_ ( .D(npu_inst_n111), .CK(
        npu_inst_pe_1_2_7_net4039), .RN(npu_inst_pe_1_2_7_n9), .Q(
        npu_inst_pe_1_2_7_int_q_weight_0_), .QN(npu_inst_pe_1_2_7_n27) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_weight_reg_1_ ( .D(npu_inst_n117), .CK(
        npu_inst_pe_1_2_7_net4039), .RN(npu_inst_pe_1_2_7_n9), .Q(
        npu_inst_pe_1_2_7_int_q_weight_1_), .QN(npu_inst_pe_1_2_7_n26) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_2_7_n113), 
        .CK(npu_inst_pe_1_2_7_net4039), .RN(npu_inst_pe_1_2_7_n9), .Q(
        npu_inst_pe_1_2_7_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_2_7_n107), 
        .CK(npu_inst_pe_1_2_7_net4039), .RN(npu_inst_pe_1_2_7_n9), .Q(
        npu_inst_pe_1_2_7_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_2_7_n112), 
        .CK(npu_inst_pe_1_2_7_net4039), .RN(npu_inst_pe_1_2_7_n10), .Q(
        npu_inst_pe_1_2_7_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_2_7_n106), 
        .CK(npu_inst_pe_1_2_7_net4039), .RN(npu_inst_pe_1_2_7_n10), .Q(
        npu_inst_pe_1_2_7_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_2_7_n111), 
        .CK(npu_inst_pe_1_2_7_net4039), .RN(npu_inst_pe_1_2_7_n10), .Q(
        npu_inst_pe_1_2_7_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_2_7_n105), 
        .CK(npu_inst_pe_1_2_7_net4039), .RN(npu_inst_pe_1_2_7_n10), .Q(
        npu_inst_pe_1_2_7_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_2_7_n110), 
        .CK(npu_inst_pe_1_2_7_net4039), .RN(npu_inst_pe_1_2_7_n10), .Q(
        npu_inst_pe_1_2_7_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_2_7_n104), 
        .CK(npu_inst_pe_1_2_7_net4039), .RN(npu_inst_pe_1_2_7_n10), .Q(
        npu_inst_pe_1_2_7_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_2_7_n109), 
        .CK(npu_inst_pe_1_2_7_net4039), .RN(npu_inst_pe_1_2_7_n10), .Q(
        npu_inst_pe_1_2_7_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_2_7_n103), 
        .CK(npu_inst_pe_1_2_7_net4039), .RN(npu_inst_pe_1_2_7_n10), .Q(
        npu_inst_pe_1_2_7_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_2_7_n108), 
        .CK(npu_inst_pe_1_2_7_net4039), .RN(npu_inst_pe_1_2_7_n10), .Q(
        npu_inst_pe_1_2_7_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_2_7_n102), 
        .CK(npu_inst_pe_1_2_7_net4039), .RN(npu_inst_pe_1_2_7_n10), .Q(
        npu_inst_pe_1_2_7_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_2_7_n86), 
        .CK(npu_inst_pe_1_2_7_net4039), .RN(npu_inst_pe_1_2_7_n10), .Q(
        npu_inst_pe_1_2_7_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_2_7_n87), 
        .CK(npu_inst_pe_1_2_7_net4039), .RN(npu_inst_pe_1_2_7_n10), .Q(
        npu_inst_pe_1_2_7_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_2_7_n88), 
        .CK(npu_inst_pe_1_2_7_net4039), .RN(npu_inst_pe_1_2_7_n11), .Q(
        npu_inst_pe_1_2_7_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_2_7_n89), 
        .CK(npu_inst_pe_1_2_7_net4039), .RN(npu_inst_pe_1_2_7_n11), .Q(
        npu_inst_pe_1_2_7_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_2_7_n90), 
        .CK(npu_inst_pe_1_2_7_net4039), .RN(npu_inst_pe_1_2_7_n11), .Q(
        npu_inst_pe_1_2_7_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_2_7_n91), 
        .CK(npu_inst_pe_1_2_7_net4039), .RN(npu_inst_pe_1_2_7_n11), .Q(
        npu_inst_pe_1_2_7_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_2_7_n92), 
        .CK(npu_inst_pe_1_2_7_net4039), .RN(npu_inst_pe_1_2_7_n11), .Q(
        npu_inst_pe_1_2_7_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_2_7_n93), 
        .CK(npu_inst_pe_1_2_7_net4039), .RN(npu_inst_pe_1_2_7_n11), .Q(
        npu_inst_pe_1_2_7_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_2_7_n94), 
        .CK(npu_inst_pe_1_2_7_net4039), .RN(npu_inst_pe_1_2_7_n11), .Q(
        npu_inst_pe_1_2_7_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_2_7_n95), 
        .CK(npu_inst_pe_1_2_7_net4039), .RN(npu_inst_pe_1_2_7_n11), .Q(
        npu_inst_pe_1_2_7_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_2_7_n96), 
        .CK(npu_inst_pe_1_2_7_net4039), .RN(npu_inst_pe_1_2_7_n11), .Q(
        npu_inst_pe_1_2_7_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_2_7_n97), 
        .CK(npu_inst_pe_1_2_7_net4039), .RN(npu_inst_pe_1_2_7_n11), .Q(
        npu_inst_pe_1_2_7_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_2_7_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_2_7_N84), .SE(1'b0), .GCK(npu_inst_pe_1_2_7_net4033) );
  CLKGATETST_X1 npu_inst_pe_1_2_7_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n64), .SE(1'b0), .GCK(npu_inst_pe_1_2_7_net4039) );
  MUX2_X1 npu_inst_pe_1_3_0_U162 ( .A(npu_inst_pe_1_3_0_n32), .B(
        npu_inst_pe_1_3_0_n29), .S(npu_inst_pe_1_3_0_n8), .Z(
        npu_inst_pe_1_3_0_N93) );
  MUX2_X1 npu_inst_pe_1_3_0_U161 ( .A(npu_inst_pe_1_3_0_n31), .B(
        npu_inst_pe_1_3_0_n30), .S(npu_inst_pe_1_3_0_n6), .Z(
        npu_inst_pe_1_3_0_n32) );
  MUX2_X1 npu_inst_pe_1_3_0_U160 ( .A(npu_inst_pe_1_3_0_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_3_0_int_q_reg_v_1__0_), .S(npu_inst_pe_1_3_0_n4), .Z(
        npu_inst_pe_1_3_0_n31) );
  MUX2_X1 npu_inst_pe_1_3_0_U159 ( .A(npu_inst_pe_1_3_0_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_3_0_int_q_reg_v_3__0_), .S(npu_inst_pe_1_3_0_n4), .Z(
        npu_inst_pe_1_3_0_n30) );
  MUX2_X1 npu_inst_pe_1_3_0_U158 ( .A(npu_inst_pe_1_3_0_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_3_0_int_q_reg_v_5__0_), .S(npu_inst_pe_1_3_0_n4), .Z(
        npu_inst_pe_1_3_0_n29) );
  MUX2_X1 npu_inst_pe_1_3_0_U157 ( .A(npu_inst_pe_1_3_0_n28), .B(
        npu_inst_pe_1_3_0_n23), .S(npu_inst_pe_1_3_0_n8), .Z(
        npu_inst_pe_1_3_0_N94) );
  MUX2_X1 npu_inst_pe_1_3_0_U156 ( .A(npu_inst_pe_1_3_0_n25), .B(
        npu_inst_pe_1_3_0_n24), .S(npu_inst_pe_1_3_0_n6), .Z(
        npu_inst_pe_1_3_0_n28) );
  MUX2_X1 npu_inst_pe_1_3_0_U155 ( .A(npu_inst_pe_1_3_0_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_3_0_int_q_reg_v_1__1_), .S(npu_inst_pe_1_3_0_n4), .Z(
        npu_inst_pe_1_3_0_n25) );
  MUX2_X1 npu_inst_pe_1_3_0_U154 ( .A(npu_inst_pe_1_3_0_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_3_0_int_q_reg_v_3__1_), .S(npu_inst_pe_1_3_0_n4), .Z(
        npu_inst_pe_1_3_0_n24) );
  MUX2_X1 npu_inst_pe_1_3_0_U153 ( .A(npu_inst_pe_1_3_0_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_3_0_int_q_reg_v_5__1_), .S(npu_inst_pe_1_3_0_n4), .Z(
        npu_inst_pe_1_3_0_n23) );
  MUX2_X1 npu_inst_pe_1_3_0_U152 ( .A(npu_inst_pe_1_3_0_n22), .B(
        npu_inst_pe_1_3_0_n19), .S(npu_inst_pe_1_3_0_n8), .Z(
        npu_inst_pe_1_3_0_o_data_h_1_) );
  MUX2_X1 npu_inst_pe_1_3_0_U151 ( .A(npu_inst_pe_1_3_0_n21), .B(
        npu_inst_pe_1_3_0_n20), .S(npu_inst_pe_1_3_0_n6), .Z(
        npu_inst_pe_1_3_0_n22) );
  MUX2_X1 npu_inst_pe_1_3_0_U150 ( .A(npu_inst_pe_1_3_0_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_3_0_int_q_reg_h_1__1_), .S(npu_inst_pe_1_3_0_n4), .Z(
        npu_inst_pe_1_3_0_n21) );
  MUX2_X1 npu_inst_pe_1_3_0_U149 ( .A(npu_inst_pe_1_3_0_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_3_0_int_q_reg_h_3__1_), .S(npu_inst_pe_1_3_0_n4), .Z(
        npu_inst_pe_1_3_0_n20) );
  MUX2_X1 npu_inst_pe_1_3_0_U148 ( .A(npu_inst_pe_1_3_0_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_3_0_int_q_reg_h_5__1_), .S(npu_inst_pe_1_3_0_n4), .Z(
        npu_inst_pe_1_3_0_n19) );
  MUX2_X1 npu_inst_pe_1_3_0_U147 ( .A(npu_inst_pe_1_3_0_n18), .B(
        npu_inst_pe_1_3_0_n15), .S(npu_inst_pe_1_3_0_n8), .Z(
        npu_inst_pe_1_3_0_o_data_h_0_) );
  MUX2_X1 npu_inst_pe_1_3_0_U146 ( .A(npu_inst_pe_1_3_0_n17), .B(
        npu_inst_pe_1_3_0_n16), .S(npu_inst_pe_1_3_0_n6), .Z(
        npu_inst_pe_1_3_0_n18) );
  MUX2_X1 npu_inst_pe_1_3_0_U145 ( .A(npu_inst_pe_1_3_0_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_3_0_int_q_reg_h_1__0_), .S(npu_inst_pe_1_3_0_n4), .Z(
        npu_inst_pe_1_3_0_n17) );
  MUX2_X1 npu_inst_pe_1_3_0_U144 ( .A(npu_inst_pe_1_3_0_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_3_0_int_q_reg_h_3__0_), .S(npu_inst_pe_1_3_0_n4), .Z(
        npu_inst_pe_1_3_0_n16) );
  MUX2_X1 npu_inst_pe_1_3_0_U143 ( .A(npu_inst_pe_1_3_0_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_3_0_int_q_reg_h_5__0_), .S(npu_inst_pe_1_3_0_n4), .Z(
        npu_inst_pe_1_3_0_n15) );
  XOR2_X1 npu_inst_pe_1_3_0_U142 ( .A(npu_inst_pe_1_3_0_int_data_0_), .B(
        npu_inst_pe_1_3_0_int_q_acc_0_), .Z(npu_inst_pe_1_3_0_N73) );
  AND2_X1 npu_inst_pe_1_3_0_U141 ( .A1(npu_inst_pe_1_3_0_int_q_acc_0_), .A2(
        npu_inst_pe_1_3_0_int_data_0_), .ZN(npu_inst_pe_1_3_0_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_3_0_U140 ( .A(npu_inst_pe_1_3_0_int_q_acc_0_), .B(
        npu_inst_pe_1_3_0_n13), .ZN(npu_inst_pe_1_3_0_N65) );
  OR2_X1 npu_inst_pe_1_3_0_U139 ( .A1(npu_inst_pe_1_3_0_n13), .A2(
        npu_inst_pe_1_3_0_int_q_acc_0_), .ZN(npu_inst_pe_1_3_0_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_3_0_U138 ( .A(npu_inst_pe_1_3_0_int_q_acc_2_), .B(
        npu_inst_pe_1_3_0_add_69_carry_2_), .Z(npu_inst_pe_1_3_0_N75) );
  AND2_X1 npu_inst_pe_1_3_0_U137 ( .A1(npu_inst_pe_1_3_0_add_69_carry_2_), 
        .A2(npu_inst_pe_1_3_0_int_q_acc_2_), .ZN(
        npu_inst_pe_1_3_0_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_3_0_U136 ( .A(npu_inst_pe_1_3_0_int_q_acc_3_), .B(
        npu_inst_pe_1_3_0_add_69_carry_3_), .Z(npu_inst_pe_1_3_0_N76) );
  AND2_X1 npu_inst_pe_1_3_0_U135 ( .A1(npu_inst_pe_1_3_0_add_69_carry_3_), 
        .A2(npu_inst_pe_1_3_0_int_q_acc_3_), .ZN(
        npu_inst_pe_1_3_0_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_3_0_U134 ( .A(npu_inst_pe_1_3_0_int_q_acc_4_), .B(
        npu_inst_pe_1_3_0_add_69_carry_4_), .Z(npu_inst_pe_1_3_0_N77) );
  AND2_X1 npu_inst_pe_1_3_0_U133 ( .A1(npu_inst_pe_1_3_0_add_69_carry_4_), 
        .A2(npu_inst_pe_1_3_0_int_q_acc_4_), .ZN(
        npu_inst_pe_1_3_0_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_3_0_U132 ( .A(npu_inst_pe_1_3_0_int_q_acc_5_), .B(
        npu_inst_pe_1_3_0_add_69_carry_5_), .Z(npu_inst_pe_1_3_0_N78) );
  AND2_X1 npu_inst_pe_1_3_0_U131 ( .A1(npu_inst_pe_1_3_0_add_69_carry_5_), 
        .A2(npu_inst_pe_1_3_0_int_q_acc_5_), .ZN(
        npu_inst_pe_1_3_0_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_3_0_U130 ( .A(npu_inst_pe_1_3_0_int_q_acc_6_), .B(
        npu_inst_pe_1_3_0_add_69_carry_6_), .Z(npu_inst_pe_1_3_0_N79) );
  AND2_X1 npu_inst_pe_1_3_0_U129 ( .A1(npu_inst_pe_1_3_0_add_69_carry_6_), 
        .A2(npu_inst_pe_1_3_0_int_q_acc_6_), .ZN(
        npu_inst_pe_1_3_0_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_3_0_U128 ( .A(npu_inst_pe_1_3_0_int_q_acc_7_), .B(
        npu_inst_pe_1_3_0_add_69_carry_7_), .Z(npu_inst_pe_1_3_0_N80) );
  XNOR2_X1 npu_inst_pe_1_3_0_U127 ( .A(npu_inst_pe_1_3_0_sub_67_carry_2_), .B(
        npu_inst_pe_1_3_0_int_q_acc_2_), .ZN(npu_inst_pe_1_3_0_N67) );
  OR2_X1 npu_inst_pe_1_3_0_U126 ( .A1(npu_inst_pe_1_3_0_int_q_acc_2_), .A2(
        npu_inst_pe_1_3_0_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_3_0_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_3_0_U125 ( .A(npu_inst_pe_1_3_0_sub_67_carry_3_), .B(
        npu_inst_pe_1_3_0_int_q_acc_3_), .ZN(npu_inst_pe_1_3_0_N68) );
  OR2_X1 npu_inst_pe_1_3_0_U124 ( .A1(npu_inst_pe_1_3_0_int_q_acc_3_), .A2(
        npu_inst_pe_1_3_0_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_3_0_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_3_0_U123 ( .A(npu_inst_pe_1_3_0_sub_67_carry_4_), .B(
        npu_inst_pe_1_3_0_int_q_acc_4_), .ZN(npu_inst_pe_1_3_0_N69) );
  OR2_X1 npu_inst_pe_1_3_0_U122 ( .A1(npu_inst_pe_1_3_0_int_q_acc_4_), .A2(
        npu_inst_pe_1_3_0_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_3_0_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_3_0_U121 ( .A(npu_inst_pe_1_3_0_sub_67_carry_5_), .B(
        npu_inst_pe_1_3_0_int_q_acc_5_), .ZN(npu_inst_pe_1_3_0_N70) );
  OR2_X1 npu_inst_pe_1_3_0_U120 ( .A1(npu_inst_pe_1_3_0_int_q_acc_5_), .A2(
        npu_inst_pe_1_3_0_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_3_0_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_3_0_U119 ( .A(npu_inst_pe_1_3_0_sub_67_carry_6_), .B(
        npu_inst_pe_1_3_0_int_q_acc_6_), .ZN(npu_inst_pe_1_3_0_N71) );
  OR2_X1 npu_inst_pe_1_3_0_U118 ( .A1(npu_inst_pe_1_3_0_int_q_acc_6_), .A2(
        npu_inst_pe_1_3_0_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_3_0_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_3_0_U117 ( .A(npu_inst_pe_1_3_0_int_q_acc_7_), .B(
        npu_inst_pe_1_3_0_sub_67_carry_7_), .ZN(npu_inst_pe_1_3_0_N72) );
  INV_X1 npu_inst_pe_1_3_0_U116 ( .A(npu_inst_n78), .ZN(npu_inst_pe_1_3_0_n7)
         );
  INV_X1 npu_inst_pe_1_3_0_U115 ( .A(npu_inst_pe_1_3_0_n7), .ZN(
        npu_inst_pe_1_3_0_n6) );
  INV_X1 npu_inst_pe_1_3_0_U114 ( .A(npu_inst_n57), .ZN(npu_inst_pe_1_3_0_n3)
         );
  AOI22_X1 npu_inst_pe_1_3_0_U113 ( .A1(npu_inst_int_data_y_4__0__0_), .A2(
        npu_inst_pe_1_3_0_n58), .B1(npu_inst_pe_1_3_0_n119), .B2(
        npu_inst_pe_1_3_0_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_3_0_n57) );
  INV_X1 npu_inst_pe_1_3_0_U112 ( .A(npu_inst_pe_1_3_0_n57), .ZN(
        npu_inst_pe_1_3_0_n108) );
  AOI22_X1 npu_inst_pe_1_3_0_U111 ( .A1(npu_inst_int_data_y_4__0__0_), .A2(
        npu_inst_pe_1_3_0_n54), .B1(npu_inst_pe_1_3_0_n118), .B2(
        npu_inst_pe_1_3_0_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_3_0_n53) );
  INV_X1 npu_inst_pe_1_3_0_U110 ( .A(npu_inst_pe_1_3_0_n53), .ZN(
        npu_inst_pe_1_3_0_n109) );
  AOI22_X1 npu_inst_pe_1_3_0_U107 ( .A1(npu_inst_int_data_y_4__0__0_), .A2(
        npu_inst_pe_1_3_0_n50), .B1(npu_inst_pe_1_3_0_n117), .B2(
        npu_inst_pe_1_3_0_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_3_0_n49) );
  INV_X1 npu_inst_pe_1_3_0_U106 ( .A(npu_inst_pe_1_3_0_n49), .ZN(
        npu_inst_pe_1_3_0_n110) );
  AOI22_X1 npu_inst_pe_1_3_0_U105 ( .A1(npu_inst_int_data_y_4__0__0_), .A2(
        npu_inst_pe_1_3_0_n46), .B1(npu_inst_pe_1_3_0_n116), .B2(
        npu_inst_pe_1_3_0_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_3_0_n45) );
  INV_X1 npu_inst_pe_1_3_0_U104 ( .A(npu_inst_pe_1_3_0_n45), .ZN(
        npu_inst_pe_1_3_0_n111) );
  AOI22_X1 npu_inst_pe_1_3_0_U103 ( .A1(npu_inst_int_data_y_4__0__0_), .A2(
        npu_inst_pe_1_3_0_n42), .B1(npu_inst_pe_1_3_0_n115), .B2(
        npu_inst_pe_1_3_0_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_3_0_n41) );
  INV_X1 npu_inst_pe_1_3_0_U102 ( .A(npu_inst_pe_1_3_0_n41), .ZN(
        npu_inst_pe_1_3_0_n112) );
  AOI22_X1 npu_inst_pe_1_3_0_U101 ( .A1(npu_inst_int_data_y_4__0__1_), .A2(
        npu_inst_pe_1_3_0_n58), .B1(npu_inst_pe_1_3_0_n119), .B2(
        npu_inst_pe_1_3_0_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_3_0_n59) );
  INV_X1 npu_inst_pe_1_3_0_U100 ( .A(npu_inst_pe_1_3_0_n59), .ZN(
        npu_inst_pe_1_3_0_n102) );
  AOI22_X1 npu_inst_pe_1_3_0_U99 ( .A1(npu_inst_int_data_y_4__0__1_), .A2(
        npu_inst_pe_1_3_0_n54), .B1(npu_inst_pe_1_3_0_n118), .B2(
        npu_inst_pe_1_3_0_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_3_0_n55) );
  INV_X1 npu_inst_pe_1_3_0_U98 ( .A(npu_inst_pe_1_3_0_n55), .ZN(
        npu_inst_pe_1_3_0_n103) );
  AOI22_X1 npu_inst_pe_1_3_0_U97 ( .A1(npu_inst_int_data_y_4__0__1_), .A2(
        npu_inst_pe_1_3_0_n50), .B1(npu_inst_pe_1_3_0_n117), .B2(
        npu_inst_pe_1_3_0_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_3_0_n51) );
  INV_X1 npu_inst_pe_1_3_0_U96 ( .A(npu_inst_pe_1_3_0_n51), .ZN(
        npu_inst_pe_1_3_0_n104) );
  AOI22_X1 npu_inst_pe_1_3_0_U95 ( .A1(npu_inst_int_data_y_4__0__1_), .A2(
        npu_inst_pe_1_3_0_n46), .B1(npu_inst_pe_1_3_0_n116), .B2(
        npu_inst_pe_1_3_0_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_3_0_n47) );
  INV_X1 npu_inst_pe_1_3_0_U94 ( .A(npu_inst_pe_1_3_0_n47), .ZN(
        npu_inst_pe_1_3_0_n105) );
  AOI22_X1 npu_inst_pe_1_3_0_U93 ( .A1(npu_inst_int_data_y_4__0__1_), .A2(
        npu_inst_pe_1_3_0_n42), .B1(npu_inst_pe_1_3_0_n115), .B2(
        npu_inst_pe_1_3_0_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_3_0_n43) );
  INV_X1 npu_inst_pe_1_3_0_U92 ( .A(npu_inst_pe_1_3_0_n43), .ZN(
        npu_inst_pe_1_3_0_n106) );
  AOI22_X1 npu_inst_pe_1_3_0_U91 ( .A1(npu_inst_pe_1_3_0_n38), .A2(
        npu_inst_int_data_y_4__0__1_), .B1(npu_inst_pe_1_3_0_n114), .B2(
        npu_inst_pe_1_3_0_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_3_0_n39) );
  INV_X1 npu_inst_pe_1_3_0_U90 ( .A(npu_inst_pe_1_3_0_n39), .ZN(
        npu_inst_pe_1_3_0_n107) );
  AOI22_X1 npu_inst_pe_1_3_0_U89 ( .A1(npu_inst_pe_1_3_0_n38), .A2(
        npu_inst_int_data_y_4__0__0_), .B1(npu_inst_pe_1_3_0_n114), .B2(
        npu_inst_pe_1_3_0_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_3_0_n37) );
  INV_X1 npu_inst_pe_1_3_0_U88 ( .A(npu_inst_pe_1_3_0_n37), .ZN(
        npu_inst_pe_1_3_0_n113) );
  NAND2_X1 npu_inst_pe_1_3_0_U87 ( .A1(npu_inst_pe_1_3_0_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_3_0_n60), .ZN(npu_inst_pe_1_3_0_n74) );
  OAI21_X1 npu_inst_pe_1_3_0_U86 ( .B1(npu_inst_pe_1_3_0_n63), .B2(
        npu_inst_pe_1_3_0_n60), .A(npu_inst_pe_1_3_0_n74), .ZN(
        npu_inst_pe_1_3_0_n97) );
  NAND2_X1 npu_inst_pe_1_3_0_U85 ( .A1(npu_inst_pe_1_3_0_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_3_0_n60), .ZN(npu_inst_pe_1_3_0_n73) );
  OAI21_X1 npu_inst_pe_1_3_0_U84 ( .B1(npu_inst_pe_1_3_0_n61), .B2(
        npu_inst_pe_1_3_0_n60), .A(npu_inst_pe_1_3_0_n73), .ZN(
        npu_inst_pe_1_3_0_n96) );
  NAND2_X1 npu_inst_pe_1_3_0_U83 ( .A1(npu_inst_pe_1_3_0_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_3_0_n56), .ZN(npu_inst_pe_1_3_0_n72) );
  OAI21_X1 npu_inst_pe_1_3_0_U82 ( .B1(npu_inst_pe_1_3_0_n63), .B2(
        npu_inst_pe_1_3_0_n56), .A(npu_inst_pe_1_3_0_n72), .ZN(
        npu_inst_pe_1_3_0_n95) );
  NAND2_X1 npu_inst_pe_1_3_0_U81 ( .A1(npu_inst_pe_1_3_0_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_3_0_n56), .ZN(npu_inst_pe_1_3_0_n71) );
  OAI21_X1 npu_inst_pe_1_3_0_U80 ( .B1(npu_inst_pe_1_3_0_n61), .B2(
        npu_inst_pe_1_3_0_n56), .A(npu_inst_pe_1_3_0_n71), .ZN(
        npu_inst_pe_1_3_0_n94) );
  NAND2_X1 npu_inst_pe_1_3_0_U79 ( .A1(npu_inst_pe_1_3_0_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_3_0_n52), .ZN(npu_inst_pe_1_3_0_n70) );
  OAI21_X1 npu_inst_pe_1_3_0_U78 ( .B1(npu_inst_pe_1_3_0_n63), .B2(
        npu_inst_pe_1_3_0_n52), .A(npu_inst_pe_1_3_0_n70), .ZN(
        npu_inst_pe_1_3_0_n93) );
  NAND2_X1 npu_inst_pe_1_3_0_U77 ( .A1(npu_inst_pe_1_3_0_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_3_0_n52), .ZN(npu_inst_pe_1_3_0_n69) );
  OAI21_X1 npu_inst_pe_1_3_0_U76 ( .B1(npu_inst_pe_1_3_0_n61), .B2(
        npu_inst_pe_1_3_0_n52), .A(npu_inst_pe_1_3_0_n69), .ZN(
        npu_inst_pe_1_3_0_n92) );
  NAND2_X1 npu_inst_pe_1_3_0_U75 ( .A1(npu_inst_pe_1_3_0_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_3_0_n48), .ZN(npu_inst_pe_1_3_0_n68) );
  OAI21_X1 npu_inst_pe_1_3_0_U74 ( .B1(npu_inst_pe_1_3_0_n63), .B2(
        npu_inst_pe_1_3_0_n48), .A(npu_inst_pe_1_3_0_n68), .ZN(
        npu_inst_pe_1_3_0_n91) );
  NAND2_X1 npu_inst_pe_1_3_0_U73 ( .A1(npu_inst_pe_1_3_0_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_3_0_n48), .ZN(npu_inst_pe_1_3_0_n67) );
  OAI21_X1 npu_inst_pe_1_3_0_U72 ( .B1(npu_inst_pe_1_3_0_n61), .B2(
        npu_inst_pe_1_3_0_n48), .A(npu_inst_pe_1_3_0_n67), .ZN(
        npu_inst_pe_1_3_0_n90) );
  NAND2_X1 npu_inst_pe_1_3_0_U71 ( .A1(npu_inst_pe_1_3_0_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_3_0_n44), .ZN(npu_inst_pe_1_3_0_n66) );
  OAI21_X1 npu_inst_pe_1_3_0_U70 ( .B1(npu_inst_pe_1_3_0_n63), .B2(
        npu_inst_pe_1_3_0_n44), .A(npu_inst_pe_1_3_0_n66), .ZN(
        npu_inst_pe_1_3_0_n89) );
  NAND2_X1 npu_inst_pe_1_3_0_U69 ( .A1(npu_inst_pe_1_3_0_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_3_0_n44), .ZN(npu_inst_pe_1_3_0_n65) );
  OAI21_X1 npu_inst_pe_1_3_0_U68 ( .B1(npu_inst_pe_1_3_0_n61), .B2(
        npu_inst_pe_1_3_0_n44), .A(npu_inst_pe_1_3_0_n65), .ZN(
        npu_inst_pe_1_3_0_n88) );
  NAND2_X1 npu_inst_pe_1_3_0_U67 ( .A1(npu_inst_pe_1_3_0_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_3_0_n40), .ZN(npu_inst_pe_1_3_0_n64) );
  OAI21_X1 npu_inst_pe_1_3_0_U66 ( .B1(npu_inst_pe_1_3_0_n63), .B2(
        npu_inst_pe_1_3_0_n40), .A(npu_inst_pe_1_3_0_n64), .ZN(
        npu_inst_pe_1_3_0_n87) );
  NAND2_X1 npu_inst_pe_1_3_0_U65 ( .A1(npu_inst_pe_1_3_0_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_3_0_n40), .ZN(npu_inst_pe_1_3_0_n62) );
  OAI21_X1 npu_inst_pe_1_3_0_U64 ( .B1(npu_inst_pe_1_3_0_n61), .B2(
        npu_inst_pe_1_3_0_n40), .A(npu_inst_pe_1_3_0_n62), .ZN(
        npu_inst_pe_1_3_0_n86) );
  AND2_X1 npu_inst_pe_1_3_0_U63 ( .A1(npu_inst_pe_1_3_0_N93), .A2(npu_inst_n57), .ZN(npu_inst_int_data_y_3__0__0_) );
  AND2_X1 npu_inst_pe_1_3_0_U62 ( .A1(npu_inst_n57), .A2(npu_inst_pe_1_3_0_N94), .ZN(npu_inst_int_data_y_3__0__1_) );
  NOR3_X1 npu_inst_pe_1_3_0_U61 ( .A1(npu_inst_pe_1_3_0_n26), .A2(npu_inst_n57), .A3(npu_inst_int_ckg[39]), .ZN(npu_inst_pe_1_3_0_n85) );
  OR2_X1 npu_inst_pe_1_3_0_U60 ( .A1(npu_inst_pe_1_3_0_n85), .A2(
        npu_inst_pe_1_3_0_n2), .ZN(npu_inst_pe_1_3_0_N84) );
  AND2_X1 npu_inst_pe_1_3_0_U59 ( .A1(npu_inst_pe_1_3_0_int_q_acc_0_), .A2(
        npu_inst_pe_1_3_0_n1), .ZN(npu_inst_int_data_res_3__0__0_) );
  AND2_X1 npu_inst_pe_1_3_0_U58 ( .A1(npu_inst_pe_1_3_0_n2), .A2(
        npu_inst_pe_1_3_0_int_q_acc_7_), .ZN(npu_inst_int_data_res_3__0__7_)
         );
  AND2_X1 npu_inst_pe_1_3_0_U57 ( .A1(npu_inst_pe_1_3_0_int_q_acc_1_), .A2(
        npu_inst_pe_1_3_0_n1), .ZN(npu_inst_int_data_res_3__0__1_) );
  AND2_X1 npu_inst_pe_1_3_0_U56 ( .A1(npu_inst_pe_1_3_0_int_q_acc_2_), .A2(
        npu_inst_pe_1_3_0_n1), .ZN(npu_inst_int_data_res_3__0__2_) );
  AND2_X1 npu_inst_pe_1_3_0_U55 ( .A1(npu_inst_pe_1_3_0_int_q_acc_3_), .A2(
        npu_inst_pe_1_3_0_n2), .ZN(npu_inst_int_data_res_3__0__3_) );
  AND2_X1 npu_inst_pe_1_3_0_U54 ( .A1(npu_inst_pe_1_3_0_int_q_acc_4_), .A2(
        npu_inst_pe_1_3_0_n2), .ZN(npu_inst_int_data_res_3__0__4_) );
  AND2_X1 npu_inst_pe_1_3_0_U53 ( .A1(npu_inst_pe_1_3_0_int_q_acc_5_), .A2(
        npu_inst_pe_1_3_0_n2), .ZN(npu_inst_int_data_res_3__0__5_) );
  AND2_X1 npu_inst_pe_1_3_0_U52 ( .A1(npu_inst_pe_1_3_0_int_q_acc_6_), .A2(
        npu_inst_pe_1_3_0_n2), .ZN(npu_inst_int_data_res_3__0__6_) );
  AOI222_X1 npu_inst_pe_1_3_0_U51 ( .A1(npu_inst_int_data_res_4__0__0_), .A2(
        npu_inst_pe_1_3_0_n1), .B1(npu_inst_pe_1_3_0_N73), .B2(
        npu_inst_pe_1_3_0_n76), .C1(npu_inst_pe_1_3_0_N65), .C2(
        npu_inst_pe_1_3_0_n77), .ZN(npu_inst_pe_1_3_0_n84) );
  INV_X1 npu_inst_pe_1_3_0_U50 ( .A(npu_inst_pe_1_3_0_n84), .ZN(
        npu_inst_pe_1_3_0_n101) );
  AOI222_X1 npu_inst_pe_1_3_0_U49 ( .A1(npu_inst_int_data_res_4__0__7_), .A2(
        npu_inst_pe_1_3_0_n1), .B1(npu_inst_pe_1_3_0_N80), .B2(
        npu_inst_pe_1_3_0_n76), .C1(npu_inst_pe_1_3_0_N72), .C2(
        npu_inst_pe_1_3_0_n77), .ZN(npu_inst_pe_1_3_0_n75) );
  INV_X1 npu_inst_pe_1_3_0_U48 ( .A(npu_inst_pe_1_3_0_n75), .ZN(
        npu_inst_pe_1_3_0_n33) );
  AOI222_X1 npu_inst_pe_1_3_0_U47 ( .A1(npu_inst_int_data_res_4__0__1_), .A2(
        npu_inst_pe_1_3_0_n1), .B1(npu_inst_pe_1_3_0_N74), .B2(
        npu_inst_pe_1_3_0_n76), .C1(npu_inst_pe_1_3_0_N66), .C2(
        npu_inst_pe_1_3_0_n77), .ZN(npu_inst_pe_1_3_0_n83) );
  INV_X1 npu_inst_pe_1_3_0_U46 ( .A(npu_inst_pe_1_3_0_n83), .ZN(
        npu_inst_pe_1_3_0_n100) );
  AOI222_X1 npu_inst_pe_1_3_0_U45 ( .A1(npu_inst_int_data_res_4__0__2_), .A2(
        npu_inst_pe_1_3_0_n1), .B1(npu_inst_pe_1_3_0_N75), .B2(
        npu_inst_pe_1_3_0_n76), .C1(npu_inst_pe_1_3_0_N67), .C2(
        npu_inst_pe_1_3_0_n77), .ZN(npu_inst_pe_1_3_0_n82) );
  INV_X1 npu_inst_pe_1_3_0_U44 ( .A(npu_inst_pe_1_3_0_n82), .ZN(
        npu_inst_pe_1_3_0_n99) );
  AOI222_X1 npu_inst_pe_1_3_0_U43 ( .A1(npu_inst_int_data_res_4__0__3_), .A2(
        npu_inst_pe_1_3_0_n1), .B1(npu_inst_pe_1_3_0_N76), .B2(
        npu_inst_pe_1_3_0_n76), .C1(npu_inst_pe_1_3_0_N68), .C2(
        npu_inst_pe_1_3_0_n77), .ZN(npu_inst_pe_1_3_0_n81) );
  INV_X1 npu_inst_pe_1_3_0_U42 ( .A(npu_inst_pe_1_3_0_n81), .ZN(
        npu_inst_pe_1_3_0_n98) );
  AOI222_X1 npu_inst_pe_1_3_0_U41 ( .A1(npu_inst_int_data_res_4__0__4_), .A2(
        npu_inst_pe_1_3_0_n1), .B1(npu_inst_pe_1_3_0_N77), .B2(
        npu_inst_pe_1_3_0_n76), .C1(npu_inst_pe_1_3_0_N69), .C2(
        npu_inst_pe_1_3_0_n77), .ZN(npu_inst_pe_1_3_0_n80) );
  INV_X1 npu_inst_pe_1_3_0_U40 ( .A(npu_inst_pe_1_3_0_n80), .ZN(
        npu_inst_pe_1_3_0_n36) );
  AOI222_X1 npu_inst_pe_1_3_0_U39 ( .A1(npu_inst_int_data_res_4__0__5_), .A2(
        npu_inst_pe_1_3_0_n1), .B1(npu_inst_pe_1_3_0_N78), .B2(
        npu_inst_pe_1_3_0_n76), .C1(npu_inst_pe_1_3_0_N70), .C2(
        npu_inst_pe_1_3_0_n77), .ZN(npu_inst_pe_1_3_0_n79) );
  INV_X1 npu_inst_pe_1_3_0_U38 ( .A(npu_inst_pe_1_3_0_n79), .ZN(
        npu_inst_pe_1_3_0_n35) );
  AOI222_X1 npu_inst_pe_1_3_0_U37 ( .A1(npu_inst_int_data_res_4__0__6_), .A2(
        npu_inst_pe_1_3_0_n1), .B1(npu_inst_pe_1_3_0_N79), .B2(
        npu_inst_pe_1_3_0_n76), .C1(npu_inst_pe_1_3_0_N71), .C2(
        npu_inst_pe_1_3_0_n77), .ZN(npu_inst_pe_1_3_0_n78) );
  INV_X1 npu_inst_pe_1_3_0_U36 ( .A(npu_inst_pe_1_3_0_n78), .ZN(
        npu_inst_pe_1_3_0_n34) );
  AND2_X1 npu_inst_pe_1_3_0_U35 ( .A1(npu_inst_pe_1_3_0_o_data_h_1_), .A2(
        npu_inst_pe_1_3_0_int_q_weight_1_), .ZN(npu_inst_pe_1_3_0_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_3_0_U34 ( .A1(npu_inst_pe_1_3_0_o_data_h_0_), .A2(
        npu_inst_pe_1_3_0_int_q_weight_1_), .ZN(npu_inst_pe_1_3_0_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_3_0_U33 ( .A(npu_inst_pe_1_3_0_int_data_1_), .ZN(
        npu_inst_pe_1_3_0_n14) );
  AOI22_X1 npu_inst_pe_1_3_0_U32 ( .A1(npu_inst_n57), .A2(
        npu_inst_int_data_y_4__0__1_), .B1(npu_inst_pe_1_3_0_n3), .B2(
        npu_inst_int_data_x_3__1__1_), .ZN(npu_inst_pe_1_3_0_n63) );
  AOI22_X1 npu_inst_pe_1_3_0_U31 ( .A1(npu_inst_n57), .A2(
        npu_inst_int_data_y_4__0__0_), .B1(npu_inst_pe_1_3_0_n3), .B2(
        npu_inst_int_data_x_3__1__0_), .ZN(npu_inst_pe_1_3_0_n61) );
  INV_X1 npu_inst_pe_1_3_0_U30 ( .A(npu_inst_pe_1_3_0_int_data_0_), .ZN(
        npu_inst_pe_1_3_0_n13) );
  INV_X1 npu_inst_pe_1_3_0_U29 ( .A(npu_inst_n70), .ZN(npu_inst_pe_1_3_0_n5)
         );
  OR3_X1 npu_inst_pe_1_3_0_U28 ( .A1(npu_inst_pe_1_3_0_n6), .A2(
        npu_inst_pe_1_3_0_n8), .A3(npu_inst_pe_1_3_0_n5), .ZN(
        npu_inst_pe_1_3_0_n56) );
  OR3_X1 npu_inst_pe_1_3_0_U27 ( .A1(npu_inst_pe_1_3_0_n5), .A2(
        npu_inst_pe_1_3_0_n8), .A3(npu_inst_pe_1_3_0_n7), .ZN(
        npu_inst_pe_1_3_0_n48) );
  INV_X1 npu_inst_pe_1_3_0_U26 ( .A(npu_inst_pe_1_3_0_n5), .ZN(
        npu_inst_pe_1_3_0_n4) );
  OR3_X1 npu_inst_pe_1_3_0_U25 ( .A1(npu_inst_pe_1_3_0_n4), .A2(
        npu_inst_pe_1_3_0_n8), .A3(npu_inst_pe_1_3_0_n7), .ZN(
        npu_inst_pe_1_3_0_n52) );
  OR3_X1 npu_inst_pe_1_3_0_U24 ( .A1(npu_inst_pe_1_3_0_n6), .A2(
        npu_inst_pe_1_3_0_n8), .A3(npu_inst_pe_1_3_0_n4), .ZN(
        npu_inst_pe_1_3_0_n60) );
  NOR2_X1 npu_inst_pe_1_3_0_U23 ( .A1(npu_inst_pe_1_3_0_n60), .A2(
        npu_inst_pe_1_3_0_n3), .ZN(npu_inst_pe_1_3_0_n58) );
  NOR2_X1 npu_inst_pe_1_3_0_U22 ( .A1(npu_inst_pe_1_3_0_n56), .A2(
        npu_inst_pe_1_3_0_n3), .ZN(npu_inst_pe_1_3_0_n54) );
  NOR2_X1 npu_inst_pe_1_3_0_U21 ( .A1(npu_inst_pe_1_3_0_n52), .A2(
        npu_inst_pe_1_3_0_n3), .ZN(npu_inst_pe_1_3_0_n50) );
  NOR2_X1 npu_inst_pe_1_3_0_U20 ( .A1(npu_inst_pe_1_3_0_n48), .A2(
        npu_inst_pe_1_3_0_n3), .ZN(npu_inst_pe_1_3_0_n46) );
  NOR2_X1 npu_inst_pe_1_3_0_U19 ( .A1(npu_inst_pe_1_3_0_n40), .A2(
        npu_inst_pe_1_3_0_n3), .ZN(npu_inst_pe_1_3_0_n38) );
  NOR2_X1 npu_inst_pe_1_3_0_U18 ( .A1(npu_inst_pe_1_3_0_n44), .A2(
        npu_inst_pe_1_3_0_n3), .ZN(npu_inst_pe_1_3_0_n42) );
  BUF_X1 npu_inst_pe_1_3_0_U17 ( .A(npu_inst_n101), .Z(npu_inst_pe_1_3_0_n8)
         );
  INV_X1 npu_inst_pe_1_3_0_U16 ( .A(npu_inst_n125), .ZN(npu_inst_pe_1_3_0_n12)
         );
  INV_X1 npu_inst_pe_1_3_0_U15 ( .A(npu_inst_pe_1_3_0_n38), .ZN(
        npu_inst_pe_1_3_0_n114) );
  INV_X1 npu_inst_pe_1_3_0_U14 ( .A(npu_inst_pe_1_3_0_n58), .ZN(
        npu_inst_pe_1_3_0_n119) );
  INV_X1 npu_inst_pe_1_3_0_U13 ( .A(npu_inst_pe_1_3_0_n54), .ZN(
        npu_inst_pe_1_3_0_n118) );
  INV_X1 npu_inst_pe_1_3_0_U12 ( .A(npu_inst_pe_1_3_0_n50), .ZN(
        npu_inst_pe_1_3_0_n117) );
  INV_X1 npu_inst_pe_1_3_0_U11 ( .A(npu_inst_pe_1_3_0_n46), .ZN(
        npu_inst_pe_1_3_0_n116) );
  INV_X1 npu_inst_pe_1_3_0_U10 ( .A(npu_inst_pe_1_3_0_n42), .ZN(
        npu_inst_pe_1_3_0_n115) );
  BUF_X1 npu_inst_pe_1_3_0_U9 ( .A(npu_inst_n26), .Z(npu_inst_pe_1_3_0_n2) );
  BUF_X1 npu_inst_pe_1_3_0_U8 ( .A(npu_inst_n26), .Z(npu_inst_pe_1_3_0_n1) );
  BUF_X1 npu_inst_pe_1_3_0_U7 ( .A(npu_inst_pe_1_3_0_n12), .Z(
        npu_inst_pe_1_3_0_n11) );
  BUF_X1 npu_inst_pe_1_3_0_U6 ( .A(npu_inst_pe_1_3_0_n12), .Z(
        npu_inst_pe_1_3_0_n10) );
  BUF_X1 npu_inst_pe_1_3_0_U5 ( .A(npu_inst_pe_1_3_0_n12), .Z(
        npu_inst_pe_1_3_0_n9) );
  NOR2_X1 npu_inst_pe_1_3_0_U4 ( .A1(npu_inst_pe_1_3_0_int_q_weight_0_), .A2(
        npu_inst_pe_1_3_0_n1), .ZN(npu_inst_pe_1_3_0_n76) );
  NOR2_X1 npu_inst_pe_1_3_0_U3 ( .A1(npu_inst_pe_1_3_0_n27), .A2(
        npu_inst_pe_1_3_0_n1), .ZN(npu_inst_pe_1_3_0_n77) );
  FA_X1 npu_inst_pe_1_3_0_sub_67_U2_1 ( .A(npu_inst_pe_1_3_0_int_q_acc_1_), 
        .B(npu_inst_pe_1_3_0_n14), .CI(npu_inst_pe_1_3_0_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_3_0_sub_67_carry_2_), .S(npu_inst_pe_1_3_0_N66) );
  FA_X1 npu_inst_pe_1_3_0_add_69_U1_1 ( .A(npu_inst_pe_1_3_0_int_q_acc_1_), 
        .B(npu_inst_pe_1_3_0_int_data_1_), .CI(
        npu_inst_pe_1_3_0_add_69_carry_1_), .CO(
        npu_inst_pe_1_3_0_add_69_carry_2_), .S(npu_inst_pe_1_3_0_N74) );
  NAND3_X1 npu_inst_pe_1_3_0_U109 ( .A1(npu_inst_pe_1_3_0_n5), .A2(
        npu_inst_pe_1_3_0_n7), .A3(npu_inst_pe_1_3_0_n8), .ZN(
        npu_inst_pe_1_3_0_n44) );
  NAND3_X1 npu_inst_pe_1_3_0_U108 ( .A1(npu_inst_pe_1_3_0_n4), .A2(
        npu_inst_pe_1_3_0_n7), .A3(npu_inst_pe_1_3_0_n8), .ZN(
        npu_inst_pe_1_3_0_n40) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_3_0_n34), .CK(
        npu_inst_pe_1_3_0_net4010), .RN(npu_inst_pe_1_3_0_n9), .Q(
        npu_inst_pe_1_3_0_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_3_0_n35), .CK(
        npu_inst_pe_1_3_0_net4010), .RN(npu_inst_pe_1_3_0_n9), .Q(
        npu_inst_pe_1_3_0_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_3_0_n36), .CK(
        npu_inst_pe_1_3_0_net4010), .RN(npu_inst_pe_1_3_0_n9), .Q(
        npu_inst_pe_1_3_0_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_3_0_n98), .CK(
        npu_inst_pe_1_3_0_net4010), .RN(npu_inst_pe_1_3_0_n9), .Q(
        npu_inst_pe_1_3_0_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_3_0_n99), .CK(
        npu_inst_pe_1_3_0_net4010), .RN(npu_inst_pe_1_3_0_n9), .Q(
        npu_inst_pe_1_3_0_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_3_0_n100), 
        .CK(npu_inst_pe_1_3_0_net4010), .RN(npu_inst_pe_1_3_0_n9), .Q(
        npu_inst_pe_1_3_0_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_3_0_n33), .CK(
        npu_inst_pe_1_3_0_net4010), .RN(npu_inst_pe_1_3_0_n9), .Q(
        npu_inst_pe_1_3_0_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_3_0_n101), 
        .CK(npu_inst_pe_1_3_0_net4010), .RN(npu_inst_pe_1_3_0_n9), .Q(
        npu_inst_pe_1_3_0_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_weight_reg_0_ ( .D(npu_inst_n111), .CK(
        npu_inst_pe_1_3_0_net4016), .RN(npu_inst_pe_1_3_0_n9), .Q(
        npu_inst_pe_1_3_0_int_q_weight_0_), .QN(npu_inst_pe_1_3_0_n27) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_weight_reg_1_ ( .D(npu_inst_n117), .CK(
        npu_inst_pe_1_3_0_net4016), .RN(npu_inst_pe_1_3_0_n9), .Q(
        npu_inst_pe_1_3_0_int_q_weight_1_), .QN(npu_inst_pe_1_3_0_n26) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_3_0_n113), 
        .CK(npu_inst_pe_1_3_0_net4016), .RN(npu_inst_pe_1_3_0_n9), .Q(
        npu_inst_pe_1_3_0_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_3_0_n107), 
        .CK(npu_inst_pe_1_3_0_net4016), .RN(npu_inst_pe_1_3_0_n9), .Q(
        npu_inst_pe_1_3_0_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_3_0_n112), 
        .CK(npu_inst_pe_1_3_0_net4016), .RN(npu_inst_pe_1_3_0_n10), .Q(
        npu_inst_pe_1_3_0_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_3_0_n106), 
        .CK(npu_inst_pe_1_3_0_net4016), .RN(npu_inst_pe_1_3_0_n10), .Q(
        npu_inst_pe_1_3_0_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_3_0_n111), 
        .CK(npu_inst_pe_1_3_0_net4016), .RN(npu_inst_pe_1_3_0_n10), .Q(
        npu_inst_pe_1_3_0_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_3_0_n105), 
        .CK(npu_inst_pe_1_3_0_net4016), .RN(npu_inst_pe_1_3_0_n10), .Q(
        npu_inst_pe_1_3_0_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_3_0_n110), 
        .CK(npu_inst_pe_1_3_0_net4016), .RN(npu_inst_pe_1_3_0_n10), .Q(
        npu_inst_pe_1_3_0_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_3_0_n104), 
        .CK(npu_inst_pe_1_3_0_net4016), .RN(npu_inst_pe_1_3_0_n10), .Q(
        npu_inst_pe_1_3_0_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_3_0_n109), 
        .CK(npu_inst_pe_1_3_0_net4016), .RN(npu_inst_pe_1_3_0_n10), .Q(
        npu_inst_pe_1_3_0_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_3_0_n103), 
        .CK(npu_inst_pe_1_3_0_net4016), .RN(npu_inst_pe_1_3_0_n10), .Q(
        npu_inst_pe_1_3_0_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_3_0_n108), 
        .CK(npu_inst_pe_1_3_0_net4016), .RN(npu_inst_pe_1_3_0_n10), .Q(
        npu_inst_pe_1_3_0_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_3_0_n102), 
        .CK(npu_inst_pe_1_3_0_net4016), .RN(npu_inst_pe_1_3_0_n10), .Q(
        npu_inst_pe_1_3_0_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_3_0_n86), 
        .CK(npu_inst_pe_1_3_0_net4016), .RN(npu_inst_pe_1_3_0_n10), .Q(
        npu_inst_pe_1_3_0_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_3_0_n87), 
        .CK(npu_inst_pe_1_3_0_net4016), .RN(npu_inst_pe_1_3_0_n10), .Q(
        npu_inst_pe_1_3_0_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_3_0_n88), 
        .CK(npu_inst_pe_1_3_0_net4016), .RN(npu_inst_pe_1_3_0_n11), .Q(
        npu_inst_pe_1_3_0_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_3_0_n89), 
        .CK(npu_inst_pe_1_3_0_net4016), .RN(npu_inst_pe_1_3_0_n11), .Q(
        npu_inst_pe_1_3_0_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_3_0_n90), 
        .CK(npu_inst_pe_1_3_0_net4016), .RN(npu_inst_pe_1_3_0_n11), .Q(
        npu_inst_pe_1_3_0_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_3_0_n91), 
        .CK(npu_inst_pe_1_3_0_net4016), .RN(npu_inst_pe_1_3_0_n11), .Q(
        npu_inst_pe_1_3_0_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_3_0_n92), 
        .CK(npu_inst_pe_1_3_0_net4016), .RN(npu_inst_pe_1_3_0_n11), .Q(
        npu_inst_pe_1_3_0_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_3_0_n93), 
        .CK(npu_inst_pe_1_3_0_net4016), .RN(npu_inst_pe_1_3_0_n11), .Q(
        npu_inst_pe_1_3_0_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_3_0_n94), 
        .CK(npu_inst_pe_1_3_0_net4016), .RN(npu_inst_pe_1_3_0_n11), .Q(
        npu_inst_pe_1_3_0_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_3_0_n95), 
        .CK(npu_inst_pe_1_3_0_net4016), .RN(npu_inst_pe_1_3_0_n11), .Q(
        npu_inst_pe_1_3_0_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_3_0_n96), 
        .CK(npu_inst_pe_1_3_0_net4016), .RN(npu_inst_pe_1_3_0_n11), .Q(
        npu_inst_pe_1_3_0_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_3_0_n97), 
        .CK(npu_inst_pe_1_3_0_net4016), .RN(npu_inst_pe_1_3_0_n11), .Q(
        npu_inst_pe_1_3_0_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_3_0_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_3_0_N84), .SE(1'b0), .GCK(npu_inst_pe_1_3_0_net4010) );
  CLKGATETST_X1 npu_inst_pe_1_3_0_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n64), .SE(1'b0), .GCK(npu_inst_pe_1_3_0_net4016) );
  MUX2_X1 npu_inst_pe_1_3_1_U162 ( .A(npu_inst_pe_1_3_1_n32), .B(
        npu_inst_pe_1_3_1_n29), .S(npu_inst_pe_1_3_1_n8), .Z(
        npu_inst_pe_1_3_1_N93) );
  MUX2_X1 npu_inst_pe_1_3_1_U161 ( .A(npu_inst_pe_1_3_1_n31), .B(
        npu_inst_pe_1_3_1_n30), .S(npu_inst_pe_1_3_1_n6), .Z(
        npu_inst_pe_1_3_1_n32) );
  MUX2_X1 npu_inst_pe_1_3_1_U160 ( .A(npu_inst_pe_1_3_1_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_3_1_int_q_reg_v_1__0_), .S(npu_inst_pe_1_3_1_n4), .Z(
        npu_inst_pe_1_3_1_n31) );
  MUX2_X1 npu_inst_pe_1_3_1_U159 ( .A(npu_inst_pe_1_3_1_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_3_1_int_q_reg_v_3__0_), .S(npu_inst_pe_1_3_1_n4), .Z(
        npu_inst_pe_1_3_1_n30) );
  MUX2_X1 npu_inst_pe_1_3_1_U158 ( .A(npu_inst_pe_1_3_1_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_3_1_int_q_reg_v_5__0_), .S(npu_inst_pe_1_3_1_n4), .Z(
        npu_inst_pe_1_3_1_n29) );
  MUX2_X1 npu_inst_pe_1_3_1_U157 ( .A(npu_inst_pe_1_3_1_n28), .B(
        npu_inst_pe_1_3_1_n23), .S(npu_inst_pe_1_3_1_n8), .Z(
        npu_inst_pe_1_3_1_N94) );
  MUX2_X1 npu_inst_pe_1_3_1_U156 ( .A(npu_inst_pe_1_3_1_n25), .B(
        npu_inst_pe_1_3_1_n24), .S(npu_inst_pe_1_3_1_n6), .Z(
        npu_inst_pe_1_3_1_n28) );
  MUX2_X1 npu_inst_pe_1_3_1_U155 ( .A(npu_inst_pe_1_3_1_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_3_1_int_q_reg_v_1__1_), .S(npu_inst_pe_1_3_1_n4), .Z(
        npu_inst_pe_1_3_1_n25) );
  MUX2_X1 npu_inst_pe_1_3_1_U154 ( .A(npu_inst_pe_1_3_1_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_3_1_int_q_reg_v_3__1_), .S(npu_inst_pe_1_3_1_n4), .Z(
        npu_inst_pe_1_3_1_n24) );
  MUX2_X1 npu_inst_pe_1_3_1_U153 ( .A(npu_inst_pe_1_3_1_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_3_1_int_q_reg_v_5__1_), .S(npu_inst_pe_1_3_1_n4), .Z(
        npu_inst_pe_1_3_1_n23) );
  MUX2_X1 npu_inst_pe_1_3_1_U152 ( .A(npu_inst_pe_1_3_1_n22), .B(
        npu_inst_pe_1_3_1_n19), .S(npu_inst_pe_1_3_1_n8), .Z(
        npu_inst_int_data_x_3__1__1_) );
  MUX2_X1 npu_inst_pe_1_3_1_U151 ( .A(npu_inst_pe_1_3_1_n21), .B(
        npu_inst_pe_1_3_1_n20), .S(npu_inst_pe_1_3_1_n6), .Z(
        npu_inst_pe_1_3_1_n22) );
  MUX2_X1 npu_inst_pe_1_3_1_U150 ( .A(npu_inst_pe_1_3_1_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_3_1_int_q_reg_h_1__1_), .S(npu_inst_pe_1_3_1_n4), .Z(
        npu_inst_pe_1_3_1_n21) );
  MUX2_X1 npu_inst_pe_1_3_1_U149 ( .A(npu_inst_pe_1_3_1_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_3_1_int_q_reg_h_3__1_), .S(npu_inst_pe_1_3_1_n4), .Z(
        npu_inst_pe_1_3_1_n20) );
  MUX2_X1 npu_inst_pe_1_3_1_U148 ( .A(npu_inst_pe_1_3_1_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_3_1_int_q_reg_h_5__1_), .S(npu_inst_pe_1_3_1_n4), .Z(
        npu_inst_pe_1_3_1_n19) );
  MUX2_X1 npu_inst_pe_1_3_1_U147 ( .A(npu_inst_pe_1_3_1_n18), .B(
        npu_inst_pe_1_3_1_n15), .S(npu_inst_pe_1_3_1_n8), .Z(
        npu_inst_int_data_x_3__1__0_) );
  MUX2_X1 npu_inst_pe_1_3_1_U146 ( .A(npu_inst_pe_1_3_1_n17), .B(
        npu_inst_pe_1_3_1_n16), .S(npu_inst_pe_1_3_1_n6), .Z(
        npu_inst_pe_1_3_1_n18) );
  MUX2_X1 npu_inst_pe_1_3_1_U145 ( .A(npu_inst_pe_1_3_1_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_3_1_int_q_reg_h_1__0_), .S(npu_inst_pe_1_3_1_n4), .Z(
        npu_inst_pe_1_3_1_n17) );
  MUX2_X1 npu_inst_pe_1_3_1_U144 ( .A(npu_inst_pe_1_3_1_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_3_1_int_q_reg_h_3__0_), .S(npu_inst_pe_1_3_1_n4), .Z(
        npu_inst_pe_1_3_1_n16) );
  MUX2_X1 npu_inst_pe_1_3_1_U143 ( .A(npu_inst_pe_1_3_1_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_3_1_int_q_reg_h_5__0_), .S(npu_inst_pe_1_3_1_n4), .Z(
        npu_inst_pe_1_3_1_n15) );
  XOR2_X1 npu_inst_pe_1_3_1_U142 ( .A(npu_inst_pe_1_3_1_int_data_0_), .B(
        npu_inst_pe_1_3_1_int_q_acc_0_), .Z(npu_inst_pe_1_3_1_N73) );
  AND2_X1 npu_inst_pe_1_3_1_U141 ( .A1(npu_inst_pe_1_3_1_int_q_acc_0_), .A2(
        npu_inst_pe_1_3_1_int_data_0_), .ZN(npu_inst_pe_1_3_1_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_3_1_U140 ( .A(npu_inst_pe_1_3_1_int_q_acc_0_), .B(
        npu_inst_pe_1_3_1_n13), .ZN(npu_inst_pe_1_3_1_N65) );
  OR2_X1 npu_inst_pe_1_3_1_U139 ( .A1(npu_inst_pe_1_3_1_n13), .A2(
        npu_inst_pe_1_3_1_int_q_acc_0_), .ZN(npu_inst_pe_1_3_1_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_3_1_U138 ( .A(npu_inst_pe_1_3_1_int_q_acc_2_), .B(
        npu_inst_pe_1_3_1_add_69_carry_2_), .Z(npu_inst_pe_1_3_1_N75) );
  AND2_X1 npu_inst_pe_1_3_1_U137 ( .A1(npu_inst_pe_1_3_1_add_69_carry_2_), 
        .A2(npu_inst_pe_1_3_1_int_q_acc_2_), .ZN(
        npu_inst_pe_1_3_1_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_3_1_U136 ( .A(npu_inst_pe_1_3_1_int_q_acc_3_), .B(
        npu_inst_pe_1_3_1_add_69_carry_3_), .Z(npu_inst_pe_1_3_1_N76) );
  AND2_X1 npu_inst_pe_1_3_1_U135 ( .A1(npu_inst_pe_1_3_1_add_69_carry_3_), 
        .A2(npu_inst_pe_1_3_1_int_q_acc_3_), .ZN(
        npu_inst_pe_1_3_1_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_3_1_U134 ( .A(npu_inst_pe_1_3_1_int_q_acc_4_), .B(
        npu_inst_pe_1_3_1_add_69_carry_4_), .Z(npu_inst_pe_1_3_1_N77) );
  AND2_X1 npu_inst_pe_1_3_1_U133 ( .A1(npu_inst_pe_1_3_1_add_69_carry_4_), 
        .A2(npu_inst_pe_1_3_1_int_q_acc_4_), .ZN(
        npu_inst_pe_1_3_1_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_3_1_U132 ( .A(npu_inst_pe_1_3_1_int_q_acc_5_), .B(
        npu_inst_pe_1_3_1_add_69_carry_5_), .Z(npu_inst_pe_1_3_1_N78) );
  AND2_X1 npu_inst_pe_1_3_1_U131 ( .A1(npu_inst_pe_1_3_1_add_69_carry_5_), 
        .A2(npu_inst_pe_1_3_1_int_q_acc_5_), .ZN(
        npu_inst_pe_1_3_1_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_3_1_U130 ( .A(npu_inst_pe_1_3_1_int_q_acc_6_), .B(
        npu_inst_pe_1_3_1_add_69_carry_6_), .Z(npu_inst_pe_1_3_1_N79) );
  AND2_X1 npu_inst_pe_1_3_1_U129 ( .A1(npu_inst_pe_1_3_1_add_69_carry_6_), 
        .A2(npu_inst_pe_1_3_1_int_q_acc_6_), .ZN(
        npu_inst_pe_1_3_1_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_3_1_U128 ( .A(npu_inst_pe_1_3_1_int_q_acc_7_), .B(
        npu_inst_pe_1_3_1_add_69_carry_7_), .Z(npu_inst_pe_1_3_1_N80) );
  XNOR2_X1 npu_inst_pe_1_3_1_U127 ( .A(npu_inst_pe_1_3_1_sub_67_carry_2_), .B(
        npu_inst_pe_1_3_1_int_q_acc_2_), .ZN(npu_inst_pe_1_3_1_N67) );
  OR2_X1 npu_inst_pe_1_3_1_U126 ( .A1(npu_inst_pe_1_3_1_int_q_acc_2_), .A2(
        npu_inst_pe_1_3_1_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_3_1_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_3_1_U125 ( .A(npu_inst_pe_1_3_1_sub_67_carry_3_), .B(
        npu_inst_pe_1_3_1_int_q_acc_3_), .ZN(npu_inst_pe_1_3_1_N68) );
  OR2_X1 npu_inst_pe_1_3_1_U124 ( .A1(npu_inst_pe_1_3_1_int_q_acc_3_), .A2(
        npu_inst_pe_1_3_1_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_3_1_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_3_1_U123 ( .A(npu_inst_pe_1_3_1_sub_67_carry_4_), .B(
        npu_inst_pe_1_3_1_int_q_acc_4_), .ZN(npu_inst_pe_1_3_1_N69) );
  OR2_X1 npu_inst_pe_1_3_1_U122 ( .A1(npu_inst_pe_1_3_1_int_q_acc_4_), .A2(
        npu_inst_pe_1_3_1_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_3_1_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_3_1_U121 ( .A(npu_inst_pe_1_3_1_sub_67_carry_5_), .B(
        npu_inst_pe_1_3_1_int_q_acc_5_), .ZN(npu_inst_pe_1_3_1_N70) );
  OR2_X1 npu_inst_pe_1_3_1_U120 ( .A1(npu_inst_pe_1_3_1_int_q_acc_5_), .A2(
        npu_inst_pe_1_3_1_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_3_1_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_3_1_U119 ( .A(npu_inst_pe_1_3_1_sub_67_carry_6_), .B(
        npu_inst_pe_1_3_1_int_q_acc_6_), .ZN(npu_inst_pe_1_3_1_N71) );
  OR2_X1 npu_inst_pe_1_3_1_U118 ( .A1(npu_inst_pe_1_3_1_int_q_acc_6_), .A2(
        npu_inst_pe_1_3_1_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_3_1_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_3_1_U117 ( .A(npu_inst_pe_1_3_1_int_q_acc_7_), .B(
        npu_inst_pe_1_3_1_sub_67_carry_7_), .ZN(npu_inst_pe_1_3_1_N72) );
  INV_X1 npu_inst_pe_1_3_1_U116 ( .A(npu_inst_n78), .ZN(npu_inst_pe_1_3_1_n7)
         );
  INV_X1 npu_inst_pe_1_3_1_U115 ( .A(npu_inst_pe_1_3_1_n7), .ZN(
        npu_inst_pe_1_3_1_n6) );
  INV_X1 npu_inst_pe_1_3_1_U114 ( .A(npu_inst_n57), .ZN(npu_inst_pe_1_3_1_n3)
         );
  AOI22_X1 npu_inst_pe_1_3_1_U113 ( .A1(npu_inst_int_data_y_4__1__0_), .A2(
        npu_inst_pe_1_3_1_n58), .B1(npu_inst_pe_1_3_1_n119), .B2(
        npu_inst_pe_1_3_1_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_3_1_n57) );
  INV_X1 npu_inst_pe_1_3_1_U112 ( .A(npu_inst_pe_1_3_1_n57), .ZN(
        npu_inst_pe_1_3_1_n108) );
  AOI22_X1 npu_inst_pe_1_3_1_U111 ( .A1(npu_inst_int_data_y_4__1__0_), .A2(
        npu_inst_pe_1_3_1_n54), .B1(npu_inst_pe_1_3_1_n118), .B2(
        npu_inst_pe_1_3_1_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_3_1_n53) );
  INV_X1 npu_inst_pe_1_3_1_U110 ( .A(npu_inst_pe_1_3_1_n53), .ZN(
        npu_inst_pe_1_3_1_n109) );
  AOI22_X1 npu_inst_pe_1_3_1_U107 ( .A1(npu_inst_int_data_y_4__1__0_), .A2(
        npu_inst_pe_1_3_1_n50), .B1(npu_inst_pe_1_3_1_n117), .B2(
        npu_inst_pe_1_3_1_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_3_1_n49) );
  INV_X1 npu_inst_pe_1_3_1_U106 ( .A(npu_inst_pe_1_3_1_n49), .ZN(
        npu_inst_pe_1_3_1_n110) );
  AOI22_X1 npu_inst_pe_1_3_1_U105 ( .A1(npu_inst_int_data_y_4__1__0_), .A2(
        npu_inst_pe_1_3_1_n46), .B1(npu_inst_pe_1_3_1_n116), .B2(
        npu_inst_pe_1_3_1_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_3_1_n45) );
  INV_X1 npu_inst_pe_1_3_1_U104 ( .A(npu_inst_pe_1_3_1_n45), .ZN(
        npu_inst_pe_1_3_1_n111) );
  AOI22_X1 npu_inst_pe_1_3_1_U103 ( .A1(npu_inst_int_data_y_4__1__0_), .A2(
        npu_inst_pe_1_3_1_n42), .B1(npu_inst_pe_1_3_1_n115), .B2(
        npu_inst_pe_1_3_1_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_3_1_n41) );
  INV_X1 npu_inst_pe_1_3_1_U102 ( .A(npu_inst_pe_1_3_1_n41), .ZN(
        npu_inst_pe_1_3_1_n112) );
  AOI22_X1 npu_inst_pe_1_3_1_U101 ( .A1(npu_inst_int_data_y_4__1__1_), .A2(
        npu_inst_pe_1_3_1_n58), .B1(npu_inst_pe_1_3_1_n119), .B2(
        npu_inst_pe_1_3_1_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_3_1_n59) );
  INV_X1 npu_inst_pe_1_3_1_U100 ( .A(npu_inst_pe_1_3_1_n59), .ZN(
        npu_inst_pe_1_3_1_n102) );
  AOI22_X1 npu_inst_pe_1_3_1_U99 ( .A1(npu_inst_int_data_y_4__1__1_), .A2(
        npu_inst_pe_1_3_1_n54), .B1(npu_inst_pe_1_3_1_n118), .B2(
        npu_inst_pe_1_3_1_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_3_1_n55) );
  INV_X1 npu_inst_pe_1_3_1_U98 ( .A(npu_inst_pe_1_3_1_n55), .ZN(
        npu_inst_pe_1_3_1_n103) );
  AOI22_X1 npu_inst_pe_1_3_1_U97 ( .A1(npu_inst_int_data_y_4__1__1_), .A2(
        npu_inst_pe_1_3_1_n50), .B1(npu_inst_pe_1_3_1_n117), .B2(
        npu_inst_pe_1_3_1_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_3_1_n51) );
  INV_X1 npu_inst_pe_1_3_1_U96 ( .A(npu_inst_pe_1_3_1_n51), .ZN(
        npu_inst_pe_1_3_1_n104) );
  AOI22_X1 npu_inst_pe_1_3_1_U95 ( .A1(npu_inst_int_data_y_4__1__1_), .A2(
        npu_inst_pe_1_3_1_n46), .B1(npu_inst_pe_1_3_1_n116), .B2(
        npu_inst_pe_1_3_1_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_3_1_n47) );
  INV_X1 npu_inst_pe_1_3_1_U94 ( .A(npu_inst_pe_1_3_1_n47), .ZN(
        npu_inst_pe_1_3_1_n105) );
  AOI22_X1 npu_inst_pe_1_3_1_U93 ( .A1(npu_inst_int_data_y_4__1__1_), .A2(
        npu_inst_pe_1_3_1_n42), .B1(npu_inst_pe_1_3_1_n115), .B2(
        npu_inst_pe_1_3_1_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_3_1_n43) );
  INV_X1 npu_inst_pe_1_3_1_U92 ( .A(npu_inst_pe_1_3_1_n43), .ZN(
        npu_inst_pe_1_3_1_n106) );
  AOI22_X1 npu_inst_pe_1_3_1_U91 ( .A1(npu_inst_pe_1_3_1_n38), .A2(
        npu_inst_int_data_y_4__1__1_), .B1(npu_inst_pe_1_3_1_n114), .B2(
        npu_inst_pe_1_3_1_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_3_1_n39) );
  INV_X1 npu_inst_pe_1_3_1_U90 ( .A(npu_inst_pe_1_3_1_n39), .ZN(
        npu_inst_pe_1_3_1_n107) );
  AOI22_X1 npu_inst_pe_1_3_1_U89 ( .A1(npu_inst_pe_1_3_1_n38), .A2(
        npu_inst_int_data_y_4__1__0_), .B1(npu_inst_pe_1_3_1_n114), .B2(
        npu_inst_pe_1_3_1_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_3_1_n37) );
  INV_X1 npu_inst_pe_1_3_1_U88 ( .A(npu_inst_pe_1_3_1_n37), .ZN(
        npu_inst_pe_1_3_1_n113) );
  NAND2_X1 npu_inst_pe_1_3_1_U87 ( .A1(npu_inst_pe_1_3_1_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_3_1_n60), .ZN(npu_inst_pe_1_3_1_n74) );
  OAI21_X1 npu_inst_pe_1_3_1_U86 ( .B1(npu_inst_pe_1_3_1_n63), .B2(
        npu_inst_pe_1_3_1_n60), .A(npu_inst_pe_1_3_1_n74), .ZN(
        npu_inst_pe_1_3_1_n97) );
  NAND2_X1 npu_inst_pe_1_3_1_U85 ( .A1(npu_inst_pe_1_3_1_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_3_1_n60), .ZN(npu_inst_pe_1_3_1_n73) );
  OAI21_X1 npu_inst_pe_1_3_1_U84 ( .B1(npu_inst_pe_1_3_1_n61), .B2(
        npu_inst_pe_1_3_1_n60), .A(npu_inst_pe_1_3_1_n73), .ZN(
        npu_inst_pe_1_3_1_n96) );
  NAND2_X1 npu_inst_pe_1_3_1_U83 ( .A1(npu_inst_pe_1_3_1_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_3_1_n56), .ZN(npu_inst_pe_1_3_1_n72) );
  OAI21_X1 npu_inst_pe_1_3_1_U82 ( .B1(npu_inst_pe_1_3_1_n63), .B2(
        npu_inst_pe_1_3_1_n56), .A(npu_inst_pe_1_3_1_n72), .ZN(
        npu_inst_pe_1_3_1_n95) );
  NAND2_X1 npu_inst_pe_1_3_1_U81 ( .A1(npu_inst_pe_1_3_1_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_3_1_n56), .ZN(npu_inst_pe_1_3_1_n71) );
  OAI21_X1 npu_inst_pe_1_3_1_U80 ( .B1(npu_inst_pe_1_3_1_n61), .B2(
        npu_inst_pe_1_3_1_n56), .A(npu_inst_pe_1_3_1_n71), .ZN(
        npu_inst_pe_1_3_1_n94) );
  NAND2_X1 npu_inst_pe_1_3_1_U79 ( .A1(npu_inst_pe_1_3_1_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_3_1_n52), .ZN(npu_inst_pe_1_3_1_n70) );
  OAI21_X1 npu_inst_pe_1_3_1_U78 ( .B1(npu_inst_pe_1_3_1_n63), .B2(
        npu_inst_pe_1_3_1_n52), .A(npu_inst_pe_1_3_1_n70), .ZN(
        npu_inst_pe_1_3_1_n93) );
  NAND2_X1 npu_inst_pe_1_3_1_U77 ( .A1(npu_inst_pe_1_3_1_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_3_1_n52), .ZN(npu_inst_pe_1_3_1_n69) );
  OAI21_X1 npu_inst_pe_1_3_1_U76 ( .B1(npu_inst_pe_1_3_1_n61), .B2(
        npu_inst_pe_1_3_1_n52), .A(npu_inst_pe_1_3_1_n69), .ZN(
        npu_inst_pe_1_3_1_n92) );
  NAND2_X1 npu_inst_pe_1_3_1_U75 ( .A1(npu_inst_pe_1_3_1_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_3_1_n48), .ZN(npu_inst_pe_1_3_1_n68) );
  OAI21_X1 npu_inst_pe_1_3_1_U74 ( .B1(npu_inst_pe_1_3_1_n63), .B2(
        npu_inst_pe_1_3_1_n48), .A(npu_inst_pe_1_3_1_n68), .ZN(
        npu_inst_pe_1_3_1_n91) );
  NAND2_X1 npu_inst_pe_1_3_1_U73 ( .A1(npu_inst_pe_1_3_1_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_3_1_n48), .ZN(npu_inst_pe_1_3_1_n67) );
  OAI21_X1 npu_inst_pe_1_3_1_U72 ( .B1(npu_inst_pe_1_3_1_n61), .B2(
        npu_inst_pe_1_3_1_n48), .A(npu_inst_pe_1_3_1_n67), .ZN(
        npu_inst_pe_1_3_1_n90) );
  NAND2_X1 npu_inst_pe_1_3_1_U71 ( .A1(npu_inst_pe_1_3_1_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_3_1_n44), .ZN(npu_inst_pe_1_3_1_n66) );
  OAI21_X1 npu_inst_pe_1_3_1_U70 ( .B1(npu_inst_pe_1_3_1_n63), .B2(
        npu_inst_pe_1_3_1_n44), .A(npu_inst_pe_1_3_1_n66), .ZN(
        npu_inst_pe_1_3_1_n89) );
  NAND2_X1 npu_inst_pe_1_3_1_U69 ( .A1(npu_inst_pe_1_3_1_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_3_1_n44), .ZN(npu_inst_pe_1_3_1_n65) );
  OAI21_X1 npu_inst_pe_1_3_1_U68 ( .B1(npu_inst_pe_1_3_1_n61), .B2(
        npu_inst_pe_1_3_1_n44), .A(npu_inst_pe_1_3_1_n65), .ZN(
        npu_inst_pe_1_3_1_n88) );
  NAND2_X1 npu_inst_pe_1_3_1_U67 ( .A1(npu_inst_pe_1_3_1_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_3_1_n40), .ZN(npu_inst_pe_1_3_1_n64) );
  OAI21_X1 npu_inst_pe_1_3_1_U66 ( .B1(npu_inst_pe_1_3_1_n63), .B2(
        npu_inst_pe_1_3_1_n40), .A(npu_inst_pe_1_3_1_n64), .ZN(
        npu_inst_pe_1_3_1_n87) );
  NAND2_X1 npu_inst_pe_1_3_1_U65 ( .A1(npu_inst_pe_1_3_1_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_3_1_n40), .ZN(npu_inst_pe_1_3_1_n62) );
  OAI21_X1 npu_inst_pe_1_3_1_U64 ( .B1(npu_inst_pe_1_3_1_n61), .B2(
        npu_inst_pe_1_3_1_n40), .A(npu_inst_pe_1_3_1_n62), .ZN(
        npu_inst_pe_1_3_1_n86) );
  AND2_X1 npu_inst_pe_1_3_1_U63 ( .A1(npu_inst_pe_1_3_1_N93), .A2(npu_inst_n57), .ZN(npu_inst_int_data_y_3__1__0_) );
  AND2_X1 npu_inst_pe_1_3_1_U62 ( .A1(npu_inst_n57), .A2(npu_inst_pe_1_3_1_N94), .ZN(npu_inst_int_data_y_3__1__1_) );
  NOR3_X1 npu_inst_pe_1_3_1_U61 ( .A1(npu_inst_pe_1_3_1_n26), .A2(npu_inst_n57), .A3(npu_inst_int_ckg[38]), .ZN(npu_inst_pe_1_3_1_n85) );
  OR2_X1 npu_inst_pe_1_3_1_U60 ( .A1(npu_inst_pe_1_3_1_n85), .A2(
        npu_inst_pe_1_3_1_n2), .ZN(npu_inst_pe_1_3_1_N84) );
  AND2_X1 npu_inst_pe_1_3_1_U59 ( .A1(npu_inst_pe_1_3_1_int_q_acc_0_), .A2(
        npu_inst_pe_1_3_1_n1), .ZN(npu_inst_int_data_res_3__1__0_) );
  AND2_X1 npu_inst_pe_1_3_1_U58 ( .A1(npu_inst_pe_1_3_1_n2), .A2(
        npu_inst_pe_1_3_1_int_q_acc_7_), .ZN(npu_inst_int_data_res_3__1__7_)
         );
  AND2_X1 npu_inst_pe_1_3_1_U57 ( .A1(npu_inst_pe_1_3_1_int_q_acc_1_), .A2(
        npu_inst_pe_1_3_1_n1), .ZN(npu_inst_int_data_res_3__1__1_) );
  AND2_X1 npu_inst_pe_1_3_1_U56 ( .A1(npu_inst_pe_1_3_1_int_q_acc_2_), .A2(
        npu_inst_pe_1_3_1_n1), .ZN(npu_inst_int_data_res_3__1__2_) );
  AND2_X1 npu_inst_pe_1_3_1_U55 ( .A1(npu_inst_pe_1_3_1_int_q_acc_3_), .A2(
        npu_inst_pe_1_3_1_n2), .ZN(npu_inst_int_data_res_3__1__3_) );
  AND2_X1 npu_inst_pe_1_3_1_U54 ( .A1(npu_inst_pe_1_3_1_int_q_acc_4_), .A2(
        npu_inst_pe_1_3_1_n2), .ZN(npu_inst_int_data_res_3__1__4_) );
  AND2_X1 npu_inst_pe_1_3_1_U53 ( .A1(npu_inst_pe_1_3_1_int_q_acc_5_), .A2(
        npu_inst_pe_1_3_1_n2), .ZN(npu_inst_int_data_res_3__1__5_) );
  AND2_X1 npu_inst_pe_1_3_1_U52 ( .A1(npu_inst_pe_1_3_1_int_q_acc_6_), .A2(
        npu_inst_pe_1_3_1_n2), .ZN(npu_inst_int_data_res_3__1__6_) );
  AOI222_X1 npu_inst_pe_1_3_1_U51 ( .A1(npu_inst_int_data_res_4__1__0_), .A2(
        npu_inst_pe_1_3_1_n1), .B1(npu_inst_pe_1_3_1_N73), .B2(
        npu_inst_pe_1_3_1_n76), .C1(npu_inst_pe_1_3_1_N65), .C2(
        npu_inst_pe_1_3_1_n77), .ZN(npu_inst_pe_1_3_1_n84) );
  INV_X1 npu_inst_pe_1_3_1_U50 ( .A(npu_inst_pe_1_3_1_n84), .ZN(
        npu_inst_pe_1_3_1_n101) );
  AOI222_X1 npu_inst_pe_1_3_1_U49 ( .A1(npu_inst_int_data_res_4__1__7_), .A2(
        npu_inst_pe_1_3_1_n1), .B1(npu_inst_pe_1_3_1_N80), .B2(
        npu_inst_pe_1_3_1_n76), .C1(npu_inst_pe_1_3_1_N72), .C2(
        npu_inst_pe_1_3_1_n77), .ZN(npu_inst_pe_1_3_1_n75) );
  INV_X1 npu_inst_pe_1_3_1_U48 ( .A(npu_inst_pe_1_3_1_n75), .ZN(
        npu_inst_pe_1_3_1_n33) );
  AOI222_X1 npu_inst_pe_1_3_1_U47 ( .A1(npu_inst_int_data_res_4__1__1_), .A2(
        npu_inst_pe_1_3_1_n1), .B1(npu_inst_pe_1_3_1_N74), .B2(
        npu_inst_pe_1_3_1_n76), .C1(npu_inst_pe_1_3_1_N66), .C2(
        npu_inst_pe_1_3_1_n77), .ZN(npu_inst_pe_1_3_1_n83) );
  INV_X1 npu_inst_pe_1_3_1_U46 ( .A(npu_inst_pe_1_3_1_n83), .ZN(
        npu_inst_pe_1_3_1_n100) );
  AOI222_X1 npu_inst_pe_1_3_1_U45 ( .A1(npu_inst_int_data_res_4__1__2_), .A2(
        npu_inst_pe_1_3_1_n1), .B1(npu_inst_pe_1_3_1_N75), .B2(
        npu_inst_pe_1_3_1_n76), .C1(npu_inst_pe_1_3_1_N67), .C2(
        npu_inst_pe_1_3_1_n77), .ZN(npu_inst_pe_1_3_1_n82) );
  INV_X1 npu_inst_pe_1_3_1_U44 ( .A(npu_inst_pe_1_3_1_n82), .ZN(
        npu_inst_pe_1_3_1_n99) );
  AOI222_X1 npu_inst_pe_1_3_1_U43 ( .A1(npu_inst_int_data_res_4__1__3_), .A2(
        npu_inst_pe_1_3_1_n1), .B1(npu_inst_pe_1_3_1_N76), .B2(
        npu_inst_pe_1_3_1_n76), .C1(npu_inst_pe_1_3_1_N68), .C2(
        npu_inst_pe_1_3_1_n77), .ZN(npu_inst_pe_1_3_1_n81) );
  INV_X1 npu_inst_pe_1_3_1_U42 ( .A(npu_inst_pe_1_3_1_n81), .ZN(
        npu_inst_pe_1_3_1_n98) );
  AOI222_X1 npu_inst_pe_1_3_1_U41 ( .A1(npu_inst_int_data_res_4__1__4_), .A2(
        npu_inst_pe_1_3_1_n1), .B1(npu_inst_pe_1_3_1_N77), .B2(
        npu_inst_pe_1_3_1_n76), .C1(npu_inst_pe_1_3_1_N69), .C2(
        npu_inst_pe_1_3_1_n77), .ZN(npu_inst_pe_1_3_1_n80) );
  INV_X1 npu_inst_pe_1_3_1_U40 ( .A(npu_inst_pe_1_3_1_n80), .ZN(
        npu_inst_pe_1_3_1_n36) );
  AOI222_X1 npu_inst_pe_1_3_1_U39 ( .A1(npu_inst_int_data_res_4__1__5_), .A2(
        npu_inst_pe_1_3_1_n1), .B1(npu_inst_pe_1_3_1_N78), .B2(
        npu_inst_pe_1_3_1_n76), .C1(npu_inst_pe_1_3_1_N70), .C2(
        npu_inst_pe_1_3_1_n77), .ZN(npu_inst_pe_1_3_1_n79) );
  INV_X1 npu_inst_pe_1_3_1_U38 ( .A(npu_inst_pe_1_3_1_n79), .ZN(
        npu_inst_pe_1_3_1_n35) );
  AOI222_X1 npu_inst_pe_1_3_1_U37 ( .A1(npu_inst_int_data_res_4__1__6_), .A2(
        npu_inst_pe_1_3_1_n1), .B1(npu_inst_pe_1_3_1_N79), .B2(
        npu_inst_pe_1_3_1_n76), .C1(npu_inst_pe_1_3_1_N71), .C2(
        npu_inst_pe_1_3_1_n77), .ZN(npu_inst_pe_1_3_1_n78) );
  INV_X1 npu_inst_pe_1_3_1_U36 ( .A(npu_inst_pe_1_3_1_n78), .ZN(
        npu_inst_pe_1_3_1_n34) );
  INV_X1 npu_inst_pe_1_3_1_U35 ( .A(npu_inst_pe_1_3_1_int_data_1_), .ZN(
        npu_inst_pe_1_3_1_n14) );
  AND2_X1 npu_inst_pe_1_3_1_U34 ( .A1(npu_inst_int_data_x_3__1__1_), .A2(
        npu_inst_pe_1_3_1_int_q_weight_1_), .ZN(npu_inst_pe_1_3_1_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_3_1_U33 ( .A1(npu_inst_int_data_x_3__1__0_), .A2(
        npu_inst_pe_1_3_1_int_q_weight_1_), .ZN(npu_inst_pe_1_3_1_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_3_1_U32 ( .A1(npu_inst_n57), .A2(
        npu_inst_int_data_y_4__1__1_), .B1(npu_inst_pe_1_3_1_n3), .B2(
        npu_inst_int_data_x_3__2__1_), .ZN(npu_inst_pe_1_3_1_n63) );
  AOI22_X1 npu_inst_pe_1_3_1_U31 ( .A1(npu_inst_n57), .A2(
        npu_inst_int_data_y_4__1__0_), .B1(npu_inst_pe_1_3_1_n3), .B2(
        npu_inst_int_data_x_3__2__0_), .ZN(npu_inst_pe_1_3_1_n61) );
  INV_X1 npu_inst_pe_1_3_1_U30 ( .A(npu_inst_pe_1_3_1_int_data_0_), .ZN(
        npu_inst_pe_1_3_1_n13) );
  INV_X1 npu_inst_pe_1_3_1_U29 ( .A(npu_inst_n70), .ZN(npu_inst_pe_1_3_1_n5)
         );
  OR3_X1 npu_inst_pe_1_3_1_U28 ( .A1(npu_inst_pe_1_3_1_n6), .A2(
        npu_inst_pe_1_3_1_n8), .A3(npu_inst_pe_1_3_1_n5), .ZN(
        npu_inst_pe_1_3_1_n56) );
  OR3_X1 npu_inst_pe_1_3_1_U27 ( .A1(npu_inst_pe_1_3_1_n5), .A2(
        npu_inst_pe_1_3_1_n8), .A3(npu_inst_pe_1_3_1_n7), .ZN(
        npu_inst_pe_1_3_1_n48) );
  INV_X1 npu_inst_pe_1_3_1_U26 ( .A(npu_inst_pe_1_3_1_n5), .ZN(
        npu_inst_pe_1_3_1_n4) );
  OR3_X1 npu_inst_pe_1_3_1_U25 ( .A1(npu_inst_pe_1_3_1_n4), .A2(
        npu_inst_pe_1_3_1_n8), .A3(npu_inst_pe_1_3_1_n7), .ZN(
        npu_inst_pe_1_3_1_n52) );
  OR3_X1 npu_inst_pe_1_3_1_U24 ( .A1(npu_inst_pe_1_3_1_n6), .A2(
        npu_inst_pe_1_3_1_n8), .A3(npu_inst_pe_1_3_1_n4), .ZN(
        npu_inst_pe_1_3_1_n60) );
  NOR2_X1 npu_inst_pe_1_3_1_U23 ( .A1(npu_inst_pe_1_3_1_n60), .A2(
        npu_inst_pe_1_3_1_n3), .ZN(npu_inst_pe_1_3_1_n58) );
  NOR2_X1 npu_inst_pe_1_3_1_U22 ( .A1(npu_inst_pe_1_3_1_n56), .A2(
        npu_inst_pe_1_3_1_n3), .ZN(npu_inst_pe_1_3_1_n54) );
  NOR2_X1 npu_inst_pe_1_3_1_U21 ( .A1(npu_inst_pe_1_3_1_n52), .A2(
        npu_inst_pe_1_3_1_n3), .ZN(npu_inst_pe_1_3_1_n50) );
  NOR2_X1 npu_inst_pe_1_3_1_U20 ( .A1(npu_inst_pe_1_3_1_n48), .A2(
        npu_inst_pe_1_3_1_n3), .ZN(npu_inst_pe_1_3_1_n46) );
  NOR2_X1 npu_inst_pe_1_3_1_U19 ( .A1(npu_inst_pe_1_3_1_n40), .A2(
        npu_inst_pe_1_3_1_n3), .ZN(npu_inst_pe_1_3_1_n38) );
  NOR2_X1 npu_inst_pe_1_3_1_U18 ( .A1(npu_inst_pe_1_3_1_n44), .A2(
        npu_inst_pe_1_3_1_n3), .ZN(npu_inst_pe_1_3_1_n42) );
  BUF_X1 npu_inst_pe_1_3_1_U17 ( .A(npu_inst_n101), .Z(npu_inst_pe_1_3_1_n8)
         );
  INV_X1 npu_inst_pe_1_3_1_U16 ( .A(npu_inst_n125), .ZN(npu_inst_pe_1_3_1_n12)
         );
  INV_X1 npu_inst_pe_1_3_1_U15 ( .A(npu_inst_pe_1_3_1_n38), .ZN(
        npu_inst_pe_1_3_1_n114) );
  INV_X1 npu_inst_pe_1_3_1_U14 ( .A(npu_inst_pe_1_3_1_n58), .ZN(
        npu_inst_pe_1_3_1_n119) );
  INV_X1 npu_inst_pe_1_3_1_U13 ( .A(npu_inst_pe_1_3_1_n54), .ZN(
        npu_inst_pe_1_3_1_n118) );
  INV_X1 npu_inst_pe_1_3_1_U12 ( .A(npu_inst_pe_1_3_1_n50), .ZN(
        npu_inst_pe_1_3_1_n117) );
  INV_X1 npu_inst_pe_1_3_1_U11 ( .A(npu_inst_pe_1_3_1_n46), .ZN(
        npu_inst_pe_1_3_1_n116) );
  INV_X1 npu_inst_pe_1_3_1_U10 ( .A(npu_inst_pe_1_3_1_n42), .ZN(
        npu_inst_pe_1_3_1_n115) );
  BUF_X1 npu_inst_pe_1_3_1_U9 ( .A(npu_inst_n26), .Z(npu_inst_pe_1_3_1_n2) );
  BUF_X1 npu_inst_pe_1_3_1_U8 ( .A(npu_inst_n26), .Z(npu_inst_pe_1_3_1_n1) );
  BUF_X1 npu_inst_pe_1_3_1_U7 ( .A(npu_inst_pe_1_3_1_n12), .Z(
        npu_inst_pe_1_3_1_n11) );
  BUF_X1 npu_inst_pe_1_3_1_U6 ( .A(npu_inst_pe_1_3_1_n12), .Z(
        npu_inst_pe_1_3_1_n10) );
  BUF_X1 npu_inst_pe_1_3_1_U5 ( .A(npu_inst_pe_1_3_1_n12), .Z(
        npu_inst_pe_1_3_1_n9) );
  NOR2_X1 npu_inst_pe_1_3_1_U4 ( .A1(npu_inst_pe_1_3_1_int_q_weight_0_), .A2(
        npu_inst_pe_1_3_1_n1), .ZN(npu_inst_pe_1_3_1_n76) );
  NOR2_X1 npu_inst_pe_1_3_1_U3 ( .A1(npu_inst_pe_1_3_1_n27), .A2(
        npu_inst_pe_1_3_1_n1), .ZN(npu_inst_pe_1_3_1_n77) );
  FA_X1 npu_inst_pe_1_3_1_sub_67_U2_1 ( .A(npu_inst_pe_1_3_1_int_q_acc_1_), 
        .B(npu_inst_pe_1_3_1_n14), .CI(npu_inst_pe_1_3_1_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_3_1_sub_67_carry_2_), .S(npu_inst_pe_1_3_1_N66) );
  FA_X1 npu_inst_pe_1_3_1_add_69_U1_1 ( .A(npu_inst_pe_1_3_1_int_q_acc_1_), 
        .B(npu_inst_pe_1_3_1_int_data_1_), .CI(
        npu_inst_pe_1_3_1_add_69_carry_1_), .CO(
        npu_inst_pe_1_3_1_add_69_carry_2_), .S(npu_inst_pe_1_3_1_N74) );
  NAND3_X1 npu_inst_pe_1_3_1_U109 ( .A1(npu_inst_pe_1_3_1_n5), .A2(
        npu_inst_pe_1_3_1_n7), .A3(npu_inst_pe_1_3_1_n8), .ZN(
        npu_inst_pe_1_3_1_n44) );
  NAND3_X1 npu_inst_pe_1_3_1_U108 ( .A1(npu_inst_pe_1_3_1_n4), .A2(
        npu_inst_pe_1_3_1_n7), .A3(npu_inst_pe_1_3_1_n8), .ZN(
        npu_inst_pe_1_3_1_n40) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_3_1_n34), .CK(
        npu_inst_pe_1_3_1_net3987), .RN(npu_inst_pe_1_3_1_n9), .Q(
        npu_inst_pe_1_3_1_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_3_1_n35), .CK(
        npu_inst_pe_1_3_1_net3987), .RN(npu_inst_pe_1_3_1_n9), .Q(
        npu_inst_pe_1_3_1_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_3_1_n36), .CK(
        npu_inst_pe_1_3_1_net3987), .RN(npu_inst_pe_1_3_1_n9), .Q(
        npu_inst_pe_1_3_1_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_3_1_n98), .CK(
        npu_inst_pe_1_3_1_net3987), .RN(npu_inst_pe_1_3_1_n9), .Q(
        npu_inst_pe_1_3_1_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_3_1_n99), .CK(
        npu_inst_pe_1_3_1_net3987), .RN(npu_inst_pe_1_3_1_n9), .Q(
        npu_inst_pe_1_3_1_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_3_1_n100), 
        .CK(npu_inst_pe_1_3_1_net3987), .RN(npu_inst_pe_1_3_1_n9), .Q(
        npu_inst_pe_1_3_1_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_3_1_n33), .CK(
        npu_inst_pe_1_3_1_net3987), .RN(npu_inst_pe_1_3_1_n9), .Q(
        npu_inst_pe_1_3_1_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_3_1_n101), 
        .CK(npu_inst_pe_1_3_1_net3987), .RN(npu_inst_pe_1_3_1_n9), .Q(
        npu_inst_pe_1_3_1_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_weight_reg_0_ ( .D(npu_inst_n111), .CK(
        npu_inst_pe_1_3_1_net3993), .RN(npu_inst_pe_1_3_1_n9), .Q(
        npu_inst_pe_1_3_1_int_q_weight_0_), .QN(npu_inst_pe_1_3_1_n27) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_weight_reg_1_ ( .D(npu_inst_n117), .CK(
        npu_inst_pe_1_3_1_net3993), .RN(npu_inst_pe_1_3_1_n9), .Q(
        npu_inst_pe_1_3_1_int_q_weight_1_), .QN(npu_inst_pe_1_3_1_n26) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_3_1_n113), 
        .CK(npu_inst_pe_1_3_1_net3993), .RN(npu_inst_pe_1_3_1_n9), .Q(
        npu_inst_pe_1_3_1_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_3_1_n107), 
        .CK(npu_inst_pe_1_3_1_net3993), .RN(npu_inst_pe_1_3_1_n9), .Q(
        npu_inst_pe_1_3_1_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_3_1_n112), 
        .CK(npu_inst_pe_1_3_1_net3993), .RN(npu_inst_pe_1_3_1_n10), .Q(
        npu_inst_pe_1_3_1_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_3_1_n106), 
        .CK(npu_inst_pe_1_3_1_net3993), .RN(npu_inst_pe_1_3_1_n10), .Q(
        npu_inst_pe_1_3_1_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_3_1_n111), 
        .CK(npu_inst_pe_1_3_1_net3993), .RN(npu_inst_pe_1_3_1_n10), .Q(
        npu_inst_pe_1_3_1_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_3_1_n105), 
        .CK(npu_inst_pe_1_3_1_net3993), .RN(npu_inst_pe_1_3_1_n10), .Q(
        npu_inst_pe_1_3_1_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_3_1_n110), 
        .CK(npu_inst_pe_1_3_1_net3993), .RN(npu_inst_pe_1_3_1_n10), .Q(
        npu_inst_pe_1_3_1_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_3_1_n104), 
        .CK(npu_inst_pe_1_3_1_net3993), .RN(npu_inst_pe_1_3_1_n10), .Q(
        npu_inst_pe_1_3_1_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_3_1_n109), 
        .CK(npu_inst_pe_1_3_1_net3993), .RN(npu_inst_pe_1_3_1_n10), .Q(
        npu_inst_pe_1_3_1_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_3_1_n103), 
        .CK(npu_inst_pe_1_3_1_net3993), .RN(npu_inst_pe_1_3_1_n10), .Q(
        npu_inst_pe_1_3_1_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_3_1_n108), 
        .CK(npu_inst_pe_1_3_1_net3993), .RN(npu_inst_pe_1_3_1_n10), .Q(
        npu_inst_pe_1_3_1_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_3_1_n102), 
        .CK(npu_inst_pe_1_3_1_net3993), .RN(npu_inst_pe_1_3_1_n10), .Q(
        npu_inst_pe_1_3_1_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_3_1_n86), 
        .CK(npu_inst_pe_1_3_1_net3993), .RN(npu_inst_pe_1_3_1_n10), .Q(
        npu_inst_pe_1_3_1_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_3_1_n87), 
        .CK(npu_inst_pe_1_3_1_net3993), .RN(npu_inst_pe_1_3_1_n10), .Q(
        npu_inst_pe_1_3_1_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_3_1_n88), 
        .CK(npu_inst_pe_1_3_1_net3993), .RN(npu_inst_pe_1_3_1_n11), .Q(
        npu_inst_pe_1_3_1_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_3_1_n89), 
        .CK(npu_inst_pe_1_3_1_net3993), .RN(npu_inst_pe_1_3_1_n11), .Q(
        npu_inst_pe_1_3_1_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_3_1_n90), 
        .CK(npu_inst_pe_1_3_1_net3993), .RN(npu_inst_pe_1_3_1_n11), .Q(
        npu_inst_pe_1_3_1_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_3_1_n91), 
        .CK(npu_inst_pe_1_3_1_net3993), .RN(npu_inst_pe_1_3_1_n11), .Q(
        npu_inst_pe_1_3_1_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_3_1_n92), 
        .CK(npu_inst_pe_1_3_1_net3993), .RN(npu_inst_pe_1_3_1_n11), .Q(
        npu_inst_pe_1_3_1_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_3_1_n93), 
        .CK(npu_inst_pe_1_3_1_net3993), .RN(npu_inst_pe_1_3_1_n11), .Q(
        npu_inst_pe_1_3_1_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_3_1_n94), 
        .CK(npu_inst_pe_1_3_1_net3993), .RN(npu_inst_pe_1_3_1_n11), .Q(
        npu_inst_pe_1_3_1_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_3_1_n95), 
        .CK(npu_inst_pe_1_3_1_net3993), .RN(npu_inst_pe_1_3_1_n11), .Q(
        npu_inst_pe_1_3_1_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_3_1_n96), 
        .CK(npu_inst_pe_1_3_1_net3993), .RN(npu_inst_pe_1_3_1_n11), .Q(
        npu_inst_pe_1_3_1_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_3_1_n97), 
        .CK(npu_inst_pe_1_3_1_net3993), .RN(npu_inst_pe_1_3_1_n11), .Q(
        npu_inst_pe_1_3_1_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_3_1_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_3_1_N84), .SE(1'b0), .GCK(npu_inst_pe_1_3_1_net3987) );
  CLKGATETST_X1 npu_inst_pe_1_3_1_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n64), .SE(1'b0), .GCK(npu_inst_pe_1_3_1_net3993) );
  MUX2_X1 npu_inst_pe_1_3_2_U162 ( .A(npu_inst_pe_1_3_2_n32), .B(
        npu_inst_pe_1_3_2_n29), .S(npu_inst_pe_1_3_2_n8), .Z(
        npu_inst_pe_1_3_2_N93) );
  MUX2_X1 npu_inst_pe_1_3_2_U161 ( .A(npu_inst_pe_1_3_2_n31), .B(
        npu_inst_pe_1_3_2_n30), .S(npu_inst_pe_1_3_2_n6), .Z(
        npu_inst_pe_1_3_2_n32) );
  MUX2_X1 npu_inst_pe_1_3_2_U160 ( .A(npu_inst_pe_1_3_2_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_3_2_int_q_reg_v_1__0_), .S(npu_inst_pe_1_3_2_n4), .Z(
        npu_inst_pe_1_3_2_n31) );
  MUX2_X1 npu_inst_pe_1_3_2_U159 ( .A(npu_inst_pe_1_3_2_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_3_2_int_q_reg_v_3__0_), .S(npu_inst_pe_1_3_2_n4), .Z(
        npu_inst_pe_1_3_2_n30) );
  MUX2_X1 npu_inst_pe_1_3_2_U158 ( .A(npu_inst_pe_1_3_2_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_3_2_int_q_reg_v_5__0_), .S(npu_inst_pe_1_3_2_n4), .Z(
        npu_inst_pe_1_3_2_n29) );
  MUX2_X1 npu_inst_pe_1_3_2_U157 ( .A(npu_inst_pe_1_3_2_n28), .B(
        npu_inst_pe_1_3_2_n23), .S(npu_inst_pe_1_3_2_n8), .Z(
        npu_inst_pe_1_3_2_N94) );
  MUX2_X1 npu_inst_pe_1_3_2_U156 ( .A(npu_inst_pe_1_3_2_n25), .B(
        npu_inst_pe_1_3_2_n24), .S(npu_inst_pe_1_3_2_n6), .Z(
        npu_inst_pe_1_3_2_n28) );
  MUX2_X1 npu_inst_pe_1_3_2_U155 ( .A(npu_inst_pe_1_3_2_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_3_2_int_q_reg_v_1__1_), .S(npu_inst_pe_1_3_2_n4), .Z(
        npu_inst_pe_1_3_2_n25) );
  MUX2_X1 npu_inst_pe_1_3_2_U154 ( .A(npu_inst_pe_1_3_2_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_3_2_int_q_reg_v_3__1_), .S(npu_inst_pe_1_3_2_n4), .Z(
        npu_inst_pe_1_3_2_n24) );
  MUX2_X1 npu_inst_pe_1_3_2_U153 ( .A(npu_inst_pe_1_3_2_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_3_2_int_q_reg_v_5__1_), .S(npu_inst_pe_1_3_2_n4), .Z(
        npu_inst_pe_1_3_2_n23) );
  MUX2_X1 npu_inst_pe_1_3_2_U152 ( .A(npu_inst_pe_1_3_2_n22), .B(
        npu_inst_pe_1_3_2_n19), .S(npu_inst_pe_1_3_2_n8), .Z(
        npu_inst_int_data_x_3__2__1_) );
  MUX2_X1 npu_inst_pe_1_3_2_U151 ( .A(npu_inst_pe_1_3_2_n21), .B(
        npu_inst_pe_1_3_2_n20), .S(npu_inst_pe_1_3_2_n6), .Z(
        npu_inst_pe_1_3_2_n22) );
  MUX2_X1 npu_inst_pe_1_3_2_U150 ( .A(npu_inst_pe_1_3_2_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_3_2_int_q_reg_h_1__1_), .S(npu_inst_pe_1_3_2_n4), .Z(
        npu_inst_pe_1_3_2_n21) );
  MUX2_X1 npu_inst_pe_1_3_2_U149 ( .A(npu_inst_pe_1_3_2_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_3_2_int_q_reg_h_3__1_), .S(npu_inst_pe_1_3_2_n4), .Z(
        npu_inst_pe_1_3_2_n20) );
  MUX2_X1 npu_inst_pe_1_3_2_U148 ( .A(npu_inst_pe_1_3_2_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_3_2_int_q_reg_h_5__1_), .S(npu_inst_pe_1_3_2_n4), .Z(
        npu_inst_pe_1_3_2_n19) );
  MUX2_X1 npu_inst_pe_1_3_2_U147 ( .A(npu_inst_pe_1_3_2_n18), .B(
        npu_inst_pe_1_3_2_n15), .S(npu_inst_pe_1_3_2_n8), .Z(
        npu_inst_int_data_x_3__2__0_) );
  MUX2_X1 npu_inst_pe_1_3_2_U146 ( .A(npu_inst_pe_1_3_2_n17), .B(
        npu_inst_pe_1_3_2_n16), .S(npu_inst_pe_1_3_2_n6), .Z(
        npu_inst_pe_1_3_2_n18) );
  MUX2_X1 npu_inst_pe_1_3_2_U145 ( .A(npu_inst_pe_1_3_2_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_3_2_int_q_reg_h_1__0_), .S(npu_inst_pe_1_3_2_n4), .Z(
        npu_inst_pe_1_3_2_n17) );
  MUX2_X1 npu_inst_pe_1_3_2_U144 ( .A(npu_inst_pe_1_3_2_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_3_2_int_q_reg_h_3__0_), .S(npu_inst_pe_1_3_2_n4), .Z(
        npu_inst_pe_1_3_2_n16) );
  MUX2_X1 npu_inst_pe_1_3_2_U143 ( .A(npu_inst_pe_1_3_2_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_3_2_int_q_reg_h_5__0_), .S(npu_inst_pe_1_3_2_n4), .Z(
        npu_inst_pe_1_3_2_n15) );
  XOR2_X1 npu_inst_pe_1_3_2_U142 ( .A(npu_inst_pe_1_3_2_int_data_0_), .B(
        npu_inst_pe_1_3_2_int_q_acc_0_), .Z(npu_inst_pe_1_3_2_N73) );
  AND2_X1 npu_inst_pe_1_3_2_U141 ( .A1(npu_inst_pe_1_3_2_int_q_acc_0_), .A2(
        npu_inst_pe_1_3_2_int_data_0_), .ZN(npu_inst_pe_1_3_2_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_3_2_U140 ( .A(npu_inst_pe_1_3_2_int_q_acc_0_), .B(
        npu_inst_pe_1_3_2_n13), .ZN(npu_inst_pe_1_3_2_N65) );
  OR2_X1 npu_inst_pe_1_3_2_U139 ( .A1(npu_inst_pe_1_3_2_n13), .A2(
        npu_inst_pe_1_3_2_int_q_acc_0_), .ZN(npu_inst_pe_1_3_2_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_3_2_U138 ( .A(npu_inst_pe_1_3_2_int_q_acc_2_), .B(
        npu_inst_pe_1_3_2_add_69_carry_2_), .Z(npu_inst_pe_1_3_2_N75) );
  AND2_X1 npu_inst_pe_1_3_2_U137 ( .A1(npu_inst_pe_1_3_2_add_69_carry_2_), 
        .A2(npu_inst_pe_1_3_2_int_q_acc_2_), .ZN(
        npu_inst_pe_1_3_2_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_3_2_U136 ( .A(npu_inst_pe_1_3_2_int_q_acc_3_), .B(
        npu_inst_pe_1_3_2_add_69_carry_3_), .Z(npu_inst_pe_1_3_2_N76) );
  AND2_X1 npu_inst_pe_1_3_2_U135 ( .A1(npu_inst_pe_1_3_2_add_69_carry_3_), 
        .A2(npu_inst_pe_1_3_2_int_q_acc_3_), .ZN(
        npu_inst_pe_1_3_2_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_3_2_U134 ( .A(npu_inst_pe_1_3_2_int_q_acc_4_), .B(
        npu_inst_pe_1_3_2_add_69_carry_4_), .Z(npu_inst_pe_1_3_2_N77) );
  AND2_X1 npu_inst_pe_1_3_2_U133 ( .A1(npu_inst_pe_1_3_2_add_69_carry_4_), 
        .A2(npu_inst_pe_1_3_2_int_q_acc_4_), .ZN(
        npu_inst_pe_1_3_2_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_3_2_U132 ( .A(npu_inst_pe_1_3_2_int_q_acc_5_), .B(
        npu_inst_pe_1_3_2_add_69_carry_5_), .Z(npu_inst_pe_1_3_2_N78) );
  AND2_X1 npu_inst_pe_1_3_2_U131 ( .A1(npu_inst_pe_1_3_2_add_69_carry_5_), 
        .A2(npu_inst_pe_1_3_2_int_q_acc_5_), .ZN(
        npu_inst_pe_1_3_2_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_3_2_U130 ( .A(npu_inst_pe_1_3_2_int_q_acc_6_), .B(
        npu_inst_pe_1_3_2_add_69_carry_6_), .Z(npu_inst_pe_1_3_2_N79) );
  AND2_X1 npu_inst_pe_1_3_2_U129 ( .A1(npu_inst_pe_1_3_2_add_69_carry_6_), 
        .A2(npu_inst_pe_1_3_2_int_q_acc_6_), .ZN(
        npu_inst_pe_1_3_2_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_3_2_U128 ( .A(npu_inst_pe_1_3_2_int_q_acc_7_), .B(
        npu_inst_pe_1_3_2_add_69_carry_7_), .Z(npu_inst_pe_1_3_2_N80) );
  XNOR2_X1 npu_inst_pe_1_3_2_U127 ( .A(npu_inst_pe_1_3_2_sub_67_carry_2_), .B(
        npu_inst_pe_1_3_2_int_q_acc_2_), .ZN(npu_inst_pe_1_3_2_N67) );
  OR2_X1 npu_inst_pe_1_3_2_U126 ( .A1(npu_inst_pe_1_3_2_int_q_acc_2_), .A2(
        npu_inst_pe_1_3_2_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_3_2_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_3_2_U125 ( .A(npu_inst_pe_1_3_2_sub_67_carry_3_), .B(
        npu_inst_pe_1_3_2_int_q_acc_3_), .ZN(npu_inst_pe_1_3_2_N68) );
  OR2_X1 npu_inst_pe_1_3_2_U124 ( .A1(npu_inst_pe_1_3_2_int_q_acc_3_), .A2(
        npu_inst_pe_1_3_2_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_3_2_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_3_2_U123 ( .A(npu_inst_pe_1_3_2_sub_67_carry_4_), .B(
        npu_inst_pe_1_3_2_int_q_acc_4_), .ZN(npu_inst_pe_1_3_2_N69) );
  OR2_X1 npu_inst_pe_1_3_2_U122 ( .A1(npu_inst_pe_1_3_2_int_q_acc_4_), .A2(
        npu_inst_pe_1_3_2_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_3_2_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_3_2_U121 ( .A(npu_inst_pe_1_3_2_sub_67_carry_5_), .B(
        npu_inst_pe_1_3_2_int_q_acc_5_), .ZN(npu_inst_pe_1_3_2_N70) );
  OR2_X1 npu_inst_pe_1_3_2_U120 ( .A1(npu_inst_pe_1_3_2_int_q_acc_5_), .A2(
        npu_inst_pe_1_3_2_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_3_2_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_3_2_U119 ( .A(npu_inst_pe_1_3_2_sub_67_carry_6_), .B(
        npu_inst_pe_1_3_2_int_q_acc_6_), .ZN(npu_inst_pe_1_3_2_N71) );
  OR2_X1 npu_inst_pe_1_3_2_U118 ( .A1(npu_inst_pe_1_3_2_int_q_acc_6_), .A2(
        npu_inst_pe_1_3_2_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_3_2_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_3_2_U117 ( .A(npu_inst_pe_1_3_2_int_q_acc_7_), .B(
        npu_inst_pe_1_3_2_sub_67_carry_7_), .ZN(npu_inst_pe_1_3_2_N72) );
  INV_X1 npu_inst_pe_1_3_2_U116 ( .A(npu_inst_n78), .ZN(npu_inst_pe_1_3_2_n7)
         );
  INV_X1 npu_inst_pe_1_3_2_U115 ( .A(npu_inst_pe_1_3_2_n7), .ZN(
        npu_inst_pe_1_3_2_n6) );
  INV_X1 npu_inst_pe_1_3_2_U114 ( .A(npu_inst_n57), .ZN(npu_inst_pe_1_3_2_n3)
         );
  AOI22_X1 npu_inst_pe_1_3_2_U113 ( .A1(npu_inst_int_data_y_4__2__0_), .A2(
        npu_inst_pe_1_3_2_n58), .B1(npu_inst_pe_1_3_2_n119), .B2(
        npu_inst_pe_1_3_2_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_3_2_n57) );
  INV_X1 npu_inst_pe_1_3_2_U112 ( .A(npu_inst_pe_1_3_2_n57), .ZN(
        npu_inst_pe_1_3_2_n108) );
  AOI22_X1 npu_inst_pe_1_3_2_U111 ( .A1(npu_inst_int_data_y_4__2__0_), .A2(
        npu_inst_pe_1_3_2_n54), .B1(npu_inst_pe_1_3_2_n118), .B2(
        npu_inst_pe_1_3_2_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_3_2_n53) );
  INV_X1 npu_inst_pe_1_3_2_U110 ( .A(npu_inst_pe_1_3_2_n53), .ZN(
        npu_inst_pe_1_3_2_n109) );
  AOI22_X1 npu_inst_pe_1_3_2_U107 ( .A1(npu_inst_int_data_y_4__2__0_), .A2(
        npu_inst_pe_1_3_2_n50), .B1(npu_inst_pe_1_3_2_n117), .B2(
        npu_inst_pe_1_3_2_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_3_2_n49) );
  INV_X1 npu_inst_pe_1_3_2_U106 ( .A(npu_inst_pe_1_3_2_n49), .ZN(
        npu_inst_pe_1_3_2_n110) );
  AOI22_X1 npu_inst_pe_1_3_2_U105 ( .A1(npu_inst_int_data_y_4__2__0_), .A2(
        npu_inst_pe_1_3_2_n46), .B1(npu_inst_pe_1_3_2_n116), .B2(
        npu_inst_pe_1_3_2_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_3_2_n45) );
  INV_X1 npu_inst_pe_1_3_2_U104 ( .A(npu_inst_pe_1_3_2_n45), .ZN(
        npu_inst_pe_1_3_2_n111) );
  AOI22_X1 npu_inst_pe_1_3_2_U103 ( .A1(npu_inst_int_data_y_4__2__0_), .A2(
        npu_inst_pe_1_3_2_n42), .B1(npu_inst_pe_1_3_2_n115), .B2(
        npu_inst_pe_1_3_2_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_3_2_n41) );
  INV_X1 npu_inst_pe_1_3_2_U102 ( .A(npu_inst_pe_1_3_2_n41), .ZN(
        npu_inst_pe_1_3_2_n112) );
  AOI22_X1 npu_inst_pe_1_3_2_U101 ( .A1(npu_inst_int_data_y_4__2__1_), .A2(
        npu_inst_pe_1_3_2_n58), .B1(npu_inst_pe_1_3_2_n119), .B2(
        npu_inst_pe_1_3_2_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_3_2_n59) );
  INV_X1 npu_inst_pe_1_3_2_U100 ( .A(npu_inst_pe_1_3_2_n59), .ZN(
        npu_inst_pe_1_3_2_n102) );
  AOI22_X1 npu_inst_pe_1_3_2_U99 ( .A1(npu_inst_int_data_y_4__2__1_), .A2(
        npu_inst_pe_1_3_2_n54), .B1(npu_inst_pe_1_3_2_n118), .B2(
        npu_inst_pe_1_3_2_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_3_2_n55) );
  INV_X1 npu_inst_pe_1_3_2_U98 ( .A(npu_inst_pe_1_3_2_n55), .ZN(
        npu_inst_pe_1_3_2_n103) );
  AOI22_X1 npu_inst_pe_1_3_2_U97 ( .A1(npu_inst_int_data_y_4__2__1_), .A2(
        npu_inst_pe_1_3_2_n50), .B1(npu_inst_pe_1_3_2_n117), .B2(
        npu_inst_pe_1_3_2_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_3_2_n51) );
  INV_X1 npu_inst_pe_1_3_2_U96 ( .A(npu_inst_pe_1_3_2_n51), .ZN(
        npu_inst_pe_1_3_2_n104) );
  AOI22_X1 npu_inst_pe_1_3_2_U95 ( .A1(npu_inst_int_data_y_4__2__1_), .A2(
        npu_inst_pe_1_3_2_n46), .B1(npu_inst_pe_1_3_2_n116), .B2(
        npu_inst_pe_1_3_2_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_3_2_n47) );
  INV_X1 npu_inst_pe_1_3_2_U94 ( .A(npu_inst_pe_1_3_2_n47), .ZN(
        npu_inst_pe_1_3_2_n105) );
  AOI22_X1 npu_inst_pe_1_3_2_U93 ( .A1(npu_inst_int_data_y_4__2__1_), .A2(
        npu_inst_pe_1_3_2_n42), .B1(npu_inst_pe_1_3_2_n115), .B2(
        npu_inst_pe_1_3_2_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_3_2_n43) );
  INV_X1 npu_inst_pe_1_3_2_U92 ( .A(npu_inst_pe_1_3_2_n43), .ZN(
        npu_inst_pe_1_3_2_n106) );
  AOI22_X1 npu_inst_pe_1_3_2_U91 ( .A1(npu_inst_pe_1_3_2_n38), .A2(
        npu_inst_int_data_y_4__2__1_), .B1(npu_inst_pe_1_3_2_n114), .B2(
        npu_inst_pe_1_3_2_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_3_2_n39) );
  INV_X1 npu_inst_pe_1_3_2_U90 ( .A(npu_inst_pe_1_3_2_n39), .ZN(
        npu_inst_pe_1_3_2_n107) );
  AOI22_X1 npu_inst_pe_1_3_2_U89 ( .A1(npu_inst_pe_1_3_2_n38), .A2(
        npu_inst_int_data_y_4__2__0_), .B1(npu_inst_pe_1_3_2_n114), .B2(
        npu_inst_pe_1_3_2_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_3_2_n37) );
  INV_X1 npu_inst_pe_1_3_2_U88 ( .A(npu_inst_pe_1_3_2_n37), .ZN(
        npu_inst_pe_1_3_2_n113) );
  NAND2_X1 npu_inst_pe_1_3_2_U87 ( .A1(npu_inst_pe_1_3_2_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_3_2_n60), .ZN(npu_inst_pe_1_3_2_n74) );
  OAI21_X1 npu_inst_pe_1_3_2_U86 ( .B1(npu_inst_pe_1_3_2_n63), .B2(
        npu_inst_pe_1_3_2_n60), .A(npu_inst_pe_1_3_2_n74), .ZN(
        npu_inst_pe_1_3_2_n97) );
  NAND2_X1 npu_inst_pe_1_3_2_U85 ( .A1(npu_inst_pe_1_3_2_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_3_2_n60), .ZN(npu_inst_pe_1_3_2_n73) );
  OAI21_X1 npu_inst_pe_1_3_2_U84 ( .B1(npu_inst_pe_1_3_2_n61), .B2(
        npu_inst_pe_1_3_2_n60), .A(npu_inst_pe_1_3_2_n73), .ZN(
        npu_inst_pe_1_3_2_n96) );
  NAND2_X1 npu_inst_pe_1_3_2_U83 ( .A1(npu_inst_pe_1_3_2_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_3_2_n56), .ZN(npu_inst_pe_1_3_2_n72) );
  OAI21_X1 npu_inst_pe_1_3_2_U82 ( .B1(npu_inst_pe_1_3_2_n63), .B2(
        npu_inst_pe_1_3_2_n56), .A(npu_inst_pe_1_3_2_n72), .ZN(
        npu_inst_pe_1_3_2_n95) );
  NAND2_X1 npu_inst_pe_1_3_2_U81 ( .A1(npu_inst_pe_1_3_2_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_3_2_n56), .ZN(npu_inst_pe_1_3_2_n71) );
  OAI21_X1 npu_inst_pe_1_3_2_U80 ( .B1(npu_inst_pe_1_3_2_n61), .B2(
        npu_inst_pe_1_3_2_n56), .A(npu_inst_pe_1_3_2_n71), .ZN(
        npu_inst_pe_1_3_2_n94) );
  NAND2_X1 npu_inst_pe_1_3_2_U79 ( .A1(npu_inst_pe_1_3_2_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_3_2_n52), .ZN(npu_inst_pe_1_3_2_n70) );
  OAI21_X1 npu_inst_pe_1_3_2_U78 ( .B1(npu_inst_pe_1_3_2_n63), .B2(
        npu_inst_pe_1_3_2_n52), .A(npu_inst_pe_1_3_2_n70), .ZN(
        npu_inst_pe_1_3_2_n93) );
  NAND2_X1 npu_inst_pe_1_3_2_U77 ( .A1(npu_inst_pe_1_3_2_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_3_2_n52), .ZN(npu_inst_pe_1_3_2_n69) );
  OAI21_X1 npu_inst_pe_1_3_2_U76 ( .B1(npu_inst_pe_1_3_2_n61), .B2(
        npu_inst_pe_1_3_2_n52), .A(npu_inst_pe_1_3_2_n69), .ZN(
        npu_inst_pe_1_3_2_n92) );
  NAND2_X1 npu_inst_pe_1_3_2_U75 ( .A1(npu_inst_pe_1_3_2_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_3_2_n48), .ZN(npu_inst_pe_1_3_2_n68) );
  OAI21_X1 npu_inst_pe_1_3_2_U74 ( .B1(npu_inst_pe_1_3_2_n63), .B2(
        npu_inst_pe_1_3_2_n48), .A(npu_inst_pe_1_3_2_n68), .ZN(
        npu_inst_pe_1_3_2_n91) );
  NAND2_X1 npu_inst_pe_1_3_2_U73 ( .A1(npu_inst_pe_1_3_2_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_3_2_n48), .ZN(npu_inst_pe_1_3_2_n67) );
  OAI21_X1 npu_inst_pe_1_3_2_U72 ( .B1(npu_inst_pe_1_3_2_n61), .B2(
        npu_inst_pe_1_3_2_n48), .A(npu_inst_pe_1_3_2_n67), .ZN(
        npu_inst_pe_1_3_2_n90) );
  NAND2_X1 npu_inst_pe_1_3_2_U71 ( .A1(npu_inst_pe_1_3_2_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_3_2_n44), .ZN(npu_inst_pe_1_3_2_n66) );
  OAI21_X1 npu_inst_pe_1_3_2_U70 ( .B1(npu_inst_pe_1_3_2_n63), .B2(
        npu_inst_pe_1_3_2_n44), .A(npu_inst_pe_1_3_2_n66), .ZN(
        npu_inst_pe_1_3_2_n89) );
  NAND2_X1 npu_inst_pe_1_3_2_U69 ( .A1(npu_inst_pe_1_3_2_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_3_2_n44), .ZN(npu_inst_pe_1_3_2_n65) );
  OAI21_X1 npu_inst_pe_1_3_2_U68 ( .B1(npu_inst_pe_1_3_2_n61), .B2(
        npu_inst_pe_1_3_2_n44), .A(npu_inst_pe_1_3_2_n65), .ZN(
        npu_inst_pe_1_3_2_n88) );
  NAND2_X1 npu_inst_pe_1_3_2_U67 ( .A1(npu_inst_pe_1_3_2_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_3_2_n40), .ZN(npu_inst_pe_1_3_2_n64) );
  OAI21_X1 npu_inst_pe_1_3_2_U66 ( .B1(npu_inst_pe_1_3_2_n63), .B2(
        npu_inst_pe_1_3_2_n40), .A(npu_inst_pe_1_3_2_n64), .ZN(
        npu_inst_pe_1_3_2_n87) );
  NAND2_X1 npu_inst_pe_1_3_2_U65 ( .A1(npu_inst_pe_1_3_2_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_3_2_n40), .ZN(npu_inst_pe_1_3_2_n62) );
  OAI21_X1 npu_inst_pe_1_3_2_U64 ( .B1(npu_inst_pe_1_3_2_n61), .B2(
        npu_inst_pe_1_3_2_n40), .A(npu_inst_pe_1_3_2_n62), .ZN(
        npu_inst_pe_1_3_2_n86) );
  AND2_X1 npu_inst_pe_1_3_2_U63 ( .A1(npu_inst_pe_1_3_2_N93), .A2(npu_inst_n57), .ZN(npu_inst_int_data_y_3__2__0_) );
  AND2_X1 npu_inst_pe_1_3_2_U62 ( .A1(npu_inst_n57), .A2(npu_inst_pe_1_3_2_N94), .ZN(npu_inst_int_data_y_3__2__1_) );
  NOR3_X1 npu_inst_pe_1_3_2_U61 ( .A1(npu_inst_pe_1_3_2_n26), .A2(npu_inst_n57), .A3(npu_inst_int_ckg[37]), .ZN(npu_inst_pe_1_3_2_n85) );
  OR2_X1 npu_inst_pe_1_3_2_U60 ( .A1(npu_inst_pe_1_3_2_n85), .A2(
        npu_inst_pe_1_3_2_n2), .ZN(npu_inst_pe_1_3_2_N84) );
  AND2_X1 npu_inst_pe_1_3_2_U59 ( .A1(npu_inst_pe_1_3_2_int_q_acc_0_), .A2(
        npu_inst_pe_1_3_2_n1), .ZN(npu_inst_int_data_res_3__2__0_) );
  AND2_X1 npu_inst_pe_1_3_2_U58 ( .A1(npu_inst_pe_1_3_2_n2), .A2(
        npu_inst_pe_1_3_2_int_q_acc_7_), .ZN(npu_inst_int_data_res_3__2__7_)
         );
  AND2_X1 npu_inst_pe_1_3_2_U57 ( .A1(npu_inst_pe_1_3_2_int_q_acc_1_), .A2(
        npu_inst_pe_1_3_2_n1), .ZN(npu_inst_int_data_res_3__2__1_) );
  AND2_X1 npu_inst_pe_1_3_2_U56 ( .A1(npu_inst_pe_1_3_2_int_q_acc_2_), .A2(
        npu_inst_pe_1_3_2_n1), .ZN(npu_inst_int_data_res_3__2__2_) );
  AND2_X1 npu_inst_pe_1_3_2_U55 ( .A1(npu_inst_pe_1_3_2_int_q_acc_3_), .A2(
        npu_inst_pe_1_3_2_n2), .ZN(npu_inst_int_data_res_3__2__3_) );
  AND2_X1 npu_inst_pe_1_3_2_U54 ( .A1(npu_inst_pe_1_3_2_int_q_acc_4_), .A2(
        npu_inst_pe_1_3_2_n2), .ZN(npu_inst_int_data_res_3__2__4_) );
  AND2_X1 npu_inst_pe_1_3_2_U53 ( .A1(npu_inst_pe_1_3_2_int_q_acc_5_), .A2(
        npu_inst_pe_1_3_2_n2), .ZN(npu_inst_int_data_res_3__2__5_) );
  AND2_X1 npu_inst_pe_1_3_2_U52 ( .A1(npu_inst_pe_1_3_2_int_q_acc_6_), .A2(
        npu_inst_pe_1_3_2_n2), .ZN(npu_inst_int_data_res_3__2__6_) );
  AOI222_X1 npu_inst_pe_1_3_2_U51 ( .A1(npu_inst_int_data_res_4__2__0_), .A2(
        npu_inst_pe_1_3_2_n1), .B1(npu_inst_pe_1_3_2_N73), .B2(
        npu_inst_pe_1_3_2_n76), .C1(npu_inst_pe_1_3_2_N65), .C2(
        npu_inst_pe_1_3_2_n77), .ZN(npu_inst_pe_1_3_2_n84) );
  INV_X1 npu_inst_pe_1_3_2_U50 ( .A(npu_inst_pe_1_3_2_n84), .ZN(
        npu_inst_pe_1_3_2_n101) );
  AOI222_X1 npu_inst_pe_1_3_2_U49 ( .A1(npu_inst_int_data_res_4__2__7_), .A2(
        npu_inst_pe_1_3_2_n1), .B1(npu_inst_pe_1_3_2_N80), .B2(
        npu_inst_pe_1_3_2_n76), .C1(npu_inst_pe_1_3_2_N72), .C2(
        npu_inst_pe_1_3_2_n77), .ZN(npu_inst_pe_1_3_2_n75) );
  INV_X1 npu_inst_pe_1_3_2_U48 ( .A(npu_inst_pe_1_3_2_n75), .ZN(
        npu_inst_pe_1_3_2_n33) );
  AOI222_X1 npu_inst_pe_1_3_2_U47 ( .A1(npu_inst_int_data_res_4__2__1_), .A2(
        npu_inst_pe_1_3_2_n1), .B1(npu_inst_pe_1_3_2_N74), .B2(
        npu_inst_pe_1_3_2_n76), .C1(npu_inst_pe_1_3_2_N66), .C2(
        npu_inst_pe_1_3_2_n77), .ZN(npu_inst_pe_1_3_2_n83) );
  INV_X1 npu_inst_pe_1_3_2_U46 ( .A(npu_inst_pe_1_3_2_n83), .ZN(
        npu_inst_pe_1_3_2_n100) );
  AOI222_X1 npu_inst_pe_1_3_2_U45 ( .A1(npu_inst_int_data_res_4__2__2_), .A2(
        npu_inst_pe_1_3_2_n1), .B1(npu_inst_pe_1_3_2_N75), .B2(
        npu_inst_pe_1_3_2_n76), .C1(npu_inst_pe_1_3_2_N67), .C2(
        npu_inst_pe_1_3_2_n77), .ZN(npu_inst_pe_1_3_2_n82) );
  INV_X1 npu_inst_pe_1_3_2_U44 ( .A(npu_inst_pe_1_3_2_n82), .ZN(
        npu_inst_pe_1_3_2_n99) );
  AOI222_X1 npu_inst_pe_1_3_2_U43 ( .A1(npu_inst_int_data_res_4__2__3_), .A2(
        npu_inst_pe_1_3_2_n1), .B1(npu_inst_pe_1_3_2_N76), .B2(
        npu_inst_pe_1_3_2_n76), .C1(npu_inst_pe_1_3_2_N68), .C2(
        npu_inst_pe_1_3_2_n77), .ZN(npu_inst_pe_1_3_2_n81) );
  INV_X1 npu_inst_pe_1_3_2_U42 ( .A(npu_inst_pe_1_3_2_n81), .ZN(
        npu_inst_pe_1_3_2_n98) );
  AOI222_X1 npu_inst_pe_1_3_2_U41 ( .A1(npu_inst_int_data_res_4__2__4_), .A2(
        npu_inst_pe_1_3_2_n1), .B1(npu_inst_pe_1_3_2_N77), .B2(
        npu_inst_pe_1_3_2_n76), .C1(npu_inst_pe_1_3_2_N69), .C2(
        npu_inst_pe_1_3_2_n77), .ZN(npu_inst_pe_1_3_2_n80) );
  INV_X1 npu_inst_pe_1_3_2_U40 ( .A(npu_inst_pe_1_3_2_n80), .ZN(
        npu_inst_pe_1_3_2_n36) );
  AOI222_X1 npu_inst_pe_1_3_2_U39 ( .A1(npu_inst_int_data_res_4__2__5_), .A2(
        npu_inst_pe_1_3_2_n1), .B1(npu_inst_pe_1_3_2_N78), .B2(
        npu_inst_pe_1_3_2_n76), .C1(npu_inst_pe_1_3_2_N70), .C2(
        npu_inst_pe_1_3_2_n77), .ZN(npu_inst_pe_1_3_2_n79) );
  INV_X1 npu_inst_pe_1_3_2_U38 ( .A(npu_inst_pe_1_3_2_n79), .ZN(
        npu_inst_pe_1_3_2_n35) );
  AOI222_X1 npu_inst_pe_1_3_2_U37 ( .A1(npu_inst_int_data_res_4__2__6_), .A2(
        npu_inst_pe_1_3_2_n1), .B1(npu_inst_pe_1_3_2_N79), .B2(
        npu_inst_pe_1_3_2_n76), .C1(npu_inst_pe_1_3_2_N71), .C2(
        npu_inst_pe_1_3_2_n77), .ZN(npu_inst_pe_1_3_2_n78) );
  INV_X1 npu_inst_pe_1_3_2_U36 ( .A(npu_inst_pe_1_3_2_n78), .ZN(
        npu_inst_pe_1_3_2_n34) );
  INV_X1 npu_inst_pe_1_3_2_U35 ( .A(npu_inst_pe_1_3_2_int_data_1_), .ZN(
        npu_inst_pe_1_3_2_n14) );
  AND2_X1 npu_inst_pe_1_3_2_U34 ( .A1(npu_inst_int_data_x_3__2__1_), .A2(
        npu_inst_pe_1_3_2_int_q_weight_1_), .ZN(npu_inst_pe_1_3_2_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_3_2_U33 ( .A1(npu_inst_int_data_x_3__2__0_), .A2(
        npu_inst_pe_1_3_2_int_q_weight_1_), .ZN(npu_inst_pe_1_3_2_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_3_2_U32 ( .A1(npu_inst_n57), .A2(
        npu_inst_int_data_y_4__2__1_), .B1(npu_inst_pe_1_3_2_n3), .B2(
        npu_inst_int_data_x_3__3__1_), .ZN(npu_inst_pe_1_3_2_n63) );
  AOI22_X1 npu_inst_pe_1_3_2_U31 ( .A1(npu_inst_n57), .A2(
        npu_inst_int_data_y_4__2__0_), .B1(npu_inst_pe_1_3_2_n3), .B2(
        npu_inst_int_data_x_3__3__0_), .ZN(npu_inst_pe_1_3_2_n61) );
  INV_X1 npu_inst_pe_1_3_2_U30 ( .A(npu_inst_pe_1_3_2_int_data_0_), .ZN(
        npu_inst_pe_1_3_2_n13) );
  INV_X1 npu_inst_pe_1_3_2_U29 ( .A(npu_inst_n70), .ZN(npu_inst_pe_1_3_2_n5)
         );
  OR3_X1 npu_inst_pe_1_3_2_U28 ( .A1(npu_inst_pe_1_3_2_n6), .A2(
        npu_inst_pe_1_3_2_n8), .A3(npu_inst_pe_1_3_2_n5), .ZN(
        npu_inst_pe_1_3_2_n56) );
  OR3_X1 npu_inst_pe_1_3_2_U27 ( .A1(npu_inst_pe_1_3_2_n5), .A2(
        npu_inst_pe_1_3_2_n8), .A3(npu_inst_pe_1_3_2_n7), .ZN(
        npu_inst_pe_1_3_2_n48) );
  INV_X1 npu_inst_pe_1_3_2_U26 ( .A(npu_inst_pe_1_3_2_n5), .ZN(
        npu_inst_pe_1_3_2_n4) );
  OR3_X1 npu_inst_pe_1_3_2_U25 ( .A1(npu_inst_pe_1_3_2_n4), .A2(
        npu_inst_pe_1_3_2_n8), .A3(npu_inst_pe_1_3_2_n7), .ZN(
        npu_inst_pe_1_3_2_n52) );
  OR3_X1 npu_inst_pe_1_3_2_U24 ( .A1(npu_inst_pe_1_3_2_n6), .A2(
        npu_inst_pe_1_3_2_n8), .A3(npu_inst_pe_1_3_2_n4), .ZN(
        npu_inst_pe_1_3_2_n60) );
  NOR2_X1 npu_inst_pe_1_3_2_U23 ( .A1(npu_inst_pe_1_3_2_n60), .A2(
        npu_inst_pe_1_3_2_n3), .ZN(npu_inst_pe_1_3_2_n58) );
  NOR2_X1 npu_inst_pe_1_3_2_U22 ( .A1(npu_inst_pe_1_3_2_n56), .A2(
        npu_inst_pe_1_3_2_n3), .ZN(npu_inst_pe_1_3_2_n54) );
  NOR2_X1 npu_inst_pe_1_3_2_U21 ( .A1(npu_inst_pe_1_3_2_n52), .A2(
        npu_inst_pe_1_3_2_n3), .ZN(npu_inst_pe_1_3_2_n50) );
  NOR2_X1 npu_inst_pe_1_3_2_U20 ( .A1(npu_inst_pe_1_3_2_n48), .A2(
        npu_inst_pe_1_3_2_n3), .ZN(npu_inst_pe_1_3_2_n46) );
  NOR2_X1 npu_inst_pe_1_3_2_U19 ( .A1(npu_inst_pe_1_3_2_n40), .A2(
        npu_inst_pe_1_3_2_n3), .ZN(npu_inst_pe_1_3_2_n38) );
  NOR2_X1 npu_inst_pe_1_3_2_U18 ( .A1(npu_inst_pe_1_3_2_n44), .A2(
        npu_inst_pe_1_3_2_n3), .ZN(npu_inst_pe_1_3_2_n42) );
  BUF_X1 npu_inst_pe_1_3_2_U17 ( .A(npu_inst_n101), .Z(npu_inst_pe_1_3_2_n8)
         );
  INV_X1 npu_inst_pe_1_3_2_U16 ( .A(npu_inst_n125), .ZN(npu_inst_pe_1_3_2_n12)
         );
  INV_X1 npu_inst_pe_1_3_2_U15 ( .A(npu_inst_pe_1_3_2_n38), .ZN(
        npu_inst_pe_1_3_2_n114) );
  INV_X1 npu_inst_pe_1_3_2_U14 ( .A(npu_inst_pe_1_3_2_n58), .ZN(
        npu_inst_pe_1_3_2_n119) );
  INV_X1 npu_inst_pe_1_3_2_U13 ( .A(npu_inst_pe_1_3_2_n54), .ZN(
        npu_inst_pe_1_3_2_n118) );
  INV_X1 npu_inst_pe_1_3_2_U12 ( .A(npu_inst_pe_1_3_2_n50), .ZN(
        npu_inst_pe_1_3_2_n117) );
  INV_X1 npu_inst_pe_1_3_2_U11 ( .A(npu_inst_pe_1_3_2_n46), .ZN(
        npu_inst_pe_1_3_2_n116) );
  INV_X1 npu_inst_pe_1_3_2_U10 ( .A(npu_inst_pe_1_3_2_n42), .ZN(
        npu_inst_pe_1_3_2_n115) );
  BUF_X1 npu_inst_pe_1_3_2_U9 ( .A(npu_inst_n25), .Z(npu_inst_pe_1_3_2_n2) );
  BUF_X1 npu_inst_pe_1_3_2_U8 ( .A(npu_inst_n25), .Z(npu_inst_pe_1_3_2_n1) );
  BUF_X1 npu_inst_pe_1_3_2_U7 ( .A(npu_inst_pe_1_3_2_n12), .Z(
        npu_inst_pe_1_3_2_n11) );
  BUF_X1 npu_inst_pe_1_3_2_U6 ( .A(npu_inst_pe_1_3_2_n12), .Z(
        npu_inst_pe_1_3_2_n10) );
  BUF_X1 npu_inst_pe_1_3_2_U5 ( .A(npu_inst_pe_1_3_2_n12), .Z(
        npu_inst_pe_1_3_2_n9) );
  NOR2_X1 npu_inst_pe_1_3_2_U4 ( .A1(npu_inst_pe_1_3_2_int_q_weight_0_), .A2(
        npu_inst_pe_1_3_2_n1), .ZN(npu_inst_pe_1_3_2_n76) );
  NOR2_X1 npu_inst_pe_1_3_2_U3 ( .A1(npu_inst_pe_1_3_2_n27), .A2(
        npu_inst_pe_1_3_2_n1), .ZN(npu_inst_pe_1_3_2_n77) );
  FA_X1 npu_inst_pe_1_3_2_sub_67_U2_1 ( .A(npu_inst_pe_1_3_2_int_q_acc_1_), 
        .B(npu_inst_pe_1_3_2_n14), .CI(npu_inst_pe_1_3_2_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_3_2_sub_67_carry_2_), .S(npu_inst_pe_1_3_2_N66) );
  FA_X1 npu_inst_pe_1_3_2_add_69_U1_1 ( .A(npu_inst_pe_1_3_2_int_q_acc_1_), 
        .B(npu_inst_pe_1_3_2_int_data_1_), .CI(
        npu_inst_pe_1_3_2_add_69_carry_1_), .CO(
        npu_inst_pe_1_3_2_add_69_carry_2_), .S(npu_inst_pe_1_3_2_N74) );
  NAND3_X1 npu_inst_pe_1_3_2_U109 ( .A1(npu_inst_pe_1_3_2_n5), .A2(
        npu_inst_pe_1_3_2_n7), .A3(npu_inst_pe_1_3_2_n8), .ZN(
        npu_inst_pe_1_3_2_n44) );
  NAND3_X1 npu_inst_pe_1_3_2_U108 ( .A1(npu_inst_pe_1_3_2_n4), .A2(
        npu_inst_pe_1_3_2_n7), .A3(npu_inst_pe_1_3_2_n8), .ZN(
        npu_inst_pe_1_3_2_n40) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_3_2_n34), .CK(
        npu_inst_pe_1_3_2_net3964), .RN(npu_inst_pe_1_3_2_n9), .Q(
        npu_inst_pe_1_3_2_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_3_2_n35), .CK(
        npu_inst_pe_1_3_2_net3964), .RN(npu_inst_pe_1_3_2_n9), .Q(
        npu_inst_pe_1_3_2_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_3_2_n36), .CK(
        npu_inst_pe_1_3_2_net3964), .RN(npu_inst_pe_1_3_2_n9), .Q(
        npu_inst_pe_1_3_2_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_3_2_n98), .CK(
        npu_inst_pe_1_3_2_net3964), .RN(npu_inst_pe_1_3_2_n9), .Q(
        npu_inst_pe_1_3_2_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_3_2_n99), .CK(
        npu_inst_pe_1_3_2_net3964), .RN(npu_inst_pe_1_3_2_n9), .Q(
        npu_inst_pe_1_3_2_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_3_2_n100), 
        .CK(npu_inst_pe_1_3_2_net3964), .RN(npu_inst_pe_1_3_2_n9), .Q(
        npu_inst_pe_1_3_2_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_3_2_n33), .CK(
        npu_inst_pe_1_3_2_net3964), .RN(npu_inst_pe_1_3_2_n9), .Q(
        npu_inst_pe_1_3_2_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_3_2_n101), 
        .CK(npu_inst_pe_1_3_2_net3964), .RN(npu_inst_pe_1_3_2_n9), .Q(
        npu_inst_pe_1_3_2_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_weight_reg_0_ ( .D(npu_inst_n111), .CK(
        npu_inst_pe_1_3_2_net3970), .RN(npu_inst_pe_1_3_2_n9), .Q(
        npu_inst_pe_1_3_2_int_q_weight_0_), .QN(npu_inst_pe_1_3_2_n27) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_weight_reg_1_ ( .D(npu_inst_n117), .CK(
        npu_inst_pe_1_3_2_net3970), .RN(npu_inst_pe_1_3_2_n9), .Q(
        npu_inst_pe_1_3_2_int_q_weight_1_), .QN(npu_inst_pe_1_3_2_n26) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_3_2_n113), 
        .CK(npu_inst_pe_1_3_2_net3970), .RN(npu_inst_pe_1_3_2_n9), .Q(
        npu_inst_pe_1_3_2_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_3_2_n107), 
        .CK(npu_inst_pe_1_3_2_net3970), .RN(npu_inst_pe_1_3_2_n9), .Q(
        npu_inst_pe_1_3_2_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_3_2_n112), 
        .CK(npu_inst_pe_1_3_2_net3970), .RN(npu_inst_pe_1_3_2_n10), .Q(
        npu_inst_pe_1_3_2_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_3_2_n106), 
        .CK(npu_inst_pe_1_3_2_net3970), .RN(npu_inst_pe_1_3_2_n10), .Q(
        npu_inst_pe_1_3_2_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_3_2_n111), 
        .CK(npu_inst_pe_1_3_2_net3970), .RN(npu_inst_pe_1_3_2_n10), .Q(
        npu_inst_pe_1_3_2_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_3_2_n105), 
        .CK(npu_inst_pe_1_3_2_net3970), .RN(npu_inst_pe_1_3_2_n10), .Q(
        npu_inst_pe_1_3_2_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_3_2_n110), 
        .CK(npu_inst_pe_1_3_2_net3970), .RN(npu_inst_pe_1_3_2_n10), .Q(
        npu_inst_pe_1_3_2_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_3_2_n104), 
        .CK(npu_inst_pe_1_3_2_net3970), .RN(npu_inst_pe_1_3_2_n10), .Q(
        npu_inst_pe_1_3_2_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_3_2_n109), 
        .CK(npu_inst_pe_1_3_2_net3970), .RN(npu_inst_pe_1_3_2_n10), .Q(
        npu_inst_pe_1_3_2_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_3_2_n103), 
        .CK(npu_inst_pe_1_3_2_net3970), .RN(npu_inst_pe_1_3_2_n10), .Q(
        npu_inst_pe_1_3_2_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_3_2_n108), 
        .CK(npu_inst_pe_1_3_2_net3970), .RN(npu_inst_pe_1_3_2_n10), .Q(
        npu_inst_pe_1_3_2_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_3_2_n102), 
        .CK(npu_inst_pe_1_3_2_net3970), .RN(npu_inst_pe_1_3_2_n10), .Q(
        npu_inst_pe_1_3_2_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_3_2_n86), 
        .CK(npu_inst_pe_1_3_2_net3970), .RN(npu_inst_pe_1_3_2_n10), .Q(
        npu_inst_pe_1_3_2_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_3_2_n87), 
        .CK(npu_inst_pe_1_3_2_net3970), .RN(npu_inst_pe_1_3_2_n10), .Q(
        npu_inst_pe_1_3_2_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_3_2_n88), 
        .CK(npu_inst_pe_1_3_2_net3970), .RN(npu_inst_pe_1_3_2_n11), .Q(
        npu_inst_pe_1_3_2_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_3_2_n89), 
        .CK(npu_inst_pe_1_3_2_net3970), .RN(npu_inst_pe_1_3_2_n11), .Q(
        npu_inst_pe_1_3_2_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_3_2_n90), 
        .CK(npu_inst_pe_1_3_2_net3970), .RN(npu_inst_pe_1_3_2_n11), .Q(
        npu_inst_pe_1_3_2_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_3_2_n91), 
        .CK(npu_inst_pe_1_3_2_net3970), .RN(npu_inst_pe_1_3_2_n11), .Q(
        npu_inst_pe_1_3_2_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_3_2_n92), 
        .CK(npu_inst_pe_1_3_2_net3970), .RN(npu_inst_pe_1_3_2_n11), .Q(
        npu_inst_pe_1_3_2_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_3_2_n93), 
        .CK(npu_inst_pe_1_3_2_net3970), .RN(npu_inst_pe_1_3_2_n11), .Q(
        npu_inst_pe_1_3_2_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_3_2_n94), 
        .CK(npu_inst_pe_1_3_2_net3970), .RN(npu_inst_pe_1_3_2_n11), .Q(
        npu_inst_pe_1_3_2_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_3_2_n95), 
        .CK(npu_inst_pe_1_3_2_net3970), .RN(npu_inst_pe_1_3_2_n11), .Q(
        npu_inst_pe_1_3_2_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_3_2_n96), 
        .CK(npu_inst_pe_1_3_2_net3970), .RN(npu_inst_pe_1_3_2_n11), .Q(
        npu_inst_pe_1_3_2_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_3_2_n97), 
        .CK(npu_inst_pe_1_3_2_net3970), .RN(npu_inst_pe_1_3_2_n11), .Q(
        npu_inst_pe_1_3_2_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_3_2_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_3_2_N84), .SE(1'b0), .GCK(npu_inst_pe_1_3_2_net3964) );
  CLKGATETST_X1 npu_inst_pe_1_3_2_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n64), .SE(1'b0), .GCK(npu_inst_pe_1_3_2_net3970) );
  MUX2_X1 npu_inst_pe_1_3_3_U162 ( .A(npu_inst_pe_1_3_3_n32), .B(
        npu_inst_pe_1_3_3_n29), .S(npu_inst_pe_1_3_3_n8), .Z(
        npu_inst_pe_1_3_3_N93) );
  MUX2_X1 npu_inst_pe_1_3_3_U161 ( .A(npu_inst_pe_1_3_3_n31), .B(
        npu_inst_pe_1_3_3_n30), .S(npu_inst_pe_1_3_3_n6), .Z(
        npu_inst_pe_1_3_3_n32) );
  MUX2_X1 npu_inst_pe_1_3_3_U160 ( .A(npu_inst_pe_1_3_3_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_3_3_int_q_reg_v_1__0_), .S(npu_inst_pe_1_3_3_n4), .Z(
        npu_inst_pe_1_3_3_n31) );
  MUX2_X1 npu_inst_pe_1_3_3_U159 ( .A(npu_inst_pe_1_3_3_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_3_3_int_q_reg_v_3__0_), .S(npu_inst_pe_1_3_3_n4), .Z(
        npu_inst_pe_1_3_3_n30) );
  MUX2_X1 npu_inst_pe_1_3_3_U158 ( .A(npu_inst_pe_1_3_3_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_3_3_int_q_reg_v_5__0_), .S(npu_inst_pe_1_3_3_n4), .Z(
        npu_inst_pe_1_3_3_n29) );
  MUX2_X1 npu_inst_pe_1_3_3_U157 ( .A(npu_inst_pe_1_3_3_n28), .B(
        npu_inst_pe_1_3_3_n23), .S(npu_inst_pe_1_3_3_n8), .Z(
        npu_inst_pe_1_3_3_N94) );
  MUX2_X1 npu_inst_pe_1_3_3_U156 ( .A(npu_inst_pe_1_3_3_n25), .B(
        npu_inst_pe_1_3_3_n24), .S(npu_inst_pe_1_3_3_n6), .Z(
        npu_inst_pe_1_3_3_n28) );
  MUX2_X1 npu_inst_pe_1_3_3_U155 ( .A(npu_inst_pe_1_3_3_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_3_3_int_q_reg_v_1__1_), .S(npu_inst_pe_1_3_3_n4), .Z(
        npu_inst_pe_1_3_3_n25) );
  MUX2_X1 npu_inst_pe_1_3_3_U154 ( .A(npu_inst_pe_1_3_3_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_3_3_int_q_reg_v_3__1_), .S(npu_inst_pe_1_3_3_n4), .Z(
        npu_inst_pe_1_3_3_n24) );
  MUX2_X1 npu_inst_pe_1_3_3_U153 ( .A(npu_inst_pe_1_3_3_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_3_3_int_q_reg_v_5__1_), .S(npu_inst_pe_1_3_3_n4), .Z(
        npu_inst_pe_1_3_3_n23) );
  MUX2_X1 npu_inst_pe_1_3_3_U152 ( .A(npu_inst_pe_1_3_3_n22), .B(
        npu_inst_pe_1_3_3_n19), .S(npu_inst_pe_1_3_3_n8), .Z(
        npu_inst_int_data_x_3__3__1_) );
  MUX2_X1 npu_inst_pe_1_3_3_U151 ( .A(npu_inst_pe_1_3_3_n21), .B(
        npu_inst_pe_1_3_3_n20), .S(npu_inst_pe_1_3_3_n6), .Z(
        npu_inst_pe_1_3_3_n22) );
  MUX2_X1 npu_inst_pe_1_3_3_U150 ( .A(npu_inst_pe_1_3_3_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_3_3_int_q_reg_h_1__1_), .S(npu_inst_pe_1_3_3_n4), .Z(
        npu_inst_pe_1_3_3_n21) );
  MUX2_X1 npu_inst_pe_1_3_3_U149 ( .A(npu_inst_pe_1_3_3_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_3_3_int_q_reg_h_3__1_), .S(npu_inst_pe_1_3_3_n4), .Z(
        npu_inst_pe_1_3_3_n20) );
  MUX2_X1 npu_inst_pe_1_3_3_U148 ( .A(npu_inst_pe_1_3_3_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_3_3_int_q_reg_h_5__1_), .S(npu_inst_pe_1_3_3_n4), .Z(
        npu_inst_pe_1_3_3_n19) );
  MUX2_X1 npu_inst_pe_1_3_3_U147 ( .A(npu_inst_pe_1_3_3_n18), .B(
        npu_inst_pe_1_3_3_n15), .S(npu_inst_pe_1_3_3_n8), .Z(
        npu_inst_int_data_x_3__3__0_) );
  MUX2_X1 npu_inst_pe_1_3_3_U146 ( .A(npu_inst_pe_1_3_3_n17), .B(
        npu_inst_pe_1_3_3_n16), .S(npu_inst_pe_1_3_3_n6), .Z(
        npu_inst_pe_1_3_3_n18) );
  MUX2_X1 npu_inst_pe_1_3_3_U145 ( .A(npu_inst_pe_1_3_3_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_3_3_int_q_reg_h_1__0_), .S(npu_inst_pe_1_3_3_n4), .Z(
        npu_inst_pe_1_3_3_n17) );
  MUX2_X1 npu_inst_pe_1_3_3_U144 ( .A(npu_inst_pe_1_3_3_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_3_3_int_q_reg_h_3__0_), .S(npu_inst_pe_1_3_3_n4), .Z(
        npu_inst_pe_1_3_3_n16) );
  MUX2_X1 npu_inst_pe_1_3_3_U143 ( .A(npu_inst_pe_1_3_3_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_3_3_int_q_reg_h_5__0_), .S(npu_inst_pe_1_3_3_n4), .Z(
        npu_inst_pe_1_3_3_n15) );
  XOR2_X1 npu_inst_pe_1_3_3_U142 ( .A(npu_inst_pe_1_3_3_int_data_0_), .B(
        npu_inst_pe_1_3_3_int_q_acc_0_), .Z(npu_inst_pe_1_3_3_N73) );
  AND2_X1 npu_inst_pe_1_3_3_U141 ( .A1(npu_inst_pe_1_3_3_int_q_acc_0_), .A2(
        npu_inst_pe_1_3_3_int_data_0_), .ZN(npu_inst_pe_1_3_3_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_3_3_U140 ( .A(npu_inst_pe_1_3_3_int_q_acc_0_), .B(
        npu_inst_pe_1_3_3_n13), .ZN(npu_inst_pe_1_3_3_N65) );
  OR2_X1 npu_inst_pe_1_3_3_U139 ( .A1(npu_inst_pe_1_3_3_n13), .A2(
        npu_inst_pe_1_3_3_int_q_acc_0_), .ZN(npu_inst_pe_1_3_3_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_3_3_U138 ( .A(npu_inst_pe_1_3_3_int_q_acc_2_), .B(
        npu_inst_pe_1_3_3_add_69_carry_2_), .Z(npu_inst_pe_1_3_3_N75) );
  AND2_X1 npu_inst_pe_1_3_3_U137 ( .A1(npu_inst_pe_1_3_3_add_69_carry_2_), 
        .A2(npu_inst_pe_1_3_3_int_q_acc_2_), .ZN(
        npu_inst_pe_1_3_3_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_3_3_U136 ( .A(npu_inst_pe_1_3_3_int_q_acc_3_), .B(
        npu_inst_pe_1_3_3_add_69_carry_3_), .Z(npu_inst_pe_1_3_3_N76) );
  AND2_X1 npu_inst_pe_1_3_3_U135 ( .A1(npu_inst_pe_1_3_3_add_69_carry_3_), 
        .A2(npu_inst_pe_1_3_3_int_q_acc_3_), .ZN(
        npu_inst_pe_1_3_3_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_3_3_U134 ( .A(npu_inst_pe_1_3_3_int_q_acc_4_), .B(
        npu_inst_pe_1_3_3_add_69_carry_4_), .Z(npu_inst_pe_1_3_3_N77) );
  AND2_X1 npu_inst_pe_1_3_3_U133 ( .A1(npu_inst_pe_1_3_3_add_69_carry_4_), 
        .A2(npu_inst_pe_1_3_3_int_q_acc_4_), .ZN(
        npu_inst_pe_1_3_3_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_3_3_U132 ( .A(npu_inst_pe_1_3_3_int_q_acc_5_), .B(
        npu_inst_pe_1_3_3_add_69_carry_5_), .Z(npu_inst_pe_1_3_3_N78) );
  AND2_X1 npu_inst_pe_1_3_3_U131 ( .A1(npu_inst_pe_1_3_3_add_69_carry_5_), 
        .A2(npu_inst_pe_1_3_3_int_q_acc_5_), .ZN(
        npu_inst_pe_1_3_3_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_3_3_U130 ( .A(npu_inst_pe_1_3_3_int_q_acc_6_), .B(
        npu_inst_pe_1_3_3_add_69_carry_6_), .Z(npu_inst_pe_1_3_3_N79) );
  AND2_X1 npu_inst_pe_1_3_3_U129 ( .A1(npu_inst_pe_1_3_3_add_69_carry_6_), 
        .A2(npu_inst_pe_1_3_3_int_q_acc_6_), .ZN(
        npu_inst_pe_1_3_3_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_3_3_U128 ( .A(npu_inst_pe_1_3_3_int_q_acc_7_), .B(
        npu_inst_pe_1_3_3_add_69_carry_7_), .Z(npu_inst_pe_1_3_3_N80) );
  XNOR2_X1 npu_inst_pe_1_3_3_U127 ( .A(npu_inst_pe_1_3_3_sub_67_carry_2_), .B(
        npu_inst_pe_1_3_3_int_q_acc_2_), .ZN(npu_inst_pe_1_3_3_N67) );
  OR2_X1 npu_inst_pe_1_3_3_U126 ( .A1(npu_inst_pe_1_3_3_int_q_acc_2_), .A2(
        npu_inst_pe_1_3_3_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_3_3_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_3_3_U125 ( .A(npu_inst_pe_1_3_3_sub_67_carry_3_), .B(
        npu_inst_pe_1_3_3_int_q_acc_3_), .ZN(npu_inst_pe_1_3_3_N68) );
  OR2_X1 npu_inst_pe_1_3_3_U124 ( .A1(npu_inst_pe_1_3_3_int_q_acc_3_), .A2(
        npu_inst_pe_1_3_3_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_3_3_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_3_3_U123 ( .A(npu_inst_pe_1_3_3_sub_67_carry_4_), .B(
        npu_inst_pe_1_3_3_int_q_acc_4_), .ZN(npu_inst_pe_1_3_3_N69) );
  OR2_X1 npu_inst_pe_1_3_3_U122 ( .A1(npu_inst_pe_1_3_3_int_q_acc_4_), .A2(
        npu_inst_pe_1_3_3_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_3_3_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_3_3_U121 ( .A(npu_inst_pe_1_3_3_sub_67_carry_5_), .B(
        npu_inst_pe_1_3_3_int_q_acc_5_), .ZN(npu_inst_pe_1_3_3_N70) );
  OR2_X1 npu_inst_pe_1_3_3_U120 ( .A1(npu_inst_pe_1_3_3_int_q_acc_5_), .A2(
        npu_inst_pe_1_3_3_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_3_3_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_3_3_U119 ( .A(npu_inst_pe_1_3_3_sub_67_carry_6_), .B(
        npu_inst_pe_1_3_3_int_q_acc_6_), .ZN(npu_inst_pe_1_3_3_N71) );
  OR2_X1 npu_inst_pe_1_3_3_U118 ( .A1(npu_inst_pe_1_3_3_int_q_acc_6_), .A2(
        npu_inst_pe_1_3_3_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_3_3_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_3_3_U117 ( .A(npu_inst_pe_1_3_3_int_q_acc_7_), .B(
        npu_inst_pe_1_3_3_sub_67_carry_7_), .ZN(npu_inst_pe_1_3_3_N72) );
  INV_X1 npu_inst_pe_1_3_3_U116 ( .A(npu_inst_n78), .ZN(npu_inst_pe_1_3_3_n7)
         );
  INV_X1 npu_inst_pe_1_3_3_U115 ( .A(npu_inst_pe_1_3_3_n7), .ZN(
        npu_inst_pe_1_3_3_n6) );
  INV_X1 npu_inst_pe_1_3_3_U114 ( .A(npu_inst_n57), .ZN(npu_inst_pe_1_3_3_n3)
         );
  AOI22_X1 npu_inst_pe_1_3_3_U113 ( .A1(npu_inst_int_data_y_4__3__0_), .A2(
        npu_inst_pe_1_3_3_n58), .B1(npu_inst_pe_1_3_3_n119), .B2(
        npu_inst_pe_1_3_3_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_3_3_n57) );
  INV_X1 npu_inst_pe_1_3_3_U112 ( .A(npu_inst_pe_1_3_3_n57), .ZN(
        npu_inst_pe_1_3_3_n108) );
  AOI22_X1 npu_inst_pe_1_3_3_U111 ( .A1(npu_inst_int_data_y_4__3__0_), .A2(
        npu_inst_pe_1_3_3_n54), .B1(npu_inst_pe_1_3_3_n118), .B2(
        npu_inst_pe_1_3_3_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_3_3_n53) );
  INV_X1 npu_inst_pe_1_3_3_U110 ( .A(npu_inst_pe_1_3_3_n53), .ZN(
        npu_inst_pe_1_3_3_n109) );
  AOI22_X1 npu_inst_pe_1_3_3_U107 ( .A1(npu_inst_int_data_y_4__3__0_), .A2(
        npu_inst_pe_1_3_3_n50), .B1(npu_inst_pe_1_3_3_n117), .B2(
        npu_inst_pe_1_3_3_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_3_3_n49) );
  INV_X1 npu_inst_pe_1_3_3_U106 ( .A(npu_inst_pe_1_3_3_n49), .ZN(
        npu_inst_pe_1_3_3_n110) );
  AOI22_X1 npu_inst_pe_1_3_3_U105 ( .A1(npu_inst_int_data_y_4__3__0_), .A2(
        npu_inst_pe_1_3_3_n46), .B1(npu_inst_pe_1_3_3_n116), .B2(
        npu_inst_pe_1_3_3_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_3_3_n45) );
  INV_X1 npu_inst_pe_1_3_3_U104 ( .A(npu_inst_pe_1_3_3_n45), .ZN(
        npu_inst_pe_1_3_3_n111) );
  AOI22_X1 npu_inst_pe_1_3_3_U103 ( .A1(npu_inst_int_data_y_4__3__0_), .A2(
        npu_inst_pe_1_3_3_n42), .B1(npu_inst_pe_1_3_3_n115), .B2(
        npu_inst_pe_1_3_3_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_3_3_n41) );
  INV_X1 npu_inst_pe_1_3_3_U102 ( .A(npu_inst_pe_1_3_3_n41), .ZN(
        npu_inst_pe_1_3_3_n112) );
  AOI22_X1 npu_inst_pe_1_3_3_U101 ( .A1(npu_inst_int_data_y_4__3__1_), .A2(
        npu_inst_pe_1_3_3_n58), .B1(npu_inst_pe_1_3_3_n119), .B2(
        npu_inst_pe_1_3_3_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_3_3_n59) );
  INV_X1 npu_inst_pe_1_3_3_U100 ( .A(npu_inst_pe_1_3_3_n59), .ZN(
        npu_inst_pe_1_3_3_n102) );
  AOI22_X1 npu_inst_pe_1_3_3_U99 ( .A1(npu_inst_int_data_y_4__3__1_), .A2(
        npu_inst_pe_1_3_3_n54), .B1(npu_inst_pe_1_3_3_n118), .B2(
        npu_inst_pe_1_3_3_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_3_3_n55) );
  INV_X1 npu_inst_pe_1_3_3_U98 ( .A(npu_inst_pe_1_3_3_n55), .ZN(
        npu_inst_pe_1_3_3_n103) );
  AOI22_X1 npu_inst_pe_1_3_3_U97 ( .A1(npu_inst_int_data_y_4__3__1_), .A2(
        npu_inst_pe_1_3_3_n50), .B1(npu_inst_pe_1_3_3_n117), .B2(
        npu_inst_pe_1_3_3_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_3_3_n51) );
  INV_X1 npu_inst_pe_1_3_3_U96 ( .A(npu_inst_pe_1_3_3_n51), .ZN(
        npu_inst_pe_1_3_3_n104) );
  AOI22_X1 npu_inst_pe_1_3_3_U95 ( .A1(npu_inst_int_data_y_4__3__1_), .A2(
        npu_inst_pe_1_3_3_n46), .B1(npu_inst_pe_1_3_3_n116), .B2(
        npu_inst_pe_1_3_3_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_3_3_n47) );
  INV_X1 npu_inst_pe_1_3_3_U94 ( .A(npu_inst_pe_1_3_3_n47), .ZN(
        npu_inst_pe_1_3_3_n105) );
  AOI22_X1 npu_inst_pe_1_3_3_U93 ( .A1(npu_inst_int_data_y_4__3__1_), .A2(
        npu_inst_pe_1_3_3_n42), .B1(npu_inst_pe_1_3_3_n115), .B2(
        npu_inst_pe_1_3_3_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_3_3_n43) );
  INV_X1 npu_inst_pe_1_3_3_U92 ( .A(npu_inst_pe_1_3_3_n43), .ZN(
        npu_inst_pe_1_3_3_n106) );
  AOI22_X1 npu_inst_pe_1_3_3_U91 ( .A1(npu_inst_pe_1_3_3_n38), .A2(
        npu_inst_int_data_y_4__3__1_), .B1(npu_inst_pe_1_3_3_n114), .B2(
        npu_inst_pe_1_3_3_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_3_3_n39) );
  INV_X1 npu_inst_pe_1_3_3_U90 ( .A(npu_inst_pe_1_3_3_n39), .ZN(
        npu_inst_pe_1_3_3_n107) );
  AOI22_X1 npu_inst_pe_1_3_3_U89 ( .A1(npu_inst_pe_1_3_3_n38), .A2(
        npu_inst_int_data_y_4__3__0_), .B1(npu_inst_pe_1_3_3_n114), .B2(
        npu_inst_pe_1_3_3_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_3_3_n37) );
  INV_X1 npu_inst_pe_1_3_3_U88 ( .A(npu_inst_pe_1_3_3_n37), .ZN(
        npu_inst_pe_1_3_3_n113) );
  NAND2_X1 npu_inst_pe_1_3_3_U87 ( .A1(npu_inst_pe_1_3_3_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_3_3_n60), .ZN(npu_inst_pe_1_3_3_n74) );
  OAI21_X1 npu_inst_pe_1_3_3_U86 ( .B1(npu_inst_pe_1_3_3_n63), .B2(
        npu_inst_pe_1_3_3_n60), .A(npu_inst_pe_1_3_3_n74), .ZN(
        npu_inst_pe_1_3_3_n97) );
  NAND2_X1 npu_inst_pe_1_3_3_U85 ( .A1(npu_inst_pe_1_3_3_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_3_3_n60), .ZN(npu_inst_pe_1_3_3_n73) );
  OAI21_X1 npu_inst_pe_1_3_3_U84 ( .B1(npu_inst_pe_1_3_3_n61), .B2(
        npu_inst_pe_1_3_3_n60), .A(npu_inst_pe_1_3_3_n73), .ZN(
        npu_inst_pe_1_3_3_n96) );
  NAND2_X1 npu_inst_pe_1_3_3_U83 ( .A1(npu_inst_pe_1_3_3_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_3_3_n56), .ZN(npu_inst_pe_1_3_3_n72) );
  OAI21_X1 npu_inst_pe_1_3_3_U82 ( .B1(npu_inst_pe_1_3_3_n63), .B2(
        npu_inst_pe_1_3_3_n56), .A(npu_inst_pe_1_3_3_n72), .ZN(
        npu_inst_pe_1_3_3_n95) );
  NAND2_X1 npu_inst_pe_1_3_3_U81 ( .A1(npu_inst_pe_1_3_3_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_3_3_n56), .ZN(npu_inst_pe_1_3_3_n71) );
  OAI21_X1 npu_inst_pe_1_3_3_U80 ( .B1(npu_inst_pe_1_3_3_n61), .B2(
        npu_inst_pe_1_3_3_n56), .A(npu_inst_pe_1_3_3_n71), .ZN(
        npu_inst_pe_1_3_3_n94) );
  NAND2_X1 npu_inst_pe_1_3_3_U79 ( .A1(npu_inst_pe_1_3_3_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_3_3_n52), .ZN(npu_inst_pe_1_3_3_n70) );
  OAI21_X1 npu_inst_pe_1_3_3_U78 ( .B1(npu_inst_pe_1_3_3_n63), .B2(
        npu_inst_pe_1_3_3_n52), .A(npu_inst_pe_1_3_3_n70), .ZN(
        npu_inst_pe_1_3_3_n93) );
  NAND2_X1 npu_inst_pe_1_3_3_U77 ( .A1(npu_inst_pe_1_3_3_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_3_3_n52), .ZN(npu_inst_pe_1_3_3_n69) );
  OAI21_X1 npu_inst_pe_1_3_3_U76 ( .B1(npu_inst_pe_1_3_3_n61), .B2(
        npu_inst_pe_1_3_3_n52), .A(npu_inst_pe_1_3_3_n69), .ZN(
        npu_inst_pe_1_3_3_n92) );
  NAND2_X1 npu_inst_pe_1_3_3_U75 ( .A1(npu_inst_pe_1_3_3_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_3_3_n48), .ZN(npu_inst_pe_1_3_3_n68) );
  OAI21_X1 npu_inst_pe_1_3_3_U74 ( .B1(npu_inst_pe_1_3_3_n63), .B2(
        npu_inst_pe_1_3_3_n48), .A(npu_inst_pe_1_3_3_n68), .ZN(
        npu_inst_pe_1_3_3_n91) );
  NAND2_X1 npu_inst_pe_1_3_3_U73 ( .A1(npu_inst_pe_1_3_3_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_3_3_n48), .ZN(npu_inst_pe_1_3_3_n67) );
  OAI21_X1 npu_inst_pe_1_3_3_U72 ( .B1(npu_inst_pe_1_3_3_n61), .B2(
        npu_inst_pe_1_3_3_n48), .A(npu_inst_pe_1_3_3_n67), .ZN(
        npu_inst_pe_1_3_3_n90) );
  NAND2_X1 npu_inst_pe_1_3_3_U71 ( .A1(npu_inst_pe_1_3_3_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_3_3_n44), .ZN(npu_inst_pe_1_3_3_n66) );
  OAI21_X1 npu_inst_pe_1_3_3_U70 ( .B1(npu_inst_pe_1_3_3_n63), .B2(
        npu_inst_pe_1_3_3_n44), .A(npu_inst_pe_1_3_3_n66), .ZN(
        npu_inst_pe_1_3_3_n89) );
  NAND2_X1 npu_inst_pe_1_3_3_U69 ( .A1(npu_inst_pe_1_3_3_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_3_3_n44), .ZN(npu_inst_pe_1_3_3_n65) );
  OAI21_X1 npu_inst_pe_1_3_3_U68 ( .B1(npu_inst_pe_1_3_3_n61), .B2(
        npu_inst_pe_1_3_3_n44), .A(npu_inst_pe_1_3_3_n65), .ZN(
        npu_inst_pe_1_3_3_n88) );
  NAND2_X1 npu_inst_pe_1_3_3_U67 ( .A1(npu_inst_pe_1_3_3_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_3_3_n40), .ZN(npu_inst_pe_1_3_3_n64) );
  OAI21_X1 npu_inst_pe_1_3_3_U66 ( .B1(npu_inst_pe_1_3_3_n63), .B2(
        npu_inst_pe_1_3_3_n40), .A(npu_inst_pe_1_3_3_n64), .ZN(
        npu_inst_pe_1_3_3_n87) );
  NAND2_X1 npu_inst_pe_1_3_3_U65 ( .A1(npu_inst_pe_1_3_3_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_3_3_n40), .ZN(npu_inst_pe_1_3_3_n62) );
  OAI21_X1 npu_inst_pe_1_3_3_U64 ( .B1(npu_inst_pe_1_3_3_n61), .B2(
        npu_inst_pe_1_3_3_n40), .A(npu_inst_pe_1_3_3_n62), .ZN(
        npu_inst_pe_1_3_3_n86) );
  AND2_X1 npu_inst_pe_1_3_3_U63 ( .A1(npu_inst_pe_1_3_3_N93), .A2(npu_inst_n57), .ZN(npu_inst_int_data_y_3__3__0_) );
  AND2_X1 npu_inst_pe_1_3_3_U62 ( .A1(npu_inst_n57), .A2(npu_inst_pe_1_3_3_N94), .ZN(npu_inst_int_data_y_3__3__1_) );
  NOR3_X1 npu_inst_pe_1_3_3_U61 ( .A1(npu_inst_pe_1_3_3_n26), .A2(npu_inst_n57), .A3(npu_inst_int_ckg[36]), .ZN(npu_inst_pe_1_3_3_n85) );
  OR2_X1 npu_inst_pe_1_3_3_U60 ( .A1(npu_inst_pe_1_3_3_n85), .A2(
        npu_inst_pe_1_3_3_n2), .ZN(npu_inst_pe_1_3_3_N84) );
  AND2_X1 npu_inst_pe_1_3_3_U59 ( .A1(npu_inst_pe_1_3_3_int_q_acc_0_), .A2(
        npu_inst_pe_1_3_3_n1), .ZN(npu_inst_int_data_res_3__3__0_) );
  AND2_X1 npu_inst_pe_1_3_3_U58 ( .A1(npu_inst_pe_1_3_3_n2), .A2(
        npu_inst_pe_1_3_3_int_q_acc_7_), .ZN(npu_inst_int_data_res_3__3__7_)
         );
  AND2_X1 npu_inst_pe_1_3_3_U57 ( .A1(npu_inst_pe_1_3_3_int_q_acc_1_), .A2(
        npu_inst_pe_1_3_3_n1), .ZN(npu_inst_int_data_res_3__3__1_) );
  AND2_X1 npu_inst_pe_1_3_3_U56 ( .A1(npu_inst_pe_1_3_3_int_q_acc_2_), .A2(
        npu_inst_pe_1_3_3_n1), .ZN(npu_inst_int_data_res_3__3__2_) );
  AND2_X1 npu_inst_pe_1_3_3_U55 ( .A1(npu_inst_pe_1_3_3_int_q_acc_3_), .A2(
        npu_inst_pe_1_3_3_n2), .ZN(npu_inst_int_data_res_3__3__3_) );
  AND2_X1 npu_inst_pe_1_3_3_U54 ( .A1(npu_inst_pe_1_3_3_int_q_acc_4_), .A2(
        npu_inst_pe_1_3_3_n2), .ZN(npu_inst_int_data_res_3__3__4_) );
  AND2_X1 npu_inst_pe_1_3_3_U53 ( .A1(npu_inst_pe_1_3_3_int_q_acc_5_), .A2(
        npu_inst_pe_1_3_3_n2), .ZN(npu_inst_int_data_res_3__3__5_) );
  AND2_X1 npu_inst_pe_1_3_3_U52 ( .A1(npu_inst_pe_1_3_3_int_q_acc_6_), .A2(
        npu_inst_pe_1_3_3_n2), .ZN(npu_inst_int_data_res_3__3__6_) );
  AOI222_X1 npu_inst_pe_1_3_3_U51 ( .A1(npu_inst_int_data_res_4__3__0_), .A2(
        npu_inst_pe_1_3_3_n1), .B1(npu_inst_pe_1_3_3_N73), .B2(
        npu_inst_pe_1_3_3_n76), .C1(npu_inst_pe_1_3_3_N65), .C2(
        npu_inst_pe_1_3_3_n77), .ZN(npu_inst_pe_1_3_3_n84) );
  INV_X1 npu_inst_pe_1_3_3_U50 ( .A(npu_inst_pe_1_3_3_n84), .ZN(
        npu_inst_pe_1_3_3_n101) );
  AOI222_X1 npu_inst_pe_1_3_3_U49 ( .A1(npu_inst_int_data_res_4__3__7_), .A2(
        npu_inst_pe_1_3_3_n1), .B1(npu_inst_pe_1_3_3_N80), .B2(
        npu_inst_pe_1_3_3_n76), .C1(npu_inst_pe_1_3_3_N72), .C2(
        npu_inst_pe_1_3_3_n77), .ZN(npu_inst_pe_1_3_3_n75) );
  INV_X1 npu_inst_pe_1_3_3_U48 ( .A(npu_inst_pe_1_3_3_n75), .ZN(
        npu_inst_pe_1_3_3_n33) );
  AOI222_X1 npu_inst_pe_1_3_3_U47 ( .A1(npu_inst_int_data_res_4__3__1_), .A2(
        npu_inst_pe_1_3_3_n1), .B1(npu_inst_pe_1_3_3_N74), .B2(
        npu_inst_pe_1_3_3_n76), .C1(npu_inst_pe_1_3_3_N66), .C2(
        npu_inst_pe_1_3_3_n77), .ZN(npu_inst_pe_1_3_3_n83) );
  INV_X1 npu_inst_pe_1_3_3_U46 ( .A(npu_inst_pe_1_3_3_n83), .ZN(
        npu_inst_pe_1_3_3_n100) );
  AOI222_X1 npu_inst_pe_1_3_3_U45 ( .A1(npu_inst_int_data_res_4__3__2_), .A2(
        npu_inst_pe_1_3_3_n1), .B1(npu_inst_pe_1_3_3_N75), .B2(
        npu_inst_pe_1_3_3_n76), .C1(npu_inst_pe_1_3_3_N67), .C2(
        npu_inst_pe_1_3_3_n77), .ZN(npu_inst_pe_1_3_3_n82) );
  INV_X1 npu_inst_pe_1_3_3_U44 ( .A(npu_inst_pe_1_3_3_n82), .ZN(
        npu_inst_pe_1_3_3_n99) );
  AOI222_X1 npu_inst_pe_1_3_3_U43 ( .A1(npu_inst_int_data_res_4__3__3_), .A2(
        npu_inst_pe_1_3_3_n1), .B1(npu_inst_pe_1_3_3_N76), .B2(
        npu_inst_pe_1_3_3_n76), .C1(npu_inst_pe_1_3_3_N68), .C2(
        npu_inst_pe_1_3_3_n77), .ZN(npu_inst_pe_1_3_3_n81) );
  INV_X1 npu_inst_pe_1_3_3_U42 ( .A(npu_inst_pe_1_3_3_n81), .ZN(
        npu_inst_pe_1_3_3_n98) );
  AOI222_X1 npu_inst_pe_1_3_3_U41 ( .A1(npu_inst_int_data_res_4__3__4_), .A2(
        npu_inst_pe_1_3_3_n1), .B1(npu_inst_pe_1_3_3_N77), .B2(
        npu_inst_pe_1_3_3_n76), .C1(npu_inst_pe_1_3_3_N69), .C2(
        npu_inst_pe_1_3_3_n77), .ZN(npu_inst_pe_1_3_3_n80) );
  INV_X1 npu_inst_pe_1_3_3_U40 ( .A(npu_inst_pe_1_3_3_n80), .ZN(
        npu_inst_pe_1_3_3_n36) );
  AOI222_X1 npu_inst_pe_1_3_3_U39 ( .A1(npu_inst_int_data_res_4__3__5_), .A2(
        npu_inst_pe_1_3_3_n1), .B1(npu_inst_pe_1_3_3_N78), .B2(
        npu_inst_pe_1_3_3_n76), .C1(npu_inst_pe_1_3_3_N70), .C2(
        npu_inst_pe_1_3_3_n77), .ZN(npu_inst_pe_1_3_3_n79) );
  INV_X1 npu_inst_pe_1_3_3_U38 ( .A(npu_inst_pe_1_3_3_n79), .ZN(
        npu_inst_pe_1_3_3_n35) );
  AOI222_X1 npu_inst_pe_1_3_3_U37 ( .A1(npu_inst_int_data_res_4__3__6_), .A2(
        npu_inst_pe_1_3_3_n1), .B1(npu_inst_pe_1_3_3_N79), .B2(
        npu_inst_pe_1_3_3_n76), .C1(npu_inst_pe_1_3_3_N71), .C2(
        npu_inst_pe_1_3_3_n77), .ZN(npu_inst_pe_1_3_3_n78) );
  INV_X1 npu_inst_pe_1_3_3_U36 ( .A(npu_inst_pe_1_3_3_n78), .ZN(
        npu_inst_pe_1_3_3_n34) );
  INV_X1 npu_inst_pe_1_3_3_U35 ( .A(npu_inst_pe_1_3_3_int_data_1_), .ZN(
        npu_inst_pe_1_3_3_n14) );
  AND2_X1 npu_inst_pe_1_3_3_U34 ( .A1(npu_inst_int_data_x_3__3__1_), .A2(
        npu_inst_pe_1_3_3_int_q_weight_1_), .ZN(npu_inst_pe_1_3_3_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_3_3_U33 ( .A1(npu_inst_int_data_x_3__3__0_), .A2(
        npu_inst_pe_1_3_3_int_q_weight_1_), .ZN(npu_inst_pe_1_3_3_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_3_3_U32 ( .A1(npu_inst_n57), .A2(
        npu_inst_int_data_y_4__3__1_), .B1(npu_inst_pe_1_3_3_n3), .B2(
        npu_inst_int_data_x_3__4__1_), .ZN(npu_inst_pe_1_3_3_n63) );
  AOI22_X1 npu_inst_pe_1_3_3_U31 ( .A1(npu_inst_n57), .A2(
        npu_inst_int_data_y_4__3__0_), .B1(npu_inst_pe_1_3_3_n3), .B2(
        npu_inst_int_data_x_3__4__0_), .ZN(npu_inst_pe_1_3_3_n61) );
  INV_X1 npu_inst_pe_1_3_3_U30 ( .A(npu_inst_pe_1_3_3_int_data_0_), .ZN(
        npu_inst_pe_1_3_3_n13) );
  INV_X1 npu_inst_pe_1_3_3_U29 ( .A(npu_inst_n70), .ZN(npu_inst_pe_1_3_3_n5)
         );
  OR3_X1 npu_inst_pe_1_3_3_U28 ( .A1(npu_inst_pe_1_3_3_n6), .A2(
        npu_inst_pe_1_3_3_n8), .A3(npu_inst_pe_1_3_3_n5), .ZN(
        npu_inst_pe_1_3_3_n56) );
  OR3_X1 npu_inst_pe_1_3_3_U27 ( .A1(npu_inst_pe_1_3_3_n5), .A2(
        npu_inst_pe_1_3_3_n8), .A3(npu_inst_pe_1_3_3_n7), .ZN(
        npu_inst_pe_1_3_3_n48) );
  INV_X1 npu_inst_pe_1_3_3_U26 ( .A(npu_inst_pe_1_3_3_n5), .ZN(
        npu_inst_pe_1_3_3_n4) );
  OR3_X1 npu_inst_pe_1_3_3_U25 ( .A1(npu_inst_pe_1_3_3_n4), .A2(
        npu_inst_pe_1_3_3_n8), .A3(npu_inst_pe_1_3_3_n7), .ZN(
        npu_inst_pe_1_3_3_n52) );
  OR3_X1 npu_inst_pe_1_3_3_U24 ( .A1(npu_inst_pe_1_3_3_n6), .A2(
        npu_inst_pe_1_3_3_n8), .A3(npu_inst_pe_1_3_3_n4), .ZN(
        npu_inst_pe_1_3_3_n60) );
  NOR2_X1 npu_inst_pe_1_3_3_U23 ( .A1(npu_inst_pe_1_3_3_n60), .A2(
        npu_inst_pe_1_3_3_n3), .ZN(npu_inst_pe_1_3_3_n58) );
  NOR2_X1 npu_inst_pe_1_3_3_U22 ( .A1(npu_inst_pe_1_3_3_n56), .A2(
        npu_inst_pe_1_3_3_n3), .ZN(npu_inst_pe_1_3_3_n54) );
  NOR2_X1 npu_inst_pe_1_3_3_U21 ( .A1(npu_inst_pe_1_3_3_n52), .A2(
        npu_inst_pe_1_3_3_n3), .ZN(npu_inst_pe_1_3_3_n50) );
  NOR2_X1 npu_inst_pe_1_3_3_U20 ( .A1(npu_inst_pe_1_3_3_n48), .A2(
        npu_inst_pe_1_3_3_n3), .ZN(npu_inst_pe_1_3_3_n46) );
  NOR2_X1 npu_inst_pe_1_3_3_U19 ( .A1(npu_inst_pe_1_3_3_n40), .A2(
        npu_inst_pe_1_3_3_n3), .ZN(npu_inst_pe_1_3_3_n38) );
  NOR2_X1 npu_inst_pe_1_3_3_U18 ( .A1(npu_inst_pe_1_3_3_n44), .A2(
        npu_inst_pe_1_3_3_n3), .ZN(npu_inst_pe_1_3_3_n42) );
  BUF_X1 npu_inst_pe_1_3_3_U17 ( .A(npu_inst_n101), .Z(npu_inst_pe_1_3_3_n8)
         );
  INV_X1 npu_inst_pe_1_3_3_U16 ( .A(npu_inst_n125), .ZN(npu_inst_pe_1_3_3_n12)
         );
  INV_X1 npu_inst_pe_1_3_3_U15 ( .A(npu_inst_pe_1_3_3_n38), .ZN(
        npu_inst_pe_1_3_3_n114) );
  INV_X1 npu_inst_pe_1_3_3_U14 ( .A(npu_inst_pe_1_3_3_n58), .ZN(
        npu_inst_pe_1_3_3_n119) );
  INV_X1 npu_inst_pe_1_3_3_U13 ( .A(npu_inst_pe_1_3_3_n54), .ZN(
        npu_inst_pe_1_3_3_n118) );
  INV_X1 npu_inst_pe_1_3_3_U12 ( .A(npu_inst_pe_1_3_3_n50), .ZN(
        npu_inst_pe_1_3_3_n117) );
  INV_X1 npu_inst_pe_1_3_3_U11 ( .A(npu_inst_pe_1_3_3_n46), .ZN(
        npu_inst_pe_1_3_3_n116) );
  INV_X1 npu_inst_pe_1_3_3_U10 ( .A(npu_inst_pe_1_3_3_n42), .ZN(
        npu_inst_pe_1_3_3_n115) );
  BUF_X1 npu_inst_pe_1_3_3_U9 ( .A(npu_inst_n25), .Z(npu_inst_pe_1_3_3_n2) );
  BUF_X1 npu_inst_pe_1_3_3_U8 ( .A(npu_inst_n25), .Z(npu_inst_pe_1_3_3_n1) );
  BUF_X1 npu_inst_pe_1_3_3_U7 ( .A(npu_inst_pe_1_3_3_n12), .Z(
        npu_inst_pe_1_3_3_n11) );
  BUF_X1 npu_inst_pe_1_3_3_U6 ( .A(npu_inst_pe_1_3_3_n12), .Z(
        npu_inst_pe_1_3_3_n10) );
  BUF_X1 npu_inst_pe_1_3_3_U5 ( .A(npu_inst_pe_1_3_3_n12), .Z(
        npu_inst_pe_1_3_3_n9) );
  NOR2_X1 npu_inst_pe_1_3_3_U4 ( .A1(npu_inst_pe_1_3_3_int_q_weight_0_), .A2(
        npu_inst_pe_1_3_3_n1), .ZN(npu_inst_pe_1_3_3_n76) );
  NOR2_X1 npu_inst_pe_1_3_3_U3 ( .A1(npu_inst_pe_1_3_3_n27), .A2(
        npu_inst_pe_1_3_3_n1), .ZN(npu_inst_pe_1_3_3_n77) );
  FA_X1 npu_inst_pe_1_3_3_sub_67_U2_1 ( .A(npu_inst_pe_1_3_3_int_q_acc_1_), 
        .B(npu_inst_pe_1_3_3_n14), .CI(npu_inst_pe_1_3_3_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_3_3_sub_67_carry_2_), .S(npu_inst_pe_1_3_3_N66) );
  FA_X1 npu_inst_pe_1_3_3_add_69_U1_1 ( .A(npu_inst_pe_1_3_3_int_q_acc_1_), 
        .B(npu_inst_pe_1_3_3_int_data_1_), .CI(
        npu_inst_pe_1_3_3_add_69_carry_1_), .CO(
        npu_inst_pe_1_3_3_add_69_carry_2_), .S(npu_inst_pe_1_3_3_N74) );
  NAND3_X1 npu_inst_pe_1_3_3_U109 ( .A1(npu_inst_pe_1_3_3_n5), .A2(
        npu_inst_pe_1_3_3_n7), .A3(npu_inst_pe_1_3_3_n8), .ZN(
        npu_inst_pe_1_3_3_n44) );
  NAND3_X1 npu_inst_pe_1_3_3_U108 ( .A1(npu_inst_pe_1_3_3_n4), .A2(
        npu_inst_pe_1_3_3_n7), .A3(npu_inst_pe_1_3_3_n8), .ZN(
        npu_inst_pe_1_3_3_n40) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_3_3_n34), .CK(
        npu_inst_pe_1_3_3_net3941), .RN(npu_inst_pe_1_3_3_n9), .Q(
        npu_inst_pe_1_3_3_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_3_3_n35), .CK(
        npu_inst_pe_1_3_3_net3941), .RN(npu_inst_pe_1_3_3_n9), .Q(
        npu_inst_pe_1_3_3_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_3_3_n36), .CK(
        npu_inst_pe_1_3_3_net3941), .RN(npu_inst_pe_1_3_3_n9), .Q(
        npu_inst_pe_1_3_3_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_3_3_n98), .CK(
        npu_inst_pe_1_3_3_net3941), .RN(npu_inst_pe_1_3_3_n9), .Q(
        npu_inst_pe_1_3_3_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_3_3_n99), .CK(
        npu_inst_pe_1_3_3_net3941), .RN(npu_inst_pe_1_3_3_n9), .Q(
        npu_inst_pe_1_3_3_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_3_3_n100), 
        .CK(npu_inst_pe_1_3_3_net3941), .RN(npu_inst_pe_1_3_3_n9), .Q(
        npu_inst_pe_1_3_3_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_3_3_n33), .CK(
        npu_inst_pe_1_3_3_net3941), .RN(npu_inst_pe_1_3_3_n9), .Q(
        npu_inst_pe_1_3_3_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_3_3_n101), 
        .CK(npu_inst_pe_1_3_3_net3941), .RN(npu_inst_pe_1_3_3_n9), .Q(
        npu_inst_pe_1_3_3_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_weight_reg_0_ ( .D(npu_inst_n111), .CK(
        npu_inst_pe_1_3_3_net3947), .RN(npu_inst_pe_1_3_3_n9), .Q(
        npu_inst_pe_1_3_3_int_q_weight_0_), .QN(npu_inst_pe_1_3_3_n27) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_weight_reg_1_ ( .D(npu_inst_n117), .CK(
        npu_inst_pe_1_3_3_net3947), .RN(npu_inst_pe_1_3_3_n9), .Q(
        npu_inst_pe_1_3_3_int_q_weight_1_), .QN(npu_inst_pe_1_3_3_n26) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_3_3_n113), 
        .CK(npu_inst_pe_1_3_3_net3947), .RN(npu_inst_pe_1_3_3_n9), .Q(
        npu_inst_pe_1_3_3_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_3_3_n107), 
        .CK(npu_inst_pe_1_3_3_net3947), .RN(npu_inst_pe_1_3_3_n9), .Q(
        npu_inst_pe_1_3_3_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_3_3_n112), 
        .CK(npu_inst_pe_1_3_3_net3947), .RN(npu_inst_pe_1_3_3_n10), .Q(
        npu_inst_pe_1_3_3_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_3_3_n106), 
        .CK(npu_inst_pe_1_3_3_net3947), .RN(npu_inst_pe_1_3_3_n10), .Q(
        npu_inst_pe_1_3_3_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_3_3_n111), 
        .CK(npu_inst_pe_1_3_3_net3947), .RN(npu_inst_pe_1_3_3_n10), .Q(
        npu_inst_pe_1_3_3_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_3_3_n105), 
        .CK(npu_inst_pe_1_3_3_net3947), .RN(npu_inst_pe_1_3_3_n10), .Q(
        npu_inst_pe_1_3_3_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_3_3_n110), 
        .CK(npu_inst_pe_1_3_3_net3947), .RN(npu_inst_pe_1_3_3_n10), .Q(
        npu_inst_pe_1_3_3_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_3_3_n104), 
        .CK(npu_inst_pe_1_3_3_net3947), .RN(npu_inst_pe_1_3_3_n10), .Q(
        npu_inst_pe_1_3_3_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_3_3_n109), 
        .CK(npu_inst_pe_1_3_3_net3947), .RN(npu_inst_pe_1_3_3_n10), .Q(
        npu_inst_pe_1_3_3_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_3_3_n103), 
        .CK(npu_inst_pe_1_3_3_net3947), .RN(npu_inst_pe_1_3_3_n10), .Q(
        npu_inst_pe_1_3_3_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_3_3_n108), 
        .CK(npu_inst_pe_1_3_3_net3947), .RN(npu_inst_pe_1_3_3_n10), .Q(
        npu_inst_pe_1_3_3_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_3_3_n102), 
        .CK(npu_inst_pe_1_3_3_net3947), .RN(npu_inst_pe_1_3_3_n10), .Q(
        npu_inst_pe_1_3_3_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_3_3_n86), 
        .CK(npu_inst_pe_1_3_3_net3947), .RN(npu_inst_pe_1_3_3_n10), .Q(
        npu_inst_pe_1_3_3_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_3_3_n87), 
        .CK(npu_inst_pe_1_3_3_net3947), .RN(npu_inst_pe_1_3_3_n10), .Q(
        npu_inst_pe_1_3_3_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_3_3_n88), 
        .CK(npu_inst_pe_1_3_3_net3947), .RN(npu_inst_pe_1_3_3_n11), .Q(
        npu_inst_pe_1_3_3_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_3_3_n89), 
        .CK(npu_inst_pe_1_3_3_net3947), .RN(npu_inst_pe_1_3_3_n11), .Q(
        npu_inst_pe_1_3_3_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_3_3_n90), 
        .CK(npu_inst_pe_1_3_3_net3947), .RN(npu_inst_pe_1_3_3_n11), .Q(
        npu_inst_pe_1_3_3_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_3_3_n91), 
        .CK(npu_inst_pe_1_3_3_net3947), .RN(npu_inst_pe_1_3_3_n11), .Q(
        npu_inst_pe_1_3_3_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_3_3_n92), 
        .CK(npu_inst_pe_1_3_3_net3947), .RN(npu_inst_pe_1_3_3_n11), .Q(
        npu_inst_pe_1_3_3_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_3_3_n93), 
        .CK(npu_inst_pe_1_3_3_net3947), .RN(npu_inst_pe_1_3_3_n11), .Q(
        npu_inst_pe_1_3_3_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_3_3_n94), 
        .CK(npu_inst_pe_1_3_3_net3947), .RN(npu_inst_pe_1_3_3_n11), .Q(
        npu_inst_pe_1_3_3_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_3_3_n95), 
        .CK(npu_inst_pe_1_3_3_net3947), .RN(npu_inst_pe_1_3_3_n11), .Q(
        npu_inst_pe_1_3_3_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_3_3_n96), 
        .CK(npu_inst_pe_1_3_3_net3947), .RN(npu_inst_pe_1_3_3_n11), .Q(
        npu_inst_pe_1_3_3_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_3_3_n97), 
        .CK(npu_inst_pe_1_3_3_net3947), .RN(npu_inst_pe_1_3_3_n11), .Q(
        npu_inst_pe_1_3_3_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_3_3_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_3_3_N84), .SE(1'b0), .GCK(npu_inst_pe_1_3_3_net3941) );
  CLKGATETST_X1 npu_inst_pe_1_3_3_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n64), .SE(1'b0), .GCK(npu_inst_pe_1_3_3_net3947) );
  MUX2_X1 npu_inst_pe_1_3_4_U161 ( .A(npu_inst_pe_1_3_4_n31), .B(
        npu_inst_pe_1_3_4_n28), .S(npu_inst_pe_1_3_4_n7), .Z(
        npu_inst_pe_1_3_4_N93) );
  MUX2_X1 npu_inst_pe_1_3_4_U160 ( .A(npu_inst_pe_1_3_4_n30), .B(
        npu_inst_pe_1_3_4_n29), .S(npu_inst_n77), .Z(npu_inst_pe_1_3_4_n31) );
  MUX2_X1 npu_inst_pe_1_3_4_U159 ( .A(npu_inst_pe_1_3_4_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_3_4_int_q_reg_v_1__0_), .S(npu_inst_pe_1_3_4_n4), .Z(
        npu_inst_pe_1_3_4_n30) );
  MUX2_X1 npu_inst_pe_1_3_4_U158 ( .A(npu_inst_pe_1_3_4_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_3_4_int_q_reg_v_3__0_), .S(npu_inst_pe_1_3_4_n4), .Z(
        npu_inst_pe_1_3_4_n29) );
  MUX2_X1 npu_inst_pe_1_3_4_U157 ( .A(npu_inst_pe_1_3_4_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_3_4_int_q_reg_v_5__0_), .S(npu_inst_pe_1_3_4_n4), .Z(
        npu_inst_pe_1_3_4_n28) );
  MUX2_X1 npu_inst_pe_1_3_4_U156 ( .A(npu_inst_pe_1_3_4_n25), .B(
        npu_inst_pe_1_3_4_n22), .S(npu_inst_pe_1_3_4_n7), .Z(
        npu_inst_pe_1_3_4_N94) );
  MUX2_X1 npu_inst_pe_1_3_4_U155 ( .A(npu_inst_pe_1_3_4_n24), .B(
        npu_inst_pe_1_3_4_n23), .S(npu_inst_n77), .Z(npu_inst_pe_1_3_4_n25) );
  MUX2_X1 npu_inst_pe_1_3_4_U154 ( .A(npu_inst_pe_1_3_4_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_3_4_int_q_reg_v_1__1_), .S(npu_inst_pe_1_3_4_n4), .Z(
        npu_inst_pe_1_3_4_n24) );
  MUX2_X1 npu_inst_pe_1_3_4_U153 ( .A(npu_inst_pe_1_3_4_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_3_4_int_q_reg_v_3__1_), .S(npu_inst_pe_1_3_4_n4), .Z(
        npu_inst_pe_1_3_4_n23) );
  MUX2_X1 npu_inst_pe_1_3_4_U152 ( .A(npu_inst_pe_1_3_4_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_3_4_int_q_reg_v_5__1_), .S(npu_inst_pe_1_3_4_n4), .Z(
        npu_inst_pe_1_3_4_n22) );
  MUX2_X1 npu_inst_pe_1_3_4_U151 ( .A(npu_inst_pe_1_3_4_n21), .B(
        npu_inst_pe_1_3_4_n18), .S(npu_inst_pe_1_3_4_n7), .Z(
        npu_inst_int_data_x_3__4__1_) );
  MUX2_X1 npu_inst_pe_1_3_4_U150 ( .A(npu_inst_pe_1_3_4_n20), .B(
        npu_inst_pe_1_3_4_n19), .S(npu_inst_n77), .Z(npu_inst_pe_1_3_4_n21) );
  MUX2_X1 npu_inst_pe_1_3_4_U149 ( .A(npu_inst_pe_1_3_4_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_3_4_int_q_reg_h_1__1_), .S(npu_inst_pe_1_3_4_n4), .Z(
        npu_inst_pe_1_3_4_n20) );
  MUX2_X1 npu_inst_pe_1_3_4_U148 ( .A(npu_inst_pe_1_3_4_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_3_4_int_q_reg_h_3__1_), .S(npu_inst_pe_1_3_4_n4), .Z(
        npu_inst_pe_1_3_4_n19) );
  MUX2_X1 npu_inst_pe_1_3_4_U147 ( .A(npu_inst_pe_1_3_4_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_3_4_int_q_reg_h_5__1_), .S(npu_inst_pe_1_3_4_n4), .Z(
        npu_inst_pe_1_3_4_n18) );
  MUX2_X1 npu_inst_pe_1_3_4_U146 ( .A(npu_inst_pe_1_3_4_n17), .B(
        npu_inst_pe_1_3_4_n14), .S(npu_inst_pe_1_3_4_n7), .Z(
        npu_inst_int_data_x_3__4__0_) );
  MUX2_X1 npu_inst_pe_1_3_4_U145 ( .A(npu_inst_pe_1_3_4_n16), .B(
        npu_inst_pe_1_3_4_n15), .S(npu_inst_n77), .Z(npu_inst_pe_1_3_4_n17) );
  MUX2_X1 npu_inst_pe_1_3_4_U144 ( .A(npu_inst_pe_1_3_4_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_3_4_int_q_reg_h_1__0_), .S(npu_inst_pe_1_3_4_n4), .Z(
        npu_inst_pe_1_3_4_n16) );
  MUX2_X1 npu_inst_pe_1_3_4_U143 ( .A(npu_inst_pe_1_3_4_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_3_4_int_q_reg_h_3__0_), .S(npu_inst_pe_1_3_4_n4), .Z(
        npu_inst_pe_1_3_4_n15) );
  MUX2_X1 npu_inst_pe_1_3_4_U142 ( .A(npu_inst_pe_1_3_4_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_3_4_int_q_reg_h_5__0_), .S(npu_inst_pe_1_3_4_n4), .Z(
        npu_inst_pe_1_3_4_n14) );
  XOR2_X1 npu_inst_pe_1_3_4_U141 ( .A(npu_inst_pe_1_3_4_int_data_0_), .B(
        npu_inst_pe_1_3_4_int_q_acc_0_), .Z(npu_inst_pe_1_3_4_N73) );
  AND2_X1 npu_inst_pe_1_3_4_U140 ( .A1(npu_inst_pe_1_3_4_int_q_acc_0_), .A2(
        npu_inst_pe_1_3_4_int_data_0_), .ZN(npu_inst_pe_1_3_4_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_3_4_U139 ( .A(npu_inst_pe_1_3_4_int_q_acc_0_), .B(
        npu_inst_pe_1_3_4_n12), .ZN(npu_inst_pe_1_3_4_N65) );
  OR2_X1 npu_inst_pe_1_3_4_U138 ( .A1(npu_inst_pe_1_3_4_n12), .A2(
        npu_inst_pe_1_3_4_int_q_acc_0_), .ZN(npu_inst_pe_1_3_4_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_3_4_U137 ( .A(npu_inst_pe_1_3_4_int_q_acc_2_), .B(
        npu_inst_pe_1_3_4_add_69_carry_2_), .Z(npu_inst_pe_1_3_4_N75) );
  AND2_X1 npu_inst_pe_1_3_4_U136 ( .A1(npu_inst_pe_1_3_4_add_69_carry_2_), 
        .A2(npu_inst_pe_1_3_4_int_q_acc_2_), .ZN(
        npu_inst_pe_1_3_4_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_3_4_U135 ( .A(npu_inst_pe_1_3_4_int_q_acc_3_), .B(
        npu_inst_pe_1_3_4_add_69_carry_3_), .Z(npu_inst_pe_1_3_4_N76) );
  AND2_X1 npu_inst_pe_1_3_4_U134 ( .A1(npu_inst_pe_1_3_4_add_69_carry_3_), 
        .A2(npu_inst_pe_1_3_4_int_q_acc_3_), .ZN(
        npu_inst_pe_1_3_4_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_3_4_U133 ( .A(npu_inst_pe_1_3_4_int_q_acc_4_), .B(
        npu_inst_pe_1_3_4_add_69_carry_4_), .Z(npu_inst_pe_1_3_4_N77) );
  AND2_X1 npu_inst_pe_1_3_4_U132 ( .A1(npu_inst_pe_1_3_4_add_69_carry_4_), 
        .A2(npu_inst_pe_1_3_4_int_q_acc_4_), .ZN(
        npu_inst_pe_1_3_4_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_3_4_U131 ( .A(npu_inst_pe_1_3_4_int_q_acc_5_), .B(
        npu_inst_pe_1_3_4_add_69_carry_5_), .Z(npu_inst_pe_1_3_4_N78) );
  AND2_X1 npu_inst_pe_1_3_4_U130 ( .A1(npu_inst_pe_1_3_4_add_69_carry_5_), 
        .A2(npu_inst_pe_1_3_4_int_q_acc_5_), .ZN(
        npu_inst_pe_1_3_4_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_3_4_U129 ( .A(npu_inst_pe_1_3_4_int_q_acc_6_), .B(
        npu_inst_pe_1_3_4_add_69_carry_6_), .Z(npu_inst_pe_1_3_4_N79) );
  AND2_X1 npu_inst_pe_1_3_4_U128 ( .A1(npu_inst_pe_1_3_4_add_69_carry_6_), 
        .A2(npu_inst_pe_1_3_4_int_q_acc_6_), .ZN(
        npu_inst_pe_1_3_4_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_3_4_U127 ( .A(npu_inst_pe_1_3_4_int_q_acc_7_), .B(
        npu_inst_pe_1_3_4_add_69_carry_7_), .Z(npu_inst_pe_1_3_4_N80) );
  XNOR2_X1 npu_inst_pe_1_3_4_U126 ( .A(npu_inst_pe_1_3_4_sub_67_carry_2_), .B(
        npu_inst_pe_1_3_4_int_q_acc_2_), .ZN(npu_inst_pe_1_3_4_N67) );
  OR2_X1 npu_inst_pe_1_3_4_U125 ( .A1(npu_inst_pe_1_3_4_int_q_acc_2_), .A2(
        npu_inst_pe_1_3_4_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_3_4_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_3_4_U124 ( .A(npu_inst_pe_1_3_4_sub_67_carry_3_), .B(
        npu_inst_pe_1_3_4_int_q_acc_3_), .ZN(npu_inst_pe_1_3_4_N68) );
  OR2_X1 npu_inst_pe_1_3_4_U123 ( .A1(npu_inst_pe_1_3_4_int_q_acc_3_), .A2(
        npu_inst_pe_1_3_4_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_3_4_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_3_4_U122 ( .A(npu_inst_pe_1_3_4_sub_67_carry_4_), .B(
        npu_inst_pe_1_3_4_int_q_acc_4_), .ZN(npu_inst_pe_1_3_4_N69) );
  OR2_X1 npu_inst_pe_1_3_4_U121 ( .A1(npu_inst_pe_1_3_4_int_q_acc_4_), .A2(
        npu_inst_pe_1_3_4_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_3_4_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_3_4_U120 ( .A(npu_inst_pe_1_3_4_sub_67_carry_5_), .B(
        npu_inst_pe_1_3_4_int_q_acc_5_), .ZN(npu_inst_pe_1_3_4_N70) );
  OR2_X1 npu_inst_pe_1_3_4_U119 ( .A1(npu_inst_pe_1_3_4_int_q_acc_5_), .A2(
        npu_inst_pe_1_3_4_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_3_4_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_3_4_U118 ( .A(npu_inst_pe_1_3_4_sub_67_carry_6_), .B(
        npu_inst_pe_1_3_4_int_q_acc_6_), .ZN(npu_inst_pe_1_3_4_N71) );
  OR2_X1 npu_inst_pe_1_3_4_U117 ( .A1(npu_inst_pe_1_3_4_int_q_acc_6_), .A2(
        npu_inst_pe_1_3_4_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_3_4_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_3_4_U116 ( .A(npu_inst_pe_1_3_4_int_q_acc_7_), .B(
        npu_inst_pe_1_3_4_sub_67_carry_7_), .ZN(npu_inst_pe_1_3_4_N72) );
  INV_X1 npu_inst_pe_1_3_4_U115 ( .A(npu_inst_n77), .ZN(npu_inst_pe_1_3_4_n6)
         );
  INV_X1 npu_inst_pe_1_3_4_U114 ( .A(npu_inst_n57), .ZN(npu_inst_pe_1_3_4_n3)
         );
  AOI22_X1 npu_inst_pe_1_3_4_U113 ( .A1(npu_inst_int_data_y_4__4__0_), .A2(
        npu_inst_pe_1_3_4_n58), .B1(npu_inst_pe_1_3_4_n118), .B2(
        npu_inst_pe_1_3_4_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_3_4_n57) );
  INV_X1 npu_inst_pe_1_3_4_U112 ( .A(npu_inst_pe_1_3_4_n57), .ZN(
        npu_inst_pe_1_3_4_n107) );
  AOI22_X1 npu_inst_pe_1_3_4_U111 ( .A1(npu_inst_int_data_y_4__4__0_), .A2(
        npu_inst_pe_1_3_4_n54), .B1(npu_inst_pe_1_3_4_n117), .B2(
        npu_inst_pe_1_3_4_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_3_4_n53) );
  INV_X1 npu_inst_pe_1_3_4_U110 ( .A(npu_inst_pe_1_3_4_n53), .ZN(
        npu_inst_pe_1_3_4_n108) );
  AOI22_X1 npu_inst_pe_1_3_4_U107 ( .A1(npu_inst_int_data_y_4__4__0_), .A2(
        npu_inst_pe_1_3_4_n50), .B1(npu_inst_pe_1_3_4_n116), .B2(
        npu_inst_pe_1_3_4_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_3_4_n49) );
  INV_X1 npu_inst_pe_1_3_4_U106 ( .A(npu_inst_pe_1_3_4_n49), .ZN(
        npu_inst_pe_1_3_4_n109) );
  AOI22_X1 npu_inst_pe_1_3_4_U105 ( .A1(npu_inst_int_data_y_4__4__0_), .A2(
        npu_inst_pe_1_3_4_n46), .B1(npu_inst_pe_1_3_4_n115), .B2(
        npu_inst_pe_1_3_4_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_3_4_n45) );
  INV_X1 npu_inst_pe_1_3_4_U104 ( .A(npu_inst_pe_1_3_4_n45), .ZN(
        npu_inst_pe_1_3_4_n110) );
  AOI22_X1 npu_inst_pe_1_3_4_U103 ( .A1(npu_inst_int_data_y_4__4__0_), .A2(
        npu_inst_pe_1_3_4_n42), .B1(npu_inst_pe_1_3_4_n114), .B2(
        npu_inst_pe_1_3_4_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_3_4_n41) );
  INV_X1 npu_inst_pe_1_3_4_U102 ( .A(npu_inst_pe_1_3_4_n41), .ZN(
        npu_inst_pe_1_3_4_n111) );
  AOI22_X1 npu_inst_pe_1_3_4_U101 ( .A1(npu_inst_int_data_y_4__4__1_), .A2(
        npu_inst_pe_1_3_4_n58), .B1(npu_inst_pe_1_3_4_n118), .B2(
        npu_inst_pe_1_3_4_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_3_4_n59) );
  INV_X1 npu_inst_pe_1_3_4_U100 ( .A(npu_inst_pe_1_3_4_n59), .ZN(
        npu_inst_pe_1_3_4_n101) );
  AOI22_X1 npu_inst_pe_1_3_4_U99 ( .A1(npu_inst_int_data_y_4__4__1_), .A2(
        npu_inst_pe_1_3_4_n54), .B1(npu_inst_pe_1_3_4_n117), .B2(
        npu_inst_pe_1_3_4_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_3_4_n55) );
  INV_X1 npu_inst_pe_1_3_4_U98 ( .A(npu_inst_pe_1_3_4_n55), .ZN(
        npu_inst_pe_1_3_4_n102) );
  AOI22_X1 npu_inst_pe_1_3_4_U97 ( .A1(npu_inst_int_data_y_4__4__1_), .A2(
        npu_inst_pe_1_3_4_n50), .B1(npu_inst_pe_1_3_4_n116), .B2(
        npu_inst_pe_1_3_4_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_3_4_n51) );
  INV_X1 npu_inst_pe_1_3_4_U96 ( .A(npu_inst_pe_1_3_4_n51), .ZN(
        npu_inst_pe_1_3_4_n103) );
  AOI22_X1 npu_inst_pe_1_3_4_U95 ( .A1(npu_inst_int_data_y_4__4__1_), .A2(
        npu_inst_pe_1_3_4_n46), .B1(npu_inst_pe_1_3_4_n115), .B2(
        npu_inst_pe_1_3_4_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_3_4_n47) );
  INV_X1 npu_inst_pe_1_3_4_U94 ( .A(npu_inst_pe_1_3_4_n47), .ZN(
        npu_inst_pe_1_3_4_n104) );
  AOI22_X1 npu_inst_pe_1_3_4_U93 ( .A1(npu_inst_int_data_y_4__4__1_), .A2(
        npu_inst_pe_1_3_4_n42), .B1(npu_inst_pe_1_3_4_n114), .B2(
        npu_inst_pe_1_3_4_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_3_4_n43) );
  INV_X1 npu_inst_pe_1_3_4_U92 ( .A(npu_inst_pe_1_3_4_n43), .ZN(
        npu_inst_pe_1_3_4_n105) );
  AOI22_X1 npu_inst_pe_1_3_4_U91 ( .A1(npu_inst_pe_1_3_4_n38), .A2(
        npu_inst_int_data_y_4__4__1_), .B1(npu_inst_pe_1_3_4_n113), .B2(
        npu_inst_pe_1_3_4_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_3_4_n39) );
  INV_X1 npu_inst_pe_1_3_4_U90 ( .A(npu_inst_pe_1_3_4_n39), .ZN(
        npu_inst_pe_1_3_4_n106) );
  AOI22_X1 npu_inst_pe_1_3_4_U89 ( .A1(npu_inst_pe_1_3_4_n38), .A2(
        npu_inst_int_data_y_4__4__0_), .B1(npu_inst_pe_1_3_4_n113), .B2(
        npu_inst_pe_1_3_4_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_3_4_n37) );
  INV_X1 npu_inst_pe_1_3_4_U88 ( .A(npu_inst_pe_1_3_4_n37), .ZN(
        npu_inst_pe_1_3_4_n112) );
  NAND2_X1 npu_inst_pe_1_3_4_U87 ( .A1(npu_inst_pe_1_3_4_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_3_4_n60), .ZN(npu_inst_pe_1_3_4_n74) );
  OAI21_X1 npu_inst_pe_1_3_4_U86 ( .B1(npu_inst_pe_1_3_4_n63), .B2(
        npu_inst_pe_1_3_4_n60), .A(npu_inst_pe_1_3_4_n74), .ZN(
        npu_inst_pe_1_3_4_n97) );
  NAND2_X1 npu_inst_pe_1_3_4_U85 ( .A1(npu_inst_pe_1_3_4_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_3_4_n60), .ZN(npu_inst_pe_1_3_4_n73) );
  OAI21_X1 npu_inst_pe_1_3_4_U84 ( .B1(npu_inst_pe_1_3_4_n61), .B2(
        npu_inst_pe_1_3_4_n60), .A(npu_inst_pe_1_3_4_n73), .ZN(
        npu_inst_pe_1_3_4_n96) );
  NAND2_X1 npu_inst_pe_1_3_4_U83 ( .A1(npu_inst_pe_1_3_4_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_3_4_n56), .ZN(npu_inst_pe_1_3_4_n72) );
  OAI21_X1 npu_inst_pe_1_3_4_U82 ( .B1(npu_inst_pe_1_3_4_n63), .B2(
        npu_inst_pe_1_3_4_n56), .A(npu_inst_pe_1_3_4_n72), .ZN(
        npu_inst_pe_1_3_4_n95) );
  NAND2_X1 npu_inst_pe_1_3_4_U81 ( .A1(npu_inst_pe_1_3_4_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_3_4_n56), .ZN(npu_inst_pe_1_3_4_n71) );
  OAI21_X1 npu_inst_pe_1_3_4_U80 ( .B1(npu_inst_pe_1_3_4_n61), .B2(
        npu_inst_pe_1_3_4_n56), .A(npu_inst_pe_1_3_4_n71), .ZN(
        npu_inst_pe_1_3_4_n94) );
  NAND2_X1 npu_inst_pe_1_3_4_U79 ( .A1(npu_inst_pe_1_3_4_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_3_4_n52), .ZN(npu_inst_pe_1_3_4_n70) );
  OAI21_X1 npu_inst_pe_1_3_4_U78 ( .B1(npu_inst_pe_1_3_4_n63), .B2(
        npu_inst_pe_1_3_4_n52), .A(npu_inst_pe_1_3_4_n70), .ZN(
        npu_inst_pe_1_3_4_n93) );
  NAND2_X1 npu_inst_pe_1_3_4_U77 ( .A1(npu_inst_pe_1_3_4_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_3_4_n52), .ZN(npu_inst_pe_1_3_4_n69) );
  OAI21_X1 npu_inst_pe_1_3_4_U76 ( .B1(npu_inst_pe_1_3_4_n61), .B2(
        npu_inst_pe_1_3_4_n52), .A(npu_inst_pe_1_3_4_n69), .ZN(
        npu_inst_pe_1_3_4_n92) );
  NAND2_X1 npu_inst_pe_1_3_4_U75 ( .A1(npu_inst_pe_1_3_4_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_3_4_n48), .ZN(npu_inst_pe_1_3_4_n68) );
  OAI21_X1 npu_inst_pe_1_3_4_U74 ( .B1(npu_inst_pe_1_3_4_n63), .B2(
        npu_inst_pe_1_3_4_n48), .A(npu_inst_pe_1_3_4_n68), .ZN(
        npu_inst_pe_1_3_4_n91) );
  NAND2_X1 npu_inst_pe_1_3_4_U73 ( .A1(npu_inst_pe_1_3_4_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_3_4_n48), .ZN(npu_inst_pe_1_3_4_n67) );
  OAI21_X1 npu_inst_pe_1_3_4_U72 ( .B1(npu_inst_pe_1_3_4_n61), .B2(
        npu_inst_pe_1_3_4_n48), .A(npu_inst_pe_1_3_4_n67), .ZN(
        npu_inst_pe_1_3_4_n90) );
  NAND2_X1 npu_inst_pe_1_3_4_U71 ( .A1(npu_inst_pe_1_3_4_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_3_4_n44), .ZN(npu_inst_pe_1_3_4_n66) );
  OAI21_X1 npu_inst_pe_1_3_4_U70 ( .B1(npu_inst_pe_1_3_4_n63), .B2(
        npu_inst_pe_1_3_4_n44), .A(npu_inst_pe_1_3_4_n66), .ZN(
        npu_inst_pe_1_3_4_n89) );
  NAND2_X1 npu_inst_pe_1_3_4_U69 ( .A1(npu_inst_pe_1_3_4_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_3_4_n44), .ZN(npu_inst_pe_1_3_4_n65) );
  OAI21_X1 npu_inst_pe_1_3_4_U68 ( .B1(npu_inst_pe_1_3_4_n61), .B2(
        npu_inst_pe_1_3_4_n44), .A(npu_inst_pe_1_3_4_n65), .ZN(
        npu_inst_pe_1_3_4_n88) );
  NAND2_X1 npu_inst_pe_1_3_4_U67 ( .A1(npu_inst_pe_1_3_4_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_3_4_n40), .ZN(npu_inst_pe_1_3_4_n64) );
  OAI21_X1 npu_inst_pe_1_3_4_U66 ( .B1(npu_inst_pe_1_3_4_n63), .B2(
        npu_inst_pe_1_3_4_n40), .A(npu_inst_pe_1_3_4_n64), .ZN(
        npu_inst_pe_1_3_4_n87) );
  NAND2_X1 npu_inst_pe_1_3_4_U65 ( .A1(npu_inst_pe_1_3_4_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_3_4_n40), .ZN(npu_inst_pe_1_3_4_n62) );
  OAI21_X1 npu_inst_pe_1_3_4_U64 ( .B1(npu_inst_pe_1_3_4_n61), .B2(
        npu_inst_pe_1_3_4_n40), .A(npu_inst_pe_1_3_4_n62), .ZN(
        npu_inst_pe_1_3_4_n86) );
  AND2_X1 npu_inst_pe_1_3_4_U63 ( .A1(npu_inst_pe_1_3_4_N93), .A2(npu_inst_n57), .ZN(npu_inst_int_data_y_3__4__0_) );
  AND2_X1 npu_inst_pe_1_3_4_U62 ( .A1(npu_inst_n57), .A2(npu_inst_pe_1_3_4_N94), .ZN(npu_inst_int_data_y_3__4__1_) );
  NOR3_X1 npu_inst_pe_1_3_4_U61 ( .A1(npu_inst_pe_1_3_4_n26), .A2(npu_inst_n57), .A3(npu_inst_int_ckg[35]), .ZN(npu_inst_pe_1_3_4_n85) );
  OR2_X1 npu_inst_pe_1_3_4_U60 ( .A1(npu_inst_pe_1_3_4_n85), .A2(
        npu_inst_pe_1_3_4_n2), .ZN(npu_inst_pe_1_3_4_N84) );
  AND2_X1 npu_inst_pe_1_3_4_U59 ( .A1(npu_inst_pe_1_3_4_int_q_acc_0_), .A2(
        npu_inst_pe_1_3_4_n1), .ZN(npu_inst_int_data_res_3__4__0_) );
  AND2_X1 npu_inst_pe_1_3_4_U58 ( .A1(npu_inst_pe_1_3_4_n2), .A2(
        npu_inst_pe_1_3_4_int_q_acc_7_), .ZN(npu_inst_int_data_res_3__4__7_)
         );
  AND2_X1 npu_inst_pe_1_3_4_U57 ( .A1(npu_inst_pe_1_3_4_int_q_acc_1_), .A2(
        npu_inst_pe_1_3_4_n1), .ZN(npu_inst_int_data_res_3__4__1_) );
  AND2_X1 npu_inst_pe_1_3_4_U56 ( .A1(npu_inst_pe_1_3_4_int_q_acc_2_), .A2(
        npu_inst_pe_1_3_4_n1), .ZN(npu_inst_int_data_res_3__4__2_) );
  AND2_X1 npu_inst_pe_1_3_4_U55 ( .A1(npu_inst_pe_1_3_4_int_q_acc_3_), .A2(
        npu_inst_pe_1_3_4_n2), .ZN(npu_inst_int_data_res_3__4__3_) );
  AND2_X1 npu_inst_pe_1_3_4_U54 ( .A1(npu_inst_pe_1_3_4_int_q_acc_4_), .A2(
        npu_inst_pe_1_3_4_n2), .ZN(npu_inst_int_data_res_3__4__4_) );
  AND2_X1 npu_inst_pe_1_3_4_U53 ( .A1(npu_inst_pe_1_3_4_int_q_acc_5_), .A2(
        npu_inst_pe_1_3_4_n2), .ZN(npu_inst_int_data_res_3__4__5_) );
  AND2_X1 npu_inst_pe_1_3_4_U52 ( .A1(npu_inst_pe_1_3_4_int_q_acc_6_), .A2(
        npu_inst_pe_1_3_4_n2), .ZN(npu_inst_int_data_res_3__4__6_) );
  AOI222_X1 npu_inst_pe_1_3_4_U51 ( .A1(npu_inst_int_data_res_4__4__0_), .A2(
        npu_inst_pe_1_3_4_n1), .B1(npu_inst_pe_1_3_4_N73), .B2(
        npu_inst_pe_1_3_4_n76), .C1(npu_inst_pe_1_3_4_N65), .C2(
        npu_inst_pe_1_3_4_n77), .ZN(npu_inst_pe_1_3_4_n84) );
  INV_X1 npu_inst_pe_1_3_4_U50 ( .A(npu_inst_pe_1_3_4_n84), .ZN(
        npu_inst_pe_1_3_4_n100) );
  AOI222_X1 npu_inst_pe_1_3_4_U49 ( .A1(npu_inst_int_data_res_4__4__7_), .A2(
        npu_inst_pe_1_3_4_n1), .B1(npu_inst_pe_1_3_4_N80), .B2(
        npu_inst_pe_1_3_4_n76), .C1(npu_inst_pe_1_3_4_N72), .C2(
        npu_inst_pe_1_3_4_n77), .ZN(npu_inst_pe_1_3_4_n75) );
  INV_X1 npu_inst_pe_1_3_4_U48 ( .A(npu_inst_pe_1_3_4_n75), .ZN(
        npu_inst_pe_1_3_4_n32) );
  AOI222_X1 npu_inst_pe_1_3_4_U47 ( .A1(npu_inst_int_data_res_4__4__1_), .A2(
        npu_inst_pe_1_3_4_n1), .B1(npu_inst_pe_1_3_4_N74), .B2(
        npu_inst_pe_1_3_4_n76), .C1(npu_inst_pe_1_3_4_N66), .C2(
        npu_inst_pe_1_3_4_n77), .ZN(npu_inst_pe_1_3_4_n83) );
  INV_X1 npu_inst_pe_1_3_4_U46 ( .A(npu_inst_pe_1_3_4_n83), .ZN(
        npu_inst_pe_1_3_4_n99) );
  AOI222_X1 npu_inst_pe_1_3_4_U45 ( .A1(npu_inst_int_data_res_4__4__2_), .A2(
        npu_inst_pe_1_3_4_n1), .B1(npu_inst_pe_1_3_4_N75), .B2(
        npu_inst_pe_1_3_4_n76), .C1(npu_inst_pe_1_3_4_N67), .C2(
        npu_inst_pe_1_3_4_n77), .ZN(npu_inst_pe_1_3_4_n82) );
  INV_X1 npu_inst_pe_1_3_4_U44 ( .A(npu_inst_pe_1_3_4_n82), .ZN(
        npu_inst_pe_1_3_4_n98) );
  AOI222_X1 npu_inst_pe_1_3_4_U43 ( .A1(npu_inst_int_data_res_4__4__3_), .A2(
        npu_inst_pe_1_3_4_n1), .B1(npu_inst_pe_1_3_4_N76), .B2(
        npu_inst_pe_1_3_4_n76), .C1(npu_inst_pe_1_3_4_N68), .C2(
        npu_inst_pe_1_3_4_n77), .ZN(npu_inst_pe_1_3_4_n81) );
  INV_X1 npu_inst_pe_1_3_4_U42 ( .A(npu_inst_pe_1_3_4_n81), .ZN(
        npu_inst_pe_1_3_4_n36) );
  AOI222_X1 npu_inst_pe_1_3_4_U41 ( .A1(npu_inst_int_data_res_4__4__4_), .A2(
        npu_inst_pe_1_3_4_n1), .B1(npu_inst_pe_1_3_4_N77), .B2(
        npu_inst_pe_1_3_4_n76), .C1(npu_inst_pe_1_3_4_N69), .C2(
        npu_inst_pe_1_3_4_n77), .ZN(npu_inst_pe_1_3_4_n80) );
  INV_X1 npu_inst_pe_1_3_4_U40 ( .A(npu_inst_pe_1_3_4_n80), .ZN(
        npu_inst_pe_1_3_4_n35) );
  AOI222_X1 npu_inst_pe_1_3_4_U39 ( .A1(npu_inst_int_data_res_4__4__5_), .A2(
        npu_inst_pe_1_3_4_n1), .B1(npu_inst_pe_1_3_4_N78), .B2(
        npu_inst_pe_1_3_4_n76), .C1(npu_inst_pe_1_3_4_N70), .C2(
        npu_inst_pe_1_3_4_n77), .ZN(npu_inst_pe_1_3_4_n79) );
  INV_X1 npu_inst_pe_1_3_4_U38 ( .A(npu_inst_pe_1_3_4_n79), .ZN(
        npu_inst_pe_1_3_4_n34) );
  AOI222_X1 npu_inst_pe_1_3_4_U37 ( .A1(npu_inst_int_data_res_4__4__6_), .A2(
        npu_inst_pe_1_3_4_n1), .B1(npu_inst_pe_1_3_4_N79), .B2(
        npu_inst_pe_1_3_4_n76), .C1(npu_inst_pe_1_3_4_N71), .C2(
        npu_inst_pe_1_3_4_n77), .ZN(npu_inst_pe_1_3_4_n78) );
  INV_X1 npu_inst_pe_1_3_4_U36 ( .A(npu_inst_pe_1_3_4_n78), .ZN(
        npu_inst_pe_1_3_4_n33) );
  INV_X1 npu_inst_pe_1_3_4_U35 ( .A(npu_inst_pe_1_3_4_int_data_1_), .ZN(
        npu_inst_pe_1_3_4_n13) );
  AND2_X1 npu_inst_pe_1_3_4_U34 ( .A1(npu_inst_int_data_x_3__4__1_), .A2(
        npu_inst_pe_1_3_4_int_q_weight_1_), .ZN(npu_inst_pe_1_3_4_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_3_4_U33 ( .A1(npu_inst_int_data_x_3__4__0_), .A2(
        npu_inst_pe_1_3_4_int_q_weight_1_), .ZN(npu_inst_pe_1_3_4_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_3_4_U32 ( .A1(npu_inst_n57), .A2(
        npu_inst_int_data_y_4__4__1_), .B1(npu_inst_pe_1_3_4_n3), .B2(
        npu_inst_int_data_x_3__5__1_), .ZN(npu_inst_pe_1_3_4_n63) );
  AOI22_X1 npu_inst_pe_1_3_4_U31 ( .A1(npu_inst_n57), .A2(
        npu_inst_int_data_y_4__4__0_), .B1(npu_inst_pe_1_3_4_n3), .B2(
        npu_inst_int_data_x_3__5__0_), .ZN(npu_inst_pe_1_3_4_n61) );
  INV_X1 npu_inst_pe_1_3_4_U30 ( .A(npu_inst_pe_1_3_4_int_data_0_), .ZN(
        npu_inst_pe_1_3_4_n12) );
  INV_X1 npu_inst_pe_1_3_4_U29 ( .A(npu_inst_n69), .ZN(npu_inst_pe_1_3_4_n5)
         );
  OR3_X1 npu_inst_pe_1_3_4_U28 ( .A1(npu_inst_n77), .A2(npu_inst_pe_1_3_4_n7), 
        .A3(npu_inst_pe_1_3_4_n5), .ZN(npu_inst_pe_1_3_4_n56) );
  OR3_X1 npu_inst_pe_1_3_4_U27 ( .A1(npu_inst_pe_1_3_4_n5), .A2(
        npu_inst_pe_1_3_4_n7), .A3(npu_inst_pe_1_3_4_n6), .ZN(
        npu_inst_pe_1_3_4_n48) );
  INV_X1 npu_inst_pe_1_3_4_U26 ( .A(npu_inst_pe_1_3_4_n5), .ZN(
        npu_inst_pe_1_3_4_n4) );
  OR3_X1 npu_inst_pe_1_3_4_U25 ( .A1(npu_inst_pe_1_3_4_n4), .A2(
        npu_inst_pe_1_3_4_n7), .A3(npu_inst_pe_1_3_4_n6), .ZN(
        npu_inst_pe_1_3_4_n52) );
  OR3_X1 npu_inst_pe_1_3_4_U24 ( .A1(npu_inst_n77), .A2(npu_inst_pe_1_3_4_n7), 
        .A3(npu_inst_pe_1_3_4_n4), .ZN(npu_inst_pe_1_3_4_n60) );
  NOR2_X1 npu_inst_pe_1_3_4_U23 ( .A1(npu_inst_pe_1_3_4_n60), .A2(
        npu_inst_pe_1_3_4_n3), .ZN(npu_inst_pe_1_3_4_n58) );
  NOR2_X1 npu_inst_pe_1_3_4_U22 ( .A1(npu_inst_pe_1_3_4_n56), .A2(
        npu_inst_pe_1_3_4_n3), .ZN(npu_inst_pe_1_3_4_n54) );
  NOR2_X1 npu_inst_pe_1_3_4_U21 ( .A1(npu_inst_pe_1_3_4_n52), .A2(
        npu_inst_pe_1_3_4_n3), .ZN(npu_inst_pe_1_3_4_n50) );
  NOR2_X1 npu_inst_pe_1_3_4_U20 ( .A1(npu_inst_pe_1_3_4_n48), .A2(
        npu_inst_pe_1_3_4_n3), .ZN(npu_inst_pe_1_3_4_n46) );
  NOR2_X1 npu_inst_pe_1_3_4_U19 ( .A1(npu_inst_pe_1_3_4_n40), .A2(
        npu_inst_pe_1_3_4_n3), .ZN(npu_inst_pe_1_3_4_n38) );
  NOR2_X1 npu_inst_pe_1_3_4_U18 ( .A1(npu_inst_pe_1_3_4_n44), .A2(
        npu_inst_pe_1_3_4_n3), .ZN(npu_inst_pe_1_3_4_n42) );
  BUF_X1 npu_inst_pe_1_3_4_U17 ( .A(npu_inst_n100), .Z(npu_inst_pe_1_3_4_n7)
         );
  INV_X1 npu_inst_pe_1_3_4_U16 ( .A(npu_inst_n124), .ZN(npu_inst_pe_1_3_4_n11)
         );
  INV_X1 npu_inst_pe_1_3_4_U15 ( .A(npu_inst_pe_1_3_4_n38), .ZN(
        npu_inst_pe_1_3_4_n113) );
  INV_X1 npu_inst_pe_1_3_4_U14 ( .A(npu_inst_pe_1_3_4_n58), .ZN(
        npu_inst_pe_1_3_4_n118) );
  INV_X1 npu_inst_pe_1_3_4_U13 ( .A(npu_inst_pe_1_3_4_n54), .ZN(
        npu_inst_pe_1_3_4_n117) );
  INV_X1 npu_inst_pe_1_3_4_U12 ( .A(npu_inst_pe_1_3_4_n50), .ZN(
        npu_inst_pe_1_3_4_n116) );
  INV_X1 npu_inst_pe_1_3_4_U11 ( .A(npu_inst_pe_1_3_4_n46), .ZN(
        npu_inst_pe_1_3_4_n115) );
  INV_X1 npu_inst_pe_1_3_4_U10 ( .A(npu_inst_pe_1_3_4_n42), .ZN(
        npu_inst_pe_1_3_4_n114) );
  BUF_X1 npu_inst_pe_1_3_4_U9 ( .A(npu_inst_n24), .Z(npu_inst_pe_1_3_4_n2) );
  BUF_X1 npu_inst_pe_1_3_4_U8 ( .A(npu_inst_n24), .Z(npu_inst_pe_1_3_4_n1) );
  BUF_X1 npu_inst_pe_1_3_4_U7 ( .A(npu_inst_pe_1_3_4_n11), .Z(
        npu_inst_pe_1_3_4_n10) );
  BUF_X1 npu_inst_pe_1_3_4_U6 ( .A(npu_inst_pe_1_3_4_n11), .Z(
        npu_inst_pe_1_3_4_n9) );
  BUF_X1 npu_inst_pe_1_3_4_U5 ( .A(npu_inst_pe_1_3_4_n11), .Z(
        npu_inst_pe_1_3_4_n8) );
  NOR2_X1 npu_inst_pe_1_3_4_U4 ( .A1(npu_inst_pe_1_3_4_int_q_weight_0_), .A2(
        npu_inst_pe_1_3_4_n1), .ZN(npu_inst_pe_1_3_4_n76) );
  NOR2_X1 npu_inst_pe_1_3_4_U3 ( .A1(npu_inst_pe_1_3_4_n27), .A2(
        npu_inst_pe_1_3_4_n1), .ZN(npu_inst_pe_1_3_4_n77) );
  FA_X1 npu_inst_pe_1_3_4_sub_67_U2_1 ( .A(npu_inst_pe_1_3_4_int_q_acc_1_), 
        .B(npu_inst_pe_1_3_4_n13), .CI(npu_inst_pe_1_3_4_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_3_4_sub_67_carry_2_), .S(npu_inst_pe_1_3_4_N66) );
  FA_X1 npu_inst_pe_1_3_4_add_69_U1_1 ( .A(npu_inst_pe_1_3_4_int_q_acc_1_), 
        .B(npu_inst_pe_1_3_4_int_data_1_), .CI(
        npu_inst_pe_1_3_4_add_69_carry_1_), .CO(
        npu_inst_pe_1_3_4_add_69_carry_2_), .S(npu_inst_pe_1_3_4_N74) );
  NAND3_X1 npu_inst_pe_1_3_4_U109 ( .A1(npu_inst_pe_1_3_4_n5), .A2(
        npu_inst_pe_1_3_4_n6), .A3(npu_inst_pe_1_3_4_n7), .ZN(
        npu_inst_pe_1_3_4_n44) );
  NAND3_X1 npu_inst_pe_1_3_4_U108 ( .A1(npu_inst_pe_1_3_4_n4), .A2(
        npu_inst_pe_1_3_4_n6), .A3(npu_inst_pe_1_3_4_n7), .ZN(
        npu_inst_pe_1_3_4_n40) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_3_4_n33), .CK(
        npu_inst_pe_1_3_4_net3918), .RN(npu_inst_pe_1_3_4_n8), .Q(
        npu_inst_pe_1_3_4_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_3_4_n34), .CK(
        npu_inst_pe_1_3_4_net3918), .RN(npu_inst_pe_1_3_4_n8), .Q(
        npu_inst_pe_1_3_4_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_3_4_n35), .CK(
        npu_inst_pe_1_3_4_net3918), .RN(npu_inst_pe_1_3_4_n8), .Q(
        npu_inst_pe_1_3_4_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_3_4_n36), .CK(
        npu_inst_pe_1_3_4_net3918), .RN(npu_inst_pe_1_3_4_n8), .Q(
        npu_inst_pe_1_3_4_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_3_4_n98), .CK(
        npu_inst_pe_1_3_4_net3918), .RN(npu_inst_pe_1_3_4_n8), .Q(
        npu_inst_pe_1_3_4_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_3_4_n99), .CK(
        npu_inst_pe_1_3_4_net3918), .RN(npu_inst_pe_1_3_4_n8), .Q(
        npu_inst_pe_1_3_4_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_3_4_n32), .CK(
        npu_inst_pe_1_3_4_net3918), .RN(npu_inst_pe_1_3_4_n8), .Q(
        npu_inst_pe_1_3_4_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_3_4_n100), 
        .CK(npu_inst_pe_1_3_4_net3918), .RN(npu_inst_pe_1_3_4_n8), .Q(
        npu_inst_pe_1_3_4_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_weight_reg_0_ ( .D(npu_inst_n110), .CK(
        npu_inst_pe_1_3_4_net3924), .RN(npu_inst_pe_1_3_4_n8), .Q(
        npu_inst_pe_1_3_4_int_q_weight_0_), .QN(npu_inst_pe_1_3_4_n27) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_weight_reg_1_ ( .D(npu_inst_n116), .CK(
        npu_inst_pe_1_3_4_net3924), .RN(npu_inst_pe_1_3_4_n8), .Q(
        npu_inst_pe_1_3_4_int_q_weight_1_), .QN(npu_inst_pe_1_3_4_n26) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_3_4_n112), 
        .CK(npu_inst_pe_1_3_4_net3924), .RN(npu_inst_pe_1_3_4_n8), .Q(
        npu_inst_pe_1_3_4_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_3_4_n106), 
        .CK(npu_inst_pe_1_3_4_net3924), .RN(npu_inst_pe_1_3_4_n8), .Q(
        npu_inst_pe_1_3_4_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_3_4_n111), 
        .CK(npu_inst_pe_1_3_4_net3924), .RN(npu_inst_pe_1_3_4_n9), .Q(
        npu_inst_pe_1_3_4_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_3_4_n105), 
        .CK(npu_inst_pe_1_3_4_net3924), .RN(npu_inst_pe_1_3_4_n9), .Q(
        npu_inst_pe_1_3_4_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_3_4_n110), 
        .CK(npu_inst_pe_1_3_4_net3924), .RN(npu_inst_pe_1_3_4_n9), .Q(
        npu_inst_pe_1_3_4_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_3_4_n104), 
        .CK(npu_inst_pe_1_3_4_net3924), .RN(npu_inst_pe_1_3_4_n9), .Q(
        npu_inst_pe_1_3_4_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_3_4_n109), 
        .CK(npu_inst_pe_1_3_4_net3924), .RN(npu_inst_pe_1_3_4_n9), .Q(
        npu_inst_pe_1_3_4_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_3_4_n103), 
        .CK(npu_inst_pe_1_3_4_net3924), .RN(npu_inst_pe_1_3_4_n9), .Q(
        npu_inst_pe_1_3_4_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_3_4_n108), 
        .CK(npu_inst_pe_1_3_4_net3924), .RN(npu_inst_pe_1_3_4_n9), .Q(
        npu_inst_pe_1_3_4_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_3_4_n102), 
        .CK(npu_inst_pe_1_3_4_net3924), .RN(npu_inst_pe_1_3_4_n9), .Q(
        npu_inst_pe_1_3_4_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_3_4_n107), 
        .CK(npu_inst_pe_1_3_4_net3924), .RN(npu_inst_pe_1_3_4_n9), .Q(
        npu_inst_pe_1_3_4_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_3_4_n101), 
        .CK(npu_inst_pe_1_3_4_net3924), .RN(npu_inst_pe_1_3_4_n9), .Q(
        npu_inst_pe_1_3_4_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_3_4_n86), 
        .CK(npu_inst_pe_1_3_4_net3924), .RN(npu_inst_pe_1_3_4_n9), .Q(
        npu_inst_pe_1_3_4_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_3_4_n87), 
        .CK(npu_inst_pe_1_3_4_net3924), .RN(npu_inst_pe_1_3_4_n9), .Q(
        npu_inst_pe_1_3_4_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_3_4_n88), 
        .CK(npu_inst_pe_1_3_4_net3924), .RN(npu_inst_pe_1_3_4_n10), .Q(
        npu_inst_pe_1_3_4_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_3_4_n89), 
        .CK(npu_inst_pe_1_3_4_net3924), .RN(npu_inst_pe_1_3_4_n10), .Q(
        npu_inst_pe_1_3_4_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_3_4_n90), 
        .CK(npu_inst_pe_1_3_4_net3924), .RN(npu_inst_pe_1_3_4_n10), .Q(
        npu_inst_pe_1_3_4_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_3_4_n91), 
        .CK(npu_inst_pe_1_3_4_net3924), .RN(npu_inst_pe_1_3_4_n10), .Q(
        npu_inst_pe_1_3_4_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_3_4_n92), 
        .CK(npu_inst_pe_1_3_4_net3924), .RN(npu_inst_pe_1_3_4_n10), .Q(
        npu_inst_pe_1_3_4_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_3_4_n93), 
        .CK(npu_inst_pe_1_3_4_net3924), .RN(npu_inst_pe_1_3_4_n10), .Q(
        npu_inst_pe_1_3_4_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_3_4_n94), 
        .CK(npu_inst_pe_1_3_4_net3924), .RN(npu_inst_pe_1_3_4_n10), .Q(
        npu_inst_pe_1_3_4_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_3_4_n95), 
        .CK(npu_inst_pe_1_3_4_net3924), .RN(npu_inst_pe_1_3_4_n10), .Q(
        npu_inst_pe_1_3_4_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_3_4_n96), 
        .CK(npu_inst_pe_1_3_4_net3924), .RN(npu_inst_pe_1_3_4_n10), .Q(
        npu_inst_pe_1_3_4_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_3_4_n97), 
        .CK(npu_inst_pe_1_3_4_net3924), .RN(npu_inst_pe_1_3_4_n10), .Q(
        npu_inst_pe_1_3_4_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_3_4_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_3_4_N84), .SE(1'b0), .GCK(npu_inst_pe_1_3_4_net3918) );
  CLKGATETST_X1 npu_inst_pe_1_3_4_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n64), .SE(1'b0), .GCK(npu_inst_pe_1_3_4_net3924) );
  MUX2_X1 npu_inst_pe_1_3_5_U162 ( .A(npu_inst_pe_1_3_5_n32), .B(
        npu_inst_pe_1_3_5_n29), .S(npu_inst_pe_1_3_5_n8), .Z(
        npu_inst_pe_1_3_5_N93) );
  MUX2_X1 npu_inst_pe_1_3_5_U161 ( .A(npu_inst_pe_1_3_5_n31), .B(
        npu_inst_pe_1_3_5_n30), .S(npu_inst_pe_1_3_5_n6), .Z(
        npu_inst_pe_1_3_5_n32) );
  MUX2_X1 npu_inst_pe_1_3_5_U160 ( .A(npu_inst_pe_1_3_5_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_3_5_int_q_reg_v_1__0_), .S(npu_inst_pe_1_3_5_n4), .Z(
        npu_inst_pe_1_3_5_n31) );
  MUX2_X1 npu_inst_pe_1_3_5_U159 ( .A(npu_inst_pe_1_3_5_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_3_5_int_q_reg_v_3__0_), .S(npu_inst_pe_1_3_5_n4), .Z(
        npu_inst_pe_1_3_5_n30) );
  MUX2_X1 npu_inst_pe_1_3_5_U158 ( .A(npu_inst_pe_1_3_5_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_3_5_int_q_reg_v_5__0_), .S(npu_inst_pe_1_3_5_n4), .Z(
        npu_inst_pe_1_3_5_n29) );
  MUX2_X1 npu_inst_pe_1_3_5_U157 ( .A(npu_inst_pe_1_3_5_n28), .B(
        npu_inst_pe_1_3_5_n23), .S(npu_inst_pe_1_3_5_n8), .Z(
        npu_inst_pe_1_3_5_N94) );
  MUX2_X1 npu_inst_pe_1_3_5_U156 ( .A(npu_inst_pe_1_3_5_n25), .B(
        npu_inst_pe_1_3_5_n24), .S(npu_inst_pe_1_3_5_n6), .Z(
        npu_inst_pe_1_3_5_n28) );
  MUX2_X1 npu_inst_pe_1_3_5_U155 ( .A(npu_inst_pe_1_3_5_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_3_5_int_q_reg_v_1__1_), .S(npu_inst_pe_1_3_5_n4), .Z(
        npu_inst_pe_1_3_5_n25) );
  MUX2_X1 npu_inst_pe_1_3_5_U154 ( .A(npu_inst_pe_1_3_5_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_3_5_int_q_reg_v_3__1_), .S(npu_inst_pe_1_3_5_n4), .Z(
        npu_inst_pe_1_3_5_n24) );
  MUX2_X1 npu_inst_pe_1_3_5_U153 ( .A(npu_inst_pe_1_3_5_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_3_5_int_q_reg_v_5__1_), .S(npu_inst_pe_1_3_5_n4), .Z(
        npu_inst_pe_1_3_5_n23) );
  MUX2_X1 npu_inst_pe_1_3_5_U152 ( .A(npu_inst_pe_1_3_5_n22), .B(
        npu_inst_pe_1_3_5_n19), .S(npu_inst_pe_1_3_5_n8), .Z(
        npu_inst_int_data_x_3__5__1_) );
  MUX2_X1 npu_inst_pe_1_3_5_U151 ( .A(npu_inst_pe_1_3_5_n21), .B(
        npu_inst_pe_1_3_5_n20), .S(npu_inst_pe_1_3_5_n6), .Z(
        npu_inst_pe_1_3_5_n22) );
  MUX2_X1 npu_inst_pe_1_3_5_U150 ( .A(npu_inst_pe_1_3_5_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_3_5_int_q_reg_h_1__1_), .S(npu_inst_pe_1_3_5_n4), .Z(
        npu_inst_pe_1_3_5_n21) );
  MUX2_X1 npu_inst_pe_1_3_5_U149 ( .A(npu_inst_pe_1_3_5_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_3_5_int_q_reg_h_3__1_), .S(npu_inst_pe_1_3_5_n4), .Z(
        npu_inst_pe_1_3_5_n20) );
  MUX2_X1 npu_inst_pe_1_3_5_U148 ( .A(npu_inst_pe_1_3_5_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_3_5_int_q_reg_h_5__1_), .S(npu_inst_pe_1_3_5_n4), .Z(
        npu_inst_pe_1_3_5_n19) );
  MUX2_X1 npu_inst_pe_1_3_5_U147 ( .A(npu_inst_pe_1_3_5_n18), .B(
        npu_inst_pe_1_3_5_n15), .S(npu_inst_pe_1_3_5_n8), .Z(
        npu_inst_int_data_x_3__5__0_) );
  MUX2_X1 npu_inst_pe_1_3_5_U146 ( .A(npu_inst_pe_1_3_5_n17), .B(
        npu_inst_pe_1_3_5_n16), .S(npu_inst_pe_1_3_5_n6), .Z(
        npu_inst_pe_1_3_5_n18) );
  MUX2_X1 npu_inst_pe_1_3_5_U145 ( .A(npu_inst_pe_1_3_5_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_3_5_int_q_reg_h_1__0_), .S(npu_inst_pe_1_3_5_n4), .Z(
        npu_inst_pe_1_3_5_n17) );
  MUX2_X1 npu_inst_pe_1_3_5_U144 ( .A(npu_inst_pe_1_3_5_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_3_5_int_q_reg_h_3__0_), .S(npu_inst_pe_1_3_5_n4), .Z(
        npu_inst_pe_1_3_5_n16) );
  MUX2_X1 npu_inst_pe_1_3_5_U143 ( .A(npu_inst_pe_1_3_5_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_3_5_int_q_reg_h_5__0_), .S(npu_inst_pe_1_3_5_n4), .Z(
        npu_inst_pe_1_3_5_n15) );
  XOR2_X1 npu_inst_pe_1_3_5_U142 ( .A(npu_inst_pe_1_3_5_int_data_0_), .B(
        npu_inst_pe_1_3_5_int_q_acc_0_), .Z(npu_inst_pe_1_3_5_N73) );
  AND2_X1 npu_inst_pe_1_3_5_U141 ( .A1(npu_inst_pe_1_3_5_int_q_acc_0_), .A2(
        npu_inst_pe_1_3_5_int_data_0_), .ZN(npu_inst_pe_1_3_5_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_3_5_U140 ( .A(npu_inst_pe_1_3_5_int_q_acc_0_), .B(
        npu_inst_pe_1_3_5_n13), .ZN(npu_inst_pe_1_3_5_N65) );
  OR2_X1 npu_inst_pe_1_3_5_U139 ( .A1(npu_inst_pe_1_3_5_n13), .A2(
        npu_inst_pe_1_3_5_int_q_acc_0_), .ZN(npu_inst_pe_1_3_5_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_3_5_U138 ( .A(npu_inst_pe_1_3_5_int_q_acc_2_), .B(
        npu_inst_pe_1_3_5_add_69_carry_2_), .Z(npu_inst_pe_1_3_5_N75) );
  AND2_X1 npu_inst_pe_1_3_5_U137 ( .A1(npu_inst_pe_1_3_5_add_69_carry_2_), 
        .A2(npu_inst_pe_1_3_5_int_q_acc_2_), .ZN(
        npu_inst_pe_1_3_5_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_3_5_U136 ( .A(npu_inst_pe_1_3_5_int_q_acc_3_), .B(
        npu_inst_pe_1_3_5_add_69_carry_3_), .Z(npu_inst_pe_1_3_5_N76) );
  AND2_X1 npu_inst_pe_1_3_5_U135 ( .A1(npu_inst_pe_1_3_5_add_69_carry_3_), 
        .A2(npu_inst_pe_1_3_5_int_q_acc_3_), .ZN(
        npu_inst_pe_1_3_5_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_3_5_U134 ( .A(npu_inst_pe_1_3_5_int_q_acc_4_), .B(
        npu_inst_pe_1_3_5_add_69_carry_4_), .Z(npu_inst_pe_1_3_5_N77) );
  AND2_X1 npu_inst_pe_1_3_5_U133 ( .A1(npu_inst_pe_1_3_5_add_69_carry_4_), 
        .A2(npu_inst_pe_1_3_5_int_q_acc_4_), .ZN(
        npu_inst_pe_1_3_5_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_3_5_U132 ( .A(npu_inst_pe_1_3_5_int_q_acc_5_), .B(
        npu_inst_pe_1_3_5_add_69_carry_5_), .Z(npu_inst_pe_1_3_5_N78) );
  AND2_X1 npu_inst_pe_1_3_5_U131 ( .A1(npu_inst_pe_1_3_5_add_69_carry_5_), 
        .A2(npu_inst_pe_1_3_5_int_q_acc_5_), .ZN(
        npu_inst_pe_1_3_5_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_3_5_U130 ( .A(npu_inst_pe_1_3_5_int_q_acc_6_), .B(
        npu_inst_pe_1_3_5_add_69_carry_6_), .Z(npu_inst_pe_1_3_5_N79) );
  AND2_X1 npu_inst_pe_1_3_5_U129 ( .A1(npu_inst_pe_1_3_5_add_69_carry_6_), 
        .A2(npu_inst_pe_1_3_5_int_q_acc_6_), .ZN(
        npu_inst_pe_1_3_5_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_3_5_U128 ( .A(npu_inst_pe_1_3_5_int_q_acc_7_), .B(
        npu_inst_pe_1_3_5_add_69_carry_7_), .Z(npu_inst_pe_1_3_5_N80) );
  XNOR2_X1 npu_inst_pe_1_3_5_U127 ( .A(npu_inst_pe_1_3_5_sub_67_carry_2_), .B(
        npu_inst_pe_1_3_5_int_q_acc_2_), .ZN(npu_inst_pe_1_3_5_N67) );
  OR2_X1 npu_inst_pe_1_3_5_U126 ( .A1(npu_inst_pe_1_3_5_int_q_acc_2_), .A2(
        npu_inst_pe_1_3_5_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_3_5_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_3_5_U125 ( .A(npu_inst_pe_1_3_5_sub_67_carry_3_), .B(
        npu_inst_pe_1_3_5_int_q_acc_3_), .ZN(npu_inst_pe_1_3_5_N68) );
  OR2_X1 npu_inst_pe_1_3_5_U124 ( .A1(npu_inst_pe_1_3_5_int_q_acc_3_), .A2(
        npu_inst_pe_1_3_5_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_3_5_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_3_5_U123 ( .A(npu_inst_pe_1_3_5_sub_67_carry_4_), .B(
        npu_inst_pe_1_3_5_int_q_acc_4_), .ZN(npu_inst_pe_1_3_5_N69) );
  OR2_X1 npu_inst_pe_1_3_5_U122 ( .A1(npu_inst_pe_1_3_5_int_q_acc_4_), .A2(
        npu_inst_pe_1_3_5_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_3_5_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_3_5_U121 ( .A(npu_inst_pe_1_3_5_sub_67_carry_5_), .B(
        npu_inst_pe_1_3_5_int_q_acc_5_), .ZN(npu_inst_pe_1_3_5_N70) );
  OR2_X1 npu_inst_pe_1_3_5_U120 ( .A1(npu_inst_pe_1_3_5_int_q_acc_5_), .A2(
        npu_inst_pe_1_3_5_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_3_5_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_3_5_U119 ( .A(npu_inst_pe_1_3_5_sub_67_carry_6_), .B(
        npu_inst_pe_1_3_5_int_q_acc_6_), .ZN(npu_inst_pe_1_3_5_N71) );
  OR2_X1 npu_inst_pe_1_3_5_U118 ( .A1(npu_inst_pe_1_3_5_int_q_acc_6_), .A2(
        npu_inst_pe_1_3_5_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_3_5_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_3_5_U117 ( .A(npu_inst_pe_1_3_5_int_q_acc_7_), .B(
        npu_inst_pe_1_3_5_sub_67_carry_7_), .ZN(npu_inst_pe_1_3_5_N72) );
  INV_X1 npu_inst_pe_1_3_5_U116 ( .A(npu_inst_n77), .ZN(npu_inst_pe_1_3_5_n7)
         );
  INV_X1 npu_inst_pe_1_3_5_U115 ( .A(npu_inst_pe_1_3_5_n7), .ZN(
        npu_inst_pe_1_3_5_n6) );
  INV_X1 npu_inst_pe_1_3_5_U114 ( .A(npu_inst_n56), .ZN(npu_inst_pe_1_3_5_n3)
         );
  AOI22_X1 npu_inst_pe_1_3_5_U113 ( .A1(npu_inst_int_data_y_4__5__0_), .A2(
        npu_inst_pe_1_3_5_n58), .B1(npu_inst_pe_1_3_5_n119), .B2(
        npu_inst_pe_1_3_5_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_3_5_n57) );
  INV_X1 npu_inst_pe_1_3_5_U112 ( .A(npu_inst_pe_1_3_5_n57), .ZN(
        npu_inst_pe_1_3_5_n108) );
  AOI22_X1 npu_inst_pe_1_3_5_U111 ( .A1(npu_inst_int_data_y_4__5__0_), .A2(
        npu_inst_pe_1_3_5_n54), .B1(npu_inst_pe_1_3_5_n118), .B2(
        npu_inst_pe_1_3_5_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_3_5_n53) );
  INV_X1 npu_inst_pe_1_3_5_U110 ( .A(npu_inst_pe_1_3_5_n53), .ZN(
        npu_inst_pe_1_3_5_n109) );
  AOI22_X1 npu_inst_pe_1_3_5_U107 ( .A1(npu_inst_int_data_y_4__5__0_), .A2(
        npu_inst_pe_1_3_5_n50), .B1(npu_inst_pe_1_3_5_n117), .B2(
        npu_inst_pe_1_3_5_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_3_5_n49) );
  INV_X1 npu_inst_pe_1_3_5_U106 ( .A(npu_inst_pe_1_3_5_n49), .ZN(
        npu_inst_pe_1_3_5_n110) );
  AOI22_X1 npu_inst_pe_1_3_5_U105 ( .A1(npu_inst_int_data_y_4__5__0_), .A2(
        npu_inst_pe_1_3_5_n46), .B1(npu_inst_pe_1_3_5_n116), .B2(
        npu_inst_pe_1_3_5_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_3_5_n45) );
  INV_X1 npu_inst_pe_1_3_5_U104 ( .A(npu_inst_pe_1_3_5_n45), .ZN(
        npu_inst_pe_1_3_5_n111) );
  AOI22_X1 npu_inst_pe_1_3_5_U103 ( .A1(npu_inst_int_data_y_4__5__0_), .A2(
        npu_inst_pe_1_3_5_n42), .B1(npu_inst_pe_1_3_5_n115), .B2(
        npu_inst_pe_1_3_5_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_3_5_n41) );
  INV_X1 npu_inst_pe_1_3_5_U102 ( .A(npu_inst_pe_1_3_5_n41), .ZN(
        npu_inst_pe_1_3_5_n112) );
  AOI22_X1 npu_inst_pe_1_3_5_U101 ( .A1(npu_inst_int_data_y_4__5__1_), .A2(
        npu_inst_pe_1_3_5_n58), .B1(npu_inst_pe_1_3_5_n119), .B2(
        npu_inst_pe_1_3_5_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_3_5_n59) );
  INV_X1 npu_inst_pe_1_3_5_U100 ( .A(npu_inst_pe_1_3_5_n59), .ZN(
        npu_inst_pe_1_3_5_n102) );
  AOI22_X1 npu_inst_pe_1_3_5_U99 ( .A1(npu_inst_int_data_y_4__5__1_), .A2(
        npu_inst_pe_1_3_5_n54), .B1(npu_inst_pe_1_3_5_n118), .B2(
        npu_inst_pe_1_3_5_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_3_5_n55) );
  INV_X1 npu_inst_pe_1_3_5_U98 ( .A(npu_inst_pe_1_3_5_n55), .ZN(
        npu_inst_pe_1_3_5_n103) );
  AOI22_X1 npu_inst_pe_1_3_5_U97 ( .A1(npu_inst_int_data_y_4__5__1_), .A2(
        npu_inst_pe_1_3_5_n50), .B1(npu_inst_pe_1_3_5_n117), .B2(
        npu_inst_pe_1_3_5_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_3_5_n51) );
  INV_X1 npu_inst_pe_1_3_5_U96 ( .A(npu_inst_pe_1_3_5_n51), .ZN(
        npu_inst_pe_1_3_5_n104) );
  AOI22_X1 npu_inst_pe_1_3_5_U95 ( .A1(npu_inst_int_data_y_4__5__1_), .A2(
        npu_inst_pe_1_3_5_n46), .B1(npu_inst_pe_1_3_5_n116), .B2(
        npu_inst_pe_1_3_5_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_3_5_n47) );
  INV_X1 npu_inst_pe_1_3_5_U94 ( .A(npu_inst_pe_1_3_5_n47), .ZN(
        npu_inst_pe_1_3_5_n105) );
  AOI22_X1 npu_inst_pe_1_3_5_U93 ( .A1(npu_inst_int_data_y_4__5__1_), .A2(
        npu_inst_pe_1_3_5_n42), .B1(npu_inst_pe_1_3_5_n115), .B2(
        npu_inst_pe_1_3_5_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_3_5_n43) );
  INV_X1 npu_inst_pe_1_3_5_U92 ( .A(npu_inst_pe_1_3_5_n43), .ZN(
        npu_inst_pe_1_3_5_n106) );
  AOI22_X1 npu_inst_pe_1_3_5_U91 ( .A1(npu_inst_pe_1_3_5_n38), .A2(
        npu_inst_int_data_y_4__5__1_), .B1(npu_inst_pe_1_3_5_n114), .B2(
        npu_inst_pe_1_3_5_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_3_5_n39) );
  INV_X1 npu_inst_pe_1_3_5_U90 ( .A(npu_inst_pe_1_3_5_n39), .ZN(
        npu_inst_pe_1_3_5_n107) );
  AOI22_X1 npu_inst_pe_1_3_5_U89 ( .A1(npu_inst_pe_1_3_5_n38), .A2(
        npu_inst_int_data_y_4__5__0_), .B1(npu_inst_pe_1_3_5_n114), .B2(
        npu_inst_pe_1_3_5_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_3_5_n37) );
  INV_X1 npu_inst_pe_1_3_5_U88 ( .A(npu_inst_pe_1_3_5_n37), .ZN(
        npu_inst_pe_1_3_5_n113) );
  NAND2_X1 npu_inst_pe_1_3_5_U87 ( .A1(npu_inst_pe_1_3_5_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_3_5_n60), .ZN(npu_inst_pe_1_3_5_n74) );
  OAI21_X1 npu_inst_pe_1_3_5_U86 ( .B1(npu_inst_pe_1_3_5_n63), .B2(
        npu_inst_pe_1_3_5_n60), .A(npu_inst_pe_1_3_5_n74), .ZN(
        npu_inst_pe_1_3_5_n97) );
  NAND2_X1 npu_inst_pe_1_3_5_U85 ( .A1(npu_inst_pe_1_3_5_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_3_5_n60), .ZN(npu_inst_pe_1_3_5_n73) );
  OAI21_X1 npu_inst_pe_1_3_5_U84 ( .B1(npu_inst_pe_1_3_5_n61), .B2(
        npu_inst_pe_1_3_5_n60), .A(npu_inst_pe_1_3_5_n73), .ZN(
        npu_inst_pe_1_3_5_n96) );
  NAND2_X1 npu_inst_pe_1_3_5_U83 ( .A1(npu_inst_pe_1_3_5_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_3_5_n56), .ZN(npu_inst_pe_1_3_5_n72) );
  OAI21_X1 npu_inst_pe_1_3_5_U82 ( .B1(npu_inst_pe_1_3_5_n63), .B2(
        npu_inst_pe_1_3_5_n56), .A(npu_inst_pe_1_3_5_n72), .ZN(
        npu_inst_pe_1_3_5_n95) );
  NAND2_X1 npu_inst_pe_1_3_5_U81 ( .A1(npu_inst_pe_1_3_5_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_3_5_n56), .ZN(npu_inst_pe_1_3_5_n71) );
  OAI21_X1 npu_inst_pe_1_3_5_U80 ( .B1(npu_inst_pe_1_3_5_n61), .B2(
        npu_inst_pe_1_3_5_n56), .A(npu_inst_pe_1_3_5_n71), .ZN(
        npu_inst_pe_1_3_5_n94) );
  NAND2_X1 npu_inst_pe_1_3_5_U79 ( .A1(npu_inst_pe_1_3_5_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_3_5_n52), .ZN(npu_inst_pe_1_3_5_n70) );
  OAI21_X1 npu_inst_pe_1_3_5_U78 ( .B1(npu_inst_pe_1_3_5_n63), .B2(
        npu_inst_pe_1_3_5_n52), .A(npu_inst_pe_1_3_5_n70), .ZN(
        npu_inst_pe_1_3_5_n93) );
  NAND2_X1 npu_inst_pe_1_3_5_U77 ( .A1(npu_inst_pe_1_3_5_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_3_5_n52), .ZN(npu_inst_pe_1_3_5_n69) );
  OAI21_X1 npu_inst_pe_1_3_5_U76 ( .B1(npu_inst_pe_1_3_5_n61), .B2(
        npu_inst_pe_1_3_5_n52), .A(npu_inst_pe_1_3_5_n69), .ZN(
        npu_inst_pe_1_3_5_n92) );
  NAND2_X1 npu_inst_pe_1_3_5_U75 ( .A1(npu_inst_pe_1_3_5_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_3_5_n48), .ZN(npu_inst_pe_1_3_5_n68) );
  OAI21_X1 npu_inst_pe_1_3_5_U74 ( .B1(npu_inst_pe_1_3_5_n63), .B2(
        npu_inst_pe_1_3_5_n48), .A(npu_inst_pe_1_3_5_n68), .ZN(
        npu_inst_pe_1_3_5_n91) );
  NAND2_X1 npu_inst_pe_1_3_5_U73 ( .A1(npu_inst_pe_1_3_5_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_3_5_n48), .ZN(npu_inst_pe_1_3_5_n67) );
  OAI21_X1 npu_inst_pe_1_3_5_U72 ( .B1(npu_inst_pe_1_3_5_n61), .B2(
        npu_inst_pe_1_3_5_n48), .A(npu_inst_pe_1_3_5_n67), .ZN(
        npu_inst_pe_1_3_5_n90) );
  NAND2_X1 npu_inst_pe_1_3_5_U71 ( .A1(npu_inst_pe_1_3_5_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_3_5_n44), .ZN(npu_inst_pe_1_3_5_n66) );
  OAI21_X1 npu_inst_pe_1_3_5_U70 ( .B1(npu_inst_pe_1_3_5_n63), .B2(
        npu_inst_pe_1_3_5_n44), .A(npu_inst_pe_1_3_5_n66), .ZN(
        npu_inst_pe_1_3_5_n89) );
  NAND2_X1 npu_inst_pe_1_3_5_U69 ( .A1(npu_inst_pe_1_3_5_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_3_5_n44), .ZN(npu_inst_pe_1_3_5_n65) );
  OAI21_X1 npu_inst_pe_1_3_5_U68 ( .B1(npu_inst_pe_1_3_5_n61), .B2(
        npu_inst_pe_1_3_5_n44), .A(npu_inst_pe_1_3_5_n65), .ZN(
        npu_inst_pe_1_3_5_n88) );
  NAND2_X1 npu_inst_pe_1_3_5_U67 ( .A1(npu_inst_pe_1_3_5_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_3_5_n40), .ZN(npu_inst_pe_1_3_5_n64) );
  OAI21_X1 npu_inst_pe_1_3_5_U66 ( .B1(npu_inst_pe_1_3_5_n63), .B2(
        npu_inst_pe_1_3_5_n40), .A(npu_inst_pe_1_3_5_n64), .ZN(
        npu_inst_pe_1_3_5_n87) );
  NAND2_X1 npu_inst_pe_1_3_5_U65 ( .A1(npu_inst_pe_1_3_5_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_3_5_n40), .ZN(npu_inst_pe_1_3_5_n62) );
  OAI21_X1 npu_inst_pe_1_3_5_U64 ( .B1(npu_inst_pe_1_3_5_n61), .B2(
        npu_inst_pe_1_3_5_n40), .A(npu_inst_pe_1_3_5_n62), .ZN(
        npu_inst_pe_1_3_5_n86) );
  AND2_X1 npu_inst_pe_1_3_5_U63 ( .A1(npu_inst_pe_1_3_5_N93), .A2(npu_inst_n56), .ZN(npu_inst_int_data_y_3__5__0_) );
  AND2_X1 npu_inst_pe_1_3_5_U62 ( .A1(npu_inst_n56), .A2(npu_inst_pe_1_3_5_N94), .ZN(npu_inst_int_data_y_3__5__1_) );
  NOR3_X1 npu_inst_pe_1_3_5_U61 ( .A1(npu_inst_pe_1_3_5_n26), .A2(npu_inst_n56), .A3(npu_inst_int_ckg[34]), .ZN(npu_inst_pe_1_3_5_n85) );
  OR2_X1 npu_inst_pe_1_3_5_U60 ( .A1(npu_inst_pe_1_3_5_n85), .A2(
        npu_inst_pe_1_3_5_n2), .ZN(npu_inst_pe_1_3_5_N84) );
  AND2_X1 npu_inst_pe_1_3_5_U59 ( .A1(npu_inst_pe_1_3_5_int_q_acc_0_), .A2(
        npu_inst_pe_1_3_5_n1), .ZN(npu_inst_int_data_res_3__5__0_) );
  AND2_X1 npu_inst_pe_1_3_5_U58 ( .A1(npu_inst_pe_1_3_5_n2), .A2(
        npu_inst_pe_1_3_5_int_q_acc_7_), .ZN(npu_inst_int_data_res_3__5__7_)
         );
  AND2_X1 npu_inst_pe_1_3_5_U57 ( .A1(npu_inst_pe_1_3_5_int_q_acc_1_), .A2(
        npu_inst_pe_1_3_5_n1), .ZN(npu_inst_int_data_res_3__5__1_) );
  AND2_X1 npu_inst_pe_1_3_5_U56 ( .A1(npu_inst_pe_1_3_5_int_q_acc_2_), .A2(
        npu_inst_pe_1_3_5_n1), .ZN(npu_inst_int_data_res_3__5__2_) );
  AND2_X1 npu_inst_pe_1_3_5_U55 ( .A1(npu_inst_pe_1_3_5_int_q_acc_3_), .A2(
        npu_inst_pe_1_3_5_n2), .ZN(npu_inst_int_data_res_3__5__3_) );
  AND2_X1 npu_inst_pe_1_3_5_U54 ( .A1(npu_inst_pe_1_3_5_int_q_acc_4_), .A2(
        npu_inst_pe_1_3_5_n2), .ZN(npu_inst_int_data_res_3__5__4_) );
  AND2_X1 npu_inst_pe_1_3_5_U53 ( .A1(npu_inst_pe_1_3_5_int_q_acc_5_), .A2(
        npu_inst_pe_1_3_5_n2), .ZN(npu_inst_int_data_res_3__5__5_) );
  AND2_X1 npu_inst_pe_1_3_5_U52 ( .A1(npu_inst_pe_1_3_5_int_q_acc_6_), .A2(
        npu_inst_pe_1_3_5_n2), .ZN(npu_inst_int_data_res_3__5__6_) );
  AOI222_X1 npu_inst_pe_1_3_5_U51 ( .A1(npu_inst_int_data_res_4__5__0_), .A2(
        npu_inst_pe_1_3_5_n1), .B1(npu_inst_pe_1_3_5_N73), .B2(
        npu_inst_pe_1_3_5_n76), .C1(npu_inst_pe_1_3_5_N65), .C2(
        npu_inst_pe_1_3_5_n77), .ZN(npu_inst_pe_1_3_5_n84) );
  INV_X1 npu_inst_pe_1_3_5_U50 ( .A(npu_inst_pe_1_3_5_n84), .ZN(
        npu_inst_pe_1_3_5_n101) );
  AOI222_X1 npu_inst_pe_1_3_5_U49 ( .A1(npu_inst_int_data_res_4__5__7_), .A2(
        npu_inst_pe_1_3_5_n1), .B1(npu_inst_pe_1_3_5_N80), .B2(
        npu_inst_pe_1_3_5_n76), .C1(npu_inst_pe_1_3_5_N72), .C2(
        npu_inst_pe_1_3_5_n77), .ZN(npu_inst_pe_1_3_5_n75) );
  INV_X1 npu_inst_pe_1_3_5_U48 ( .A(npu_inst_pe_1_3_5_n75), .ZN(
        npu_inst_pe_1_3_5_n33) );
  AOI222_X1 npu_inst_pe_1_3_5_U47 ( .A1(npu_inst_int_data_res_4__5__1_), .A2(
        npu_inst_pe_1_3_5_n1), .B1(npu_inst_pe_1_3_5_N74), .B2(
        npu_inst_pe_1_3_5_n76), .C1(npu_inst_pe_1_3_5_N66), .C2(
        npu_inst_pe_1_3_5_n77), .ZN(npu_inst_pe_1_3_5_n83) );
  INV_X1 npu_inst_pe_1_3_5_U46 ( .A(npu_inst_pe_1_3_5_n83), .ZN(
        npu_inst_pe_1_3_5_n100) );
  AOI222_X1 npu_inst_pe_1_3_5_U45 ( .A1(npu_inst_int_data_res_4__5__2_), .A2(
        npu_inst_pe_1_3_5_n1), .B1(npu_inst_pe_1_3_5_N75), .B2(
        npu_inst_pe_1_3_5_n76), .C1(npu_inst_pe_1_3_5_N67), .C2(
        npu_inst_pe_1_3_5_n77), .ZN(npu_inst_pe_1_3_5_n82) );
  INV_X1 npu_inst_pe_1_3_5_U44 ( .A(npu_inst_pe_1_3_5_n82), .ZN(
        npu_inst_pe_1_3_5_n99) );
  AOI222_X1 npu_inst_pe_1_3_5_U43 ( .A1(npu_inst_int_data_res_4__5__3_), .A2(
        npu_inst_pe_1_3_5_n1), .B1(npu_inst_pe_1_3_5_N76), .B2(
        npu_inst_pe_1_3_5_n76), .C1(npu_inst_pe_1_3_5_N68), .C2(
        npu_inst_pe_1_3_5_n77), .ZN(npu_inst_pe_1_3_5_n81) );
  INV_X1 npu_inst_pe_1_3_5_U42 ( .A(npu_inst_pe_1_3_5_n81), .ZN(
        npu_inst_pe_1_3_5_n98) );
  AOI222_X1 npu_inst_pe_1_3_5_U41 ( .A1(npu_inst_int_data_res_4__5__4_), .A2(
        npu_inst_pe_1_3_5_n1), .B1(npu_inst_pe_1_3_5_N77), .B2(
        npu_inst_pe_1_3_5_n76), .C1(npu_inst_pe_1_3_5_N69), .C2(
        npu_inst_pe_1_3_5_n77), .ZN(npu_inst_pe_1_3_5_n80) );
  INV_X1 npu_inst_pe_1_3_5_U40 ( .A(npu_inst_pe_1_3_5_n80), .ZN(
        npu_inst_pe_1_3_5_n36) );
  AOI222_X1 npu_inst_pe_1_3_5_U39 ( .A1(npu_inst_int_data_res_4__5__5_), .A2(
        npu_inst_pe_1_3_5_n1), .B1(npu_inst_pe_1_3_5_N78), .B2(
        npu_inst_pe_1_3_5_n76), .C1(npu_inst_pe_1_3_5_N70), .C2(
        npu_inst_pe_1_3_5_n77), .ZN(npu_inst_pe_1_3_5_n79) );
  INV_X1 npu_inst_pe_1_3_5_U38 ( .A(npu_inst_pe_1_3_5_n79), .ZN(
        npu_inst_pe_1_3_5_n35) );
  AOI222_X1 npu_inst_pe_1_3_5_U37 ( .A1(npu_inst_int_data_res_4__5__6_), .A2(
        npu_inst_pe_1_3_5_n1), .B1(npu_inst_pe_1_3_5_N79), .B2(
        npu_inst_pe_1_3_5_n76), .C1(npu_inst_pe_1_3_5_N71), .C2(
        npu_inst_pe_1_3_5_n77), .ZN(npu_inst_pe_1_3_5_n78) );
  INV_X1 npu_inst_pe_1_3_5_U36 ( .A(npu_inst_pe_1_3_5_n78), .ZN(
        npu_inst_pe_1_3_5_n34) );
  INV_X1 npu_inst_pe_1_3_5_U35 ( .A(npu_inst_pe_1_3_5_int_data_1_), .ZN(
        npu_inst_pe_1_3_5_n14) );
  AND2_X1 npu_inst_pe_1_3_5_U34 ( .A1(npu_inst_int_data_x_3__5__1_), .A2(
        npu_inst_pe_1_3_5_int_q_weight_1_), .ZN(npu_inst_pe_1_3_5_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_3_5_U33 ( .A1(npu_inst_int_data_x_3__5__0_), .A2(
        npu_inst_pe_1_3_5_int_q_weight_1_), .ZN(npu_inst_pe_1_3_5_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_3_5_U32 ( .A1(npu_inst_n56), .A2(
        npu_inst_int_data_y_4__5__1_), .B1(npu_inst_pe_1_3_5_n3), .B2(
        npu_inst_int_data_x_3__6__1_), .ZN(npu_inst_pe_1_3_5_n63) );
  AOI22_X1 npu_inst_pe_1_3_5_U31 ( .A1(npu_inst_n56), .A2(
        npu_inst_int_data_y_4__5__0_), .B1(npu_inst_pe_1_3_5_n3), .B2(
        npu_inst_int_data_x_3__6__0_), .ZN(npu_inst_pe_1_3_5_n61) );
  INV_X1 npu_inst_pe_1_3_5_U30 ( .A(npu_inst_pe_1_3_5_int_data_0_), .ZN(
        npu_inst_pe_1_3_5_n13) );
  INV_X1 npu_inst_pe_1_3_5_U29 ( .A(npu_inst_n69), .ZN(npu_inst_pe_1_3_5_n5)
         );
  OR3_X1 npu_inst_pe_1_3_5_U28 ( .A1(npu_inst_pe_1_3_5_n6), .A2(
        npu_inst_pe_1_3_5_n8), .A3(npu_inst_pe_1_3_5_n5), .ZN(
        npu_inst_pe_1_3_5_n56) );
  OR3_X1 npu_inst_pe_1_3_5_U27 ( .A1(npu_inst_pe_1_3_5_n5), .A2(
        npu_inst_pe_1_3_5_n8), .A3(npu_inst_pe_1_3_5_n7), .ZN(
        npu_inst_pe_1_3_5_n48) );
  INV_X1 npu_inst_pe_1_3_5_U26 ( .A(npu_inst_pe_1_3_5_n5), .ZN(
        npu_inst_pe_1_3_5_n4) );
  OR3_X1 npu_inst_pe_1_3_5_U25 ( .A1(npu_inst_pe_1_3_5_n4), .A2(
        npu_inst_pe_1_3_5_n8), .A3(npu_inst_pe_1_3_5_n7), .ZN(
        npu_inst_pe_1_3_5_n52) );
  OR3_X1 npu_inst_pe_1_3_5_U24 ( .A1(npu_inst_pe_1_3_5_n6), .A2(
        npu_inst_pe_1_3_5_n8), .A3(npu_inst_pe_1_3_5_n4), .ZN(
        npu_inst_pe_1_3_5_n60) );
  NOR2_X1 npu_inst_pe_1_3_5_U23 ( .A1(npu_inst_pe_1_3_5_n60), .A2(
        npu_inst_pe_1_3_5_n3), .ZN(npu_inst_pe_1_3_5_n58) );
  NOR2_X1 npu_inst_pe_1_3_5_U22 ( .A1(npu_inst_pe_1_3_5_n56), .A2(
        npu_inst_pe_1_3_5_n3), .ZN(npu_inst_pe_1_3_5_n54) );
  NOR2_X1 npu_inst_pe_1_3_5_U21 ( .A1(npu_inst_pe_1_3_5_n52), .A2(
        npu_inst_pe_1_3_5_n3), .ZN(npu_inst_pe_1_3_5_n50) );
  NOR2_X1 npu_inst_pe_1_3_5_U20 ( .A1(npu_inst_pe_1_3_5_n48), .A2(
        npu_inst_pe_1_3_5_n3), .ZN(npu_inst_pe_1_3_5_n46) );
  NOR2_X1 npu_inst_pe_1_3_5_U19 ( .A1(npu_inst_pe_1_3_5_n40), .A2(
        npu_inst_pe_1_3_5_n3), .ZN(npu_inst_pe_1_3_5_n38) );
  NOR2_X1 npu_inst_pe_1_3_5_U18 ( .A1(npu_inst_pe_1_3_5_n44), .A2(
        npu_inst_pe_1_3_5_n3), .ZN(npu_inst_pe_1_3_5_n42) );
  BUF_X1 npu_inst_pe_1_3_5_U17 ( .A(npu_inst_n100), .Z(npu_inst_pe_1_3_5_n8)
         );
  INV_X1 npu_inst_pe_1_3_5_U16 ( .A(npu_inst_n124), .ZN(npu_inst_pe_1_3_5_n12)
         );
  INV_X1 npu_inst_pe_1_3_5_U15 ( .A(npu_inst_pe_1_3_5_n38), .ZN(
        npu_inst_pe_1_3_5_n114) );
  INV_X1 npu_inst_pe_1_3_5_U14 ( .A(npu_inst_pe_1_3_5_n58), .ZN(
        npu_inst_pe_1_3_5_n119) );
  INV_X1 npu_inst_pe_1_3_5_U13 ( .A(npu_inst_pe_1_3_5_n54), .ZN(
        npu_inst_pe_1_3_5_n118) );
  INV_X1 npu_inst_pe_1_3_5_U12 ( .A(npu_inst_pe_1_3_5_n50), .ZN(
        npu_inst_pe_1_3_5_n117) );
  INV_X1 npu_inst_pe_1_3_5_U11 ( .A(npu_inst_pe_1_3_5_n46), .ZN(
        npu_inst_pe_1_3_5_n116) );
  INV_X1 npu_inst_pe_1_3_5_U10 ( .A(npu_inst_pe_1_3_5_n42), .ZN(
        npu_inst_pe_1_3_5_n115) );
  BUF_X1 npu_inst_pe_1_3_5_U9 ( .A(npu_inst_n24), .Z(npu_inst_pe_1_3_5_n2) );
  BUF_X1 npu_inst_pe_1_3_5_U8 ( .A(npu_inst_n24), .Z(npu_inst_pe_1_3_5_n1) );
  BUF_X1 npu_inst_pe_1_3_5_U7 ( .A(npu_inst_pe_1_3_5_n12), .Z(
        npu_inst_pe_1_3_5_n11) );
  BUF_X1 npu_inst_pe_1_3_5_U6 ( .A(npu_inst_pe_1_3_5_n12), .Z(
        npu_inst_pe_1_3_5_n10) );
  BUF_X1 npu_inst_pe_1_3_5_U5 ( .A(npu_inst_pe_1_3_5_n12), .Z(
        npu_inst_pe_1_3_5_n9) );
  NOR2_X1 npu_inst_pe_1_3_5_U4 ( .A1(npu_inst_pe_1_3_5_int_q_weight_0_), .A2(
        npu_inst_pe_1_3_5_n1), .ZN(npu_inst_pe_1_3_5_n76) );
  NOR2_X1 npu_inst_pe_1_3_5_U3 ( .A1(npu_inst_pe_1_3_5_n27), .A2(
        npu_inst_pe_1_3_5_n1), .ZN(npu_inst_pe_1_3_5_n77) );
  FA_X1 npu_inst_pe_1_3_5_sub_67_U2_1 ( .A(npu_inst_pe_1_3_5_int_q_acc_1_), 
        .B(npu_inst_pe_1_3_5_n14), .CI(npu_inst_pe_1_3_5_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_3_5_sub_67_carry_2_), .S(npu_inst_pe_1_3_5_N66) );
  FA_X1 npu_inst_pe_1_3_5_add_69_U1_1 ( .A(npu_inst_pe_1_3_5_int_q_acc_1_), 
        .B(npu_inst_pe_1_3_5_int_data_1_), .CI(
        npu_inst_pe_1_3_5_add_69_carry_1_), .CO(
        npu_inst_pe_1_3_5_add_69_carry_2_), .S(npu_inst_pe_1_3_5_N74) );
  NAND3_X1 npu_inst_pe_1_3_5_U109 ( .A1(npu_inst_pe_1_3_5_n5), .A2(
        npu_inst_pe_1_3_5_n7), .A3(npu_inst_pe_1_3_5_n8), .ZN(
        npu_inst_pe_1_3_5_n44) );
  NAND3_X1 npu_inst_pe_1_3_5_U108 ( .A1(npu_inst_pe_1_3_5_n4), .A2(
        npu_inst_pe_1_3_5_n7), .A3(npu_inst_pe_1_3_5_n8), .ZN(
        npu_inst_pe_1_3_5_n40) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_3_5_n34), .CK(
        npu_inst_pe_1_3_5_net3895), .RN(npu_inst_pe_1_3_5_n9), .Q(
        npu_inst_pe_1_3_5_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_3_5_n35), .CK(
        npu_inst_pe_1_3_5_net3895), .RN(npu_inst_pe_1_3_5_n9), .Q(
        npu_inst_pe_1_3_5_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_3_5_n36), .CK(
        npu_inst_pe_1_3_5_net3895), .RN(npu_inst_pe_1_3_5_n9), .Q(
        npu_inst_pe_1_3_5_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_3_5_n98), .CK(
        npu_inst_pe_1_3_5_net3895), .RN(npu_inst_pe_1_3_5_n9), .Q(
        npu_inst_pe_1_3_5_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_3_5_n99), .CK(
        npu_inst_pe_1_3_5_net3895), .RN(npu_inst_pe_1_3_5_n9), .Q(
        npu_inst_pe_1_3_5_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_3_5_n100), 
        .CK(npu_inst_pe_1_3_5_net3895), .RN(npu_inst_pe_1_3_5_n9), .Q(
        npu_inst_pe_1_3_5_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_3_5_n33), .CK(
        npu_inst_pe_1_3_5_net3895), .RN(npu_inst_pe_1_3_5_n9), .Q(
        npu_inst_pe_1_3_5_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_3_5_n101), 
        .CK(npu_inst_pe_1_3_5_net3895), .RN(npu_inst_pe_1_3_5_n9), .Q(
        npu_inst_pe_1_3_5_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_weight_reg_0_ ( .D(npu_inst_n110), .CK(
        npu_inst_pe_1_3_5_net3901), .RN(npu_inst_pe_1_3_5_n9), .Q(
        npu_inst_pe_1_3_5_int_q_weight_0_), .QN(npu_inst_pe_1_3_5_n27) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_weight_reg_1_ ( .D(npu_inst_n116), .CK(
        npu_inst_pe_1_3_5_net3901), .RN(npu_inst_pe_1_3_5_n9), .Q(
        npu_inst_pe_1_3_5_int_q_weight_1_), .QN(npu_inst_pe_1_3_5_n26) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_3_5_n113), 
        .CK(npu_inst_pe_1_3_5_net3901), .RN(npu_inst_pe_1_3_5_n9), .Q(
        npu_inst_pe_1_3_5_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_3_5_n107), 
        .CK(npu_inst_pe_1_3_5_net3901), .RN(npu_inst_pe_1_3_5_n9), .Q(
        npu_inst_pe_1_3_5_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_3_5_n112), 
        .CK(npu_inst_pe_1_3_5_net3901), .RN(npu_inst_pe_1_3_5_n10), .Q(
        npu_inst_pe_1_3_5_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_3_5_n106), 
        .CK(npu_inst_pe_1_3_5_net3901), .RN(npu_inst_pe_1_3_5_n10), .Q(
        npu_inst_pe_1_3_5_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_3_5_n111), 
        .CK(npu_inst_pe_1_3_5_net3901), .RN(npu_inst_pe_1_3_5_n10), .Q(
        npu_inst_pe_1_3_5_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_3_5_n105), 
        .CK(npu_inst_pe_1_3_5_net3901), .RN(npu_inst_pe_1_3_5_n10), .Q(
        npu_inst_pe_1_3_5_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_3_5_n110), 
        .CK(npu_inst_pe_1_3_5_net3901), .RN(npu_inst_pe_1_3_5_n10), .Q(
        npu_inst_pe_1_3_5_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_3_5_n104), 
        .CK(npu_inst_pe_1_3_5_net3901), .RN(npu_inst_pe_1_3_5_n10), .Q(
        npu_inst_pe_1_3_5_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_3_5_n109), 
        .CK(npu_inst_pe_1_3_5_net3901), .RN(npu_inst_pe_1_3_5_n10), .Q(
        npu_inst_pe_1_3_5_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_3_5_n103), 
        .CK(npu_inst_pe_1_3_5_net3901), .RN(npu_inst_pe_1_3_5_n10), .Q(
        npu_inst_pe_1_3_5_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_3_5_n108), 
        .CK(npu_inst_pe_1_3_5_net3901), .RN(npu_inst_pe_1_3_5_n10), .Q(
        npu_inst_pe_1_3_5_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_3_5_n102), 
        .CK(npu_inst_pe_1_3_5_net3901), .RN(npu_inst_pe_1_3_5_n10), .Q(
        npu_inst_pe_1_3_5_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_3_5_n86), 
        .CK(npu_inst_pe_1_3_5_net3901), .RN(npu_inst_pe_1_3_5_n10), .Q(
        npu_inst_pe_1_3_5_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_3_5_n87), 
        .CK(npu_inst_pe_1_3_5_net3901), .RN(npu_inst_pe_1_3_5_n10), .Q(
        npu_inst_pe_1_3_5_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_3_5_n88), 
        .CK(npu_inst_pe_1_3_5_net3901), .RN(npu_inst_pe_1_3_5_n11), .Q(
        npu_inst_pe_1_3_5_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_3_5_n89), 
        .CK(npu_inst_pe_1_3_5_net3901), .RN(npu_inst_pe_1_3_5_n11), .Q(
        npu_inst_pe_1_3_5_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_3_5_n90), 
        .CK(npu_inst_pe_1_3_5_net3901), .RN(npu_inst_pe_1_3_5_n11), .Q(
        npu_inst_pe_1_3_5_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_3_5_n91), 
        .CK(npu_inst_pe_1_3_5_net3901), .RN(npu_inst_pe_1_3_5_n11), .Q(
        npu_inst_pe_1_3_5_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_3_5_n92), 
        .CK(npu_inst_pe_1_3_5_net3901), .RN(npu_inst_pe_1_3_5_n11), .Q(
        npu_inst_pe_1_3_5_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_3_5_n93), 
        .CK(npu_inst_pe_1_3_5_net3901), .RN(npu_inst_pe_1_3_5_n11), .Q(
        npu_inst_pe_1_3_5_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_3_5_n94), 
        .CK(npu_inst_pe_1_3_5_net3901), .RN(npu_inst_pe_1_3_5_n11), .Q(
        npu_inst_pe_1_3_5_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_3_5_n95), 
        .CK(npu_inst_pe_1_3_5_net3901), .RN(npu_inst_pe_1_3_5_n11), .Q(
        npu_inst_pe_1_3_5_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_3_5_n96), 
        .CK(npu_inst_pe_1_3_5_net3901), .RN(npu_inst_pe_1_3_5_n11), .Q(
        npu_inst_pe_1_3_5_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_3_5_n97), 
        .CK(npu_inst_pe_1_3_5_net3901), .RN(npu_inst_pe_1_3_5_n11), .Q(
        npu_inst_pe_1_3_5_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_3_5_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_3_5_N84), .SE(1'b0), .GCK(npu_inst_pe_1_3_5_net3895) );
  CLKGATETST_X1 npu_inst_pe_1_3_5_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n64), .SE(1'b0), .GCK(npu_inst_pe_1_3_5_net3901) );
  MUX2_X1 npu_inst_pe_1_3_6_U162 ( .A(npu_inst_pe_1_3_6_n32), .B(
        npu_inst_pe_1_3_6_n29), .S(npu_inst_pe_1_3_6_n8), .Z(
        npu_inst_pe_1_3_6_N93) );
  MUX2_X1 npu_inst_pe_1_3_6_U161 ( .A(npu_inst_pe_1_3_6_n31), .B(
        npu_inst_pe_1_3_6_n30), .S(npu_inst_pe_1_3_6_n6), .Z(
        npu_inst_pe_1_3_6_n32) );
  MUX2_X1 npu_inst_pe_1_3_6_U160 ( .A(npu_inst_pe_1_3_6_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_3_6_int_q_reg_v_1__0_), .S(npu_inst_pe_1_3_6_n4), .Z(
        npu_inst_pe_1_3_6_n31) );
  MUX2_X1 npu_inst_pe_1_3_6_U159 ( .A(npu_inst_pe_1_3_6_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_3_6_int_q_reg_v_3__0_), .S(npu_inst_pe_1_3_6_n4), .Z(
        npu_inst_pe_1_3_6_n30) );
  MUX2_X1 npu_inst_pe_1_3_6_U158 ( .A(npu_inst_pe_1_3_6_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_3_6_int_q_reg_v_5__0_), .S(npu_inst_pe_1_3_6_n4), .Z(
        npu_inst_pe_1_3_6_n29) );
  MUX2_X1 npu_inst_pe_1_3_6_U157 ( .A(npu_inst_pe_1_3_6_n28), .B(
        npu_inst_pe_1_3_6_n23), .S(npu_inst_pe_1_3_6_n8), .Z(
        npu_inst_pe_1_3_6_N94) );
  MUX2_X1 npu_inst_pe_1_3_6_U156 ( .A(npu_inst_pe_1_3_6_n25), .B(
        npu_inst_pe_1_3_6_n24), .S(npu_inst_pe_1_3_6_n6), .Z(
        npu_inst_pe_1_3_6_n28) );
  MUX2_X1 npu_inst_pe_1_3_6_U155 ( .A(npu_inst_pe_1_3_6_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_3_6_int_q_reg_v_1__1_), .S(npu_inst_pe_1_3_6_n4), .Z(
        npu_inst_pe_1_3_6_n25) );
  MUX2_X1 npu_inst_pe_1_3_6_U154 ( .A(npu_inst_pe_1_3_6_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_3_6_int_q_reg_v_3__1_), .S(npu_inst_pe_1_3_6_n4), .Z(
        npu_inst_pe_1_3_6_n24) );
  MUX2_X1 npu_inst_pe_1_3_6_U153 ( .A(npu_inst_pe_1_3_6_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_3_6_int_q_reg_v_5__1_), .S(npu_inst_pe_1_3_6_n4), .Z(
        npu_inst_pe_1_3_6_n23) );
  MUX2_X1 npu_inst_pe_1_3_6_U152 ( .A(npu_inst_pe_1_3_6_n22), .B(
        npu_inst_pe_1_3_6_n19), .S(npu_inst_pe_1_3_6_n8), .Z(
        npu_inst_int_data_x_3__6__1_) );
  MUX2_X1 npu_inst_pe_1_3_6_U151 ( .A(npu_inst_pe_1_3_6_n21), .B(
        npu_inst_pe_1_3_6_n20), .S(npu_inst_pe_1_3_6_n6), .Z(
        npu_inst_pe_1_3_6_n22) );
  MUX2_X1 npu_inst_pe_1_3_6_U150 ( .A(npu_inst_pe_1_3_6_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_3_6_int_q_reg_h_1__1_), .S(npu_inst_pe_1_3_6_n4), .Z(
        npu_inst_pe_1_3_6_n21) );
  MUX2_X1 npu_inst_pe_1_3_6_U149 ( .A(npu_inst_pe_1_3_6_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_3_6_int_q_reg_h_3__1_), .S(npu_inst_pe_1_3_6_n4), .Z(
        npu_inst_pe_1_3_6_n20) );
  MUX2_X1 npu_inst_pe_1_3_6_U148 ( .A(npu_inst_pe_1_3_6_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_3_6_int_q_reg_h_5__1_), .S(npu_inst_pe_1_3_6_n4), .Z(
        npu_inst_pe_1_3_6_n19) );
  MUX2_X1 npu_inst_pe_1_3_6_U147 ( .A(npu_inst_pe_1_3_6_n18), .B(
        npu_inst_pe_1_3_6_n15), .S(npu_inst_pe_1_3_6_n8), .Z(
        npu_inst_int_data_x_3__6__0_) );
  MUX2_X1 npu_inst_pe_1_3_6_U146 ( .A(npu_inst_pe_1_3_6_n17), .B(
        npu_inst_pe_1_3_6_n16), .S(npu_inst_pe_1_3_6_n6), .Z(
        npu_inst_pe_1_3_6_n18) );
  MUX2_X1 npu_inst_pe_1_3_6_U145 ( .A(npu_inst_pe_1_3_6_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_3_6_int_q_reg_h_1__0_), .S(npu_inst_pe_1_3_6_n4), .Z(
        npu_inst_pe_1_3_6_n17) );
  MUX2_X1 npu_inst_pe_1_3_6_U144 ( .A(npu_inst_pe_1_3_6_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_3_6_int_q_reg_h_3__0_), .S(npu_inst_pe_1_3_6_n4), .Z(
        npu_inst_pe_1_3_6_n16) );
  MUX2_X1 npu_inst_pe_1_3_6_U143 ( .A(npu_inst_pe_1_3_6_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_3_6_int_q_reg_h_5__0_), .S(npu_inst_pe_1_3_6_n4), .Z(
        npu_inst_pe_1_3_6_n15) );
  XOR2_X1 npu_inst_pe_1_3_6_U142 ( .A(npu_inst_pe_1_3_6_int_data_0_), .B(
        npu_inst_pe_1_3_6_int_q_acc_0_), .Z(npu_inst_pe_1_3_6_N73) );
  AND2_X1 npu_inst_pe_1_3_6_U141 ( .A1(npu_inst_pe_1_3_6_int_q_acc_0_), .A2(
        npu_inst_pe_1_3_6_int_data_0_), .ZN(npu_inst_pe_1_3_6_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_3_6_U140 ( .A(npu_inst_pe_1_3_6_int_q_acc_0_), .B(
        npu_inst_pe_1_3_6_n13), .ZN(npu_inst_pe_1_3_6_N65) );
  OR2_X1 npu_inst_pe_1_3_6_U139 ( .A1(npu_inst_pe_1_3_6_n13), .A2(
        npu_inst_pe_1_3_6_int_q_acc_0_), .ZN(npu_inst_pe_1_3_6_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_3_6_U138 ( .A(npu_inst_pe_1_3_6_int_q_acc_2_), .B(
        npu_inst_pe_1_3_6_add_69_carry_2_), .Z(npu_inst_pe_1_3_6_N75) );
  AND2_X1 npu_inst_pe_1_3_6_U137 ( .A1(npu_inst_pe_1_3_6_add_69_carry_2_), 
        .A2(npu_inst_pe_1_3_6_int_q_acc_2_), .ZN(
        npu_inst_pe_1_3_6_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_3_6_U136 ( .A(npu_inst_pe_1_3_6_int_q_acc_3_), .B(
        npu_inst_pe_1_3_6_add_69_carry_3_), .Z(npu_inst_pe_1_3_6_N76) );
  AND2_X1 npu_inst_pe_1_3_6_U135 ( .A1(npu_inst_pe_1_3_6_add_69_carry_3_), 
        .A2(npu_inst_pe_1_3_6_int_q_acc_3_), .ZN(
        npu_inst_pe_1_3_6_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_3_6_U134 ( .A(npu_inst_pe_1_3_6_int_q_acc_4_), .B(
        npu_inst_pe_1_3_6_add_69_carry_4_), .Z(npu_inst_pe_1_3_6_N77) );
  AND2_X1 npu_inst_pe_1_3_6_U133 ( .A1(npu_inst_pe_1_3_6_add_69_carry_4_), 
        .A2(npu_inst_pe_1_3_6_int_q_acc_4_), .ZN(
        npu_inst_pe_1_3_6_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_3_6_U132 ( .A(npu_inst_pe_1_3_6_int_q_acc_5_), .B(
        npu_inst_pe_1_3_6_add_69_carry_5_), .Z(npu_inst_pe_1_3_6_N78) );
  AND2_X1 npu_inst_pe_1_3_6_U131 ( .A1(npu_inst_pe_1_3_6_add_69_carry_5_), 
        .A2(npu_inst_pe_1_3_6_int_q_acc_5_), .ZN(
        npu_inst_pe_1_3_6_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_3_6_U130 ( .A(npu_inst_pe_1_3_6_int_q_acc_6_), .B(
        npu_inst_pe_1_3_6_add_69_carry_6_), .Z(npu_inst_pe_1_3_6_N79) );
  AND2_X1 npu_inst_pe_1_3_6_U129 ( .A1(npu_inst_pe_1_3_6_add_69_carry_6_), 
        .A2(npu_inst_pe_1_3_6_int_q_acc_6_), .ZN(
        npu_inst_pe_1_3_6_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_3_6_U128 ( .A(npu_inst_pe_1_3_6_int_q_acc_7_), .B(
        npu_inst_pe_1_3_6_add_69_carry_7_), .Z(npu_inst_pe_1_3_6_N80) );
  XNOR2_X1 npu_inst_pe_1_3_6_U127 ( .A(npu_inst_pe_1_3_6_sub_67_carry_2_), .B(
        npu_inst_pe_1_3_6_int_q_acc_2_), .ZN(npu_inst_pe_1_3_6_N67) );
  OR2_X1 npu_inst_pe_1_3_6_U126 ( .A1(npu_inst_pe_1_3_6_int_q_acc_2_), .A2(
        npu_inst_pe_1_3_6_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_3_6_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_3_6_U125 ( .A(npu_inst_pe_1_3_6_sub_67_carry_3_), .B(
        npu_inst_pe_1_3_6_int_q_acc_3_), .ZN(npu_inst_pe_1_3_6_N68) );
  OR2_X1 npu_inst_pe_1_3_6_U124 ( .A1(npu_inst_pe_1_3_6_int_q_acc_3_), .A2(
        npu_inst_pe_1_3_6_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_3_6_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_3_6_U123 ( .A(npu_inst_pe_1_3_6_sub_67_carry_4_), .B(
        npu_inst_pe_1_3_6_int_q_acc_4_), .ZN(npu_inst_pe_1_3_6_N69) );
  OR2_X1 npu_inst_pe_1_3_6_U122 ( .A1(npu_inst_pe_1_3_6_int_q_acc_4_), .A2(
        npu_inst_pe_1_3_6_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_3_6_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_3_6_U121 ( .A(npu_inst_pe_1_3_6_sub_67_carry_5_), .B(
        npu_inst_pe_1_3_6_int_q_acc_5_), .ZN(npu_inst_pe_1_3_6_N70) );
  OR2_X1 npu_inst_pe_1_3_6_U120 ( .A1(npu_inst_pe_1_3_6_int_q_acc_5_), .A2(
        npu_inst_pe_1_3_6_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_3_6_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_3_6_U119 ( .A(npu_inst_pe_1_3_6_sub_67_carry_6_), .B(
        npu_inst_pe_1_3_6_int_q_acc_6_), .ZN(npu_inst_pe_1_3_6_N71) );
  OR2_X1 npu_inst_pe_1_3_6_U118 ( .A1(npu_inst_pe_1_3_6_int_q_acc_6_), .A2(
        npu_inst_pe_1_3_6_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_3_6_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_3_6_U117 ( .A(npu_inst_pe_1_3_6_int_q_acc_7_), .B(
        npu_inst_pe_1_3_6_sub_67_carry_7_), .ZN(npu_inst_pe_1_3_6_N72) );
  INV_X1 npu_inst_pe_1_3_6_U116 ( .A(npu_inst_n77), .ZN(npu_inst_pe_1_3_6_n7)
         );
  INV_X1 npu_inst_pe_1_3_6_U115 ( .A(npu_inst_pe_1_3_6_n7), .ZN(
        npu_inst_pe_1_3_6_n6) );
  INV_X1 npu_inst_pe_1_3_6_U114 ( .A(npu_inst_n56), .ZN(npu_inst_pe_1_3_6_n3)
         );
  AOI22_X1 npu_inst_pe_1_3_6_U113 ( .A1(npu_inst_int_data_y_4__6__0_), .A2(
        npu_inst_pe_1_3_6_n58), .B1(npu_inst_pe_1_3_6_n119), .B2(
        npu_inst_pe_1_3_6_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_3_6_n57) );
  INV_X1 npu_inst_pe_1_3_6_U112 ( .A(npu_inst_pe_1_3_6_n57), .ZN(
        npu_inst_pe_1_3_6_n108) );
  AOI22_X1 npu_inst_pe_1_3_6_U111 ( .A1(npu_inst_int_data_y_4__6__0_), .A2(
        npu_inst_pe_1_3_6_n54), .B1(npu_inst_pe_1_3_6_n118), .B2(
        npu_inst_pe_1_3_6_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_3_6_n53) );
  INV_X1 npu_inst_pe_1_3_6_U110 ( .A(npu_inst_pe_1_3_6_n53), .ZN(
        npu_inst_pe_1_3_6_n109) );
  AOI22_X1 npu_inst_pe_1_3_6_U107 ( .A1(npu_inst_int_data_y_4__6__0_), .A2(
        npu_inst_pe_1_3_6_n50), .B1(npu_inst_pe_1_3_6_n117), .B2(
        npu_inst_pe_1_3_6_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_3_6_n49) );
  INV_X1 npu_inst_pe_1_3_6_U106 ( .A(npu_inst_pe_1_3_6_n49), .ZN(
        npu_inst_pe_1_3_6_n110) );
  AOI22_X1 npu_inst_pe_1_3_6_U105 ( .A1(npu_inst_int_data_y_4__6__0_), .A2(
        npu_inst_pe_1_3_6_n46), .B1(npu_inst_pe_1_3_6_n116), .B2(
        npu_inst_pe_1_3_6_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_3_6_n45) );
  INV_X1 npu_inst_pe_1_3_6_U104 ( .A(npu_inst_pe_1_3_6_n45), .ZN(
        npu_inst_pe_1_3_6_n111) );
  AOI22_X1 npu_inst_pe_1_3_6_U103 ( .A1(npu_inst_int_data_y_4__6__0_), .A2(
        npu_inst_pe_1_3_6_n42), .B1(npu_inst_pe_1_3_6_n115), .B2(
        npu_inst_pe_1_3_6_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_3_6_n41) );
  INV_X1 npu_inst_pe_1_3_6_U102 ( .A(npu_inst_pe_1_3_6_n41), .ZN(
        npu_inst_pe_1_3_6_n112) );
  AOI22_X1 npu_inst_pe_1_3_6_U101 ( .A1(npu_inst_int_data_y_4__6__1_), .A2(
        npu_inst_pe_1_3_6_n58), .B1(npu_inst_pe_1_3_6_n119), .B2(
        npu_inst_pe_1_3_6_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_3_6_n59) );
  INV_X1 npu_inst_pe_1_3_6_U100 ( .A(npu_inst_pe_1_3_6_n59), .ZN(
        npu_inst_pe_1_3_6_n102) );
  AOI22_X1 npu_inst_pe_1_3_6_U99 ( .A1(npu_inst_int_data_y_4__6__1_), .A2(
        npu_inst_pe_1_3_6_n54), .B1(npu_inst_pe_1_3_6_n118), .B2(
        npu_inst_pe_1_3_6_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_3_6_n55) );
  INV_X1 npu_inst_pe_1_3_6_U98 ( .A(npu_inst_pe_1_3_6_n55), .ZN(
        npu_inst_pe_1_3_6_n103) );
  AOI22_X1 npu_inst_pe_1_3_6_U97 ( .A1(npu_inst_int_data_y_4__6__1_), .A2(
        npu_inst_pe_1_3_6_n50), .B1(npu_inst_pe_1_3_6_n117), .B2(
        npu_inst_pe_1_3_6_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_3_6_n51) );
  INV_X1 npu_inst_pe_1_3_6_U96 ( .A(npu_inst_pe_1_3_6_n51), .ZN(
        npu_inst_pe_1_3_6_n104) );
  AOI22_X1 npu_inst_pe_1_3_6_U95 ( .A1(npu_inst_int_data_y_4__6__1_), .A2(
        npu_inst_pe_1_3_6_n46), .B1(npu_inst_pe_1_3_6_n116), .B2(
        npu_inst_pe_1_3_6_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_3_6_n47) );
  INV_X1 npu_inst_pe_1_3_6_U94 ( .A(npu_inst_pe_1_3_6_n47), .ZN(
        npu_inst_pe_1_3_6_n105) );
  AOI22_X1 npu_inst_pe_1_3_6_U93 ( .A1(npu_inst_int_data_y_4__6__1_), .A2(
        npu_inst_pe_1_3_6_n42), .B1(npu_inst_pe_1_3_6_n115), .B2(
        npu_inst_pe_1_3_6_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_3_6_n43) );
  INV_X1 npu_inst_pe_1_3_6_U92 ( .A(npu_inst_pe_1_3_6_n43), .ZN(
        npu_inst_pe_1_3_6_n106) );
  AOI22_X1 npu_inst_pe_1_3_6_U91 ( .A1(npu_inst_pe_1_3_6_n38), .A2(
        npu_inst_int_data_y_4__6__1_), .B1(npu_inst_pe_1_3_6_n114), .B2(
        npu_inst_pe_1_3_6_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_3_6_n39) );
  INV_X1 npu_inst_pe_1_3_6_U90 ( .A(npu_inst_pe_1_3_6_n39), .ZN(
        npu_inst_pe_1_3_6_n107) );
  AOI22_X1 npu_inst_pe_1_3_6_U89 ( .A1(npu_inst_pe_1_3_6_n38), .A2(
        npu_inst_int_data_y_4__6__0_), .B1(npu_inst_pe_1_3_6_n114), .B2(
        npu_inst_pe_1_3_6_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_3_6_n37) );
  INV_X1 npu_inst_pe_1_3_6_U88 ( .A(npu_inst_pe_1_3_6_n37), .ZN(
        npu_inst_pe_1_3_6_n113) );
  NAND2_X1 npu_inst_pe_1_3_6_U87 ( .A1(npu_inst_pe_1_3_6_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_3_6_n60), .ZN(npu_inst_pe_1_3_6_n74) );
  OAI21_X1 npu_inst_pe_1_3_6_U86 ( .B1(npu_inst_pe_1_3_6_n63), .B2(
        npu_inst_pe_1_3_6_n60), .A(npu_inst_pe_1_3_6_n74), .ZN(
        npu_inst_pe_1_3_6_n97) );
  NAND2_X1 npu_inst_pe_1_3_6_U85 ( .A1(npu_inst_pe_1_3_6_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_3_6_n60), .ZN(npu_inst_pe_1_3_6_n73) );
  OAI21_X1 npu_inst_pe_1_3_6_U84 ( .B1(npu_inst_pe_1_3_6_n61), .B2(
        npu_inst_pe_1_3_6_n60), .A(npu_inst_pe_1_3_6_n73), .ZN(
        npu_inst_pe_1_3_6_n96) );
  NAND2_X1 npu_inst_pe_1_3_6_U83 ( .A1(npu_inst_pe_1_3_6_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_3_6_n56), .ZN(npu_inst_pe_1_3_6_n72) );
  OAI21_X1 npu_inst_pe_1_3_6_U82 ( .B1(npu_inst_pe_1_3_6_n63), .B2(
        npu_inst_pe_1_3_6_n56), .A(npu_inst_pe_1_3_6_n72), .ZN(
        npu_inst_pe_1_3_6_n95) );
  NAND2_X1 npu_inst_pe_1_3_6_U81 ( .A1(npu_inst_pe_1_3_6_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_3_6_n56), .ZN(npu_inst_pe_1_3_6_n71) );
  OAI21_X1 npu_inst_pe_1_3_6_U80 ( .B1(npu_inst_pe_1_3_6_n61), .B2(
        npu_inst_pe_1_3_6_n56), .A(npu_inst_pe_1_3_6_n71), .ZN(
        npu_inst_pe_1_3_6_n94) );
  NAND2_X1 npu_inst_pe_1_3_6_U79 ( .A1(npu_inst_pe_1_3_6_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_3_6_n52), .ZN(npu_inst_pe_1_3_6_n70) );
  OAI21_X1 npu_inst_pe_1_3_6_U78 ( .B1(npu_inst_pe_1_3_6_n63), .B2(
        npu_inst_pe_1_3_6_n52), .A(npu_inst_pe_1_3_6_n70), .ZN(
        npu_inst_pe_1_3_6_n93) );
  NAND2_X1 npu_inst_pe_1_3_6_U77 ( .A1(npu_inst_pe_1_3_6_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_3_6_n52), .ZN(npu_inst_pe_1_3_6_n69) );
  OAI21_X1 npu_inst_pe_1_3_6_U76 ( .B1(npu_inst_pe_1_3_6_n61), .B2(
        npu_inst_pe_1_3_6_n52), .A(npu_inst_pe_1_3_6_n69), .ZN(
        npu_inst_pe_1_3_6_n92) );
  NAND2_X1 npu_inst_pe_1_3_6_U75 ( .A1(npu_inst_pe_1_3_6_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_3_6_n48), .ZN(npu_inst_pe_1_3_6_n68) );
  OAI21_X1 npu_inst_pe_1_3_6_U74 ( .B1(npu_inst_pe_1_3_6_n63), .B2(
        npu_inst_pe_1_3_6_n48), .A(npu_inst_pe_1_3_6_n68), .ZN(
        npu_inst_pe_1_3_6_n91) );
  NAND2_X1 npu_inst_pe_1_3_6_U73 ( .A1(npu_inst_pe_1_3_6_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_3_6_n48), .ZN(npu_inst_pe_1_3_6_n67) );
  OAI21_X1 npu_inst_pe_1_3_6_U72 ( .B1(npu_inst_pe_1_3_6_n61), .B2(
        npu_inst_pe_1_3_6_n48), .A(npu_inst_pe_1_3_6_n67), .ZN(
        npu_inst_pe_1_3_6_n90) );
  NAND2_X1 npu_inst_pe_1_3_6_U71 ( .A1(npu_inst_pe_1_3_6_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_3_6_n44), .ZN(npu_inst_pe_1_3_6_n66) );
  OAI21_X1 npu_inst_pe_1_3_6_U70 ( .B1(npu_inst_pe_1_3_6_n63), .B2(
        npu_inst_pe_1_3_6_n44), .A(npu_inst_pe_1_3_6_n66), .ZN(
        npu_inst_pe_1_3_6_n89) );
  NAND2_X1 npu_inst_pe_1_3_6_U69 ( .A1(npu_inst_pe_1_3_6_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_3_6_n44), .ZN(npu_inst_pe_1_3_6_n65) );
  OAI21_X1 npu_inst_pe_1_3_6_U68 ( .B1(npu_inst_pe_1_3_6_n61), .B2(
        npu_inst_pe_1_3_6_n44), .A(npu_inst_pe_1_3_6_n65), .ZN(
        npu_inst_pe_1_3_6_n88) );
  NAND2_X1 npu_inst_pe_1_3_6_U67 ( .A1(npu_inst_pe_1_3_6_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_3_6_n40), .ZN(npu_inst_pe_1_3_6_n64) );
  OAI21_X1 npu_inst_pe_1_3_6_U66 ( .B1(npu_inst_pe_1_3_6_n63), .B2(
        npu_inst_pe_1_3_6_n40), .A(npu_inst_pe_1_3_6_n64), .ZN(
        npu_inst_pe_1_3_6_n87) );
  NAND2_X1 npu_inst_pe_1_3_6_U65 ( .A1(npu_inst_pe_1_3_6_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_3_6_n40), .ZN(npu_inst_pe_1_3_6_n62) );
  OAI21_X1 npu_inst_pe_1_3_6_U64 ( .B1(npu_inst_pe_1_3_6_n61), .B2(
        npu_inst_pe_1_3_6_n40), .A(npu_inst_pe_1_3_6_n62), .ZN(
        npu_inst_pe_1_3_6_n86) );
  AND2_X1 npu_inst_pe_1_3_6_U63 ( .A1(npu_inst_pe_1_3_6_N93), .A2(npu_inst_n56), .ZN(npu_inst_int_data_y_3__6__0_) );
  AND2_X1 npu_inst_pe_1_3_6_U62 ( .A1(npu_inst_n56), .A2(npu_inst_pe_1_3_6_N94), .ZN(npu_inst_int_data_y_3__6__1_) );
  NOR3_X1 npu_inst_pe_1_3_6_U61 ( .A1(npu_inst_pe_1_3_6_n26), .A2(npu_inst_n56), .A3(npu_inst_int_ckg[33]), .ZN(npu_inst_pe_1_3_6_n85) );
  OR2_X1 npu_inst_pe_1_3_6_U60 ( .A1(npu_inst_pe_1_3_6_n85), .A2(
        npu_inst_pe_1_3_6_n2), .ZN(npu_inst_pe_1_3_6_N84) );
  AND2_X1 npu_inst_pe_1_3_6_U59 ( .A1(npu_inst_pe_1_3_6_int_q_acc_0_), .A2(
        npu_inst_pe_1_3_6_n1), .ZN(npu_inst_int_data_res_3__6__0_) );
  AND2_X1 npu_inst_pe_1_3_6_U58 ( .A1(npu_inst_pe_1_3_6_n2), .A2(
        npu_inst_pe_1_3_6_int_q_acc_7_), .ZN(npu_inst_int_data_res_3__6__7_)
         );
  AND2_X1 npu_inst_pe_1_3_6_U57 ( .A1(npu_inst_pe_1_3_6_int_q_acc_1_), .A2(
        npu_inst_pe_1_3_6_n1), .ZN(npu_inst_int_data_res_3__6__1_) );
  AND2_X1 npu_inst_pe_1_3_6_U56 ( .A1(npu_inst_pe_1_3_6_int_q_acc_2_), .A2(
        npu_inst_pe_1_3_6_n1), .ZN(npu_inst_int_data_res_3__6__2_) );
  AND2_X1 npu_inst_pe_1_3_6_U55 ( .A1(npu_inst_pe_1_3_6_int_q_acc_3_), .A2(
        npu_inst_pe_1_3_6_n2), .ZN(npu_inst_int_data_res_3__6__3_) );
  AND2_X1 npu_inst_pe_1_3_6_U54 ( .A1(npu_inst_pe_1_3_6_int_q_acc_4_), .A2(
        npu_inst_pe_1_3_6_n2), .ZN(npu_inst_int_data_res_3__6__4_) );
  AND2_X1 npu_inst_pe_1_3_6_U53 ( .A1(npu_inst_pe_1_3_6_int_q_acc_5_), .A2(
        npu_inst_pe_1_3_6_n2), .ZN(npu_inst_int_data_res_3__6__5_) );
  AND2_X1 npu_inst_pe_1_3_6_U52 ( .A1(npu_inst_pe_1_3_6_int_q_acc_6_), .A2(
        npu_inst_pe_1_3_6_n2), .ZN(npu_inst_int_data_res_3__6__6_) );
  AOI222_X1 npu_inst_pe_1_3_6_U51 ( .A1(npu_inst_int_data_res_4__6__0_), .A2(
        npu_inst_pe_1_3_6_n1), .B1(npu_inst_pe_1_3_6_N73), .B2(
        npu_inst_pe_1_3_6_n76), .C1(npu_inst_pe_1_3_6_N65), .C2(
        npu_inst_pe_1_3_6_n77), .ZN(npu_inst_pe_1_3_6_n84) );
  INV_X1 npu_inst_pe_1_3_6_U50 ( .A(npu_inst_pe_1_3_6_n84), .ZN(
        npu_inst_pe_1_3_6_n101) );
  AOI222_X1 npu_inst_pe_1_3_6_U49 ( .A1(npu_inst_int_data_res_4__6__7_), .A2(
        npu_inst_pe_1_3_6_n1), .B1(npu_inst_pe_1_3_6_N80), .B2(
        npu_inst_pe_1_3_6_n76), .C1(npu_inst_pe_1_3_6_N72), .C2(
        npu_inst_pe_1_3_6_n77), .ZN(npu_inst_pe_1_3_6_n75) );
  INV_X1 npu_inst_pe_1_3_6_U48 ( .A(npu_inst_pe_1_3_6_n75), .ZN(
        npu_inst_pe_1_3_6_n33) );
  AOI222_X1 npu_inst_pe_1_3_6_U47 ( .A1(npu_inst_int_data_res_4__6__1_), .A2(
        npu_inst_pe_1_3_6_n1), .B1(npu_inst_pe_1_3_6_N74), .B2(
        npu_inst_pe_1_3_6_n76), .C1(npu_inst_pe_1_3_6_N66), .C2(
        npu_inst_pe_1_3_6_n77), .ZN(npu_inst_pe_1_3_6_n83) );
  INV_X1 npu_inst_pe_1_3_6_U46 ( .A(npu_inst_pe_1_3_6_n83), .ZN(
        npu_inst_pe_1_3_6_n100) );
  AOI222_X1 npu_inst_pe_1_3_6_U45 ( .A1(npu_inst_int_data_res_4__6__2_), .A2(
        npu_inst_pe_1_3_6_n1), .B1(npu_inst_pe_1_3_6_N75), .B2(
        npu_inst_pe_1_3_6_n76), .C1(npu_inst_pe_1_3_6_N67), .C2(
        npu_inst_pe_1_3_6_n77), .ZN(npu_inst_pe_1_3_6_n82) );
  INV_X1 npu_inst_pe_1_3_6_U44 ( .A(npu_inst_pe_1_3_6_n82), .ZN(
        npu_inst_pe_1_3_6_n99) );
  AOI222_X1 npu_inst_pe_1_3_6_U43 ( .A1(npu_inst_int_data_res_4__6__3_), .A2(
        npu_inst_pe_1_3_6_n1), .B1(npu_inst_pe_1_3_6_N76), .B2(
        npu_inst_pe_1_3_6_n76), .C1(npu_inst_pe_1_3_6_N68), .C2(
        npu_inst_pe_1_3_6_n77), .ZN(npu_inst_pe_1_3_6_n81) );
  INV_X1 npu_inst_pe_1_3_6_U42 ( .A(npu_inst_pe_1_3_6_n81), .ZN(
        npu_inst_pe_1_3_6_n98) );
  AOI222_X1 npu_inst_pe_1_3_6_U41 ( .A1(npu_inst_int_data_res_4__6__4_), .A2(
        npu_inst_pe_1_3_6_n1), .B1(npu_inst_pe_1_3_6_N77), .B2(
        npu_inst_pe_1_3_6_n76), .C1(npu_inst_pe_1_3_6_N69), .C2(
        npu_inst_pe_1_3_6_n77), .ZN(npu_inst_pe_1_3_6_n80) );
  INV_X1 npu_inst_pe_1_3_6_U40 ( .A(npu_inst_pe_1_3_6_n80), .ZN(
        npu_inst_pe_1_3_6_n36) );
  AOI222_X1 npu_inst_pe_1_3_6_U39 ( .A1(npu_inst_int_data_res_4__6__5_), .A2(
        npu_inst_pe_1_3_6_n1), .B1(npu_inst_pe_1_3_6_N78), .B2(
        npu_inst_pe_1_3_6_n76), .C1(npu_inst_pe_1_3_6_N70), .C2(
        npu_inst_pe_1_3_6_n77), .ZN(npu_inst_pe_1_3_6_n79) );
  INV_X1 npu_inst_pe_1_3_6_U38 ( .A(npu_inst_pe_1_3_6_n79), .ZN(
        npu_inst_pe_1_3_6_n35) );
  AOI222_X1 npu_inst_pe_1_3_6_U37 ( .A1(npu_inst_int_data_res_4__6__6_), .A2(
        npu_inst_pe_1_3_6_n1), .B1(npu_inst_pe_1_3_6_N79), .B2(
        npu_inst_pe_1_3_6_n76), .C1(npu_inst_pe_1_3_6_N71), .C2(
        npu_inst_pe_1_3_6_n77), .ZN(npu_inst_pe_1_3_6_n78) );
  INV_X1 npu_inst_pe_1_3_6_U36 ( .A(npu_inst_pe_1_3_6_n78), .ZN(
        npu_inst_pe_1_3_6_n34) );
  INV_X1 npu_inst_pe_1_3_6_U35 ( .A(npu_inst_pe_1_3_6_int_data_1_), .ZN(
        npu_inst_pe_1_3_6_n14) );
  AND2_X1 npu_inst_pe_1_3_6_U34 ( .A1(npu_inst_int_data_x_3__6__1_), .A2(
        npu_inst_pe_1_3_6_int_q_weight_1_), .ZN(npu_inst_pe_1_3_6_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_3_6_U33 ( .A1(npu_inst_int_data_x_3__6__0_), .A2(
        npu_inst_pe_1_3_6_int_q_weight_1_), .ZN(npu_inst_pe_1_3_6_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_3_6_U32 ( .A1(npu_inst_n56), .A2(
        npu_inst_int_data_y_4__6__1_), .B1(npu_inst_pe_1_3_6_n3), .B2(
        npu_inst_int_data_x_3__7__1_), .ZN(npu_inst_pe_1_3_6_n63) );
  AOI22_X1 npu_inst_pe_1_3_6_U31 ( .A1(npu_inst_n56), .A2(
        npu_inst_int_data_y_4__6__0_), .B1(npu_inst_pe_1_3_6_n3), .B2(
        npu_inst_int_data_x_3__7__0_), .ZN(npu_inst_pe_1_3_6_n61) );
  INV_X1 npu_inst_pe_1_3_6_U30 ( .A(npu_inst_pe_1_3_6_int_data_0_), .ZN(
        npu_inst_pe_1_3_6_n13) );
  INV_X1 npu_inst_pe_1_3_6_U29 ( .A(npu_inst_n69), .ZN(npu_inst_pe_1_3_6_n5)
         );
  OR3_X1 npu_inst_pe_1_3_6_U28 ( .A1(npu_inst_pe_1_3_6_n6), .A2(
        npu_inst_pe_1_3_6_n8), .A3(npu_inst_pe_1_3_6_n5), .ZN(
        npu_inst_pe_1_3_6_n56) );
  OR3_X1 npu_inst_pe_1_3_6_U27 ( .A1(npu_inst_pe_1_3_6_n5), .A2(
        npu_inst_pe_1_3_6_n8), .A3(npu_inst_pe_1_3_6_n7), .ZN(
        npu_inst_pe_1_3_6_n48) );
  INV_X1 npu_inst_pe_1_3_6_U26 ( .A(npu_inst_pe_1_3_6_n5), .ZN(
        npu_inst_pe_1_3_6_n4) );
  OR3_X1 npu_inst_pe_1_3_6_U25 ( .A1(npu_inst_pe_1_3_6_n4), .A2(
        npu_inst_pe_1_3_6_n8), .A3(npu_inst_pe_1_3_6_n7), .ZN(
        npu_inst_pe_1_3_6_n52) );
  OR3_X1 npu_inst_pe_1_3_6_U24 ( .A1(npu_inst_pe_1_3_6_n6), .A2(
        npu_inst_pe_1_3_6_n8), .A3(npu_inst_pe_1_3_6_n4), .ZN(
        npu_inst_pe_1_3_6_n60) );
  NOR2_X1 npu_inst_pe_1_3_6_U23 ( .A1(npu_inst_pe_1_3_6_n60), .A2(
        npu_inst_pe_1_3_6_n3), .ZN(npu_inst_pe_1_3_6_n58) );
  NOR2_X1 npu_inst_pe_1_3_6_U22 ( .A1(npu_inst_pe_1_3_6_n56), .A2(
        npu_inst_pe_1_3_6_n3), .ZN(npu_inst_pe_1_3_6_n54) );
  NOR2_X1 npu_inst_pe_1_3_6_U21 ( .A1(npu_inst_pe_1_3_6_n52), .A2(
        npu_inst_pe_1_3_6_n3), .ZN(npu_inst_pe_1_3_6_n50) );
  NOR2_X1 npu_inst_pe_1_3_6_U20 ( .A1(npu_inst_pe_1_3_6_n48), .A2(
        npu_inst_pe_1_3_6_n3), .ZN(npu_inst_pe_1_3_6_n46) );
  NOR2_X1 npu_inst_pe_1_3_6_U19 ( .A1(npu_inst_pe_1_3_6_n40), .A2(
        npu_inst_pe_1_3_6_n3), .ZN(npu_inst_pe_1_3_6_n38) );
  NOR2_X1 npu_inst_pe_1_3_6_U18 ( .A1(npu_inst_pe_1_3_6_n44), .A2(
        npu_inst_pe_1_3_6_n3), .ZN(npu_inst_pe_1_3_6_n42) );
  BUF_X1 npu_inst_pe_1_3_6_U17 ( .A(npu_inst_n100), .Z(npu_inst_pe_1_3_6_n8)
         );
  INV_X1 npu_inst_pe_1_3_6_U16 ( .A(npu_inst_n124), .ZN(npu_inst_pe_1_3_6_n12)
         );
  INV_X1 npu_inst_pe_1_3_6_U15 ( .A(npu_inst_pe_1_3_6_n38), .ZN(
        npu_inst_pe_1_3_6_n114) );
  INV_X1 npu_inst_pe_1_3_6_U14 ( .A(npu_inst_pe_1_3_6_n58), .ZN(
        npu_inst_pe_1_3_6_n119) );
  INV_X1 npu_inst_pe_1_3_6_U13 ( .A(npu_inst_pe_1_3_6_n54), .ZN(
        npu_inst_pe_1_3_6_n118) );
  INV_X1 npu_inst_pe_1_3_6_U12 ( .A(npu_inst_pe_1_3_6_n50), .ZN(
        npu_inst_pe_1_3_6_n117) );
  INV_X1 npu_inst_pe_1_3_6_U11 ( .A(npu_inst_pe_1_3_6_n46), .ZN(
        npu_inst_pe_1_3_6_n116) );
  INV_X1 npu_inst_pe_1_3_6_U10 ( .A(npu_inst_pe_1_3_6_n42), .ZN(
        npu_inst_pe_1_3_6_n115) );
  BUF_X1 npu_inst_pe_1_3_6_U9 ( .A(npu_inst_n23), .Z(npu_inst_pe_1_3_6_n2) );
  BUF_X1 npu_inst_pe_1_3_6_U8 ( .A(npu_inst_n23), .Z(npu_inst_pe_1_3_6_n1) );
  BUF_X1 npu_inst_pe_1_3_6_U7 ( .A(npu_inst_pe_1_3_6_n12), .Z(
        npu_inst_pe_1_3_6_n11) );
  BUF_X1 npu_inst_pe_1_3_6_U6 ( .A(npu_inst_pe_1_3_6_n12), .Z(
        npu_inst_pe_1_3_6_n10) );
  BUF_X1 npu_inst_pe_1_3_6_U5 ( .A(npu_inst_pe_1_3_6_n12), .Z(
        npu_inst_pe_1_3_6_n9) );
  NOR2_X1 npu_inst_pe_1_3_6_U4 ( .A1(npu_inst_pe_1_3_6_int_q_weight_0_), .A2(
        npu_inst_pe_1_3_6_n1), .ZN(npu_inst_pe_1_3_6_n76) );
  NOR2_X1 npu_inst_pe_1_3_6_U3 ( .A1(npu_inst_pe_1_3_6_n27), .A2(
        npu_inst_pe_1_3_6_n1), .ZN(npu_inst_pe_1_3_6_n77) );
  FA_X1 npu_inst_pe_1_3_6_sub_67_U2_1 ( .A(npu_inst_pe_1_3_6_int_q_acc_1_), 
        .B(npu_inst_pe_1_3_6_n14), .CI(npu_inst_pe_1_3_6_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_3_6_sub_67_carry_2_), .S(npu_inst_pe_1_3_6_N66) );
  FA_X1 npu_inst_pe_1_3_6_add_69_U1_1 ( .A(npu_inst_pe_1_3_6_int_q_acc_1_), 
        .B(npu_inst_pe_1_3_6_int_data_1_), .CI(
        npu_inst_pe_1_3_6_add_69_carry_1_), .CO(
        npu_inst_pe_1_3_6_add_69_carry_2_), .S(npu_inst_pe_1_3_6_N74) );
  NAND3_X1 npu_inst_pe_1_3_6_U109 ( .A1(npu_inst_pe_1_3_6_n5), .A2(
        npu_inst_pe_1_3_6_n7), .A3(npu_inst_pe_1_3_6_n8), .ZN(
        npu_inst_pe_1_3_6_n44) );
  NAND3_X1 npu_inst_pe_1_3_6_U108 ( .A1(npu_inst_pe_1_3_6_n4), .A2(
        npu_inst_pe_1_3_6_n7), .A3(npu_inst_pe_1_3_6_n8), .ZN(
        npu_inst_pe_1_3_6_n40) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_3_6_n34), .CK(
        npu_inst_pe_1_3_6_net3872), .RN(npu_inst_pe_1_3_6_n9), .Q(
        npu_inst_pe_1_3_6_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_3_6_n35), .CK(
        npu_inst_pe_1_3_6_net3872), .RN(npu_inst_pe_1_3_6_n9), .Q(
        npu_inst_pe_1_3_6_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_3_6_n36), .CK(
        npu_inst_pe_1_3_6_net3872), .RN(npu_inst_pe_1_3_6_n9), .Q(
        npu_inst_pe_1_3_6_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_3_6_n98), .CK(
        npu_inst_pe_1_3_6_net3872), .RN(npu_inst_pe_1_3_6_n9), .Q(
        npu_inst_pe_1_3_6_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_3_6_n99), .CK(
        npu_inst_pe_1_3_6_net3872), .RN(npu_inst_pe_1_3_6_n9), .Q(
        npu_inst_pe_1_3_6_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_3_6_n100), 
        .CK(npu_inst_pe_1_3_6_net3872), .RN(npu_inst_pe_1_3_6_n9), .Q(
        npu_inst_pe_1_3_6_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_3_6_n33), .CK(
        npu_inst_pe_1_3_6_net3872), .RN(npu_inst_pe_1_3_6_n9), .Q(
        npu_inst_pe_1_3_6_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_3_6_n101), 
        .CK(npu_inst_pe_1_3_6_net3872), .RN(npu_inst_pe_1_3_6_n9), .Q(
        npu_inst_pe_1_3_6_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_weight_reg_0_ ( .D(npu_inst_n110), .CK(
        npu_inst_pe_1_3_6_net3878), .RN(npu_inst_pe_1_3_6_n9), .Q(
        npu_inst_pe_1_3_6_int_q_weight_0_), .QN(npu_inst_pe_1_3_6_n27) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_weight_reg_1_ ( .D(npu_inst_n116), .CK(
        npu_inst_pe_1_3_6_net3878), .RN(npu_inst_pe_1_3_6_n9), .Q(
        npu_inst_pe_1_3_6_int_q_weight_1_), .QN(npu_inst_pe_1_3_6_n26) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_3_6_n113), 
        .CK(npu_inst_pe_1_3_6_net3878), .RN(npu_inst_pe_1_3_6_n9), .Q(
        npu_inst_pe_1_3_6_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_3_6_n107), 
        .CK(npu_inst_pe_1_3_6_net3878), .RN(npu_inst_pe_1_3_6_n9), .Q(
        npu_inst_pe_1_3_6_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_3_6_n112), 
        .CK(npu_inst_pe_1_3_6_net3878), .RN(npu_inst_pe_1_3_6_n10), .Q(
        npu_inst_pe_1_3_6_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_3_6_n106), 
        .CK(npu_inst_pe_1_3_6_net3878), .RN(npu_inst_pe_1_3_6_n10), .Q(
        npu_inst_pe_1_3_6_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_3_6_n111), 
        .CK(npu_inst_pe_1_3_6_net3878), .RN(npu_inst_pe_1_3_6_n10), .Q(
        npu_inst_pe_1_3_6_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_3_6_n105), 
        .CK(npu_inst_pe_1_3_6_net3878), .RN(npu_inst_pe_1_3_6_n10), .Q(
        npu_inst_pe_1_3_6_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_3_6_n110), 
        .CK(npu_inst_pe_1_3_6_net3878), .RN(npu_inst_pe_1_3_6_n10), .Q(
        npu_inst_pe_1_3_6_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_3_6_n104), 
        .CK(npu_inst_pe_1_3_6_net3878), .RN(npu_inst_pe_1_3_6_n10), .Q(
        npu_inst_pe_1_3_6_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_3_6_n109), 
        .CK(npu_inst_pe_1_3_6_net3878), .RN(npu_inst_pe_1_3_6_n10), .Q(
        npu_inst_pe_1_3_6_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_3_6_n103), 
        .CK(npu_inst_pe_1_3_6_net3878), .RN(npu_inst_pe_1_3_6_n10), .Q(
        npu_inst_pe_1_3_6_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_3_6_n108), 
        .CK(npu_inst_pe_1_3_6_net3878), .RN(npu_inst_pe_1_3_6_n10), .Q(
        npu_inst_pe_1_3_6_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_3_6_n102), 
        .CK(npu_inst_pe_1_3_6_net3878), .RN(npu_inst_pe_1_3_6_n10), .Q(
        npu_inst_pe_1_3_6_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_3_6_n86), 
        .CK(npu_inst_pe_1_3_6_net3878), .RN(npu_inst_pe_1_3_6_n10), .Q(
        npu_inst_pe_1_3_6_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_3_6_n87), 
        .CK(npu_inst_pe_1_3_6_net3878), .RN(npu_inst_pe_1_3_6_n10), .Q(
        npu_inst_pe_1_3_6_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_3_6_n88), 
        .CK(npu_inst_pe_1_3_6_net3878), .RN(npu_inst_pe_1_3_6_n11), .Q(
        npu_inst_pe_1_3_6_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_3_6_n89), 
        .CK(npu_inst_pe_1_3_6_net3878), .RN(npu_inst_pe_1_3_6_n11), .Q(
        npu_inst_pe_1_3_6_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_3_6_n90), 
        .CK(npu_inst_pe_1_3_6_net3878), .RN(npu_inst_pe_1_3_6_n11), .Q(
        npu_inst_pe_1_3_6_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_3_6_n91), 
        .CK(npu_inst_pe_1_3_6_net3878), .RN(npu_inst_pe_1_3_6_n11), .Q(
        npu_inst_pe_1_3_6_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_3_6_n92), 
        .CK(npu_inst_pe_1_3_6_net3878), .RN(npu_inst_pe_1_3_6_n11), .Q(
        npu_inst_pe_1_3_6_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_3_6_n93), 
        .CK(npu_inst_pe_1_3_6_net3878), .RN(npu_inst_pe_1_3_6_n11), .Q(
        npu_inst_pe_1_3_6_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_3_6_n94), 
        .CK(npu_inst_pe_1_3_6_net3878), .RN(npu_inst_pe_1_3_6_n11), .Q(
        npu_inst_pe_1_3_6_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_3_6_n95), 
        .CK(npu_inst_pe_1_3_6_net3878), .RN(npu_inst_pe_1_3_6_n11), .Q(
        npu_inst_pe_1_3_6_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_3_6_n96), 
        .CK(npu_inst_pe_1_3_6_net3878), .RN(npu_inst_pe_1_3_6_n11), .Q(
        npu_inst_pe_1_3_6_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_3_6_n97), 
        .CK(npu_inst_pe_1_3_6_net3878), .RN(npu_inst_pe_1_3_6_n11), .Q(
        npu_inst_pe_1_3_6_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_3_6_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_3_6_N84), .SE(1'b0), .GCK(npu_inst_pe_1_3_6_net3872) );
  CLKGATETST_X1 npu_inst_pe_1_3_6_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n64), .SE(1'b0), .GCK(npu_inst_pe_1_3_6_net3878) );
  MUX2_X1 npu_inst_pe_1_3_7_U162 ( .A(npu_inst_pe_1_3_7_n32), .B(
        npu_inst_pe_1_3_7_n29), .S(npu_inst_pe_1_3_7_n8), .Z(
        npu_inst_pe_1_3_7_N93) );
  MUX2_X1 npu_inst_pe_1_3_7_U161 ( .A(npu_inst_pe_1_3_7_n31), .B(
        npu_inst_pe_1_3_7_n30), .S(npu_inst_pe_1_3_7_n6), .Z(
        npu_inst_pe_1_3_7_n32) );
  MUX2_X1 npu_inst_pe_1_3_7_U160 ( .A(npu_inst_pe_1_3_7_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_3_7_int_q_reg_v_1__0_), .S(npu_inst_pe_1_3_7_n4), .Z(
        npu_inst_pe_1_3_7_n31) );
  MUX2_X1 npu_inst_pe_1_3_7_U159 ( .A(npu_inst_pe_1_3_7_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_3_7_int_q_reg_v_3__0_), .S(npu_inst_pe_1_3_7_n4), .Z(
        npu_inst_pe_1_3_7_n30) );
  MUX2_X1 npu_inst_pe_1_3_7_U158 ( .A(npu_inst_pe_1_3_7_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_3_7_int_q_reg_v_5__0_), .S(npu_inst_pe_1_3_7_n4), .Z(
        npu_inst_pe_1_3_7_n29) );
  MUX2_X1 npu_inst_pe_1_3_7_U157 ( .A(npu_inst_pe_1_3_7_n28), .B(
        npu_inst_pe_1_3_7_n23), .S(npu_inst_pe_1_3_7_n8), .Z(
        npu_inst_pe_1_3_7_N94) );
  MUX2_X1 npu_inst_pe_1_3_7_U156 ( .A(npu_inst_pe_1_3_7_n25), .B(
        npu_inst_pe_1_3_7_n24), .S(npu_inst_pe_1_3_7_n6), .Z(
        npu_inst_pe_1_3_7_n28) );
  MUX2_X1 npu_inst_pe_1_3_7_U155 ( .A(npu_inst_pe_1_3_7_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_3_7_int_q_reg_v_1__1_), .S(npu_inst_pe_1_3_7_n4), .Z(
        npu_inst_pe_1_3_7_n25) );
  MUX2_X1 npu_inst_pe_1_3_7_U154 ( .A(npu_inst_pe_1_3_7_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_3_7_int_q_reg_v_3__1_), .S(npu_inst_pe_1_3_7_n4), .Z(
        npu_inst_pe_1_3_7_n24) );
  MUX2_X1 npu_inst_pe_1_3_7_U153 ( .A(npu_inst_pe_1_3_7_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_3_7_int_q_reg_v_5__1_), .S(npu_inst_pe_1_3_7_n4), .Z(
        npu_inst_pe_1_3_7_n23) );
  MUX2_X1 npu_inst_pe_1_3_7_U152 ( .A(npu_inst_pe_1_3_7_n22), .B(
        npu_inst_pe_1_3_7_n19), .S(npu_inst_pe_1_3_7_n8), .Z(
        npu_inst_int_data_x_3__7__1_) );
  MUX2_X1 npu_inst_pe_1_3_7_U151 ( .A(npu_inst_pe_1_3_7_n21), .B(
        npu_inst_pe_1_3_7_n20), .S(npu_inst_pe_1_3_7_n6), .Z(
        npu_inst_pe_1_3_7_n22) );
  MUX2_X1 npu_inst_pe_1_3_7_U150 ( .A(npu_inst_pe_1_3_7_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_3_7_int_q_reg_h_1__1_), .S(npu_inst_pe_1_3_7_n4), .Z(
        npu_inst_pe_1_3_7_n21) );
  MUX2_X1 npu_inst_pe_1_3_7_U149 ( .A(npu_inst_pe_1_3_7_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_3_7_int_q_reg_h_3__1_), .S(npu_inst_pe_1_3_7_n4), .Z(
        npu_inst_pe_1_3_7_n20) );
  MUX2_X1 npu_inst_pe_1_3_7_U148 ( .A(npu_inst_pe_1_3_7_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_3_7_int_q_reg_h_5__1_), .S(npu_inst_pe_1_3_7_n4), .Z(
        npu_inst_pe_1_3_7_n19) );
  MUX2_X1 npu_inst_pe_1_3_7_U147 ( .A(npu_inst_pe_1_3_7_n18), .B(
        npu_inst_pe_1_3_7_n15), .S(npu_inst_pe_1_3_7_n8), .Z(
        npu_inst_int_data_x_3__7__0_) );
  MUX2_X1 npu_inst_pe_1_3_7_U146 ( .A(npu_inst_pe_1_3_7_n17), .B(
        npu_inst_pe_1_3_7_n16), .S(npu_inst_pe_1_3_7_n6), .Z(
        npu_inst_pe_1_3_7_n18) );
  MUX2_X1 npu_inst_pe_1_3_7_U145 ( .A(npu_inst_pe_1_3_7_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_3_7_int_q_reg_h_1__0_), .S(npu_inst_pe_1_3_7_n4), .Z(
        npu_inst_pe_1_3_7_n17) );
  MUX2_X1 npu_inst_pe_1_3_7_U144 ( .A(npu_inst_pe_1_3_7_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_3_7_int_q_reg_h_3__0_), .S(npu_inst_pe_1_3_7_n4), .Z(
        npu_inst_pe_1_3_7_n16) );
  MUX2_X1 npu_inst_pe_1_3_7_U143 ( .A(npu_inst_pe_1_3_7_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_3_7_int_q_reg_h_5__0_), .S(npu_inst_pe_1_3_7_n4), .Z(
        npu_inst_pe_1_3_7_n15) );
  XOR2_X1 npu_inst_pe_1_3_7_U142 ( .A(npu_inst_pe_1_3_7_int_data_0_), .B(
        npu_inst_pe_1_3_7_int_q_acc_0_), .Z(npu_inst_pe_1_3_7_N73) );
  AND2_X1 npu_inst_pe_1_3_7_U141 ( .A1(npu_inst_pe_1_3_7_int_q_acc_0_), .A2(
        npu_inst_pe_1_3_7_int_data_0_), .ZN(npu_inst_pe_1_3_7_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_3_7_U140 ( .A(npu_inst_pe_1_3_7_int_q_acc_0_), .B(
        npu_inst_pe_1_3_7_n13), .ZN(npu_inst_pe_1_3_7_N65) );
  OR2_X1 npu_inst_pe_1_3_7_U139 ( .A1(npu_inst_pe_1_3_7_n13), .A2(
        npu_inst_pe_1_3_7_int_q_acc_0_), .ZN(npu_inst_pe_1_3_7_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_3_7_U138 ( .A(npu_inst_pe_1_3_7_int_q_acc_2_), .B(
        npu_inst_pe_1_3_7_add_69_carry_2_), .Z(npu_inst_pe_1_3_7_N75) );
  AND2_X1 npu_inst_pe_1_3_7_U137 ( .A1(npu_inst_pe_1_3_7_add_69_carry_2_), 
        .A2(npu_inst_pe_1_3_7_int_q_acc_2_), .ZN(
        npu_inst_pe_1_3_7_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_3_7_U136 ( .A(npu_inst_pe_1_3_7_int_q_acc_3_), .B(
        npu_inst_pe_1_3_7_add_69_carry_3_), .Z(npu_inst_pe_1_3_7_N76) );
  AND2_X1 npu_inst_pe_1_3_7_U135 ( .A1(npu_inst_pe_1_3_7_add_69_carry_3_), 
        .A2(npu_inst_pe_1_3_7_int_q_acc_3_), .ZN(
        npu_inst_pe_1_3_7_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_3_7_U134 ( .A(npu_inst_pe_1_3_7_int_q_acc_4_), .B(
        npu_inst_pe_1_3_7_add_69_carry_4_), .Z(npu_inst_pe_1_3_7_N77) );
  AND2_X1 npu_inst_pe_1_3_7_U133 ( .A1(npu_inst_pe_1_3_7_add_69_carry_4_), 
        .A2(npu_inst_pe_1_3_7_int_q_acc_4_), .ZN(
        npu_inst_pe_1_3_7_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_3_7_U132 ( .A(npu_inst_pe_1_3_7_int_q_acc_5_), .B(
        npu_inst_pe_1_3_7_add_69_carry_5_), .Z(npu_inst_pe_1_3_7_N78) );
  AND2_X1 npu_inst_pe_1_3_7_U131 ( .A1(npu_inst_pe_1_3_7_add_69_carry_5_), 
        .A2(npu_inst_pe_1_3_7_int_q_acc_5_), .ZN(
        npu_inst_pe_1_3_7_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_3_7_U130 ( .A(npu_inst_pe_1_3_7_int_q_acc_6_), .B(
        npu_inst_pe_1_3_7_add_69_carry_6_), .Z(npu_inst_pe_1_3_7_N79) );
  AND2_X1 npu_inst_pe_1_3_7_U129 ( .A1(npu_inst_pe_1_3_7_add_69_carry_6_), 
        .A2(npu_inst_pe_1_3_7_int_q_acc_6_), .ZN(
        npu_inst_pe_1_3_7_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_3_7_U128 ( .A(npu_inst_pe_1_3_7_int_q_acc_7_), .B(
        npu_inst_pe_1_3_7_add_69_carry_7_), .Z(npu_inst_pe_1_3_7_N80) );
  XNOR2_X1 npu_inst_pe_1_3_7_U127 ( .A(npu_inst_pe_1_3_7_sub_67_carry_2_), .B(
        npu_inst_pe_1_3_7_int_q_acc_2_), .ZN(npu_inst_pe_1_3_7_N67) );
  OR2_X1 npu_inst_pe_1_3_7_U126 ( .A1(npu_inst_pe_1_3_7_int_q_acc_2_), .A2(
        npu_inst_pe_1_3_7_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_3_7_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_3_7_U125 ( .A(npu_inst_pe_1_3_7_sub_67_carry_3_), .B(
        npu_inst_pe_1_3_7_int_q_acc_3_), .ZN(npu_inst_pe_1_3_7_N68) );
  OR2_X1 npu_inst_pe_1_3_7_U124 ( .A1(npu_inst_pe_1_3_7_int_q_acc_3_), .A2(
        npu_inst_pe_1_3_7_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_3_7_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_3_7_U123 ( .A(npu_inst_pe_1_3_7_sub_67_carry_4_), .B(
        npu_inst_pe_1_3_7_int_q_acc_4_), .ZN(npu_inst_pe_1_3_7_N69) );
  OR2_X1 npu_inst_pe_1_3_7_U122 ( .A1(npu_inst_pe_1_3_7_int_q_acc_4_), .A2(
        npu_inst_pe_1_3_7_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_3_7_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_3_7_U121 ( .A(npu_inst_pe_1_3_7_sub_67_carry_5_), .B(
        npu_inst_pe_1_3_7_int_q_acc_5_), .ZN(npu_inst_pe_1_3_7_N70) );
  OR2_X1 npu_inst_pe_1_3_7_U120 ( .A1(npu_inst_pe_1_3_7_int_q_acc_5_), .A2(
        npu_inst_pe_1_3_7_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_3_7_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_3_7_U119 ( .A(npu_inst_pe_1_3_7_sub_67_carry_6_), .B(
        npu_inst_pe_1_3_7_int_q_acc_6_), .ZN(npu_inst_pe_1_3_7_N71) );
  OR2_X1 npu_inst_pe_1_3_7_U118 ( .A1(npu_inst_pe_1_3_7_int_q_acc_6_), .A2(
        npu_inst_pe_1_3_7_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_3_7_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_3_7_U117 ( .A(npu_inst_pe_1_3_7_int_q_acc_7_), .B(
        npu_inst_pe_1_3_7_sub_67_carry_7_), .ZN(npu_inst_pe_1_3_7_N72) );
  INV_X1 npu_inst_pe_1_3_7_U116 ( .A(npu_inst_n77), .ZN(npu_inst_pe_1_3_7_n7)
         );
  INV_X1 npu_inst_pe_1_3_7_U115 ( .A(npu_inst_pe_1_3_7_n7), .ZN(
        npu_inst_pe_1_3_7_n6) );
  INV_X1 npu_inst_pe_1_3_7_U114 ( .A(npu_inst_n56), .ZN(npu_inst_pe_1_3_7_n3)
         );
  AOI22_X1 npu_inst_pe_1_3_7_U113 ( .A1(npu_inst_int_data_y_4__7__0_), .A2(
        npu_inst_pe_1_3_7_n58), .B1(npu_inst_pe_1_3_7_n119), .B2(
        npu_inst_pe_1_3_7_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_3_7_n57) );
  INV_X1 npu_inst_pe_1_3_7_U112 ( .A(npu_inst_pe_1_3_7_n57), .ZN(
        npu_inst_pe_1_3_7_n108) );
  AOI22_X1 npu_inst_pe_1_3_7_U111 ( .A1(npu_inst_int_data_y_4__7__0_), .A2(
        npu_inst_pe_1_3_7_n54), .B1(npu_inst_pe_1_3_7_n118), .B2(
        npu_inst_pe_1_3_7_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_3_7_n53) );
  INV_X1 npu_inst_pe_1_3_7_U110 ( .A(npu_inst_pe_1_3_7_n53), .ZN(
        npu_inst_pe_1_3_7_n109) );
  AOI22_X1 npu_inst_pe_1_3_7_U107 ( .A1(npu_inst_int_data_y_4__7__0_), .A2(
        npu_inst_pe_1_3_7_n50), .B1(npu_inst_pe_1_3_7_n117), .B2(
        npu_inst_pe_1_3_7_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_3_7_n49) );
  INV_X1 npu_inst_pe_1_3_7_U106 ( .A(npu_inst_pe_1_3_7_n49), .ZN(
        npu_inst_pe_1_3_7_n110) );
  AOI22_X1 npu_inst_pe_1_3_7_U105 ( .A1(npu_inst_int_data_y_4__7__0_), .A2(
        npu_inst_pe_1_3_7_n46), .B1(npu_inst_pe_1_3_7_n116), .B2(
        npu_inst_pe_1_3_7_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_3_7_n45) );
  INV_X1 npu_inst_pe_1_3_7_U104 ( .A(npu_inst_pe_1_3_7_n45), .ZN(
        npu_inst_pe_1_3_7_n111) );
  AOI22_X1 npu_inst_pe_1_3_7_U103 ( .A1(npu_inst_int_data_y_4__7__0_), .A2(
        npu_inst_pe_1_3_7_n42), .B1(npu_inst_pe_1_3_7_n115), .B2(
        npu_inst_pe_1_3_7_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_3_7_n41) );
  INV_X1 npu_inst_pe_1_3_7_U102 ( .A(npu_inst_pe_1_3_7_n41), .ZN(
        npu_inst_pe_1_3_7_n112) );
  AOI22_X1 npu_inst_pe_1_3_7_U101 ( .A1(npu_inst_int_data_y_4__7__1_), .A2(
        npu_inst_pe_1_3_7_n58), .B1(npu_inst_pe_1_3_7_n119), .B2(
        npu_inst_pe_1_3_7_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_3_7_n59) );
  INV_X1 npu_inst_pe_1_3_7_U100 ( .A(npu_inst_pe_1_3_7_n59), .ZN(
        npu_inst_pe_1_3_7_n102) );
  AOI22_X1 npu_inst_pe_1_3_7_U99 ( .A1(npu_inst_int_data_y_4__7__1_), .A2(
        npu_inst_pe_1_3_7_n54), .B1(npu_inst_pe_1_3_7_n118), .B2(
        npu_inst_pe_1_3_7_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_3_7_n55) );
  INV_X1 npu_inst_pe_1_3_7_U98 ( .A(npu_inst_pe_1_3_7_n55), .ZN(
        npu_inst_pe_1_3_7_n103) );
  AOI22_X1 npu_inst_pe_1_3_7_U97 ( .A1(npu_inst_int_data_y_4__7__1_), .A2(
        npu_inst_pe_1_3_7_n50), .B1(npu_inst_pe_1_3_7_n117), .B2(
        npu_inst_pe_1_3_7_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_3_7_n51) );
  INV_X1 npu_inst_pe_1_3_7_U96 ( .A(npu_inst_pe_1_3_7_n51), .ZN(
        npu_inst_pe_1_3_7_n104) );
  AOI22_X1 npu_inst_pe_1_3_7_U95 ( .A1(npu_inst_int_data_y_4__7__1_), .A2(
        npu_inst_pe_1_3_7_n46), .B1(npu_inst_pe_1_3_7_n116), .B2(
        npu_inst_pe_1_3_7_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_3_7_n47) );
  INV_X1 npu_inst_pe_1_3_7_U94 ( .A(npu_inst_pe_1_3_7_n47), .ZN(
        npu_inst_pe_1_3_7_n105) );
  AOI22_X1 npu_inst_pe_1_3_7_U93 ( .A1(npu_inst_int_data_y_4__7__1_), .A2(
        npu_inst_pe_1_3_7_n42), .B1(npu_inst_pe_1_3_7_n115), .B2(
        npu_inst_pe_1_3_7_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_3_7_n43) );
  INV_X1 npu_inst_pe_1_3_7_U92 ( .A(npu_inst_pe_1_3_7_n43), .ZN(
        npu_inst_pe_1_3_7_n106) );
  AOI22_X1 npu_inst_pe_1_3_7_U91 ( .A1(npu_inst_pe_1_3_7_n38), .A2(
        npu_inst_int_data_y_4__7__1_), .B1(npu_inst_pe_1_3_7_n114), .B2(
        npu_inst_pe_1_3_7_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_3_7_n39) );
  INV_X1 npu_inst_pe_1_3_7_U90 ( .A(npu_inst_pe_1_3_7_n39), .ZN(
        npu_inst_pe_1_3_7_n107) );
  AOI22_X1 npu_inst_pe_1_3_7_U89 ( .A1(npu_inst_pe_1_3_7_n38), .A2(
        npu_inst_int_data_y_4__7__0_), .B1(npu_inst_pe_1_3_7_n114), .B2(
        npu_inst_pe_1_3_7_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_3_7_n37) );
  INV_X1 npu_inst_pe_1_3_7_U88 ( .A(npu_inst_pe_1_3_7_n37), .ZN(
        npu_inst_pe_1_3_7_n113) );
  AND2_X1 npu_inst_pe_1_3_7_U87 ( .A1(npu_inst_pe_1_3_7_N93), .A2(npu_inst_n56), .ZN(npu_inst_int_data_y_3__7__0_) );
  AND2_X1 npu_inst_pe_1_3_7_U86 ( .A1(npu_inst_n56), .A2(npu_inst_pe_1_3_7_N94), .ZN(npu_inst_int_data_y_3__7__1_) );
  NOR3_X1 npu_inst_pe_1_3_7_U85 ( .A1(npu_inst_pe_1_3_7_n26), .A2(npu_inst_n56), .A3(npu_inst_int_ckg[32]), .ZN(npu_inst_pe_1_3_7_n85) );
  OR2_X1 npu_inst_pe_1_3_7_U84 ( .A1(npu_inst_pe_1_3_7_n85), .A2(
        npu_inst_pe_1_3_7_n2), .ZN(npu_inst_pe_1_3_7_N84) );
  AND2_X1 npu_inst_pe_1_3_7_U83 ( .A1(npu_inst_pe_1_3_7_int_q_acc_0_), .A2(
        npu_inst_pe_1_3_7_n1), .ZN(npu_inst_int_data_res_3__7__0_) );
  AND2_X1 npu_inst_pe_1_3_7_U82 ( .A1(npu_inst_pe_1_3_7_n2), .A2(
        npu_inst_pe_1_3_7_int_q_acc_7_), .ZN(npu_inst_int_data_res_3__7__7_)
         );
  AND2_X1 npu_inst_pe_1_3_7_U81 ( .A1(npu_inst_pe_1_3_7_int_q_acc_1_), .A2(
        npu_inst_pe_1_3_7_n1), .ZN(npu_inst_int_data_res_3__7__1_) );
  AND2_X1 npu_inst_pe_1_3_7_U80 ( .A1(npu_inst_pe_1_3_7_int_q_acc_2_), .A2(
        npu_inst_pe_1_3_7_n1), .ZN(npu_inst_int_data_res_3__7__2_) );
  AND2_X1 npu_inst_pe_1_3_7_U79 ( .A1(npu_inst_pe_1_3_7_int_q_acc_3_), .A2(
        npu_inst_pe_1_3_7_n2), .ZN(npu_inst_int_data_res_3__7__3_) );
  AND2_X1 npu_inst_pe_1_3_7_U78 ( .A1(npu_inst_pe_1_3_7_int_q_acc_4_), .A2(
        npu_inst_pe_1_3_7_n2), .ZN(npu_inst_int_data_res_3__7__4_) );
  AND2_X1 npu_inst_pe_1_3_7_U77 ( .A1(npu_inst_pe_1_3_7_int_q_acc_5_), .A2(
        npu_inst_pe_1_3_7_n2), .ZN(npu_inst_int_data_res_3__7__5_) );
  AND2_X1 npu_inst_pe_1_3_7_U76 ( .A1(npu_inst_pe_1_3_7_int_q_acc_6_), .A2(
        npu_inst_pe_1_3_7_n2), .ZN(npu_inst_int_data_res_3__7__6_) );
  AOI222_X1 npu_inst_pe_1_3_7_U75 ( .A1(npu_inst_int_data_res_4__7__0_), .A2(
        npu_inst_pe_1_3_7_n1), .B1(npu_inst_pe_1_3_7_N73), .B2(
        npu_inst_pe_1_3_7_n76), .C1(npu_inst_pe_1_3_7_N65), .C2(
        npu_inst_pe_1_3_7_n77), .ZN(npu_inst_pe_1_3_7_n84) );
  INV_X1 npu_inst_pe_1_3_7_U74 ( .A(npu_inst_pe_1_3_7_n84), .ZN(
        npu_inst_pe_1_3_7_n101) );
  AOI222_X1 npu_inst_pe_1_3_7_U73 ( .A1(npu_inst_int_data_res_4__7__7_), .A2(
        npu_inst_pe_1_3_7_n1), .B1(npu_inst_pe_1_3_7_N80), .B2(
        npu_inst_pe_1_3_7_n76), .C1(npu_inst_pe_1_3_7_N72), .C2(
        npu_inst_pe_1_3_7_n77), .ZN(npu_inst_pe_1_3_7_n75) );
  INV_X1 npu_inst_pe_1_3_7_U72 ( .A(npu_inst_pe_1_3_7_n75), .ZN(
        npu_inst_pe_1_3_7_n33) );
  AOI222_X1 npu_inst_pe_1_3_7_U71 ( .A1(npu_inst_int_data_res_4__7__1_), .A2(
        npu_inst_pe_1_3_7_n1), .B1(npu_inst_pe_1_3_7_N74), .B2(
        npu_inst_pe_1_3_7_n76), .C1(npu_inst_pe_1_3_7_N66), .C2(
        npu_inst_pe_1_3_7_n77), .ZN(npu_inst_pe_1_3_7_n83) );
  INV_X1 npu_inst_pe_1_3_7_U70 ( .A(npu_inst_pe_1_3_7_n83), .ZN(
        npu_inst_pe_1_3_7_n100) );
  AOI222_X1 npu_inst_pe_1_3_7_U69 ( .A1(npu_inst_int_data_res_4__7__2_), .A2(
        npu_inst_pe_1_3_7_n1), .B1(npu_inst_pe_1_3_7_N75), .B2(
        npu_inst_pe_1_3_7_n76), .C1(npu_inst_pe_1_3_7_N67), .C2(
        npu_inst_pe_1_3_7_n77), .ZN(npu_inst_pe_1_3_7_n82) );
  INV_X1 npu_inst_pe_1_3_7_U68 ( .A(npu_inst_pe_1_3_7_n82), .ZN(
        npu_inst_pe_1_3_7_n99) );
  AOI222_X1 npu_inst_pe_1_3_7_U67 ( .A1(npu_inst_int_data_res_4__7__3_), .A2(
        npu_inst_pe_1_3_7_n1), .B1(npu_inst_pe_1_3_7_N76), .B2(
        npu_inst_pe_1_3_7_n76), .C1(npu_inst_pe_1_3_7_N68), .C2(
        npu_inst_pe_1_3_7_n77), .ZN(npu_inst_pe_1_3_7_n81) );
  INV_X1 npu_inst_pe_1_3_7_U66 ( .A(npu_inst_pe_1_3_7_n81), .ZN(
        npu_inst_pe_1_3_7_n98) );
  AOI222_X1 npu_inst_pe_1_3_7_U65 ( .A1(npu_inst_int_data_res_4__7__4_), .A2(
        npu_inst_pe_1_3_7_n1), .B1(npu_inst_pe_1_3_7_N77), .B2(
        npu_inst_pe_1_3_7_n76), .C1(npu_inst_pe_1_3_7_N69), .C2(
        npu_inst_pe_1_3_7_n77), .ZN(npu_inst_pe_1_3_7_n80) );
  INV_X1 npu_inst_pe_1_3_7_U64 ( .A(npu_inst_pe_1_3_7_n80), .ZN(
        npu_inst_pe_1_3_7_n36) );
  AOI222_X1 npu_inst_pe_1_3_7_U63 ( .A1(npu_inst_int_data_res_4__7__5_), .A2(
        npu_inst_pe_1_3_7_n1), .B1(npu_inst_pe_1_3_7_N78), .B2(
        npu_inst_pe_1_3_7_n76), .C1(npu_inst_pe_1_3_7_N70), .C2(
        npu_inst_pe_1_3_7_n77), .ZN(npu_inst_pe_1_3_7_n79) );
  INV_X1 npu_inst_pe_1_3_7_U62 ( .A(npu_inst_pe_1_3_7_n79), .ZN(
        npu_inst_pe_1_3_7_n35) );
  AOI222_X1 npu_inst_pe_1_3_7_U61 ( .A1(npu_inst_int_data_res_4__7__6_), .A2(
        npu_inst_pe_1_3_7_n1), .B1(npu_inst_pe_1_3_7_N79), .B2(
        npu_inst_pe_1_3_7_n76), .C1(npu_inst_pe_1_3_7_N71), .C2(
        npu_inst_pe_1_3_7_n77), .ZN(npu_inst_pe_1_3_7_n78) );
  INV_X1 npu_inst_pe_1_3_7_U60 ( .A(npu_inst_pe_1_3_7_n78), .ZN(
        npu_inst_pe_1_3_7_n34) );
  INV_X1 npu_inst_pe_1_3_7_U59 ( .A(npu_inst_pe_1_3_7_int_data_1_), .ZN(
        npu_inst_pe_1_3_7_n14) );
  AND2_X1 npu_inst_pe_1_3_7_U58 ( .A1(npu_inst_int_data_x_3__7__1_), .A2(
        npu_inst_pe_1_3_7_int_q_weight_1_), .ZN(npu_inst_pe_1_3_7_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_3_7_U57 ( .A1(npu_inst_int_data_x_3__7__0_), .A2(
        npu_inst_pe_1_3_7_int_q_weight_1_), .ZN(npu_inst_pe_1_3_7_int_data_0_)
         );
  NAND2_X1 npu_inst_pe_1_3_7_U56 ( .A1(npu_inst_pe_1_3_7_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_3_7_n60), .ZN(npu_inst_pe_1_3_7_n74) );
  OAI21_X1 npu_inst_pe_1_3_7_U55 ( .B1(npu_inst_pe_1_3_7_n63), .B2(
        npu_inst_pe_1_3_7_n60), .A(npu_inst_pe_1_3_7_n74), .ZN(
        npu_inst_pe_1_3_7_n97) );
  NAND2_X1 npu_inst_pe_1_3_7_U54 ( .A1(npu_inst_pe_1_3_7_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_3_7_n60), .ZN(npu_inst_pe_1_3_7_n73) );
  OAI21_X1 npu_inst_pe_1_3_7_U53 ( .B1(npu_inst_pe_1_3_7_n61), .B2(
        npu_inst_pe_1_3_7_n60), .A(npu_inst_pe_1_3_7_n73), .ZN(
        npu_inst_pe_1_3_7_n96) );
  NAND2_X1 npu_inst_pe_1_3_7_U52 ( .A1(npu_inst_pe_1_3_7_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_3_7_n56), .ZN(npu_inst_pe_1_3_7_n72) );
  OAI21_X1 npu_inst_pe_1_3_7_U51 ( .B1(npu_inst_pe_1_3_7_n63), .B2(
        npu_inst_pe_1_3_7_n56), .A(npu_inst_pe_1_3_7_n72), .ZN(
        npu_inst_pe_1_3_7_n95) );
  NAND2_X1 npu_inst_pe_1_3_7_U50 ( .A1(npu_inst_pe_1_3_7_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_3_7_n56), .ZN(npu_inst_pe_1_3_7_n71) );
  OAI21_X1 npu_inst_pe_1_3_7_U49 ( .B1(npu_inst_pe_1_3_7_n61), .B2(
        npu_inst_pe_1_3_7_n56), .A(npu_inst_pe_1_3_7_n71), .ZN(
        npu_inst_pe_1_3_7_n94) );
  NAND2_X1 npu_inst_pe_1_3_7_U48 ( .A1(npu_inst_pe_1_3_7_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_3_7_n52), .ZN(npu_inst_pe_1_3_7_n70) );
  OAI21_X1 npu_inst_pe_1_3_7_U47 ( .B1(npu_inst_pe_1_3_7_n63), .B2(
        npu_inst_pe_1_3_7_n52), .A(npu_inst_pe_1_3_7_n70), .ZN(
        npu_inst_pe_1_3_7_n93) );
  NAND2_X1 npu_inst_pe_1_3_7_U46 ( .A1(npu_inst_pe_1_3_7_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_3_7_n52), .ZN(npu_inst_pe_1_3_7_n69) );
  OAI21_X1 npu_inst_pe_1_3_7_U45 ( .B1(npu_inst_pe_1_3_7_n61), .B2(
        npu_inst_pe_1_3_7_n52), .A(npu_inst_pe_1_3_7_n69), .ZN(
        npu_inst_pe_1_3_7_n92) );
  NAND2_X1 npu_inst_pe_1_3_7_U44 ( .A1(npu_inst_pe_1_3_7_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_3_7_n48), .ZN(npu_inst_pe_1_3_7_n68) );
  OAI21_X1 npu_inst_pe_1_3_7_U43 ( .B1(npu_inst_pe_1_3_7_n63), .B2(
        npu_inst_pe_1_3_7_n48), .A(npu_inst_pe_1_3_7_n68), .ZN(
        npu_inst_pe_1_3_7_n91) );
  NAND2_X1 npu_inst_pe_1_3_7_U42 ( .A1(npu_inst_pe_1_3_7_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_3_7_n48), .ZN(npu_inst_pe_1_3_7_n67) );
  OAI21_X1 npu_inst_pe_1_3_7_U41 ( .B1(npu_inst_pe_1_3_7_n61), .B2(
        npu_inst_pe_1_3_7_n48), .A(npu_inst_pe_1_3_7_n67), .ZN(
        npu_inst_pe_1_3_7_n90) );
  NAND2_X1 npu_inst_pe_1_3_7_U40 ( .A1(npu_inst_pe_1_3_7_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_3_7_n44), .ZN(npu_inst_pe_1_3_7_n66) );
  OAI21_X1 npu_inst_pe_1_3_7_U39 ( .B1(npu_inst_pe_1_3_7_n63), .B2(
        npu_inst_pe_1_3_7_n44), .A(npu_inst_pe_1_3_7_n66), .ZN(
        npu_inst_pe_1_3_7_n89) );
  NAND2_X1 npu_inst_pe_1_3_7_U38 ( .A1(npu_inst_pe_1_3_7_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_3_7_n44), .ZN(npu_inst_pe_1_3_7_n65) );
  OAI21_X1 npu_inst_pe_1_3_7_U37 ( .B1(npu_inst_pe_1_3_7_n61), .B2(
        npu_inst_pe_1_3_7_n44), .A(npu_inst_pe_1_3_7_n65), .ZN(
        npu_inst_pe_1_3_7_n88) );
  NAND2_X1 npu_inst_pe_1_3_7_U36 ( .A1(npu_inst_pe_1_3_7_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_3_7_n40), .ZN(npu_inst_pe_1_3_7_n64) );
  OAI21_X1 npu_inst_pe_1_3_7_U35 ( .B1(npu_inst_pe_1_3_7_n63), .B2(
        npu_inst_pe_1_3_7_n40), .A(npu_inst_pe_1_3_7_n64), .ZN(
        npu_inst_pe_1_3_7_n87) );
  NAND2_X1 npu_inst_pe_1_3_7_U34 ( .A1(npu_inst_pe_1_3_7_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_3_7_n40), .ZN(npu_inst_pe_1_3_7_n62) );
  OAI21_X1 npu_inst_pe_1_3_7_U33 ( .B1(npu_inst_pe_1_3_7_n61), .B2(
        npu_inst_pe_1_3_7_n40), .A(npu_inst_pe_1_3_7_n62), .ZN(
        npu_inst_pe_1_3_7_n86) );
  INV_X1 npu_inst_pe_1_3_7_U32 ( .A(npu_inst_pe_1_3_7_int_data_0_), .ZN(
        npu_inst_pe_1_3_7_n13) );
  INV_X1 npu_inst_pe_1_3_7_U31 ( .A(npu_inst_n69), .ZN(npu_inst_pe_1_3_7_n5)
         );
  AOI22_X1 npu_inst_pe_1_3_7_U30 ( .A1(npu_inst_n56), .A2(
        npu_inst_int_data_y_4__7__1_), .B1(npu_inst_pe_1_3_7_n3), .B2(
        int_i_data_h_npu[9]), .ZN(npu_inst_pe_1_3_7_n63) );
  AOI22_X1 npu_inst_pe_1_3_7_U29 ( .A1(npu_inst_n56), .A2(
        npu_inst_int_data_y_4__7__0_), .B1(npu_inst_pe_1_3_7_n3), .B2(
        int_i_data_h_npu[8]), .ZN(npu_inst_pe_1_3_7_n61) );
  OR3_X1 npu_inst_pe_1_3_7_U28 ( .A1(npu_inst_pe_1_3_7_n6), .A2(
        npu_inst_pe_1_3_7_n8), .A3(npu_inst_pe_1_3_7_n5), .ZN(
        npu_inst_pe_1_3_7_n56) );
  OR3_X1 npu_inst_pe_1_3_7_U27 ( .A1(npu_inst_pe_1_3_7_n5), .A2(
        npu_inst_pe_1_3_7_n8), .A3(npu_inst_pe_1_3_7_n7), .ZN(
        npu_inst_pe_1_3_7_n48) );
  INV_X1 npu_inst_pe_1_3_7_U26 ( .A(npu_inst_pe_1_3_7_n5), .ZN(
        npu_inst_pe_1_3_7_n4) );
  OR3_X1 npu_inst_pe_1_3_7_U25 ( .A1(npu_inst_pe_1_3_7_n4), .A2(
        npu_inst_pe_1_3_7_n8), .A3(npu_inst_pe_1_3_7_n7), .ZN(
        npu_inst_pe_1_3_7_n52) );
  OR3_X1 npu_inst_pe_1_3_7_U24 ( .A1(npu_inst_pe_1_3_7_n6), .A2(
        npu_inst_pe_1_3_7_n8), .A3(npu_inst_pe_1_3_7_n4), .ZN(
        npu_inst_pe_1_3_7_n60) );
  NOR2_X1 npu_inst_pe_1_3_7_U23 ( .A1(npu_inst_pe_1_3_7_n60), .A2(
        npu_inst_pe_1_3_7_n3), .ZN(npu_inst_pe_1_3_7_n58) );
  NOR2_X1 npu_inst_pe_1_3_7_U22 ( .A1(npu_inst_pe_1_3_7_n56), .A2(
        npu_inst_pe_1_3_7_n3), .ZN(npu_inst_pe_1_3_7_n54) );
  NOR2_X1 npu_inst_pe_1_3_7_U21 ( .A1(npu_inst_pe_1_3_7_n52), .A2(
        npu_inst_pe_1_3_7_n3), .ZN(npu_inst_pe_1_3_7_n50) );
  NOR2_X1 npu_inst_pe_1_3_7_U20 ( .A1(npu_inst_pe_1_3_7_n48), .A2(
        npu_inst_pe_1_3_7_n3), .ZN(npu_inst_pe_1_3_7_n46) );
  NOR2_X1 npu_inst_pe_1_3_7_U19 ( .A1(npu_inst_pe_1_3_7_n40), .A2(
        npu_inst_pe_1_3_7_n3), .ZN(npu_inst_pe_1_3_7_n38) );
  NOR2_X1 npu_inst_pe_1_3_7_U18 ( .A1(npu_inst_pe_1_3_7_n44), .A2(
        npu_inst_pe_1_3_7_n3), .ZN(npu_inst_pe_1_3_7_n42) );
  BUF_X1 npu_inst_pe_1_3_7_U17 ( .A(npu_inst_n100), .Z(npu_inst_pe_1_3_7_n8)
         );
  INV_X1 npu_inst_pe_1_3_7_U16 ( .A(npu_inst_n124), .ZN(npu_inst_pe_1_3_7_n12)
         );
  INV_X1 npu_inst_pe_1_3_7_U15 ( .A(npu_inst_pe_1_3_7_n38), .ZN(
        npu_inst_pe_1_3_7_n114) );
  INV_X1 npu_inst_pe_1_3_7_U14 ( .A(npu_inst_pe_1_3_7_n58), .ZN(
        npu_inst_pe_1_3_7_n119) );
  INV_X1 npu_inst_pe_1_3_7_U13 ( .A(npu_inst_pe_1_3_7_n54), .ZN(
        npu_inst_pe_1_3_7_n118) );
  INV_X1 npu_inst_pe_1_3_7_U12 ( .A(npu_inst_pe_1_3_7_n50), .ZN(
        npu_inst_pe_1_3_7_n117) );
  INV_X1 npu_inst_pe_1_3_7_U11 ( .A(npu_inst_pe_1_3_7_n46), .ZN(
        npu_inst_pe_1_3_7_n116) );
  INV_X1 npu_inst_pe_1_3_7_U10 ( .A(npu_inst_pe_1_3_7_n42), .ZN(
        npu_inst_pe_1_3_7_n115) );
  BUF_X1 npu_inst_pe_1_3_7_U9 ( .A(npu_inst_n23), .Z(npu_inst_pe_1_3_7_n2) );
  BUF_X1 npu_inst_pe_1_3_7_U8 ( .A(npu_inst_n23), .Z(npu_inst_pe_1_3_7_n1) );
  BUF_X1 npu_inst_pe_1_3_7_U7 ( .A(npu_inst_pe_1_3_7_n12), .Z(
        npu_inst_pe_1_3_7_n11) );
  BUF_X1 npu_inst_pe_1_3_7_U6 ( .A(npu_inst_pe_1_3_7_n12), .Z(
        npu_inst_pe_1_3_7_n10) );
  BUF_X1 npu_inst_pe_1_3_7_U5 ( .A(npu_inst_pe_1_3_7_n12), .Z(
        npu_inst_pe_1_3_7_n9) );
  NOR2_X1 npu_inst_pe_1_3_7_U4 ( .A1(npu_inst_pe_1_3_7_int_q_weight_0_), .A2(
        npu_inst_pe_1_3_7_n1), .ZN(npu_inst_pe_1_3_7_n76) );
  NOR2_X1 npu_inst_pe_1_3_7_U3 ( .A1(npu_inst_pe_1_3_7_n27), .A2(
        npu_inst_pe_1_3_7_n1), .ZN(npu_inst_pe_1_3_7_n77) );
  FA_X1 npu_inst_pe_1_3_7_sub_67_U2_1 ( .A(npu_inst_pe_1_3_7_int_q_acc_1_), 
        .B(npu_inst_pe_1_3_7_n14), .CI(npu_inst_pe_1_3_7_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_3_7_sub_67_carry_2_), .S(npu_inst_pe_1_3_7_N66) );
  FA_X1 npu_inst_pe_1_3_7_add_69_U1_1 ( .A(npu_inst_pe_1_3_7_int_q_acc_1_), 
        .B(npu_inst_pe_1_3_7_int_data_1_), .CI(
        npu_inst_pe_1_3_7_add_69_carry_1_), .CO(
        npu_inst_pe_1_3_7_add_69_carry_2_), .S(npu_inst_pe_1_3_7_N74) );
  NAND3_X1 npu_inst_pe_1_3_7_U109 ( .A1(npu_inst_pe_1_3_7_n5), .A2(
        npu_inst_pe_1_3_7_n7), .A3(npu_inst_pe_1_3_7_n8), .ZN(
        npu_inst_pe_1_3_7_n44) );
  NAND3_X1 npu_inst_pe_1_3_7_U108 ( .A1(npu_inst_pe_1_3_7_n4), .A2(
        npu_inst_pe_1_3_7_n7), .A3(npu_inst_pe_1_3_7_n8), .ZN(
        npu_inst_pe_1_3_7_n40) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_3_7_n34), .CK(
        npu_inst_pe_1_3_7_net3849), .RN(npu_inst_pe_1_3_7_n9), .Q(
        npu_inst_pe_1_3_7_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_3_7_n35), .CK(
        npu_inst_pe_1_3_7_net3849), .RN(npu_inst_pe_1_3_7_n9), .Q(
        npu_inst_pe_1_3_7_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_3_7_n36), .CK(
        npu_inst_pe_1_3_7_net3849), .RN(npu_inst_pe_1_3_7_n9), .Q(
        npu_inst_pe_1_3_7_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_3_7_n98), .CK(
        npu_inst_pe_1_3_7_net3849), .RN(npu_inst_pe_1_3_7_n9), .Q(
        npu_inst_pe_1_3_7_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_3_7_n99), .CK(
        npu_inst_pe_1_3_7_net3849), .RN(npu_inst_pe_1_3_7_n9), .Q(
        npu_inst_pe_1_3_7_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_3_7_n100), 
        .CK(npu_inst_pe_1_3_7_net3849), .RN(npu_inst_pe_1_3_7_n9), .Q(
        npu_inst_pe_1_3_7_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_3_7_n33), .CK(
        npu_inst_pe_1_3_7_net3849), .RN(npu_inst_pe_1_3_7_n9), .Q(
        npu_inst_pe_1_3_7_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_3_7_n101), 
        .CK(npu_inst_pe_1_3_7_net3849), .RN(npu_inst_pe_1_3_7_n9), .Q(
        npu_inst_pe_1_3_7_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_weight_reg_0_ ( .D(npu_inst_n110), .CK(
        npu_inst_pe_1_3_7_net3855), .RN(npu_inst_pe_1_3_7_n9), .Q(
        npu_inst_pe_1_3_7_int_q_weight_0_), .QN(npu_inst_pe_1_3_7_n27) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_weight_reg_1_ ( .D(npu_inst_n116), .CK(
        npu_inst_pe_1_3_7_net3855), .RN(npu_inst_pe_1_3_7_n9), .Q(
        npu_inst_pe_1_3_7_int_q_weight_1_), .QN(npu_inst_pe_1_3_7_n26) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_3_7_n113), 
        .CK(npu_inst_pe_1_3_7_net3855), .RN(npu_inst_pe_1_3_7_n9), .Q(
        npu_inst_pe_1_3_7_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_3_7_n107), 
        .CK(npu_inst_pe_1_3_7_net3855), .RN(npu_inst_pe_1_3_7_n9), .Q(
        npu_inst_pe_1_3_7_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_3_7_n112), 
        .CK(npu_inst_pe_1_3_7_net3855), .RN(npu_inst_pe_1_3_7_n10), .Q(
        npu_inst_pe_1_3_7_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_3_7_n106), 
        .CK(npu_inst_pe_1_3_7_net3855), .RN(npu_inst_pe_1_3_7_n10), .Q(
        npu_inst_pe_1_3_7_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_3_7_n111), 
        .CK(npu_inst_pe_1_3_7_net3855), .RN(npu_inst_pe_1_3_7_n10), .Q(
        npu_inst_pe_1_3_7_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_3_7_n105), 
        .CK(npu_inst_pe_1_3_7_net3855), .RN(npu_inst_pe_1_3_7_n10), .Q(
        npu_inst_pe_1_3_7_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_3_7_n110), 
        .CK(npu_inst_pe_1_3_7_net3855), .RN(npu_inst_pe_1_3_7_n10), .Q(
        npu_inst_pe_1_3_7_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_3_7_n104), 
        .CK(npu_inst_pe_1_3_7_net3855), .RN(npu_inst_pe_1_3_7_n10), .Q(
        npu_inst_pe_1_3_7_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_3_7_n109), 
        .CK(npu_inst_pe_1_3_7_net3855), .RN(npu_inst_pe_1_3_7_n10), .Q(
        npu_inst_pe_1_3_7_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_3_7_n103), 
        .CK(npu_inst_pe_1_3_7_net3855), .RN(npu_inst_pe_1_3_7_n10), .Q(
        npu_inst_pe_1_3_7_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_3_7_n108), 
        .CK(npu_inst_pe_1_3_7_net3855), .RN(npu_inst_pe_1_3_7_n10), .Q(
        npu_inst_pe_1_3_7_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_3_7_n102), 
        .CK(npu_inst_pe_1_3_7_net3855), .RN(npu_inst_pe_1_3_7_n10), .Q(
        npu_inst_pe_1_3_7_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_3_7_n86), 
        .CK(npu_inst_pe_1_3_7_net3855), .RN(npu_inst_pe_1_3_7_n10), .Q(
        npu_inst_pe_1_3_7_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_3_7_n87), 
        .CK(npu_inst_pe_1_3_7_net3855), .RN(npu_inst_pe_1_3_7_n10), .Q(
        npu_inst_pe_1_3_7_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_3_7_n88), 
        .CK(npu_inst_pe_1_3_7_net3855), .RN(npu_inst_pe_1_3_7_n11), .Q(
        npu_inst_pe_1_3_7_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_3_7_n89), 
        .CK(npu_inst_pe_1_3_7_net3855), .RN(npu_inst_pe_1_3_7_n11), .Q(
        npu_inst_pe_1_3_7_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_3_7_n90), 
        .CK(npu_inst_pe_1_3_7_net3855), .RN(npu_inst_pe_1_3_7_n11), .Q(
        npu_inst_pe_1_3_7_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_3_7_n91), 
        .CK(npu_inst_pe_1_3_7_net3855), .RN(npu_inst_pe_1_3_7_n11), .Q(
        npu_inst_pe_1_3_7_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_3_7_n92), 
        .CK(npu_inst_pe_1_3_7_net3855), .RN(npu_inst_pe_1_3_7_n11), .Q(
        npu_inst_pe_1_3_7_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_3_7_n93), 
        .CK(npu_inst_pe_1_3_7_net3855), .RN(npu_inst_pe_1_3_7_n11), .Q(
        npu_inst_pe_1_3_7_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_3_7_n94), 
        .CK(npu_inst_pe_1_3_7_net3855), .RN(npu_inst_pe_1_3_7_n11), .Q(
        npu_inst_pe_1_3_7_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_3_7_n95), 
        .CK(npu_inst_pe_1_3_7_net3855), .RN(npu_inst_pe_1_3_7_n11), .Q(
        npu_inst_pe_1_3_7_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_3_7_n96), 
        .CK(npu_inst_pe_1_3_7_net3855), .RN(npu_inst_pe_1_3_7_n11), .Q(
        npu_inst_pe_1_3_7_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_3_7_n97), 
        .CK(npu_inst_pe_1_3_7_net3855), .RN(npu_inst_pe_1_3_7_n11), .Q(
        npu_inst_pe_1_3_7_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_3_7_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_3_7_N84), .SE(1'b0), .GCK(npu_inst_pe_1_3_7_net3849) );
  CLKGATETST_X1 npu_inst_pe_1_3_7_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n63), .SE(1'b0), .GCK(npu_inst_pe_1_3_7_net3855) );
  MUX2_X1 npu_inst_pe_1_4_0_U162 ( .A(npu_inst_pe_1_4_0_n32), .B(
        npu_inst_pe_1_4_0_n29), .S(npu_inst_pe_1_4_0_n8), .Z(
        npu_inst_pe_1_4_0_N93) );
  MUX2_X1 npu_inst_pe_1_4_0_U161 ( .A(npu_inst_pe_1_4_0_n31), .B(
        npu_inst_pe_1_4_0_n30), .S(npu_inst_pe_1_4_0_n6), .Z(
        npu_inst_pe_1_4_0_n32) );
  MUX2_X1 npu_inst_pe_1_4_0_U160 ( .A(npu_inst_pe_1_4_0_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_4_0_int_q_reg_v_1__0_), .S(npu_inst_pe_1_4_0_n4), .Z(
        npu_inst_pe_1_4_0_n31) );
  MUX2_X1 npu_inst_pe_1_4_0_U159 ( .A(npu_inst_pe_1_4_0_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_4_0_int_q_reg_v_3__0_), .S(npu_inst_pe_1_4_0_n4), .Z(
        npu_inst_pe_1_4_0_n30) );
  MUX2_X1 npu_inst_pe_1_4_0_U158 ( .A(npu_inst_pe_1_4_0_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_4_0_int_q_reg_v_5__0_), .S(npu_inst_pe_1_4_0_n4), .Z(
        npu_inst_pe_1_4_0_n29) );
  MUX2_X1 npu_inst_pe_1_4_0_U157 ( .A(npu_inst_pe_1_4_0_n28), .B(
        npu_inst_pe_1_4_0_n23), .S(npu_inst_pe_1_4_0_n8), .Z(
        npu_inst_pe_1_4_0_N94) );
  MUX2_X1 npu_inst_pe_1_4_0_U156 ( .A(npu_inst_pe_1_4_0_n25), .B(
        npu_inst_pe_1_4_0_n24), .S(npu_inst_pe_1_4_0_n6), .Z(
        npu_inst_pe_1_4_0_n28) );
  MUX2_X1 npu_inst_pe_1_4_0_U155 ( .A(npu_inst_pe_1_4_0_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_4_0_int_q_reg_v_1__1_), .S(npu_inst_pe_1_4_0_n4), .Z(
        npu_inst_pe_1_4_0_n25) );
  MUX2_X1 npu_inst_pe_1_4_0_U154 ( .A(npu_inst_pe_1_4_0_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_4_0_int_q_reg_v_3__1_), .S(npu_inst_pe_1_4_0_n4), .Z(
        npu_inst_pe_1_4_0_n24) );
  MUX2_X1 npu_inst_pe_1_4_0_U153 ( .A(npu_inst_pe_1_4_0_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_4_0_int_q_reg_v_5__1_), .S(npu_inst_pe_1_4_0_n4), .Z(
        npu_inst_pe_1_4_0_n23) );
  MUX2_X1 npu_inst_pe_1_4_0_U152 ( .A(npu_inst_pe_1_4_0_n22), .B(
        npu_inst_pe_1_4_0_n19), .S(npu_inst_pe_1_4_0_n8), .Z(
        npu_inst_pe_1_4_0_o_data_h_1_) );
  MUX2_X1 npu_inst_pe_1_4_0_U151 ( .A(npu_inst_pe_1_4_0_n21), .B(
        npu_inst_pe_1_4_0_n20), .S(npu_inst_pe_1_4_0_n6), .Z(
        npu_inst_pe_1_4_0_n22) );
  MUX2_X1 npu_inst_pe_1_4_0_U150 ( .A(npu_inst_pe_1_4_0_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_4_0_int_q_reg_h_1__1_), .S(npu_inst_pe_1_4_0_n4), .Z(
        npu_inst_pe_1_4_0_n21) );
  MUX2_X1 npu_inst_pe_1_4_0_U149 ( .A(npu_inst_pe_1_4_0_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_4_0_int_q_reg_h_3__1_), .S(npu_inst_pe_1_4_0_n4), .Z(
        npu_inst_pe_1_4_0_n20) );
  MUX2_X1 npu_inst_pe_1_4_0_U148 ( .A(npu_inst_pe_1_4_0_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_4_0_int_q_reg_h_5__1_), .S(npu_inst_pe_1_4_0_n4), .Z(
        npu_inst_pe_1_4_0_n19) );
  MUX2_X1 npu_inst_pe_1_4_0_U147 ( .A(npu_inst_pe_1_4_0_n18), .B(
        npu_inst_pe_1_4_0_n15), .S(npu_inst_pe_1_4_0_n8), .Z(
        npu_inst_pe_1_4_0_o_data_h_0_) );
  MUX2_X1 npu_inst_pe_1_4_0_U146 ( .A(npu_inst_pe_1_4_0_n17), .B(
        npu_inst_pe_1_4_0_n16), .S(npu_inst_pe_1_4_0_n6), .Z(
        npu_inst_pe_1_4_0_n18) );
  MUX2_X1 npu_inst_pe_1_4_0_U145 ( .A(npu_inst_pe_1_4_0_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_4_0_int_q_reg_h_1__0_), .S(npu_inst_pe_1_4_0_n4), .Z(
        npu_inst_pe_1_4_0_n17) );
  MUX2_X1 npu_inst_pe_1_4_0_U144 ( .A(npu_inst_pe_1_4_0_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_4_0_int_q_reg_h_3__0_), .S(npu_inst_pe_1_4_0_n4), .Z(
        npu_inst_pe_1_4_0_n16) );
  MUX2_X1 npu_inst_pe_1_4_0_U143 ( .A(npu_inst_pe_1_4_0_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_4_0_int_q_reg_h_5__0_), .S(npu_inst_pe_1_4_0_n4), .Z(
        npu_inst_pe_1_4_0_n15) );
  XOR2_X1 npu_inst_pe_1_4_0_U142 ( .A(npu_inst_pe_1_4_0_int_data_0_), .B(
        npu_inst_pe_1_4_0_int_q_acc_0_), .Z(npu_inst_pe_1_4_0_N73) );
  AND2_X1 npu_inst_pe_1_4_0_U141 ( .A1(npu_inst_pe_1_4_0_int_q_acc_0_), .A2(
        npu_inst_pe_1_4_0_int_data_0_), .ZN(npu_inst_pe_1_4_0_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_4_0_U140 ( .A(npu_inst_pe_1_4_0_int_q_acc_0_), .B(
        npu_inst_pe_1_4_0_n13), .ZN(npu_inst_pe_1_4_0_N65) );
  OR2_X1 npu_inst_pe_1_4_0_U139 ( .A1(npu_inst_pe_1_4_0_n13), .A2(
        npu_inst_pe_1_4_0_int_q_acc_0_), .ZN(npu_inst_pe_1_4_0_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_4_0_U138 ( .A(npu_inst_pe_1_4_0_int_q_acc_2_), .B(
        npu_inst_pe_1_4_0_add_69_carry_2_), .Z(npu_inst_pe_1_4_0_N75) );
  AND2_X1 npu_inst_pe_1_4_0_U137 ( .A1(npu_inst_pe_1_4_0_add_69_carry_2_), 
        .A2(npu_inst_pe_1_4_0_int_q_acc_2_), .ZN(
        npu_inst_pe_1_4_0_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_4_0_U136 ( .A(npu_inst_pe_1_4_0_int_q_acc_3_), .B(
        npu_inst_pe_1_4_0_add_69_carry_3_), .Z(npu_inst_pe_1_4_0_N76) );
  AND2_X1 npu_inst_pe_1_4_0_U135 ( .A1(npu_inst_pe_1_4_0_add_69_carry_3_), 
        .A2(npu_inst_pe_1_4_0_int_q_acc_3_), .ZN(
        npu_inst_pe_1_4_0_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_4_0_U134 ( .A(npu_inst_pe_1_4_0_int_q_acc_4_), .B(
        npu_inst_pe_1_4_0_add_69_carry_4_), .Z(npu_inst_pe_1_4_0_N77) );
  AND2_X1 npu_inst_pe_1_4_0_U133 ( .A1(npu_inst_pe_1_4_0_add_69_carry_4_), 
        .A2(npu_inst_pe_1_4_0_int_q_acc_4_), .ZN(
        npu_inst_pe_1_4_0_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_4_0_U132 ( .A(npu_inst_pe_1_4_0_int_q_acc_5_), .B(
        npu_inst_pe_1_4_0_add_69_carry_5_), .Z(npu_inst_pe_1_4_0_N78) );
  AND2_X1 npu_inst_pe_1_4_0_U131 ( .A1(npu_inst_pe_1_4_0_add_69_carry_5_), 
        .A2(npu_inst_pe_1_4_0_int_q_acc_5_), .ZN(
        npu_inst_pe_1_4_0_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_4_0_U130 ( .A(npu_inst_pe_1_4_0_int_q_acc_6_), .B(
        npu_inst_pe_1_4_0_add_69_carry_6_), .Z(npu_inst_pe_1_4_0_N79) );
  AND2_X1 npu_inst_pe_1_4_0_U129 ( .A1(npu_inst_pe_1_4_0_add_69_carry_6_), 
        .A2(npu_inst_pe_1_4_0_int_q_acc_6_), .ZN(
        npu_inst_pe_1_4_0_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_4_0_U128 ( .A(npu_inst_pe_1_4_0_int_q_acc_7_), .B(
        npu_inst_pe_1_4_0_add_69_carry_7_), .Z(npu_inst_pe_1_4_0_N80) );
  XNOR2_X1 npu_inst_pe_1_4_0_U127 ( .A(npu_inst_pe_1_4_0_sub_67_carry_2_), .B(
        npu_inst_pe_1_4_0_int_q_acc_2_), .ZN(npu_inst_pe_1_4_0_N67) );
  OR2_X1 npu_inst_pe_1_4_0_U126 ( .A1(npu_inst_pe_1_4_0_int_q_acc_2_), .A2(
        npu_inst_pe_1_4_0_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_4_0_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_4_0_U125 ( .A(npu_inst_pe_1_4_0_sub_67_carry_3_), .B(
        npu_inst_pe_1_4_0_int_q_acc_3_), .ZN(npu_inst_pe_1_4_0_N68) );
  OR2_X1 npu_inst_pe_1_4_0_U124 ( .A1(npu_inst_pe_1_4_0_int_q_acc_3_), .A2(
        npu_inst_pe_1_4_0_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_4_0_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_4_0_U123 ( .A(npu_inst_pe_1_4_0_sub_67_carry_4_), .B(
        npu_inst_pe_1_4_0_int_q_acc_4_), .ZN(npu_inst_pe_1_4_0_N69) );
  OR2_X1 npu_inst_pe_1_4_0_U122 ( .A1(npu_inst_pe_1_4_0_int_q_acc_4_), .A2(
        npu_inst_pe_1_4_0_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_4_0_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_4_0_U121 ( .A(npu_inst_pe_1_4_0_sub_67_carry_5_), .B(
        npu_inst_pe_1_4_0_int_q_acc_5_), .ZN(npu_inst_pe_1_4_0_N70) );
  OR2_X1 npu_inst_pe_1_4_0_U120 ( .A1(npu_inst_pe_1_4_0_int_q_acc_5_), .A2(
        npu_inst_pe_1_4_0_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_4_0_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_4_0_U119 ( .A(npu_inst_pe_1_4_0_sub_67_carry_6_), .B(
        npu_inst_pe_1_4_0_int_q_acc_6_), .ZN(npu_inst_pe_1_4_0_N71) );
  OR2_X1 npu_inst_pe_1_4_0_U118 ( .A1(npu_inst_pe_1_4_0_int_q_acc_6_), .A2(
        npu_inst_pe_1_4_0_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_4_0_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_4_0_U117 ( .A(npu_inst_pe_1_4_0_int_q_acc_7_), .B(
        npu_inst_pe_1_4_0_sub_67_carry_7_), .ZN(npu_inst_pe_1_4_0_N72) );
  INV_X1 npu_inst_pe_1_4_0_U116 ( .A(npu_inst_n77), .ZN(npu_inst_pe_1_4_0_n7)
         );
  INV_X1 npu_inst_pe_1_4_0_U115 ( .A(npu_inst_pe_1_4_0_n7), .ZN(
        npu_inst_pe_1_4_0_n6) );
  INV_X1 npu_inst_pe_1_4_0_U114 ( .A(npu_inst_n56), .ZN(npu_inst_pe_1_4_0_n3)
         );
  AOI22_X1 npu_inst_pe_1_4_0_U113 ( .A1(npu_inst_int_data_y_5__0__0_), .A2(
        npu_inst_pe_1_4_0_n58), .B1(npu_inst_pe_1_4_0_n119), .B2(
        npu_inst_pe_1_4_0_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_4_0_n57) );
  INV_X1 npu_inst_pe_1_4_0_U112 ( .A(npu_inst_pe_1_4_0_n57), .ZN(
        npu_inst_pe_1_4_0_n108) );
  AOI22_X1 npu_inst_pe_1_4_0_U111 ( .A1(npu_inst_int_data_y_5__0__0_), .A2(
        npu_inst_pe_1_4_0_n54), .B1(npu_inst_pe_1_4_0_n118), .B2(
        npu_inst_pe_1_4_0_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_4_0_n53) );
  INV_X1 npu_inst_pe_1_4_0_U110 ( .A(npu_inst_pe_1_4_0_n53), .ZN(
        npu_inst_pe_1_4_0_n109) );
  AOI22_X1 npu_inst_pe_1_4_0_U107 ( .A1(npu_inst_int_data_y_5__0__0_), .A2(
        npu_inst_pe_1_4_0_n50), .B1(npu_inst_pe_1_4_0_n117), .B2(
        npu_inst_pe_1_4_0_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_4_0_n49) );
  INV_X1 npu_inst_pe_1_4_0_U106 ( .A(npu_inst_pe_1_4_0_n49), .ZN(
        npu_inst_pe_1_4_0_n110) );
  AOI22_X1 npu_inst_pe_1_4_0_U105 ( .A1(npu_inst_int_data_y_5__0__0_), .A2(
        npu_inst_pe_1_4_0_n46), .B1(npu_inst_pe_1_4_0_n116), .B2(
        npu_inst_pe_1_4_0_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_4_0_n45) );
  INV_X1 npu_inst_pe_1_4_0_U104 ( .A(npu_inst_pe_1_4_0_n45), .ZN(
        npu_inst_pe_1_4_0_n111) );
  AOI22_X1 npu_inst_pe_1_4_0_U103 ( .A1(npu_inst_int_data_y_5__0__0_), .A2(
        npu_inst_pe_1_4_0_n42), .B1(npu_inst_pe_1_4_0_n115), .B2(
        npu_inst_pe_1_4_0_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_4_0_n41) );
  INV_X1 npu_inst_pe_1_4_0_U102 ( .A(npu_inst_pe_1_4_0_n41), .ZN(
        npu_inst_pe_1_4_0_n112) );
  AOI22_X1 npu_inst_pe_1_4_0_U101 ( .A1(npu_inst_int_data_y_5__0__1_), .A2(
        npu_inst_pe_1_4_0_n58), .B1(npu_inst_pe_1_4_0_n119), .B2(
        npu_inst_pe_1_4_0_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_4_0_n59) );
  INV_X1 npu_inst_pe_1_4_0_U100 ( .A(npu_inst_pe_1_4_0_n59), .ZN(
        npu_inst_pe_1_4_0_n102) );
  AOI22_X1 npu_inst_pe_1_4_0_U99 ( .A1(npu_inst_int_data_y_5__0__1_), .A2(
        npu_inst_pe_1_4_0_n54), .B1(npu_inst_pe_1_4_0_n118), .B2(
        npu_inst_pe_1_4_0_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_4_0_n55) );
  INV_X1 npu_inst_pe_1_4_0_U98 ( .A(npu_inst_pe_1_4_0_n55), .ZN(
        npu_inst_pe_1_4_0_n103) );
  AOI22_X1 npu_inst_pe_1_4_0_U97 ( .A1(npu_inst_int_data_y_5__0__1_), .A2(
        npu_inst_pe_1_4_0_n50), .B1(npu_inst_pe_1_4_0_n117), .B2(
        npu_inst_pe_1_4_0_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_4_0_n51) );
  INV_X1 npu_inst_pe_1_4_0_U96 ( .A(npu_inst_pe_1_4_0_n51), .ZN(
        npu_inst_pe_1_4_0_n104) );
  AOI22_X1 npu_inst_pe_1_4_0_U95 ( .A1(npu_inst_int_data_y_5__0__1_), .A2(
        npu_inst_pe_1_4_0_n46), .B1(npu_inst_pe_1_4_0_n116), .B2(
        npu_inst_pe_1_4_0_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_4_0_n47) );
  INV_X1 npu_inst_pe_1_4_0_U94 ( .A(npu_inst_pe_1_4_0_n47), .ZN(
        npu_inst_pe_1_4_0_n105) );
  AOI22_X1 npu_inst_pe_1_4_0_U93 ( .A1(npu_inst_int_data_y_5__0__1_), .A2(
        npu_inst_pe_1_4_0_n42), .B1(npu_inst_pe_1_4_0_n115), .B2(
        npu_inst_pe_1_4_0_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_4_0_n43) );
  INV_X1 npu_inst_pe_1_4_0_U92 ( .A(npu_inst_pe_1_4_0_n43), .ZN(
        npu_inst_pe_1_4_0_n106) );
  AOI22_X1 npu_inst_pe_1_4_0_U91 ( .A1(npu_inst_pe_1_4_0_n38), .A2(
        npu_inst_int_data_y_5__0__1_), .B1(npu_inst_pe_1_4_0_n114), .B2(
        npu_inst_pe_1_4_0_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_4_0_n39) );
  INV_X1 npu_inst_pe_1_4_0_U90 ( .A(npu_inst_pe_1_4_0_n39), .ZN(
        npu_inst_pe_1_4_0_n107) );
  AOI22_X1 npu_inst_pe_1_4_0_U89 ( .A1(npu_inst_pe_1_4_0_n38), .A2(
        npu_inst_int_data_y_5__0__0_), .B1(npu_inst_pe_1_4_0_n114), .B2(
        npu_inst_pe_1_4_0_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_4_0_n37) );
  INV_X1 npu_inst_pe_1_4_0_U88 ( .A(npu_inst_pe_1_4_0_n37), .ZN(
        npu_inst_pe_1_4_0_n113) );
  NOR3_X1 npu_inst_pe_1_4_0_U87 ( .A1(npu_inst_pe_1_4_0_n26), .A2(npu_inst_n56), .A3(npu_inst_int_ckg[31]), .ZN(npu_inst_pe_1_4_0_n85) );
  OR2_X1 npu_inst_pe_1_4_0_U86 ( .A1(npu_inst_pe_1_4_0_n85), .A2(
        npu_inst_pe_1_4_0_n2), .ZN(npu_inst_pe_1_4_0_N84) );
  NAND2_X1 npu_inst_pe_1_4_0_U85 ( .A1(npu_inst_pe_1_4_0_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_4_0_n60), .ZN(npu_inst_pe_1_4_0_n74) );
  OAI21_X1 npu_inst_pe_1_4_0_U84 ( .B1(npu_inst_pe_1_4_0_n63), .B2(
        npu_inst_pe_1_4_0_n60), .A(npu_inst_pe_1_4_0_n74), .ZN(
        npu_inst_pe_1_4_0_n97) );
  NAND2_X1 npu_inst_pe_1_4_0_U83 ( .A1(npu_inst_pe_1_4_0_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_4_0_n60), .ZN(npu_inst_pe_1_4_0_n73) );
  OAI21_X1 npu_inst_pe_1_4_0_U82 ( .B1(npu_inst_pe_1_4_0_n61), .B2(
        npu_inst_pe_1_4_0_n60), .A(npu_inst_pe_1_4_0_n73), .ZN(
        npu_inst_pe_1_4_0_n96) );
  NAND2_X1 npu_inst_pe_1_4_0_U81 ( .A1(npu_inst_pe_1_4_0_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_4_0_n56), .ZN(npu_inst_pe_1_4_0_n72) );
  OAI21_X1 npu_inst_pe_1_4_0_U80 ( .B1(npu_inst_pe_1_4_0_n63), .B2(
        npu_inst_pe_1_4_0_n56), .A(npu_inst_pe_1_4_0_n72), .ZN(
        npu_inst_pe_1_4_0_n95) );
  NAND2_X1 npu_inst_pe_1_4_0_U79 ( .A1(npu_inst_pe_1_4_0_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_4_0_n56), .ZN(npu_inst_pe_1_4_0_n71) );
  OAI21_X1 npu_inst_pe_1_4_0_U78 ( .B1(npu_inst_pe_1_4_0_n61), .B2(
        npu_inst_pe_1_4_0_n56), .A(npu_inst_pe_1_4_0_n71), .ZN(
        npu_inst_pe_1_4_0_n94) );
  NAND2_X1 npu_inst_pe_1_4_0_U77 ( .A1(npu_inst_pe_1_4_0_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_4_0_n52), .ZN(npu_inst_pe_1_4_0_n70) );
  OAI21_X1 npu_inst_pe_1_4_0_U76 ( .B1(npu_inst_pe_1_4_0_n63), .B2(
        npu_inst_pe_1_4_0_n52), .A(npu_inst_pe_1_4_0_n70), .ZN(
        npu_inst_pe_1_4_0_n93) );
  NAND2_X1 npu_inst_pe_1_4_0_U75 ( .A1(npu_inst_pe_1_4_0_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_4_0_n52), .ZN(npu_inst_pe_1_4_0_n69) );
  OAI21_X1 npu_inst_pe_1_4_0_U74 ( .B1(npu_inst_pe_1_4_0_n61), .B2(
        npu_inst_pe_1_4_0_n52), .A(npu_inst_pe_1_4_0_n69), .ZN(
        npu_inst_pe_1_4_0_n92) );
  NAND2_X1 npu_inst_pe_1_4_0_U73 ( .A1(npu_inst_pe_1_4_0_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_4_0_n48), .ZN(npu_inst_pe_1_4_0_n68) );
  OAI21_X1 npu_inst_pe_1_4_0_U72 ( .B1(npu_inst_pe_1_4_0_n63), .B2(
        npu_inst_pe_1_4_0_n48), .A(npu_inst_pe_1_4_0_n68), .ZN(
        npu_inst_pe_1_4_0_n91) );
  NAND2_X1 npu_inst_pe_1_4_0_U71 ( .A1(npu_inst_pe_1_4_0_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_4_0_n48), .ZN(npu_inst_pe_1_4_0_n67) );
  OAI21_X1 npu_inst_pe_1_4_0_U70 ( .B1(npu_inst_pe_1_4_0_n61), .B2(
        npu_inst_pe_1_4_0_n48), .A(npu_inst_pe_1_4_0_n67), .ZN(
        npu_inst_pe_1_4_0_n90) );
  NAND2_X1 npu_inst_pe_1_4_0_U69 ( .A1(npu_inst_pe_1_4_0_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_4_0_n44), .ZN(npu_inst_pe_1_4_0_n66) );
  OAI21_X1 npu_inst_pe_1_4_0_U68 ( .B1(npu_inst_pe_1_4_0_n63), .B2(
        npu_inst_pe_1_4_0_n44), .A(npu_inst_pe_1_4_0_n66), .ZN(
        npu_inst_pe_1_4_0_n89) );
  NAND2_X1 npu_inst_pe_1_4_0_U67 ( .A1(npu_inst_pe_1_4_0_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_4_0_n44), .ZN(npu_inst_pe_1_4_0_n65) );
  OAI21_X1 npu_inst_pe_1_4_0_U66 ( .B1(npu_inst_pe_1_4_0_n61), .B2(
        npu_inst_pe_1_4_0_n44), .A(npu_inst_pe_1_4_0_n65), .ZN(
        npu_inst_pe_1_4_0_n88) );
  NAND2_X1 npu_inst_pe_1_4_0_U65 ( .A1(npu_inst_pe_1_4_0_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_4_0_n40), .ZN(npu_inst_pe_1_4_0_n64) );
  OAI21_X1 npu_inst_pe_1_4_0_U64 ( .B1(npu_inst_pe_1_4_0_n63), .B2(
        npu_inst_pe_1_4_0_n40), .A(npu_inst_pe_1_4_0_n64), .ZN(
        npu_inst_pe_1_4_0_n87) );
  NAND2_X1 npu_inst_pe_1_4_0_U63 ( .A1(npu_inst_pe_1_4_0_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_4_0_n40), .ZN(npu_inst_pe_1_4_0_n62) );
  OAI21_X1 npu_inst_pe_1_4_0_U62 ( .B1(npu_inst_pe_1_4_0_n61), .B2(
        npu_inst_pe_1_4_0_n40), .A(npu_inst_pe_1_4_0_n62), .ZN(
        npu_inst_pe_1_4_0_n86) );
  AND2_X1 npu_inst_pe_1_4_0_U61 ( .A1(npu_inst_pe_1_4_0_N93), .A2(npu_inst_n56), .ZN(npu_inst_int_data_y_4__0__0_) );
  AND2_X1 npu_inst_pe_1_4_0_U60 ( .A1(npu_inst_n56), .A2(npu_inst_pe_1_4_0_N94), .ZN(npu_inst_int_data_y_4__0__1_) );
  AND2_X1 npu_inst_pe_1_4_0_U59 ( .A1(npu_inst_pe_1_4_0_int_q_acc_0_), .A2(
        npu_inst_pe_1_4_0_n1), .ZN(npu_inst_int_data_res_4__0__0_) );
  AND2_X1 npu_inst_pe_1_4_0_U58 ( .A1(npu_inst_pe_1_4_0_n2), .A2(
        npu_inst_pe_1_4_0_int_q_acc_7_), .ZN(npu_inst_int_data_res_4__0__7_)
         );
  AND2_X1 npu_inst_pe_1_4_0_U57 ( .A1(npu_inst_pe_1_4_0_int_q_acc_1_), .A2(
        npu_inst_pe_1_4_0_n1), .ZN(npu_inst_int_data_res_4__0__1_) );
  AND2_X1 npu_inst_pe_1_4_0_U56 ( .A1(npu_inst_pe_1_4_0_int_q_acc_2_), .A2(
        npu_inst_pe_1_4_0_n1), .ZN(npu_inst_int_data_res_4__0__2_) );
  AND2_X1 npu_inst_pe_1_4_0_U55 ( .A1(npu_inst_pe_1_4_0_int_q_acc_3_), .A2(
        npu_inst_pe_1_4_0_n2), .ZN(npu_inst_int_data_res_4__0__3_) );
  AND2_X1 npu_inst_pe_1_4_0_U54 ( .A1(npu_inst_pe_1_4_0_int_q_acc_4_), .A2(
        npu_inst_pe_1_4_0_n2), .ZN(npu_inst_int_data_res_4__0__4_) );
  AND2_X1 npu_inst_pe_1_4_0_U53 ( .A1(npu_inst_pe_1_4_0_int_q_acc_5_), .A2(
        npu_inst_pe_1_4_0_n2), .ZN(npu_inst_int_data_res_4__0__5_) );
  AND2_X1 npu_inst_pe_1_4_0_U52 ( .A1(npu_inst_pe_1_4_0_int_q_acc_6_), .A2(
        npu_inst_pe_1_4_0_n2), .ZN(npu_inst_int_data_res_4__0__6_) );
  AOI222_X1 npu_inst_pe_1_4_0_U51 ( .A1(npu_inst_int_data_res_5__0__0_), .A2(
        npu_inst_pe_1_4_0_n1), .B1(npu_inst_pe_1_4_0_N73), .B2(
        npu_inst_pe_1_4_0_n76), .C1(npu_inst_pe_1_4_0_N65), .C2(
        npu_inst_pe_1_4_0_n77), .ZN(npu_inst_pe_1_4_0_n84) );
  INV_X1 npu_inst_pe_1_4_0_U50 ( .A(npu_inst_pe_1_4_0_n84), .ZN(
        npu_inst_pe_1_4_0_n101) );
  AOI222_X1 npu_inst_pe_1_4_0_U49 ( .A1(npu_inst_int_data_res_5__0__7_), .A2(
        npu_inst_pe_1_4_0_n1), .B1(npu_inst_pe_1_4_0_N80), .B2(
        npu_inst_pe_1_4_0_n76), .C1(npu_inst_pe_1_4_0_N72), .C2(
        npu_inst_pe_1_4_0_n77), .ZN(npu_inst_pe_1_4_0_n75) );
  INV_X1 npu_inst_pe_1_4_0_U48 ( .A(npu_inst_pe_1_4_0_n75), .ZN(
        npu_inst_pe_1_4_0_n33) );
  AOI222_X1 npu_inst_pe_1_4_0_U47 ( .A1(npu_inst_int_data_res_5__0__1_), .A2(
        npu_inst_pe_1_4_0_n1), .B1(npu_inst_pe_1_4_0_N74), .B2(
        npu_inst_pe_1_4_0_n76), .C1(npu_inst_pe_1_4_0_N66), .C2(
        npu_inst_pe_1_4_0_n77), .ZN(npu_inst_pe_1_4_0_n83) );
  INV_X1 npu_inst_pe_1_4_0_U46 ( .A(npu_inst_pe_1_4_0_n83), .ZN(
        npu_inst_pe_1_4_0_n100) );
  AOI222_X1 npu_inst_pe_1_4_0_U45 ( .A1(npu_inst_int_data_res_5__0__2_), .A2(
        npu_inst_pe_1_4_0_n1), .B1(npu_inst_pe_1_4_0_N75), .B2(
        npu_inst_pe_1_4_0_n76), .C1(npu_inst_pe_1_4_0_N67), .C2(
        npu_inst_pe_1_4_0_n77), .ZN(npu_inst_pe_1_4_0_n82) );
  INV_X1 npu_inst_pe_1_4_0_U44 ( .A(npu_inst_pe_1_4_0_n82), .ZN(
        npu_inst_pe_1_4_0_n99) );
  AOI222_X1 npu_inst_pe_1_4_0_U43 ( .A1(npu_inst_int_data_res_5__0__3_), .A2(
        npu_inst_pe_1_4_0_n1), .B1(npu_inst_pe_1_4_0_N76), .B2(
        npu_inst_pe_1_4_0_n76), .C1(npu_inst_pe_1_4_0_N68), .C2(
        npu_inst_pe_1_4_0_n77), .ZN(npu_inst_pe_1_4_0_n81) );
  INV_X1 npu_inst_pe_1_4_0_U42 ( .A(npu_inst_pe_1_4_0_n81), .ZN(
        npu_inst_pe_1_4_0_n98) );
  AOI222_X1 npu_inst_pe_1_4_0_U41 ( .A1(npu_inst_int_data_res_5__0__4_), .A2(
        npu_inst_pe_1_4_0_n1), .B1(npu_inst_pe_1_4_0_N77), .B2(
        npu_inst_pe_1_4_0_n76), .C1(npu_inst_pe_1_4_0_N69), .C2(
        npu_inst_pe_1_4_0_n77), .ZN(npu_inst_pe_1_4_0_n80) );
  INV_X1 npu_inst_pe_1_4_0_U40 ( .A(npu_inst_pe_1_4_0_n80), .ZN(
        npu_inst_pe_1_4_0_n36) );
  AOI222_X1 npu_inst_pe_1_4_0_U39 ( .A1(npu_inst_int_data_res_5__0__5_), .A2(
        npu_inst_pe_1_4_0_n1), .B1(npu_inst_pe_1_4_0_N78), .B2(
        npu_inst_pe_1_4_0_n76), .C1(npu_inst_pe_1_4_0_N70), .C2(
        npu_inst_pe_1_4_0_n77), .ZN(npu_inst_pe_1_4_0_n79) );
  INV_X1 npu_inst_pe_1_4_0_U38 ( .A(npu_inst_pe_1_4_0_n79), .ZN(
        npu_inst_pe_1_4_0_n35) );
  AOI222_X1 npu_inst_pe_1_4_0_U37 ( .A1(npu_inst_int_data_res_5__0__6_), .A2(
        npu_inst_pe_1_4_0_n1), .B1(npu_inst_pe_1_4_0_N79), .B2(
        npu_inst_pe_1_4_0_n76), .C1(npu_inst_pe_1_4_0_N71), .C2(
        npu_inst_pe_1_4_0_n77), .ZN(npu_inst_pe_1_4_0_n78) );
  INV_X1 npu_inst_pe_1_4_0_U36 ( .A(npu_inst_pe_1_4_0_n78), .ZN(
        npu_inst_pe_1_4_0_n34) );
  AND2_X1 npu_inst_pe_1_4_0_U35 ( .A1(npu_inst_pe_1_4_0_o_data_h_1_), .A2(
        npu_inst_pe_1_4_0_int_q_weight_1_), .ZN(npu_inst_pe_1_4_0_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_4_0_U34 ( .A1(npu_inst_pe_1_4_0_o_data_h_0_), .A2(
        npu_inst_pe_1_4_0_int_q_weight_1_), .ZN(npu_inst_pe_1_4_0_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_4_0_U33 ( .A(npu_inst_pe_1_4_0_int_data_1_), .ZN(
        npu_inst_pe_1_4_0_n14) );
  AOI22_X1 npu_inst_pe_1_4_0_U32 ( .A1(npu_inst_n56), .A2(
        npu_inst_int_data_y_5__0__1_), .B1(npu_inst_pe_1_4_0_n3), .B2(
        npu_inst_int_data_x_4__1__1_), .ZN(npu_inst_pe_1_4_0_n63) );
  AOI22_X1 npu_inst_pe_1_4_0_U31 ( .A1(npu_inst_n56), .A2(
        npu_inst_int_data_y_5__0__0_), .B1(npu_inst_pe_1_4_0_n3), .B2(
        npu_inst_int_data_x_4__1__0_), .ZN(npu_inst_pe_1_4_0_n61) );
  INV_X1 npu_inst_pe_1_4_0_U30 ( .A(npu_inst_pe_1_4_0_int_data_0_), .ZN(
        npu_inst_pe_1_4_0_n13) );
  INV_X1 npu_inst_pe_1_4_0_U29 ( .A(npu_inst_n69), .ZN(npu_inst_pe_1_4_0_n5)
         );
  OR3_X1 npu_inst_pe_1_4_0_U28 ( .A1(npu_inst_pe_1_4_0_n6), .A2(
        npu_inst_pe_1_4_0_n8), .A3(npu_inst_pe_1_4_0_n5), .ZN(
        npu_inst_pe_1_4_0_n56) );
  OR3_X1 npu_inst_pe_1_4_0_U27 ( .A1(npu_inst_pe_1_4_0_n5), .A2(
        npu_inst_pe_1_4_0_n8), .A3(npu_inst_pe_1_4_0_n7), .ZN(
        npu_inst_pe_1_4_0_n48) );
  INV_X1 npu_inst_pe_1_4_0_U26 ( .A(npu_inst_pe_1_4_0_n5), .ZN(
        npu_inst_pe_1_4_0_n4) );
  OR3_X1 npu_inst_pe_1_4_0_U25 ( .A1(npu_inst_pe_1_4_0_n4), .A2(
        npu_inst_pe_1_4_0_n8), .A3(npu_inst_pe_1_4_0_n7), .ZN(
        npu_inst_pe_1_4_0_n52) );
  OR3_X1 npu_inst_pe_1_4_0_U24 ( .A1(npu_inst_pe_1_4_0_n6), .A2(
        npu_inst_pe_1_4_0_n8), .A3(npu_inst_pe_1_4_0_n4), .ZN(
        npu_inst_pe_1_4_0_n60) );
  NOR2_X1 npu_inst_pe_1_4_0_U23 ( .A1(npu_inst_pe_1_4_0_n60), .A2(
        npu_inst_pe_1_4_0_n3), .ZN(npu_inst_pe_1_4_0_n58) );
  NOR2_X1 npu_inst_pe_1_4_0_U22 ( .A1(npu_inst_pe_1_4_0_n56), .A2(
        npu_inst_pe_1_4_0_n3), .ZN(npu_inst_pe_1_4_0_n54) );
  NOR2_X1 npu_inst_pe_1_4_0_U21 ( .A1(npu_inst_pe_1_4_0_n52), .A2(
        npu_inst_pe_1_4_0_n3), .ZN(npu_inst_pe_1_4_0_n50) );
  NOR2_X1 npu_inst_pe_1_4_0_U20 ( .A1(npu_inst_pe_1_4_0_n48), .A2(
        npu_inst_pe_1_4_0_n3), .ZN(npu_inst_pe_1_4_0_n46) );
  NOR2_X1 npu_inst_pe_1_4_0_U19 ( .A1(npu_inst_pe_1_4_0_n40), .A2(
        npu_inst_pe_1_4_0_n3), .ZN(npu_inst_pe_1_4_0_n38) );
  NOR2_X1 npu_inst_pe_1_4_0_U18 ( .A1(npu_inst_pe_1_4_0_n44), .A2(
        npu_inst_pe_1_4_0_n3), .ZN(npu_inst_pe_1_4_0_n42) );
  BUF_X1 npu_inst_pe_1_4_0_U17 ( .A(npu_inst_n99), .Z(npu_inst_pe_1_4_0_n8) );
  INV_X1 npu_inst_pe_1_4_0_U16 ( .A(npu_inst_n124), .ZN(npu_inst_pe_1_4_0_n12)
         );
  INV_X1 npu_inst_pe_1_4_0_U15 ( .A(npu_inst_pe_1_4_0_n38), .ZN(
        npu_inst_pe_1_4_0_n114) );
  INV_X1 npu_inst_pe_1_4_0_U14 ( .A(npu_inst_pe_1_4_0_n58), .ZN(
        npu_inst_pe_1_4_0_n119) );
  INV_X1 npu_inst_pe_1_4_0_U13 ( .A(npu_inst_pe_1_4_0_n54), .ZN(
        npu_inst_pe_1_4_0_n118) );
  INV_X1 npu_inst_pe_1_4_0_U12 ( .A(npu_inst_pe_1_4_0_n50), .ZN(
        npu_inst_pe_1_4_0_n117) );
  INV_X1 npu_inst_pe_1_4_0_U11 ( .A(npu_inst_pe_1_4_0_n46), .ZN(
        npu_inst_pe_1_4_0_n116) );
  INV_X1 npu_inst_pe_1_4_0_U10 ( .A(npu_inst_pe_1_4_0_n42), .ZN(
        npu_inst_pe_1_4_0_n115) );
  BUF_X1 npu_inst_pe_1_4_0_U9 ( .A(npu_inst_n22), .Z(npu_inst_pe_1_4_0_n2) );
  BUF_X1 npu_inst_pe_1_4_0_U8 ( .A(npu_inst_n22), .Z(npu_inst_pe_1_4_0_n1) );
  BUF_X1 npu_inst_pe_1_4_0_U7 ( .A(npu_inst_pe_1_4_0_n12), .Z(
        npu_inst_pe_1_4_0_n11) );
  BUF_X1 npu_inst_pe_1_4_0_U6 ( .A(npu_inst_pe_1_4_0_n12), .Z(
        npu_inst_pe_1_4_0_n10) );
  BUF_X1 npu_inst_pe_1_4_0_U5 ( .A(npu_inst_pe_1_4_0_n12), .Z(
        npu_inst_pe_1_4_0_n9) );
  NOR2_X1 npu_inst_pe_1_4_0_U4 ( .A1(npu_inst_pe_1_4_0_int_q_weight_0_), .A2(
        npu_inst_pe_1_4_0_n1), .ZN(npu_inst_pe_1_4_0_n76) );
  NOR2_X1 npu_inst_pe_1_4_0_U3 ( .A1(npu_inst_pe_1_4_0_n27), .A2(
        npu_inst_pe_1_4_0_n1), .ZN(npu_inst_pe_1_4_0_n77) );
  FA_X1 npu_inst_pe_1_4_0_sub_67_U2_1 ( .A(npu_inst_pe_1_4_0_int_q_acc_1_), 
        .B(npu_inst_pe_1_4_0_n14), .CI(npu_inst_pe_1_4_0_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_4_0_sub_67_carry_2_), .S(npu_inst_pe_1_4_0_N66) );
  FA_X1 npu_inst_pe_1_4_0_add_69_U1_1 ( .A(npu_inst_pe_1_4_0_int_q_acc_1_), 
        .B(npu_inst_pe_1_4_0_int_data_1_), .CI(
        npu_inst_pe_1_4_0_add_69_carry_1_), .CO(
        npu_inst_pe_1_4_0_add_69_carry_2_), .S(npu_inst_pe_1_4_0_N74) );
  NAND3_X1 npu_inst_pe_1_4_0_U109 ( .A1(npu_inst_pe_1_4_0_n5), .A2(
        npu_inst_pe_1_4_0_n7), .A3(npu_inst_pe_1_4_0_n8), .ZN(
        npu_inst_pe_1_4_0_n44) );
  NAND3_X1 npu_inst_pe_1_4_0_U108 ( .A1(npu_inst_pe_1_4_0_n4), .A2(
        npu_inst_pe_1_4_0_n7), .A3(npu_inst_pe_1_4_0_n8), .ZN(
        npu_inst_pe_1_4_0_n40) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_4_0_n34), .CK(
        npu_inst_pe_1_4_0_net3826), .RN(npu_inst_pe_1_4_0_n9), .Q(
        npu_inst_pe_1_4_0_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_4_0_n35), .CK(
        npu_inst_pe_1_4_0_net3826), .RN(npu_inst_pe_1_4_0_n9), .Q(
        npu_inst_pe_1_4_0_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_4_0_n36), .CK(
        npu_inst_pe_1_4_0_net3826), .RN(npu_inst_pe_1_4_0_n9), .Q(
        npu_inst_pe_1_4_0_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_4_0_n98), .CK(
        npu_inst_pe_1_4_0_net3826), .RN(npu_inst_pe_1_4_0_n9), .Q(
        npu_inst_pe_1_4_0_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_4_0_n99), .CK(
        npu_inst_pe_1_4_0_net3826), .RN(npu_inst_pe_1_4_0_n9), .Q(
        npu_inst_pe_1_4_0_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_4_0_n100), 
        .CK(npu_inst_pe_1_4_0_net3826), .RN(npu_inst_pe_1_4_0_n9), .Q(
        npu_inst_pe_1_4_0_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_4_0_n33), .CK(
        npu_inst_pe_1_4_0_net3826), .RN(npu_inst_pe_1_4_0_n9), .Q(
        npu_inst_pe_1_4_0_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_4_0_n101), 
        .CK(npu_inst_pe_1_4_0_net3826), .RN(npu_inst_pe_1_4_0_n9), .Q(
        npu_inst_pe_1_4_0_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_weight_reg_0_ ( .D(npu_inst_n110), .CK(
        npu_inst_pe_1_4_0_net3832), .RN(npu_inst_pe_1_4_0_n9), .Q(
        npu_inst_pe_1_4_0_int_q_weight_0_), .QN(npu_inst_pe_1_4_0_n27) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_weight_reg_1_ ( .D(npu_inst_n116), .CK(
        npu_inst_pe_1_4_0_net3832), .RN(npu_inst_pe_1_4_0_n9), .Q(
        npu_inst_pe_1_4_0_int_q_weight_1_), .QN(npu_inst_pe_1_4_0_n26) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_4_0_n113), 
        .CK(npu_inst_pe_1_4_0_net3832), .RN(npu_inst_pe_1_4_0_n9), .Q(
        npu_inst_pe_1_4_0_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_4_0_n107), 
        .CK(npu_inst_pe_1_4_0_net3832), .RN(npu_inst_pe_1_4_0_n9), .Q(
        npu_inst_pe_1_4_0_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_4_0_n112), 
        .CK(npu_inst_pe_1_4_0_net3832), .RN(npu_inst_pe_1_4_0_n10), .Q(
        npu_inst_pe_1_4_0_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_4_0_n106), 
        .CK(npu_inst_pe_1_4_0_net3832), .RN(npu_inst_pe_1_4_0_n10), .Q(
        npu_inst_pe_1_4_0_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_4_0_n111), 
        .CK(npu_inst_pe_1_4_0_net3832), .RN(npu_inst_pe_1_4_0_n10), .Q(
        npu_inst_pe_1_4_0_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_4_0_n105), 
        .CK(npu_inst_pe_1_4_0_net3832), .RN(npu_inst_pe_1_4_0_n10), .Q(
        npu_inst_pe_1_4_0_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_4_0_n110), 
        .CK(npu_inst_pe_1_4_0_net3832), .RN(npu_inst_pe_1_4_0_n10), .Q(
        npu_inst_pe_1_4_0_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_4_0_n104), 
        .CK(npu_inst_pe_1_4_0_net3832), .RN(npu_inst_pe_1_4_0_n10), .Q(
        npu_inst_pe_1_4_0_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_4_0_n109), 
        .CK(npu_inst_pe_1_4_0_net3832), .RN(npu_inst_pe_1_4_0_n10), .Q(
        npu_inst_pe_1_4_0_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_4_0_n103), 
        .CK(npu_inst_pe_1_4_0_net3832), .RN(npu_inst_pe_1_4_0_n10), .Q(
        npu_inst_pe_1_4_0_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_4_0_n108), 
        .CK(npu_inst_pe_1_4_0_net3832), .RN(npu_inst_pe_1_4_0_n10), .Q(
        npu_inst_pe_1_4_0_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_4_0_n102), 
        .CK(npu_inst_pe_1_4_0_net3832), .RN(npu_inst_pe_1_4_0_n10), .Q(
        npu_inst_pe_1_4_0_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_4_0_n86), 
        .CK(npu_inst_pe_1_4_0_net3832), .RN(npu_inst_pe_1_4_0_n10), .Q(
        npu_inst_pe_1_4_0_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_4_0_n87), 
        .CK(npu_inst_pe_1_4_0_net3832), .RN(npu_inst_pe_1_4_0_n10), .Q(
        npu_inst_pe_1_4_0_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_4_0_n88), 
        .CK(npu_inst_pe_1_4_0_net3832), .RN(npu_inst_pe_1_4_0_n11), .Q(
        npu_inst_pe_1_4_0_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_4_0_n89), 
        .CK(npu_inst_pe_1_4_0_net3832), .RN(npu_inst_pe_1_4_0_n11), .Q(
        npu_inst_pe_1_4_0_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_4_0_n90), 
        .CK(npu_inst_pe_1_4_0_net3832), .RN(npu_inst_pe_1_4_0_n11), .Q(
        npu_inst_pe_1_4_0_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_4_0_n91), 
        .CK(npu_inst_pe_1_4_0_net3832), .RN(npu_inst_pe_1_4_0_n11), .Q(
        npu_inst_pe_1_4_0_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_4_0_n92), 
        .CK(npu_inst_pe_1_4_0_net3832), .RN(npu_inst_pe_1_4_0_n11), .Q(
        npu_inst_pe_1_4_0_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_4_0_n93), 
        .CK(npu_inst_pe_1_4_0_net3832), .RN(npu_inst_pe_1_4_0_n11), .Q(
        npu_inst_pe_1_4_0_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_4_0_n94), 
        .CK(npu_inst_pe_1_4_0_net3832), .RN(npu_inst_pe_1_4_0_n11), .Q(
        npu_inst_pe_1_4_0_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_4_0_n95), 
        .CK(npu_inst_pe_1_4_0_net3832), .RN(npu_inst_pe_1_4_0_n11), .Q(
        npu_inst_pe_1_4_0_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_4_0_n96), 
        .CK(npu_inst_pe_1_4_0_net3832), .RN(npu_inst_pe_1_4_0_n11), .Q(
        npu_inst_pe_1_4_0_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_4_0_n97), 
        .CK(npu_inst_pe_1_4_0_net3832), .RN(npu_inst_pe_1_4_0_n11), .Q(
        npu_inst_pe_1_4_0_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_4_0_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_4_0_N84), .SE(1'b0), .GCK(npu_inst_pe_1_4_0_net3826) );
  CLKGATETST_X1 npu_inst_pe_1_4_0_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n63), .SE(1'b0), .GCK(npu_inst_pe_1_4_0_net3832) );
  MUX2_X1 npu_inst_pe_1_4_1_U162 ( .A(npu_inst_pe_1_4_1_n32), .B(
        npu_inst_pe_1_4_1_n29), .S(npu_inst_pe_1_4_1_n8), .Z(
        npu_inst_pe_1_4_1_N93) );
  MUX2_X1 npu_inst_pe_1_4_1_U161 ( .A(npu_inst_pe_1_4_1_n31), .B(
        npu_inst_pe_1_4_1_n30), .S(npu_inst_pe_1_4_1_n6), .Z(
        npu_inst_pe_1_4_1_n32) );
  MUX2_X1 npu_inst_pe_1_4_1_U160 ( .A(npu_inst_pe_1_4_1_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_4_1_int_q_reg_v_1__0_), .S(npu_inst_pe_1_4_1_n4), .Z(
        npu_inst_pe_1_4_1_n31) );
  MUX2_X1 npu_inst_pe_1_4_1_U159 ( .A(npu_inst_pe_1_4_1_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_4_1_int_q_reg_v_3__0_), .S(npu_inst_pe_1_4_1_n4), .Z(
        npu_inst_pe_1_4_1_n30) );
  MUX2_X1 npu_inst_pe_1_4_1_U158 ( .A(npu_inst_pe_1_4_1_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_4_1_int_q_reg_v_5__0_), .S(npu_inst_pe_1_4_1_n4), .Z(
        npu_inst_pe_1_4_1_n29) );
  MUX2_X1 npu_inst_pe_1_4_1_U157 ( .A(npu_inst_pe_1_4_1_n28), .B(
        npu_inst_pe_1_4_1_n23), .S(npu_inst_pe_1_4_1_n8), .Z(
        npu_inst_pe_1_4_1_N94) );
  MUX2_X1 npu_inst_pe_1_4_1_U156 ( .A(npu_inst_pe_1_4_1_n25), .B(
        npu_inst_pe_1_4_1_n24), .S(npu_inst_pe_1_4_1_n6), .Z(
        npu_inst_pe_1_4_1_n28) );
  MUX2_X1 npu_inst_pe_1_4_1_U155 ( .A(npu_inst_pe_1_4_1_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_4_1_int_q_reg_v_1__1_), .S(npu_inst_pe_1_4_1_n4), .Z(
        npu_inst_pe_1_4_1_n25) );
  MUX2_X1 npu_inst_pe_1_4_1_U154 ( .A(npu_inst_pe_1_4_1_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_4_1_int_q_reg_v_3__1_), .S(npu_inst_pe_1_4_1_n4), .Z(
        npu_inst_pe_1_4_1_n24) );
  MUX2_X1 npu_inst_pe_1_4_1_U153 ( .A(npu_inst_pe_1_4_1_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_4_1_int_q_reg_v_5__1_), .S(npu_inst_pe_1_4_1_n4), .Z(
        npu_inst_pe_1_4_1_n23) );
  MUX2_X1 npu_inst_pe_1_4_1_U152 ( .A(npu_inst_pe_1_4_1_n22), .B(
        npu_inst_pe_1_4_1_n19), .S(npu_inst_pe_1_4_1_n8), .Z(
        npu_inst_int_data_x_4__1__1_) );
  MUX2_X1 npu_inst_pe_1_4_1_U151 ( .A(npu_inst_pe_1_4_1_n21), .B(
        npu_inst_pe_1_4_1_n20), .S(npu_inst_pe_1_4_1_n6), .Z(
        npu_inst_pe_1_4_1_n22) );
  MUX2_X1 npu_inst_pe_1_4_1_U150 ( .A(npu_inst_pe_1_4_1_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_4_1_int_q_reg_h_1__1_), .S(npu_inst_pe_1_4_1_n4), .Z(
        npu_inst_pe_1_4_1_n21) );
  MUX2_X1 npu_inst_pe_1_4_1_U149 ( .A(npu_inst_pe_1_4_1_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_4_1_int_q_reg_h_3__1_), .S(npu_inst_pe_1_4_1_n4), .Z(
        npu_inst_pe_1_4_1_n20) );
  MUX2_X1 npu_inst_pe_1_4_1_U148 ( .A(npu_inst_pe_1_4_1_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_4_1_int_q_reg_h_5__1_), .S(npu_inst_pe_1_4_1_n4), .Z(
        npu_inst_pe_1_4_1_n19) );
  MUX2_X1 npu_inst_pe_1_4_1_U147 ( .A(npu_inst_pe_1_4_1_n18), .B(
        npu_inst_pe_1_4_1_n15), .S(npu_inst_pe_1_4_1_n8), .Z(
        npu_inst_int_data_x_4__1__0_) );
  MUX2_X1 npu_inst_pe_1_4_1_U146 ( .A(npu_inst_pe_1_4_1_n17), .B(
        npu_inst_pe_1_4_1_n16), .S(npu_inst_pe_1_4_1_n6), .Z(
        npu_inst_pe_1_4_1_n18) );
  MUX2_X1 npu_inst_pe_1_4_1_U145 ( .A(npu_inst_pe_1_4_1_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_4_1_int_q_reg_h_1__0_), .S(npu_inst_pe_1_4_1_n4), .Z(
        npu_inst_pe_1_4_1_n17) );
  MUX2_X1 npu_inst_pe_1_4_1_U144 ( .A(npu_inst_pe_1_4_1_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_4_1_int_q_reg_h_3__0_), .S(npu_inst_pe_1_4_1_n4), .Z(
        npu_inst_pe_1_4_1_n16) );
  MUX2_X1 npu_inst_pe_1_4_1_U143 ( .A(npu_inst_pe_1_4_1_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_4_1_int_q_reg_h_5__0_), .S(npu_inst_pe_1_4_1_n4), .Z(
        npu_inst_pe_1_4_1_n15) );
  XOR2_X1 npu_inst_pe_1_4_1_U142 ( .A(npu_inst_pe_1_4_1_int_data_0_), .B(
        npu_inst_pe_1_4_1_int_q_acc_0_), .Z(npu_inst_pe_1_4_1_N73) );
  AND2_X1 npu_inst_pe_1_4_1_U141 ( .A1(npu_inst_pe_1_4_1_int_q_acc_0_), .A2(
        npu_inst_pe_1_4_1_int_data_0_), .ZN(npu_inst_pe_1_4_1_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_4_1_U140 ( .A(npu_inst_pe_1_4_1_int_q_acc_0_), .B(
        npu_inst_pe_1_4_1_n13), .ZN(npu_inst_pe_1_4_1_N65) );
  OR2_X1 npu_inst_pe_1_4_1_U139 ( .A1(npu_inst_pe_1_4_1_n13), .A2(
        npu_inst_pe_1_4_1_int_q_acc_0_), .ZN(npu_inst_pe_1_4_1_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_4_1_U138 ( .A(npu_inst_pe_1_4_1_int_q_acc_2_), .B(
        npu_inst_pe_1_4_1_add_69_carry_2_), .Z(npu_inst_pe_1_4_1_N75) );
  AND2_X1 npu_inst_pe_1_4_1_U137 ( .A1(npu_inst_pe_1_4_1_add_69_carry_2_), 
        .A2(npu_inst_pe_1_4_1_int_q_acc_2_), .ZN(
        npu_inst_pe_1_4_1_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_4_1_U136 ( .A(npu_inst_pe_1_4_1_int_q_acc_3_), .B(
        npu_inst_pe_1_4_1_add_69_carry_3_), .Z(npu_inst_pe_1_4_1_N76) );
  AND2_X1 npu_inst_pe_1_4_1_U135 ( .A1(npu_inst_pe_1_4_1_add_69_carry_3_), 
        .A2(npu_inst_pe_1_4_1_int_q_acc_3_), .ZN(
        npu_inst_pe_1_4_1_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_4_1_U134 ( .A(npu_inst_pe_1_4_1_int_q_acc_4_), .B(
        npu_inst_pe_1_4_1_add_69_carry_4_), .Z(npu_inst_pe_1_4_1_N77) );
  AND2_X1 npu_inst_pe_1_4_1_U133 ( .A1(npu_inst_pe_1_4_1_add_69_carry_4_), 
        .A2(npu_inst_pe_1_4_1_int_q_acc_4_), .ZN(
        npu_inst_pe_1_4_1_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_4_1_U132 ( .A(npu_inst_pe_1_4_1_int_q_acc_5_), .B(
        npu_inst_pe_1_4_1_add_69_carry_5_), .Z(npu_inst_pe_1_4_1_N78) );
  AND2_X1 npu_inst_pe_1_4_1_U131 ( .A1(npu_inst_pe_1_4_1_add_69_carry_5_), 
        .A2(npu_inst_pe_1_4_1_int_q_acc_5_), .ZN(
        npu_inst_pe_1_4_1_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_4_1_U130 ( .A(npu_inst_pe_1_4_1_int_q_acc_6_), .B(
        npu_inst_pe_1_4_1_add_69_carry_6_), .Z(npu_inst_pe_1_4_1_N79) );
  AND2_X1 npu_inst_pe_1_4_1_U129 ( .A1(npu_inst_pe_1_4_1_add_69_carry_6_), 
        .A2(npu_inst_pe_1_4_1_int_q_acc_6_), .ZN(
        npu_inst_pe_1_4_1_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_4_1_U128 ( .A(npu_inst_pe_1_4_1_int_q_acc_7_), .B(
        npu_inst_pe_1_4_1_add_69_carry_7_), .Z(npu_inst_pe_1_4_1_N80) );
  XNOR2_X1 npu_inst_pe_1_4_1_U127 ( .A(npu_inst_pe_1_4_1_sub_67_carry_2_), .B(
        npu_inst_pe_1_4_1_int_q_acc_2_), .ZN(npu_inst_pe_1_4_1_N67) );
  OR2_X1 npu_inst_pe_1_4_1_U126 ( .A1(npu_inst_pe_1_4_1_int_q_acc_2_), .A2(
        npu_inst_pe_1_4_1_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_4_1_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_4_1_U125 ( .A(npu_inst_pe_1_4_1_sub_67_carry_3_), .B(
        npu_inst_pe_1_4_1_int_q_acc_3_), .ZN(npu_inst_pe_1_4_1_N68) );
  OR2_X1 npu_inst_pe_1_4_1_U124 ( .A1(npu_inst_pe_1_4_1_int_q_acc_3_), .A2(
        npu_inst_pe_1_4_1_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_4_1_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_4_1_U123 ( .A(npu_inst_pe_1_4_1_sub_67_carry_4_), .B(
        npu_inst_pe_1_4_1_int_q_acc_4_), .ZN(npu_inst_pe_1_4_1_N69) );
  OR2_X1 npu_inst_pe_1_4_1_U122 ( .A1(npu_inst_pe_1_4_1_int_q_acc_4_), .A2(
        npu_inst_pe_1_4_1_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_4_1_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_4_1_U121 ( .A(npu_inst_pe_1_4_1_sub_67_carry_5_), .B(
        npu_inst_pe_1_4_1_int_q_acc_5_), .ZN(npu_inst_pe_1_4_1_N70) );
  OR2_X1 npu_inst_pe_1_4_1_U120 ( .A1(npu_inst_pe_1_4_1_int_q_acc_5_), .A2(
        npu_inst_pe_1_4_1_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_4_1_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_4_1_U119 ( .A(npu_inst_pe_1_4_1_sub_67_carry_6_), .B(
        npu_inst_pe_1_4_1_int_q_acc_6_), .ZN(npu_inst_pe_1_4_1_N71) );
  OR2_X1 npu_inst_pe_1_4_1_U118 ( .A1(npu_inst_pe_1_4_1_int_q_acc_6_), .A2(
        npu_inst_pe_1_4_1_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_4_1_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_4_1_U117 ( .A(npu_inst_pe_1_4_1_int_q_acc_7_), .B(
        npu_inst_pe_1_4_1_sub_67_carry_7_), .ZN(npu_inst_pe_1_4_1_N72) );
  INV_X1 npu_inst_pe_1_4_1_U116 ( .A(npu_inst_n77), .ZN(npu_inst_pe_1_4_1_n7)
         );
  INV_X1 npu_inst_pe_1_4_1_U115 ( .A(npu_inst_pe_1_4_1_n7), .ZN(
        npu_inst_pe_1_4_1_n6) );
  INV_X1 npu_inst_pe_1_4_1_U114 ( .A(npu_inst_n56), .ZN(npu_inst_pe_1_4_1_n3)
         );
  AOI22_X1 npu_inst_pe_1_4_1_U113 ( .A1(npu_inst_int_data_y_5__1__0_), .A2(
        npu_inst_pe_1_4_1_n58), .B1(npu_inst_pe_1_4_1_n119), .B2(
        npu_inst_pe_1_4_1_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_4_1_n57) );
  INV_X1 npu_inst_pe_1_4_1_U112 ( .A(npu_inst_pe_1_4_1_n57), .ZN(
        npu_inst_pe_1_4_1_n108) );
  AOI22_X1 npu_inst_pe_1_4_1_U111 ( .A1(npu_inst_int_data_y_5__1__0_), .A2(
        npu_inst_pe_1_4_1_n54), .B1(npu_inst_pe_1_4_1_n118), .B2(
        npu_inst_pe_1_4_1_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_4_1_n53) );
  INV_X1 npu_inst_pe_1_4_1_U110 ( .A(npu_inst_pe_1_4_1_n53), .ZN(
        npu_inst_pe_1_4_1_n109) );
  AOI22_X1 npu_inst_pe_1_4_1_U107 ( .A1(npu_inst_int_data_y_5__1__0_), .A2(
        npu_inst_pe_1_4_1_n50), .B1(npu_inst_pe_1_4_1_n117), .B2(
        npu_inst_pe_1_4_1_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_4_1_n49) );
  INV_X1 npu_inst_pe_1_4_1_U106 ( .A(npu_inst_pe_1_4_1_n49), .ZN(
        npu_inst_pe_1_4_1_n110) );
  AOI22_X1 npu_inst_pe_1_4_1_U105 ( .A1(npu_inst_int_data_y_5__1__0_), .A2(
        npu_inst_pe_1_4_1_n46), .B1(npu_inst_pe_1_4_1_n116), .B2(
        npu_inst_pe_1_4_1_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_4_1_n45) );
  INV_X1 npu_inst_pe_1_4_1_U104 ( .A(npu_inst_pe_1_4_1_n45), .ZN(
        npu_inst_pe_1_4_1_n111) );
  AOI22_X1 npu_inst_pe_1_4_1_U103 ( .A1(npu_inst_int_data_y_5__1__0_), .A2(
        npu_inst_pe_1_4_1_n42), .B1(npu_inst_pe_1_4_1_n115), .B2(
        npu_inst_pe_1_4_1_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_4_1_n41) );
  INV_X1 npu_inst_pe_1_4_1_U102 ( .A(npu_inst_pe_1_4_1_n41), .ZN(
        npu_inst_pe_1_4_1_n112) );
  AOI22_X1 npu_inst_pe_1_4_1_U101 ( .A1(npu_inst_int_data_y_5__1__1_), .A2(
        npu_inst_pe_1_4_1_n58), .B1(npu_inst_pe_1_4_1_n119), .B2(
        npu_inst_pe_1_4_1_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_4_1_n59) );
  INV_X1 npu_inst_pe_1_4_1_U100 ( .A(npu_inst_pe_1_4_1_n59), .ZN(
        npu_inst_pe_1_4_1_n102) );
  AOI22_X1 npu_inst_pe_1_4_1_U99 ( .A1(npu_inst_int_data_y_5__1__1_), .A2(
        npu_inst_pe_1_4_1_n54), .B1(npu_inst_pe_1_4_1_n118), .B2(
        npu_inst_pe_1_4_1_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_4_1_n55) );
  INV_X1 npu_inst_pe_1_4_1_U98 ( .A(npu_inst_pe_1_4_1_n55), .ZN(
        npu_inst_pe_1_4_1_n103) );
  AOI22_X1 npu_inst_pe_1_4_1_U97 ( .A1(npu_inst_int_data_y_5__1__1_), .A2(
        npu_inst_pe_1_4_1_n50), .B1(npu_inst_pe_1_4_1_n117), .B2(
        npu_inst_pe_1_4_1_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_4_1_n51) );
  INV_X1 npu_inst_pe_1_4_1_U96 ( .A(npu_inst_pe_1_4_1_n51), .ZN(
        npu_inst_pe_1_4_1_n104) );
  AOI22_X1 npu_inst_pe_1_4_1_U95 ( .A1(npu_inst_int_data_y_5__1__1_), .A2(
        npu_inst_pe_1_4_1_n46), .B1(npu_inst_pe_1_4_1_n116), .B2(
        npu_inst_pe_1_4_1_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_4_1_n47) );
  INV_X1 npu_inst_pe_1_4_1_U94 ( .A(npu_inst_pe_1_4_1_n47), .ZN(
        npu_inst_pe_1_4_1_n105) );
  AOI22_X1 npu_inst_pe_1_4_1_U93 ( .A1(npu_inst_int_data_y_5__1__1_), .A2(
        npu_inst_pe_1_4_1_n42), .B1(npu_inst_pe_1_4_1_n115), .B2(
        npu_inst_pe_1_4_1_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_4_1_n43) );
  INV_X1 npu_inst_pe_1_4_1_U92 ( .A(npu_inst_pe_1_4_1_n43), .ZN(
        npu_inst_pe_1_4_1_n106) );
  AOI22_X1 npu_inst_pe_1_4_1_U91 ( .A1(npu_inst_pe_1_4_1_n38), .A2(
        npu_inst_int_data_y_5__1__1_), .B1(npu_inst_pe_1_4_1_n114), .B2(
        npu_inst_pe_1_4_1_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_4_1_n39) );
  INV_X1 npu_inst_pe_1_4_1_U90 ( .A(npu_inst_pe_1_4_1_n39), .ZN(
        npu_inst_pe_1_4_1_n107) );
  AOI22_X1 npu_inst_pe_1_4_1_U89 ( .A1(npu_inst_pe_1_4_1_n38), .A2(
        npu_inst_int_data_y_5__1__0_), .B1(npu_inst_pe_1_4_1_n114), .B2(
        npu_inst_pe_1_4_1_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_4_1_n37) );
  INV_X1 npu_inst_pe_1_4_1_U88 ( .A(npu_inst_pe_1_4_1_n37), .ZN(
        npu_inst_pe_1_4_1_n113) );
  NAND2_X1 npu_inst_pe_1_4_1_U87 ( .A1(npu_inst_pe_1_4_1_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_4_1_n60), .ZN(npu_inst_pe_1_4_1_n74) );
  OAI21_X1 npu_inst_pe_1_4_1_U86 ( .B1(npu_inst_pe_1_4_1_n63), .B2(
        npu_inst_pe_1_4_1_n60), .A(npu_inst_pe_1_4_1_n74), .ZN(
        npu_inst_pe_1_4_1_n97) );
  NAND2_X1 npu_inst_pe_1_4_1_U85 ( .A1(npu_inst_pe_1_4_1_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_4_1_n60), .ZN(npu_inst_pe_1_4_1_n73) );
  OAI21_X1 npu_inst_pe_1_4_1_U84 ( .B1(npu_inst_pe_1_4_1_n61), .B2(
        npu_inst_pe_1_4_1_n60), .A(npu_inst_pe_1_4_1_n73), .ZN(
        npu_inst_pe_1_4_1_n96) );
  NAND2_X1 npu_inst_pe_1_4_1_U83 ( .A1(npu_inst_pe_1_4_1_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_4_1_n56), .ZN(npu_inst_pe_1_4_1_n72) );
  OAI21_X1 npu_inst_pe_1_4_1_U82 ( .B1(npu_inst_pe_1_4_1_n63), .B2(
        npu_inst_pe_1_4_1_n56), .A(npu_inst_pe_1_4_1_n72), .ZN(
        npu_inst_pe_1_4_1_n95) );
  NAND2_X1 npu_inst_pe_1_4_1_U81 ( .A1(npu_inst_pe_1_4_1_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_4_1_n56), .ZN(npu_inst_pe_1_4_1_n71) );
  OAI21_X1 npu_inst_pe_1_4_1_U80 ( .B1(npu_inst_pe_1_4_1_n61), .B2(
        npu_inst_pe_1_4_1_n56), .A(npu_inst_pe_1_4_1_n71), .ZN(
        npu_inst_pe_1_4_1_n94) );
  NAND2_X1 npu_inst_pe_1_4_1_U79 ( .A1(npu_inst_pe_1_4_1_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_4_1_n52), .ZN(npu_inst_pe_1_4_1_n70) );
  OAI21_X1 npu_inst_pe_1_4_1_U78 ( .B1(npu_inst_pe_1_4_1_n63), .B2(
        npu_inst_pe_1_4_1_n52), .A(npu_inst_pe_1_4_1_n70), .ZN(
        npu_inst_pe_1_4_1_n93) );
  NAND2_X1 npu_inst_pe_1_4_1_U77 ( .A1(npu_inst_pe_1_4_1_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_4_1_n52), .ZN(npu_inst_pe_1_4_1_n69) );
  OAI21_X1 npu_inst_pe_1_4_1_U76 ( .B1(npu_inst_pe_1_4_1_n61), .B2(
        npu_inst_pe_1_4_1_n52), .A(npu_inst_pe_1_4_1_n69), .ZN(
        npu_inst_pe_1_4_1_n92) );
  NAND2_X1 npu_inst_pe_1_4_1_U75 ( .A1(npu_inst_pe_1_4_1_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_4_1_n48), .ZN(npu_inst_pe_1_4_1_n68) );
  OAI21_X1 npu_inst_pe_1_4_1_U74 ( .B1(npu_inst_pe_1_4_1_n63), .B2(
        npu_inst_pe_1_4_1_n48), .A(npu_inst_pe_1_4_1_n68), .ZN(
        npu_inst_pe_1_4_1_n91) );
  NAND2_X1 npu_inst_pe_1_4_1_U73 ( .A1(npu_inst_pe_1_4_1_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_4_1_n48), .ZN(npu_inst_pe_1_4_1_n67) );
  OAI21_X1 npu_inst_pe_1_4_1_U72 ( .B1(npu_inst_pe_1_4_1_n61), .B2(
        npu_inst_pe_1_4_1_n48), .A(npu_inst_pe_1_4_1_n67), .ZN(
        npu_inst_pe_1_4_1_n90) );
  NAND2_X1 npu_inst_pe_1_4_1_U71 ( .A1(npu_inst_pe_1_4_1_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_4_1_n44), .ZN(npu_inst_pe_1_4_1_n66) );
  OAI21_X1 npu_inst_pe_1_4_1_U70 ( .B1(npu_inst_pe_1_4_1_n63), .B2(
        npu_inst_pe_1_4_1_n44), .A(npu_inst_pe_1_4_1_n66), .ZN(
        npu_inst_pe_1_4_1_n89) );
  NAND2_X1 npu_inst_pe_1_4_1_U69 ( .A1(npu_inst_pe_1_4_1_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_4_1_n44), .ZN(npu_inst_pe_1_4_1_n65) );
  OAI21_X1 npu_inst_pe_1_4_1_U68 ( .B1(npu_inst_pe_1_4_1_n61), .B2(
        npu_inst_pe_1_4_1_n44), .A(npu_inst_pe_1_4_1_n65), .ZN(
        npu_inst_pe_1_4_1_n88) );
  NAND2_X1 npu_inst_pe_1_4_1_U67 ( .A1(npu_inst_pe_1_4_1_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_4_1_n40), .ZN(npu_inst_pe_1_4_1_n64) );
  OAI21_X1 npu_inst_pe_1_4_1_U66 ( .B1(npu_inst_pe_1_4_1_n63), .B2(
        npu_inst_pe_1_4_1_n40), .A(npu_inst_pe_1_4_1_n64), .ZN(
        npu_inst_pe_1_4_1_n87) );
  NAND2_X1 npu_inst_pe_1_4_1_U65 ( .A1(npu_inst_pe_1_4_1_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_4_1_n40), .ZN(npu_inst_pe_1_4_1_n62) );
  OAI21_X1 npu_inst_pe_1_4_1_U64 ( .B1(npu_inst_pe_1_4_1_n61), .B2(
        npu_inst_pe_1_4_1_n40), .A(npu_inst_pe_1_4_1_n62), .ZN(
        npu_inst_pe_1_4_1_n86) );
  AND2_X1 npu_inst_pe_1_4_1_U63 ( .A1(npu_inst_pe_1_4_1_N93), .A2(npu_inst_n56), .ZN(npu_inst_int_data_y_4__1__0_) );
  AND2_X1 npu_inst_pe_1_4_1_U62 ( .A1(npu_inst_n56), .A2(npu_inst_pe_1_4_1_N94), .ZN(npu_inst_int_data_y_4__1__1_) );
  NOR3_X1 npu_inst_pe_1_4_1_U61 ( .A1(npu_inst_pe_1_4_1_n26), .A2(npu_inst_n56), .A3(npu_inst_int_ckg[30]), .ZN(npu_inst_pe_1_4_1_n85) );
  OR2_X1 npu_inst_pe_1_4_1_U60 ( .A1(npu_inst_pe_1_4_1_n85), .A2(
        npu_inst_pe_1_4_1_n2), .ZN(npu_inst_pe_1_4_1_N84) );
  AND2_X1 npu_inst_pe_1_4_1_U59 ( .A1(npu_inst_pe_1_4_1_int_q_acc_0_), .A2(
        npu_inst_pe_1_4_1_n1), .ZN(npu_inst_int_data_res_4__1__0_) );
  AND2_X1 npu_inst_pe_1_4_1_U58 ( .A1(npu_inst_pe_1_4_1_n2), .A2(
        npu_inst_pe_1_4_1_int_q_acc_7_), .ZN(npu_inst_int_data_res_4__1__7_)
         );
  AND2_X1 npu_inst_pe_1_4_1_U57 ( .A1(npu_inst_pe_1_4_1_int_q_acc_1_), .A2(
        npu_inst_pe_1_4_1_n1), .ZN(npu_inst_int_data_res_4__1__1_) );
  AND2_X1 npu_inst_pe_1_4_1_U56 ( .A1(npu_inst_pe_1_4_1_int_q_acc_2_), .A2(
        npu_inst_pe_1_4_1_n1), .ZN(npu_inst_int_data_res_4__1__2_) );
  AND2_X1 npu_inst_pe_1_4_1_U55 ( .A1(npu_inst_pe_1_4_1_int_q_acc_3_), .A2(
        npu_inst_pe_1_4_1_n2), .ZN(npu_inst_int_data_res_4__1__3_) );
  AND2_X1 npu_inst_pe_1_4_1_U54 ( .A1(npu_inst_pe_1_4_1_int_q_acc_4_), .A2(
        npu_inst_pe_1_4_1_n2), .ZN(npu_inst_int_data_res_4__1__4_) );
  AND2_X1 npu_inst_pe_1_4_1_U53 ( .A1(npu_inst_pe_1_4_1_int_q_acc_5_), .A2(
        npu_inst_pe_1_4_1_n2), .ZN(npu_inst_int_data_res_4__1__5_) );
  AND2_X1 npu_inst_pe_1_4_1_U52 ( .A1(npu_inst_pe_1_4_1_int_q_acc_6_), .A2(
        npu_inst_pe_1_4_1_n2), .ZN(npu_inst_int_data_res_4__1__6_) );
  AOI222_X1 npu_inst_pe_1_4_1_U51 ( .A1(npu_inst_int_data_res_5__1__0_), .A2(
        npu_inst_pe_1_4_1_n1), .B1(npu_inst_pe_1_4_1_N73), .B2(
        npu_inst_pe_1_4_1_n76), .C1(npu_inst_pe_1_4_1_N65), .C2(
        npu_inst_pe_1_4_1_n77), .ZN(npu_inst_pe_1_4_1_n84) );
  INV_X1 npu_inst_pe_1_4_1_U50 ( .A(npu_inst_pe_1_4_1_n84), .ZN(
        npu_inst_pe_1_4_1_n101) );
  AOI222_X1 npu_inst_pe_1_4_1_U49 ( .A1(npu_inst_int_data_res_5__1__7_), .A2(
        npu_inst_pe_1_4_1_n1), .B1(npu_inst_pe_1_4_1_N80), .B2(
        npu_inst_pe_1_4_1_n76), .C1(npu_inst_pe_1_4_1_N72), .C2(
        npu_inst_pe_1_4_1_n77), .ZN(npu_inst_pe_1_4_1_n75) );
  INV_X1 npu_inst_pe_1_4_1_U48 ( .A(npu_inst_pe_1_4_1_n75), .ZN(
        npu_inst_pe_1_4_1_n33) );
  AOI222_X1 npu_inst_pe_1_4_1_U47 ( .A1(npu_inst_int_data_res_5__1__1_), .A2(
        npu_inst_pe_1_4_1_n1), .B1(npu_inst_pe_1_4_1_N74), .B2(
        npu_inst_pe_1_4_1_n76), .C1(npu_inst_pe_1_4_1_N66), .C2(
        npu_inst_pe_1_4_1_n77), .ZN(npu_inst_pe_1_4_1_n83) );
  INV_X1 npu_inst_pe_1_4_1_U46 ( .A(npu_inst_pe_1_4_1_n83), .ZN(
        npu_inst_pe_1_4_1_n100) );
  AOI222_X1 npu_inst_pe_1_4_1_U45 ( .A1(npu_inst_int_data_res_5__1__2_), .A2(
        npu_inst_pe_1_4_1_n1), .B1(npu_inst_pe_1_4_1_N75), .B2(
        npu_inst_pe_1_4_1_n76), .C1(npu_inst_pe_1_4_1_N67), .C2(
        npu_inst_pe_1_4_1_n77), .ZN(npu_inst_pe_1_4_1_n82) );
  INV_X1 npu_inst_pe_1_4_1_U44 ( .A(npu_inst_pe_1_4_1_n82), .ZN(
        npu_inst_pe_1_4_1_n99) );
  AOI222_X1 npu_inst_pe_1_4_1_U43 ( .A1(npu_inst_int_data_res_5__1__3_), .A2(
        npu_inst_pe_1_4_1_n1), .B1(npu_inst_pe_1_4_1_N76), .B2(
        npu_inst_pe_1_4_1_n76), .C1(npu_inst_pe_1_4_1_N68), .C2(
        npu_inst_pe_1_4_1_n77), .ZN(npu_inst_pe_1_4_1_n81) );
  INV_X1 npu_inst_pe_1_4_1_U42 ( .A(npu_inst_pe_1_4_1_n81), .ZN(
        npu_inst_pe_1_4_1_n98) );
  AOI222_X1 npu_inst_pe_1_4_1_U41 ( .A1(npu_inst_int_data_res_5__1__4_), .A2(
        npu_inst_pe_1_4_1_n1), .B1(npu_inst_pe_1_4_1_N77), .B2(
        npu_inst_pe_1_4_1_n76), .C1(npu_inst_pe_1_4_1_N69), .C2(
        npu_inst_pe_1_4_1_n77), .ZN(npu_inst_pe_1_4_1_n80) );
  INV_X1 npu_inst_pe_1_4_1_U40 ( .A(npu_inst_pe_1_4_1_n80), .ZN(
        npu_inst_pe_1_4_1_n36) );
  AOI222_X1 npu_inst_pe_1_4_1_U39 ( .A1(npu_inst_int_data_res_5__1__5_), .A2(
        npu_inst_pe_1_4_1_n1), .B1(npu_inst_pe_1_4_1_N78), .B2(
        npu_inst_pe_1_4_1_n76), .C1(npu_inst_pe_1_4_1_N70), .C2(
        npu_inst_pe_1_4_1_n77), .ZN(npu_inst_pe_1_4_1_n79) );
  INV_X1 npu_inst_pe_1_4_1_U38 ( .A(npu_inst_pe_1_4_1_n79), .ZN(
        npu_inst_pe_1_4_1_n35) );
  AOI222_X1 npu_inst_pe_1_4_1_U37 ( .A1(npu_inst_int_data_res_5__1__6_), .A2(
        npu_inst_pe_1_4_1_n1), .B1(npu_inst_pe_1_4_1_N79), .B2(
        npu_inst_pe_1_4_1_n76), .C1(npu_inst_pe_1_4_1_N71), .C2(
        npu_inst_pe_1_4_1_n77), .ZN(npu_inst_pe_1_4_1_n78) );
  INV_X1 npu_inst_pe_1_4_1_U36 ( .A(npu_inst_pe_1_4_1_n78), .ZN(
        npu_inst_pe_1_4_1_n34) );
  INV_X1 npu_inst_pe_1_4_1_U35 ( .A(npu_inst_pe_1_4_1_int_data_1_), .ZN(
        npu_inst_pe_1_4_1_n14) );
  AND2_X1 npu_inst_pe_1_4_1_U34 ( .A1(npu_inst_int_data_x_4__1__1_), .A2(
        npu_inst_pe_1_4_1_int_q_weight_1_), .ZN(npu_inst_pe_1_4_1_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_4_1_U33 ( .A1(npu_inst_int_data_x_4__1__0_), .A2(
        npu_inst_pe_1_4_1_int_q_weight_1_), .ZN(npu_inst_pe_1_4_1_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_4_1_U32 ( .A1(npu_inst_n56), .A2(
        npu_inst_int_data_y_5__1__1_), .B1(npu_inst_pe_1_4_1_n3), .B2(
        npu_inst_int_data_x_4__2__1_), .ZN(npu_inst_pe_1_4_1_n63) );
  AOI22_X1 npu_inst_pe_1_4_1_U31 ( .A1(npu_inst_n56), .A2(
        npu_inst_int_data_y_5__1__0_), .B1(npu_inst_pe_1_4_1_n3), .B2(
        npu_inst_int_data_x_4__2__0_), .ZN(npu_inst_pe_1_4_1_n61) );
  INV_X1 npu_inst_pe_1_4_1_U30 ( .A(npu_inst_pe_1_4_1_int_data_0_), .ZN(
        npu_inst_pe_1_4_1_n13) );
  INV_X1 npu_inst_pe_1_4_1_U29 ( .A(npu_inst_n69), .ZN(npu_inst_pe_1_4_1_n5)
         );
  OR3_X1 npu_inst_pe_1_4_1_U28 ( .A1(npu_inst_pe_1_4_1_n6), .A2(
        npu_inst_pe_1_4_1_n8), .A3(npu_inst_pe_1_4_1_n5), .ZN(
        npu_inst_pe_1_4_1_n56) );
  OR3_X1 npu_inst_pe_1_4_1_U27 ( .A1(npu_inst_pe_1_4_1_n5), .A2(
        npu_inst_pe_1_4_1_n8), .A3(npu_inst_pe_1_4_1_n7), .ZN(
        npu_inst_pe_1_4_1_n48) );
  INV_X1 npu_inst_pe_1_4_1_U26 ( .A(npu_inst_pe_1_4_1_n5), .ZN(
        npu_inst_pe_1_4_1_n4) );
  OR3_X1 npu_inst_pe_1_4_1_U25 ( .A1(npu_inst_pe_1_4_1_n4), .A2(
        npu_inst_pe_1_4_1_n8), .A3(npu_inst_pe_1_4_1_n7), .ZN(
        npu_inst_pe_1_4_1_n52) );
  OR3_X1 npu_inst_pe_1_4_1_U24 ( .A1(npu_inst_pe_1_4_1_n6), .A2(
        npu_inst_pe_1_4_1_n8), .A3(npu_inst_pe_1_4_1_n4), .ZN(
        npu_inst_pe_1_4_1_n60) );
  NOR2_X1 npu_inst_pe_1_4_1_U23 ( .A1(npu_inst_pe_1_4_1_n60), .A2(
        npu_inst_pe_1_4_1_n3), .ZN(npu_inst_pe_1_4_1_n58) );
  NOR2_X1 npu_inst_pe_1_4_1_U22 ( .A1(npu_inst_pe_1_4_1_n56), .A2(
        npu_inst_pe_1_4_1_n3), .ZN(npu_inst_pe_1_4_1_n54) );
  NOR2_X1 npu_inst_pe_1_4_1_U21 ( .A1(npu_inst_pe_1_4_1_n52), .A2(
        npu_inst_pe_1_4_1_n3), .ZN(npu_inst_pe_1_4_1_n50) );
  NOR2_X1 npu_inst_pe_1_4_1_U20 ( .A1(npu_inst_pe_1_4_1_n48), .A2(
        npu_inst_pe_1_4_1_n3), .ZN(npu_inst_pe_1_4_1_n46) );
  NOR2_X1 npu_inst_pe_1_4_1_U19 ( .A1(npu_inst_pe_1_4_1_n40), .A2(
        npu_inst_pe_1_4_1_n3), .ZN(npu_inst_pe_1_4_1_n38) );
  NOR2_X1 npu_inst_pe_1_4_1_U18 ( .A1(npu_inst_pe_1_4_1_n44), .A2(
        npu_inst_pe_1_4_1_n3), .ZN(npu_inst_pe_1_4_1_n42) );
  BUF_X1 npu_inst_pe_1_4_1_U17 ( .A(npu_inst_n99), .Z(npu_inst_pe_1_4_1_n8) );
  INV_X1 npu_inst_pe_1_4_1_U16 ( .A(npu_inst_n124), .ZN(npu_inst_pe_1_4_1_n12)
         );
  INV_X1 npu_inst_pe_1_4_1_U15 ( .A(npu_inst_pe_1_4_1_n38), .ZN(
        npu_inst_pe_1_4_1_n114) );
  INV_X1 npu_inst_pe_1_4_1_U14 ( .A(npu_inst_pe_1_4_1_n58), .ZN(
        npu_inst_pe_1_4_1_n119) );
  INV_X1 npu_inst_pe_1_4_1_U13 ( .A(npu_inst_pe_1_4_1_n54), .ZN(
        npu_inst_pe_1_4_1_n118) );
  INV_X1 npu_inst_pe_1_4_1_U12 ( .A(npu_inst_pe_1_4_1_n50), .ZN(
        npu_inst_pe_1_4_1_n117) );
  INV_X1 npu_inst_pe_1_4_1_U11 ( .A(npu_inst_pe_1_4_1_n46), .ZN(
        npu_inst_pe_1_4_1_n116) );
  INV_X1 npu_inst_pe_1_4_1_U10 ( .A(npu_inst_pe_1_4_1_n42), .ZN(
        npu_inst_pe_1_4_1_n115) );
  BUF_X1 npu_inst_pe_1_4_1_U9 ( .A(npu_inst_n22), .Z(npu_inst_pe_1_4_1_n2) );
  BUF_X1 npu_inst_pe_1_4_1_U8 ( .A(npu_inst_n22), .Z(npu_inst_pe_1_4_1_n1) );
  BUF_X1 npu_inst_pe_1_4_1_U7 ( .A(npu_inst_pe_1_4_1_n12), .Z(
        npu_inst_pe_1_4_1_n11) );
  BUF_X1 npu_inst_pe_1_4_1_U6 ( .A(npu_inst_pe_1_4_1_n12), .Z(
        npu_inst_pe_1_4_1_n10) );
  BUF_X1 npu_inst_pe_1_4_1_U5 ( .A(npu_inst_pe_1_4_1_n12), .Z(
        npu_inst_pe_1_4_1_n9) );
  NOR2_X1 npu_inst_pe_1_4_1_U4 ( .A1(npu_inst_pe_1_4_1_int_q_weight_0_), .A2(
        npu_inst_pe_1_4_1_n1), .ZN(npu_inst_pe_1_4_1_n76) );
  NOR2_X1 npu_inst_pe_1_4_1_U3 ( .A1(npu_inst_pe_1_4_1_n27), .A2(
        npu_inst_pe_1_4_1_n1), .ZN(npu_inst_pe_1_4_1_n77) );
  FA_X1 npu_inst_pe_1_4_1_sub_67_U2_1 ( .A(npu_inst_pe_1_4_1_int_q_acc_1_), 
        .B(npu_inst_pe_1_4_1_n14), .CI(npu_inst_pe_1_4_1_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_4_1_sub_67_carry_2_), .S(npu_inst_pe_1_4_1_N66) );
  FA_X1 npu_inst_pe_1_4_1_add_69_U1_1 ( .A(npu_inst_pe_1_4_1_int_q_acc_1_), 
        .B(npu_inst_pe_1_4_1_int_data_1_), .CI(
        npu_inst_pe_1_4_1_add_69_carry_1_), .CO(
        npu_inst_pe_1_4_1_add_69_carry_2_), .S(npu_inst_pe_1_4_1_N74) );
  NAND3_X1 npu_inst_pe_1_4_1_U109 ( .A1(npu_inst_pe_1_4_1_n5), .A2(
        npu_inst_pe_1_4_1_n7), .A3(npu_inst_pe_1_4_1_n8), .ZN(
        npu_inst_pe_1_4_1_n44) );
  NAND3_X1 npu_inst_pe_1_4_1_U108 ( .A1(npu_inst_pe_1_4_1_n4), .A2(
        npu_inst_pe_1_4_1_n7), .A3(npu_inst_pe_1_4_1_n8), .ZN(
        npu_inst_pe_1_4_1_n40) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_4_1_n34), .CK(
        npu_inst_pe_1_4_1_net3803), .RN(npu_inst_pe_1_4_1_n9), .Q(
        npu_inst_pe_1_4_1_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_4_1_n35), .CK(
        npu_inst_pe_1_4_1_net3803), .RN(npu_inst_pe_1_4_1_n9), .Q(
        npu_inst_pe_1_4_1_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_4_1_n36), .CK(
        npu_inst_pe_1_4_1_net3803), .RN(npu_inst_pe_1_4_1_n9), .Q(
        npu_inst_pe_1_4_1_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_4_1_n98), .CK(
        npu_inst_pe_1_4_1_net3803), .RN(npu_inst_pe_1_4_1_n9), .Q(
        npu_inst_pe_1_4_1_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_4_1_n99), .CK(
        npu_inst_pe_1_4_1_net3803), .RN(npu_inst_pe_1_4_1_n9), .Q(
        npu_inst_pe_1_4_1_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_4_1_n100), 
        .CK(npu_inst_pe_1_4_1_net3803), .RN(npu_inst_pe_1_4_1_n9), .Q(
        npu_inst_pe_1_4_1_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_4_1_n33), .CK(
        npu_inst_pe_1_4_1_net3803), .RN(npu_inst_pe_1_4_1_n9), .Q(
        npu_inst_pe_1_4_1_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_4_1_n101), 
        .CK(npu_inst_pe_1_4_1_net3803), .RN(npu_inst_pe_1_4_1_n9), .Q(
        npu_inst_pe_1_4_1_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_weight_reg_0_ ( .D(npu_inst_n110), .CK(
        npu_inst_pe_1_4_1_net3809), .RN(npu_inst_pe_1_4_1_n9), .Q(
        npu_inst_pe_1_4_1_int_q_weight_0_), .QN(npu_inst_pe_1_4_1_n27) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_weight_reg_1_ ( .D(npu_inst_n116), .CK(
        npu_inst_pe_1_4_1_net3809), .RN(npu_inst_pe_1_4_1_n9), .Q(
        npu_inst_pe_1_4_1_int_q_weight_1_), .QN(npu_inst_pe_1_4_1_n26) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_4_1_n113), 
        .CK(npu_inst_pe_1_4_1_net3809), .RN(npu_inst_pe_1_4_1_n9), .Q(
        npu_inst_pe_1_4_1_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_4_1_n107), 
        .CK(npu_inst_pe_1_4_1_net3809), .RN(npu_inst_pe_1_4_1_n9), .Q(
        npu_inst_pe_1_4_1_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_4_1_n112), 
        .CK(npu_inst_pe_1_4_1_net3809), .RN(npu_inst_pe_1_4_1_n10), .Q(
        npu_inst_pe_1_4_1_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_4_1_n106), 
        .CK(npu_inst_pe_1_4_1_net3809), .RN(npu_inst_pe_1_4_1_n10), .Q(
        npu_inst_pe_1_4_1_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_4_1_n111), 
        .CK(npu_inst_pe_1_4_1_net3809), .RN(npu_inst_pe_1_4_1_n10), .Q(
        npu_inst_pe_1_4_1_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_4_1_n105), 
        .CK(npu_inst_pe_1_4_1_net3809), .RN(npu_inst_pe_1_4_1_n10), .Q(
        npu_inst_pe_1_4_1_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_4_1_n110), 
        .CK(npu_inst_pe_1_4_1_net3809), .RN(npu_inst_pe_1_4_1_n10), .Q(
        npu_inst_pe_1_4_1_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_4_1_n104), 
        .CK(npu_inst_pe_1_4_1_net3809), .RN(npu_inst_pe_1_4_1_n10), .Q(
        npu_inst_pe_1_4_1_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_4_1_n109), 
        .CK(npu_inst_pe_1_4_1_net3809), .RN(npu_inst_pe_1_4_1_n10), .Q(
        npu_inst_pe_1_4_1_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_4_1_n103), 
        .CK(npu_inst_pe_1_4_1_net3809), .RN(npu_inst_pe_1_4_1_n10), .Q(
        npu_inst_pe_1_4_1_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_4_1_n108), 
        .CK(npu_inst_pe_1_4_1_net3809), .RN(npu_inst_pe_1_4_1_n10), .Q(
        npu_inst_pe_1_4_1_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_4_1_n102), 
        .CK(npu_inst_pe_1_4_1_net3809), .RN(npu_inst_pe_1_4_1_n10), .Q(
        npu_inst_pe_1_4_1_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_4_1_n86), 
        .CK(npu_inst_pe_1_4_1_net3809), .RN(npu_inst_pe_1_4_1_n10), .Q(
        npu_inst_pe_1_4_1_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_4_1_n87), 
        .CK(npu_inst_pe_1_4_1_net3809), .RN(npu_inst_pe_1_4_1_n10), .Q(
        npu_inst_pe_1_4_1_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_4_1_n88), 
        .CK(npu_inst_pe_1_4_1_net3809), .RN(npu_inst_pe_1_4_1_n11), .Q(
        npu_inst_pe_1_4_1_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_4_1_n89), 
        .CK(npu_inst_pe_1_4_1_net3809), .RN(npu_inst_pe_1_4_1_n11), .Q(
        npu_inst_pe_1_4_1_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_4_1_n90), 
        .CK(npu_inst_pe_1_4_1_net3809), .RN(npu_inst_pe_1_4_1_n11), .Q(
        npu_inst_pe_1_4_1_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_4_1_n91), 
        .CK(npu_inst_pe_1_4_1_net3809), .RN(npu_inst_pe_1_4_1_n11), .Q(
        npu_inst_pe_1_4_1_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_4_1_n92), 
        .CK(npu_inst_pe_1_4_1_net3809), .RN(npu_inst_pe_1_4_1_n11), .Q(
        npu_inst_pe_1_4_1_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_4_1_n93), 
        .CK(npu_inst_pe_1_4_1_net3809), .RN(npu_inst_pe_1_4_1_n11), .Q(
        npu_inst_pe_1_4_1_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_4_1_n94), 
        .CK(npu_inst_pe_1_4_1_net3809), .RN(npu_inst_pe_1_4_1_n11), .Q(
        npu_inst_pe_1_4_1_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_4_1_n95), 
        .CK(npu_inst_pe_1_4_1_net3809), .RN(npu_inst_pe_1_4_1_n11), .Q(
        npu_inst_pe_1_4_1_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_4_1_n96), 
        .CK(npu_inst_pe_1_4_1_net3809), .RN(npu_inst_pe_1_4_1_n11), .Q(
        npu_inst_pe_1_4_1_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_4_1_n97), 
        .CK(npu_inst_pe_1_4_1_net3809), .RN(npu_inst_pe_1_4_1_n11), .Q(
        npu_inst_pe_1_4_1_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_4_1_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_4_1_N84), .SE(1'b0), .GCK(npu_inst_pe_1_4_1_net3803) );
  CLKGATETST_X1 npu_inst_pe_1_4_1_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n63), .SE(1'b0), .GCK(npu_inst_pe_1_4_1_net3809) );
  MUX2_X1 npu_inst_pe_1_4_2_U162 ( .A(npu_inst_pe_1_4_2_n32), .B(
        npu_inst_pe_1_4_2_n29), .S(npu_inst_pe_1_4_2_n8), .Z(
        npu_inst_pe_1_4_2_N93) );
  MUX2_X1 npu_inst_pe_1_4_2_U161 ( .A(npu_inst_pe_1_4_2_n31), .B(
        npu_inst_pe_1_4_2_n30), .S(npu_inst_pe_1_4_2_n6), .Z(
        npu_inst_pe_1_4_2_n32) );
  MUX2_X1 npu_inst_pe_1_4_2_U160 ( .A(npu_inst_pe_1_4_2_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_4_2_int_q_reg_v_1__0_), .S(npu_inst_pe_1_4_2_n4), .Z(
        npu_inst_pe_1_4_2_n31) );
  MUX2_X1 npu_inst_pe_1_4_2_U159 ( .A(npu_inst_pe_1_4_2_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_4_2_int_q_reg_v_3__0_), .S(npu_inst_pe_1_4_2_n4), .Z(
        npu_inst_pe_1_4_2_n30) );
  MUX2_X1 npu_inst_pe_1_4_2_U158 ( .A(npu_inst_pe_1_4_2_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_4_2_int_q_reg_v_5__0_), .S(npu_inst_pe_1_4_2_n4), .Z(
        npu_inst_pe_1_4_2_n29) );
  MUX2_X1 npu_inst_pe_1_4_2_U157 ( .A(npu_inst_pe_1_4_2_n28), .B(
        npu_inst_pe_1_4_2_n23), .S(npu_inst_pe_1_4_2_n8), .Z(
        npu_inst_pe_1_4_2_N94) );
  MUX2_X1 npu_inst_pe_1_4_2_U156 ( .A(npu_inst_pe_1_4_2_n25), .B(
        npu_inst_pe_1_4_2_n24), .S(npu_inst_pe_1_4_2_n6), .Z(
        npu_inst_pe_1_4_2_n28) );
  MUX2_X1 npu_inst_pe_1_4_2_U155 ( .A(npu_inst_pe_1_4_2_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_4_2_int_q_reg_v_1__1_), .S(npu_inst_pe_1_4_2_n4), .Z(
        npu_inst_pe_1_4_2_n25) );
  MUX2_X1 npu_inst_pe_1_4_2_U154 ( .A(npu_inst_pe_1_4_2_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_4_2_int_q_reg_v_3__1_), .S(npu_inst_pe_1_4_2_n4), .Z(
        npu_inst_pe_1_4_2_n24) );
  MUX2_X1 npu_inst_pe_1_4_2_U153 ( .A(npu_inst_pe_1_4_2_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_4_2_int_q_reg_v_5__1_), .S(npu_inst_pe_1_4_2_n4), .Z(
        npu_inst_pe_1_4_2_n23) );
  MUX2_X1 npu_inst_pe_1_4_2_U152 ( .A(npu_inst_pe_1_4_2_n22), .B(
        npu_inst_pe_1_4_2_n19), .S(npu_inst_pe_1_4_2_n8), .Z(
        npu_inst_int_data_x_4__2__1_) );
  MUX2_X1 npu_inst_pe_1_4_2_U151 ( .A(npu_inst_pe_1_4_2_n21), .B(
        npu_inst_pe_1_4_2_n20), .S(npu_inst_pe_1_4_2_n6), .Z(
        npu_inst_pe_1_4_2_n22) );
  MUX2_X1 npu_inst_pe_1_4_2_U150 ( .A(npu_inst_pe_1_4_2_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_4_2_int_q_reg_h_1__1_), .S(npu_inst_pe_1_4_2_n4), .Z(
        npu_inst_pe_1_4_2_n21) );
  MUX2_X1 npu_inst_pe_1_4_2_U149 ( .A(npu_inst_pe_1_4_2_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_4_2_int_q_reg_h_3__1_), .S(npu_inst_pe_1_4_2_n4), .Z(
        npu_inst_pe_1_4_2_n20) );
  MUX2_X1 npu_inst_pe_1_4_2_U148 ( .A(npu_inst_pe_1_4_2_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_4_2_int_q_reg_h_5__1_), .S(npu_inst_pe_1_4_2_n4), .Z(
        npu_inst_pe_1_4_2_n19) );
  MUX2_X1 npu_inst_pe_1_4_2_U147 ( .A(npu_inst_pe_1_4_2_n18), .B(
        npu_inst_pe_1_4_2_n15), .S(npu_inst_pe_1_4_2_n8), .Z(
        npu_inst_int_data_x_4__2__0_) );
  MUX2_X1 npu_inst_pe_1_4_2_U146 ( .A(npu_inst_pe_1_4_2_n17), .B(
        npu_inst_pe_1_4_2_n16), .S(npu_inst_pe_1_4_2_n6), .Z(
        npu_inst_pe_1_4_2_n18) );
  MUX2_X1 npu_inst_pe_1_4_2_U145 ( .A(npu_inst_pe_1_4_2_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_4_2_int_q_reg_h_1__0_), .S(npu_inst_pe_1_4_2_n4), .Z(
        npu_inst_pe_1_4_2_n17) );
  MUX2_X1 npu_inst_pe_1_4_2_U144 ( .A(npu_inst_pe_1_4_2_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_4_2_int_q_reg_h_3__0_), .S(npu_inst_pe_1_4_2_n4), .Z(
        npu_inst_pe_1_4_2_n16) );
  MUX2_X1 npu_inst_pe_1_4_2_U143 ( .A(npu_inst_pe_1_4_2_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_4_2_int_q_reg_h_5__0_), .S(npu_inst_pe_1_4_2_n4), .Z(
        npu_inst_pe_1_4_2_n15) );
  XOR2_X1 npu_inst_pe_1_4_2_U142 ( .A(npu_inst_pe_1_4_2_int_data_0_), .B(
        npu_inst_pe_1_4_2_int_q_acc_0_), .Z(npu_inst_pe_1_4_2_N73) );
  AND2_X1 npu_inst_pe_1_4_2_U141 ( .A1(npu_inst_pe_1_4_2_int_q_acc_0_), .A2(
        npu_inst_pe_1_4_2_int_data_0_), .ZN(npu_inst_pe_1_4_2_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_4_2_U140 ( .A(npu_inst_pe_1_4_2_int_q_acc_0_), .B(
        npu_inst_pe_1_4_2_n13), .ZN(npu_inst_pe_1_4_2_N65) );
  OR2_X1 npu_inst_pe_1_4_2_U139 ( .A1(npu_inst_pe_1_4_2_n13), .A2(
        npu_inst_pe_1_4_2_int_q_acc_0_), .ZN(npu_inst_pe_1_4_2_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_4_2_U138 ( .A(npu_inst_pe_1_4_2_int_q_acc_2_), .B(
        npu_inst_pe_1_4_2_add_69_carry_2_), .Z(npu_inst_pe_1_4_2_N75) );
  AND2_X1 npu_inst_pe_1_4_2_U137 ( .A1(npu_inst_pe_1_4_2_add_69_carry_2_), 
        .A2(npu_inst_pe_1_4_2_int_q_acc_2_), .ZN(
        npu_inst_pe_1_4_2_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_4_2_U136 ( .A(npu_inst_pe_1_4_2_int_q_acc_3_), .B(
        npu_inst_pe_1_4_2_add_69_carry_3_), .Z(npu_inst_pe_1_4_2_N76) );
  AND2_X1 npu_inst_pe_1_4_2_U135 ( .A1(npu_inst_pe_1_4_2_add_69_carry_3_), 
        .A2(npu_inst_pe_1_4_2_int_q_acc_3_), .ZN(
        npu_inst_pe_1_4_2_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_4_2_U134 ( .A(npu_inst_pe_1_4_2_int_q_acc_4_), .B(
        npu_inst_pe_1_4_2_add_69_carry_4_), .Z(npu_inst_pe_1_4_2_N77) );
  AND2_X1 npu_inst_pe_1_4_2_U133 ( .A1(npu_inst_pe_1_4_2_add_69_carry_4_), 
        .A2(npu_inst_pe_1_4_2_int_q_acc_4_), .ZN(
        npu_inst_pe_1_4_2_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_4_2_U132 ( .A(npu_inst_pe_1_4_2_int_q_acc_5_), .B(
        npu_inst_pe_1_4_2_add_69_carry_5_), .Z(npu_inst_pe_1_4_2_N78) );
  AND2_X1 npu_inst_pe_1_4_2_U131 ( .A1(npu_inst_pe_1_4_2_add_69_carry_5_), 
        .A2(npu_inst_pe_1_4_2_int_q_acc_5_), .ZN(
        npu_inst_pe_1_4_2_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_4_2_U130 ( .A(npu_inst_pe_1_4_2_int_q_acc_6_), .B(
        npu_inst_pe_1_4_2_add_69_carry_6_), .Z(npu_inst_pe_1_4_2_N79) );
  AND2_X1 npu_inst_pe_1_4_2_U129 ( .A1(npu_inst_pe_1_4_2_add_69_carry_6_), 
        .A2(npu_inst_pe_1_4_2_int_q_acc_6_), .ZN(
        npu_inst_pe_1_4_2_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_4_2_U128 ( .A(npu_inst_pe_1_4_2_int_q_acc_7_), .B(
        npu_inst_pe_1_4_2_add_69_carry_7_), .Z(npu_inst_pe_1_4_2_N80) );
  XNOR2_X1 npu_inst_pe_1_4_2_U127 ( .A(npu_inst_pe_1_4_2_sub_67_carry_2_), .B(
        npu_inst_pe_1_4_2_int_q_acc_2_), .ZN(npu_inst_pe_1_4_2_N67) );
  OR2_X1 npu_inst_pe_1_4_2_U126 ( .A1(npu_inst_pe_1_4_2_int_q_acc_2_), .A2(
        npu_inst_pe_1_4_2_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_4_2_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_4_2_U125 ( .A(npu_inst_pe_1_4_2_sub_67_carry_3_), .B(
        npu_inst_pe_1_4_2_int_q_acc_3_), .ZN(npu_inst_pe_1_4_2_N68) );
  OR2_X1 npu_inst_pe_1_4_2_U124 ( .A1(npu_inst_pe_1_4_2_int_q_acc_3_), .A2(
        npu_inst_pe_1_4_2_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_4_2_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_4_2_U123 ( .A(npu_inst_pe_1_4_2_sub_67_carry_4_), .B(
        npu_inst_pe_1_4_2_int_q_acc_4_), .ZN(npu_inst_pe_1_4_2_N69) );
  OR2_X1 npu_inst_pe_1_4_2_U122 ( .A1(npu_inst_pe_1_4_2_int_q_acc_4_), .A2(
        npu_inst_pe_1_4_2_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_4_2_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_4_2_U121 ( .A(npu_inst_pe_1_4_2_sub_67_carry_5_), .B(
        npu_inst_pe_1_4_2_int_q_acc_5_), .ZN(npu_inst_pe_1_4_2_N70) );
  OR2_X1 npu_inst_pe_1_4_2_U120 ( .A1(npu_inst_pe_1_4_2_int_q_acc_5_), .A2(
        npu_inst_pe_1_4_2_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_4_2_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_4_2_U119 ( .A(npu_inst_pe_1_4_2_sub_67_carry_6_), .B(
        npu_inst_pe_1_4_2_int_q_acc_6_), .ZN(npu_inst_pe_1_4_2_N71) );
  OR2_X1 npu_inst_pe_1_4_2_U118 ( .A1(npu_inst_pe_1_4_2_int_q_acc_6_), .A2(
        npu_inst_pe_1_4_2_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_4_2_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_4_2_U117 ( .A(npu_inst_pe_1_4_2_int_q_acc_7_), .B(
        npu_inst_pe_1_4_2_sub_67_carry_7_), .ZN(npu_inst_pe_1_4_2_N72) );
  INV_X1 npu_inst_pe_1_4_2_U116 ( .A(npu_inst_n77), .ZN(npu_inst_pe_1_4_2_n7)
         );
  INV_X1 npu_inst_pe_1_4_2_U115 ( .A(npu_inst_pe_1_4_2_n7), .ZN(
        npu_inst_pe_1_4_2_n6) );
  INV_X1 npu_inst_pe_1_4_2_U114 ( .A(npu_inst_n56), .ZN(npu_inst_pe_1_4_2_n3)
         );
  AOI22_X1 npu_inst_pe_1_4_2_U113 ( .A1(npu_inst_int_data_y_5__2__0_), .A2(
        npu_inst_pe_1_4_2_n58), .B1(npu_inst_pe_1_4_2_n119), .B2(
        npu_inst_pe_1_4_2_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_4_2_n57) );
  INV_X1 npu_inst_pe_1_4_2_U112 ( .A(npu_inst_pe_1_4_2_n57), .ZN(
        npu_inst_pe_1_4_2_n108) );
  AOI22_X1 npu_inst_pe_1_4_2_U111 ( .A1(npu_inst_int_data_y_5__2__0_), .A2(
        npu_inst_pe_1_4_2_n54), .B1(npu_inst_pe_1_4_2_n118), .B2(
        npu_inst_pe_1_4_2_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_4_2_n53) );
  INV_X1 npu_inst_pe_1_4_2_U110 ( .A(npu_inst_pe_1_4_2_n53), .ZN(
        npu_inst_pe_1_4_2_n109) );
  AOI22_X1 npu_inst_pe_1_4_2_U107 ( .A1(npu_inst_int_data_y_5__2__0_), .A2(
        npu_inst_pe_1_4_2_n50), .B1(npu_inst_pe_1_4_2_n117), .B2(
        npu_inst_pe_1_4_2_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_4_2_n49) );
  INV_X1 npu_inst_pe_1_4_2_U106 ( .A(npu_inst_pe_1_4_2_n49), .ZN(
        npu_inst_pe_1_4_2_n110) );
  AOI22_X1 npu_inst_pe_1_4_2_U105 ( .A1(npu_inst_int_data_y_5__2__0_), .A2(
        npu_inst_pe_1_4_2_n46), .B1(npu_inst_pe_1_4_2_n116), .B2(
        npu_inst_pe_1_4_2_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_4_2_n45) );
  INV_X1 npu_inst_pe_1_4_2_U104 ( .A(npu_inst_pe_1_4_2_n45), .ZN(
        npu_inst_pe_1_4_2_n111) );
  AOI22_X1 npu_inst_pe_1_4_2_U103 ( .A1(npu_inst_int_data_y_5__2__0_), .A2(
        npu_inst_pe_1_4_2_n42), .B1(npu_inst_pe_1_4_2_n115), .B2(
        npu_inst_pe_1_4_2_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_4_2_n41) );
  INV_X1 npu_inst_pe_1_4_2_U102 ( .A(npu_inst_pe_1_4_2_n41), .ZN(
        npu_inst_pe_1_4_2_n112) );
  AOI22_X1 npu_inst_pe_1_4_2_U101 ( .A1(npu_inst_int_data_y_5__2__1_), .A2(
        npu_inst_pe_1_4_2_n58), .B1(npu_inst_pe_1_4_2_n119), .B2(
        npu_inst_pe_1_4_2_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_4_2_n59) );
  INV_X1 npu_inst_pe_1_4_2_U100 ( .A(npu_inst_pe_1_4_2_n59), .ZN(
        npu_inst_pe_1_4_2_n102) );
  AOI22_X1 npu_inst_pe_1_4_2_U99 ( .A1(npu_inst_int_data_y_5__2__1_), .A2(
        npu_inst_pe_1_4_2_n54), .B1(npu_inst_pe_1_4_2_n118), .B2(
        npu_inst_pe_1_4_2_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_4_2_n55) );
  INV_X1 npu_inst_pe_1_4_2_U98 ( .A(npu_inst_pe_1_4_2_n55), .ZN(
        npu_inst_pe_1_4_2_n103) );
  AOI22_X1 npu_inst_pe_1_4_2_U97 ( .A1(npu_inst_int_data_y_5__2__1_), .A2(
        npu_inst_pe_1_4_2_n50), .B1(npu_inst_pe_1_4_2_n117), .B2(
        npu_inst_pe_1_4_2_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_4_2_n51) );
  INV_X1 npu_inst_pe_1_4_2_U96 ( .A(npu_inst_pe_1_4_2_n51), .ZN(
        npu_inst_pe_1_4_2_n104) );
  AOI22_X1 npu_inst_pe_1_4_2_U95 ( .A1(npu_inst_int_data_y_5__2__1_), .A2(
        npu_inst_pe_1_4_2_n46), .B1(npu_inst_pe_1_4_2_n116), .B2(
        npu_inst_pe_1_4_2_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_4_2_n47) );
  INV_X1 npu_inst_pe_1_4_2_U94 ( .A(npu_inst_pe_1_4_2_n47), .ZN(
        npu_inst_pe_1_4_2_n105) );
  AOI22_X1 npu_inst_pe_1_4_2_U93 ( .A1(npu_inst_int_data_y_5__2__1_), .A2(
        npu_inst_pe_1_4_2_n42), .B1(npu_inst_pe_1_4_2_n115), .B2(
        npu_inst_pe_1_4_2_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_4_2_n43) );
  INV_X1 npu_inst_pe_1_4_2_U92 ( .A(npu_inst_pe_1_4_2_n43), .ZN(
        npu_inst_pe_1_4_2_n106) );
  AOI22_X1 npu_inst_pe_1_4_2_U91 ( .A1(npu_inst_pe_1_4_2_n38), .A2(
        npu_inst_int_data_y_5__2__1_), .B1(npu_inst_pe_1_4_2_n114), .B2(
        npu_inst_pe_1_4_2_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_4_2_n39) );
  INV_X1 npu_inst_pe_1_4_2_U90 ( .A(npu_inst_pe_1_4_2_n39), .ZN(
        npu_inst_pe_1_4_2_n107) );
  AOI22_X1 npu_inst_pe_1_4_2_U89 ( .A1(npu_inst_pe_1_4_2_n38), .A2(
        npu_inst_int_data_y_5__2__0_), .B1(npu_inst_pe_1_4_2_n114), .B2(
        npu_inst_pe_1_4_2_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_4_2_n37) );
  INV_X1 npu_inst_pe_1_4_2_U88 ( .A(npu_inst_pe_1_4_2_n37), .ZN(
        npu_inst_pe_1_4_2_n113) );
  NAND2_X1 npu_inst_pe_1_4_2_U87 ( .A1(npu_inst_pe_1_4_2_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_4_2_n60), .ZN(npu_inst_pe_1_4_2_n74) );
  OAI21_X1 npu_inst_pe_1_4_2_U86 ( .B1(npu_inst_pe_1_4_2_n63), .B2(
        npu_inst_pe_1_4_2_n60), .A(npu_inst_pe_1_4_2_n74), .ZN(
        npu_inst_pe_1_4_2_n97) );
  NAND2_X1 npu_inst_pe_1_4_2_U85 ( .A1(npu_inst_pe_1_4_2_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_4_2_n60), .ZN(npu_inst_pe_1_4_2_n73) );
  OAI21_X1 npu_inst_pe_1_4_2_U84 ( .B1(npu_inst_pe_1_4_2_n61), .B2(
        npu_inst_pe_1_4_2_n60), .A(npu_inst_pe_1_4_2_n73), .ZN(
        npu_inst_pe_1_4_2_n96) );
  NAND2_X1 npu_inst_pe_1_4_2_U83 ( .A1(npu_inst_pe_1_4_2_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_4_2_n56), .ZN(npu_inst_pe_1_4_2_n72) );
  OAI21_X1 npu_inst_pe_1_4_2_U82 ( .B1(npu_inst_pe_1_4_2_n63), .B2(
        npu_inst_pe_1_4_2_n56), .A(npu_inst_pe_1_4_2_n72), .ZN(
        npu_inst_pe_1_4_2_n95) );
  NAND2_X1 npu_inst_pe_1_4_2_U81 ( .A1(npu_inst_pe_1_4_2_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_4_2_n56), .ZN(npu_inst_pe_1_4_2_n71) );
  OAI21_X1 npu_inst_pe_1_4_2_U80 ( .B1(npu_inst_pe_1_4_2_n61), .B2(
        npu_inst_pe_1_4_2_n56), .A(npu_inst_pe_1_4_2_n71), .ZN(
        npu_inst_pe_1_4_2_n94) );
  NAND2_X1 npu_inst_pe_1_4_2_U79 ( .A1(npu_inst_pe_1_4_2_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_4_2_n52), .ZN(npu_inst_pe_1_4_2_n70) );
  OAI21_X1 npu_inst_pe_1_4_2_U78 ( .B1(npu_inst_pe_1_4_2_n63), .B2(
        npu_inst_pe_1_4_2_n52), .A(npu_inst_pe_1_4_2_n70), .ZN(
        npu_inst_pe_1_4_2_n93) );
  NAND2_X1 npu_inst_pe_1_4_2_U77 ( .A1(npu_inst_pe_1_4_2_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_4_2_n52), .ZN(npu_inst_pe_1_4_2_n69) );
  OAI21_X1 npu_inst_pe_1_4_2_U76 ( .B1(npu_inst_pe_1_4_2_n61), .B2(
        npu_inst_pe_1_4_2_n52), .A(npu_inst_pe_1_4_2_n69), .ZN(
        npu_inst_pe_1_4_2_n92) );
  NAND2_X1 npu_inst_pe_1_4_2_U75 ( .A1(npu_inst_pe_1_4_2_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_4_2_n48), .ZN(npu_inst_pe_1_4_2_n68) );
  OAI21_X1 npu_inst_pe_1_4_2_U74 ( .B1(npu_inst_pe_1_4_2_n63), .B2(
        npu_inst_pe_1_4_2_n48), .A(npu_inst_pe_1_4_2_n68), .ZN(
        npu_inst_pe_1_4_2_n91) );
  NAND2_X1 npu_inst_pe_1_4_2_U73 ( .A1(npu_inst_pe_1_4_2_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_4_2_n48), .ZN(npu_inst_pe_1_4_2_n67) );
  OAI21_X1 npu_inst_pe_1_4_2_U72 ( .B1(npu_inst_pe_1_4_2_n61), .B2(
        npu_inst_pe_1_4_2_n48), .A(npu_inst_pe_1_4_2_n67), .ZN(
        npu_inst_pe_1_4_2_n90) );
  NAND2_X1 npu_inst_pe_1_4_2_U71 ( .A1(npu_inst_pe_1_4_2_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_4_2_n44), .ZN(npu_inst_pe_1_4_2_n66) );
  OAI21_X1 npu_inst_pe_1_4_2_U70 ( .B1(npu_inst_pe_1_4_2_n63), .B2(
        npu_inst_pe_1_4_2_n44), .A(npu_inst_pe_1_4_2_n66), .ZN(
        npu_inst_pe_1_4_2_n89) );
  NAND2_X1 npu_inst_pe_1_4_2_U69 ( .A1(npu_inst_pe_1_4_2_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_4_2_n44), .ZN(npu_inst_pe_1_4_2_n65) );
  OAI21_X1 npu_inst_pe_1_4_2_U68 ( .B1(npu_inst_pe_1_4_2_n61), .B2(
        npu_inst_pe_1_4_2_n44), .A(npu_inst_pe_1_4_2_n65), .ZN(
        npu_inst_pe_1_4_2_n88) );
  NAND2_X1 npu_inst_pe_1_4_2_U67 ( .A1(npu_inst_pe_1_4_2_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_4_2_n40), .ZN(npu_inst_pe_1_4_2_n64) );
  OAI21_X1 npu_inst_pe_1_4_2_U66 ( .B1(npu_inst_pe_1_4_2_n63), .B2(
        npu_inst_pe_1_4_2_n40), .A(npu_inst_pe_1_4_2_n64), .ZN(
        npu_inst_pe_1_4_2_n87) );
  NAND2_X1 npu_inst_pe_1_4_2_U65 ( .A1(npu_inst_pe_1_4_2_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_4_2_n40), .ZN(npu_inst_pe_1_4_2_n62) );
  OAI21_X1 npu_inst_pe_1_4_2_U64 ( .B1(npu_inst_pe_1_4_2_n61), .B2(
        npu_inst_pe_1_4_2_n40), .A(npu_inst_pe_1_4_2_n62), .ZN(
        npu_inst_pe_1_4_2_n86) );
  AND2_X1 npu_inst_pe_1_4_2_U63 ( .A1(npu_inst_pe_1_4_2_N93), .A2(npu_inst_n56), .ZN(npu_inst_int_data_y_4__2__0_) );
  AND2_X1 npu_inst_pe_1_4_2_U62 ( .A1(npu_inst_n56), .A2(npu_inst_pe_1_4_2_N94), .ZN(npu_inst_int_data_y_4__2__1_) );
  NOR3_X1 npu_inst_pe_1_4_2_U61 ( .A1(npu_inst_pe_1_4_2_n26), .A2(npu_inst_n56), .A3(npu_inst_int_ckg[29]), .ZN(npu_inst_pe_1_4_2_n85) );
  OR2_X1 npu_inst_pe_1_4_2_U60 ( .A1(npu_inst_pe_1_4_2_n85), .A2(
        npu_inst_pe_1_4_2_n2), .ZN(npu_inst_pe_1_4_2_N84) );
  AND2_X1 npu_inst_pe_1_4_2_U59 ( .A1(npu_inst_pe_1_4_2_int_q_acc_0_), .A2(
        npu_inst_pe_1_4_2_n1), .ZN(npu_inst_int_data_res_4__2__0_) );
  AND2_X1 npu_inst_pe_1_4_2_U58 ( .A1(npu_inst_pe_1_4_2_n2), .A2(
        npu_inst_pe_1_4_2_int_q_acc_7_), .ZN(npu_inst_int_data_res_4__2__7_)
         );
  AND2_X1 npu_inst_pe_1_4_2_U57 ( .A1(npu_inst_pe_1_4_2_int_q_acc_1_), .A2(
        npu_inst_pe_1_4_2_n1), .ZN(npu_inst_int_data_res_4__2__1_) );
  AND2_X1 npu_inst_pe_1_4_2_U56 ( .A1(npu_inst_pe_1_4_2_int_q_acc_2_), .A2(
        npu_inst_pe_1_4_2_n1), .ZN(npu_inst_int_data_res_4__2__2_) );
  AND2_X1 npu_inst_pe_1_4_2_U55 ( .A1(npu_inst_pe_1_4_2_int_q_acc_3_), .A2(
        npu_inst_pe_1_4_2_n2), .ZN(npu_inst_int_data_res_4__2__3_) );
  AND2_X1 npu_inst_pe_1_4_2_U54 ( .A1(npu_inst_pe_1_4_2_int_q_acc_4_), .A2(
        npu_inst_pe_1_4_2_n2), .ZN(npu_inst_int_data_res_4__2__4_) );
  AND2_X1 npu_inst_pe_1_4_2_U53 ( .A1(npu_inst_pe_1_4_2_int_q_acc_5_), .A2(
        npu_inst_pe_1_4_2_n2), .ZN(npu_inst_int_data_res_4__2__5_) );
  AND2_X1 npu_inst_pe_1_4_2_U52 ( .A1(npu_inst_pe_1_4_2_int_q_acc_6_), .A2(
        npu_inst_pe_1_4_2_n2), .ZN(npu_inst_int_data_res_4__2__6_) );
  AOI222_X1 npu_inst_pe_1_4_2_U51 ( .A1(npu_inst_int_data_res_5__2__0_), .A2(
        npu_inst_pe_1_4_2_n1), .B1(npu_inst_pe_1_4_2_N73), .B2(
        npu_inst_pe_1_4_2_n76), .C1(npu_inst_pe_1_4_2_N65), .C2(
        npu_inst_pe_1_4_2_n77), .ZN(npu_inst_pe_1_4_2_n84) );
  INV_X1 npu_inst_pe_1_4_2_U50 ( .A(npu_inst_pe_1_4_2_n84), .ZN(
        npu_inst_pe_1_4_2_n101) );
  AOI222_X1 npu_inst_pe_1_4_2_U49 ( .A1(npu_inst_int_data_res_5__2__7_), .A2(
        npu_inst_pe_1_4_2_n1), .B1(npu_inst_pe_1_4_2_N80), .B2(
        npu_inst_pe_1_4_2_n76), .C1(npu_inst_pe_1_4_2_N72), .C2(
        npu_inst_pe_1_4_2_n77), .ZN(npu_inst_pe_1_4_2_n75) );
  INV_X1 npu_inst_pe_1_4_2_U48 ( .A(npu_inst_pe_1_4_2_n75), .ZN(
        npu_inst_pe_1_4_2_n33) );
  AOI222_X1 npu_inst_pe_1_4_2_U47 ( .A1(npu_inst_int_data_res_5__2__1_), .A2(
        npu_inst_pe_1_4_2_n1), .B1(npu_inst_pe_1_4_2_N74), .B2(
        npu_inst_pe_1_4_2_n76), .C1(npu_inst_pe_1_4_2_N66), .C2(
        npu_inst_pe_1_4_2_n77), .ZN(npu_inst_pe_1_4_2_n83) );
  INV_X1 npu_inst_pe_1_4_2_U46 ( .A(npu_inst_pe_1_4_2_n83), .ZN(
        npu_inst_pe_1_4_2_n100) );
  AOI222_X1 npu_inst_pe_1_4_2_U45 ( .A1(npu_inst_int_data_res_5__2__2_), .A2(
        npu_inst_pe_1_4_2_n1), .B1(npu_inst_pe_1_4_2_N75), .B2(
        npu_inst_pe_1_4_2_n76), .C1(npu_inst_pe_1_4_2_N67), .C2(
        npu_inst_pe_1_4_2_n77), .ZN(npu_inst_pe_1_4_2_n82) );
  INV_X1 npu_inst_pe_1_4_2_U44 ( .A(npu_inst_pe_1_4_2_n82), .ZN(
        npu_inst_pe_1_4_2_n99) );
  AOI222_X1 npu_inst_pe_1_4_2_U43 ( .A1(npu_inst_int_data_res_5__2__3_), .A2(
        npu_inst_pe_1_4_2_n1), .B1(npu_inst_pe_1_4_2_N76), .B2(
        npu_inst_pe_1_4_2_n76), .C1(npu_inst_pe_1_4_2_N68), .C2(
        npu_inst_pe_1_4_2_n77), .ZN(npu_inst_pe_1_4_2_n81) );
  INV_X1 npu_inst_pe_1_4_2_U42 ( .A(npu_inst_pe_1_4_2_n81), .ZN(
        npu_inst_pe_1_4_2_n98) );
  AOI222_X1 npu_inst_pe_1_4_2_U41 ( .A1(npu_inst_int_data_res_5__2__4_), .A2(
        npu_inst_pe_1_4_2_n1), .B1(npu_inst_pe_1_4_2_N77), .B2(
        npu_inst_pe_1_4_2_n76), .C1(npu_inst_pe_1_4_2_N69), .C2(
        npu_inst_pe_1_4_2_n77), .ZN(npu_inst_pe_1_4_2_n80) );
  INV_X1 npu_inst_pe_1_4_2_U40 ( .A(npu_inst_pe_1_4_2_n80), .ZN(
        npu_inst_pe_1_4_2_n36) );
  AOI222_X1 npu_inst_pe_1_4_2_U39 ( .A1(npu_inst_int_data_res_5__2__5_), .A2(
        npu_inst_pe_1_4_2_n1), .B1(npu_inst_pe_1_4_2_N78), .B2(
        npu_inst_pe_1_4_2_n76), .C1(npu_inst_pe_1_4_2_N70), .C2(
        npu_inst_pe_1_4_2_n77), .ZN(npu_inst_pe_1_4_2_n79) );
  INV_X1 npu_inst_pe_1_4_2_U38 ( .A(npu_inst_pe_1_4_2_n79), .ZN(
        npu_inst_pe_1_4_2_n35) );
  AOI222_X1 npu_inst_pe_1_4_2_U37 ( .A1(npu_inst_int_data_res_5__2__6_), .A2(
        npu_inst_pe_1_4_2_n1), .B1(npu_inst_pe_1_4_2_N79), .B2(
        npu_inst_pe_1_4_2_n76), .C1(npu_inst_pe_1_4_2_N71), .C2(
        npu_inst_pe_1_4_2_n77), .ZN(npu_inst_pe_1_4_2_n78) );
  INV_X1 npu_inst_pe_1_4_2_U36 ( .A(npu_inst_pe_1_4_2_n78), .ZN(
        npu_inst_pe_1_4_2_n34) );
  INV_X1 npu_inst_pe_1_4_2_U35 ( .A(npu_inst_pe_1_4_2_int_data_1_), .ZN(
        npu_inst_pe_1_4_2_n14) );
  AND2_X1 npu_inst_pe_1_4_2_U34 ( .A1(npu_inst_int_data_x_4__2__1_), .A2(
        npu_inst_pe_1_4_2_int_q_weight_1_), .ZN(npu_inst_pe_1_4_2_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_4_2_U33 ( .A1(npu_inst_int_data_x_4__2__0_), .A2(
        npu_inst_pe_1_4_2_int_q_weight_1_), .ZN(npu_inst_pe_1_4_2_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_4_2_U32 ( .A1(npu_inst_n56), .A2(
        npu_inst_int_data_y_5__2__1_), .B1(npu_inst_pe_1_4_2_n3), .B2(
        npu_inst_int_data_x_4__3__1_), .ZN(npu_inst_pe_1_4_2_n63) );
  AOI22_X1 npu_inst_pe_1_4_2_U31 ( .A1(npu_inst_n56), .A2(
        npu_inst_int_data_y_5__2__0_), .B1(npu_inst_pe_1_4_2_n3), .B2(
        npu_inst_int_data_x_4__3__0_), .ZN(npu_inst_pe_1_4_2_n61) );
  INV_X1 npu_inst_pe_1_4_2_U30 ( .A(npu_inst_pe_1_4_2_int_data_0_), .ZN(
        npu_inst_pe_1_4_2_n13) );
  INV_X1 npu_inst_pe_1_4_2_U29 ( .A(npu_inst_n69), .ZN(npu_inst_pe_1_4_2_n5)
         );
  OR3_X1 npu_inst_pe_1_4_2_U28 ( .A1(npu_inst_pe_1_4_2_n6), .A2(
        npu_inst_pe_1_4_2_n8), .A3(npu_inst_pe_1_4_2_n5), .ZN(
        npu_inst_pe_1_4_2_n56) );
  OR3_X1 npu_inst_pe_1_4_2_U27 ( .A1(npu_inst_pe_1_4_2_n5), .A2(
        npu_inst_pe_1_4_2_n8), .A3(npu_inst_pe_1_4_2_n7), .ZN(
        npu_inst_pe_1_4_2_n48) );
  INV_X1 npu_inst_pe_1_4_2_U26 ( .A(npu_inst_pe_1_4_2_n5), .ZN(
        npu_inst_pe_1_4_2_n4) );
  OR3_X1 npu_inst_pe_1_4_2_U25 ( .A1(npu_inst_pe_1_4_2_n4), .A2(
        npu_inst_pe_1_4_2_n8), .A3(npu_inst_pe_1_4_2_n7), .ZN(
        npu_inst_pe_1_4_2_n52) );
  OR3_X1 npu_inst_pe_1_4_2_U24 ( .A1(npu_inst_pe_1_4_2_n6), .A2(
        npu_inst_pe_1_4_2_n8), .A3(npu_inst_pe_1_4_2_n4), .ZN(
        npu_inst_pe_1_4_2_n60) );
  NOR2_X1 npu_inst_pe_1_4_2_U23 ( .A1(npu_inst_pe_1_4_2_n60), .A2(
        npu_inst_pe_1_4_2_n3), .ZN(npu_inst_pe_1_4_2_n58) );
  NOR2_X1 npu_inst_pe_1_4_2_U22 ( .A1(npu_inst_pe_1_4_2_n56), .A2(
        npu_inst_pe_1_4_2_n3), .ZN(npu_inst_pe_1_4_2_n54) );
  NOR2_X1 npu_inst_pe_1_4_2_U21 ( .A1(npu_inst_pe_1_4_2_n52), .A2(
        npu_inst_pe_1_4_2_n3), .ZN(npu_inst_pe_1_4_2_n50) );
  NOR2_X1 npu_inst_pe_1_4_2_U20 ( .A1(npu_inst_pe_1_4_2_n48), .A2(
        npu_inst_pe_1_4_2_n3), .ZN(npu_inst_pe_1_4_2_n46) );
  NOR2_X1 npu_inst_pe_1_4_2_U19 ( .A1(npu_inst_pe_1_4_2_n40), .A2(
        npu_inst_pe_1_4_2_n3), .ZN(npu_inst_pe_1_4_2_n38) );
  NOR2_X1 npu_inst_pe_1_4_2_U18 ( .A1(npu_inst_pe_1_4_2_n44), .A2(
        npu_inst_pe_1_4_2_n3), .ZN(npu_inst_pe_1_4_2_n42) );
  BUF_X1 npu_inst_pe_1_4_2_U17 ( .A(npu_inst_n99), .Z(npu_inst_pe_1_4_2_n8) );
  INV_X1 npu_inst_pe_1_4_2_U16 ( .A(npu_inst_n124), .ZN(npu_inst_pe_1_4_2_n12)
         );
  INV_X1 npu_inst_pe_1_4_2_U15 ( .A(npu_inst_pe_1_4_2_n38), .ZN(
        npu_inst_pe_1_4_2_n114) );
  INV_X1 npu_inst_pe_1_4_2_U14 ( .A(npu_inst_pe_1_4_2_n58), .ZN(
        npu_inst_pe_1_4_2_n119) );
  INV_X1 npu_inst_pe_1_4_2_U13 ( .A(npu_inst_pe_1_4_2_n54), .ZN(
        npu_inst_pe_1_4_2_n118) );
  INV_X1 npu_inst_pe_1_4_2_U12 ( .A(npu_inst_pe_1_4_2_n50), .ZN(
        npu_inst_pe_1_4_2_n117) );
  INV_X1 npu_inst_pe_1_4_2_U11 ( .A(npu_inst_pe_1_4_2_n46), .ZN(
        npu_inst_pe_1_4_2_n116) );
  INV_X1 npu_inst_pe_1_4_2_U10 ( .A(npu_inst_pe_1_4_2_n42), .ZN(
        npu_inst_pe_1_4_2_n115) );
  BUF_X1 npu_inst_pe_1_4_2_U9 ( .A(npu_inst_n21), .Z(npu_inst_pe_1_4_2_n2) );
  BUF_X1 npu_inst_pe_1_4_2_U8 ( .A(npu_inst_n21), .Z(npu_inst_pe_1_4_2_n1) );
  BUF_X1 npu_inst_pe_1_4_2_U7 ( .A(npu_inst_pe_1_4_2_n12), .Z(
        npu_inst_pe_1_4_2_n11) );
  BUF_X1 npu_inst_pe_1_4_2_U6 ( .A(npu_inst_pe_1_4_2_n12), .Z(
        npu_inst_pe_1_4_2_n10) );
  BUF_X1 npu_inst_pe_1_4_2_U5 ( .A(npu_inst_pe_1_4_2_n12), .Z(
        npu_inst_pe_1_4_2_n9) );
  NOR2_X1 npu_inst_pe_1_4_2_U4 ( .A1(npu_inst_pe_1_4_2_int_q_weight_0_), .A2(
        npu_inst_pe_1_4_2_n1), .ZN(npu_inst_pe_1_4_2_n76) );
  NOR2_X1 npu_inst_pe_1_4_2_U3 ( .A1(npu_inst_pe_1_4_2_n27), .A2(
        npu_inst_pe_1_4_2_n1), .ZN(npu_inst_pe_1_4_2_n77) );
  FA_X1 npu_inst_pe_1_4_2_sub_67_U2_1 ( .A(npu_inst_pe_1_4_2_int_q_acc_1_), 
        .B(npu_inst_pe_1_4_2_n14), .CI(npu_inst_pe_1_4_2_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_4_2_sub_67_carry_2_), .S(npu_inst_pe_1_4_2_N66) );
  FA_X1 npu_inst_pe_1_4_2_add_69_U1_1 ( .A(npu_inst_pe_1_4_2_int_q_acc_1_), 
        .B(npu_inst_pe_1_4_2_int_data_1_), .CI(
        npu_inst_pe_1_4_2_add_69_carry_1_), .CO(
        npu_inst_pe_1_4_2_add_69_carry_2_), .S(npu_inst_pe_1_4_2_N74) );
  NAND3_X1 npu_inst_pe_1_4_2_U109 ( .A1(npu_inst_pe_1_4_2_n5), .A2(
        npu_inst_pe_1_4_2_n7), .A3(npu_inst_pe_1_4_2_n8), .ZN(
        npu_inst_pe_1_4_2_n44) );
  NAND3_X1 npu_inst_pe_1_4_2_U108 ( .A1(npu_inst_pe_1_4_2_n4), .A2(
        npu_inst_pe_1_4_2_n7), .A3(npu_inst_pe_1_4_2_n8), .ZN(
        npu_inst_pe_1_4_2_n40) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_4_2_n34), .CK(
        npu_inst_pe_1_4_2_net3780), .RN(npu_inst_pe_1_4_2_n9), .Q(
        npu_inst_pe_1_4_2_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_4_2_n35), .CK(
        npu_inst_pe_1_4_2_net3780), .RN(npu_inst_pe_1_4_2_n9), .Q(
        npu_inst_pe_1_4_2_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_4_2_n36), .CK(
        npu_inst_pe_1_4_2_net3780), .RN(npu_inst_pe_1_4_2_n9), .Q(
        npu_inst_pe_1_4_2_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_4_2_n98), .CK(
        npu_inst_pe_1_4_2_net3780), .RN(npu_inst_pe_1_4_2_n9), .Q(
        npu_inst_pe_1_4_2_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_4_2_n99), .CK(
        npu_inst_pe_1_4_2_net3780), .RN(npu_inst_pe_1_4_2_n9), .Q(
        npu_inst_pe_1_4_2_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_4_2_n100), 
        .CK(npu_inst_pe_1_4_2_net3780), .RN(npu_inst_pe_1_4_2_n9), .Q(
        npu_inst_pe_1_4_2_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_4_2_n33), .CK(
        npu_inst_pe_1_4_2_net3780), .RN(npu_inst_pe_1_4_2_n9), .Q(
        npu_inst_pe_1_4_2_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_4_2_n101), 
        .CK(npu_inst_pe_1_4_2_net3780), .RN(npu_inst_pe_1_4_2_n9), .Q(
        npu_inst_pe_1_4_2_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_weight_reg_0_ ( .D(npu_inst_n110), .CK(
        npu_inst_pe_1_4_2_net3786), .RN(npu_inst_pe_1_4_2_n9), .Q(
        npu_inst_pe_1_4_2_int_q_weight_0_), .QN(npu_inst_pe_1_4_2_n27) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_weight_reg_1_ ( .D(npu_inst_n116), .CK(
        npu_inst_pe_1_4_2_net3786), .RN(npu_inst_pe_1_4_2_n9), .Q(
        npu_inst_pe_1_4_2_int_q_weight_1_), .QN(npu_inst_pe_1_4_2_n26) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_4_2_n113), 
        .CK(npu_inst_pe_1_4_2_net3786), .RN(npu_inst_pe_1_4_2_n9), .Q(
        npu_inst_pe_1_4_2_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_4_2_n107), 
        .CK(npu_inst_pe_1_4_2_net3786), .RN(npu_inst_pe_1_4_2_n9), .Q(
        npu_inst_pe_1_4_2_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_4_2_n112), 
        .CK(npu_inst_pe_1_4_2_net3786), .RN(npu_inst_pe_1_4_2_n10), .Q(
        npu_inst_pe_1_4_2_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_4_2_n106), 
        .CK(npu_inst_pe_1_4_2_net3786), .RN(npu_inst_pe_1_4_2_n10), .Q(
        npu_inst_pe_1_4_2_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_4_2_n111), 
        .CK(npu_inst_pe_1_4_2_net3786), .RN(npu_inst_pe_1_4_2_n10), .Q(
        npu_inst_pe_1_4_2_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_4_2_n105), 
        .CK(npu_inst_pe_1_4_2_net3786), .RN(npu_inst_pe_1_4_2_n10), .Q(
        npu_inst_pe_1_4_2_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_4_2_n110), 
        .CK(npu_inst_pe_1_4_2_net3786), .RN(npu_inst_pe_1_4_2_n10), .Q(
        npu_inst_pe_1_4_2_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_4_2_n104), 
        .CK(npu_inst_pe_1_4_2_net3786), .RN(npu_inst_pe_1_4_2_n10), .Q(
        npu_inst_pe_1_4_2_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_4_2_n109), 
        .CK(npu_inst_pe_1_4_2_net3786), .RN(npu_inst_pe_1_4_2_n10), .Q(
        npu_inst_pe_1_4_2_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_4_2_n103), 
        .CK(npu_inst_pe_1_4_2_net3786), .RN(npu_inst_pe_1_4_2_n10), .Q(
        npu_inst_pe_1_4_2_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_4_2_n108), 
        .CK(npu_inst_pe_1_4_2_net3786), .RN(npu_inst_pe_1_4_2_n10), .Q(
        npu_inst_pe_1_4_2_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_4_2_n102), 
        .CK(npu_inst_pe_1_4_2_net3786), .RN(npu_inst_pe_1_4_2_n10), .Q(
        npu_inst_pe_1_4_2_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_4_2_n86), 
        .CK(npu_inst_pe_1_4_2_net3786), .RN(npu_inst_pe_1_4_2_n10), .Q(
        npu_inst_pe_1_4_2_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_4_2_n87), 
        .CK(npu_inst_pe_1_4_2_net3786), .RN(npu_inst_pe_1_4_2_n10), .Q(
        npu_inst_pe_1_4_2_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_4_2_n88), 
        .CK(npu_inst_pe_1_4_2_net3786), .RN(npu_inst_pe_1_4_2_n11), .Q(
        npu_inst_pe_1_4_2_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_4_2_n89), 
        .CK(npu_inst_pe_1_4_2_net3786), .RN(npu_inst_pe_1_4_2_n11), .Q(
        npu_inst_pe_1_4_2_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_4_2_n90), 
        .CK(npu_inst_pe_1_4_2_net3786), .RN(npu_inst_pe_1_4_2_n11), .Q(
        npu_inst_pe_1_4_2_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_4_2_n91), 
        .CK(npu_inst_pe_1_4_2_net3786), .RN(npu_inst_pe_1_4_2_n11), .Q(
        npu_inst_pe_1_4_2_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_4_2_n92), 
        .CK(npu_inst_pe_1_4_2_net3786), .RN(npu_inst_pe_1_4_2_n11), .Q(
        npu_inst_pe_1_4_2_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_4_2_n93), 
        .CK(npu_inst_pe_1_4_2_net3786), .RN(npu_inst_pe_1_4_2_n11), .Q(
        npu_inst_pe_1_4_2_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_4_2_n94), 
        .CK(npu_inst_pe_1_4_2_net3786), .RN(npu_inst_pe_1_4_2_n11), .Q(
        npu_inst_pe_1_4_2_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_4_2_n95), 
        .CK(npu_inst_pe_1_4_2_net3786), .RN(npu_inst_pe_1_4_2_n11), .Q(
        npu_inst_pe_1_4_2_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_4_2_n96), 
        .CK(npu_inst_pe_1_4_2_net3786), .RN(npu_inst_pe_1_4_2_n11), .Q(
        npu_inst_pe_1_4_2_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_4_2_n97), 
        .CK(npu_inst_pe_1_4_2_net3786), .RN(npu_inst_pe_1_4_2_n11), .Q(
        npu_inst_pe_1_4_2_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_4_2_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_4_2_N84), .SE(1'b0), .GCK(npu_inst_pe_1_4_2_net3780) );
  CLKGATETST_X1 npu_inst_pe_1_4_2_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n63), .SE(1'b0), .GCK(npu_inst_pe_1_4_2_net3786) );
  MUX2_X1 npu_inst_pe_1_4_3_U162 ( .A(npu_inst_pe_1_4_3_n32), .B(
        npu_inst_pe_1_4_3_n29), .S(npu_inst_pe_1_4_3_n8), .Z(
        npu_inst_pe_1_4_3_N93) );
  MUX2_X1 npu_inst_pe_1_4_3_U161 ( .A(npu_inst_pe_1_4_3_n31), .B(
        npu_inst_pe_1_4_3_n30), .S(npu_inst_pe_1_4_3_n6), .Z(
        npu_inst_pe_1_4_3_n32) );
  MUX2_X1 npu_inst_pe_1_4_3_U160 ( .A(npu_inst_pe_1_4_3_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_4_3_int_q_reg_v_1__0_), .S(npu_inst_pe_1_4_3_n4), .Z(
        npu_inst_pe_1_4_3_n31) );
  MUX2_X1 npu_inst_pe_1_4_3_U159 ( .A(npu_inst_pe_1_4_3_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_4_3_int_q_reg_v_3__0_), .S(npu_inst_pe_1_4_3_n4), .Z(
        npu_inst_pe_1_4_3_n30) );
  MUX2_X1 npu_inst_pe_1_4_3_U158 ( .A(npu_inst_pe_1_4_3_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_4_3_int_q_reg_v_5__0_), .S(npu_inst_pe_1_4_3_n4), .Z(
        npu_inst_pe_1_4_3_n29) );
  MUX2_X1 npu_inst_pe_1_4_3_U157 ( .A(npu_inst_pe_1_4_3_n28), .B(
        npu_inst_pe_1_4_3_n23), .S(npu_inst_pe_1_4_3_n8), .Z(
        npu_inst_pe_1_4_3_N94) );
  MUX2_X1 npu_inst_pe_1_4_3_U156 ( .A(npu_inst_pe_1_4_3_n25), .B(
        npu_inst_pe_1_4_3_n24), .S(npu_inst_pe_1_4_3_n6), .Z(
        npu_inst_pe_1_4_3_n28) );
  MUX2_X1 npu_inst_pe_1_4_3_U155 ( .A(npu_inst_pe_1_4_3_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_4_3_int_q_reg_v_1__1_), .S(npu_inst_pe_1_4_3_n4), .Z(
        npu_inst_pe_1_4_3_n25) );
  MUX2_X1 npu_inst_pe_1_4_3_U154 ( .A(npu_inst_pe_1_4_3_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_4_3_int_q_reg_v_3__1_), .S(npu_inst_pe_1_4_3_n4), .Z(
        npu_inst_pe_1_4_3_n24) );
  MUX2_X1 npu_inst_pe_1_4_3_U153 ( .A(npu_inst_pe_1_4_3_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_4_3_int_q_reg_v_5__1_), .S(npu_inst_pe_1_4_3_n4), .Z(
        npu_inst_pe_1_4_3_n23) );
  MUX2_X1 npu_inst_pe_1_4_3_U152 ( .A(npu_inst_pe_1_4_3_n22), .B(
        npu_inst_pe_1_4_3_n19), .S(npu_inst_pe_1_4_3_n8), .Z(
        npu_inst_int_data_x_4__3__1_) );
  MUX2_X1 npu_inst_pe_1_4_3_U151 ( .A(npu_inst_pe_1_4_3_n21), .B(
        npu_inst_pe_1_4_3_n20), .S(npu_inst_pe_1_4_3_n6), .Z(
        npu_inst_pe_1_4_3_n22) );
  MUX2_X1 npu_inst_pe_1_4_3_U150 ( .A(npu_inst_pe_1_4_3_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_4_3_int_q_reg_h_1__1_), .S(npu_inst_pe_1_4_3_n4), .Z(
        npu_inst_pe_1_4_3_n21) );
  MUX2_X1 npu_inst_pe_1_4_3_U149 ( .A(npu_inst_pe_1_4_3_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_4_3_int_q_reg_h_3__1_), .S(npu_inst_pe_1_4_3_n4), .Z(
        npu_inst_pe_1_4_3_n20) );
  MUX2_X1 npu_inst_pe_1_4_3_U148 ( .A(npu_inst_pe_1_4_3_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_4_3_int_q_reg_h_5__1_), .S(npu_inst_pe_1_4_3_n4), .Z(
        npu_inst_pe_1_4_3_n19) );
  MUX2_X1 npu_inst_pe_1_4_3_U147 ( .A(npu_inst_pe_1_4_3_n18), .B(
        npu_inst_pe_1_4_3_n15), .S(npu_inst_pe_1_4_3_n8), .Z(
        npu_inst_int_data_x_4__3__0_) );
  MUX2_X1 npu_inst_pe_1_4_3_U146 ( .A(npu_inst_pe_1_4_3_n17), .B(
        npu_inst_pe_1_4_3_n16), .S(npu_inst_pe_1_4_3_n6), .Z(
        npu_inst_pe_1_4_3_n18) );
  MUX2_X1 npu_inst_pe_1_4_3_U145 ( .A(npu_inst_pe_1_4_3_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_4_3_int_q_reg_h_1__0_), .S(npu_inst_pe_1_4_3_n4), .Z(
        npu_inst_pe_1_4_3_n17) );
  MUX2_X1 npu_inst_pe_1_4_3_U144 ( .A(npu_inst_pe_1_4_3_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_4_3_int_q_reg_h_3__0_), .S(npu_inst_pe_1_4_3_n4), .Z(
        npu_inst_pe_1_4_3_n16) );
  MUX2_X1 npu_inst_pe_1_4_3_U143 ( .A(npu_inst_pe_1_4_3_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_4_3_int_q_reg_h_5__0_), .S(npu_inst_pe_1_4_3_n4), .Z(
        npu_inst_pe_1_4_3_n15) );
  XOR2_X1 npu_inst_pe_1_4_3_U142 ( .A(npu_inst_pe_1_4_3_int_data_0_), .B(
        npu_inst_pe_1_4_3_int_q_acc_0_), .Z(npu_inst_pe_1_4_3_N73) );
  AND2_X1 npu_inst_pe_1_4_3_U141 ( .A1(npu_inst_pe_1_4_3_int_q_acc_0_), .A2(
        npu_inst_pe_1_4_3_int_data_0_), .ZN(npu_inst_pe_1_4_3_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_4_3_U140 ( .A(npu_inst_pe_1_4_3_int_q_acc_0_), .B(
        npu_inst_pe_1_4_3_n13), .ZN(npu_inst_pe_1_4_3_N65) );
  OR2_X1 npu_inst_pe_1_4_3_U139 ( .A1(npu_inst_pe_1_4_3_n13), .A2(
        npu_inst_pe_1_4_3_int_q_acc_0_), .ZN(npu_inst_pe_1_4_3_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_4_3_U138 ( .A(npu_inst_pe_1_4_3_int_q_acc_2_), .B(
        npu_inst_pe_1_4_3_add_69_carry_2_), .Z(npu_inst_pe_1_4_3_N75) );
  AND2_X1 npu_inst_pe_1_4_3_U137 ( .A1(npu_inst_pe_1_4_3_add_69_carry_2_), 
        .A2(npu_inst_pe_1_4_3_int_q_acc_2_), .ZN(
        npu_inst_pe_1_4_3_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_4_3_U136 ( .A(npu_inst_pe_1_4_3_int_q_acc_3_), .B(
        npu_inst_pe_1_4_3_add_69_carry_3_), .Z(npu_inst_pe_1_4_3_N76) );
  AND2_X1 npu_inst_pe_1_4_3_U135 ( .A1(npu_inst_pe_1_4_3_add_69_carry_3_), 
        .A2(npu_inst_pe_1_4_3_int_q_acc_3_), .ZN(
        npu_inst_pe_1_4_3_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_4_3_U134 ( .A(npu_inst_pe_1_4_3_int_q_acc_4_), .B(
        npu_inst_pe_1_4_3_add_69_carry_4_), .Z(npu_inst_pe_1_4_3_N77) );
  AND2_X1 npu_inst_pe_1_4_3_U133 ( .A1(npu_inst_pe_1_4_3_add_69_carry_4_), 
        .A2(npu_inst_pe_1_4_3_int_q_acc_4_), .ZN(
        npu_inst_pe_1_4_3_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_4_3_U132 ( .A(npu_inst_pe_1_4_3_int_q_acc_5_), .B(
        npu_inst_pe_1_4_3_add_69_carry_5_), .Z(npu_inst_pe_1_4_3_N78) );
  AND2_X1 npu_inst_pe_1_4_3_U131 ( .A1(npu_inst_pe_1_4_3_add_69_carry_5_), 
        .A2(npu_inst_pe_1_4_3_int_q_acc_5_), .ZN(
        npu_inst_pe_1_4_3_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_4_3_U130 ( .A(npu_inst_pe_1_4_3_int_q_acc_6_), .B(
        npu_inst_pe_1_4_3_add_69_carry_6_), .Z(npu_inst_pe_1_4_3_N79) );
  AND2_X1 npu_inst_pe_1_4_3_U129 ( .A1(npu_inst_pe_1_4_3_add_69_carry_6_), 
        .A2(npu_inst_pe_1_4_3_int_q_acc_6_), .ZN(
        npu_inst_pe_1_4_3_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_4_3_U128 ( .A(npu_inst_pe_1_4_3_int_q_acc_7_), .B(
        npu_inst_pe_1_4_3_add_69_carry_7_), .Z(npu_inst_pe_1_4_3_N80) );
  XNOR2_X1 npu_inst_pe_1_4_3_U127 ( .A(npu_inst_pe_1_4_3_sub_67_carry_2_), .B(
        npu_inst_pe_1_4_3_int_q_acc_2_), .ZN(npu_inst_pe_1_4_3_N67) );
  OR2_X1 npu_inst_pe_1_4_3_U126 ( .A1(npu_inst_pe_1_4_3_int_q_acc_2_), .A2(
        npu_inst_pe_1_4_3_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_4_3_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_4_3_U125 ( .A(npu_inst_pe_1_4_3_sub_67_carry_3_), .B(
        npu_inst_pe_1_4_3_int_q_acc_3_), .ZN(npu_inst_pe_1_4_3_N68) );
  OR2_X1 npu_inst_pe_1_4_3_U124 ( .A1(npu_inst_pe_1_4_3_int_q_acc_3_), .A2(
        npu_inst_pe_1_4_3_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_4_3_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_4_3_U123 ( .A(npu_inst_pe_1_4_3_sub_67_carry_4_), .B(
        npu_inst_pe_1_4_3_int_q_acc_4_), .ZN(npu_inst_pe_1_4_3_N69) );
  OR2_X1 npu_inst_pe_1_4_3_U122 ( .A1(npu_inst_pe_1_4_3_int_q_acc_4_), .A2(
        npu_inst_pe_1_4_3_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_4_3_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_4_3_U121 ( .A(npu_inst_pe_1_4_3_sub_67_carry_5_), .B(
        npu_inst_pe_1_4_3_int_q_acc_5_), .ZN(npu_inst_pe_1_4_3_N70) );
  OR2_X1 npu_inst_pe_1_4_3_U120 ( .A1(npu_inst_pe_1_4_3_int_q_acc_5_), .A2(
        npu_inst_pe_1_4_3_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_4_3_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_4_3_U119 ( .A(npu_inst_pe_1_4_3_sub_67_carry_6_), .B(
        npu_inst_pe_1_4_3_int_q_acc_6_), .ZN(npu_inst_pe_1_4_3_N71) );
  OR2_X1 npu_inst_pe_1_4_3_U118 ( .A1(npu_inst_pe_1_4_3_int_q_acc_6_), .A2(
        npu_inst_pe_1_4_3_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_4_3_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_4_3_U117 ( .A(npu_inst_pe_1_4_3_int_q_acc_7_), .B(
        npu_inst_pe_1_4_3_sub_67_carry_7_), .ZN(npu_inst_pe_1_4_3_N72) );
  INV_X1 npu_inst_pe_1_4_3_U116 ( .A(npu_inst_n77), .ZN(npu_inst_pe_1_4_3_n7)
         );
  INV_X1 npu_inst_pe_1_4_3_U115 ( .A(npu_inst_pe_1_4_3_n7), .ZN(
        npu_inst_pe_1_4_3_n6) );
  INV_X1 npu_inst_pe_1_4_3_U114 ( .A(npu_inst_n56), .ZN(npu_inst_pe_1_4_3_n3)
         );
  AOI22_X1 npu_inst_pe_1_4_3_U113 ( .A1(npu_inst_int_data_y_5__3__0_), .A2(
        npu_inst_pe_1_4_3_n58), .B1(npu_inst_pe_1_4_3_n119), .B2(
        npu_inst_pe_1_4_3_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_4_3_n57) );
  INV_X1 npu_inst_pe_1_4_3_U112 ( .A(npu_inst_pe_1_4_3_n57), .ZN(
        npu_inst_pe_1_4_3_n108) );
  AOI22_X1 npu_inst_pe_1_4_3_U111 ( .A1(npu_inst_int_data_y_5__3__0_), .A2(
        npu_inst_pe_1_4_3_n54), .B1(npu_inst_pe_1_4_3_n118), .B2(
        npu_inst_pe_1_4_3_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_4_3_n53) );
  INV_X1 npu_inst_pe_1_4_3_U110 ( .A(npu_inst_pe_1_4_3_n53), .ZN(
        npu_inst_pe_1_4_3_n109) );
  AOI22_X1 npu_inst_pe_1_4_3_U107 ( .A1(npu_inst_int_data_y_5__3__0_), .A2(
        npu_inst_pe_1_4_3_n50), .B1(npu_inst_pe_1_4_3_n117), .B2(
        npu_inst_pe_1_4_3_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_4_3_n49) );
  INV_X1 npu_inst_pe_1_4_3_U106 ( .A(npu_inst_pe_1_4_3_n49), .ZN(
        npu_inst_pe_1_4_3_n110) );
  AOI22_X1 npu_inst_pe_1_4_3_U105 ( .A1(npu_inst_int_data_y_5__3__0_), .A2(
        npu_inst_pe_1_4_3_n46), .B1(npu_inst_pe_1_4_3_n116), .B2(
        npu_inst_pe_1_4_3_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_4_3_n45) );
  INV_X1 npu_inst_pe_1_4_3_U104 ( .A(npu_inst_pe_1_4_3_n45), .ZN(
        npu_inst_pe_1_4_3_n111) );
  AOI22_X1 npu_inst_pe_1_4_3_U103 ( .A1(npu_inst_int_data_y_5__3__0_), .A2(
        npu_inst_pe_1_4_3_n42), .B1(npu_inst_pe_1_4_3_n115), .B2(
        npu_inst_pe_1_4_3_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_4_3_n41) );
  INV_X1 npu_inst_pe_1_4_3_U102 ( .A(npu_inst_pe_1_4_3_n41), .ZN(
        npu_inst_pe_1_4_3_n112) );
  AOI22_X1 npu_inst_pe_1_4_3_U101 ( .A1(npu_inst_int_data_y_5__3__1_), .A2(
        npu_inst_pe_1_4_3_n58), .B1(npu_inst_pe_1_4_3_n119), .B2(
        npu_inst_pe_1_4_3_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_4_3_n59) );
  INV_X1 npu_inst_pe_1_4_3_U100 ( .A(npu_inst_pe_1_4_3_n59), .ZN(
        npu_inst_pe_1_4_3_n102) );
  AOI22_X1 npu_inst_pe_1_4_3_U99 ( .A1(npu_inst_int_data_y_5__3__1_), .A2(
        npu_inst_pe_1_4_3_n54), .B1(npu_inst_pe_1_4_3_n118), .B2(
        npu_inst_pe_1_4_3_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_4_3_n55) );
  INV_X1 npu_inst_pe_1_4_3_U98 ( .A(npu_inst_pe_1_4_3_n55), .ZN(
        npu_inst_pe_1_4_3_n103) );
  AOI22_X1 npu_inst_pe_1_4_3_U97 ( .A1(npu_inst_int_data_y_5__3__1_), .A2(
        npu_inst_pe_1_4_3_n50), .B1(npu_inst_pe_1_4_3_n117), .B2(
        npu_inst_pe_1_4_3_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_4_3_n51) );
  INV_X1 npu_inst_pe_1_4_3_U96 ( .A(npu_inst_pe_1_4_3_n51), .ZN(
        npu_inst_pe_1_4_3_n104) );
  AOI22_X1 npu_inst_pe_1_4_3_U95 ( .A1(npu_inst_int_data_y_5__3__1_), .A2(
        npu_inst_pe_1_4_3_n46), .B1(npu_inst_pe_1_4_3_n116), .B2(
        npu_inst_pe_1_4_3_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_4_3_n47) );
  INV_X1 npu_inst_pe_1_4_3_U94 ( .A(npu_inst_pe_1_4_3_n47), .ZN(
        npu_inst_pe_1_4_3_n105) );
  AOI22_X1 npu_inst_pe_1_4_3_U93 ( .A1(npu_inst_int_data_y_5__3__1_), .A2(
        npu_inst_pe_1_4_3_n42), .B1(npu_inst_pe_1_4_3_n115), .B2(
        npu_inst_pe_1_4_3_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_4_3_n43) );
  INV_X1 npu_inst_pe_1_4_3_U92 ( .A(npu_inst_pe_1_4_3_n43), .ZN(
        npu_inst_pe_1_4_3_n106) );
  AOI22_X1 npu_inst_pe_1_4_3_U91 ( .A1(npu_inst_pe_1_4_3_n38), .A2(
        npu_inst_int_data_y_5__3__1_), .B1(npu_inst_pe_1_4_3_n114), .B2(
        npu_inst_pe_1_4_3_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_4_3_n39) );
  INV_X1 npu_inst_pe_1_4_3_U90 ( .A(npu_inst_pe_1_4_3_n39), .ZN(
        npu_inst_pe_1_4_3_n107) );
  AOI22_X1 npu_inst_pe_1_4_3_U89 ( .A1(npu_inst_pe_1_4_3_n38), .A2(
        npu_inst_int_data_y_5__3__0_), .B1(npu_inst_pe_1_4_3_n114), .B2(
        npu_inst_pe_1_4_3_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_4_3_n37) );
  INV_X1 npu_inst_pe_1_4_3_U88 ( .A(npu_inst_pe_1_4_3_n37), .ZN(
        npu_inst_pe_1_4_3_n113) );
  NAND2_X1 npu_inst_pe_1_4_3_U87 ( .A1(npu_inst_pe_1_4_3_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_4_3_n60), .ZN(npu_inst_pe_1_4_3_n74) );
  OAI21_X1 npu_inst_pe_1_4_3_U86 ( .B1(npu_inst_pe_1_4_3_n63), .B2(
        npu_inst_pe_1_4_3_n60), .A(npu_inst_pe_1_4_3_n74), .ZN(
        npu_inst_pe_1_4_3_n97) );
  NAND2_X1 npu_inst_pe_1_4_3_U85 ( .A1(npu_inst_pe_1_4_3_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_4_3_n60), .ZN(npu_inst_pe_1_4_3_n73) );
  OAI21_X1 npu_inst_pe_1_4_3_U84 ( .B1(npu_inst_pe_1_4_3_n61), .B2(
        npu_inst_pe_1_4_3_n60), .A(npu_inst_pe_1_4_3_n73), .ZN(
        npu_inst_pe_1_4_3_n96) );
  NAND2_X1 npu_inst_pe_1_4_3_U83 ( .A1(npu_inst_pe_1_4_3_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_4_3_n56), .ZN(npu_inst_pe_1_4_3_n72) );
  OAI21_X1 npu_inst_pe_1_4_3_U82 ( .B1(npu_inst_pe_1_4_3_n63), .B2(
        npu_inst_pe_1_4_3_n56), .A(npu_inst_pe_1_4_3_n72), .ZN(
        npu_inst_pe_1_4_3_n95) );
  NAND2_X1 npu_inst_pe_1_4_3_U81 ( .A1(npu_inst_pe_1_4_3_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_4_3_n56), .ZN(npu_inst_pe_1_4_3_n71) );
  OAI21_X1 npu_inst_pe_1_4_3_U80 ( .B1(npu_inst_pe_1_4_3_n61), .B2(
        npu_inst_pe_1_4_3_n56), .A(npu_inst_pe_1_4_3_n71), .ZN(
        npu_inst_pe_1_4_3_n94) );
  NAND2_X1 npu_inst_pe_1_4_3_U79 ( .A1(npu_inst_pe_1_4_3_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_4_3_n52), .ZN(npu_inst_pe_1_4_3_n70) );
  OAI21_X1 npu_inst_pe_1_4_3_U78 ( .B1(npu_inst_pe_1_4_3_n63), .B2(
        npu_inst_pe_1_4_3_n52), .A(npu_inst_pe_1_4_3_n70), .ZN(
        npu_inst_pe_1_4_3_n93) );
  NAND2_X1 npu_inst_pe_1_4_3_U77 ( .A1(npu_inst_pe_1_4_3_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_4_3_n52), .ZN(npu_inst_pe_1_4_3_n69) );
  OAI21_X1 npu_inst_pe_1_4_3_U76 ( .B1(npu_inst_pe_1_4_3_n61), .B2(
        npu_inst_pe_1_4_3_n52), .A(npu_inst_pe_1_4_3_n69), .ZN(
        npu_inst_pe_1_4_3_n92) );
  NAND2_X1 npu_inst_pe_1_4_3_U75 ( .A1(npu_inst_pe_1_4_3_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_4_3_n48), .ZN(npu_inst_pe_1_4_3_n68) );
  OAI21_X1 npu_inst_pe_1_4_3_U74 ( .B1(npu_inst_pe_1_4_3_n63), .B2(
        npu_inst_pe_1_4_3_n48), .A(npu_inst_pe_1_4_3_n68), .ZN(
        npu_inst_pe_1_4_3_n91) );
  NAND2_X1 npu_inst_pe_1_4_3_U73 ( .A1(npu_inst_pe_1_4_3_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_4_3_n48), .ZN(npu_inst_pe_1_4_3_n67) );
  OAI21_X1 npu_inst_pe_1_4_3_U72 ( .B1(npu_inst_pe_1_4_3_n61), .B2(
        npu_inst_pe_1_4_3_n48), .A(npu_inst_pe_1_4_3_n67), .ZN(
        npu_inst_pe_1_4_3_n90) );
  NAND2_X1 npu_inst_pe_1_4_3_U71 ( .A1(npu_inst_pe_1_4_3_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_4_3_n44), .ZN(npu_inst_pe_1_4_3_n66) );
  OAI21_X1 npu_inst_pe_1_4_3_U70 ( .B1(npu_inst_pe_1_4_3_n63), .B2(
        npu_inst_pe_1_4_3_n44), .A(npu_inst_pe_1_4_3_n66), .ZN(
        npu_inst_pe_1_4_3_n89) );
  NAND2_X1 npu_inst_pe_1_4_3_U69 ( .A1(npu_inst_pe_1_4_3_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_4_3_n44), .ZN(npu_inst_pe_1_4_3_n65) );
  OAI21_X1 npu_inst_pe_1_4_3_U68 ( .B1(npu_inst_pe_1_4_3_n61), .B2(
        npu_inst_pe_1_4_3_n44), .A(npu_inst_pe_1_4_3_n65), .ZN(
        npu_inst_pe_1_4_3_n88) );
  NAND2_X1 npu_inst_pe_1_4_3_U67 ( .A1(npu_inst_pe_1_4_3_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_4_3_n40), .ZN(npu_inst_pe_1_4_3_n64) );
  OAI21_X1 npu_inst_pe_1_4_3_U66 ( .B1(npu_inst_pe_1_4_3_n63), .B2(
        npu_inst_pe_1_4_3_n40), .A(npu_inst_pe_1_4_3_n64), .ZN(
        npu_inst_pe_1_4_3_n87) );
  NAND2_X1 npu_inst_pe_1_4_3_U65 ( .A1(npu_inst_pe_1_4_3_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_4_3_n40), .ZN(npu_inst_pe_1_4_3_n62) );
  OAI21_X1 npu_inst_pe_1_4_3_U64 ( .B1(npu_inst_pe_1_4_3_n61), .B2(
        npu_inst_pe_1_4_3_n40), .A(npu_inst_pe_1_4_3_n62), .ZN(
        npu_inst_pe_1_4_3_n86) );
  AND2_X1 npu_inst_pe_1_4_3_U63 ( .A1(npu_inst_pe_1_4_3_N93), .A2(npu_inst_n56), .ZN(npu_inst_int_data_y_4__3__0_) );
  AND2_X1 npu_inst_pe_1_4_3_U62 ( .A1(npu_inst_n56), .A2(npu_inst_pe_1_4_3_N94), .ZN(npu_inst_int_data_y_4__3__1_) );
  NOR3_X1 npu_inst_pe_1_4_3_U61 ( .A1(npu_inst_pe_1_4_3_n26), .A2(npu_inst_n56), .A3(npu_inst_int_ckg[28]), .ZN(npu_inst_pe_1_4_3_n85) );
  OR2_X1 npu_inst_pe_1_4_3_U60 ( .A1(npu_inst_pe_1_4_3_n85), .A2(
        npu_inst_pe_1_4_3_n2), .ZN(npu_inst_pe_1_4_3_N84) );
  AND2_X1 npu_inst_pe_1_4_3_U59 ( .A1(npu_inst_pe_1_4_3_int_q_acc_0_), .A2(
        npu_inst_pe_1_4_3_n1), .ZN(npu_inst_int_data_res_4__3__0_) );
  AND2_X1 npu_inst_pe_1_4_3_U58 ( .A1(npu_inst_pe_1_4_3_n2), .A2(
        npu_inst_pe_1_4_3_int_q_acc_7_), .ZN(npu_inst_int_data_res_4__3__7_)
         );
  AND2_X1 npu_inst_pe_1_4_3_U57 ( .A1(npu_inst_pe_1_4_3_int_q_acc_1_), .A2(
        npu_inst_pe_1_4_3_n1), .ZN(npu_inst_int_data_res_4__3__1_) );
  AND2_X1 npu_inst_pe_1_4_3_U56 ( .A1(npu_inst_pe_1_4_3_int_q_acc_2_), .A2(
        npu_inst_pe_1_4_3_n1), .ZN(npu_inst_int_data_res_4__3__2_) );
  AND2_X1 npu_inst_pe_1_4_3_U55 ( .A1(npu_inst_pe_1_4_3_int_q_acc_3_), .A2(
        npu_inst_pe_1_4_3_n2), .ZN(npu_inst_int_data_res_4__3__3_) );
  AND2_X1 npu_inst_pe_1_4_3_U54 ( .A1(npu_inst_pe_1_4_3_int_q_acc_4_), .A2(
        npu_inst_pe_1_4_3_n2), .ZN(npu_inst_int_data_res_4__3__4_) );
  AND2_X1 npu_inst_pe_1_4_3_U53 ( .A1(npu_inst_pe_1_4_3_int_q_acc_5_), .A2(
        npu_inst_pe_1_4_3_n2), .ZN(npu_inst_int_data_res_4__3__5_) );
  AND2_X1 npu_inst_pe_1_4_3_U52 ( .A1(npu_inst_pe_1_4_3_int_q_acc_6_), .A2(
        npu_inst_pe_1_4_3_n2), .ZN(npu_inst_int_data_res_4__3__6_) );
  AOI222_X1 npu_inst_pe_1_4_3_U51 ( .A1(npu_inst_int_data_res_5__3__0_), .A2(
        npu_inst_pe_1_4_3_n1), .B1(npu_inst_pe_1_4_3_N73), .B2(
        npu_inst_pe_1_4_3_n76), .C1(npu_inst_pe_1_4_3_N65), .C2(
        npu_inst_pe_1_4_3_n77), .ZN(npu_inst_pe_1_4_3_n84) );
  INV_X1 npu_inst_pe_1_4_3_U50 ( .A(npu_inst_pe_1_4_3_n84), .ZN(
        npu_inst_pe_1_4_3_n101) );
  AOI222_X1 npu_inst_pe_1_4_3_U49 ( .A1(npu_inst_int_data_res_5__3__7_), .A2(
        npu_inst_pe_1_4_3_n1), .B1(npu_inst_pe_1_4_3_N80), .B2(
        npu_inst_pe_1_4_3_n76), .C1(npu_inst_pe_1_4_3_N72), .C2(
        npu_inst_pe_1_4_3_n77), .ZN(npu_inst_pe_1_4_3_n75) );
  INV_X1 npu_inst_pe_1_4_3_U48 ( .A(npu_inst_pe_1_4_3_n75), .ZN(
        npu_inst_pe_1_4_3_n33) );
  AOI222_X1 npu_inst_pe_1_4_3_U47 ( .A1(npu_inst_int_data_res_5__3__1_), .A2(
        npu_inst_pe_1_4_3_n1), .B1(npu_inst_pe_1_4_3_N74), .B2(
        npu_inst_pe_1_4_3_n76), .C1(npu_inst_pe_1_4_3_N66), .C2(
        npu_inst_pe_1_4_3_n77), .ZN(npu_inst_pe_1_4_3_n83) );
  INV_X1 npu_inst_pe_1_4_3_U46 ( .A(npu_inst_pe_1_4_3_n83), .ZN(
        npu_inst_pe_1_4_3_n100) );
  AOI222_X1 npu_inst_pe_1_4_3_U45 ( .A1(npu_inst_int_data_res_5__3__2_), .A2(
        npu_inst_pe_1_4_3_n1), .B1(npu_inst_pe_1_4_3_N75), .B2(
        npu_inst_pe_1_4_3_n76), .C1(npu_inst_pe_1_4_3_N67), .C2(
        npu_inst_pe_1_4_3_n77), .ZN(npu_inst_pe_1_4_3_n82) );
  INV_X1 npu_inst_pe_1_4_3_U44 ( .A(npu_inst_pe_1_4_3_n82), .ZN(
        npu_inst_pe_1_4_3_n99) );
  AOI222_X1 npu_inst_pe_1_4_3_U43 ( .A1(npu_inst_int_data_res_5__3__3_), .A2(
        npu_inst_pe_1_4_3_n1), .B1(npu_inst_pe_1_4_3_N76), .B2(
        npu_inst_pe_1_4_3_n76), .C1(npu_inst_pe_1_4_3_N68), .C2(
        npu_inst_pe_1_4_3_n77), .ZN(npu_inst_pe_1_4_3_n81) );
  INV_X1 npu_inst_pe_1_4_3_U42 ( .A(npu_inst_pe_1_4_3_n81), .ZN(
        npu_inst_pe_1_4_3_n98) );
  AOI222_X1 npu_inst_pe_1_4_3_U41 ( .A1(npu_inst_int_data_res_5__3__4_), .A2(
        npu_inst_pe_1_4_3_n1), .B1(npu_inst_pe_1_4_3_N77), .B2(
        npu_inst_pe_1_4_3_n76), .C1(npu_inst_pe_1_4_3_N69), .C2(
        npu_inst_pe_1_4_3_n77), .ZN(npu_inst_pe_1_4_3_n80) );
  INV_X1 npu_inst_pe_1_4_3_U40 ( .A(npu_inst_pe_1_4_3_n80), .ZN(
        npu_inst_pe_1_4_3_n36) );
  AOI222_X1 npu_inst_pe_1_4_3_U39 ( .A1(npu_inst_int_data_res_5__3__5_), .A2(
        npu_inst_pe_1_4_3_n1), .B1(npu_inst_pe_1_4_3_N78), .B2(
        npu_inst_pe_1_4_3_n76), .C1(npu_inst_pe_1_4_3_N70), .C2(
        npu_inst_pe_1_4_3_n77), .ZN(npu_inst_pe_1_4_3_n79) );
  INV_X1 npu_inst_pe_1_4_3_U38 ( .A(npu_inst_pe_1_4_3_n79), .ZN(
        npu_inst_pe_1_4_3_n35) );
  AOI222_X1 npu_inst_pe_1_4_3_U37 ( .A1(npu_inst_int_data_res_5__3__6_), .A2(
        npu_inst_pe_1_4_3_n1), .B1(npu_inst_pe_1_4_3_N79), .B2(
        npu_inst_pe_1_4_3_n76), .C1(npu_inst_pe_1_4_3_N71), .C2(
        npu_inst_pe_1_4_3_n77), .ZN(npu_inst_pe_1_4_3_n78) );
  INV_X1 npu_inst_pe_1_4_3_U36 ( .A(npu_inst_pe_1_4_3_n78), .ZN(
        npu_inst_pe_1_4_3_n34) );
  INV_X1 npu_inst_pe_1_4_3_U35 ( .A(npu_inst_pe_1_4_3_int_data_1_), .ZN(
        npu_inst_pe_1_4_3_n14) );
  AND2_X1 npu_inst_pe_1_4_3_U34 ( .A1(npu_inst_int_data_x_4__3__1_), .A2(
        npu_inst_pe_1_4_3_int_q_weight_1_), .ZN(npu_inst_pe_1_4_3_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_4_3_U33 ( .A1(npu_inst_int_data_x_4__3__0_), .A2(
        npu_inst_pe_1_4_3_int_q_weight_1_), .ZN(npu_inst_pe_1_4_3_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_4_3_U32 ( .A1(npu_inst_n56), .A2(
        npu_inst_int_data_y_5__3__1_), .B1(npu_inst_pe_1_4_3_n3), .B2(
        npu_inst_int_data_x_4__4__1_), .ZN(npu_inst_pe_1_4_3_n63) );
  AOI22_X1 npu_inst_pe_1_4_3_U31 ( .A1(npu_inst_n56), .A2(
        npu_inst_int_data_y_5__3__0_), .B1(npu_inst_pe_1_4_3_n3), .B2(
        npu_inst_int_data_x_4__4__0_), .ZN(npu_inst_pe_1_4_3_n61) );
  INV_X1 npu_inst_pe_1_4_3_U30 ( .A(npu_inst_pe_1_4_3_int_data_0_), .ZN(
        npu_inst_pe_1_4_3_n13) );
  INV_X1 npu_inst_pe_1_4_3_U29 ( .A(npu_inst_n69), .ZN(npu_inst_pe_1_4_3_n5)
         );
  OR3_X1 npu_inst_pe_1_4_3_U28 ( .A1(npu_inst_pe_1_4_3_n6), .A2(
        npu_inst_pe_1_4_3_n8), .A3(npu_inst_pe_1_4_3_n5), .ZN(
        npu_inst_pe_1_4_3_n56) );
  OR3_X1 npu_inst_pe_1_4_3_U27 ( .A1(npu_inst_pe_1_4_3_n5), .A2(
        npu_inst_pe_1_4_3_n8), .A3(npu_inst_pe_1_4_3_n7), .ZN(
        npu_inst_pe_1_4_3_n48) );
  INV_X1 npu_inst_pe_1_4_3_U26 ( .A(npu_inst_pe_1_4_3_n5), .ZN(
        npu_inst_pe_1_4_3_n4) );
  OR3_X1 npu_inst_pe_1_4_3_U25 ( .A1(npu_inst_pe_1_4_3_n4), .A2(
        npu_inst_pe_1_4_3_n8), .A3(npu_inst_pe_1_4_3_n7), .ZN(
        npu_inst_pe_1_4_3_n52) );
  OR3_X1 npu_inst_pe_1_4_3_U24 ( .A1(npu_inst_pe_1_4_3_n6), .A2(
        npu_inst_pe_1_4_3_n8), .A3(npu_inst_pe_1_4_3_n4), .ZN(
        npu_inst_pe_1_4_3_n60) );
  NOR2_X1 npu_inst_pe_1_4_3_U23 ( .A1(npu_inst_pe_1_4_3_n60), .A2(
        npu_inst_pe_1_4_3_n3), .ZN(npu_inst_pe_1_4_3_n58) );
  NOR2_X1 npu_inst_pe_1_4_3_U22 ( .A1(npu_inst_pe_1_4_3_n56), .A2(
        npu_inst_pe_1_4_3_n3), .ZN(npu_inst_pe_1_4_3_n54) );
  NOR2_X1 npu_inst_pe_1_4_3_U21 ( .A1(npu_inst_pe_1_4_3_n52), .A2(
        npu_inst_pe_1_4_3_n3), .ZN(npu_inst_pe_1_4_3_n50) );
  NOR2_X1 npu_inst_pe_1_4_3_U20 ( .A1(npu_inst_pe_1_4_3_n48), .A2(
        npu_inst_pe_1_4_3_n3), .ZN(npu_inst_pe_1_4_3_n46) );
  NOR2_X1 npu_inst_pe_1_4_3_U19 ( .A1(npu_inst_pe_1_4_3_n40), .A2(
        npu_inst_pe_1_4_3_n3), .ZN(npu_inst_pe_1_4_3_n38) );
  NOR2_X1 npu_inst_pe_1_4_3_U18 ( .A1(npu_inst_pe_1_4_3_n44), .A2(
        npu_inst_pe_1_4_3_n3), .ZN(npu_inst_pe_1_4_3_n42) );
  BUF_X1 npu_inst_pe_1_4_3_U17 ( .A(npu_inst_n99), .Z(npu_inst_pe_1_4_3_n8) );
  INV_X1 npu_inst_pe_1_4_3_U16 ( .A(npu_inst_n124), .ZN(npu_inst_pe_1_4_3_n12)
         );
  INV_X1 npu_inst_pe_1_4_3_U15 ( .A(npu_inst_pe_1_4_3_n38), .ZN(
        npu_inst_pe_1_4_3_n114) );
  INV_X1 npu_inst_pe_1_4_3_U14 ( .A(npu_inst_pe_1_4_3_n58), .ZN(
        npu_inst_pe_1_4_3_n119) );
  INV_X1 npu_inst_pe_1_4_3_U13 ( .A(npu_inst_pe_1_4_3_n54), .ZN(
        npu_inst_pe_1_4_3_n118) );
  INV_X1 npu_inst_pe_1_4_3_U12 ( .A(npu_inst_pe_1_4_3_n50), .ZN(
        npu_inst_pe_1_4_3_n117) );
  INV_X1 npu_inst_pe_1_4_3_U11 ( .A(npu_inst_pe_1_4_3_n46), .ZN(
        npu_inst_pe_1_4_3_n116) );
  INV_X1 npu_inst_pe_1_4_3_U10 ( .A(npu_inst_pe_1_4_3_n42), .ZN(
        npu_inst_pe_1_4_3_n115) );
  BUF_X1 npu_inst_pe_1_4_3_U9 ( .A(npu_inst_n21), .Z(npu_inst_pe_1_4_3_n2) );
  BUF_X1 npu_inst_pe_1_4_3_U8 ( .A(npu_inst_n21), .Z(npu_inst_pe_1_4_3_n1) );
  BUF_X1 npu_inst_pe_1_4_3_U7 ( .A(npu_inst_pe_1_4_3_n12), .Z(
        npu_inst_pe_1_4_3_n11) );
  BUF_X1 npu_inst_pe_1_4_3_U6 ( .A(npu_inst_pe_1_4_3_n12), .Z(
        npu_inst_pe_1_4_3_n10) );
  BUF_X1 npu_inst_pe_1_4_3_U5 ( .A(npu_inst_pe_1_4_3_n12), .Z(
        npu_inst_pe_1_4_3_n9) );
  NOR2_X1 npu_inst_pe_1_4_3_U4 ( .A1(npu_inst_pe_1_4_3_int_q_weight_0_), .A2(
        npu_inst_pe_1_4_3_n1), .ZN(npu_inst_pe_1_4_3_n76) );
  NOR2_X1 npu_inst_pe_1_4_3_U3 ( .A1(npu_inst_pe_1_4_3_n27), .A2(
        npu_inst_pe_1_4_3_n1), .ZN(npu_inst_pe_1_4_3_n77) );
  FA_X1 npu_inst_pe_1_4_3_sub_67_U2_1 ( .A(npu_inst_pe_1_4_3_int_q_acc_1_), 
        .B(npu_inst_pe_1_4_3_n14), .CI(npu_inst_pe_1_4_3_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_4_3_sub_67_carry_2_), .S(npu_inst_pe_1_4_3_N66) );
  FA_X1 npu_inst_pe_1_4_3_add_69_U1_1 ( .A(npu_inst_pe_1_4_3_int_q_acc_1_), 
        .B(npu_inst_pe_1_4_3_int_data_1_), .CI(
        npu_inst_pe_1_4_3_add_69_carry_1_), .CO(
        npu_inst_pe_1_4_3_add_69_carry_2_), .S(npu_inst_pe_1_4_3_N74) );
  NAND3_X1 npu_inst_pe_1_4_3_U109 ( .A1(npu_inst_pe_1_4_3_n5), .A2(
        npu_inst_pe_1_4_3_n7), .A3(npu_inst_pe_1_4_3_n8), .ZN(
        npu_inst_pe_1_4_3_n44) );
  NAND3_X1 npu_inst_pe_1_4_3_U108 ( .A1(npu_inst_pe_1_4_3_n4), .A2(
        npu_inst_pe_1_4_3_n7), .A3(npu_inst_pe_1_4_3_n8), .ZN(
        npu_inst_pe_1_4_3_n40) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_4_3_n34), .CK(
        npu_inst_pe_1_4_3_net3757), .RN(npu_inst_pe_1_4_3_n9), .Q(
        npu_inst_pe_1_4_3_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_4_3_n35), .CK(
        npu_inst_pe_1_4_3_net3757), .RN(npu_inst_pe_1_4_3_n9), .Q(
        npu_inst_pe_1_4_3_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_4_3_n36), .CK(
        npu_inst_pe_1_4_3_net3757), .RN(npu_inst_pe_1_4_3_n9), .Q(
        npu_inst_pe_1_4_3_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_4_3_n98), .CK(
        npu_inst_pe_1_4_3_net3757), .RN(npu_inst_pe_1_4_3_n9), .Q(
        npu_inst_pe_1_4_3_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_4_3_n99), .CK(
        npu_inst_pe_1_4_3_net3757), .RN(npu_inst_pe_1_4_3_n9), .Q(
        npu_inst_pe_1_4_3_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_4_3_n100), 
        .CK(npu_inst_pe_1_4_3_net3757), .RN(npu_inst_pe_1_4_3_n9), .Q(
        npu_inst_pe_1_4_3_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_4_3_n33), .CK(
        npu_inst_pe_1_4_3_net3757), .RN(npu_inst_pe_1_4_3_n9), .Q(
        npu_inst_pe_1_4_3_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_4_3_n101), 
        .CK(npu_inst_pe_1_4_3_net3757), .RN(npu_inst_pe_1_4_3_n9), .Q(
        npu_inst_pe_1_4_3_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_weight_reg_0_ ( .D(npu_inst_n110), .CK(
        npu_inst_pe_1_4_3_net3763), .RN(npu_inst_pe_1_4_3_n9), .Q(
        npu_inst_pe_1_4_3_int_q_weight_0_), .QN(npu_inst_pe_1_4_3_n27) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_weight_reg_1_ ( .D(npu_inst_n116), .CK(
        npu_inst_pe_1_4_3_net3763), .RN(npu_inst_pe_1_4_3_n9), .Q(
        npu_inst_pe_1_4_3_int_q_weight_1_), .QN(npu_inst_pe_1_4_3_n26) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_4_3_n113), 
        .CK(npu_inst_pe_1_4_3_net3763), .RN(npu_inst_pe_1_4_3_n9), .Q(
        npu_inst_pe_1_4_3_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_4_3_n107), 
        .CK(npu_inst_pe_1_4_3_net3763), .RN(npu_inst_pe_1_4_3_n9), .Q(
        npu_inst_pe_1_4_3_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_4_3_n112), 
        .CK(npu_inst_pe_1_4_3_net3763), .RN(npu_inst_pe_1_4_3_n10), .Q(
        npu_inst_pe_1_4_3_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_4_3_n106), 
        .CK(npu_inst_pe_1_4_3_net3763), .RN(npu_inst_pe_1_4_3_n10), .Q(
        npu_inst_pe_1_4_3_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_4_3_n111), 
        .CK(npu_inst_pe_1_4_3_net3763), .RN(npu_inst_pe_1_4_3_n10), .Q(
        npu_inst_pe_1_4_3_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_4_3_n105), 
        .CK(npu_inst_pe_1_4_3_net3763), .RN(npu_inst_pe_1_4_3_n10), .Q(
        npu_inst_pe_1_4_3_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_4_3_n110), 
        .CK(npu_inst_pe_1_4_3_net3763), .RN(npu_inst_pe_1_4_3_n10), .Q(
        npu_inst_pe_1_4_3_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_4_3_n104), 
        .CK(npu_inst_pe_1_4_3_net3763), .RN(npu_inst_pe_1_4_3_n10), .Q(
        npu_inst_pe_1_4_3_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_4_3_n109), 
        .CK(npu_inst_pe_1_4_3_net3763), .RN(npu_inst_pe_1_4_3_n10), .Q(
        npu_inst_pe_1_4_3_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_4_3_n103), 
        .CK(npu_inst_pe_1_4_3_net3763), .RN(npu_inst_pe_1_4_3_n10), .Q(
        npu_inst_pe_1_4_3_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_4_3_n108), 
        .CK(npu_inst_pe_1_4_3_net3763), .RN(npu_inst_pe_1_4_3_n10), .Q(
        npu_inst_pe_1_4_3_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_4_3_n102), 
        .CK(npu_inst_pe_1_4_3_net3763), .RN(npu_inst_pe_1_4_3_n10), .Q(
        npu_inst_pe_1_4_3_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_4_3_n86), 
        .CK(npu_inst_pe_1_4_3_net3763), .RN(npu_inst_pe_1_4_3_n10), .Q(
        npu_inst_pe_1_4_3_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_4_3_n87), 
        .CK(npu_inst_pe_1_4_3_net3763), .RN(npu_inst_pe_1_4_3_n10), .Q(
        npu_inst_pe_1_4_3_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_4_3_n88), 
        .CK(npu_inst_pe_1_4_3_net3763), .RN(npu_inst_pe_1_4_3_n11), .Q(
        npu_inst_pe_1_4_3_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_4_3_n89), 
        .CK(npu_inst_pe_1_4_3_net3763), .RN(npu_inst_pe_1_4_3_n11), .Q(
        npu_inst_pe_1_4_3_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_4_3_n90), 
        .CK(npu_inst_pe_1_4_3_net3763), .RN(npu_inst_pe_1_4_3_n11), .Q(
        npu_inst_pe_1_4_3_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_4_3_n91), 
        .CK(npu_inst_pe_1_4_3_net3763), .RN(npu_inst_pe_1_4_3_n11), .Q(
        npu_inst_pe_1_4_3_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_4_3_n92), 
        .CK(npu_inst_pe_1_4_3_net3763), .RN(npu_inst_pe_1_4_3_n11), .Q(
        npu_inst_pe_1_4_3_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_4_3_n93), 
        .CK(npu_inst_pe_1_4_3_net3763), .RN(npu_inst_pe_1_4_3_n11), .Q(
        npu_inst_pe_1_4_3_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_4_3_n94), 
        .CK(npu_inst_pe_1_4_3_net3763), .RN(npu_inst_pe_1_4_3_n11), .Q(
        npu_inst_pe_1_4_3_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_4_3_n95), 
        .CK(npu_inst_pe_1_4_3_net3763), .RN(npu_inst_pe_1_4_3_n11), .Q(
        npu_inst_pe_1_4_3_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_4_3_n96), 
        .CK(npu_inst_pe_1_4_3_net3763), .RN(npu_inst_pe_1_4_3_n11), .Q(
        npu_inst_pe_1_4_3_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_4_3_n97), 
        .CK(npu_inst_pe_1_4_3_net3763), .RN(npu_inst_pe_1_4_3_n11), .Q(
        npu_inst_pe_1_4_3_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_4_3_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_4_3_N84), .SE(1'b0), .GCK(npu_inst_pe_1_4_3_net3757) );
  CLKGATETST_X1 npu_inst_pe_1_4_3_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n63), .SE(1'b0), .GCK(npu_inst_pe_1_4_3_net3763) );
  MUX2_X1 npu_inst_pe_1_4_4_U162 ( .A(npu_inst_pe_1_4_4_n32), .B(
        npu_inst_pe_1_4_4_n29), .S(npu_inst_pe_1_4_4_n8), .Z(
        npu_inst_pe_1_4_4_N93) );
  MUX2_X1 npu_inst_pe_1_4_4_U161 ( .A(npu_inst_pe_1_4_4_n31), .B(
        npu_inst_pe_1_4_4_n30), .S(npu_inst_pe_1_4_4_n6), .Z(
        npu_inst_pe_1_4_4_n32) );
  MUX2_X1 npu_inst_pe_1_4_4_U160 ( .A(npu_inst_pe_1_4_4_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_4_4_int_q_reg_v_1__0_), .S(npu_inst_pe_1_4_4_n4), .Z(
        npu_inst_pe_1_4_4_n31) );
  MUX2_X1 npu_inst_pe_1_4_4_U159 ( .A(npu_inst_pe_1_4_4_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_4_4_int_q_reg_v_3__0_), .S(npu_inst_pe_1_4_4_n4), .Z(
        npu_inst_pe_1_4_4_n30) );
  MUX2_X1 npu_inst_pe_1_4_4_U158 ( .A(npu_inst_pe_1_4_4_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_4_4_int_q_reg_v_5__0_), .S(npu_inst_pe_1_4_4_n4), .Z(
        npu_inst_pe_1_4_4_n29) );
  MUX2_X1 npu_inst_pe_1_4_4_U157 ( .A(npu_inst_pe_1_4_4_n28), .B(
        npu_inst_pe_1_4_4_n23), .S(npu_inst_pe_1_4_4_n8), .Z(
        npu_inst_pe_1_4_4_N94) );
  MUX2_X1 npu_inst_pe_1_4_4_U156 ( .A(npu_inst_pe_1_4_4_n25), .B(
        npu_inst_pe_1_4_4_n24), .S(npu_inst_pe_1_4_4_n6), .Z(
        npu_inst_pe_1_4_4_n28) );
  MUX2_X1 npu_inst_pe_1_4_4_U155 ( .A(npu_inst_pe_1_4_4_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_4_4_int_q_reg_v_1__1_), .S(npu_inst_pe_1_4_4_n4), .Z(
        npu_inst_pe_1_4_4_n25) );
  MUX2_X1 npu_inst_pe_1_4_4_U154 ( .A(npu_inst_pe_1_4_4_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_4_4_int_q_reg_v_3__1_), .S(npu_inst_pe_1_4_4_n4), .Z(
        npu_inst_pe_1_4_4_n24) );
  MUX2_X1 npu_inst_pe_1_4_4_U153 ( .A(npu_inst_pe_1_4_4_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_4_4_int_q_reg_v_5__1_), .S(npu_inst_pe_1_4_4_n4), .Z(
        npu_inst_pe_1_4_4_n23) );
  MUX2_X1 npu_inst_pe_1_4_4_U152 ( .A(npu_inst_pe_1_4_4_n22), .B(
        npu_inst_pe_1_4_4_n19), .S(npu_inst_pe_1_4_4_n8), .Z(
        npu_inst_int_data_x_4__4__1_) );
  MUX2_X1 npu_inst_pe_1_4_4_U151 ( .A(npu_inst_pe_1_4_4_n21), .B(
        npu_inst_pe_1_4_4_n20), .S(npu_inst_pe_1_4_4_n6), .Z(
        npu_inst_pe_1_4_4_n22) );
  MUX2_X1 npu_inst_pe_1_4_4_U150 ( .A(npu_inst_pe_1_4_4_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_4_4_int_q_reg_h_1__1_), .S(npu_inst_pe_1_4_4_n4), .Z(
        npu_inst_pe_1_4_4_n21) );
  MUX2_X1 npu_inst_pe_1_4_4_U149 ( .A(npu_inst_pe_1_4_4_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_4_4_int_q_reg_h_3__1_), .S(npu_inst_pe_1_4_4_n4), .Z(
        npu_inst_pe_1_4_4_n20) );
  MUX2_X1 npu_inst_pe_1_4_4_U148 ( .A(npu_inst_pe_1_4_4_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_4_4_int_q_reg_h_5__1_), .S(npu_inst_pe_1_4_4_n4), .Z(
        npu_inst_pe_1_4_4_n19) );
  MUX2_X1 npu_inst_pe_1_4_4_U147 ( .A(npu_inst_pe_1_4_4_n18), .B(
        npu_inst_pe_1_4_4_n15), .S(npu_inst_pe_1_4_4_n8), .Z(
        npu_inst_int_data_x_4__4__0_) );
  MUX2_X1 npu_inst_pe_1_4_4_U146 ( .A(npu_inst_pe_1_4_4_n17), .B(
        npu_inst_pe_1_4_4_n16), .S(npu_inst_pe_1_4_4_n6), .Z(
        npu_inst_pe_1_4_4_n18) );
  MUX2_X1 npu_inst_pe_1_4_4_U145 ( .A(npu_inst_pe_1_4_4_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_4_4_int_q_reg_h_1__0_), .S(npu_inst_pe_1_4_4_n4), .Z(
        npu_inst_pe_1_4_4_n17) );
  MUX2_X1 npu_inst_pe_1_4_4_U144 ( .A(npu_inst_pe_1_4_4_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_4_4_int_q_reg_h_3__0_), .S(npu_inst_pe_1_4_4_n4), .Z(
        npu_inst_pe_1_4_4_n16) );
  MUX2_X1 npu_inst_pe_1_4_4_U143 ( .A(npu_inst_pe_1_4_4_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_4_4_int_q_reg_h_5__0_), .S(npu_inst_pe_1_4_4_n4), .Z(
        npu_inst_pe_1_4_4_n15) );
  XOR2_X1 npu_inst_pe_1_4_4_U142 ( .A(npu_inst_pe_1_4_4_int_data_0_), .B(
        npu_inst_pe_1_4_4_int_q_acc_0_), .Z(npu_inst_pe_1_4_4_N73) );
  AND2_X1 npu_inst_pe_1_4_4_U141 ( .A1(npu_inst_pe_1_4_4_int_q_acc_0_), .A2(
        npu_inst_pe_1_4_4_int_data_0_), .ZN(npu_inst_pe_1_4_4_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_4_4_U140 ( .A(npu_inst_pe_1_4_4_int_q_acc_0_), .B(
        npu_inst_pe_1_4_4_n13), .ZN(npu_inst_pe_1_4_4_N65) );
  OR2_X1 npu_inst_pe_1_4_4_U139 ( .A1(npu_inst_pe_1_4_4_n13), .A2(
        npu_inst_pe_1_4_4_int_q_acc_0_), .ZN(npu_inst_pe_1_4_4_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_4_4_U138 ( .A(npu_inst_pe_1_4_4_int_q_acc_2_), .B(
        npu_inst_pe_1_4_4_add_69_carry_2_), .Z(npu_inst_pe_1_4_4_N75) );
  AND2_X1 npu_inst_pe_1_4_4_U137 ( .A1(npu_inst_pe_1_4_4_add_69_carry_2_), 
        .A2(npu_inst_pe_1_4_4_int_q_acc_2_), .ZN(
        npu_inst_pe_1_4_4_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_4_4_U136 ( .A(npu_inst_pe_1_4_4_int_q_acc_3_), .B(
        npu_inst_pe_1_4_4_add_69_carry_3_), .Z(npu_inst_pe_1_4_4_N76) );
  AND2_X1 npu_inst_pe_1_4_4_U135 ( .A1(npu_inst_pe_1_4_4_add_69_carry_3_), 
        .A2(npu_inst_pe_1_4_4_int_q_acc_3_), .ZN(
        npu_inst_pe_1_4_4_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_4_4_U134 ( .A(npu_inst_pe_1_4_4_int_q_acc_4_), .B(
        npu_inst_pe_1_4_4_add_69_carry_4_), .Z(npu_inst_pe_1_4_4_N77) );
  AND2_X1 npu_inst_pe_1_4_4_U133 ( .A1(npu_inst_pe_1_4_4_add_69_carry_4_), 
        .A2(npu_inst_pe_1_4_4_int_q_acc_4_), .ZN(
        npu_inst_pe_1_4_4_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_4_4_U132 ( .A(npu_inst_pe_1_4_4_int_q_acc_5_), .B(
        npu_inst_pe_1_4_4_add_69_carry_5_), .Z(npu_inst_pe_1_4_4_N78) );
  AND2_X1 npu_inst_pe_1_4_4_U131 ( .A1(npu_inst_pe_1_4_4_add_69_carry_5_), 
        .A2(npu_inst_pe_1_4_4_int_q_acc_5_), .ZN(
        npu_inst_pe_1_4_4_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_4_4_U130 ( .A(npu_inst_pe_1_4_4_int_q_acc_6_), .B(
        npu_inst_pe_1_4_4_add_69_carry_6_), .Z(npu_inst_pe_1_4_4_N79) );
  AND2_X1 npu_inst_pe_1_4_4_U129 ( .A1(npu_inst_pe_1_4_4_add_69_carry_6_), 
        .A2(npu_inst_pe_1_4_4_int_q_acc_6_), .ZN(
        npu_inst_pe_1_4_4_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_4_4_U128 ( .A(npu_inst_pe_1_4_4_int_q_acc_7_), .B(
        npu_inst_pe_1_4_4_add_69_carry_7_), .Z(npu_inst_pe_1_4_4_N80) );
  XNOR2_X1 npu_inst_pe_1_4_4_U127 ( .A(npu_inst_pe_1_4_4_sub_67_carry_2_), .B(
        npu_inst_pe_1_4_4_int_q_acc_2_), .ZN(npu_inst_pe_1_4_4_N67) );
  OR2_X1 npu_inst_pe_1_4_4_U126 ( .A1(npu_inst_pe_1_4_4_int_q_acc_2_), .A2(
        npu_inst_pe_1_4_4_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_4_4_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_4_4_U125 ( .A(npu_inst_pe_1_4_4_sub_67_carry_3_), .B(
        npu_inst_pe_1_4_4_int_q_acc_3_), .ZN(npu_inst_pe_1_4_4_N68) );
  OR2_X1 npu_inst_pe_1_4_4_U124 ( .A1(npu_inst_pe_1_4_4_int_q_acc_3_), .A2(
        npu_inst_pe_1_4_4_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_4_4_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_4_4_U123 ( .A(npu_inst_pe_1_4_4_sub_67_carry_4_), .B(
        npu_inst_pe_1_4_4_int_q_acc_4_), .ZN(npu_inst_pe_1_4_4_N69) );
  OR2_X1 npu_inst_pe_1_4_4_U122 ( .A1(npu_inst_pe_1_4_4_int_q_acc_4_), .A2(
        npu_inst_pe_1_4_4_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_4_4_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_4_4_U121 ( .A(npu_inst_pe_1_4_4_sub_67_carry_5_), .B(
        npu_inst_pe_1_4_4_int_q_acc_5_), .ZN(npu_inst_pe_1_4_4_N70) );
  OR2_X1 npu_inst_pe_1_4_4_U120 ( .A1(npu_inst_pe_1_4_4_int_q_acc_5_), .A2(
        npu_inst_pe_1_4_4_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_4_4_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_4_4_U119 ( .A(npu_inst_pe_1_4_4_sub_67_carry_6_), .B(
        npu_inst_pe_1_4_4_int_q_acc_6_), .ZN(npu_inst_pe_1_4_4_N71) );
  OR2_X1 npu_inst_pe_1_4_4_U118 ( .A1(npu_inst_pe_1_4_4_int_q_acc_6_), .A2(
        npu_inst_pe_1_4_4_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_4_4_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_4_4_U117 ( .A(npu_inst_pe_1_4_4_int_q_acc_7_), .B(
        npu_inst_pe_1_4_4_sub_67_carry_7_), .ZN(npu_inst_pe_1_4_4_N72) );
  INV_X1 npu_inst_pe_1_4_4_U116 ( .A(npu_inst_n77), .ZN(npu_inst_pe_1_4_4_n7)
         );
  INV_X1 npu_inst_pe_1_4_4_U115 ( .A(npu_inst_pe_1_4_4_n7), .ZN(
        npu_inst_pe_1_4_4_n6) );
  INV_X1 npu_inst_pe_1_4_4_U114 ( .A(npu_inst_n55), .ZN(npu_inst_pe_1_4_4_n3)
         );
  AOI22_X1 npu_inst_pe_1_4_4_U113 ( .A1(npu_inst_int_data_y_5__4__0_), .A2(
        npu_inst_pe_1_4_4_n58), .B1(npu_inst_pe_1_4_4_n119), .B2(
        npu_inst_pe_1_4_4_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_4_4_n57) );
  INV_X1 npu_inst_pe_1_4_4_U112 ( .A(npu_inst_pe_1_4_4_n57), .ZN(
        npu_inst_pe_1_4_4_n108) );
  AOI22_X1 npu_inst_pe_1_4_4_U111 ( .A1(npu_inst_int_data_y_5__4__0_), .A2(
        npu_inst_pe_1_4_4_n54), .B1(npu_inst_pe_1_4_4_n118), .B2(
        npu_inst_pe_1_4_4_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_4_4_n53) );
  INV_X1 npu_inst_pe_1_4_4_U110 ( .A(npu_inst_pe_1_4_4_n53), .ZN(
        npu_inst_pe_1_4_4_n109) );
  AOI22_X1 npu_inst_pe_1_4_4_U107 ( .A1(npu_inst_int_data_y_5__4__0_), .A2(
        npu_inst_pe_1_4_4_n50), .B1(npu_inst_pe_1_4_4_n117), .B2(
        npu_inst_pe_1_4_4_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_4_4_n49) );
  INV_X1 npu_inst_pe_1_4_4_U106 ( .A(npu_inst_pe_1_4_4_n49), .ZN(
        npu_inst_pe_1_4_4_n110) );
  AOI22_X1 npu_inst_pe_1_4_4_U105 ( .A1(npu_inst_int_data_y_5__4__0_), .A2(
        npu_inst_pe_1_4_4_n46), .B1(npu_inst_pe_1_4_4_n116), .B2(
        npu_inst_pe_1_4_4_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_4_4_n45) );
  INV_X1 npu_inst_pe_1_4_4_U104 ( .A(npu_inst_pe_1_4_4_n45), .ZN(
        npu_inst_pe_1_4_4_n111) );
  AOI22_X1 npu_inst_pe_1_4_4_U103 ( .A1(npu_inst_int_data_y_5__4__0_), .A2(
        npu_inst_pe_1_4_4_n42), .B1(npu_inst_pe_1_4_4_n115), .B2(
        npu_inst_pe_1_4_4_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_4_4_n41) );
  INV_X1 npu_inst_pe_1_4_4_U102 ( .A(npu_inst_pe_1_4_4_n41), .ZN(
        npu_inst_pe_1_4_4_n112) );
  AOI22_X1 npu_inst_pe_1_4_4_U101 ( .A1(npu_inst_int_data_y_5__4__1_), .A2(
        npu_inst_pe_1_4_4_n58), .B1(npu_inst_pe_1_4_4_n119), .B2(
        npu_inst_pe_1_4_4_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_4_4_n59) );
  INV_X1 npu_inst_pe_1_4_4_U100 ( .A(npu_inst_pe_1_4_4_n59), .ZN(
        npu_inst_pe_1_4_4_n102) );
  AOI22_X1 npu_inst_pe_1_4_4_U99 ( .A1(npu_inst_int_data_y_5__4__1_), .A2(
        npu_inst_pe_1_4_4_n54), .B1(npu_inst_pe_1_4_4_n118), .B2(
        npu_inst_pe_1_4_4_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_4_4_n55) );
  INV_X1 npu_inst_pe_1_4_4_U98 ( .A(npu_inst_pe_1_4_4_n55), .ZN(
        npu_inst_pe_1_4_4_n103) );
  AOI22_X1 npu_inst_pe_1_4_4_U97 ( .A1(npu_inst_int_data_y_5__4__1_), .A2(
        npu_inst_pe_1_4_4_n50), .B1(npu_inst_pe_1_4_4_n117), .B2(
        npu_inst_pe_1_4_4_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_4_4_n51) );
  INV_X1 npu_inst_pe_1_4_4_U96 ( .A(npu_inst_pe_1_4_4_n51), .ZN(
        npu_inst_pe_1_4_4_n104) );
  AOI22_X1 npu_inst_pe_1_4_4_U95 ( .A1(npu_inst_int_data_y_5__4__1_), .A2(
        npu_inst_pe_1_4_4_n46), .B1(npu_inst_pe_1_4_4_n116), .B2(
        npu_inst_pe_1_4_4_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_4_4_n47) );
  INV_X1 npu_inst_pe_1_4_4_U94 ( .A(npu_inst_pe_1_4_4_n47), .ZN(
        npu_inst_pe_1_4_4_n105) );
  AOI22_X1 npu_inst_pe_1_4_4_U93 ( .A1(npu_inst_int_data_y_5__4__1_), .A2(
        npu_inst_pe_1_4_4_n42), .B1(npu_inst_pe_1_4_4_n115), .B2(
        npu_inst_pe_1_4_4_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_4_4_n43) );
  INV_X1 npu_inst_pe_1_4_4_U92 ( .A(npu_inst_pe_1_4_4_n43), .ZN(
        npu_inst_pe_1_4_4_n106) );
  AOI22_X1 npu_inst_pe_1_4_4_U91 ( .A1(npu_inst_pe_1_4_4_n38), .A2(
        npu_inst_int_data_y_5__4__1_), .B1(npu_inst_pe_1_4_4_n114), .B2(
        npu_inst_pe_1_4_4_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_4_4_n39) );
  INV_X1 npu_inst_pe_1_4_4_U90 ( .A(npu_inst_pe_1_4_4_n39), .ZN(
        npu_inst_pe_1_4_4_n107) );
  AOI22_X1 npu_inst_pe_1_4_4_U89 ( .A1(npu_inst_pe_1_4_4_n38), .A2(
        npu_inst_int_data_y_5__4__0_), .B1(npu_inst_pe_1_4_4_n114), .B2(
        npu_inst_pe_1_4_4_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_4_4_n37) );
  INV_X1 npu_inst_pe_1_4_4_U88 ( .A(npu_inst_pe_1_4_4_n37), .ZN(
        npu_inst_pe_1_4_4_n113) );
  NOR3_X1 npu_inst_pe_1_4_4_U87 ( .A1(npu_inst_pe_1_4_4_n26), .A2(npu_inst_n55), .A3(npu_inst_int_ckg[27]), .ZN(npu_inst_pe_1_4_4_n85) );
  OR2_X1 npu_inst_pe_1_4_4_U86 ( .A1(npu_inst_pe_1_4_4_n85), .A2(
        npu_inst_pe_1_4_4_n2), .ZN(npu_inst_pe_1_4_4_N84) );
  NAND2_X1 npu_inst_pe_1_4_4_U85 ( .A1(npu_inst_pe_1_4_4_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_4_4_n60), .ZN(npu_inst_pe_1_4_4_n74) );
  OAI21_X1 npu_inst_pe_1_4_4_U84 ( .B1(npu_inst_pe_1_4_4_n63), .B2(
        npu_inst_pe_1_4_4_n60), .A(npu_inst_pe_1_4_4_n74), .ZN(
        npu_inst_pe_1_4_4_n97) );
  NAND2_X1 npu_inst_pe_1_4_4_U83 ( .A1(npu_inst_pe_1_4_4_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_4_4_n60), .ZN(npu_inst_pe_1_4_4_n73) );
  OAI21_X1 npu_inst_pe_1_4_4_U82 ( .B1(npu_inst_pe_1_4_4_n61), .B2(
        npu_inst_pe_1_4_4_n60), .A(npu_inst_pe_1_4_4_n73), .ZN(
        npu_inst_pe_1_4_4_n96) );
  NAND2_X1 npu_inst_pe_1_4_4_U81 ( .A1(npu_inst_pe_1_4_4_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_4_4_n56), .ZN(npu_inst_pe_1_4_4_n72) );
  OAI21_X1 npu_inst_pe_1_4_4_U80 ( .B1(npu_inst_pe_1_4_4_n63), .B2(
        npu_inst_pe_1_4_4_n56), .A(npu_inst_pe_1_4_4_n72), .ZN(
        npu_inst_pe_1_4_4_n95) );
  NAND2_X1 npu_inst_pe_1_4_4_U79 ( .A1(npu_inst_pe_1_4_4_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_4_4_n56), .ZN(npu_inst_pe_1_4_4_n71) );
  OAI21_X1 npu_inst_pe_1_4_4_U78 ( .B1(npu_inst_pe_1_4_4_n61), .B2(
        npu_inst_pe_1_4_4_n56), .A(npu_inst_pe_1_4_4_n71), .ZN(
        npu_inst_pe_1_4_4_n94) );
  NAND2_X1 npu_inst_pe_1_4_4_U77 ( .A1(npu_inst_pe_1_4_4_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_4_4_n52), .ZN(npu_inst_pe_1_4_4_n70) );
  OAI21_X1 npu_inst_pe_1_4_4_U76 ( .B1(npu_inst_pe_1_4_4_n63), .B2(
        npu_inst_pe_1_4_4_n52), .A(npu_inst_pe_1_4_4_n70), .ZN(
        npu_inst_pe_1_4_4_n93) );
  NAND2_X1 npu_inst_pe_1_4_4_U75 ( .A1(npu_inst_pe_1_4_4_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_4_4_n52), .ZN(npu_inst_pe_1_4_4_n69) );
  OAI21_X1 npu_inst_pe_1_4_4_U74 ( .B1(npu_inst_pe_1_4_4_n61), .B2(
        npu_inst_pe_1_4_4_n52), .A(npu_inst_pe_1_4_4_n69), .ZN(
        npu_inst_pe_1_4_4_n92) );
  NAND2_X1 npu_inst_pe_1_4_4_U73 ( .A1(npu_inst_pe_1_4_4_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_4_4_n48), .ZN(npu_inst_pe_1_4_4_n68) );
  OAI21_X1 npu_inst_pe_1_4_4_U72 ( .B1(npu_inst_pe_1_4_4_n63), .B2(
        npu_inst_pe_1_4_4_n48), .A(npu_inst_pe_1_4_4_n68), .ZN(
        npu_inst_pe_1_4_4_n91) );
  NAND2_X1 npu_inst_pe_1_4_4_U71 ( .A1(npu_inst_pe_1_4_4_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_4_4_n48), .ZN(npu_inst_pe_1_4_4_n67) );
  OAI21_X1 npu_inst_pe_1_4_4_U70 ( .B1(npu_inst_pe_1_4_4_n61), .B2(
        npu_inst_pe_1_4_4_n48), .A(npu_inst_pe_1_4_4_n67), .ZN(
        npu_inst_pe_1_4_4_n90) );
  NAND2_X1 npu_inst_pe_1_4_4_U69 ( .A1(npu_inst_pe_1_4_4_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_4_4_n44), .ZN(npu_inst_pe_1_4_4_n66) );
  OAI21_X1 npu_inst_pe_1_4_4_U68 ( .B1(npu_inst_pe_1_4_4_n63), .B2(
        npu_inst_pe_1_4_4_n44), .A(npu_inst_pe_1_4_4_n66), .ZN(
        npu_inst_pe_1_4_4_n89) );
  NAND2_X1 npu_inst_pe_1_4_4_U67 ( .A1(npu_inst_pe_1_4_4_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_4_4_n44), .ZN(npu_inst_pe_1_4_4_n65) );
  OAI21_X1 npu_inst_pe_1_4_4_U66 ( .B1(npu_inst_pe_1_4_4_n61), .B2(
        npu_inst_pe_1_4_4_n44), .A(npu_inst_pe_1_4_4_n65), .ZN(
        npu_inst_pe_1_4_4_n88) );
  NAND2_X1 npu_inst_pe_1_4_4_U65 ( .A1(npu_inst_pe_1_4_4_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_4_4_n40), .ZN(npu_inst_pe_1_4_4_n64) );
  OAI21_X1 npu_inst_pe_1_4_4_U64 ( .B1(npu_inst_pe_1_4_4_n63), .B2(
        npu_inst_pe_1_4_4_n40), .A(npu_inst_pe_1_4_4_n64), .ZN(
        npu_inst_pe_1_4_4_n87) );
  NAND2_X1 npu_inst_pe_1_4_4_U63 ( .A1(npu_inst_pe_1_4_4_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_4_4_n40), .ZN(npu_inst_pe_1_4_4_n62) );
  OAI21_X1 npu_inst_pe_1_4_4_U62 ( .B1(npu_inst_pe_1_4_4_n61), .B2(
        npu_inst_pe_1_4_4_n40), .A(npu_inst_pe_1_4_4_n62), .ZN(
        npu_inst_pe_1_4_4_n86) );
  AND2_X1 npu_inst_pe_1_4_4_U61 ( .A1(npu_inst_pe_1_4_4_N93), .A2(npu_inst_n55), .ZN(npu_inst_int_data_y_4__4__0_) );
  AND2_X1 npu_inst_pe_1_4_4_U60 ( .A1(npu_inst_n55), .A2(npu_inst_pe_1_4_4_N94), .ZN(npu_inst_int_data_y_4__4__1_) );
  AND2_X1 npu_inst_pe_1_4_4_U59 ( .A1(npu_inst_pe_1_4_4_int_q_acc_0_), .A2(
        npu_inst_pe_1_4_4_n1), .ZN(npu_inst_int_data_res_4__4__0_) );
  AND2_X1 npu_inst_pe_1_4_4_U58 ( .A1(npu_inst_pe_1_4_4_n2), .A2(
        npu_inst_pe_1_4_4_int_q_acc_7_), .ZN(npu_inst_int_data_res_4__4__7_)
         );
  AND2_X1 npu_inst_pe_1_4_4_U57 ( .A1(npu_inst_pe_1_4_4_int_q_acc_1_), .A2(
        npu_inst_pe_1_4_4_n1), .ZN(npu_inst_int_data_res_4__4__1_) );
  AND2_X1 npu_inst_pe_1_4_4_U56 ( .A1(npu_inst_pe_1_4_4_int_q_acc_2_), .A2(
        npu_inst_pe_1_4_4_n1), .ZN(npu_inst_int_data_res_4__4__2_) );
  AND2_X1 npu_inst_pe_1_4_4_U55 ( .A1(npu_inst_pe_1_4_4_int_q_acc_3_), .A2(
        npu_inst_pe_1_4_4_n2), .ZN(npu_inst_int_data_res_4__4__3_) );
  AND2_X1 npu_inst_pe_1_4_4_U54 ( .A1(npu_inst_pe_1_4_4_int_q_acc_4_), .A2(
        npu_inst_pe_1_4_4_n2), .ZN(npu_inst_int_data_res_4__4__4_) );
  AND2_X1 npu_inst_pe_1_4_4_U53 ( .A1(npu_inst_pe_1_4_4_int_q_acc_5_), .A2(
        npu_inst_pe_1_4_4_n2), .ZN(npu_inst_int_data_res_4__4__5_) );
  AND2_X1 npu_inst_pe_1_4_4_U52 ( .A1(npu_inst_pe_1_4_4_int_q_acc_6_), .A2(
        npu_inst_pe_1_4_4_n2), .ZN(npu_inst_int_data_res_4__4__6_) );
  AOI222_X1 npu_inst_pe_1_4_4_U51 ( .A1(npu_inst_int_data_res_5__4__0_), .A2(
        npu_inst_pe_1_4_4_n1), .B1(npu_inst_pe_1_4_4_N73), .B2(
        npu_inst_pe_1_4_4_n76), .C1(npu_inst_pe_1_4_4_N65), .C2(
        npu_inst_pe_1_4_4_n77), .ZN(npu_inst_pe_1_4_4_n84) );
  INV_X1 npu_inst_pe_1_4_4_U50 ( .A(npu_inst_pe_1_4_4_n84), .ZN(
        npu_inst_pe_1_4_4_n101) );
  AOI222_X1 npu_inst_pe_1_4_4_U49 ( .A1(npu_inst_int_data_res_5__4__7_), .A2(
        npu_inst_pe_1_4_4_n1), .B1(npu_inst_pe_1_4_4_N80), .B2(
        npu_inst_pe_1_4_4_n76), .C1(npu_inst_pe_1_4_4_N72), .C2(
        npu_inst_pe_1_4_4_n77), .ZN(npu_inst_pe_1_4_4_n75) );
  INV_X1 npu_inst_pe_1_4_4_U48 ( .A(npu_inst_pe_1_4_4_n75), .ZN(
        npu_inst_pe_1_4_4_n33) );
  AOI222_X1 npu_inst_pe_1_4_4_U47 ( .A1(npu_inst_int_data_res_5__4__1_), .A2(
        npu_inst_pe_1_4_4_n1), .B1(npu_inst_pe_1_4_4_N74), .B2(
        npu_inst_pe_1_4_4_n76), .C1(npu_inst_pe_1_4_4_N66), .C2(
        npu_inst_pe_1_4_4_n77), .ZN(npu_inst_pe_1_4_4_n83) );
  INV_X1 npu_inst_pe_1_4_4_U46 ( .A(npu_inst_pe_1_4_4_n83), .ZN(
        npu_inst_pe_1_4_4_n100) );
  AOI222_X1 npu_inst_pe_1_4_4_U45 ( .A1(npu_inst_int_data_res_5__4__2_), .A2(
        npu_inst_pe_1_4_4_n1), .B1(npu_inst_pe_1_4_4_N75), .B2(
        npu_inst_pe_1_4_4_n76), .C1(npu_inst_pe_1_4_4_N67), .C2(
        npu_inst_pe_1_4_4_n77), .ZN(npu_inst_pe_1_4_4_n82) );
  INV_X1 npu_inst_pe_1_4_4_U44 ( .A(npu_inst_pe_1_4_4_n82), .ZN(
        npu_inst_pe_1_4_4_n99) );
  AOI222_X1 npu_inst_pe_1_4_4_U43 ( .A1(npu_inst_int_data_res_5__4__3_), .A2(
        npu_inst_pe_1_4_4_n1), .B1(npu_inst_pe_1_4_4_N76), .B2(
        npu_inst_pe_1_4_4_n76), .C1(npu_inst_pe_1_4_4_N68), .C2(
        npu_inst_pe_1_4_4_n77), .ZN(npu_inst_pe_1_4_4_n81) );
  INV_X1 npu_inst_pe_1_4_4_U42 ( .A(npu_inst_pe_1_4_4_n81), .ZN(
        npu_inst_pe_1_4_4_n98) );
  AOI222_X1 npu_inst_pe_1_4_4_U41 ( .A1(npu_inst_int_data_res_5__4__4_), .A2(
        npu_inst_pe_1_4_4_n1), .B1(npu_inst_pe_1_4_4_N77), .B2(
        npu_inst_pe_1_4_4_n76), .C1(npu_inst_pe_1_4_4_N69), .C2(
        npu_inst_pe_1_4_4_n77), .ZN(npu_inst_pe_1_4_4_n80) );
  INV_X1 npu_inst_pe_1_4_4_U40 ( .A(npu_inst_pe_1_4_4_n80), .ZN(
        npu_inst_pe_1_4_4_n36) );
  AOI222_X1 npu_inst_pe_1_4_4_U39 ( .A1(npu_inst_int_data_res_5__4__5_), .A2(
        npu_inst_pe_1_4_4_n1), .B1(npu_inst_pe_1_4_4_N78), .B2(
        npu_inst_pe_1_4_4_n76), .C1(npu_inst_pe_1_4_4_N70), .C2(
        npu_inst_pe_1_4_4_n77), .ZN(npu_inst_pe_1_4_4_n79) );
  INV_X1 npu_inst_pe_1_4_4_U38 ( .A(npu_inst_pe_1_4_4_n79), .ZN(
        npu_inst_pe_1_4_4_n35) );
  AOI222_X1 npu_inst_pe_1_4_4_U37 ( .A1(npu_inst_int_data_res_5__4__6_), .A2(
        npu_inst_pe_1_4_4_n1), .B1(npu_inst_pe_1_4_4_N79), .B2(
        npu_inst_pe_1_4_4_n76), .C1(npu_inst_pe_1_4_4_N71), .C2(
        npu_inst_pe_1_4_4_n77), .ZN(npu_inst_pe_1_4_4_n78) );
  INV_X1 npu_inst_pe_1_4_4_U36 ( .A(npu_inst_pe_1_4_4_n78), .ZN(
        npu_inst_pe_1_4_4_n34) );
  INV_X1 npu_inst_pe_1_4_4_U35 ( .A(npu_inst_pe_1_4_4_int_data_1_), .ZN(
        npu_inst_pe_1_4_4_n14) );
  AND2_X1 npu_inst_pe_1_4_4_U34 ( .A1(npu_inst_int_data_x_4__4__1_), .A2(
        npu_inst_pe_1_4_4_int_q_weight_1_), .ZN(npu_inst_pe_1_4_4_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_4_4_U33 ( .A1(npu_inst_int_data_x_4__4__0_), .A2(
        npu_inst_pe_1_4_4_int_q_weight_1_), .ZN(npu_inst_pe_1_4_4_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_4_4_U32 ( .A1(npu_inst_n55), .A2(
        npu_inst_int_data_y_5__4__1_), .B1(npu_inst_pe_1_4_4_n3), .B2(
        npu_inst_int_data_x_4__5__1_), .ZN(npu_inst_pe_1_4_4_n63) );
  AOI22_X1 npu_inst_pe_1_4_4_U31 ( .A1(npu_inst_n55), .A2(
        npu_inst_int_data_y_5__4__0_), .B1(npu_inst_pe_1_4_4_n3), .B2(
        npu_inst_int_data_x_4__5__0_), .ZN(npu_inst_pe_1_4_4_n61) );
  INV_X1 npu_inst_pe_1_4_4_U30 ( .A(npu_inst_pe_1_4_4_int_data_0_), .ZN(
        npu_inst_pe_1_4_4_n13) );
  INV_X1 npu_inst_pe_1_4_4_U29 ( .A(npu_inst_n69), .ZN(npu_inst_pe_1_4_4_n5)
         );
  OR3_X1 npu_inst_pe_1_4_4_U28 ( .A1(npu_inst_pe_1_4_4_n6), .A2(
        npu_inst_pe_1_4_4_n8), .A3(npu_inst_pe_1_4_4_n5), .ZN(
        npu_inst_pe_1_4_4_n56) );
  OR3_X1 npu_inst_pe_1_4_4_U27 ( .A1(npu_inst_pe_1_4_4_n5), .A2(
        npu_inst_pe_1_4_4_n8), .A3(npu_inst_pe_1_4_4_n7), .ZN(
        npu_inst_pe_1_4_4_n48) );
  INV_X1 npu_inst_pe_1_4_4_U26 ( .A(npu_inst_pe_1_4_4_n5), .ZN(
        npu_inst_pe_1_4_4_n4) );
  OR3_X1 npu_inst_pe_1_4_4_U25 ( .A1(npu_inst_pe_1_4_4_n4), .A2(
        npu_inst_pe_1_4_4_n8), .A3(npu_inst_pe_1_4_4_n7), .ZN(
        npu_inst_pe_1_4_4_n52) );
  OR3_X1 npu_inst_pe_1_4_4_U24 ( .A1(npu_inst_pe_1_4_4_n6), .A2(
        npu_inst_pe_1_4_4_n8), .A3(npu_inst_pe_1_4_4_n4), .ZN(
        npu_inst_pe_1_4_4_n60) );
  NOR2_X1 npu_inst_pe_1_4_4_U23 ( .A1(npu_inst_pe_1_4_4_n60), .A2(
        npu_inst_pe_1_4_4_n3), .ZN(npu_inst_pe_1_4_4_n58) );
  NOR2_X1 npu_inst_pe_1_4_4_U22 ( .A1(npu_inst_pe_1_4_4_n56), .A2(
        npu_inst_pe_1_4_4_n3), .ZN(npu_inst_pe_1_4_4_n54) );
  NOR2_X1 npu_inst_pe_1_4_4_U21 ( .A1(npu_inst_pe_1_4_4_n52), .A2(
        npu_inst_pe_1_4_4_n3), .ZN(npu_inst_pe_1_4_4_n50) );
  NOR2_X1 npu_inst_pe_1_4_4_U20 ( .A1(npu_inst_pe_1_4_4_n48), .A2(
        npu_inst_pe_1_4_4_n3), .ZN(npu_inst_pe_1_4_4_n46) );
  NOR2_X1 npu_inst_pe_1_4_4_U19 ( .A1(npu_inst_pe_1_4_4_n40), .A2(
        npu_inst_pe_1_4_4_n3), .ZN(npu_inst_pe_1_4_4_n38) );
  NOR2_X1 npu_inst_pe_1_4_4_U18 ( .A1(npu_inst_pe_1_4_4_n44), .A2(
        npu_inst_pe_1_4_4_n3), .ZN(npu_inst_pe_1_4_4_n42) );
  BUF_X1 npu_inst_pe_1_4_4_U17 ( .A(npu_inst_n98), .Z(npu_inst_pe_1_4_4_n8) );
  INV_X1 npu_inst_pe_1_4_4_U16 ( .A(npu_inst_n124), .ZN(npu_inst_pe_1_4_4_n12)
         );
  INV_X1 npu_inst_pe_1_4_4_U15 ( .A(npu_inst_pe_1_4_4_n38), .ZN(
        npu_inst_pe_1_4_4_n114) );
  INV_X1 npu_inst_pe_1_4_4_U14 ( .A(npu_inst_pe_1_4_4_n58), .ZN(
        npu_inst_pe_1_4_4_n119) );
  INV_X1 npu_inst_pe_1_4_4_U13 ( .A(npu_inst_pe_1_4_4_n54), .ZN(
        npu_inst_pe_1_4_4_n118) );
  INV_X1 npu_inst_pe_1_4_4_U12 ( .A(npu_inst_pe_1_4_4_n50), .ZN(
        npu_inst_pe_1_4_4_n117) );
  INV_X1 npu_inst_pe_1_4_4_U11 ( .A(npu_inst_pe_1_4_4_n46), .ZN(
        npu_inst_pe_1_4_4_n116) );
  INV_X1 npu_inst_pe_1_4_4_U10 ( .A(npu_inst_pe_1_4_4_n42), .ZN(
        npu_inst_pe_1_4_4_n115) );
  BUF_X1 npu_inst_pe_1_4_4_U9 ( .A(npu_inst_n20), .Z(npu_inst_pe_1_4_4_n2) );
  BUF_X1 npu_inst_pe_1_4_4_U8 ( .A(npu_inst_n20), .Z(npu_inst_pe_1_4_4_n1) );
  BUF_X1 npu_inst_pe_1_4_4_U7 ( .A(npu_inst_pe_1_4_4_n12), .Z(
        npu_inst_pe_1_4_4_n11) );
  BUF_X1 npu_inst_pe_1_4_4_U6 ( .A(npu_inst_pe_1_4_4_n12), .Z(
        npu_inst_pe_1_4_4_n10) );
  BUF_X1 npu_inst_pe_1_4_4_U5 ( .A(npu_inst_pe_1_4_4_n12), .Z(
        npu_inst_pe_1_4_4_n9) );
  NOR2_X1 npu_inst_pe_1_4_4_U4 ( .A1(npu_inst_pe_1_4_4_int_q_weight_0_), .A2(
        npu_inst_pe_1_4_4_n1), .ZN(npu_inst_pe_1_4_4_n76) );
  NOR2_X1 npu_inst_pe_1_4_4_U3 ( .A1(npu_inst_pe_1_4_4_n27), .A2(
        npu_inst_pe_1_4_4_n1), .ZN(npu_inst_pe_1_4_4_n77) );
  FA_X1 npu_inst_pe_1_4_4_sub_67_U2_1 ( .A(npu_inst_pe_1_4_4_int_q_acc_1_), 
        .B(npu_inst_pe_1_4_4_n14), .CI(npu_inst_pe_1_4_4_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_4_4_sub_67_carry_2_), .S(npu_inst_pe_1_4_4_N66) );
  FA_X1 npu_inst_pe_1_4_4_add_69_U1_1 ( .A(npu_inst_pe_1_4_4_int_q_acc_1_), 
        .B(npu_inst_pe_1_4_4_int_data_1_), .CI(
        npu_inst_pe_1_4_4_add_69_carry_1_), .CO(
        npu_inst_pe_1_4_4_add_69_carry_2_), .S(npu_inst_pe_1_4_4_N74) );
  NAND3_X1 npu_inst_pe_1_4_4_U109 ( .A1(npu_inst_pe_1_4_4_n5), .A2(
        npu_inst_pe_1_4_4_n7), .A3(npu_inst_pe_1_4_4_n8), .ZN(
        npu_inst_pe_1_4_4_n44) );
  NAND3_X1 npu_inst_pe_1_4_4_U108 ( .A1(npu_inst_pe_1_4_4_n4), .A2(
        npu_inst_pe_1_4_4_n7), .A3(npu_inst_pe_1_4_4_n8), .ZN(
        npu_inst_pe_1_4_4_n40) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_4_4_n34), .CK(
        npu_inst_pe_1_4_4_net3734), .RN(npu_inst_pe_1_4_4_n9), .Q(
        npu_inst_pe_1_4_4_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_4_4_n35), .CK(
        npu_inst_pe_1_4_4_net3734), .RN(npu_inst_pe_1_4_4_n9), .Q(
        npu_inst_pe_1_4_4_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_4_4_n36), .CK(
        npu_inst_pe_1_4_4_net3734), .RN(npu_inst_pe_1_4_4_n9), .Q(
        npu_inst_pe_1_4_4_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_4_4_n98), .CK(
        npu_inst_pe_1_4_4_net3734), .RN(npu_inst_pe_1_4_4_n9), .Q(
        npu_inst_pe_1_4_4_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_4_4_n99), .CK(
        npu_inst_pe_1_4_4_net3734), .RN(npu_inst_pe_1_4_4_n9), .Q(
        npu_inst_pe_1_4_4_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_4_4_n100), 
        .CK(npu_inst_pe_1_4_4_net3734), .RN(npu_inst_pe_1_4_4_n9), .Q(
        npu_inst_pe_1_4_4_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_4_4_n33), .CK(
        npu_inst_pe_1_4_4_net3734), .RN(npu_inst_pe_1_4_4_n9), .Q(
        npu_inst_pe_1_4_4_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_4_4_n101), 
        .CK(npu_inst_pe_1_4_4_net3734), .RN(npu_inst_pe_1_4_4_n9), .Q(
        npu_inst_pe_1_4_4_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_weight_reg_0_ ( .D(npu_inst_n110), .CK(
        npu_inst_pe_1_4_4_net3740), .RN(npu_inst_pe_1_4_4_n9), .Q(
        npu_inst_pe_1_4_4_int_q_weight_0_), .QN(npu_inst_pe_1_4_4_n27) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_weight_reg_1_ ( .D(npu_inst_n116), .CK(
        npu_inst_pe_1_4_4_net3740), .RN(npu_inst_pe_1_4_4_n9), .Q(
        npu_inst_pe_1_4_4_int_q_weight_1_), .QN(npu_inst_pe_1_4_4_n26) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_4_4_n113), 
        .CK(npu_inst_pe_1_4_4_net3740), .RN(npu_inst_pe_1_4_4_n9), .Q(
        npu_inst_pe_1_4_4_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_4_4_n107), 
        .CK(npu_inst_pe_1_4_4_net3740), .RN(npu_inst_pe_1_4_4_n9), .Q(
        npu_inst_pe_1_4_4_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_4_4_n112), 
        .CK(npu_inst_pe_1_4_4_net3740), .RN(npu_inst_pe_1_4_4_n10), .Q(
        npu_inst_pe_1_4_4_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_4_4_n106), 
        .CK(npu_inst_pe_1_4_4_net3740), .RN(npu_inst_pe_1_4_4_n10), .Q(
        npu_inst_pe_1_4_4_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_4_4_n111), 
        .CK(npu_inst_pe_1_4_4_net3740), .RN(npu_inst_pe_1_4_4_n10), .Q(
        npu_inst_pe_1_4_4_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_4_4_n105), 
        .CK(npu_inst_pe_1_4_4_net3740), .RN(npu_inst_pe_1_4_4_n10), .Q(
        npu_inst_pe_1_4_4_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_4_4_n110), 
        .CK(npu_inst_pe_1_4_4_net3740), .RN(npu_inst_pe_1_4_4_n10), .Q(
        npu_inst_pe_1_4_4_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_4_4_n104), 
        .CK(npu_inst_pe_1_4_4_net3740), .RN(npu_inst_pe_1_4_4_n10), .Q(
        npu_inst_pe_1_4_4_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_4_4_n109), 
        .CK(npu_inst_pe_1_4_4_net3740), .RN(npu_inst_pe_1_4_4_n10), .Q(
        npu_inst_pe_1_4_4_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_4_4_n103), 
        .CK(npu_inst_pe_1_4_4_net3740), .RN(npu_inst_pe_1_4_4_n10), .Q(
        npu_inst_pe_1_4_4_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_4_4_n108), 
        .CK(npu_inst_pe_1_4_4_net3740), .RN(npu_inst_pe_1_4_4_n10), .Q(
        npu_inst_pe_1_4_4_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_4_4_n102), 
        .CK(npu_inst_pe_1_4_4_net3740), .RN(npu_inst_pe_1_4_4_n10), .Q(
        npu_inst_pe_1_4_4_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_4_4_n86), 
        .CK(npu_inst_pe_1_4_4_net3740), .RN(npu_inst_pe_1_4_4_n10), .Q(
        npu_inst_pe_1_4_4_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_4_4_n87), 
        .CK(npu_inst_pe_1_4_4_net3740), .RN(npu_inst_pe_1_4_4_n10), .Q(
        npu_inst_pe_1_4_4_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_4_4_n88), 
        .CK(npu_inst_pe_1_4_4_net3740), .RN(npu_inst_pe_1_4_4_n11), .Q(
        npu_inst_pe_1_4_4_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_4_4_n89), 
        .CK(npu_inst_pe_1_4_4_net3740), .RN(npu_inst_pe_1_4_4_n11), .Q(
        npu_inst_pe_1_4_4_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_4_4_n90), 
        .CK(npu_inst_pe_1_4_4_net3740), .RN(npu_inst_pe_1_4_4_n11), .Q(
        npu_inst_pe_1_4_4_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_4_4_n91), 
        .CK(npu_inst_pe_1_4_4_net3740), .RN(npu_inst_pe_1_4_4_n11), .Q(
        npu_inst_pe_1_4_4_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_4_4_n92), 
        .CK(npu_inst_pe_1_4_4_net3740), .RN(npu_inst_pe_1_4_4_n11), .Q(
        npu_inst_pe_1_4_4_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_4_4_n93), 
        .CK(npu_inst_pe_1_4_4_net3740), .RN(npu_inst_pe_1_4_4_n11), .Q(
        npu_inst_pe_1_4_4_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_4_4_n94), 
        .CK(npu_inst_pe_1_4_4_net3740), .RN(npu_inst_pe_1_4_4_n11), .Q(
        npu_inst_pe_1_4_4_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_4_4_n95), 
        .CK(npu_inst_pe_1_4_4_net3740), .RN(npu_inst_pe_1_4_4_n11), .Q(
        npu_inst_pe_1_4_4_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_4_4_n96), 
        .CK(npu_inst_pe_1_4_4_net3740), .RN(npu_inst_pe_1_4_4_n11), .Q(
        npu_inst_pe_1_4_4_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_4_4_n97), 
        .CK(npu_inst_pe_1_4_4_net3740), .RN(npu_inst_pe_1_4_4_n11), .Q(
        npu_inst_pe_1_4_4_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_4_4_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_4_4_N84), .SE(1'b0), .GCK(npu_inst_pe_1_4_4_net3734) );
  CLKGATETST_X1 npu_inst_pe_1_4_4_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n63), .SE(1'b0), .GCK(npu_inst_pe_1_4_4_net3740) );
  MUX2_X1 npu_inst_pe_1_4_5_U162 ( .A(npu_inst_pe_1_4_5_n32), .B(
        npu_inst_pe_1_4_5_n29), .S(npu_inst_pe_1_4_5_n8), .Z(
        npu_inst_pe_1_4_5_N93) );
  MUX2_X1 npu_inst_pe_1_4_5_U161 ( .A(npu_inst_pe_1_4_5_n31), .B(
        npu_inst_pe_1_4_5_n30), .S(npu_inst_pe_1_4_5_n6), .Z(
        npu_inst_pe_1_4_5_n32) );
  MUX2_X1 npu_inst_pe_1_4_5_U160 ( .A(npu_inst_pe_1_4_5_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_4_5_int_q_reg_v_1__0_), .S(npu_inst_pe_1_4_5_n4), .Z(
        npu_inst_pe_1_4_5_n31) );
  MUX2_X1 npu_inst_pe_1_4_5_U159 ( .A(npu_inst_pe_1_4_5_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_4_5_int_q_reg_v_3__0_), .S(npu_inst_pe_1_4_5_n4), .Z(
        npu_inst_pe_1_4_5_n30) );
  MUX2_X1 npu_inst_pe_1_4_5_U158 ( .A(npu_inst_pe_1_4_5_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_4_5_int_q_reg_v_5__0_), .S(npu_inst_pe_1_4_5_n4), .Z(
        npu_inst_pe_1_4_5_n29) );
  MUX2_X1 npu_inst_pe_1_4_5_U157 ( .A(npu_inst_pe_1_4_5_n28), .B(
        npu_inst_pe_1_4_5_n23), .S(npu_inst_pe_1_4_5_n8), .Z(
        npu_inst_pe_1_4_5_N94) );
  MUX2_X1 npu_inst_pe_1_4_5_U156 ( .A(npu_inst_pe_1_4_5_n25), .B(
        npu_inst_pe_1_4_5_n24), .S(npu_inst_pe_1_4_5_n6), .Z(
        npu_inst_pe_1_4_5_n28) );
  MUX2_X1 npu_inst_pe_1_4_5_U155 ( .A(npu_inst_pe_1_4_5_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_4_5_int_q_reg_v_1__1_), .S(npu_inst_pe_1_4_5_n4), .Z(
        npu_inst_pe_1_4_5_n25) );
  MUX2_X1 npu_inst_pe_1_4_5_U154 ( .A(npu_inst_pe_1_4_5_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_4_5_int_q_reg_v_3__1_), .S(npu_inst_pe_1_4_5_n4), .Z(
        npu_inst_pe_1_4_5_n24) );
  MUX2_X1 npu_inst_pe_1_4_5_U153 ( .A(npu_inst_pe_1_4_5_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_4_5_int_q_reg_v_5__1_), .S(npu_inst_pe_1_4_5_n4), .Z(
        npu_inst_pe_1_4_5_n23) );
  MUX2_X1 npu_inst_pe_1_4_5_U152 ( .A(npu_inst_pe_1_4_5_n22), .B(
        npu_inst_pe_1_4_5_n19), .S(npu_inst_pe_1_4_5_n8), .Z(
        npu_inst_int_data_x_4__5__1_) );
  MUX2_X1 npu_inst_pe_1_4_5_U151 ( .A(npu_inst_pe_1_4_5_n21), .B(
        npu_inst_pe_1_4_5_n20), .S(npu_inst_pe_1_4_5_n6), .Z(
        npu_inst_pe_1_4_5_n22) );
  MUX2_X1 npu_inst_pe_1_4_5_U150 ( .A(npu_inst_pe_1_4_5_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_4_5_int_q_reg_h_1__1_), .S(npu_inst_pe_1_4_5_n4), .Z(
        npu_inst_pe_1_4_5_n21) );
  MUX2_X1 npu_inst_pe_1_4_5_U149 ( .A(npu_inst_pe_1_4_5_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_4_5_int_q_reg_h_3__1_), .S(npu_inst_pe_1_4_5_n4), .Z(
        npu_inst_pe_1_4_5_n20) );
  MUX2_X1 npu_inst_pe_1_4_5_U148 ( .A(npu_inst_pe_1_4_5_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_4_5_int_q_reg_h_5__1_), .S(npu_inst_pe_1_4_5_n4), .Z(
        npu_inst_pe_1_4_5_n19) );
  MUX2_X1 npu_inst_pe_1_4_5_U147 ( .A(npu_inst_pe_1_4_5_n18), .B(
        npu_inst_pe_1_4_5_n15), .S(npu_inst_pe_1_4_5_n8), .Z(
        npu_inst_int_data_x_4__5__0_) );
  MUX2_X1 npu_inst_pe_1_4_5_U146 ( .A(npu_inst_pe_1_4_5_n17), .B(
        npu_inst_pe_1_4_5_n16), .S(npu_inst_pe_1_4_5_n6), .Z(
        npu_inst_pe_1_4_5_n18) );
  MUX2_X1 npu_inst_pe_1_4_5_U145 ( .A(npu_inst_pe_1_4_5_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_4_5_int_q_reg_h_1__0_), .S(npu_inst_pe_1_4_5_n4), .Z(
        npu_inst_pe_1_4_5_n17) );
  MUX2_X1 npu_inst_pe_1_4_5_U144 ( .A(npu_inst_pe_1_4_5_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_4_5_int_q_reg_h_3__0_), .S(npu_inst_pe_1_4_5_n4), .Z(
        npu_inst_pe_1_4_5_n16) );
  MUX2_X1 npu_inst_pe_1_4_5_U143 ( .A(npu_inst_pe_1_4_5_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_4_5_int_q_reg_h_5__0_), .S(npu_inst_pe_1_4_5_n4), .Z(
        npu_inst_pe_1_4_5_n15) );
  XOR2_X1 npu_inst_pe_1_4_5_U142 ( .A(npu_inst_pe_1_4_5_int_data_0_), .B(
        npu_inst_pe_1_4_5_int_q_acc_0_), .Z(npu_inst_pe_1_4_5_N73) );
  AND2_X1 npu_inst_pe_1_4_5_U141 ( .A1(npu_inst_pe_1_4_5_int_q_acc_0_), .A2(
        npu_inst_pe_1_4_5_int_data_0_), .ZN(npu_inst_pe_1_4_5_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_4_5_U140 ( .A(npu_inst_pe_1_4_5_int_q_acc_0_), .B(
        npu_inst_pe_1_4_5_n13), .ZN(npu_inst_pe_1_4_5_N65) );
  OR2_X1 npu_inst_pe_1_4_5_U139 ( .A1(npu_inst_pe_1_4_5_n13), .A2(
        npu_inst_pe_1_4_5_int_q_acc_0_), .ZN(npu_inst_pe_1_4_5_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_4_5_U138 ( .A(npu_inst_pe_1_4_5_int_q_acc_2_), .B(
        npu_inst_pe_1_4_5_add_69_carry_2_), .Z(npu_inst_pe_1_4_5_N75) );
  AND2_X1 npu_inst_pe_1_4_5_U137 ( .A1(npu_inst_pe_1_4_5_add_69_carry_2_), 
        .A2(npu_inst_pe_1_4_5_int_q_acc_2_), .ZN(
        npu_inst_pe_1_4_5_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_4_5_U136 ( .A(npu_inst_pe_1_4_5_int_q_acc_3_), .B(
        npu_inst_pe_1_4_5_add_69_carry_3_), .Z(npu_inst_pe_1_4_5_N76) );
  AND2_X1 npu_inst_pe_1_4_5_U135 ( .A1(npu_inst_pe_1_4_5_add_69_carry_3_), 
        .A2(npu_inst_pe_1_4_5_int_q_acc_3_), .ZN(
        npu_inst_pe_1_4_5_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_4_5_U134 ( .A(npu_inst_pe_1_4_5_int_q_acc_4_), .B(
        npu_inst_pe_1_4_5_add_69_carry_4_), .Z(npu_inst_pe_1_4_5_N77) );
  AND2_X1 npu_inst_pe_1_4_5_U133 ( .A1(npu_inst_pe_1_4_5_add_69_carry_4_), 
        .A2(npu_inst_pe_1_4_5_int_q_acc_4_), .ZN(
        npu_inst_pe_1_4_5_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_4_5_U132 ( .A(npu_inst_pe_1_4_5_int_q_acc_5_), .B(
        npu_inst_pe_1_4_5_add_69_carry_5_), .Z(npu_inst_pe_1_4_5_N78) );
  AND2_X1 npu_inst_pe_1_4_5_U131 ( .A1(npu_inst_pe_1_4_5_add_69_carry_5_), 
        .A2(npu_inst_pe_1_4_5_int_q_acc_5_), .ZN(
        npu_inst_pe_1_4_5_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_4_5_U130 ( .A(npu_inst_pe_1_4_5_int_q_acc_6_), .B(
        npu_inst_pe_1_4_5_add_69_carry_6_), .Z(npu_inst_pe_1_4_5_N79) );
  AND2_X1 npu_inst_pe_1_4_5_U129 ( .A1(npu_inst_pe_1_4_5_add_69_carry_6_), 
        .A2(npu_inst_pe_1_4_5_int_q_acc_6_), .ZN(
        npu_inst_pe_1_4_5_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_4_5_U128 ( .A(npu_inst_pe_1_4_5_int_q_acc_7_), .B(
        npu_inst_pe_1_4_5_add_69_carry_7_), .Z(npu_inst_pe_1_4_5_N80) );
  XNOR2_X1 npu_inst_pe_1_4_5_U127 ( .A(npu_inst_pe_1_4_5_sub_67_carry_2_), .B(
        npu_inst_pe_1_4_5_int_q_acc_2_), .ZN(npu_inst_pe_1_4_5_N67) );
  OR2_X1 npu_inst_pe_1_4_5_U126 ( .A1(npu_inst_pe_1_4_5_int_q_acc_2_), .A2(
        npu_inst_pe_1_4_5_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_4_5_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_4_5_U125 ( .A(npu_inst_pe_1_4_5_sub_67_carry_3_), .B(
        npu_inst_pe_1_4_5_int_q_acc_3_), .ZN(npu_inst_pe_1_4_5_N68) );
  OR2_X1 npu_inst_pe_1_4_5_U124 ( .A1(npu_inst_pe_1_4_5_int_q_acc_3_), .A2(
        npu_inst_pe_1_4_5_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_4_5_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_4_5_U123 ( .A(npu_inst_pe_1_4_5_sub_67_carry_4_), .B(
        npu_inst_pe_1_4_5_int_q_acc_4_), .ZN(npu_inst_pe_1_4_5_N69) );
  OR2_X1 npu_inst_pe_1_4_5_U122 ( .A1(npu_inst_pe_1_4_5_int_q_acc_4_), .A2(
        npu_inst_pe_1_4_5_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_4_5_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_4_5_U121 ( .A(npu_inst_pe_1_4_5_sub_67_carry_5_), .B(
        npu_inst_pe_1_4_5_int_q_acc_5_), .ZN(npu_inst_pe_1_4_5_N70) );
  OR2_X1 npu_inst_pe_1_4_5_U120 ( .A1(npu_inst_pe_1_4_5_int_q_acc_5_), .A2(
        npu_inst_pe_1_4_5_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_4_5_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_4_5_U119 ( .A(npu_inst_pe_1_4_5_sub_67_carry_6_), .B(
        npu_inst_pe_1_4_5_int_q_acc_6_), .ZN(npu_inst_pe_1_4_5_N71) );
  OR2_X1 npu_inst_pe_1_4_5_U118 ( .A1(npu_inst_pe_1_4_5_int_q_acc_6_), .A2(
        npu_inst_pe_1_4_5_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_4_5_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_4_5_U117 ( .A(npu_inst_pe_1_4_5_int_q_acc_7_), .B(
        npu_inst_pe_1_4_5_sub_67_carry_7_), .ZN(npu_inst_pe_1_4_5_N72) );
  INV_X1 npu_inst_pe_1_4_5_U116 ( .A(npu_inst_n77), .ZN(npu_inst_pe_1_4_5_n7)
         );
  INV_X1 npu_inst_pe_1_4_5_U115 ( .A(npu_inst_pe_1_4_5_n7), .ZN(
        npu_inst_pe_1_4_5_n6) );
  INV_X1 npu_inst_pe_1_4_5_U114 ( .A(npu_inst_n55), .ZN(npu_inst_pe_1_4_5_n3)
         );
  AOI22_X1 npu_inst_pe_1_4_5_U113 ( .A1(npu_inst_int_data_y_5__5__0_), .A2(
        npu_inst_pe_1_4_5_n58), .B1(npu_inst_pe_1_4_5_n119), .B2(
        npu_inst_pe_1_4_5_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_4_5_n57) );
  INV_X1 npu_inst_pe_1_4_5_U112 ( .A(npu_inst_pe_1_4_5_n57), .ZN(
        npu_inst_pe_1_4_5_n108) );
  AOI22_X1 npu_inst_pe_1_4_5_U111 ( .A1(npu_inst_int_data_y_5__5__0_), .A2(
        npu_inst_pe_1_4_5_n54), .B1(npu_inst_pe_1_4_5_n118), .B2(
        npu_inst_pe_1_4_5_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_4_5_n53) );
  INV_X1 npu_inst_pe_1_4_5_U110 ( .A(npu_inst_pe_1_4_5_n53), .ZN(
        npu_inst_pe_1_4_5_n109) );
  AOI22_X1 npu_inst_pe_1_4_5_U107 ( .A1(npu_inst_int_data_y_5__5__0_), .A2(
        npu_inst_pe_1_4_5_n50), .B1(npu_inst_pe_1_4_5_n117), .B2(
        npu_inst_pe_1_4_5_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_4_5_n49) );
  INV_X1 npu_inst_pe_1_4_5_U106 ( .A(npu_inst_pe_1_4_5_n49), .ZN(
        npu_inst_pe_1_4_5_n110) );
  AOI22_X1 npu_inst_pe_1_4_5_U105 ( .A1(npu_inst_int_data_y_5__5__0_), .A2(
        npu_inst_pe_1_4_5_n46), .B1(npu_inst_pe_1_4_5_n116), .B2(
        npu_inst_pe_1_4_5_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_4_5_n45) );
  INV_X1 npu_inst_pe_1_4_5_U104 ( .A(npu_inst_pe_1_4_5_n45), .ZN(
        npu_inst_pe_1_4_5_n111) );
  AOI22_X1 npu_inst_pe_1_4_5_U103 ( .A1(npu_inst_int_data_y_5__5__0_), .A2(
        npu_inst_pe_1_4_5_n42), .B1(npu_inst_pe_1_4_5_n115), .B2(
        npu_inst_pe_1_4_5_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_4_5_n41) );
  INV_X1 npu_inst_pe_1_4_5_U102 ( .A(npu_inst_pe_1_4_5_n41), .ZN(
        npu_inst_pe_1_4_5_n112) );
  AOI22_X1 npu_inst_pe_1_4_5_U101 ( .A1(npu_inst_int_data_y_5__5__1_), .A2(
        npu_inst_pe_1_4_5_n58), .B1(npu_inst_pe_1_4_5_n119), .B2(
        npu_inst_pe_1_4_5_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_4_5_n59) );
  INV_X1 npu_inst_pe_1_4_5_U100 ( .A(npu_inst_pe_1_4_5_n59), .ZN(
        npu_inst_pe_1_4_5_n102) );
  AOI22_X1 npu_inst_pe_1_4_5_U99 ( .A1(npu_inst_int_data_y_5__5__1_), .A2(
        npu_inst_pe_1_4_5_n54), .B1(npu_inst_pe_1_4_5_n118), .B2(
        npu_inst_pe_1_4_5_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_4_5_n55) );
  INV_X1 npu_inst_pe_1_4_5_U98 ( .A(npu_inst_pe_1_4_5_n55), .ZN(
        npu_inst_pe_1_4_5_n103) );
  AOI22_X1 npu_inst_pe_1_4_5_U97 ( .A1(npu_inst_int_data_y_5__5__1_), .A2(
        npu_inst_pe_1_4_5_n50), .B1(npu_inst_pe_1_4_5_n117), .B2(
        npu_inst_pe_1_4_5_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_4_5_n51) );
  INV_X1 npu_inst_pe_1_4_5_U96 ( .A(npu_inst_pe_1_4_5_n51), .ZN(
        npu_inst_pe_1_4_5_n104) );
  AOI22_X1 npu_inst_pe_1_4_5_U95 ( .A1(npu_inst_int_data_y_5__5__1_), .A2(
        npu_inst_pe_1_4_5_n46), .B1(npu_inst_pe_1_4_5_n116), .B2(
        npu_inst_pe_1_4_5_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_4_5_n47) );
  INV_X1 npu_inst_pe_1_4_5_U94 ( .A(npu_inst_pe_1_4_5_n47), .ZN(
        npu_inst_pe_1_4_5_n105) );
  AOI22_X1 npu_inst_pe_1_4_5_U93 ( .A1(npu_inst_int_data_y_5__5__1_), .A2(
        npu_inst_pe_1_4_5_n42), .B1(npu_inst_pe_1_4_5_n115), .B2(
        npu_inst_pe_1_4_5_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_4_5_n43) );
  INV_X1 npu_inst_pe_1_4_5_U92 ( .A(npu_inst_pe_1_4_5_n43), .ZN(
        npu_inst_pe_1_4_5_n106) );
  AOI22_X1 npu_inst_pe_1_4_5_U91 ( .A1(npu_inst_pe_1_4_5_n38), .A2(
        npu_inst_int_data_y_5__5__1_), .B1(npu_inst_pe_1_4_5_n114), .B2(
        npu_inst_pe_1_4_5_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_4_5_n39) );
  INV_X1 npu_inst_pe_1_4_5_U90 ( .A(npu_inst_pe_1_4_5_n39), .ZN(
        npu_inst_pe_1_4_5_n107) );
  AOI22_X1 npu_inst_pe_1_4_5_U89 ( .A1(npu_inst_pe_1_4_5_n38), .A2(
        npu_inst_int_data_y_5__5__0_), .B1(npu_inst_pe_1_4_5_n114), .B2(
        npu_inst_pe_1_4_5_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_4_5_n37) );
  INV_X1 npu_inst_pe_1_4_5_U88 ( .A(npu_inst_pe_1_4_5_n37), .ZN(
        npu_inst_pe_1_4_5_n113) );
  NAND2_X1 npu_inst_pe_1_4_5_U87 ( .A1(npu_inst_pe_1_4_5_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_4_5_n60), .ZN(npu_inst_pe_1_4_5_n74) );
  OAI21_X1 npu_inst_pe_1_4_5_U86 ( .B1(npu_inst_pe_1_4_5_n63), .B2(
        npu_inst_pe_1_4_5_n60), .A(npu_inst_pe_1_4_5_n74), .ZN(
        npu_inst_pe_1_4_5_n97) );
  NAND2_X1 npu_inst_pe_1_4_5_U85 ( .A1(npu_inst_pe_1_4_5_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_4_5_n60), .ZN(npu_inst_pe_1_4_5_n73) );
  OAI21_X1 npu_inst_pe_1_4_5_U84 ( .B1(npu_inst_pe_1_4_5_n61), .B2(
        npu_inst_pe_1_4_5_n60), .A(npu_inst_pe_1_4_5_n73), .ZN(
        npu_inst_pe_1_4_5_n96) );
  NAND2_X1 npu_inst_pe_1_4_5_U83 ( .A1(npu_inst_pe_1_4_5_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_4_5_n56), .ZN(npu_inst_pe_1_4_5_n72) );
  OAI21_X1 npu_inst_pe_1_4_5_U82 ( .B1(npu_inst_pe_1_4_5_n63), .B2(
        npu_inst_pe_1_4_5_n56), .A(npu_inst_pe_1_4_5_n72), .ZN(
        npu_inst_pe_1_4_5_n95) );
  NAND2_X1 npu_inst_pe_1_4_5_U81 ( .A1(npu_inst_pe_1_4_5_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_4_5_n56), .ZN(npu_inst_pe_1_4_5_n71) );
  OAI21_X1 npu_inst_pe_1_4_5_U80 ( .B1(npu_inst_pe_1_4_5_n61), .B2(
        npu_inst_pe_1_4_5_n56), .A(npu_inst_pe_1_4_5_n71), .ZN(
        npu_inst_pe_1_4_5_n94) );
  NAND2_X1 npu_inst_pe_1_4_5_U79 ( .A1(npu_inst_pe_1_4_5_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_4_5_n52), .ZN(npu_inst_pe_1_4_5_n70) );
  OAI21_X1 npu_inst_pe_1_4_5_U78 ( .B1(npu_inst_pe_1_4_5_n63), .B2(
        npu_inst_pe_1_4_5_n52), .A(npu_inst_pe_1_4_5_n70), .ZN(
        npu_inst_pe_1_4_5_n93) );
  NAND2_X1 npu_inst_pe_1_4_5_U77 ( .A1(npu_inst_pe_1_4_5_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_4_5_n52), .ZN(npu_inst_pe_1_4_5_n69) );
  OAI21_X1 npu_inst_pe_1_4_5_U76 ( .B1(npu_inst_pe_1_4_5_n61), .B2(
        npu_inst_pe_1_4_5_n52), .A(npu_inst_pe_1_4_5_n69), .ZN(
        npu_inst_pe_1_4_5_n92) );
  NAND2_X1 npu_inst_pe_1_4_5_U75 ( .A1(npu_inst_pe_1_4_5_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_4_5_n48), .ZN(npu_inst_pe_1_4_5_n68) );
  OAI21_X1 npu_inst_pe_1_4_5_U74 ( .B1(npu_inst_pe_1_4_5_n63), .B2(
        npu_inst_pe_1_4_5_n48), .A(npu_inst_pe_1_4_5_n68), .ZN(
        npu_inst_pe_1_4_5_n91) );
  NAND2_X1 npu_inst_pe_1_4_5_U73 ( .A1(npu_inst_pe_1_4_5_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_4_5_n48), .ZN(npu_inst_pe_1_4_5_n67) );
  OAI21_X1 npu_inst_pe_1_4_5_U72 ( .B1(npu_inst_pe_1_4_5_n61), .B2(
        npu_inst_pe_1_4_5_n48), .A(npu_inst_pe_1_4_5_n67), .ZN(
        npu_inst_pe_1_4_5_n90) );
  NAND2_X1 npu_inst_pe_1_4_5_U71 ( .A1(npu_inst_pe_1_4_5_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_4_5_n44), .ZN(npu_inst_pe_1_4_5_n66) );
  OAI21_X1 npu_inst_pe_1_4_5_U70 ( .B1(npu_inst_pe_1_4_5_n63), .B2(
        npu_inst_pe_1_4_5_n44), .A(npu_inst_pe_1_4_5_n66), .ZN(
        npu_inst_pe_1_4_5_n89) );
  NAND2_X1 npu_inst_pe_1_4_5_U69 ( .A1(npu_inst_pe_1_4_5_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_4_5_n44), .ZN(npu_inst_pe_1_4_5_n65) );
  OAI21_X1 npu_inst_pe_1_4_5_U68 ( .B1(npu_inst_pe_1_4_5_n61), .B2(
        npu_inst_pe_1_4_5_n44), .A(npu_inst_pe_1_4_5_n65), .ZN(
        npu_inst_pe_1_4_5_n88) );
  NAND2_X1 npu_inst_pe_1_4_5_U67 ( .A1(npu_inst_pe_1_4_5_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_4_5_n40), .ZN(npu_inst_pe_1_4_5_n64) );
  OAI21_X1 npu_inst_pe_1_4_5_U66 ( .B1(npu_inst_pe_1_4_5_n63), .B2(
        npu_inst_pe_1_4_5_n40), .A(npu_inst_pe_1_4_5_n64), .ZN(
        npu_inst_pe_1_4_5_n87) );
  NAND2_X1 npu_inst_pe_1_4_5_U65 ( .A1(npu_inst_pe_1_4_5_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_4_5_n40), .ZN(npu_inst_pe_1_4_5_n62) );
  OAI21_X1 npu_inst_pe_1_4_5_U64 ( .B1(npu_inst_pe_1_4_5_n61), .B2(
        npu_inst_pe_1_4_5_n40), .A(npu_inst_pe_1_4_5_n62), .ZN(
        npu_inst_pe_1_4_5_n86) );
  AND2_X1 npu_inst_pe_1_4_5_U63 ( .A1(npu_inst_pe_1_4_5_N93), .A2(npu_inst_n55), .ZN(npu_inst_int_data_y_4__5__0_) );
  AND2_X1 npu_inst_pe_1_4_5_U62 ( .A1(npu_inst_n55), .A2(npu_inst_pe_1_4_5_N94), .ZN(npu_inst_int_data_y_4__5__1_) );
  NOR3_X1 npu_inst_pe_1_4_5_U61 ( .A1(npu_inst_pe_1_4_5_n26), .A2(npu_inst_n55), .A3(npu_inst_int_ckg[26]), .ZN(npu_inst_pe_1_4_5_n85) );
  OR2_X1 npu_inst_pe_1_4_5_U60 ( .A1(npu_inst_pe_1_4_5_n85), .A2(
        npu_inst_pe_1_4_5_n2), .ZN(npu_inst_pe_1_4_5_N84) );
  AND2_X1 npu_inst_pe_1_4_5_U59 ( .A1(npu_inst_pe_1_4_5_int_q_acc_0_), .A2(
        npu_inst_pe_1_4_5_n1), .ZN(npu_inst_int_data_res_4__5__0_) );
  AND2_X1 npu_inst_pe_1_4_5_U58 ( .A1(npu_inst_pe_1_4_5_n2), .A2(
        npu_inst_pe_1_4_5_int_q_acc_7_), .ZN(npu_inst_int_data_res_4__5__7_)
         );
  AND2_X1 npu_inst_pe_1_4_5_U57 ( .A1(npu_inst_pe_1_4_5_int_q_acc_1_), .A2(
        npu_inst_pe_1_4_5_n1), .ZN(npu_inst_int_data_res_4__5__1_) );
  AND2_X1 npu_inst_pe_1_4_5_U56 ( .A1(npu_inst_pe_1_4_5_int_q_acc_2_), .A2(
        npu_inst_pe_1_4_5_n1), .ZN(npu_inst_int_data_res_4__5__2_) );
  AND2_X1 npu_inst_pe_1_4_5_U55 ( .A1(npu_inst_pe_1_4_5_int_q_acc_3_), .A2(
        npu_inst_pe_1_4_5_n2), .ZN(npu_inst_int_data_res_4__5__3_) );
  AND2_X1 npu_inst_pe_1_4_5_U54 ( .A1(npu_inst_pe_1_4_5_int_q_acc_4_), .A2(
        npu_inst_pe_1_4_5_n2), .ZN(npu_inst_int_data_res_4__5__4_) );
  AND2_X1 npu_inst_pe_1_4_5_U53 ( .A1(npu_inst_pe_1_4_5_int_q_acc_5_), .A2(
        npu_inst_pe_1_4_5_n2), .ZN(npu_inst_int_data_res_4__5__5_) );
  AND2_X1 npu_inst_pe_1_4_5_U52 ( .A1(npu_inst_pe_1_4_5_int_q_acc_6_), .A2(
        npu_inst_pe_1_4_5_n2), .ZN(npu_inst_int_data_res_4__5__6_) );
  AOI222_X1 npu_inst_pe_1_4_5_U51 ( .A1(npu_inst_int_data_res_5__5__0_), .A2(
        npu_inst_pe_1_4_5_n1), .B1(npu_inst_pe_1_4_5_N73), .B2(
        npu_inst_pe_1_4_5_n76), .C1(npu_inst_pe_1_4_5_N65), .C2(
        npu_inst_pe_1_4_5_n77), .ZN(npu_inst_pe_1_4_5_n84) );
  INV_X1 npu_inst_pe_1_4_5_U50 ( .A(npu_inst_pe_1_4_5_n84), .ZN(
        npu_inst_pe_1_4_5_n101) );
  AOI222_X1 npu_inst_pe_1_4_5_U49 ( .A1(npu_inst_int_data_res_5__5__7_), .A2(
        npu_inst_pe_1_4_5_n1), .B1(npu_inst_pe_1_4_5_N80), .B2(
        npu_inst_pe_1_4_5_n76), .C1(npu_inst_pe_1_4_5_N72), .C2(
        npu_inst_pe_1_4_5_n77), .ZN(npu_inst_pe_1_4_5_n75) );
  INV_X1 npu_inst_pe_1_4_5_U48 ( .A(npu_inst_pe_1_4_5_n75), .ZN(
        npu_inst_pe_1_4_5_n33) );
  AOI222_X1 npu_inst_pe_1_4_5_U47 ( .A1(npu_inst_int_data_res_5__5__1_), .A2(
        npu_inst_pe_1_4_5_n1), .B1(npu_inst_pe_1_4_5_N74), .B2(
        npu_inst_pe_1_4_5_n76), .C1(npu_inst_pe_1_4_5_N66), .C2(
        npu_inst_pe_1_4_5_n77), .ZN(npu_inst_pe_1_4_5_n83) );
  INV_X1 npu_inst_pe_1_4_5_U46 ( .A(npu_inst_pe_1_4_5_n83), .ZN(
        npu_inst_pe_1_4_5_n100) );
  AOI222_X1 npu_inst_pe_1_4_5_U45 ( .A1(npu_inst_int_data_res_5__5__2_), .A2(
        npu_inst_pe_1_4_5_n1), .B1(npu_inst_pe_1_4_5_N75), .B2(
        npu_inst_pe_1_4_5_n76), .C1(npu_inst_pe_1_4_5_N67), .C2(
        npu_inst_pe_1_4_5_n77), .ZN(npu_inst_pe_1_4_5_n82) );
  INV_X1 npu_inst_pe_1_4_5_U44 ( .A(npu_inst_pe_1_4_5_n82), .ZN(
        npu_inst_pe_1_4_5_n99) );
  AOI222_X1 npu_inst_pe_1_4_5_U43 ( .A1(npu_inst_int_data_res_5__5__3_), .A2(
        npu_inst_pe_1_4_5_n1), .B1(npu_inst_pe_1_4_5_N76), .B2(
        npu_inst_pe_1_4_5_n76), .C1(npu_inst_pe_1_4_5_N68), .C2(
        npu_inst_pe_1_4_5_n77), .ZN(npu_inst_pe_1_4_5_n81) );
  INV_X1 npu_inst_pe_1_4_5_U42 ( .A(npu_inst_pe_1_4_5_n81), .ZN(
        npu_inst_pe_1_4_5_n98) );
  AOI222_X1 npu_inst_pe_1_4_5_U41 ( .A1(npu_inst_int_data_res_5__5__4_), .A2(
        npu_inst_pe_1_4_5_n1), .B1(npu_inst_pe_1_4_5_N77), .B2(
        npu_inst_pe_1_4_5_n76), .C1(npu_inst_pe_1_4_5_N69), .C2(
        npu_inst_pe_1_4_5_n77), .ZN(npu_inst_pe_1_4_5_n80) );
  INV_X1 npu_inst_pe_1_4_5_U40 ( .A(npu_inst_pe_1_4_5_n80), .ZN(
        npu_inst_pe_1_4_5_n36) );
  AOI222_X1 npu_inst_pe_1_4_5_U39 ( .A1(npu_inst_int_data_res_5__5__5_), .A2(
        npu_inst_pe_1_4_5_n1), .B1(npu_inst_pe_1_4_5_N78), .B2(
        npu_inst_pe_1_4_5_n76), .C1(npu_inst_pe_1_4_5_N70), .C2(
        npu_inst_pe_1_4_5_n77), .ZN(npu_inst_pe_1_4_5_n79) );
  INV_X1 npu_inst_pe_1_4_5_U38 ( .A(npu_inst_pe_1_4_5_n79), .ZN(
        npu_inst_pe_1_4_5_n35) );
  AOI222_X1 npu_inst_pe_1_4_5_U37 ( .A1(npu_inst_int_data_res_5__5__6_), .A2(
        npu_inst_pe_1_4_5_n1), .B1(npu_inst_pe_1_4_5_N79), .B2(
        npu_inst_pe_1_4_5_n76), .C1(npu_inst_pe_1_4_5_N71), .C2(
        npu_inst_pe_1_4_5_n77), .ZN(npu_inst_pe_1_4_5_n78) );
  INV_X1 npu_inst_pe_1_4_5_U36 ( .A(npu_inst_pe_1_4_5_n78), .ZN(
        npu_inst_pe_1_4_5_n34) );
  INV_X1 npu_inst_pe_1_4_5_U35 ( .A(npu_inst_pe_1_4_5_int_data_1_), .ZN(
        npu_inst_pe_1_4_5_n14) );
  AND2_X1 npu_inst_pe_1_4_5_U34 ( .A1(npu_inst_int_data_x_4__5__1_), .A2(
        npu_inst_pe_1_4_5_int_q_weight_1_), .ZN(npu_inst_pe_1_4_5_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_4_5_U33 ( .A1(npu_inst_int_data_x_4__5__0_), .A2(
        npu_inst_pe_1_4_5_int_q_weight_1_), .ZN(npu_inst_pe_1_4_5_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_4_5_U32 ( .A1(npu_inst_n55), .A2(
        npu_inst_int_data_y_5__5__1_), .B1(npu_inst_pe_1_4_5_n3), .B2(
        npu_inst_int_data_x_4__6__1_), .ZN(npu_inst_pe_1_4_5_n63) );
  AOI22_X1 npu_inst_pe_1_4_5_U31 ( .A1(npu_inst_n55), .A2(
        npu_inst_int_data_y_5__5__0_), .B1(npu_inst_pe_1_4_5_n3), .B2(
        npu_inst_int_data_x_4__6__0_), .ZN(npu_inst_pe_1_4_5_n61) );
  INV_X1 npu_inst_pe_1_4_5_U30 ( .A(npu_inst_pe_1_4_5_int_data_0_), .ZN(
        npu_inst_pe_1_4_5_n13) );
  INV_X1 npu_inst_pe_1_4_5_U29 ( .A(npu_inst_n69), .ZN(npu_inst_pe_1_4_5_n5)
         );
  OR3_X1 npu_inst_pe_1_4_5_U28 ( .A1(npu_inst_pe_1_4_5_n6), .A2(
        npu_inst_pe_1_4_5_n8), .A3(npu_inst_pe_1_4_5_n5), .ZN(
        npu_inst_pe_1_4_5_n56) );
  OR3_X1 npu_inst_pe_1_4_5_U27 ( .A1(npu_inst_pe_1_4_5_n5), .A2(
        npu_inst_pe_1_4_5_n8), .A3(npu_inst_pe_1_4_5_n7), .ZN(
        npu_inst_pe_1_4_5_n48) );
  INV_X1 npu_inst_pe_1_4_5_U26 ( .A(npu_inst_pe_1_4_5_n5), .ZN(
        npu_inst_pe_1_4_5_n4) );
  OR3_X1 npu_inst_pe_1_4_5_U25 ( .A1(npu_inst_pe_1_4_5_n4), .A2(
        npu_inst_pe_1_4_5_n8), .A3(npu_inst_pe_1_4_5_n7), .ZN(
        npu_inst_pe_1_4_5_n52) );
  OR3_X1 npu_inst_pe_1_4_5_U24 ( .A1(npu_inst_pe_1_4_5_n6), .A2(
        npu_inst_pe_1_4_5_n8), .A3(npu_inst_pe_1_4_5_n4), .ZN(
        npu_inst_pe_1_4_5_n60) );
  NOR2_X1 npu_inst_pe_1_4_5_U23 ( .A1(npu_inst_pe_1_4_5_n60), .A2(
        npu_inst_pe_1_4_5_n3), .ZN(npu_inst_pe_1_4_5_n58) );
  NOR2_X1 npu_inst_pe_1_4_5_U22 ( .A1(npu_inst_pe_1_4_5_n56), .A2(
        npu_inst_pe_1_4_5_n3), .ZN(npu_inst_pe_1_4_5_n54) );
  NOR2_X1 npu_inst_pe_1_4_5_U21 ( .A1(npu_inst_pe_1_4_5_n52), .A2(
        npu_inst_pe_1_4_5_n3), .ZN(npu_inst_pe_1_4_5_n50) );
  NOR2_X1 npu_inst_pe_1_4_5_U20 ( .A1(npu_inst_pe_1_4_5_n48), .A2(
        npu_inst_pe_1_4_5_n3), .ZN(npu_inst_pe_1_4_5_n46) );
  NOR2_X1 npu_inst_pe_1_4_5_U19 ( .A1(npu_inst_pe_1_4_5_n40), .A2(
        npu_inst_pe_1_4_5_n3), .ZN(npu_inst_pe_1_4_5_n38) );
  NOR2_X1 npu_inst_pe_1_4_5_U18 ( .A1(npu_inst_pe_1_4_5_n44), .A2(
        npu_inst_pe_1_4_5_n3), .ZN(npu_inst_pe_1_4_5_n42) );
  BUF_X1 npu_inst_pe_1_4_5_U17 ( .A(npu_inst_n98), .Z(npu_inst_pe_1_4_5_n8) );
  INV_X1 npu_inst_pe_1_4_5_U16 ( .A(npu_inst_n124), .ZN(npu_inst_pe_1_4_5_n12)
         );
  INV_X1 npu_inst_pe_1_4_5_U15 ( .A(npu_inst_pe_1_4_5_n38), .ZN(
        npu_inst_pe_1_4_5_n114) );
  INV_X1 npu_inst_pe_1_4_5_U14 ( .A(npu_inst_pe_1_4_5_n58), .ZN(
        npu_inst_pe_1_4_5_n119) );
  INV_X1 npu_inst_pe_1_4_5_U13 ( .A(npu_inst_pe_1_4_5_n54), .ZN(
        npu_inst_pe_1_4_5_n118) );
  INV_X1 npu_inst_pe_1_4_5_U12 ( .A(npu_inst_pe_1_4_5_n50), .ZN(
        npu_inst_pe_1_4_5_n117) );
  INV_X1 npu_inst_pe_1_4_5_U11 ( .A(npu_inst_pe_1_4_5_n46), .ZN(
        npu_inst_pe_1_4_5_n116) );
  INV_X1 npu_inst_pe_1_4_5_U10 ( .A(npu_inst_pe_1_4_5_n42), .ZN(
        npu_inst_pe_1_4_5_n115) );
  BUF_X1 npu_inst_pe_1_4_5_U9 ( .A(npu_inst_n20), .Z(npu_inst_pe_1_4_5_n2) );
  BUF_X1 npu_inst_pe_1_4_5_U8 ( .A(npu_inst_n20), .Z(npu_inst_pe_1_4_5_n1) );
  BUF_X1 npu_inst_pe_1_4_5_U7 ( .A(npu_inst_pe_1_4_5_n12), .Z(
        npu_inst_pe_1_4_5_n11) );
  BUF_X1 npu_inst_pe_1_4_5_U6 ( .A(npu_inst_pe_1_4_5_n12), .Z(
        npu_inst_pe_1_4_5_n10) );
  BUF_X1 npu_inst_pe_1_4_5_U5 ( .A(npu_inst_pe_1_4_5_n12), .Z(
        npu_inst_pe_1_4_5_n9) );
  NOR2_X1 npu_inst_pe_1_4_5_U4 ( .A1(npu_inst_pe_1_4_5_int_q_weight_0_), .A2(
        npu_inst_pe_1_4_5_n1), .ZN(npu_inst_pe_1_4_5_n76) );
  NOR2_X1 npu_inst_pe_1_4_5_U3 ( .A1(npu_inst_pe_1_4_5_n27), .A2(
        npu_inst_pe_1_4_5_n1), .ZN(npu_inst_pe_1_4_5_n77) );
  FA_X1 npu_inst_pe_1_4_5_sub_67_U2_1 ( .A(npu_inst_pe_1_4_5_int_q_acc_1_), 
        .B(npu_inst_pe_1_4_5_n14), .CI(npu_inst_pe_1_4_5_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_4_5_sub_67_carry_2_), .S(npu_inst_pe_1_4_5_N66) );
  FA_X1 npu_inst_pe_1_4_5_add_69_U1_1 ( .A(npu_inst_pe_1_4_5_int_q_acc_1_), 
        .B(npu_inst_pe_1_4_5_int_data_1_), .CI(
        npu_inst_pe_1_4_5_add_69_carry_1_), .CO(
        npu_inst_pe_1_4_5_add_69_carry_2_), .S(npu_inst_pe_1_4_5_N74) );
  NAND3_X1 npu_inst_pe_1_4_5_U109 ( .A1(npu_inst_pe_1_4_5_n5), .A2(
        npu_inst_pe_1_4_5_n7), .A3(npu_inst_pe_1_4_5_n8), .ZN(
        npu_inst_pe_1_4_5_n44) );
  NAND3_X1 npu_inst_pe_1_4_5_U108 ( .A1(npu_inst_pe_1_4_5_n4), .A2(
        npu_inst_pe_1_4_5_n7), .A3(npu_inst_pe_1_4_5_n8), .ZN(
        npu_inst_pe_1_4_5_n40) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_4_5_n34), .CK(
        npu_inst_pe_1_4_5_net3711), .RN(npu_inst_pe_1_4_5_n9), .Q(
        npu_inst_pe_1_4_5_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_4_5_n35), .CK(
        npu_inst_pe_1_4_5_net3711), .RN(npu_inst_pe_1_4_5_n9), .Q(
        npu_inst_pe_1_4_5_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_4_5_n36), .CK(
        npu_inst_pe_1_4_5_net3711), .RN(npu_inst_pe_1_4_5_n9), .Q(
        npu_inst_pe_1_4_5_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_4_5_n98), .CK(
        npu_inst_pe_1_4_5_net3711), .RN(npu_inst_pe_1_4_5_n9), .Q(
        npu_inst_pe_1_4_5_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_4_5_n99), .CK(
        npu_inst_pe_1_4_5_net3711), .RN(npu_inst_pe_1_4_5_n9), .Q(
        npu_inst_pe_1_4_5_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_4_5_n100), 
        .CK(npu_inst_pe_1_4_5_net3711), .RN(npu_inst_pe_1_4_5_n9), .Q(
        npu_inst_pe_1_4_5_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_4_5_n33), .CK(
        npu_inst_pe_1_4_5_net3711), .RN(npu_inst_pe_1_4_5_n9), .Q(
        npu_inst_pe_1_4_5_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_4_5_n101), 
        .CK(npu_inst_pe_1_4_5_net3711), .RN(npu_inst_pe_1_4_5_n9), .Q(
        npu_inst_pe_1_4_5_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_weight_reg_0_ ( .D(npu_inst_n110), .CK(
        npu_inst_pe_1_4_5_net3717), .RN(npu_inst_pe_1_4_5_n9), .Q(
        npu_inst_pe_1_4_5_int_q_weight_0_), .QN(npu_inst_pe_1_4_5_n27) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_weight_reg_1_ ( .D(npu_inst_n116), .CK(
        npu_inst_pe_1_4_5_net3717), .RN(npu_inst_pe_1_4_5_n9), .Q(
        npu_inst_pe_1_4_5_int_q_weight_1_), .QN(npu_inst_pe_1_4_5_n26) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_4_5_n113), 
        .CK(npu_inst_pe_1_4_5_net3717), .RN(npu_inst_pe_1_4_5_n9), .Q(
        npu_inst_pe_1_4_5_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_4_5_n107), 
        .CK(npu_inst_pe_1_4_5_net3717), .RN(npu_inst_pe_1_4_5_n9), .Q(
        npu_inst_pe_1_4_5_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_4_5_n112), 
        .CK(npu_inst_pe_1_4_5_net3717), .RN(npu_inst_pe_1_4_5_n10), .Q(
        npu_inst_pe_1_4_5_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_4_5_n106), 
        .CK(npu_inst_pe_1_4_5_net3717), .RN(npu_inst_pe_1_4_5_n10), .Q(
        npu_inst_pe_1_4_5_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_4_5_n111), 
        .CK(npu_inst_pe_1_4_5_net3717), .RN(npu_inst_pe_1_4_5_n10), .Q(
        npu_inst_pe_1_4_5_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_4_5_n105), 
        .CK(npu_inst_pe_1_4_5_net3717), .RN(npu_inst_pe_1_4_5_n10), .Q(
        npu_inst_pe_1_4_5_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_4_5_n110), 
        .CK(npu_inst_pe_1_4_5_net3717), .RN(npu_inst_pe_1_4_5_n10), .Q(
        npu_inst_pe_1_4_5_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_4_5_n104), 
        .CK(npu_inst_pe_1_4_5_net3717), .RN(npu_inst_pe_1_4_5_n10), .Q(
        npu_inst_pe_1_4_5_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_4_5_n109), 
        .CK(npu_inst_pe_1_4_5_net3717), .RN(npu_inst_pe_1_4_5_n10), .Q(
        npu_inst_pe_1_4_5_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_4_5_n103), 
        .CK(npu_inst_pe_1_4_5_net3717), .RN(npu_inst_pe_1_4_5_n10), .Q(
        npu_inst_pe_1_4_5_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_4_5_n108), 
        .CK(npu_inst_pe_1_4_5_net3717), .RN(npu_inst_pe_1_4_5_n10), .Q(
        npu_inst_pe_1_4_5_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_4_5_n102), 
        .CK(npu_inst_pe_1_4_5_net3717), .RN(npu_inst_pe_1_4_5_n10), .Q(
        npu_inst_pe_1_4_5_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_4_5_n86), 
        .CK(npu_inst_pe_1_4_5_net3717), .RN(npu_inst_pe_1_4_5_n10), .Q(
        npu_inst_pe_1_4_5_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_4_5_n87), 
        .CK(npu_inst_pe_1_4_5_net3717), .RN(npu_inst_pe_1_4_5_n10), .Q(
        npu_inst_pe_1_4_5_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_4_5_n88), 
        .CK(npu_inst_pe_1_4_5_net3717), .RN(npu_inst_pe_1_4_5_n11), .Q(
        npu_inst_pe_1_4_5_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_4_5_n89), 
        .CK(npu_inst_pe_1_4_5_net3717), .RN(npu_inst_pe_1_4_5_n11), .Q(
        npu_inst_pe_1_4_5_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_4_5_n90), 
        .CK(npu_inst_pe_1_4_5_net3717), .RN(npu_inst_pe_1_4_5_n11), .Q(
        npu_inst_pe_1_4_5_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_4_5_n91), 
        .CK(npu_inst_pe_1_4_5_net3717), .RN(npu_inst_pe_1_4_5_n11), .Q(
        npu_inst_pe_1_4_5_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_4_5_n92), 
        .CK(npu_inst_pe_1_4_5_net3717), .RN(npu_inst_pe_1_4_5_n11), .Q(
        npu_inst_pe_1_4_5_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_4_5_n93), 
        .CK(npu_inst_pe_1_4_5_net3717), .RN(npu_inst_pe_1_4_5_n11), .Q(
        npu_inst_pe_1_4_5_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_4_5_n94), 
        .CK(npu_inst_pe_1_4_5_net3717), .RN(npu_inst_pe_1_4_5_n11), .Q(
        npu_inst_pe_1_4_5_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_4_5_n95), 
        .CK(npu_inst_pe_1_4_5_net3717), .RN(npu_inst_pe_1_4_5_n11), .Q(
        npu_inst_pe_1_4_5_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_4_5_n96), 
        .CK(npu_inst_pe_1_4_5_net3717), .RN(npu_inst_pe_1_4_5_n11), .Q(
        npu_inst_pe_1_4_5_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_4_5_n97), 
        .CK(npu_inst_pe_1_4_5_net3717), .RN(npu_inst_pe_1_4_5_n11), .Q(
        npu_inst_pe_1_4_5_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_4_5_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_4_5_N84), .SE(1'b0), .GCK(npu_inst_pe_1_4_5_net3711) );
  CLKGATETST_X1 npu_inst_pe_1_4_5_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n63), .SE(1'b0), .GCK(npu_inst_pe_1_4_5_net3717) );
  MUX2_X1 npu_inst_pe_1_4_6_U162 ( .A(npu_inst_pe_1_4_6_n32), .B(
        npu_inst_pe_1_4_6_n29), .S(npu_inst_pe_1_4_6_n8), .Z(
        npu_inst_pe_1_4_6_N93) );
  MUX2_X1 npu_inst_pe_1_4_6_U161 ( .A(npu_inst_pe_1_4_6_n31), .B(
        npu_inst_pe_1_4_6_n30), .S(npu_inst_pe_1_4_6_n6), .Z(
        npu_inst_pe_1_4_6_n32) );
  MUX2_X1 npu_inst_pe_1_4_6_U160 ( .A(npu_inst_pe_1_4_6_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_4_6_int_q_reg_v_1__0_), .S(npu_inst_pe_1_4_6_n4), .Z(
        npu_inst_pe_1_4_6_n31) );
  MUX2_X1 npu_inst_pe_1_4_6_U159 ( .A(npu_inst_pe_1_4_6_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_4_6_int_q_reg_v_3__0_), .S(npu_inst_pe_1_4_6_n4), .Z(
        npu_inst_pe_1_4_6_n30) );
  MUX2_X1 npu_inst_pe_1_4_6_U158 ( .A(npu_inst_pe_1_4_6_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_4_6_int_q_reg_v_5__0_), .S(npu_inst_pe_1_4_6_n4), .Z(
        npu_inst_pe_1_4_6_n29) );
  MUX2_X1 npu_inst_pe_1_4_6_U157 ( .A(npu_inst_pe_1_4_6_n28), .B(
        npu_inst_pe_1_4_6_n23), .S(npu_inst_pe_1_4_6_n8), .Z(
        npu_inst_pe_1_4_6_N94) );
  MUX2_X1 npu_inst_pe_1_4_6_U156 ( .A(npu_inst_pe_1_4_6_n25), .B(
        npu_inst_pe_1_4_6_n24), .S(npu_inst_pe_1_4_6_n6), .Z(
        npu_inst_pe_1_4_6_n28) );
  MUX2_X1 npu_inst_pe_1_4_6_U155 ( .A(npu_inst_pe_1_4_6_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_4_6_int_q_reg_v_1__1_), .S(npu_inst_pe_1_4_6_n4), .Z(
        npu_inst_pe_1_4_6_n25) );
  MUX2_X1 npu_inst_pe_1_4_6_U154 ( .A(npu_inst_pe_1_4_6_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_4_6_int_q_reg_v_3__1_), .S(npu_inst_pe_1_4_6_n4), .Z(
        npu_inst_pe_1_4_6_n24) );
  MUX2_X1 npu_inst_pe_1_4_6_U153 ( .A(npu_inst_pe_1_4_6_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_4_6_int_q_reg_v_5__1_), .S(npu_inst_pe_1_4_6_n4), .Z(
        npu_inst_pe_1_4_6_n23) );
  MUX2_X1 npu_inst_pe_1_4_6_U152 ( .A(npu_inst_pe_1_4_6_n22), .B(
        npu_inst_pe_1_4_6_n19), .S(npu_inst_pe_1_4_6_n8), .Z(
        npu_inst_int_data_x_4__6__1_) );
  MUX2_X1 npu_inst_pe_1_4_6_U151 ( .A(npu_inst_pe_1_4_6_n21), .B(
        npu_inst_pe_1_4_6_n20), .S(npu_inst_pe_1_4_6_n6), .Z(
        npu_inst_pe_1_4_6_n22) );
  MUX2_X1 npu_inst_pe_1_4_6_U150 ( .A(npu_inst_pe_1_4_6_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_4_6_int_q_reg_h_1__1_), .S(npu_inst_pe_1_4_6_n4), .Z(
        npu_inst_pe_1_4_6_n21) );
  MUX2_X1 npu_inst_pe_1_4_6_U149 ( .A(npu_inst_pe_1_4_6_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_4_6_int_q_reg_h_3__1_), .S(npu_inst_pe_1_4_6_n4), .Z(
        npu_inst_pe_1_4_6_n20) );
  MUX2_X1 npu_inst_pe_1_4_6_U148 ( .A(npu_inst_pe_1_4_6_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_4_6_int_q_reg_h_5__1_), .S(npu_inst_pe_1_4_6_n4), .Z(
        npu_inst_pe_1_4_6_n19) );
  MUX2_X1 npu_inst_pe_1_4_6_U147 ( .A(npu_inst_pe_1_4_6_n18), .B(
        npu_inst_pe_1_4_6_n15), .S(npu_inst_pe_1_4_6_n8), .Z(
        npu_inst_int_data_x_4__6__0_) );
  MUX2_X1 npu_inst_pe_1_4_6_U146 ( .A(npu_inst_pe_1_4_6_n17), .B(
        npu_inst_pe_1_4_6_n16), .S(npu_inst_pe_1_4_6_n6), .Z(
        npu_inst_pe_1_4_6_n18) );
  MUX2_X1 npu_inst_pe_1_4_6_U145 ( .A(npu_inst_pe_1_4_6_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_4_6_int_q_reg_h_1__0_), .S(npu_inst_pe_1_4_6_n4), .Z(
        npu_inst_pe_1_4_6_n17) );
  MUX2_X1 npu_inst_pe_1_4_6_U144 ( .A(npu_inst_pe_1_4_6_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_4_6_int_q_reg_h_3__0_), .S(npu_inst_pe_1_4_6_n4), .Z(
        npu_inst_pe_1_4_6_n16) );
  MUX2_X1 npu_inst_pe_1_4_6_U143 ( .A(npu_inst_pe_1_4_6_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_4_6_int_q_reg_h_5__0_), .S(npu_inst_pe_1_4_6_n4), .Z(
        npu_inst_pe_1_4_6_n15) );
  XOR2_X1 npu_inst_pe_1_4_6_U142 ( .A(npu_inst_pe_1_4_6_int_data_0_), .B(
        npu_inst_pe_1_4_6_int_q_acc_0_), .Z(npu_inst_pe_1_4_6_N73) );
  AND2_X1 npu_inst_pe_1_4_6_U141 ( .A1(npu_inst_pe_1_4_6_int_q_acc_0_), .A2(
        npu_inst_pe_1_4_6_int_data_0_), .ZN(npu_inst_pe_1_4_6_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_4_6_U140 ( .A(npu_inst_pe_1_4_6_int_q_acc_0_), .B(
        npu_inst_pe_1_4_6_n13), .ZN(npu_inst_pe_1_4_6_N65) );
  OR2_X1 npu_inst_pe_1_4_6_U139 ( .A1(npu_inst_pe_1_4_6_n13), .A2(
        npu_inst_pe_1_4_6_int_q_acc_0_), .ZN(npu_inst_pe_1_4_6_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_4_6_U138 ( .A(npu_inst_pe_1_4_6_int_q_acc_2_), .B(
        npu_inst_pe_1_4_6_add_69_carry_2_), .Z(npu_inst_pe_1_4_6_N75) );
  AND2_X1 npu_inst_pe_1_4_6_U137 ( .A1(npu_inst_pe_1_4_6_add_69_carry_2_), 
        .A2(npu_inst_pe_1_4_6_int_q_acc_2_), .ZN(
        npu_inst_pe_1_4_6_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_4_6_U136 ( .A(npu_inst_pe_1_4_6_int_q_acc_3_), .B(
        npu_inst_pe_1_4_6_add_69_carry_3_), .Z(npu_inst_pe_1_4_6_N76) );
  AND2_X1 npu_inst_pe_1_4_6_U135 ( .A1(npu_inst_pe_1_4_6_add_69_carry_3_), 
        .A2(npu_inst_pe_1_4_6_int_q_acc_3_), .ZN(
        npu_inst_pe_1_4_6_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_4_6_U134 ( .A(npu_inst_pe_1_4_6_int_q_acc_4_), .B(
        npu_inst_pe_1_4_6_add_69_carry_4_), .Z(npu_inst_pe_1_4_6_N77) );
  AND2_X1 npu_inst_pe_1_4_6_U133 ( .A1(npu_inst_pe_1_4_6_add_69_carry_4_), 
        .A2(npu_inst_pe_1_4_6_int_q_acc_4_), .ZN(
        npu_inst_pe_1_4_6_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_4_6_U132 ( .A(npu_inst_pe_1_4_6_int_q_acc_5_), .B(
        npu_inst_pe_1_4_6_add_69_carry_5_), .Z(npu_inst_pe_1_4_6_N78) );
  AND2_X1 npu_inst_pe_1_4_6_U131 ( .A1(npu_inst_pe_1_4_6_add_69_carry_5_), 
        .A2(npu_inst_pe_1_4_6_int_q_acc_5_), .ZN(
        npu_inst_pe_1_4_6_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_4_6_U130 ( .A(npu_inst_pe_1_4_6_int_q_acc_6_), .B(
        npu_inst_pe_1_4_6_add_69_carry_6_), .Z(npu_inst_pe_1_4_6_N79) );
  AND2_X1 npu_inst_pe_1_4_6_U129 ( .A1(npu_inst_pe_1_4_6_add_69_carry_6_), 
        .A2(npu_inst_pe_1_4_6_int_q_acc_6_), .ZN(
        npu_inst_pe_1_4_6_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_4_6_U128 ( .A(npu_inst_pe_1_4_6_int_q_acc_7_), .B(
        npu_inst_pe_1_4_6_add_69_carry_7_), .Z(npu_inst_pe_1_4_6_N80) );
  XNOR2_X1 npu_inst_pe_1_4_6_U127 ( .A(npu_inst_pe_1_4_6_sub_67_carry_2_), .B(
        npu_inst_pe_1_4_6_int_q_acc_2_), .ZN(npu_inst_pe_1_4_6_N67) );
  OR2_X1 npu_inst_pe_1_4_6_U126 ( .A1(npu_inst_pe_1_4_6_int_q_acc_2_), .A2(
        npu_inst_pe_1_4_6_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_4_6_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_4_6_U125 ( .A(npu_inst_pe_1_4_6_sub_67_carry_3_), .B(
        npu_inst_pe_1_4_6_int_q_acc_3_), .ZN(npu_inst_pe_1_4_6_N68) );
  OR2_X1 npu_inst_pe_1_4_6_U124 ( .A1(npu_inst_pe_1_4_6_int_q_acc_3_), .A2(
        npu_inst_pe_1_4_6_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_4_6_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_4_6_U123 ( .A(npu_inst_pe_1_4_6_sub_67_carry_4_), .B(
        npu_inst_pe_1_4_6_int_q_acc_4_), .ZN(npu_inst_pe_1_4_6_N69) );
  OR2_X1 npu_inst_pe_1_4_6_U122 ( .A1(npu_inst_pe_1_4_6_int_q_acc_4_), .A2(
        npu_inst_pe_1_4_6_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_4_6_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_4_6_U121 ( .A(npu_inst_pe_1_4_6_sub_67_carry_5_), .B(
        npu_inst_pe_1_4_6_int_q_acc_5_), .ZN(npu_inst_pe_1_4_6_N70) );
  OR2_X1 npu_inst_pe_1_4_6_U120 ( .A1(npu_inst_pe_1_4_6_int_q_acc_5_), .A2(
        npu_inst_pe_1_4_6_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_4_6_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_4_6_U119 ( .A(npu_inst_pe_1_4_6_sub_67_carry_6_), .B(
        npu_inst_pe_1_4_6_int_q_acc_6_), .ZN(npu_inst_pe_1_4_6_N71) );
  OR2_X1 npu_inst_pe_1_4_6_U118 ( .A1(npu_inst_pe_1_4_6_int_q_acc_6_), .A2(
        npu_inst_pe_1_4_6_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_4_6_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_4_6_U117 ( .A(npu_inst_pe_1_4_6_int_q_acc_7_), .B(
        npu_inst_pe_1_4_6_sub_67_carry_7_), .ZN(npu_inst_pe_1_4_6_N72) );
  INV_X1 npu_inst_pe_1_4_6_U116 ( .A(npu_inst_n77), .ZN(npu_inst_pe_1_4_6_n7)
         );
  INV_X1 npu_inst_pe_1_4_6_U115 ( .A(npu_inst_pe_1_4_6_n7), .ZN(
        npu_inst_pe_1_4_6_n6) );
  INV_X1 npu_inst_pe_1_4_6_U114 ( .A(npu_inst_n55), .ZN(npu_inst_pe_1_4_6_n3)
         );
  AOI22_X1 npu_inst_pe_1_4_6_U113 ( .A1(npu_inst_int_data_y_5__6__0_), .A2(
        npu_inst_pe_1_4_6_n58), .B1(npu_inst_pe_1_4_6_n119), .B2(
        npu_inst_pe_1_4_6_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_4_6_n57) );
  INV_X1 npu_inst_pe_1_4_6_U112 ( .A(npu_inst_pe_1_4_6_n57), .ZN(
        npu_inst_pe_1_4_6_n108) );
  AOI22_X1 npu_inst_pe_1_4_6_U111 ( .A1(npu_inst_int_data_y_5__6__0_), .A2(
        npu_inst_pe_1_4_6_n54), .B1(npu_inst_pe_1_4_6_n118), .B2(
        npu_inst_pe_1_4_6_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_4_6_n53) );
  INV_X1 npu_inst_pe_1_4_6_U110 ( .A(npu_inst_pe_1_4_6_n53), .ZN(
        npu_inst_pe_1_4_6_n109) );
  AOI22_X1 npu_inst_pe_1_4_6_U107 ( .A1(npu_inst_int_data_y_5__6__0_), .A2(
        npu_inst_pe_1_4_6_n50), .B1(npu_inst_pe_1_4_6_n117), .B2(
        npu_inst_pe_1_4_6_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_4_6_n49) );
  INV_X1 npu_inst_pe_1_4_6_U106 ( .A(npu_inst_pe_1_4_6_n49), .ZN(
        npu_inst_pe_1_4_6_n110) );
  AOI22_X1 npu_inst_pe_1_4_6_U105 ( .A1(npu_inst_int_data_y_5__6__0_), .A2(
        npu_inst_pe_1_4_6_n46), .B1(npu_inst_pe_1_4_6_n116), .B2(
        npu_inst_pe_1_4_6_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_4_6_n45) );
  INV_X1 npu_inst_pe_1_4_6_U104 ( .A(npu_inst_pe_1_4_6_n45), .ZN(
        npu_inst_pe_1_4_6_n111) );
  AOI22_X1 npu_inst_pe_1_4_6_U103 ( .A1(npu_inst_int_data_y_5__6__0_), .A2(
        npu_inst_pe_1_4_6_n42), .B1(npu_inst_pe_1_4_6_n115), .B2(
        npu_inst_pe_1_4_6_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_4_6_n41) );
  INV_X1 npu_inst_pe_1_4_6_U102 ( .A(npu_inst_pe_1_4_6_n41), .ZN(
        npu_inst_pe_1_4_6_n112) );
  AOI22_X1 npu_inst_pe_1_4_6_U101 ( .A1(npu_inst_int_data_y_5__6__1_), .A2(
        npu_inst_pe_1_4_6_n58), .B1(npu_inst_pe_1_4_6_n119), .B2(
        npu_inst_pe_1_4_6_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_4_6_n59) );
  INV_X1 npu_inst_pe_1_4_6_U100 ( .A(npu_inst_pe_1_4_6_n59), .ZN(
        npu_inst_pe_1_4_6_n102) );
  AOI22_X1 npu_inst_pe_1_4_6_U99 ( .A1(npu_inst_int_data_y_5__6__1_), .A2(
        npu_inst_pe_1_4_6_n54), .B1(npu_inst_pe_1_4_6_n118), .B2(
        npu_inst_pe_1_4_6_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_4_6_n55) );
  INV_X1 npu_inst_pe_1_4_6_U98 ( .A(npu_inst_pe_1_4_6_n55), .ZN(
        npu_inst_pe_1_4_6_n103) );
  AOI22_X1 npu_inst_pe_1_4_6_U97 ( .A1(npu_inst_int_data_y_5__6__1_), .A2(
        npu_inst_pe_1_4_6_n50), .B1(npu_inst_pe_1_4_6_n117), .B2(
        npu_inst_pe_1_4_6_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_4_6_n51) );
  INV_X1 npu_inst_pe_1_4_6_U96 ( .A(npu_inst_pe_1_4_6_n51), .ZN(
        npu_inst_pe_1_4_6_n104) );
  AOI22_X1 npu_inst_pe_1_4_6_U95 ( .A1(npu_inst_int_data_y_5__6__1_), .A2(
        npu_inst_pe_1_4_6_n46), .B1(npu_inst_pe_1_4_6_n116), .B2(
        npu_inst_pe_1_4_6_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_4_6_n47) );
  INV_X1 npu_inst_pe_1_4_6_U94 ( .A(npu_inst_pe_1_4_6_n47), .ZN(
        npu_inst_pe_1_4_6_n105) );
  AOI22_X1 npu_inst_pe_1_4_6_U93 ( .A1(npu_inst_int_data_y_5__6__1_), .A2(
        npu_inst_pe_1_4_6_n42), .B1(npu_inst_pe_1_4_6_n115), .B2(
        npu_inst_pe_1_4_6_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_4_6_n43) );
  INV_X1 npu_inst_pe_1_4_6_U92 ( .A(npu_inst_pe_1_4_6_n43), .ZN(
        npu_inst_pe_1_4_6_n106) );
  AOI22_X1 npu_inst_pe_1_4_6_U91 ( .A1(npu_inst_pe_1_4_6_n38), .A2(
        npu_inst_int_data_y_5__6__1_), .B1(npu_inst_pe_1_4_6_n114), .B2(
        npu_inst_pe_1_4_6_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_4_6_n39) );
  INV_X1 npu_inst_pe_1_4_6_U90 ( .A(npu_inst_pe_1_4_6_n39), .ZN(
        npu_inst_pe_1_4_6_n107) );
  AOI22_X1 npu_inst_pe_1_4_6_U89 ( .A1(npu_inst_pe_1_4_6_n38), .A2(
        npu_inst_int_data_y_5__6__0_), .B1(npu_inst_pe_1_4_6_n114), .B2(
        npu_inst_pe_1_4_6_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_4_6_n37) );
  INV_X1 npu_inst_pe_1_4_6_U88 ( .A(npu_inst_pe_1_4_6_n37), .ZN(
        npu_inst_pe_1_4_6_n113) );
  NAND2_X1 npu_inst_pe_1_4_6_U87 ( .A1(npu_inst_pe_1_4_6_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_4_6_n60), .ZN(npu_inst_pe_1_4_6_n74) );
  OAI21_X1 npu_inst_pe_1_4_6_U86 ( .B1(npu_inst_pe_1_4_6_n63), .B2(
        npu_inst_pe_1_4_6_n60), .A(npu_inst_pe_1_4_6_n74), .ZN(
        npu_inst_pe_1_4_6_n97) );
  NAND2_X1 npu_inst_pe_1_4_6_U85 ( .A1(npu_inst_pe_1_4_6_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_4_6_n60), .ZN(npu_inst_pe_1_4_6_n73) );
  OAI21_X1 npu_inst_pe_1_4_6_U84 ( .B1(npu_inst_pe_1_4_6_n61), .B2(
        npu_inst_pe_1_4_6_n60), .A(npu_inst_pe_1_4_6_n73), .ZN(
        npu_inst_pe_1_4_6_n96) );
  NAND2_X1 npu_inst_pe_1_4_6_U83 ( .A1(npu_inst_pe_1_4_6_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_4_6_n56), .ZN(npu_inst_pe_1_4_6_n72) );
  OAI21_X1 npu_inst_pe_1_4_6_U82 ( .B1(npu_inst_pe_1_4_6_n63), .B2(
        npu_inst_pe_1_4_6_n56), .A(npu_inst_pe_1_4_6_n72), .ZN(
        npu_inst_pe_1_4_6_n95) );
  NAND2_X1 npu_inst_pe_1_4_6_U81 ( .A1(npu_inst_pe_1_4_6_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_4_6_n56), .ZN(npu_inst_pe_1_4_6_n71) );
  OAI21_X1 npu_inst_pe_1_4_6_U80 ( .B1(npu_inst_pe_1_4_6_n61), .B2(
        npu_inst_pe_1_4_6_n56), .A(npu_inst_pe_1_4_6_n71), .ZN(
        npu_inst_pe_1_4_6_n94) );
  NAND2_X1 npu_inst_pe_1_4_6_U79 ( .A1(npu_inst_pe_1_4_6_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_4_6_n52), .ZN(npu_inst_pe_1_4_6_n70) );
  OAI21_X1 npu_inst_pe_1_4_6_U78 ( .B1(npu_inst_pe_1_4_6_n63), .B2(
        npu_inst_pe_1_4_6_n52), .A(npu_inst_pe_1_4_6_n70), .ZN(
        npu_inst_pe_1_4_6_n93) );
  NAND2_X1 npu_inst_pe_1_4_6_U77 ( .A1(npu_inst_pe_1_4_6_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_4_6_n52), .ZN(npu_inst_pe_1_4_6_n69) );
  OAI21_X1 npu_inst_pe_1_4_6_U76 ( .B1(npu_inst_pe_1_4_6_n61), .B2(
        npu_inst_pe_1_4_6_n52), .A(npu_inst_pe_1_4_6_n69), .ZN(
        npu_inst_pe_1_4_6_n92) );
  NAND2_X1 npu_inst_pe_1_4_6_U75 ( .A1(npu_inst_pe_1_4_6_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_4_6_n48), .ZN(npu_inst_pe_1_4_6_n68) );
  OAI21_X1 npu_inst_pe_1_4_6_U74 ( .B1(npu_inst_pe_1_4_6_n63), .B2(
        npu_inst_pe_1_4_6_n48), .A(npu_inst_pe_1_4_6_n68), .ZN(
        npu_inst_pe_1_4_6_n91) );
  NAND2_X1 npu_inst_pe_1_4_6_U73 ( .A1(npu_inst_pe_1_4_6_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_4_6_n48), .ZN(npu_inst_pe_1_4_6_n67) );
  OAI21_X1 npu_inst_pe_1_4_6_U72 ( .B1(npu_inst_pe_1_4_6_n61), .B2(
        npu_inst_pe_1_4_6_n48), .A(npu_inst_pe_1_4_6_n67), .ZN(
        npu_inst_pe_1_4_6_n90) );
  NAND2_X1 npu_inst_pe_1_4_6_U71 ( .A1(npu_inst_pe_1_4_6_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_4_6_n44), .ZN(npu_inst_pe_1_4_6_n66) );
  OAI21_X1 npu_inst_pe_1_4_6_U70 ( .B1(npu_inst_pe_1_4_6_n63), .B2(
        npu_inst_pe_1_4_6_n44), .A(npu_inst_pe_1_4_6_n66), .ZN(
        npu_inst_pe_1_4_6_n89) );
  NAND2_X1 npu_inst_pe_1_4_6_U69 ( .A1(npu_inst_pe_1_4_6_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_4_6_n44), .ZN(npu_inst_pe_1_4_6_n65) );
  OAI21_X1 npu_inst_pe_1_4_6_U68 ( .B1(npu_inst_pe_1_4_6_n61), .B2(
        npu_inst_pe_1_4_6_n44), .A(npu_inst_pe_1_4_6_n65), .ZN(
        npu_inst_pe_1_4_6_n88) );
  NAND2_X1 npu_inst_pe_1_4_6_U67 ( .A1(npu_inst_pe_1_4_6_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_4_6_n40), .ZN(npu_inst_pe_1_4_6_n64) );
  OAI21_X1 npu_inst_pe_1_4_6_U66 ( .B1(npu_inst_pe_1_4_6_n63), .B2(
        npu_inst_pe_1_4_6_n40), .A(npu_inst_pe_1_4_6_n64), .ZN(
        npu_inst_pe_1_4_6_n87) );
  NAND2_X1 npu_inst_pe_1_4_6_U65 ( .A1(npu_inst_pe_1_4_6_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_4_6_n40), .ZN(npu_inst_pe_1_4_6_n62) );
  OAI21_X1 npu_inst_pe_1_4_6_U64 ( .B1(npu_inst_pe_1_4_6_n61), .B2(
        npu_inst_pe_1_4_6_n40), .A(npu_inst_pe_1_4_6_n62), .ZN(
        npu_inst_pe_1_4_6_n86) );
  AND2_X1 npu_inst_pe_1_4_6_U63 ( .A1(npu_inst_pe_1_4_6_N93), .A2(npu_inst_n55), .ZN(npu_inst_int_data_y_4__6__0_) );
  AND2_X1 npu_inst_pe_1_4_6_U62 ( .A1(npu_inst_n55), .A2(npu_inst_pe_1_4_6_N94), .ZN(npu_inst_int_data_y_4__6__1_) );
  NOR3_X1 npu_inst_pe_1_4_6_U61 ( .A1(npu_inst_pe_1_4_6_n26), .A2(npu_inst_n55), .A3(npu_inst_int_ckg[25]), .ZN(npu_inst_pe_1_4_6_n85) );
  OR2_X1 npu_inst_pe_1_4_6_U60 ( .A1(npu_inst_pe_1_4_6_n85), .A2(
        npu_inst_pe_1_4_6_n2), .ZN(npu_inst_pe_1_4_6_N84) );
  AND2_X1 npu_inst_pe_1_4_6_U59 ( .A1(npu_inst_pe_1_4_6_int_q_acc_0_), .A2(
        npu_inst_pe_1_4_6_n1), .ZN(npu_inst_int_data_res_4__6__0_) );
  AND2_X1 npu_inst_pe_1_4_6_U58 ( .A1(npu_inst_pe_1_4_6_n2), .A2(
        npu_inst_pe_1_4_6_int_q_acc_7_), .ZN(npu_inst_int_data_res_4__6__7_)
         );
  AND2_X1 npu_inst_pe_1_4_6_U57 ( .A1(npu_inst_pe_1_4_6_int_q_acc_1_), .A2(
        npu_inst_pe_1_4_6_n1), .ZN(npu_inst_int_data_res_4__6__1_) );
  AND2_X1 npu_inst_pe_1_4_6_U56 ( .A1(npu_inst_pe_1_4_6_int_q_acc_2_), .A2(
        npu_inst_pe_1_4_6_n1), .ZN(npu_inst_int_data_res_4__6__2_) );
  AND2_X1 npu_inst_pe_1_4_6_U55 ( .A1(npu_inst_pe_1_4_6_int_q_acc_3_), .A2(
        npu_inst_pe_1_4_6_n2), .ZN(npu_inst_int_data_res_4__6__3_) );
  AND2_X1 npu_inst_pe_1_4_6_U54 ( .A1(npu_inst_pe_1_4_6_int_q_acc_4_), .A2(
        npu_inst_pe_1_4_6_n2), .ZN(npu_inst_int_data_res_4__6__4_) );
  AND2_X1 npu_inst_pe_1_4_6_U53 ( .A1(npu_inst_pe_1_4_6_int_q_acc_5_), .A2(
        npu_inst_pe_1_4_6_n2), .ZN(npu_inst_int_data_res_4__6__5_) );
  AND2_X1 npu_inst_pe_1_4_6_U52 ( .A1(npu_inst_pe_1_4_6_int_q_acc_6_), .A2(
        npu_inst_pe_1_4_6_n2), .ZN(npu_inst_int_data_res_4__6__6_) );
  AOI222_X1 npu_inst_pe_1_4_6_U51 ( .A1(npu_inst_int_data_res_5__6__0_), .A2(
        npu_inst_pe_1_4_6_n1), .B1(npu_inst_pe_1_4_6_N73), .B2(
        npu_inst_pe_1_4_6_n76), .C1(npu_inst_pe_1_4_6_N65), .C2(
        npu_inst_pe_1_4_6_n77), .ZN(npu_inst_pe_1_4_6_n84) );
  INV_X1 npu_inst_pe_1_4_6_U50 ( .A(npu_inst_pe_1_4_6_n84), .ZN(
        npu_inst_pe_1_4_6_n101) );
  AOI222_X1 npu_inst_pe_1_4_6_U49 ( .A1(npu_inst_int_data_res_5__6__7_), .A2(
        npu_inst_pe_1_4_6_n1), .B1(npu_inst_pe_1_4_6_N80), .B2(
        npu_inst_pe_1_4_6_n76), .C1(npu_inst_pe_1_4_6_N72), .C2(
        npu_inst_pe_1_4_6_n77), .ZN(npu_inst_pe_1_4_6_n75) );
  INV_X1 npu_inst_pe_1_4_6_U48 ( .A(npu_inst_pe_1_4_6_n75), .ZN(
        npu_inst_pe_1_4_6_n33) );
  AOI222_X1 npu_inst_pe_1_4_6_U47 ( .A1(npu_inst_int_data_res_5__6__1_), .A2(
        npu_inst_pe_1_4_6_n1), .B1(npu_inst_pe_1_4_6_N74), .B2(
        npu_inst_pe_1_4_6_n76), .C1(npu_inst_pe_1_4_6_N66), .C2(
        npu_inst_pe_1_4_6_n77), .ZN(npu_inst_pe_1_4_6_n83) );
  INV_X1 npu_inst_pe_1_4_6_U46 ( .A(npu_inst_pe_1_4_6_n83), .ZN(
        npu_inst_pe_1_4_6_n100) );
  AOI222_X1 npu_inst_pe_1_4_6_U45 ( .A1(npu_inst_int_data_res_5__6__2_), .A2(
        npu_inst_pe_1_4_6_n1), .B1(npu_inst_pe_1_4_6_N75), .B2(
        npu_inst_pe_1_4_6_n76), .C1(npu_inst_pe_1_4_6_N67), .C2(
        npu_inst_pe_1_4_6_n77), .ZN(npu_inst_pe_1_4_6_n82) );
  INV_X1 npu_inst_pe_1_4_6_U44 ( .A(npu_inst_pe_1_4_6_n82), .ZN(
        npu_inst_pe_1_4_6_n99) );
  AOI222_X1 npu_inst_pe_1_4_6_U43 ( .A1(npu_inst_int_data_res_5__6__3_), .A2(
        npu_inst_pe_1_4_6_n1), .B1(npu_inst_pe_1_4_6_N76), .B2(
        npu_inst_pe_1_4_6_n76), .C1(npu_inst_pe_1_4_6_N68), .C2(
        npu_inst_pe_1_4_6_n77), .ZN(npu_inst_pe_1_4_6_n81) );
  INV_X1 npu_inst_pe_1_4_6_U42 ( .A(npu_inst_pe_1_4_6_n81), .ZN(
        npu_inst_pe_1_4_6_n98) );
  AOI222_X1 npu_inst_pe_1_4_6_U41 ( .A1(npu_inst_int_data_res_5__6__4_), .A2(
        npu_inst_pe_1_4_6_n1), .B1(npu_inst_pe_1_4_6_N77), .B2(
        npu_inst_pe_1_4_6_n76), .C1(npu_inst_pe_1_4_6_N69), .C2(
        npu_inst_pe_1_4_6_n77), .ZN(npu_inst_pe_1_4_6_n80) );
  INV_X1 npu_inst_pe_1_4_6_U40 ( .A(npu_inst_pe_1_4_6_n80), .ZN(
        npu_inst_pe_1_4_6_n36) );
  AOI222_X1 npu_inst_pe_1_4_6_U39 ( .A1(npu_inst_int_data_res_5__6__5_), .A2(
        npu_inst_pe_1_4_6_n1), .B1(npu_inst_pe_1_4_6_N78), .B2(
        npu_inst_pe_1_4_6_n76), .C1(npu_inst_pe_1_4_6_N70), .C2(
        npu_inst_pe_1_4_6_n77), .ZN(npu_inst_pe_1_4_6_n79) );
  INV_X1 npu_inst_pe_1_4_6_U38 ( .A(npu_inst_pe_1_4_6_n79), .ZN(
        npu_inst_pe_1_4_6_n35) );
  AOI222_X1 npu_inst_pe_1_4_6_U37 ( .A1(npu_inst_int_data_res_5__6__6_), .A2(
        npu_inst_pe_1_4_6_n1), .B1(npu_inst_pe_1_4_6_N79), .B2(
        npu_inst_pe_1_4_6_n76), .C1(npu_inst_pe_1_4_6_N71), .C2(
        npu_inst_pe_1_4_6_n77), .ZN(npu_inst_pe_1_4_6_n78) );
  INV_X1 npu_inst_pe_1_4_6_U36 ( .A(npu_inst_pe_1_4_6_n78), .ZN(
        npu_inst_pe_1_4_6_n34) );
  INV_X1 npu_inst_pe_1_4_6_U35 ( .A(npu_inst_pe_1_4_6_int_data_1_), .ZN(
        npu_inst_pe_1_4_6_n14) );
  AND2_X1 npu_inst_pe_1_4_6_U34 ( .A1(npu_inst_int_data_x_4__6__1_), .A2(
        npu_inst_pe_1_4_6_int_q_weight_1_), .ZN(npu_inst_pe_1_4_6_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_4_6_U33 ( .A1(npu_inst_int_data_x_4__6__0_), .A2(
        npu_inst_pe_1_4_6_int_q_weight_1_), .ZN(npu_inst_pe_1_4_6_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_4_6_U32 ( .A1(npu_inst_n55), .A2(
        npu_inst_int_data_y_5__6__1_), .B1(npu_inst_pe_1_4_6_n3), .B2(
        npu_inst_int_data_x_4__7__1_), .ZN(npu_inst_pe_1_4_6_n63) );
  AOI22_X1 npu_inst_pe_1_4_6_U31 ( .A1(npu_inst_n55), .A2(
        npu_inst_int_data_y_5__6__0_), .B1(npu_inst_pe_1_4_6_n3), .B2(
        npu_inst_int_data_x_4__7__0_), .ZN(npu_inst_pe_1_4_6_n61) );
  INV_X1 npu_inst_pe_1_4_6_U30 ( .A(npu_inst_pe_1_4_6_int_data_0_), .ZN(
        npu_inst_pe_1_4_6_n13) );
  INV_X1 npu_inst_pe_1_4_6_U29 ( .A(npu_inst_n69), .ZN(npu_inst_pe_1_4_6_n5)
         );
  OR3_X1 npu_inst_pe_1_4_6_U28 ( .A1(npu_inst_pe_1_4_6_n6), .A2(
        npu_inst_pe_1_4_6_n8), .A3(npu_inst_pe_1_4_6_n5), .ZN(
        npu_inst_pe_1_4_6_n56) );
  OR3_X1 npu_inst_pe_1_4_6_U27 ( .A1(npu_inst_pe_1_4_6_n5), .A2(
        npu_inst_pe_1_4_6_n8), .A3(npu_inst_pe_1_4_6_n7), .ZN(
        npu_inst_pe_1_4_6_n48) );
  INV_X1 npu_inst_pe_1_4_6_U26 ( .A(npu_inst_pe_1_4_6_n5), .ZN(
        npu_inst_pe_1_4_6_n4) );
  OR3_X1 npu_inst_pe_1_4_6_U25 ( .A1(npu_inst_pe_1_4_6_n4), .A2(
        npu_inst_pe_1_4_6_n8), .A3(npu_inst_pe_1_4_6_n7), .ZN(
        npu_inst_pe_1_4_6_n52) );
  OR3_X1 npu_inst_pe_1_4_6_U24 ( .A1(npu_inst_pe_1_4_6_n6), .A2(
        npu_inst_pe_1_4_6_n8), .A3(npu_inst_pe_1_4_6_n4), .ZN(
        npu_inst_pe_1_4_6_n60) );
  NOR2_X1 npu_inst_pe_1_4_6_U23 ( .A1(npu_inst_pe_1_4_6_n60), .A2(
        npu_inst_pe_1_4_6_n3), .ZN(npu_inst_pe_1_4_6_n58) );
  NOR2_X1 npu_inst_pe_1_4_6_U22 ( .A1(npu_inst_pe_1_4_6_n56), .A2(
        npu_inst_pe_1_4_6_n3), .ZN(npu_inst_pe_1_4_6_n54) );
  NOR2_X1 npu_inst_pe_1_4_6_U21 ( .A1(npu_inst_pe_1_4_6_n52), .A2(
        npu_inst_pe_1_4_6_n3), .ZN(npu_inst_pe_1_4_6_n50) );
  NOR2_X1 npu_inst_pe_1_4_6_U20 ( .A1(npu_inst_pe_1_4_6_n48), .A2(
        npu_inst_pe_1_4_6_n3), .ZN(npu_inst_pe_1_4_6_n46) );
  NOR2_X1 npu_inst_pe_1_4_6_U19 ( .A1(npu_inst_pe_1_4_6_n40), .A2(
        npu_inst_pe_1_4_6_n3), .ZN(npu_inst_pe_1_4_6_n38) );
  NOR2_X1 npu_inst_pe_1_4_6_U18 ( .A1(npu_inst_pe_1_4_6_n44), .A2(
        npu_inst_pe_1_4_6_n3), .ZN(npu_inst_pe_1_4_6_n42) );
  BUF_X1 npu_inst_pe_1_4_6_U17 ( .A(npu_inst_n98), .Z(npu_inst_pe_1_4_6_n8) );
  INV_X1 npu_inst_pe_1_4_6_U16 ( .A(npu_inst_n124), .ZN(npu_inst_pe_1_4_6_n12)
         );
  INV_X1 npu_inst_pe_1_4_6_U15 ( .A(npu_inst_pe_1_4_6_n38), .ZN(
        npu_inst_pe_1_4_6_n114) );
  INV_X1 npu_inst_pe_1_4_6_U14 ( .A(npu_inst_pe_1_4_6_n58), .ZN(
        npu_inst_pe_1_4_6_n119) );
  INV_X1 npu_inst_pe_1_4_6_U13 ( .A(npu_inst_pe_1_4_6_n54), .ZN(
        npu_inst_pe_1_4_6_n118) );
  INV_X1 npu_inst_pe_1_4_6_U12 ( .A(npu_inst_pe_1_4_6_n50), .ZN(
        npu_inst_pe_1_4_6_n117) );
  INV_X1 npu_inst_pe_1_4_6_U11 ( .A(npu_inst_pe_1_4_6_n46), .ZN(
        npu_inst_pe_1_4_6_n116) );
  INV_X1 npu_inst_pe_1_4_6_U10 ( .A(npu_inst_pe_1_4_6_n42), .ZN(
        npu_inst_pe_1_4_6_n115) );
  BUF_X1 npu_inst_pe_1_4_6_U9 ( .A(npu_inst_n19), .Z(npu_inst_pe_1_4_6_n2) );
  BUF_X1 npu_inst_pe_1_4_6_U8 ( .A(npu_inst_n19), .Z(npu_inst_pe_1_4_6_n1) );
  BUF_X1 npu_inst_pe_1_4_6_U7 ( .A(npu_inst_pe_1_4_6_n12), .Z(
        npu_inst_pe_1_4_6_n11) );
  BUF_X1 npu_inst_pe_1_4_6_U6 ( .A(npu_inst_pe_1_4_6_n12), .Z(
        npu_inst_pe_1_4_6_n10) );
  BUF_X1 npu_inst_pe_1_4_6_U5 ( .A(npu_inst_pe_1_4_6_n12), .Z(
        npu_inst_pe_1_4_6_n9) );
  NOR2_X1 npu_inst_pe_1_4_6_U4 ( .A1(npu_inst_pe_1_4_6_int_q_weight_0_), .A2(
        npu_inst_pe_1_4_6_n1), .ZN(npu_inst_pe_1_4_6_n76) );
  NOR2_X1 npu_inst_pe_1_4_6_U3 ( .A1(npu_inst_pe_1_4_6_n27), .A2(
        npu_inst_pe_1_4_6_n1), .ZN(npu_inst_pe_1_4_6_n77) );
  FA_X1 npu_inst_pe_1_4_6_sub_67_U2_1 ( .A(npu_inst_pe_1_4_6_int_q_acc_1_), 
        .B(npu_inst_pe_1_4_6_n14), .CI(npu_inst_pe_1_4_6_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_4_6_sub_67_carry_2_), .S(npu_inst_pe_1_4_6_N66) );
  FA_X1 npu_inst_pe_1_4_6_add_69_U1_1 ( .A(npu_inst_pe_1_4_6_int_q_acc_1_), 
        .B(npu_inst_pe_1_4_6_int_data_1_), .CI(
        npu_inst_pe_1_4_6_add_69_carry_1_), .CO(
        npu_inst_pe_1_4_6_add_69_carry_2_), .S(npu_inst_pe_1_4_6_N74) );
  NAND3_X1 npu_inst_pe_1_4_6_U109 ( .A1(npu_inst_pe_1_4_6_n5), .A2(
        npu_inst_pe_1_4_6_n7), .A3(npu_inst_pe_1_4_6_n8), .ZN(
        npu_inst_pe_1_4_6_n44) );
  NAND3_X1 npu_inst_pe_1_4_6_U108 ( .A1(npu_inst_pe_1_4_6_n4), .A2(
        npu_inst_pe_1_4_6_n7), .A3(npu_inst_pe_1_4_6_n8), .ZN(
        npu_inst_pe_1_4_6_n40) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_4_6_n34), .CK(
        npu_inst_pe_1_4_6_net3688), .RN(npu_inst_pe_1_4_6_n9), .Q(
        npu_inst_pe_1_4_6_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_4_6_n35), .CK(
        npu_inst_pe_1_4_6_net3688), .RN(npu_inst_pe_1_4_6_n9), .Q(
        npu_inst_pe_1_4_6_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_4_6_n36), .CK(
        npu_inst_pe_1_4_6_net3688), .RN(npu_inst_pe_1_4_6_n9), .Q(
        npu_inst_pe_1_4_6_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_4_6_n98), .CK(
        npu_inst_pe_1_4_6_net3688), .RN(npu_inst_pe_1_4_6_n9), .Q(
        npu_inst_pe_1_4_6_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_4_6_n99), .CK(
        npu_inst_pe_1_4_6_net3688), .RN(npu_inst_pe_1_4_6_n9), .Q(
        npu_inst_pe_1_4_6_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_4_6_n100), 
        .CK(npu_inst_pe_1_4_6_net3688), .RN(npu_inst_pe_1_4_6_n9), .Q(
        npu_inst_pe_1_4_6_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_4_6_n33), .CK(
        npu_inst_pe_1_4_6_net3688), .RN(npu_inst_pe_1_4_6_n9), .Q(
        npu_inst_pe_1_4_6_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_4_6_n101), 
        .CK(npu_inst_pe_1_4_6_net3688), .RN(npu_inst_pe_1_4_6_n9), .Q(
        npu_inst_pe_1_4_6_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_weight_reg_0_ ( .D(npu_inst_n110), .CK(
        npu_inst_pe_1_4_6_net3694), .RN(npu_inst_pe_1_4_6_n9), .Q(
        npu_inst_pe_1_4_6_int_q_weight_0_), .QN(npu_inst_pe_1_4_6_n27) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_weight_reg_1_ ( .D(npu_inst_n116), .CK(
        npu_inst_pe_1_4_6_net3694), .RN(npu_inst_pe_1_4_6_n9), .Q(
        npu_inst_pe_1_4_6_int_q_weight_1_), .QN(npu_inst_pe_1_4_6_n26) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_4_6_n113), 
        .CK(npu_inst_pe_1_4_6_net3694), .RN(npu_inst_pe_1_4_6_n9), .Q(
        npu_inst_pe_1_4_6_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_4_6_n107), 
        .CK(npu_inst_pe_1_4_6_net3694), .RN(npu_inst_pe_1_4_6_n9), .Q(
        npu_inst_pe_1_4_6_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_4_6_n112), 
        .CK(npu_inst_pe_1_4_6_net3694), .RN(npu_inst_pe_1_4_6_n10), .Q(
        npu_inst_pe_1_4_6_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_4_6_n106), 
        .CK(npu_inst_pe_1_4_6_net3694), .RN(npu_inst_pe_1_4_6_n10), .Q(
        npu_inst_pe_1_4_6_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_4_6_n111), 
        .CK(npu_inst_pe_1_4_6_net3694), .RN(npu_inst_pe_1_4_6_n10), .Q(
        npu_inst_pe_1_4_6_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_4_6_n105), 
        .CK(npu_inst_pe_1_4_6_net3694), .RN(npu_inst_pe_1_4_6_n10), .Q(
        npu_inst_pe_1_4_6_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_4_6_n110), 
        .CK(npu_inst_pe_1_4_6_net3694), .RN(npu_inst_pe_1_4_6_n10), .Q(
        npu_inst_pe_1_4_6_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_4_6_n104), 
        .CK(npu_inst_pe_1_4_6_net3694), .RN(npu_inst_pe_1_4_6_n10), .Q(
        npu_inst_pe_1_4_6_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_4_6_n109), 
        .CK(npu_inst_pe_1_4_6_net3694), .RN(npu_inst_pe_1_4_6_n10), .Q(
        npu_inst_pe_1_4_6_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_4_6_n103), 
        .CK(npu_inst_pe_1_4_6_net3694), .RN(npu_inst_pe_1_4_6_n10), .Q(
        npu_inst_pe_1_4_6_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_4_6_n108), 
        .CK(npu_inst_pe_1_4_6_net3694), .RN(npu_inst_pe_1_4_6_n10), .Q(
        npu_inst_pe_1_4_6_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_4_6_n102), 
        .CK(npu_inst_pe_1_4_6_net3694), .RN(npu_inst_pe_1_4_6_n10), .Q(
        npu_inst_pe_1_4_6_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_4_6_n86), 
        .CK(npu_inst_pe_1_4_6_net3694), .RN(npu_inst_pe_1_4_6_n10), .Q(
        npu_inst_pe_1_4_6_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_4_6_n87), 
        .CK(npu_inst_pe_1_4_6_net3694), .RN(npu_inst_pe_1_4_6_n10), .Q(
        npu_inst_pe_1_4_6_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_4_6_n88), 
        .CK(npu_inst_pe_1_4_6_net3694), .RN(npu_inst_pe_1_4_6_n11), .Q(
        npu_inst_pe_1_4_6_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_4_6_n89), 
        .CK(npu_inst_pe_1_4_6_net3694), .RN(npu_inst_pe_1_4_6_n11), .Q(
        npu_inst_pe_1_4_6_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_4_6_n90), 
        .CK(npu_inst_pe_1_4_6_net3694), .RN(npu_inst_pe_1_4_6_n11), .Q(
        npu_inst_pe_1_4_6_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_4_6_n91), 
        .CK(npu_inst_pe_1_4_6_net3694), .RN(npu_inst_pe_1_4_6_n11), .Q(
        npu_inst_pe_1_4_6_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_4_6_n92), 
        .CK(npu_inst_pe_1_4_6_net3694), .RN(npu_inst_pe_1_4_6_n11), .Q(
        npu_inst_pe_1_4_6_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_4_6_n93), 
        .CK(npu_inst_pe_1_4_6_net3694), .RN(npu_inst_pe_1_4_6_n11), .Q(
        npu_inst_pe_1_4_6_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_4_6_n94), 
        .CK(npu_inst_pe_1_4_6_net3694), .RN(npu_inst_pe_1_4_6_n11), .Q(
        npu_inst_pe_1_4_6_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_4_6_n95), 
        .CK(npu_inst_pe_1_4_6_net3694), .RN(npu_inst_pe_1_4_6_n11), .Q(
        npu_inst_pe_1_4_6_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_4_6_n96), 
        .CK(npu_inst_pe_1_4_6_net3694), .RN(npu_inst_pe_1_4_6_n11), .Q(
        npu_inst_pe_1_4_6_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_4_6_n97), 
        .CK(npu_inst_pe_1_4_6_net3694), .RN(npu_inst_pe_1_4_6_n11), .Q(
        npu_inst_pe_1_4_6_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_4_6_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_4_6_N84), .SE(1'b0), .GCK(npu_inst_pe_1_4_6_net3688) );
  CLKGATETST_X1 npu_inst_pe_1_4_6_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n63), .SE(1'b0), .GCK(npu_inst_pe_1_4_6_net3694) );
  MUX2_X1 npu_inst_pe_1_4_7_U162 ( .A(npu_inst_pe_1_4_7_n32), .B(
        npu_inst_pe_1_4_7_n29), .S(npu_inst_pe_1_4_7_n8), .Z(
        npu_inst_pe_1_4_7_N93) );
  MUX2_X1 npu_inst_pe_1_4_7_U161 ( .A(npu_inst_pe_1_4_7_n31), .B(
        npu_inst_pe_1_4_7_n30), .S(npu_inst_pe_1_4_7_n6), .Z(
        npu_inst_pe_1_4_7_n32) );
  MUX2_X1 npu_inst_pe_1_4_7_U160 ( .A(npu_inst_pe_1_4_7_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_4_7_int_q_reg_v_1__0_), .S(npu_inst_pe_1_4_7_n4), .Z(
        npu_inst_pe_1_4_7_n31) );
  MUX2_X1 npu_inst_pe_1_4_7_U159 ( .A(npu_inst_pe_1_4_7_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_4_7_int_q_reg_v_3__0_), .S(npu_inst_pe_1_4_7_n4), .Z(
        npu_inst_pe_1_4_7_n30) );
  MUX2_X1 npu_inst_pe_1_4_7_U158 ( .A(npu_inst_pe_1_4_7_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_4_7_int_q_reg_v_5__0_), .S(npu_inst_pe_1_4_7_n4), .Z(
        npu_inst_pe_1_4_7_n29) );
  MUX2_X1 npu_inst_pe_1_4_7_U157 ( .A(npu_inst_pe_1_4_7_n28), .B(
        npu_inst_pe_1_4_7_n23), .S(npu_inst_pe_1_4_7_n8), .Z(
        npu_inst_pe_1_4_7_N94) );
  MUX2_X1 npu_inst_pe_1_4_7_U156 ( .A(npu_inst_pe_1_4_7_n25), .B(
        npu_inst_pe_1_4_7_n24), .S(npu_inst_pe_1_4_7_n6), .Z(
        npu_inst_pe_1_4_7_n28) );
  MUX2_X1 npu_inst_pe_1_4_7_U155 ( .A(npu_inst_pe_1_4_7_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_4_7_int_q_reg_v_1__1_), .S(npu_inst_pe_1_4_7_n4), .Z(
        npu_inst_pe_1_4_7_n25) );
  MUX2_X1 npu_inst_pe_1_4_7_U154 ( .A(npu_inst_pe_1_4_7_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_4_7_int_q_reg_v_3__1_), .S(npu_inst_pe_1_4_7_n4), .Z(
        npu_inst_pe_1_4_7_n24) );
  MUX2_X1 npu_inst_pe_1_4_7_U153 ( .A(npu_inst_pe_1_4_7_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_4_7_int_q_reg_v_5__1_), .S(npu_inst_pe_1_4_7_n4), .Z(
        npu_inst_pe_1_4_7_n23) );
  MUX2_X1 npu_inst_pe_1_4_7_U152 ( .A(npu_inst_pe_1_4_7_n22), .B(
        npu_inst_pe_1_4_7_n19), .S(npu_inst_pe_1_4_7_n8), .Z(
        npu_inst_int_data_x_4__7__1_) );
  MUX2_X1 npu_inst_pe_1_4_7_U151 ( .A(npu_inst_pe_1_4_7_n21), .B(
        npu_inst_pe_1_4_7_n20), .S(npu_inst_pe_1_4_7_n6), .Z(
        npu_inst_pe_1_4_7_n22) );
  MUX2_X1 npu_inst_pe_1_4_7_U150 ( .A(npu_inst_pe_1_4_7_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_4_7_int_q_reg_h_1__1_), .S(npu_inst_pe_1_4_7_n4), .Z(
        npu_inst_pe_1_4_7_n21) );
  MUX2_X1 npu_inst_pe_1_4_7_U149 ( .A(npu_inst_pe_1_4_7_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_4_7_int_q_reg_h_3__1_), .S(npu_inst_pe_1_4_7_n4), .Z(
        npu_inst_pe_1_4_7_n20) );
  MUX2_X1 npu_inst_pe_1_4_7_U148 ( .A(npu_inst_pe_1_4_7_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_4_7_int_q_reg_h_5__1_), .S(npu_inst_pe_1_4_7_n4), .Z(
        npu_inst_pe_1_4_7_n19) );
  MUX2_X1 npu_inst_pe_1_4_7_U147 ( .A(npu_inst_pe_1_4_7_n18), .B(
        npu_inst_pe_1_4_7_n15), .S(npu_inst_pe_1_4_7_n8), .Z(
        npu_inst_int_data_x_4__7__0_) );
  MUX2_X1 npu_inst_pe_1_4_7_U146 ( .A(npu_inst_pe_1_4_7_n17), .B(
        npu_inst_pe_1_4_7_n16), .S(npu_inst_pe_1_4_7_n6), .Z(
        npu_inst_pe_1_4_7_n18) );
  MUX2_X1 npu_inst_pe_1_4_7_U145 ( .A(npu_inst_pe_1_4_7_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_4_7_int_q_reg_h_1__0_), .S(npu_inst_pe_1_4_7_n4), .Z(
        npu_inst_pe_1_4_7_n17) );
  MUX2_X1 npu_inst_pe_1_4_7_U144 ( .A(npu_inst_pe_1_4_7_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_4_7_int_q_reg_h_3__0_), .S(npu_inst_pe_1_4_7_n4), .Z(
        npu_inst_pe_1_4_7_n16) );
  MUX2_X1 npu_inst_pe_1_4_7_U143 ( .A(npu_inst_pe_1_4_7_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_4_7_int_q_reg_h_5__0_), .S(npu_inst_pe_1_4_7_n4), .Z(
        npu_inst_pe_1_4_7_n15) );
  XOR2_X1 npu_inst_pe_1_4_7_U142 ( .A(npu_inst_pe_1_4_7_int_data_0_), .B(
        npu_inst_pe_1_4_7_int_q_acc_0_), .Z(npu_inst_pe_1_4_7_N73) );
  AND2_X1 npu_inst_pe_1_4_7_U141 ( .A1(npu_inst_pe_1_4_7_int_q_acc_0_), .A2(
        npu_inst_pe_1_4_7_int_data_0_), .ZN(npu_inst_pe_1_4_7_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_4_7_U140 ( .A(npu_inst_pe_1_4_7_int_q_acc_0_), .B(
        npu_inst_pe_1_4_7_n13), .ZN(npu_inst_pe_1_4_7_N65) );
  OR2_X1 npu_inst_pe_1_4_7_U139 ( .A1(npu_inst_pe_1_4_7_n13), .A2(
        npu_inst_pe_1_4_7_int_q_acc_0_), .ZN(npu_inst_pe_1_4_7_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_4_7_U138 ( .A(npu_inst_pe_1_4_7_int_q_acc_2_), .B(
        npu_inst_pe_1_4_7_add_69_carry_2_), .Z(npu_inst_pe_1_4_7_N75) );
  AND2_X1 npu_inst_pe_1_4_7_U137 ( .A1(npu_inst_pe_1_4_7_add_69_carry_2_), 
        .A2(npu_inst_pe_1_4_7_int_q_acc_2_), .ZN(
        npu_inst_pe_1_4_7_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_4_7_U136 ( .A(npu_inst_pe_1_4_7_int_q_acc_3_), .B(
        npu_inst_pe_1_4_7_add_69_carry_3_), .Z(npu_inst_pe_1_4_7_N76) );
  AND2_X1 npu_inst_pe_1_4_7_U135 ( .A1(npu_inst_pe_1_4_7_add_69_carry_3_), 
        .A2(npu_inst_pe_1_4_7_int_q_acc_3_), .ZN(
        npu_inst_pe_1_4_7_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_4_7_U134 ( .A(npu_inst_pe_1_4_7_int_q_acc_4_), .B(
        npu_inst_pe_1_4_7_add_69_carry_4_), .Z(npu_inst_pe_1_4_7_N77) );
  AND2_X1 npu_inst_pe_1_4_7_U133 ( .A1(npu_inst_pe_1_4_7_add_69_carry_4_), 
        .A2(npu_inst_pe_1_4_7_int_q_acc_4_), .ZN(
        npu_inst_pe_1_4_7_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_4_7_U132 ( .A(npu_inst_pe_1_4_7_int_q_acc_5_), .B(
        npu_inst_pe_1_4_7_add_69_carry_5_), .Z(npu_inst_pe_1_4_7_N78) );
  AND2_X1 npu_inst_pe_1_4_7_U131 ( .A1(npu_inst_pe_1_4_7_add_69_carry_5_), 
        .A2(npu_inst_pe_1_4_7_int_q_acc_5_), .ZN(
        npu_inst_pe_1_4_7_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_4_7_U130 ( .A(npu_inst_pe_1_4_7_int_q_acc_6_), .B(
        npu_inst_pe_1_4_7_add_69_carry_6_), .Z(npu_inst_pe_1_4_7_N79) );
  AND2_X1 npu_inst_pe_1_4_7_U129 ( .A1(npu_inst_pe_1_4_7_add_69_carry_6_), 
        .A2(npu_inst_pe_1_4_7_int_q_acc_6_), .ZN(
        npu_inst_pe_1_4_7_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_4_7_U128 ( .A(npu_inst_pe_1_4_7_int_q_acc_7_), .B(
        npu_inst_pe_1_4_7_add_69_carry_7_), .Z(npu_inst_pe_1_4_7_N80) );
  XNOR2_X1 npu_inst_pe_1_4_7_U127 ( .A(npu_inst_pe_1_4_7_sub_67_carry_2_), .B(
        npu_inst_pe_1_4_7_int_q_acc_2_), .ZN(npu_inst_pe_1_4_7_N67) );
  OR2_X1 npu_inst_pe_1_4_7_U126 ( .A1(npu_inst_pe_1_4_7_int_q_acc_2_), .A2(
        npu_inst_pe_1_4_7_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_4_7_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_4_7_U125 ( .A(npu_inst_pe_1_4_7_sub_67_carry_3_), .B(
        npu_inst_pe_1_4_7_int_q_acc_3_), .ZN(npu_inst_pe_1_4_7_N68) );
  OR2_X1 npu_inst_pe_1_4_7_U124 ( .A1(npu_inst_pe_1_4_7_int_q_acc_3_), .A2(
        npu_inst_pe_1_4_7_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_4_7_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_4_7_U123 ( .A(npu_inst_pe_1_4_7_sub_67_carry_4_), .B(
        npu_inst_pe_1_4_7_int_q_acc_4_), .ZN(npu_inst_pe_1_4_7_N69) );
  OR2_X1 npu_inst_pe_1_4_7_U122 ( .A1(npu_inst_pe_1_4_7_int_q_acc_4_), .A2(
        npu_inst_pe_1_4_7_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_4_7_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_4_7_U121 ( .A(npu_inst_pe_1_4_7_sub_67_carry_5_), .B(
        npu_inst_pe_1_4_7_int_q_acc_5_), .ZN(npu_inst_pe_1_4_7_N70) );
  OR2_X1 npu_inst_pe_1_4_7_U120 ( .A1(npu_inst_pe_1_4_7_int_q_acc_5_), .A2(
        npu_inst_pe_1_4_7_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_4_7_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_4_7_U119 ( .A(npu_inst_pe_1_4_7_sub_67_carry_6_), .B(
        npu_inst_pe_1_4_7_int_q_acc_6_), .ZN(npu_inst_pe_1_4_7_N71) );
  OR2_X1 npu_inst_pe_1_4_7_U118 ( .A1(npu_inst_pe_1_4_7_int_q_acc_6_), .A2(
        npu_inst_pe_1_4_7_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_4_7_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_4_7_U117 ( .A(npu_inst_pe_1_4_7_int_q_acc_7_), .B(
        npu_inst_pe_1_4_7_sub_67_carry_7_), .ZN(npu_inst_pe_1_4_7_N72) );
  INV_X1 npu_inst_pe_1_4_7_U116 ( .A(npu_inst_n77), .ZN(npu_inst_pe_1_4_7_n7)
         );
  INV_X1 npu_inst_pe_1_4_7_U115 ( .A(npu_inst_pe_1_4_7_n7), .ZN(
        npu_inst_pe_1_4_7_n6) );
  INV_X1 npu_inst_pe_1_4_7_U114 ( .A(npu_inst_n55), .ZN(npu_inst_pe_1_4_7_n3)
         );
  AOI22_X1 npu_inst_pe_1_4_7_U113 ( .A1(npu_inst_int_data_y_5__7__0_), .A2(
        npu_inst_pe_1_4_7_n58), .B1(npu_inst_pe_1_4_7_n119), .B2(
        npu_inst_pe_1_4_7_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_4_7_n57) );
  INV_X1 npu_inst_pe_1_4_7_U112 ( .A(npu_inst_pe_1_4_7_n57), .ZN(
        npu_inst_pe_1_4_7_n108) );
  AOI22_X1 npu_inst_pe_1_4_7_U111 ( .A1(npu_inst_int_data_y_5__7__0_), .A2(
        npu_inst_pe_1_4_7_n54), .B1(npu_inst_pe_1_4_7_n118), .B2(
        npu_inst_pe_1_4_7_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_4_7_n53) );
  INV_X1 npu_inst_pe_1_4_7_U110 ( .A(npu_inst_pe_1_4_7_n53), .ZN(
        npu_inst_pe_1_4_7_n109) );
  AOI22_X1 npu_inst_pe_1_4_7_U107 ( .A1(npu_inst_int_data_y_5__7__0_), .A2(
        npu_inst_pe_1_4_7_n50), .B1(npu_inst_pe_1_4_7_n117), .B2(
        npu_inst_pe_1_4_7_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_4_7_n49) );
  INV_X1 npu_inst_pe_1_4_7_U106 ( .A(npu_inst_pe_1_4_7_n49), .ZN(
        npu_inst_pe_1_4_7_n110) );
  AOI22_X1 npu_inst_pe_1_4_7_U105 ( .A1(npu_inst_int_data_y_5__7__0_), .A2(
        npu_inst_pe_1_4_7_n46), .B1(npu_inst_pe_1_4_7_n116), .B2(
        npu_inst_pe_1_4_7_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_4_7_n45) );
  INV_X1 npu_inst_pe_1_4_7_U104 ( .A(npu_inst_pe_1_4_7_n45), .ZN(
        npu_inst_pe_1_4_7_n111) );
  AOI22_X1 npu_inst_pe_1_4_7_U103 ( .A1(npu_inst_int_data_y_5__7__0_), .A2(
        npu_inst_pe_1_4_7_n42), .B1(npu_inst_pe_1_4_7_n115), .B2(
        npu_inst_pe_1_4_7_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_4_7_n41) );
  INV_X1 npu_inst_pe_1_4_7_U102 ( .A(npu_inst_pe_1_4_7_n41), .ZN(
        npu_inst_pe_1_4_7_n112) );
  AOI22_X1 npu_inst_pe_1_4_7_U101 ( .A1(npu_inst_int_data_y_5__7__1_), .A2(
        npu_inst_pe_1_4_7_n58), .B1(npu_inst_pe_1_4_7_n119), .B2(
        npu_inst_pe_1_4_7_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_4_7_n59) );
  INV_X1 npu_inst_pe_1_4_7_U100 ( .A(npu_inst_pe_1_4_7_n59), .ZN(
        npu_inst_pe_1_4_7_n102) );
  AOI22_X1 npu_inst_pe_1_4_7_U99 ( .A1(npu_inst_int_data_y_5__7__1_), .A2(
        npu_inst_pe_1_4_7_n54), .B1(npu_inst_pe_1_4_7_n118), .B2(
        npu_inst_pe_1_4_7_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_4_7_n55) );
  INV_X1 npu_inst_pe_1_4_7_U98 ( .A(npu_inst_pe_1_4_7_n55), .ZN(
        npu_inst_pe_1_4_7_n103) );
  AOI22_X1 npu_inst_pe_1_4_7_U97 ( .A1(npu_inst_int_data_y_5__7__1_), .A2(
        npu_inst_pe_1_4_7_n50), .B1(npu_inst_pe_1_4_7_n117), .B2(
        npu_inst_pe_1_4_7_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_4_7_n51) );
  INV_X1 npu_inst_pe_1_4_7_U96 ( .A(npu_inst_pe_1_4_7_n51), .ZN(
        npu_inst_pe_1_4_7_n104) );
  AOI22_X1 npu_inst_pe_1_4_7_U95 ( .A1(npu_inst_int_data_y_5__7__1_), .A2(
        npu_inst_pe_1_4_7_n46), .B1(npu_inst_pe_1_4_7_n116), .B2(
        npu_inst_pe_1_4_7_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_4_7_n47) );
  INV_X1 npu_inst_pe_1_4_7_U94 ( .A(npu_inst_pe_1_4_7_n47), .ZN(
        npu_inst_pe_1_4_7_n105) );
  AOI22_X1 npu_inst_pe_1_4_7_U93 ( .A1(npu_inst_int_data_y_5__7__1_), .A2(
        npu_inst_pe_1_4_7_n42), .B1(npu_inst_pe_1_4_7_n115), .B2(
        npu_inst_pe_1_4_7_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_4_7_n43) );
  INV_X1 npu_inst_pe_1_4_7_U92 ( .A(npu_inst_pe_1_4_7_n43), .ZN(
        npu_inst_pe_1_4_7_n106) );
  AOI22_X1 npu_inst_pe_1_4_7_U91 ( .A1(npu_inst_pe_1_4_7_n38), .A2(
        npu_inst_int_data_y_5__7__1_), .B1(npu_inst_pe_1_4_7_n114), .B2(
        npu_inst_pe_1_4_7_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_4_7_n39) );
  INV_X1 npu_inst_pe_1_4_7_U90 ( .A(npu_inst_pe_1_4_7_n39), .ZN(
        npu_inst_pe_1_4_7_n107) );
  AOI22_X1 npu_inst_pe_1_4_7_U89 ( .A1(npu_inst_pe_1_4_7_n38), .A2(
        npu_inst_int_data_y_5__7__0_), .B1(npu_inst_pe_1_4_7_n114), .B2(
        npu_inst_pe_1_4_7_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_4_7_n37) );
  INV_X1 npu_inst_pe_1_4_7_U88 ( .A(npu_inst_pe_1_4_7_n37), .ZN(
        npu_inst_pe_1_4_7_n113) );
  AND2_X1 npu_inst_pe_1_4_7_U87 ( .A1(npu_inst_pe_1_4_7_N93), .A2(npu_inst_n55), .ZN(npu_inst_int_data_y_4__7__0_) );
  AND2_X1 npu_inst_pe_1_4_7_U86 ( .A1(npu_inst_n55), .A2(npu_inst_pe_1_4_7_N94), .ZN(npu_inst_int_data_y_4__7__1_) );
  NOR3_X1 npu_inst_pe_1_4_7_U85 ( .A1(npu_inst_pe_1_4_7_n26), .A2(npu_inst_n55), .A3(npu_inst_int_ckg[24]), .ZN(npu_inst_pe_1_4_7_n85) );
  OR2_X1 npu_inst_pe_1_4_7_U84 ( .A1(npu_inst_pe_1_4_7_n85), .A2(
        npu_inst_pe_1_4_7_n2), .ZN(npu_inst_pe_1_4_7_N84) );
  AND2_X1 npu_inst_pe_1_4_7_U83 ( .A1(npu_inst_pe_1_4_7_int_q_acc_0_), .A2(
        npu_inst_pe_1_4_7_n1), .ZN(npu_inst_int_data_res_4__7__0_) );
  AND2_X1 npu_inst_pe_1_4_7_U82 ( .A1(npu_inst_pe_1_4_7_n2), .A2(
        npu_inst_pe_1_4_7_int_q_acc_7_), .ZN(npu_inst_int_data_res_4__7__7_)
         );
  AND2_X1 npu_inst_pe_1_4_7_U81 ( .A1(npu_inst_pe_1_4_7_int_q_acc_1_), .A2(
        npu_inst_pe_1_4_7_n1), .ZN(npu_inst_int_data_res_4__7__1_) );
  AND2_X1 npu_inst_pe_1_4_7_U80 ( .A1(npu_inst_pe_1_4_7_int_q_acc_2_), .A2(
        npu_inst_pe_1_4_7_n1), .ZN(npu_inst_int_data_res_4__7__2_) );
  AND2_X1 npu_inst_pe_1_4_7_U79 ( .A1(npu_inst_pe_1_4_7_int_q_acc_3_), .A2(
        npu_inst_pe_1_4_7_n2), .ZN(npu_inst_int_data_res_4__7__3_) );
  AND2_X1 npu_inst_pe_1_4_7_U78 ( .A1(npu_inst_pe_1_4_7_int_q_acc_4_), .A2(
        npu_inst_pe_1_4_7_n2), .ZN(npu_inst_int_data_res_4__7__4_) );
  AND2_X1 npu_inst_pe_1_4_7_U77 ( .A1(npu_inst_pe_1_4_7_int_q_acc_5_), .A2(
        npu_inst_pe_1_4_7_n2), .ZN(npu_inst_int_data_res_4__7__5_) );
  AND2_X1 npu_inst_pe_1_4_7_U76 ( .A1(npu_inst_pe_1_4_7_int_q_acc_6_), .A2(
        npu_inst_pe_1_4_7_n2), .ZN(npu_inst_int_data_res_4__7__6_) );
  AOI222_X1 npu_inst_pe_1_4_7_U75 ( .A1(npu_inst_int_data_res_5__7__0_), .A2(
        npu_inst_pe_1_4_7_n1), .B1(npu_inst_pe_1_4_7_N73), .B2(
        npu_inst_pe_1_4_7_n76), .C1(npu_inst_pe_1_4_7_N65), .C2(
        npu_inst_pe_1_4_7_n77), .ZN(npu_inst_pe_1_4_7_n84) );
  INV_X1 npu_inst_pe_1_4_7_U74 ( .A(npu_inst_pe_1_4_7_n84), .ZN(
        npu_inst_pe_1_4_7_n101) );
  AOI222_X1 npu_inst_pe_1_4_7_U73 ( .A1(npu_inst_int_data_res_5__7__7_), .A2(
        npu_inst_pe_1_4_7_n1), .B1(npu_inst_pe_1_4_7_N80), .B2(
        npu_inst_pe_1_4_7_n76), .C1(npu_inst_pe_1_4_7_N72), .C2(
        npu_inst_pe_1_4_7_n77), .ZN(npu_inst_pe_1_4_7_n75) );
  INV_X1 npu_inst_pe_1_4_7_U72 ( .A(npu_inst_pe_1_4_7_n75), .ZN(
        npu_inst_pe_1_4_7_n33) );
  AOI222_X1 npu_inst_pe_1_4_7_U71 ( .A1(npu_inst_int_data_res_5__7__1_), .A2(
        npu_inst_pe_1_4_7_n1), .B1(npu_inst_pe_1_4_7_N74), .B2(
        npu_inst_pe_1_4_7_n76), .C1(npu_inst_pe_1_4_7_N66), .C2(
        npu_inst_pe_1_4_7_n77), .ZN(npu_inst_pe_1_4_7_n83) );
  INV_X1 npu_inst_pe_1_4_7_U70 ( .A(npu_inst_pe_1_4_7_n83), .ZN(
        npu_inst_pe_1_4_7_n100) );
  AOI222_X1 npu_inst_pe_1_4_7_U69 ( .A1(npu_inst_int_data_res_5__7__2_), .A2(
        npu_inst_pe_1_4_7_n1), .B1(npu_inst_pe_1_4_7_N75), .B2(
        npu_inst_pe_1_4_7_n76), .C1(npu_inst_pe_1_4_7_N67), .C2(
        npu_inst_pe_1_4_7_n77), .ZN(npu_inst_pe_1_4_7_n82) );
  INV_X1 npu_inst_pe_1_4_7_U68 ( .A(npu_inst_pe_1_4_7_n82), .ZN(
        npu_inst_pe_1_4_7_n99) );
  AOI222_X1 npu_inst_pe_1_4_7_U67 ( .A1(npu_inst_int_data_res_5__7__3_), .A2(
        npu_inst_pe_1_4_7_n1), .B1(npu_inst_pe_1_4_7_N76), .B2(
        npu_inst_pe_1_4_7_n76), .C1(npu_inst_pe_1_4_7_N68), .C2(
        npu_inst_pe_1_4_7_n77), .ZN(npu_inst_pe_1_4_7_n81) );
  INV_X1 npu_inst_pe_1_4_7_U66 ( .A(npu_inst_pe_1_4_7_n81), .ZN(
        npu_inst_pe_1_4_7_n98) );
  AOI222_X1 npu_inst_pe_1_4_7_U65 ( .A1(npu_inst_int_data_res_5__7__4_), .A2(
        npu_inst_pe_1_4_7_n1), .B1(npu_inst_pe_1_4_7_N77), .B2(
        npu_inst_pe_1_4_7_n76), .C1(npu_inst_pe_1_4_7_N69), .C2(
        npu_inst_pe_1_4_7_n77), .ZN(npu_inst_pe_1_4_7_n80) );
  INV_X1 npu_inst_pe_1_4_7_U64 ( .A(npu_inst_pe_1_4_7_n80), .ZN(
        npu_inst_pe_1_4_7_n36) );
  AOI222_X1 npu_inst_pe_1_4_7_U63 ( .A1(npu_inst_int_data_res_5__7__5_), .A2(
        npu_inst_pe_1_4_7_n1), .B1(npu_inst_pe_1_4_7_N78), .B2(
        npu_inst_pe_1_4_7_n76), .C1(npu_inst_pe_1_4_7_N70), .C2(
        npu_inst_pe_1_4_7_n77), .ZN(npu_inst_pe_1_4_7_n79) );
  INV_X1 npu_inst_pe_1_4_7_U62 ( .A(npu_inst_pe_1_4_7_n79), .ZN(
        npu_inst_pe_1_4_7_n35) );
  AOI222_X1 npu_inst_pe_1_4_7_U61 ( .A1(npu_inst_int_data_res_5__7__6_), .A2(
        npu_inst_pe_1_4_7_n1), .B1(npu_inst_pe_1_4_7_N79), .B2(
        npu_inst_pe_1_4_7_n76), .C1(npu_inst_pe_1_4_7_N71), .C2(
        npu_inst_pe_1_4_7_n77), .ZN(npu_inst_pe_1_4_7_n78) );
  INV_X1 npu_inst_pe_1_4_7_U60 ( .A(npu_inst_pe_1_4_7_n78), .ZN(
        npu_inst_pe_1_4_7_n34) );
  INV_X1 npu_inst_pe_1_4_7_U59 ( .A(npu_inst_pe_1_4_7_int_data_1_), .ZN(
        npu_inst_pe_1_4_7_n14) );
  AND2_X1 npu_inst_pe_1_4_7_U58 ( .A1(npu_inst_int_data_x_4__7__1_), .A2(
        npu_inst_pe_1_4_7_int_q_weight_1_), .ZN(npu_inst_pe_1_4_7_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_4_7_U57 ( .A1(npu_inst_int_data_x_4__7__0_), .A2(
        npu_inst_pe_1_4_7_int_q_weight_1_), .ZN(npu_inst_pe_1_4_7_int_data_0_)
         );
  NAND2_X1 npu_inst_pe_1_4_7_U56 ( .A1(npu_inst_pe_1_4_7_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_4_7_n60), .ZN(npu_inst_pe_1_4_7_n74) );
  OAI21_X1 npu_inst_pe_1_4_7_U55 ( .B1(npu_inst_pe_1_4_7_n63), .B2(
        npu_inst_pe_1_4_7_n60), .A(npu_inst_pe_1_4_7_n74), .ZN(
        npu_inst_pe_1_4_7_n97) );
  NAND2_X1 npu_inst_pe_1_4_7_U54 ( .A1(npu_inst_pe_1_4_7_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_4_7_n60), .ZN(npu_inst_pe_1_4_7_n73) );
  OAI21_X1 npu_inst_pe_1_4_7_U53 ( .B1(npu_inst_pe_1_4_7_n61), .B2(
        npu_inst_pe_1_4_7_n60), .A(npu_inst_pe_1_4_7_n73), .ZN(
        npu_inst_pe_1_4_7_n96) );
  NAND2_X1 npu_inst_pe_1_4_7_U52 ( .A1(npu_inst_pe_1_4_7_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_4_7_n56), .ZN(npu_inst_pe_1_4_7_n72) );
  OAI21_X1 npu_inst_pe_1_4_7_U51 ( .B1(npu_inst_pe_1_4_7_n63), .B2(
        npu_inst_pe_1_4_7_n56), .A(npu_inst_pe_1_4_7_n72), .ZN(
        npu_inst_pe_1_4_7_n95) );
  NAND2_X1 npu_inst_pe_1_4_7_U50 ( .A1(npu_inst_pe_1_4_7_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_4_7_n56), .ZN(npu_inst_pe_1_4_7_n71) );
  OAI21_X1 npu_inst_pe_1_4_7_U49 ( .B1(npu_inst_pe_1_4_7_n61), .B2(
        npu_inst_pe_1_4_7_n56), .A(npu_inst_pe_1_4_7_n71), .ZN(
        npu_inst_pe_1_4_7_n94) );
  NAND2_X1 npu_inst_pe_1_4_7_U48 ( .A1(npu_inst_pe_1_4_7_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_4_7_n52), .ZN(npu_inst_pe_1_4_7_n70) );
  OAI21_X1 npu_inst_pe_1_4_7_U47 ( .B1(npu_inst_pe_1_4_7_n63), .B2(
        npu_inst_pe_1_4_7_n52), .A(npu_inst_pe_1_4_7_n70), .ZN(
        npu_inst_pe_1_4_7_n93) );
  NAND2_X1 npu_inst_pe_1_4_7_U46 ( .A1(npu_inst_pe_1_4_7_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_4_7_n52), .ZN(npu_inst_pe_1_4_7_n69) );
  OAI21_X1 npu_inst_pe_1_4_7_U45 ( .B1(npu_inst_pe_1_4_7_n61), .B2(
        npu_inst_pe_1_4_7_n52), .A(npu_inst_pe_1_4_7_n69), .ZN(
        npu_inst_pe_1_4_7_n92) );
  NAND2_X1 npu_inst_pe_1_4_7_U44 ( .A1(npu_inst_pe_1_4_7_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_4_7_n48), .ZN(npu_inst_pe_1_4_7_n68) );
  OAI21_X1 npu_inst_pe_1_4_7_U43 ( .B1(npu_inst_pe_1_4_7_n63), .B2(
        npu_inst_pe_1_4_7_n48), .A(npu_inst_pe_1_4_7_n68), .ZN(
        npu_inst_pe_1_4_7_n91) );
  NAND2_X1 npu_inst_pe_1_4_7_U42 ( .A1(npu_inst_pe_1_4_7_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_4_7_n48), .ZN(npu_inst_pe_1_4_7_n67) );
  OAI21_X1 npu_inst_pe_1_4_7_U41 ( .B1(npu_inst_pe_1_4_7_n61), .B2(
        npu_inst_pe_1_4_7_n48), .A(npu_inst_pe_1_4_7_n67), .ZN(
        npu_inst_pe_1_4_7_n90) );
  NAND2_X1 npu_inst_pe_1_4_7_U40 ( .A1(npu_inst_pe_1_4_7_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_4_7_n44), .ZN(npu_inst_pe_1_4_7_n66) );
  OAI21_X1 npu_inst_pe_1_4_7_U39 ( .B1(npu_inst_pe_1_4_7_n63), .B2(
        npu_inst_pe_1_4_7_n44), .A(npu_inst_pe_1_4_7_n66), .ZN(
        npu_inst_pe_1_4_7_n89) );
  NAND2_X1 npu_inst_pe_1_4_7_U38 ( .A1(npu_inst_pe_1_4_7_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_4_7_n44), .ZN(npu_inst_pe_1_4_7_n65) );
  OAI21_X1 npu_inst_pe_1_4_7_U37 ( .B1(npu_inst_pe_1_4_7_n61), .B2(
        npu_inst_pe_1_4_7_n44), .A(npu_inst_pe_1_4_7_n65), .ZN(
        npu_inst_pe_1_4_7_n88) );
  NAND2_X1 npu_inst_pe_1_4_7_U36 ( .A1(npu_inst_pe_1_4_7_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_4_7_n40), .ZN(npu_inst_pe_1_4_7_n64) );
  OAI21_X1 npu_inst_pe_1_4_7_U35 ( .B1(npu_inst_pe_1_4_7_n63), .B2(
        npu_inst_pe_1_4_7_n40), .A(npu_inst_pe_1_4_7_n64), .ZN(
        npu_inst_pe_1_4_7_n87) );
  NAND2_X1 npu_inst_pe_1_4_7_U34 ( .A1(npu_inst_pe_1_4_7_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_4_7_n40), .ZN(npu_inst_pe_1_4_7_n62) );
  OAI21_X1 npu_inst_pe_1_4_7_U33 ( .B1(npu_inst_pe_1_4_7_n61), .B2(
        npu_inst_pe_1_4_7_n40), .A(npu_inst_pe_1_4_7_n62), .ZN(
        npu_inst_pe_1_4_7_n86) );
  INV_X1 npu_inst_pe_1_4_7_U32 ( .A(npu_inst_pe_1_4_7_int_data_0_), .ZN(
        npu_inst_pe_1_4_7_n13) );
  INV_X1 npu_inst_pe_1_4_7_U31 ( .A(npu_inst_n69), .ZN(npu_inst_pe_1_4_7_n5)
         );
  AOI22_X1 npu_inst_pe_1_4_7_U30 ( .A1(npu_inst_n55), .A2(
        npu_inst_int_data_y_5__7__1_), .B1(npu_inst_pe_1_4_7_n3), .B2(
        int_i_data_h_npu[7]), .ZN(npu_inst_pe_1_4_7_n63) );
  AOI22_X1 npu_inst_pe_1_4_7_U29 ( .A1(npu_inst_n55), .A2(
        npu_inst_int_data_y_5__7__0_), .B1(npu_inst_pe_1_4_7_n3), .B2(
        int_i_data_h_npu[6]), .ZN(npu_inst_pe_1_4_7_n61) );
  OR3_X1 npu_inst_pe_1_4_7_U28 ( .A1(npu_inst_pe_1_4_7_n6), .A2(
        npu_inst_pe_1_4_7_n8), .A3(npu_inst_pe_1_4_7_n5), .ZN(
        npu_inst_pe_1_4_7_n56) );
  OR3_X1 npu_inst_pe_1_4_7_U27 ( .A1(npu_inst_pe_1_4_7_n5), .A2(
        npu_inst_pe_1_4_7_n8), .A3(npu_inst_pe_1_4_7_n7), .ZN(
        npu_inst_pe_1_4_7_n48) );
  INV_X1 npu_inst_pe_1_4_7_U26 ( .A(npu_inst_pe_1_4_7_n5), .ZN(
        npu_inst_pe_1_4_7_n4) );
  OR3_X1 npu_inst_pe_1_4_7_U25 ( .A1(npu_inst_pe_1_4_7_n4), .A2(
        npu_inst_pe_1_4_7_n8), .A3(npu_inst_pe_1_4_7_n7), .ZN(
        npu_inst_pe_1_4_7_n52) );
  OR3_X1 npu_inst_pe_1_4_7_U24 ( .A1(npu_inst_pe_1_4_7_n6), .A2(
        npu_inst_pe_1_4_7_n8), .A3(npu_inst_pe_1_4_7_n4), .ZN(
        npu_inst_pe_1_4_7_n60) );
  NOR2_X1 npu_inst_pe_1_4_7_U23 ( .A1(npu_inst_pe_1_4_7_n60), .A2(
        npu_inst_pe_1_4_7_n3), .ZN(npu_inst_pe_1_4_7_n58) );
  NOR2_X1 npu_inst_pe_1_4_7_U22 ( .A1(npu_inst_pe_1_4_7_n56), .A2(
        npu_inst_pe_1_4_7_n3), .ZN(npu_inst_pe_1_4_7_n54) );
  NOR2_X1 npu_inst_pe_1_4_7_U21 ( .A1(npu_inst_pe_1_4_7_n52), .A2(
        npu_inst_pe_1_4_7_n3), .ZN(npu_inst_pe_1_4_7_n50) );
  NOR2_X1 npu_inst_pe_1_4_7_U20 ( .A1(npu_inst_pe_1_4_7_n48), .A2(
        npu_inst_pe_1_4_7_n3), .ZN(npu_inst_pe_1_4_7_n46) );
  NOR2_X1 npu_inst_pe_1_4_7_U19 ( .A1(npu_inst_pe_1_4_7_n40), .A2(
        npu_inst_pe_1_4_7_n3), .ZN(npu_inst_pe_1_4_7_n38) );
  NOR2_X1 npu_inst_pe_1_4_7_U18 ( .A1(npu_inst_pe_1_4_7_n44), .A2(
        npu_inst_pe_1_4_7_n3), .ZN(npu_inst_pe_1_4_7_n42) );
  BUF_X1 npu_inst_pe_1_4_7_U17 ( .A(npu_inst_n98), .Z(npu_inst_pe_1_4_7_n8) );
  INV_X1 npu_inst_pe_1_4_7_U16 ( .A(npu_inst_n124), .ZN(npu_inst_pe_1_4_7_n12)
         );
  INV_X1 npu_inst_pe_1_4_7_U15 ( .A(npu_inst_pe_1_4_7_n38), .ZN(
        npu_inst_pe_1_4_7_n114) );
  INV_X1 npu_inst_pe_1_4_7_U14 ( .A(npu_inst_pe_1_4_7_n58), .ZN(
        npu_inst_pe_1_4_7_n119) );
  INV_X1 npu_inst_pe_1_4_7_U13 ( .A(npu_inst_pe_1_4_7_n54), .ZN(
        npu_inst_pe_1_4_7_n118) );
  INV_X1 npu_inst_pe_1_4_7_U12 ( .A(npu_inst_pe_1_4_7_n50), .ZN(
        npu_inst_pe_1_4_7_n117) );
  INV_X1 npu_inst_pe_1_4_7_U11 ( .A(npu_inst_pe_1_4_7_n46), .ZN(
        npu_inst_pe_1_4_7_n116) );
  INV_X1 npu_inst_pe_1_4_7_U10 ( .A(npu_inst_pe_1_4_7_n42), .ZN(
        npu_inst_pe_1_4_7_n115) );
  BUF_X1 npu_inst_pe_1_4_7_U9 ( .A(npu_inst_n19), .Z(npu_inst_pe_1_4_7_n2) );
  BUF_X1 npu_inst_pe_1_4_7_U8 ( .A(npu_inst_n19), .Z(npu_inst_pe_1_4_7_n1) );
  BUF_X1 npu_inst_pe_1_4_7_U7 ( .A(npu_inst_pe_1_4_7_n12), .Z(
        npu_inst_pe_1_4_7_n11) );
  BUF_X1 npu_inst_pe_1_4_7_U6 ( .A(npu_inst_pe_1_4_7_n12), .Z(
        npu_inst_pe_1_4_7_n10) );
  BUF_X1 npu_inst_pe_1_4_7_U5 ( .A(npu_inst_pe_1_4_7_n12), .Z(
        npu_inst_pe_1_4_7_n9) );
  NOR2_X1 npu_inst_pe_1_4_7_U4 ( .A1(npu_inst_pe_1_4_7_int_q_weight_0_), .A2(
        npu_inst_pe_1_4_7_n1), .ZN(npu_inst_pe_1_4_7_n76) );
  NOR2_X1 npu_inst_pe_1_4_7_U3 ( .A1(npu_inst_pe_1_4_7_n27), .A2(
        npu_inst_pe_1_4_7_n1), .ZN(npu_inst_pe_1_4_7_n77) );
  FA_X1 npu_inst_pe_1_4_7_sub_67_U2_1 ( .A(npu_inst_pe_1_4_7_int_q_acc_1_), 
        .B(npu_inst_pe_1_4_7_n14), .CI(npu_inst_pe_1_4_7_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_4_7_sub_67_carry_2_), .S(npu_inst_pe_1_4_7_N66) );
  FA_X1 npu_inst_pe_1_4_7_add_69_U1_1 ( .A(npu_inst_pe_1_4_7_int_q_acc_1_), 
        .B(npu_inst_pe_1_4_7_int_data_1_), .CI(
        npu_inst_pe_1_4_7_add_69_carry_1_), .CO(
        npu_inst_pe_1_4_7_add_69_carry_2_), .S(npu_inst_pe_1_4_7_N74) );
  NAND3_X1 npu_inst_pe_1_4_7_U109 ( .A1(npu_inst_pe_1_4_7_n5), .A2(
        npu_inst_pe_1_4_7_n7), .A3(npu_inst_pe_1_4_7_n8), .ZN(
        npu_inst_pe_1_4_7_n44) );
  NAND3_X1 npu_inst_pe_1_4_7_U108 ( .A1(npu_inst_pe_1_4_7_n4), .A2(
        npu_inst_pe_1_4_7_n7), .A3(npu_inst_pe_1_4_7_n8), .ZN(
        npu_inst_pe_1_4_7_n40) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_4_7_n34), .CK(
        npu_inst_pe_1_4_7_net3665), .RN(npu_inst_pe_1_4_7_n9), .Q(
        npu_inst_pe_1_4_7_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_4_7_n35), .CK(
        npu_inst_pe_1_4_7_net3665), .RN(npu_inst_pe_1_4_7_n9), .Q(
        npu_inst_pe_1_4_7_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_4_7_n36), .CK(
        npu_inst_pe_1_4_7_net3665), .RN(npu_inst_pe_1_4_7_n9), .Q(
        npu_inst_pe_1_4_7_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_4_7_n98), .CK(
        npu_inst_pe_1_4_7_net3665), .RN(npu_inst_pe_1_4_7_n9), .Q(
        npu_inst_pe_1_4_7_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_4_7_n99), .CK(
        npu_inst_pe_1_4_7_net3665), .RN(npu_inst_pe_1_4_7_n9), .Q(
        npu_inst_pe_1_4_7_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_4_7_n100), 
        .CK(npu_inst_pe_1_4_7_net3665), .RN(npu_inst_pe_1_4_7_n9), .Q(
        npu_inst_pe_1_4_7_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_4_7_n33), .CK(
        npu_inst_pe_1_4_7_net3665), .RN(npu_inst_pe_1_4_7_n9), .Q(
        npu_inst_pe_1_4_7_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_4_7_n101), 
        .CK(npu_inst_pe_1_4_7_net3665), .RN(npu_inst_pe_1_4_7_n9), .Q(
        npu_inst_pe_1_4_7_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_weight_reg_0_ ( .D(npu_inst_n110), .CK(
        npu_inst_pe_1_4_7_net3671), .RN(npu_inst_pe_1_4_7_n9), .Q(
        npu_inst_pe_1_4_7_int_q_weight_0_), .QN(npu_inst_pe_1_4_7_n27) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_weight_reg_1_ ( .D(npu_inst_n116), .CK(
        npu_inst_pe_1_4_7_net3671), .RN(npu_inst_pe_1_4_7_n9), .Q(
        npu_inst_pe_1_4_7_int_q_weight_1_), .QN(npu_inst_pe_1_4_7_n26) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_4_7_n113), 
        .CK(npu_inst_pe_1_4_7_net3671), .RN(npu_inst_pe_1_4_7_n9), .Q(
        npu_inst_pe_1_4_7_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_4_7_n107), 
        .CK(npu_inst_pe_1_4_7_net3671), .RN(npu_inst_pe_1_4_7_n9), .Q(
        npu_inst_pe_1_4_7_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_4_7_n112), 
        .CK(npu_inst_pe_1_4_7_net3671), .RN(npu_inst_pe_1_4_7_n10), .Q(
        npu_inst_pe_1_4_7_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_4_7_n106), 
        .CK(npu_inst_pe_1_4_7_net3671), .RN(npu_inst_pe_1_4_7_n10), .Q(
        npu_inst_pe_1_4_7_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_4_7_n111), 
        .CK(npu_inst_pe_1_4_7_net3671), .RN(npu_inst_pe_1_4_7_n10), .Q(
        npu_inst_pe_1_4_7_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_4_7_n105), 
        .CK(npu_inst_pe_1_4_7_net3671), .RN(npu_inst_pe_1_4_7_n10), .Q(
        npu_inst_pe_1_4_7_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_4_7_n110), 
        .CK(npu_inst_pe_1_4_7_net3671), .RN(npu_inst_pe_1_4_7_n10), .Q(
        npu_inst_pe_1_4_7_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_4_7_n104), 
        .CK(npu_inst_pe_1_4_7_net3671), .RN(npu_inst_pe_1_4_7_n10), .Q(
        npu_inst_pe_1_4_7_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_4_7_n109), 
        .CK(npu_inst_pe_1_4_7_net3671), .RN(npu_inst_pe_1_4_7_n10), .Q(
        npu_inst_pe_1_4_7_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_4_7_n103), 
        .CK(npu_inst_pe_1_4_7_net3671), .RN(npu_inst_pe_1_4_7_n10), .Q(
        npu_inst_pe_1_4_7_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_4_7_n108), 
        .CK(npu_inst_pe_1_4_7_net3671), .RN(npu_inst_pe_1_4_7_n10), .Q(
        npu_inst_pe_1_4_7_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_4_7_n102), 
        .CK(npu_inst_pe_1_4_7_net3671), .RN(npu_inst_pe_1_4_7_n10), .Q(
        npu_inst_pe_1_4_7_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_4_7_n86), 
        .CK(npu_inst_pe_1_4_7_net3671), .RN(npu_inst_pe_1_4_7_n10), .Q(
        npu_inst_pe_1_4_7_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_4_7_n87), 
        .CK(npu_inst_pe_1_4_7_net3671), .RN(npu_inst_pe_1_4_7_n10), .Q(
        npu_inst_pe_1_4_7_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_4_7_n88), 
        .CK(npu_inst_pe_1_4_7_net3671), .RN(npu_inst_pe_1_4_7_n11), .Q(
        npu_inst_pe_1_4_7_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_4_7_n89), 
        .CK(npu_inst_pe_1_4_7_net3671), .RN(npu_inst_pe_1_4_7_n11), .Q(
        npu_inst_pe_1_4_7_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_4_7_n90), 
        .CK(npu_inst_pe_1_4_7_net3671), .RN(npu_inst_pe_1_4_7_n11), .Q(
        npu_inst_pe_1_4_7_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_4_7_n91), 
        .CK(npu_inst_pe_1_4_7_net3671), .RN(npu_inst_pe_1_4_7_n11), .Q(
        npu_inst_pe_1_4_7_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_4_7_n92), 
        .CK(npu_inst_pe_1_4_7_net3671), .RN(npu_inst_pe_1_4_7_n11), .Q(
        npu_inst_pe_1_4_7_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_4_7_n93), 
        .CK(npu_inst_pe_1_4_7_net3671), .RN(npu_inst_pe_1_4_7_n11), .Q(
        npu_inst_pe_1_4_7_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_4_7_n94), 
        .CK(npu_inst_pe_1_4_7_net3671), .RN(npu_inst_pe_1_4_7_n11), .Q(
        npu_inst_pe_1_4_7_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_4_7_n95), 
        .CK(npu_inst_pe_1_4_7_net3671), .RN(npu_inst_pe_1_4_7_n11), .Q(
        npu_inst_pe_1_4_7_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_4_7_n96), 
        .CK(npu_inst_pe_1_4_7_net3671), .RN(npu_inst_pe_1_4_7_n11), .Q(
        npu_inst_pe_1_4_7_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_4_7_n97), 
        .CK(npu_inst_pe_1_4_7_net3671), .RN(npu_inst_pe_1_4_7_n11), .Q(
        npu_inst_pe_1_4_7_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_4_7_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_4_7_N84), .SE(1'b0), .GCK(npu_inst_pe_1_4_7_net3665) );
  CLKGATETST_X1 npu_inst_pe_1_4_7_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n63), .SE(1'b0), .GCK(npu_inst_pe_1_4_7_net3671) );
  MUX2_X1 npu_inst_pe_1_5_0_U161 ( .A(npu_inst_pe_1_5_0_n31), .B(
        npu_inst_pe_1_5_0_n28), .S(npu_inst_pe_1_5_0_n7), .Z(
        npu_inst_pe_1_5_0_N93) );
  MUX2_X1 npu_inst_pe_1_5_0_U160 ( .A(npu_inst_pe_1_5_0_n30), .B(
        npu_inst_pe_1_5_0_n29), .S(npu_inst_n76), .Z(npu_inst_pe_1_5_0_n31) );
  MUX2_X1 npu_inst_pe_1_5_0_U159 ( .A(npu_inst_pe_1_5_0_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_5_0_int_q_reg_v_1__0_), .S(npu_inst_pe_1_5_0_n4), .Z(
        npu_inst_pe_1_5_0_n30) );
  MUX2_X1 npu_inst_pe_1_5_0_U158 ( .A(npu_inst_pe_1_5_0_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_5_0_int_q_reg_v_3__0_), .S(npu_inst_pe_1_5_0_n4), .Z(
        npu_inst_pe_1_5_0_n29) );
  MUX2_X1 npu_inst_pe_1_5_0_U157 ( .A(npu_inst_pe_1_5_0_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_5_0_int_q_reg_v_5__0_), .S(npu_inst_pe_1_5_0_n4), .Z(
        npu_inst_pe_1_5_0_n28) );
  MUX2_X1 npu_inst_pe_1_5_0_U156 ( .A(npu_inst_pe_1_5_0_n25), .B(
        npu_inst_pe_1_5_0_n22), .S(npu_inst_pe_1_5_0_n7), .Z(
        npu_inst_pe_1_5_0_N94) );
  MUX2_X1 npu_inst_pe_1_5_0_U155 ( .A(npu_inst_pe_1_5_0_n24), .B(
        npu_inst_pe_1_5_0_n23), .S(npu_inst_n76), .Z(npu_inst_pe_1_5_0_n25) );
  MUX2_X1 npu_inst_pe_1_5_0_U154 ( .A(npu_inst_pe_1_5_0_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_5_0_int_q_reg_v_1__1_), .S(npu_inst_pe_1_5_0_n4), .Z(
        npu_inst_pe_1_5_0_n24) );
  MUX2_X1 npu_inst_pe_1_5_0_U153 ( .A(npu_inst_pe_1_5_0_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_5_0_int_q_reg_v_3__1_), .S(npu_inst_pe_1_5_0_n4), .Z(
        npu_inst_pe_1_5_0_n23) );
  MUX2_X1 npu_inst_pe_1_5_0_U152 ( .A(npu_inst_pe_1_5_0_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_5_0_int_q_reg_v_5__1_), .S(npu_inst_pe_1_5_0_n4), .Z(
        npu_inst_pe_1_5_0_n22) );
  MUX2_X1 npu_inst_pe_1_5_0_U151 ( .A(npu_inst_pe_1_5_0_n21), .B(
        npu_inst_pe_1_5_0_n18), .S(npu_inst_pe_1_5_0_n7), .Z(
        npu_inst_pe_1_5_0_o_data_h_1_) );
  MUX2_X1 npu_inst_pe_1_5_0_U150 ( .A(npu_inst_pe_1_5_0_n20), .B(
        npu_inst_pe_1_5_0_n19), .S(npu_inst_n76), .Z(npu_inst_pe_1_5_0_n21) );
  MUX2_X1 npu_inst_pe_1_5_0_U149 ( .A(npu_inst_pe_1_5_0_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_5_0_int_q_reg_h_1__1_), .S(npu_inst_pe_1_5_0_n4), .Z(
        npu_inst_pe_1_5_0_n20) );
  MUX2_X1 npu_inst_pe_1_5_0_U148 ( .A(npu_inst_pe_1_5_0_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_5_0_int_q_reg_h_3__1_), .S(npu_inst_pe_1_5_0_n4), .Z(
        npu_inst_pe_1_5_0_n19) );
  MUX2_X1 npu_inst_pe_1_5_0_U147 ( .A(npu_inst_pe_1_5_0_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_5_0_int_q_reg_h_5__1_), .S(npu_inst_pe_1_5_0_n4), .Z(
        npu_inst_pe_1_5_0_n18) );
  MUX2_X1 npu_inst_pe_1_5_0_U146 ( .A(npu_inst_pe_1_5_0_n17), .B(
        npu_inst_pe_1_5_0_n14), .S(npu_inst_pe_1_5_0_n7), .Z(
        npu_inst_pe_1_5_0_o_data_h_0_) );
  MUX2_X1 npu_inst_pe_1_5_0_U145 ( .A(npu_inst_pe_1_5_0_n16), .B(
        npu_inst_pe_1_5_0_n15), .S(npu_inst_n76), .Z(npu_inst_pe_1_5_0_n17) );
  MUX2_X1 npu_inst_pe_1_5_0_U144 ( .A(npu_inst_pe_1_5_0_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_5_0_int_q_reg_h_1__0_), .S(npu_inst_pe_1_5_0_n4), .Z(
        npu_inst_pe_1_5_0_n16) );
  MUX2_X1 npu_inst_pe_1_5_0_U143 ( .A(npu_inst_pe_1_5_0_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_5_0_int_q_reg_h_3__0_), .S(npu_inst_pe_1_5_0_n4), .Z(
        npu_inst_pe_1_5_0_n15) );
  MUX2_X1 npu_inst_pe_1_5_0_U142 ( .A(npu_inst_pe_1_5_0_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_5_0_int_q_reg_h_5__0_), .S(npu_inst_pe_1_5_0_n4), .Z(
        npu_inst_pe_1_5_0_n14) );
  XOR2_X1 npu_inst_pe_1_5_0_U141 ( .A(npu_inst_pe_1_5_0_int_data_0_), .B(
        npu_inst_pe_1_5_0_int_q_acc_0_), .Z(npu_inst_pe_1_5_0_N73) );
  AND2_X1 npu_inst_pe_1_5_0_U140 ( .A1(npu_inst_pe_1_5_0_int_q_acc_0_), .A2(
        npu_inst_pe_1_5_0_int_data_0_), .ZN(npu_inst_pe_1_5_0_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_5_0_U139 ( .A(npu_inst_pe_1_5_0_int_q_acc_0_), .B(
        npu_inst_pe_1_5_0_n12), .ZN(npu_inst_pe_1_5_0_N65) );
  OR2_X1 npu_inst_pe_1_5_0_U138 ( .A1(npu_inst_pe_1_5_0_n12), .A2(
        npu_inst_pe_1_5_0_int_q_acc_0_), .ZN(npu_inst_pe_1_5_0_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_5_0_U137 ( .A(npu_inst_pe_1_5_0_int_q_acc_2_), .B(
        npu_inst_pe_1_5_0_add_69_carry_2_), .Z(npu_inst_pe_1_5_0_N75) );
  AND2_X1 npu_inst_pe_1_5_0_U136 ( .A1(npu_inst_pe_1_5_0_add_69_carry_2_), 
        .A2(npu_inst_pe_1_5_0_int_q_acc_2_), .ZN(
        npu_inst_pe_1_5_0_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_5_0_U135 ( .A(npu_inst_pe_1_5_0_int_q_acc_3_), .B(
        npu_inst_pe_1_5_0_add_69_carry_3_), .Z(npu_inst_pe_1_5_0_N76) );
  AND2_X1 npu_inst_pe_1_5_0_U134 ( .A1(npu_inst_pe_1_5_0_add_69_carry_3_), 
        .A2(npu_inst_pe_1_5_0_int_q_acc_3_), .ZN(
        npu_inst_pe_1_5_0_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_5_0_U133 ( .A(npu_inst_pe_1_5_0_int_q_acc_4_), .B(
        npu_inst_pe_1_5_0_add_69_carry_4_), .Z(npu_inst_pe_1_5_0_N77) );
  AND2_X1 npu_inst_pe_1_5_0_U132 ( .A1(npu_inst_pe_1_5_0_add_69_carry_4_), 
        .A2(npu_inst_pe_1_5_0_int_q_acc_4_), .ZN(
        npu_inst_pe_1_5_0_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_5_0_U131 ( .A(npu_inst_pe_1_5_0_int_q_acc_5_), .B(
        npu_inst_pe_1_5_0_add_69_carry_5_), .Z(npu_inst_pe_1_5_0_N78) );
  AND2_X1 npu_inst_pe_1_5_0_U130 ( .A1(npu_inst_pe_1_5_0_add_69_carry_5_), 
        .A2(npu_inst_pe_1_5_0_int_q_acc_5_), .ZN(
        npu_inst_pe_1_5_0_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_5_0_U129 ( .A(npu_inst_pe_1_5_0_int_q_acc_6_), .B(
        npu_inst_pe_1_5_0_add_69_carry_6_), .Z(npu_inst_pe_1_5_0_N79) );
  AND2_X1 npu_inst_pe_1_5_0_U128 ( .A1(npu_inst_pe_1_5_0_add_69_carry_6_), 
        .A2(npu_inst_pe_1_5_0_int_q_acc_6_), .ZN(
        npu_inst_pe_1_5_0_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_5_0_U127 ( .A(npu_inst_pe_1_5_0_int_q_acc_7_), .B(
        npu_inst_pe_1_5_0_add_69_carry_7_), .Z(npu_inst_pe_1_5_0_N80) );
  XNOR2_X1 npu_inst_pe_1_5_0_U126 ( .A(npu_inst_pe_1_5_0_sub_67_carry_2_), .B(
        npu_inst_pe_1_5_0_int_q_acc_2_), .ZN(npu_inst_pe_1_5_0_N67) );
  OR2_X1 npu_inst_pe_1_5_0_U125 ( .A1(npu_inst_pe_1_5_0_int_q_acc_2_), .A2(
        npu_inst_pe_1_5_0_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_5_0_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_5_0_U124 ( .A(npu_inst_pe_1_5_0_sub_67_carry_3_), .B(
        npu_inst_pe_1_5_0_int_q_acc_3_), .ZN(npu_inst_pe_1_5_0_N68) );
  OR2_X1 npu_inst_pe_1_5_0_U123 ( .A1(npu_inst_pe_1_5_0_int_q_acc_3_), .A2(
        npu_inst_pe_1_5_0_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_5_0_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_5_0_U122 ( .A(npu_inst_pe_1_5_0_sub_67_carry_4_), .B(
        npu_inst_pe_1_5_0_int_q_acc_4_), .ZN(npu_inst_pe_1_5_0_N69) );
  OR2_X1 npu_inst_pe_1_5_0_U121 ( .A1(npu_inst_pe_1_5_0_int_q_acc_4_), .A2(
        npu_inst_pe_1_5_0_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_5_0_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_5_0_U120 ( .A(npu_inst_pe_1_5_0_sub_67_carry_5_), .B(
        npu_inst_pe_1_5_0_int_q_acc_5_), .ZN(npu_inst_pe_1_5_0_N70) );
  OR2_X1 npu_inst_pe_1_5_0_U119 ( .A1(npu_inst_pe_1_5_0_int_q_acc_5_), .A2(
        npu_inst_pe_1_5_0_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_5_0_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_5_0_U118 ( .A(npu_inst_pe_1_5_0_sub_67_carry_6_), .B(
        npu_inst_pe_1_5_0_int_q_acc_6_), .ZN(npu_inst_pe_1_5_0_N71) );
  OR2_X1 npu_inst_pe_1_5_0_U117 ( .A1(npu_inst_pe_1_5_0_int_q_acc_6_), .A2(
        npu_inst_pe_1_5_0_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_5_0_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_5_0_U116 ( .A(npu_inst_pe_1_5_0_int_q_acc_7_), .B(
        npu_inst_pe_1_5_0_sub_67_carry_7_), .ZN(npu_inst_pe_1_5_0_N72) );
  INV_X1 npu_inst_pe_1_5_0_U115 ( .A(npu_inst_n76), .ZN(npu_inst_pe_1_5_0_n6)
         );
  INV_X1 npu_inst_pe_1_5_0_U114 ( .A(npu_inst_n55), .ZN(npu_inst_pe_1_5_0_n3)
         );
  AOI22_X1 npu_inst_pe_1_5_0_U113 ( .A1(npu_inst_int_data_y_6__0__0_), .A2(
        npu_inst_pe_1_5_0_n58), .B1(npu_inst_pe_1_5_0_n118), .B2(
        npu_inst_pe_1_5_0_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_5_0_n57) );
  INV_X1 npu_inst_pe_1_5_0_U112 ( .A(npu_inst_pe_1_5_0_n57), .ZN(
        npu_inst_pe_1_5_0_n107) );
  AOI22_X1 npu_inst_pe_1_5_0_U111 ( .A1(npu_inst_int_data_y_6__0__0_), .A2(
        npu_inst_pe_1_5_0_n54), .B1(npu_inst_pe_1_5_0_n117), .B2(
        npu_inst_pe_1_5_0_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_5_0_n53) );
  INV_X1 npu_inst_pe_1_5_0_U110 ( .A(npu_inst_pe_1_5_0_n53), .ZN(
        npu_inst_pe_1_5_0_n108) );
  AOI22_X1 npu_inst_pe_1_5_0_U107 ( .A1(npu_inst_int_data_y_6__0__0_), .A2(
        npu_inst_pe_1_5_0_n50), .B1(npu_inst_pe_1_5_0_n116), .B2(
        npu_inst_pe_1_5_0_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_5_0_n49) );
  INV_X1 npu_inst_pe_1_5_0_U106 ( .A(npu_inst_pe_1_5_0_n49), .ZN(
        npu_inst_pe_1_5_0_n109) );
  AOI22_X1 npu_inst_pe_1_5_0_U105 ( .A1(npu_inst_int_data_y_6__0__0_), .A2(
        npu_inst_pe_1_5_0_n46), .B1(npu_inst_pe_1_5_0_n115), .B2(
        npu_inst_pe_1_5_0_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_5_0_n45) );
  INV_X1 npu_inst_pe_1_5_0_U104 ( .A(npu_inst_pe_1_5_0_n45), .ZN(
        npu_inst_pe_1_5_0_n110) );
  AOI22_X1 npu_inst_pe_1_5_0_U103 ( .A1(npu_inst_int_data_y_6__0__0_), .A2(
        npu_inst_pe_1_5_0_n42), .B1(npu_inst_pe_1_5_0_n114), .B2(
        npu_inst_pe_1_5_0_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_5_0_n41) );
  INV_X1 npu_inst_pe_1_5_0_U102 ( .A(npu_inst_pe_1_5_0_n41), .ZN(
        npu_inst_pe_1_5_0_n111) );
  AOI22_X1 npu_inst_pe_1_5_0_U101 ( .A1(npu_inst_int_data_y_6__0__1_), .A2(
        npu_inst_pe_1_5_0_n58), .B1(npu_inst_pe_1_5_0_n118), .B2(
        npu_inst_pe_1_5_0_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_5_0_n59) );
  INV_X1 npu_inst_pe_1_5_0_U100 ( .A(npu_inst_pe_1_5_0_n59), .ZN(
        npu_inst_pe_1_5_0_n101) );
  AOI22_X1 npu_inst_pe_1_5_0_U99 ( .A1(npu_inst_int_data_y_6__0__1_), .A2(
        npu_inst_pe_1_5_0_n54), .B1(npu_inst_pe_1_5_0_n117), .B2(
        npu_inst_pe_1_5_0_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_5_0_n55) );
  INV_X1 npu_inst_pe_1_5_0_U98 ( .A(npu_inst_pe_1_5_0_n55), .ZN(
        npu_inst_pe_1_5_0_n102) );
  AOI22_X1 npu_inst_pe_1_5_0_U97 ( .A1(npu_inst_int_data_y_6__0__1_), .A2(
        npu_inst_pe_1_5_0_n50), .B1(npu_inst_pe_1_5_0_n116), .B2(
        npu_inst_pe_1_5_0_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_5_0_n51) );
  INV_X1 npu_inst_pe_1_5_0_U96 ( .A(npu_inst_pe_1_5_0_n51), .ZN(
        npu_inst_pe_1_5_0_n103) );
  AOI22_X1 npu_inst_pe_1_5_0_U95 ( .A1(npu_inst_int_data_y_6__0__1_), .A2(
        npu_inst_pe_1_5_0_n46), .B1(npu_inst_pe_1_5_0_n115), .B2(
        npu_inst_pe_1_5_0_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_5_0_n47) );
  INV_X1 npu_inst_pe_1_5_0_U94 ( .A(npu_inst_pe_1_5_0_n47), .ZN(
        npu_inst_pe_1_5_0_n104) );
  AOI22_X1 npu_inst_pe_1_5_0_U93 ( .A1(npu_inst_int_data_y_6__0__1_), .A2(
        npu_inst_pe_1_5_0_n42), .B1(npu_inst_pe_1_5_0_n114), .B2(
        npu_inst_pe_1_5_0_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_5_0_n43) );
  INV_X1 npu_inst_pe_1_5_0_U92 ( .A(npu_inst_pe_1_5_0_n43), .ZN(
        npu_inst_pe_1_5_0_n105) );
  AOI22_X1 npu_inst_pe_1_5_0_U91 ( .A1(npu_inst_pe_1_5_0_n38), .A2(
        npu_inst_int_data_y_6__0__1_), .B1(npu_inst_pe_1_5_0_n113), .B2(
        npu_inst_pe_1_5_0_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_5_0_n39) );
  INV_X1 npu_inst_pe_1_5_0_U90 ( .A(npu_inst_pe_1_5_0_n39), .ZN(
        npu_inst_pe_1_5_0_n106) );
  AOI22_X1 npu_inst_pe_1_5_0_U89 ( .A1(npu_inst_pe_1_5_0_n38), .A2(
        npu_inst_int_data_y_6__0__0_), .B1(npu_inst_pe_1_5_0_n113), .B2(
        npu_inst_pe_1_5_0_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_5_0_n37) );
  INV_X1 npu_inst_pe_1_5_0_U88 ( .A(npu_inst_pe_1_5_0_n37), .ZN(
        npu_inst_pe_1_5_0_n112) );
  NAND2_X1 npu_inst_pe_1_5_0_U87 ( .A1(npu_inst_pe_1_5_0_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_5_0_n60), .ZN(npu_inst_pe_1_5_0_n74) );
  OAI21_X1 npu_inst_pe_1_5_0_U86 ( .B1(npu_inst_pe_1_5_0_n63), .B2(
        npu_inst_pe_1_5_0_n60), .A(npu_inst_pe_1_5_0_n74), .ZN(
        npu_inst_pe_1_5_0_n97) );
  NAND2_X1 npu_inst_pe_1_5_0_U85 ( .A1(npu_inst_pe_1_5_0_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_5_0_n60), .ZN(npu_inst_pe_1_5_0_n73) );
  OAI21_X1 npu_inst_pe_1_5_0_U84 ( .B1(npu_inst_pe_1_5_0_n61), .B2(
        npu_inst_pe_1_5_0_n60), .A(npu_inst_pe_1_5_0_n73), .ZN(
        npu_inst_pe_1_5_0_n96) );
  NAND2_X1 npu_inst_pe_1_5_0_U83 ( .A1(npu_inst_pe_1_5_0_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_5_0_n56), .ZN(npu_inst_pe_1_5_0_n72) );
  OAI21_X1 npu_inst_pe_1_5_0_U82 ( .B1(npu_inst_pe_1_5_0_n63), .B2(
        npu_inst_pe_1_5_0_n56), .A(npu_inst_pe_1_5_0_n72), .ZN(
        npu_inst_pe_1_5_0_n95) );
  NAND2_X1 npu_inst_pe_1_5_0_U81 ( .A1(npu_inst_pe_1_5_0_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_5_0_n56), .ZN(npu_inst_pe_1_5_0_n71) );
  OAI21_X1 npu_inst_pe_1_5_0_U80 ( .B1(npu_inst_pe_1_5_0_n61), .B2(
        npu_inst_pe_1_5_0_n56), .A(npu_inst_pe_1_5_0_n71), .ZN(
        npu_inst_pe_1_5_0_n94) );
  NAND2_X1 npu_inst_pe_1_5_0_U79 ( .A1(npu_inst_pe_1_5_0_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_5_0_n52), .ZN(npu_inst_pe_1_5_0_n70) );
  OAI21_X1 npu_inst_pe_1_5_0_U78 ( .B1(npu_inst_pe_1_5_0_n63), .B2(
        npu_inst_pe_1_5_0_n52), .A(npu_inst_pe_1_5_0_n70), .ZN(
        npu_inst_pe_1_5_0_n93) );
  NAND2_X1 npu_inst_pe_1_5_0_U77 ( .A1(npu_inst_pe_1_5_0_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_5_0_n52), .ZN(npu_inst_pe_1_5_0_n69) );
  OAI21_X1 npu_inst_pe_1_5_0_U76 ( .B1(npu_inst_pe_1_5_0_n61), .B2(
        npu_inst_pe_1_5_0_n52), .A(npu_inst_pe_1_5_0_n69), .ZN(
        npu_inst_pe_1_5_0_n92) );
  NAND2_X1 npu_inst_pe_1_5_0_U75 ( .A1(npu_inst_pe_1_5_0_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_5_0_n48), .ZN(npu_inst_pe_1_5_0_n68) );
  OAI21_X1 npu_inst_pe_1_5_0_U74 ( .B1(npu_inst_pe_1_5_0_n63), .B2(
        npu_inst_pe_1_5_0_n48), .A(npu_inst_pe_1_5_0_n68), .ZN(
        npu_inst_pe_1_5_0_n91) );
  NAND2_X1 npu_inst_pe_1_5_0_U73 ( .A1(npu_inst_pe_1_5_0_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_5_0_n48), .ZN(npu_inst_pe_1_5_0_n67) );
  OAI21_X1 npu_inst_pe_1_5_0_U72 ( .B1(npu_inst_pe_1_5_0_n61), .B2(
        npu_inst_pe_1_5_0_n48), .A(npu_inst_pe_1_5_0_n67), .ZN(
        npu_inst_pe_1_5_0_n90) );
  NAND2_X1 npu_inst_pe_1_5_0_U71 ( .A1(npu_inst_pe_1_5_0_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_5_0_n44), .ZN(npu_inst_pe_1_5_0_n66) );
  OAI21_X1 npu_inst_pe_1_5_0_U70 ( .B1(npu_inst_pe_1_5_0_n63), .B2(
        npu_inst_pe_1_5_0_n44), .A(npu_inst_pe_1_5_0_n66), .ZN(
        npu_inst_pe_1_5_0_n89) );
  NAND2_X1 npu_inst_pe_1_5_0_U69 ( .A1(npu_inst_pe_1_5_0_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_5_0_n44), .ZN(npu_inst_pe_1_5_0_n65) );
  OAI21_X1 npu_inst_pe_1_5_0_U68 ( .B1(npu_inst_pe_1_5_0_n61), .B2(
        npu_inst_pe_1_5_0_n44), .A(npu_inst_pe_1_5_0_n65), .ZN(
        npu_inst_pe_1_5_0_n88) );
  NAND2_X1 npu_inst_pe_1_5_0_U67 ( .A1(npu_inst_pe_1_5_0_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_5_0_n40), .ZN(npu_inst_pe_1_5_0_n64) );
  OAI21_X1 npu_inst_pe_1_5_0_U66 ( .B1(npu_inst_pe_1_5_0_n63), .B2(
        npu_inst_pe_1_5_0_n40), .A(npu_inst_pe_1_5_0_n64), .ZN(
        npu_inst_pe_1_5_0_n87) );
  NAND2_X1 npu_inst_pe_1_5_0_U65 ( .A1(npu_inst_pe_1_5_0_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_5_0_n40), .ZN(npu_inst_pe_1_5_0_n62) );
  OAI21_X1 npu_inst_pe_1_5_0_U64 ( .B1(npu_inst_pe_1_5_0_n61), .B2(
        npu_inst_pe_1_5_0_n40), .A(npu_inst_pe_1_5_0_n62), .ZN(
        npu_inst_pe_1_5_0_n86) );
  AND2_X1 npu_inst_pe_1_5_0_U63 ( .A1(npu_inst_pe_1_5_0_N93), .A2(npu_inst_n55), .ZN(npu_inst_int_data_y_5__0__0_) );
  AND2_X1 npu_inst_pe_1_5_0_U62 ( .A1(npu_inst_n55), .A2(npu_inst_pe_1_5_0_N94), .ZN(npu_inst_int_data_y_5__0__1_) );
  NOR3_X1 npu_inst_pe_1_5_0_U61 ( .A1(npu_inst_pe_1_5_0_n26), .A2(npu_inst_n55), .A3(npu_inst_int_ckg[23]), .ZN(npu_inst_pe_1_5_0_n85) );
  OR2_X1 npu_inst_pe_1_5_0_U60 ( .A1(npu_inst_pe_1_5_0_n85), .A2(
        npu_inst_pe_1_5_0_n2), .ZN(npu_inst_pe_1_5_0_N84) );
  AND2_X1 npu_inst_pe_1_5_0_U59 ( .A1(npu_inst_pe_1_5_0_int_q_acc_0_), .A2(
        npu_inst_pe_1_5_0_n1), .ZN(npu_inst_int_data_res_5__0__0_) );
  AND2_X1 npu_inst_pe_1_5_0_U58 ( .A1(npu_inst_pe_1_5_0_n2), .A2(
        npu_inst_pe_1_5_0_int_q_acc_7_), .ZN(npu_inst_int_data_res_5__0__7_)
         );
  AND2_X1 npu_inst_pe_1_5_0_U57 ( .A1(npu_inst_pe_1_5_0_int_q_acc_1_), .A2(
        npu_inst_pe_1_5_0_n1), .ZN(npu_inst_int_data_res_5__0__1_) );
  AND2_X1 npu_inst_pe_1_5_0_U56 ( .A1(npu_inst_pe_1_5_0_int_q_acc_2_), .A2(
        npu_inst_pe_1_5_0_n1), .ZN(npu_inst_int_data_res_5__0__2_) );
  AND2_X1 npu_inst_pe_1_5_0_U55 ( .A1(npu_inst_pe_1_5_0_int_q_acc_3_), .A2(
        npu_inst_pe_1_5_0_n2), .ZN(npu_inst_int_data_res_5__0__3_) );
  AND2_X1 npu_inst_pe_1_5_0_U54 ( .A1(npu_inst_pe_1_5_0_int_q_acc_4_), .A2(
        npu_inst_pe_1_5_0_n2), .ZN(npu_inst_int_data_res_5__0__4_) );
  AND2_X1 npu_inst_pe_1_5_0_U53 ( .A1(npu_inst_pe_1_5_0_int_q_acc_5_), .A2(
        npu_inst_pe_1_5_0_n2), .ZN(npu_inst_int_data_res_5__0__5_) );
  AND2_X1 npu_inst_pe_1_5_0_U52 ( .A1(npu_inst_pe_1_5_0_int_q_acc_6_), .A2(
        npu_inst_pe_1_5_0_n2), .ZN(npu_inst_int_data_res_5__0__6_) );
  AOI222_X1 npu_inst_pe_1_5_0_U51 ( .A1(npu_inst_int_data_res_6__0__0_), .A2(
        npu_inst_pe_1_5_0_n1), .B1(npu_inst_pe_1_5_0_N73), .B2(
        npu_inst_pe_1_5_0_n76), .C1(npu_inst_pe_1_5_0_N65), .C2(
        npu_inst_pe_1_5_0_n77), .ZN(npu_inst_pe_1_5_0_n84) );
  INV_X1 npu_inst_pe_1_5_0_U50 ( .A(npu_inst_pe_1_5_0_n84), .ZN(
        npu_inst_pe_1_5_0_n100) );
  AOI222_X1 npu_inst_pe_1_5_0_U49 ( .A1(npu_inst_int_data_res_6__0__7_), .A2(
        npu_inst_pe_1_5_0_n1), .B1(npu_inst_pe_1_5_0_N80), .B2(
        npu_inst_pe_1_5_0_n76), .C1(npu_inst_pe_1_5_0_N72), .C2(
        npu_inst_pe_1_5_0_n77), .ZN(npu_inst_pe_1_5_0_n75) );
  INV_X1 npu_inst_pe_1_5_0_U48 ( .A(npu_inst_pe_1_5_0_n75), .ZN(
        npu_inst_pe_1_5_0_n32) );
  AOI222_X1 npu_inst_pe_1_5_0_U47 ( .A1(npu_inst_int_data_res_6__0__1_), .A2(
        npu_inst_pe_1_5_0_n1), .B1(npu_inst_pe_1_5_0_N74), .B2(
        npu_inst_pe_1_5_0_n76), .C1(npu_inst_pe_1_5_0_N66), .C2(
        npu_inst_pe_1_5_0_n77), .ZN(npu_inst_pe_1_5_0_n83) );
  INV_X1 npu_inst_pe_1_5_0_U46 ( .A(npu_inst_pe_1_5_0_n83), .ZN(
        npu_inst_pe_1_5_0_n99) );
  AOI222_X1 npu_inst_pe_1_5_0_U45 ( .A1(npu_inst_int_data_res_6__0__2_), .A2(
        npu_inst_pe_1_5_0_n1), .B1(npu_inst_pe_1_5_0_N75), .B2(
        npu_inst_pe_1_5_0_n76), .C1(npu_inst_pe_1_5_0_N67), .C2(
        npu_inst_pe_1_5_0_n77), .ZN(npu_inst_pe_1_5_0_n82) );
  INV_X1 npu_inst_pe_1_5_0_U44 ( .A(npu_inst_pe_1_5_0_n82), .ZN(
        npu_inst_pe_1_5_0_n98) );
  AOI222_X1 npu_inst_pe_1_5_0_U43 ( .A1(npu_inst_int_data_res_6__0__3_), .A2(
        npu_inst_pe_1_5_0_n1), .B1(npu_inst_pe_1_5_0_N76), .B2(
        npu_inst_pe_1_5_0_n76), .C1(npu_inst_pe_1_5_0_N68), .C2(
        npu_inst_pe_1_5_0_n77), .ZN(npu_inst_pe_1_5_0_n81) );
  INV_X1 npu_inst_pe_1_5_0_U42 ( .A(npu_inst_pe_1_5_0_n81), .ZN(
        npu_inst_pe_1_5_0_n36) );
  AOI222_X1 npu_inst_pe_1_5_0_U41 ( .A1(npu_inst_int_data_res_6__0__4_), .A2(
        npu_inst_pe_1_5_0_n1), .B1(npu_inst_pe_1_5_0_N77), .B2(
        npu_inst_pe_1_5_0_n76), .C1(npu_inst_pe_1_5_0_N69), .C2(
        npu_inst_pe_1_5_0_n77), .ZN(npu_inst_pe_1_5_0_n80) );
  INV_X1 npu_inst_pe_1_5_0_U40 ( .A(npu_inst_pe_1_5_0_n80), .ZN(
        npu_inst_pe_1_5_0_n35) );
  AOI222_X1 npu_inst_pe_1_5_0_U39 ( .A1(npu_inst_int_data_res_6__0__5_), .A2(
        npu_inst_pe_1_5_0_n1), .B1(npu_inst_pe_1_5_0_N78), .B2(
        npu_inst_pe_1_5_0_n76), .C1(npu_inst_pe_1_5_0_N70), .C2(
        npu_inst_pe_1_5_0_n77), .ZN(npu_inst_pe_1_5_0_n79) );
  INV_X1 npu_inst_pe_1_5_0_U38 ( .A(npu_inst_pe_1_5_0_n79), .ZN(
        npu_inst_pe_1_5_0_n34) );
  AOI222_X1 npu_inst_pe_1_5_0_U37 ( .A1(npu_inst_int_data_res_6__0__6_), .A2(
        npu_inst_pe_1_5_0_n1), .B1(npu_inst_pe_1_5_0_N79), .B2(
        npu_inst_pe_1_5_0_n76), .C1(npu_inst_pe_1_5_0_N71), .C2(
        npu_inst_pe_1_5_0_n77), .ZN(npu_inst_pe_1_5_0_n78) );
  INV_X1 npu_inst_pe_1_5_0_U36 ( .A(npu_inst_pe_1_5_0_n78), .ZN(
        npu_inst_pe_1_5_0_n33) );
  AND2_X1 npu_inst_pe_1_5_0_U35 ( .A1(npu_inst_pe_1_5_0_o_data_h_1_), .A2(
        npu_inst_pe_1_5_0_int_q_weight_1_), .ZN(npu_inst_pe_1_5_0_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_5_0_U34 ( .A1(npu_inst_pe_1_5_0_o_data_h_0_), .A2(
        npu_inst_pe_1_5_0_int_q_weight_1_), .ZN(npu_inst_pe_1_5_0_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_5_0_U33 ( .A(npu_inst_pe_1_5_0_int_data_1_), .ZN(
        npu_inst_pe_1_5_0_n13) );
  AOI22_X1 npu_inst_pe_1_5_0_U32 ( .A1(npu_inst_n55), .A2(
        npu_inst_int_data_y_6__0__1_), .B1(npu_inst_pe_1_5_0_n3), .B2(
        npu_inst_int_data_x_5__1__1_), .ZN(npu_inst_pe_1_5_0_n63) );
  AOI22_X1 npu_inst_pe_1_5_0_U31 ( .A1(npu_inst_n55), .A2(
        npu_inst_int_data_y_6__0__0_), .B1(npu_inst_pe_1_5_0_n3), .B2(
        npu_inst_int_data_x_5__1__0_), .ZN(npu_inst_pe_1_5_0_n61) );
  INV_X1 npu_inst_pe_1_5_0_U30 ( .A(npu_inst_pe_1_5_0_int_data_0_), .ZN(
        npu_inst_pe_1_5_0_n12) );
  INV_X1 npu_inst_pe_1_5_0_U29 ( .A(npu_inst_n68), .ZN(npu_inst_pe_1_5_0_n5)
         );
  OR3_X1 npu_inst_pe_1_5_0_U28 ( .A1(npu_inst_n76), .A2(npu_inst_pe_1_5_0_n7), 
        .A3(npu_inst_pe_1_5_0_n5), .ZN(npu_inst_pe_1_5_0_n56) );
  OR3_X1 npu_inst_pe_1_5_0_U27 ( .A1(npu_inst_pe_1_5_0_n5), .A2(
        npu_inst_pe_1_5_0_n7), .A3(npu_inst_pe_1_5_0_n6), .ZN(
        npu_inst_pe_1_5_0_n48) );
  INV_X1 npu_inst_pe_1_5_0_U26 ( .A(npu_inst_pe_1_5_0_n5), .ZN(
        npu_inst_pe_1_5_0_n4) );
  OR3_X1 npu_inst_pe_1_5_0_U25 ( .A1(npu_inst_pe_1_5_0_n4), .A2(
        npu_inst_pe_1_5_0_n7), .A3(npu_inst_pe_1_5_0_n6), .ZN(
        npu_inst_pe_1_5_0_n52) );
  OR3_X1 npu_inst_pe_1_5_0_U24 ( .A1(npu_inst_n76), .A2(npu_inst_pe_1_5_0_n7), 
        .A3(npu_inst_pe_1_5_0_n4), .ZN(npu_inst_pe_1_5_0_n60) );
  NOR2_X1 npu_inst_pe_1_5_0_U23 ( .A1(npu_inst_pe_1_5_0_n60), .A2(
        npu_inst_pe_1_5_0_n3), .ZN(npu_inst_pe_1_5_0_n58) );
  NOR2_X1 npu_inst_pe_1_5_0_U22 ( .A1(npu_inst_pe_1_5_0_n56), .A2(
        npu_inst_pe_1_5_0_n3), .ZN(npu_inst_pe_1_5_0_n54) );
  NOR2_X1 npu_inst_pe_1_5_0_U21 ( .A1(npu_inst_pe_1_5_0_n52), .A2(
        npu_inst_pe_1_5_0_n3), .ZN(npu_inst_pe_1_5_0_n50) );
  NOR2_X1 npu_inst_pe_1_5_0_U20 ( .A1(npu_inst_pe_1_5_0_n48), .A2(
        npu_inst_pe_1_5_0_n3), .ZN(npu_inst_pe_1_5_0_n46) );
  NOR2_X1 npu_inst_pe_1_5_0_U19 ( .A1(npu_inst_pe_1_5_0_n40), .A2(
        npu_inst_pe_1_5_0_n3), .ZN(npu_inst_pe_1_5_0_n38) );
  NOR2_X1 npu_inst_pe_1_5_0_U18 ( .A1(npu_inst_pe_1_5_0_n44), .A2(
        npu_inst_pe_1_5_0_n3), .ZN(npu_inst_pe_1_5_0_n42) );
  BUF_X1 npu_inst_pe_1_5_0_U17 ( .A(npu_inst_n97), .Z(npu_inst_pe_1_5_0_n7) );
  INV_X1 npu_inst_pe_1_5_0_U16 ( .A(npu_inst_n123), .ZN(npu_inst_pe_1_5_0_n11)
         );
  INV_X1 npu_inst_pe_1_5_0_U15 ( .A(npu_inst_pe_1_5_0_n38), .ZN(
        npu_inst_pe_1_5_0_n113) );
  INV_X1 npu_inst_pe_1_5_0_U14 ( .A(npu_inst_pe_1_5_0_n58), .ZN(
        npu_inst_pe_1_5_0_n118) );
  INV_X1 npu_inst_pe_1_5_0_U13 ( .A(npu_inst_pe_1_5_0_n54), .ZN(
        npu_inst_pe_1_5_0_n117) );
  INV_X1 npu_inst_pe_1_5_0_U12 ( .A(npu_inst_pe_1_5_0_n50), .ZN(
        npu_inst_pe_1_5_0_n116) );
  INV_X1 npu_inst_pe_1_5_0_U11 ( .A(npu_inst_pe_1_5_0_n46), .ZN(
        npu_inst_pe_1_5_0_n115) );
  INV_X1 npu_inst_pe_1_5_0_U10 ( .A(npu_inst_pe_1_5_0_n42), .ZN(
        npu_inst_pe_1_5_0_n114) );
  BUF_X1 npu_inst_pe_1_5_0_U9 ( .A(npu_inst_n18), .Z(npu_inst_pe_1_5_0_n2) );
  BUF_X1 npu_inst_pe_1_5_0_U8 ( .A(npu_inst_n18), .Z(npu_inst_pe_1_5_0_n1) );
  BUF_X1 npu_inst_pe_1_5_0_U7 ( .A(npu_inst_pe_1_5_0_n11), .Z(
        npu_inst_pe_1_5_0_n10) );
  BUF_X1 npu_inst_pe_1_5_0_U6 ( .A(npu_inst_pe_1_5_0_n11), .Z(
        npu_inst_pe_1_5_0_n9) );
  BUF_X1 npu_inst_pe_1_5_0_U5 ( .A(npu_inst_pe_1_5_0_n11), .Z(
        npu_inst_pe_1_5_0_n8) );
  NOR2_X1 npu_inst_pe_1_5_0_U4 ( .A1(npu_inst_pe_1_5_0_int_q_weight_0_), .A2(
        npu_inst_pe_1_5_0_n1), .ZN(npu_inst_pe_1_5_0_n76) );
  NOR2_X1 npu_inst_pe_1_5_0_U3 ( .A1(npu_inst_pe_1_5_0_n27), .A2(
        npu_inst_pe_1_5_0_n1), .ZN(npu_inst_pe_1_5_0_n77) );
  FA_X1 npu_inst_pe_1_5_0_sub_67_U2_1 ( .A(npu_inst_pe_1_5_0_int_q_acc_1_), 
        .B(npu_inst_pe_1_5_0_n13), .CI(npu_inst_pe_1_5_0_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_5_0_sub_67_carry_2_), .S(npu_inst_pe_1_5_0_N66) );
  FA_X1 npu_inst_pe_1_5_0_add_69_U1_1 ( .A(npu_inst_pe_1_5_0_int_q_acc_1_), 
        .B(npu_inst_pe_1_5_0_int_data_1_), .CI(
        npu_inst_pe_1_5_0_add_69_carry_1_), .CO(
        npu_inst_pe_1_5_0_add_69_carry_2_), .S(npu_inst_pe_1_5_0_N74) );
  NAND3_X1 npu_inst_pe_1_5_0_U109 ( .A1(npu_inst_pe_1_5_0_n5), .A2(
        npu_inst_pe_1_5_0_n6), .A3(npu_inst_pe_1_5_0_n7), .ZN(
        npu_inst_pe_1_5_0_n44) );
  NAND3_X1 npu_inst_pe_1_5_0_U108 ( .A1(npu_inst_pe_1_5_0_n4), .A2(
        npu_inst_pe_1_5_0_n6), .A3(npu_inst_pe_1_5_0_n7), .ZN(
        npu_inst_pe_1_5_0_n40) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_5_0_n33), .CK(
        npu_inst_pe_1_5_0_net3642), .RN(npu_inst_pe_1_5_0_n8), .Q(
        npu_inst_pe_1_5_0_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_5_0_n34), .CK(
        npu_inst_pe_1_5_0_net3642), .RN(npu_inst_pe_1_5_0_n8), .Q(
        npu_inst_pe_1_5_0_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_5_0_n35), .CK(
        npu_inst_pe_1_5_0_net3642), .RN(npu_inst_pe_1_5_0_n8), .Q(
        npu_inst_pe_1_5_0_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_5_0_n36), .CK(
        npu_inst_pe_1_5_0_net3642), .RN(npu_inst_pe_1_5_0_n8), .Q(
        npu_inst_pe_1_5_0_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_5_0_n98), .CK(
        npu_inst_pe_1_5_0_net3642), .RN(npu_inst_pe_1_5_0_n8), .Q(
        npu_inst_pe_1_5_0_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_5_0_n99), .CK(
        npu_inst_pe_1_5_0_net3642), .RN(npu_inst_pe_1_5_0_n8), .Q(
        npu_inst_pe_1_5_0_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_5_0_n32), .CK(
        npu_inst_pe_1_5_0_net3642), .RN(npu_inst_pe_1_5_0_n8), .Q(
        npu_inst_pe_1_5_0_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_5_0_n100), 
        .CK(npu_inst_pe_1_5_0_net3642), .RN(npu_inst_pe_1_5_0_n8), .Q(
        npu_inst_pe_1_5_0_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_weight_reg_0_ ( .D(npu_inst_n109), .CK(
        npu_inst_pe_1_5_0_net3648), .RN(npu_inst_pe_1_5_0_n8), .Q(
        npu_inst_pe_1_5_0_int_q_weight_0_), .QN(npu_inst_pe_1_5_0_n27) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_weight_reg_1_ ( .D(npu_inst_n115), .CK(
        npu_inst_pe_1_5_0_net3648), .RN(npu_inst_pe_1_5_0_n8), .Q(
        npu_inst_pe_1_5_0_int_q_weight_1_), .QN(npu_inst_pe_1_5_0_n26) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_5_0_n112), 
        .CK(npu_inst_pe_1_5_0_net3648), .RN(npu_inst_pe_1_5_0_n8), .Q(
        npu_inst_pe_1_5_0_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_5_0_n106), 
        .CK(npu_inst_pe_1_5_0_net3648), .RN(npu_inst_pe_1_5_0_n8), .Q(
        npu_inst_pe_1_5_0_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_5_0_n111), 
        .CK(npu_inst_pe_1_5_0_net3648), .RN(npu_inst_pe_1_5_0_n9), .Q(
        npu_inst_pe_1_5_0_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_5_0_n105), 
        .CK(npu_inst_pe_1_5_0_net3648), .RN(npu_inst_pe_1_5_0_n9), .Q(
        npu_inst_pe_1_5_0_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_5_0_n110), 
        .CK(npu_inst_pe_1_5_0_net3648), .RN(npu_inst_pe_1_5_0_n9), .Q(
        npu_inst_pe_1_5_0_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_5_0_n104), 
        .CK(npu_inst_pe_1_5_0_net3648), .RN(npu_inst_pe_1_5_0_n9), .Q(
        npu_inst_pe_1_5_0_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_5_0_n109), 
        .CK(npu_inst_pe_1_5_0_net3648), .RN(npu_inst_pe_1_5_0_n9), .Q(
        npu_inst_pe_1_5_0_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_5_0_n103), 
        .CK(npu_inst_pe_1_5_0_net3648), .RN(npu_inst_pe_1_5_0_n9), .Q(
        npu_inst_pe_1_5_0_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_5_0_n108), 
        .CK(npu_inst_pe_1_5_0_net3648), .RN(npu_inst_pe_1_5_0_n9), .Q(
        npu_inst_pe_1_5_0_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_5_0_n102), 
        .CK(npu_inst_pe_1_5_0_net3648), .RN(npu_inst_pe_1_5_0_n9), .Q(
        npu_inst_pe_1_5_0_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_5_0_n107), 
        .CK(npu_inst_pe_1_5_0_net3648), .RN(npu_inst_pe_1_5_0_n9), .Q(
        npu_inst_pe_1_5_0_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_5_0_n101), 
        .CK(npu_inst_pe_1_5_0_net3648), .RN(npu_inst_pe_1_5_0_n9), .Q(
        npu_inst_pe_1_5_0_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_5_0_n86), 
        .CK(npu_inst_pe_1_5_0_net3648), .RN(npu_inst_pe_1_5_0_n9), .Q(
        npu_inst_pe_1_5_0_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_5_0_n87), 
        .CK(npu_inst_pe_1_5_0_net3648), .RN(npu_inst_pe_1_5_0_n9), .Q(
        npu_inst_pe_1_5_0_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_5_0_n88), 
        .CK(npu_inst_pe_1_5_0_net3648), .RN(npu_inst_pe_1_5_0_n10), .Q(
        npu_inst_pe_1_5_0_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_5_0_n89), 
        .CK(npu_inst_pe_1_5_0_net3648), .RN(npu_inst_pe_1_5_0_n10), .Q(
        npu_inst_pe_1_5_0_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_5_0_n90), 
        .CK(npu_inst_pe_1_5_0_net3648), .RN(npu_inst_pe_1_5_0_n10), .Q(
        npu_inst_pe_1_5_0_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_5_0_n91), 
        .CK(npu_inst_pe_1_5_0_net3648), .RN(npu_inst_pe_1_5_0_n10), .Q(
        npu_inst_pe_1_5_0_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_5_0_n92), 
        .CK(npu_inst_pe_1_5_0_net3648), .RN(npu_inst_pe_1_5_0_n10), .Q(
        npu_inst_pe_1_5_0_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_5_0_n93), 
        .CK(npu_inst_pe_1_5_0_net3648), .RN(npu_inst_pe_1_5_0_n10), .Q(
        npu_inst_pe_1_5_0_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_5_0_n94), 
        .CK(npu_inst_pe_1_5_0_net3648), .RN(npu_inst_pe_1_5_0_n10), .Q(
        npu_inst_pe_1_5_0_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_5_0_n95), 
        .CK(npu_inst_pe_1_5_0_net3648), .RN(npu_inst_pe_1_5_0_n10), .Q(
        npu_inst_pe_1_5_0_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_5_0_n96), 
        .CK(npu_inst_pe_1_5_0_net3648), .RN(npu_inst_pe_1_5_0_n10), .Q(
        npu_inst_pe_1_5_0_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_5_0_n97), 
        .CK(npu_inst_pe_1_5_0_net3648), .RN(npu_inst_pe_1_5_0_n10), .Q(
        npu_inst_pe_1_5_0_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_5_0_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_5_0_N84), .SE(1'b0), .GCK(npu_inst_pe_1_5_0_net3642) );
  CLKGATETST_X1 npu_inst_pe_1_5_0_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n63), .SE(1'b0), .GCK(npu_inst_pe_1_5_0_net3648) );
  MUX2_X1 npu_inst_pe_1_5_1_U162 ( .A(npu_inst_pe_1_5_1_n32), .B(
        npu_inst_pe_1_5_1_n29), .S(npu_inst_pe_1_5_1_n8), .Z(
        npu_inst_pe_1_5_1_N93) );
  MUX2_X1 npu_inst_pe_1_5_1_U161 ( .A(npu_inst_pe_1_5_1_n31), .B(
        npu_inst_pe_1_5_1_n30), .S(npu_inst_pe_1_5_1_n6), .Z(
        npu_inst_pe_1_5_1_n32) );
  MUX2_X1 npu_inst_pe_1_5_1_U160 ( .A(npu_inst_pe_1_5_1_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_5_1_int_q_reg_v_1__0_), .S(npu_inst_pe_1_5_1_n4), .Z(
        npu_inst_pe_1_5_1_n31) );
  MUX2_X1 npu_inst_pe_1_5_1_U159 ( .A(npu_inst_pe_1_5_1_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_5_1_int_q_reg_v_3__0_), .S(npu_inst_pe_1_5_1_n4), .Z(
        npu_inst_pe_1_5_1_n30) );
  MUX2_X1 npu_inst_pe_1_5_1_U158 ( .A(npu_inst_pe_1_5_1_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_5_1_int_q_reg_v_5__0_), .S(npu_inst_pe_1_5_1_n4), .Z(
        npu_inst_pe_1_5_1_n29) );
  MUX2_X1 npu_inst_pe_1_5_1_U157 ( .A(npu_inst_pe_1_5_1_n28), .B(
        npu_inst_pe_1_5_1_n23), .S(npu_inst_pe_1_5_1_n8), .Z(
        npu_inst_pe_1_5_1_N94) );
  MUX2_X1 npu_inst_pe_1_5_1_U156 ( .A(npu_inst_pe_1_5_1_n25), .B(
        npu_inst_pe_1_5_1_n24), .S(npu_inst_pe_1_5_1_n6), .Z(
        npu_inst_pe_1_5_1_n28) );
  MUX2_X1 npu_inst_pe_1_5_1_U155 ( .A(npu_inst_pe_1_5_1_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_5_1_int_q_reg_v_1__1_), .S(npu_inst_pe_1_5_1_n4), .Z(
        npu_inst_pe_1_5_1_n25) );
  MUX2_X1 npu_inst_pe_1_5_1_U154 ( .A(npu_inst_pe_1_5_1_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_5_1_int_q_reg_v_3__1_), .S(npu_inst_pe_1_5_1_n4), .Z(
        npu_inst_pe_1_5_1_n24) );
  MUX2_X1 npu_inst_pe_1_5_1_U153 ( .A(npu_inst_pe_1_5_1_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_5_1_int_q_reg_v_5__1_), .S(npu_inst_pe_1_5_1_n4), .Z(
        npu_inst_pe_1_5_1_n23) );
  MUX2_X1 npu_inst_pe_1_5_1_U152 ( .A(npu_inst_pe_1_5_1_n22), .B(
        npu_inst_pe_1_5_1_n19), .S(npu_inst_pe_1_5_1_n8), .Z(
        npu_inst_int_data_x_5__1__1_) );
  MUX2_X1 npu_inst_pe_1_5_1_U151 ( .A(npu_inst_pe_1_5_1_n21), .B(
        npu_inst_pe_1_5_1_n20), .S(npu_inst_pe_1_5_1_n6), .Z(
        npu_inst_pe_1_5_1_n22) );
  MUX2_X1 npu_inst_pe_1_5_1_U150 ( .A(npu_inst_pe_1_5_1_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_5_1_int_q_reg_h_1__1_), .S(npu_inst_pe_1_5_1_n4), .Z(
        npu_inst_pe_1_5_1_n21) );
  MUX2_X1 npu_inst_pe_1_5_1_U149 ( .A(npu_inst_pe_1_5_1_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_5_1_int_q_reg_h_3__1_), .S(npu_inst_pe_1_5_1_n4), .Z(
        npu_inst_pe_1_5_1_n20) );
  MUX2_X1 npu_inst_pe_1_5_1_U148 ( .A(npu_inst_pe_1_5_1_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_5_1_int_q_reg_h_5__1_), .S(npu_inst_pe_1_5_1_n4), .Z(
        npu_inst_pe_1_5_1_n19) );
  MUX2_X1 npu_inst_pe_1_5_1_U147 ( .A(npu_inst_pe_1_5_1_n18), .B(
        npu_inst_pe_1_5_1_n15), .S(npu_inst_pe_1_5_1_n8), .Z(
        npu_inst_int_data_x_5__1__0_) );
  MUX2_X1 npu_inst_pe_1_5_1_U146 ( .A(npu_inst_pe_1_5_1_n17), .B(
        npu_inst_pe_1_5_1_n16), .S(npu_inst_pe_1_5_1_n6), .Z(
        npu_inst_pe_1_5_1_n18) );
  MUX2_X1 npu_inst_pe_1_5_1_U145 ( .A(npu_inst_pe_1_5_1_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_5_1_int_q_reg_h_1__0_), .S(npu_inst_pe_1_5_1_n4), .Z(
        npu_inst_pe_1_5_1_n17) );
  MUX2_X1 npu_inst_pe_1_5_1_U144 ( .A(npu_inst_pe_1_5_1_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_5_1_int_q_reg_h_3__0_), .S(npu_inst_pe_1_5_1_n4), .Z(
        npu_inst_pe_1_5_1_n16) );
  MUX2_X1 npu_inst_pe_1_5_1_U143 ( .A(npu_inst_pe_1_5_1_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_5_1_int_q_reg_h_5__0_), .S(npu_inst_pe_1_5_1_n4), .Z(
        npu_inst_pe_1_5_1_n15) );
  XOR2_X1 npu_inst_pe_1_5_1_U142 ( .A(npu_inst_pe_1_5_1_int_data_0_), .B(
        npu_inst_pe_1_5_1_int_q_acc_0_), .Z(npu_inst_pe_1_5_1_N73) );
  AND2_X1 npu_inst_pe_1_5_1_U141 ( .A1(npu_inst_pe_1_5_1_int_q_acc_0_), .A2(
        npu_inst_pe_1_5_1_int_data_0_), .ZN(npu_inst_pe_1_5_1_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_5_1_U140 ( .A(npu_inst_pe_1_5_1_int_q_acc_0_), .B(
        npu_inst_pe_1_5_1_n13), .ZN(npu_inst_pe_1_5_1_N65) );
  OR2_X1 npu_inst_pe_1_5_1_U139 ( .A1(npu_inst_pe_1_5_1_n13), .A2(
        npu_inst_pe_1_5_1_int_q_acc_0_), .ZN(npu_inst_pe_1_5_1_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_5_1_U138 ( .A(npu_inst_pe_1_5_1_int_q_acc_2_), .B(
        npu_inst_pe_1_5_1_add_69_carry_2_), .Z(npu_inst_pe_1_5_1_N75) );
  AND2_X1 npu_inst_pe_1_5_1_U137 ( .A1(npu_inst_pe_1_5_1_add_69_carry_2_), 
        .A2(npu_inst_pe_1_5_1_int_q_acc_2_), .ZN(
        npu_inst_pe_1_5_1_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_5_1_U136 ( .A(npu_inst_pe_1_5_1_int_q_acc_3_), .B(
        npu_inst_pe_1_5_1_add_69_carry_3_), .Z(npu_inst_pe_1_5_1_N76) );
  AND2_X1 npu_inst_pe_1_5_1_U135 ( .A1(npu_inst_pe_1_5_1_add_69_carry_3_), 
        .A2(npu_inst_pe_1_5_1_int_q_acc_3_), .ZN(
        npu_inst_pe_1_5_1_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_5_1_U134 ( .A(npu_inst_pe_1_5_1_int_q_acc_4_), .B(
        npu_inst_pe_1_5_1_add_69_carry_4_), .Z(npu_inst_pe_1_5_1_N77) );
  AND2_X1 npu_inst_pe_1_5_1_U133 ( .A1(npu_inst_pe_1_5_1_add_69_carry_4_), 
        .A2(npu_inst_pe_1_5_1_int_q_acc_4_), .ZN(
        npu_inst_pe_1_5_1_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_5_1_U132 ( .A(npu_inst_pe_1_5_1_int_q_acc_5_), .B(
        npu_inst_pe_1_5_1_add_69_carry_5_), .Z(npu_inst_pe_1_5_1_N78) );
  AND2_X1 npu_inst_pe_1_5_1_U131 ( .A1(npu_inst_pe_1_5_1_add_69_carry_5_), 
        .A2(npu_inst_pe_1_5_1_int_q_acc_5_), .ZN(
        npu_inst_pe_1_5_1_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_5_1_U130 ( .A(npu_inst_pe_1_5_1_int_q_acc_6_), .B(
        npu_inst_pe_1_5_1_add_69_carry_6_), .Z(npu_inst_pe_1_5_1_N79) );
  AND2_X1 npu_inst_pe_1_5_1_U129 ( .A1(npu_inst_pe_1_5_1_add_69_carry_6_), 
        .A2(npu_inst_pe_1_5_1_int_q_acc_6_), .ZN(
        npu_inst_pe_1_5_1_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_5_1_U128 ( .A(npu_inst_pe_1_5_1_int_q_acc_7_), .B(
        npu_inst_pe_1_5_1_add_69_carry_7_), .Z(npu_inst_pe_1_5_1_N80) );
  XNOR2_X1 npu_inst_pe_1_5_1_U127 ( .A(npu_inst_pe_1_5_1_sub_67_carry_2_), .B(
        npu_inst_pe_1_5_1_int_q_acc_2_), .ZN(npu_inst_pe_1_5_1_N67) );
  OR2_X1 npu_inst_pe_1_5_1_U126 ( .A1(npu_inst_pe_1_5_1_int_q_acc_2_), .A2(
        npu_inst_pe_1_5_1_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_5_1_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_5_1_U125 ( .A(npu_inst_pe_1_5_1_sub_67_carry_3_), .B(
        npu_inst_pe_1_5_1_int_q_acc_3_), .ZN(npu_inst_pe_1_5_1_N68) );
  OR2_X1 npu_inst_pe_1_5_1_U124 ( .A1(npu_inst_pe_1_5_1_int_q_acc_3_), .A2(
        npu_inst_pe_1_5_1_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_5_1_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_5_1_U123 ( .A(npu_inst_pe_1_5_1_sub_67_carry_4_), .B(
        npu_inst_pe_1_5_1_int_q_acc_4_), .ZN(npu_inst_pe_1_5_1_N69) );
  OR2_X1 npu_inst_pe_1_5_1_U122 ( .A1(npu_inst_pe_1_5_1_int_q_acc_4_), .A2(
        npu_inst_pe_1_5_1_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_5_1_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_5_1_U121 ( .A(npu_inst_pe_1_5_1_sub_67_carry_5_), .B(
        npu_inst_pe_1_5_1_int_q_acc_5_), .ZN(npu_inst_pe_1_5_1_N70) );
  OR2_X1 npu_inst_pe_1_5_1_U120 ( .A1(npu_inst_pe_1_5_1_int_q_acc_5_), .A2(
        npu_inst_pe_1_5_1_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_5_1_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_5_1_U119 ( .A(npu_inst_pe_1_5_1_sub_67_carry_6_), .B(
        npu_inst_pe_1_5_1_int_q_acc_6_), .ZN(npu_inst_pe_1_5_1_N71) );
  OR2_X1 npu_inst_pe_1_5_1_U118 ( .A1(npu_inst_pe_1_5_1_int_q_acc_6_), .A2(
        npu_inst_pe_1_5_1_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_5_1_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_5_1_U117 ( .A(npu_inst_pe_1_5_1_int_q_acc_7_), .B(
        npu_inst_pe_1_5_1_sub_67_carry_7_), .ZN(npu_inst_pe_1_5_1_N72) );
  INV_X1 npu_inst_pe_1_5_1_U116 ( .A(npu_inst_n76), .ZN(npu_inst_pe_1_5_1_n7)
         );
  INV_X1 npu_inst_pe_1_5_1_U115 ( .A(npu_inst_pe_1_5_1_n7), .ZN(
        npu_inst_pe_1_5_1_n6) );
  INV_X1 npu_inst_pe_1_5_1_U114 ( .A(npu_inst_n55), .ZN(npu_inst_pe_1_5_1_n3)
         );
  AOI22_X1 npu_inst_pe_1_5_1_U113 ( .A1(npu_inst_int_data_y_6__1__0_), .A2(
        npu_inst_pe_1_5_1_n58), .B1(npu_inst_pe_1_5_1_n119), .B2(
        npu_inst_pe_1_5_1_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_5_1_n57) );
  INV_X1 npu_inst_pe_1_5_1_U112 ( .A(npu_inst_pe_1_5_1_n57), .ZN(
        npu_inst_pe_1_5_1_n108) );
  AOI22_X1 npu_inst_pe_1_5_1_U111 ( .A1(npu_inst_int_data_y_6__1__0_), .A2(
        npu_inst_pe_1_5_1_n54), .B1(npu_inst_pe_1_5_1_n118), .B2(
        npu_inst_pe_1_5_1_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_5_1_n53) );
  INV_X1 npu_inst_pe_1_5_1_U110 ( .A(npu_inst_pe_1_5_1_n53), .ZN(
        npu_inst_pe_1_5_1_n109) );
  AOI22_X1 npu_inst_pe_1_5_1_U107 ( .A1(npu_inst_int_data_y_6__1__0_), .A2(
        npu_inst_pe_1_5_1_n50), .B1(npu_inst_pe_1_5_1_n117), .B2(
        npu_inst_pe_1_5_1_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_5_1_n49) );
  INV_X1 npu_inst_pe_1_5_1_U106 ( .A(npu_inst_pe_1_5_1_n49), .ZN(
        npu_inst_pe_1_5_1_n110) );
  AOI22_X1 npu_inst_pe_1_5_1_U105 ( .A1(npu_inst_int_data_y_6__1__0_), .A2(
        npu_inst_pe_1_5_1_n46), .B1(npu_inst_pe_1_5_1_n116), .B2(
        npu_inst_pe_1_5_1_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_5_1_n45) );
  INV_X1 npu_inst_pe_1_5_1_U104 ( .A(npu_inst_pe_1_5_1_n45), .ZN(
        npu_inst_pe_1_5_1_n111) );
  AOI22_X1 npu_inst_pe_1_5_1_U103 ( .A1(npu_inst_int_data_y_6__1__0_), .A2(
        npu_inst_pe_1_5_1_n42), .B1(npu_inst_pe_1_5_1_n115), .B2(
        npu_inst_pe_1_5_1_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_5_1_n41) );
  INV_X1 npu_inst_pe_1_5_1_U102 ( .A(npu_inst_pe_1_5_1_n41), .ZN(
        npu_inst_pe_1_5_1_n112) );
  AOI22_X1 npu_inst_pe_1_5_1_U101 ( .A1(npu_inst_int_data_y_6__1__1_), .A2(
        npu_inst_pe_1_5_1_n58), .B1(npu_inst_pe_1_5_1_n119), .B2(
        npu_inst_pe_1_5_1_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_5_1_n59) );
  INV_X1 npu_inst_pe_1_5_1_U100 ( .A(npu_inst_pe_1_5_1_n59), .ZN(
        npu_inst_pe_1_5_1_n102) );
  AOI22_X1 npu_inst_pe_1_5_1_U99 ( .A1(npu_inst_int_data_y_6__1__1_), .A2(
        npu_inst_pe_1_5_1_n54), .B1(npu_inst_pe_1_5_1_n118), .B2(
        npu_inst_pe_1_5_1_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_5_1_n55) );
  INV_X1 npu_inst_pe_1_5_1_U98 ( .A(npu_inst_pe_1_5_1_n55), .ZN(
        npu_inst_pe_1_5_1_n103) );
  AOI22_X1 npu_inst_pe_1_5_1_U97 ( .A1(npu_inst_int_data_y_6__1__1_), .A2(
        npu_inst_pe_1_5_1_n50), .B1(npu_inst_pe_1_5_1_n117), .B2(
        npu_inst_pe_1_5_1_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_5_1_n51) );
  INV_X1 npu_inst_pe_1_5_1_U96 ( .A(npu_inst_pe_1_5_1_n51), .ZN(
        npu_inst_pe_1_5_1_n104) );
  AOI22_X1 npu_inst_pe_1_5_1_U95 ( .A1(npu_inst_int_data_y_6__1__1_), .A2(
        npu_inst_pe_1_5_1_n46), .B1(npu_inst_pe_1_5_1_n116), .B2(
        npu_inst_pe_1_5_1_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_5_1_n47) );
  INV_X1 npu_inst_pe_1_5_1_U94 ( .A(npu_inst_pe_1_5_1_n47), .ZN(
        npu_inst_pe_1_5_1_n105) );
  AOI22_X1 npu_inst_pe_1_5_1_U93 ( .A1(npu_inst_int_data_y_6__1__1_), .A2(
        npu_inst_pe_1_5_1_n42), .B1(npu_inst_pe_1_5_1_n115), .B2(
        npu_inst_pe_1_5_1_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_5_1_n43) );
  INV_X1 npu_inst_pe_1_5_1_U92 ( .A(npu_inst_pe_1_5_1_n43), .ZN(
        npu_inst_pe_1_5_1_n106) );
  AOI22_X1 npu_inst_pe_1_5_1_U91 ( .A1(npu_inst_pe_1_5_1_n38), .A2(
        npu_inst_int_data_y_6__1__1_), .B1(npu_inst_pe_1_5_1_n114), .B2(
        npu_inst_pe_1_5_1_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_5_1_n39) );
  INV_X1 npu_inst_pe_1_5_1_U90 ( .A(npu_inst_pe_1_5_1_n39), .ZN(
        npu_inst_pe_1_5_1_n107) );
  AOI22_X1 npu_inst_pe_1_5_1_U89 ( .A1(npu_inst_pe_1_5_1_n38), .A2(
        npu_inst_int_data_y_6__1__0_), .B1(npu_inst_pe_1_5_1_n114), .B2(
        npu_inst_pe_1_5_1_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_5_1_n37) );
  INV_X1 npu_inst_pe_1_5_1_U88 ( .A(npu_inst_pe_1_5_1_n37), .ZN(
        npu_inst_pe_1_5_1_n113) );
  NAND2_X1 npu_inst_pe_1_5_1_U87 ( .A1(npu_inst_pe_1_5_1_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_5_1_n60), .ZN(npu_inst_pe_1_5_1_n74) );
  OAI21_X1 npu_inst_pe_1_5_1_U86 ( .B1(npu_inst_pe_1_5_1_n63), .B2(
        npu_inst_pe_1_5_1_n60), .A(npu_inst_pe_1_5_1_n74), .ZN(
        npu_inst_pe_1_5_1_n97) );
  NAND2_X1 npu_inst_pe_1_5_1_U85 ( .A1(npu_inst_pe_1_5_1_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_5_1_n60), .ZN(npu_inst_pe_1_5_1_n73) );
  OAI21_X1 npu_inst_pe_1_5_1_U84 ( .B1(npu_inst_pe_1_5_1_n61), .B2(
        npu_inst_pe_1_5_1_n60), .A(npu_inst_pe_1_5_1_n73), .ZN(
        npu_inst_pe_1_5_1_n96) );
  NAND2_X1 npu_inst_pe_1_5_1_U83 ( .A1(npu_inst_pe_1_5_1_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_5_1_n56), .ZN(npu_inst_pe_1_5_1_n72) );
  OAI21_X1 npu_inst_pe_1_5_1_U82 ( .B1(npu_inst_pe_1_5_1_n63), .B2(
        npu_inst_pe_1_5_1_n56), .A(npu_inst_pe_1_5_1_n72), .ZN(
        npu_inst_pe_1_5_1_n95) );
  NAND2_X1 npu_inst_pe_1_5_1_U81 ( .A1(npu_inst_pe_1_5_1_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_5_1_n56), .ZN(npu_inst_pe_1_5_1_n71) );
  OAI21_X1 npu_inst_pe_1_5_1_U80 ( .B1(npu_inst_pe_1_5_1_n61), .B2(
        npu_inst_pe_1_5_1_n56), .A(npu_inst_pe_1_5_1_n71), .ZN(
        npu_inst_pe_1_5_1_n94) );
  NAND2_X1 npu_inst_pe_1_5_1_U79 ( .A1(npu_inst_pe_1_5_1_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_5_1_n52), .ZN(npu_inst_pe_1_5_1_n70) );
  OAI21_X1 npu_inst_pe_1_5_1_U78 ( .B1(npu_inst_pe_1_5_1_n63), .B2(
        npu_inst_pe_1_5_1_n52), .A(npu_inst_pe_1_5_1_n70), .ZN(
        npu_inst_pe_1_5_1_n93) );
  NAND2_X1 npu_inst_pe_1_5_1_U77 ( .A1(npu_inst_pe_1_5_1_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_5_1_n52), .ZN(npu_inst_pe_1_5_1_n69) );
  OAI21_X1 npu_inst_pe_1_5_1_U76 ( .B1(npu_inst_pe_1_5_1_n61), .B2(
        npu_inst_pe_1_5_1_n52), .A(npu_inst_pe_1_5_1_n69), .ZN(
        npu_inst_pe_1_5_1_n92) );
  NAND2_X1 npu_inst_pe_1_5_1_U75 ( .A1(npu_inst_pe_1_5_1_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_5_1_n48), .ZN(npu_inst_pe_1_5_1_n68) );
  OAI21_X1 npu_inst_pe_1_5_1_U74 ( .B1(npu_inst_pe_1_5_1_n63), .B2(
        npu_inst_pe_1_5_1_n48), .A(npu_inst_pe_1_5_1_n68), .ZN(
        npu_inst_pe_1_5_1_n91) );
  NAND2_X1 npu_inst_pe_1_5_1_U73 ( .A1(npu_inst_pe_1_5_1_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_5_1_n48), .ZN(npu_inst_pe_1_5_1_n67) );
  OAI21_X1 npu_inst_pe_1_5_1_U72 ( .B1(npu_inst_pe_1_5_1_n61), .B2(
        npu_inst_pe_1_5_1_n48), .A(npu_inst_pe_1_5_1_n67), .ZN(
        npu_inst_pe_1_5_1_n90) );
  NAND2_X1 npu_inst_pe_1_5_1_U71 ( .A1(npu_inst_pe_1_5_1_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_5_1_n44), .ZN(npu_inst_pe_1_5_1_n66) );
  OAI21_X1 npu_inst_pe_1_5_1_U70 ( .B1(npu_inst_pe_1_5_1_n63), .B2(
        npu_inst_pe_1_5_1_n44), .A(npu_inst_pe_1_5_1_n66), .ZN(
        npu_inst_pe_1_5_1_n89) );
  NAND2_X1 npu_inst_pe_1_5_1_U69 ( .A1(npu_inst_pe_1_5_1_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_5_1_n44), .ZN(npu_inst_pe_1_5_1_n65) );
  OAI21_X1 npu_inst_pe_1_5_1_U68 ( .B1(npu_inst_pe_1_5_1_n61), .B2(
        npu_inst_pe_1_5_1_n44), .A(npu_inst_pe_1_5_1_n65), .ZN(
        npu_inst_pe_1_5_1_n88) );
  NAND2_X1 npu_inst_pe_1_5_1_U67 ( .A1(npu_inst_pe_1_5_1_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_5_1_n40), .ZN(npu_inst_pe_1_5_1_n64) );
  OAI21_X1 npu_inst_pe_1_5_1_U66 ( .B1(npu_inst_pe_1_5_1_n63), .B2(
        npu_inst_pe_1_5_1_n40), .A(npu_inst_pe_1_5_1_n64), .ZN(
        npu_inst_pe_1_5_1_n87) );
  NAND2_X1 npu_inst_pe_1_5_1_U65 ( .A1(npu_inst_pe_1_5_1_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_5_1_n40), .ZN(npu_inst_pe_1_5_1_n62) );
  OAI21_X1 npu_inst_pe_1_5_1_U64 ( .B1(npu_inst_pe_1_5_1_n61), .B2(
        npu_inst_pe_1_5_1_n40), .A(npu_inst_pe_1_5_1_n62), .ZN(
        npu_inst_pe_1_5_1_n86) );
  AND2_X1 npu_inst_pe_1_5_1_U63 ( .A1(npu_inst_pe_1_5_1_N93), .A2(npu_inst_n55), .ZN(npu_inst_int_data_y_5__1__0_) );
  AND2_X1 npu_inst_pe_1_5_1_U62 ( .A1(npu_inst_n55), .A2(npu_inst_pe_1_5_1_N94), .ZN(npu_inst_int_data_y_5__1__1_) );
  NOR3_X1 npu_inst_pe_1_5_1_U61 ( .A1(npu_inst_pe_1_5_1_n26), .A2(npu_inst_n55), .A3(npu_inst_int_ckg[22]), .ZN(npu_inst_pe_1_5_1_n85) );
  OR2_X1 npu_inst_pe_1_5_1_U60 ( .A1(npu_inst_pe_1_5_1_n85), .A2(
        npu_inst_pe_1_5_1_n2), .ZN(npu_inst_pe_1_5_1_N84) );
  AND2_X1 npu_inst_pe_1_5_1_U59 ( .A1(npu_inst_pe_1_5_1_int_q_acc_0_), .A2(
        npu_inst_pe_1_5_1_n1), .ZN(npu_inst_int_data_res_5__1__0_) );
  AND2_X1 npu_inst_pe_1_5_1_U58 ( .A1(npu_inst_pe_1_5_1_n2), .A2(
        npu_inst_pe_1_5_1_int_q_acc_7_), .ZN(npu_inst_int_data_res_5__1__7_)
         );
  AND2_X1 npu_inst_pe_1_5_1_U57 ( .A1(npu_inst_pe_1_5_1_int_q_acc_1_), .A2(
        npu_inst_pe_1_5_1_n1), .ZN(npu_inst_int_data_res_5__1__1_) );
  AND2_X1 npu_inst_pe_1_5_1_U56 ( .A1(npu_inst_pe_1_5_1_int_q_acc_2_), .A2(
        npu_inst_pe_1_5_1_n1), .ZN(npu_inst_int_data_res_5__1__2_) );
  AND2_X1 npu_inst_pe_1_5_1_U55 ( .A1(npu_inst_pe_1_5_1_int_q_acc_3_), .A2(
        npu_inst_pe_1_5_1_n2), .ZN(npu_inst_int_data_res_5__1__3_) );
  AND2_X1 npu_inst_pe_1_5_1_U54 ( .A1(npu_inst_pe_1_5_1_int_q_acc_4_), .A2(
        npu_inst_pe_1_5_1_n2), .ZN(npu_inst_int_data_res_5__1__4_) );
  AND2_X1 npu_inst_pe_1_5_1_U53 ( .A1(npu_inst_pe_1_5_1_int_q_acc_5_), .A2(
        npu_inst_pe_1_5_1_n2), .ZN(npu_inst_int_data_res_5__1__5_) );
  AND2_X1 npu_inst_pe_1_5_1_U52 ( .A1(npu_inst_pe_1_5_1_int_q_acc_6_), .A2(
        npu_inst_pe_1_5_1_n2), .ZN(npu_inst_int_data_res_5__1__6_) );
  AOI222_X1 npu_inst_pe_1_5_1_U51 ( .A1(npu_inst_int_data_res_6__1__0_), .A2(
        npu_inst_pe_1_5_1_n1), .B1(npu_inst_pe_1_5_1_N73), .B2(
        npu_inst_pe_1_5_1_n76), .C1(npu_inst_pe_1_5_1_N65), .C2(
        npu_inst_pe_1_5_1_n77), .ZN(npu_inst_pe_1_5_1_n84) );
  INV_X1 npu_inst_pe_1_5_1_U50 ( .A(npu_inst_pe_1_5_1_n84), .ZN(
        npu_inst_pe_1_5_1_n101) );
  AOI222_X1 npu_inst_pe_1_5_1_U49 ( .A1(npu_inst_int_data_res_6__1__7_), .A2(
        npu_inst_pe_1_5_1_n1), .B1(npu_inst_pe_1_5_1_N80), .B2(
        npu_inst_pe_1_5_1_n76), .C1(npu_inst_pe_1_5_1_N72), .C2(
        npu_inst_pe_1_5_1_n77), .ZN(npu_inst_pe_1_5_1_n75) );
  INV_X1 npu_inst_pe_1_5_1_U48 ( .A(npu_inst_pe_1_5_1_n75), .ZN(
        npu_inst_pe_1_5_1_n33) );
  AOI222_X1 npu_inst_pe_1_5_1_U47 ( .A1(npu_inst_int_data_res_6__1__1_), .A2(
        npu_inst_pe_1_5_1_n1), .B1(npu_inst_pe_1_5_1_N74), .B2(
        npu_inst_pe_1_5_1_n76), .C1(npu_inst_pe_1_5_1_N66), .C2(
        npu_inst_pe_1_5_1_n77), .ZN(npu_inst_pe_1_5_1_n83) );
  INV_X1 npu_inst_pe_1_5_1_U46 ( .A(npu_inst_pe_1_5_1_n83), .ZN(
        npu_inst_pe_1_5_1_n100) );
  AOI222_X1 npu_inst_pe_1_5_1_U45 ( .A1(npu_inst_int_data_res_6__1__2_), .A2(
        npu_inst_pe_1_5_1_n1), .B1(npu_inst_pe_1_5_1_N75), .B2(
        npu_inst_pe_1_5_1_n76), .C1(npu_inst_pe_1_5_1_N67), .C2(
        npu_inst_pe_1_5_1_n77), .ZN(npu_inst_pe_1_5_1_n82) );
  INV_X1 npu_inst_pe_1_5_1_U44 ( .A(npu_inst_pe_1_5_1_n82), .ZN(
        npu_inst_pe_1_5_1_n99) );
  AOI222_X1 npu_inst_pe_1_5_1_U43 ( .A1(npu_inst_int_data_res_6__1__3_), .A2(
        npu_inst_pe_1_5_1_n1), .B1(npu_inst_pe_1_5_1_N76), .B2(
        npu_inst_pe_1_5_1_n76), .C1(npu_inst_pe_1_5_1_N68), .C2(
        npu_inst_pe_1_5_1_n77), .ZN(npu_inst_pe_1_5_1_n81) );
  INV_X1 npu_inst_pe_1_5_1_U42 ( .A(npu_inst_pe_1_5_1_n81), .ZN(
        npu_inst_pe_1_5_1_n98) );
  AOI222_X1 npu_inst_pe_1_5_1_U41 ( .A1(npu_inst_int_data_res_6__1__4_), .A2(
        npu_inst_pe_1_5_1_n1), .B1(npu_inst_pe_1_5_1_N77), .B2(
        npu_inst_pe_1_5_1_n76), .C1(npu_inst_pe_1_5_1_N69), .C2(
        npu_inst_pe_1_5_1_n77), .ZN(npu_inst_pe_1_5_1_n80) );
  INV_X1 npu_inst_pe_1_5_1_U40 ( .A(npu_inst_pe_1_5_1_n80), .ZN(
        npu_inst_pe_1_5_1_n36) );
  AOI222_X1 npu_inst_pe_1_5_1_U39 ( .A1(npu_inst_int_data_res_6__1__5_), .A2(
        npu_inst_pe_1_5_1_n1), .B1(npu_inst_pe_1_5_1_N78), .B2(
        npu_inst_pe_1_5_1_n76), .C1(npu_inst_pe_1_5_1_N70), .C2(
        npu_inst_pe_1_5_1_n77), .ZN(npu_inst_pe_1_5_1_n79) );
  INV_X1 npu_inst_pe_1_5_1_U38 ( .A(npu_inst_pe_1_5_1_n79), .ZN(
        npu_inst_pe_1_5_1_n35) );
  AOI222_X1 npu_inst_pe_1_5_1_U37 ( .A1(npu_inst_int_data_res_6__1__6_), .A2(
        npu_inst_pe_1_5_1_n1), .B1(npu_inst_pe_1_5_1_N79), .B2(
        npu_inst_pe_1_5_1_n76), .C1(npu_inst_pe_1_5_1_N71), .C2(
        npu_inst_pe_1_5_1_n77), .ZN(npu_inst_pe_1_5_1_n78) );
  INV_X1 npu_inst_pe_1_5_1_U36 ( .A(npu_inst_pe_1_5_1_n78), .ZN(
        npu_inst_pe_1_5_1_n34) );
  INV_X1 npu_inst_pe_1_5_1_U35 ( .A(npu_inst_pe_1_5_1_int_data_1_), .ZN(
        npu_inst_pe_1_5_1_n14) );
  AND2_X1 npu_inst_pe_1_5_1_U34 ( .A1(npu_inst_int_data_x_5__1__1_), .A2(
        npu_inst_pe_1_5_1_int_q_weight_1_), .ZN(npu_inst_pe_1_5_1_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_5_1_U33 ( .A1(npu_inst_int_data_x_5__1__0_), .A2(
        npu_inst_pe_1_5_1_int_q_weight_1_), .ZN(npu_inst_pe_1_5_1_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_5_1_U32 ( .A1(npu_inst_n55), .A2(
        npu_inst_int_data_y_6__1__1_), .B1(npu_inst_pe_1_5_1_n3), .B2(
        npu_inst_int_data_x_5__2__1_), .ZN(npu_inst_pe_1_5_1_n63) );
  AOI22_X1 npu_inst_pe_1_5_1_U31 ( .A1(npu_inst_n55), .A2(
        npu_inst_int_data_y_6__1__0_), .B1(npu_inst_pe_1_5_1_n3), .B2(
        npu_inst_int_data_x_5__2__0_), .ZN(npu_inst_pe_1_5_1_n61) );
  INV_X1 npu_inst_pe_1_5_1_U30 ( .A(npu_inst_pe_1_5_1_int_data_0_), .ZN(
        npu_inst_pe_1_5_1_n13) );
  INV_X1 npu_inst_pe_1_5_1_U29 ( .A(npu_inst_n68), .ZN(npu_inst_pe_1_5_1_n5)
         );
  OR3_X1 npu_inst_pe_1_5_1_U28 ( .A1(npu_inst_pe_1_5_1_n6), .A2(
        npu_inst_pe_1_5_1_n8), .A3(npu_inst_pe_1_5_1_n5), .ZN(
        npu_inst_pe_1_5_1_n56) );
  OR3_X1 npu_inst_pe_1_5_1_U27 ( .A1(npu_inst_pe_1_5_1_n5), .A2(
        npu_inst_pe_1_5_1_n8), .A3(npu_inst_pe_1_5_1_n7), .ZN(
        npu_inst_pe_1_5_1_n48) );
  INV_X1 npu_inst_pe_1_5_1_U26 ( .A(npu_inst_pe_1_5_1_n5), .ZN(
        npu_inst_pe_1_5_1_n4) );
  OR3_X1 npu_inst_pe_1_5_1_U25 ( .A1(npu_inst_pe_1_5_1_n4), .A2(
        npu_inst_pe_1_5_1_n8), .A3(npu_inst_pe_1_5_1_n7), .ZN(
        npu_inst_pe_1_5_1_n52) );
  OR3_X1 npu_inst_pe_1_5_1_U24 ( .A1(npu_inst_pe_1_5_1_n6), .A2(
        npu_inst_pe_1_5_1_n8), .A3(npu_inst_pe_1_5_1_n4), .ZN(
        npu_inst_pe_1_5_1_n60) );
  NOR2_X1 npu_inst_pe_1_5_1_U23 ( .A1(npu_inst_pe_1_5_1_n60), .A2(
        npu_inst_pe_1_5_1_n3), .ZN(npu_inst_pe_1_5_1_n58) );
  NOR2_X1 npu_inst_pe_1_5_1_U22 ( .A1(npu_inst_pe_1_5_1_n56), .A2(
        npu_inst_pe_1_5_1_n3), .ZN(npu_inst_pe_1_5_1_n54) );
  NOR2_X1 npu_inst_pe_1_5_1_U21 ( .A1(npu_inst_pe_1_5_1_n52), .A2(
        npu_inst_pe_1_5_1_n3), .ZN(npu_inst_pe_1_5_1_n50) );
  NOR2_X1 npu_inst_pe_1_5_1_U20 ( .A1(npu_inst_pe_1_5_1_n48), .A2(
        npu_inst_pe_1_5_1_n3), .ZN(npu_inst_pe_1_5_1_n46) );
  NOR2_X1 npu_inst_pe_1_5_1_U19 ( .A1(npu_inst_pe_1_5_1_n40), .A2(
        npu_inst_pe_1_5_1_n3), .ZN(npu_inst_pe_1_5_1_n38) );
  NOR2_X1 npu_inst_pe_1_5_1_U18 ( .A1(npu_inst_pe_1_5_1_n44), .A2(
        npu_inst_pe_1_5_1_n3), .ZN(npu_inst_pe_1_5_1_n42) );
  BUF_X1 npu_inst_pe_1_5_1_U17 ( .A(npu_inst_n97), .Z(npu_inst_pe_1_5_1_n8) );
  INV_X1 npu_inst_pe_1_5_1_U16 ( .A(npu_inst_n123), .ZN(npu_inst_pe_1_5_1_n12)
         );
  INV_X1 npu_inst_pe_1_5_1_U15 ( .A(npu_inst_pe_1_5_1_n38), .ZN(
        npu_inst_pe_1_5_1_n114) );
  INV_X1 npu_inst_pe_1_5_1_U14 ( .A(npu_inst_pe_1_5_1_n58), .ZN(
        npu_inst_pe_1_5_1_n119) );
  INV_X1 npu_inst_pe_1_5_1_U13 ( .A(npu_inst_pe_1_5_1_n54), .ZN(
        npu_inst_pe_1_5_1_n118) );
  INV_X1 npu_inst_pe_1_5_1_U12 ( .A(npu_inst_pe_1_5_1_n50), .ZN(
        npu_inst_pe_1_5_1_n117) );
  INV_X1 npu_inst_pe_1_5_1_U11 ( .A(npu_inst_pe_1_5_1_n46), .ZN(
        npu_inst_pe_1_5_1_n116) );
  INV_X1 npu_inst_pe_1_5_1_U10 ( .A(npu_inst_pe_1_5_1_n42), .ZN(
        npu_inst_pe_1_5_1_n115) );
  BUF_X1 npu_inst_pe_1_5_1_U9 ( .A(npu_inst_n18), .Z(npu_inst_pe_1_5_1_n2) );
  BUF_X1 npu_inst_pe_1_5_1_U8 ( .A(npu_inst_n18), .Z(npu_inst_pe_1_5_1_n1) );
  BUF_X1 npu_inst_pe_1_5_1_U7 ( .A(npu_inst_pe_1_5_1_n12), .Z(
        npu_inst_pe_1_5_1_n11) );
  BUF_X1 npu_inst_pe_1_5_1_U6 ( .A(npu_inst_pe_1_5_1_n12), .Z(
        npu_inst_pe_1_5_1_n10) );
  BUF_X1 npu_inst_pe_1_5_1_U5 ( .A(npu_inst_pe_1_5_1_n12), .Z(
        npu_inst_pe_1_5_1_n9) );
  NOR2_X1 npu_inst_pe_1_5_1_U4 ( .A1(npu_inst_pe_1_5_1_int_q_weight_0_), .A2(
        npu_inst_pe_1_5_1_n1), .ZN(npu_inst_pe_1_5_1_n76) );
  NOR2_X1 npu_inst_pe_1_5_1_U3 ( .A1(npu_inst_pe_1_5_1_n27), .A2(
        npu_inst_pe_1_5_1_n1), .ZN(npu_inst_pe_1_5_1_n77) );
  FA_X1 npu_inst_pe_1_5_1_sub_67_U2_1 ( .A(npu_inst_pe_1_5_1_int_q_acc_1_), 
        .B(npu_inst_pe_1_5_1_n14), .CI(npu_inst_pe_1_5_1_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_5_1_sub_67_carry_2_), .S(npu_inst_pe_1_5_1_N66) );
  FA_X1 npu_inst_pe_1_5_1_add_69_U1_1 ( .A(npu_inst_pe_1_5_1_int_q_acc_1_), 
        .B(npu_inst_pe_1_5_1_int_data_1_), .CI(
        npu_inst_pe_1_5_1_add_69_carry_1_), .CO(
        npu_inst_pe_1_5_1_add_69_carry_2_), .S(npu_inst_pe_1_5_1_N74) );
  NAND3_X1 npu_inst_pe_1_5_1_U109 ( .A1(npu_inst_pe_1_5_1_n5), .A2(
        npu_inst_pe_1_5_1_n7), .A3(npu_inst_pe_1_5_1_n8), .ZN(
        npu_inst_pe_1_5_1_n44) );
  NAND3_X1 npu_inst_pe_1_5_1_U108 ( .A1(npu_inst_pe_1_5_1_n4), .A2(
        npu_inst_pe_1_5_1_n7), .A3(npu_inst_pe_1_5_1_n8), .ZN(
        npu_inst_pe_1_5_1_n40) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_5_1_n34), .CK(
        npu_inst_pe_1_5_1_net3619), .RN(npu_inst_pe_1_5_1_n9), .Q(
        npu_inst_pe_1_5_1_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_5_1_n35), .CK(
        npu_inst_pe_1_5_1_net3619), .RN(npu_inst_pe_1_5_1_n9), .Q(
        npu_inst_pe_1_5_1_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_5_1_n36), .CK(
        npu_inst_pe_1_5_1_net3619), .RN(npu_inst_pe_1_5_1_n9), .Q(
        npu_inst_pe_1_5_1_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_5_1_n98), .CK(
        npu_inst_pe_1_5_1_net3619), .RN(npu_inst_pe_1_5_1_n9), .Q(
        npu_inst_pe_1_5_1_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_5_1_n99), .CK(
        npu_inst_pe_1_5_1_net3619), .RN(npu_inst_pe_1_5_1_n9), .Q(
        npu_inst_pe_1_5_1_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_5_1_n100), 
        .CK(npu_inst_pe_1_5_1_net3619), .RN(npu_inst_pe_1_5_1_n9), .Q(
        npu_inst_pe_1_5_1_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_5_1_n33), .CK(
        npu_inst_pe_1_5_1_net3619), .RN(npu_inst_pe_1_5_1_n9), .Q(
        npu_inst_pe_1_5_1_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_5_1_n101), 
        .CK(npu_inst_pe_1_5_1_net3619), .RN(npu_inst_pe_1_5_1_n9), .Q(
        npu_inst_pe_1_5_1_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_weight_reg_0_ ( .D(npu_inst_n109), .CK(
        npu_inst_pe_1_5_1_net3625), .RN(npu_inst_pe_1_5_1_n9), .Q(
        npu_inst_pe_1_5_1_int_q_weight_0_), .QN(npu_inst_pe_1_5_1_n27) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_weight_reg_1_ ( .D(npu_inst_n115), .CK(
        npu_inst_pe_1_5_1_net3625), .RN(npu_inst_pe_1_5_1_n9), .Q(
        npu_inst_pe_1_5_1_int_q_weight_1_), .QN(npu_inst_pe_1_5_1_n26) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_5_1_n113), 
        .CK(npu_inst_pe_1_5_1_net3625), .RN(npu_inst_pe_1_5_1_n9), .Q(
        npu_inst_pe_1_5_1_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_5_1_n107), 
        .CK(npu_inst_pe_1_5_1_net3625), .RN(npu_inst_pe_1_5_1_n9), .Q(
        npu_inst_pe_1_5_1_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_5_1_n112), 
        .CK(npu_inst_pe_1_5_1_net3625), .RN(npu_inst_pe_1_5_1_n10), .Q(
        npu_inst_pe_1_5_1_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_5_1_n106), 
        .CK(npu_inst_pe_1_5_1_net3625), .RN(npu_inst_pe_1_5_1_n10), .Q(
        npu_inst_pe_1_5_1_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_5_1_n111), 
        .CK(npu_inst_pe_1_5_1_net3625), .RN(npu_inst_pe_1_5_1_n10), .Q(
        npu_inst_pe_1_5_1_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_5_1_n105), 
        .CK(npu_inst_pe_1_5_1_net3625), .RN(npu_inst_pe_1_5_1_n10), .Q(
        npu_inst_pe_1_5_1_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_5_1_n110), 
        .CK(npu_inst_pe_1_5_1_net3625), .RN(npu_inst_pe_1_5_1_n10), .Q(
        npu_inst_pe_1_5_1_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_5_1_n104), 
        .CK(npu_inst_pe_1_5_1_net3625), .RN(npu_inst_pe_1_5_1_n10), .Q(
        npu_inst_pe_1_5_1_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_5_1_n109), 
        .CK(npu_inst_pe_1_5_1_net3625), .RN(npu_inst_pe_1_5_1_n10), .Q(
        npu_inst_pe_1_5_1_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_5_1_n103), 
        .CK(npu_inst_pe_1_5_1_net3625), .RN(npu_inst_pe_1_5_1_n10), .Q(
        npu_inst_pe_1_5_1_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_5_1_n108), 
        .CK(npu_inst_pe_1_5_1_net3625), .RN(npu_inst_pe_1_5_1_n10), .Q(
        npu_inst_pe_1_5_1_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_5_1_n102), 
        .CK(npu_inst_pe_1_5_1_net3625), .RN(npu_inst_pe_1_5_1_n10), .Q(
        npu_inst_pe_1_5_1_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_5_1_n86), 
        .CK(npu_inst_pe_1_5_1_net3625), .RN(npu_inst_pe_1_5_1_n10), .Q(
        npu_inst_pe_1_5_1_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_5_1_n87), 
        .CK(npu_inst_pe_1_5_1_net3625), .RN(npu_inst_pe_1_5_1_n10), .Q(
        npu_inst_pe_1_5_1_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_5_1_n88), 
        .CK(npu_inst_pe_1_5_1_net3625), .RN(npu_inst_pe_1_5_1_n11), .Q(
        npu_inst_pe_1_5_1_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_5_1_n89), 
        .CK(npu_inst_pe_1_5_1_net3625), .RN(npu_inst_pe_1_5_1_n11), .Q(
        npu_inst_pe_1_5_1_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_5_1_n90), 
        .CK(npu_inst_pe_1_5_1_net3625), .RN(npu_inst_pe_1_5_1_n11), .Q(
        npu_inst_pe_1_5_1_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_5_1_n91), 
        .CK(npu_inst_pe_1_5_1_net3625), .RN(npu_inst_pe_1_5_1_n11), .Q(
        npu_inst_pe_1_5_1_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_5_1_n92), 
        .CK(npu_inst_pe_1_5_1_net3625), .RN(npu_inst_pe_1_5_1_n11), .Q(
        npu_inst_pe_1_5_1_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_5_1_n93), 
        .CK(npu_inst_pe_1_5_1_net3625), .RN(npu_inst_pe_1_5_1_n11), .Q(
        npu_inst_pe_1_5_1_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_5_1_n94), 
        .CK(npu_inst_pe_1_5_1_net3625), .RN(npu_inst_pe_1_5_1_n11), .Q(
        npu_inst_pe_1_5_1_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_5_1_n95), 
        .CK(npu_inst_pe_1_5_1_net3625), .RN(npu_inst_pe_1_5_1_n11), .Q(
        npu_inst_pe_1_5_1_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_5_1_n96), 
        .CK(npu_inst_pe_1_5_1_net3625), .RN(npu_inst_pe_1_5_1_n11), .Q(
        npu_inst_pe_1_5_1_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_5_1_n97), 
        .CK(npu_inst_pe_1_5_1_net3625), .RN(npu_inst_pe_1_5_1_n11), .Q(
        npu_inst_pe_1_5_1_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_5_1_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_5_1_N84), .SE(1'b0), .GCK(npu_inst_pe_1_5_1_net3619) );
  CLKGATETST_X1 npu_inst_pe_1_5_1_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n63), .SE(1'b0), .GCK(npu_inst_pe_1_5_1_net3625) );
  MUX2_X1 npu_inst_pe_1_5_2_U162 ( .A(npu_inst_pe_1_5_2_n32), .B(
        npu_inst_pe_1_5_2_n29), .S(npu_inst_pe_1_5_2_n8), .Z(
        npu_inst_pe_1_5_2_N93) );
  MUX2_X1 npu_inst_pe_1_5_2_U161 ( .A(npu_inst_pe_1_5_2_n31), .B(
        npu_inst_pe_1_5_2_n30), .S(npu_inst_pe_1_5_2_n6), .Z(
        npu_inst_pe_1_5_2_n32) );
  MUX2_X1 npu_inst_pe_1_5_2_U160 ( .A(npu_inst_pe_1_5_2_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_5_2_int_q_reg_v_1__0_), .S(npu_inst_pe_1_5_2_n4), .Z(
        npu_inst_pe_1_5_2_n31) );
  MUX2_X1 npu_inst_pe_1_5_2_U159 ( .A(npu_inst_pe_1_5_2_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_5_2_int_q_reg_v_3__0_), .S(npu_inst_pe_1_5_2_n4), .Z(
        npu_inst_pe_1_5_2_n30) );
  MUX2_X1 npu_inst_pe_1_5_2_U158 ( .A(npu_inst_pe_1_5_2_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_5_2_int_q_reg_v_5__0_), .S(npu_inst_pe_1_5_2_n4), .Z(
        npu_inst_pe_1_5_2_n29) );
  MUX2_X1 npu_inst_pe_1_5_2_U157 ( .A(npu_inst_pe_1_5_2_n28), .B(
        npu_inst_pe_1_5_2_n23), .S(npu_inst_pe_1_5_2_n8), .Z(
        npu_inst_pe_1_5_2_N94) );
  MUX2_X1 npu_inst_pe_1_5_2_U156 ( .A(npu_inst_pe_1_5_2_n25), .B(
        npu_inst_pe_1_5_2_n24), .S(npu_inst_pe_1_5_2_n6), .Z(
        npu_inst_pe_1_5_2_n28) );
  MUX2_X1 npu_inst_pe_1_5_2_U155 ( .A(npu_inst_pe_1_5_2_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_5_2_int_q_reg_v_1__1_), .S(npu_inst_pe_1_5_2_n4), .Z(
        npu_inst_pe_1_5_2_n25) );
  MUX2_X1 npu_inst_pe_1_5_2_U154 ( .A(npu_inst_pe_1_5_2_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_5_2_int_q_reg_v_3__1_), .S(npu_inst_pe_1_5_2_n4), .Z(
        npu_inst_pe_1_5_2_n24) );
  MUX2_X1 npu_inst_pe_1_5_2_U153 ( .A(npu_inst_pe_1_5_2_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_5_2_int_q_reg_v_5__1_), .S(npu_inst_pe_1_5_2_n4), .Z(
        npu_inst_pe_1_5_2_n23) );
  MUX2_X1 npu_inst_pe_1_5_2_U152 ( .A(npu_inst_pe_1_5_2_n22), .B(
        npu_inst_pe_1_5_2_n19), .S(npu_inst_pe_1_5_2_n8), .Z(
        npu_inst_int_data_x_5__2__1_) );
  MUX2_X1 npu_inst_pe_1_5_2_U151 ( .A(npu_inst_pe_1_5_2_n21), .B(
        npu_inst_pe_1_5_2_n20), .S(npu_inst_pe_1_5_2_n6), .Z(
        npu_inst_pe_1_5_2_n22) );
  MUX2_X1 npu_inst_pe_1_5_2_U150 ( .A(npu_inst_pe_1_5_2_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_5_2_int_q_reg_h_1__1_), .S(npu_inst_pe_1_5_2_n4), .Z(
        npu_inst_pe_1_5_2_n21) );
  MUX2_X1 npu_inst_pe_1_5_2_U149 ( .A(npu_inst_pe_1_5_2_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_5_2_int_q_reg_h_3__1_), .S(npu_inst_pe_1_5_2_n4), .Z(
        npu_inst_pe_1_5_2_n20) );
  MUX2_X1 npu_inst_pe_1_5_2_U148 ( .A(npu_inst_pe_1_5_2_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_5_2_int_q_reg_h_5__1_), .S(npu_inst_pe_1_5_2_n4), .Z(
        npu_inst_pe_1_5_2_n19) );
  MUX2_X1 npu_inst_pe_1_5_2_U147 ( .A(npu_inst_pe_1_5_2_n18), .B(
        npu_inst_pe_1_5_2_n15), .S(npu_inst_pe_1_5_2_n8), .Z(
        npu_inst_int_data_x_5__2__0_) );
  MUX2_X1 npu_inst_pe_1_5_2_U146 ( .A(npu_inst_pe_1_5_2_n17), .B(
        npu_inst_pe_1_5_2_n16), .S(npu_inst_pe_1_5_2_n6), .Z(
        npu_inst_pe_1_5_2_n18) );
  MUX2_X1 npu_inst_pe_1_5_2_U145 ( .A(npu_inst_pe_1_5_2_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_5_2_int_q_reg_h_1__0_), .S(npu_inst_pe_1_5_2_n4), .Z(
        npu_inst_pe_1_5_2_n17) );
  MUX2_X1 npu_inst_pe_1_5_2_U144 ( .A(npu_inst_pe_1_5_2_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_5_2_int_q_reg_h_3__0_), .S(npu_inst_pe_1_5_2_n4), .Z(
        npu_inst_pe_1_5_2_n16) );
  MUX2_X1 npu_inst_pe_1_5_2_U143 ( .A(npu_inst_pe_1_5_2_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_5_2_int_q_reg_h_5__0_), .S(npu_inst_pe_1_5_2_n4), .Z(
        npu_inst_pe_1_5_2_n15) );
  XOR2_X1 npu_inst_pe_1_5_2_U142 ( .A(npu_inst_pe_1_5_2_int_data_0_), .B(
        npu_inst_pe_1_5_2_int_q_acc_0_), .Z(npu_inst_pe_1_5_2_N73) );
  AND2_X1 npu_inst_pe_1_5_2_U141 ( .A1(npu_inst_pe_1_5_2_int_q_acc_0_), .A2(
        npu_inst_pe_1_5_2_int_data_0_), .ZN(npu_inst_pe_1_5_2_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_5_2_U140 ( .A(npu_inst_pe_1_5_2_int_q_acc_0_), .B(
        npu_inst_pe_1_5_2_n13), .ZN(npu_inst_pe_1_5_2_N65) );
  OR2_X1 npu_inst_pe_1_5_2_U139 ( .A1(npu_inst_pe_1_5_2_n13), .A2(
        npu_inst_pe_1_5_2_int_q_acc_0_), .ZN(npu_inst_pe_1_5_2_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_5_2_U138 ( .A(npu_inst_pe_1_5_2_int_q_acc_2_), .B(
        npu_inst_pe_1_5_2_add_69_carry_2_), .Z(npu_inst_pe_1_5_2_N75) );
  AND2_X1 npu_inst_pe_1_5_2_U137 ( .A1(npu_inst_pe_1_5_2_add_69_carry_2_), 
        .A2(npu_inst_pe_1_5_2_int_q_acc_2_), .ZN(
        npu_inst_pe_1_5_2_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_5_2_U136 ( .A(npu_inst_pe_1_5_2_int_q_acc_3_), .B(
        npu_inst_pe_1_5_2_add_69_carry_3_), .Z(npu_inst_pe_1_5_2_N76) );
  AND2_X1 npu_inst_pe_1_5_2_U135 ( .A1(npu_inst_pe_1_5_2_add_69_carry_3_), 
        .A2(npu_inst_pe_1_5_2_int_q_acc_3_), .ZN(
        npu_inst_pe_1_5_2_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_5_2_U134 ( .A(npu_inst_pe_1_5_2_int_q_acc_4_), .B(
        npu_inst_pe_1_5_2_add_69_carry_4_), .Z(npu_inst_pe_1_5_2_N77) );
  AND2_X1 npu_inst_pe_1_5_2_U133 ( .A1(npu_inst_pe_1_5_2_add_69_carry_4_), 
        .A2(npu_inst_pe_1_5_2_int_q_acc_4_), .ZN(
        npu_inst_pe_1_5_2_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_5_2_U132 ( .A(npu_inst_pe_1_5_2_int_q_acc_5_), .B(
        npu_inst_pe_1_5_2_add_69_carry_5_), .Z(npu_inst_pe_1_5_2_N78) );
  AND2_X1 npu_inst_pe_1_5_2_U131 ( .A1(npu_inst_pe_1_5_2_add_69_carry_5_), 
        .A2(npu_inst_pe_1_5_2_int_q_acc_5_), .ZN(
        npu_inst_pe_1_5_2_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_5_2_U130 ( .A(npu_inst_pe_1_5_2_int_q_acc_6_), .B(
        npu_inst_pe_1_5_2_add_69_carry_6_), .Z(npu_inst_pe_1_5_2_N79) );
  AND2_X1 npu_inst_pe_1_5_2_U129 ( .A1(npu_inst_pe_1_5_2_add_69_carry_6_), 
        .A2(npu_inst_pe_1_5_2_int_q_acc_6_), .ZN(
        npu_inst_pe_1_5_2_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_5_2_U128 ( .A(npu_inst_pe_1_5_2_int_q_acc_7_), .B(
        npu_inst_pe_1_5_2_add_69_carry_7_), .Z(npu_inst_pe_1_5_2_N80) );
  XNOR2_X1 npu_inst_pe_1_5_2_U127 ( .A(npu_inst_pe_1_5_2_sub_67_carry_2_), .B(
        npu_inst_pe_1_5_2_int_q_acc_2_), .ZN(npu_inst_pe_1_5_2_N67) );
  OR2_X1 npu_inst_pe_1_5_2_U126 ( .A1(npu_inst_pe_1_5_2_int_q_acc_2_), .A2(
        npu_inst_pe_1_5_2_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_5_2_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_5_2_U125 ( .A(npu_inst_pe_1_5_2_sub_67_carry_3_), .B(
        npu_inst_pe_1_5_2_int_q_acc_3_), .ZN(npu_inst_pe_1_5_2_N68) );
  OR2_X1 npu_inst_pe_1_5_2_U124 ( .A1(npu_inst_pe_1_5_2_int_q_acc_3_), .A2(
        npu_inst_pe_1_5_2_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_5_2_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_5_2_U123 ( .A(npu_inst_pe_1_5_2_sub_67_carry_4_), .B(
        npu_inst_pe_1_5_2_int_q_acc_4_), .ZN(npu_inst_pe_1_5_2_N69) );
  OR2_X1 npu_inst_pe_1_5_2_U122 ( .A1(npu_inst_pe_1_5_2_int_q_acc_4_), .A2(
        npu_inst_pe_1_5_2_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_5_2_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_5_2_U121 ( .A(npu_inst_pe_1_5_2_sub_67_carry_5_), .B(
        npu_inst_pe_1_5_2_int_q_acc_5_), .ZN(npu_inst_pe_1_5_2_N70) );
  OR2_X1 npu_inst_pe_1_5_2_U120 ( .A1(npu_inst_pe_1_5_2_int_q_acc_5_), .A2(
        npu_inst_pe_1_5_2_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_5_2_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_5_2_U119 ( .A(npu_inst_pe_1_5_2_sub_67_carry_6_), .B(
        npu_inst_pe_1_5_2_int_q_acc_6_), .ZN(npu_inst_pe_1_5_2_N71) );
  OR2_X1 npu_inst_pe_1_5_2_U118 ( .A1(npu_inst_pe_1_5_2_int_q_acc_6_), .A2(
        npu_inst_pe_1_5_2_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_5_2_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_5_2_U117 ( .A(npu_inst_pe_1_5_2_int_q_acc_7_), .B(
        npu_inst_pe_1_5_2_sub_67_carry_7_), .ZN(npu_inst_pe_1_5_2_N72) );
  INV_X1 npu_inst_pe_1_5_2_U116 ( .A(npu_inst_n76), .ZN(npu_inst_pe_1_5_2_n7)
         );
  INV_X1 npu_inst_pe_1_5_2_U115 ( .A(npu_inst_pe_1_5_2_n7), .ZN(
        npu_inst_pe_1_5_2_n6) );
  INV_X1 npu_inst_pe_1_5_2_U114 ( .A(npu_inst_n55), .ZN(npu_inst_pe_1_5_2_n3)
         );
  AOI22_X1 npu_inst_pe_1_5_2_U113 ( .A1(npu_inst_int_data_y_6__2__0_), .A2(
        npu_inst_pe_1_5_2_n58), .B1(npu_inst_pe_1_5_2_n119), .B2(
        npu_inst_pe_1_5_2_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_5_2_n57) );
  INV_X1 npu_inst_pe_1_5_2_U112 ( .A(npu_inst_pe_1_5_2_n57), .ZN(
        npu_inst_pe_1_5_2_n108) );
  AOI22_X1 npu_inst_pe_1_5_2_U111 ( .A1(npu_inst_int_data_y_6__2__0_), .A2(
        npu_inst_pe_1_5_2_n54), .B1(npu_inst_pe_1_5_2_n118), .B2(
        npu_inst_pe_1_5_2_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_5_2_n53) );
  INV_X1 npu_inst_pe_1_5_2_U110 ( .A(npu_inst_pe_1_5_2_n53), .ZN(
        npu_inst_pe_1_5_2_n109) );
  AOI22_X1 npu_inst_pe_1_5_2_U107 ( .A1(npu_inst_int_data_y_6__2__0_), .A2(
        npu_inst_pe_1_5_2_n50), .B1(npu_inst_pe_1_5_2_n117), .B2(
        npu_inst_pe_1_5_2_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_5_2_n49) );
  INV_X1 npu_inst_pe_1_5_2_U106 ( .A(npu_inst_pe_1_5_2_n49), .ZN(
        npu_inst_pe_1_5_2_n110) );
  AOI22_X1 npu_inst_pe_1_5_2_U105 ( .A1(npu_inst_int_data_y_6__2__0_), .A2(
        npu_inst_pe_1_5_2_n46), .B1(npu_inst_pe_1_5_2_n116), .B2(
        npu_inst_pe_1_5_2_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_5_2_n45) );
  INV_X1 npu_inst_pe_1_5_2_U104 ( .A(npu_inst_pe_1_5_2_n45), .ZN(
        npu_inst_pe_1_5_2_n111) );
  AOI22_X1 npu_inst_pe_1_5_2_U103 ( .A1(npu_inst_int_data_y_6__2__0_), .A2(
        npu_inst_pe_1_5_2_n42), .B1(npu_inst_pe_1_5_2_n115), .B2(
        npu_inst_pe_1_5_2_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_5_2_n41) );
  INV_X1 npu_inst_pe_1_5_2_U102 ( .A(npu_inst_pe_1_5_2_n41), .ZN(
        npu_inst_pe_1_5_2_n112) );
  AOI22_X1 npu_inst_pe_1_5_2_U101 ( .A1(npu_inst_int_data_y_6__2__1_), .A2(
        npu_inst_pe_1_5_2_n58), .B1(npu_inst_pe_1_5_2_n119), .B2(
        npu_inst_pe_1_5_2_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_5_2_n59) );
  INV_X1 npu_inst_pe_1_5_2_U100 ( .A(npu_inst_pe_1_5_2_n59), .ZN(
        npu_inst_pe_1_5_2_n102) );
  AOI22_X1 npu_inst_pe_1_5_2_U99 ( .A1(npu_inst_int_data_y_6__2__1_), .A2(
        npu_inst_pe_1_5_2_n54), .B1(npu_inst_pe_1_5_2_n118), .B2(
        npu_inst_pe_1_5_2_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_5_2_n55) );
  INV_X1 npu_inst_pe_1_5_2_U98 ( .A(npu_inst_pe_1_5_2_n55), .ZN(
        npu_inst_pe_1_5_2_n103) );
  AOI22_X1 npu_inst_pe_1_5_2_U97 ( .A1(npu_inst_int_data_y_6__2__1_), .A2(
        npu_inst_pe_1_5_2_n50), .B1(npu_inst_pe_1_5_2_n117), .B2(
        npu_inst_pe_1_5_2_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_5_2_n51) );
  INV_X1 npu_inst_pe_1_5_2_U96 ( .A(npu_inst_pe_1_5_2_n51), .ZN(
        npu_inst_pe_1_5_2_n104) );
  AOI22_X1 npu_inst_pe_1_5_2_U95 ( .A1(npu_inst_int_data_y_6__2__1_), .A2(
        npu_inst_pe_1_5_2_n46), .B1(npu_inst_pe_1_5_2_n116), .B2(
        npu_inst_pe_1_5_2_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_5_2_n47) );
  INV_X1 npu_inst_pe_1_5_2_U94 ( .A(npu_inst_pe_1_5_2_n47), .ZN(
        npu_inst_pe_1_5_2_n105) );
  AOI22_X1 npu_inst_pe_1_5_2_U93 ( .A1(npu_inst_int_data_y_6__2__1_), .A2(
        npu_inst_pe_1_5_2_n42), .B1(npu_inst_pe_1_5_2_n115), .B2(
        npu_inst_pe_1_5_2_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_5_2_n43) );
  INV_X1 npu_inst_pe_1_5_2_U92 ( .A(npu_inst_pe_1_5_2_n43), .ZN(
        npu_inst_pe_1_5_2_n106) );
  AOI22_X1 npu_inst_pe_1_5_2_U91 ( .A1(npu_inst_pe_1_5_2_n38), .A2(
        npu_inst_int_data_y_6__2__1_), .B1(npu_inst_pe_1_5_2_n114), .B2(
        npu_inst_pe_1_5_2_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_5_2_n39) );
  INV_X1 npu_inst_pe_1_5_2_U90 ( .A(npu_inst_pe_1_5_2_n39), .ZN(
        npu_inst_pe_1_5_2_n107) );
  AOI22_X1 npu_inst_pe_1_5_2_U89 ( .A1(npu_inst_pe_1_5_2_n38), .A2(
        npu_inst_int_data_y_6__2__0_), .B1(npu_inst_pe_1_5_2_n114), .B2(
        npu_inst_pe_1_5_2_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_5_2_n37) );
  INV_X1 npu_inst_pe_1_5_2_U88 ( .A(npu_inst_pe_1_5_2_n37), .ZN(
        npu_inst_pe_1_5_2_n113) );
  NAND2_X1 npu_inst_pe_1_5_2_U87 ( .A1(npu_inst_pe_1_5_2_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_5_2_n60), .ZN(npu_inst_pe_1_5_2_n74) );
  OAI21_X1 npu_inst_pe_1_5_2_U86 ( .B1(npu_inst_pe_1_5_2_n63), .B2(
        npu_inst_pe_1_5_2_n60), .A(npu_inst_pe_1_5_2_n74), .ZN(
        npu_inst_pe_1_5_2_n97) );
  NAND2_X1 npu_inst_pe_1_5_2_U85 ( .A1(npu_inst_pe_1_5_2_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_5_2_n60), .ZN(npu_inst_pe_1_5_2_n73) );
  OAI21_X1 npu_inst_pe_1_5_2_U84 ( .B1(npu_inst_pe_1_5_2_n61), .B2(
        npu_inst_pe_1_5_2_n60), .A(npu_inst_pe_1_5_2_n73), .ZN(
        npu_inst_pe_1_5_2_n96) );
  NAND2_X1 npu_inst_pe_1_5_2_U83 ( .A1(npu_inst_pe_1_5_2_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_5_2_n56), .ZN(npu_inst_pe_1_5_2_n72) );
  OAI21_X1 npu_inst_pe_1_5_2_U82 ( .B1(npu_inst_pe_1_5_2_n63), .B2(
        npu_inst_pe_1_5_2_n56), .A(npu_inst_pe_1_5_2_n72), .ZN(
        npu_inst_pe_1_5_2_n95) );
  NAND2_X1 npu_inst_pe_1_5_2_U81 ( .A1(npu_inst_pe_1_5_2_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_5_2_n56), .ZN(npu_inst_pe_1_5_2_n71) );
  OAI21_X1 npu_inst_pe_1_5_2_U80 ( .B1(npu_inst_pe_1_5_2_n61), .B2(
        npu_inst_pe_1_5_2_n56), .A(npu_inst_pe_1_5_2_n71), .ZN(
        npu_inst_pe_1_5_2_n94) );
  NAND2_X1 npu_inst_pe_1_5_2_U79 ( .A1(npu_inst_pe_1_5_2_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_5_2_n52), .ZN(npu_inst_pe_1_5_2_n70) );
  OAI21_X1 npu_inst_pe_1_5_2_U78 ( .B1(npu_inst_pe_1_5_2_n63), .B2(
        npu_inst_pe_1_5_2_n52), .A(npu_inst_pe_1_5_2_n70), .ZN(
        npu_inst_pe_1_5_2_n93) );
  NAND2_X1 npu_inst_pe_1_5_2_U77 ( .A1(npu_inst_pe_1_5_2_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_5_2_n52), .ZN(npu_inst_pe_1_5_2_n69) );
  OAI21_X1 npu_inst_pe_1_5_2_U76 ( .B1(npu_inst_pe_1_5_2_n61), .B2(
        npu_inst_pe_1_5_2_n52), .A(npu_inst_pe_1_5_2_n69), .ZN(
        npu_inst_pe_1_5_2_n92) );
  NAND2_X1 npu_inst_pe_1_5_2_U75 ( .A1(npu_inst_pe_1_5_2_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_5_2_n48), .ZN(npu_inst_pe_1_5_2_n68) );
  OAI21_X1 npu_inst_pe_1_5_2_U74 ( .B1(npu_inst_pe_1_5_2_n63), .B2(
        npu_inst_pe_1_5_2_n48), .A(npu_inst_pe_1_5_2_n68), .ZN(
        npu_inst_pe_1_5_2_n91) );
  NAND2_X1 npu_inst_pe_1_5_2_U73 ( .A1(npu_inst_pe_1_5_2_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_5_2_n48), .ZN(npu_inst_pe_1_5_2_n67) );
  OAI21_X1 npu_inst_pe_1_5_2_U72 ( .B1(npu_inst_pe_1_5_2_n61), .B2(
        npu_inst_pe_1_5_2_n48), .A(npu_inst_pe_1_5_2_n67), .ZN(
        npu_inst_pe_1_5_2_n90) );
  NAND2_X1 npu_inst_pe_1_5_2_U71 ( .A1(npu_inst_pe_1_5_2_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_5_2_n44), .ZN(npu_inst_pe_1_5_2_n66) );
  OAI21_X1 npu_inst_pe_1_5_2_U70 ( .B1(npu_inst_pe_1_5_2_n63), .B2(
        npu_inst_pe_1_5_2_n44), .A(npu_inst_pe_1_5_2_n66), .ZN(
        npu_inst_pe_1_5_2_n89) );
  NAND2_X1 npu_inst_pe_1_5_2_U69 ( .A1(npu_inst_pe_1_5_2_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_5_2_n44), .ZN(npu_inst_pe_1_5_2_n65) );
  OAI21_X1 npu_inst_pe_1_5_2_U68 ( .B1(npu_inst_pe_1_5_2_n61), .B2(
        npu_inst_pe_1_5_2_n44), .A(npu_inst_pe_1_5_2_n65), .ZN(
        npu_inst_pe_1_5_2_n88) );
  NAND2_X1 npu_inst_pe_1_5_2_U67 ( .A1(npu_inst_pe_1_5_2_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_5_2_n40), .ZN(npu_inst_pe_1_5_2_n64) );
  OAI21_X1 npu_inst_pe_1_5_2_U66 ( .B1(npu_inst_pe_1_5_2_n63), .B2(
        npu_inst_pe_1_5_2_n40), .A(npu_inst_pe_1_5_2_n64), .ZN(
        npu_inst_pe_1_5_2_n87) );
  NAND2_X1 npu_inst_pe_1_5_2_U65 ( .A1(npu_inst_pe_1_5_2_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_5_2_n40), .ZN(npu_inst_pe_1_5_2_n62) );
  OAI21_X1 npu_inst_pe_1_5_2_U64 ( .B1(npu_inst_pe_1_5_2_n61), .B2(
        npu_inst_pe_1_5_2_n40), .A(npu_inst_pe_1_5_2_n62), .ZN(
        npu_inst_pe_1_5_2_n86) );
  AND2_X1 npu_inst_pe_1_5_2_U63 ( .A1(npu_inst_pe_1_5_2_N93), .A2(npu_inst_n55), .ZN(npu_inst_int_data_y_5__2__0_) );
  AND2_X1 npu_inst_pe_1_5_2_U62 ( .A1(npu_inst_n55), .A2(npu_inst_pe_1_5_2_N94), .ZN(npu_inst_int_data_y_5__2__1_) );
  NOR3_X1 npu_inst_pe_1_5_2_U61 ( .A1(npu_inst_pe_1_5_2_n26), .A2(npu_inst_n55), .A3(npu_inst_int_ckg[21]), .ZN(npu_inst_pe_1_5_2_n85) );
  OR2_X1 npu_inst_pe_1_5_2_U60 ( .A1(npu_inst_pe_1_5_2_n85), .A2(
        npu_inst_pe_1_5_2_n2), .ZN(npu_inst_pe_1_5_2_N84) );
  AND2_X1 npu_inst_pe_1_5_2_U59 ( .A1(npu_inst_pe_1_5_2_int_q_acc_0_), .A2(
        npu_inst_pe_1_5_2_n1), .ZN(npu_inst_int_data_res_5__2__0_) );
  AND2_X1 npu_inst_pe_1_5_2_U58 ( .A1(npu_inst_pe_1_5_2_n2), .A2(
        npu_inst_pe_1_5_2_int_q_acc_7_), .ZN(npu_inst_int_data_res_5__2__7_)
         );
  AND2_X1 npu_inst_pe_1_5_2_U57 ( .A1(npu_inst_pe_1_5_2_int_q_acc_1_), .A2(
        npu_inst_pe_1_5_2_n1), .ZN(npu_inst_int_data_res_5__2__1_) );
  AND2_X1 npu_inst_pe_1_5_2_U56 ( .A1(npu_inst_pe_1_5_2_int_q_acc_2_), .A2(
        npu_inst_pe_1_5_2_n1), .ZN(npu_inst_int_data_res_5__2__2_) );
  AND2_X1 npu_inst_pe_1_5_2_U55 ( .A1(npu_inst_pe_1_5_2_int_q_acc_3_), .A2(
        npu_inst_pe_1_5_2_n2), .ZN(npu_inst_int_data_res_5__2__3_) );
  AND2_X1 npu_inst_pe_1_5_2_U54 ( .A1(npu_inst_pe_1_5_2_int_q_acc_4_), .A2(
        npu_inst_pe_1_5_2_n2), .ZN(npu_inst_int_data_res_5__2__4_) );
  AND2_X1 npu_inst_pe_1_5_2_U53 ( .A1(npu_inst_pe_1_5_2_int_q_acc_5_), .A2(
        npu_inst_pe_1_5_2_n2), .ZN(npu_inst_int_data_res_5__2__5_) );
  AND2_X1 npu_inst_pe_1_5_2_U52 ( .A1(npu_inst_pe_1_5_2_int_q_acc_6_), .A2(
        npu_inst_pe_1_5_2_n2), .ZN(npu_inst_int_data_res_5__2__6_) );
  AOI222_X1 npu_inst_pe_1_5_2_U51 ( .A1(npu_inst_int_data_res_6__2__0_), .A2(
        npu_inst_pe_1_5_2_n1), .B1(npu_inst_pe_1_5_2_N73), .B2(
        npu_inst_pe_1_5_2_n76), .C1(npu_inst_pe_1_5_2_N65), .C2(
        npu_inst_pe_1_5_2_n77), .ZN(npu_inst_pe_1_5_2_n84) );
  INV_X1 npu_inst_pe_1_5_2_U50 ( .A(npu_inst_pe_1_5_2_n84), .ZN(
        npu_inst_pe_1_5_2_n101) );
  AOI222_X1 npu_inst_pe_1_5_2_U49 ( .A1(npu_inst_int_data_res_6__2__7_), .A2(
        npu_inst_pe_1_5_2_n1), .B1(npu_inst_pe_1_5_2_N80), .B2(
        npu_inst_pe_1_5_2_n76), .C1(npu_inst_pe_1_5_2_N72), .C2(
        npu_inst_pe_1_5_2_n77), .ZN(npu_inst_pe_1_5_2_n75) );
  INV_X1 npu_inst_pe_1_5_2_U48 ( .A(npu_inst_pe_1_5_2_n75), .ZN(
        npu_inst_pe_1_5_2_n33) );
  AOI222_X1 npu_inst_pe_1_5_2_U47 ( .A1(npu_inst_int_data_res_6__2__1_), .A2(
        npu_inst_pe_1_5_2_n1), .B1(npu_inst_pe_1_5_2_N74), .B2(
        npu_inst_pe_1_5_2_n76), .C1(npu_inst_pe_1_5_2_N66), .C2(
        npu_inst_pe_1_5_2_n77), .ZN(npu_inst_pe_1_5_2_n83) );
  INV_X1 npu_inst_pe_1_5_2_U46 ( .A(npu_inst_pe_1_5_2_n83), .ZN(
        npu_inst_pe_1_5_2_n100) );
  AOI222_X1 npu_inst_pe_1_5_2_U45 ( .A1(npu_inst_int_data_res_6__2__2_), .A2(
        npu_inst_pe_1_5_2_n1), .B1(npu_inst_pe_1_5_2_N75), .B2(
        npu_inst_pe_1_5_2_n76), .C1(npu_inst_pe_1_5_2_N67), .C2(
        npu_inst_pe_1_5_2_n77), .ZN(npu_inst_pe_1_5_2_n82) );
  INV_X1 npu_inst_pe_1_5_2_U44 ( .A(npu_inst_pe_1_5_2_n82), .ZN(
        npu_inst_pe_1_5_2_n99) );
  AOI222_X1 npu_inst_pe_1_5_2_U43 ( .A1(npu_inst_int_data_res_6__2__3_), .A2(
        npu_inst_pe_1_5_2_n1), .B1(npu_inst_pe_1_5_2_N76), .B2(
        npu_inst_pe_1_5_2_n76), .C1(npu_inst_pe_1_5_2_N68), .C2(
        npu_inst_pe_1_5_2_n77), .ZN(npu_inst_pe_1_5_2_n81) );
  INV_X1 npu_inst_pe_1_5_2_U42 ( .A(npu_inst_pe_1_5_2_n81), .ZN(
        npu_inst_pe_1_5_2_n98) );
  AOI222_X1 npu_inst_pe_1_5_2_U41 ( .A1(npu_inst_int_data_res_6__2__4_), .A2(
        npu_inst_pe_1_5_2_n1), .B1(npu_inst_pe_1_5_2_N77), .B2(
        npu_inst_pe_1_5_2_n76), .C1(npu_inst_pe_1_5_2_N69), .C2(
        npu_inst_pe_1_5_2_n77), .ZN(npu_inst_pe_1_5_2_n80) );
  INV_X1 npu_inst_pe_1_5_2_U40 ( .A(npu_inst_pe_1_5_2_n80), .ZN(
        npu_inst_pe_1_5_2_n36) );
  AOI222_X1 npu_inst_pe_1_5_2_U39 ( .A1(npu_inst_int_data_res_6__2__5_), .A2(
        npu_inst_pe_1_5_2_n1), .B1(npu_inst_pe_1_5_2_N78), .B2(
        npu_inst_pe_1_5_2_n76), .C1(npu_inst_pe_1_5_2_N70), .C2(
        npu_inst_pe_1_5_2_n77), .ZN(npu_inst_pe_1_5_2_n79) );
  INV_X1 npu_inst_pe_1_5_2_U38 ( .A(npu_inst_pe_1_5_2_n79), .ZN(
        npu_inst_pe_1_5_2_n35) );
  AOI222_X1 npu_inst_pe_1_5_2_U37 ( .A1(npu_inst_int_data_res_6__2__6_), .A2(
        npu_inst_pe_1_5_2_n1), .B1(npu_inst_pe_1_5_2_N79), .B2(
        npu_inst_pe_1_5_2_n76), .C1(npu_inst_pe_1_5_2_N71), .C2(
        npu_inst_pe_1_5_2_n77), .ZN(npu_inst_pe_1_5_2_n78) );
  INV_X1 npu_inst_pe_1_5_2_U36 ( .A(npu_inst_pe_1_5_2_n78), .ZN(
        npu_inst_pe_1_5_2_n34) );
  INV_X1 npu_inst_pe_1_5_2_U35 ( .A(npu_inst_pe_1_5_2_int_data_1_), .ZN(
        npu_inst_pe_1_5_2_n14) );
  AND2_X1 npu_inst_pe_1_5_2_U34 ( .A1(npu_inst_int_data_x_5__2__1_), .A2(
        npu_inst_pe_1_5_2_int_q_weight_1_), .ZN(npu_inst_pe_1_5_2_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_5_2_U33 ( .A1(npu_inst_int_data_x_5__2__0_), .A2(
        npu_inst_pe_1_5_2_int_q_weight_1_), .ZN(npu_inst_pe_1_5_2_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_5_2_U32 ( .A1(npu_inst_n55), .A2(
        npu_inst_int_data_y_6__2__1_), .B1(npu_inst_pe_1_5_2_n3), .B2(
        npu_inst_int_data_x_5__3__1_), .ZN(npu_inst_pe_1_5_2_n63) );
  AOI22_X1 npu_inst_pe_1_5_2_U31 ( .A1(npu_inst_n55), .A2(
        npu_inst_int_data_y_6__2__0_), .B1(npu_inst_pe_1_5_2_n3), .B2(
        npu_inst_int_data_x_5__3__0_), .ZN(npu_inst_pe_1_5_2_n61) );
  INV_X1 npu_inst_pe_1_5_2_U30 ( .A(npu_inst_pe_1_5_2_int_data_0_), .ZN(
        npu_inst_pe_1_5_2_n13) );
  INV_X1 npu_inst_pe_1_5_2_U29 ( .A(npu_inst_n68), .ZN(npu_inst_pe_1_5_2_n5)
         );
  OR3_X1 npu_inst_pe_1_5_2_U28 ( .A1(npu_inst_pe_1_5_2_n6), .A2(
        npu_inst_pe_1_5_2_n8), .A3(npu_inst_pe_1_5_2_n5), .ZN(
        npu_inst_pe_1_5_2_n56) );
  OR3_X1 npu_inst_pe_1_5_2_U27 ( .A1(npu_inst_pe_1_5_2_n5), .A2(
        npu_inst_pe_1_5_2_n8), .A3(npu_inst_pe_1_5_2_n7), .ZN(
        npu_inst_pe_1_5_2_n48) );
  INV_X1 npu_inst_pe_1_5_2_U26 ( .A(npu_inst_pe_1_5_2_n5), .ZN(
        npu_inst_pe_1_5_2_n4) );
  OR3_X1 npu_inst_pe_1_5_2_U25 ( .A1(npu_inst_pe_1_5_2_n4), .A2(
        npu_inst_pe_1_5_2_n8), .A3(npu_inst_pe_1_5_2_n7), .ZN(
        npu_inst_pe_1_5_2_n52) );
  OR3_X1 npu_inst_pe_1_5_2_U24 ( .A1(npu_inst_pe_1_5_2_n6), .A2(
        npu_inst_pe_1_5_2_n8), .A3(npu_inst_pe_1_5_2_n4), .ZN(
        npu_inst_pe_1_5_2_n60) );
  NOR2_X1 npu_inst_pe_1_5_2_U23 ( .A1(npu_inst_pe_1_5_2_n60), .A2(
        npu_inst_pe_1_5_2_n3), .ZN(npu_inst_pe_1_5_2_n58) );
  NOR2_X1 npu_inst_pe_1_5_2_U22 ( .A1(npu_inst_pe_1_5_2_n56), .A2(
        npu_inst_pe_1_5_2_n3), .ZN(npu_inst_pe_1_5_2_n54) );
  NOR2_X1 npu_inst_pe_1_5_2_U21 ( .A1(npu_inst_pe_1_5_2_n52), .A2(
        npu_inst_pe_1_5_2_n3), .ZN(npu_inst_pe_1_5_2_n50) );
  NOR2_X1 npu_inst_pe_1_5_2_U20 ( .A1(npu_inst_pe_1_5_2_n48), .A2(
        npu_inst_pe_1_5_2_n3), .ZN(npu_inst_pe_1_5_2_n46) );
  NOR2_X1 npu_inst_pe_1_5_2_U19 ( .A1(npu_inst_pe_1_5_2_n40), .A2(
        npu_inst_pe_1_5_2_n3), .ZN(npu_inst_pe_1_5_2_n38) );
  NOR2_X1 npu_inst_pe_1_5_2_U18 ( .A1(npu_inst_pe_1_5_2_n44), .A2(
        npu_inst_pe_1_5_2_n3), .ZN(npu_inst_pe_1_5_2_n42) );
  BUF_X1 npu_inst_pe_1_5_2_U17 ( .A(npu_inst_n97), .Z(npu_inst_pe_1_5_2_n8) );
  INV_X1 npu_inst_pe_1_5_2_U16 ( .A(npu_inst_n123), .ZN(npu_inst_pe_1_5_2_n12)
         );
  INV_X1 npu_inst_pe_1_5_2_U15 ( .A(npu_inst_pe_1_5_2_n38), .ZN(
        npu_inst_pe_1_5_2_n114) );
  INV_X1 npu_inst_pe_1_5_2_U14 ( .A(npu_inst_pe_1_5_2_n58), .ZN(
        npu_inst_pe_1_5_2_n119) );
  INV_X1 npu_inst_pe_1_5_2_U13 ( .A(npu_inst_pe_1_5_2_n54), .ZN(
        npu_inst_pe_1_5_2_n118) );
  INV_X1 npu_inst_pe_1_5_2_U12 ( .A(npu_inst_pe_1_5_2_n50), .ZN(
        npu_inst_pe_1_5_2_n117) );
  INV_X1 npu_inst_pe_1_5_2_U11 ( .A(npu_inst_pe_1_5_2_n46), .ZN(
        npu_inst_pe_1_5_2_n116) );
  INV_X1 npu_inst_pe_1_5_2_U10 ( .A(npu_inst_pe_1_5_2_n42), .ZN(
        npu_inst_pe_1_5_2_n115) );
  BUF_X1 npu_inst_pe_1_5_2_U9 ( .A(npu_inst_n17), .Z(npu_inst_pe_1_5_2_n2) );
  BUF_X1 npu_inst_pe_1_5_2_U8 ( .A(npu_inst_n17), .Z(npu_inst_pe_1_5_2_n1) );
  BUF_X1 npu_inst_pe_1_5_2_U7 ( .A(npu_inst_pe_1_5_2_n12), .Z(
        npu_inst_pe_1_5_2_n11) );
  BUF_X1 npu_inst_pe_1_5_2_U6 ( .A(npu_inst_pe_1_5_2_n12), .Z(
        npu_inst_pe_1_5_2_n10) );
  BUF_X1 npu_inst_pe_1_5_2_U5 ( .A(npu_inst_pe_1_5_2_n12), .Z(
        npu_inst_pe_1_5_2_n9) );
  NOR2_X1 npu_inst_pe_1_5_2_U4 ( .A1(npu_inst_pe_1_5_2_int_q_weight_0_), .A2(
        npu_inst_pe_1_5_2_n1), .ZN(npu_inst_pe_1_5_2_n76) );
  NOR2_X1 npu_inst_pe_1_5_2_U3 ( .A1(npu_inst_pe_1_5_2_n27), .A2(
        npu_inst_pe_1_5_2_n1), .ZN(npu_inst_pe_1_5_2_n77) );
  FA_X1 npu_inst_pe_1_5_2_sub_67_U2_1 ( .A(npu_inst_pe_1_5_2_int_q_acc_1_), 
        .B(npu_inst_pe_1_5_2_n14), .CI(npu_inst_pe_1_5_2_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_5_2_sub_67_carry_2_), .S(npu_inst_pe_1_5_2_N66) );
  FA_X1 npu_inst_pe_1_5_2_add_69_U1_1 ( .A(npu_inst_pe_1_5_2_int_q_acc_1_), 
        .B(npu_inst_pe_1_5_2_int_data_1_), .CI(
        npu_inst_pe_1_5_2_add_69_carry_1_), .CO(
        npu_inst_pe_1_5_2_add_69_carry_2_), .S(npu_inst_pe_1_5_2_N74) );
  NAND3_X1 npu_inst_pe_1_5_2_U109 ( .A1(npu_inst_pe_1_5_2_n5), .A2(
        npu_inst_pe_1_5_2_n7), .A3(npu_inst_pe_1_5_2_n8), .ZN(
        npu_inst_pe_1_5_2_n44) );
  NAND3_X1 npu_inst_pe_1_5_2_U108 ( .A1(npu_inst_pe_1_5_2_n4), .A2(
        npu_inst_pe_1_5_2_n7), .A3(npu_inst_pe_1_5_2_n8), .ZN(
        npu_inst_pe_1_5_2_n40) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_5_2_n34), .CK(
        npu_inst_pe_1_5_2_net3596), .RN(npu_inst_pe_1_5_2_n9), .Q(
        npu_inst_pe_1_5_2_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_5_2_n35), .CK(
        npu_inst_pe_1_5_2_net3596), .RN(npu_inst_pe_1_5_2_n9), .Q(
        npu_inst_pe_1_5_2_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_5_2_n36), .CK(
        npu_inst_pe_1_5_2_net3596), .RN(npu_inst_pe_1_5_2_n9), .Q(
        npu_inst_pe_1_5_2_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_5_2_n98), .CK(
        npu_inst_pe_1_5_2_net3596), .RN(npu_inst_pe_1_5_2_n9), .Q(
        npu_inst_pe_1_5_2_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_5_2_n99), .CK(
        npu_inst_pe_1_5_2_net3596), .RN(npu_inst_pe_1_5_2_n9), .Q(
        npu_inst_pe_1_5_2_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_5_2_n100), 
        .CK(npu_inst_pe_1_5_2_net3596), .RN(npu_inst_pe_1_5_2_n9), .Q(
        npu_inst_pe_1_5_2_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_5_2_n33), .CK(
        npu_inst_pe_1_5_2_net3596), .RN(npu_inst_pe_1_5_2_n9), .Q(
        npu_inst_pe_1_5_2_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_5_2_n101), 
        .CK(npu_inst_pe_1_5_2_net3596), .RN(npu_inst_pe_1_5_2_n9), .Q(
        npu_inst_pe_1_5_2_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_weight_reg_0_ ( .D(npu_inst_n109), .CK(
        npu_inst_pe_1_5_2_net3602), .RN(npu_inst_pe_1_5_2_n9), .Q(
        npu_inst_pe_1_5_2_int_q_weight_0_), .QN(npu_inst_pe_1_5_2_n27) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_weight_reg_1_ ( .D(npu_inst_n115), .CK(
        npu_inst_pe_1_5_2_net3602), .RN(npu_inst_pe_1_5_2_n9), .Q(
        npu_inst_pe_1_5_2_int_q_weight_1_), .QN(npu_inst_pe_1_5_2_n26) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_5_2_n113), 
        .CK(npu_inst_pe_1_5_2_net3602), .RN(npu_inst_pe_1_5_2_n9), .Q(
        npu_inst_pe_1_5_2_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_5_2_n107), 
        .CK(npu_inst_pe_1_5_2_net3602), .RN(npu_inst_pe_1_5_2_n9), .Q(
        npu_inst_pe_1_5_2_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_5_2_n112), 
        .CK(npu_inst_pe_1_5_2_net3602), .RN(npu_inst_pe_1_5_2_n10), .Q(
        npu_inst_pe_1_5_2_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_5_2_n106), 
        .CK(npu_inst_pe_1_5_2_net3602), .RN(npu_inst_pe_1_5_2_n10), .Q(
        npu_inst_pe_1_5_2_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_5_2_n111), 
        .CK(npu_inst_pe_1_5_2_net3602), .RN(npu_inst_pe_1_5_2_n10), .Q(
        npu_inst_pe_1_5_2_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_5_2_n105), 
        .CK(npu_inst_pe_1_5_2_net3602), .RN(npu_inst_pe_1_5_2_n10), .Q(
        npu_inst_pe_1_5_2_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_5_2_n110), 
        .CK(npu_inst_pe_1_5_2_net3602), .RN(npu_inst_pe_1_5_2_n10), .Q(
        npu_inst_pe_1_5_2_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_5_2_n104), 
        .CK(npu_inst_pe_1_5_2_net3602), .RN(npu_inst_pe_1_5_2_n10), .Q(
        npu_inst_pe_1_5_2_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_5_2_n109), 
        .CK(npu_inst_pe_1_5_2_net3602), .RN(npu_inst_pe_1_5_2_n10), .Q(
        npu_inst_pe_1_5_2_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_5_2_n103), 
        .CK(npu_inst_pe_1_5_2_net3602), .RN(npu_inst_pe_1_5_2_n10), .Q(
        npu_inst_pe_1_5_2_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_5_2_n108), 
        .CK(npu_inst_pe_1_5_2_net3602), .RN(npu_inst_pe_1_5_2_n10), .Q(
        npu_inst_pe_1_5_2_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_5_2_n102), 
        .CK(npu_inst_pe_1_5_2_net3602), .RN(npu_inst_pe_1_5_2_n10), .Q(
        npu_inst_pe_1_5_2_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_5_2_n86), 
        .CK(npu_inst_pe_1_5_2_net3602), .RN(npu_inst_pe_1_5_2_n10), .Q(
        npu_inst_pe_1_5_2_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_5_2_n87), 
        .CK(npu_inst_pe_1_5_2_net3602), .RN(npu_inst_pe_1_5_2_n10), .Q(
        npu_inst_pe_1_5_2_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_5_2_n88), 
        .CK(npu_inst_pe_1_5_2_net3602), .RN(npu_inst_pe_1_5_2_n11), .Q(
        npu_inst_pe_1_5_2_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_5_2_n89), 
        .CK(npu_inst_pe_1_5_2_net3602), .RN(npu_inst_pe_1_5_2_n11), .Q(
        npu_inst_pe_1_5_2_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_5_2_n90), 
        .CK(npu_inst_pe_1_5_2_net3602), .RN(npu_inst_pe_1_5_2_n11), .Q(
        npu_inst_pe_1_5_2_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_5_2_n91), 
        .CK(npu_inst_pe_1_5_2_net3602), .RN(npu_inst_pe_1_5_2_n11), .Q(
        npu_inst_pe_1_5_2_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_5_2_n92), 
        .CK(npu_inst_pe_1_5_2_net3602), .RN(npu_inst_pe_1_5_2_n11), .Q(
        npu_inst_pe_1_5_2_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_5_2_n93), 
        .CK(npu_inst_pe_1_5_2_net3602), .RN(npu_inst_pe_1_5_2_n11), .Q(
        npu_inst_pe_1_5_2_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_5_2_n94), 
        .CK(npu_inst_pe_1_5_2_net3602), .RN(npu_inst_pe_1_5_2_n11), .Q(
        npu_inst_pe_1_5_2_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_5_2_n95), 
        .CK(npu_inst_pe_1_5_2_net3602), .RN(npu_inst_pe_1_5_2_n11), .Q(
        npu_inst_pe_1_5_2_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_5_2_n96), 
        .CK(npu_inst_pe_1_5_2_net3602), .RN(npu_inst_pe_1_5_2_n11), .Q(
        npu_inst_pe_1_5_2_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_5_2_n97), 
        .CK(npu_inst_pe_1_5_2_net3602), .RN(npu_inst_pe_1_5_2_n11), .Q(
        npu_inst_pe_1_5_2_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_5_2_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_5_2_N84), .SE(1'b0), .GCK(npu_inst_pe_1_5_2_net3596) );
  CLKGATETST_X1 npu_inst_pe_1_5_2_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n62), .SE(1'b0), .GCK(npu_inst_pe_1_5_2_net3602) );
  MUX2_X1 npu_inst_pe_1_5_3_U162 ( .A(npu_inst_pe_1_5_3_n32), .B(
        npu_inst_pe_1_5_3_n29), .S(npu_inst_pe_1_5_3_n8), .Z(
        npu_inst_pe_1_5_3_N93) );
  MUX2_X1 npu_inst_pe_1_5_3_U161 ( .A(npu_inst_pe_1_5_3_n31), .B(
        npu_inst_pe_1_5_3_n30), .S(npu_inst_pe_1_5_3_n6), .Z(
        npu_inst_pe_1_5_3_n32) );
  MUX2_X1 npu_inst_pe_1_5_3_U160 ( .A(npu_inst_pe_1_5_3_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_5_3_int_q_reg_v_1__0_), .S(npu_inst_pe_1_5_3_n4), .Z(
        npu_inst_pe_1_5_3_n31) );
  MUX2_X1 npu_inst_pe_1_5_3_U159 ( .A(npu_inst_pe_1_5_3_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_5_3_int_q_reg_v_3__0_), .S(npu_inst_pe_1_5_3_n4), .Z(
        npu_inst_pe_1_5_3_n30) );
  MUX2_X1 npu_inst_pe_1_5_3_U158 ( .A(npu_inst_pe_1_5_3_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_5_3_int_q_reg_v_5__0_), .S(npu_inst_pe_1_5_3_n4), .Z(
        npu_inst_pe_1_5_3_n29) );
  MUX2_X1 npu_inst_pe_1_5_3_U157 ( .A(npu_inst_pe_1_5_3_n28), .B(
        npu_inst_pe_1_5_3_n23), .S(npu_inst_pe_1_5_3_n8), .Z(
        npu_inst_pe_1_5_3_N94) );
  MUX2_X1 npu_inst_pe_1_5_3_U156 ( .A(npu_inst_pe_1_5_3_n25), .B(
        npu_inst_pe_1_5_3_n24), .S(npu_inst_pe_1_5_3_n6), .Z(
        npu_inst_pe_1_5_3_n28) );
  MUX2_X1 npu_inst_pe_1_5_3_U155 ( .A(npu_inst_pe_1_5_3_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_5_3_int_q_reg_v_1__1_), .S(npu_inst_pe_1_5_3_n4), .Z(
        npu_inst_pe_1_5_3_n25) );
  MUX2_X1 npu_inst_pe_1_5_3_U154 ( .A(npu_inst_pe_1_5_3_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_5_3_int_q_reg_v_3__1_), .S(npu_inst_pe_1_5_3_n4), .Z(
        npu_inst_pe_1_5_3_n24) );
  MUX2_X1 npu_inst_pe_1_5_3_U153 ( .A(npu_inst_pe_1_5_3_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_5_3_int_q_reg_v_5__1_), .S(npu_inst_pe_1_5_3_n4), .Z(
        npu_inst_pe_1_5_3_n23) );
  MUX2_X1 npu_inst_pe_1_5_3_U152 ( .A(npu_inst_pe_1_5_3_n22), .B(
        npu_inst_pe_1_5_3_n19), .S(npu_inst_pe_1_5_3_n8), .Z(
        npu_inst_int_data_x_5__3__1_) );
  MUX2_X1 npu_inst_pe_1_5_3_U151 ( .A(npu_inst_pe_1_5_3_n21), .B(
        npu_inst_pe_1_5_3_n20), .S(npu_inst_pe_1_5_3_n6), .Z(
        npu_inst_pe_1_5_3_n22) );
  MUX2_X1 npu_inst_pe_1_5_3_U150 ( .A(npu_inst_pe_1_5_3_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_5_3_int_q_reg_h_1__1_), .S(npu_inst_pe_1_5_3_n4), .Z(
        npu_inst_pe_1_5_3_n21) );
  MUX2_X1 npu_inst_pe_1_5_3_U149 ( .A(npu_inst_pe_1_5_3_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_5_3_int_q_reg_h_3__1_), .S(npu_inst_pe_1_5_3_n4), .Z(
        npu_inst_pe_1_5_3_n20) );
  MUX2_X1 npu_inst_pe_1_5_3_U148 ( .A(npu_inst_pe_1_5_3_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_5_3_int_q_reg_h_5__1_), .S(npu_inst_pe_1_5_3_n4), .Z(
        npu_inst_pe_1_5_3_n19) );
  MUX2_X1 npu_inst_pe_1_5_3_U147 ( .A(npu_inst_pe_1_5_3_n18), .B(
        npu_inst_pe_1_5_3_n15), .S(npu_inst_pe_1_5_3_n8), .Z(
        npu_inst_int_data_x_5__3__0_) );
  MUX2_X1 npu_inst_pe_1_5_3_U146 ( .A(npu_inst_pe_1_5_3_n17), .B(
        npu_inst_pe_1_5_3_n16), .S(npu_inst_pe_1_5_3_n6), .Z(
        npu_inst_pe_1_5_3_n18) );
  MUX2_X1 npu_inst_pe_1_5_3_U145 ( .A(npu_inst_pe_1_5_3_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_5_3_int_q_reg_h_1__0_), .S(npu_inst_pe_1_5_3_n4), .Z(
        npu_inst_pe_1_5_3_n17) );
  MUX2_X1 npu_inst_pe_1_5_3_U144 ( .A(npu_inst_pe_1_5_3_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_5_3_int_q_reg_h_3__0_), .S(npu_inst_pe_1_5_3_n4), .Z(
        npu_inst_pe_1_5_3_n16) );
  MUX2_X1 npu_inst_pe_1_5_3_U143 ( .A(npu_inst_pe_1_5_3_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_5_3_int_q_reg_h_5__0_), .S(npu_inst_pe_1_5_3_n4), .Z(
        npu_inst_pe_1_5_3_n15) );
  XOR2_X1 npu_inst_pe_1_5_3_U142 ( .A(npu_inst_pe_1_5_3_int_data_0_), .B(
        npu_inst_pe_1_5_3_int_q_acc_0_), .Z(npu_inst_pe_1_5_3_N73) );
  AND2_X1 npu_inst_pe_1_5_3_U141 ( .A1(npu_inst_pe_1_5_3_int_q_acc_0_), .A2(
        npu_inst_pe_1_5_3_int_data_0_), .ZN(npu_inst_pe_1_5_3_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_5_3_U140 ( .A(npu_inst_pe_1_5_3_int_q_acc_0_), .B(
        npu_inst_pe_1_5_3_n13), .ZN(npu_inst_pe_1_5_3_N65) );
  OR2_X1 npu_inst_pe_1_5_3_U139 ( .A1(npu_inst_pe_1_5_3_n13), .A2(
        npu_inst_pe_1_5_3_int_q_acc_0_), .ZN(npu_inst_pe_1_5_3_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_5_3_U138 ( .A(npu_inst_pe_1_5_3_int_q_acc_2_), .B(
        npu_inst_pe_1_5_3_add_69_carry_2_), .Z(npu_inst_pe_1_5_3_N75) );
  AND2_X1 npu_inst_pe_1_5_3_U137 ( .A1(npu_inst_pe_1_5_3_add_69_carry_2_), 
        .A2(npu_inst_pe_1_5_3_int_q_acc_2_), .ZN(
        npu_inst_pe_1_5_3_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_5_3_U136 ( .A(npu_inst_pe_1_5_3_int_q_acc_3_), .B(
        npu_inst_pe_1_5_3_add_69_carry_3_), .Z(npu_inst_pe_1_5_3_N76) );
  AND2_X1 npu_inst_pe_1_5_3_U135 ( .A1(npu_inst_pe_1_5_3_add_69_carry_3_), 
        .A2(npu_inst_pe_1_5_3_int_q_acc_3_), .ZN(
        npu_inst_pe_1_5_3_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_5_3_U134 ( .A(npu_inst_pe_1_5_3_int_q_acc_4_), .B(
        npu_inst_pe_1_5_3_add_69_carry_4_), .Z(npu_inst_pe_1_5_3_N77) );
  AND2_X1 npu_inst_pe_1_5_3_U133 ( .A1(npu_inst_pe_1_5_3_add_69_carry_4_), 
        .A2(npu_inst_pe_1_5_3_int_q_acc_4_), .ZN(
        npu_inst_pe_1_5_3_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_5_3_U132 ( .A(npu_inst_pe_1_5_3_int_q_acc_5_), .B(
        npu_inst_pe_1_5_3_add_69_carry_5_), .Z(npu_inst_pe_1_5_3_N78) );
  AND2_X1 npu_inst_pe_1_5_3_U131 ( .A1(npu_inst_pe_1_5_3_add_69_carry_5_), 
        .A2(npu_inst_pe_1_5_3_int_q_acc_5_), .ZN(
        npu_inst_pe_1_5_3_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_5_3_U130 ( .A(npu_inst_pe_1_5_3_int_q_acc_6_), .B(
        npu_inst_pe_1_5_3_add_69_carry_6_), .Z(npu_inst_pe_1_5_3_N79) );
  AND2_X1 npu_inst_pe_1_5_3_U129 ( .A1(npu_inst_pe_1_5_3_add_69_carry_6_), 
        .A2(npu_inst_pe_1_5_3_int_q_acc_6_), .ZN(
        npu_inst_pe_1_5_3_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_5_3_U128 ( .A(npu_inst_pe_1_5_3_int_q_acc_7_), .B(
        npu_inst_pe_1_5_3_add_69_carry_7_), .Z(npu_inst_pe_1_5_3_N80) );
  XNOR2_X1 npu_inst_pe_1_5_3_U127 ( .A(npu_inst_pe_1_5_3_sub_67_carry_2_), .B(
        npu_inst_pe_1_5_3_int_q_acc_2_), .ZN(npu_inst_pe_1_5_3_N67) );
  OR2_X1 npu_inst_pe_1_5_3_U126 ( .A1(npu_inst_pe_1_5_3_int_q_acc_2_), .A2(
        npu_inst_pe_1_5_3_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_5_3_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_5_3_U125 ( .A(npu_inst_pe_1_5_3_sub_67_carry_3_), .B(
        npu_inst_pe_1_5_3_int_q_acc_3_), .ZN(npu_inst_pe_1_5_3_N68) );
  OR2_X1 npu_inst_pe_1_5_3_U124 ( .A1(npu_inst_pe_1_5_3_int_q_acc_3_), .A2(
        npu_inst_pe_1_5_3_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_5_3_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_5_3_U123 ( .A(npu_inst_pe_1_5_3_sub_67_carry_4_), .B(
        npu_inst_pe_1_5_3_int_q_acc_4_), .ZN(npu_inst_pe_1_5_3_N69) );
  OR2_X1 npu_inst_pe_1_5_3_U122 ( .A1(npu_inst_pe_1_5_3_int_q_acc_4_), .A2(
        npu_inst_pe_1_5_3_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_5_3_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_5_3_U121 ( .A(npu_inst_pe_1_5_3_sub_67_carry_5_), .B(
        npu_inst_pe_1_5_3_int_q_acc_5_), .ZN(npu_inst_pe_1_5_3_N70) );
  OR2_X1 npu_inst_pe_1_5_3_U120 ( .A1(npu_inst_pe_1_5_3_int_q_acc_5_), .A2(
        npu_inst_pe_1_5_3_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_5_3_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_5_3_U119 ( .A(npu_inst_pe_1_5_3_sub_67_carry_6_), .B(
        npu_inst_pe_1_5_3_int_q_acc_6_), .ZN(npu_inst_pe_1_5_3_N71) );
  OR2_X1 npu_inst_pe_1_5_3_U118 ( .A1(npu_inst_pe_1_5_3_int_q_acc_6_), .A2(
        npu_inst_pe_1_5_3_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_5_3_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_5_3_U117 ( .A(npu_inst_pe_1_5_3_int_q_acc_7_), .B(
        npu_inst_pe_1_5_3_sub_67_carry_7_), .ZN(npu_inst_pe_1_5_3_N72) );
  INV_X1 npu_inst_pe_1_5_3_U116 ( .A(npu_inst_n76), .ZN(npu_inst_pe_1_5_3_n7)
         );
  INV_X1 npu_inst_pe_1_5_3_U115 ( .A(npu_inst_pe_1_5_3_n7), .ZN(
        npu_inst_pe_1_5_3_n6) );
  INV_X1 npu_inst_pe_1_5_3_U114 ( .A(npu_inst_n54), .ZN(npu_inst_pe_1_5_3_n3)
         );
  AOI22_X1 npu_inst_pe_1_5_3_U113 ( .A1(npu_inst_int_data_y_6__3__0_), .A2(
        npu_inst_pe_1_5_3_n58), .B1(npu_inst_pe_1_5_3_n119), .B2(
        npu_inst_pe_1_5_3_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_5_3_n57) );
  INV_X1 npu_inst_pe_1_5_3_U112 ( .A(npu_inst_pe_1_5_3_n57), .ZN(
        npu_inst_pe_1_5_3_n108) );
  AOI22_X1 npu_inst_pe_1_5_3_U111 ( .A1(npu_inst_int_data_y_6__3__0_), .A2(
        npu_inst_pe_1_5_3_n54), .B1(npu_inst_pe_1_5_3_n118), .B2(
        npu_inst_pe_1_5_3_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_5_3_n53) );
  INV_X1 npu_inst_pe_1_5_3_U110 ( .A(npu_inst_pe_1_5_3_n53), .ZN(
        npu_inst_pe_1_5_3_n109) );
  AOI22_X1 npu_inst_pe_1_5_3_U107 ( .A1(npu_inst_int_data_y_6__3__0_), .A2(
        npu_inst_pe_1_5_3_n50), .B1(npu_inst_pe_1_5_3_n117), .B2(
        npu_inst_pe_1_5_3_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_5_3_n49) );
  INV_X1 npu_inst_pe_1_5_3_U106 ( .A(npu_inst_pe_1_5_3_n49), .ZN(
        npu_inst_pe_1_5_3_n110) );
  AOI22_X1 npu_inst_pe_1_5_3_U105 ( .A1(npu_inst_int_data_y_6__3__0_), .A2(
        npu_inst_pe_1_5_3_n46), .B1(npu_inst_pe_1_5_3_n116), .B2(
        npu_inst_pe_1_5_3_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_5_3_n45) );
  INV_X1 npu_inst_pe_1_5_3_U104 ( .A(npu_inst_pe_1_5_3_n45), .ZN(
        npu_inst_pe_1_5_3_n111) );
  AOI22_X1 npu_inst_pe_1_5_3_U103 ( .A1(npu_inst_int_data_y_6__3__0_), .A2(
        npu_inst_pe_1_5_3_n42), .B1(npu_inst_pe_1_5_3_n115), .B2(
        npu_inst_pe_1_5_3_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_5_3_n41) );
  INV_X1 npu_inst_pe_1_5_3_U102 ( .A(npu_inst_pe_1_5_3_n41), .ZN(
        npu_inst_pe_1_5_3_n112) );
  AOI22_X1 npu_inst_pe_1_5_3_U101 ( .A1(npu_inst_int_data_y_6__3__1_), .A2(
        npu_inst_pe_1_5_3_n58), .B1(npu_inst_pe_1_5_3_n119), .B2(
        npu_inst_pe_1_5_3_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_5_3_n59) );
  INV_X1 npu_inst_pe_1_5_3_U100 ( .A(npu_inst_pe_1_5_3_n59), .ZN(
        npu_inst_pe_1_5_3_n102) );
  AOI22_X1 npu_inst_pe_1_5_3_U99 ( .A1(npu_inst_int_data_y_6__3__1_), .A2(
        npu_inst_pe_1_5_3_n54), .B1(npu_inst_pe_1_5_3_n118), .B2(
        npu_inst_pe_1_5_3_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_5_3_n55) );
  INV_X1 npu_inst_pe_1_5_3_U98 ( .A(npu_inst_pe_1_5_3_n55), .ZN(
        npu_inst_pe_1_5_3_n103) );
  AOI22_X1 npu_inst_pe_1_5_3_U97 ( .A1(npu_inst_int_data_y_6__3__1_), .A2(
        npu_inst_pe_1_5_3_n50), .B1(npu_inst_pe_1_5_3_n117), .B2(
        npu_inst_pe_1_5_3_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_5_3_n51) );
  INV_X1 npu_inst_pe_1_5_3_U96 ( .A(npu_inst_pe_1_5_3_n51), .ZN(
        npu_inst_pe_1_5_3_n104) );
  AOI22_X1 npu_inst_pe_1_5_3_U95 ( .A1(npu_inst_int_data_y_6__3__1_), .A2(
        npu_inst_pe_1_5_3_n46), .B1(npu_inst_pe_1_5_3_n116), .B2(
        npu_inst_pe_1_5_3_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_5_3_n47) );
  INV_X1 npu_inst_pe_1_5_3_U94 ( .A(npu_inst_pe_1_5_3_n47), .ZN(
        npu_inst_pe_1_5_3_n105) );
  AOI22_X1 npu_inst_pe_1_5_3_U93 ( .A1(npu_inst_int_data_y_6__3__1_), .A2(
        npu_inst_pe_1_5_3_n42), .B1(npu_inst_pe_1_5_3_n115), .B2(
        npu_inst_pe_1_5_3_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_5_3_n43) );
  INV_X1 npu_inst_pe_1_5_3_U92 ( .A(npu_inst_pe_1_5_3_n43), .ZN(
        npu_inst_pe_1_5_3_n106) );
  AOI22_X1 npu_inst_pe_1_5_3_U91 ( .A1(npu_inst_pe_1_5_3_n38), .A2(
        npu_inst_int_data_y_6__3__1_), .B1(npu_inst_pe_1_5_3_n114), .B2(
        npu_inst_pe_1_5_3_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_5_3_n39) );
  INV_X1 npu_inst_pe_1_5_3_U90 ( .A(npu_inst_pe_1_5_3_n39), .ZN(
        npu_inst_pe_1_5_3_n107) );
  AOI22_X1 npu_inst_pe_1_5_3_U89 ( .A1(npu_inst_pe_1_5_3_n38), .A2(
        npu_inst_int_data_y_6__3__0_), .B1(npu_inst_pe_1_5_3_n114), .B2(
        npu_inst_pe_1_5_3_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_5_3_n37) );
  INV_X1 npu_inst_pe_1_5_3_U88 ( .A(npu_inst_pe_1_5_3_n37), .ZN(
        npu_inst_pe_1_5_3_n113) );
  NAND2_X1 npu_inst_pe_1_5_3_U87 ( .A1(npu_inst_pe_1_5_3_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_5_3_n60), .ZN(npu_inst_pe_1_5_3_n74) );
  OAI21_X1 npu_inst_pe_1_5_3_U86 ( .B1(npu_inst_pe_1_5_3_n63), .B2(
        npu_inst_pe_1_5_3_n60), .A(npu_inst_pe_1_5_3_n74), .ZN(
        npu_inst_pe_1_5_3_n97) );
  NAND2_X1 npu_inst_pe_1_5_3_U85 ( .A1(npu_inst_pe_1_5_3_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_5_3_n60), .ZN(npu_inst_pe_1_5_3_n73) );
  OAI21_X1 npu_inst_pe_1_5_3_U84 ( .B1(npu_inst_pe_1_5_3_n61), .B2(
        npu_inst_pe_1_5_3_n60), .A(npu_inst_pe_1_5_3_n73), .ZN(
        npu_inst_pe_1_5_3_n96) );
  NAND2_X1 npu_inst_pe_1_5_3_U83 ( .A1(npu_inst_pe_1_5_3_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_5_3_n56), .ZN(npu_inst_pe_1_5_3_n72) );
  OAI21_X1 npu_inst_pe_1_5_3_U82 ( .B1(npu_inst_pe_1_5_3_n63), .B2(
        npu_inst_pe_1_5_3_n56), .A(npu_inst_pe_1_5_3_n72), .ZN(
        npu_inst_pe_1_5_3_n95) );
  NAND2_X1 npu_inst_pe_1_5_3_U81 ( .A1(npu_inst_pe_1_5_3_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_5_3_n56), .ZN(npu_inst_pe_1_5_3_n71) );
  OAI21_X1 npu_inst_pe_1_5_3_U80 ( .B1(npu_inst_pe_1_5_3_n61), .B2(
        npu_inst_pe_1_5_3_n56), .A(npu_inst_pe_1_5_3_n71), .ZN(
        npu_inst_pe_1_5_3_n94) );
  NAND2_X1 npu_inst_pe_1_5_3_U79 ( .A1(npu_inst_pe_1_5_3_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_5_3_n52), .ZN(npu_inst_pe_1_5_3_n70) );
  OAI21_X1 npu_inst_pe_1_5_3_U78 ( .B1(npu_inst_pe_1_5_3_n63), .B2(
        npu_inst_pe_1_5_3_n52), .A(npu_inst_pe_1_5_3_n70), .ZN(
        npu_inst_pe_1_5_3_n93) );
  NAND2_X1 npu_inst_pe_1_5_3_U77 ( .A1(npu_inst_pe_1_5_3_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_5_3_n52), .ZN(npu_inst_pe_1_5_3_n69) );
  OAI21_X1 npu_inst_pe_1_5_3_U76 ( .B1(npu_inst_pe_1_5_3_n61), .B2(
        npu_inst_pe_1_5_3_n52), .A(npu_inst_pe_1_5_3_n69), .ZN(
        npu_inst_pe_1_5_3_n92) );
  NAND2_X1 npu_inst_pe_1_5_3_U75 ( .A1(npu_inst_pe_1_5_3_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_5_3_n48), .ZN(npu_inst_pe_1_5_3_n68) );
  OAI21_X1 npu_inst_pe_1_5_3_U74 ( .B1(npu_inst_pe_1_5_3_n63), .B2(
        npu_inst_pe_1_5_3_n48), .A(npu_inst_pe_1_5_3_n68), .ZN(
        npu_inst_pe_1_5_3_n91) );
  NAND2_X1 npu_inst_pe_1_5_3_U73 ( .A1(npu_inst_pe_1_5_3_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_5_3_n48), .ZN(npu_inst_pe_1_5_3_n67) );
  OAI21_X1 npu_inst_pe_1_5_3_U72 ( .B1(npu_inst_pe_1_5_3_n61), .B2(
        npu_inst_pe_1_5_3_n48), .A(npu_inst_pe_1_5_3_n67), .ZN(
        npu_inst_pe_1_5_3_n90) );
  NAND2_X1 npu_inst_pe_1_5_3_U71 ( .A1(npu_inst_pe_1_5_3_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_5_3_n44), .ZN(npu_inst_pe_1_5_3_n66) );
  OAI21_X1 npu_inst_pe_1_5_3_U70 ( .B1(npu_inst_pe_1_5_3_n63), .B2(
        npu_inst_pe_1_5_3_n44), .A(npu_inst_pe_1_5_3_n66), .ZN(
        npu_inst_pe_1_5_3_n89) );
  NAND2_X1 npu_inst_pe_1_5_3_U69 ( .A1(npu_inst_pe_1_5_3_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_5_3_n44), .ZN(npu_inst_pe_1_5_3_n65) );
  OAI21_X1 npu_inst_pe_1_5_3_U68 ( .B1(npu_inst_pe_1_5_3_n61), .B2(
        npu_inst_pe_1_5_3_n44), .A(npu_inst_pe_1_5_3_n65), .ZN(
        npu_inst_pe_1_5_3_n88) );
  NAND2_X1 npu_inst_pe_1_5_3_U67 ( .A1(npu_inst_pe_1_5_3_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_5_3_n40), .ZN(npu_inst_pe_1_5_3_n64) );
  OAI21_X1 npu_inst_pe_1_5_3_U66 ( .B1(npu_inst_pe_1_5_3_n63), .B2(
        npu_inst_pe_1_5_3_n40), .A(npu_inst_pe_1_5_3_n64), .ZN(
        npu_inst_pe_1_5_3_n87) );
  NAND2_X1 npu_inst_pe_1_5_3_U65 ( .A1(npu_inst_pe_1_5_3_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_5_3_n40), .ZN(npu_inst_pe_1_5_3_n62) );
  OAI21_X1 npu_inst_pe_1_5_3_U64 ( .B1(npu_inst_pe_1_5_3_n61), .B2(
        npu_inst_pe_1_5_3_n40), .A(npu_inst_pe_1_5_3_n62), .ZN(
        npu_inst_pe_1_5_3_n86) );
  AND2_X1 npu_inst_pe_1_5_3_U63 ( .A1(npu_inst_pe_1_5_3_N93), .A2(npu_inst_n54), .ZN(npu_inst_int_data_y_5__3__0_) );
  AND2_X1 npu_inst_pe_1_5_3_U62 ( .A1(npu_inst_n54), .A2(npu_inst_pe_1_5_3_N94), .ZN(npu_inst_int_data_y_5__3__1_) );
  NOR3_X1 npu_inst_pe_1_5_3_U61 ( .A1(npu_inst_pe_1_5_3_n26), .A2(npu_inst_n54), .A3(npu_inst_int_ckg[20]), .ZN(npu_inst_pe_1_5_3_n85) );
  OR2_X1 npu_inst_pe_1_5_3_U60 ( .A1(npu_inst_pe_1_5_3_n85), .A2(
        npu_inst_pe_1_5_3_n2), .ZN(npu_inst_pe_1_5_3_N84) );
  AND2_X1 npu_inst_pe_1_5_3_U59 ( .A1(npu_inst_pe_1_5_3_int_q_acc_0_), .A2(
        npu_inst_pe_1_5_3_n1), .ZN(npu_inst_int_data_res_5__3__0_) );
  AND2_X1 npu_inst_pe_1_5_3_U58 ( .A1(npu_inst_pe_1_5_3_n2), .A2(
        npu_inst_pe_1_5_3_int_q_acc_7_), .ZN(npu_inst_int_data_res_5__3__7_)
         );
  AND2_X1 npu_inst_pe_1_5_3_U57 ( .A1(npu_inst_pe_1_5_3_int_q_acc_1_), .A2(
        npu_inst_pe_1_5_3_n1), .ZN(npu_inst_int_data_res_5__3__1_) );
  AND2_X1 npu_inst_pe_1_5_3_U56 ( .A1(npu_inst_pe_1_5_3_int_q_acc_2_), .A2(
        npu_inst_pe_1_5_3_n1), .ZN(npu_inst_int_data_res_5__3__2_) );
  AND2_X1 npu_inst_pe_1_5_3_U55 ( .A1(npu_inst_pe_1_5_3_int_q_acc_3_), .A2(
        npu_inst_pe_1_5_3_n2), .ZN(npu_inst_int_data_res_5__3__3_) );
  AND2_X1 npu_inst_pe_1_5_3_U54 ( .A1(npu_inst_pe_1_5_3_int_q_acc_4_), .A2(
        npu_inst_pe_1_5_3_n2), .ZN(npu_inst_int_data_res_5__3__4_) );
  AND2_X1 npu_inst_pe_1_5_3_U53 ( .A1(npu_inst_pe_1_5_3_int_q_acc_5_), .A2(
        npu_inst_pe_1_5_3_n2), .ZN(npu_inst_int_data_res_5__3__5_) );
  AND2_X1 npu_inst_pe_1_5_3_U52 ( .A1(npu_inst_pe_1_5_3_int_q_acc_6_), .A2(
        npu_inst_pe_1_5_3_n2), .ZN(npu_inst_int_data_res_5__3__6_) );
  AOI222_X1 npu_inst_pe_1_5_3_U51 ( .A1(npu_inst_int_data_res_6__3__0_), .A2(
        npu_inst_pe_1_5_3_n1), .B1(npu_inst_pe_1_5_3_N73), .B2(
        npu_inst_pe_1_5_3_n76), .C1(npu_inst_pe_1_5_3_N65), .C2(
        npu_inst_pe_1_5_3_n77), .ZN(npu_inst_pe_1_5_3_n84) );
  INV_X1 npu_inst_pe_1_5_3_U50 ( .A(npu_inst_pe_1_5_3_n84), .ZN(
        npu_inst_pe_1_5_3_n101) );
  AOI222_X1 npu_inst_pe_1_5_3_U49 ( .A1(npu_inst_int_data_res_6__3__7_), .A2(
        npu_inst_pe_1_5_3_n1), .B1(npu_inst_pe_1_5_3_N80), .B2(
        npu_inst_pe_1_5_3_n76), .C1(npu_inst_pe_1_5_3_N72), .C2(
        npu_inst_pe_1_5_3_n77), .ZN(npu_inst_pe_1_5_3_n75) );
  INV_X1 npu_inst_pe_1_5_3_U48 ( .A(npu_inst_pe_1_5_3_n75), .ZN(
        npu_inst_pe_1_5_3_n33) );
  AOI222_X1 npu_inst_pe_1_5_3_U47 ( .A1(npu_inst_int_data_res_6__3__1_), .A2(
        npu_inst_pe_1_5_3_n1), .B1(npu_inst_pe_1_5_3_N74), .B2(
        npu_inst_pe_1_5_3_n76), .C1(npu_inst_pe_1_5_3_N66), .C2(
        npu_inst_pe_1_5_3_n77), .ZN(npu_inst_pe_1_5_3_n83) );
  INV_X1 npu_inst_pe_1_5_3_U46 ( .A(npu_inst_pe_1_5_3_n83), .ZN(
        npu_inst_pe_1_5_3_n100) );
  AOI222_X1 npu_inst_pe_1_5_3_U45 ( .A1(npu_inst_int_data_res_6__3__2_), .A2(
        npu_inst_pe_1_5_3_n1), .B1(npu_inst_pe_1_5_3_N75), .B2(
        npu_inst_pe_1_5_3_n76), .C1(npu_inst_pe_1_5_3_N67), .C2(
        npu_inst_pe_1_5_3_n77), .ZN(npu_inst_pe_1_5_3_n82) );
  INV_X1 npu_inst_pe_1_5_3_U44 ( .A(npu_inst_pe_1_5_3_n82), .ZN(
        npu_inst_pe_1_5_3_n99) );
  AOI222_X1 npu_inst_pe_1_5_3_U43 ( .A1(npu_inst_int_data_res_6__3__3_), .A2(
        npu_inst_pe_1_5_3_n1), .B1(npu_inst_pe_1_5_3_N76), .B2(
        npu_inst_pe_1_5_3_n76), .C1(npu_inst_pe_1_5_3_N68), .C2(
        npu_inst_pe_1_5_3_n77), .ZN(npu_inst_pe_1_5_3_n81) );
  INV_X1 npu_inst_pe_1_5_3_U42 ( .A(npu_inst_pe_1_5_3_n81), .ZN(
        npu_inst_pe_1_5_3_n98) );
  AOI222_X1 npu_inst_pe_1_5_3_U41 ( .A1(npu_inst_int_data_res_6__3__4_), .A2(
        npu_inst_pe_1_5_3_n1), .B1(npu_inst_pe_1_5_3_N77), .B2(
        npu_inst_pe_1_5_3_n76), .C1(npu_inst_pe_1_5_3_N69), .C2(
        npu_inst_pe_1_5_3_n77), .ZN(npu_inst_pe_1_5_3_n80) );
  INV_X1 npu_inst_pe_1_5_3_U40 ( .A(npu_inst_pe_1_5_3_n80), .ZN(
        npu_inst_pe_1_5_3_n36) );
  AOI222_X1 npu_inst_pe_1_5_3_U39 ( .A1(npu_inst_int_data_res_6__3__5_), .A2(
        npu_inst_pe_1_5_3_n1), .B1(npu_inst_pe_1_5_3_N78), .B2(
        npu_inst_pe_1_5_3_n76), .C1(npu_inst_pe_1_5_3_N70), .C2(
        npu_inst_pe_1_5_3_n77), .ZN(npu_inst_pe_1_5_3_n79) );
  INV_X1 npu_inst_pe_1_5_3_U38 ( .A(npu_inst_pe_1_5_3_n79), .ZN(
        npu_inst_pe_1_5_3_n35) );
  AOI222_X1 npu_inst_pe_1_5_3_U37 ( .A1(npu_inst_int_data_res_6__3__6_), .A2(
        npu_inst_pe_1_5_3_n1), .B1(npu_inst_pe_1_5_3_N79), .B2(
        npu_inst_pe_1_5_3_n76), .C1(npu_inst_pe_1_5_3_N71), .C2(
        npu_inst_pe_1_5_3_n77), .ZN(npu_inst_pe_1_5_3_n78) );
  INV_X1 npu_inst_pe_1_5_3_U36 ( .A(npu_inst_pe_1_5_3_n78), .ZN(
        npu_inst_pe_1_5_3_n34) );
  INV_X1 npu_inst_pe_1_5_3_U35 ( .A(npu_inst_pe_1_5_3_int_data_1_), .ZN(
        npu_inst_pe_1_5_3_n14) );
  AND2_X1 npu_inst_pe_1_5_3_U34 ( .A1(npu_inst_int_data_x_5__3__1_), .A2(
        npu_inst_pe_1_5_3_int_q_weight_1_), .ZN(npu_inst_pe_1_5_3_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_5_3_U33 ( .A1(npu_inst_int_data_x_5__3__0_), .A2(
        npu_inst_pe_1_5_3_int_q_weight_1_), .ZN(npu_inst_pe_1_5_3_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_5_3_U32 ( .A1(npu_inst_n54), .A2(
        npu_inst_int_data_y_6__3__1_), .B1(npu_inst_pe_1_5_3_n3), .B2(
        npu_inst_int_data_x_5__4__1_), .ZN(npu_inst_pe_1_5_3_n63) );
  AOI22_X1 npu_inst_pe_1_5_3_U31 ( .A1(npu_inst_n54), .A2(
        npu_inst_int_data_y_6__3__0_), .B1(npu_inst_pe_1_5_3_n3), .B2(
        npu_inst_int_data_x_5__4__0_), .ZN(npu_inst_pe_1_5_3_n61) );
  INV_X1 npu_inst_pe_1_5_3_U30 ( .A(npu_inst_pe_1_5_3_int_data_0_), .ZN(
        npu_inst_pe_1_5_3_n13) );
  INV_X1 npu_inst_pe_1_5_3_U29 ( .A(npu_inst_n68), .ZN(npu_inst_pe_1_5_3_n5)
         );
  OR3_X1 npu_inst_pe_1_5_3_U28 ( .A1(npu_inst_pe_1_5_3_n6), .A2(
        npu_inst_pe_1_5_3_n8), .A3(npu_inst_pe_1_5_3_n5), .ZN(
        npu_inst_pe_1_5_3_n56) );
  OR3_X1 npu_inst_pe_1_5_3_U27 ( .A1(npu_inst_pe_1_5_3_n5), .A2(
        npu_inst_pe_1_5_3_n8), .A3(npu_inst_pe_1_5_3_n7), .ZN(
        npu_inst_pe_1_5_3_n48) );
  INV_X1 npu_inst_pe_1_5_3_U26 ( .A(npu_inst_pe_1_5_3_n5), .ZN(
        npu_inst_pe_1_5_3_n4) );
  OR3_X1 npu_inst_pe_1_5_3_U25 ( .A1(npu_inst_pe_1_5_3_n4), .A2(
        npu_inst_pe_1_5_3_n8), .A3(npu_inst_pe_1_5_3_n7), .ZN(
        npu_inst_pe_1_5_3_n52) );
  OR3_X1 npu_inst_pe_1_5_3_U24 ( .A1(npu_inst_pe_1_5_3_n6), .A2(
        npu_inst_pe_1_5_3_n8), .A3(npu_inst_pe_1_5_3_n4), .ZN(
        npu_inst_pe_1_5_3_n60) );
  NOR2_X1 npu_inst_pe_1_5_3_U23 ( .A1(npu_inst_pe_1_5_3_n60), .A2(
        npu_inst_pe_1_5_3_n3), .ZN(npu_inst_pe_1_5_3_n58) );
  NOR2_X1 npu_inst_pe_1_5_3_U22 ( .A1(npu_inst_pe_1_5_3_n56), .A2(
        npu_inst_pe_1_5_3_n3), .ZN(npu_inst_pe_1_5_3_n54) );
  NOR2_X1 npu_inst_pe_1_5_3_U21 ( .A1(npu_inst_pe_1_5_3_n52), .A2(
        npu_inst_pe_1_5_3_n3), .ZN(npu_inst_pe_1_5_3_n50) );
  NOR2_X1 npu_inst_pe_1_5_3_U20 ( .A1(npu_inst_pe_1_5_3_n48), .A2(
        npu_inst_pe_1_5_3_n3), .ZN(npu_inst_pe_1_5_3_n46) );
  NOR2_X1 npu_inst_pe_1_5_3_U19 ( .A1(npu_inst_pe_1_5_3_n40), .A2(
        npu_inst_pe_1_5_3_n3), .ZN(npu_inst_pe_1_5_3_n38) );
  NOR2_X1 npu_inst_pe_1_5_3_U18 ( .A1(npu_inst_pe_1_5_3_n44), .A2(
        npu_inst_pe_1_5_3_n3), .ZN(npu_inst_pe_1_5_3_n42) );
  BUF_X1 npu_inst_pe_1_5_3_U17 ( .A(npu_inst_n97), .Z(npu_inst_pe_1_5_3_n8) );
  INV_X1 npu_inst_pe_1_5_3_U16 ( .A(npu_inst_n123), .ZN(npu_inst_pe_1_5_3_n12)
         );
  INV_X1 npu_inst_pe_1_5_3_U15 ( .A(npu_inst_pe_1_5_3_n38), .ZN(
        npu_inst_pe_1_5_3_n114) );
  INV_X1 npu_inst_pe_1_5_3_U14 ( .A(npu_inst_pe_1_5_3_n58), .ZN(
        npu_inst_pe_1_5_3_n119) );
  INV_X1 npu_inst_pe_1_5_3_U13 ( .A(npu_inst_pe_1_5_3_n54), .ZN(
        npu_inst_pe_1_5_3_n118) );
  INV_X1 npu_inst_pe_1_5_3_U12 ( .A(npu_inst_pe_1_5_3_n50), .ZN(
        npu_inst_pe_1_5_3_n117) );
  INV_X1 npu_inst_pe_1_5_3_U11 ( .A(npu_inst_pe_1_5_3_n46), .ZN(
        npu_inst_pe_1_5_3_n116) );
  INV_X1 npu_inst_pe_1_5_3_U10 ( .A(npu_inst_pe_1_5_3_n42), .ZN(
        npu_inst_pe_1_5_3_n115) );
  BUF_X1 npu_inst_pe_1_5_3_U9 ( .A(npu_inst_n17), .Z(npu_inst_pe_1_5_3_n2) );
  BUF_X1 npu_inst_pe_1_5_3_U8 ( .A(npu_inst_n17), .Z(npu_inst_pe_1_5_3_n1) );
  BUF_X1 npu_inst_pe_1_5_3_U7 ( .A(npu_inst_pe_1_5_3_n12), .Z(
        npu_inst_pe_1_5_3_n11) );
  BUF_X1 npu_inst_pe_1_5_3_U6 ( .A(npu_inst_pe_1_5_3_n12), .Z(
        npu_inst_pe_1_5_3_n10) );
  BUF_X1 npu_inst_pe_1_5_3_U5 ( .A(npu_inst_pe_1_5_3_n12), .Z(
        npu_inst_pe_1_5_3_n9) );
  NOR2_X1 npu_inst_pe_1_5_3_U4 ( .A1(npu_inst_pe_1_5_3_int_q_weight_0_), .A2(
        npu_inst_pe_1_5_3_n1), .ZN(npu_inst_pe_1_5_3_n76) );
  NOR2_X1 npu_inst_pe_1_5_3_U3 ( .A1(npu_inst_pe_1_5_3_n27), .A2(
        npu_inst_pe_1_5_3_n1), .ZN(npu_inst_pe_1_5_3_n77) );
  FA_X1 npu_inst_pe_1_5_3_sub_67_U2_1 ( .A(npu_inst_pe_1_5_3_int_q_acc_1_), 
        .B(npu_inst_pe_1_5_3_n14), .CI(npu_inst_pe_1_5_3_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_5_3_sub_67_carry_2_), .S(npu_inst_pe_1_5_3_N66) );
  FA_X1 npu_inst_pe_1_5_3_add_69_U1_1 ( .A(npu_inst_pe_1_5_3_int_q_acc_1_), 
        .B(npu_inst_pe_1_5_3_int_data_1_), .CI(
        npu_inst_pe_1_5_3_add_69_carry_1_), .CO(
        npu_inst_pe_1_5_3_add_69_carry_2_), .S(npu_inst_pe_1_5_3_N74) );
  NAND3_X1 npu_inst_pe_1_5_3_U109 ( .A1(npu_inst_pe_1_5_3_n5), .A2(
        npu_inst_pe_1_5_3_n7), .A3(npu_inst_pe_1_5_3_n8), .ZN(
        npu_inst_pe_1_5_3_n44) );
  NAND3_X1 npu_inst_pe_1_5_3_U108 ( .A1(npu_inst_pe_1_5_3_n4), .A2(
        npu_inst_pe_1_5_3_n7), .A3(npu_inst_pe_1_5_3_n8), .ZN(
        npu_inst_pe_1_5_3_n40) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_5_3_n34), .CK(
        npu_inst_pe_1_5_3_net3573), .RN(npu_inst_pe_1_5_3_n9), .Q(
        npu_inst_pe_1_5_3_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_5_3_n35), .CK(
        npu_inst_pe_1_5_3_net3573), .RN(npu_inst_pe_1_5_3_n9), .Q(
        npu_inst_pe_1_5_3_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_5_3_n36), .CK(
        npu_inst_pe_1_5_3_net3573), .RN(npu_inst_pe_1_5_3_n9), .Q(
        npu_inst_pe_1_5_3_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_5_3_n98), .CK(
        npu_inst_pe_1_5_3_net3573), .RN(npu_inst_pe_1_5_3_n9), .Q(
        npu_inst_pe_1_5_3_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_5_3_n99), .CK(
        npu_inst_pe_1_5_3_net3573), .RN(npu_inst_pe_1_5_3_n9), .Q(
        npu_inst_pe_1_5_3_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_5_3_n100), 
        .CK(npu_inst_pe_1_5_3_net3573), .RN(npu_inst_pe_1_5_3_n9), .Q(
        npu_inst_pe_1_5_3_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_5_3_n33), .CK(
        npu_inst_pe_1_5_3_net3573), .RN(npu_inst_pe_1_5_3_n9), .Q(
        npu_inst_pe_1_5_3_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_5_3_n101), 
        .CK(npu_inst_pe_1_5_3_net3573), .RN(npu_inst_pe_1_5_3_n9), .Q(
        npu_inst_pe_1_5_3_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_weight_reg_0_ ( .D(npu_inst_n109), .CK(
        npu_inst_pe_1_5_3_net3579), .RN(npu_inst_pe_1_5_3_n9), .Q(
        npu_inst_pe_1_5_3_int_q_weight_0_), .QN(npu_inst_pe_1_5_3_n27) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_weight_reg_1_ ( .D(npu_inst_n115), .CK(
        npu_inst_pe_1_5_3_net3579), .RN(npu_inst_pe_1_5_3_n9), .Q(
        npu_inst_pe_1_5_3_int_q_weight_1_), .QN(npu_inst_pe_1_5_3_n26) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_5_3_n113), 
        .CK(npu_inst_pe_1_5_3_net3579), .RN(npu_inst_pe_1_5_3_n9), .Q(
        npu_inst_pe_1_5_3_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_5_3_n107), 
        .CK(npu_inst_pe_1_5_3_net3579), .RN(npu_inst_pe_1_5_3_n9), .Q(
        npu_inst_pe_1_5_3_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_5_3_n112), 
        .CK(npu_inst_pe_1_5_3_net3579), .RN(npu_inst_pe_1_5_3_n10), .Q(
        npu_inst_pe_1_5_3_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_5_3_n106), 
        .CK(npu_inst_pe_1_5_3_net3579), .RN(npu_inst_pe_1_5_3_n10), .Q(
        npu_inst_pe_1_5_3_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_5_3_n111), 
        .CK(npu_inst_pe_1_5_3_net3579), .RN(npu_inst_pe_1_5_3_n10), .Q(
        npu_inst_pe_1_5_3_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_5_3_n105), 
        .CK(npu_inst_pe_1_5_3_net3579), .RN(npu_inst_pe_1_5_3_n10), .Q(
        npu_inst_pe_1_5_3_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_5_3_n110), 
        .CK(npu_inst_pe_1_5_3_net3579), .RN(npu_inst_pe_1_5_3_n10), .Q(
        npu_inst_pe_1_5_3_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_5_3_n104), 
        .CK(npu_inst_pe_1_5_3_net3579), .RN(npu_inst_pe_1_5_3_n10), .Q(
        npu_inst_pe_1_5_3_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_5_3_n109), 
        .CK(npu_inst_pe_1_5_3_net3579), .RN(npu_inst_pe_1_5_3_n10), .Q(
        npu_inst_pe_1_5_3_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_5_3_n103), 
        .CK(npu_inst_pe_1_5_3_net3579), .RN(npu_inst_pe_1_5_3_n10), .Q(
        npu_inst_pe_1_5_3_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_5_3_n108), 
        .CK(npu_inst_pe_1_5_3_net3579), .RN(npu_inst_pe_1_5_3_n10), .Q(
        npu_inst_pe_1_5_3_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_5_3_n102), 
        .CK(npu_inst_pe_1_5_3_net3579), .RN(npu_inst_pe_1_5_3_n10), .Q(
        npu_inst_pe_1_5_3_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_5_3_n86), 
        .CK(npu_inst_pe_1_5_3_net3579), .RN(npu_inst_pe_1_5_3_n10), .Q(
        npu_inst_pe_1_5_3_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_5_3_n87), 
        .CK(npu_inst_pe_1_5_3_net3579), .RN(npu_inst_pe_1_5_3_n10), .Q(
        npu_inst_pe_1_5_3_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_5_3_n88), 
        .CK(npu_inst_pe_1_5_3_net3579), .RN(npu_inst_pe_1_5_3_n11), .Q(
        npu_inst_pe_1_5_3_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_5_3_n89), 
        .CK(npu_inst_pe_1_5_3_net3579), .RN(npu_inst_pe_1_5_3_n11), .Q(
        npu_inst_pe_1_5_3_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_5_3_n90), 
        .CK(npu_inst_pe_1_5_3_net3579), .RN(npu_inst_pe_1_5_3_n11), .Q(
        npu_inst_pe_1_5_3_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_5_3_n91), 
        .CK(npu_inst_pe_1_5_3_net3579), .RN(npu_inst_pe_1_5_3_n11), .Q(
        npu_inst_pe_1_5_3_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_5_3_n92), 
        .CK(npu_inst_pe_1_5_3_net3579), .RN(npu_inst_pe_1_5_3_n11), .Q(
        npu_inst_pe_1_5_3_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_5_3_n93), 
        .CK(npu_inst_pe_1_5_3_net3579), .RN(npu_inst_pe_1_5_3_n11), .Q(
        npu_inst_pe_1_5_3_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_5_3_n94), 
        .CK(npu_inst_pe_1_5_3_net3579), .RN(npu_inst_pe_1_5_3_n11), .Q(
        npu_inst_pe_1_5_3_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_5_3_n95), 
        .CK(npu_inst_pe_1_5_3_net3579), .RN(npu_inst_pe_1_5_3_n11), .Q(
        npu_inst_pe_1_5_3_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_5_3_n96), 
        .CK(npu_inst_pe_1_5_3_net3579), .RN(npu_inst_pe_1_5_3_n11), .Q(
        npu_inst_pe_1_5_3_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_5_3_n97), 
        .CK(npu_inst_pe_1_5_3_net3579), .RN(npu_inst_pe_1_5_3_n11), .Q(
        npu_inst_pe_1_5_3_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_5_3_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_5_3_N84), .SE(1'b0), .GCK(npu_inst_pe_1_5_3_net3573) );
  CLKGATETST_X1 npu_inst_pe_1_5_3_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n62), .SE(1'b0), .GCK(npu_inst_pe_1_5_3_net3579) );
  MUX2_X1 npu_inst_pe_1_5_4_U162 ( .A(npu_inst_pe_1_5_4_n32), .B(
        npu_inst_pe_1_5_4_n29), .S(npu_inst_pe_1_5_4_n8), .Z(
        npu_inst_pe_1_5_4_N93) );
  MUX2_X1 npu_inst_pe_1_5_4_U161 ( .A(npu_inst_pe_1_5_4_n31), .B(
        npu_inst_pe_1_5_4_n30), .S(npu_inst_pe_1_5_4_n6), .Z(
        npu_inst_pe_1_5_4_n32) );
  MUX2_X1 npu_inst_pe_1_5_4_U160 ( .A(npu_inst_pe_1_5_4_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_5_4_int_q_reg_v_1__0_), .S(npu_inst_pe_1_5_4_n4), .Z(
        npu_inst_pe_1_5_4_n31) );
  MUX2_X1 npu_inst_pe_1_5_4_U159 ( .A(npu_inst_pe_1_5_4_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_5_4_int_q_reg_v_3__0_), .S(npu_inst_pe_1_5_4_n4), .Z(
        npu_inst_pe_1_5_4_n30) );
  MUX2_X1 npu_inst_pe_1_5_4_U158 ( .A(npu_inst_pe_1_5_4_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_5_4_int_q_reg_v_5__0_), .S(npu_inst_pe_1_5_4_n4), .Z(
        npu_inst_pe_1_5_4_n29) );
  MUX2_X1 npu_inst_pe_1_5_4_U157 ( .A(npu_inst_pe_1_5_4_n28), .B(
        npu_inst_pe_1_5_4_n23), .S(npu_inst_pe_1_5_4_n8), .Z(
        npu_inst_pe_1_5_4_N94) );
  MUX2_X1 npu_inst_pe_1_5_4_U156 ( .A(npu_inst_pe_1_5_4_n25), .B(
        npu_inst_pe_1_5_4_n24), .S(npu_inst_pe_1_5_4_n6), .Z(
        npu_inst_pe_1_5_4_n28) );
  MUX2_X1 npu_inst_pe_1_5_4_U155 ( .A(npu_inst_pe_1_5_4_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_5_4_int_q_reg_v_1__1_), .S(npu_inst_pe_1_5_4_n4), .Z(
        npu_inst_pe_1_5_4_n25) );
  MUX2_X1 npu_inst_pe_1_5_4_U154 ( .A(npu_inst_pe_1_5_4_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_5_4_int_q_reg_v_3__1_), .S(npu_inst_pe_1_5_4_n4), .Z(
        npu_inst_pe_1_5_4_n24) );
  MUX2_X1 npu_inst_pe_1_5_4_U153 ( .A(npu_inst_pe_1_5_4_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_5_4_int_q_reg_v_5__1_), .S(npu_inst_pe_1_5_4_n4), .Z(
        npu_inst_pe_1_5_4_n23) );
  MUX2_X1 npu_inst_pe_1_5_4_U152 ( .A(npu_inst_pe_1_5_4_n22), .B(
        npu_inst_pe_1_5_4_n19), .S(npu_inst_pe_1_5_4_n8), .Z(
        npu_inst_int_data_x_5__4__1_) );
  MUX2_X1 npu_inst_pe_1_5_4_U151 ( .A(npu_inst_pe_1_5_4_n21), .B(
        npu_inst_pe_1_5_4_n20), .S(npu_inst_pe_1_5_4_n6), .Z(
        npu_inst_pe_1_5_4_n22) );
  MUX2_X1 npu_inst_pe_1_5_4_U150 ( .A(npu_inst_pe_1_5_4_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_5_4_int_q_reg_h_1__1_), .S(npu_inst_pe_1_5_4_n4), .Z(
        npu_inst_pe_1_5_4_n21) );
  MUX2_X1 npu_inst_pe_1_5_4_U149 ( .A(npu_inst_pe_1_5_4_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_5_4_int_q_reg_h_3__1_), .S(npu_inst_pe_1_5_4_n4), .Z(
        npu_inst_pe_1_5_4_n20) );
  MUX2_X1 npu_inst_pe_1_5_4_U148 ( .A(npu_inst_pe_1_5_4_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_5_4_int_q_reg_h_5__1_), .S(npu_inst_pe_1_5_4_n4), .Z(
        npu_inst_pe_1_5_4_n19) );
  MUX2_X1 npu_inst_pe_1_5_4_U147 ( .A(npu_inst_pe_1_5_4_n18), .B(
        npu_inst_pe_1_5_4_n15), .S(npu_inst_pe_1_5_4_n8), .Z(
        npu_inst_int_data_x_5__4__0_) );
  MUX2_X1 npu_inst_pe_1_5_4_U146 ( .A(npu_inst_pe_1_5_4_n17), .B(
        npu_inst_pe_1_5_4_n16), .S(npu_inst_pe_1_5_4_n6), .Z(
        npu_inst_pe_1_5_4_n18) );
  MUX2_X1 npu_inst_pe_1_5_4_U145 ( .A(npu_inst_pe_1_5_4_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_5_4_int_q_reg_h_1__0_), .S(npu_inst_pe_1_5_4_n4), .Z(
        npu_inst_pe_1_5_4_n17) );
  MUX2_X1 npu_inst_pe_1_5_4_U144 ( .A(npu_inst_pe_1_5_4_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_5_4_int_q_reg_h_3__0_), .S(npu_inst_pe_1_5_4_n4), .Z(
        npu_inst_pe_1_5_4_n16) );
  MUX2_X1 npu_inst_pe_1_5_4_U143 ( .A(npu_inst_pe_1_5_4_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_5_4_int_q_reg_h_5__0_), .S(npu_inst_pe_1_5_4_n4), .Z(
        npu_inst_pe_1_5_4_n15) );
  XOR2_X1 npu_inst_pe_1_5_4_U142 ( .A(npu_inst_pe_1_5_4_int_data_0_), .B(
        npu_inst_pe_1_5_4_int_q_acc_0_), .Z(npu_inst_pe_1_5_4_N73) );
  AND2_X1 npu_inst_pe_1_5_4_U141 ( .A1(npu_inst_pe_1_5_4_int_q_acc_0_), .A2(
        npu_inst_pe_1_5_4_int_data_0_), .ZN(npu_inst_pe_1_5_4_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_5_4_U140 ( .A(npu_inst_pe_1_5_4_int_q_acc_0_), .B(
        npu_inst_pe_1_5_4_n13), .ZN(npu_inst_pe_1_5_4_N65) );
  OR2_X1 npu_inst_pe_1_5_4_U139 ( .A1(npu_inst_pe_1_5_4_n13), .A2(
        npu_inst_pe_1_5_4_int_q_acc_0_), .ZN(npu_inst_pe_1_5_4_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_5_4_U138 ( .A(npu_inst_pe_1_5_4_int_q_acc_2_), .B(
        npu_inst_pe_1_5_4_add_69_carry_2_), .Z(npu_inst_pe_1_5_4_N75) );
  AND2_X1 npu_inst_pe_1_5_4_U137 ( .A1(npu_inst_pe_1_5_4_add_69_carry_2_), 
        .A2(npu_inst_pe_1_5_4_int_q_acc_2_), .ZN(
        npu_inst_pe_1_5_4_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_5_4_U136 ( .A(npu_inst_pe_1_5_4_int_q_acc_3_), .B(
        npu_inst_pe_1_5_4_add_69_carry_3_), .Z(npu_inst_pe_1_5_4_N76) );
  AND2_X1 npu_inst_pe_1_5_4_U135 ( .A1(npu_inst_pe_1_5_4_add_69_carry_3_), 
        .A2(npu_inst_pe_1_5_4_int_q_acc_3_), .ZN(
        npu_inst_pe_1_5_4_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_5_4_U134 ( .A(npu_inst_pe_1_5_4_int_q_acc_4_), .B(
        npu_inst_pe_1_5_4_add_69_carry_4_), .Z(npu_inst_pe_1_5_4_N77) );
  AND2_X1 npu_inst_pe_1_5_4_U133 ( .A1(npu_inst_pe_1_5_4_add_69_carry_4_), 
        .A2(npu_inst_pe_1_5_4_int_q_acc_4_), .ZN(
        npu_inst_pe_1_5_4_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_5_4_U132 ( .A(npu_inst_pe_1_5_4_int_q_acc_5_), .B(
        npu_inst_pe_1_5_4_add_69_carry_5_), .Z(npu_inst_pe_1_5_4_N78) );
  AND2_X1 npu_inst_pe_1_5_4_U131 ( .A1(npu_inst_pe_1_5_4_add_69_carry_5_), 
        .A2(npu_inst_pe_1_5_4_int_q_acc_5_), .ZN(
        npu_inst_pe_1_5_4_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_5_4_U130 ( .A(npu_inst_pe_1_5_4_int_q_acc_6_), .B(
        npu_inst_pe_1_5_4_add_69_carry_6_), .Z(npu_inst_pe_1_5_4_N79) );
  AND2_X1 npu_inst_pe_1_5_4_U129 ( .A1(npu_inst_pe_1_5_4_add_69_carry_6_), 
        .A2(npu_inst_pe_1_5_4_int_q_acc_6_), .ZN(
        npu_inst_pe_1_5_4_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_5_4_U128 ( .A(npu_inst_pe_1_5_4_int_q_acc_7_), .B(
        npu_inst_pe_1_5_4_add_69_carry_7_), .Z(npu_inst_pe_1_5_4_N80) );
  XNOR2_X1 npu_inst_pe_1_5_4_U127 ( .A(npu_inst_pe_1_5_4_sub_67_carry_2_), .B(
        npu_inst_pe_1_5_4_int_q_acc_2_), .ZN(npu_inst_pe_1_5_4_N67) );
  OR2_X1 npu_inst_pe_1_5_4_U126 ( .A1(npu_inst_pe_1_5_4_int_q_acc_2_), .A2(
        npu_inst_pe_1_5_4_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_5_4_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_5_4_U125 ( .A(npu_inst_pe_1_5_4_sub_67_carry_3_), .B(
        npu_inst_pe_1_5_4_int_q_acc_3_), .ZN(npu_inst_pe_1_5_4_N68) );
  OR2_X1 npu_inst_pe_1_5_4_U124 ( .A1(npu_inst_pe_1_5_4_int_q_acc_3_), .A2(
        npu_inst_pe_1_5_4_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_5_4_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_5_4_U123 ( .A(npu_inst_pe_1_5_4_sub_67_carry_4_), .B(
        npu_inst_pe_1_5_4_int_q_acc_4_), .ZN(npu_inst_pe_1_5_4_N69) );
  OR2_X1 npu_inst_pe_1_5_4_U122 ( .A1(npu_inst_pe_1_5_4_int_q_acc_4_), .A2(
        npu_inst_pe_1_5_4_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_5_4_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_5_4_U121 ( .A(npu_inst_pe_1_5_4_sub_67_carry_5_), .B(
        npu_inst_pe_1_5_4_int_q_acc_5_), .ZN(npu_inst_pe_1_5_4_N70) );
  OR2_X1 npu_inst_pe_1_5_4_U120 ( .A1(npu_inst_pe_1_5_4_int_q_acc_5_), .A2(
        npu_inst_pe_1_5_4_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_5_4_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_5_4_U119 ( .A(npu_inst_pe_1_5_4_sub_67_carry_6_), .B(
        npu_inst_pe_1_5_4_int_q_acc_6_), .ZN(npu_inst_pe_1_5_4_N71) );
  OR2_X1 npu_inst_pe_1_5_4_U118 ( .A1(npu_inst_pe_1_5_4_int_q_acc_6_), .A2(
        npu_inst_pe_1_5_4_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_5_4_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_5_4_U117 ( .A(npu_inst_pe_1_5_4_int_q_acc_7_), .B(
        npu_inst_pe_1_5_4_sub_67_carry_7_), .ZN(npu_inst_pe_1_5_4_N72) );
  INV_X1 npu_inst_pe_1_5_4_U116 ( .A(npu_inst_n76), .ZN(npu_inst_pe_1_5_4_n7)
         );
  INV_X1 npu_inst_pe_1_5_4_U115 ( .A(npu_inst_pe_1_5_4_n7), .ZN(
        npu_inst_pe_1_5_4_n6) );
  INV_X1 npu_inst_pe_1_5_4_U114 ( .A(npu_inst_n54), .ZN(npu_inst_pe_1_5_4_n3)
         );
  AOI22_X1 npu_inst_pe_1_5_4_U113 ( .A1(npu_inst_int_data_y_6__4__0_), .A2(
        npu_inst_pe_1_5_4_n58), .B1(npu_inst_pe_1_5_4_n119), .B2(
        npu_inst_pe_1_5_4_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_5_4_n57) );
  INV_X1 npu_inst_pe_1_5_4_U112 ( .A(npu_inst_pe_1_5_4_n57), .ZN(
        npu_inst_pe_1_5_4_n108) );
  AOI22_X1 npu_inst_pe_1_5_4_U111 ( .A1(npu_inst_int_data_y_6__4__0_), .A2(
        npu_inst_pe_1_5_4_n54), .B1(npu_inst_pe_1_5_4_n118), .B2(
        npu_inst_pe_1_5_4_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_5_4_n53) );
  INV_X1 npu_inst_pe_1_5_4_U110 ( .A(npu_inst_pe_1_5_4_n53), .ZN(
        npu_inst_pe_1_5_4_n109) );
  AOI22_X1 npu_inst_pe_1_5_4_U107 ( .A1(npu_inst_int_data_y_6__4__0_), .A2(
        npu_inst_pe_1_5_4_n50), .B1(npu_inst_pe_1_5_4_n117), .B2(
        npu_inst_pe_1_5_4_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_5_4_n49) );
  INV_X1 npu_inst_pe_1_5_4_U106 ( .A(npu_inst_pe_1_5_4_n49), .ZN(
        npu_inst_pe_1_5_4_n110) );
  AOI22_X1 npu_inst_pe_1_5_4_U105 ( .A1(npu_inst_int_data_y_6__4__0_), .A2(
        npu_inst_pe_1_5_4_n46), .B1(npu_inst_pe_1_5_4_n116), .B2(
        npu_inst_pe_1_5_4_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_5_4_n45) );
  INV_X1 npu_inst_pe_1_5_4_U104 ( .A(npu_inst_pe_1_5_4_n45), .ZN(
        npu_inst_pe_1_5_4_n111) );
  AOI22_X1 npu_inst_pe_1_5_4_U103 ( .A1(npu_inst_int_data_y_6__4__0_), .A2(
        npu_inst_pe_1_5_4_n42), .B1(npu_inst_pe_1_5_4_n115), .B2(
        npu_inst_pe_1_5_4_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_5_4_n41) );
  INV_X1 npu_inst_pe_1_5_4_U102 ( .A(npu_inst_pe_1_5_4_n41), .ZN(
        npu_inst_pe_1_5_4_n112) );
  AOI22_X1 npu_inst_pe_1_5_4_U101 ( .A1(npu_inst_int_data_y_6__4__1_), .A2(
        npu_inst_pe_1_5_4_n58), .B1(npu_inst_pe_1_5_4_n119), .B2(
        npu_inst_pe_1_5_4_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_5_4_n59) );
  INV_X1 npu_inst_pe_1_5_4_U100 ( .A(npu_inst_pe_1_5_4_n59), .ZN(
        npu_inst_pe_1_5_4_n102) );
  AOI22_X1 npu_inst_pe_1_5_4_U99 ( .A1(npu_inst_int_data_y_6__4__1_), .A2(
        npu_inst_pe_1_5_4_n54), .B1(npu_inst_pe_1_5_4_n118), .B2(
        npu_inst_pe_1_5_4_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_5_4_n55) );
  INV_X1 npu_inst_pe_1_5_4_U98 ( .A(npu_inst_pe_1_5_4_n55), .ZN(
        npu_inst_pe_1_5_4_n103) );
  AOI22_X1 npu_inst_pe_1_5_4_U97 ( .A1(npu_inst_int_data_y_6__4__1_), .A2(
        npu_inst_pe_1_5_4_n50), .B1(npu_inst_pe_1_5_4_n117), .B2(
        npu_inst_pe_1_5_4_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_5_4_n51) );
  INV_X1 npu_inst_pe_1_5_4_U96 ( .A(npu_inst_pe_1_5_4_n51), .ZN(
        npu_inst_pe_1_5_4_n104) );
  AOI22_X1 npu_inst_pe_1_5_4_U95 ( .A1(npu_inst_int_data_y_6__4__1_), .A2(
        npu_inst_pe_1_5_4_n46), .B1(npu_inst_pe_1_5_4_n116), .B2(
        npu_inst_pe_1_5_4_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_5_4_n47) );
  INV_X1 npu_inst_pe_1_5_4_U94 ( .A(npu_inst_pe_1_5_4_n47), .ZN(
        npu_inst_pe_1_5_4_n105) );
  AOI22_X1 npu_inst_pe_1_5_4_U93 ( .A1(npu_inst_int_data_y_6__4__1_), .A2(
        npu_inst_pe_1_5_4_n42), .B1(npu_inst_pe_1_5_4_n115), .B2(
        npu_inst_pe_1_5_4_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_5_4_n43) );
  INV_X1 npu_inst_pe_1_5_4_U92 ( .A(npu_inst_pe_1_5_4_n43), .ZN(
        npu_inst_pe_1_5_4_n106) );
  AOI22_X1 npu_inst_pe_1_5_4_U91 ( .A1(npu_inst_pe_1_5_4_n38), .A2(
        npu_inst_int_data_y_6__4__1_), .B1(npu_inst_pe_1_5_4_n114), .B2(
        npu_inst_pe_1_5_4_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_5_4_n39) );
  INV_X1 npu_inst_pe_1_5_4_U90 ( .A(npu_inst_pe_1_5_4_n39), .ZN(
        npu_inst_pe_1_5_4_n107) );
  AOI22_X1 npu_inst_pe_1_5_4_U89 ( .A1(npu_inst_pe_1_5_4_n38), .A2(
        npu_inst_int_data_y_6__4__0_), .B1(npu_inst_pe_1_5_4_n114), .B2(
        npu_inst_pe_1_5_4_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_5_4_n37) );
  INV_X1 npu_inst_pe_1_5_4_U88 ( .A(npu_inst_pe_1_5_4_n37), .ZN(
        npu_inst_pe_1_5_4_n113) );
  NAND2_X1 npu_inst_pe_1_5_4_U87 ( .A1(npu_inst_pe_1_5_4_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_5_4_n60), .ZN(npu_inst_pe_1_5_4_n74) );
  OAI21_X1 npu_inst_pe_1_5_4_U86 ( .B1(npu_inst_pe_1_5_4_n63), .B2(
        npu_inst_pe_1_5_4_n60), .A(npu_inst_pe_1_5_4_n74), .ZN(
        npu_inst_pe_1_5_4_n97) );
  NAND2_X1 npu_inst_pe_1_5_4_U85 ( .A1(npu_inst_pe_1_5_4_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_5_4_n60), .ZN(npu_inst_pe_1_5_4_n73) );
  OAI21_X1 npu_inst_pe_1_5_4_U84 ( .B1(npu_inst_pe_1_5_4_n61), .B2(
        npu_inst_pe_1_5_4_n60), .A(npu_inst_pe_1_5_4_n73), .ZN(
        npu_inst_pe_1_5_4_n96) );
  NAND2_X1 npu_inst_pe_1_5_4_U83 ( .A1(npu_inst_pe_1_5_4_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_5_4_n56), .ZN(npu_inst_pe_1_5_4_n72) );
  OAI21_X1 npu_inst_pe_1_5_4_U82 ( .B1(npu_inst_pe_1_5_4_n63), .B2(
        npu_inst_pe_1_5_4_n56), .A(npu_inst_pe_1_5_4_n72), .ZN(
        npu_inst_pe_1_5_4_n95) );
  NAND2_X1 npu_inst_pe_1_5_4_U81 ( .A1(npu_inst_pe_1_5_4_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_5_4_n56), .ZN(npu_inst_pe_1_5_4_n71) );
  OAI21_X1 npu_inst_pe_1_5_4_U80 ( .B1(npu_inst_pe_1_5_4_n61), .B2(
        npu_inst_pe_1_5_4_n56), .A(npu_inst_pe_1_5_4_n71), .ZN(
        npu_inst_pe_1_5_4_n94) );
  NAND2_X1 npu_inst_pe_1_5_4_U79 ( .A1(npu_inst_pe_1_5_4_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_5_4_n52), .ZN(npu_inst_pe_1_5_4_n70) );
  OAI21_X1 npu_inst_pe_1_5_4_U78 ( .B1(npu_inst_pe_1_5_4_n63), .B2(
        npu_inst_pe_1_5_4_n52), .A(npu_inst_pe_1_5_4_n70), .ZN(
        npu_inst_pe_1_5_4_n93) );
  NAND2_X1 npu_inst_pe_1_5_4_U77 ( .A1(npu_inst_pe_1_5_4_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_5_4_n52), .ZN(npu_inst_pe_1_5_4_n69) );
  OAI21_X1 npu_inst_pe_1_5_4_U76 ( .B1(npu_inst_pe_1_5_4_n61), .B2(
        npu_inst_pe_1_5_4_n52), .A(npu_inst_pe_1_5_4_n69), .ZN(
        npu_inst_pe_1_5_4_n92) );
  NAND2_X1 npu_inst_pe_1_5_4_U75 ( .A1(npu_inst_pe_1_5_4_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_5_4_n48), .ZN(npu_inst_pe_1_5_4_n68) );
  OAI21_X1 npu_inst_pe_1_5_4_U74 ( .B1(npu_inst_pe_1_5_4_n63), .B2(
        npu_inst_pe_1_5_4_n48), .A(npu_inst_pe_1_5_4_n68), .ZN(
        npu_inst_pe_1_5_4_n91) );
  NAND2_X1 npu_inst_pe_1_5_4_U73 ( .A1(npu_inst_pe_1_5_4_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_5_4_n48), .ZN(npu_inst_pe_1_5_4_n67) );
  OAI21_X1 npu_inst_pe_1_5_4_U72 ( .B1(npu_inst_pe_1_5_4_n61), .B2(
        npu_inst_pe_1_5_4_n48), .A(npu_inst_pe_1_5_4_n67), .ZN(
        npu_inst_pe_1_5_4_n90) );
  NAND2_X1 npu_inst_pe_1_5_4_U71 ( .A1(npu_inst_pe_1_5_4_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_5_4_n44), .ZN(npu_inst_pe_1_5_4_n66) );
  OAI21_X1 npu_inst_pe_1_5_4_U70 ( .B1(npu_inst_pe_1_5_4_n63), .B2(
        npu_inst_pe_1_5_4_n44), .A(npu_inst_pe_1_5_4_n66), .ZN(
        npu_inst_pe_1_5_4_n89) );
  NAND2_X1 npu_inst_pe_1_5_4_U69 ( .A1(npu_inst_pe_1_5_4_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_5_4_n44), .ZN(npu_inst_pe_1_5_4_n65) );
  OAI21_X1 npu_inst_pe_1_5_4_U68 ( .B1(npu_inst_pe_1_5_4_n61), .B2(
        npu_inst_pe_1_5_4_n44), .A(npu_inst_pe_1_5_4_n65), .ZN(
        npu_inst_pe_1_5_4_n88) );
  NAND2_X1 npu_inst_pe_1_5_4_U67 ( .A1(npu_inst_pe_1_5_4_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_5_4_n40), .ZN(npu_inst_pe_1_5_4_n64) );
  OAI21_X1 npu_inst_pe_1_5_4_U66 ( .B1(npu_inst_pe_1_5_4_n63), .B2(
        npu_inst_pe_1_5_4_n40), .A(npu_inst_pe_1_5_4_n64), .ZN(
        npu_inst_pe_1_5_4_n87) );
  NAND2_X1 npu_inst_pe_1_5_4_U65 ( .A1(npu_inst_pe_1_5_4_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_5_4_n40), .ZN(npu_inst_pe_1_5_4_n62) );
  OAI21_X1 npu_inst_pe_1_5_4_U64 ( .B1(npu_inst_pe_1_5_4_n61), .B2(
        npu_inst_pe_1_5_4_n40), .A(npu_inst_pe_1_5_4_n62), .ZN(
        npu_inst_pe_1_5_4_n86) );
  AND2_X1 npu_inst_pe_1_5_4_U63 ( .A1(npu_inst_pe_1_5_4_N93), .A2(npu_inst_n54), .ZN(npu_inst_int_data_y_5__4__0_) );
  AND2_X1 npu_inst_pe_1_5_4_U62 ( .A1(npu_inst_n54), .A2(npu_inst_pe_1_5_4_N94), .ZN(npu_inst_int_data_y_5__4__1_) );
  NOR3_X1 npu_inst_pe_1_5_4_U61 ( .A1(npu_inst_pe_1_5_4_n26), .A2(npu_inst_n54), .A3(npu_inst_int_ckg[19]), .ZN(npu_inst_pe_1_5_4_n85) );
  OR2_X1 npu_inst_pe_1_5_4_U60 ( .A1(npu_inst_pe_1_5_4_n85), .A2(
        npu_inst_pe_1_5_4_n2), .ZN(npu_inst_pe_1_5_4_N84) );
  AND2_X1 npu_inst_pe_1_5_4_U59 ( .A1(npu_inst_pe_1_5_4_int_q_acc_0_), .A2(
        npu_inst_pe_1_5_4_n1), .ZN(npu_inst_int_data_res_5__4__0_) );
  AND2_X1 npu_inst_pe_1_5_4_U58 ( .A1(npu_inst_pe_1_5_4_n2), .A2(
        npu_inst_pe_1_5_4_int_q_acc_7_), .ZN(npu_inst_int_data_res_5__4__7_)
         );
  AND2_X1 npu_inst_pe_1_5_4_U57 ( .A1(npu_inst_pe_1_5_4_int_q_acc_1_), .A2(
        npu_inst_pe_1_5_4_n1), .ZN(npu_inst_int_data_res_5__4__1_) );
  AND2_X1 npu_inst_pe_1_5_4_U56 ( .A1(npu_inst_pe_1_5_4_int_q_acc_2_), .A2(
        npu_inst_pe_1_5_4_n1), .ZN(npu_inst_int_data_res_5__4__2_) );
  AND2_X1 npu_inst_pe_1_5_4_U55 ( .A1(npu_inst_pe_1_5_4_int_q_acc_3_), .A2(
        npu_inst_pe_1_5_4_n2), .ZN(npu_inst_int_data_res_5__4__3_) );
  AND2_X1 npu_inst_pe_1_5_4_U54 ( .A1(npu_inst_pe_1_5_4_int_q_acc_4_), .A2(
        npu_inst_pe_1_5_4_n2), .ZN(npu_inst_int_data_res_5__4__4_) );
  AND2_X1 npu_inst_pe_1_5_4_U53 ( .A1(npu_inst_pe_1_5_4_int_q_acc_5_), .A2(
        npu_inst_pe_1_5_4_n2), .ZN(npu_inst_int_data_res_5__4__5_) );
  AND2_X1 npu_inst_pe_1_5_4_U52 ( .A1(npu_inst_pe_1_5_4_int_q_acc_6_), .A2(
        npu_inst_pe_1_5_4_n2), .ZN(npu_inst_int_data_res_5__4__6_) );
  AOI222_X1 npu_inst_pe_1_5_4_U51 ( .A1(npu_inst_int_data_res_6__4__0_), .A2(
        npu_inst_pe_1_5_4_n1), .B1(npu_inst_pe_1_5_4_N73), .B2(
        npu_inst_pe_1_5_4_n76), .C1(npu_inst_pe_1_5_4_N65), .C2(
        npu_inst_pe_1_5_4_n77), .ZN(npu_inst_pe_1_5_4_n84) );
  INV_X1 npu_inst_pe_1_5_4_U50 ( .A(npu_inst_pe_1_5_4_n84), .ZN(
        npu_inst_pe_1_5_4_n101) );
  AOI222_X1 npu_inst_pe_1_5_4_U49 ( .A1(npu_inst_int_data_res_6__4__7_), .A2(
        npu_inst_pe_1_5_4_n1), .B1(npu_inst_pe_1_5_4_N80), .B2(
        npu_inst_pe_1_5_4_n76), .C1(npu_inst_pe_1_5_4_N72), .C2(
        npu_inst_pe_1_5_4_n77), .ZN(npu_inst_pe_1_5_4_n75) );
  INV_X1 npu_inst_pe_1_5_4_U48 ( .A(npu_inst_pe_1_5_4_n75), .ZN(
        npu_inst_pe_1_5_4_n33) );
  AOI222_X1 npu_inst_pe_1_5_4_U47 ( .A1(npu_inst_int_data_res_6__4__1_), .A2(
        npu_inst_pe_1_5_4_n1), .B1(npu_inst_pe_1_5_4_N74), .B2(
        npu_inst_pe_1_5_4_n76), .C1(npu_inst_pe_1_5_4_N66), .C2(
        npu_inst_pe_1_5_4_n77), .ZN(npu_inst_pe_1_5_4_n83) );
  INV_X1 npu_inst_pe_1_5_4_U46 ( .A(npu_inst_pe_1_5_4_n83), .ZN(
        npu_inst_pe_1_5_4_n100) );
  AOI222_X1 npu_inst_pe_1_5_4_U45 ( .A1(npu_inst_int_data_res_6__4__2_), .A2(
        npu_inst_pe_1_5_4_n1), .B1(npu_inst_pe_1_5_4_N75), .B2(
        npu_inst_pe_1_5_4_n76), .C1(npu_inst_pe_1_5_4_N67), .C2(
        npu_inst_pe_1_5_4_n77), .ZN(npu_inst_pe_1_5_4_n82) );
  INV_X1 npu_inst_pe_1_5_4_U44 ( .A(npu_inst_pe_1_5_4_n82), .ZN(
        npu_inst_pe_1_5_4_n99) );
  AOI222_X1 npu_inst_pe_1_5_4_U43 ( .A1(npu_inst_int_data_res_6__4__3_), .A2(
        npu_inst_pe_1_5_4_n1), .B1(npu_inst_pe_1_5_4_N76), .B2(
        npu_inst_pe_1_5_4_n76), .C1(npu_inst_pe_1_5_4_N68), .C2(
        npu_inst_pe_1_5_4_n77), .ZN(npu_inst_pe_1_5_4_n81) );
  INV_X1 npu_inst_pe_1_5_4_U42 ( .A(npu_inst_pe_1_5_4_n81), .ZN(
        npu_inst_pe_1_5_4_n98) );
  AOI222_X1 npu_inst_pe_1_5_4_U41 ( .A1(npu_inst_int_data_res_6__4__4_), .A2(
        npu_inst_pe_1_5_4_n1), .B1(npu_inst_pe_1_5_4_N77), .B2(
        npu_inst_pe_1_5_4_n76), .C1(npu_inst_pe_1_5_4_N69), .C2(
        npu_inst_pe_1_5_4_n77), .ZN(npu_inst_pe_1_5_4_n80) );
  INV_X1 npu_inst_pe_1_5_4_U40 ( .A(npu_inst_pe_1_5_4_n80), .ZN(
        npu_inst_pe_1_5_4_n36) );
  AOI222_X1 npu_inst_pe_1_5_4_U39 ( .A1(npu_inst_int_data_res_6__4__5_), .A2(
        npu_inst_pe_1_5_4_n1), .B1(npu_inst_pe_1_5_4_N78), .B2(
        npu_inst_pe_1_5_4_n76), .C1(npu_inst_pe_1_5_4_N70), .C2(
        npu_inst_pe_1_5_4_n77), .ZN(npu_inst_pe_1_5_4_n79) );
  INV_X1 npu_inst_pe_1_5_4_U38 ( .A(npu_inst_pe_1_5_4_n79), .ZN(
        npu_inst_pe_1_5_4_n35) );
  AOI222_X1 npu_inst_pe_1_5_4_U37 ( .A1(npu_inst_int_data_res_6__4__6_), .A2(
        npu_inst_pe_1_5_4_n1), .B1(npu_inst_pe_1_5_4_N79), .B2(
        npu_inst_pe_1_5_4_n76), .C1(npu_inst_pe_1_5_4_N71), .C2(
        npu_inst_pe_1_5_4_n77), .ZN(npu_inst_pe_1_5_4_n78) );
  INV_X1 npu_inst_pe_1_5_4_U36 ( .A(npu_inst_pe_1_5_4_n78), .ZN(
        npu_inst_pe_1_5_4_n34) );
  INV_X1 npu_inst_pe_1_5_4_U35 ( .A(npu_inst_pe_1_5_4_int_data_1_), .ZN(
        npu_inst_pe_1_5_4_n14) );
  AND2_X1 npu_inst_pe_1_5_4_U34 ( .A1(npu_inst_int_data_x_5__4__1_), .A2(
        npu_inst_pe_1_5_4_int_q_weight_1_), .ZN(npu_inst_pe_1_5_4_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_5_4_U33 ( .A1(npu_inst_int_data_x_5__4__0_), .A2(
        npu_inst_pe_1_5_4_int_q_weight_1_), .ZN(npu_inst_pe_1_5_4_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_5_4_U32 ( .A1(npu_inst_n54), .A2(
        npu_inst_int_data_y_6__4__1_), .B1(npu_inst_pe_1_5_4_n3), .B2(
        npu_inst_int_data_x_5__5__1_), .ZN(npu_inst_pe_1_5_4_n63) );
  AOI22_X1 npu_inst_pe_1_5_4_U31 ( .A1(npu_inst_n54), .A2(
        npu_inst_int_data_y_6__4__0_), .B1(npu_inst_pe_1_5_4_n3), .B2(
        npu_inst_int_data_x_5__5__0_), .ZN(npu_inst_pe_1_5_4_n61) );
  INV_X1 npu_inst_pe_1_5_4_U30 ( .A(npu_inst_pe_1_5_4_int_data_0_), .ZN(
        npu_inst_pe_1_5_4_n13) );
  INV_X1 npu_inst_pe_1_5_4_U29 ( .A(npu_inst_n68), .ZN(npu_inst_pe_1_5_4_n5)
         );
  OR3_X1 npu_inst_pe_1_5_4_U28 ( .A1(npu_inst_pe_1_5_4_n6), .A2(
        npu_inst_pe_1_5_4_n8), .A3(npu_inst_pe_1_5_4_n5), .ZN(
        npu_inst_pe_1_5_4_n56) );
  OR3_X1 npu_inst_pe_1_5_4_U27 ( .A1(npu_inst_pe_1_5_4_n5), .A2(
        npu_inst_pe_1_5_4_n8), .A3(npu_inst_pe_1_5_4_n7), .ZN(
        npu_inst_pe_1_5_4_n48) );
  INV_X1 npu_inst_pe_1_5_4_U26 ( .A(npu_inst_pe_1_5_4_n5), .ZN(
        npu_inst_pe_1_5_4_n4) );
  OR3_X1 npu_inst_pe_1_5_4_U25 ( .A1(npu_inst_pe_1_5_4_n4), .A2(
        npu_inst_pe_1_5_4_n8), .A3(npu_inst_pe_1_5_4_n7), .ZN(
        npu_inst_pe_1_5_4_n52) );
  OR3_X1 npu_inst_pe_1_5_4_U24 ( .A1(npu_inst_pe_1_5_4_n6), .A2(
        npu_inst_pe_1_5_4_n8), .A3(npu_inst_pe_1_5_4_n4), .ZN(
        npu_inst_pe_1_5_4_n60) );
  NOR2_X1 npu_inst_pe_1_5_4_U23 ( .A1(npu_inst_pe_1_5_4_n60), .A2(
        npu_inst_pe_1_5_4_n3), .ZN(npu_inst_pe_1_5_4_n58) );
  NOR2_X1 npu_inst_pe_1_5_4_U22 ( .A1(npu_inst_pe_1_5_4_n56), .A2(
        npu_inst_pe_1_5_4_n3), .ZN(npu_inst_pe_1_5_4_n54) );
  NOR2_X1 npu_inst_pe_1_5_4_U21 ( .A1(npu_inst_pe_1_5_4_n52), .A2(
        npu_inst_pe_1_5_4_n3), .ZN(npu_inst_pe_1_5_4_n50) );
  NOR2_X1 npu_inst_pe_1_5_4_U20 ( .A1(npu_inst_pe_1_5_4_n48), .A2(
        npu_inst_pe_1_5_4_n3), .ZN(npu_inst_pe_1_5_4_n46) );
  NOR2_X1 npu_inst_pe_1_5_4_U19 ( .A1(npu_inst_pe_1_5_4_n40), .A2(
        npu_inst_pe_1_5_4_n3), .ZN(npu_inst_pe_1_5_4_n38) );
  NOR2_X1 npu_inst_pe_1_5_4_U18 ( .A1(npu_inst_pe_1_5_4_n44), .A2(
        npu_inst_pe_1_5_4_n3), .ZN(npu_inst_pe_1_5_4_n42) );
  BUF_X1 npu_inst_pe_1_5_4_U17 ( .A(npu_inst_n96), .Z(npu_inst_pe_1_5_4_n8) );
  INV_X1 npu_inst_pe_1_5_4_U16 ( .A(npu_inst_n123), .ZN(npu_inst_pe_1_5_4_n12)
         );
  INV_X1 npu_inst_pe_1_5_4_U15 ( .A(npu_inst_pe_1_5_4_n38), .ZN(
        npu_inst_pe_1_5_4_n114) );
  INV_X1 npu_inst_pe_1_5_4_U14 ( .A(npu_inst_pe_1_5_4_n58), .ZN(
        npu_inst_pe_1_5_4_n119) );
  INV_X1 npu_inst_pe_1_5_4_U13 ( .A(npu_inst_pe_1_5_4_n54), .ZN(
        npu_inst_pe_1_5_4_n118) );
  INV_X1 npu_inst_pe_1_5_4_U12 ( .A(npu_inst_pe_1_5_4_n50), .ZN(
        npu_inst_pe_1_5_4_n117) );
  INV_X1 npu_inst_pe_1_5_4_U11 ( .A(npu_inst_pe_1_5_4_n46), .ZN(
        npu_inst_pe_1_5_4_n116) );
  INV_X1 npu_inst_pe_1_5_4_U10 ( .A(npu_inst_pe_1_5_4_n42), .ZN(
        npu_inst_pe_1_5_4_n115) );
  BUF_X1 npu_inst_pe_1_5_4_U9 ( .A(npu_inst_n16), .Z(npu_inst_pe_1_5_4_n2) );
  BUF_X1 npu_inst_pe_1_5_4_U8 ( .A(npu_inst_n16), .Z(npu_inst_pe_1_5_4_n1) );
  BUF_X1 npu_inst_pe_1_5_4_U7 ( .A(npu_inst_pe_1_5_4_n12), .Z(
        npu_inst_pe_1_5_4_n11) );
  BUF_X1 npu_inst_pe_1_5_4_U6 ( .A(npu_inst_pe_1_5_4_n12), .Z(
        npu_inst_pe_1_5_4_n10) );
  BUF_X1 npu_inst_pe_1_5_4_U5 ( .A(npu_inst_pe_1_5_4_n12), .Z(
        npu_inst_pe_1_5_4_n9) );
  NOR2_X1 npu_inst_pe_1_5_4_U4 ( .A1(npu_inst_pe_1_5_4_int_q_weight_0_), .A2(
        npu_inst_pe_1_5_4_n1), .ZN(npu_inst_pe_1_5_4_n76) );
  NOR2_X1 npu_inst_pe_1_5_4_U3 ( .A1(npu_inst_pe_1_5_4_n27), .A2(
        npu_inst_pe_1_5_4_n1), .ZN(npu_inst_pe_1_5_4_n77) );
  FA_X1 npu_inst_pe_1_5_4_sub_67_U2_1 ( .A(npu_inst_pe_1_5_4_int_q_acc_1_), 
        .B(npu_inst_pe_1_5_4_n14), .CI(npu_inst_pe_1_5_4_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_5_4_sub_67_carry_2_), .S(npu_inst_pe_1_5_4_N66) );
  FA_X1 npu_inst_pe_1_5_4_add_69_U1_1 ( .A(npu_inst_pe_1_5_4_int_q_acc_1_), 
        .B(npu_inst_pe_1_5_4_int_data_1_), .CI(
        npu_inst_pe_1_5_4_add_69_carry_1_), .CO(
        npu_inst_pe_1_5_4_add_69_carry_2_), .S(npu_inst_pe_1_5_4_N74) );
  NAND3_X1 npu_inst_pe_1_5_4_U109 ( .A1(npu_inst_pe_1_5_4_n5), .A2(
        npu_inst_pe_1_5_4_n7), .A3(npu_inst_pe_1_5_4_n8), .ZN(
        npu_inst_pe_1_5_4_n44) );
  NAND3_X1 npu_inst_pe_1_5_4_U108 ( .A1(npu_inst_pe_1_5_4_n4), .A2(
        npu_inst_pe_1_5_4_n7), .A3(npu_inst_pe_1_5_4_n8), .ZN(
        npu_inst_pe_1_5_4_n40) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_5_4_n34), .CK(
        npu_inst_pe_1_5_4_net3550), .RN(npu_inst_pe_1_5_4_n9), .Q(
        npu_inst_pe_1_5_4_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_5_4_n35), .CK(
        npu_inst_pe_1_5_4_net3550), .RN(npu_inst_pe_1_5_4_n9), .Q(
        npu_inst_pe_1_5_4_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_5_4_n36), .CK(
        npu_inst_pe_1_5_4_net3550), .RN(npu_inst_pe_1_5_4_n9), .Q(
        npu_inst_pe_1_5_4_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_5_4_n98), .CK(
        npu_inst_pe_1_5_4_net3550), .RN(npu_inst_pe_1_5_4_n9), .Q(
        npu_inst_pe_1_5_4_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_5_4_n99), .CK(
        npu_inst_pe_1_5_4_net3550), .RN(npu_inst_pe_1_5_4_n9), .Q(
        npu_inst_pe_1_5_4_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_5_4_n100), 
        .CK(npu_inst_pe_1_5_4_net3550), .RN(npu_inst_pe_1_5_4_n9), .Q(
        npu_inst_pe_1_5_4_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_5_4_n33), .CK(
        npu_inst_pe_1_5_4_net3550), .RN(npu_inst_pe_1_5_4_n9), .Q(
        npu_inst_pe_1_5_4_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_5_4_n101), 
        .CK(npu_inst_pe_1_5_4_net3550), .RN(npu_inst_pe_1_5_4_n9), .Q(
        npu_inst_pe_1_5_4_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_weight_reg_0_ ( .D(npu_inst_n109), .CK(
        npu_inst_pe_1_5_4_net3556), .RN(npu_inst_pe_1_5_4_n9), .Q(
        npu_inst_pe_1_5_4_int_q_weight_0_), .QN(npu_inst_pe_1_5_4_n27) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_weight_reg_1_ ( .D(npu_inst_n115), .CK(
        npu_inst_pe_1_5_4_net3556), .RN(npu_inst_pe_1_5_4_n9), .Q(
        npu_inst_pe_1_5_4_int_q_weight_1_), .QN(npu_inst_pe_1_5_4_n26) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_5_4_n113), 
        .CK(npu_inst_pe_1_5_4_net3556), .RN(npu_inst_pe_1_5_4_n9), .Q(
        npu_inst_pe_1_5_4_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_5_4_n107), 
        .CK(npu_inst_pe_1_5_4_net3556), .RN(npu_inst_pe_1_5_4_n9), .Q(
        npu_inst_pe_1_5_4_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_5_4_n112), 
        .CK(npu_inst_pe_1_5_4_net3556), .RN(npu_inst_pe_1_5_4_n10), .Q(
        npu_inst_pe_1_5_4_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_5_4_n106), 
        .CK(npu_inst_pe_1_5_4_net3556), .RN(npu_inst_pe_1_5_4_n10), .Q(
        npu_inst_pe_1_5_4_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_5_4_n111), 
        .CK(npu_inst_pe_1_5_4_net3556), .RN(npu_inst_pe_1_5_4_n10), .Q(
        npu_inst_pe_1_5_4_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_5_4_n105), 
        .CK(npu_inst_pe_1_5_4_net3556), .RN(npu_inst_pe_1_5_4_n10), .Q(
        npu_inst_pe_1_5_4_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_5_4_n110), 
        .CK(npu_inst_pe_1_5_4_net3556), .RN(npu_inst_pe_1_5_4_n10), .Q(
        npu_inst_pe_1_5_4_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_5_4_n104), 
        .CK(npu_inst_pe_1_5_4_net3556), .RN(npu_inst_pe_1_5_4_n10), .Q(
        npu_inst_pe_1_5_4_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_5_4_n109), 
        .CK(npu_inst_pe_1_5_4_net3556), .RN(npu_inst_pe_1_5_4_n10), .Q(
        npu_inst_pe_1_5_4_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_5_4_n103), 
        .CK(npu_inst_pe_1_5_4_net3556), .RN(npu_inst_pe_1_5_4_n10), .Q(
        npu_inst_pe_1_5_4_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_5_4_n108), 
        .CK(npu_inst_pe_1_5_4_net3556), .RN(npu_inst_pe_1_5_4_n10), .Q(
        npu_inst_pe_1_5_4_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_5_4_n102), 
        .CK(npu_inst_pe_1_5_4_net3556), .RN(npu_inst_pe_1_5_4_n10), .Q(
        npu_inst_pe_1_5_4_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_5_4_n86), 
        .CK(npu_inst_pe_1_5_4_net3556), .RN(npu_inst_pe_1_5_4_n10), .Q(
        npu_inst_pe_1_5_4_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_5_4_n87), 
        .CK(npu_inst_pe_1_5_4_net3556), .RN(npu_inst_pe_1_5_4_n10), .Q(
        npu_inst_pe_1_5_4_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_5_4_n88), 
        .CK(npu_inst_pe_1_5_4_net3556), .RN(npu_inst_pe_1_5_4_n11), .Q(
        npu_inst_pe_1_5_4_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_5_4_n89), 
        .CK(npu_inst_pe_1_5_4_net3556), .RN(npu_inst_pe_1_5_4_n11), .Q(
        npu_inst_pe_1_5_4_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_5_4_n90), 
        .CK(npu_inst_pe_1_5_4_net3556), .RN(npu_inst_pe_1_5_4_n11), .Q(
        npu_inst_pe_1_5_4_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_5_4_n91), 
        .CK(npu_inst_pe_1_5_4_net3556), .RN(npu_inst_pe_1_5_4_n11), .Q(
        npu_inst_pe_1_5_4_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_5_4_n92), 
        .CK(npu_inst_pe_1_5_4_net3556), .RN(npu_inst_pe_1_5_4_n11), .Q(
        npu_inst_pe_1_5_4_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_5_4_n93), 
        .CK(npu_inst_pe_1_5_4_net3556), .RN(npu_inst_pe_1_5_4_n11), .Q(
        npu_inst_pe_1_5_4_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_5_4_n94), 
        .CK(npu_inst_pe_1_5_4_net3556), .RN(npu_inst_pe_1_5_4_n11), .Q(
        npu_inst_pe_1_5_4_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_5_4_n95), 
        .CK(npu_inst_pe_1_5_4_net3556), .RN(npu_inst_pe_1_5_4_n11), .Q(
        npu_inst_pe_1_5_4_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_5_4_n96), 
        .CK(npu_inst_pe_1_5_4_net3556), .RN(npu_inst_pe_1_5_4_n11), .Q(
        npu_inst_pe_1_5_4_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_5_4_n97), 
        .CK(npu_inst_pe_1_5_4_net3556), .RN(npu_inst_pe_1_5_4_n11), .Q(
        npu_inst_pe_1_5_4_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_5_4_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_5_4_N84), .SE(1'b0), .GCK(npu_inst_pe_1_5_4_net3550) );
  CLKGATETST_X1 npu_inst_pe_1_5_4_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n62), .SE(1'b0), .GCK(npu_inst_pe_1_5_4_net3556) );
  MUX2_X1 npu_inst_pe_1_5_5_U162 ( .A(npu_inst_pe_1_5_5_n32), .B(
        npu_inst_pe_1_5_5_n29), .S(npu_inst_pe_1_5_5_n8), .Z(
        npu_inst_pe_1_5_5_N93) );
  MUX2_X1 npu_inst_pe_1_5_5_U161 ( .A(npu_inst_pe_1_5_5_n31), .B(
        npu_inst_pe_1_5_5_n30), .S(npu_inst_pe_1_5_5_n6), .Z(
        npu_inst_pe_1_5_5_n32) );
  MUX2_X1 npu_inst_pe_1_5_5_U160 ( .A(npu_inst_pe_1_5_5_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_5_5_int_q_reg_v_1__0_), .S(npu_inst_pe_1_5_5_n4), .Z(
        npu_inst_pe_1_5_5_n31) );
  MUX2_X1 npu_inst_pe_1_5_5_U159 ( .A(npu_inst_pe_1_5_5_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_5_5_int_q_reg_v_3__0_), .S(npu_inst_pe_1_5_5_n4), .Z(
        npu_inst_pe_1_5_5_n30) );
  MUX2_X1 npu_inst_pe_1_5_5_U158 ( .A(npu_inst_pe_1_5_5_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_5_5_int_q_reg_v_5__0_), .S(npu_inst_pe_1_5_5_n4), .Z(
        npu_inst_pe_1_5_5_n29) );
  MUX2_X1 npu_inst_pe_1_5_5_U157 ( .A(npu_inst_pe_1_5_5_n28), .B(
        npu_inst_pe_1_5_5_n23), .S(npu_inst_pe_1_5_5_n8), .Z(
        npu_inst_pe_1_5_5_N94) );
  MUX2_X1 npu_inst_pe_1_5_5_U156 ( .A(npu_inst_pe_1_5_5_n25), .B(
        npu_inst_pe_1_5_5_n24), .S(npu_inst_pe_1_5_5_n6), .Z(
        npu_inst_pe_1_5_5_n28) );
  MUX2_X1 npu_inst_pe_1_5_5_U155 ( .A(npu_inst_pe_1_5_5_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_5_5_int_q_reg_v_1__1_), .S(npu_inst_pe_1_5_5_n4), .Z(
        npu_inst_pe_1_5_5_n25) );
  MUX2_X1 npu_inst_pe_1_5_5_U154 ( .A(npu_inst_pe_1_5_5_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_5_5_int_q_reg_v_3__1_), .S(npu_inst_pe_1_5_5_n4), .Z(
        npu_inst_pe_1_5_5_n24) );
  MUX2_X1 npu_inst_pe_1_5_5_U153 ( .A(npu_inst_pe_1_5_5_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_5_5_int_q_reg_v_5__1_), .S(npu_inst_pe_1_5_5_n4), .Z(
        npu_inst_pe_1_5_5_n23) );
  MUX2_X1 npu_inst_pe_1_5_5_U152 ( .A(npu_inst_pe_1_5_5_n22), .B(
        npu_inst_pe_1_5_5_n19), .S(npu_inst_pe_1_5_5_n8), .Z(
        npu_inst_int_data_x_5__5__1_) );
  MUX2_X1 npu_inst_pe_1_5_5_U151 ( .A(npu_inst_pe_1_5_5_n21), .B(
        npu_inst_pe_1_5_5_n20), .S(npu_inst_pe_1_5_5_n6), .Z(
        npu_inst_pe_1_5_5_n22) );
  MUX2_X1 npu_inst_pe_1_5_5_U150 ( .A(npu_inst_pe_1_5_5_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_5_5_int_q_reg_h_1__1_), .S(npu_inst_pe_1_5_5_n4), .Z(
        npu_inst_pe_1_5_5_n21) );
  MUX2_X1 npu_inst_pe_1_5_5_U149 ( .A(npu_inst_pe_1_5_5_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_5_5_int_q_reg_h_3__1_), .S(npu_inst_pe_1_5_5_n4), .Z(
        npu_inst_pe_1_5_5_n20) );
  MUX2_X1 npu_inst_pe_1_5_5_U148 ( .A(npu_inst_pe_1_5_5_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_5_5_int_q_reg_h_5__1_), .S(npu_inst_pe_1_5_5_n4), .Z(
        npu_inst_pe_1_5_5_n19) );
  MUX2_X1 npu_inst_pe_1_5_5_U147 ( .A(npu_inst_pe_1_5_5_n18), .B(
        npu_inst_pe_1_5_5_n15), .S(npu_inst_pe_1_5_5_n8), .Z(
        npu_inst_int_data_x_5__5__0_) );
  MUX2_X1 npu_inst_pe_1_5_5_U146 ( .A(npu_inst_pe_1_5_5_n17), .B(
        npu_inst_pe_1_5_5_n16), .S(npu_inst_pe_1_5_5_n6), .Z(
        npu_inst_pe_1_5_5_n18) );
  MUX2_X1 npu_inst_pe_1_5_5_U145 ( .A(npu_inst_pe_1_5_5_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_5_5_int_q_reg_h_1__0_), .S(npu_inst_pe_1_5_5_n4), .Z(
        npu_inst_pe_1_5_5_n17) );
  MUX2_X1 npu_inst_pe_1_5_5_U144 ( .A(npu_inst_pe_1_5_5_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_5_5_int_q_reg_h_3__0_), .S(npu_inst_pe_1_5_5_n4), .Z(
        npu_inst_pe_1_5_5_n16) );
  MUX2_X1 npu_inst_pe_1_5_5_U143 ( .A(npu_inst_pe_1_5_5_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_5_5_int_q_reg_h_5__0_), .S(npu_inst_pe_1_5_5_n4), .Z(
        npu_inst_pe_1_5_5_n15) );
  XOR2_X1 npu_inst_pe_1_5_5_U142 ( .A(npu_inst_pe_1_5_5_int_data_0_), .B(
        npu_inst_pe_1_5_5_int_q_acc_0_), .Z(npu_inst_pe_1_5_5_N73) );
  AND2_X1 npu_inst_pe_1_5_5_U141 ( .A1(npu_inst_pe_1_5_5_int_q_acc_0_), .A2(
        npu_inst_pe_1_5_5_int_data_0_), .ZN(npu_inst_pe_1_5_5_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_5_5_U140 ( .A(npu_inst_pe_1_5_5_int_q_acc_0_), .B(
        npu_inst_pe_1_5_5_n13), .ZN(npu_inst_pe_1_5_5_N65) );
  OR2_X1 npu_inst_pe_1_5_5_U139 ( .A1(npu_inst_pe_1_5_5_n13), .A2(
        npu_inst_pe_1_5_5_int_q_acc_0_), .ZN(npu_inst_pe_1_5_5_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_5_5_U138 ( .A(npu_inst_pe_1_5_5_int_q_acc_2_), .B(
        npu_inst_pe_1_5_5_add_69_carry_2_), .Z(npu_inst_pe_1_5_5_N75) );
  AND2_X1 npu_inst_pe_1_5_5_U137 ( .A1(npu_inst_pe_1_5_5_add_69_carry_2_), 
        .A2(npu_inst_pe_1_5_5_int_q_acc_2_), .ZN(
        npu_inst_pe_1_5_5_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_5_5_U136 ( .A(npu_inst_pe_1_5_5_int_q_acc_3_), .B(
        npu_inst_pe_1_5_5_add_69_carry_3_), .Z(npu_inst_pe_1_5_5_N76) );
  AND2_X1 npu_inst_pe_1_5_5_U135 ( .A1(npu_inst_pe_1_5_5_add_69_carry_3_), 
        .A2(npu_inst_pe_1_5_5_int_q_acc_3_), .ZN(
        npu_inst_pe_1_5_5_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_5_5_U134 ( .A(npu_inst_pe_1_5_5_int_q_acc_4_), .B(
        npu_inst_pe_1_5_5_add_69_carry_4_), .Z(npu_inst_pe_1_5_5_N77) );
  AND2_X1 npu_inst_pe_1_5_5_U133 ( .A1(npu_inst_pe_1_5_5_add_69_carry_4_), 
        .A2(npu_inst_pe_1_5_5_int_q_acc_4_), .ZN(
        npu_inst_pe_1_5_5_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_5_5_U132 ( .A(npu_inst_pe_1_5_5_int_q_acc_5_), .B(
        npu_inst_pe_1_5_5_add_69_carry_5_), .Z(npu_inst_pe_1_5_5_N78) );
  AND2_X1 npu_inst_pe_1_5_5_U131 ( .A1(npu_inst_pe_1_5_5_add_69_carry_5_), 
        .A2(npu_inst_pe_1_5_5_int_q_acc_5_), .ZN(
        npu_inst_pe_1_5_5_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_5_5_U130 ( .A(npu_inst_pe_1_5_5_int_q_acc_6_), .B(
        npu_inst_pe_1_5_5_add_69_carry_6_), .Z(npu_inst_pe_1_5_5_N79) );
  AND2_X1 npu_inst_pe_1_5_5_U129 ( .A1(npu_inst_pe_1_5_5_add_69_carry_6_), 
        .A2(npu_inst_pe_1_5_5_int_q_acc_6_), .ZN(
        npu_inst_pe_1_5_5_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_5_5_U128 ( .A(npu_inst_pe_1_5_5_int_q_acc_7_), .B(
        npu_inst_pe_1_5_5_add_69_carry_7_), .Z(npu_inst_pe_1_5_5_N80) );
  XNOR2_X1 npu_inst_pe_1_5_5_U127 ( .A(npu_inst_pe_1_5_5_sub_67_carry_2_), .B(
        npu_inst_pe_1_5_5_int_q_acc_2_), .ZN(npu_inst_pe_1_5_5_N67) );
  OR2_X1 npu_inst_pe_1_5_5_U126 ( .A1(npu_inst_pe_1_5_5_int_q_acc_2_), .A2(
        npu_inst_pe_1_5_5_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_5_5_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_5_5_U125 ( .A(npu_inst_pe_1_5_5_sub_67_carry_3_), .B(
        npu_inst_pe_1_5_5_int_q_acc_3_), .ZN(npu_inst_pe_1_5_5_N68) );
  OR2_X1 npu_inst_pe_1_5_5_U124 ( .A1(npu_inst_pe_1_5_5_int_q_acc_3_), .A2(
        npu_inst_pe_1_5_5_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_5_5_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_5_5_U123 ( .A(npu_inst_pe_1_5_5_sub_67_carry_4_), .B(
        npu_inst_pe_1_5_5_int_q_acc_4_), .ZN(npu_inst_pe_1_5_5_N69) );
  OR2_X1 npu_inst_pe_1_5_5_U122 ( .A1(npu_inst_pe_1_5_5_int_q_acc_4_), .A2(
        npu_inst_pe_1_5_5_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_5_5_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_5_5_U121 ( .A(npu_inst_pe_1_5_5_sub_67_carry_5_), .B(
        npu_inst_pe_1_5_5_int_q_acc_5_), .ZN(npu_inst_pe_1_5_5_N70) );
  OR2_X1 npu_inst_pe_1_5_5_U120 ( .A1(npu_inst_pe_1_5_5_int_q_acc_5_), .A2(
        npu_inst_pe_1_5_5_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_5_5_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_5_5_U119 ( .A(npu_inst_pe_1_5_5_sub_67_carry_6_), .B(
        npu_inst_pe_1_5_5_int_q_acc_6_), .ZN(npu_inst_pe_1_5_5_N71) );
  OR2_X1 npu_inst_pe_1_5_5_U118 ( .A1(npu_inst_pe_1_5_5_int_q_acc_6_), .A2(
        npu_inst_pe_1_5_5_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_5_5_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_5_5_U117 ( .A(npu_inst_pe_1_5_5_int_q_acc_7_), .B(
        npu_inst_pe_1_5_5_sub_67_carry_7_), .ZN(npu_inst_pe_1_5_5_N72) );
  INV_X1 npu_inst_pe_1_5_5_U116 ( .A(npu_inst_n76), .ZN(npu_inst_pe_1_5_5_n7)
         );
  INV_X1 npu_inst_pe_1_5_5_U115 ( .A(npu_inst_pe_1_5_5_n7), .ZN(
        npu_inst_pe_1_5_5_n6) );
  INV_X1 npu_inst_pe_1_5_5_U114 ( .A(npu_inst_n54), .ZN(npu_inst_pe_1_5_5_n3)
         );
  AOI22_X1 npu_inst_pe_1_5_5_U113 ( .A1(npu_inst_int_data_y_6__5__0_), .A2(
        npu_inst_pe_1_5_5_n58), .B1(npu_inst_pe_1_5_5_n119), .B2(
        npu_inst_pe_1_5_5_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_5_5_n57) );
  INV_X1 npu_inst_pe_1_5_5_U112 ( .A(npu_inst_pe_1_5_5_n57), .ZN(
        npu_inst_pe_1_5_5_n108) );
  AOI22_X1 npu_inst_pe_1_5_5_U111 ( .A1(npu_inst_int_data_y_6__5__0_), .A2(
        npu_inst_pe_1_5_5_n54), .B1(npu_inst_pe_1_5_5_n118), .B2(
        npu_inst_pe_1_5_5_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_5_5_n53) );
  INV_X1 npu_inst_pe_1_5_5_U110 ( .A(npu_inst_pe_1_5_5_n53), .ZN(
        npu_inst_pe_1_5_5_n109) );
  AOI22_X1 npu_inst_pe_1_5_5_U107 ( .A1(npu_inst_int_data_y_6__5__0_), .A2(
        npu_inst_pe_1_5_5_n50), .B1(npu_inst_pe_1_5_5_n117), .B2(
        npu_inst_pe_1_5_5_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_5_5_n49) );
  INV_X1 npu_inst_pe_1_5_5_U106 ( .A(npu_inst_pe_1_5_5_n49), .ZN(
        npu_inst_pe_1_5_5_n110) );
  AOI22_X1 npu_inst_pe_1_5_5_U105 ( .A1(npu_inst_int_data_y_6__5__0_), .A2(
        npu_inst_pe_1_5_5_n46), .B1(npu_inst_pe_1_5_5_n116), .B2(
        npu_inst_pe_1_5_5_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_5_5_n45) );
  INV_X1 npu_inst_pe_1_5_5_U104 ( .A(npu_inst_pe_1_5_5_n45), .ZN(
        npu_inst_pe_1_5_5_n111) );
  AOI22_X1 npu_inst_pe_1_5_5_U103 ( .A1(npu_inst_int_data_y_6__5__0_), .A2(
        npu_inst_pe_1_5_5_n42), .B1(npu_inst_pe_1_5_5_n115), .B2(
        npu_inst_pe_1_5_5_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_5_5_n41) );
  INV_X1 npu_inst_pe_1_5_5_U102 ( .A(npu_inst_pe_1_5_5_n41), .ZN(
        npu_inst_pe_1_5_5_n112) );
  AOI22_X1 npu_inst_pe_1_5_5_U101 ( .A1(npu_inst_int_data_y_6__5__1_), .A2(
        npu_inst_pe_1_5_5_n58), .B1(npu_inst_pe_1_5_5_n119), .B2(
        npu_inst_pe_1_5_5_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_5_5_n59) );
  INV_X1 npu_inst_pe_1_5_5_U100 ( .A(npu_inst_pe_1_5_5_n59), .ZN(
        npu_inst_pe_1_5_5_n102) );
  AOI22_X1 npu_inst_pe_1_5_5_U99 ( .A1(npu_inst_int_data_y_6__5__1_), .A2(
        npu_inst_pe_1_5_5_n54), .B1(npu_inst_pe_1_5_5_n118), .B2(
        npu_inst_pe_1_5_5_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_5_5_n55) );
  INV_X1 npu_inst_pe_1_5_5_U98 ( .A(npu_inst_pe_1_5_5_n55), .ZN(
        npu_inst_pe_1_5_5_n103) );
  AOI22_X1 npu_inst_pe_1_5_5_U97 ( .A1(npu_inst_int_data_y_6__5__1_), .A2(
        npu_inst_pe_1_5_5_n50), .B1(npu_inst_pe_1_5_5_n117), .B2(
        npu_inst_pe_1_5_5_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_5_5_n51) );
  INV_X1 npu_inst_pe_1_5_5_U96 ( .A(npu_inst_pe_1_5_5_n51), .ZN(
        npu_inst_pe_1_5_5_n104) );
  AOI22_X1 npu_inst_pe_1_5_5_U95 ( .A1(npu_inst_int_data_y_6__5__1_), .A2(
        npu_inst_pe_1_5_5_n46), .B1(npu_inst_pe_1_5_5_n116), .B2(
        npu_inst_pe_1_5_5_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_5_5_n47) );
  INV_X1 npu_inst_pe_1_5_5_U94 ( .A(npu_inst_pe_1_5_5_n47), .ZN(
        npu_inst_pe_1_5_5_n105) );
  AOI22_X1 npu_inst_pe_1_5_5_U93 ( .A1(npu_inst_int_data_y_6__5__1_), .A2(
        npu_inst_pe_1_5_5_n42), .B1(npu_inst_pe_1_5_5_n115), .B2(
        npu_inst_pe_1_5_5_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_5_5_n43) );
  INV_X1 npu_inst_pe_1_5_5_U92 ( .A(npu_inst_pe_1_5_5_n43), .ZN(
        npu_inst_pe_1_5_5_n106) );
  AOI22_X1 npu_inst_pe_1_5_5_U91 ( .A1(npu_inst_pe_1_5_5_n38), .A2(
        npu_inst_int_data_y_6__5__1_), .B1(npu_inst_pe_1_5_5_n114), .B2(
        npu_inst_pe_1_5_5_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_5_5_n39) );
  INV_X1 npu_inst_pe_1_5_5_U90 ( .A(npu_inst_pe_1_5_5_n39), .ZN(
        npu_inst_pe_1_5_5_n107) );
  AOI22_X1 npu_inst_pe_1_5_5_U89 ( .A1(npu_inst_pe_1_5_5_n38), .A2(
        npu_inst_int_data_y_6__5__0_), .B1(npu_inst_pe_1_5_5_n114), .B2(
        npu_inst_pe_1_5_5_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_5_5_n37) );
  INV_X1 npu_inst_pe_1_5_5_U88 ( .A(npu_inst_pe_1_5_5_n37), .ZN(
        npu_inst_pe_1_5_5_n113) );
  NAND2_X1 npu_inst_pe_1_5_5_U87 ( .A1(npu_inst_pe_1_5_5_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_5_5_n60), .ZN(npu_inst_pe_1_5_5_n74) );
  OAI21_X1 npu_inst_pe_1_5_5_U86 ( .B1(npu_inst_pe_1_5_5_n63), .B2(
        npu_inst_pe_1_5_5_n60), .A(npu_inst_pe_1_5_5_n74), .ZN(
        npu_inst_pe_1_5_5_n97) );
  NAND2_X1 npu_inst_pe_1_5_5_U85 ( .A1(npu_inst_pe_1_5_5_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_5_5_n60), .ZN(npu_inst_pe_1_5_5_n73) );
  OAI21_X1 npu_inst_pe_1_5_5_U84 ( .B1(npu_inst_pe_1_5_5_n61), .B2(
        npu_inst_pe_1_5_5_n60), .A(npu_inst_pe_1_5_5_n73), .ZN(
        npu_inst_pe_1_5_5_n96) );
  NAND2_X1 npu_inst_pe_1_5_5_U83 ( .A1(npu_inst_pe_1_5_5_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_5_5_n56), .ZN(npu_inst_pe_1_5_5_n72) );
  OAI21_X1 npu_inst_pe_1_5_5_U82 ( .B1(npu_inst_pe_1_5_5_n63), .B2(
        npu_inst_pe_1_5_5_n56), .A(npu_inst_pe_1_5_5_n72), .ZN(
        npu_inst_pe_1_5_5_n95) );
  NAND2_X1 npu_inst_pe_1_5_5_U81 ( .A1(npu_inst_pe_1_5_5_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_5_5_n56), .ZN(npu_inst_pe_1_5_5_n71) );
  OAI21_X1 npu_inst_pe_1_5_5_U80 ( .B1(npu_inst_pe_1_5_5_n61), .B2(
        npu_inst_pe_1_5_5_n56), .A(npu_inst_pe_1_5_5_n71), .ZN(
        npu_inst_pe_1_5_5_n94) );
  NAND2_X1 npu_inst_pe_1_5_5_U79 ( .A1(npu_inst_pe_1_5_5_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_5_5_n52), .ZN(npu_inst_pe_1_5_5_n70) );
  OAI21_X1 npu_inst_pe_1_5_5_U78 ( .B1(npu_inst_pe_1_5_5_n63), .B2(
        npu_inst_pe_1_5_5_n52), .A(npu_inst_pe_1_5_5_n70), .ZN(
        npu_inst_pe_1_5_5_n93) );
  NAND2_X1 npu_inst_pe_1_5_5_U77 ( .A1(npu_inst_pe_1_5_5_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_5_5_n52), .ZN(npu_inst_pe_1_5_5_n69) );
  OAI21_X1 npu_inst_pe_1_5_5_U76 ( .B1(npu_inst_pe_1_5_5_n61), .B2(
        npu_inst_pe_1_5_5_n52), .A(npu_inst_pe_1_5_5_n69), .ZN(
        npu_inst_pe_1_5_5_n92) );
  NAND2_X1 npu_inst_pe_1_5_5_U75 ( .A1(npu_inst_pe_1_5_5_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_5_5_n48), .ZN(npu_inst_pe_1_5_5_n68) );
  OAI21_X1 npu_inst_pe_1_5_5_U74 ( .B1(npu_inst_pe_1_5_5_n63), .B2(
        npu_inst_pe_1_5_5_n48), .A(npu_inst_pe_1_5_5_n68), .ZN(
        npu_inst_pe_1_5_5_n91) );
  NAND2_X1 npu_inst_pe_1_5_5_U73 ( .A1(npu_inst_pe_1_5_5_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_5_5_n48), .ZN(npu_inst_pe_1_5_5_n67) );
  OAI21_X1 npu_inst_pe_1_5_5_U72 ( .B1(npu_inst_pe_1_5_5_n61), .B2(
        npu_inst_pe_1_5_5_n48), .A(npu_inst_pe_1_5_5_n67), .ZN(
        npu_inst_pe_1_5_5_n90) );
  NAND2_X1 npu_inst_pe_1_5_5_U71 ( .A1(npu_inst_pe_1_5_5_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_5_5_n44), .ZN(npu_inst_pe_1_5_5_n66) );
  OAI21_X1 npu_inst_pe_1_5_5_U70 ( .B1(npu_inst_pe_1_5_5_n63), .B2(
        npu_inst_pe_1_5_5_n44), .A(npu_inst_pe_1_5_5_n66), .ZN(
        npu_inst_pe_1_5_5_n89) );
  NAND2_X1 npu_inst_pe_1_5_5_U69 ( .A1(npu_inst_pe_1_5_5_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_5_5_n44), .ZN(npu_inst_pe_1_5_5_n65) );
  OAI21_X1 npu_inst_pe_1_5_5_U68 ( .B1(npu_inst_pe_1_5_5_n61), .B2(
        npu_inst_pe_1_5_5_n44), .A(npu_inst_pe_1_5_5_n65), .ZN(
        npu_inst_pe_1_5_5_n88) );
  NAND2_X1 npu_inst_pe_1_5_5_U67 ( .A1(npu_inst_pe_1_5_5_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_5_5_n40), .ZN(npu_inst_pe_1_5_5_n64) );
  OAI21_X1 npu_inst_pe_1_5_5_U66 ( .B1(npu_inst_pe_1_5_5_n63), .B2(
        npu_inst_pe_1_5_5_n40), .A(npu_inst_pe_1_5_5_n64), .ZN(
        npu_inst_pe_1_5_5_n87) );
  NAND2_X1 npu_inst_pe_1_5_5_U65 ( .A1(npu_inst_pe_1_5_5_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_5_5_n40), .ZN(npu_inst_pe_1_5_5_n62) );
  OAI21_X1 npu_inst_pe_1_5_5_U64 ( .B1(npu_inst_pe_1_5_5_n61), .B2(
        npu_inst_pe_1_5_5_n40), .A(npu_inst_pe_1_5_5_n62), .ZN(
        npu_inst_pe_1_5_5_n86) );
  AND2_X1 npu_inst_pe_1_5_5_U63 ( .A1(npu_inst_pe_1_5_5_N93), .A2(npu_inst_n54), .ZN(npu_inst_int_data_y_5__5__0_) );
  AND2_X1 npu_inst_pe_1_5_5_U62 ( .A1(npu_inst_n54), .A2(npu_inst_pe_1_5_5_N94), .ZN(npu_inst_int_data_y_5__5__1_) );
  NOR3_X1 npu_inst_pe_1_5_5_U61 ( .A1(npu_inst_pe_1_5_5_n26), .A2(npu_inst_n54), .A3(npu_inst_int_ckg[18]), .ZN(npu_inst_pe_1_5_5_n85) );
  OR2_X1 npu_inst_pe_1_5_5_U60 ( .A1(npu_inst_pe_1_5_5_n85), .A2(
        npu_inst_pe_1_5_5_n2), .ZN(npu_inst_pe_1_5_5_N84) );
  AND2_X1 npu_inst_pe_1_5_5_U59 ( .A1(npu_inst_pe_1_5_5_int_q_acc_0_), .A2(
        npu_inst_pe_1_5_5_n1), .ZN(npu_inst_int_data_res_5__5__0_) );
  AND2_X1 npu_inst_pe_1_5_5_U58 ( .A1(npu_inst_pe_1_5_5_n2), .A2(
        npu_inst_pe_1_5_5_int_q_acc_7_), .ZN(npu_inst_int_data_res_5__5__7_)
         );
  AND2_X1 npu_inst_pe_1_5_5_U57 ( .A1(npu_inst_pe_1_5_5_int_q_acc_1_), .A2(
        npu_inst_pe_1_5_5_n1), .ZN(npu_inst_int_data_res_5__5__1_) );
  AND2_X1 npu_inst_pe_1_5_5_U56 ( .A1(npu_inst_pe_1_5_5_int_q_acc_2_), .A2(
        npu_inst_pe_1_5_5_n1), .ZN(npu_inst_int_data_res_5__5__2_) );
  AND2_X1 npu_inst_pe_1_5_5_U55 ( .A1(npu_inst_pe_1_5_5_int_q_acc_3_), .A2(
        npu_inst_pe_1_5_5_n2), .ZN(npu_inst_int_data_res_5__5__3_) );
  AND2_X1 npu_inst_pe_1_5_5_U54 ( .A1(npu_inst_pe_1_5_5_int_q_acc_4_), .A2(
        npu_inst_pe_1_5_5_n2), .ZN(npu_inst_int_data_res_5__5__4_) );
  AND2_X1 npu_inst_pe_1_5_5_U53 ( .A1(npu_inst_pe_1_5_5_int_q_acc_5_), .A2(
        npu_inst_pe_1_5_5_n2), .ZN(npu_inst_int_data_res_5__5__5_) );
  AND2_X1 npu_inst_pe_1_5_5_U52 ( .A1(npu_inst_pe_1_5_5_int_q_acc_6_), .A2(
        npu_inst_pe_1_5_5_n2), .ZN(npu_inst_int_data_res_5__5__6_) );
  AOI222_X1 npu_inst_pe_1_5_5_U51 ( .A1(npu_inst_int_data_res_6__5__0_), .A2(
        npu_inst_pe_1_5_5_n1), .B1(npu_inst_pe_1_5_5_N73), .B2(
        npu_inst_pe_1_5_5_n76), .C1(npu_inst_pe_1_5_5_N65), .C2(
        npu_inst_pe_1_5_5_n77), .ZN(npu_inst_pe_1_5_5_n84) );
  INV_X1 npu_inst_pe_1_5_5_U50 ( .A(npu_inst_pe_1_5_5_n84), .ZN(
        npu_inst_pe_1_5_5_n101) );
  AOI222_X1 npu_inst_pe_1_5_5_U49 ( .A1(npu_inst_int_data_res_6__5__7_), .A2(
        npu_inst_pe_1_5_5_n1), .B1(npu_inst_pe_1_5_5_N80), .B2(
        npu_inst_pe_1_5_5_n76), .C1(npu_inst_pe_1_5_5_N72), .C2(
        npu_inst_pe_1_5_5_n77), .ZN(npu_inst_pe_1_5_5_n75) );
  INV_X1 npu_inst_pe_1_5_5_U48 ( .A(npu_inst_pe_1_5_5_n75), .ZN(
        npu_inst_pe_1_5_5_n33) );
  AOI222_X1 npu_inst_pe_1_5_5_U47 ( .A1(npu_inst_int_data_res_6__5__1_), .A2(
        npu_inst_pe_1_5_5_n1), .B1(npu_inst_pe_1_5_5_N74), .B2(
        npu_inst_pe_1_5_5_n76), .C1(npu_inst_pe_1_5_5_N66), .C2(
        npu_inst_pe_1_5_5_n77), .ZN(npu_inst_pe_1_5_5_n83) );
  INV_X1 npu_inst_pe_1_5_5_U46 ( .A(npu_inst_pe_1_5_5_n83), .ZN(
        npu_inst_pe_1_5_5_n100) );
  AOI222_X1 npu_inst_pe_1_5_5_U45 ( .A1(npu_inst_int_data_res_6__5__2_), .A2(
        npu_inst_pe_1_5_5_n1), .B1(npu_inst_pe_1_5_5_N75), .B2(
        npu_inst_pe_1_5_5_n76), .C1(npu_inst_pe_1_5_5_N67), .C2(
        npu_inst_pe_1_5_5_n77), .ZN(npu_inst_pe_1_5_5_n82) );
  INV_X1 npu_inst_pe_1_5_5_U44 ( .A(npu_inst_pe_1_5_5_n82), .ZN(
        npu_inst_pe_1_5_5_n99) );
  AOI222_X1 npu_inst_pe_1_5_5_U43 ( .A1(npu_inst_int_data_res_6__5__3_), .A2(
        npu_inst_pe_1_5_5_n1), .B1(npu_inst_pe_1_5_5_N76), .B2(
        npu_inst_pe_1_5_5_n76), .C1(npu_inst_pe_1_5_5_N68), .C2(
        npu_inst_pe_1_5_5_n77), .ZN(npu_inst_pe_1_5_5_n81) );
  INV_X1 npu_inst_pe_1_5_5_U42 ( .A(npu_inst_pe_1_5_5_n81), .ZN(
        npu_inst_pe_1_5_5_n98) );
  AOI222_X1 npu_inst_pe_1_5_5_U41 ( .A1(npu_inst_int_data_res_6__5__4_), .A2(
        npu_inst_pe_1_5_5_n1), .B1(npu_inst_pe_1_5_5_N77), .B2(
        npu_inst_pe_1_5_5_n76), .C1(npu_inst_pe_1_5_5_N69), .C2(
        npu_inst_pe_1_5_5_n77), .ZN(npu_inst_pe_1_5_5_n80) );
  INV_X1 npu_inst_pe_1_5_5_U40 ( .A(npu_inst_pe_1_5_5_n80), .ZN(
        npu_inst_pe_1_5_5_n36) );
  AOI222_X1 npu_inst_pe_1_5_5_U39 ( .A1(npu_inst_int_data_res_6__5__5_), .A2(
        npu_inst_pe_1_5_5_n1), .B1(npu_inst_pe_1_5_5_N78), .B2(
        npu_inst_pe_1_5_5_n76), .C1(npu_inst_pe_1_5_5_N70), .C2(
        npu_inst_pe_1_5_5_n77), .ZN(npu_inst_pe_1_5_5_n79) );
  INV_X1 npu_inst_pe_1_5_5_U38 ( .A(npu_inst_pe_1_5_5_n79), .ZN(
        npu_inst_pe_1_5_5_n35) );
  AOI222_X1 npu_inst_pe_1_5_5_U37 ( .A1(npu_inst_int_data_res_6__5__6_), .A2(
        npu_inst_pe_1_5_5_n1), .B1(npu_inst_pe_1_5_5_N79), .B2(
        npu_inst_pe_1_5_5_n76), .C1(npu_inst_pe_1_5_5_N71), .C2(
        npu_inst_pe_1_5_5_n77), .ZN(npu_inst_pe_1_5_5_n78) );
  INV_X1 npu_inst_pe_1_5_5_U36 ( .A(npu_inst_pe_1_5_5_n78), .ZN(
        npu_inst_pe_1_5_5_n34) );
  INV_X1 npu_inst_pe_1_5_5_U35 ( .A(npu_inst_pe_1_5_5_int_data_1_), .ZN(
        npu_inst_pe_1_5_5_n14) );
  AND2_X1 npu_inst_pe_1_5_5_U34 ( .A1(npu_inst_int_data_x_5__5__1_), .A2(
        npu_inst_pe_1_5_5_int_q_weight_1_), .ZN(npu_inst_pe_1_5_5_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_5_5_U33 ( .A1(npu_inst_int_data_x_5__5__0_), .A2(
        npu_inst_pe_1_5_5_int_q_weight_1_), .ZN(npu_inst_pe_1_5_5_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_5_5_U32 ( .A1(npu_inst_n54), .A2(
        npu_inst_int_data_y_6__5__1_), .B1(npu_inst_pe_1_5_5_n3), .B2(
        npu_inst_int_data_x_5__6__1_), .ZN(npu_inst_pe_1_5_5_n63) );
  AOI22_X1 npu_inst_pe_1_5_5_U31 ( .A1(npu_inst_n54), .A2(
        npu_inst_int_data_y_6__5__0_), .B1(npu_inst_pe_1_5_5_n3), .B2(
        npu_inst_int_data_x_5__6__0_), .ZN(npu_inst_pe_1_5_5_n61) );
  INV_X1 npu_inst_pe_1_5_5_U30 ( .A(npu_inst_pe_1_5_5_int_data_0_), .ZN(
        npu_inst_pe_1_5_5_n13) );
  INV_X1 npu_inst_pe_1_5_5_U29 ( .A(npu_inst_n68), .ZN(npu_inst_pe_1_5_5_n5)
         );
  OR3_X1 npu_inst_pe_1_5_5_U28 ( .A1(npu_inst_pe_1_5_5_n6), .A2(
        npu_inst_pe_1_5_5_n8), .A3(npu_inst_pe_1_5_5_n5), .ZN(
        npu_inst_pe_1_5_5_n56) );
  OR3_X1 npu_inst_pe_1_5_5_U27 ( .A1(npu_inst_pe_1_5_5_n5), .A2(
        npu_inst_pe_1_5_5_n8), .A3(npu_inst_pe_1_5_5_n7), .ZN(
        npu_inst_pe_1_5_5_n48) );
  INV_X1 npu_inst_pe_1_5_5_U26 ( .A(npu_inst_pe_1_5_5_n5), .ZN(
        npu_inst_pe_1_5_5_n4) );
  OR3_X1 npu_inst_pe_1_5_5_U25 ( .A1(npu_inst_pe_1_5_5_n4), .A2(
        npu_inst_pe_1_5_5_n8), .A3(npu_inst_pe_1_5_5_n7), .ZN(
        npu_inst_pe_1_5_5_n52) );
  OR3_X1 npu_inst_pe_1_5_5_U24 ( .A1(npu_inst_pe_1_5_5_n6), .A2(
        npu_inst_pe_1_5_5_n8), .A3(npu_inst_pe_1_5_5_n4), .ZN(
        npu_inst_pe_1_5_5_n60) );
  NOR2_X1 npu_inst_pe_1_5_5_U23 ( .A1(npu_inst_pe_1_5_5_n60), .A2(
        npu_inst_pe_1_5_5_n3), .ZN(npu_inst_pe_1_5_5_n58) );
  NOR2_X1 npu_inst_pe_1_5_5_U22 ( .A1(npu_inst_pe_1_5_5_n56), .A2(
        npu_inst_pe_1_5_5_n3), .ZN(npu_inst_pe_1_5_5_n54) );
  NOR2_X1 npu_inst_pe_1_5_5_U21 ( .A1(npu_inst_pe_1_5_5_n52), .A2(
        npu_inst_pe_1_5_5_n3), .ZN(npu_inst_pe_1_5_5_n50) );
  NOR2_X1 npu_inst_pe_1_5_5_U20 ( .A1(npu_inst_pe_1_5_5_n48), .A2(
        npu_inst_pe_1_5_5_n3), .ZN(npu_inst_pe_1_5_5_n46) );
  NOR2_X1 npu_inst_pe_1_5_5_U19 ( .A1(npu_inst_pe_1_5_5_n40), .A2(
        npu_inst_pe_1_5_5_n3), .ZN(npu_inst_pe_1_5_5_n38) );
  NOR2_X1 npu_inst_pe_1_5_5_U18 ( .A1(npu_inst_pe_1_5_5_n44), .A2(
        npu_inst_pe_1_5_5_n3), .ZN(npu_inst_pe_1_5_5_n42) );
  BUF_X1 npu_inst_pe_1_5_5_U17 ( .A(npu_inst_n96), .Z(npu_inst_pe_1_5_5_n8) );
  INV_X1 npu_inst_pe_1_5_5_U16 ( .A(npu_inst_n123), .ZN(npu_inst_pe_1_5_5_n12)
         );
  INV_X1 npu_inst_pe_1_5_5_U15 ( .A(npu_inst_pe_1_5_5_n38), .ZN(
        npu_inst_pe_1_5_5_n114) );
  INV_X1 npu_inst_pe_1_5_5_U14 ( .A(npu_inst_pe_1_5_5_n58), .ZN(
        npu_inst_pe_1_5_5_n119) );
  INV_X1 npu_inst_pe_1_5_5_U13 ( .A(npu_inst_pe_1_5_5_n54), .ZN(
        npu_inst_pe_1_5_5_n118) );
  INV_X1 npu_inst_pe_1_5_5_U12 ( .A(npu_inst_pe_1_5_5_n50), .ZN(
        npu_inst_pe_1_5_5_n117) );
  INV_X1 npu_inst_pe_1_5_5_U11 ( .A(npu_inst_pe_1_5_5_n46), .ZN(
        npu_inst_pe_1_5_5_n116) );
  INV_X1 npu_inst_pe_1_5_5_U10 ( .A(npu_inst_pe_1_5_5_n42), .ZN(
        npu_inst_pe_1_5_5_n115) );
  BUF_X1 npu_inst_pe_1_5_5_U9 ( .A(npu_inst_n16), .Z(npu_inst_pe_1_5_5_n2) );
  BUF_X1 npu_inst_pe_1_5_5_U8 ( .A(npu_inst_n16), .Z(npu_inst_pe_1_5_5_n1) );
  BUF_X1 npu_inst_pe_1_5_5_U7 ( .A(npu_inst_pe_1_5_5_n12), .Z(
        npu_inst_pe_1_5_5_n11) );
  BUF_X1 npu_inst_pe_1_5_5_U6 ( .A(npu_inst_pe_1_5_5_n12), .Z(
        npu_inst_pe_1_5_5_n10) );
  BUF_X1 npu_inst_pe_1_5_5_U5 ( .A(npu_inst_pe_1_5_5_n12), .Z(
        npu_inst_pe_1_5_5_n9) );
  NOR2_X1 npu_inst_pe_1_5_5_U4 ( .A1(npu_inst_pe_1_5_5_int_q_weight_0_), .A2(
        npu_inst_pe_1_5_5_n1), .ZN(npu_inst_pe_1_5_5_n76) );
  NOR2_X1 npu_inst_pe_1_5_5_U3 ( .A1(npu_inst_pe_1_5_5_n27), .A2(
        npu_inst_pe_1_5_5_n1), .ZN(npu_inst_pe_1_5_5_n77) );
  FA_X1 npu_inst_pe_1_5_5_sub_67_U2_1 ( .A(npu_inst_pe_1_5_5_int_q_acc_1_), 
        .B(npu_inst_pe_1_5_5_n14), .CI(npu_inst_pe_1_5_5_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_5_5_sub_67_carry_2_), .S(npu_inst_pe_1_5_5_N66) );
  FA_X1 npu_inst_pe_1_5_5_add_69_U1_1 ( .A(npu_inst_pe_1_5_5_int_q_acc_1_), 
        .B(npu_inst_pe_1_5_5_int_data_1_), .CI(
        npu_inst_pe_1_5_5_add_69_carry_1_), .CO(
        npu_inst_pe_1_5_5_add_69_carry_2_), .S(npu_inst_pe_1_5_5_N74) );
  NAND3_X1 npu_inst_pe_1_5_5_U109 ( .A1(npu_inst_pe_1_5_5_n5), .A2(
        npu_inst_pe_1_5_5_n7), .A3(npu_inst_pe_1_5_5_n8), .ZN(
        npu_inst_pe_1_5_5_n44) );
  NAND3_X1 npu_inst_pe_1_5_5_U108 ( .A1(npu_inst_pe_1_5_5_n4), .A2(
        npu_inst_pe_1_5_5_n7), .A3(npu_inst_pe_1_5_5_n8), .ZN(
        npu_inst_pe_1_5_5_n40) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_5_5_n34), .CK(
        npu_inst_pe_1_5_5_net3527), .RN(npu_inst_pe_1_5_5_n9), .Q(
        npu_inst_pe_1_5_5_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_5_5_n35), .CK(
        npu_inst_pe_1_5_5_net3527), .RN(npu_inst_pe_1_5_5_n9), .Q(
        npu_inst_pe_1_5_5_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_5_5_n36), .CK(
        npu_inst_pe_1_5_5_net3527), .RN(npu_inst_pe_1_5_5_n9), .Q(
        npu_inst_pe_1_5_5_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_5_5_n98), .CK(
        npu_inst_pe_1_5_5_net3527), .RN(npu_inst_pe_1_5_5_n9), .Q(
        npu_inst_pe_1_5_5_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_5_5_n99), .CK(
        npu_inst_pe_1_5_5_net3527), .RN(npu_inst_pe_1_5_5_n9), .Q(
        npu_inst_pe_1_5_5_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_5_5_n100), 
        .CK(npu_inst_pe_1_5_5_net3527), .RN(npu_inst_pe_1_5_5_n9), .Q(
        npu_inst_pe_1_5_5_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_5_5_n33), .CK(
        npu_inst_pe_1_5_5_net3527), .RN(npu_inst_pe_1_5_5_n9), .Q(
        npu_inst_pe_1_5_5_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_5_5_n101), 
        .CK(npu_inst_pe_1_5_5_net3527), .RN(npu_inst_pe_1_5_5_n9), .Q(
        npu_inst_pe_1_5_5_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_weight_reg_0_ ( .D(npu_inst_n109), .CK(
        npu_inst_pe_1_5_5_net3533), .RN(npu_inst_pe_1_5_5_n9), .Q(
        npu_inst_pe_1_5_5_int_q_weight_0_), .QN(npu_inst_pe_1_5_5_n27) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_weight_reg_1_ ( .D(npu_inst_n115), .CK(
        npu_inst_pe_1_5_5_net3533), .RN(npu_inst_pe_1_5_5_n9), .Q(
        npu_inst_pe_1_5_5_int_q_weight_1_), .QN(npu_inst_pe_1_5_5_n26) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_5_5_n113), 
        .CK(npu_inst_pe_1_5_5_net3533), .RN(npu_inst_pe_1_5_5_n9), .Q(
        npu_inst_pe_1_5_5_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_5_5_n107), 
        .CK(npu_inst_pe_1_5_5_net3533), .RN(npu_inst_pe_1_5_5_n9), .Q(
        npu_inst_pe_1_5_5_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_5_5_n112), 
        .CK(npu_inst_pe_1_5_5_net3533), .RN(npu_inst_pe_1_5_5_n10), .Q(
        npu_inst_pe_1_5_5_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_5_5_n106), 
        .CK(npu_inst_pe_1_5_5_net3533), .RN(npu_inst_pe_1_5_5_n10), .Q(
        npu_inst_pe_1_5_5_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_5_5_n111), 
        .CK(npu_inst_pe_1_5_5_net3533), .RN(npu_inst_pe_1_5_5_n10), .Q(
        npu_inst_pe_1_5_5_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_5_5_n105), 
        .CK(npu_inst_pe_1_5_5_net3533), .RN(npu_inst_pe_1_5_5_n10), .Q(
        npu_inst_pe_1_5_5_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_5_5_n110), 
        .CK(npu_inst_pe_1_5_5_net3533), .RN(npu_inst_pe_1_5_5_n10), .Q(
        npu_inst_pe_1_5_5_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_5_5_n104), 
        .CK(npu_inst_pe_1_5_5_net3533), .RN(npu_inst_pe_1_5_5_n10), .Q(
        npu_inst_pe_1_5_5_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_5_5_n109), 
        .CK(npu_inst_pe_1_5_5_net3533), .RN(npu_inst_pe_1_5_5_n10), .Q(
        npu_inst_pe_1_5_5_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_5_5_n103), 
        .CK(npu_inst_pe_1_5_5_net3533), .RN(npu_inst_pe_1_5_5_n10), .Q(
        npu_inst_pe_1_5_5_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_5_5_n108), 
        .CK(npu_inst_pe_1_5_5_net3533), .RN(npu_inst_pe_1_5_5_n10), .Q(
        npu_inst_pe_1_5_5_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_5_5_n102), 
        .CK(npu_inst_pe_1_5_5_net3533), .RN(npu_inst_pe_1_5_5_n10), .Q(
        npu_inst_pe_1_5_5_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_5_5_n86), 
        .CK(npu_inst_pe_1_5_5_net3533), .RN(npu_inst_pe_1_5_5_n10), .Q(
        npu_inst_pe_1_5_5_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_5_5_n87), 
        .CK(npu_inst_pe_1_5_5_net3533), .RN(npu_inst_pe_1_5_5_n10), .Q(
        npu_inst_pe_1_5_5_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_5_5_n88), 
        .CK(npu_inst_pe_1_5_5_net3533), .RN(npu_inst_pe_1_5_5_n11), .Q(
        npu_inst_pe_1_5_5_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_5_5_n89), 
        .CK(npu_inst_pe_1_5_5_net3533), .RN(npu_inst_pe_1_5_5_n11), .Q(
        npu_inst_pe_1_5_5_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_5_5_n90), 
        .CK(npu_inst_pe_1_5_5_net3533), .RN(npu_inst_pe_1_5_5_n11), .Q(
        npu_inst_pe_1_5_5_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_5_5_n91), 
        .CK(npu_inst_pe_1_5_5_net3533), .RN(npu_inst_pe_1_5_5_n11), .Q(
        npu_inst_pe_1_5_5_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_5_5_n92), 
        .CK(npu_inst_pe_1_5_5_net3533), .RN(npu_inst_pe_1_5_5_n11), .Q(
        npu_inst_pe_1_5_5_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_5_5_n93), 
        .CK(npu_inst_pe_1_5_5_net3533), .RN(npu_inst_pe_1_5_5_n11), .Q(
        npu_inst_pe_1_5_5_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_5_5_n94), 
        .CK(npu_inst_pe_1_5_5_net3533), .RN(npu_inst_pe_1_5_5_n11), .Q(
        npu_inst_pe_1_5_5_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_5_5_n95), 
        .CK(npu_inst_pe_1_5_5_net3533), .RN(npu_inst_pe_1_5_5_n11), .Q(
        npu_inst_pe_1_5_5_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_5_5_n96), 
        .CK(npu_inst_pe_1_5_5_net3533), .RN(npu_inst_pe_1_5_5_n11), .Q(
        npu_inst_pe_1_5_5_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_5_5_n97), 
        .CK(npu_inst_pe_1_5_5_net3533), .RN(npu_inst_pe_1_5_5_n11), .Q(
        npu_inst_pe_1_5_5_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_5_5_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_5_5_N84), .SE(1'b0), .GCK(npu_inst_pe_1_5_5_net3527) );
  CLKGATETST_X1 npu_inst_pe_1_5_5_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n62), .SE(1'b0), .GCK(npu_inst_pe_1_5_5_net3533) );
  MUX2_X1 npu_inst_pe_1_5_6_U162 ( .A(npu_inst_pe_1_5_6_n32), .B(
        npu_inst_pe_1_5_6_n29), .S(npu_inst_pe_1_5_6_n8), .Z(
        npu_inst_pe_1_5_6_N93) );
  MUX2_X1 npu_inst_pe_1_5_6_U161 ( .A(npu_inst_pe_1_5_6_n31), .B(
        npu_inst_pe_1_5_6_n30), .S(npu_inst_pe_1_5_6_n6), .Z(
        npu_inst_pe_1_5_6_n32) );
  MUX2_X1 npu_inst_pe_1_5_6_U160 ( .A(npu_inst_pe_1_5_6_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_5_6_int_q_reg_v_1__0_), .S(npu_inst_pe_1_5_6_n4), .Z(
        npu_inst_pe_1_5_6_n31) );
  MUX2_X1 npu_inst_pe_1_5_6_U159 ( .A(npu_inst_pe_1_5_6_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_5_6_int_q_reg_v_3__0_), .S(npu_inst_pe_1_5_6_n4), .Z(
        npu_inst_pe_1_5_6_n30) );
  MUX2_X1 npu_inst_pe_1_5_6_U158 ( .A(npu_inst_pe_1_5_6_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_5_6_int_q_reg_v_5__0_), .S(npu_inst_pe_1_5_6_n4), .Z(
        npu_inst_pe_1_5_6_n29) );
  MUX2_X1 npu_inst_pe_1_5_6_U157 ( .A(npu_inst_pe_1_5_6_n28), .B(
        npu_inst_pe_1_5_6_n23), .S(npu_inst_pe_1_5_6_n8), .Z(
        npu_inst_pe_1_5_6_N94) );
  MUX2_X1 npu_inst_pe_1_5_6_U156 ( .A(npu_inst_pe_1_5_6_n25), .B(
        npu_inst_pe_1_5_6_n24), .S(npu_inst_pe_1_5_6_n6), .Z(
        npu_inst_pe_1_5_6_n28) );
  MUX2_X1 npu_inst_pe_1_5_6_U155 ( .A(npu_inst_pe_1_5_6_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_5_6_int_q_reg_v_1__1_), .S(npu_inst_pe_1_5_6_n4), .Z(
        npu_inst_pe_1_5_6_n25) );
  MUX2_X1 npu_inst_pe_1_5_6_U154 ( .A(npu_inst_pe_1_5_6_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_5_6_int_q_reg_v_3__1_), .S(npu_inst_pe_1_5_6_n4), .Z(
        npu_inst_pe_1_5_6_n24) );
  MUX2_X1 npu_inst_pe_1_5_6_U153 ( .A(npu_inst_pe_1_5_6_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_5_6_int_q_reg_v_5__1_), .S(npu_inst_pe_1_5_6_n4), .Z(
        npu_inst_pe_1_5_6_n23) );
  MUX2_X1 npu_inst_pe_1_5_6_U152 ( .A(npu_inst_pe_1_5_6_n22), .B(
        npu_inst_pe_1_5_6_n19), .S(npu_inst_pe_1_5_6_n8), .Z(
        npu_inst_int_data_x_5__6__1_) );
  MUX2_X1 npu_inst_pe_1_5_6_U151 ( .A(npu_inst_pe_1_5_6_n21), .B(
        npu_inst_pe_1_5_6_n20), .S(npu_inst_pe_1_5_6_n6), .Z(
        npu_inst_pe_1_5_6_n22) );
  MUX2_X1 npu_inst_pe_1_5_6_U150 ( .A(npu_inst_pe_1_5_6_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_5_6_int_q_reg_h_1__1_), .S(npu_inst_pe_1_5_6_n4), .Z(
        npu_inst_pe_1_5_6_n21) );
  MUX2_X1 npu_inst_pe_1_5_6_U149 ( .A(npu_inst_pe_1_5_6_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_5_6_int_q_reg_h_3__1_), .S(npu_inst_pe_1_5_6_n4), .Z(
        npu_inst_pe_1_5_6_n20) );
  MUX2_X1 npu_inst_pe_1_5_6_U148 ( .A(npu_inst_pe_1_5_6_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_5_6_int_q_reg_h_5__1_), .S(npu_inst_pe_1_5_6_n4), .Z(
        npu_inst_pe_1_5_6_n19) );
  MUX2_X1 npu_inst_pe_1_5_6_U147 ( .A(npu_inst_pe_1_5_6_n18), .B(
        npu_inst_pe_1_5_6_n15), .S(npu_inst_pe_1_5_6_n8), .Z(
        npu_inst_int_data_x_5__6__0_) );
  MUX2_X1 npu_inst_pe_1_5_6_U146 ( .A(npu_inst_pe_1_5_6_n17), .B(
        npu_inst_pe_1_5_6_n16), .S(npu_inst_pe_1_5_6_n6), .Z(
        npu_inst_pe_1_5_6_n18) );
  MUX2_X1 npu_inst_pe_1_5_6_U145 ( .A(npu_inst_pe_1_5_6_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_5_6_int_q_reg_h_1__0_), .S(npu_inst_pe_1_5_6_n4), .Z(
        npu_inst_pe_1_5_6_n17) );
  MUX2_X1 npu_inst_pe_1_5_6_U144 ( .A(npu_inst_pe_1_5_6_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_5_6_int_q_reg_h_3__0_), .S(npu_inst_pe_1_5_6_n4), .Z(
        npu_inst_pe_1_5_6_n16) );
  MUX2_X1 npu_inst_pe_1_5_6_U143 ( .A(npu_inst_pe_1_5_6_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_5_6_int_q_reg_h_5__0_), .S(npu_inst_pe_1_5_6_n4), .Z(
        npu_inst_pe_1_5_6_n15) );
  XOR2_X1 npu_inst_pe_1_5_6_U142 ( .A(npu_inst_pe_1_5_6_int_data_0_), .B(
        npu_inst_pe_1_5_6_int_q_acc_0_), .Z(npu_inst_pe_1_5_6_N73) );
  AND2_X1 npu_inst_pe_1_5_6_U141 ( .A1(npu_inst_pe_1_5_6_int_q_acc_0_), .A2(
        npu_inst_pe_1_5_6_int_data_0_), .ZN(npu_inst_pe_1_5_6_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_5_6_U140 ( .A(npu_inst_pe_1_5_6_int_q_acc_0_), .B(
        npu_inst_pe_1_5_6_n13), .ZN(npu_inst_pe_1_5_6_N65) );
  OR2_X1 npu_inst_pe_1_5_6_U139 ( .A1(npu_inst_pe_1_5_6_n13), .A2(
        npu_inst_pe_1_5_6_int_q_acc_0_), .ZN(npu_inst_pe_1_5_6_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_5_6_U138 ( .A(npu_inst_pe_1_5_6_int_q_acc_2_), .B(
        npu_inst_pe_1_5_6_add_69_carry_2_), .Z(npu_inst_pe_1_5_6_N75) );
  AND2_X1 npu_inst_pe_1_5_6_U137 ( .A1(npu_inst_pe_1_5_6_add_69_carry_2_), 
        .A2(npu_inst_pe_1_5_6_int_q_acc_2_), .ZN(
        npu_inst_pe_1_5_6_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_5_6_U136 ( .A(npu_inst_pe_1_5_6_int_q_acc_3_), .B(
        npu_inst_pe_1_5_6_add_69_carry_3_), .Z(npu_inst_pe_1_5_6_N76) );
  AND2_X1 npu_inst_pe_1_5_6_U135 ( .A1(npu_inst_pe_1_5_6_add_69_carry_3_), 
        .A2(npu_inst_pe_1_5_6_int_q_acc_3_), .ZN(
        npu_inst_pe_1_5_6_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_5_6_U134 ( .A(npu_inst_pe_1_5_6_int_q_acc_4_), .B(
        npu_inst_pe_1_5_6_add_69_carry_4_), .Z(npu_inst_pe_1_5_6_N77) );
  AND2_X1 npu_inst_pe_1_5_6_U133 ( .A1(npu_inst_pe_1_5_6_add_69_carry_4_), 
        .A2(npu_inst_pe_1_5_6_int_q_acc_4_), .ZN(
        npu_inst_pe_1_5_6_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_5_6_U132 ( .A(npu_inst_pe_1_5_6_int_q_acc_5_), .B(
        npu_inst_pe_1_5_6_add_69_carry_5_), .Z(npu_inst_pe_1_5_6_N78) );
  AND2_X1 npu_inst_pe_1_5_6_U131 ( .A1(npu_inst_pe_1_5_6_add_69_carry_5_), 
        .A2(npu_inst_pe_1_5_6_int_q_acc_5_), .ZN(
        npu_inst_pe_1_5_6_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_5_6_U130 ( .A(npu_inst_pe_1_5_6_int_q_acc_6_), .B(
        npu_inst_pe_1_5_6_add_69_carry_6_), .Z(npu_inst_pe_1_5_6_N79) );
  AND2_X1 npu_inst_pe_1_5_6_U129 ( .A1(npu_inst_pe_1_5_6_add_69_carry_6_), 
        .A2(npu_inst_pe_1_5_6_int_q_acc_6_), .ZN(
        npu_inst_pe_1_5_6_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_5_6_U128 ( .A(npu_inst_pe_1_5_6_int_q_acc_7_), .B(
        npu_inst_pe_1_5_6_add_69_carry_7_), .Z(npu_inst_pe_1_5_6_N80) );
  XNOR2_X1 npu_inst_pe_1_5_6_U127 ( .A(npu_inst_pe_1_5_6_sub_67_carry_2_), .B(
        npu_inst_pe_1_5_6_int_q_acc_2_), .ZN(npu_inst_pe_1_5_6_N67) );
  OR2_X1 npu_inst_pe_1_5_6_U126 ( .A1(npu_inst_pe_1_5_6_int_q_acc_2_), .A2(
        npu_inst_pe_1_5_6_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_5_6_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_5_6_U125 ( .A(npu_inst_pe_1_5_6_sub_67_carry_3_), .B(
        npu_inst_pe_1_5_6_int_q_acc_3_), .ZN(npu_inst_pe_1_5_6_N68) );
  OR2_X1 npu_inst_pe_1_5_6_U124 ( .A1(npu_inst_pe_1_5_6_int_q_acc_3_), .A2(
        npu_inst_pe_1_5_6_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_5_6_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_5_6_U123 ( .A(npu_inst_pe_1_5_6_sub_67_carry_4_), .B(
        npu_inst_pe_1_5_6_int_q_acc_4_), .ZN(npu_inst_pe_1_5_6_N69) );
  OR2_X1 npu_inst_pe_1_5_6_U122 ( .A1(npu_inst_pe_1_5_6_int_q_acc_4_), .A2(
        npu_inst_pe_1_5_6_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_5_6_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_5_6_U121 ( .A(npu_inst_pe_1_5_6_sub_67_carry_5_), .B(
        npu_inst_pe_1_5_6_int_q_acc_5_), .ZN(npu_inst_pe_1_5_6_N70) );
  OR2_X1 npu_inst_pe_1_5_6_U120 ( .A1(npu_inst_pe_1_5_6_int_q_acc_5_), .A2(
        npu_inst_pe_1_5_6_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_5_6_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_5_6_U119 ( .A(npu_inst_pe_1_5_6_sub_67_carry_6_), .B(
        npu_inst_pe_1_5_6_int_q_acc_6_), .ZN(npu_inst_pe_1_5_6_N71) );
  OR2_X1 npu_inst_pe_1_5_6_U118 ( .A1(npu_inst_pe_1_5_6_int_q_acc_6_), .A2(
        npu_inst_pe_1_5_6_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_5_6_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_5_6_U117 ( .A(npu_inst_pe_1_5_6_int_q_acc_7_), .B(
        npu_inst_pe_1_5_6_sub_67_carry_7_), .ZN(npu_inst_pe_1_5_6_N72) );
  INV_X1 npu_inst_pe_1_5_6_U116 ( .A(npu_inst_n76), .ZN(npu_inst_pe_1_5_6_n7)
         );
  INV_X1 npu_inst_pe_1_5_6_U115 ( .A(npu_inst_pe_1_5_6_n7), .ZN(
        npu_inst_pe_1_5_6_n6) );
  INV_X1 npu_inst_pe_1_5_6_U114 ( .A(npu_inst_n54), .ZN(npu_inst_pe_1_5_6_n3)
         );
  AOI22_X1 npu_inst_pe_1_5_6_U113 ( .A1(npu_inst_int_data_y_6__6__0_), .A2(
        npu_inst_pe_1_5_6_n58), .B1(npu_inst_pe_1_5_6_n119), .B2(
        npu_inst_pe_1_5_6_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_5_6_n57) );
  INV_X1 npu_inst_pe_1_5_6_U112 ( .A(npu_inst_pe_1_5_6_n57), .ZN(
        npu_inst_pe_1_5_6_n108) );
  AOI22_X1 npu_inst_pe_1_5_6_U111 ( .A1(npu_inst_int_data_y_6__6__0_), .A2(
        npu_inst_pe_1_5_6_n54), .B1(npu_inst_pe_1_5_6_n118), .B2(
        npu_inst_pe_1_5_6_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_5_6_n53) );
  INV_X1 npu_inst_pe_1_5_6_U110 ( .A(npu_inst_pe_1_5_6_n53), .ZN(
        npu_inst_pe_1_5_6_n109) );
  AOI22_X1 npu_inst_pe_1_5_6_U107 ( .A1(npu_inst_int_data_y_6__6__0_), .A2(
        npu_inst_pe_1_5_6_n50), .B1(npu_inst_pe_1_5_6_n117), .B2(
        npu_inst_pe_1_5_6_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_5_6_n49) );
  INV_X1 npu_inst_pe_1_5_6_U106 ( .A(npu_inst_pe_1_5_6_n49), .ZN(
        npu_inst_pe_1_5_6_n110) );
  AOI22_X1 npu_inst_pe_1_5_6_U105 ( .A1(npu_inst_int_data_y_6__6__0_), .A2(
        npu_inst_pe_1_5_6_n46), .B1(npu_inst_pe_1_5_6_n116), .B2(
        npu_inst_pe_1_5_6_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_5_6_n45) );
  INV_X1 npu_inst_pe_1_5_6_U104 ( .A(npu_inst_pe_1_5_6_n45), .ZN(
        npu_inst_pe_1_5_6_n111) );
  AOI22_X1 npu_inst_pe_1_5_6_U103 ( .A1(npu_inst_int_data_y_6__6__0_), .A2(
        npu_inst_pe_1_5_6_n42), .B1(npu_inst_pe_1_5_6_n115), .B2(
        npu_inst_pe_1_5_6_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_5_6_n41) );
  INV_X1 npu_inst_pe_1_5_6_U102 ( .A(npu_inst_pe_1_5_6_n41), .ZN(
        npu_inst_pe_1_5_6_n112) );
  AOI22_X1 npu_inst_pe_1_5_6_U101 ( .A1(npu_inst_int_data_y_6__6__1_), .A2(
        npu_inst_pe_1_5_6_n58), .B1(npu_inst_pe_1_5_6_n119), .B2(
        npu_inst_pe_1_5_6_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_5_6_n59) );
  INV_X1 npu_inst_pe_1_5_6_U100 ( .A(npu_inst_pe_1_5_6_n59), .ZN(
        npu_inst_pe_1_5_6_n102) );
  AOI22_X1 npu_inst_pe_1_5_6_U99 ( .A1(npu_inst_int_data_y_6__6__1_), .A2(
        npu_inst_pe_1_5_6_n54), .B1(npu_inst_pe_1_5_6_n118), .B2(
        npu_inst_pe_1_5_6_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_5_6_n55) );
  INV_X1 npu_inst_pe_1_5_6_U98 ( .A(npu_inst_pe_1_5_6_n55), .ZN(
        npu_inst_pe_1_5_6_n103) );
  AOI22_X1 npu_inst_pe_1_5_6_U97 ( .A1(npu_inst_int_data_y_6__6__1_), .A2(
        npu_inst_pe_1_5_6_n50), .B1(npu_inst_pe_1_5_6_n117), .B2(
        npu_inst_pe_1_5_6_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_5_6_n51) );
  INV_X1 npu_inst_pe_1_5_6_U96 ( .A(npu_inst_pe_1_5_6_n51), .ZN(
        npu_inst_pe_1_5_6_n104) );
  AOI22_X1 npu_inst_pe_1_5_6_U95 ( .A1(npu_inst_int_data_y_6__6__1_), .A2(
        npu_inst_pe_1_5_6_n46), .B1(npu_inst_pe_1_5_6_n116), .B2(
        npu_inst_pe_1_5_6_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_5_6_n47) );
  INV_X1 npu_inst_pe_1_5_6_U94 ( .A(npu_inst_pe_1_5_6_n47), .ZN(
        npu_inst_pe_1_5_6_n105) );
  AOI22_X1 npu_inst_pe_1_5_6_U93 ( .A1(npu_inst_int_data_y_6__6__1_), .A2(
        npu_inst_pe_1_5_6_n42), .B1(npu_inst_pe_1_5_6_n115), .B2(
        npu_inst_pe_1_5_6_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_5_6_n43) );
  INV_X1 npu_inst_pe_1_5_6_U92 ( .A(npu_inst_pe_1_5_6_n43), .ZN(
        npu_inst_pe_1_5_6_n106) );
  AOI22_X1 npu_inst_pe_1_5_6_U91 ( .A1(npu_inst_pe_1_5_6_n38), .A2(
        npu_inst_int_data_y_6__6__1_), .B1(npu_inst_pe_1_5_6_n114), .B2(
        npu_inst_pe_1_5_6_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_5_6_n39) );
  INV_X1 npu_inst_pe_1_5_6_U90 ( .A(npu_inst_pe_1_5_6_n39), .ZN(
        npu_inst_pe_1_5_6_n107) );
  AOI22_X1 npu_inst_pe_1_5_6_U89 ( .A1(npu_inst_pe_1_5_6_n38), .A2(
        npu_inst_int_data_y_6__6__0_), .B1(npu_inst_pe_1_5_6_n114), .B2(
        npu_inst_pe_1_5_6_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_5_6_n37) );
  INV_X1 npu_inst_pe_1_5_6_U88 ( .A(npu_inst_pe_1_5_6_n37), .ZN(
        npu_inst_pe_1_5_6_n113) );
  NAND2_X1 npu_inst_pe_1_5_6_U87 ( .A1(npu_inst_pe_1_5_6_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_5_6_n60), .ZN(npu_inst_pe_1_5_6_n74) );
  OAI21_X1 npu_inst_pe_1_5_6_U86 ( .B1(npu_inst_pe_1_5_6_n63), .B2(
        npu_inst_pe_1_5_6_n60), .A(npu_inst_pe_1_5_6_n74), .ZN(
        npu_inst_pe_1_5_6_n97) );
  NAND2_X1 npu_inst_pe_1_5_6_U85 ( .A1(npu_inst_pe_1_5_6_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_5_6_n60), .ZN(npu_inst_pe_1_5_6_n73) );
  OAI21_X1 npu_inst_pe_1_5_6_U84 ( .B1(npu_inst_pe_1_5_6_n61), .B2(
        npu_inst_pe_1_5_6_n60), .A(npu_inst_pe_1_5_6_n73), .ZN(
        npu_inst_pe_1_5_6_n96) );
  NAND2_X1 npu_inst_pe_1_5_6_U83 ( .A1(npu_inst_pe_1_5_6_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_5_6_n56), .ZN(npu_inst_pe_1_5_6_n72) );
  OAI21_X1 npu_inst_pe_1_5_6_U82 ( .B1(npu_inst_pe_1_5_6_n63), .B2(
        npu_inst_pe_1_5_6_n56), .A(npu_inst_pe_1_5_6_n72), .ZN(
        npu_inst_pe_1_5_6_n95) );
  NAND2_X1 npu_inst_pe_1_5_6_U81 ( .A1(npu_inst_pe_1_5_6_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_5_6_n56), .ZN(npu_inst_pe_1_5_6_n71) );
  OAI21_X1 npu_inst_pe_1_5_6_U80 ( .B1(npu_inst_pe_1_5_6_n61), .B2(
        npu_inst_pe_1_5_6_n56), .A(npu_inst_pe_1_5_6_n71), .ZN(
        npu_inst_pe_1_5_6_n94) );
  NAND2_X1 npu_inst_pe_1_5_6_U79 ( .A1(npu_inst_pe_1_5_6_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_5_6_n52), .ZN(npu_inst_pe_1_5_6_n70) );
  OAI21_X1 npu_inst_pe_1_5_6_U78 ( .B1(npu_inst_pe_1_5_6_n63), .B2(
        npu_inst_pe_1_5_6_n52), .A(npu_inst_pe_1_5_6_n70), .ZN(
        npu_inst_pe_1_5_6_n93) );
  NAND2_X1 npu_inst_pe_1_5_6_U77 ( .A1(npu_inst_pe_1_5_6_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_5_6_n52), .ZN(npu_inst_pe_1_5_6_n69) );
  OAI21_X1 npu_inst_pe_1_5_6_U76 ( .B1(npu_inst_pe_1_5_6_n61), .B2(
        npu_inst_pe_1_5_6_n52), .A(npu_inst_pe_1_5_6_n69), .ZN(
        npu_inst_pe_1_5_6_n92) );
  NAND2_X1 npu_inst_pe_1_5_6_U75 ( .A1(npu_inst_pe_1_5_6_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_5_6_n48), .ZN(npu_inst_pe_1_5_6_n68) );
  OAI21_X1 npu_inst_pe_1_5_6_U74 ( .B1(npu_inst_pe_1_5_6_n63), .B2(
        npu_inst_pe_1_5_6_n48), .A(npu_inst_pe_1_5_6_n68), .ZN(
        npu_inst_pe_1_5_6_n91) );
  NAND2_X1 npu_inst_pe_1_5_6_U73 ( .A1(npu_inst_pe_1_5_6_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_5_6_n48), .ZN(npu_inst_pe_1_5_6_n67) );
  OAI21_X1 npu_inst_pe_1_5_6_U72 ( .B1(npu_inst_pe_1_5_6_n61), .B2(
        npu_inst_pe_1_5_6_n48), .A(npu_inst_pe_1_5_6_n67), .ZN(
        npu_inst_pe_1_5_6_n90) );
  NAND2_X1 npu_inst_pe_1_5_6_U71 ( .A1(npu_inst_pe_1_5_6_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_5_6_n44), .ZN(npu_inst_pe_1_5_6_n66) );
  OAI21_X1 npu_inst_pe_1_5_6_U70 ( .B1(npu_inst_pe_1_5_6_n63), .B2(
        npu_inst_pe_1_5_6_n44), .A(npu_inst_pe_1_5_6_n66), .ZN(
        npu_inst_pe_1_5_6_n89) );
  NAND2_X1 npu_inst_pe_1_5_6_U69 ( .A1(npu_inst_pe_1_5_6_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_5_6_n44), .ZN(npu_inst_pe_1_5_6_n65) );
  OAI21_X1 npu_inst_pe_1_5_6_U68 ( .B1(npu_inst_pe_1_5_6_n61), .B2(
        npu_inst_pe_1_5_6_n44), .A(npu_inst_pe_1_5_6_n65), .ZN(
        npu_inst_pe_1_5_6_n88) );
  NAND2_X1 npu_inst_pe_1_5_6_U67 ( .A1(npu_inst_pe_1_5_6_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_5_6_n40), .ZN(npu_inst_pe_1_5_6_n64) );
  OAI21_X1 npu_inst_pe_1_5_6_U66 ( .B1(npu_inst_pe_1_5_6_n63), .B2(
        npu_inst_pe_1_5_6_n40), .A(npu_inst_pe_1_5_6_n64), .ZN(
        npu_inst_pe_1_5_6_n87) );
  NAND2_X1 npu_inst_pe_1_5_6_U65 ( .A1(npu_inst_pe_1_5_6_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_5_6_n40), .ZN(npu_inst_pe_1_5_6_n62) );
  OAI21_X1 npu_inst_pe_1_5_6_U64 ( .B1(npu_inst_pe_1_5_6_n61), .B2(
        npu_inst_pe_1_5_6_n40), .A(npu_inst_pe_1_5_6_n62), .ZN(
        npu_inst_pe_1_5_6_n86) );
  AND2_X1 npu_inst_pe_1_5_6_U63 ( .A1(npu_inst_pe_1_5_6_N93), .A2(npu_inst_n54), .ZN(npu_inst_int_data_y_5__6__0_) );
  AND2_X1 npu_inst_pe_1_5_6_U62 ( .A1(npu_inst_n54), .A2(npu_inst_pe_1_5_6_N94), .ZN(npu_inst_int_data_y_5__6__1_) );
  NOR3_X1 npu_inst_pe_1_5_6_U61 ( .A1(npu_inst_pe_1_5_6_n26), .A2(npu_inst_n54), .A3(npu_inst_int_ckg[17]), .ZN(npu_inst_pe_1_5_6_n85) );
  OR2_X1 npu_inst_pe_1_5_6_U60 ( .A1(npu_inst_pe_1_5_6_n85), .A2(
        npu_inst_pe_1_5_6_n2), .ZN(npu_inst_pe_1_5_6_N84) );
  AND2_X1 npu_inst_pe_1_5_6_U59 ( .A1(npu_inst_pe_1_5_6_int_q_acc_0_), .A2(
        npu_inst_pe_1_5_6_n1), .ZN(npu_inst_int_data_res_5__6__0_) );
  AND2_X1 npu_inst_pe_1_5_6_U58 ( .A1(npu_inst_pe_1_5_6_n2), .A2(
        npu_inst_pe_1_5_6_int_q_acc_7_), .ZN(npu_inst_int_data_res_5__6__7_)
         );
  AND2_X1 npu_inst_pe_1_5_6_U57 ( .A1(npu_inst_pe_1_5_6_int_q_acc_1_), .A2(
        npu_inst_pe_1_5_6_n1), .ZN(npu_inst_int_data_res_5__6__1_) );
  AND2_X1 npu_inst_pe_1_5_6_U56 ( .A1(npu_inst_pe_1_5_6_int_q_acc_2_), .A2(
        npu_inst_pe_1_5_6_n1), .ZN(npu_inst_int_data_res_5__6__2_) );
  AND2_X1 npu_inst_pe_1_5_6_U55 ( .A1(npu_inst_pe_1_5_6_int_q_acc_3_), .A2(
        npu_inst_pe_1_5_6_n2), .ZN(npu_inst_int_data_res_5__6__3_) );
  AND2_X1 npu_inst_pe_1_5_6_U54 ( .A1(npu_inst_pe_1_5_6_int_q_acc_4_), .A2(
        npu_inst_pe_1_5_6_n2), .ZN(npu_inst_int_data_res_5__6__4_) );
  AND2_X1 npu_inst_pe_1_5_6_U53 ( .A1(npu_inst_pe_1_5_6_int_q_acc_5_), .A2(
        npu_inst_pe_1_5_6_n2), .ZN(npu_inst_int_data_res_5__6__5_) );
  AND2_X1 npu_inst_pe_1_5_6_U52 ( .A1(npu_inst_pe_1_5_6_int_q_acc_6_), .A2(
        npu_inst_pe_1_5_6_n2), .ZN(npu_inst_int_data_res_5__6__6_) );
  AOI222_X1 npu_inst_pe_1_5_6_U51 ( .A1(npu_inst_int_data_res_6__6__0_), .A2(
        npu_inst_pe_1_5_6_n1), .B1(npu_inst_pe_1_5_6_N73), .B2(
        npu_inst_pe_1_5_6_n76), .C1(npu_inst_pe_1_5_6_N65), .C2(
        npu_inst_pe_1_5_6_n77), .ZN(npu_inst_pe_1_5_6_n84) );
  INV_X1 npu_inst_pe_1_5_6_U50 ( .A(npu_inst_pe_1_5_6_n84), .ZN(
        npu_inst_pe_1_5_6_n101) );
  AOI222_X1 npu_inst_pe_1_5_6_U49 ( .A1(npu_inst_int_data_res_6__6__7_), .A2(
        npu_inst_pe_1_5_6_n1), .B1(npu_inst_pe_1_5_6_N80), .B2(
        npu_inst_pe_1_5_6_n76), .C1(npu_inst_pe_1_5_6_N72), .C2(
        npu_inst_pe_1_5_6_n77), .ZN(npu_inst_pe_1_5_6_n75) );
  INV_X1 npu_inst_pe_1_5_6_U48 ( .A(npu_inst_pe_1_5_6_n75), .ZN(
        npu_inst_pe_1_5_6_n33) );
  AOI222_X1 npu_inst_pe_1_5_6_U47 ( .A1(npu_inst_int_data_res_6__6__1_), .A2(
        npu_inst_pe_1_5_6_n1), .B1(npu_inst_pe_1_5_6_N74), .B2(
        npu_inst_pe_1_5_6_n76), .C1(npu_inst_pe_1_5_6_N66), .C2(
        npu_inst_pe_1_5_6_n77), .ZN(npu_inst_pe_1_5_6_n83) );
  INV_X1 npu_inst_pe_1_5_6_U46 ( .A(npu_inst_pe_1_5_6_n83), .ZN(
        npu_inst_pe_1_5_6_n100) );
  AOI222_X1 npu_inst_pe_1_5_6_U45 ( .A1(npu_inst_int_data_res_6__6__2_), .A2(
        npu_inst_pe_1_5_6_n1), .B1(npu_inst_pe_1_5_6_N75), .B2(
        npu_inst_pe_1_5_6_n76), .C1(npu_inst_pe_1_5_6_N67), .C2(
        npu_inst_pe_1_5_6_n77), .ZN(npu_inst_pe_1_5_6_n82) );
  INV_X1 npu_inst_pe_1_5_6_U44 ( .A(npu_inst_pe_1_5_6_n82), .ZN(
        npu_inst_pe_1_5_6_n99) );
  AOI222_X1 npu_inst_pe_1_5_6_U43 ( .A1(npu_inst_int_data_res_6__6__3_), .A2(
        npu_inst_pe_1_5_6_n1), .B1(npu_inst_pe_1_5_6_N76), .B2(
        npu_inst_pe_1_5_6_n76), .C1(npu_inst_pe_1_5_6_N68), .C2(
        npu_inst_pe_1_5_6_n77), .ZN(npu_inst_pe_1_5_6_n81) );
  INV_X1 npu_inst_pe_1_5_6_U42 ( .A(npu_inst_pe_1_5_6_n81), .ZN(
        npu_inst_pe_1_5_6_n98) );
  AOI222_X1 npu_inst_pe_1_5_6_U41 ( .A1(npu_inst_int_data_res_6__6__4_), .A2(
        npu_inst_pe_1_5_6_n1), .B1(npu_inst_pe_1_5_6_N77), .B2(
        npu_inst_pe_1_5_6_n76), .C1(npu_inst_pe_1_5_6_N69), .C2(
        npu_inst_pe_1_5_6_n77), .ZN(npu_inst_pe_1_5_6_n80) );
  INV_X1 npu_inst_pe_1_5_6_U40 ( .A(npu_inst_pe_1_5_6_n80), .ZN(
        npu_inst_pe_1_5_6_n36) );
  AOI222_X1 npu_inst_pe_1_5_6_U39 ( .A1(npu_inst_int_data_res_6__6__5_), .A2(
        npu_inst_pe_1_5_6_n1), .B1(npu_inst_pe_1_5_6_N78), .B2(
        npu_inst_pe_1_5_6_n76), .C1(npu_inst_pe_1_5_6_N70), .C2(
        npu_inst_pe_1_5_6_n77), .ZN(npu_inst_pe_1_5_6_n79) );
  INV_X1 npu_inst_pe_1_5_6_U38 ( .A(npu_inst_pe_1_5_6_n79), .ZN(
        npu_inst_pe_1_5_6_n35) );
  AOI222_X1 npu_inst_pe_1_5_6_U37 ( .A1(npu_inst_int_data_res_6__6__6_), .A2(
        npu_inst_pe_1_5_6_n1), .B1(npu_inst_pe_1_5_6_N79), .B2(
        npu_inst_pe_1_5_6_n76), .C1(npu_inst_pe_1_5_6_N71), .C2(
        npu_inst_pe_1_5_6_n77), .ZN(npu_inst_pe_1_5_6_n78) );
  INV_X1 npu_inst_pe_1_5_6_U36 ( .A(npu_inst_pe_1_5_6_n78), .ZN(
        npu_inst_pe_1_5_6_n34) );
  INV_X1 npu_inst_pe_1_5_6_U35 ( .A(npu_inst_pe_1_5_6_int_data_1_), .ZN(
        npu_inst_pe_1_5_6_n14) );
  AND2_X1 npu_inst_pe_1_5_6_U34 ( .A1(npu_inst_int_data_x_5__6__1_), .A2(
        npu_inst_pe_1_5_6_int_q_weight_1_), .ZN(npu_inst_pe_1_5_6_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_5_6_U33 ( .A1(npu_inst_int_data_x_5__6__0_), .A2(
        npu_inst_pe_1_5_6_int_q_weight_1_), .ZN(npu_inst_pe_1_5_6_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_5_6_U32 ( .A1(npu_inst_n54), .A2(
        npu_inst_int_data_y_6__6__1_), .B1(npu_inst_pe_1_5_6_n3), .B2(
        npu_inst_int_data_x_5__7__1_), .ZN(npu_inst_pe_1_5_6_n63) );
  AOI22_X1 npu_inst_pe_1_5_6_U31 ( .A1(npu_inst_n54), .A2(
        npu_inst_int_data_y_6__6__0_), .B1(npu_inst_pe_1_5_6_n3), .B2(
        npu_inst_int_data_x_5__7__0_), .ZN(npu_inst_pe_1_5_6_n61) );
  INV_X1 npu_inst_pe_1_5_6_U30 ( .A(npu_inst_pe_1_5_6_int_data_0_), .ZN(
        npu_inst_pe_1_5_6_n13) );
  INV_X1 npu_inst_pe_1_5_6_U29 ( .A(npu_inst_n68), .ZN(npu_inst_pe_1_5_6_n5)
         );
  OR3_X1 npu_inst_pe_1_5_6_U28 ( .A1(npu_inst_pe_1_5_6_n6), .A2(
        npu_inst_pe_1_5_6_n8), .A3(npu_inst_pe_1_5_6_n5), .ZN(
        npu_inst_pe_1_5_6_n56) );
  OR3_X1 npu_inst_pe_1_5_6_U27 ( .A1(npu_inst_pe_1_5_6_n5), .A2(
        npu_inst_pe_1_5_6_n8), .A3(npu_inst_pe_1_5_6_n7), .ZN(
        npu_inst_pe_1_5_6_n48) );
  INV_X1 npu_inst_pe_1_5_6_U26 ( .A(npu_inst_pe_1_5_6_n5), .ZN(
        npu_inst_pe_1_5_6_n4) );
  OR3_X1 npu_inst_pe_1_5_6_U25 ( .A1(npu_inst_pe_1_5_6_n4), .A2(
        npu_inst_pe_1_5_6_n8), .A3(npu_inst_pe_1_5_6_n7), .ZN(
        npu_inst_pe_1_5_6_n52) );
  OR3_X1 npu_inst_pe_1_5_6_U24 ( .A1(npu_inst_pe_1_5_6_n6), .A2(
        npu_inst_pe_1_5_6_n8), .A3(npu_inst_pe_1_5_6_n4), .ZN(
        npu_inst_pe_1_5_6_n60) );
  NOR2_X1 npu_inst_pe_1_5_6_U23 ( .A1(npu_inst_pe_1_5_6_n60), .A2(
        npu_inst_pe_1_5_6_n3), .ZN(npu_inst_pe_1_5_6_n58) );
  NOR2_X1 npu_inst_pe_1_5_6_U22 ( .A1(npu_inst_pe_1_5_6_n56), .A2(
        npu_inst_pe_1_5_6_n3), .ZN(npu_inst_pe_1_5_6_n54) );
  NOR2_X1 npu_inst_pe_1_5_6_U21 ( .A1(npu_inst_pe_1_5_6_n52), .A2(
        npu_inst_pe_1_5_6_n3), .ZN(npu_inst_pe_1_5_6_n50) );
  NOR2_X1 npu_inst_pe_1_5_6_U20 ( .A1(npu_inst_pe_1_5_6_n48), .A2(
        npu_inst_pe_1_5_6_n3), .ZN(npu_inst_pe_1_5_6_n46) );
  NOR2_X1 npu_inst_pe_1_5_6_U19 ( .A1(npu_inst_pe_1_5_6_n40), .A2(
        npu_inst_pe_1_5_6_n3), .ZN(npu_inst_pe_1_5_6_n38) );
  NOR2_X1 npu_inst_pe_1_5_6_U18 ( .A1(npu_inst_pe_1_5_6_n44), .A2(
        npu_inst_pe_1_5_6_n3), .ZN(npu_inst_pe_1_5_6_n42) );
  BUF_X1 npu_inst_pe_1_5_6_U17 ( .A(npu_inst_n96), .Z(npu_inst_pe_1_5_6_n8) );
  INV_X1 npu_inst_pe_1_5_6_U16 ( .A(npu_inst_n123), .ZN(npu_inst_pe_1_5_6_n12)
         );
  INV_X1 npu_inst_pe_1_5_6_U15 ( .A(npu_inst_pe_1_5_6_n38), .ZN(
        npu_inst_pe_1_5_6_n114) );
  INV_X1 npu_inst_pe_1_5_6_U14 ( .A(npu_inst_pe_1_5_6_n58), .ZN(
        npu_inst_pe_1_5_6_n119) );
  INV_X1 npu_inst_pe_1_5_6_U13 ( .A(npu_inst_pe_1_5_6_n54), .ZN(
        npu_inst_pe_1_5_6_n118) );
  INV_X1 npu_inst_pe_1_5_6_U12 ( .A(npu_inst_pe_1_5_6_n50), .ZN(
        npu_inst_pe_1_5_6_n117) );
  INV_X1 npu_inst_pe_1_5_6_U11 ( .A(npu_inst_pe_1_5_6_n46), .ZN(
        npu_inst_pe_1_5_6_n116) );
  INV_X1 npu_inst_pe_1_5_6_U10 ( .A(npu_inst_pe_1_5_6_n42), .ZN(
        npu_inst_pe_1_5_6_n115) );
  BUF_X1 npu_inst_pe_1_5_6_U9 ( .A(npu_inst_n15), .Z(npu_inst_pe_1_5_6_n2) );
  BUF_X1 npu_inst_pe_1_5_6_U8 ( .A(npu_inst_n15), .Z(npu_inst_pe_1_5_6_n1) );
  BUF_X1 npu_inst_pe_1_5_6_U7 ( .A(npu_inst_pe_1_5_6_n12), .Z(
        npu_inst_pe_1_5_6_n11) );
  BUF_X1 npu_inst_pe_1_5_6_U6 ( .A(npu_inst_pe_1_5_6_n12), .Z(
        npu_inst_pe_1_5_6_n10) );
  BUF_X1 npu_inst_pe_1_5_6_U5 ( .A(npu_inst_pe_1_5_6_n12), .Z(
        npu_inst_pe_1_5_6_n9) );
  NOR2_X1 npu_inst_pe_1_5_6_U4 ( .A1(npu_inst_pe_1_5_6_int_q_weight_0_), .A2(
        npu_inst_pe_1_5_6_n1), .ZN(npu_inst_pe_1_5_6_n76) );
  NOR2_X1 npu_inst_pe_1_5_6_U3 ( .A1(npu_inst_pe_1_5_6_n27), .A2(
        npu_inst_pe_1_5_6_n1), .ZN(npu_inst_pe_1_5_6_n77) );
  FA_X1 npu_inst_pe_1_5_6_sub_67_U2_1 ( .A(npu_inst_pe_1_5_6_int_q_acc_1_), 
        .B(npu_inst_pe_1_5_6_n14), .CI(npu_inst_pe_1_5_6_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_5_6_sub_67_carry_2_), .S(npu_inst_pe_1_5_6_N66) );
  FA_X1 npu_inst_pe_1_5_6_add_69_U1_1 ( .A(npu_inst_pe_1_5_6_int_q_acc_1_), 
        .B(npu_inst_pe_1_5_6_int_data_1_), .CI(
        npu_inst_pe_1_5_6_add_69_carry_1_), .CO(
        npu_inst_pe_1_5_6_add_69_carry_2_), .S(npu_inst_pe_1_5_6_N74) );
  NAND3_X1 npu_inst_pe_1_5_6_U109 ( .A1(npu_inst_pe_1_5_6_n5), .A2(
        npu_inst_pe_1_5_6_n7), .A3(npu_inst_pe_1_5_6_n8), .ZN(
        npu_inst_pe_1_5_6_n44) );
  NAND3_X1 npu_inst_pe_1_5_6_U108 ( .A1(npu_inst_pe_1_5_6_n4), .A2(
        npu_inst_pe_1_5_6_n7), .A3(npu_inst_pe_1_5_6_n8), .ZN(
        npu_inst_pe_1_5_6_n40) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_5_6_n34), .CK(
        npu_inst_pe_1_5_6_net3504), .RN(npu_inst_pe_1_5_6_n9), .Q(
        npu_inst_pe_1_5_6_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_5_6_n35), .CK(
        npu_inst_pe_1_5_6_net3504), .RN(npu_inst_pe_1_5_6_n9), .Q(
        npu_inst_pe_1_5_6_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_5_6_n36), .CK(
        npu_inst_pe_1_5_6_net3504), .RN(npu_inst_pe_1_5_6_n9), .Q(
        npu_inst_pe_1_5_6_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_5_6_n98), .CK(
        npu_inst_pe_1_5_6_net3504), .RN(npu_inst_pe_1_5_6_n9), .Q(
        npu_inst_pe_1_5_6_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_5_6_n99), .CK(
        npu_inst_pe_1_5_6_net3504), .RN(npu_inst_pe_1_5_6_n9), .Q(
        npu_inst_pe_1_5_6_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_5_6_n100), 
        .CK(npu_inst_pe_1_5_6_net3504), .RN(npu_inst_pe_1_5_6_n9), .Q(
        npu_inst_pe_1_5_6_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_5_6_n33), .CK(
        npu_inst_pe_1_5_6_net3504), .RN(npu_inst_pe_1_5_6_n9), .Q(
        npu_inst_pe_1_5_6_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_5_6_n101), 
        .CK(npu_inst_pe_1_5_6_net3504), .RN(npu_inst_pe_1_5_6_n9), .Q(
        npu_inst_pe_1_5_6_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_weight_reg_0_ ( .D(npu_inst_n109), .CK(
        npu_inst_pe_1_5_6_net3510), .RN(npu_inst_pe_1_5_6_n9), .Q(
        npu_inst_pe_1_5_6_int_q_weight_0_), .QN(npu_inst_pe_1_5_6_n27) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_weight_reg_1_ ( .D(npu_inst_n115), .CK(
        npu_inst_pe_1_5_6_net3510), .RN(npu_inst_pe_1_5_6_n9), .Q(
        npu_inst_pe_1_5_6_int_q_weight_1_), .QN(npu_inst_pe_1_5_6_n26) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_5_6_n113), 
        .CK(npu_inst_pe_1_5_6_net3510), .RN(npu_inst_pe_1_5_6_n9), .Q(
        npu_inst_pe_1_5_6_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_5_6_n107), 
        .CK(npu_inst_pe_1_5_6_net3510), .RN(npu_inst_pe_1_5_6_n9), .Q(
        npu_inst_pe_1_5_6_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_5_6_n112), 
        .CK(npu_inst_pe_1_5_6_net3510), .RN(npu_inst_pe_1_5_6_n10), .Q(
        npu_inst_pe_1_5_6_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_5_6_n106), 
        .CK(npu_inst_pe_1_5_6_net3510), .RN(npu_inst_pe_1_5_6_n10), .Q(
        npu_inst_pe_1_5_6_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_5_6_n111), 
        .CK(npu_inst_pe_1_5_6_net3510), .RN(npu_inst_pe_1_5_6_n10), .Q(
        npu_inst_pe_1_5_6_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_5_6_n105), 
        .CK(npu_inst_pe_1_5_6_net3510), .RN(npu_inst_pe_1_5_6_n10), .Q(
        npu_inst_pe_1_5_6_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_5_6_n110), 
        .CK(npu_inst_pe_1_5_6_net3510), .RN(npu_inst_pe_1_5_6_n10), .Q(
        npu_inst_pe_1_5_6_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_5_6_n104), 
        .CK(npu_inst_pe_1_5_6_net3510), .RN(npu_inst_pe_1_5_6_n10), .Q(
        npu_inst_pe_1_5_6_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_5_6_n109), 
        .CK(npu_inst_pe_1_5_6_net3510), .RN(npu_inst_pe_1_5_6_n10), .Q(
        npu_inst_pe_1_5_6_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_5_6_n103), 
        .CK(npu_inst_pe_1_5_6_net3510), .RN(npu_inst_pe_1_5_6_n10), .Q(
        npu_inst_pe_1_5_6_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_5_6_n108), 
        .CK(npu_inst_pe_1_5_6_net3510), .RN(npu_inst_pe_1_5_6_n10), .Q(
        npu_inst_pe_1_5_6_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_5_6_n102), 
        .CK(npu_inst_pe_1_5_6_net3510), .RN(npu_inst_pe_1_5_6_n10), .Q(
        npu_inst_pe_1_5_6_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_5_6_n86), 
        .CK(npu_inst_pe_1_5_6_net3510), .RN(npu_inst_pe_1_5_6_n10), .Q(
        npu_inst_pe_1_5_6_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_5_6_n87), 
        .CK(npu_inst_pe_1_5_6_net3510), .RN(npu_inst_pe_1_5_6_n10), .Q(
        npu_inst_pe_1_5_6_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_5_6_n88), 
        .CK(npu_inst_pe_1_5_6_net3510), .RN(npu_inst_pe_1_5_6_n11), .Q(
        npu_inst_pe_1_5_6_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_5_6_n89), 
        .CK(npu_inst_pe_1_5_6_net3510), .RN(npu_inst_pe_1_5_6_n11), .Q(
        npu_inst_pe_1_5_6_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_5_6_n90), 
        .CK(npu_inst_pe_1_5_6_net3510), .RN(npu_inst_pe_1_5_6_n11), .Q(
        npu_inst_pe_1_5_6_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_5_6_n91), 
        .CK(npu_inst_pe_1_5_6_net3510), .RN(npu_inst_pe_1_5_6_n11), .Q(
        npu_inst_pe_1_5_6_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_5_6_n92), 
        .CK(npu_inst_pe_1_5_6_net3510), .RN(npu_inst_pe_1_5_6_n11), .Q(
        npu_inst_pe_1_5_6_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_5_6_n93), 
        .CK(npu_inst_pe_1_5_6_net3510), .RN(npu_inst_pe_1_5_6_n11), .Q(
        npu_inst_pe_1_5_6_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_5_6_n94), 
        .CK(npu_inst_pe_1_5_6_net3510), .RN(npu_inst_pe_1_5_6_n11), .Q(
        npu_inst_pe_1_5_6_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_5_6_n95), 
        .CK(npu_inst_pe_1_5_6_net3510), .RN(npu_inst_pe_1_5_6_n11), .Q(
        npu_inst_pe_1_5_6_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_5_6_n96), 
        .CK(npu_inst_pe_1_5_6_net3510), .RN(npu_inst_pe_1_5_6_n11), .Q(
        npu_inst_pe_1_5_6_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_5_6_n97), 
        .CK(npu_inst_pe_1_5_6_net3510), .RN(npu_inst_pe_1_5_6_n11), .Q(
        npu_inst_pe_1_5_6_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_5_6_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_5_6_N84), .SE(1'b0), .GCK(npu_inst_pe_1_5_6_net3504) );
  CLKGATETST_X1 npu_inst_pe_1_5_6_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n62), .SE(1'b0), .GCK(npu_inst_pe_1_5_6_net3510) );
  MUX2_X1 npu_inst_pe_1_5_7_U162 ( .A(npu_inst_pe_1_5_7_n32), .B(
        npu_inst_pe_1_5_7_n29), .S(npu_inst_pe_1_5_7_n8), .Z(
        npu_inst_pe_1_5_7_N93) );
  MUX2_X1 npu_inst_pe_1_5_7_U161 ( .A(npu_inst_pe_1_5_7_n31), .B(
        npu_inst_pe_1_5_7_n30), .S(npu_inst_pe_1_5_7_n6), .Z(
        npu_inst_pe_1_5_7_n32) );
  MUX2_X1 npu_inst_pe_1_5_7_U160 ( .A(npu_inst_pe_1_5_7_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_5_7_int_q_reg_v_1__0_), .S(npu_inst_pe_1_5_7_n4), .Z(
        npu_inst_pe_1_5_7_n31) );
  MUX2_X1 npu_inst_pe_1_5_7_U159 ( .A(npu_inst_pe_1_5_7_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_5_7_int_q_reg_v_3__0_), .S(npu_inst_pe_1_5_7_n4), .Z(
        npu_inst_pe_1_5_7_n30) );
  MUX2_X1 npu_inst_pe_1_5_7_U158 ( .A(npu_inst_pe_1_5_7_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_5_7_int_q_reg_v_5__0_), .S(npu_inst_pe_1_5_7_n4), .Z(
        npu_inst_pe_1_5_7_n29) );
  MUX2_X1 npu_inst_pe_1_5_7_U157 ( .A(npu_inst_pe_1_5_7_n28), .B(
        npu_inst_pe_1_5_7_n23), .S(npu_inst_pe_1_5_7_n8), .Z(
        npu_inst_pe_1_5_7_N94) );
  MUX2_X1 npu_inst_pe_1_5_7_U156 ( .A(npu_inst_pe_1_5_7_n25), .B(
        npu_inst_pe_1_5_7_n24), .S(npu_inst_pe_1_5_7_n6), .Z(
        npu_inst_pe_1_5_7_n28) );
  MUX2_X1 npu_inst_pe_1_5_7_U155 ( .A(npu_inst_pe_1_5_7_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_5_7_int_q_reg_v_1__1_), .S(npu_inst_pe_1_5_7_n4), .Z(
        npu_inst_pe_1_5_7_n25) );
  MUX2_X1 npu_inst_pe_1_5_7_U154 ( .A(npu_inst_pe_1_5_7_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_5_7_int_q_reg_v_3__1_), .S(npu_inst_pe_1_5_7_n4), .Z(
        npu_inst_pe_1_5_7_n24) );
  MUX2_X1 npu_inst_pe_1_5_7_U153 ( .A(npu_inst_pe_1_5_7_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_5_7_int_q_reg_v_5__1_), .S(npu_inst_pe_1_5_7_n4), .Z(
        npu_inst_pe_1_5_7_n23) );
  MUX2_X1 npu_inst_pe_1_5_7_U152 ( .A(npu_inst_pe_1_5_7_n22), .B(
        npu_inst_pe_1_5_7_n19), .S(npu_inst_pe_1_5_7_n8), .Z(
        npu_inst_int_data_x_5__7__1_) );
  MUX2_X1 npu_inst_pe_1_5_7_U151 ( .A(npu_inst_pe_1_5_7_n21), .B(
        npu_inst_pe_1_5_7_n20), .S(npu_inst_pe_1_5_7_n6), .Z(
        npu_inst_pe_1_5_7_n22) );
  MUX2_X1 npu_inst_pe_1_5_7_U150 ( .A(npu_inst_pe_1_5_7_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_5_7_int_q_reg_h_1__1_), .S(npu_inst_pe_1_5_7_n4), .Z(
        npu_inst_pe_1_5_7_n21) );
  MUX2_X1 npu_inst_pe_1_5_7_U149 ( .A(npu_inst_pe_1_5_7_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_5_7_int_q_reg_h_3__1_), .S(npu_inst_pe_1_5_7_n4), .Z(
        npu_inst_pe_1_5_7_n20) );
  MUX2_X1 npu_inst_pe_1_5_7_U148 ( .A(npu_inst_pe_1_5_7_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_5_7_int_q_reg_h_5__1_), .S(npu_inst_pe_1_5_7_n4), .Z(
        npu_inst_pe_1_5_7_n19) );
  MUX2_X1 npu_inst_pe_1_5_7_U147 ( .A(npu_inst_pe_1_5_7_n18), .B(
        npu_inst_pe_1_5_7_n15), .S(npu_inst_pe_1_5_7_n8), .Z(
        npu_inst_int_data_x_5__7__0_) );
  MUX2_X1 npu_inst_pe_1_5_7_U146 ( .A(npu_inst_pe_1_5_7_n17), .B(
        npu_inst_pe_1_5_7_n16), .S(npu_inst_pe_1_5_7_n6), .Z(
        npu_inst_pe_1_5_7_n18) );
  MUX2_X1 npu_inst_pe_1_5_7_U145 ( .A(npu_inst_pe_1_5_7_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_5_7_int_q_reg_h_1__0_), .S(npu_inst_pe_1_5_7_n4), .Z(
        npu_inst_pe_1_5_7_n17) );
  MUX2_X1 npu_inst_pe_1_5_7_U144 ( .A(npu_inst_pe_1_5_7_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_5_7_int_q_reg_h_3__0_), .S(npu_inst_pe_1_5_7_n4), .Z(
        npu_inst_pe_1_5_7_n16) );
  MUX2_X1 npu_inst_pe_1_5_7_U143 ( .A(npu_inst_pe_1_5_7_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_5_7_int_q_reg_h_5__0_), .S(npu_inst_pe_1_5_7_n4), .Z(
        npu_inst_pe_1_5_7_n15) );
  XOR2_X1 npu_inst_pe_1_5_7_U142 ( .A(npu_inst_pe_1_5_7_int_data_0_), .B(
        npu_inst_pe_1_5_7_int_q_acc_0_), .Z(npu_inst_pe_1_5_7_N73) );
  AND2_X1 npu_inst_pe_1_5_7_U141 ( .A1(npu_inst_pe_1_5_7_int_q_acc_0_), .A2(
        npu_inst_pe_1_5_7_int_data_0_), .ZN(npu_inst_pe_1_5_7_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_5_7_U140 ( .A(npu_inst_pe_1_5_7_int_q_acc_0_), .B(
        npu_inst_pe_1_5_7_n13), .ZN(npu_inst_pe_1_5_7_N65) );
  OR2_X1 npu_inst_pe_1_5_7_U139 ( .A1(npu_inst_pe_1_5_7_n13), .A2(
        npu_inst_pe_1_5_7_int_q_acc_0_), .ZN(npu_inst_pe_1_5_7_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_5_7_U138 ( .A(npu_inst_pe_1_5_7_int_q_acc_2_), .B(
        npu_inst_pe_1_5_7_add_69_carry_2_), .Z(npu_inst_pe_1_5_7_N75) );
  AND2_X1 npu_inst_pe_1_5_7_U137 ( .A1(npu_inst_pe_1_5_7_add_69_carry_2_), 
        .A2(npu_inst_pe_1_5_7_int_q_acc_2_), .ZN(
        npu_inst_pe_1_5_7_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_5_7_U136 ( .A(npu_inst_pe_1_5_7_int_q_acc_3_), .B(
        npu_inst_pe_1_5_7_add_69_carry_3_), .Z(npu_inst_pe_1_5_7_N76) );
  AND2_X1 npu_inst_pe_1_5_7_U135 ( .A1(npu_inst_pe_1_5_7_add_69_carry_3_), 
        .A2(npu_inst_pe_1_5_7_int_q_acc_3_), .ZN(
        npu_inst_pe_1_5_7_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_5_7_U134 ( .A(npu_inst_pe_1_5_7_int_q_acc_4_), .B(
        npu_inst_pe_1_5_7_add_69_carry_4_), .Z(npu_inst_pe_1_5_7_N77) );
  AND2_X1 npu_inst_pe_1_5_7_U133 ( .A1(npu_inst_pe_1_5_7_add_69_carry_4_), 
        .A2(npu_inst_pe_1_5_7_int_q_acc_4_), .ZN(
        npu_inst_pe_1_5_7_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_5_7_U132 ( .A(npu_inst_pe_1_5_7_int_q_acc_5_), .B(
        npu_inst_pe_1_5_7_add_69_carry_5_), .Z(npu_inst_pe_1_5_7_N78) );
  AND2_X1 npu_inst_pe_1_5_7_U131 ( .A1(npu_inst_pe_1_5_7_add_69_carry_5_), 
        .A2(npu_inst_pe_1_5_7_int_q_acc_5_), .ZN(
        npu_inst_pe_1_5_7_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_5_7_U130 ( .A(npu_inst_pe_1_5_7_int_q_acc_6_), .B(
        npu_inst_pe_1_5_7_add_69_carry_6_), .Z(npu_inst_pe_1_5_7_N79) );
  AND2_X1 npu_inst_pe_1_5_7_U129 ( .A1(npu_inst_pe_1_5_7_add_69_carry_6_), 
        .A2(npu_inst_pe_1_5_7_int_q_acc_6_), .ZN(
        npu_inst_pe_1_5_7_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_5_7_U128 ( .A(npu_inst_pe_1_5_7_int_q_acc_7_), .B(
        npu_inst_pe_1_5_7_add_69_carry_7_), .Z(npu_inst_pe_1_5_7_N80) );
  XNOR2_X1 npu_inst_pe_1_5_7_U127 ( .A(npu_inst_pe_1_5_7_sub_67_carry_2_), .B(
        npu_inst_pe_1_5_7_int_q_acc_2_), .ZN(npu_inst_pe_1_5_7_N67) );
  OR2_X1 npu_inst_pe_1_5_7_U126 ( .A1(npu_inst_pe_1_5_7_int_q_acc_2_), .A2(
        npu_inst_pe_1_5_7_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_5_7_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_5_7_U125 ( .A(npu_inst_pe_1_5_7_sub_67_carry_3_), .B(
        npu_inst_pe_1_5_7_int_q_acc_3_), .ZN(npu_inst_pe_1_5_7_N68) );
  OR2_X1 npu_inst_pe_1_5_7_U124 ( .A1(npu_inst_pe_1_5_7_int_q_acc_3_), .A2(
        npu_inst_pe_1_5_7_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_5_7_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_5_7_U123 ( .A(npu_inst_pe_1_5_7_sub_67_carry_4_), .B(
        npu_inst_pe_1_5_7_int_q_acc_4_), .ZN(npu_inst_pe_1_5_7_N69) );
  OR2_X1 npu_inst_pe_1_5_7_U122 ( .A1(npu_inst_pe_1_5_7_int_q_acc_4_), .A2(
        npu_inst_pe_1_5_7_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_5_7_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_5_7_U121 ( .A(npu_inst_pe_1_5_7_sub_67_carry_5_), .B(
        npu_inst_pe_1_5_7_int_q_acc_5_), .ZN(npu_inst_pe_1_5_7_N70) );
  OR2_X1 npu_inst_pe_1_5_7_U120 ( .A1(npu_inst_pe_1_5_7_int_q_acc_5_), .A2(
        npu_inst_pe_1_5_7_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_5_7_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_5_7_U119 ( .A(npu_inst_pe_1_5_7_sub_67_carry_6_), .B(
        npu_inst_pe_1_5_7_int_q_acc_6_), .ZN(npu_inst_pe_1_5_7_N71) );
  OR2_X1 npu_inst_pe_1_5_7_U118 ( .A1(npu_inst_pe_1_5_7_int_q_acc_6_), .A2(
        npu_inst_pe_1_5_7_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_5_7_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_5_7_U117 ( .A(npu_inst_pe_1_5_7_int_q_acc_7_), .B(
        npu_inst_pe_1_5_7_sub_67_carry_7_), .ZN(npu_inst_pe_1_5_7_N72) );
  INV_X1 npu_inst_pe_1_5_7_U116 ( .A(npu_inst_n76), .ZN(npu_inst_pe_1_5_7_n7)
         );
  INV_X1 npu_inst_pe_1_5_7_U115 ( .A(npu_inst_pe_1_5_7_n7), .ZN(
        npu_inst_pe_1_5_7_n6) );
  INV_X1 npu_inst_pe_1_5_7_U114 ( .A(npu_inst_n54), .ZN(npu_inst_pe_1_5_7_n3)
         );
  AOI22_X1 npu_inst_pe_1_5_7_U113 ( .A1(npu_inst_int_data_y_6__7__0_), .A2(
        npu_inst_pe_1_5_7_n58), .B1(npu_inst_pe_1_5_7_n119), .B2(
        npu_inst_pe_1_5_7_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_5_7_n57) );
  INV_X1 npu_inst_pe_1_5_7_U112 ( .A(npu_inst_pe_1_5_7_n57), .ZN(
        npu_inst_pe_1_5_7_n108) );
  AOI22_X1 npu_inst_pe_1_5_7_U111 ( .A1(npu_inst_int_data_y_6__7__0_), .A2(
        npu_inst_pe_1_5_7_n54), .B1(npu_inst_pe_1_5_7_n118), .B2(
        npu_inst_pe_1_5_7_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_5_7_n53) );
  INV_X1 npu_inst_pe_1_5_7_U110 ( .A(npu_inst_pe_1_5_7_n53), .ZN(
        npu_inst_pe_1_5_7_n109) );
  AOI22_X1 npu_inst_pe_1_5_7_U107 ( .A1(npu_inst_int_data_y_6__7__0_), .A2(
        npu_inst_pe_1_5_7_n50), .B1(npu_inst_pe_1_5_7_n117), .B2(
        npu_inst_pe_1_5_7_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_5_7_n49) );
  INV_X1 npu_inst_pe_1_5_7_U106 ( .A(npu_inst_pe_1_5_7_n49), .ZN(
        npu_inst_pe_1_5_7_n110) );
  AOI22_X1 npu_inst_pe_1_5_7_U105 ( .A1(npu_inst_int_data_y_6__7__0_), .A2(
        npu_inst_pe_1_5_7_n46), .B1(npu_inst_pe_1_5_7_n116), .B2(
        npu_inst_pe_1_5_7_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_5_7_n45) );
  INV_X1 npu_inst_pe_1_5_7_U104 ( .A(npu_inst_pe_1_5_7_n45), .ZN(
        npu_inst_pe_1_5_7_n111) );
  AOI22_X1 npu_inst_pe_1_5_7_U103 ( .A1(npu_inst_int_data_y_6__7__0_), .A2(
        npu_inst_pe_1_5_7_n42), .B1(npu_inst_pe_1_5_7_n115), .B2(
        npu_inst_pe_1_5_7_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_5_7_n41) );
  INV_X1 npu_inst_pe_1_5_7_U102 ( .A(npu_inst_pe_1_5_7_n41), .ZN(
        npu_inst_pe_1_5_7_n112) );
  AOI22_X1 npu_inst_pe_1_5_7_U101 ( .A1(npu_inst_int_data_y_6__7__1_), .A2(
        npu_inst_pe_1_5_7_n58), .B1(npu_inst_pe_1_5_7_n119), .B2(
        npu_inst_pe_1_5_7_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_5_7_n59) );
  INV_X1 npu_inst_pe_1_5_7_U100 ( .A(npu_inst_pe_1_5_7_n59), .ZN(
        npu_inst_pe_1_5_7_n102) );
  AOI22_X1 npu_inst_pe_1_5_7_U99 ( .A1(npu_inst_int_data_y_6__7__1_), .A2(
        npu_inst_pe_1_5_7_n54), .B1(npu_inst_pe_1_5_7_n118), .B2(
        npu_inst_pe_1_5_7_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_5_7_n55) );
  INV_X1 npu_inst_pe_1_5_7_U98 ( .A(npu_inst_pe_1_5_7_n55), .ZN(
        npu_inst_pe_1_5_7_n103) );
  AOI22_X1 npu_inst_pe_1_5_7_U97 ( .A1(npu_inst_int_data_y_6__7__1_), .A2(
        npu_inst_pe_1_5_7_n50), .B1(npu_inst_pe_1_5_7_n117), .B2(
        npu_inst_pe_1_5_7_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_5_7_n51) );
  INV_X1 npu_inst_pe_1_5_7_U96 ( .A(npu_inst_pe_1_5_7_n51), .ZN(
        npu_inst_pe_1_5_7_n104) );
  AOI22_X1 npu_inst_pe_1_5_7_U95 ( .A1(npu_inst_int_data_y_6__7__1_), .A2(
        npu_inst_pe_1_5_7_n46), .B1(npu_inst_pe_1_5_7_n116), .B2(
        npu_inst_pe_1_5_7_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_5_7_n47) );
  INV_X1 npu_inst_pe_1_5_7_U94 ( .A(npu_inst_pe_1_5_7_n47), .ZN(
        npu_inst_pe_1_5_7_n105) );
  AOI22_X1 npu_inst_pe_1_5_7_U93 ( .A1(npu_inst_int_data_y_6__7__1_), .A2(
        npu_inst_pe_1_5_7_n42), .B1(npu_inst_pe_1_5_7_n115), .B2(
        npu_inst_pe_1_5_7_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_5_7_n43) );
  INV_X1 npu_inst_pe_1_5_7_U92 ( .A(npu_inst_pe_1_5_7_n43), .ZN(
        npu_inst_pe_1_5_7_n106) );
  AOI22_X1 npu_inst_pe_1_5_7_U91 ( .A1(npu_inst_pe_1_5_7_n38), .A2(
        npu_inst_int_data_y_6__7__1_), .B1(npu_inst_pe_1_5_7_n114), .B2(
        npu_inst_pe_1_5_7_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_5_7_n39) );
  INV_X1 npu_inst_pe_1_5_7_U90 ( .A(npu_inst_pe_1_5_7_n39), .ZN(
        npu_inst_pe_1_5_7_n107) );
  AOI22_X1 npu_inst_pe_1_5_7_U89 ( .A1(npu_inst_pe_1_5_7_n38), .A2(
        npu_inst_int_data_y_6__7__0_), .B1(npu_inst_pe_1_5_7_n114), .B2(
        npu_inst_pe_1_5_7_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_5_7_n37) );
  INV_X1 npu_inst_pe_1_5_7_U88 ( .A(npu_inst_pe_1_5_7_n37), .ZN(
        npu_inst_pe_1_5_7_n113) );
  AND2_X1 npu_inst_pe_1_5_7_U87 ( .A1(npu_inst_pe_1_5_7_N93), .A2(npu_inst_n54), .ZN(npu_inst_int_data_y_5__7__0_) );
  AND2_X1 npu_inst_pe_1_5_7_U86 ( .A1(npu_inst_n54), .A2(npu_inst_pe_1_5_7_N94), .ZN(npu_inst_int_data_y_5__7__1_) );
  NOR3_X1 npu_inst_pe_1_5_7_U85 ( .A1(npu_inst_pe_1_5_7_n26), .A2(npu_inst_n54), .A3(npu_inst_int_ckg[16]), .ZN(npu_inst_pe_1_5_7_n85) );
  OR2_X1 npu_inst_pe_1_5_7_U84 ( .A1(npu_inst_pe_1_5_7_n85), .A2(
        npu_inst_pe_1_5_7_n2), .ZN(npu_inst_pe_1_5_7_N84) );
  AND2_X1 npu_inst_pe_1_5_7_U83 ( .A1(npu_inst_pe_1_5_7_int_q_acc_0_), .A2(
        npu_inst_pe_1_5_7_n1), .ZN(npu_inst_int_data_res_5__7__0_) );
  AND2_X1 npu_inst_pe_1_5_7_U82 ( .A1(npu_inst_pe_1_5_7_n2), .A2(
        npu_inst_pe_1_5_7_int_q_acc_7_), .ZN(npu_inst_int_data_res_5__7__7_)
         );
  AND2_X1 npu_inst_pe_1_5_7_U81 ( .A1(npu_inst_pe_1_5_7_int_q_acc_1_), .A2(
        npu_inst_pe_1_5_7_n1), .ZN(npu_inst_int_data_res_5__7__1_) );
  AND2_X1 npu_inst_pe_1_5_7_U80 ( .A1(npu_inst_pe_1_5_7_int_q_acc_2_), .A2(
        npu_inst_pe_1_5_7_n1), .ZN(npu_inst_int_data_res_5__7__2_) );
  AND2_X1 npu_inst_pe_1_5_7_U79 ( .A1(npu_inst_pe_1_5_7_int_q_acc_3_), .A2(
        npu_inst_pe_1_5_7_n2), .ZN(npu_inst_int_data_res_5__7__3_) );
  AND2_X1 npu_inst_pe_1_5_7_U78 ( .A1(npu_inst_pe_1_5_7_int_q_acc_4_), .A2(
        npu_inst_pe_1_5_7_n2), .ZN(npu_inst_int_data_res_5__7__4_) );
  AND2_X1 npu_inst_pe_1_5_7_U77 ( .A1(npu_inst_pe_1_5_7_int_q_acc_5_), .A2(
        npu_inst_pe_1_5_7_n2), .ZN(npu_inst_int_data_res_5__7__5_) );
  AND2_X1 npu_inst_pe_1_5_7_U76 ( .A1(npu_inst_pe_1_5_7_int_q_acc_6_), .A2(
        npu_inst_pe_1_5_7_n2), .ZN(npu_inst_int_data_res_5__7__6_) );
  AOI222_X1 npu_inst_pe_1_5_7_U75 ( .A1(npu_inst_int_data_res_6__7__0_), .A2(
        npu_inst_pe_1_5_7_n1), .B1(npu_inst_pe_1_5_7_N73), .B2(
        npu_inst_pe_1_5_7_n76), .C1(npu_inst_pe_1_5_7_N65), .C2(
        npu_inst_pe_1_5_7_n77), .ZN(npu_inst_pe_1_5_7_n84) );
  INV_X1 npu_inst_pe_1_5_7_U74 ( .A(npu_inst_pe_1_5_7_n84), .ZN(
        npu_inst_pe_1_5_7_n101) );
  AOI222_X1 npu_inst_pe_1_5_7_U73 ( .A1(npu_inst_int_data_res_6__7__7_), .A2(
        npu_inst_pe_1_5_7_n1), .B1(npu_inst_pe_1_5_7_N80), .B2(
        npu_inst_pe_1_5_7_n76), .C1(npu_inst_pe_1_5_7_N72), .C2(
        npu_inst_pe_1_5_7_n77), .ZN(npu_inst_pe_1_5_7_n75) );
  INV_X1 npu_inst_pe_1_5_7_U72 ( .A(npu_inst_pe_1_5_7_n75), .ZN(
        npu_inst_pe_1_5_7_n33) );
  AOI222_X1 npu_inst_pe_1_5_7_U71 ( .A1(npu_inst_int_data_res_6__7__1_), .A2(
        npu_inst_pe_1_5_7_n1), .B1(npu_inst_pe_1_5_7_N74), .B2(
        npu_inst_pe_1_5_7_n76), .C1(npu_inst_pe_1_5_7_N66), .C2(
        npu_inst_pe_1_5_7_n77), .ZN(npu_inst_pe_1_5_7_n83) );
  INV_X1 npu_inst_pe_1_5_7_U70 ( .A(npu_inst_pe_1_5_7_n83), .ZN(
        npu_inst_pe_1_5_7_n100) );
  AOI222_X1 npu_inst_pe_1_5_7_U69 ( .A1(npu_inst_int_data_res_6__7__2_), .A2(
        npu_inst_pe_1_5_7_n1), .B1(npu_inst_pe_1_5_7_N75), .B2(
        npu_inst_pe_1_5_7_n76), .C1(npu_inst_pe_1_5_7_N67), .C2(
        npu_inst_pe_1_5_7_n77), .ZN(npu_inst_pe_1_5_7_n82) );
  INV_X1 npu_inst_pe_1_5_7_U68 ( .A(npu_inst_pe_1_5_7_n82), .ZN(
        npu_inst_pe_1_5_7_n99) );
  AOI222_X1 npu_inst_pe_1_5_7_U67 ( .A1(npu_inst_int_data_res_6__7__3_), .A2(
        npu_inst_pe_1_5_7_n1), .B1(npu_inst_pe_1_5_7_N76), .B2(
        npu_inst_pe_1_5_7_n76), .C1(npu_inst_pe_1_5_7_N68), .C2(
        npu_inst_pe_1_5_7_n77), .ZN(npu_inst_pe_1_5_7_n81) );
  INV_X1 npu_inst_pe_1_5_7_U66 ( .A(npu_inst_pe_1_5_7_n81), .ZN(
        npu_inst_pe_1_5_7_n98) );
  AOI222_X1 npu_inst_pe_1_5_7_U65 ( .A1(npu_inst_int_data_res_6__7__4_), .A2(
        npu_inst_pe_1_5_7_n1), .B1(npu_inst_pe_1_5_7_N77), .B2(
        npu_inst_pe_1_5_7_n76), .C1(npu_inst_pe_1_5_7_N69), .C2(
        npu_inst_pe_1_5_7_n77), .ZN(npu_inst_pe_1_5_7_n80) );
  INV_X1 npu_inst_pe_1_5_7_U64 ( .A(npu_inst_pe_1_5_7_n80), .ZN(
        npu_inst_pe_1_5_7_n36) );
  AOI222_X1 npu_inst_pe_1_5_7_U63 ( .A1(npu_inst_int_data_res_6__7__5_), .A2(
        npu_inst_pe_1_5_7_n1), .B1(npu_inst_pe_1_5_7_N78), .B2(
        npu_inst_pe_1_5_7_n76), .C1(npu_inst_pe_1_5_7_N70), .C2(
        npu_inst_pe_1_5_7_n77), .ZN(npu_inst_pe_1_5_7_n79) );
  INV_X1 npu_inst_pe_1_5_7_U62 ( .A(npu_inst_pe_1_5_7_n79), .ZN(
        npu_inst_pe_1_5_7_n35) );
  AOI222_X1 npu_inst_pe_1_5_7_U61 ( .A1(npu_inst_int_data_res_6__7__6_), .A2(
        npu_inst_pe_1_5_7_n1), .B1(npu_inst_pe_1_5_7_N79), .B2(
        npu_inst_pe_1_5_7_n76), .C1(npu_inst_pe_1_5_7_N71), .C2(
        npu_inst_pe_1_5_7_n77), .ZN(npu_inst_pe_1_5_7_n78) );
  INV_X1 npu_inst_pe_1_5_7_U60 ( .A(npu_inst_pe_1_5_7_n78), .ZN(
        npu_inst_pe_1_5_7_n34) );
  INV_X1 npu_inst_pe_1_5_7_U59 ( .A(npu_inst_pe_1_5_7_int_data_1_), .ZN(
        npu_inst_pe_1_5_7_n14) );
  AND2_X1 npu_inst_pe_1_5_7_U58 ( .A1(npu_inst_int_data_x_5__7__1_), .A2(
        npu_inst_pe_1_5_7_int_q_weight_1_), .ZN(npu_inst_pe_1_5_7_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_5_7_U57 ( .A1(npu_inst_int_data_x_5__7__0_), .A2(
        npu_inst_pe_1_5_7_int_q_weight_1_), .ZN(npu_inst_pe_1_5_7_int_data_0_)
         );
  NAND2_X1 npu_inst_pe_1_5_7_U56 ( .A1(npu_inst_pe_1_5_7_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_5_7_n60), .ZN(npu_inst_pe_1_5_7_n74) );
  OAI21_X1 npu_inst_pe_1_5_7_U55 ( .B1(npu_inst_pe_1_5_7_n63), .B2(
        npu_inst_pe_1_5_7_n60), .A(npu_inst_pe_1_5_7_n74), .ZN(
        npu_inst_pe_1_5_7_n97) );
  NAND2_X1 npu_inst_pe_1_5_7_U54 ( .A1(npu_inst_pe_1_5_7_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_5_7_n60), .ZN(npu_inst_pe_1_5_7_n73) );
  OAI21_X1 npu_inst_pe_1_5_7_U53 ( .B1(npu_inst_pe_1_5_7_n61), .B2(
        npu_inst_pe_1_5_7_n60), .A(npu_inst_pe_1_5_7_n73), .ZN(
        npu_inst_pe_1_5_7_n96) );
  NAND2_X1 npu_inst_pe_1_5_7_U52 ( .A1(npu_inst_pe_1_5_7_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_5_7_n56), .ZN(npu_inst_pe_1_5_7_n72) );
  OAI21_X1 npu_inst_pe_1_5_7_U51 ( .B1(npu_inst_pe_1_5_7_n63), .B2(
        npu_inst_pe_1_5_7_n56), .A(npu_inst_pe_1_5_7_n72), .ZN(
        npu_inst_pe_1_5_7_n95) );
  NAND2_X1 npu_inst_pe_1_5_7_U50 ( .A1(npu_inst_pe_1_5_7_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_5_7_n56), .ZN(npu_inst_pe_1_5_7_n71) );
  OAI21_X1 npu_inst_pe_1_5_7_U49 ( .B1(npu_inst_pe_1_5_7_n61), .B2(
        npu_inst_pe_1_5_7_n56), .A(npu_inst_pe_1_5_7_n71), .ZN(
        npu_inst_pe_1_5_7_n94) );
  NAND2_X1 npu_inst_pe_1_5_7_U48 ( .A1(npu_inst_pe_1_5_7_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_5_7_n52), .ZN(npu_inst_pe_1_5_7_n70) );
  OAI21_X1 npu_inst_pe_1_5_7_U47 ( .B1(npu_inst_pe_1_5_7_n63), .B2(
        npu_inst_pe_1_5_7_n52), .A(npu_inst_pe_1_5_7_n70), .ZN(
        npu_inst_pe_1_5_7_n93) );
  NAND2_X1 npu_inst_pe_1_5_7_U46 ( .A1(npu_inst_pe_1_5_7_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_5_7_n52), .ZN(npu_inst_pe_1_5_7_n69) );
  OAI21_X1 npu_inst_pe_1_5_7_U45 ( .B1(npu_inst_pe_1_5_7_n61), .B2(
        npu_inst_pe_1_5_7_n52), .A(npu_inst_pe_1_5_7_n69), .ZN(
        npu_inst_pe_1_5_7_n92) );
  NAND2_X1 npu_inst_pe_1_5_7_U44 ( .A1(npu_inst_pe_1_5_7_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_5_7_n48), .ZN(npu_inst_pe_1_5_7_n68) );
  OAI21_X1 npu_inst_pe_1_5_7_U43 ( .B1(npu_inst_pe_1_5_7_n63), .B2(
        npu_inst_pe_1_5_7_n48), .A(npu_inst_pe_1_5_7_n68), .ZN(
        npu_inst_pe_1_5_7_n91) );
  NAND2_X1 npu_inst_pe_1_5_7_U42 ( .A1(npu_inst_pe_1_5_7_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_5_7_n48), .ZN(npu_inst_pe_1_5_7_n67) );
  OAI21_X1 npu_inst_pe_1_5_7_U41 ( .B1(npu_inst_pe_1_5_7_n61), .B2(
        npu_inst_pe_1_5_7_n48), .A(npu_inst_pe_1_5_7_n67), .ZN(
        npu_inst_pe_1_5_7_n90) );
  NAND2_X1 npu_inst_pe_1_5_7_U40 ( .A1(npu_inst_pe_1_5_7_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_5_7_n44), .ZN(npu_inst_pe_1_5_7_n66) );
  OAI21_X1 npu_inst_pe_1_5_7_U39 ( .B1(npu_inst_pe_1_5_7_n63), .B2(
        npu_inst_pe_1_5_7_n44), .A(npu_inst_pe_1_5_7_n66), .ZN(
        npu_inst_pe_1_5_7_n89) );
  NAND2_X1 npu_inst_pe_1_5_7_U38 ( .A1(npu_inst_pe_1_5_7_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_5_7_n44), .ZN(npu_inst_pe_1_5_7_n65) );
  OAI21_X1 npu_inst_pe_1_5_7_U37 ( .B1(npu_inst_pe_1_5_7_n61), .B2(
        npu_inst_pe_1_5_7_n44), .A(npu_inst_pe_1_5_7_n65), .ZN(
        npu_inst_pe_1_5_7_n88) );
  NAND2_X1 npu_inst_pe_1_5_7_U36 ( .A1(npu_inst_pe_1_5_7_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_5_7_n40), .ZN(npu_inst_pe_1_5_7_n64) );
  OAI21_X1 npu_inst_pe_1_5_7_U35 ( .B1(npu_inst_pe_1_5_7_n63), .B2(
        npu_inst_pe_1_5_7_n40), .A(npu_inst_pe_1_5_7_n64), .ZN(
        npu_inst_pe_1_5_7_n87) );
  NAND2_X1 npu_inst_pe_1_5_7_U34 ( .A1(npu_inst_pe_1_5_7_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_5_7_n40), .ZN(npu_inst_pe_1_5_7_n62) );
  OAI21_X1 npu_inst_pe_1_5_7_U33 ( .B1(npu_inst_pe_1_5_7_n61), .B2(
        npu_inst_pe_1_5_7_n40), .A(npu_inst_pe_1_5_7_n62), .ZN(
        npu_inst_pe_1_5_7_n86) );
  INV_X1 npu_inst_pe_1_5_7_U32 ( .A(npu_inst_pe_1_5_7_int_data_0_), .ZN(
        npu_inst_pe_1_5_7_n13) );
  INV_X1 npu_inst_pe_1_5_7_U31 ( .A(npu_inst_n68), .ZN(npu_inst_pe_1_5_7_n5)
         );
  AOI22_X1 npu_inst_pe_1_5_7_U30 ( .A1(npu_inst_n54), .A2(
        npu_inst_int_data_y_6__7__1_), .B1(npu_inst_pe_1_5_7_n3), .B2(
        int_i_data_h_npu[5]), .ZN(npu_inst_pe_1_5_7_n63) );
  AOI22_X1 npu_inst_pe_1_5_7_U29 ( .A1(npu_inst_n54), .A2(
        npu_inst_int_data_y_6__7__0_), .B1(npu_inst_pe_1_5_7_n3), .B2(
        int_i_data_h_npu[4]), .ZN(npu_inst_pe_1_5_7_n61) );
  OR3_X1 npu_inst_pe_1_5_7_U28 ( .A1(npu_inst_pe_1_5_7_n6), .A2(
        npu_inst_pe_1_5_7_n8), .A3(npu_inst_pe_1_5_7_n5), .ZN(
        npu_inst_pe_1_5_7_n56) );
  OR3_X1 npu_inst_pe_1_5_7_U27 ( .A1(npu_inst_pe_1_5_7_n5), .A2(
        npu_inst_pe_1_5_7_n8), .A3(npu_inst_pe_1_5_7_n7), .ZN(
        npu_inst_pe_1_5_7_n48) );
  INV_X1 npu_inst_pe_1_5_7_U26 ( .A(npu_inst_pe_1_5_7_n5), .ZN(
        npu_inst_pe_1_5_7_n4) );
  OR3_X1 npu_inst_pe_1_5_7_U25 ( .A1(npu_inst_pe_1_5_7_n4), .A2(
        npu_inst_pe_1_5_7_n8), .A3(npu_inst_pe_1_5_7_n7), .ZN(
        npu_inst_pe_1_5_7_n52) );
  OR3_X1 npu_inst_pe_1_5_7_U24 ( .A1(npu_inst_pe_1_5_7_n6), .A2(
        npu_inst_pe_1_5_7_n8), .A3(npu_inst_pe_1_5_7_n4), .ZN(
        npu_inst_pe_1_5_7_n60) );
  NOR2_X1 npu_inst_pe_1_5_7_U23 ( .A1(npu_inst_pe_1_5_7_n60), .A2(
        npu_inst_pe_1_5_7_n3), .ZN(npu_inst_pe_1_5_7_n58) );
  NOR2_X1 npu_inst_pe_1_5_7_U22 ( .A1(npu_inst_pe_1_5_7_n56), .A2(
        npu_inst_pe_1_5_7_n3), .ZN(npu_inst_pe_1_5_7_n54) );
  NOR2_X1 npu_inst_pe_1_5_7_U21 ( .A1(npu_inst_pe_1_5_7_n52), .A2(
        npu_inst_pe_1_5_7_n3), .ZN(npu_inst_pe_1_5_7_n50) );
  NOR2_X1 npu_inst_pe_1_5_7_U20 ( .A1(npu_inst_pe_1_5_7_n48), .A2(
        npu_inst_pe_1_5_7_n3), .ZN(npu_inst_pe_1_5_7_n46) );
  NOR2_X1 npu_inst_pe_1_5_7_U19 ( .A1(npu_inst_pe_1_5_7_n40), .A2(
        npu_inst_pe_1_5_7_n3), .ZN(npu_inst_pe_1_5_7_n38) );
  NOR2_X1 npu_inst_pe_1_5_7_U18 ( .A1(npu_inst_pe_1_5_7_n44), .A2(
        npu_inst_pe_1_5_7_n3), .ZN(npu_inst_pe_1_5_7_n42) );
  BUF_X1 npu_inst_pe_1_5_7_U17 ( .A(npu_inst_n96), .Z(npu_inst_pe_1_5_7_n8) );
  INV_X1 npu_inst_pe_1_5_7_U16 ( .A(npu_inst_n123), .ZN(npu_inst_pe_1_5_7_n12)
         );
  INV_X1 npu_inst_pe_1_5_7_U15 ( .A(npu_inst_pe_1_5_7_n38), .ZN(
        npu_inst_pe_1_5_7_n114) );
  INV_X1 npu_inst_pe_1_5_7_U14 ( .A(npu_inst_pe_1_5_7_n58), .ZN(
        npu_inst_pe_1_5_7_n119) );
  INV_X1 npu_inst_pe_1_5_7_U13 ( .A(npu_inst_pe_1_5_7_n54), .ZN(
        npu_inst_pe_1_5_7_n118) );
  INV_X1 npu_inst_pe_1_5_7_U12 ( .A(npu_inst_pe_1_5_7_n50), .ZN(
        npu_inst_pe_1_5_7_n117) );
  INV_X1 npu_inst_pe_1_5_7_U11 ( .A(npu_inst_pe_1_5_7_n46), .ZN(
        npu_inst_pe_1_5_7_n116) );
  INV_X1 npu_inst_pe_1_5_7_U10 ( .A(npu_inst_pe_1_5_7_n42), .ZN(
        npu_inst_pe_1_5_7_n115) );
  BUF_X1 npu_inst_pe_1_5_7_U9 ( .A(npu_inst_n15), .Z(npu_inst_pe_1_5_7_n2) );
  BUF_X1 npu_inst_pe_1_5_7_U8 ( .A(npu_inst_n15), .Z(npu_inst_pe_1_5_7_n1) );
  BUF_X1 npu_inst_pe_1_5_7_U7 ( .A(npu_inst_pe_1_5_7_n12), .Z(
        npu_inst_pe_1_5_7_n11) );
  BUF_X1 npu_inst_pe_1_5_7_U6 ( .A(npu_inst_pe_1_5_7_n12), .Z(
        npu_inst_pe_1_5_7_n10) );
  BUF_X1 npu_inst_pe_1_5_7_U5 ( .A(npu_inst_pe_1_5_7_n12), .Z(
        npu_inst_pe_1_5_7_n9) );
  NOR2_X1 npu_inst_pe_1_5_7_U4 ( .A1(npu_inst_pe_1_5_7_int_q_weight_0_), .A2(
        npu_inst_pe_1_5_7_n1), .ZN(npu_inst_pe_1_5_7_n76) );
  NOR2_X1 npu_inst_pe_1_5_7_U3 ( .A1(npu_inst_pe_1_5_7_n27), .A2(
        npu_inst_pe_1_5_7_n1), .ZN(npu_inst_pe_1_5_7_n77) );
  FA_X1 npu_inst_pe_1_5_7_sub_67_U2_1 ( .A(npu_inst_pe_1_5_7_int_q_acc_1_), 
        .B(npu_inst_pe_1_5_7_n14), .CI(npu_inst_pe_1_5_7_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_5_7_sub_67_carry_2_), .S(npu_inst_pe_1_5_7_N66) );
  FA_X1 npu_inst_pe_1_5_7_add_69_U1_1 ( .A(npu_inst_pe_1_5_7_int_q_acc_1_), 
        .B(npu_inst_pe_1_5_7_int_data_1_), .CI(
        npu_inst_pe_1_5_7_add_69_carry_1_), .CO(
        npu_inst_pe_1_5_7_add_69_carry_2_), .S(npu_inst_pe_1_5_7_N74) );
  NAND3_X1 npu_inst_pe_1_5_7_U109 ( .A1(npu_inst_pe_1_5_7_n5), .A2(
        npu_inst_pe_1_5_7_n7), .A3(npu_inst_pe_1_5_7_n8), .ZN(
        npu_inst_pe_1_5_7_n44) );
  NAND3_X1 npu_inst_pe_1_5_7_U108 ( .A1(npu_inst_pe_1_5_7_n4), .A2(
        npu_inst_pe_1_5_7_n7), .A3(npu_inst_pe_1_5_7_n8), .ZN(
        npu_inst_pe_1_5_7_n40) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_5_7_n34), .CK(
        npu_inst_pe_1_5_7_net3481), .RN(npu_inst_pe_1_5_7_n9), .Q(
        npu_inst_pe_1_5_7_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_5_7_n35), .CK(
        npu_inst_pe_1_5_7_net3481), .RN(npu_inst_pe_1_5_7_n9), .Q(
        npu_inst_pe_1_5_7_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_5_7_n36), .CK(
        npu_inst_pe_1_5_7_net3481), .RN(npu_inst_pe_1_5_7_n9), .Q(
        npu_inst_pe_1_5_7_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_5_7_n98), .CK(
        npu_inst_pe_1_5_7_net3481), .RN(npu_inst_pe_1_5_7_n9), .Q(
        npu_inst_pe_1_5_7_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_5_7_n99), .CK(
        npu_inst_pe_1_5_7_net3481), .RN(npu_inst_pe_1_5_7_n9), .Q(
        npu_inst_pe_1_5_7_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_5_7_n100), 
        .CK(npu_inst_pe_1_5_7_net3481), .RN(npu_inst_pe_1_5_7_n9), .Q(
        npu_inst_pe_1_5_7_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_5_7_n33), .CK(
        npu_inst_pe_1_5_7_net3481), .RN(npu_inst_pe_1_5_7_n9), .Q(
        npu_inst_pe_1_5_7_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_5_7_n101), 
        .CK(npu_inst_pe_1_5_7_net3481), .RN(npu_inst_pe_1_5_7_n9), .Q(
        npu_inst_pe_1_5_7_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_weight_reg_0_ ( .D(npu_inst_n109), .CK(
        npu_inst_pe_1_5_7_net3487), .RN(npu_inst_pe_1_5_7_n9), .Q(
        npu_inst_pe_1_5_7_int_q_weight_0_), .QN(npu_inst_pe_1_5_7_n27) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_weight_reg_1_ ( .D(npu_inst_n115), .CK(
        npu_inst_pe_1_5_7_net3487), .RN(npu_inst_pe_1_5_7_n9), .Q(
        npu_inst_pe_1_5_7_int_q_weight_1_), .QN(npu_inst_pe_1_5_7_n26) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_5_7_n113), 
        .CK(npu_inst_pe_1_5_7_net3487), .RN(npu_inst_pe_1_5_7_n9), .Q(
        npu_inst_pe_1_5_7_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_5_7_n107), 
        .CK(npu_inst_pe_1_5_7_net3487), .RN(npu_inst_pe_1_5_7_n9), .Q(
        npu_inst_pe_1_5_7_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_5_7_n112), 
        .CK(npu_inst_pe_1_5_7_net3487), .RN(npu_inst_pe_1_5_7_n10), .Q(
        npu_inst_pe_1_5_7_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_5_7_n106), 
        .CK(npu_inst_pe_1_5_7_net3487), .RN(npu_inst_pe_1_5_7_n10), .Q(
        npu_inst_pe_1_5_7_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_5_7_n111), 
        .CK(npu_inst_pe_1_5_7_net3487), .RN(npu_inst_pe_1_5_7_n10), .Q(
        npu_inst_pe_1_5_7_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_5_7_n105), 
        .CK(npu_inst_pe_1_5_7_net3487), .RN(npu_inst_pe_1_5_7_n10), .Q(
        npu_inst_pe_1_5_7_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_5_7_n110), 
        .CK(npu_inst_pe_1_5_7_net3487), .RN(npu_inst_pe_1_5_7_n10), .Q(
        npu_inst_pe_1_5_7_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_5_7_n104), 
        .CK(npu_inst_pe_1_5_7_net3487), .RN(npu_inst_pe_1_5_7_n10), .Q(
        npu_inst_pe_1_5_7_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_5_7_n109), 
        .CK(npu_inst_pe_1_5_7_net3487), .RN(npu_inst_pe_1_5_7_n10), .Q(
        npu_inst_pe_1_5_7_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_5_7_n103), 
        .CK(npu_inst_pe_1_5_7_net3487), .RN(npu_inst_pe_1_5_7_n10), .Q(
        npu_inst_pe_1_5_7_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_5_7_n108), 
        .CK(npu_inst_pe_1_5_7_net3487), .RN(npu_inst_pe_1_5_7_n10), .Q(
        npu_inst_pe_1_5_7_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_5_7_n102), 
        .CK(npu_inst_pe_1_5_7_net3487), .RN(npu_inst_pe_1_5_7_n10), .Q(
        npu_inst_pe_1_5_7_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_5_7_n86), 
        .CK(npu_inst_pe_1_5_7_net3487), .RN(npu_inst_pe_1_5_7_n10), .Q(
        npu_inst_pe_1_5_7_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_5_7_n87), 
        .CK(npu_inst_pe_1_5_7_net3487), .RN(npu_inst_pe_1_5_7_n10), .Q(
        npu_inst_pe_1_5_7_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_5_7_n88), 
        .CK(npu_inst_pe_1_5_7_net3487), .RN(npu_inst_pe_1_5_7_n11), .Q(
        npu_inst_pe_1_5_7_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_5_7_n89), 
        .CK(npu_inst_pe_1_5_7_net3487), .RN(npu_inst_pe_1_5_7_n11), .Q(
        npu_inst_pe_1_5_7_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_5_7_n90), 
        .CK(npu_inst_pe_1_5_7_net3487), .RN(npu_inst_pe_1_5_7_n11), .Q(
        npu_inst_pe_1_5_7_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_5_7_n91), 
        .CK(npu_inst_pe_1_5_7_net3487), .RN(npu_inst_pe_1_5_7_n11), .Q(
        npu_inst_pe_1_5_7_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_5_7_n92), 
        .CK(npu_inst_pe_1_5_7_net3487), .RN(npu_inst_pe_1_5_7_n11), .Q(
        npu_inst_pe_1_5_7_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_5_7_n93), 
        .CK(npu_inst_pe_1_5_7_net3487), .RN(npu_inst_pe_1_5_7_n11), .Q(
        npu_inst_pe_1_5_7_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_5_7_n94), 
        .CK(npu_inst_pe_1_5_7_net3487), .RN(npu_inst_pe_1_5_7_n11), .Q(
        npu_inst_pe_1_5_7_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_5_7_n95), 
        .CK(npu_inst_pe_1_5_7_net3487), .RN(npu_inst_pe_1_5_7_n11), .Q(
        npu_inst_pe_1_5_7_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_5_7_n96), 
        .CK(npu_inst_pe_1_5_7_net3487), .RN(npu_inst_pe_1_5_7_n11), .Q(
        npu_inst_pe_1_5_7_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_5_7_n97), 
        .CK(npu_inst_pe_1_5_7_net3487), .RN(npu_inst_pe_1_5_7_n11), .Q(
        npu_inst_pe_1_5_7_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_5_7_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_5_7_N84), .SE(1'b0), .GCK(npu_inst_pe_1_5_7_net3481) );
  CLKGATETST_X1 npu_inst_pe_1_5_7_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n62), .SE(1'b0), .GCK(npu_inst_pe_1_5_7_net3487) );
  MUX2_X1 npu_inst_pe_1_6_0_U162 ( .A(npu_inst_pe_1_6_0_n32), .B(
        npu_inst_pe_1_6_0_n29), .S(npu_inst_pe_1_6_0_n8), .Z(
        npu_inst_pe_1_6_0_N93) );
  MUX2_X1 npu_inst_pe_1_6_0_U161 ( .A(npu_inst_pe_1_6_0_n31), .B(
        npu_inst_pe_1_6_0_n30), .S(npu_inst_pe_1_6_0_n6), .Z(
        npu_inst_pe_1_6_0_n32) );
  MUX2_X1 npu_inst_pe_1_6_0_U160 ( .A(npu_inst_pe_1_6_0_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_6_0_int_q_reg_v_1__0_), .S(npu_inst_pe_1_6_0_n4), .Z(
        npu_inst_pe_1_6_0_n31) );
  MUX2_X1 npu_inst_pe_1_6_0_U159 ( .A(npu_inst_pe_1_6_0_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_6_0_int_q_reg_v_3__0_), .S(npu_inst_pe_1_6_0_n4), .Z(
        npu_inst_pe_1_6_0_n30) );
  MUX2_X1 npu_inst_pe_1_6_0_U158 ( .A(npu_inst_pe_1_6_0_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_6_0_int_q_reg_v_5__0_), .S(npu_inst_pe_1_6_0_n4), .Z(
        npu_inst_pe_1_6_0_n29) );
  MUX2_X1 npu_inst_pe_1_6_0_U157 ( .A(npu_inst_pe_1_6_0_n28), .B(
        npu_inst_pe_1_6_0_n23), .S(npu_inst_pe_1_6_0_n8), .Z(
        npu_inst_pe_1_6_0_N94) );
  MUX2_X1 npu_inst_pe_1_6_0_U156 ( .A(npu_inst_pe_1_6_0_n25), .B(
        npu_inst_pe_1_6_0_n24), .S(npu_inst_pe_1_6_0_n6), .Z(
        npu_inst_pe_1_6_0_n28) );
  MUX2_X1 npu_inst_pe_1_6_0_U155 ( .A(npu_inst_pe_1_6_0_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_6_0_int_q_reg_v_1__1_), .S(npu_inst_pe_1_6_0_n4), .Z(
        npu_inst_pe_1_6_0_n25) );
  MUX2_X1 npu_inst_pe_1_6_0_U154 ( .A(npu_inst_pe_1_6_0_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_6_0_int_q_reg_v_3__1_), .S(npu_inst_pe_1_6_0_n4), .Z(
        npu_inst_pe_1_6_0_n24) );
  MUX2_X1 npu_inst_pe_1_6_0_U153 ( .A(npu_inst_pe_1_6_0_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_6_0_int_q_reg_v_5__1_), .S(npu_inst_pe_1_6_0_n4), .Z(
        npu_inst_pe_1_6_0_n23) );
  MUX2_X1 npu_inst_pe_1_6_0_U152 ( .A(npu_inst_pe_1_6_0_n22), .B(
        npu_inst_pe_1_6_0_n19), .S(npu_inst_pe_1_6_0_n8), .Z(
        npu_inst_pe_1_6_0_o_data_h_1_) );
  MUX2_X1 npu_inst_pe_1_6_0_U151 ( .A(npu_inst_pe_1_6_0_n21), .B(
        npu_inst_pe_1_6_0_n20), .S(npu_inst_pe_1_6_0_n6), .Z(
        npu_inst_pe_1_6_0_n22) );
  MUX2_X1 npu_inst_pe_1_6_0_U150 ( .A(npu_inst_pe_1_6_0_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_6_0_int_q_reg_h_1__1_), .S(npu_inst_pe_1_6_0_n4), .Z(
        npu_inst_pe_1_6_0_n21) );
  MUX2_X1 npu_inst_pe_1_6_0_U149 ( .A(npu_inst_pe_1_6_0_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_6_0_int_q_reg_h_3__1_), .S(npu_inst_pe_1_6_0_n4), .Z(
        npu_inst_pe_1_6_0_n20) );
  MUX2_X1 npu_inst_pe_1_6_0_U148 ( .A(npu_inst_pe_1_6_0_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_6_0_int_q_reg_h_5__1_), .S(npu_inst_pe_1_6_0_n4), .Z(
        npu_inst_pe_1_6_0_n19) );
  MUX2_X1 npu_inst_pe_1_6_0_U147 ( .A(npu_inst_pe_1_6_0_n18), .B(
        npu_inst_pe_1_6_0_n15), .S(npu_inst_pe_1_6_0_n8), .Z(
        npu_inst_pe_1_6_0_o_data_h_0_) );
  MUX2_X1 npu_inst_pe_1_6_0_U146 ( .A(npu_inst_pe_1_6_0_n17), .B(
        npu_inst_pe_1_6_0_n16), .S(npu_inst_pe_1_6_0_n6), .Z(
        npu_inst_pe_1_6_0_n18) );
  MUX2_X1 npu_inst_pe_1_6_0_U145 ( .A(npu_inst_pe_1_6_0_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_6_0_int_q_reg_h_1__0_), .S(npu_inst_pe_1_6_0_n4), .Z(
        npu_inst_pe_1_6_0_n17) );
  MUX2_X1 npu_inst_pe_1_6_0_U144 ( .A(npu_inst_pe_1_6_0_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_6_0_int_q_reg_h_3__0_), .S(npu_inst_pe_1_6_0_n4), .Z(
        npu_inst_pe_1_6_0_n16) );
  MUX2_X1 npu_inst_pe_1_6_0_U143 ( .A(npu_inst_pe_1_6_0_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_6_0_int_q_reg_h_5__0_), .S(npu_inst_pe_1_6_0_n4), .Z(
        npu_inst_pe_1_6_0_n15) );
  XOR2_X1 npu_inst_pe_1_6_0_U142 ( .A(npu_inst_pe_1_6_0_int_data_0_), .B(
        npu_inst_pe_1_6_0_int_q_acc_0_), .Z(npu_inst_pe_1_6_0_N73) );
  AND2_X1 npu_inst_pe_1_6_0_U141 ( .A1(npu_inst_pe_1_6_0_int_q_acc_0_), .A2(
        npu_inst_pe_1_6_0_int_data_0_), .ZN(npu_inst_pe_1_6_0_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_6_0_U140 ( .A(npu_inst_pe_1_6_0_int_q_acc_0_), .B(
        npu_inst_pe_1_6_0_n13), .ZN(npu_inst_pe_1_6_0_N65) );
  OR2_X1 npu_inst_pe_1_6_0_U139 ( .A1(npu_inst_pe_1_6_0_n13), .A2(
        npu_inst_pe_1_6_0_int_q_acc_0_), .ZN(npu_inst_pe_1_6_0_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_6_0_U138 ( .A(npu_inst_pe_1_6_0_int_q_acc_2_), .B(
        npu_inst_pe_1_6_0_add_69_carry_2_), .Z(npu_inst_pe_1_6_0_N75) );
  AND2_X1 npu_inst_pe_1_6_0_U137 ( .A1(npu_inst_pe_1_6_0_add_69_carry_2_), 
        .A2(npu_inst_pe_1_6_0_int_q_acc_2_), .ZN(
        npu_inst_pe_1_6_0_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_6_0_U136 ( .A(npu_inst_pe_1_6_0_int_q_acc_3_), .B(
        npu_inst_pe_1_6_0_add_69_carry_3_), .Z(npu_inst_pe_1_6_0_N76) );
  AND2_X1 npu_inst_pe_1_6_0_U135 ( .A1(npu_inst_pe_1_6_0_add_69_carry_3_), 
        .A2(npu_inst_pe_1_6_0_int_q_acc_3_), .ZN(
        npu_inst_pe_1_6_0_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_6_0_U134 ( .A(npu_inst_pe_1_6_0_int_q_acc_4_), .B(
        npu_inst_pe_1_6_0_add_69_carry_4_), .Z(npu_inst_pe_1_6_0_N77) );
  AND2_X1 npu_inst_pe_1_6_0_U133 ( .A1(npu_inst_pe_1_6_0_add_69_carry_4_), 
        .A2(npu_inst_pe_1_6_0_int_q_acc_4_), .ZN(
        npu_inst_pe_1_6_0_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_6_0_U132 ( .A(npu_inst_pe_1_6_0_int_q_acc_5_), .B(
        npu_inst_pe_1_6_0_add_69_carry_5_), .Z(npu_inst_pe_1_6_0_N78) );
  AND2_X1 npu_inst_pe_1_6_0_U131 ( .A1(npu_inst_pe_1_6_0_add_69_carry_5_), 
        .A2(npu_inst_pe_1_6_0_int_q_acc_5_), .ZN(
        npu_inst_pe_1_6_0_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_6_0_U130 ( .A(npu_inst_pe_1_6_0_int_q_acc_6_), .B(
        npu_inst_pe_1_6_0_add_69_carry_6_), .Z(npu_inst_pe_1_6_0_N79) );
  AND2_X1 npu_inst_pe_1_6_0_U129 ( .A1(npu_inst_pe_1_6_0_add_69_carry_6_), 
        .A2(npu_inst_pe_1_6_0_int_q_acc_6_), .ZN(
        npu_inst_pe_1_6_0_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_6_0_U128 ( .A(npu_inst_pe_1_6_0_int_q_acc_7_), .B(
        npu_inst_pe_1_6_0_add_69_carry_7_), .Z(npu_inst_pe_1_6_0_N80) );
  XNOR2_X1 npu_inst_pe_1_6_0_U127 ( .A(npu_inst_pe_1_6_0_sub_67_carry_2_), .B(
        npu_inst_pe_1_6_0_int_q_acc_2_), .ZN(npu_inst_pe_1_6_0_N67) );
  OR2_X1 npu_inst_pe_1_6_0_U126 ( .A1(npu_inst_pe_1_6_0_int_q_acc_2_), .A2(
        npu_inst_pe_1_6_0_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_6_0_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_6_0_U125 ( .A(npu_inst_pe_1_6_0_sub_67_carry_3_), .B(
        npu_inst_pe_1_6_0_int_q_acc_3_), .ZN(npu_inst_pe_1_6_0_N68) );
  OR2_X1 npu_inst_pe_1_6_0_U124 ( .A1(npu_inst_pe_1_6_0_int_q_acc_3_), .A2(
        npu_inst_pe_1_6_0_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_6_0_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_6_0_U123 ( .A(npu_inst_pe_1_6_0_sub_67_carry_4_), .B(
        npu_inst_pe_1_6_0_int_q_acc_4_), .ZN(npu_inst_pe_1_6_0_N69) );
  OR2_X1 npu_inst_pe_1_6_0_U122 ( .A1(npu_inst_pe_1_6_0_int_q_acc_4_), .A2(
        npu_inst_pe_1_6_0_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_6_0_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_6_0_U121 ( .A(npu_inst_pe_1_6_0_sub_67_carry_5_), .B(
        npu_inst_pe_1_6_0_int_q_acc_5_), .ZN(npu_inst_pe_1_6_0_N70) );
  OR2_X1 npu_inst_pe_1_6_0_U120 ( .A1(npu_inst_pe_1_6_0_int_q_acc_5_), .A2(
        npu_inst_pe_1_6_0_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_6_0_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_6_0_U119 ( .A(npu_inst_pe_1_6_0_sub_67_carry_6_), .B(
        npu_inst_pe_1_6_0_int_q_acc_6_), .ZN(npu_inst_pe_1_6_0_N71) );
  OR2_X1 npu_inst_pe_1_6_0_U118 ( .A1(npu_inst_pe_1_6_0_int_q_acc_6_), .A2(
        npu_inst_pe_1_6_0_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_6_0_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_6_0_U117 ( .A(npu_inst_pe_1_6_0_int_q_acc_7_), .B(
        npu_inst_pe_1_6_0_sub_67_carry_7_), .ZN(npu_inst_pe_1_6_0_N72) );
  INV_X1 npu_inst_pe_1_6_0_U116 ( .A(npu_inst_n76), .ZN(npu_inst_pe_1_6_0_n7)
         );
  INV_X1 npu_inst_pe_1_6_0_U115 ( .A(npu_inst_pe_1_6_0_n7), .ZN(
        npu_inst_pe_1_6_0_n6) );
  INV_X1 npu_inst_pe_1_6_0_U114 ( .A(npu_inst_n54), .ZN(npu_inst_pe_1_6_0_n3)
         );
  AOI22_X1 npu_inst_pe_1_6_0_U113 ( .A1(npu_inst_int_data_y_7__0__0_), .A2(
        npu_inst_pe_1_6_0_n58), .B1(npu_inst_pe_1_6_0_n119), .B2(
        npu_inst_pe_1_6_0_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_6_0_n57) );
  INV_X1 npu_inst_pe_1_6_0_U112 ( .A(npu_inst_pe_1_6_0_n57), .ZN(
        npu_inst_pe_1_6_0_n108) );
  AOI22_X1 npu_inst_pe_1_6_0_U111 ( .A1(npu_inst_int_data_y_7__0__0_), .A2(
        npu_inst_pe_1_6_0_n54), .B1(npu_inst_pe_1_6_0_n118), .B2(
        npu_inst_pe_1_6_0_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_6_0_n53) );
  INV_X1 npu_inst_pe_1_6_0_U110 ( .A(npu_inst_pe_1_6_0_n53), .ZN(
        npu_inst_pe_1_6_0_n109) );
  AOI22_X1 npu_inst_pe_1_6_0_U107 ( .A1(npu_inst_int_data_y_7__0__0_), .A2(
        npu_inst_pe_1_6_0_n50), .B1(npu_inst_pe_1_6_0_n117), .B2(
        npu_inst_pe_1_6_0_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_6_0_n49) );
  INV_X1 npu_inst_pe_1_6_0_U106 ( .A(npu_inst_pe_1_6_0_n49), .ZN(
        npu_inst_pe_1_6_0_n110) );
  AOI22_X1 npu_inst_pe_1_6_0_U105 ( .A1(npu_inst_int_data_y_7__0__0_), .A2(
        npu_inst_pe_1_6_0_n46), .B1(npu_inst_pe_1_6_0_n116), .B2(
        npu_inst_pe_1_6_0_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_6_0_n45) );
  INV_X1 npu_inst_pe_1_6_0_U104 ( .A(npu_inst_pe_1_6_0_n45), .ZN(
        npu_inst_pe_1_6_0_n111) );
  AOI22_X1 npu_inst_pe_1_6_0_U103 ( .A1(npu_inst_int_data_y_7__0__0_), .A2(
        npu_inst_pe_1_6_0_n42), .B1(npu_inst_pe_1_6_0_n115), .B2(
        npu_inst_pe_1_6_0_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_6_0_n41) );
  INV_X1 npu_inst_pe_1_6_0_U102 ( .A(npu_inst_pe_1_6_0_n41), .ZN(
        npu_inst_pe_1_6_0_n112) );
  AOI22_X1 npu_inst_pe_1_6_0_U101 ( .A1(npu_inst_int_data_y_7__0__1_), .A2(
        npu_inst_pe_1_6_0_n58), .B1(npu_inst_pe_1_6_0_n119), .B2(
        npu_inst_pe_1_6_0_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_6_0_n59) );
  INV_X1 npu_inst_pe_1_6_0_U100 ( .A(npu_inst_pe_1_6_0_n59), .ZN(
        npu_inst_pe_1_6_0_n102) );
  AOI22_X1 npu_inst_pe_1_6_0_U99 ( .A1(npu_inst_int_data_y_7__0__1_), .A2(
        npu_inst_pe_1_6_0_n54), .B1(npu_inst_pe_1_6_0_n118), .B2(
        npu_inst_pe_1_6_0_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_6_0_n55) );
  INV_X1 npu_inst_pe_1_6_0_U98 ( .A(npu_inst_pe_1_6_0_n55), .ZN(
        npu_inst_pe_1_6_0_n103) );
  AOI22_X1 npu_inst_pe_1_6_0_U97 ( .A1(npu_inst_int_data_y_7__0__1_), .A2(
        npu_inst_pe_1_6_0_n50), .B1(npu_inst_pe_1_6_0_n117), .B2(
        npu_inst_pe_1_6_0_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_6_0_n51) );
  INV_X1 npu_inst_pe_1_6_0_U96 ( .A(npu_inst_pe_1_6_0_n51), .ZN(
        npu_inst_pe_1_6_0_n104) );
  AOI22_X1 npu_inst_pe_1_6_0_U95 ( .A1(npu_inst_int_data_y_7__0__1_), .A2(
        npu_inst_pe_1_6_0_n46), .B1(npu_inst_pe_1_6_0_n116), .B2(
        npu_inst_pe_1_6_0_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_6_0_n47) );
  INV_X1 npu_inst_pe_1_6_0_U94 ( .A(npu_inst_pe_1_6_0_n47), .ZN(
        npu_inst_pe_1_6_0_n105) );
  AOI22_X1 npu_inst_pe_1_6_0_U93 ( .A1(npu_inst_int_data_y_7__0__1_), .A2(
        npu_inst_pe_1_6_0_n42), .B1(npu_inst_pe_1_6_0_n115), .B2(
        npu_inst_pe_1_6_0_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_6_0_n43) );
  INV_X1 npu_inst_pe_1_6_0_U92 ( .A(npu_inst_pe_1_6_0_n43), .ZN(
        npu_inst_pe_1_6_0_n106) );
  AOI22_X1 npu_inst_pe_1_6_0_U91 ( .A1(npu_inst_pe_1_6_0_n38), .A2(
        npu_inst_int_data_y_7__0__1_), .B1(npu_inst_pe_1_6_0_n114), .B2(
        npu_inst_pe_1_6_0_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_6_0_n39) );
  INV_X1 npu_inst_pe_1_6_0_U90 ( .A(npu_inst_pe_1_6_0_n39), .ZN(
        npu_inst_pe_1_6_0_n107) );
  AOI22_X1 npu_inst_pe_1_6_0_U89 ( .A1(npu_inst_pe_1_6_0_n38), .A2(
        npu_inst_int_data_y_7__0__0_), .B1(npu_inst_pe_1_6_0_n114), .B2(
        npu_inst_pe_1_6_0_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_6_0_n37) );
  INV_X1 npu_inst_pe_1_6_0_U88 ( .A(npu_inst_pe_1_6_0_n37), .ZN(
        npu_inst_pe_1_6_0_n113) );
  NAND2_X1 npu_inst_pe_1_6_0_U87 ( .A1(npu_inst_pe_1_6_0_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_6_0_n60), .ZN(npu_inst_pe_1_6_0_n74) );
  OAI21_X1 npu_inst_pe_1_6_0_U86 ( .B1(npu_inst_pe_1_6_0_n63), .B2(
        npu_inst_pe_1_6_0_n60), .A(npu_inst_pe_1_6_0_n74), .ZN(
        npu_inst_pe_1_6_0_n97) );
  NAND2_X1 npu_inst_pe_1_6_0_U85 ( .A1(npu_inst_pe_1_6_0_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_6_0_n60), .ZN(npu_inst_pe_1_6_0_n73) );
  OAI21_X1 npu_inst_pe_1_6_0_U84 ( .B1(npu_inst_pe_1_6_0_n61), .B2(
        npu_inst_pe_1_6_0_n60), .A(npu_inst_pe_1_6_0_n73), .ZN(
        npu_inst_pe_1_6_0_n96) );
  NAND2_X1 npu_inst_pe_1_6_0_U83 ( .A1(npu_inst_pe_1_6_0_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_6_0_n56), .ZN(npu_inst_pe_1_6_0_n72) );
  OAI21_X1 npu_inst_pe_1_6_0_U82 ( .B1(npu_inst_pe_1_6_0_n63), .B2(
        npu_inst_pe_1_6_0_n56), .A(npu_inst_pe_1_6_0_n72), .ZN(
        npu_inst_pe_1_6_0_n95) );
  NAND2_X1 npu_inst_pe_1_6_0_U81 ( .A1(npu_inst_pe_1_6_0_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_6_0_n56), .ZN(npu_inst_pe_1_6_0_n71) );
  OAI21_X1 npu_inst_pe_1_6_0_U80 ( .B1(npu_inst_pe_1_6_0_n61), .B2(
        npu_inst_pe_1_6_0_n56), .A(npu_inst_pe_1_6_0_n71), .ZN(
        npu_inst_pe_1_6_0_n94) );
  NAND2_X1 npu_inst_pe_1_6_0_U79 ( .A1(npu_inst_pe_1_6_0_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_6_0_n52), .ZN(npu_inst_pe_1_6_0_n70) );
  OAI21_X1 npu_inst_pe_1_6_0_U78 ( .B1(npu_inst_pe_1_6_0_n63), .B2(
        npu_inst_pe_1_6_0_n52), .A(npu_inst_pe_1_6_0_n70), .ZN(
        npu_inst_pe_1_6_0_n93) );
  NAND2_X1 npu_inst_pe_1_6_0_U77 ( .A1(npu_inst_pe_1_6_0_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_6_0_n52), .ZN(npu_inst_pe_1_6_0_n69) );
  OAI21_X1 npu_inst_pe_1_6_0_U76 ( .B1(npu_inst_pe_1_6_0_n61), .B2(
        npu_inst_pe_1_6_0_n52), .A(npu_inst_pe_1_6_0_n69), .ZN(
        npu_inst_pe_1_6_0_n92) );
  NAND2_X1 npu_inst_pe_1_6_0_U75 ( .A1(npu_inst_pe_1_6_0_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_6_0_n48), .ZN(npu_inst_pe_1_6_0_n68) );
  OAI21_X1 npu_inst_pe_1_6_0_U74 ( .B1(npu_inst_pe_1_6_0_n63), .B2(
        npu_inst_pe_1_6_0_n48), .A(npu_inst_pe_1_6_0_n68), .ZN(
        npu_inst_pe_1_6_0_n91) );
  NAND2_X1 npu_inst_pe_1_6_0_U73 ( .A1(npu_inst_pe_1_6_0_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_6_0_n48), .ZN(npu_inst_pe_1_6_0_n67) );
  OAI21_X1 npu_inst_pe_1_6_0_U72 ( .B1(npu_inst_pe_1_6_0_n61), .B2(
        npu_inst_pe_1_6_0_n48), .A(npu_inst_pe_1_6_0_n67), .ZN(
        npu_inst_pe_1_6_0_n90) );
  NAND2_X1 npu_inst_pe_1_6_0_U71 ( .A1(npu_inst_pe_1_6_0_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_6_0_n44), .ZN(npu_inst_pe_1_6_0_n66) );
  OAI21_X1 npu_inst_pe_1_6_0_U70 ( .B1(npu_inst_pe_1_6_0_n63), .B2(
        npu_inst_pe_1_6_0_n44), .A(npu_inst_pe_1_6_0_n66), .ZN(
        npu_inst_pe_1_6_0_n89) );
  NAND2_X1 npu_inst_pe_1_6_0_U69 ( .A1(npu_inst_pe_1_6_0_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_6_0_n44), .ZN(npu_inst_pe_1_6_0_n65) );
  OAI21_X1 npu_inst_pe_1_6_0_U68 ( .B1(npu_inst_pe_1_6_0_n61), .B2(
        npu_inst_pe_1_6_0_n44), .A(npu_inst_pe_1_6_0_n65), .ZN(
        npu_inst_pe_1_6_0_n88) );
  NAND2_X1 npu_inst_pe_1_6_0_U67 ( .A1(npu_inst_pe_1_6_0_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_6_0_n40), .ZN(npu_inst_pe_1_6_0_n64) );
  OAI21_X1 npu_inst_pe_1_6_0_U66 ( .B1(npu_inst_pe_1_6_0_n63), .B2(
        npu_inst_pe_1_6_0_n40), .A(npu_inst_pe_1_6_0_n64), .ZN(
        npu_inst_pe_1_6_0_n87) );
  NAND2_X1 npu_inst_pe_1_6_0_U65 ( .A1(npu_inst_pe_1_6_0_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_6_0_n40), .ZN(npu_inst_pe_1_6_0_n62) );
  OAI21_X1 npu_inst_pe_1_6_0_U64 ( .B1(npu_inst_pe_1_6_0_n61), .B2(
        npu_inst_pe_1_6_0_n40), .A(npu_inst_pe_1_6_0_n62), .ZN(
        npu_inst_pe_1_6_0_n86) );
  AND2_X1 npu_inst_pe_1_6_0_U63 ( .A1(npu_inst_pe_1_6_0_N93), .A2(npu_inst_n54), .ZN(npu_inst_int_data_y_6__0__0_) );
  AND2_X1 npu_inst_pe_1_6_0_U62 ( .A1(npu_inst_n54), .A2(npu_inst_pe_1_6_0_N94), .ZN(npu_inst_int_data_y_6__0__1_) );
  NOR3_X1 npu_inst_pe_1_6_0_U61 ( .A1(npu_inst_pe_1_6_0_n26), .A2(npu_inst_n54), .A3(npu_inst_int_ckg[15]), .ZN(npu_inst_pe_1_6_0_n85) );
  OR2_X1 npu_inst_pe_1_6_0_U60 ( .A1(npu_inst_pe_1_6_0_n85), .A2(
        npu_inst_pe_1_6_0_n2), .ZN(npu_inst_pe_1_6_0_N84) );
  AND2_X1 npu_inst_pe_1_6_0_U59 ( .A1(npu_inst_pe_1_6_0_int_q_acc_0_), .A2(
        npu_inst_pe_1_6_0_n1), .ZN(npu_inst_int_data_res_6__0__0_) );
  AND2_X1 npu_inst_pe_1_6_0_U58 ( .A1(npu_inst_pe_1_6_0_n2), .A2(
        npu_inst_pe_1_6_0_int_q_acc_7_), .ZN(npu_inst_int_data_res_6__0__7_)
         );
  AND2_X1 npu_inst_pe_1_6_0_U57 ( .A1(npu_inst_pe_1_6_0_int_q_acc_1_), .A2(
        npu_inst_pe_1_6_0_n1), .ZN(npu_inst_int_data_res_6__0__1_) );
  AND2_X1 npu_inst_pe_1_6_0_U56 ( .A1(npu_inst_pe_1_6_0_int_q_acc_2_), .A2(
        npu_inst_pe_1_6_0_n1), .ZN(npu_inst_int_data_res_6__0__2_) );
  AND2_X1 npu_inst_pe_1_6_0_U55 ( .A1(npu_inst_pe_1_6_0_int_q_acc_3_), .A2(
        npu_inst_pe_1_6_0_n2), .ZN(npu_inst_int_data_res_6__0__3_) );
  AND2_X1 npu_inst_pe_1_6_0_U54 ( .A1(npu_inst_pe_1_6_0_int_q_acc_4_), .A2(
        npu_inst_pe_1_6_0_n2), .ZN(npu_inst_int_data_res_6__0__4_) );
  AND2_X1 npu_inst_pe_1_6_0_U53 ( .A1(npu_inst_pe_1_6_0_int_q_acc_5_), .A2(
        npu_inst_pe_1_6_0_n2), .ZN(npu_inst_int_data_res_6__0__5_) );
  AND2_X1 npu_inst_pe_1_6_0_U52 ( .A1(npu_inst_pe_1_6_0_int_q_acc_6_), .A2(
        npu_inst_pe_1_6_0_n2), .ZN(npu_inst_int_data_res_6__0__6_) );
  AOI222_X1 npu_inst_pe_1_6_0_U51 ( .A1(npu_inst_int_data_res_7__0__0_), .A2(
        npu_inst_pe_1_6_0_n1), .B1(npu_inst_pe_1_6_0_N73), .B2(
        npu_inst_pe_1_6_0_n76), .C1(npu_inst_pe_1_6_0_N65), .C2(
        npu_inst_pe_1_6_0_n77), .ZN(npu_inst_pe_1_6_0_n84) );
  INV_X1 npu_inst_pe_1_6_0_U50 ( .A(npu_inst_pe_1_6_0_n84), .ZN(
        npu_inst_pe_1_6_0_n101) );
  AOI222_X1 npu_inst_pe_1_6_0_U49 ( .A1(npu_inst_int_data_res_7__0__7_), .A2(
        npu_inst_pe_1_6_0_n1), .B1(npu_inst_pe_1_6_0_N80), .B2(
        npu_inst_pe_1_6_0_n76), .C1(npu_inst_pe_1_6_0_N72), .C2(
        npu_inst_pe_1_6_0_n77), .ZN(npu_inst_pe_1_6_0_n75) );
  INV_X1 npu_inst_pe_1_6_0_U48 ( .A(npu_inst_pe_1_6_0_n75), .ZN(
        npu_inst_pe_1_6_0_n33) );
  AOI222_X1 npu_inst_pe_1_6_0_U47 ( .A1(npu_inst_int_data_res_7__0__1_), .A2(
        npu_inst_pe_1_6_0_n1), .B1(npu_inst_pe_1_6_0_N74), .B2(
        npu_inst_pe_1_6_0_n76), .C1(npu_inst_pe_1_6_0_N66), .C2(
        npu_inst_pe_1_6_0_n77), .ZN(npu_inst_pe_1_6_0_n83) );
  INV_X1 npu_inst_pe_1_6_0_U46 ( .A(npu_inst_pe_1_6_0_n83), .ZN(
        npu_inst_pe_1_6_0_n100) );
  AOI222_X1 npu_inst_pe_1_6_0_U45 ( .A1(npu_inst_int_data_res_7__0__2_), .A2(
        npu_inst_pe_1_6_0_n1), .B1(npu_inst_pe_1_6_0_N75), .B2(
        npu_inst_pe_1_6_0_n76), .C1(npu_inst_pe_1_6_0_N67), .C2(
        npu_inst_pe_1_6_0_n77), .ZN(npu_inst_pe_1_6_0_n82) );
  INV_X1 npu_inst_pe_1_6_0_U44 ( .A(npu_inst_pe_1_6_0_n82), .ZN(
        npu_inst_pe_1_6_0_n99) );
  AOI222_X1 npu_inst_pe_1_6_0_U43 ( .A1(npu_inst_int_data_res_7__0__3_), .A2(
        npu_inst_pe_1_6_0_n1), .B1(npu_inst_pe_1_6_0_N76), .B2(
        npu_inst_pe_1_6_0_n76), .C1(npu_inst_pe_1_6_0_N68), .C2(
        npu_inst_pe_1_6_0_n77), .ZN(npu_inst_pe_1_6_0_n81) );
  INV_X1 npu_inst_pe_1_6_0_U42 ( .A(npu_inst_pe_1_6_0_n81), .ZN(
        npu_inst_pe_1_6_0_n98) );
  AOI222_X1 npu_inst_pe_1_6_0_U41 ( .A1(npu_inst_int_data_res_7__0__4_), .A2(
        npu_inst_pe_1_6_0_n1), .B1(npu_inst_pe_1_6_0_N77), .B2(
        npu_inst_pe_1_6_0_n76), .C1(npu_inst_pe_1_6_0_N69), .C2(
        npu_inst_pe_1_6_0_n77), .ZN(npu_inst_pe_1_6_0_n80) );
  INV_X1 npu_inst_pe_1_6_0_U40 ( .A(npu_inst_pe_1_6_0_n80), .ZN(
        npu_inst_pe_1_6_0_n36) );
  AOI222_X1 npu_inst_pe_1_6_0_U39 ( .A1(npu_inst_int_data_res_7__0__5_), .A2(
        npu_inst_pe_1_6_0_n1), .B1(npu_inst_pe_1_6_0_N78), .B2(
        npu_inst_pe_1_6_0_n76), .C1(npu_inst_pe_1_6_0_N70), .C2(
        npu_inst_pe_1_6_0_n77), .ZN(npu_inst_pe_1_6_0_n79) );
  INV_X1 npu_inst_pe_1_6_0_U38 ( .A(npu_inst_pe_1_6_0_n79), .ZN(
        npu_inst_pe_1_6_0_n35) );
  AOI222_X1 npu_inst_pe_1_6_0_U37 ( .A1(npu_inst_int_data_res_7__0__6_), .A2(
        npu_inst_pe_1_6_0_n1), .B1(npu_inst_pe_1_6_0_N79), .B2(
        npu_inst_pe_1_6_0_n76), .C1(npu_inst_pe_1_6_0_N71), .C2(
        npu_inst_pe_1_6_0_n77), .ZN(npu_inst_pe_1_6_0_n78) );
  INV_X1 npu_inst_pe_1_6_0_U36 ( .A(npu_inst_pe_1_6_0_n78), .ZN(
        npu_inst_pe_1_6_0_n34) );
  AND2_X1 npu_inst_pe_1_6_0_U35 ( .A1(npu_inst_pe_1_6_0_o_data_h_1_), .A2(
        npu_inst_pe_1_6_0_int_q_weight_1_), .ZN(npu_inst_pe_1_6_0_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_6_0_U34 ( .A1(npu_inst_pe_1_6_0_o_data_h_0_), .A2(
        npu_inst_pe_1_6_0_int_q_weight_1_), .ZN(npu_inst_pe_1_6_0_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_6_0_U33 ( .A(npu_inst_pe_1_6_0_int_data_1_), .ZN(
        npu_inst_pe_1_6_0_n14) );
  AOI22_X1 npu_inst_pe_1_6_0_U32 ( .A1(npu_inst_n54), .A2(
        npu_inst_int_data_y_7__0__1_), .B1(npu_inst_pe_1_6_0_n3), .B2(
        npu_inst_int_data_x_6__1__1_), .ZN(npu_inst_pe_1_6_0_n63) );
  AOI22_X1 npu_inst_pe_1_6_0_U31 ( .A1(npu_inst_n54), .A2(
        npu_inst_int_data_y_7__0__0_), .B1(npu_inst_pe_1_6_0_n3), .B2(
        npu_inst_int_data_x_6__1__0_), .ZN(npu_inst_pe_1_6_0_n61) );
  INV_X1 npu_inst_pe_1_6_0_U30 ( .A(npu_inst_pe_1_6_0_int_data_0_), .ZN(
        npu_inst_pe_1_6_0_n13) );
  INV_X1 npu_inst_pe_1_6_0_U29 ( .A(npu_inst_n68), .ZN(npu_inst_pe_1_6_0_n5)
         );
  OR3_X1 npu_inst_pe_1_6_0_U28 ( .A1(npu_inst_pe_1_6_0_n6), .A2(
        npu_inst_pe_1_6_0_n8), .A3(npu_inst_pe_1_6_0_n5), .ZN(
        npu_inst_pe_1_6_0_n56) );
  OR3_X1 npu_inst_pe_1_6_0_U27 ( .A1(npu_inst_pe_1_6_0_n5), .A2(
        npu_inst_pe_1_6_0_n8), .A3(npu_inst_pe_1_6_0_n7), .ZN(
        npu_inst_pe_1_6_0_n48) );
  INV_X1 npu_inst_pe_1_6_0_U26 ( .A(npu_inst_pe_1_6_0_n5), .ZN(
        npu_inst_pe_1_6_0_n4) );
  OR3_X1 npu_inst_pe_1_6_0_U25 ( .A1(npu_inst_pe_1_6_0_n4), .A2(
        npu_inst_pe_1_6_0_n8), .A3(npu_inst_pe_1_6_0_n7), .ZN(
        npu_inst_pe_1_6_0_n52) );
  OR3_X1 npu_inst_pe_1_6_0_U24 ( .A1(npu_inst_pe_1_6_0_n6), .A2(
        npu_inst_pe_1_6_0_n8), .A3(npu_inst_pe_1_6_0_n4), .ZN(
        npu_inst_pe_1_6_0_n60) );
  NOR2_X1 npu_inst_pe_1_6_0_U23 ( .A1(npu_inst_pe_1_6_0_n60), .A2(
        npu_inst_pe_1_6_0_n3), .ZN(npu_inst_pe_1_6_0_n58) );
  NOR2_X1 npu_inst_pe_1_6_0_U22 ( .A1(npu_inst_pe_1_6_0_n56), .A2(
        npu_inst_pe_1_6_0_n3), .ZN(npu_inst_pe_1_6_0_n54) );
  NOR2_X1 npu_inst_pe_1_6_0_U21 ( .A1(npu_inst_pe_1_6_0_n52), .A2(
        npu_inst_pe_1_6_0_n3), .ZN(npu_inst_pe_1_6_0_n50) );
  NOR2_X1 npu_inst_pe_1_6_0_U20 ( .A1(npu_inst_pe_1_6_0_n48), .A2(
        npu_inst_pe_1_6_0_n3), .ZN(npu_inst_pe_1_6_0_n46) );
  NOR2_X1 npu_inst_pe_1_6_0_U19 ( .A1(npu_inst_pe_1_6_0_n40), .A2(
        npu_inst_pe_1_6_0_n3), .ZN(npu_inst_pe_1_6_0_n38) );
  NOR2_X1 npu_inst_pe_1_6_0_U18 ( .A1(npu_inst_pe_1_6_0_n44), .A2(
        npu_inst_pe_1_6_0_n3), .ZN(npu_inst_pe_1_6_0_n42) );
  BUF_X1 npu_inst_pe_1_6_0_U17 ( .A(npu_inst_n95), .Z(npu_inst_pe_1_6_0_n8) );
  INV_X1 npu_inst_pe_1_6_0_U16 ( .A(npu_inst_n123), .ZN(npu_inst_pe_1_6_0_n12)
         );
  INV_X1 npu_inst_pe_1_6_0_U15 ( .A(npu_inst_pe_1_6_0_n38), .ZN(
        npu_inst_pe_1_6_0_n114) );
  INV_X1 npu_inst_pe_1_6_0_U14 ( .A(npu_inst_pe_1_6_0_n58), .ZN(
        npu_inst_pe_1_6_0_n119) );
  INV_X1 npu_inst_pe_1_6_0_U13 ( .A(npu_inst_pe_1_6_0_n54), .ZN(
        npu_inst_pe_1_6_0_n118) );
  INV_X1 npu_inst_pe_1_6_0_U12 ( .A(npu_inst_pe_1_6_0_n50), .ZN(
        npu_inst_pe_1_6_0_n117) );
  INV_X1 npu_inst_pe_1_6_0_U11 ( .A(npu_inst_pe_1_6_0_n46), .ZN(
        npu_inst_pe_1_6_0_n116) );
  INV_X1 npu_inst_pe_1_6_0_U10 ( .A(npu_inst_pe_1_6_0_n42), .ZN(
        npu_inst_pe_1_6_0_n115) );
  BUF_X1 npu_inst_pe_1_6_0_U9 ( .A(npu_inst_n14), .Z(npu_inst_pe_1_6_0_n2) );
  BUF_X1 npu_inst_pe_1_6_0_U8 ( .A(npu_inst_n14), .Z(npu_inst_pe_1_6_0_n1) );
  BUF_X1 npu_inst_pe_1_6_0_U7 ( .A(npu_inst_pe_1_6_0_n12), .Z(
        npu_inst_pe_1_6_0_n11) );
  BUF_X1 npu_inst_pe_1_6_0_U6 ( .A(npu_inst_pe_1_6_0_n12), .Z(
        npu_inst_pe_1_6_0_n10) );
  BUF_X1 npu_inst_pe_1_6_0_U5 ( .A(npu_inst_pe_1_6_0_n12), .Z(
        npu_inst_pe_1_6_0_n9) );
  NOR2_X1 npu_inst_pe_1_6_0_U4 ( .A1(npu_inst_pe_1_6_0_int_q_weight_0_), .A2(
        npu_inst_pe_1_6_0_n1), .ZN(npu_inst_pe_1_6_0_n76) );
  NOR2_X1 npu_inst_pe_1_6_0_U3 ( .A1(npu_inst_pe_1_6_0_n27), .A2(
        npu_inst_pe_1_6_0_n1), .ZN(npu_inst_pe_1_6_0_n77) );
  FA_X1 npu_inst_pe_1_6_0_sub_67_U2_1 ( .A(npu_inst_pe_1_6_0_int_q_acc_1_), 
        .B(npu_inst_pe_1_6_0_n14), .CI(npu_inst_pe_1_6_0_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_6_0_sub_67_carry_2_), .S(npu_inst_pe_1_6_0_N66) );
  FA_X1 npu_inst_pe_1_6_0_add_69_U1_1 ( .A(npu_inst_pe_1_6_0_int_q_acc_1_), 
        .B(npu_inst_pe_1_6_0_int_data_1_), .CI(
        npu_inst_pe_1_6_0_add_69_carry_1_), .CO(
        npu_inst_pe_1_6_0_add_69_carry_2_), .S(npu_inst_pe_1_6_0_N74) );
  NAND3_X1 npu_inst_pe_1_6_0_U109 ( .A1(npu_inst_pe_1_6_0_n5), .A2(
        npu_inst_pe_1_6_0_n7), .A3(npu_inst_pe_1_6_0_n8), .ZN(
        npu_inst_pe_1_6_0_n44) );
  NAND3_X1 npu_inst_pe_1_6_0_U108 ( .A1(npu_inst_pe_1_6_0_n4), .A2(
        npu_inst_pe_1_6_0_n7), .A3(npu_inst_pe_1_6_0_n8), .ZN(
        npu_inst_pe_1_6_0_n40) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_6_0_n34), .CK(
        npu_inst_pe_1_6_0_net3458), .RN(npu_inst_pe_1_6_0_n9), .Q(
        npu_inst_pe_1_6_0_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_6_0_n35), .CK(
        npu_inst_pe_1_6_0_net3458), .RN(npu_inst_pe_1_6_0_n9), .Q(
        npu_inst_pe_1_6_0_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_6_0_n36), .CK(
        npu_inst_pe_1_6_0_net3458), .RN(npu_inst_pe_1_6_0_n9), .Q(
        npu_inst_pe_1_6_0_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_6_0_n98), .CK(
        npu_inst_pe_1_6_0_net3458), .RN(npu_inst_pe_1_6_0_n9), .Q(
        npu_inst_pe_1_6_0_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_6_0_n99), .CK(
        npu_inst_pe_1_6_0_net3458), .RN(npu_inst_pe_1_6_0_n9), .Q(
        npu_inst_pe_1_6_0_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_6_0_n100), 
        .CK(npu_inst_pe_1_6_0_net3458), .RN(npu_inst_pe_1_6_0_n9), .Q(
        npu_inst_pe_1_6_0_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_6_0_n33), .CK(
        npu_inst_pe_1_6_0_net3458), .RN(npu_inst_pe_1_6_0_n9), .Q(
        npu_inst_pe_1_6_0_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_6_0_n101), 
        .CK(npu_inst_pe_1_6_0_net3458), .RN(npu_inst_pe_1_6_0_n9), .Q(
        npu_inst_pe_1_6_0_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_weight_reg_0_ ( .D(npu_inst_n109), .CK(
        npu_inst_pe_1_6_0_net3464), .RN(npu_inst_pe_1_6_0_n9), .Q(
        npu_inst_pe_1_6_0_int_q_weight_0_), .QN(npu_inst_pe_1_6_0_n27) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_weight_reg_1_ ( .D(npu_inst_n115), .CK(
        npu_inst_pe_1_6_0_net3464), .RN(npu_inst_pe_1_6_0_n9), .Q(
        npu_inst_pe_1_6_0_int_q_weight_1_), .QN(npu_inst_pe_1_6_0_n26) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_6_0_n113), 
        .CK(npu_inst_pe_1_6_0_net3464), .RN(npu_inst_pe_1_6_0_n9), .Q(
        npu_inst_pe_1_6_0_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_6_0_n107), 
        .CK(npu_inst_pe_1_6_0_net3464), .RN(npu_inst_pe_1_6_0_n9), .Q(
        npu_inst_pe_1_6_0_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_6_0_n112), 
        .CK(npu_inst_pe_1_6_0_net3464), .RN(npu_inst_pe_1_6_0_n10), .Q(
        npu_inst_pe_1_6_0_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_6_0_n106), 
        .CK(npu_inst_pe_1_6_0_net3464), .RN(npu_inst_pe_1_6_0_n10), .Q(
        npu_inst_pe_1_6_0_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_6_0_n111), 
        .CK(npu_inst_pe_1_6_0_net3464), .RN(npu_inst_pe_1_6_0_n10), .Q(
        npu_inst_pe_1_6_0_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_6_0_n105), 
        .CK(npu_inst_pe_1_6_0_net3464), .RN(npu_inst_pe_1_6_0_n10), .Q(
        npu_inst_pe_1_6_0_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_6_0_n110), 
        .CK(npu_inst_pe_1_6_0_net3464), .RN(npu_inst_pe_1_6_0_n10), .Q(
        npu_inst_pe_1_6_0_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_6_0_n104), 
        .CK(npu_inst_pe_1_6_0_net3464), .RN(npu_inst_pe_1_6_0_n10), .Q(
        npu_inst_pe_1_6_0_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_6_0_n109), 
        .CK(npu_inst_pe_1_6_0_net3464), .RN(npu_inst_pe_1_6_0_n10), .Q(
        npu_inst_pe_1_6_0_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_6_0_n103), 
        .CK(npu_inst_pe_1_6_0_net3464), .RN(npu_inst_pe_1_6_0_n10), .Q(
        npu_inst_pe_1_6_0_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_6_0_n108), 
        .CK(npu_inst_pe_1_6_0_net3464), .RN(npu_inst_pe_1_6_0_n10), .Q(
        npu_inst_pe_1_6_0_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_6_0_n102), 
        .CK(npu_inst_pe_1_6_0_net3464), .RN(npu_inst_pe_1_6_0_n10), .Q(
        npu_inst_pe_1_6_0_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_6_0_n86), 
        .CK(npu_inst_pe_1_6_0_net3464), .RN(npu_inst_pe_1_6_0_n10), .Q(
        npu_inst_pe_1_6_0_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_6_0_n87), 
        .CK(npu_inst_pe_1_6_0_net3464), .RN(npu_inst_pe_1_6_0_n10), .Q(
        npu_inst_pe_1_6_0_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_6_0_n88), 
        .CK(npu_inst_pe_1_6_0_net3464), .RN(npu_inst_pe_1_6_0_n11), .Q(
        npu_inst_pe_1_6_0_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_6_0_n89), 
        .CK(npu_inst_pe_1_6_0_net3464), .RN(npu_inst_pe_1_6_0_n11), .Q(
        npu_inst_pe_1_6_0_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_6_0_n90), 
        .CK(npu_inst_pe_1_6_0_net3464), .RN(npu_inst_pe_1_6_0_n11), .Q(
        npu_inst_pe_1_6_0_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_6_0_n91), 
        .CK(npu_inst_pe_1_6_0_net3464), .RN(npu_inst_pe_1_6_0_n11), .Q(
        npu_inst_pe_1_6_0_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_6_0_n92), 
        .CK(npu_inst_pe_1_6_0_net3464), .RN(npu_inst_pe_1_6_0_n11), .Q(
        npu_inst_pe_1_6_0_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_6_0_n93), 
        .CK(npu_inst_pe_1_6_0_net3464), .RN(npu_inst_pe_1_6_0_n11), .Q(
        npu_inst_pe_1_6_0_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_6_0_n94), 
        .CK(npu_inst_pe_1_6_0_net3464), .RN(npu_inst_pe_1_6_0_n11), .Q(
        npu_inst_pe_1_6_0_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_6_0_n95), 
        .CK(npu_inst_pe_1_6_0_net3464), .RN(npu_inst_pe_1_6_0_n11), .Q(
        npu_inst_pe_1_6_0_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_6_0_n96), 
        .CK(npu_inst_pe_1_6_0_net3464), .RN(npu_inst_pe_1_6_0_n11), .Q(
        npu_inst_pe_1_6_0_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_6_0_n97), 
        .CK(npu_inst_pe_1_6_0_net3464), .RN(npu_inst_pe_1_6_0_n11), .Q(
        npu_inst_pe_1_6_0_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_6_0_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_6_0_N84), .SE(1'b0), .GCK(npu_inst_pe_1_6_0_net3458) );
  CLKGATETST_X1 npu_inst_pe_1_6_0_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n62), .SE(1'b0), .GCK(npu_inst_pe_1_6_0_net3464) );
  MUX2_X1 npu_inst_pe_1_6_1_U162 ( .A(npu_inst_pe_1_6_1_n32), .B(
        npu_inst_pe_1_6_1_n29), .S(npu_inst_pe_1_6_1_n8), .Z(
        npu_inst_pe_1_6_1_N93) );
  MUX2_X1 npu_inst_pe_1_6_1_U161 ( .A(npu_inst_pe_1_6_1_n31), .B(
        npu_inst_pe_1_6_1_n30), .S(npu_inst_pe_1_6_1_n6), .Z(
        npu_inst_pe_1_6_1_n32) );
  MUX2_X1 npu_inst_pe_1_6_1_U160 ( .A(npu_inst_pe_1_6_1_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_6_1_int_q_reg_v_1__0_), .S(npu_inst_pe_1_6_1_n4), .Z(
        npu_inst_pe_1_6_1_n31) );
  MUX2_X1 npu_inst_pe_1_6_1_U159 ( .A(npu_inst_pe_1_6_1_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_6_1_int_q_reg_v_3__0_), .S(npu_inst_pe_1_6_1_n4), .Z(
        npu_inst_pe_1_6_1_n30) );
  MUX2_X1 npu_inst_pe_1_6_1_U158 ( .A(npu_inst_pe_1_6_1_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_6_1_int_q_reg_v_5__0_), .S(npu_inst_pe_1_6_1_n4), .Z(
        npu_inst_pe_1_6_1_n29) );
  MUX2_X1 npu_inst_pe_1_6_1_U157 ( .A(npu_inst_pe_1_6_1_n28), .B(
        npu_inst_pe_1_6_1_n23), .S(npu_inst_pe_1_6_1_n8), .Z(
        npu_inst_pe_1_6_1_N94) );
  MUX2_X1 npu_inst_pe_1_6_1_U156 ( .A(npu_inst_pe_1_6_1_n25), .B(
        npu_inst_pe_1_6_1_n24), .S(npu_inst_pe_1_6_1_n6), .Z(
        npu_inst_pe_1_6_1_n28) );
  MUX2_X1 npu_inst_pe_1_6_1_U155 ( .A(npu_inst_pe_1_6_1_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_6_1_int_q_reg_v_1__1_), .S(npu_inst_pe_1_6_1_n4), .Z(
        npu_inst_pe_1_6_1_n25) );
  MUX2_X1 npu_inst_pe_1_6_1_U154 ( .A(npu_inst_pe_1_6_1_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_6_1_int_q_reg_v_3__1_), .S(npu_inst_pe_1_6_1_n4), .Z(
        npu_inst_pe_1_6_1_n24) );
  MUX2_X1 npu_inst_pe_1_6_1_U153 ( .A(npu_inst_pe_1_6_1_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_6_1_int_q_reg_v_5__1_), .S(npu_inst_pe_1_6_1_n4), .Z(
        npu_inst_pe_1_6_1_n23) );
  MUX2_X1 npu_inst_pe_1_6_1_U152 ( .A(npu_inst_pe_1_6_1_n22), .B(
        npu_inst_pe_1_6_1_n19), .S(npu_inst_pe_1_6_1_n8), .Z(
        npu_inst_int_data_x_6__1__1_) );
  MUX2_X1 npu_inst_pe_1_6_1_U151 ( .A(npu_inst_pe_1_6_1_n21), .B(
        npu_inst_pe_1_6_1_n20), .S(npu_inst_pe_1_6_1_n6), .Z(
        npu_inst_pe_1_6_1_n22) );
  MUX2_X1 npu_inst_pe_1_6_1_U150 ( .A(npu_inst_pe_1_6_1_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_6_1_int_q_reg_h_1__1_), .S(npu_inst_pe_1_6_1_n4), .Z(
        npu_inst_pe_1_6_1_n21) );
  MUX2_X1 npu_inst_pe_1_6_1_U149 ( .A(npu_inst_pe_1_6_1_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_6_1_int_q_reg_h_3__1_), .S(npu_inst_pe_1_6_1_n4), .Z(
        npu_inst_pe_1_6_1_n20) );
  MUX2_X1 npu_inst_pe_1_6_1_U148 ( .A(npu_inst_pe_1_6_1_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_6_1_int_q_reg_h_5__1_), .S(npu_inst_pe_1_6_1_n4), .Z(
        npu_inst_pe_1_6_1_n19) );
  MUX2_X1 npu_inst_pe_1_6_1_U147 ( .A(npu_inst_pe_1_6_1_n18), .B(
        npu_inst_pe_1_6_1_n15), .S(npu_inst_pe_1_6_1_n8), .Z(
        npu_inst_int_data_x_6__1__0_) );
  MUX2_X1 npu_inst_pe_1_6_1_U146 ( .A(npu_inst_pe_1_6_1_n17), .B(
        npu_inst_pe_1_6_1_n16), .S(npu_inst_pe_1_6_1_n6), .Z(
        npu_inst_pe_1_6_1_n18) );
  MUX2_X1 npu_inst_pe_1_6_1_U145 ( .A(npu_inst_pe_1_6_1_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_6_1_int_q_reg_h_1__0_), .S(npu_inst_pe_1_6_1_n4), .Z(
        npu_inst_pe_1_6_1_n17) );
  MUX2_X1 npu_inst_pe_1_6_1_U144 ( .A(npu_inst_pe_1_6_1_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_6_1_int_q_reg_h_3__0_), .S(npu_inst_pe_1_6_1_n4), .Z(
        npu_inst_pe_1_6_1_n16) );
  MUX2_X1 npu_inst_pe_1_6_1_U143 ( .A(npu_inst_pe_1_6_1_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_6_1_int_q_reg_h_5__0_), .S(npu_inst_pe_1_6_1_n4), .Z(
        npu_inst_pe_1_6_1_n15) );
  XOR2_X1 npu_inst_pe_1_6_1_U142 ( .A(npu_inst_pe_1_6_1_int_data_0_), .B(
        npu_inst_pe_1_6_1_int_q_acc_0_), .Z(npu_inst_pe_1_6_1_N73) );
  AND2_X1 npu_inst_pe_1_6_1_U141 ( .A1(npu_inst_pe_1_6_1_int_q_acc_0_), .A2(
        npu_inst_pe_1_6_1_int_data_0_), .ZN(npu_inst_pe_1_6_1_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_6_1_U140 ( .A(npu_inst_pe_1_6_1_int_q_acc_0_), .B(
        npu_inst_pe_1_6_1_n13), .ZN(npu_inst_pe_1_6_1_N65) );
  OR2_X1 npu_inst_pe_1_6_1_U139 ( .A1(npu_inst_pe_1_6_1_n13), .A2(
        npu_inst_pe_1_6_1_int_q_acc_0_), .ZN(npu_inst_pe_1_6_1_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_6_1_U138 ( .A(npu_inst_pe_1_6_1_int_q_acc_2_), .B(
        npu_inst_pe_1_6_1_add_69_carry_2_), .Z(npu_inst_pe_1_6_1_N75) );
  AND2_X1 npu_inst_pe_1_6_1_U137 ( .A1(npu_inst_pe_1_6_1_add_69_carry_2_), 
        .A2(npu_inst_pe_1_6_1_int_q_acc_2_), .ZN(
        npu_inst_pe_1_6_1_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_6_1_U136 ( .A(npu_inst_pe_1_6_1_int_q_acc_3_), .B(
        npu_inst_pe_1_6_1_add_69_carry_3_), .Z(npu_inst_pe_1_6_1_N76) );
  AND2_X1 npu_inst_pe_1_6_1_U135 ( .A1(npu_inst_pe_1_6_1_add_69_carry_3_), 
        .A2(npu_inst_pe_1_6_1_int_q_acc_3_), .ZN(
        npu_inst_pe_1_6_1_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_6_1_U134 ( .A(npu_inst_pe_1_6_1_int_q_acc_4_), .B(
        npu_inst_pe_1_6_1_add_69_carry_4_), .Z(npu_inst_pe_1_6_1_N77) );
  AND2_X1 npu_inst_pe_1_6_1_U133 ( .A1(npu_inst_pe_1_6_1_add_69_carry_4_), 
        .A2(npu_inst_pe_1_6_1_int_q_acc_4_), .ZN(
        npu_inst_pe_1_6_1_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_6_1_U132 ( .A(npu_inst_pe_1_6_1_int_q_acc_5_), .B(
        npu_inst_pe_1_6_1_add_69_carry_5_), .Z(npu_inst_pe_1_6_1_N78) );
  AND2_X1 npu_inst_pe_1_6_1_U131 ( .A1(npu_inst_pe_1_6_1_add_69_carry_5_), 
        .A2(npu_inst_pe_1_6_1_int_q_acc_5_), .ZN(
        npu_inst_pe_1_6_1_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_6_1_U130 ( .A(npu_inst_pe_1_6_1_int_q_acc_6_), .B(
        npu_inst_pe_1_6_1_add_69_carry_6_), .Z(npu_inst_pe_1_6_1_N79) );
  AND2_X1 npu_inst_pe_1_6_1_U129 ( .A1(npu_inst_pe_1_6_1_add_69_carry_6_), 
        .A2(npu_inst_pe_1_6_1_int_q_acc_6_), .ZN(
        npu_inst_pe_1_6_1_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_6_1_U128 ( .A(npu_inst_pe_1_6_1_int_q_acc_7_), .B(
        npu_inst_pe_1_6_1_add_69_carry_7_), .Z(npu_inst_pe_1_6_1_N80) );
  XNOR2_X1 npu_inst_pe_1_6_1_U127 ( .A(npu_inst_pe_1_6_1_sub_67_carry_2_), .B(
        npu_inst_pe_1_6_1_int_q_acc_2_), .ZN(npu_inst_pe_1_6_1_N67) );
  OR2_X1 npu_inst_pe_1_6_1_U126 ( .A1(npu_inst_pe_1_6_1_int_q_acc_2_), .A2(
        npu_inst_pe_1_6_1_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_6_1_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_6_1_U125 ( .A(npu_inst_pe_1_6_1_sub_67_carry_3_), .B(
        npu_inst_pe_1_6_1_int_q_acc_3_), .ZN(npu_inst_pe_1_6_1_N68) );
  OR2_X1 npu_inst_pe_1_6_1_U124 ( .A1(npu_inst_pe_1_6_1_int_q_acc_3_), .A2(
        npu_inst_pe_1_6_1_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_6_1_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_6_1_U123 ( .A(npu_inst_pe_1_6_1_sub_67_carry_4_), .B(
        npu_inst_pe_1_6_1_int_q_acc_4_), .ZN(npu_inst_pe_1_6_1_N69) );
  OR2_X1 npu_inst_pe_1_6_1_U122 ( .A1(npu_inst_pe_1_6_1_int_q_acc_4_), .A2(
        npu_inst_pe_1_6_1_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_6_1_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_6_1_U121 ( .A(npu_inst_pe_1_6_1_sub_67_carry_5_), .B(
        npu_inst_pe_1_6_1_int_q_acc_5_), .ZN(npu_inst_pe_1_6_1_N70) );
  OR2_X1 npu_inst_pe_1_6_1_U120 ( .A1(npu_inst_pe_1_6_1_int_q_acc_5_), .A2(
        npu_inst_pe_1_6_1_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_6_1_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_6_1_U119 ( .A(npu_inst_pe_1_6_1_sub_67_carry_6_), .B(
        npu_inst_pe_1_6_1_int_q_acc_6_), .ZN(npu_inst_pe_1_6_1_N71) );
  OR2_X1 npu_inst_pe_1_6_1_U118 ( .A1(npu_inst_pe_1_6_1_int_q_acc_6_), .A2(
        npu_inst_pe_1_6_1_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_6_1_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_6_1_U117 ( .A(npu_inst_pe_1_6_1_int_q_acc_7_), .B(
        npu_inst_pe_1_6_1_sub_67_carry_7_), .ZN(npu_inst_pe_1_6_1_N72) );
  INV_X1 npu_inst_pe_1_6_1_U116 ( .A(npu_inst_n76), .ZN(npu_inst_pe_1_6_1_n7)
         );
  INV_X1 npu_inst_pe_1_6_1_U115 ( .A(npu_inst_pe_1_6_1_n7), .ZN(
        npu_inst_pe_1_6_1_n6) );
  INV_X1 npu_inst_pe_1_6_1_U114 ( .A(npu_inst_n54), .ZN(npu_inst_pe_1_6_1_n3)
         );
  AOI22_X1 npu_inst_pe_1_6_1_U113 ( .A1(npu_inst_int_data_y_7__1__0_), .A2(
        npu_inst_pe_1_6_1_n58), .B1(npu_inst_pe_1_6_1_n119), .B2(
        npu_inst_pe_1_6_1_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_6_1_n57) );
  INV_X1 npu_inst_pe_1_6_1_U112 ( .A(npu_inst_pe_1_6_1_n57), .ZN(
        npu_inst_pe_1_6_1_n108) );
  AOI22_X1 npu_inst_pe_1_6_1_U111 ( .A1(npu_inst_int_data_y_7__1__0_), .A2(
        npu_inst_pe_1_6_1_n54), .B1(npu_inst_pe_1_6_1_n118), .B2(
        npu_inst_pe_1_6_1_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_6_1_n53) );
  INV_X1 npu_inst_pe_1_6_1_U110 ( .A(npu_inst_pe_1_6_1_n53), .ZN(
        npu_inst_pe_1_6_1_n109) );
  AOI22_X1 npu_inst_pe_1_6_1_U107 ( .A1(npu_inst_int_data_y_7__1__0_), .A2(
        npu_inst_pe_1_6_1_n50), .B1(npu_inst_pe_1_6_1_n117), .B2(
        npu_inst_pe_1_6_1_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_6_1_n49) );
  INV_X1 npu_inst_pe_1_6_1_U106 ( .A(npu_inst_pe_1_6_1_n49), .ZN(
        npu_inst_pe_1_6_1_n110) );
  AOI22_X1 npu_inst_pe_1_6_1_U105 ( .A1(npu_inst_int_data_y_7__1__0_), .A2(
        npu_inst_pe_1_6_1_n46), .B1(npu_inst_pe_1_6_1_n116), .B2(
        npu_inst_pe_1_6_1_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_6_1_n45) );
  INV_X1 npu_inst_pe_1_6_1_U104 ( .A(npu_inst_pe_1_6_1_n45), .ZN(
        npu_inst_pe_1_6_1_n111) );
  AOI22_X1 npu_inst_pe_1_6_1_U103 ( .A1(npu_inst_int_data_y_7__1__0_), .A2(
        npu_inst_pe_1_6_1_n42), .B1(npu_inst_pe_1_6_1_n115), .B2(
        npu_inst_pe_1_6_1_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_6_1_n41) );
  INV_X1 npu_inst_pe_1_6_1_U102 ( .A(npu_inst_pe_1_6_1_n41), .ZN(
        npu_inst_pe_1_6_1_n112) );
  AOI22_X1 npu_inst_pe_1_6_1_U101 ( .A1(npu_inst_int_data_y_7__1__1_), .A2(
        npu_inst_pe_1_6_1_n58), .B1(npu_inst_pe_1_6_1_n119), .B2(
        npu_inst_pe_1_6_1_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_6_1_n59) );
  INV_X1 npu_inst_pe_1_6_1_U100 ( .A(npu_inst_pe_1_6_1_n59), .ZN(
        npu_inst_pe_1_6_1_n102) );
  AOI22_X1 npu_inst_pe_1_6_1_U99 ( .A1(npu_inst_int_data_y_7__1__1_), .A2(
        npu_inst_pe_1_6_1_n54), .B1(npu_inst_pe_1_6_1_n118), .B2(
        npu_inst_pe_1_6_1_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_6_1_n55) );
  INV_X1 npu_inst_pe_1_6_1_U98 ( .A(npu_inst_pe_1_6_1_n55), .ZN(
        npu_inst_pe_1_6_1_n103) );
  AOI22_X1 npu_inst_pe_1_6_1_U97 ( .A1(npu_inst_int_data_y_7__1__1_), .A2(
        npu_inst_pe_1_6_1_n50), .B1(npu_inst_pe_1_6_1_n117), .B2(
        npu_inst_pe_1_6_1_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_6_1_n51) );
  INV_X1 npu_inst_pe_1_6_1_U96 ( .A(npu_inst_pe_1_6_1_n51), .ZN(
        npu_inst_pe_1_6_1_n104) );
  AOI22_X1 npu_inst_pe_1_6_1_U95 ( .A1(npu_inst_int_data_y_7__1__1_), .A2(
        npu_inst_pe_1_6_1_n46), .B1(npu_inst_pe_1_6_1_n116), .B2(
        npu_inst_pe_1_6_1_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_6_1_n47) );
  INV_X1 npu_inst_pe_1_6_1_U94 ( .A(npu_inst_pe_1_6_1_n47), .ZN(
        npu_inst_pe_1_6_1_n105) );
  AOI22_X1 npu_inst_pe_1_6_1_U93 ( .A1(npu_inst_int_data_y_7__1__1_), .A2(
        npu_inst_pe_1_6_1_n42), .B1(npu_inst_pe_1_6_1_n115), .B2(
        npu_inst_pe_1_6_1_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_6_1_n43) );
  INV_X1 npu_inst_pe_1_6_1_U92 ( .A(npu_inst_pe_1_6_1_n43), .ZN(
        npu_inst_pe_1_6_1_n106) );
  AOI22_X1 npu_inst_pe_1_6_1_U91 ( .A1(npu_inst_pe_1_6_1_n38), .A2(
        npu_inst_int_data_y_7__1__1_), .B1(npu_inst_pe_1_6_1_n114), .B2(
        npu_inst_pe_1_6_1_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_6_1_n39) );
  INV_X1 npu_inst_pe_1_6_1_U90 ( .A(npu_inst_pe_1_6_1_n39), .ZN(
        npu_inst_pe_1_6_1_n107) );
  AOI22_X1 npu_inst_pe_1_6_1_U89 ( .A1(npu_inst_pe_1_6_1_n38), .A2(
        npu_inst_int_data_y_7__1__0_), .B1(npu_inst_pe_1_6_1_n114), .B2(
        npu_inst_pe_1_6_1_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_6_1_n37) );
  INV_X1 npu_inst_pe_1_6_1_U88 ( .A(npu_inst_pe_1_6_1_n37), .ZN(
        npu_inst_pe_1_6_1_n113) );
  NAND2_X1 npu_inst_pe_1_6_1_U87 ( .A1(npu_inst_pe_1_6_1_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_6_1_n60), .ZN(npu_inst_pe_1_6_1_n74) );
  OAI21_X1 npu_inst_pe_1_6_1_U86 ( .B1(npu_inst_pe_1_6_1_n63), .B2(
        npu_inst_pe_1_6_1_n60), .A(npu_inst_pe_1_6_1_n74), .ZN(
        npu_inst_pe_1_6_1_n97) );
  NAND2_X1 npu_inst_pe_1_6_1_U85 ( .A1(npu_inst_pe_1_6_1_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_6_1_n60), .ZN(npu_inst_pe_1_6_1_n73) );
  OAI21_X1 npu_inst_pe_1_6_1_U84 ( .B1(npu_inst_pe_1_6_1_n61), .B2(
        npu_inst_pe_1_6_1_n60), .A(npu_inst_pe_1_6_1_n73), .ZN(
        npu_inst_pe_1_6_1_n96) );
  NAND2_X1 npu_inst_pe_1_6_1_U83 ( .A1(npu_inst_pe_1_6_1_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_6_1_n56), .ZN(npu_inst_pe_1_6_1_n72) );
  OAI21_X1 npu_inst_pe_1_6_1_U82 ( .B1(npu_inst_pe_1_6_1_n63), .B2(
        npu_inst_pe_1_6_1_n56), .A(npu_inst_pe_1_6_1_n72), .ZN(
        npu_inst_pe_1_6_1_n95) );
  NAND2_X1 npu_inst_pe_1_6_1_U81 ( .A1(npu_inst_pe_1_6_1_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_6_1_n56), .ZN(npu_inst_pe_1_6_1_n71) );
  OAI21_X1 npu_inst_pe_1_6_1_U80 ( .B1(npu_inst_pe_1_6_1_n61), .B2(
        npu_inst_pe_1_6_1_n56), .A(npu_inst_pe_1_6_1_n71), .ZN(
        npu_inst_pe_1_6_1_n94) );
  NAND2_X1 npu_inst_pe_1_6_1_U79 ( .A1(npu_inst_pe_1_6_1_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_6_1_n52), .ZN(npu_inst_pe_1_6_1_n70) );
  OAI21_X1 npu_inst_pe_1_6_1_U78 ( .B1(npu_inst_pe_1_6_1_n63), .B2(
        npu_inst_pe_1_6_1_n52), .A(npu_inst_pe_1_6_1_n70), .ZN(
        npu_inst_pe_1_6_1_n93) );
  NAND2_X1 npu_inst_pe_1_6_1_U77 ( .A1(npu_inst_pe_1_6_1_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_6_1_n52), .ZN(npu_inst_pe_1_6_1_n69) );
  OAI21_X1 npu_inst_pe_1_6_1_U76 ( .B1(npu_inst_pe_1_6_1_n61), .B2(
        npu_inst_pe_1_6_1_n52), .A(npu_inst_pe_1_6_1_n69), .ZN(
        npu_inst_pe_1_6_1_n92) );
  NAND2_X1 npu_inst_pe_1_6_1_U75 ( .A1(npu_inst_pe_1_6_1_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_6_1_n48), .ZN(npu_inst_pe_1_6_1_n68) );
  OAI21_X1 npu_inst_pe_1_6_1_U74 ( .B1(npu_inst_pe_1_6_1_n63), .B2(
        npu_inst_pe_1_6_1_n48), .A(npu_inst_pe_1_6_1_n68), .ZN(
        npu_inst_pe_1_6_1_n91) );
  NAND2_X1 npu_inst_pe_1_6_1_U73 ( .A1(npu_inst_pe_1_6_1_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_6_1_n48), .ZN(npu_inst_pe_1_6_1_n67) );
  OAI21_X1 npu_inst_pe_1_6_1_U72 ( .B1(npu_inst_pe_1_6_1_n61), .B2(
        npu_inst_pe_1_6_1_n48), .A(npu_inst_pe_1_6_1_n67), .ZN(
        npu_inst_pe_1_6_1_n90) );
  NAND2_X1 npu_inst_pe_1_6_1_U71 ( .A1(npu_inst_pe_1_6_1_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_6_1_n44), .ZN(npu_inst_pe_1_6_1_n66) );
  OAI21_X1 npu_inst_pe_1_6_1_U70 ( .B1(npu_inst_pe_1_6_1_n63), .B2(
        npu_inst_pe_1_6_1_n44), .A(npu_inst_pe_1_6_1_n66), .ZN(
        npu_inst_pe_1_6_1_n89) );
  NAND2_X1 npu_inst_pe_1_6_1_U69 ( .A1(npu_inst_pe_1_6_1_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_6_1_n44), .ZN(npu_inst_pe_1_6_1_n65) );
  OAI21_X1 npu_inst_pe_1_6_1_U68 ( .B1(npu_inst_pe_1_6_1_n61), .B2(
        npu_inst_pe_1_6_1_n44), .A(npu_inst_pe_1_6_1_n65), .ZN(
        npu_inst_pe_1_6_1_n88) );
  NAND2_X1 npu_inst_pe_1_6_1_U67 ( .A1(npu_inst_pe_1_6_1_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_6_1_n40), .ZN(npu_inst_pe_1_6_1_n64) );
  OAI21_X1 npu_inst_pe_1_6_1_U66 ( .B1(npu_inst_pe_1_6_1_n63), .B2(
        npu_inst_pe_1_6_1_n40), .A(npu_inst_pe_1_6_1_n64), .ZN(
        npu_inst_pe_1_6_1_n87) );
  NAND2_X1 npu_inst_pe_1_6_1_U65 ( .A1(npu_inst_pe_1_6_1_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_6_1_n40), .ZN(npu_inst_pe_1_6_1_n62) );
  OAI21_X1 npu_inst_pe_1_6_1_U64 ( .B1(npu_inst_pe_1_6_1_n61), .B2(
        npu_inst_pe_1_6_1_n40), .A(npu_inst_pe_1_6_1_n62), .ZN(
        npu_inst_pe_1_6_1_n86) );
  AND2_X1 npu_inst_pe_1_6_1_U63 ( .A1(npu_inst_pe_1_6_1_N93), .A2(npu_inst_n54), .ZN(npu_inst_int_data_y_6__1__0_) );
  AND2_X1 npu_inst_pe_1_6_1_U62 ( .A1(npu_inst_n54), .A2(npu_inst_pe_1_6_1_N94), .ZN(npu_inst_int_data_y_6__1__1_) );
  NOR3_X1 npu_inst_pe_1_6_1_U61 ( .A1(npu_inst_pe_1_6_1_n26), .A2(npu_inst_n54), .A3(npu_inst_int_ckg[14]), .ZN(npu_inst_pe_1_6_1_n85) );
  OR2_X1 npu_inst_pe_1_6_1_U60 ( .A1(npu_inst_pe_1_6_1_n85), .A2(
        npu_inst_pe_1_6_1_n2), .ZN(npu_inst_pe_1_6_1_N84) );
  AND2_X1 npu_inst_pe_1_6_1_U59 ( .A1(npu_inst_pe_1_6_1_int_q_acc_0_), .A2(
        npu_inst_pe_1_6_1_n1), .ZN(npu_inst_int_data_res_6__1__0_) );
  AND2_X1 npu_inst_pe_1_6_1_U58 ( .A1(npu_inst_pe_1_6_1_n2), .A2(
        npu_inst_pe_1_6_1_int_q_acc_7_), .ZN(npu_inst_int_data_res_6__1__7_)
         );
  AND2_X1 npu_inst_pe_1_6_1_U57 ( .A1(npu_inst_pe_1_6_1_int_q_acc_1_), .A2(
        npu_inst_pe_1_6_1_n1), .ZN(npu_inst_int_data_res_6__1__1_) );
  AND2_X1 npu_inst_pe_1_6_1_U56 ( .A1(npu_inst_pe_1_6_1_int_q_acc_2_), .A2(
        npu_inst_pe_1_6_1_n1), .ZN(npu_inst_int_data_res_6__1__2_) );
  AND2_X1 npu_inst_pe_1_6_1_U55 ( .A1(npu_inst_pe_1_6_1_int_q_acc_3_), .A2(
        npu_inst_pe_1_6_1_n2), .ZN(npu_inst_int_data_res_6__1__3_) );
  AND2_X1 npu_inst_pe_1_6_1_U54 ( .A1(npu_inst_pe_1_6_1_int_q_acc_4_), .A2(
        npu_inst_pe_1_6_1_n2), .ZN(npu_inst_int_data_res_6__1__4_) );
  AND2_X1 npu_inst_pe_1_6_1_U53 ( .A1(npu_inst_pe_1_6_1_int_q_acc_5_), .A2(
        npu_inst_pe_1_6_1_n2), .ZN(npu_inst_int_data_res_6__1__5_) );
  AND2_X1 npu_inst_pe_1_6_1_U52 ( .A1(npu_inst_pe_1_6_1_int_q_acc_6_), .A2(
        npu_inst_pe_1_6_1_n2), .ZN(npu_inst_int_data_res_6__1__6_) );
  AOI222_X1 npu_inst_pe_1_6_1_U51 ( .A1(npu_inst_int_data_res_7__1__0_), .A2(
        npu_inst_pe_1_6_1_n1), .B1(npu_inst_pe_1_6_1_N73), .B2(
        npu_inst_pe_1_6_1_n76), .C1(npu_inst_pe_1_6_1_N65), .C2(
        npu_inst_pe_1_6_1_n77), .ZN(npu_inst_pe_1_6_1_n84) );
  INV_X1 npu_inst_pe_1_6_1_U50 ( .A(npu_inst_pe_1_6_1_n84), .ZN(
        npu_inst_pe_1_6_1_n101) );
  AOI222_X1 npu_inst_pe_1_6_1_U49 ( .A1(npu_inst_int_data_res_7__1__7_), .A2(
        npu_inst_pe_1_6_1_n1), .B1(npu_inst_pe_1_6_1_N80), .B2(
        npu_inst_pe_1_6_1_n76), .C1(npu_inst_pe_1_6_1_N72), .C2(
        npu_inst_pe_1_6_1_n77), .ZN(npu_inst_pe_1_6_1_n75) );
  INV_X1 npu_inst_pe_1_6_1_U48 ( .A(npu_inst_pe_1_6_1_n75), .ZN(
        npu_inst_pe_1_6_1_n33) );
  AOI222_X1 npu_inst_pe_1_6_1_U47 ( .A1(npu_inst_int_data_res_7__1__1_), .A2(
        npu_inst_pe_1_6_1_n1), .B1(npu_inst_pe_1_6_1_N74), .B2(
        npu_inst_pe_1_6_1_n76), .C1(npu_inst_pe_1_6_1_N66), .C2(
        npu_inst_pe_1_6_1_n77), .ZN(npu_inst_pe_1_6_1_n83) );
  INV_X1 npu_inst_pe_1_6_1_U46 ( .A(npu_inst_pe_1_6_1_n83), .ZN(
        npu_inst_pe_1_6_1_n100) );
  AOI222_X1 npu_inst_pe_1_6_1_U45 ( .A1(npu_inst_int_data_res_7__1__2_), .A2(
        npu_inst_pe_1_6_1_n1), .B1(npu_inst_pe_1_6_1_N75), .B2(
        npu_inst_pe_1_6_1_n76), .C1(npu_inst_pe_1_6_1_N67), .C2(
        npu_inst_pe_1_6_1_n77), .ZN(npu_inst_pe_1_6_1_n82) );
  INV_X1 npu_inst_pe_1_6_1_U44 ( .A(npu_inst_pe_1_6_1_n82), .ZN(
        npu_inst_pe_1_6_1_n99) );
  AOI222_X1 npu_inst_pe_1_6_1_U43 ( .A1(npu_inst_int_data_res_7__1__3_), .A2(
        npu_inst_pe_1_6_1_n1), .B1(npu_inst_pe_1_6_1_N76), .B2(
        npu_inst_pe_1_6_1_n76), .C1(npu_inst_pe_1_6_1_N68), .C2(
        npu_inst_pe_1_6_1_n77), .ZN(npu_inst_pe_1_6_1_n81) );
  INV_X1 npu_inst_pe_1_6_1_U42 ( .A(npu_inst_pe_1_6_1_n81), .ZN(
        npu_inst_pe_1_6_1_n98) );
  AOI222_X1 npu_inst_pe_1_6_1_U41 ( .A1(npu_inst_int_data_res_7__1__4_), .A2(
        npu_inst_pe_1_6_1_n1), .B1(npu_inst_pe_1_6_1_N77), .B2(
        npu_inst_pe_1_6_1_n76), .C1(npu_inst_pe_1_6_1_N69), .C2(
        npu_inst_pe_1_6_1_n77), .ZN(npu_inst_pe_1_6_1_n80) );
  INV_X1 npu_inst_pe_1_6_1_U40 ( .A(npu_inst_pe_1_6_1_n80), .ZN(
        npu_inst_pe_1_6_1_n36) );
  AOI222_X1 npu_inst_pe_1_6_1_U39 ( .A1(npu_inst_int_data_res_7__1__5_), .A2(
        npu_inst_pe_1_6_1_n1), .B1(npu_inst_pe_1_6_1_N78), .B2(
        npu_inst_pe_1_6_1_n76), .C1(npu_inst_pe_1_6_1_N70), .C2(
        npu_inst_pe_1_6_1_n77), .ZN(npu_inst_pe_1_6_1_n79) );
  INV_X1 npu_inst_pe_1_6_1_U38 ( .A(npu_inst_pe_1_6_1_n79), .ZN(
        npu_inst_pe_1_6_1_n35) );
  AOI222_X1 npu_inst_pe_1_6_1_U37 ( .A1(npu_inst_int_data_res_7__1__6_), .A2(
        npu_inst_pe_1_6_1_n1), .B1(npu_inst_pe_1_6_1_N79), .B2(
        npu_inst_pe_1_6_1_n76), .C1(npu_inst_pe_1_6_1_N71), .C2(
        npu_inst_pe_1_6_1_n77), .ZN(npu_inst_pe_1_6_1_n78) );
  INV_X1 npu_inst_pe_1_6_1_U36 ( .A(npu_inst_pe_1_6_1_n78), .ZN(
        npu_inst_pe_1_6_1_n34) );
  INV_X1 npu_inst_pe_1_6_1_U35 ( .A(npu_inst_pe_1_6_1_int_data_1_), .ZN(
        npu_inst_pe_1_6_1_n14) );
  AND2_X1 npu_inst_pe_1_6_1_U34 ( .A1(npu_inst_int_data_x_6__1__1_), .A2(
        npu_inst_pe_1_6_1_int_q_weight_1_), .ZN(npu_inst_pe_1_6_1_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_6_1_U33 ( .A1(npu_inst_int_data_x_6__1__0_), .A2(
        npu_inst_pe_1_6_1_int_q_weight_1_), .ZN(npu_inst_pe_1_6_1_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_6_1_U32 ( .A1(npu_inst_n54), .A2(
        npu_inst_int_data_y_7__1__1_), .B1(npu_inst_pe_1_6_1_n3), .B2(
        npu_inst_int_data_x_6__2__1_), .ZN(npu_inst_pe_1_6_1_n63) );
  AOI22_X1 npu_inst_pe_1_6_1_U31 ( .A1(npu_inst_n54), .A2(
        npu_inst_int_data_y_7__1__0_), .B1(npu_inst_pe_1_6_1_n3), .B2(
        npu_inst_int_data_x_6__2__0_), .ZN(npu_inst_pe_1_6_1_n61) );
  INV_X1 npu_inst_pe_1_6_1_U30 ( .A(npu_inst_pe_1_6_1_int_data_0_), .ZN(
        npu_inst_pe_1_6_1_n13) );
  INV_X1 npu_inst_pe_1_6_1_U29 ( .A(npu_inst_n68), .ZN(npu_inst_pe_1_6_1_n5)
         );
  OR3_X1 npu_inst_pe_1_6_1_U28 ( .A1(npu_inst_pe_1_6_1_n6), .A2(
        npu_inst_pe_1_6_1_n8), .A3(npu_inst_pe_1_6_1_n5), .ZN(
        npu_inst_pe_1_6_1_n56) );
  OR3_X1 npu_inst_pe_1_6_1_U27 ( .A1(npu_inst_pe_1_6_1_n5), .A2(
        npu_inst_pe_1_6_1_n8), .A3(npu_inst_pe_1_6_1_n7), .ZN(
        npu_inst_pe_1_6_1_n48) );
  INV_X1 npu_inst_pe_1_6_1_U26 ( .A(npu_inst_pe_1_6_1_n5), .ZN(
        npu_inst_pe_1_6_1_n4) );
  OR3_X1 npu_inst_pe_1_6_1_U25 ( .A1(npu_inst_pe_1_6_1_n4), .A2(
        npu_inst_pe_1_6_1_n8), .A3(npu_inst_pe_1_6_1_n7), .ZN(
        npu_inst_pe_1_6_1_n52) );
  OR3_X1 npu_inst_pe_1_6_1_U24 ( .A1(npu_inst_pe_1_6_1_n6), .A2(
        npu_inst_pe_1_6_1_n8), .A3(npu_inst_pe_1_6_1_n4), .ZN(
        npu_inst_pe_1_6_1_n60) );
  NOR2_X1 npu_inst_pe_1_6_1_U23 ( .A1(npu_inst_pe_1_6_1_n60), .A2(
        npu_inst_pe_1_6_1_n3), .ZN(npu_inst_pe_1_6_1_n58) );
  NOR2_X1 npu_inst_pe_1_6_1_U22 ( .A1(npu_inst_pe_1_6_1_n56), .A2(
        npu_inst_pe_1_6_1_n3), .ZN(npu_inst_pe_1_6_1_n54) );
  NOR2_X1 npu_inst_pe_1_6_1_U21 ( .A1(npu_inst_pe_1_6_1_n52), .A2(
        npu_inst_pe_1_6_1_n3), .ZN(npu_inst_pe_1_6_1_n50) );
  NOR2_X1 npu_inst_pe_1_6_1_U20 ( .A1(npu_inst_pe_1_6_1_n48), .A2(
        npu_inst_pe_1_6_1_n3), .ZN(npu_inst_pe_1_6_1_n46) );
  NOR2_X1 npu_inst_pe_1_6_1_U19 ( .A1(npu_inst_pe_1_6_1_n40), .A2(
        npu_inst_pe_1_6_1_n3), .ZN(npu_inst_pe_1_6_1_n38) );
  NOR2_X1 npu_inst_pe_1_6_1_U18 ( .A1(npu_inst_pe_1_6_1_n44), .A2(
        npu_inst_pe_1_6_1_n3), .ZN(npu_inst_pe_1_6_1_n42) );
  BUF_X1 npu_inst_pe_1_6_1_U17 ( .A(npu_inst_n95), .Z(npu_inst_pe_1_6_1_n8) );
  INV_X1 npu_inst_pe_1_6_1_U16 ( .A(npu_inst_n123), .ZN(npu_inst_pe_1_6_1_n12)
         );
  INV_X1 npu_inst_pe_1_6_1_U15 ( .A(npu_inst_pe_1_6_1_n38), .ZN(
        npu_inst_pe_1_6_1_n114) );
  INV_X1 npu_inst_pe_1_6_1_U14 ( .A(npu_inst_pe_1_6_1_n58), .ZN(
        npu_inst_pe_1_6_1_n119) );
  INV_X1 npu_inst_pe_1_6_1_U13 ( .A(npu_inst_pe_1_6_1_n54), .ZN(
        npu_inst_pe_1_6_1_n118) );
  INV_X1 npu_inst_pe_1_6_1_U12 ( .A(npu_inst_pe_1_6_1_n50), .ZN(
        npu_inst_pe_1_6_1_n117) );
  INV_X1 npu_inst_pe_1_6_1_U11 ( .A(npu_inst_pe_1_6_1_n46), .ZN(
        npu_inst_pe_1_6_1_n116) );
  INV_X1 npu_inst_pe_1_6_1_U10 ( .A(npu_inst_pe_1_6_1_n42), .ZN(
        npu_inst_pe_1_6_1_n115) );
  BUF_X1 npu_inst_pe_1_6_1_U9 ( .A(npu_inst_n14), .Z(npu_inst_pe_1_6_1_n2) );
  BUF_X1 npu_inst_pe_1_6_1_U8 ( .A(npu_inst_n14), .Z(npu_inst_pe_1_6_1_n1) );
  BUF_X1 npu_inst_pe_1_6_1_U7 ( .A(npu_inst_pe_1_6_1_n12), .Z(
        npu_inst_pe_1_6_1_n11) );
  BUF_X1 npu_inst_pe_1_6_1_U6 ( .A(npu_inst_pe_1_6_1_n12), .Z(
        npu_inst_pe_1_6_1_n10) );
  BUF_X1 npu_inst_pe_1_6_1_U5 ( .A(npu_inst_pe_1_6_1_n12), .Z(
        npu_inst_pe_1_6_1_n9) );
  NOR2_X1 npu_inst_pe_1_6_1_U4 ( .A1(npu_inst_pe_1_6_1_int_q_weight_0_), .A2(
        npu_inst_pe_1_6_1_n1), .ZN(npu_inst_pe_1_6_1_n76) );
  NOR2_X1 npu_inst_pe_1_6_1_U3 ( .A1(npu_inst_pe_1_6_1_n27), .A2(
        npu_inst_pe_1_6_1_n1), .ZN(npu_inst_pe_1_6_1_n77) );
  FA_X1 npu_inst_pe_1_6_1_sub_67_U2_1 ( .A(npu_inst_pe_1_6_1_int_q_acc_1_), 
        .B(npu_inst_pe_1_6_1_n14), .CI(npu_inst_pe_1_6_1_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_6_1_sub_67_carry_2_), .S(npu_inst_pe_1_6_1_N66) );
  FA_X1 npu_inst_pe_1_6_1_add_69_U1_1 ( .A(npu_inst_pe_1_6_1_int_q_acc_1_), 
        .B(npu_inst_pe_1_6_1_int_data_1_), .CI(
        npu_inst_pe_1_6_1_add_69_carry_1_), .CO(
        npu_inst_pe_1_6_1_add_69_carry_2_), .S(npu_inst_pe_1_6_1_N74) );
  NAND3_X1 npu_inst_pe_1_6_1_U109 ( .A1(npu_inst_pe_1_6_1_n5), .A2(
        npu_inst_pe_1_6_1_n7), .A3(npu_inst_pe_1_6_1_n8), .ZN(
        npu_inst_pe_1_6_1_n44) );
  NAND3_X1 npu_inst_pe_1_6_1_U108 ( .A1(npu_inst_pe_1_6_1_n4), .A2(
        npu_inst_pe_1_6_1_n7), .A3(npu_inst_pe_1_6_1_n8), .ZN(
        npu_inst_pe_1_6_1_n40) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_6_1_n34), .CK(
        npu_inst_pe_1_6_1_net3435), .RN(npu_inst_pe_1_6_1_n9), .Q(
        npu_inst_pe_1_6_1_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_6_1_n35), .CK(
        npu_inst_pe_1_6_1_net3435), .RN(npu_inst_pe_1_6_1_n9), .Q(
        npu_inst_pe_1_6_1_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_6_1_n36), .CK(
        npu_inst_pe_1_6_1_net3435), .RN(npu_inst_pe_1_6_1_n9), .Q(
        npu_inst_pe_1_6_1_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_6_1_n98), .CK(
        npu_inst_pe_1_6_1_net3435), .RN(npu_inst_pe_1_6_1_n9), .Q(
        npu_inst_pe_1_6_1_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_6_1_n99), .CK(
        npu_inst_pe_1_6_1_net3435), .RN(npu_inst_pe_1_6_1_n9), .Q(
        npu_inst_pe_1_6_1_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_6_1_n100), 
        .CK(npu_inst_pe_1_6_1_net3435), .RN(npu_inst_pe_1_6_1_n9), .Q(
        npu_inst_pe_1_6_1_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_6_1_n33), .CK(
        npu_inst_pe_1_6_1_net3435), .RN(npu_inst_pe_1_6_1_n9), .Q(
        npu_inst_pe_1_6_1_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_6_1_n101), 
        .CK(npu_inst_pe_1_6_1_net3435), .RN(npu_inst_pe_1_6_1_n9), .Q(
        npu_inst_pe_1_6_1_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_weight_reg_0_ ( .D(npu_inst_n109), .CK(
        npu_inst_pe_1_6_1_net3441), .RN(npu_inst_pe_1_6_1_n9), .Q(
        npu_inst_pe_1_6_1_int_q_weight_0_), .QN(npu_inst_pe_1_6_1_n27) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_weight_reg_1_ ( .D(npu_inst_n115), .CK(
        npu_inst_pe_1_6_1_net3441), .RN(npu_inst_pe_1_6_1_n9), .Q(
        npu_inst_pe_1_6_1_int_q_weight_1_), .QN(npu_inst_pe_1_6_1_n26) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_6_1_n113), 
        .CK(npu_inst_pe_1_6_1_net3441), .RN(npu_inst_pe_1_6_1_n9), .Q(
        npu_inst_pe_1_6_1_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_6_1_n107), 
        .CK(npu_inst_pe_1_6_1_net3441), .RN(npu_inst_pe_1_6_1_n9), .Q(
        npu_inst_pe_1_6_1_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_6_1_n112), 
        .CK(npu_inst_pe_1_6_1_net3441), .RN(npu_inst_pe_1_6_1_n10), .Q(
        npu_inst_pe_1_6_1_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_6_1_n106), 
        .CK(npu_inst_pe_1_6_1_net3441), .RN(npu_inst_pe_1_6_1_n10), .Q(
        npu_inst_pe_1_6_1_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_6_1_n111), 
        .CK(npu_inst_pe_1_6_1_net3441), .RN(npu_inst_pe_1_6_1_n10), .Q(
        npu_inst_pe_1_6_1_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_6_1_n105), 
        .CK(npu_inst_pe_1_6_1_net3441), .RN(npu_inst_pe_1_6_1_n10), .Q(
        npu_inst_pe_1_6_1_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_6_1_n110), 
        .CK(npu_inst_pe_1_6_1_net3441), .RN(npu_inst_pe_1_6_1_n10), .Q(
        npu_inst_pe_1_6_1_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_6_1_n104), 
        .CK(npu_inst_pe_1_6_1_net3441), .RN(npu_inst_pe_1_6_1_n10), .Q(
        npu_inst_pe_1_6_1_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_6_1_n109), 
        .CK(npu_inst_pe_1_6_1_net3441), .RN(npu_inst_pe_1_6_1_n10), .Q(
        npu_inst_pe_1_6_1_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_6_1_n103), 
        .CK(npu_inst_pe_1_6_1_net3441), .RN(npu_inst_pe_1_6_1_n10), .Q(
        npu_inst_pe_1_6_1_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_6_1_n108), 
        .CK(npu_inst_pe_1_6_1_net3441), .RN(npu_inst_pe_1_6_1_n10), .Q(
        npu_inst_pe_1_6_1_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_6_1_n102), 
        .CK(npu_inst_pe_1_6_1_net3441), .RN(npu_inst_pe_1_6_1_n10), .Q(
        npu_inst_pe_1_6_1_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_6_1_n86), 
        .CK(npu_inst_pe_1_6_1_net3441), .RN(npu_inst_pe_1_6_1_n10), .Q(
        npu_inst_pe_1_6_1_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_6_1_n87), 
        .CK(npu_inst_pe_1_6_1_net3441), .RN(npu_inst_pe_1_6_1_n10), .Q(
        npu_inst_pe_1_6_1_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_6_1_n88), 
        .CK(npu_inst_pe_1_6_1_net3441), .RN(npu_inst_pe_1_6_1_n11), .Q(
        npu_inst_pe_1_6_1_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_6_1_n89), 
        .CK(npu_inst_pe_1_6_1_net3441), .RN(npu_inst_pe_1_6_1_n11), .Q(
        npu_inst_pe_1_6_1_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_6_1_n90), 
        .CK(npu_inst_pe_1_6_1_net3441), .RN(npu_inst_pe_1_6_1_n11), .Q(
        npu_inst_pe_1_6_1_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_6_1_n91), 
        .CK(npu_inst_pe_1_6_1_net3441), .RN(npu_inst_pe_1_6_1_n11), .Q(
        npu_inst_pe_1_6_1_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_6_1_n92), 
        .CK(npu_inst_pe_1_6_1_net3441), .RN(npu_inst_pe_1_6_1_n11), .Q(
        npu_inst_pe_1_6_1_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_6_1_n93), 
        .CK(npu_inst_pe_1_6_1_net3441), .RN(npu_inst_pe_1_6_1_n11), .Q(
        npu_inst_pe_1_6_1_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_6_1_n94), 
        .CK(npu_inst_pe_1_6_1_net3441), .RN(npu_inst_pe_1_6_1_n11), .Q(
        npu_inst_pe_1_6_1_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_6_1_n95), 
        .CK(npu_inst_pe_1_6_1_net3441), .RN(npu_inst_pe_1_6_1_n11), .Q(
        npu_inst_pe_1_6_1_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_6_1_n96), 
        .CK(npu_inst_pe_1_6_1_net3441), .RN(npu_inst_pe_1_6_1_n11), .Q(
        npu_inst_pe_1_6_1_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_6_1_n97), 
        .CK(npu_inst_pe_1_6_1_net3441), .RN(npu_inst_pe_1_6_1_n11), .Q(
        npu_inst_pe_1_6_1_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_6_1_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_6_1_N84), .SE(1'b0), .GCK(npu_inst_pe_1_6_1_net3435) );
  CLKGATETST_X1 npu_inst_pe_1_6_1_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n62), .SE(1'b0), .GCK(npu_inst_pe_1_6_1_net3441) );
  MUX2_X1 npu_inst_pe_1_6_2_U162 ( .A(npu_inst_pe_1_6_2_n32), .B(
        npu_inst_pe_1_6_2_n29), .S(npu_inst_pe_1_6_2_n8), .Z(
        npu_inst_pe_1_6_2_N93) );
  MUX2_X1 npu_inst_pe_1_6_2_U161 ( .A(npu_inst_pe_1_6_2_n31), .B(
        npu_inst_pe_1_6_2_n30), .S(npu_inst_pe_1_6_2_n6), .Z(
        npu_inst_pe_1_6_2_n32) );
  MUX2_X1 npu_inst_pe_1_6_2_U160 ( .A(npu_inst_pe_1_6_2_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_6_2_int_q_reg_v_1__0_), .S(npu_inst_pe_1_6_2_n4), .Z(
        npu_inst_pe_1_6_2_n31) );
  MUX2_X1 npu_inst_pe_1_6_2_U159 ( .A(npu_inst_pe_1_6_2_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_6_2_int_q_reg_v_3__0_), .S(npu_inst_pe_1_6_2_n4), .Z(
        npu_inst_pe_1_6_2_n30) );
  MUX2_X1 npu_inst_pe_1_6_2_U158 ( .A(npu_inst_pe_1_6_2_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_6_2_int_q_reg_v_5__0_), .S(npu_inst_pe_1_6_2_n4), .Z(
        npu_inst_pe_1_6_2_n29) );
  MUX2_X1 npu_inst_pe_1_6_2_U157 ( .A(npu_inst_pe_1_6_2_n28), .B(
        npu_inst_pe_1_6_2_n23), .S(npu_inst_pe_1_6_2_n8), .Z(
        npu_inst_pe_1_6_2_N94) );
  MUX2_X1 npu_inst_pe_1_6_2_U156 ( .A(npu_inst_pe_1_6_2_n25), .B(
        npu_inst_pe_1_6_2_n24), .S(npu_inst_pe_1_6_2_n6), .Z(
        npu_inst_pe_1_6_2_n28) );
  MUX2_X1 npu_inst_pe_1_6_2_U155 ( .A(npu_inst_pe_1_6_2_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_6_2_int_q_reg_v_1__1_), .S(npu_inst_pe_1_6_2_n4), .Z(
        npu_inst_pe_1_6_2_n25) );
  MUX2_X1 npu_inst_pe_1_6_2_U154 ( .A(npu_inst_pe_1_6_2_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_6_2_int_q_reg_v_3__1_), .S(npu_inst_pe_1_6_2_n4), .Z(
        npu_inst_pe_1_6_2_n24) );
  MUX2_X1 npu_inst_pe_1_6_2_U153 ( .A(npu_inst_pe_1_6_2_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_6_2_int_q_reg_v_5__1_), .S(npu_inst_pe_1_6_2_n4), .Z(
        npu_inst_pe_1_6_2_n23) );
  MUX2_X1 npu_inst_pe_1_6_2_U152 ( .A(npu_inst_pe_1_6_2_n22), .B(
        npu_inst_pe_1_6_2_n19), .S(npu_inst_pe_1_6_2_n8), .Z(
        npu_inst_int_data_x_6__2__1_) );
  MUX2_X1 npu_inst_pe_1_6_2_U151 ( .A(npu_inst_pe_1_6_2_n21), .B(
        npu_inst_pe_1_6_2_n20), .S(npu_inst_pe_1_6_2_n6), .Z(
        npu_inst_pe_1_6_2_n22) );
  MUX2_X1 npu_inst_pe_1_6_2_U150 ( .A(npu_inst_pe_1_6_2_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_6_2_int_q_reg_h_1__1_), .S(npu_inst_pe_1_6_2_n4), .Z(
        npu_inst_pe_1_6_2_n21) );
  MUX2_X1 npu_inst_pe_1_6_2_U149 ( .A(npu_inst_pe_1_6_2_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_6_2_int_q_reg_h_3__1_), .S(npu_inst_pe_1_6_2_n4), .Z(
        npu_inst_pe_1_6_2_n20) );
  MUX2_X1 npu_inst_pe_1_6_2_U148 ( .A(npu_inst_pe_1_6_2_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_6_2_int_q_reg_h_5__1_), .S(npu_inst_pe_1_6_2_n4), .Z(
        npu_inst_pe_1_6_2_n19) );
  MUX2_X1 npu_inst_pe_1_6_2_U147 ( .A(npu_inst_pe_1_6_2_n18), .B(
        npu_inst_pe_1_6_2_n15), .S(npu_inst_pe_1_6_2_n8), .Z(
        npu_inst_int_data_x_6__2__0_) );
  MUX2_X1 npu_inst_pe_1_6_2_U146 ( .A(npu_inst_pe_1_6_2_n17), .B(
        npu_inst_pe_1_6_2_n16), .S(npu_inst_pe_1_6_2_n6), .Z(
        npu_inst_pe_1_6_2_n18) );
  MUX2_X1 npu_inst_pe_1_6_2_U145 ( .A(npu_inst_pe_1_6_2_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_6_2_int_q_reg_h_1__0_), .S(npu_inst_pe_1_6_2_n4), .Z(
        npu_inst_pe_1_6_2_n17) );
  MUX2_X1 npu_inst_pe_1_6_2_U144 ( .A(npu_inst_pe_1_6_2_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_6_2_int_q_reg_h_3__0_), .S(npu_inst_pe_1_6_2_n4), .Z(
        npu_inst_pe_1_6_2_n16) );
  MUX2_X1 npu_inst_pe_1_6_2_U143 ( .A(npu_inst_pe_1_6_2_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_6_2_int_q_reg_h_5__0_), .S(npu_inst_pe_1_6_2_n4), .Z(
        npu_inst_pe_1_6_2_n15) );
  XOR2_X1 npu_inst_pe_1_6_2_U142 ( .A(npu_inst_pe_1_6_2_int_data_0_), .B(
        npu_inst_pe_1_6_2_int_q_acc_0_), .Z(npu_inst_pe_1_6_2_N73) );
  AND2_X1 npu_inst_pe_1_6_2_U141 ( .A1(npu_inst_pe_1_6_2_int_q_acc_0_), .A2(
        npu_inst_pe_1_6_2_int_data_0_), .ZN(npu_inst_pe_1_6_2_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_6_2_U140 ( .A(npu_inst_pe_1_6_2_int_q_acc_0_), .B(
        npu_inst_pe_1_6_2_n13), .ZN(npu_inst_pe_1_6_2_N65) );
  OR2_X1 npu_inst_pe_1_6_2_U139 ( .A1(npu_inst_pe_1_6_2_n13), .A2(
        npu_inst_pe_1_6_2_int_q_acc_0_), .ZN(npu_inst_pe_1_6_2_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_6_2_U138 ( .A(npu_inst_pe_1_6_2_int_q_acc_2_), .B(
        npu_inst_pe_1_6_2_add_69_carry_2_), .Z(npu_inst_pe_1_6_2_N75) );
  AND2_X1 npu_inst_pe_1_6_2_U137 ( .A1(npu_inst_pe_1_6_2_add_69_carry_2_), 
        .A2(npu_inst_pe_1_6_2_int_q_acc_2_), .ZN(
        npu_inst_pe_1_6_2_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_6_2_U136 ( .A(npu_inst_pe_1_6_2_int_q_acc_3_), .B(
        npu_inst_pe_1_6_2_add_69_carry_3_), .Z(npu_inst_pe_1_6_2_N76) );
  AND2_X1 npu_inst_pe_1_6_2_U135 ( .A1(npu_inst_pe_1_6_2_add_69_carry_3_), 
        .A2(npu_inst_pe_1_6_2_int_q_acc_3_), .ZN(
        npu_inst_pe_1_6_2_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_6_2_U134 ( .A(npu_inst_pe_1_6_2_int_q_acc_4_), .B(
        npu_inst_pe_1_6_2_add_69_carry_4_), .Z(npu_inst_pe_1_6_2_N77) );
  AND2_X1 npu_inst_pe_1_6_2_U133 ( .A1(npu_inst_pe_1_6_2_add_69_carry_4_), 
        .A2(npu_inst_pe_1_6_2_int_q_acc_4_), .ZN(
        npu_inst_pe_1_6_2_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_6_2_U132 ( .A(npu_inst_pe_1_6_2_int_q_acc_5_), .B(
        npu_inst_pe_1_6_2_add_69_carry_5_), .Z(npu_inst_pe_1_6_2_N78) );
  AND2_X1 npu_inst_pe_1_6_2_U131 ( .A1(npu_inst_pe_1_6_2_add_69_carry_5_), 
        .A2(npu_inst_pe_1_6_2_int_q_acc_5_), .ZN(
        npu_inst_pe_1_6_2_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_6_2_U130 ( .A(npu_inst_pe_1_6_2_int_q_acc_6_), .B(
        npu_inst_pe_1_6_2_add_69_carry_6_), .Z(npu_inst_pe_1_6_2_N79) );
  AND2_X1 npu_inst_pe_1_6_2_U129 ( .A1(npu_inst_pe_1_6_2_add_69_carry_6_), 
        .A2(npu_inst_pe_1_6_2_int_q_acc_6_), .ZN(
        npu_inst_pe_1_6_2_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_6_2_U128 ( .A(npu_inst_pe_1_6_2_int_q_acc_7_), .B(
        npu_inst_pe_1_6_2_add_69_carry_7_), .Z(npu_inst_pe_1_6_2_N80) );
  XNOR2_X1 npu_inst_pe_1_6_2_U127 ( .A(npu_inst_pe_1_6_2_sub_67_carry_2_), .B(
        npu_inst_pe_1_6_2_int_q_acc_2_), .ZN(npu_inst_pe_1_6_2_N67) );
  OR2_X1 npu_inst_pe_1_6_2_U126 ( .A1(npu_inst_pe_1_6_2_int_q_acc_2_), .A2(
        npu_inst_pe_1_6_2_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_6_2_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_6_2_U125 ( .A(npu_inst_pe_1_6_2_sub_67_carry_3_), .B(
        npu_inst_pe_1_6_2_int_q_acc_3_), .ZN(npu_inst_pe_1_6_2_N68) );
  OR2_X1 npu_inst_pe_1_6_2_U124 ( .A1(npu_inst_pe_1_6_2_int_q_acc_3_), .A2(
        npu_inst_pe_1_6_2_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_6_2_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_6_2_U123 ( .A(npu_inst_pe_1_6_2_sub_67_carry_4_), .B(
        npu_inst_pe_1_6_2_int_q_acc_4_), .ZN(npu_inst_pe_1_6_2_N69) );
  OR2_X1 npu_inst_pe_1_6_2_U122 ( .A1(npu_inst_pe_1_6_2_int_q_acc_4_), .A2(
        npu_inst_pe_1_6_2_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_6_2_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_6_2_U121 ( .A(npu_inst_pe_1_6_2_sub_67_carry_5_), .B(
        npu_inst_pe_1_6_2_int_q_acc_5_), .ZN(npu_inst_pe_1_6_2_N70) );
  OR2_X1 npu_inst_pe_1_6_2_U120 ( .A1(npu_inst_pe_1_6_2_int_q_acc_5_), .A2(
        npu_inst_pe_1_6_2_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_6_2_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_6_2_U119 ( .A(npu_inst_pe_1_6_2_sub_67_carry_6_), .B(
        npu_inst_pe_1_6_2_int_q_acc_6_), .ZN(npu_inst_pe_1_6_2_N71) );
  OR2_X1 npu_inst_pe_1_6_2_U118 ( .A1(npu_inst_pe_1_6_2_int_q_acc_6_), .A2(
        npu_inst_pe_1_6_2_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_6_2_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_6_2_U117 ( .A(npu_inst_pe_1_6_2_int_q_acc_7_), .B(
        npu_inst_pe_1_6_2_sub_67_carry_7_), .ZN(npu_inst_pe_1_6_2_N72) );
  INV_X1 npu_inst_pe_1_6_2_U116 ( .A(npu_inst_n76), .ZN(npu_inst_pe_1_6_2_n7)
         );
  INV_X1 npu_inst_pe_1_6_2_U115 ( .A(npu_inst_pe_1_6_2_n7), .ZN(
        npu_inst_pe_1_6_2_n6) );
  INV_X1 npu_inst_pe_1_6_2_U114 ( .A(npu_inst_n53), .ZN(npu_inst_pe_1_6_2_n3)
         );
  AOI22_X1 npu_inst_pe_1_6_2_U113 ( .A1(npu_inst_int_data_y_7__2__0_), .A2(
        npu_inst_pe_1_6_2_n58), .B1(npu_inst_pe_1_6_2_n119), .B2(
        npu_inst_pe_1_6_2_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_6_2_n57) );
  INV_X1 npu_inst_pe_1_6_2_U112 ( .A(npu_inst_pe_1_6_2_n57), .ZN(
        npu_inst_pe_1_6_2_n108) );
  AOI22_X1 npu_inst_pe_1_6_2_U111 ( .A1(npu_inst_int_data_y_7__2__0_), .A2(
        npu_inst_pe_1_6_2_n54), .B1(npu_inst_pe_1_6_2_n118), .B2(
        npu_inst_pe_1_6_2_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_6_2_n53) );
  INV_X1 npu_inst_pe_1_6_2_U110 ( .A(npu_inst_pe_1_6_2_n53), .ZN(
        npu_inst_pe_1_6_2_n109) );
  AOI22_X1 npu_inst_pe_1_6_2_U107 ( .A1(npu_inst_int_data_y_7__2__0_), .A2(
        npu_inst_pe_1_6_2_n50), .B1(npu_inst_pe_1_6_2_n117), .B2(
        npu_inst_pe_1_6_2_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_6_2_n49) );
  INV_X1 npu_inst_pe_1_6_2_U106 ( .A(npu_inst_pe_1_6_2_n49), .ZN(
        npu_inst_pe_1_6_2_n110) );
  AOI22_X1 npu_inst_pe_1_6_2_U105 ( .A1(npu_inst_int_data_y_7__2__0_), .A2(
        npu_inst_pe_1_6_2_n46), .B1(npu_inst_pe_1_6_2_n116), .B2(
        npu_inst_pe_1_6_2_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_6_2_n45) );
  INV_X1 npu_inst_pe_1_6_2_U104 ( .A(npu_inst_pe_1_6_2_n45), .ZN(
        npu_inst_pe_1_6_2_n111) );
  AOI22_X1 npu_inst_pe_1_6_2_U103 ( .A1(npu_inst_int_data_y_7__2__0_), .A2(
        npu_inst_pe_1_6_2_n42), .B1(npu_inst_pe_1_6_2_n115), .B2(
        npu_inst_pe_1_6_2_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_6_2_n41) );
  INV_X1 npu_inst_pe_1_6_2_U102 ( .A(npu_inst_pe_1_6_2_n41), .ZN(
        npu_inst_pe_1_6_2_n112) );
  AOI22_X1 npu_inst_pe_1_6_2_U101 ( .A1(npu_inst_int_data_y_7__2__1_), .A2(
        npu_inst_pe_1_6_2_n58), .B1(npu_inst_pe_1_6_2_n119), .B2(
        npu_inst_pe_1_6_2_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_6_2_n59) );
  INV_X1 npu_inst_pe_1_6_2_U100 ( .A(npu_inst_pe_1_6_2_n59), .ZN(
        npu_inst_pe_1_6_2_n102) );
  AOI22_X1 npu_inst_pe_1_6_2_U99 ( .A1(npu_inst_int_data_y_7__2__1_), .A2(
        npu_inst_pe_1_6_2_n54), .B1(npu_inst_pe_1_6_2_n118), .B2(
        npu_inst_pe_1_6_2_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_6_2_n55) );
  INV_X1 npu_inst_pe_1_6_2_U98 ( .A(npu_inst_pe_1_6_2_n55), .ZN(
        npu_inst_pe_1_6_2_n103) );
  AOI22_X1 npu_inst_pe_1_6_2_U97 ( .A1(npu_inst_int_data_y_7__2__1_), .A2(
        npu_inst_pe_1_6_2_n50), .B1(npu_inst_pe_1_6_2_n117), .B2(
        npu_inst_pe_1_6_2_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_6_2_n51) );
  INV_X1 npu_inst_pe_1_6_2_U96 ( .A(npu_inst_pe_1_6_2_n51), .ZN(
        npu_inst_pe_1_6_2_n104) );
  AOI22_X1 npu_inst_pe_1_6_2_U95 ( .A1(npu_inst_int_data_y_7__2__1_), .A2(
        npu_inst_pe_1_6_2_n46), .B1(npu_inst_pe_1_6_2_n116), .B2(
        npu_inst_pe_1_6_2_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_6_2_n47) );
  INV_X1 npu_inst_pe_1_6_2_U94 ( .A(npu_inst_pe_1_6_2_n47), .ZN(
        npu_inst_pe_1_6_2_n105) );
  AOI22_X1 npu_inst_pe_1_6_2_U93 ( .A1(npu_inst_int_data_y_7__2__1_), .A2(
        npu_inst_pe_1_6_2_n42), .B1(npu_inst_pe_1_6_2_n115), .B2(
        npu_inst_pe_1_6_2_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_6_2_n43) );
  INV_X1 npu_inst_pe_1_6_2_U92 ( .A(npu_inst_pe_1_6_2_n43), .ZN(
        npu_inst_pe_1_6_2_n106) );
  AOI22_X1 npu_inst_pe_1_6_2_U91 ( .A1(npu_inst_pe_1_6_2_n38), .A2(
        npu_inst_int_data_y_7__2__1_), .B1(npu_inst_pe_1_6_2_n114), .B2(
        npu_inst_pe_1_6_2_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_6_2_n39) );
  INV_X1 npu_inst_pe_1_6_2_U90 ( .A(npu_inst_pe_1_6_2_n39), .ZN(
        npu_inst_pe_1_6_2_n107) );
  AOI22_X1 npu_inst_pe_1_6_2_U89 ( .A1(npu_inst_pe_1_6_2_n38), .A2(
        npu_inst_int_data_y_7__2__0_), .B1(npu_inst_pe_1_6_2_n114), .B2(
        npu_inst_pe_1_6_2_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_6_2_n37) );
  INV_X1 npu_inst_pe_1_6_2_U88 ( .A(npu_inst_pe_1_6_2_n37), .ZN(
        npu_inst_pe_1_6_2_n113) );
  NAND2_X1 npu_inst_pe_1_6_2_U87 ( .A1(npu_inst_pe_1_6_2_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_6_2_n60), .ZN(npu_inst_pe_1_6_2_n74) );
  OAI21_X1 npu_inst_pe_1_6_2_U86 ( .B1(npu_inst_pe_1_6_2_n63), .B2(
        npu_inst_pe_1_6_2_n60), .A(npu_inst_pe_1_6_2_n74), .ZN(
        npu_inst_pe_1_6_2_n97) );
  NAND2_X1 npu_inst_pe_1_6_2_U85 ( .A1(npu_inst_pe_1_6_2_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_6_2_n60), .ZN(npu_inst_pe_1_6_2_n73) );
  OAI21_X1 npu_inst_pe_1_6_2_U84 ( .B1(npu_inst_pe_1_6_2_n61), .B2(
        npu_inst_pe_1_6_2_n60), .A(npu_inst_pe_1_6_2_n73), .ZN(
        npu_inst_pe_1_6_2_n96) );
  NAND2_X1 npu_inst_pe_1_6_2_U83 ( .A1(npu_inst_pe_1_6_2_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_6_2_n56), .ZN(npu_inst_pe_1_6_2_n72) );
  OAI21_X1 npu_inst_pe_1_6_2_U82 ( .B1(npu_inst_pe_1_6_2_n63), .B2(
        npu_inst_pe_1_6_2_n56), .A(npu_inst_pe_1_6_2_n72), .ZN(
        npu_inst_pe_1_6_2_n95) );
  NAND2_X1 npu_inst_pe_1_6_2_U81 ( .A1(npu_inst_pe_1_6_2_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_6_2_n56), .ZN(npu_inst_pe_1_6_2_n71) );
  OAI21_X1 npu_inst_pe_1_6_2_U80 ( .B1(npu_inst_pe_1_6_2_n61), .B2(
        npu_inst_pe_1_6_2_n56), .A(npu_inst_pe_1_6_2_n71), .ZN(
        npu_inst_pe_1_6_2_n94) );
  NAND2_X1 npu_inst_pe_1_6_2_U79 ( .A1(npu_inst_pe_1_6_2_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_6_2_n52), .ZN(npu_inst_pe_1_6_2_n70) );
  OAI21_X1 npu_inst_pe_1_6_2_U78 ( .B1(npu_inst_pe_1_6_2_n63), .B2(
        npu_inst_pe_1_6_2_n52), .A(npu_inst_pe_1_6_2_n70), .ZN(
        npu_inst_pe_1_6_2_n93) );
  NAND2_X1 npu_inst_pe_1_6_2_U77 ( .A1(npu_inst_pe_1_6_2_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_6_2_n52), .ZN(npu_inst_pe_1_6_2_n69) );
  OAI21_X1 npu_inst_pe_1_6_2_U76 ( .B1(npu_inst_pe_1_6_2_n61), .B2(
        npu_inst_pe_1_6_2_n52), .A(npu_inst_pe_1_6_2_n69), .ZN(
        npu_inst_pe_1_6_2_n92) );
  NAND2_X1 npu_inst_pe_1_6_2_U75 ( .A1(npu_inst_pe_1_6_2_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_6_2_n48), .ZN(npu_inst_pe_1_6_2_n68) );
  OAI21_X1 npu_inst_pe_1_6_2_U74 ( .B1(npu_inst_pe_1_6_2_n63), .B2(
        npu_inst_pe_1_6_2_n48), .A(npu_inst_pe_1_6_2_n68), .ZN(
        npu_inst_pe_1_6_2_n91) );
  NAND2_X1 npu_inst_pe_1_6_2_U73 ( .A1(npu_inst_pe_1_6_2_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_6_2_n48), .ZN(npu_inst_pe_1_6_2_n67) );
  OAI21_X1 npu_inst_pe_1_6_2_U72 ( .B1(npu_inst_pe_1_6_2_n61), .B2(
        npu_inst_pe_1_6_2_n48), .A(npu_inst_pe_1_6_2_n67), .ZN(
        npu_inst_pe_1_6_2_n90) );
  NAND2_X1 npu_inst_pe_1_6_2_U71 ( .A1(npu_inst_pe_1_6_2_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_6_2_n44), .ZN(npu_inst_pe_1_6_2_n66) );
  OAI21_X1 npu_inst_pe_1_6_2_U70 ( .B1(npu_inst_pe_1_6_2_n63), .B2(
        npu_inst_pe_1_6_2_n44), .A(npu_inst_pe_1_6_2_n66), .ZN(
        npu_inst_pe_1_6_2_n89) );
  NAND2_X1 npu_inst_pe_1_6_2_U69 ( .A1(npu_inst_pe_1_6_2_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_6_2_n44), .ZN(npu_inst_pe_1_6_2_n65) );
  OAI21_X1 npu_inst_pe_1_6_2_U68 ( .B1(npu_inst_pe_1_6_2_n61), .B2(
        npu_inst_pe_1_6_2_n44), .A(npu_inst_pe_1_6_2_n65), .ZN(
        npu_inst_pe_1_6_2_n88) );
  NAND2_X1 npu_inst_pe_1_6_2_U67 ( .A1(npu_inst_pe_1_6_2_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_6_2_n40), .ZN(npu_inst_pe_1_6_2_n64) );
  OAI21_X1 npu_inst_pe_1_6_2_U66 ( .B1(npu_inst_pe_1_6_2_n63), .B2(
        npu_inst_pe_1_6_2_n40), .A(npu_inst_pe_1_6_2_n64), .ZN(
        npu_inst_pe_1_6_2_n87) );
  NAND2_X1 npu_inst_pe_1_6_2_U65 ( .A1(npu_inst_pe_1_6_2_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_6_2_n40), .ZN(npu_inst_pe_1_6_2_n62) );
  OAI21_X1 npu_inst_pe_1_6_2_U64 ( .B1(npu_inst_pe_1_6_2_n61), .B2(
        npu_inst_pe_1_6_2_n40), .A(npu_inst_pe_1_6_2_n62), .ZN(
        npu_inst_pe_1_6_2_n86) );
  AND2_X1 npu_inst_pe_1_6_2_U63 ( .A1(npu_inst_pe_1_6_2_N93), .A2(npu_inst_n53), .ZN(npu_inst_int_data_y_6__2__0_) );
  AND2_X1 npu_inst_pe_1_6_2_U62 ( .A1(npu_inst_n53), .A2(npu_inst_pe_1_6_2_N94), .ZN(npu_inst_int_data_y_6__2__1_) );
  NOR3_X1 npu_inst_pe_1_6_2_U61 ( .A1(npu_inst_pe_1_6_2_n26), .A2(npu_inst_n53), .A3(npu_inst_int_ckg[13]), .ZN(npu_inst_pe_1_6_2_n85) );
  OR2_X1 npu_inst_pe_1_6_2_U60 ( .A1(npu_inst_pe_1_6_2_n85), .A2(
        npu_inst_pe_1_6_2_n2), .ZN(npu_inst_pe_1_6_2_N84) );
  AND2_X1 npu_inst_pe_1_6_2_U59 ( .A1(npu_inst_pe_1_6_2_int_q_acc_0_), .A2(
        npu_inst_pe_1_6_2_n1), .ZN(npu_inst_int_data_res_6__2__0_) );
  AND2_X1 npu_inst_pe_1_6_2_U58 ( .A1(npu_inst_pe_1_6_2_n2), .A2(
        npu_inst_pe_1_6_2_int_q_acc_7_), .ZN(npu_inst_int_data_res_6__2__7_)
         );
  AND2_X1 npu_inst_pe_1_6_2_U57 ( .A1(npu_inst_pe_1_6_2_int_q_acc_1_), .A2(
        npu_inst_pe_1_6_2_n1), .ZN(npu_inst_int_data_res_6__2__1_) );
  AND2_X1 npu_inst_pe_1_6_2_U56 ( .A1(npu_inst_pe_1_6_2_int_q_acc_2_), .A2(
        npu_inst_pe_1_6_2_n1), .ZN(npu_inst_int_data_res_6__2__2_) );
  AND2_X1 npu_inst_pe_1_6_2_U55 ( .A1(npu_inst_pe_1_6_2_int_q_acc_3_), .A2(
        npu_inst_pe_1_6_2_n2), .ZN(npu_inst_int_data_res_6__2__3_) );
  AND2_X1 npu_inst_pe_1_6_2_U54 ( .A1(npu_inst_pe_1_6_2_int_q_acc_4_), .A2(
        npu_inst_pe_1_6_2_n2), .ZN(npu_inst_int_data_res_6__2__4_) );
  AND2_X1 npu_inst_pe_1_6_2_U53 ( .A1(npu_inst_pe_1_6_2_int_q_acc_5_), .A2(
        npu_inst_pe_1_6_2_n2), .ZN(npu_inst_int_data_res_6__2__5_) );
  AND2_X1 npu_inst_pe_1_6_2_U52 ( .A1(npu_inst_pe_1_6_2_int_q_acc_6_), .A2(
        npu_inst_pe_1_6_2_n2), .ZN(npu_inst_int_data_res_6__2__6_) );
  AOI222_X1 npu_inst_pe_1_6_2_U51 ( .A1(npu_inst_int_data_res_7__2__0_), .A2(
        npu_inst_pe_1_6_2_n1), .B1(npu_inst_pe_1_6_2_N73), .B2(
        npu_inst_pe_1_6_2_n76), .C1(npu_inst_pe_1_6_2_N65), .C2(
        npu_inst_pe_1_6_2_n77), .ZN(npu_inst_pe_1_6_2_n84) );
  INV_X1 npu_inst_pe_1_6_2_U50 ( .A(npu_inst_pe_1_6_2_n84), .ZN(
        npu_inst_pe_1_6_2_n101) );
  AOI222_X1 npu_inst_pe_1_6_2_U49 ( .A1(npu_inst_int_data_res_7__2__7_), .A2(
        npu_inst_pe_1_6_2_n1), .B1(npu_inst_pe_1_6_2_N80), .B2(
        npu_inst_pe_1_6_2_n76), .C1(npu_inst_pe_1_6_2_N72), .C2(
        npu_inst_pe_1_6_2_n77), .ZN(npu_inst_pe_1_6_2_n75) );
  INV_X1 npu_inst_pe_1_6_2_U48 ( .A(npu_inst_pe_1_6_2_n75), .ZN(
        npu_inst_pe_1_6_2_n33) );
  AOI222_X1 npu_inst_pe_1_6_2_U47 ( .A1(npu_inst_int_data_res_7__2__1_), .A2(
        npu_inst_pe_1_6_2_n1), .B1(npu_inst_pe_1_6_2_N74), .B2(
        npu_inst_pe_1_6_2_n76), .C1(npu_inst_pe_1_6_2_N66), .C2(
        npu_inst_pe_1_6_2_n77), .ZN(npu_inst_pe_1_6_2_n83) );
  INV_X1 npu_inst_pe_1_6_2_U46 ( .A(npu_inst_pe_1_6_2_n83), .ZN(
        npu_inst_pe_1_6_2_n100) );
  AOI222_X1 npu_inst_pe_1_6_2_U45 ( .A1(npu_inst_int_data_res_7__2__2_), .A2(
        npu_inst_pe_1_6_2_n1), .B1(npu_inst_pe_1_6_2_N75), .B2(
        npu_inst_pe_1_6_2_n76), .C1(npu_inst_pe_1_6_2_N67), .C2(
        npu_inst_pe_1_6_2_n77), .ZN(npu_inst_pe_1_6_2_n82) );
  INV_X1 npu_inst_pe_1_6_2_U44 ( .A(npu_inst_pe_1_6_2_n82), .ZN(
        npu_inst_pe_1_6_2_n99) );
  AOI222_X1 npu_inst_pe_1_6_2_U43 ( .A1(npu_inst_int_data_res_7__2__3_), .A2(
        npu_inst_pe_1_6_2_n1), .B1(npu_inst_pe_1_6_2_N76), .B2(
        npu_inst_pe_1_6_2_n76), .C1(npu_inst_pe_1_6_2_N68), .C2(
        npu_inst_pe_1_6_2_n77), .ZN(npu_inst_pe_1_6_2_n81) );
  INV_X1 npu_inst_pe_1_6_2_U42 ( .A(npu_inst_pe_1_6_2_n81), .ZN(
        npu_inst_pe_1_6_2_n98) );
  AOI222_X1 npu_inst_pe_1_6_2_U41 ( .A1(npu_inst_int_data_res_7__2__4_), .A2(
        npu_inst_pe_1_6_2_n1), .B1(npu_inst_pe_1_6_2_N77), .B2(
        npu_inst_pe_1_6_2_n76), .C1(npu_inst_pe_1_6_2_N69), .C2(
        npu_inst_pe_1_6_2_n77), .ZN(npu_inst_pe_1_6_2_n80) );
  INV_X1 npu_inst_pe_1_6_2_U40 ( .A(npu_inst_pe_1_6_2_n80), .ZN(
        npu_inst_pe_1_6_2_n36) );
  AOI222_X1 npu_inst_pe_1_6_2_U39 ( .A1(npu_inst_int_data_res_7__2__5_), .A2(
        npu_inst_pe_1_6_2_n1), .B1(npu_inst_pe_1_6_2_N78), .B2(
        npu_inst_pe_1_6_2_n76), .C1(npu_inst_pe_1_6_2_N70), .C2(
        npu_inst_pe_1_6_2_n77), .ZN(npu_inst_pe_1_6_2_n79) );
  INV_X1 npu_inst_pe_1_6_2_U38 ( .A(npu_inst_pe_1_6_2_n79), .ZN(
        npu_inst_pe_1_6_2_n35) );
  AOI222_X1 npu_inst_pe_1_6_2_U37 ( .A1(npu_inst_int_data_res_7__2__6_), .A2(
        npu_inst_pe_1_6_2_n1), .B1(npu_inst_pe_1_6_2_N79), .B2(
        npu_inst_pe_1_6_2_n76), .C1(npu_inst_pe_1_6_2_N71), .C2(
        npu_inst_pe_1_6_2_n77), .ZN(npu_inst_pe_1_6_2_n78) );
  INV_X1 npu_inst_pe_1_6_2_U36 ( .A(npu_inst_pe_1_6_2_n78), .ZN(
        npu_inst_pe_1_6_2_n34) );
  INV_X1 npu_inst_pe_1_6_2_U35 ( .A(npu_inst_pe_1_6_2_int_data_1_), .ZN(
        npu_inst_pe_1_6_2_n14) );
  AND2_X1 npu_inst_pe_1_6_2_U34 ( .A1(npu_inst_int_data_x_6__2__1_), .A2(
        npu_inst_pe_1_6_2_int_q_weight_1_), .ZN(npu_inst_pe_1_6_2_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_6_2_U33 ( .A1(npu_inst_int_data_x_6__2__0_), .A2(
        npu_inst_pe_1_6_2_int_q_weight_1_), .ZN(npu_inst_pe_1_6_2_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_6_2_U32 ( .A1(npu_inst_n53), .A2(
        npu_inst_int_data_y_7__2__1_), .B1(npu_inst_pe_1_6_2_n3), .B2(
        npu_inst_int_data_x_6__3__1_), .ZN(npu_inst_pe_1_6_2_n63) );
  AOI22_X1 npu_inst_pe_1_6_2_U31 ( .A1(npu_inst_n53), .A2(
        npu_inst_int_data_y_7__2__0_), .B1(npu_inst_pe_1_6_2_n3), .B2(
        npu_inst_int_data_x_6__3__0_), .ZN(npu_inst_pe_1_6_2_n61) );
  INV_X1 npu_inst_pe_1_6_2_U30 ( .A(npu_inst_pe_1_6_2_int_data_0_), .ZN(
        npu_inst_pe_1_6_2_n13) );
  INV_X1 npu_inst_pe_1_6_2_U29 ( .A(npu_inst_n68), .ZN(npu_inst_pe_1_6_2_n5)
         );
  OR3_X1 npu_inst_pe_1_6_2_U28 ( .A1(npu_inst_pe_1_6_2_n6), .A2(
        npu_inst_pe_1_6_2_n8), .A3(npu_inst_pe_1_6_2_n5), .ZN(
        npu_inst_pe_1_6_2_n56) );
  OR3_X1 npu_inst_pe_1_6_2_U27 ( .A1(npu_inst_pe_1_6_2_n5), .A2(
        npu_inst_pe_1_6_2_n8), .A3(npu_inst_pe_1_6_2_n7), .ZN(
        npu_inst_pe_1_6_2_n48) );
  INV_X1 npu_inst_pe_1_6_2_U26 ( .A(npu_inst_pe_1_6_2_n5), .ZN(
        npu_inst_pe_1_6_2_n4) );
  OR3_X1 npu_inst_pe_1_6_2_U25 ( .A1(npu_inst_pe_1_6_2_n4), .A2(
        npu_inst_pe_1_6_2_n8), .A3(npu_inst_pe_1_6_2_n7), .ZN(
        npu_inst_pe_1_6_2_n52) );
  OR3_X1 npu_inst_pe_1_6_2_U24 ( .A1(npu_inst_pe_1_6_2_n6), .A2(
        npu_inst_pe_1_6_2_n8), .A3(npu_inst_pe_1_6_2_n4), .ZN(
        npu_inst_pe_1_6_2_n60) );
  NOR2_X1 npu_inst_pe_1_6_2_U23 ( .A1(npu_inst_pe_1_6_2_n60), .A2(
        npu_inst_pe_1_6_2_n3), .ZN(npu_inst_pe_1_6_2_n58) );
  NOR2_X1 npu_inst_pe_1_6_2_U22 ( .A1(npu_inst_pe_1_6_2_n56), .A2(
        npu_inst_pe_1_6_2_n3), .ZN(npu_inst_pe_1_6_2_n54) );
  NOR2_X1 npu_inst_pe_1_6_2_U21 ( .A1(npu_inst_pe_1_6_2_n52), .A2(
        npu_inst_pe_1_6_2_n3), .ZN(npu_inst_pe_1_6_2_n50) );
  NOR2_X1 npu_inst_pe_1_6_2_U20 ( .A1(npu_inst_pe_1_6_2_n48), .A2(
        npu_inst_pe_1_6_2_n3), .ZN(npu_inst_pe_1_6_2_n46) );
  NOR2_X1 npu_inst_pe_1_6_2_U19 ( .A1(npu_inst_pe_1_6_2_n40), .A2(
        npu_inst_pe_1_6_2_n3), .ZN(npu_inst_pe_1_6_2_n38) );
  NOR2_X1 npu_inst_pe_1_6_2_U18 ( .A1(npu_inst_pe_1_6_2_n44), .A2(
        npu_inst_pe_1_6_2_n3), .ZN(npu_inst_pe_1_6_2_n42) );
  BUF_X1 npu_inst_pe_1_6_2_U17 ( .A(npu_inst_n95), .Z(npu_inst_pe_1_6_2_n8) );
  INV_X1 npu_inst_pe_1_6_2_U16 ( .A(npu_inst_n123), .ZN(npu_inst_pe_1_6_2_n12)
         );
  INV_X1 npu_inst_pe_1_6_2_U15 ( .A(npu_inst_pe_1_6_2_n38), .ZN(
        npu_inst_pe_1_6_2_n114) );
  INV_X1 npu_inst_pe_1_6_2_U14 ( .A(npu_inst_pe_1_6_2_n58), .ZN(
        npu_inst_pe_1_6_2_n119) );
  INV_X1 npu_inst_pe_1_6_2_U13 ( .A(npu_inst_pe_1_6_2_n54), .ZN(
        npu_inst_pe_1_6_2_n118) );
  INV_X1 npu_inst_pe_1_6_2_U12 ( .A(npu_inst_pe_1_6_2_n50), .ZN(
        npu_inst_pe_1_6_2_n117) );
  INV_X1 npu_inst_pe_1_6_2_U11 ( .A(npu_inst_pe_1_6_2_n46), .ZN(
        npu_inst_pe_1_6_2_n116) );
  INV_X1 npu_inst_pe_1_6_2_U10 ( .A(npu_inst_pe_1_6_2_n42), .ZN(
        npu_inst_pe_1_6_2_n115) );
  BUF_X1 npu_inst_pe_1_6_2_U9 ( .A(npu_inst_n13), .Z(npu_inst_pe_1_6_2_n2) );
  BUF_X1 npu_inst_pe_1_6_2_U8 ( .A(npu_inst_n13), .Z(npu_inst_pe_1_6_2_n1) );
  BUF_X1 npu_inst_pe_1_6_2_U7 ( .A(npu_inst_pe_1_6_2_n12), .Z(
        npu_inst_pe_1_6_2_n11) );
  BUF_X1 npu_inst_pe_1_6_2_U6 ( .A(npu_inst_pe_1_6_2_n12), .Z(
        npu_inst_pe_1_6_2_n10) );
  BUF_X1 npu_inst_pe_1_6_2_U5 ( .A(npu_inst_pe_1_6_2_n12), .Z(
        npu_inst_pe_1_6_2_n9) );
  NOR2_X1 npu_inst_pe_1_6_2_U4 ( .A1(npu_inst_pe_1_6_2_int_q_weight_0_), .A2(
        npu_inst_pe_1_6_2_n1), .ZN(npu_inst_pe_1_6_2_n76) );
  NOR2_X1 npu_inst_pe_1_6_2_U3 ( .A1(npu_inst_pe_1_6_2_n27), .A2(
        npu_inst_pe_1_6_2_n1), .ZN(npu_inst_pe_1_6_2_n77) );
  FA_X1 npu_inst_pe_1_6_2_sub_67_U2_1 ( .A(npu_inst_pe_1_6_2_int_q_acc_1_), 
        .B(npu_inst_pe_1_6_2_n14), .CI(npu_inst_pe_1_6_2_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_6_2_sub_67_carry_2_), .S(npu_inst_pe_1_6_2_N66) );
  FA_X1 npu_inst_pe_1_6_2_add_69_U1_1 ( .A(npu_inst_pe_1_6_2_int_q_acc_1_), 
        .B(npu_inst_pe_1_6_2_int_data_1_), .CI(
        npu_inst_pe_1_6_2_add_69_carry_1_), .CO(
        npu_inst_pe_1_6_2_add_69_carry_2_), .S(npu_inst_pe_1_6_2_N74) );
  NAND3_X1 npu_inst_pe_1_6_2_U109 ( .A1(npu_inst_pe_1_6_2_n5), .A2(
        npu_inst_pe_1_6_2_n7), .A3(npu_inst_pe_1_6_2_n8), .ZN(
        npu_inst_pe_1_6_2_n44) );
  NAND3_X1 npu_inst_pe_1_6_2_U108 ( .A1(npu_inst_pe_1_6_2_n4), .A2(
        npu_inst_pe_1_6_2_n7), .A3(npu_inst_pe_1_6_2_n8), .ZN(
        npu_inst_pe_1_6_2_n40) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_6_2_n34), .CK(
        npu_inst_pe_1_6_2_net3412), .RN(npu_inst_pe_1_6_2_n9), .Q(
        npu_inst_pe_1_6_2_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_6_2_n35), .CK(
        npu_inst_pe_1_6_2_net3412), .RN(npu_inst_pe_1_6_2_n9), .Q(
        npu_inst_pe_1_6_2_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_6_2_n36), .CK(
        npu_inst_pe_1_6_2_net3412), .RN(npu_inst_pe_1_6_2_n9), .Q(
        npu_inst_pe_1_6_2_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_6_2_n98), .CK(
        npu_inst_pe_1_6_2_net3412), .RN(npu_inst_pe_1_6_2_n9), .Q(
        npu_inst_pe_1_6_2_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_6_2_n99), .CK(
        npu_inst_pe_1_6_2_net3412), .RN(npu_inst_pe_1_6_2_n9), .Q(
        npu_inst_pe_1_6_2_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_6_2_n100), 
        .CK(npu_inst_pe_1_6_2_net3412), .RN(npu_inst_pe_1_6_2_n9), .Q(
        npu_inst_pe_1_6_2_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_6_2_n33), .CK(
        npu_inst_pe_1_6_2_net3412), .RN(npu_inst_pe_1_6_2_n9), .Q(
        npu_inst_pe_1_6_2_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_6_2_n101), 
        .CK(npu_inst_pe_1_6_2_net3412), .RN(npu_inst_pe_1_6_2_n9), .Q(
        npu_inst_pe_1_6_2_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_weight_reg_0_ ( .D(npu_inst_n109), .CK(
        npu_inst_pe_1_6_2_net3418), .RN(npu_inst_pe_1_6_2_n9), .Q(
        npu_inst_pe_1_6_2_int_q_weight_0_), .QN(npu_inst_pe_1_6_2_n27) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_weight_reg_1_ ( .D(npu_inst_n115), .CK(
        npu_inst_pe_1_6_2_net3418), .RN(npu_inst_pe_1_6_2_n9), .Q(
        npu_inst_pe_1_6_2_int_q_weight_1_), .QN(npu_inst_pe_1_6_2_n26) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_6_2_n113), 
        .CK(npu_inst_pe_1_6_2_net3418), .RN(npu_inst_pe_1_6_2_n9), .Q(
        npu_inst_pe_1_6_2_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_6_2_n107), 
        .CK(npu_inst_pe_1_6_2_net3418), .RN(npu_inst_pe_1_6_2_n9), .Q(
        npu_inst_pe_1_6_2_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_6_2_n112), 
        .CK(npu_inst_pe_1_6_2_net3418), .RN(npu_inst_pe_1_6_2_n10), .Q(
        npu_inst_pe_1_6_2_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_6_2_n106), 
        .CK(npu_inst_pe_1_6_2_net3418), .RN(npu_inst_pe_1_6_2_n10), .Q(
        npu_inst_pe_1_6_2_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_6_2_n111), 
        .CK(npu_inst_pe_1_6_2_net3418), .RN(npu_inst_pe_1_6_2_n10), .Q(
        npu_inst_pe_1_6_2_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_6_2_n105), 
        .CK(npu_inst_pe_1_6_2_net3418), .RN(npu_inst_pe_1_6_2_n10), .Q(
        npu_inst_pe_1_6_2_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_6_2_n110), 
        .CK(npu_inst_pe_1_6_2_net3418), .RN(npu_inst_pe_1_6_2_n10), .Q(
        npu_inst_pe_1_6_2_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_6_2_n104), 
        .CK(npu_inst_pe_1_6_2_net3418), .RN(npu_inst_pe_1_6_2_n10), .Q(
        npu_inst_pe_1_6_2_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_6_2_n109), 
        .CK(npu_inst_pe_1_6_2_net3418), .RN(npu_inst_pe_1_6_2_n10), .Q(
        npu_inst_pe_1_6_2_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_6_2_n103), 
        .CK(npu_inst_pe_1_6_2_net3418), .RN(npu_inst_pe_1_6_2_n10), .Q(
        npu_inst_pe_1_6_2_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_6_2_n108), 
        .CK(npu_inst_pe_1_6_2_net3418), .RN(npu_inst_pe_1_6_2_n10), .Q(
        npu_inst_pe_1_6_2_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_6_2_n102), 
        .CK(npu_inst_pe_1_6_2_net3418), .RN(npu_inst_pe_1_6_2_n10), .Q(
        npu_inst_pe_1_6_2_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_6_2_n86), 
        .CK(npu_inst_pe_1_6_2_net3418), .RN(npu_inst_pe_1_6_2_n10), .Q(
        npu_inst_pe_1_6_2_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_6_2_n87), 
        .CK(npu_inst_pe_1_6_2_net3418), .RN(npu_inst_pe_1_6_2_n10), .Q(
        npu_inst_pe_1_6_2_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_6_2_n88), 
        .CK(npu_inst_pe_1_6_2_net3418), .RN(npu_inst_pe_1_6_2_n11), .Q(
        npu_inst_pe_1_6_2_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_6_2_n89), 
        .CK(npu_inst_pe_1_6_2_net3418), .RN(npu_inst_pe_1_6_2_n11), .Q(
        npu_inst_pe_1_6_2_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_6_2_n90), 
        .CK(npu_inst_pe_1_6_2_net3418), .RN(npu_inst_pe_1_6_2_n11), .Q(
        npu_inst_pe_1_6_2_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_6_2_n91), 
        .CK(npu_inst_pe_1_6_2_net3418), .RN(npu_inst_pe_1_6_2_n11), .Q(
        npu_inst_pe_1_6_2_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_6_2_n92), 
        .CK(npu_inst_pe_1_6_2_net3418), .RN(npu_inst_pe_1_6_2_n11), .Q(
        npu_inst_pe_1_6_2_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_6_2_n93), 
        .CK(npu_inst_pe_1_6_2_net3418), .RN(npu_inst_pe_1_6_2_n11), .Q(
        npu_inst_pe_1_6_2_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_6_2_n94), 
        .CK(npu_inst_pe_1_6_2_net3418), .RN(npu_inst_pe_1_6_2_n11), .Q(
        npu_inst_pe_1_6_2_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_6_2_n95), 
        .CK(npu_inst_pe_1_6_2_net3418), .RN(npu_inst_pe_1_6_2_n11), .Q(
        npu_inst_pe_1_6_2_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_6_2_n96), 
        .CK(npu_inst_pe_1_6_2_net3418), .RN(npu_inst_pe_1_6_2_n11), .Q(
        npu_inst_pe_1_6_2_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_6_2_n97), 
        .CK(npu_inst_pe_1_6_2_net3418), .RN(npu_inst_pe_1_6_2_n11), .Q(
        npu_inst_pe_1_6_2_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_6_2_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_6_2_N84), .SE(1'b0), .GCK(npu_inst_pe_1_6_2_net3412) );
  CLKGATETST_X1 npu_inst_pe_1_6_2_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n62), .SE(1'b0), .GCK(npu_inst_pe_1_6_2_net3418) );
  MUX2_X1 npu_inst_pe_1_6_3_U162 ( .A(npu_inst_pe_1_6_3_n32), .B(
        npu_inst_pe_1_6_3_n29), .S(npu_inst_pe_1_6_3_n8), .Z(
        npu_inst_pe_1_6_3_N93) );
  MUX2_X1 npu_inst_pe_1_6_3_U161 ( .A(npu_inst_pe_1_6_3_n31), .B(
        npu_inst_pe_1_6_3_n30), .S(npu_inst_pe_1_6_3_n6), .Z(
        npu_inst_pe_1_6_3_n32) );
  MUX2_X1 npu_inst_pe_1_6_3_U160 ( .A(npu_inst_pe_1_6_3_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_6_3_int_q_reg_v_1__0_), .S(npu_inst_pe_1_6_3_n4), .Z(
        npu_inst_pe_1_6_3_n31) );
  MUX2_X1 npu_inst_pe_1_6_3_U159 ( .A(npu_inst_pe_1_6_3_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_6_3_int_q_reg_v_3__0_), .S(npu_inst_pe_1_6_3_n4), .Z(
        npu_inst_pe_1_6_3_n30) );
  MUX2_X1 npu_inst_pe_1_6_3_U158 ( .A(npu_inst_pe_1_6_3_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_6_3_int_q_reg_v_5__0_), .S(npu_inst_pe_1_6_3_n4), .Z(
        npu_inst_pe_1_6_3_n29) );
  MUX2_X1 npu_inst_pe_1_6_3_U157 ( .A(npu_inst_pe_1_6_3_n28), .B(
        npu_inst_pe_1_6_3_n23), .S(npu_inst_pe_1_6_3_n8), .Z(
        npu_inst_pe_1_6_3_N94) );
  MUX2_X1 npu_inst_pe_1_6_3_U156 ( .A(npu_inst_pe_1_6_3_n25), .B(
        npu_inst_pe_1_6_3_n24), .S(npu_inst_pe_1_6_3_n6), .Z(
        npu_inst_pe_1_6_3_n28) );
  MUX2_X1 npu_inst_pe_1_6_3_U155 ( .A(npu_inst_pe_1_6_3_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_6_3_int_q_reg_v_1__1_), .S(npu_inst_pe_1_6_3_n4), .Z(
        npu_inst_pe_1_6_3_n25) );
  MUX2_X1 npu_inst_pe_1_6_3_U154 ( .A(npu_inst_pe_1_6_3_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_6_3_int_q_reg_v_3__1_), .S(npu_inst_pe_1_6_3_n4), .Z(
        npu_inst_pe_1_6_3_n24) );
  MUX2_X1 npu_inst_pe_1_6_3_U153 ( .A(npu_inst_pe_1_6_3_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_6_3_int_q_reg_v_5__1_), .S(npu_inst_pe_1_6_3_n4), .Z(
        npu_inst_pe_1_6_3_n23) );
  MUX2_X1 npu_inst_pe_1_6_3_U152 ( .A(npu_inst_pe_1_6_3_n22), .B(
        npu_inst_pe_1_6_3_n19), .S(npu_inst_pe_1_6_3_n8), .Z(
        npu_inst_int_data_x_6__3__1_) );
  MUX2_X1 npu_inst_pe_1_6_3_U151 ( .A(npu_inst_pe_1_6_3_n21), .B(
        npu_inst_pe_1_6_3_n20), .S(npu_inst_pe_1_6_3_n6), .Z(
        npu_inst_pe_1_6_3_n22) );
  MUX2_X1 npu_inst_pe_1_6_3_U150 ( .A(npu_inst_pe_1_6_3_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_6_3_int_q_reg_h_1__1_), .S(npu_inst_pe_1_6_3_n4), .Z(
        npu_inst_pe_1_6_3_n21) );
  MUX2_X1 npu_inst_pe_1_6_3_U149 ( .A(npu_inst_pe_1_6_3_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_6_3_int_q_reg_h_3__1_), .S(npu_inst_pe_1_6_3_n4), .Z(
        npu_inst_pe_1_6_3_n20) );
  MUX2_X1 npu_inst_pe_1_6_3_U148 ( .A(npu_inst_pe_1_6_3_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_6_3_int_q_reg_h_5__1_), .S(npu_inst_pe_1_6_3_n4), .Z(
        npu_inst_pe_1_6_3_n19) );
  MUX2_X1 npu_inst_pe_1_6_3_U147 ( .A(npu_inst_pe_1_6_3_n18), .B(
        npu_inst_pe_1_6_3_n15), .S(npu_inst_pe_1_6_3_n8), .Z(
        npu_inst_int_data_x_6__3__0_) );
  MUX2_X1 npu_inst_pe_1_6_3_U146 ( .A(npu_inst_pe_1_6_3_n17), .B(
        npu_inst_pe_1_6_3_n16), .S(npu_inst_pe_1_6_3_n6), .Z(
        npu_inst_pe_1_6_3_n18) );
  MUX2_X1 npu_inst_pe_1_6_3_U145 ( .A(npu_inst_pe_1_6_3_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_6_3_int_q_reg_h_1__0_), .S(npu_inst_pe_1_6_3_n4), .Z(
        npu_inst_pe_1_6_3_n17) );
  MUX2_X1 npu_inst_pe_1_6_3_U144 ( .A(npu_inst_pe_1_6_3_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_6_3_int_q_reg_h_3__0_), .S(npu_inst_pe_1_6_3_n4), .Z(
        npu_inst_pe_1_6_3_n16) );
  MUX2_X1 npu_inst_pe_1_6_3_U143 ( .A(npu_inst_pe_1_6_3_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_6_3_int_q_reg_h_5__0_), .S(npu_inst_pe_1_6_3_n4), .Z(
        npu_inst_pe_1_6_3_n15) );
  XOR2_X1 npu_inst_pe_1_6_3_U142 ( .A(npu_inst_pe_1_6_3_int_data_0_), .B(
        npu_inst_pe_1_6_3_int_q_acc_0_), .Z(npu_inst_pe_1_6_3_N73) );
  AND2_X1 npu_inst_pe_1_6_3_U141 ( .A1(npu_inst_pe_1_6_3_int_q_acc_0_), .A2(
        npu_inst_pe_1_6_3_int_data_0_), .ZN(npu_inst_pe_1_6_3_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_6_3_U140 ( .A(npu_inst_pe_1_6_3_int_q_acc_0_), .B(
        npu_inst_pe_1_6_3_n13), .ZN(npu_inst_pe_1_6_3_N65) );
  OR2_X1 npu_inst_pe_1_6_3_U139 ( .A1(npu_inst_pe_1_6_3_n13), .A2(
        npu_inst_pe_1_6_3_int_q_acc_0_), .ZN(npu_inst_pe_1_6_3_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_6_3_U138 ( .A(npu_inst_pe_1_6_3_int_q_acc_2_), .B(
        npu_inst_pe_1_6_3_add_69_carry_2_), .Z(npu_inst_pe_1_6_3_N75) );
  AND2_X1 npu_inst_pe_1_6_3_U137 ( .A1(npu_inst_pe_1_6_3_add_69_carry_2_), 
        .A2(npu_inst_pe_1_6_3_int_q_acc_2_), .ZN(
        npu_inst_pe_1_6_3_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_6_3_U136 ( .A(npu_inst_pe_1_6_3_int_q_acc_3_), .B(
        npu_inst_pe_1_6_3_add_69_carry_3_), .Z(npu_inst_pe_1_6_3_N76) );
  AND2_X1 npu_inst_pe_1_6_3_U135 ( .A1(npu_inst_pe_1_6_3_add_69_carry_3_), 
        .A2(npu_inst_pe_1_6_3_int_q_acc_3_), .ZN(
        npu_inst_pe_1_6_3_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_6_3_U134 ( .A(npu_inst_pe_1_6_3_int_q_acc_4_), .B(
        npu_inst_pe_1_6_3_add_69_carry_4_), .Z(npu_inst_pe_1_6_3_N77) );
  AND2_X1 npu_inst_pe_1_6_3_U133 ( .A1(npu_inst_pe_1_6_3_add_69_carry_4_), 
        .A2(npu_inst_pe_1_6_3_int_q_acc_4_), .ZN(
        npu_inst_pe_1_6_3_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_6_3_U132 ( .A(npu_inst_pe_1_6_3_int_q_acc_5_), .B(
        npu_inst_pe_1_6_3_add_69_carry_5_), .Z(npu_inst_pe_1_6_3_N78) );
  AND2_X1 npu_inst_pe_1_6_3_U131 ( .A1(npu_inst_pe_1_6_3_add_69_carry_5_), 
        .A2(npu_inst_pe_1_6_3_int_q_acc_5_), .ZN(
        npu_inst_pe_1_6_3_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_6_3_U130 ( .A(npu_inst_pe_1_6_3_int_q_acc_6_), .B(
        npu_inst_pe_1_6_3_add_69_carry_6_), .Z(npu_inst_pe_1_6_3_N79) );
  AND2_X1 npu_inst_pe_1_6_3_U129 ( .A1(npu_inst_pe_1_6_3_add_69_carry_6_), 
        .A2(npu_inst_pe_1_6_3_int_q_acc_6_), .ZN(
        npu_inst_pe_1_6_3_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_6_3_U128 ( .A(npu_inst_pe_1_6_3_int_q_acc_7_), .B(
        npu_inst_pe_1_6_3_add_69_carry_7_), .Z(npu_inst_pe_1_6_3_N80) );
  XNOR2_X1 npu_inst_pe_1_6_3_U127 ( .A(npu_inst_pe_1_6_3_sub_67_carry_2_), .B(
        npu_inst_pe_1_6_3_int_q_acc_2_), .ZN(npu_inst_pe_1_6_3_N67) );
  OR2_X1 npu_inst_pe_1_6_3_U126 ( .A1(npu_inst_pe_1_6_3_int_q_acc_2_), .A2(
        npu_inst_pe_1_6_3_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_6_3_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_6_3_U125 ( .A(npu_inst_pe_1_6_3_sub_67_carry_3_), .B(
        npu_inst_pe_1_6_3_int_q_acc_3_), .ZN(npu_inst_pe_1_6_3_N68) );
  OR2_X1 npu_inst_pe_1_6_3_U124 ( .A1(npu_inst_pe_1_6_3_int_q_acc_3_), .A2(
        npu_inst_pe_1_6_3_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_6_3_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_6_3_U123 ( .A(npu_inst_pe_1_6_3_sub_67_carry_4_), .B(
        npu_inst_pe_1_6_3_int_q_acc_4_), .ZN(npu_inst_pe_1_6_3_N69) );
  OR2_X1 npu_inst_pe_1_6_3_U122 ( .A1(npu_inst_pe_1_6_3_int_q_acc_4_), .A2(
        npu_inst_pe_1_6_3_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_6_3_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_6_3_U121 ( .A(npu_inst_pe_1_6_3_sub_67_carry_5_), .B(
        npu_inst_pe_1_6_3_int_q_acc_5_), .ZN(npu_inst_pe_1_6_3_N70) );
  OR2_X1 npu_inst_pe_1_6_3_U120 ( .A1(npu_inst_pe_1_6_3_int_q_acc_5_), .A2(
        npu_inst_pe_1_6_3_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_6_3_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_6_3_U119 ( .A(npu_inst_pe_1_6_3_sub_67_carry_6_), .B(
        npu_inst_pe_1_6_3_int_q_acc_6_), .ZN(npu_inst_pe_1_6_3_N71) );
  OR2_X1 npu_inst_pe_1_6_3_U118 ( .A1(npu_inst_pe_1_6_3_int_q_acc_6_), .A2(
        npu_inst_pe_1_6_3_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_6_3_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_6_3_U117 ( .A(npu_inst_pe_1_6_3_int_q_acc_7_), .B(
        npu_inst_pe_1_6_3_sub_67_carry_7_), .ZN(npu_inst_pe_1_6_3_N72) );
  INV_X1 npu_inst_pe_1_6_3_U116 ( .A(npu_inst_n76), .ZN(npu_inst_pe_1_6_3_n7)
         );
  INV_X1 npu_inst_pe_1_6_3_U115 ( .A(npu_inst_pe_1_6_3_n7), .ZN(
        npu_inst_pe_1_6_3_n6) );
  INV_X1 npu_inst_pe_1_6_3_U114 ( .A(npu_inst_n53), .ZN(npu_inst_pe_1_6_3_n3)
         );
  AOI22_X1 npu_inst_pe_1_6_3_U113 ( .A1(npu_inst_int_data_y_7__3__0_), .A2(
        npu_inst_pe_1_6_3_n58), .B1(npu_inst_pe_1_6_3_n119), .B2(
        npu_inst_pe_1_6_3_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_6_3_n57) );
  INV_X1 npu_inst_pe_1_6_3_U112 ( .A(npu_inst_pe_1_6_3_n57), .ZN(
        npu_inst_pe_1_6_3_n108) );
  AOI22_X1 npu_inst_pe_1_6_3_U111 ( .A1(npu_inst_int_data_y_7__3__0_), .A2(
        npu_inst_pe_1_6_3_n54), .B1(npu_inst_pe_1_6_3_n118), .B2(
        npu_inst_pe_1_6_3_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_6_3_n53) );
  INV_X1 npu_inst_pe_1_6_3_U110 ( .A(npu_inst_pe_1_6_3_n53), .ZN(
        npu_inst_pe_1_6_3_n109) );
  AOI22_X1 npu_inst_pe_1_6_3_U107 ( .A1(npu_inst_int_data_y_7__3__0_), .A2(
        npu_inst_pe_1_6_3_n50), .B1(npu_inst_pe_1_6_3_n117), .B2(
        npu_inst_pe_1_6_3_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_6_3_n49) );
  INV_X1 npu_inst_pe_1_6_3_U106 ( .A(npu_inst_pe_1_6_3_n49), .ZN(
        npu_inst_pe_1_6_3_n110) );
  AOI22_X1 npu_inst_pe_1_6_3_U105 ( .A1(npu_inst_int_data_y_7__3__0_), .A2(
        npu_inst_pe_1_6_3_n46), .B1(npu_inst_pe_1_6_3_n116), .B2(
        npu_inst_pe_1_6_3_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_6_3_n45) );
  INV_X1 npu_inst_pe_1_6_3_U104 ( .A(npu_inst_pe_1_6_3_n45), .ZN(
        npu_inst_pe_1_6_3_n111) );
  AOI22_X1 npu_inst_pe_1_6_3_U103 ( .A1(npu_inst_int_data_y_7__3__0_), .A2(
        npu_inst_pe_1_6_3_n42), .B1(npu_inst_pe_1_6_3_n115), .B2(
        npu_inst_pe_1_6_3_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_6_3_n41) );
  INV_X1 npu_inst_pe_1_6_3_U102 ( .A(npu_inst_pe_1_6_3_n41), .ZN(
        npu_inst_pe_1_6_3_n112) );
  AOI22_X1 npu_inst_pe_1_6_3_U101 ( .A1(npu_inst_int_data_y_7__3__1_), .A2(
        npu_inst_pe_1_6_3_n58), .B1(npu_inst_pe_1_6_3_n119), .B2(
        npu_inst_pe_1_6_3_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_6_3_n59) );
  INV_X1 npu_inst_pe_1_6_3_U100 ( .A(npu_inst_pe_1_6_3_n59), .ZN(
        npu_inst_pe_1_6_3_n102) );
  AOI22_X1 npu_inst_pe_1_6_3_U99 ( .A1(npu_inst_int_data_y_7__3__1_), .A2(
        npu_inst_pe_1_6_3_n54), .B1(npu_inst_pe_1_6_3_n118), .B2(
        npu_inst_pe_1_6_3_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_6_3_n55) );
  INV_X1 npu_inst_pe_1_6_3_U98 ( .A(npu_inst_pe_1_6_3_n55), .ZN(
        npu_inst_pe_1_6_3_n103) );
  AOI22_X1 npu_inst_pe_1_6_3_U97 ( .A1(npu_inst_int_data_y_7__3__1_), .A2(
        npu_inst_pe_1_6_3_n50), .B1(npu_inst_pe_1_6_3_n117), .B2(
        npu_inst_pe_1_6_3_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_6_3_n51) );
  INV_X1 npu_inst_pe_1_6_3_U96 ( .A(npu_inst_pe_1_6_3_n51), .ZN(
        npu_inst_pe_1_6_3_n104) );
  AOI22_X1 npu_inst_pe_1_6_3_U95 ( .A1(npu_inst_int_data_y_7__3__1_), .A2(
        npu_inst_pe_1_6_3_n46), .B1(npu_inst_pe_1_6_3_n116), .B2(
        npu_inst_pe_1_6_3_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_6_3_n47) );
  INV_X1 npu_inst_pe_1_6_3_U94 ( .A(npu_inst_pe_1_6_3_n47), .ZN(
        npu_inst_pe_1_6_3_n105) );
  AOI22_X1 npu_inst_pe_1_6_3_U93 ( .A1(npu_inst_int_data_y_7__3__1_), .A2(
        npu_inst_pe_1_6_3_n42), .B1(npu_inst_pe_1_6_3_n115), .B2(
        npu_inst_pe_1_6_3_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_6_3_n43) );
  INV_X1 npu_inst_pe_1_6_3_U92 ( .A(npu_inst_pe_1_6_3_n43), .ZN(
        npu_inst_pe_1_6_3_n106) );
  AOI22_X1 npu_inst_pe_1_6_3_U91 ( .A1(npu_inst_pe_1_6_3_n38), .A2(
        npu_inst_int_data_y_7__3__1_), .B1(npu_inst_pe_1_6_3_n114), .B2(
        npu_inst_pe_1_6_3_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_6_3_n39) );
  INV_X1 npu_inst_pe_1_6_3_U90 ( .A(npu_inst_pe_1_6_3_n39), .ZN(
        npu_inst_pe_1_6_3_n107) );
  AOI22_X1 npu_inst_pe_1_6_3_U89 ( .A1(npu_inst_pe_1_6_3_n38), .A2(
        npu_inst_int_data_y_7__3__0_), .B1(npu_inst_pe_1_6_3_n114), .B2(
        npu_inst_pe_1_6_3_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_6_3_n37) );
  INV_X1 npu_inst_pe_1_6_3_U88 ( .A(npu_inst_pe_1_6_3_n37), .ZN(
        npu_inst_pe_1_6_3_n113) );
  NAND2_X1 npu_inst_pe_1_6_3_U87 ( .A1(npu_inst_pe_1_6_3_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_6_3_n60), .ZN(npu_inst_pe_1_6_3_n74) );
  OAI21_X1 npu_inst_pe_1_6_3_U86 ( .B1(npu_inst_pe_1_6_3_n63), .B2(
        npu_inst_pe_1_6_3_n60), .A(npu_inst_pe_1_6_3_n74), .ZN(
        npu_inst_pe_1_6_3_n97) );
  NAND2_X1 npu_inst_pe_1_6_3_U85 ( .A1(npu_inst_pe_1_6_3_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_6_3_n60), .ZN(npu_inst_pe_1_6_3_n73) );
  OAI21_X1 npu_inst_pe_1_6_3_U84 ( .B1(npu_inst_pe_1_6_3_n61), .B2(
        npu_inst_pe_1_6_3_n60), .A(npu_inst_pe_1_6_3_n73), .ZN(
        npu_inst_pe_1_6_3_n96) );
  NAND2_X1 npu_inst_pe_1_6_3_U83 ( .A1(npu_inst_pe_1_6_3_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_6_3_n56), .ZN(npu_inst_pe_1_6_3_n72) );
  OAI21_X1 npu_inst_pe_1_6_3_U82 ( .B1(npu_inst_pe_1_6_3_n63), .B2(
        npu_inst_pe_1_6_3_n56), .A(npu_inst_pe_1_6_3_n72), .ZN(
        npu_inst_pe_1_6_3_n95) );
  NAND2_X1 npu_inst_pe_1_6_3_U81 ( .A1(npu_inst_pe_1_6_3_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_6_3_n56), .ZN(npu_inst_pe_1_6_3_n71) );
  OAI21_X1 npu_inst_pe_1_6_3_U80 ( .B1(npu_inst_pe_1_6_3_n61), .B2(
        npu_inst_pe_1_6_3_n56), .A(npu_inst_pe_1_6_3_n71), .ZN(
        npu_inst_pe_1_6_3_n94) );
  NAND2_X1 npu_inst_pe_1_6_3_U79 ( .A1(npu_inst_pe_1_6_3_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_6_3_n52), .ZN(npu_inst_pe_1_6_3_n70) );
  OAI21_X1 npu_inst_pe_1_6_3_U78 ( .B1(npu_inst_pe_1_6_3_n63), .B2(
        npu_inst_pe_1_6_3_n52), .A(npu_inst_pe_1_6_3_n70), .ZN(
        npu_inst_pe_1_6_3_n93) );
  NAND2_X1 npu_inst_pe_1_6_3_U77 ( .A1(npu_inst_pe_1_6_3_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_6_3_n52), .ZN(npu_inst_pe_1_6_3_n69) );
  OAI21_X1 npu_inst_pe_1_6_3_U76 ( .B1(npu_inst_pe_1_6_3_n61), .B2(
        npu_inst_pe_1_6_3_n52), .A(npu_inst_pe_1_6_3_n69), .ZN(
        npu_inst_pe_1_6_3_n92) );
  NAND2_X1 npu_inst_pe_1_6_3_U75 ( .A1(npu_inst_pe_1_6_3_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_6_3_n48), .ZN(npu_inst_pe_1_6_3_n68) );
  OAI21_X1 npu_inst_pe_1_6_3_U74 ( .B1(npu_inst_pe_1_6_3_n63), .B2(
        npu_inst_pe_1_6_3_n48), .A(npu_inst_pe_1_6_3_n68), .ZN(
        npu_inst_pe_1_6_3_n91) );
  NAND2_X1 npu_inst_pe_1_6_3_U73 ( .A1(npu_inst_pe_1_6_3_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_6_3_n48), .ZN(npu_inst_pe_1_6_3_n67) );
  OAI21_X1 npu_inst_pe_1_6_3_U72 ( .B1(npu_inst_pe_1_6_3_n61), .B2(
        npu_inst_pe_1_6_3_n48), .A(npu_inst_pe_1_6_3_n67), .ZN(
        npu_inst_pe_1_6_3_n90) );
  NAND2_X1 npu_inst_pe_1_6_3_U71 ( .A1(npu_inst_pe_1_6_3_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_6_3_n44), .ZN(npu_inst_pe_1_6_3_n66) );
  OAI21_X1 npu_inst_pe_1_6_3_U70 ( .B1(npu_inst_pe_1_6_3_n63), .B2(
        npu_inst_pe_1_6_3_n44), .A(npu_inst_pe_1_6_3_n66), .ZN(
        npu_inst_pe_1_6_3_n89) );
  NAND2_X1 npu_inst_pe_1_6_3_U69 ( .A1(npu_inst_pe_1_6_3_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_6_3_n44), .ZN(npu_inst_pe_1_6_3_n65) );
  OAI21_X1 npu_inst_pe_1_6_3_U68 ( .B1(npu_inst_pe_1_6_3_n61), .B2(
        npu_inst_pe_1_6_3_n44), .A(npu_inst_pe_1_6_3_n65), .ZN(
        npu_inst_pe_1_6_3_n88) );
  NAND2_X1 npu_inst_pe_1_6_3_U67 ( .A1(npu_inst_pe_1_6_3_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_6_3_n40), .ZN(npu_inst_pe_1_6_3_n64) );
  OAI21_X1 npu_inst_pe_1_6_3_U66 ( .B1(npu_inst_pe_1_6_3_n63), .B2(
        npu_inst_pe_1_6_3_n40), .A(npu_inst_pe_1_6_3_n64), .ZN(
        npu_inst_pe_1_6_3_n87) );
  NAND2_X1 npu_inst_pe_1_6_3_U65 ( .A1(npu_inst_pe_1_6_3_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_6_3_n40), .ZN(npu_inst_pe_1_6_3_n62) );
  OAI21_X1 npu_inst_pe_1_6_3_U64 ( .B1(npu_inst_pe_1_6_3_n61), .B2(
        npu_inst_pe_1_6_3_n40), .A(npu_inst_pe_1_6_3_n62), .ZN(
        npu_inst_pe_1_6_3_n86) );
  AND2_X1 npu_inst_pe_1_6_3_U63 ( .A1(npu_inst_pe_1_6_3_N93), .A2(npu_inst_n53), .ZN(npu_inst_int_data_y_6__3__0_) );
  AND2_X1 npu_inst_pe_1_6_3_U62 ( .A1(npu_inst_n53), .A2(npu_inst_pe_1_6_3_N94), .ZN(npu_inst_int_data_y_6__3__1_) );
  NOR3_X1 npu_inst_pe_1_6_3_U61 ( .A1(npu_inst_pe_1_6_3_n26), .A2(npu_inst_n53), .A3(npu_inst_int_ckg[12]), .ZN(npu_inst_pe_1_6_3_n85) );
  OR2_X1 npu_inst_pe_1_6_3_U60 ( .A1(npu_inst_pe_1_6_3_n85), .A2(
        npu_inst_pe_1_6_3_n2), .ZN(npu_inst_pe_1_6_3_N84) );
  AND2_X1 npu_inst_pe_1_6_3_U59 ( .A1(npu_inst_pe_1_6_3_int_q_acc_0_), .A2(
        npu_inst_pe_1_6_3_n1), .ZN(npu_inst_int_data_res_6__3__0_) );
  AND2_X1 npu_inst_pe_1_6_3_U58 ( .A1(npu_inst_pe_1_6_3_n2), .A2(
        npu_inst_pe_1_6_3_int_q_acc_7_), .ZN(npu_inst_int_data_res_6__3__7_)
         );
  AND2_X1 npu_inst_pe_1_6_3_U57 ( .A1(npu_inst_pe_1_6_3_int_q_acc_1_), .A2(
        npu_inst_pe_1_6_3_n1), .ZN(npu_inst_int_data_res_6__3__1_) );
  AND2_X1 npu_inst_pe_1_6_3_U56 ( .A1(npu_inst_pe_1_6_3_int_q_acc_2_), .A2(
        npu_inst_pe_1_6_3_n1), .ZN(npu_inst_int_data_res_6__3__2_) );
  AND2_X1 npu_inst_pe_1_6_3_U55 ( .A1(npu_inst_pe_1_6_3_int_q_acc_3_), .A2(
        npu_inst_pe_1_6_3_n2), .ZN(npu_inst_int_data_res_6__3__3_) );
  AND2_X1 npu_inst_pe_1_6_3_U54 ( .A1(npu_inst_pe_1_6_3_int_q_acc_4_), .A2(
        npu_inst_pe_1_6_3_n2), .ZN(npu_inst_int_data_res_6__3__4_) );
  AND2_X1 npu_inst_pe_1_6_3_U53 ( .A1(npu_inst_pe_1_6_3_int_q_acc_5_), .A2(
        npu_inst_pe_1_6_3_n2), .ZN(npu_inst_int_data_res_6__3__5_) );
  AND2_X1 npu_inst_pe_1_6_3_U52 ( .A1(npu_inst_pe_1_6_3_int_q_acc_6_), .A2(
        npu_inst_pe_1_6_3_n2), .ZN(npu_inst_int_data_res_6__3__6_) );
  AOI222_X1 npu_inst_pe_1_6_3_U51 ( .A1(npu_inst_int_data_res_7__3__0_), .A2(
        npu_inst_pe_1_6_3_n1), .B1(npu_inst_pe_1_6_3_N73), .B2(
        npu_inst_pe_1_6_3_n76), .C1(npu_inst_pe_1_6_3_N65), .C2(
        npu_inst_pe_1_6_3_n77), .ZN(npu_inst_pe_1_6_3_n84) );
  INV_X1 npu_inst_pe_1_6_3_U50 ( .A(npu_inst_pe_1_6_3_n84), .ZN(
        npu_inst_pe_1_6_3_n101) );
  AOI222_X1 npu_inst_pe_1_6_3_U49 ( .A1(npu_inst_int_data_res_7__3__7_), .A2(
        npu_inst_pe_1_6_3_n1), .B1(npu_inst_pe_1_6_3_N80), .B2(
        npu_inst_pe_1_6_3_n76), .C1(npu_inst_pe_1_6_3_N72), .C2(
        npu_inst_pe_1_6_3_n77), .ZN(npu_inst_pe_1_6_3_n75) );
  INV_X1 npu_inst_pe_1_6_3_U48 ( .A(npu_inst_pe_1_6_3_n75), .ZN(
        npu_inst_pe_1_6_3_n33) );
  AOI222_X1 npu_inst_pe_1_6_3_U47 ( .A1(npu_inst_int_data_res_7__3__1_), .A2(
        npu_inst_pe_1_6_3_n1), .B1(npu_inst_pe_1_6_3_N74), .B2(
        npu_inst_pe_1_6_3_n76), .C1(npu_inst_pe_1_6_3_N66), .C2(
        npu_inst_pe_1_6_3_n77), .ZN(npu_inst_pe_1_6_3_n83) );
  INV_X1 npu_inst_pe_1_6_3_U46 ( .A(npu_inst_pe_1_6_3_n83), .ZN(
        npu_inst_pe_1_6_3_n100) );
  AOI222_X1 npu_inst_pe_1_6_3_U45 ( .A1(npu_inst_int_data_res_7__3__2_), .A2(
        npu_inst_pe_1_6_3_n1), .B1(npu_inst_pe_1_6_3_N75), .B2(
        npu_inst_pe_1_6_3_n76), .C1(npu_inst_pe_1_6_3_N67), .C2(
        npu_inst_pe_1_6_3_n77), .ZN(npu_inst_pe_1_6_3_n82) );
  INV_X1 npu_inst_pe_1_6_3_U44 ( .A(npu_inst_pe_1_6_3_n82), .ZN(
        npu_inst_pe_1_6_3_n99) );
  AOI222_X1 npu_inst_pe_1_6_3_U43 ( .A1(npu_inst_int_data_res_7__3__3_), .A2(
        npu_inst_pe_1_6_3_n1), .B1(npu_inst_pe_1_6_3_N76), .B2(
        npu_inst_pe_1_6_3_n76), .C1(npu_inst_pe_1_6_3_N68), .C2(
        npu_inst_pe_1_6_3_n77), .ZN(npu_inst_pe_1_6_3_n81) );
  INV_X1 npu_inst_pe_1_6_3_U42 ( .A(npu_inst_pe_1_6_3_n81), .ZN(
        npu_inst_pe_1_6_3_n98) );
  AOI222_X1 npu_inst_pe_1_6_3_U41 ( .A1(npu_inst_int_data_res_7__3__4_), .A2(
        npu_inst_pe_1_6_3_n1), .B1(npu_inst_pe_1_6_3_N77), .B2(
        npu_inst_pe_1_6_3_n76), .C1(npu_inst_pe_1_6_3_N69), .C2(
        npu_inst_pe_1_6_3_n77), .ZN(npu_inst_pe_1_6_3_n80) );
  INV_X1 npu_inst_pe_1_6_3_U40 ( .A(npu_inst_pe_1_6_3_n80), .ZN(
        npu_inst_pe_1_6_3_n36) );
  AOI222_X1 npu_inst_pe_1_6_3_U39 ( .A1(npu_inst_int_data_res_7__3__5_), .A2(
        npu_inst_pe_1_6_3_n1), .B1(npu_inst_pe_1_6_3_N78), .B2(
        npu_inst_pe_1_6_3_n76), .C1(npu_inst_pe_1_6_3_N70), .C2(
        npu_inst_pe_1_6_3_n77), .ZN(npu_inst_pe_1_6_3_n79) );
  INV_X1 npu_inst_pe_1_6_3_U38 ( .A(npu_inst_pe_1_6_3_n79), .ZN(
        npu_inst_pe_1_6_3_n35) );
  AOI222_X1 npu_inst_pe_1_6_3_U37 ( .A1(npu_inst_int_data_res_7__3__6_), .A2(
        npu_inst_pe_1_6_3_n1), .B1(npu_inst_pe_1_6_3_N79), .B2(
        npu_inst_pe_1_6_3_n76), .C1(npu_inst_pe_1_6_3_N71), .C2(
        npu_inst_pe_1_6_3_n77), .ZN(npu_inst_pe_1_6_3_n78) );
  INV_X1 npu_inst_pe_1_6_3_U36 ( .A(npu_inst_pe_1_6_3_n78), .ZN(
        npu_inst_pe_1_6_3_n34) );
  INV_X1 npu_inst_pe_1_6_3_U35 ( .A(npu_inst_pe_1_6_3_int_data_1_), .ZN(
        npu_inst_pe_1_6_3_n14) );
  AND2_X1 npu_inst_pe_1_6_3_U34 ( .A1(npu_inst_int_data_x_6__3__1_), .A2(
        npu_inst_pe_1_6_3_int_q_weight_1_), .ZN(npu_inst_pe_1_6_3_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_6_3_U33 ( .A1(npu_inst_int_data_x_6__3__0_), .A2(
        npu_inst_pe_1_6_3_int_q_weight_1_), .ZN(npu_inst_pe_1_6_3_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_6_3_U32 ( .A1(npu_inst_n53), .A2(
        npu_inst_int_data_y_7__3__1_), .B1(npu_inst_pe_1_6_3_n3), .B2(
        npu_inst_int_data_x_6__4__1_), .ZN(npu_inst_pe_1_6_3_n63) );
  AOI22_X1 npu_inst_pe_1_6_3_U31 ( .A1(npu_inst_n53), .A2(
        npu_inst_int_data_y_7__3__0_), .B1(npu_inst_pe_1_6_3_n3), .B2(
        npu_inst_int_data_x_6__4__0_), .ZN(npu_inst_pe_1_6_3_n61) );
  INV_X1 npu_inst_pe_1_6_3_U30 ( .A(npu_inst_pe_1_6_3_int_data_0_), .ZN(
        npu_inst_pe_1_6_3_n13) );
  INV_X1 npu_inst_pe_1_6_3_U29 ( .A(npu_inst_n68), .ZN(npu_inst_pe_1_6_3_n5)
         );
  OR3_X1 npu_inst_pe_1_6_3_U28 ( .A1(npu_inst_pe_1_6_3_n6), .A2(
        npu_inst_pe_1_6_3_n8), .A3(npu_inst_pe_1_6_3_n5), .ZN(
        npu_inst_pe_1_6_3_n56) );
  OR3_X1 npu_inst_pe_1_6_3_U27 ( .A1(npu_inst_pe_1_6_3_n5), .A2(
        npu_inst_pe_1_6_3_n8), .A3(npu_inst_pe_1_6_3_n7), .ZN(
        npu_inst_pe_1_6_3_n48) );
  INV_X1 npu_inst_pe_1_6_3_U26 ( .A(npu_inst_pe_1_6_3_n5), .ZN(
        npu_inst_pe_1_6_3_n4) );
  OR3_X1 npu_inst_pe_1_6_3_U25 ( .A1(npu_inst_pe_1_6_3_n4), .A2(
        npu_inst_pe_1_6_3_n8), .A3(npu_inst_pe_1_6_3_n7), .ZN(
        npu_inst_pe_1_6_3_n52) );
  OR3_X1 npu_inst_pe_1_6_3_U24 ( .A1(npu_inst_pe_1_6_3_n6), .A2(
        npu_inst_pe_1_6_3_n8), .A3(npu_inst_pe_1_6_3_n4), .ZN(
        npu_inst_pe_1_6_3_n60) );
  NOR2_X1 npu_inst_pe_1_6_3_U23 ( .A1(npu_inst_pe_1_6_3_n60), .A2(
        npu_inst_pe_1_6_3_n3), .ZN(npu_inst_pe_1_6_3_n58) );
  NOR2_X1 npu_inst_pe_1_6_3_U22 ( .A1(npu_inst_pe_1_6_3_n56), .A2(
        npu_inst_pe_1_6_3_n3), .ZN(npu_inst_pe_1_6_3_n54) );
  NOR2_X1 npu_inst_pe_1_6_3_U21 ( .A1(npu_inst_pe_1_6_3_n52), .A2(
        npu_inst_pe_1_6_3_n3), .ZN(npu_inst_pe_1_6_3_n50) );
  NOR2_X1 npu_inst_pe_1_6_3_U20 ( .A1(npu_inst_pe_1_6_3_n48), .A2(
        npu_inst_pe_1_6_3_n3), .ZN(npu_inst_pe_1_6_3_n46) );
  NOR2_X1 npu_inst_pe_1_6_3_U19 ( .A1(npu_inst_pe_1_6_3_n40), .A2(
        npu_inst_pe_1_6_3_n3), .ZN(npu_inst_pe_1_6_3_n38) );
  NOR2_X1 npu_inst_pe_1_6_3_U18 ( .A1(npu_inst_pe_1_6_3_n44), .A2(
        npu_inst_pe_1_6_3_n3), .ZN(npu_inst_pe_1_6_3_n42) );
  BUF_X1 npu_inst_pe_1_6_3_U17 ( .A(npu_inst_n95), .Z(npu_inst_pe_1_6_3_n8) );
  INV_X1 npu_inst_pe_1_6_3_U16 ( .A(npu_inst_n123), .ZN(npu_inst_pe_1_6_3_n12)
         );
  INV_X1 npu_inst_pe_1_6_3_U15 ( .A(npu_inst_pe_1_6_3_n38), .ZN(
        npu_inst_pe_1_6_3_n114) );
  INV_X1 npu_inst_pe_1_6_3_U14 ( .A(npu_inst_pe_1_6_3_n58), .ZN(
        npu_inst_pe_1_6_3_n119) );
  INV_X1 npu_inst_pe_1_6_3_U13 ( .A(npu_inst_pe_1_6_3_n54), .ZN(
        npu_inst_pe_1_6_3_n118) );
  INV_X1 npu_inst_pe_1_6_3_U12 ( .A(npu_inst_pe_1_6_3_n50), .ZN(
        npu_inst_pe_1_6_3_n117) );
  INV_X1 npu_inst_pe_1_6_3_U11 ( .A(npu_inst_pe_1_6_3_n46), .ZN(
        npu_inst_pe_1_6_3_n116) );
  INV_X1 npu_inst_pe_1_6_3_U10 ( .A(npu_inst_pe_1_6_3_n42), .ZN(
        npu_inst_pe_1_6_3_n115) );
  BUF_X1 npu_inst_pe_1_6_3_U9 ( .A(npu_inst_n13), .Z(npu_inst_pe_1_6_3_n2) );
  BUF_X1 npu_inst_pe_1_6_3_U8 ( .A(npu_inst_n13), .Z(npu_inst_pe_1_6_3_n1) );
  BUF_X1 npu_inst_pe_1_6_3_U7 ( .A(npu_inst_pe_1_6_3_n12), .Z(
        npu_inst_pe_1_6_3_n11) );
  BUF_X1 npu_inst_pe_1_6_3_U6 ( .A(npu_inst_pe_1_6_3_n12), .Z(
        npu_inst_pe_1_6_3_n10) );
  BUF_X1 npu_inst_pe_1_6_3_U5 ( .A(npu_inst_pe_1_6_3_n12), .Z(
        npu_inst_pe_1_6_3_n9) );
  NOR2_X1 npu_inst_pe_1_6_3_U4 ( .A1(npu_inst_pe_1_6_3_int_q_weight_0_), .A2(
        npu_inst_pe_1_6_3_n1), .ZN(npu_inst_pe_1_6_3_n76) );
  NOR2_X1 npu_inst_pe_1_6_3_U3 ( .A1(npu_inst_pe_1_6_3_n27), .A2(
        npu_inst_pe_1_6_3_n1), .ZN(npu_inst_pe_1_6_3_n77) );
  FA_X1 npu_inst_pe_1_6_3_sub_67_U2_1 ( .A(npu_inst_pe_1_6_3_int_q_acc_1_), 
        .B(npu_inst_pe_1_6_3_n14), .CI(npu_inst_pe_1_6_3_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_6_3_sub_67_carry_2_), .S(npu_inst_pe_1_6_3_N66) );
  FA_X1 npu_inst_pe_1_6_3_add_69_U1_1 ( .A(npu_inst_pe_1_6_3_int_q_acc_1_), 
        .B(npu_inst_pe_1_6_3_int_data_1_), .CI(
        npu_inst_pe_1_6_3_add_69_carry_1_), .CO(
        npu_inst_pe_1_6_3_add_69_carry_2_), .S(npu_inst_pe_1_6_3_N74) );
  NAND3_X1 npu_inst_pe_1_6_3_U109 ( .A1(npu_inst_pe_1_6_3_n5), .A2(
        npu_inst_pe_1_6_3_n7), .A3(npu_inst_pe_1_6_3_n8), .ZN(
        npu_inst_pe_1_6_3_n44) );
  NAND3_X1 npu_inst_pe_1_6_3_U108 ( .A1(npu_inst_pe_1_6_3_n4), .A2(
        npu_inst_pe_1_6_3_n7), .A3(npu_inst_pe_1_6_3_n8), .ZN(
        npu_inst_pe_1_6_3_n40) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_6_3_n34), .CK(
        npu_inst_pe_1_6_3_net3389), .RN(npu_inst_pe_1_6_3_n9), .Q(
        npu_inst_pe_1_6_3_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_6_3_n35), .CK(
        npu_inst_pe_1_6_3_net3389), .RN(npu_inst_pe_1_6_3_n9), .Q(
        npu_inst_pe_1_6_3_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_6_3_n36), .CK(
        npu_inst_pe_1_6_3_net3389), .RN(npu_inst_pe_1_6_3_n9), .Q(
        npu_inst_pe_1_6_3_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_6_3_n98), .CK(
        npu_inst_pe_1_6_3_net3389), .RN(npu_inst_pe_1_6_3_n9), .Q(
        npu_inst_pe_1_6_3_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_6_3_n99), .CK(
        npu_inst_pe_1_6_3_net3389), .RN(npu_inst_pe_1_6_3_n9), .Q(
        npu_inst_pe_1_6_3_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_6_3_n100), 
        .CK(npu_inst_pe_1_6_3_net3389), .RN(npu_inst_pe_1_6_3_n9), .Q(
        npu_inst_pe_1_6_3_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_6_3_n33), .CK(
        npu_inst_pe_1_6_3_net3389), .RN(npu_inst_pe_1_6_3_n9), .Q(
        npu_inst_pe_1_6_3_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_6_3_n101), 
        .CK(npu_inst_pe_1_6_3_net3389), .RN(npu_inst_pe_1_6_3_n9), .Q(
        npu_inst_pe_1_6_3_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_weight_reg_0_ ( .D(npu_inst_n109), .CK(
        npu_inst_pe_1_6_3_net3395), .RN(npu_inst_pe_1_6_3_n9), .Q(
        npu_inst_pe_1_6_3_int_q_weight_0_), .QN(npu_inst_pe_1_6_3_n27) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_weight_reg_1_ ( .D(npu_inst_n115), .CK(
        npu_inst_pe_1_6_3_net3395), .RN(npu_inst_pe_1_6_3_n9), .Q(
        npu_inst_pe_1_6_3_int_q_weight_1_), .QN(npu_inst_pe_1_6_3_n26) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_6_3_n113), 
        .CK(npu_inst_pe_1_6_3_net3395), .RN(npu_inst_pe_1_6_3_n9), .Q(
        npu_inst_pe_1_6_3_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_6_3_n107), 
        .CK(npu_inst_pe_1_6_3_net3395), .RN(npu_inst_pe_1_6_3_n9), .Q(
        npu_inst_pe_1_6_3_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_6_3_n112), 
        .CK(npu_inst_pe_1_6_3_net3395), .RN(npu_inst_pe_1_6_3_n10), .Q(
        npu_inst_pe_1_6_3_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_6_3_n106), 
        .CK(npu_inst_pe_1_6_3_net3395), .RN(npu_inst_pe_1_6_3_n10), .Q(
        npu_inst_pe_1_6_3_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_6_3_n111), 
        .CK(npu_inst_pe_1_6_3_net3395), .RN(npu_inst_pe_1_6_3_n10), .Q(
        npu_inst_pe_1_6_3_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_6_3_n105), 
        .CK(npu_inst_pe_1_6_3_net3395), .RN(npu_inst_pe_1_6_3_n10), .Q(
        npu_inst_pe_1_6_3_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_6_3_n110), 
        .CK(npu_inst_pe_1_6_3_net3395), .RN(npu_inst_pe_1_6_3_n10), .Q(
        npu_inst_pe_1_6_3_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_6_3_n104), 
        .CK(npu_inst_pe_1_6_3_net3395), .RN(npu_inst_pe_1_6_3_n10), .Q(
        npu_inst_pe_1_6_3_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_6_3_n109), 
        .CK(npu_inst_pe_1_6_3_net3395), .RN(npu_inst_pe_1_6_3_n10), .Q(
        npu_inst_pe_1_6_3_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_6_3_n103), 
        .CK(npu_inst_pe_1_6_3_net3395), .RN(npu_inst_pe_1_6_3_n10), .Q(
        npu_inst_pe_1_6_3_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_6_3_n108), 
        .CK(npu_inst_pe_1_6_3_net3395), .RN(npu_inst_pe_1_6_3_n10), .Q(
        npu_inst_pe_1_6_3_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_6_3_n102), 
        .CK(npu_inst_pe_1_6_3_net3395), .RN(npu_inst_pe_1_6_3_n10), .Q(
        npu_inst_pe_1_6_3_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_6_3_n86), 
        .CK(npu_inst_pe_1_6_3_net3395), .RN(npu_inst_pe_1_6_3_n10), .Q(
        npu_inst_pe_1_6_3_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_6_3_n87), 
        .CK(npu_inst_pe_1_6_3_net3395), .RN(npu_inst_pe_1_6_3_n10), .Q(
        npu_inst_pe_1_6_3_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_6_3_n88), 
        .CK(npu_inst_pe_1_6_3_net3395), .RN(npu_inst_pe_1_6_3_n11), .Q(
        npu_inst_pe_1_6_3_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_6_3_n89), 
        .CK(npu_inst_pe_1_6_3_net3395), .RN(npu_inst_pe_1_6_3_n11), .Q(
        npu_inst_pe_1_6_3_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_6_3_n90), 
        .CK(npu_inst_pe_1_6_3_net3395), .RN(npu_inst_pe_1_6_3_n11), .Q(
        npu_inst_pe_1_6_3_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_6_3_n91), 
        .CK(npu_inst_pe_1_6_3_net3395), .RN(npu_inst_pe_1_6_3_n11), .Q(
        npu_inst_pe_1_6_3_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_6_3_n92), 
        .CK(npu_inst_pe_1_6_3_net3395), .RN(npu_inst_pe_1_6_3_n11), .Q(
        npu_inst_pe_1_6_3_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_6_3_n93), 
        .CK(npu_inst_pe_1_6_3_net3395), .RN(npu_inst_pe_1_6_3_n11), .Q(
        npu_inst_pe_1_6_3_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_6_3_n94), 
        .CK(npu_inst_pe_1_6_3_net3395), .RN(npu_inst_pe_1_6_3_n11), .Q(
        npu_inst_pe_1_6_3_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_6_3_n95), 
        .CK(npu_inst_pe_1_6_3_net3395), .RN(npu_inst_pe_1_6_3_n11), .Q(
        npu_inst_pe_1_6_3_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_6_3_n96), 
        .CK(npu_inst_pe_1_6_3_net3395), .RN(npu_inst_pe_1_6_3_n11), .Q(
        npu_inst_pe_1_6_3_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_6_3_n97), 
        .CK(npu_inst_pe_1_6_3_net3395), .RN(npu_inst_pe_1_6_3_n11), .Q(
        npu_inst_pe_1_6_3_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_6_3_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_6_3_N84), .SE(1'b0), .GCK(npu_inst_pe_1_6_3_net3389) );
  CLKGATETST_X1 npu_inst_pe_1_6_3_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n62), .SE(1'b0), .GCK(npu_inst_pe_1_6_3_net3395) );
  MUX2_X1 npu_inst_pe_1_6_4_U161 ( .A(npu_inst_pe_1_6_4_n31), .B(
        npu_inst_pe_1_6_4_n28), .S(npu_inst_pe_1_6_4_n7), .Z(
        npu_inst_pe_1_6_4_N93) );
  MUX2_X1 npu_inst_pe_1_6_4_U160 ( .A(npu_inst_pe_1_6_4_n30), .B(
        npu_inst_pe_1_6_4_n29), .S(npu_inst_n75), .Z(npu_inst_pe_1_6_4_n31) );
  MUX2_X1 npu_inst_pe_1_6_4_U159 ( .A(npu_inst_pe_1_6_4_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_6_4_int_q_reg_v_1__0_), .S(npu_inst_pe_1_6_4_n4), .Z(
        npu_inst_pe_1_6_4_n30) );
  MUX2_X1 npu_inst_pe_1_6_4_U158 ( .A(npu_inst_pe_1_6_4_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_6_4_int_q_reg_v_3__0_), .S(npu_inst_pe_1_6_4_n4), .Z(
        npu_inst_pe_1_6_4_n29) );
  MUX2_X1 npu_inst_pe_1_6_4_U157 ( .A(npu_inst_pe_1_6_4_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_6_4_int_q_reg_v_5__0_), .S(npu_inst_pe_1_6_4_n4), .Z(
        npu_inst_pe_1_6_4_n28) );
  MUX2_X1 npu_inst_pe_1_6_4_U156 ( .A(npu_inst_pe_1_6_4_n25), .B(
        npu_inst_pe_1_6_4_n22), .S(npu_inst_pe_1_6_4_n7), .Z(
        npu_inst_pe_1_6_4_N94) );
  MUX2_X1 npu_inst_pe_1_6_4_U155 ( .A(npu_inst_pe_1_6_4_n24), .B(
        npu_inst_pe_1_6_4_n23), .S(npu_inst_n75), .Z(npu_inst_pe_1_6_4_n25) );
  MUX2_X1 npu_inst_pe_1_6_4_U154 ( .A(npu_inst_pe_1_6_4_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_6_4_int_q_reg_v_1__1_), .S(npu_inst_pe_1_6_4_n4), .Z(
        npu_inst_pe_1_6_4_n24) );
  MUX2_X1 npu_inst_pe_1_6_4_U153 ( .A(npu_inst_pe_1_6_4_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_6_4_int_q_reg_v_3__1_), .S(npu_inst_pe_1_6_4_n4), .Z(
        npu_inst_pe_1_6_4_n23) );
  MUX2_X1 npu_inst_pe_1_6_4_U152 ( .A(npu_inst_pe_1_6_4_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_6_4_int_q_reg_v_5__1_), .S(npu_inst_pe_1_6_4_n4), .Z(
        npu_inst_pe_1_6_4_n22) );
  MUX2_X1 npu_inst_pe_1_6_4_U151 ( .A(npu_inst_pe_1_6_4_n21), .B(
        npu_inst_pe_1_6_4_n18), .S(npu_inst_pe_1_6_4_n7), .Z(
        npu_inst_int_data_x_6__4__1_) );
  MUX2_X1 npu_inst_pe_1_6_4_U150 ( .A(npu_inst_pe_1_6_4_n20), .B(
        npu_inst_pe_1_6_4_n19), .S(npu_inst_n75), .Z(npu_inst_pe_1_6_4_n21) );
  MUX2_X1 npu_inst_pe_1_6_4_U149 ( .A(npu_inst_pe_1_6_4_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_6_4_int_q_reg_h_1__1_), .S(npu_inst_pe_1_6_4_n4), .Z(
        npu_inst_pe_1_6_4_n20) );
  MUX2_X1 npu_inst_pe_1_6_4_U148 ( .A(npu_inst_pe_1_6_4_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_6_4_int_q_reg_h_3__1_), .S(npu_inst_pe_1_6_4_n4), .Z(
        npu_inst_pe_1_6_4_n19) );
  MUX2_X1 npu_inst_pe_1_6_4_U147 ( .A(npu_inst_pe_1_6_4_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_6_4_int_q_reg_h_5__1_), .S(npu_inst_pe_1_6_4_n4), .Z(
        npu_inst_pe_1_6_4_n18) );
  MUX2_X1 npu_inst_pe_1_6_4_U146 ( .A(npu_inst_pe_1_6_4_n17), .B(
        npu_inst_pe_1_6_4_n14), .S(npu_inst_pe_1_6_4_n7), .Z(
        npu_inst_int_data_x_6__4__0_) );
  MUX2_X1 npu_inst_pe_1_6_4_U145 ( .A(npu_inst_pe_1_6_4_n16), .B(
        npu_inst_pe_1_6_4_n15), .S(npu_inst_n75), .Z(npu_inst_pe_1_6_4_n17) );
  MUX2_X1 npu_inst_pe_1_6_4_U144 ( .A(npu_inst_pe_1_6_4_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_6_4_int_q_reg_h_1__0_), .S(npu_inst_pe_1_6_4_n4), .Z(
        npu_inst_pe_1_6_4_n16) );
  MUX2_X1 npu_inst_pe_1_6_4_U143 ( .A(npu_inst_pe_1_6_4_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_6_4_int_q_reg_h_3__0_), .S(npu_inst_pe_1_6_4_n4), .Z(
        npu_inst_pe_1_6_4_n15) );
  MUX2_X1 npu_inst_pe_1_6_4_U142 ( .A(npu_inst_pe_1_6_4_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_6_4_int_q_reg_h_5__0_), .S(npu_inst_pe_1_6_4_n4), .Z(
        npu_inst_pe_1_6_4_n14) );
  XOR2_X1 npu_inst_pe_1_6_4_U141 ( .A(npu_inst_pe_1_6_4_int_data_0_), .B(
        npu_inst_pe_1_6_4_int_q_acc_0_), .Z(npu_inst_pe_1_6_4_N73) );
  AND2_X1 npu_inst_pe_1_6_4_U140 ( .A1(npu_inst_pe_1_6_4_int_q_acc_0_), .A2(
        npu_inst_pe_1_6_4_int_data_0_), .ZN(npu_inst_pe_1_6_4_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_6_4_U139 ( .A(npu_inst_pe_1_6_4_int_q_acc_0_), .B(
        npu_inst_pe_1_6_4_n12), .ZN(npu_inst_pe_1_6_4_N65) );
  OR2_X1 npu_inst_pe_1_6_4_U138 ( .A1(npu_inst_pe_1_6_4_n12), .A2(
        npu_inst_pe_1_6_4_int_q_acc_0_), .ZN(npu_inst_pe_1_6_4_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_6_4_U137 ( .A(npu_inst_pe_1_6_4_int_q_acc_2_), .B(
        npu_inst_pe_1_6_4_add_69_carry_2_), .Z(npu_inst_pe_1_6_4_N75) );
  AND2_X1 npu_inst_pe_1_6_4_U136 ( .A1(npu_inst_pe_1_6_4_add_69_carry_2_), 
        .A2(npu_inst_pe_1_6_4_int_q_acc_2_), .ZN(
        npu_inst_pe_1_6_4_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_6_4_U135 ( .A(npu_inst_pe_1_6_4_int_q_acc_3_), .B(
        npu_inst_pe_1_6_4_add_69_carry_3_), .Z(npu_inst_pe_1_6_4_N76) );
  AND2_X1 npu_inst_pe_1_6_4_U134 ( .A1(npu_inst_pe_1_6_4_add_69_carry_3_), 
        .A2(npu_inst_pe_1_6_4_int_q_acc_3_), .ZN(
        npu_inst_pe_1_6_4_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_6_4_U133 ( .A(npu_inst_pe_1_6_4_int_q_acc_4_), .B(
        npu_inst_pe_1_6_4_add_69_carry_4_), .Z(npu_inst_pe_1_6_4_N77) );
  AND2_X1 npu_inst_pe_1_6_4_U132 ( .A1(npu_inst_pe_1_6_4_add_69_carry_4_), 
        .A2(npu_inst_pe_1_6_4_int_q_acc_4_), .ZN(
        npu_inst_pe_1_6_4_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_6_4_U131 ( .A(npu_inst_pe_1_6_4_int_q_acc_5_), .B(
        npu_inst_pe_1_6_4_add_69_carry_5_), .Z(npu_inst_pe_1_6_4_N78) );
  AND2_X1 npu_inst_pe_1_6_4_U130 ( .A1(npu_inst_pe_1_6_4_add_69_carry_5_), 
        .A2(npu_inst_pe_1_6_4_int_q_acc_5_), .ZN(
        npu_inst_pe_1_6_4_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_6_4_U129 ( .A(npu_inst_pe_1_6_4_int_q_acc_6_), .B(
        npu_inst_pe_1_6_4_add_69_carry_6_), .Z(npu_inst_pe_1_6_4_N79) );
  AND2_X1 npu_inst_pe_1_6_4_U128 ( .A1(npu_inst_pe_1_6_4_add_69_carry_6_), 
        .A2(npu_inst_pe_1_6_4_int_q_acc_6_), .ZN(
        npu_inst_pe_1_6_4_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_6_4_U127 ( .A(npu_inst_pe_1_6_4_int_q_acc_7_), .B(
        npu_inst_pe_1_6_4_add_69_carry_7_), .Z(npu_inst_pe_1_6_4_N80) );
  XNOR2_X1 npu_inst_pe_1_6_4_U126 ( .A(npu_inst_pe_1_6_4_sub_67_carry_2_), .B(
        npu_inst_pe_1_6_4_int_q_acc_2_), .ZN(npu_inst_pe_1_6_4_N67) );
  OR2_X1 npu_inst_pe_1_6_4_U125 ( .A1(npu_inst_pe_1_6_4_int_q_acc_2_), .A2(
        npu_inst_pe_1_6_4_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_6_4_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_6_4_U124 ( .A(npu_inst_pe_1_6_4_sub_67_carry_3_), .B(
        npu_inst_pe_1_6_4_int_q_acc_3_), .ZN(npu_inst_pe_1_6_4_N68) );
  OR2_X1 npu_inst_pe_1_6_4_U123 ( .A1(npu_inst_pe_1_6_4_int_q_acc_3_), .A2(
        npu_inst_pe_1_6_4_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_6_4_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_6_4_U122 ( .A(npu_inst_pe_1_6_4_sub_67_carry_4_), .B(
        npu_inst_pe_1_6_4_int_q_acc_4_), .ZN(npu_inst_pe_1_6_4_N69) );
  OR2_X1 npu_inst_pe_1_6_4_U121 ( .A1(npu_inst_pe_1_6_4_int_q_acc_4_), .A2(
        npu_inst_pe_1_6_4_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_6_4_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_6_4_U120 ( .A(npu_inst_pe_1_6_4_sub_67_carry_5_), .B(
        npu_inst_pe_1_6_4_int_q_acc_5_), .ZN(npu_inst_pe_1_6_4_N70) );
  OR2_X1 npu_inst_pe_1_6_4_U119 ( .A1(npu_inst_pe_1_6_4_int_q_acc_5_), .A2(
        npu_inst_pe_1_6_4_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_6_4_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_6_4_U118 ( .A(npu_inst_pe_1_6_4_sub_67_carry_6_), .B(
        npu_inst_pe_1_6_4_int_q_acc_6_), .ZN(npu_inst_pe_1_6_4_N71) );
  OR2_X1 npu_inst_pe_1_6_4_U117 ( .A1(npu_inst_pe_1_6_4_int_q_acc_6_), .A2(
        npu_inst_pe_1_6_4_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_6_4_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_6_4_U116 ( .A(npu_inst_pe_1_6_4_int_q_acc_7_), .B(
        npu_inst_pe_1_6_4_sub_67_carry_7_), .ZN(npu_inst_pe_1_6_4_N72) );
  INV_X1 npu_inst_pe_1_6_4_U115 ( .A(npu_inst_n75), .ZN(npu_inst_pe_1_6_4_n6)
         );
  INV_X1 npu_inst_pe_1_6_4_U114 ( .A(npu_inst_n53), .ZN(npu_inst_pe_1_6_4_n3)
         );
  AOI22_X1 npu_inst_pe_1_6_4_U113 ( .A1(npu_inst_int_data_y_7__4__0_), .A2(
        npu_inst_pe_1_6_4_n58), .B1(npu_inst_pe_1_6_4_n118), .B2(
        npu_inst_pe_1_6_4_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_6_4_n57) );
  INV_X1 npu_inst_pe_1_6_4_U112 ( .A(npu_inst_pe_1_6_4_n57), .ZN(
        npu_inst_pe_1_6_4_n107) );
  AOI22_X1 npu_inst_pe_1_6_4_U111 ( .A1(npu_inst_int_data_y_7__4__0_), .A2(
        npu_inst_pe_1_6_4_n54), .B1(npu_inst_pe_1_6_4_n117), .B2(
        npu_inst_pe_1_6_4_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_6_4_n53) );
  INV_X1 npu_inst_pe_1_6_4_U110 ( .A(npu_inst_pe_1_6_4_n53), .ZN(
        npu_inst_pe_1_6_4_n108) );
  AOI22_X1 npu_inst_pe_1_6_4_U107 ( .A1(npu_inst_int_data_y_7__4__0_), .A2(
        npu_inst_pe_1_6_4_n50), .B1(npu_inst_pe_1_6_4_n116), .B2(
        npu_inst_pe_1_6_4_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_6_4_n49) );
  INV_X1 npu_inst_pe_1_6_4_U106 ( .A(npu_inst_pe_1_6_4_n49), .ZN(
        npu_inst_pe_1_6_4_n109) );
  AOI22_X1 npu_inst_pe_1_6_4_U105 ( .A1(npu_inst_int_data_y_7__4__0_), .A2(
        npu_inst_pe_1_6_4_n46), .B1(npu_inst_pe_1_6_4_n115), .B2(
        npu_inst_pe_1_6_4_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_6_4_n45) );
  INV_X1 npu_inst_pe_1_6_4_U104 ( .A(npu_inst_pe_1_6_4_n45), .ZN(
        npu_inst_pe_1_6_4_n110) );
  AOI22_X1 npu_inst_pe_1_6_4_U103 ( .A1(npu_inst_int_data_y_7__4__0_), .A2(
        npu_inst_pe_1_6_4_n42), .B1(npu_inst_pe_1_6_4_n114), .B2(
        npu_inst_pe_1_6_4_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_6_4_n41) );
  INV_X1 npu_inst_pe_1_6_4_U102 ( .A(npu_inst_pe_1_6_4_n41), .ZN(
        npu_inst_pe_1_6_4_n111) );
  AOI22_X1 npu_inst_pe_1_6_4_U101 ( .A1(npu_inst_int_data_y_7__4__1_), .A2(
        npu_inst_pe_1_6_4_n58), .B1(npu_inst_pe_1_6_4_n118), .B2(
        npu_inst_pe_1_6_4_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_6_4_n59) );
  INV_X1 npu_inst_pe_1_6_4_U100 ( .A(npu_inst_pe_1_6_4_n59), .ZN(
        npu_inst_pe_1_6_4_n101) );
  AOI22_X1 npu_inst_pe_1_6_4_U99 ( .A1(npu_inst_int_data_y_7__4__1_), .A2(
        npu_inst_pe_1_6_4_n54), .B1(npu_inst_pe_1_6_4_n117), .B2(
        npu_inst_pe_1_6_4_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_6_4_n55) );
  INV_X1 npu_inst_pe_1_6_4_U98 ( .A(npu_inst_pe_1_6_4_n55), .ZN(
        npu_inst_pe_1_6_4_n102) );
  AOI22_X1 npu_inst_pe_1_6_4_U97 ( .A1(npu_inst_int_data_y_7__4__1_), .A2(
        npu_inst_pe_1_6_4_n50), .B1(npu_inst_pe_1_6_4_n116), .B2(
        npu_inst_pe_1_6_4_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_6_4_n51) );
  INV_X1 npu_inst_pe_1_6_4_U96 ( .A(npu_inst_pe_1_6_4_n51), .ZN(
        npu_inst_pe_1_6_4_n103) );
  AOI22_X1 npu_inst_pe_1_6_4_U95 ( .A1(npu_inst_int_data_y_7__4__1_), .A2(
        npu_inst_pe_1_6_4_n46), .B1(npu_inst_pe_1_6_4_n115), .B2(
        npu_inst_pe_1_6_4_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_6_4_n47) );
  INV_X1 npu_inst_pe_1_6_4_U94 ( .A(npu_inst_pe_1_6_4_n47), .ZN(
        npu_inst_pe_1_6_4_n104) );
  AOI22_X1 npu_inst_pe_1_6_4_U93 ( .A1(npu_inst_int_data_y_7__4__1_), .A2(
        npu_inst_pe_1_6_4_n42), .B1(npu_inst_pe_1_6_4_n114), .B2(
        npu_inst_pe_1_6_4_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_6_4_n43) );
  INV_X1 npu_inst_pe_1_6_4_U92 ( .A(npu_inst_pe_1_6_4_n43), .ZN(
        npu_inst_pe_1_6_4_n105) );
  AOI22_X1 npu_inst_pe_1_6_4_U91 ( .A1(npu_inst_pe_1_6_4_n38), .A2(
        npu_inst_int_data_y_7__4__1_), .B1(npu_inst_pe_1_6_4_n113), .B2(
        npu_inst_pe_1_6_4_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_6_4_n39) );
  INV_X1 npu_inst_pe_1_6_4_U90 ( .A(npu_inst_pe_1_6_4_n39), .ZN(
        npu_inst_pe_1_6_4_n106) );
  AOI22_X1 npu_inst_pe_1_6_4_U89 ( .A1(npu_inst_pe_1_6_4_n38), .A2(
        npu_inst_int_data_y_7__4__0_), .B1(npu_inst_pe_1_6_4_n113), .B2(
        npu_inst_pe_1_6_4_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_6_4_n37) );
  INV_X1 npu_inst_pe_1_6_4_U88 ( .A(npu_inst_pe_1_6_4_n37), .ZN(
        npu_inst_pe_1_6_4_n112) );
  NAND2_X1 npu_inst_pe_1_6_4_U87 ( .A1(npu_inst_pe_1_6_4_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_6_4_n60), .ZN(npu_inst_pe_1_6_4_n74) );
  OAI21_X1 npu_inst_pe_1_6_4_U86 ( .B1(npu_inst_pe_1_6_4_n63), .B2(
        npu_inst_pe_1_6_4_n60), .A(npu_inst_pe_1_6_4_n74), .ZN(
        npu_inst_pe_1_6_4_n97) );
  NAND2_X1 npu_inst_pe_1_6_4_U85 ( .A1(npu_inst_pe_1_6_4_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_6_4_n60), .ZN(npu_inst_pe_1_6_4_n73) );
  OAI21_X1 npu_inst_pe_1_6_4_U84 ( .B1(npu_inst_pe_1_6_4_n61), .B2(
        npu_inst_pe_1_6_4_n60), .A(npu_inst_pe_1_6_4_n73), .ZN(
        npu_inst_pe_1_6_4_n96) );
  NAND2_X1 npu_inst_pe_1_6_4_U83 ( .A1(npu_inst_pe_1_6_4_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_6_4_n56), .ZN(npu_inst_pe_1_6_4_n72) );
  OAI21_X1 npu_inst_pe_1_6_4_U82 ( .B1(npu_inst_pe_1_6_4_n63), .B2(
        npu_inst_pe_1_6_4_n56), .A(npu_inst_pe_1_6_4_n72), .ZN(
        npu_inst_pe_1_6_4_n95) );
  NAND2_X1 npu_inst_pe_1_6_4_U81 ( .A1(npu_inst_pe_1_6_4_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_6_4_n56), .ZN(npu_inst_pe_1_6_4_n71) );
  OAI21_X1 npu_inst_pe_1_6_4_U80 ( .B1(npu_inst_pe_1_6_4_n61), .B2(
        npu_inst_pe_1_6_4_n56), .A(npu_inst_pe_1_6_4_n71), .ZN(
        npu_inst_pe_1_6_4_n94) );
  NAND2_X1 npu_inst_pe_1_6_4_U79 ( .A1(npu_inst_pe_1_6_4_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_6_4_n52), .ZN(npu_inst_pe_1_6_4_n70) );
  OAI21_X1 npu_inst_pe_1_6_4_U78 ( .B1(npu_inst_pe_1_6_4_n63), .B2(
        npu_inst_pe_1_6_4_n52), .A(npu_inst_pe_1_6_4_n70), .ZN(
        npu_inst_pe_1_6_4_n93) );
  NAND2_X1 npu_inst_pe_1_6_4_U77 ( .A1(npu_inst_pe_1_6_4_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_6_4_n52), .ZN(npu_inst_pe_1_6_4_n69) );
  OAI21_X1 npu_inst_pe_1_6_4_U76 ( .B1(npu_inst_pe_1_6_4_n61), .B2(
        npu_inst_pe_1_6_4_n52), .A(npu_inst_pe_1_6_4_n69), .ZN(
        npu_inst_pe_1_6_4_n92) );
  NAND2_X1 npu_inst_pe_1_6_4_U75 ( .A1(npu_inst_pe_1_6_4_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_6_4_n48), .ZN(npu_inst_pe_1_6_4_n68) );
  OAI21_X1 npu_inst_pe_1_6_4_U74 ( .B1(npu_inst_pe_1_6_4_n63), .B2(
        npu_inst_pe_1_6_4_n48), .A(npu_inst_pe_1_6_4_n68), .ZN(
        npu_inst_pe_1_6_4_n91) );
  NAND2_X1 npu_inst_pe_1_6_4_U73 ( .A1(npu_inst_pe_1_6_4_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_6_4_n48), .ZN(npu_inst_pe_1_6_4_n67) );
  OAI21_X1 npu_inst_pe_1_6_4_U72 ( .B1(npu_inst_pe_1_6_4_n61), .B2(
        npu_inst_pe_1_6_4_n48), .A(npu_inst_pe_1_6_4_n67), .ZN(
        npu_inst_pe_1_6_4_n90) );
  NAND2_X1 npu_inst_pe_1_6_4_U71 ( .A1(npu_inst_pe_1_6_4_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_6_4_n44), .ZN(npu_inst_pe_1_6_4_n66) );
  OAI21_X1 npu_inst_pe_1_6_4_U70 ( .B1(npu_inst_pe_1_6_4_n63), .B2(
        npu_inst_pe_1_6_4_n44), .A(npu_inst_pe_1_6_4_n66), .ZN(
        npu_inst_pe_1_6_4_n89) );
  NAND2_X1 npu_inst_pe_1_6_4_U69 ( .A1(npu_inst_pe_1_6_4_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_6_4_n44), .ZN(npu_inst_pe_1_6_4_n65) );
  OAI21_X1 npu_inst_pe_1_6_4_U68 ( .B1(npu_inst_pe_1_6_4_n61), .B2(
        npu_inst_pe_1_6_4_n44), .A(npu_inst_pe_1_6_4_n65), .ZN(
        npu_inst_pe_1_6_4_n88) );
  NAND2_X1 npu_inst_pe_1_6_4_U67 ( .A1(npu_inst_pe_1_6_4_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_6_4_n40), .ZN(npu_inst_pe_1_6_4_n64) );
  OAI21_X1 npu_inst_pe_1_6_4_U66 ( .B1(npu_inst_pe_1_6_4_n63), .B2(
        npu_inst_pe_1_6_4_n40), .A(npu_inst_pe_1_6_4_n64), .ZN(
        npu_inst_pe_1_6_4_n87) );
  NAND2_X1 npu_inst_pe_1_6_4_U65 ( .A1(npu_inst_pe_1_6_4_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_6_4_n40), .ZN(npu_inst_pe_1_6_4_n62) );
  OAI21_X1 npu_inst_pe_1_6_4_U64 ( .B1(npu_inst_pe_1_6_4_n61), .B2(
        npu_inst_pe_1_6_4_n40), .A(npu_inst_pe_1_6_4_n62), .ZN(
        npu_inst_pe_1_6_4_n86) );
  AND2_X1 npu_inst_pe_1_6_4_U63 ( .A1(npu_inst_pe_1_6_4_N93), .A2(npu_inst_n53), .ZN(npu_inst_int_data_y_6__4__0_) );
  AND2_X1 npu_inst_pe_1_6_4_U62 ( .A1(npu_inst_n53), .A2(npu_inst_pe_1_6_4_N94), .ZN(npu_inst_int_data_y_6__4__1_) );
  NOR3_X1 npu_inst_pe_1_6_4_U61 ( .A1(npu_inst_pe_1_6_4_n26), .A2(npu_inst_n53), .A3(npu_inst_int_ckg[11]), .ZN(npu_inst_pe_1_6_4_n85) );
  OR2_X1 npu_inst_pe_1_6_4_U60 ( .A1(npu_inst_pe_1_6_4_n85), .A2(
        npu_inst_pe_1_6_4_n2), .ZN(npu_inst_pe_1_6_4_N84) );
  AND2_X1 npu_inst_pe_1_6_4_U59 ( .A1(npu_inst_pe_1_6_4_int_q_acc_0_), .A2(
        npu_inst_pe_1_6_4_n1), .ZN(npu_inst_int_data_res_6__4__0_) );
  AND2_X1 npu_inst_pe_1_6_4_U58 ( .A1(npu_inst_pe_1_6_4_n2), .A2(
        npu_inst_pe_1_6_4_int_q_acc_7_), .ZN(npu_inst_int_data_res_6__4__7_)
         );
  AND2_X1 npu_inst_pe_1_6_4_U57 ( .A1(npu_inst_pe_1_6_4_int_q_acc_1_), .A2(
        npu_inst_pe_1_6_4_n1), .ZN(npu_inst_int_data_res_6__4__1_) );
  AND2_X1 npu_inst_pe_1_6_4_U56 ( .A1(npu_inst_pe_1_6_4_int_q_acc_2_), .A2(
        npu_inst_pe_1_6_4_n1), .ZN(npu_inst_int_data_res_6__4__2_) );
  AND2_X1 npu_inst_pe_1_6_4_U55 ( .A1(npu_inst_pe_1_6_4_int_q_acc_3_), .A2(
        npu_inst_pe_1_6_4_n2), .ZN(npu_inst_int_data_res_6__4__3_) );
  AND2_X1 npu_inst_pe_1_6_4_U54 ( .A1(npu_inst_pe_1_6_4_int_q_acc_4_), .A2(
        npu_inst_pe_1_6_4_n2), .ZN(npu_inst_int_data_res_6__4__4_) );
  AND2_X1 npu_inst_pe_1_6_4_U53 ( .A1(npu_inst_pe_1_6_4_int_q_acc_5_), .A2(
        npu_inst_pe_1_6_4_n2), .ZN(npu_inst_int_data_res_6__4__5_) );
  AND2_X1 npu_inst_pe_1_6_4_U52 ( .A1(npu_inst_pe_1_6_4_int_q_acc_6_), .A2(
        npu_inst_pe_1_6_4_n2), .ZN(npu_inst_int_data_res_6__4__6_) );
  AOI222_X1 npu_inst_pe_1_6_4_U51 ( .A1(npu_inst_int_data_res_7__4__0_), .A2(
        npu_inst_pe_1_6_4_n1), .B1(npu_inst_pe_1_6_4_N73), .B2(
        npu_inst_pe_1_6_4_n76), .C1(npu_inst_pe_1_6_4_N65), .C2(
        npu_inst_pe_1_6_4_n77), .ZN(npu_inst_pe_1_6_4_n84) );
  INV_X1 npu_inst_pe_1_6_4_U50 ( .A(npu_inst_pe_1_6_4_n84), .ZN(
        npu_inst_pe_1_6_4_n100) );
  AOI222_X1 npu_inst_pe_1_6_4_U49 ( .A1(npu_inst_int_data_res_7__4__7_), .A2(
        npu_inst_pe_1_6_4_n1), .B1(npu_inst_pe_1_6_4_N80), .B2(
        npu_inst_pe_1_6_4_n76), .C1(npu_inst_pe_1_6_4_N72), .C2(
        npu_inst_pe_1_6_4_n77), .ZN(npu_inst_pe_1_6_4_n75) );
  INV_X1 npu_inst_pe_1_6_4_U48 ( .A(npu_inst_pe_1_6_4_n75), .ZN(
        npu_inst_pe_1_6_4_n32) );
  AOI222_X1 npu_inst_pe_1_6_4_U47 ( .A1(npu_inst_int_data_res_7__4__1_), .A2(
        npu_inst_pe_1_6_4_n1), .B1(npu_inst_pe_1_6_4_N74), .B2(
        npu_inst_pe_1_6_4_n76), .C1(npu_inst_pe_1_6_4_N66), .C2(
        npu_inst_pe_1_6_4_n77), .ZN(npu_inst_pe_1_6_4_n83) );
  INV_X1 npu_inst_pe_1_6_4_U46 ( .A(npu_inst_pe_1_6_4_n83), .ZN(
        npu_inst_pe_1_6_4_n99) );
  AOI222_X1 npu_inst_pe_1_6_4_U45 ( .A1(npu_inst_int_data_res_7__4__2_), .A2(
        npu_inst_pe_1_6_4_n1), .B1(npu_inst_pe_1_6_4_N75), .B2(
        npu_inst_pe_1_6_4_n76), .C1(npu_inst_pe_1_6_4_N67), .C2(
        npu_inst_pe_1_6_4_n77), .ZN(npu_inst_pe_1_6_4_n82) );
  INV_X1 npu_inst_pe_1_6_4_U44 ( .A(npu_inst_pe_1_6_4_n82), .ZN(
        npu_inst_pe_1_6_4_n98) );
  AOI222_X1 npu_inst_pe_1_6_4_U43 ( .A1(npu_inst_int_data_res_7__4__3_), .A2(
        npu_inst_pe_1_6_4_n1), .B1(npu_inst_pe_1_6_4_N76), .B2(
        npu_inst_pe_1_6_4_n76), .C1(npu_inst_pe_1_6_4_N68), .C2(
        npu_inst_pe_1_6_4_n77), .ZN(npu_inst_pe_1_6_4_n81) );
  INV_X1 npu_inst_pe_1_6_4_U42 ( .A(npu_inst_pe_1_6_4_n81), .ZN(
        npu_inst_pe_1_6_4_n36) );
  AOI222_X1 npu_inst_pe_1_6_4_U41 ( .A1(npu_inst_int_data_res_7__4__4_), .A2(
        npu_inst_pe_1_6_4_n1), .B1(npu_inst_pe_1_6_4_N77), .B2(
        npu_inst_pe_1_6_4_n76), .C1(npu_inst_pe_1_6_4_N69), .C2(
        npu_inst_pe_1_6_4_n77), .ZN(npu_inst_pe_1_6_4_n80) );
  INV_X1 npu_inst_pe_1_6_4_U40 ( .A(npu_inst_pe_1_6_4_n80), .ZN(
        npu_inst_pe_1_6_4_n35) );
  AOI222_X1 npu_inst_pe_1_6_4_U39 ( .A1(npu_inst_int_data_res_7__4__5_), .A2(
        npu_inst_pe_1_6_4_n1), .B1(npu_inst_pe_1_6_4_N78), .B2(
        npu_inst_pe_1_6_4_n76), .C1(npu_inst_pe_1_6_4_N70), .C2(
        npu_inst_pe_1_6_4_n77), .ZN(npu_inst_pe_1_6_4_n79) );
  INV_X1 npu_inst_pe_1_6_4_U38 ( .A(npu_inst_pe_1_6_4_n79), .ZN(
        npu_inst_pe_1_6_4_n34) );
  AOI222_X1 npu_inst_pe_1_6_4_U37 ( .A1(npu_inst_int_data_res_7__4__6_), .A2(
        npu_inst_pe_1_6_4_n1), .B1(npu_inst_pe_1_6_4_N79), .B2(
        npu_inst_pe_1_6_4_n76), .C1(npu_inst_pe_1_6_4_N71), .C2(
        npu_inst_pe_1_6_4_n77), .ZN(npu_inst_pe_1_6_4_n78) );
  INV_X1 npu_inst_pe_1_6_4_U36 ( .A(npu_inst_pe_1_6_4_n78), .ZN(
        npu_inst_pe_1_6_4_n33) );
  INV_X1 npu_inst_pe_1_6_4_U35 ( .A(npu_inst_pe_1_6_4_int_data_1_), .ZN(
        npu_inst_pe_1_6_4_n13) );
  AND2_X1 npu_inst_pe_1_6_4_U34 ( .A1(npu_inst_int_data_x_6__4__1_), .A2(
        npu_inst_pe_1_6_4_int_q_weight_1_), .ZN(npu_inst_pe_1_6_4_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_6_4_U33 ( .A1(npu_inst_int_data_x_6__4__0_), .A2(
        npu_inst_pe_1_6_4_int_q_weight_1_), .ZN(npu_inst_pe_1_6_4_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_6_4_U32 ( .A1(npu_inst_n53), .A2(
        npu_inst_int_data_y_7__4__1_), .B1(npu_inst_pe_1_6_4_n3), .B2(
        npu_inst_int_data_x_6__5__1_), .ZN(npu_inst_pe_1_6_4_n63) );
  AOI22_X1 npu_inst_pe_1_6_4_U31 ( .A1(npu_inst_n53), .A2(
        npu_inst_int_data_y_7__4__0_), .B1(npu_inst_pe_1_6_4_n3), .B2(
        npu_inst_int_data_x_6__5__0_), .ZN(npu_inst_pe_1_6_4_n61) );
  INV_X1 npu_inst_pe_1_6_4_U30 ( .A(npu_inst_pe_1_6_4_int_data_0_), .ZN(
        npu_inst_pe_1_6_4_n12) );
  INV_X1 npu_inst_pe_1_6_4_U29 ( .A(npu_inst_n67), .ZN(npu_inst_pe_1_6_4_n5)
         );
  OR3_X1 npu_inst_pe_1_6_4_U28 ( .A1(npu_inst_n75), .A2(npu_inst_pe_1_6_4_n7), 
        .A3(npu_inst_pe_1_6_4_n5), .ZN(npu_inst_pe_1_6_4_n56) );
  OR3_X1 npu_inst_pe_1_6_4_U27 ( .A1(npu_inst_pe_1_6_4_n5), .A2(
        npu_inst_pe_1_6_4_n7), .A3(npu_inst_pe_1_6_4_n6), .ZN(
        npu_inst_pe_1_6_4_n48) );
  INV_X1 npu_inst_pe_1_6_4_U26 ( .A(npu_inst_pe_1_6_4_n5), .ZN(
        npu_inst_pe_1_6_4_n4) );
  OR3_X1 npu_inst_pe_1_6_4_U25 ( .A1(npu_inst_pe_1_6_4_n4), .A2(
        npu_inst_pe_1_6_4_n7), .A3(npu_inst_pe_1_6_4_n6), .ZN(
        npu_inst_pe_1_6_4_n52) );
  OR3_X1 npu_inst_pe_1_6_4_U24 ( .A1(npu_inst_n75), .A2(npu_inst_pe_1_6_4_n7), 
        .A3(npu_inst_pe_1_6_4_n4), .ZN(npu_inst_pe_1_6_4_n60) );
  NOR2_X1 npu_inst_pe_1_6_4_U23 ( .A1(npu_inst_pe_1_6_4_n60), .A2(
        npu_inst_pe_1_6_4_n3), .ZN(npu_inst_pe_1_6_4_n58) );
  NOR2_X1 npu_inst_pe_1_6_4_U22 ( .A1(npu_inst_pe_1_6_4_n56), .A2(
        npu_inst_pe_1_6_4_n3), .ZN(npu_inst_pe_1_6_4_n54) );
  NOR2_X1 npu_inst_pe_1_6_4_U21 ( .A1(npu_inst_pe_1_6_4_n52), .A2(
        npu_inst_pe_1_6_4_n3), .ZN(npu_inst_pe_1_6_4_n50) );
  NOR2_X1 npu_inst_pe_1_6_4_U20 ( .A1(npu_inst_pe_1_6_4_n48), .A2(
        npu_inst_pe_1_6_4_n3), .ZN(npu_inst_pe_1_6_4_n46) );
  NOR2_X1 npu_inst_pe_1_6_4_U19 ( .A1(npu_inst_pe_1_6_4_n40), .A2(
        npu_inst_pe_1_6_4_n3), .ZN(npu_inst_pe_1_6_4_n38) );
  NOR2_X1 npu_inst_pe_1_6_4_U18 ( .A1(npu_inst_pe_1_6_4_n44), .A2(
        npu_inst_pe_1_6_4_n3), .ZN(npu_inst_pe_1_6_4_n42) );
  BUF_X1 npu_inst_pe_1_6_4_U17 ( .A(npu_inst_n94), .Z(npu_inst_pe_1_6_4_n7) );
  INV_X1 npu_inst_pe_1_6_4_U16 ( .A(npu_inst_n122), .ZN(npu_inst_pe_1_6_4_n11)
         );
  INV_X1 npu_inst_pe_1_6_4_U15 ( .A(npu_inst_pe_1_6_4_n38), .ZN(
        npu_inst_pe_1_6_4_n113) );
  INV_X1 npu_inst_pe_1_6_4_U14 ( .A(npu_inst_pe_1_6_4_n58), .ZN(
        npu_inst_pe_1_6_4_n118) );
  INV_X1 npu_inst_pe_1_6_4_U13 ( .A(npu_inst_pe_1_6_4_n54), .ZN(
        npu_inst_pe_1_6_4_n117) );
  INV_X1 npu_inst_pe_1_6_4_U12 ( .A(npu_inst_pe_1_6_4_n50), .ZN(
        npu_inst_pe_1_6_4_n116) );
  INV_X1 npu_inst_pe_1_6_4_U11 ( .A(npu_inst_pe_1_6_4_n46), .ZN(
        npu_inst_pe_1_6_4_n115) );
  INV_X1 npu_inst_pe_1_6_4_U10 ( .A(npu_inst_pe_1_6_4_n42), .ZN(
        npu_inst_pe_1_6_4_n114) );
  BUF_X1 npu_inst_pe_1_6_4_U9 ( .A(npu_inst_n12), .Z(npu_inst_pe_1_6_4_n2) );
  BUF_X1 npu_inst_pe_1_6_4_U8 ( .A(npu_inst_n12), .Z(npu_inst_pe_1_6_4_n1) );
  BUF_X1 npu_inst_pe_1_6_4_U7 ( .A(npu_inst_pe_1_6_4_n11), .Z(
        npu_inst_pe_1_6_4_n10) );
  BUF_X1 npu_inst_pe_1_6_4_U6 ( .A(npu_inst_pe_1_6_4_n11), .Z(
        npu_inst_pe_1_6_4_n9) );
  BUF_X1 npu_inst_pe_1_6_4_U5 ( .A(npu_inst_pe_1_6_4_n11), .Z(
        npu_inst_pe_1_6_4_n8) );
  NOR2_X1 npu_inst_pe_1_6_4_U4 ( .A1(npu_inst_pe_1_6_4_int_q_weight_0_), .A2(
        npu_inst_pe_1_6_4_n1), .ZN(npu_inst_pe_1_6_4_n76) );
  NOR2_X1 npu_inst_pe_1_6_4_U3 ( .A1(npu_inst_pe_1_6_4_n27), .A2(
        npu_inst_pe_1_6_4_n1), .ZN(npu_inst_pe_1_6_4_n77) );
  FA_X1 npu_inst_pe_1_6_4_sub_67_U2_1 ( .A(npu_inst_pe_1_6_4_int_q_acc_1_), 
        .B(npu_inst_pe_1_6_4_n13), .CI(npu_inst_pe_1_6_4_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_6_4_sub_67_carry_2_), .S(npu_inst_pe_1_6_4_N66) );
  FA_X1 npu_inst_pe_1_6_4_add_69_U1_1 ( .A(npu_inst_pe_1_6_4_int_q_acc_1_), 
        .B(npu_inst_pe_1_6_4_int_data_1_), .CI(
        npu_inst_pe_1_6_4_add_69_carry_1_), .CO(
        npu_inst_pe_1_6_4_add_69_carry_2_), .S(npu_inst_pe_1_6_4_N74) );
  NAND3_X1 npu_inst_pe_1_6_4_U109 ( .A1(npu_inst_pe_1_6_4_n5), .A2(
        npu_inst_pe_1_6_4_n6), .A3(npu_inst_pe_1_6_4_n7), .ZN(
        npu_inst_pe_1_6_4_n44) );
  NAND3_X1 npu_inst_pe_1_6_4_U108 ( .A1(npu_inst_pe_1_6_4_n4), .A2(
        npu_inst_pe_1_6_4_n6), .A3(npu_inst_pe_1_6_4_n7), .ZN(
        npu_inst_pe_1_6_4_n40) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_6_4_n33), .CK(
        npu_inst_pe_1_6_4_net3366), .RN(npu_inst_pe_1_6_4_n8), .Q(
        npu_inst_pe_1_6_4_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_6_4_n34), .CK(
        npu_inst_pe_1_6_4_net3366), .RN(npu_inst_pe_1_6_4_n8), .Q(
        npu_inst_pe_1_6_4_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_6_4_n35), .CK(
        npu_inst_pe_1_6_4_net3366), .RN(npu_inst_pe_1_6_4_n8), .Q(
        npu_inst_pe_1_6_4_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_6_4_n36), .CK(
        npu_inst_pe_1_6_4_net3366), .RN(npu_inst_pe_1_6_4_n8), .Q(
        npu_inst_pe_1_6_4_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_6_4_n98), .CK(
        npu_inst_pe_1_6_4_net3366), .RN(npu_inst_pe_1_6_4_n8), .Q(
        npu_inst_pe_1_6_4_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_6_4_n99), .CK(
        npu_inst_pe_1_6_4_net3366), .RN(npu_inst_pe_1_6_4_n8), .Q(
        npu_inst_pe_1_6_4_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_6_4_n32), .CK(
        npu_inst_pe_1_6_4_net3366), .RN(npu_inst_pe_1_6_4_n8), .Q(
        npu_inst_pe_1_6_4_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_6_4_n100), 
        .CK(npu_inst_pe_1_6_4_net3366), .RN(npu_inst_pe_1_6_4_n8), .Q(
        npu_inst_pe_1_6_4_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_weight_reg_0_ ( .D(npu_inst_n108), .CK(
        npu_inst_pe_1_6_4_net3372), .RN(npu_inst_pe_1_6_4_n8), .Q(
        npu_inst_pe_1_6_4_int_q_weight_0_), .QN(npu_inst_pe_1_6_4_n27) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_weight_reg_1_ ( .D(npu_inst_n114), .CK(
        npu_inst_pe_1_6_4_net3372), .RN(npu_inst_pe_1_6_4_n8), .Q(
        npu_inst_pe_1_6_4_int_q_weight_1_), .QN(npu_inst_pe_1_6_4_n26) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_6_4_n112), 
        .CK(npu_inst_pe_1_6_4_net3372), .RN(npu_inst_pe_1_6_4_n8), .Q(
        npu_inst_pe_1_6_4_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_6_4_n106), 
        .CK(npu_inst_pe_1_6_4_net3372), .RN(npu_inst_pe_1_6_4_n8), .Q(
        npu_inst_pe_1_6_4_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_6_4_n111), 
        .CK(npu_inst_pe_1_6_4_net3372), .RN(npu_inst_pe_1_6_4_n9), .Q(
        npu_inst_pe_1_6_4_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_6_4_n105), 
        .CK(npu_inst_pe_1_6_4_net3372), .RN(npu_inst_pe_1_6_4_n9), .Q(
        npu_inst_pe_1_6_4_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_6_4_n110), 
        .CK(npu_inst_pe_1_6_4_net3372), .RN(npu_inst_pe_1_6_4_n9), .Q(
        npu_inst_pe_1_6_4_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_6_4_n104), 
        .CK(npu_inst_pe_1_6_4_net3372), .RN(npu_inst_pe_1_6_4_n9), .Q(
        npu_inst_pe_1_6_4_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_6_4_n109), 
        .CK(npu_inst_pe_1_6_4_net3372), .RN(npu_inst_pe_1_6_4_n9), .Q(
        npu_inst_pe_1_6_4_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_6_4_n103), 
        .CK(npu_inst_pe_1_6_4_net3372), .RN(npu_inst_pe_1_6_4_n9), .Q(
        npu_inst_pe_1_6_4_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_6_4_n108), 
        .CK(npu_inst_pe_1_6_4_net3372), .RN(npu_inst_pe_1_6_4_n9), .Q(
        npu_inst_pe_1_6_4_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_6_4_n102), 
        .CK(npu_inst_pe_1_6_4_net3372), .RN(npu_inst_pe_1_6_4_n9), .Q(
        npu_inst_pe_1_6_4_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_6_4_n107), 
        .CK(npu_inst_pe_1_6_4_net3372), .RN(npu_inst_pe_1_6_4_n9), .Q(
        npu_inst_pe_1_6_4_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_6_4_n101), 
        .CK(npu_inst_pe_1_6_4_net3372), .RN(npu_inst_pe_1_6_4_n9), .Q(
        npu_inst_pe_1_6_4_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_6_4_n86), 
        .CK(npu_inst_pe_1_6_4_net3372), .RN(npu_inst_pe_1_6_4_n9), .Q(
        npu_inst_pe_1_6_4_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_6_4_n87), 
        .CK(npu_inst_pe_1_6_4_net3372), .RN(npu_inst_pe_1_6_4_n9), .Q(
        npu_inst_pe_1_6_4_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_6_4_n88), 
        .CK(npu_inst_pe_1_6_4_net3372), .RN(npu_inst_pe_1_6_4_n10), .Q(
        npu_inst_pe_1_6_4_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_6_4_n89), 
        .CK(npu_inst_pe_1_6_4_net3372), .RN(npu_inst_pe_1_6_4_n10), .Q(
        npu_inst_pe_1_6_4_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_6_4_n90), 
        .CK(npu_inst_pe_1_6_4_net3372), .RN(npu_inst_pe_1_6_4_n10), .Q(
        npu_inst_pe_1_6_4_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_6_4_n91), 
        .CK(npu_inst_pe_1_6_4_net3372), .RN(npu_inst_pe_1_6_4_n10), .Q(
        npu_inst_pe_1_6_4_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_6_4_n92), 
        .CK(npu_inst_pe_1_6_4_net3372), .RN(npu_inst_pe_1_6_4_n10), .Q(
        npu_inst_pe_1_6_4_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_6_4_n93), 
        .CK(npu_inst_pe_1_6_4_net3372), .RN(npu_inst_pe_1_6_4_n10), .Q(
        npu_inst_pe_1_6_4_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_6_4_n94), 
        .CK(npu_inst_pe_1_6_4_net3372), .RN(npu_inst_pe_1_6_4_n10), .Q(
        npu_inst_pe_1_6_4_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_6_4_n95), 
        .CK(npu_inst_pe_1_6_4_net3372), .RN(npu_inst_pe_1_6_4_n10), .Q(
        npu_inst_pe_1_6_4_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_6_4_n96), 
        .CK(npu_inst_pe_1_6_4_net3372), .RN(npu_inst_pe_1_6_4_n10), .Q(
        npu_inst_pe_1_6_4_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_6_4_n97), 
        .CK(npu_inst_pe_1_6_4_net3372), .RN(npu_inst_pe_1_6_4_n10), .Q(
        npu_inst_pe_1_6_4_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_6_4_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_6_4_N84), .SE(1'b0), .GCK(npu_inst_pe_1_6_4_net3366) );
  CLKGATETST_X1 npu_inst_pe_1_6_4_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n62), .SE(1'b0), .GCK(npu_inst_pe_1_6_4_net3372) );
  MUX2_X1 npu_inst_pe_1_6_5_U162 ( .A(npu_inst_pe_1_6_5_n32), .B(
        npu_inst_pe_1_6_5_n29), .S(npu_inst_pe_1_6_5_n8), .Z(
        npu_inst_pe_1_6_5_N93) );
  MUX2_X1 npu_inst_pe_1_6_5_U161 ( .A(npu_inst_pe_1_6_5_n31), .B(
        npu_inst_pe_1_6_5_n30), .S(npu_inst_pe_1_6_5_n6), .Z(
        npu_inst_pe_1_6_5_n32) );
  MUX2_X1 npu_inst_pe_1_6_5_U160 ( .A(npu_inst_pe_1_6_5_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_6_5_int_q_reg_v_1__0_), .S(npu_inst_pe_1_6_5_n4), .Z(
        npu_inst_pe_1_6_5_n31) );
  MUX2_X1 npu_inst_pe_1_6_5_U159 ( .A(npu_inst_pe_1_6_5_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_6_5_int_q_reg_v_3__0_), .S(npu_inst_pe_1_6_5_n4), .Z(
        npu_inst_pe_1_6_5_n30) );
  MUX2_X1 npu_inst_pe_1_6_5_U158 ( .A(npu_inst_pe_1_6_5_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_6_5_int_q_reg_v_5__0_), .S(npu_inst_pe_1_6_5_n4), .Z(
        npu_inst_pe_1_6_5_n29) );
  MUX2_X1 npu_inst_pe_1_6_5_U157 ( .A(npu_inst_pe_1_6_5_n28), .B(
        npu_inst_pe_1_6_5_n23), .S(npu_inst_pe_1_6_5_n8), .Z(
        npu_inst_pe_1_6_5_N94) );
  MUX2_X1 npu_inst_pe_1_6_5_U156 ( .A(npu_inst_pe_1_6_5_n25), .B(
        npu_inst_pe_1_6_5_n24), .S(npu_inst_pe_1_6_5_n6), .Z(
        npu_inst_pe_1_6_5_n28) );
  MUX2_X1 npu_inst_pe_1_6_5_U155 ( .A(npu_inst_pe_1_6_5_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_6_5_int_q_reg_v_1__1_), .S(npu_inst_pe_1_6_5_n4), .Z(
        npu_inst_pe_1_6_5_n25) );
  MUX2_X1 npu_inst_pe_1_6_5_U154 ( .A(npu_inst_pe_1_6_5_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_6_5_int_q_reg_v_3__1_), .S(npu_inst_pe_1_6_5_n4), .Z(
        npu_inst_pe_1_6_5_n24) );
  MUX2_X1 npu_inst_pe_1_6_5_U153 ( .A(npu_inst_pe_1_6_5_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_6_5_int_q_reg_v_5__1_), .S(npu_inst_pe_1_6_5_n4), .Z(
        npu_inst_pe_1_6_5_n23) );
  MUX2_X1 npu_inst_pe_1_6_5_U152 ( .A(npu_inst_pe_1_6_5_n22), .B(
        npu_inst_pe_1_6_5_n19), .S(npu_inst_pe_1_6_5_n8), .Z(
        npu_inst_int_data_x_6__5__1_) );
  MUX2_X1 npu_inst_pe_1_6_5_U151 ( .A(npu_inst_pe_1_6_5_n21), .B(
        npu_inst_pe_1_6_5_n20), .S(npu_inst_pe_1_6_5_n6), .Z(
        npu_inst_pe_1_6_5_n22) );
  MUX2_X1 npu_inst_pe_1_6_5_U150 ( .A(npu_inst_pe_1_6_5_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_6_5_int_q_reg_h_1__1_), .S(npu_inst_pe_1_6_5_n4), .Z(
        npu_inst_pe_1_6_5_n21) );
  MUX2_X1 npu_inst_pe_1_6_5_U149 ( .A(npu_inst_pe_1_6_5_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_6_5_int_q_reg_h_3__1_), .S(npu_inst_pe_1_6_5_n4), .Z(
        npu_inst_pe_1_6_5_n20) );
  MUX2_X1 npu_inst_pe_1_6_5_U148 ( .A(npu_inst_pe_1_6_5_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_6_5_int_q_reg_h_5__1_), .S(npu_inst_pe_1_6_5_n4), .Z(
        npu_inst_pe_1_6_5_n19) );
  MUX2_X1 npu_inst_pe_1_6_5_U147 ( .A(npu_inst_pe_1_6_5_n18), .B(
        npu_inst_pe_1_6_5_n15), .S(npu_inst_pe_1_6_5_n8), .Z(
        npu_inst_int_data_x_6__5__0_) );
  MUX2_X1 npu_inst_pe_1_6_5_U146 ( .A(npu_inst_pe_1_6_5_n17), .B(
        npu_inst_pe_1_6_5_n16), .S(npu_inst_pe_1_6_5_n6), .Z(
        npu_inst_pe_1_6_5_n18) );
  MUX2_X1 npu_inst_pe_1_6_5_U145 ( .A(npu_inst_pe_1_6_5_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_6_5_int_q_reg_h_1__0_), .S(npu_inst_pe_1_6_5_n4), .Z(
        npu_inst_pe_1_6_5_n17) );
  MUX2_X1 npu_inst_pe_1_6_5_U144 ( .A(npu_inst_pe_1_6_5_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_6_5_int_q_reg_h_3__0_), .S(npu_inst_pe_1_6_5_n4), .Z(
        npu_inst_pe_1_6_5_n16) );
  MUX2_X1 npu_inst_pe_1_6_5_U143 ( .A(npu_inst_pe_1_6_5_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_6_5_int_q_reg_h_5__0_), .S(npu_inst_pe_1_6_5_n4), .Z(
        npu_inst_pe_1_6_5_n15) );
  XOR2_X1 npu_inst_pe_1_6_5_U142 ( .A(npu_inst_pe_1_6_5_int_data_0_), .B(
        npu_inst_pe_1_6_5_int_q_acc_0_), .Z(npu_inst_pe_1_6_5_N73) );
  AND2_X1 npu_inst_pe_1_6_5_U141 ( .A1(npu_inst_pe_1_6_5_int_q_acc_0_), .A2(
        npu_inst_pe_1_6_5_int_data_0_), .ZN(npu_inst_pe_1_6_5_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_6_5_U140 ( .A(npu_inst_pe_1_6_5_int_q_acc_0_), .B(
        npu_inst_pe_1_6_5_n13), .ZN(npu_inst_pe_1_6_5_N65) );
  OR2_X1 npu_inst_pe_1_6_5_U139 ( .A1(npu_inst_pe_1_6_5_n13), .A2(
        npu_inst_pe_1_6_5_int_q_acc_0_), .ZN(npu_inst_pe_1_6_5_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_6_5_U138 ( .A(npu_inst_pe_1_6_5_int_q_acc_2_), .B(
        npu_inst_pe_1_6_5_add_69_carry_2_), .Z(npu_inst_pe_1_6_5_N75) );
  AND2_X1 npu_inst_pe_1_6_5_U137 ( .A1(npu_inst_pe_1_6_5_add_69_carry_2_), 
        .A2(npu_inst_pe_1_6_5_int_q_acc_2_), .ZN(
        npu_inst_pe_1_6_5_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_6_5_U136 ( .A(npu_inst_pe_1_6_5_int_q_acc_3_), .B(
        npu_inst_pe_1_6_5_add_69_carry_3_), .Z(npu_inst_pe_1_6_5_N76) );
  AND2_X1 npu_inst_pe_1_6_5_U135 ( .A1(npu_inst_pe_1_6_5_add_69_carry_3_), 
        .A2(npu_inst_pe_1_6_5_int_q_acc_3_), .ZN(
        npu_inst_pe_1_6_5_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_6_5_U134 ( .A(npu_inst_pe_1_6_5_int_q_acc_4_), .B(
        npu_inst_pe_1_6_5_add_69_carry_4_), .Z(npu_inst_pe_1_6_5_N77) );
  AND2_X1 npu_inst_pe_1_6_5_U133 ( .A1(npu_inst_pe_1_6_5_add_69_carry_4_), 
        .A2(npu_inst_pe_1_6_5_int_q_acc_4_), .ZN(
        npu_inst_pe_1_6_5_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_6_5_U132 ( .A(npu_inst_pe_1_6_5_int_q_acc_5_), .B(
        npu_inst_pe_1_6_5_add_69_carry_5_), .Z(npu_inst_pe_1_6_5_N78) );
  AND2_X1 npu_inst_pe_1_6_5_U131 ( .A1(npu_inst_pe_1_6_5_add_69_carry_5_), 
        .A2(npu_inst_pe_1_6_5_int_q_acc_5_), .ZN(
        npu_inst_pe_1_6_5_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_6_5_U130 ( .A(npu_inst_pe_1_6_5_int_q_acc_6_), .B(
        npu_inst_pe_1_6_5_add_69_carry_6_), .Z(npu_inst_pe_1_6_5_N79) );
  AND2_X1 npu_inst_pe_1_6_5_U129 ( .A1(npu_inst_pe_1_6_5_add_69_carry_6_), 
        .A2(npu_inst_pe_1_6_5_int_q_acc_6_), .ZN(
        npu_inst_pe_1_6_5_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_6_5_U128 ( .A(npu_inst_pe_1_6_5_int_q_acc_7_), .B(
        npu_inst_pe_1_6_5_add_69_carry_7_), .Z(npu_inst_pe_1_6_5_N80) );
  XNOR2_X1 npu_inst_pe_1_6_5_U127 ( .A(npu_inst_pe_1_6_5_sub_67_carry_2_), .B(
        npu_inst_pe_1_6_5_int_q_acc_2_), .ZN(npu_inst_pe_1_6_5_N67) );
  OR2_X1 npu_inst_pe_1_6_5_U126 ( .A1(npu_inst_pe_1_6_5_int_q_acc_2_), .A2(
        npu_inst_pe_1_6_5_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_6_5_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_6_5_U125 ( .A(npu_inst_pe_1_6_5_sub_67_carry_3_), .B(
        npu_inst_pe_1_6_5_int_q_acc_3_), .ZN(npu_inst_pe_1_6_5_N68) );
  OR2_X1 npu_inst_pe_1_6_5_U124 ( .A1(npu_inst_pe_1_6_5_int_q_acc_3_), .A2(
        npu_inst_pe_1_6_5_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_6_5_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_6_5_U123 ( .A(npu_inst_pe_1_6_5_sub_67_carry_4_), .B(
        npu_inst_pe_1_6_5_int_q_acc_4_), .ZN(npu_inst_pe_1_6_5_N69) );
  OR2_X1 npu_inst_pe_1_6_5_U122 ( .A1(npu_inst_pe_1_6_5_int_q_acc_4_), .A2(
        npu_inst_pe_1_6_5_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_6_5_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_6_5_U121 ( .A(npu_inst_pe_1_6_5_sub_67_carry_5_), .B(
        npu_inst_pe_1_6_5_int_q_acc_5_), .ZN(npu_inst_pe_1_6_5_N70) );
  OR2_X1 npu_inst_pe_1_6_5_U120 ( .A1(npu_inst_pe_1_6_5_int_q_acc_5_), .A2(
        npu_inst_pe_1_6_5_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_6_5_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_6_5_U119 ( .A(npu_inst_pe_1_6_5_sub_67_carry_6_), .B(
        npu_inst_pe_1_6_5_int_q_acc_6_), .ZN(npu_inst_pe_1_6_5_N71) );
  OR2_X1 npu_inst_pe_1_6_5_U118 ( .A1(npu_inst_pe_1_6_5_int_q_acc_6_), .A2(
        npu_inst_pe_1_6_5_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_6_5_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_6_5_U117 ( .A(npu_inst_pe_1_6_5_int_q_acc_7_), .B(
        npu_inst_pe_1_6_5_sub_67_carry_7_), .ZN(npu_inst_pe_1_6_5_N72) );
  INV_X1 npu_inst_pe_1_6_5_U116 ( .A(npu_inst_n75), .ZN(npu_inst_pe_1_6_5_n7)
         );
  INV_X1 npu_inst_pe_1_6_5_U115 ( .A(npu_inst_pe_1_6_5_n7), .ZN(
        npu_inst_pe_1_6_5_n6) );
  INV_X1 npu_inst_pe_1_6_5_U114 ( .A(npu_inst_n53), .ZN(npu_inst_pe_1_6_5_n3)
         );
  AOI22_X1 npu_inst_pe_1_6_5_U113 ( .A1(npu_inst_int_data_y_7__5__0_), .A2(
        npu_inst_pe_1_6_5_n58), .B1(npu_inst_pe_1_6_5_n119), .B2(
        npu_inst_pe_1_6_5_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_6_5_n57) );
  INV_X1 npu_inst_pe_1_6_5_U112 ( .A(npu_inst_pe_1_6_5_n57), .ZN(
        npu_inst_pe_1_6_5_n108) );
  AOI22_X1 npu_inst_pe_1_6_5_U111 ( .A1(npu_inst_int_data_y_7__5__0_), .A2(
        npu_inst_pe_1_6_5_n54), .B1(npu_inst_pe_1_6_5_n118), .B2(
        npu_inst_pe_1_6_5_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_6_5_n53) );
  INV_X1 npu_inst_pe_1_6_5_U110 ( .A(npu_inst_pe_1_6_5_n53), .ZN(
        npu_inst_pe_1_6_5_n109) );
  AOI22_X1 npu_inst_pe_1_6_5_U107 ( .A1(npu_inst_int_data_y_7__5__0_), .A2(
        npu_inst_pe_1_6_5_n50), .B1(npu_inst_pe_1_6_5_n117), .B2(
        npu_inst_pe_1_6_5_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_6_5_n49) );
  INV_X1 npu_inst_pe_1_6_5_U106 ( .A(npu_inst_pe_1_6_5_n49), .ZN(
        npu_inst_pe_1_6_5_n110) );
  AOI22_X1 npu_inst_pe_1_6_5_U105 ( .A1(npu_inst_int_data_y_7__5__0_), .A2(
        npu_inst_pe_1_6_5_n46), .B1(npu_inst_pe_1_6_5_n116), .B2(
        npu_inst_pe_1_6_5_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_6_5_n45) );
  INV_X1 npu_inst_pe_1_6_5_U104 ( .A(npu_inst_pe_1_6_5_n45), .ZN(
        npu_inst_pe_1_6_5_n111) );
  AOI22_X1 npu_inst_pe_1_6_5_U103 ( .A1(npu_inst_int_data_y_7__5__0_), .A2(
        npu_inst_pe_1_6_5_n42), .B1(npu_inst_pe_1_6_5_n115), .B2(
        npu_inst_pe_1_6_5_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_6_5_n41) );
  INV_X1 npu_inst_pe_1_6_5_U102 ( .A(npu_inst_pe_1_6_5_n41), .ZN(
        npu_inst_pe_1_6_5_n112) );
  AOI22_X1 npu_inst_pe_1_6_5_U101 ( .A1(npu_inst_int_data_y_7__5__1_), .A2(
        npu_inst_pe_1_6_5_n58), .B1(npu_inst_pe_1_6_5_n119), .B2(
        npu_inst_pe_1_6_5_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_6_5_n59) );
  INV_X1 npu_inst_pe_1_6_5_U100 ( .A(npu_inst_pe_1_6_5_n59), .ZN(
        npu_inst_pe_1_6_5_n102) );
  AOI22_X1 npu_inst_pe_1_6_5_U99 ( .A1(npu_inst_int_data_y_7__5__1_), .A2(
        npu_inst_pe_1_6_5_n54), .B1(npu_inst_pe_1_6_5_n118), .B2(
        npu_inst_pe_1_6_5_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_6_5_n55) );
  INV_X1 npu_inst_pe_1_6_5_U98 ( .A(npu_inst_pe_1_6_5_n55), .ZN(
        npu_inst_pe_1_6_5_n103) );
  AOI22_X1 npu_inst_pe_1_6_5_U97 ( .A1(npu_inst_int_data_y_7__5__1_), .A2(
        npu_inst_pe_1_6_5_n50), .B1(npu_inst_pe_1_6_5_n117), .B2(
        npu_inst_pe_1_6_5_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_6_5_n51) );
  INV_X1 npu_inst_pe_1_6_5_U96 ( .A(npu_inst_pe_1_6_5_n51), .ZN(
        npu_inst_pe_1_6_5_n104) );
  AOI22_X1 npu_inst_pe_1_6_5_U95 ( .A1(npu_inst_int_data_y_7__5__1_), .A2(
        npu_inst_pe_1_6_5_n46), .B1(npu_inst_pe_1_6_5_n116), .B2(
        npu_inst_pe_1_6_5_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_6_5_n47) );
  INV_X1 npu_inst_pe_1_6_5_U94 ( .A(npu_inst_pe_1_6_5_n47), .ZN(
        npu_inst_pe_1_6_5_n105) );
  AOI22_X1 npu_inst_pe_1_6_5_U93 ( .A1(npu_inst_int_data_y_7__5__1_), .A2(
        npu_inst_pe_1_6_5_n42), .B1(npu_inst_pe_1_6_5_n115), .B2(
        npu_inst_pe_1_6_5_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_6_5_n43) );
  INV_X1 npu_inst_pe_1_6_5_U92 ( .A(npu_inst_pe_1_6_5_n43), .ZN(
        npu_inst_pe_1_6_5_n106) );
  AOI22_X1 npu_inst_pe_1_6_5_U91 ( .A1(npu_inst_pe_1_6_5_n38), .A2(
        npu_inst_int_data_y_7__5__1_), .B1(npu_inst_pe_1_6_5_n114), .B2(
        npu_inst_pe_1_6_5_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_6_5_n39) );
  INV_X1 npu_inst_pe_1_6_5_U90 ( .A(npu_inst_pe_1_6_5_n39), .ZN(
        npu_inst_pe_1_6_5_n107) );
  AOI22_X1 npu_inst_pe_1_6_5_U89 ( .A1(npu_inst_pe_1_6_5_n38), .A2(
        npu_inst_int_data_y_7__5__0_), .B1(npu_inst_pe_1_6_5_n114), .B2(
        npu_inst_pe_1_6_5_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_6_5_n37) );
  INV_X1 npu_inst_pe_1_6_5_U88 ( .A(npu_inst_pe_1_6_5_n37), .ZN(
        npu_inst_pe_1_6_5_n113) );
  NAND2_X1 npu_inst_pe_1_6_5_U87 ( .A1(npu_inst_pe_1_6_5_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_6_5_n60), .ZN(npu_inst_pe_1_6_5_n74) );
  OAI21_X1 npu_inst_pe_1_6_5_U86 ( .B1(npu_inst_pe_1_6_5_n63), .B2(
        npu_inst_pe_1_6_5_n60), .A(npu_inst_pe_1_6_5_n74), .ZN(
        npu_inst_pe_1_6_5_n97) );
  NAND2_X1 npu_inst_pe_1_6_5_U85 ( .A1(npu_inst_pe_1_6_5_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_6_5_n60), .ZN(npu_inst_pe_1_6_5_n73) );
  OAI21_X1 npu_inst_pe_1_6_5_U84 ( .B1(npu_inst_pe_1_6_5_n61), .B2(
        npu_inst_pe_1_6_5_n60), .A(npu_inst_pe_1_6_5_n73), .ZN(
        npu_inst_pe_1_6_5_n96) );
  NAND2_X1 npu_inst_pe_1_6_5_U83 ( .A1(npu_inst_pe_1_6_5_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_6_5_n56), .ZN(npu_inst_pe_1_6_5_n72) );
  OAI21_X1 npu_inst_pe_1_6_5_U82 ( .B1(npu_inst_pe_1_6_5_n63), .B2(
        npu_inst_pe_1_6_5_n56), .A(npu_inst_pe_1_6_5_n72), .ZN(
        npu_inst_pe_1_6_5_n95) );
  NAND2_X1 npu_inst_pe_1_6_5_U81 ( .A1(npu_inst_pe_1_6_5_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_6_5_n56), .ZN(npu_inst_pe_1_6_5_n71) );
  OAI21_X1 npu_inst_pe_1_6_5_U80 ( .B1(npu_inst_pe_1_6_5_n61), .B2(
        npu_inst_pe_1_6_5_n56), .A(npu_inst_pe_1_6_5_n71), .ZN(
        npu_inst_pe_1_6_5_n94) );
  NAND2_X1 npu_inst_pe_1_6_5_U79 ( .A1(npu_inst_pe_1_6_5_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_6_5_n52), .ZN(npu_inst_pe_1_6_5_n70) );
  OAI21_X1 npu_inst_pe_1_6_5_U78 ( .B1(npu_inst_pe_1_6_5_n63), .B2(
        npu_inst_pe_1_6_5_n52), .A(npu_inst_pe_1_6_5_n70), .ZN(
        npu_inst_pe_1_6_5_n93) );
  NAND2_X1 npu_inst_pe_1_6_5_U77 ( .A1(npu_inst_pe_1_6_5_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_6_5_n52), .ZN(npu_inst_pe_1_6_5_n69) );
  OAI21_X1 npu_inst_pe_1_6_5_U76 ( .B1(npu_inst_pe_1_6_5_n61), .B2(
        npu_inst_pe_1_6_5_n52), .A(npu_inst_pe_1_6_5_n69), .ZN(
        npu_inst_pe_1_6_5_n92) );
  NAND2_X1 npu_inst_pe_1_6_5_U75 ( .A1(npu_inst_pe_1_6_5_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_6_5_n48), .ZN(npu_inst_pe_1_6_5_n68) );
  OAI21_X1 npu_inst_pe_1_6_5_U74 ( .B1(npu_inst_pe_1_6_5_n63), .B2(
        npu_inst_pe_1_6_5_n48), .A(npu_inst_pe_1_6_5_n68), .ZN(
        npu_inst_pe_1_6_5_n91) );
  NAND2_X1 npu_inst_pe_1_6_5_U73 ( .A1(npu_inst_pe_1_6_5_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_6_5_n48), .ZN(npu_inst_pe_1_6_5_n67) );
  OAI21_X1 npu_inst_pe_1_6_5_U72 ( .B1(npu_inst_pe_1_6_5_n61), .B2(
        npu_inst_pe_1_6_5_n48), .A(npu_inst_pe_1_6_5_n67), .ZN(
        npu_inst_pe_1_6_5_n90) );
  NAND2_X1 npu_inst_pe_1_6_5_U71 ( .A1(npu_inst_pe_1_6_5_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_6_5_n44), .ZN(npu_inst_pe_1_6_5_n66) );
  OAI21_X1 npu_inst_pe_1_6_5_U70 ( .B1(npu_inst_pe_1_6_5_n63), .B2(
        npu_inst_pe_1_6_5_n44), .A(npu_inst_pe_1_6_5_n66), .ZN(
        npu_inst_pe_1_6_5_n89) );
  NAND2_X1 npu_inst_pe_1_6_5_U69 ( .A1(npu_inst_pe_1_6_5_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_6_5_n44), .ZN(npu_inst_pe_1_6_5_n65) );
  OAI21_X1 npu_inst_pe_1_6_5_U68 ( .B1(npu_inst_pe_1_6_5_n61), .B2(
        npu_inst_pe_1_6_5_n44), .A(npu_inst_pe_1_6_5_n65), .ZN(
        npu_inst_pe_1_6_5_n88) );
  NAND2_X1 npu_inst_pe_1_6_5_U67 ( .A1(npu_inst_pe_1_6_5_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_6_5_n40), .ZN(npu_inst_pe_1_6_5_n64) );
  OAI21_X1 npu_inst_pe_1_6_5_U66 ( .B1(npu_inst_pe_1_6_5_n63), .B2(
        npu_inst_pe_1_6_5_n40), .A(npu_inst_pe_1_6_5_n64), .ZN(
        npu_inst_pe_1_6_5_n87) );
  NAND2_X1 npu_inst_pe_1_6_5_U65 ( .A1(npu_inst_pe_1_6_5_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_6_5_n40), .ZN(npu_inst_pe_1_6_5_n62) );
  OAI21_X1 npu_inst_pe_1_6_5_U64 ( .B1(npu_inst_pe_1_6_5_n61), .B2(
        npu_inst_pe_1_6_5_n40), .A(npu_inst_pe_1_6_5_n62), .ZN(
        npu_inst_pe_1_6_5_n86) );
  AND2_X1 npu_inst_pe_1_6_5_U63 ( .A1(npu_inst_pe_1_6_5_N93), .A2(npu_inst_n53), .ZN(npu_inst_int_data_y_6__5__0_) );
  AND2_X1 npu_inst_pe_1_6_5_U62 ( .A1(npu_inst_n53), .A2(npu_inst_pe_1_6_5_N94), .ZN(npu_inst_int_data_y_6__5__1_) );
  NOR3_X1 npu_inst_pe_1_6_5_U61 ( .A1(npu_inst_pe_1_6_5_n26), .A2(npu_inst_n53), .A3(npu_inst_int_ckg[10]), .ZN(npu_inst_pe_1_6_5_n85) );
  OR2_X1 npu_inst_pe_1_6_5_U60 ( .A1(npu_inst_pe_1_6_5_n85), .A2(
        npu_inst_pe_1_6_5_n2), .ZN(npu_inst_pe_1_6_5_N84) );
  AND2_X1 npu_inst_pe_1_6_5_U59 ( .A1(npu_inst_pe_1_6_5_int_q_acc_0_), .A2(
        npu_inst_pe_1_6_5_n1), .ZN(npu_inst_int_data_res_6__5__0_) );
  AND2_X1 npu_inst_pe_1_6_5_U58 ( .A1(npu_inst_pe_1_6_5_n2), .A2(
        npu_inst_pe_1_6_5_int_q_acc_7_), .ZN(npu_inst_int_data_res_6__5__7_)
         );
  AND2_X1 npu_inst_pe_1_6_5_U57 ( .A1(npu_inst_pe_1_6_5_int_q_acc_1_), .A2(
        npu_inst_pe_1_6_5_n1), .ZN(npu_inst_int_data_res_6__5__1_) );
  AND2_X1 npu_inst_pe_1_6_5_U56 ( .A1(npu_inst_pe_1_6_5_int_q_acc_2_), .A2(
        npu_inst_pe_1_6_5_n1), .ZN(npu_inst_int_data_res_6__5__2_) );
  AND2_X1 npu_inst_pe_1_6_5_U55 ( .A1(npu_inst_pe_1_6_5_int_q_acc_3_), .A2(
        npu_inst_pe_1_6_5_n2), .ZN(npu_inst_int_data_res_6__5__3_) );
  AND2_X1 npu_inst_pe_1_6_5_U54 ( .A1(npu_inst_pe_1_6_5_int_q_acc_4_), .A2(
        npu_inst_pe_1_6_5_n2), .ZN(npu_inst_int_data_res_6__5__4_) );
  AND2_X1 npu_inst_pe_1_6_5_U53 ( .A1(npu_inst_pe_1_6_5_int_q_acc_5_), .A2(
        npu_inst_pe_1_6_5_n2), .ZN(npu_inst_int_data_res_6__5__5_) );
  AND2_X1 npu_inst_pe_1_6_5_U52 ( .A1(npu_inst_pe_1_6_5_int_q_acc_6_), .A2(
        npu_inst_pe_1_6_5_n2), .ZN(npu_inst_int_data_res_6__5__6_) );
  AOI222_X1 npu_inst_pe_1_6_5_U51 ( .A1(npu_inst_int_data_res_7__5__0_), .A2(
        npu_inst_pe_1_6_5_n1), .B1(npu_inst_pe_1_6_5_N73), .B2(
        npu_inst_pe_1_6_5_n76), .C1(npu_inst_pe_1_6_5_N65), .C2(
        npu_inst_pe_1_6_5_n77), .ZN(npu_inst_pe_1_6_5_n84) );
  INV_X1 npu_inst_pe_1_6_5_U50 ( .A(npu_inst_pe_1_6_5_n84), .ZN(
        npu_inst_pe_1_6_5_n101) );
  AOI222_X1 npu_inst_pe_1_6_5_U49 ( .A1(npu_inst_int_data_res_7__5__7_), .A2(
        npu_inst_pe_1_6_5_n1), .B1(npu_inst_pe_1_6_5_N80), .B2(
        npu_inst_pe_1_6_5_n76), .C1(npu_inst_pe_1_6_5_N72), .C2(
        npu_inst_pe_1_6_5_n77), .ZN(npu_inst_pe_1_6_5_n75) );
  INV_X1 npu_inst_pe_1_6_5_U48 ( .A(npu_inst_pe_1_6_5_n75), .ZN(
        npu_inst_pe_1_6_5_n33) );
  AOI222_X1 npu_inst_pe_1_6_5_U47 ( .A1(npu_inst_int_data_res_7__5__1_), .A2(
        npu_inst_pe_1_6_5_n1), .B1(npu_inst_pe_1_6_5_N74), .B2(
        npu_inst_pe_1_6_5_n76), .C1(npu_inst_pe_1_6_5_N66), .C2(
        npu_inst_pe_1_6_5_n77), .ZN(npu_inst_pe_1_6_5_n83) );
  INV_X1 npu_inst_pe_1_6_5_U46 ( .A(npu_inst_pe_1_6_5_n83), .ZN(
        npu_inst_pe_1_6_5_n100) );
  AOI222_X1 npu_inst_pe_1_6_5_U45 ( .A1(npu_inst_int_data_res_7__5__2_), .A2(
        npu_inst_pe_1_6_5_n1), .B1(npu_inst_pe_1_6_5_N75), .B2(
        npu_inst_pe_1_6_5_n76), .C1(npu_inst_pe_1_6_5_N67), .C2(
        npu_inst_pe_1_6_5_n77), .ZN(npu_inst_pe_1_6_5_n82) );
  INV_X1 npu_inst_pe_1_6_5_U44 ( .A(npu_inst_pe_1_6_5_n82), .ZN(
        npu_inst_pe_1_6_5_n99) );
  AOI222_X1 npu_inst_pe_1_6_5_U43 ( .A1(npu_inst_int_data_res_7__5__3_), .A2(
        npu_inst_pe_1_6_5_n1), .B1(npu_inst_pe_1_6_5_N76), .B2(
        npu_inst_pe_1_6_5_n76), .C1(npu_inst_pe_1_6_5_N68), .C2(
        npu_inst_pe_1_6_5_n77), .ZN(npu_inst_pe_1_6_5_n81) );
  INV_X1 npu_inst_pe_1_6_5_U42 ( .A(npu_inst_pe_1_6_5_n81), .ZN(
        npu_inst_pe_1_6_5_n98) );
  AOI222_X1 npu_inst_pe_1_6_5_U41 ( .A1(npu_inst_int_data_res_7__5__4_), .A2(
        npu_inst_pe_1_6_5_n1), .B1(npu_inst_pe_1_6_5_N77), .B2(
        npu_inst_pe_1_6_5_n76), .C1(npu_inst_pe_1_6_5_N69), .C2(
        npu_inst_pe_1_6_5_n77), .ZN(npu_inst_pe_1_6_5_n80) );
  INV_X1 npu_inst_pe_1_6_5_U40 ( .A(npu_inst_pe_1_6_5_n80), .ZN(
        npu_inst_pe_1_6_5_n36) );
  AOI222_X1 npu_inst_pe_1_6_5_U39 ( .A1(npu_inst_int_data_res_7__5__5_), .A2(
        npu_inst_pe_1_6_5_n1), .B1(npu_inst_pe_1_6_5_N78), .B2(
        npu_inst_pe_1_6_5_n76), .C1(npu_inst_pe_1_6_5_N70), .C2(
        npu_inst_pe_1_6_5_n77), .ZN(npu_inst_pe_1_6_5_n79) );
  INV_X1 npu_inst_pe_1_6_5_U38 ( .A(npu_inst_pe_1_6_5_n79), .ZN(
        npu_inst_pe_1_6_5_n35) );
  AOI222_X1 npu_inst_pe_1_6_5_U37 ( .A1(npu_inst_int_data_res_7__5__6_), .A2(
        npu_inst_pe_1_6_5_n1), .B1(npu_inst_pe_1_6_5_N79), .B2(
        npu_inst_pe_1_6_5_n76), .C1(npu_inst_pe_1_6_5_N71), .C2(
        npu_inst_pe_1_6_5_n77), .ZN(npu_inst_pe_1_6_5_n78) );
  INV_X1 npu_inst_pe_1_6_5_U36 ( .A(npu_inst_pe_1_6_5_n78), .ZN(
        npu_inst_pe_1_6_5_n34) );
  INV_X1 npu_inst_pe_1_6_5_U35 ( .A(npu_inst_pe_1_6_5_int_data_1_), .ZN(
        npu_inst_pe_1_6_5_n14) );
  AND2_X1 npu_inst_pe_1_6_5_U34 ( .A1(npu_inst_int_data_x_6__5__1_), .A2(
        npu_inst_pe_1_6_5_int_q_weight_1_), .ZN(npu_inst_pe_1_6_5_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_6_5_U33 ( .A1(npu_inst_int_data_x_6__5__0_), .A2(
        npu_inst_pe_1_6_5_int_q_weight_1_), .ZN(npu_inst_pe_1_6_5_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_6_5_U32 ( .A1(npu_inst_n53), .A2(
        npu_inst_int_data_y_7__5__1_), .B1(npu_inst_pe_1_6_5_n3), .B2(
        npu_inst_int_data_x_6__6__1_), .ZN(npu_inst_pe_1_6_5_n63) );
  AOI22_X1 npu_inst_pe_1_6_5_U31 ( .A1(npu_inst_n53), .A2(
        npu_inst_int_data_y_7__5__0_), .B1(npu_inst_pe_1_6_5_n3), .B2(
        npu_inst_int_data_x_6__6__0_), .ZN(npu_inst_pe_1_6_5_n61) );
  INV_X1 npu_inst_pe_1_6_5_U30 ( .A(npu_inst_pe_1_6_5_int_data_0_), .ZN(
        npu_inst_pe_1_6_5_n13) );
  INV_X1 npu_inst_pe_1_6_5_U29 ( .A(npu_inst_n67), .ZN(npu_inst_pe_1_6_5_n5)
         );
  OR3_X1 npu_inst_pe_1_6_5_U28 ( .A1(npu_inst_pe_1_6_5_n6), .A2(
        npu_inst_pe_1_6_5_n8), .A3(npu_inst_pe_1_6_5_n5), .ZN(
        npu_inst_pe_1_6_5_n56) );
  OR3_X1 npu_inst_pe_1_6_5_U27 ( .A1(npu_inst_pe_1_6_5_n5), .A2(
        npu_inst_pe_1_6_5_n8), .A3(npu_inst_pe_1_6_5_n7), .ZN(
        npu_inst_pe_1_6_5_n48) );
  INV_X1 npu_inst_pe_1_6_5_U26 ( .A(npu_inst_pe_1_6_5_n5), .ZN(
        npu_inst_pe_1_6_5_n4) );
  OR3_X1 npu_inst_pe_1_6_5_U25 ( .A1(npu_inst_pe_1_6_5_n4), .A2(
        npu_inst_pe_1_6_5_n8), .A3(npu_inst_pe_1_6_5_n7), .ZN(
        npu_inst_pe_1_6_5_n52) );
  OR3_X1 npu_inst_pe_1_6_5_U24 ( .A1(npu_inst_pe_1_6_5_n6), .A2(
        npu_inst_pe_1_6_5_n8), .A3(npu_inst_pe_1_6_5_n4), .ZN(
        npu_inst_pe_1_6_5_n60) );
  NOR2_X1 npu_inst_pe_1_6_5_U23 ( .A1(npu_inst_pe_1_6_5_n60), .A2(
        npu_inst_pe_1_6_5_n3), .ZN(npu_inst_pe_1_6_5_n58) );
  NOR2_X1 npu_inst_pe_1_6_5_U22 ( .A1(npu_inst_pe_1_6_5_n56), .A2(
        npu_inst_pe_1_6_5_n3), .ZN(npu_inst_pe_1_6_5_n54) );
  NOR2_X1 npu_inst_pe_1_6_5_U21 ( .A1(npu_inst_pe_1_6_5_n52), .A2(
        npu_inst_pe_1_6_5_n3), .ZN(npu_inst_pe_1_6_5_n50) );
  NOR2_X1 npu_inst_pe_1_6_5_U20 ( .A1(npu_inst_pe_1_6_5_n48), .A2(
        npu_inst_pe_1_6_5_n3), .ZN(npu_inst_pe_1_6_5_n46) );
  NOR2_X1 npu_inst_pe_1_6_5_U19 ( .A1(npu_inst_pe_1_6_5_n40), .A2(
        npu_inst_pe_1_6_5_n3), .ZN(npu_inst_pe_1_6_5_n38) );
  NOR2_X1 npu_inst_pe_1_6_5_U18 ( .A1(npu_inst_pe_1_6_5_n44), .A2(
        npu_inst_pe_1_6_5_n3), .ZN(npu_inst_pe_1_6_5_n42) );
  BUF_X1 npu_inst_pe_1_6_5_U17 ( .A(npu_inst_n94), .Z(npu_inst_pe_1_6_5_n8) );
  INV_X1 npu_inst_pe_1_6_5_U16 ( .A(npu_inst_n122), .ZN(npu_inst_pe_1_6_5_n12)
         );
  INV_X1 npu_inst_pe_1_6_5_U15 ( .A(npu_inst_pe_1_6_5_n38), .ZN(
        npu_inst_pe_1_6_5_n114) );
  INV_X1 npu_inst_pe_1_6_5_U14 ( .A(npu_inst_pe_1_6_5_n58), .ZN(
        npu_inst_pe_1_6_5_n119) );
  INV_X1 npu_inst_pe_1_6_5_U13 ( .A(npu_inst_pe_1_6_5_n54), .ZN(
        npu_inst_pe_1_6_5_n118) );
  INV_X1 npu_inst_pe_1_6_5_U12 ( .A(npu_inst_pe_1_6_5_n50), .ZN(
        npu_inst_pe_1_6_5_n117) );
  INV_X1 npu_inst_pe_1_6_5_U11 ( .A(npu_inst_pe_1_6_5_n46), .ZN(
        npu_inst_pe_1_6_5_n116) );
  INV_X1 npu_inst_pe_1_6_5_U10 ( .A(npu_inst_pe_1_6_5_n42), .ZN(
        npu_inst_pe_1_6_5_n115) );
  BUF_X1 npu_inst_pe_1_6_5_U9 ( .A(npu_inst_n12), .Z(npu_inst_pe_1_6_5_n2) );
  BUF_X1 npu_inst_pe_1_6_5_U8 ( .A(npu_inst_n12), .Z(npu_inst_pe_1_6_5_n1) );
  BUF_X1 npu_inst_pe_1_6_5_U7 ( .A(npu_inst_pe_1_6_5_n12), .Z(
        npu_inst_pe_1_6_5_n11) );
  BUF_X1 npu_inst_pe_1_6_5_U6 ( .A(npu_inst_pe_1_6_5_n12), .Z(
        npu_inst_pe_1_6_5_n10) );
  BUF_X1 npu_inst_pe_1_6_5_U5 ( .A(npu_inst_pe_1_6_5_n12), .Z(
        npu_inst_pe_1_6_5_n9) );
  NOR2_X1 npu_inst_pe_1_6_5_U4 ( .A1(npu_inst_pe_1_6_5_int_q_weight_0_), .A2(
        npu_inst_pe_1_6_5_n1), .ZN(npu_inst_pe_1_6_5_n76) );
  NOR2_X1 npu_inst_pe_1_6_5_U3 ( .A1(npu_inst_pe_1_6_5_n27), .A2(
        npu_inst_pe_1_6_5_n1), .ZN(npu_inst_pe_1_6_5_n77) );
  FA_X1 npu_inst_pe_1_6_5_sub_67_U2_1 ( .A(npu_inst_pe_1_6_5_int_q_acc_1_), 
        .B(npu_inst_pe_1_6_5_n14), .CI(npu_inst_pe_1_6_5_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_6_5_sub_67_carry_2_), .S(npu_inst_pe_1_6_5_N66) );
  FA_X1 npu_inst_pe_1_6_5_add_69_U1_1 ( .A(npu_inst_pe_1_6_5_int_q_acc_1_), 
        .B(npu_inst_pe_1_6_5_int_data_1_), .CI(
        npu_inst_pe_1_6_5_add_69_carry_1_), .CO(
        npu_inst_pe_1_6_5_add_69_carry_2_), .S(npu_inst_pe_1_6_5_N74) );
  NAND3_X1 npu_inst_pe_1_6_5_U109 ( .A1(npu_inst_pe_1_6_5_n5), .A2(
        npu_inst_pe_1_6_5_n7), .A3(npu_inst_pe_1_6_5_n8), .ZN(
        npu_inst_pe_1_6_5_n44) );
  NAND3_X1 npu_inst_pe_1_6_5_U108 ( .A1(npu_inst_pe_1_6_5_n4), .A2(
        npu_inst_pe_1_6_5_n7), .A3(npu_inst_pe_1_6_5_n8), .ZN(
        npu_inst_pe_1_6_5_n40) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_6_5_n34), .CK(
        npu_inst_pe_1_6_5_net3343), .RN(npu_inst_pe_1_6_5_n9), .Q(
        npu_inst_pe_1_6_5_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_6_5_n35), .CK(
        npu_inst_pe_1_6_5_net3343), .RN(npu_inst_pe_1_6_5_n9), .Q(
        npu_inst_pe_1_6_5_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_6_5_n36), .CK(
        npu_inst_pe_1_6_5_net3343), .RN(npu_inst_pe_1_6_5_n9), .Q(
        npu_inst_pe_1_6_5_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_6_5_n98), .CK(
        npu_inst_pe_1_6_5_net3343), .RN(npu_inst_pe_1_6_5_n9), .Q(
        npu_inst_pe_1_6_5_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_6_5_n99), .CK(
        npu_inst_pe_1_6_5_net3343), .RN(npu_inst_pe_1_6_5_n9), .Q(
        npu_inst_pe_1_6_5_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_6_5_n100), 
        .CK(npu_inst_pe_1_6_5_net3343), .RN(npu_inst_pe_1_6_5_n9), .Q(
        npu_inst_pe_1_6_5_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_6_5_n33), .CK(
        npu_inst_pe_1_6_5_net3343), .RN(npu_inst_pe_1_6_5_n9), .Q(
        npu_inst_pe_1_6_5_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_6_5_n101), 
        .CK(npu_inst_pe_1_6_5_net3343), .RN(npu_inst_pe_1_6_5_n9), .Q(
        npu_inst_pe_1_6_5_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_weight_reg_0_ ( .D(npu_inst_n108), .CK(
        npu_inst_pe_1_6_5_net3349), .RN(npu_inst_pe_1_6_5_n9), .Q(
        npu_inst_pe_1_6_5_int_q_weight_0_), .QN(npu_inst_pe_1_6_5_n27) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_weight_reg_1_ ( .D(npu_inst_n114), .CK(
        npu_inst_pe_1_6_5_net3349), .RN(npu_inst_pe_1_6_5_n9), .Q(
        npu_inst_pe_1_6_5_int_q_weight_1_), .QN(npu_inst_pe_1_6_5_n26) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_6_5_n113), 
        .CK(npu_inst_pe_1_6_5_net3349), .RN(npu_inst_pe_1_6_5_n9), .Q(
        npu_inst_pe_1_6_5_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_6_5_n107), 
        .CK(npu_inst_pe_1_6_5_net3349), .RN(npu_inst_pe_1_6_5_n9), .Q(
        npu_inst_pe_1_6_5_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_6_5_n112), 
        .CK(npu_inst_pe_1_6_5_net3349), .RN(npu_inst_pe_1_6_5_n10), .Q(
        npu_inst_pe_1_6_5_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_6_5_n106), 
        .CK(npu_inst_pe_1_6_5_net3349), .RN(npu_inst_pe_1_6_5_n10), .Q(
        npu_inst_pe_1_6_5_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_6_5_n111), 
        .CK(npu_inst_pe_1_6_5_net3349), .RN(npu_inst_pe_1_6_5_n10), .Q(
        npu_inst_pe_1_6_5_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_6_5_n105), 
        .CK(npu_inst_pe_1_6_5_net3349), .RN(npu_inst_pe_1_6_5_n10), .Q(
        npu_inst_pe_1_6_5_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_6_5_n110), 
        .CK(npu_inst_pe_1_6_5_net3349), .RN(npu_inst_pe_1_6_5_n10), .Q(
        npu_inst_pe_1_6_5_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_6_5_n104), 
        .CK(npu_inst_pe_1_6_5_net3349), .RN(npu_inst_pe_1_6_5_n10), .Q(
        npu_inst_pe_1_6_5_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_6_5_n109), 
        .CK(npu_inst_pe_1_6_5_net3349), .RN(npu_inst_pe_1_6_5_n10), .Q(
        npu_inst_pe_1_6_5_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_6_5_n103), 
        .CK(npu_inst_pe_1_6_5_net3349), .RN(npu_inst_pe_1_6_5_n10), .Q(
        npu_inst_pe_1_6_5_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_6_5_n108), 
        .CK(npu_inst_pe_1_6_5_net3349), .RN(npu_inst_pe_1_6_5_n10), .Q(
        npu_inst_pe_1_6_5_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_6_5_n102), 
        .CK(npu_inst_pe_1_6_5_net3349), .RN(npu_inst_pe_1_6_5_n10), .Q(
        npu_inst_pe_1_6_5_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_6_5_n86), 
        .CK(npu_inst_pe_1_6_5_net3349), .RN(npu_inst_pe_1_6_5_n10), .Q(
        npu_inst_pe_1_6_5_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_6_5_n87), 
        .CK(npu_inst_pe_1_6_5_net3349), .RN(npu_inst_pe_1_6_5_n10), .Q(
        npu_inst_pe_1_6_5_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_6_5_n88), 
        .CK(npu_inst_pe_1_6_5_net3349), .RN(npu_inst_pe_1_6_5_n11), .Q(
        npu_inst_pe_1_6_5_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_6_5_n89), 
        .CK(npu_inst_pe_1_6_5_net3349), .RN(npu_inst_pe_1_6_5_n11), .Q(
        npu_inst_pe_1_6_5_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_6_5_n90), 
        .CK(npu_inst_pe_1_6_5_net3349), .RN(npu_inst_pe_1_6_5_n11), .Q(
        npu_inst_pe_1_6_5_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_6_5_n91), 
        .CK(npu_inst_pe_1_6_5_net3349), .RN(npu_inst_pe_1_6_5_n11), .Q(
        npu_inst_pe_1_6_5_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_6_5_n92), 
        .CK(npu_inst_pe_1_6_5_net3349), .RN(npu_inst_pe_1_6_5_n11), .Q(
        npu_inst_pe_1_6_5_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_6_5_n93), 
        .CK(npu_inst_pe_1_6_5_net3349), .RN(npu_inst_pe_1_6_5_n11), .Q(
        npu_inst_pe_1_6_5_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_6_5_n94), 
        .CK(npu_inst_pe_1_6_5_net3349), .RN(npu_inst_pe_1_6_5_n11), .Q(
        npu_inst_pe_1_6_5_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_6_5_n95), 
        .CK(npu_inst_pe_1_6_5_net3349), .RN(npu_inst_pe_1_6_5_n11), .Q(
        npu_inst_pe_1_6_5_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_6_5_n96), 
        .CK(npu_inst_pe_1_6_5_net3349), .RN(npu_inst_pe_1_6_5_n11), .Q(
        npu_inst_pe_1_6_5_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_6_5_n97), 
        .CK(npu_inst_pe_1_6_5_net3349), .RN(npu_inst_pe_1_6_5_n11), .Q(
        npu_inst_pe_1_6_5_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_6_5_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_6_5_N84), .SE(1'b0), .GCK(npu_inst_pe_1_6_5_net3343) );
  CLKGATETST_X1 npu_inst_pe_1_6_5_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n61), .SE(1'b0), .GCK(npu_inst_pe_1_6_5_net3349) );
  MUX2_X1 npu_inst_pe_1_6_6_U162 ( .A(npu_inst_pe_1_6_6_n32), .B(
        npu_inst_pe_1_6_6_n29), .S(npu_inst_pe_1_6_6_n8), .Z(
        npu_inst_pe_1_6_6_N93) );
  MUX2_X1 npu_inst_pe_1_6_6_U161 ( .A(npu_inst_pe_1_6_6_n31), .B(
        npu_inst_pe_1_6_6_n30), .S(npu_inst_pe_1_6_6_n6), .Z(
        npu_inst_pe_1_6_6_n32) );
  MUX2_X1 npu_inst_pe_1_6_6_U160 ( .A(npu_inst_pe_1_6_6_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_6_6_int_q_reg_v_1__0_), .S(npu_inst_pe_1_6_6_n4), .Z(
        npu_inst_pe_1_6_6_n31) );
  MUX2_X1 npu_inst_pe_1_6_6_U159 ( .A(npu_inst_pe_1_6_6_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_6_6_int_q_reg_v_3__0_), .S(npu_inst_pe_1_6_6_n4), .Z(
        npu_inst_pe_1_6_6_n30) );
  MUX2_X1 npu_inst_pe_1_6_6_U158 ( .A(npu_inst_pe_1_6_6_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_6_6_int_q_reg_v_5__0_), .S(npu_inst_pe_1_6_6_n4), .Z(
        npu_inst_pe_1_6_6_n29) );
  MUX2_X1 npu_inst_pe_1_6_6_U157 ( .A(npu_inst_pe_1_6_6_n28), .B(
        npu_inst_pe_1_6_6_n23), .S(npu_inst_pe_1_6_6_n8), .Z(
        npu_inst_pe_1_6_6_N94) );
  MUX2_X1 npu_inst_pe_1_6_6_U156 ( .A(npu_inst_pe_1_6_6_n25), .B(
        npu_inst_pe_1_6_6_n24), .S(npu_inst_pe_1_6_6_n6), .Z(
        npu_inst_pe_1_6_6_n28) );
  MUX2_X1 npu_inst_pe_1_6_6_U155 ( .A(npu_inst_pe_1_6_6_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_6_6_int_q_reg_v_1__1_), .S(npu_inst_pe_1_6_6_n4), .Z(
        npu_inst_pe_1_6_6_n25) );
  MUX2_X1 npu_inst_pe_1_6_6_U154 ( .A(npu_inst_pe_1_6_6_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_6_6_int_q_reg_v_3__1_), .S(npu_inst_pe_1_6_6_n4), .Z(
        npu_inst_pe_1_6_6_n24) );
  MUX2_X1 npu_inst_pe_1_6_6_U153 ( .A(npu_inst_pe_1_6_6_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_6_6_int_q_reg_v_5__1_), .S(npu_inst_pe_1_6_6_n4), .Z(
        npu_inst_pe_1_6_6_n23) );
  MUX2_X1 npu_inst_pe_1_6_6_U152 ( .A(npu_inst_pe_1_6_6_n22), .B(
        npu_inst_pe_1_6_6_n19), .S(npu_inst_pe_1_6_6_n8), .Z(
        npu_inst_int_data_x_6__6__1_) );
  MUX2_X1 npu_inst_pe_1_6_6_U151 ( .A(npu_inst_pe_1_6_6_n21), .B(
        npu_inst_pe_1_6_6_n20), .S(npu_inst_pe_1_6_6_n6), .Z(
        npu_inst_pe_1_6_6_n22) );
  MUX2_X1 npu_inst_pe_1_6_6_U150 ( .A(npu_inst_pe_1_6_6_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_6_6_int_q_reg_h_1__1_), .S(npu_inst_pe_1_6_6_n4), .Z(
        npu_inst_pe_1_6_6_n21) );
  MUX2_X1 npu_inst_pe_1_6_6_U149 ( .A(npu_inst_pe_1_6_6_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_6_6_int_q_reg_h_3__1_), .S(npu_inst_pe_1_6_6_n4), .Z(
        npu_inst_pe_1_6_6_n20) );
  MUX2_X1 npu_inst_pe_1_6_6_U148 ( .A(npu_inst_pe_1_6_6_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_6_6_int_q_reg_h_5__1_), .S(npu_inst_pe_1_6_6_n4), .Z(
        npu_inst_pe_1_6_6_n19) );
  MUX2_X1 npu_inst_pe_1_6_6_U147 ( .A(npu_inst_pe_1_6_6_n18), .B(
        npu_inst_pe_1_6_6_n15), .S(npu_inst_pe_1_6_6_n8), .Z(
        npu_inst_int_data_x_6__6__0_) );
  MUX2_X1 npu_inst_pe_1_6_6_U146 ( .A(npu_inst_pe_1_6_6_n17), .B(
        npu_inst_pe_1_6_6_n16), .S(npu_inst_pe_1_6_6_n6), .Z(
        npu_inst_pe_1_6_6_n18) );
  MUX2_X1 npu_inst_pe_1_6_6_U145 ( .A(npu_inst_pe_1_6_6_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_6_6_int_q_reg_h_1__0_), .S(npu_inst_pe_1_6_6_n4), .Z(
        npu_inst_pe_1_6_6_n17) );
  MUX2_X1 npu_inst_pe_1_6_6_U144 ( .A(npu_inst_pe_1_6_6_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_6_6_int_q_reg_h_3__0_), .S(npu_inst_pe_1_6_6_n4), .Z(
        npu_inst_pe_1_6_6_n16) );
  MUX2_X1 npu_inst_pe_1_6_6_U143 ( .A(npu_inst_pe_1_6_6_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_6_6_int_q_reg_h_5__0_), .S(npu_inst_pe_1_6_6_n4), .Z(
        npu_inst_pe_1_6_6_n15) );
  XOR2_X1 npu_inst_pe_1_6_6_U142 ( .A(npu_inst_pe_1_6_6_int_data_0_), .B(
        npu_inst_pe_1_6_6_int_q_acc_0_), .Z(npu_inst_pe_1_6_6_N73) );
  AND2_X1 npu_inst_pe_1_6_6_U141 ( .A1(npu_inst_pe_1_6_6_int_q_acc_0_), .A2(
        npu_inst_pe_1_6_6_int_data_0_), .ZN(npu_inst_pe_1_6_6_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_6_6_U140 ( .A(npu_inst_pe_1_6_6_int_q_acc_0_), .B(
        npu_inst_pe_1_6_6_n13), .ZN(npu_inst_pe_1_6_6_N65) );
  OR2_X1 npu_inst_pe_1_6_6_U139 ( .A1(npu_inst_pe_1_6_6_n13), .A2(
        npu_inst_pe_1_6_6_int_q_acc_0_), .ZN(npu_inst_pe_1_6_6_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_6_6_U138 ( .A(npu_inst_pe_1_6_6_int_q_acc_2_), .B(
        npu_inst_pe_1_6_6_add_69_carry_2_), .Z(npu_inst_pe_1_6_6_N75) );
  AND2_X1 npu_inst_pe_1_6_6_U137 ( .A1(npu_inst_pe_1_6_6_add_69_carry_2_), 
        .A2(npu_inst_pe_1_6_6_int_q_acc_2_), .ZN(
        npu_inst_pe_1_6_6_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_6_6_U136 ( .A(npu_inst_pe_1_6_6_int_q_acc_3_), .B(
        npu_inst_pe_1_6_6_add_69_carry_3_), .Z(npu_inst_pe_1_6_6_N76) );
  AND2_X1 npu_inst_pe_1_6_6_U135 ( .A1(npu_inst_pe_1_6_6_add_69_carry_3_), 
        .A2(npu_inst_pe_1_6_6_int_q_acc_3_), .ZN(
        npu_inst_pe_1_6_6_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_6_6_U134 ( .A(npu_inst_pe_1_6_6_int_q_acc_4_), .B(
        npu_inst_pe_1_6_6_add_69_carry_4_), .Z(npu_inst_pe_1_6_6_N77) );
  AND2_X1 npu_inst_pe_1_6_6_U133 ( .A1(npu_inst_pe_1_6_6_add_69_carry_4_), 
        .A2(npu_inst_pe_1_6_6_int_q_acc_4_), .ZN(
        npu_inst_pe_1_6_6_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_6_6_U132 ( .A(npu_inst_pe_1_6_6_int_q_acc_5_), .B(
        npu_inst_pe_1_6_6_add_69_carry_5_), .Z(npu_inst_pe_1_6_6_N78) );
  AND2_X1 npu_inst_pe_1_6_6_U131 ( .A1(npu_inst_pe_1_6_6_add_69_carry_5_), 
        .A2(npu_inst_pe_1_6_6_int_q_acc_5_), .ZN(
        npu_inst_pe_1_6_6_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_6_6_U130 ( .A(npu_inst_pe_1_6_6_int_q_acc_6_), .B(
        npu_inst_pe_1_6_6_add_69_carry_6_), .Z(npu_inst_pe_1_6_6_N79) );
  AND2_X1 npu_inst_pe_1_6_6_U129 ( .A1(npu_inst_pe_1_6_6_add_69_carry_6_), 
        .A2(npu_inst_pe_1_6_6_int_q_acc_6_), .ZN(
        npu_inst_pe_1_6_6_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_6_6_U128 ( .A(npu_inst_pe_1_6_6_int_q_acc_7_), .B(
        npu_inst_pe_1_6_6_add_69_carry_7_), .Z(npu_inst_pe_1_6_6_N80) );
  XNOR2_X1 npu_inst_pe_1_6_6_U127 ( .A(npu_inst_pe_1_6_6_sub_67_carry_2_), .B(
        npu_inst_pe_1_6_6_int_q_acc_2_), .ZN(npu_inst_pe_1_6_6_N67) );
  OR2_X1 npu_inst_pe_1_6_6_U126 ( .A1(npu_inst_pe_1_6_6_int_q_acc_2_), .A2(
        npu_inst_pe_1_6_6_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_6_6_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_6_6_U125 ( .A(npu_inst_pe_1_6_6_sub_67_carry_3_), .B(
        npu_inst_pe_1_6_6_int_q_acc_3_), .ZN(npu_inst_pe_1_6_6_N68) );
  OR2_X1 npu_inst_pe_1_6_6_U124 ( .A1(npu_inst_pe_1_6_6_int_q_acc_3_), .A2(
        npu_inst_pe_1_6_6_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_6_6_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_6_6_U123 ( .A(npu_inst_pe_1_6_6_sub_67_carry_4_), .B(
        npu_inst_pe_1_6_6_int_q_acc_4_), .ZN(npu_inst_pe_1_6_6_N69) );
  OR2_X1 npu_inst_pe_1_6_6_U122 ( .A1(npu_inst_pe_1_6_6_int_q_acc_4_), .A2(
        npu_inst_pe_1_6_6_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_6_6_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_6_6_U121 ( .A(npu_inst_pe_1_6_6_sub_67_carry_5_), .B(
        npu_inst_pe_1_6_6_int_q_acc_5_), .ZN(npu_inst_pe_1_6_6_N70) );
  OR2_X1 npu_inst_pe_1_6_6_U120 ( .A1(npu_inst_pe_1_6_6_int_q_acc_5_), .A2(
        npu_inst_pe_1_6_6_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_6_6_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_6_6_U119 ( .A(npu_inst_pe_1_6_6_sub_67_carry_6_), .B(
        npu_inst_pe_1_6_6_int_q_acc_6_), .ZN(npu_inst_pe_1_6_6_N71) );
  OR2_X1 npu_inst_pe_1_6_6_U118 ( .A1(npu_inst_pe_1_6_6_int_q_acc_6_), .A2(
        npu_inst_pe_1_6_6_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_6_6_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_6_6_U117 ( .A(npu_inst_pe_1_6_6_int_q_acc_7_), .B(
        npu_inst_pe_1_6_6_sub_67_carry_7_), .ZN(npu_inst_pe_1_6_6_N72) );
  INV_X1 npu_inst_pe_1_6_6_U116 ( .A(npu_inst_n75), .ZN(npu_inst_pe_1_6_6_n7)
         );
  INV_X1 npu_inst_pe_1_6_6_U115 ( .A(npu_inst_pe_1_6_6_n7), .ZN(
        npu_inst_pe_1_6_6_n6) );
  INV_X1 npu_inst_pe_1_6_6_U114 ( .A(npu_inst_n53), .ZN(npu_inst_pe_1_6_6_n3)
         );
  AOI22_X1 npu_inst_pe_1_6_6_U113 ( .A1(npu_inst_int_data_y_7__6__0_), .A2(
        npu_inst_pe_1_6_6_n58), .B1(npu_inst_pe_1_6_6_n119), .B2(
        npu_inst_pe_1_6_6_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_6_6_n57) );
  INV_X1 npu_inst_pe_1_6_6_U112 ( .A(npu_inst_pe_1_6_6_n57), .ZN(
        npu_inst_pe_1_6_6_n108) );
  AOI22_X1 npu_inst_pe_1_6_6_U111 ( .A1(npu_inst_int_data_y_7__6__0_), .A2(
        npu_inst_pe_1_6_6_n54), .B1(npu_inst_pe_1_6_6_n118), .B2(
        npu_inst_pe_1_6_6_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_6_6_n53) );
  INV_X1 npu_inst_pe_1_6_6_U110 ( .A(npu_inst_pe_1_6_6_n53), .ZN(
        npu_inst_pe_1_6_6_n109) );
  AOI22_X1 npu_inst_pe_1_6_6_U107 ( .A1(npu_inst_int_data_y_7__6__0_), .A2(
        npu_inst_pe_1_6_6_n50), .B1(npu_inst_pe_1_6_6_n117), .B2(
        npu_inst_pe_1_6_6_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_6_6_n49) );
  INV_X1 npu_inst_pe_1_6_6_U106 ( .A(npu_inst_pe_1_6_6_n49), .ZN(
        npu_inst_pe_1_6_6_n110) );
  AOI22_X1 npu_inst_pe_1_6_6_U105 ( .A1(npu_inst_int_data_y_7__6__0_), .A2(
        npu_inst_pe_1_6_6_n46), .B1(npu_inst_pe_1_6_6_n116), .B2(
        npu_inst_pe_1_6_6_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_6_6_n45) );
  INV_X1 npu_inst_pe_1_6_6_U104 ( .A(npu_inst_pe_1_6_6_n45), .ZN(
        npu_inst_pe_1_6_6_n111) );
  AOI22_X1 npu_inst_pe_1_6_6_U103 ( .A1(npu_inst_int_data_y_7__6__0_), .A2(
        npu_inst_pe_1_6_6_n42), .B1(npu_inst_pe_1_6_6_n115), .B2(
        npu_inst_pe_1_6_6_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_6_6_n41) );
  INV_X1 npu_inst_pe_1_6_6_U102 ( .A(npu_inst_pe_1_6_6_n41), .ZN(
        npu_inst_pe_1_6_6_n112) );
  AOI22_X1 npu_inst_pe_1_6_6_U101 ( .A1(npu_inst_int_data_y_7__6__1_), .A2(
        npu_inst_pe_1_6_6_n58), .B1(npu_inst_pe_1_6_6_n119), .B2(
        npu_inst_pe_1_6_6_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_6_6_n59) );
  INV_X1 npu_inst_pe_1_6_6_U100 ( .A(npu_inst_pe_1_6_6_n59), .ZN(
        npu_inst_pe_1_6_6_n102) );
  AOI22_X1 npu_inst_pe_1_6_6_U99 ( .A1(npu_inst_int_data_y_7__6__1_), .A2(
        npu_inst_pe_1_6_6_n54), .B1(npu_inst_pe_1_6_6_n118), .B2(
        npu_inst_pe_1_6_6_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_6_6_n55) );
  INV_X1 npu_inst_pe_1_6_6_U98 ( .A(npu_inst_pe_1_6_6_n55), .ZN(
        npu_inst_pe_1_6_6_n103) );
  AOI22_X1 npu_inst_pe_1_6_6_U97 ( .A1(npu_inst_int_data_y_7__6__1_), .A2(
        npu_inst_pe_1_6_6_n50), .B1(npu_inst_pe_1_6_6_n117), .B2(
        npu_inst_pe_1_6_6_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_6_6_n51) );
  INV_X1 npu_inst_pe_1_6_6_U96 ( .A(npu_inst_pe_1_6_6_n51), .ZN(
        npu_inst_pe_1_6_6_n104) );
  AOI22_X1 npu_inst_pe_1_6_6_U95 ( .A1(npu_inst_int_data_y_7__6__1_), .A2(
        npu_inst_pe_1_6_6_n46), .B1(npu_inst_pe_1_6_6_n116), .B2(
        npu_inst_pe_1_6_6_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_6_6_n47) );
  INV_X1 npu_inst_pe_1_6_6_U94 ( .A(npu_inst_pe_1_6_6_n47), .ZN(
        npu_inst_pe_1_6_6_n105) );
  AOI22_X1 npu_inst_pe_1_6_6_U93 ( .A1(npu_inst_int_data_y_7__6__1_), .A2(
        npu_inst_pe_1_6_6_n42), .B1(npu_inst_pe_1_6_6_n115), .B2(
        npu_inst_pe_1_6_6_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_6_6_n43) );
  INV_X1 npu_inst_pe_1_6_6_U92 ( .A(npu_inst_pe_1_6_6_n43), .ZN(
        npu_inst_pe_1_6_6_n106) );
  AOI22_X1 npu_inst_pe_1_6_6_U91 ( .A1(npu_inst_pe_1_6_6_n38), .A2(
        npu_inst_int_data_y_7__6__1_), .B1(npu_inst_pe_1_6_6_n114), .B2(
        npu_inst_pe_1_6_6_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_6_6_n39) );
  INV_X1 npu_inst_pe_1_6_6_U90 ( .A(npu_inst_pe_1_6_6_n39), .ZN(
        npu_inst_pe_1_6_6_n107) );
  AOI22_X1 npu_inst_pe_1_6_6_U89 ( .A1(npu_inst_pe_1_6_6_n38), .A2(
        npu_inst_int_data_y_7__6__0_), .B1(npu_inst_pe_1_6_6_n114), .B2(
        npu_inst_pe_1_6_6_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_6_6_n37) );
  INV_X1 npu_inst_pe_1_6_6_U88 ( .A(npu_inst_pe_1_6_6_n37), .ZN(
        npu_inst_pe_1_6_6_n113) );
  NAND2_X1 npu_inst_pe_1_6_6_U87 ( .A1(npu_inst_pe_1_6_6_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_6_6_n60), .ZN(npu_inst_pe_1_6_6_n74) );
  OAI21_X1 npu_inst_pe_1_6_6_U86 ( .B1(npu_inst_pe_1_6_6_n63), .B2(
        npu_inst_pe_1_6_6_n60), .A(npu_inst_pe_1_6_6_n74), .ZN(
        npu_inst_pe_1_6_6_n97) );
  NAND2_X1 npu_inst_pe_1_6_6_U85 ( .A1(npu_inst_pe_1_6_6_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_6_6_n60), .ZN(npu_inst_pe_1_6_6_n73) );
  OAI21_X1 npu_inst_pe_1_6_6_U84 ( .B1(npu_inst_pe_1_6_6_n61), .B2(
        npu_inst_pe_1_6_6_n60), .A(npu_inst_pe_1_6_6_n73), .ZN(
        npu_inst_pe_1_6_6_n96) );
  NAND2_X1 npu_inst_pe_1_6_6_U83 ( .A1(npu_inst_pe_1_6_6_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_6_6_n56), .ZN(npu_inst_pe_1_6_6_n72) );
  OAI21_X1 npu_inst_pe_1_6_6_U82 ( .B1(npu_inst_pe_1_6_6_n63), .B2(
        npu_inst_pe_1_6_6_n56), .A(npu_inst_pe_1_6_6_n72), .ZN(
        npu_inst_pe_1_6_6_n95) );
  NAND2_X1 npu_inst_pe_1_6_6_U81 ( .A1(npu_inst_pe_1_6_6_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_6_6_n56), .ZN(npu_inst_pe_1_6_6_n71) );
  OAI21_X1 npu_inst_pe_1_6_6_U80 ( .B1(npu_inst_pe_1_6_6_n61), .B2(
        npu_inst_pe_1_6_6_n56), .A(npu_inst_pe_1_6_6_n71), .ZN(
        npu_inst_pe_1_6_6_n94) );
  NAND2_X1 npu_inst_pe_1_6_6_U79 ( .A1(npu_inst_pe_1_6_6_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_6_6_n52), .ZN(npu_inst_pe_1_6_6_n70) );
  OAI21_X1 npu_inst_pe_1_6_6_U78 ( .B1(npu_inst_pe_1_6_6_n63), .B2(
        npu_inst_pe_1_6_6_n52), .A(npu_inst_pe_1_6_6_n70), .ZN(
        npu_inst_pe_1_6_6_n93) );
  NAND2_X1 npu_inst_pe_1_6_6_U77 ( .A1(npu_inst_pe_1_6_6_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_6_6_n52), .ZN(npu_inst_pe_1_6_6_n69) );
  OAI21_X1 npu_inst_pe_1_6_6_U76 ( .B1(npu_inst_pe_1_6_6_n61), .B2(
        npu_inst_pe_1_6_6_n52), .A(npu_inst_pe_1_6_6_n69), .ZN(
        npu_inst_pe_1_6_6_n92) );
  NAND2_X1 npu_inst_pe_1_6_6_U75 ( .A1(npu_inst_pe_1_6_6_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_6_6_n48), .ZN(npu_inst_pe_1_6_6_n68) );
  OAI21_X1 npu_inst_pe_1_6_6_U74 ( .B1(npu_inst_pe_1_6_6_n63), .B2(
        npu_inst_pe_1_6_6_n48), .A(npu_inst_pe_1_6_6_n68), .ZN(
        npu_inst_pe_1_6_6_n91) );
  NAND2_X1 npu_inst_pe_1_6_6_U73 ( .A1(npu_inst_pe_1_6_6_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_6_6_n48), .ZN(npu_inst_pe_1_6_6_n67) );
  OAI21_X1 npu_inst_pe_1_6_6_U72 ( .B1(npu_inst_pe_1_6_6_n61), .B2(
        npu_inst_pe_1_6_6_n48), .A(npu_inst_pe_1_6_6_n67), .ZN(
        npu_inst_pe_1_6_6_n90) );
  NAND2_X1 npu_inst_pe_1_6_6_U71 ( .A1(npu_inst_pe_1_6_6_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_6_6_n44), .ZN(npu_inst_pe_1_6_6_n66) );
  OAI21_X1 npu_inst_pe_1_6_6_U70 ( .B1(npu_inst_pe_1_6_6_n63), .B2(
        npu_inst_pe_1_6_6_n44), .A(npu_inst_pe_1_6_6_n66), .ZN(
        npu_inst_pe_1_6_6_n89) );
  NAND2_X1 npu_inst_pe_1_6_6_U69 ( .A1(npu_inst_pe_1_6_6_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_6_6_n44), .ZN(npu_inst_pe_1_6_6_n65) );
  OAI21_X1 npu_inst_pe_1_6_6_U68 ( .B1(npu_inst_pe_1_6_6_n61), .B2(
        npu_inst_pe_1_6_6_n44), .A(npu_inst_pe_1_6_6_n65), .ZN(
        npu_inst_pe_1_6_6_n88) );
  NAND2_X1 npu_inst_pe_1_6_6_U67 ( .A1(npu_inst_pe_1_6_6_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_6_6_n40), .ZN(npu_inst_pe_1_6_6_n64) );
  OAI21_X1 npu_inst_pe_1_6_6_U66 ( .B1(npu_inst_pe_1_6_6_n63), .B2(
        npu_inst_pe_1_6_6_n40), .A(npu_inst_pe_1_6_6_n64), .ZN(
        npu_inst_pe_1_6_6_n87) );
  NAND2_X1 npu_inst_pe_1_6_6_U65 ( .A1(npu_inst_pe_1_6_6_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_6_6_n40), .ZN(npu_inst_pe_1_6_6_n62) );
  OAI21_X1 npu_inst_pe_1_6_6_U64 ( .B1(npu_inst_pe_1_6_6_n61), .B2(
        npu_inst_pe_1_6_6_n40), .A(npu_inst_pe_1_6_6_n62), .ZN(
        npu_inst_pe_1_6_6_n86) );
  AND2_X1 npu_inst_pe_1_6_6_U63 ( .A1(npu_inst_pe_1_6_6_N93), .A2(npu_inst_n53), .ZN(npu_inst_int_data_y_6__6__0_) );
  AND2_X1 npu_inst_pe_1_6_6_U62 ( .A1(npu_inst_n53), .A2(npu_inst_pe_1_6_6_N94), .ZN(npu_inst_int_data_y_6__6__1_) );
  NOR3_X1 npu_inst_pe_1_6_6_U61 ( .A1(npu_inst_pe_1_6_6_n26), .A2(npu_inst_n53), .A3(npu_inst_int_ckg[9]), .ZN(npu_inst_pe_1_6_6_n85) );
  OR2_X1 npu_inst_pe_1_6_6_U60 ( .A1(npu_inst_pe_1_6_6_n85), .A2(
        npu_inst_pe_1_6_6_n2), .ZN(npu_inst_pe_1_6_6_N84) );
  AND2_X1 npu_inst_pe_1_6_6_U59 ( .A1(npu_inst_pe_1_6_6_int_q_acc_0_), .A2(
        npu_inst_pe_1_6_6_n1), .ZN(npu_inst_int_data_res_6__6__0_) );
  AND2_X1 npu_inst_pe_1_6_6_U58 ( .A1(npu_inst_pe_1_6_6_n2), .A2(
        npu_inst_pe_1_6_6_int_q_acc_7_), .ZN(npu_inst_int_data_res_6__6__7_)
         );
  AND2_X1 npu_inst_pe_1_6_6_U57 ( .A1(npu_inst_pe_1_6_6_int_q_acc_1_), .A2(
        npu_inst_pe_1_6_6_n1), .ZN(npu_inst_int_data_res_6__6__1_) );
  AND2_X1 npu_inst_pe_1_6_6_U56 ( .A1(npu_inst_pe_1_6_6_int_q_acc_2_), .A2(
        npu_inst_pe_1_6_6_n1), .ZN(npu_inst_int_data_res_6__6__2_) );
  AND2_X1 npu_inst_pe_1_6_6_U55 ( .A1(npu_inst_pe_1_6_6_int_q_acc_3_), .A2(
        npu_inst_pe_1_6_6_n2), .ZN(npu_inst_int_data_res_6__6__3_) );
  AND2_X1 npu_inst_pe_1_6_6_U54 ( .A1(npu_inst_pe_1_6_6_int_q_acc_4_), .A2(
        npu_inst_pe_1_6_6_n2), .ZN(npu_inst_int_data_res_6__6__4_) );
  AND2_X1 npu_inst_pe_1_6_6_U53 ( .A1(npu_inst_pe_1_6_6_int_q_acc_5_), .A2(
        npu_inst_pe_1_6_6_n2), .ZN(npu_inst_int_data_res_6__6__5_) );
  AND2_X1 npu_inst_pe_1_6_6_U52 ( .A1(npu_inst_pe_1_6_6_int_q_acc_6_), .A2(
        npu_inst_pe_1_6_6_n2), .ZN(npu_inst_int_data_res_6__6__6_) );
  AOI222_X1 npu_inst_pe_1_6_6_U51 ( .A1(npu_inst_int_data_res_7__6__0_), .A2(
        npu_inst_pe_1_6_6_n1), .B1(npu_inst_pe_1_6_6_N73), .B2(
        npu_inst_pe_1_6_6_n76), .C1(npu_inst_pe_1_6_6_N65), .C2(
        npu_inst_pe_1_6_6_n77), .ZN(npu_inst_pe_1_6_6_n84) );
  INV_X1 npu_inst_pe_1_6_6_U50 ( .A(npu_inst_pe_1_6_6_n84), .ZN(
        npu_inst_pe_1_6_6_n101) );
  AOI222_X1 npu_inst_pe_1_6_6_U49 ( .A1(npu_inst_int_data_res_7__6__7_), .A2(
        npu_inst_pe_1_6_6_n1), .B1(npu_inst_pe_1_6_6_N80), .B2(
        npu_inst_pe_1_6_6_n76), .C1(npu_inst_pe_1_6_6_N72), .C2(
        npu_inst_pe_1_6_6_n77), .ZN(npu_inst_pe_1_6_6_n75) );
  INV_X1 npu_inst_pe_1_6_6_U48 ( .A(npu_inst_pe_1_6_6_n75), .ZN(
        npu_inst_pe_1_6_6_n33) );
  AOI222_X1 npu_inst_pe_1_6_6_U47 ( .A1(npu_inst_int_data_res_7__6__1_), .A2(
        npu_inst_pe_1_6_6_n1), .B1(npu_inst_pe_1_6_6_N74), .B2(
        npu_inst_pe_1_6_6_n76), .C1(npu_inst_pe_1_6_6_N66), .C2(
        npu_inst_pe_1_6_6_n77), .ZN(npu_inst_pe_1_6_6_n83) );
  INV_X1 npu_inst_pe_1_6_6_U46 ( .A(npu_inst_pe_1_6_6_n83), .ZN(
        npu_inst_pe_1_6_6_n100) );
  AOI222_X1 npu_inst_pe_1_6_6_U45 ( .A1(npu_inst_int_data_res_7__6__2_), .A2(
        npu_inst_pe_1_6_6_n1), .B1(npu_inst_pe_1_6_6_N75), .B2(
        npu_inst_pe_1_6_6_n76), .C1(npu_inst_pe_1_6_6_N67), .C2(
        npu_inst_pe_1_6_6_n77), .ZN(npu_inst_pe_1_6_6_n82) );
  INV_X1 npu_inst_pe_1_6_6_U44 ( .A(npu_inst_pe_1_6_6_n82), .ZN(
        npu_inst_pe_1_6_6_n99) );
  AOI222_X1 npu_inst_pe_1_6_6_U43 ( .A1(npu_inst_int_data_res_7__6__3_), .A2(
        npu_inst_pe_1_6_6_n1), .B1(npu_inst_pe_1_6_6_N76), .B2(
        npu_inst_pe_1_6_6_n76), .C1(npu_inst_pe_1_6_6_N68), .C2(
        npu_inst_pe_1_6_6_n77), .ZN(npu_inst_pe_1_6_6_n81) );
  INV_X1 npu_inst_pe_1_6_6_U42 ( .A(npu_inst_pe_1_6_6_n81), .ZN(
        npu_inst_pe_1_6_6_n98) );
  AOI222_X1 npu_inst_pe_1_6_6_U41 ( .A1(npu_inst_int_data_res_7__6__4_), .A2(
        npu_inst_pe_1_6_6_n1), .B1(npu_inst_pe_1_6_6_N77), .B2(
        npu_inst_pe_1_6_6_n76), .C1(npu_inst_pe_1_6_6_N69), .C2(
        npu_inst_pe_1_6_6_n77), .ZN(npu_inst_pe_1_6_6_n80) );
  INV_X1 npu_inst_pe_1_6_6_U40 ( .A(npu_inst_pe_1_6_6_n80), .ZN(
        npu_inst_pe_1_6_6_n36) );
  AOI222_X1 npu_inst_pe_1_6_6_U39 ( .A1(npu_inst_int_data_res_7__6__5_), .A2(
        npu_inst_pe_1_6_6_n1), .B1(npu_inst_pe_1_6_6_N78), .B2(
        npu_inst_pe_1_6_6_n76), .C1(npu_inst_pe_1_6_6_N70), .C2(
        npu_inst_pe_1_6_6_n77), .ZN(npu_inst_pe_1_6_6_n79) );
  INV_X1 npu_inst_pe_1_6_6_U38 ( .A(npu_inst_pe_1_6_6_n79), .ZN(
        npu_inst_pe_1_6_6_n35) );
  AOI222_X1 npu_inst_pe_1_6_6_U37 ( .A1(npu_inst_int_data_res_7__6__6_), .A2(
        npu_inst_pe_1_6_6_n1), .B1(npu_inst_pe_1_6_6_N79), .B2(
        npu_inst_pe_1_6_6_n76), .C1(npu_inst_pe_1_6_6_N71), .C2(
        npu_inst_pe_1_6_6_n77), .ZN(npu_inst_pe_1_6_6_n78) );
  INV_X1 npu_inst_pe_1_6_6_U36 ( .A(npu_inst_pe_1_6_6_n78), .ZN(
        npu_inst_pe_1_6_6_n34) );
  INV_X1 npu_inst_pe_1_6_6_U35 ( .A(npu_inst_pe_1_6_6_int_data_1_), .ZN(
        npu_inst_pe_1_6_6_n14) );
  AND2_X1 npu_inst_pe_1_6_6_U34 ( .A1(npu_inst_int_data_x_6__6__1_), .A2(
        npu_inst_pe_1_6_6_int_q_weight_1_), .ZN(npu_inst_pe_1_6_6_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_6_6_U33 ( .A1(npu_inst_int_data_x_6__6__0_), .A2(
        npu_inst_pe_1_6_6_int_q_weight_1_), .ZN(npu_inst_pe_1_6_6_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_6_6_U32 ( .A1(npu_inst_n53), .A2(
        npu_inst_int_data_y_7__6__1_), .B1(npu_inst_pe_1_6_6_n3), .B2(
        npu_inst_int_data_x_6__7__1_), .ZN(npu_inst_pe_1_6_6_n63) );
  AOI22_X1 npu_inst_pe_1_6_6_U31 ( .A1(npu_inst_n53), .A2(
        npu_inst_int_data_y_7__6__0_), .B1(npu_inst_pe_1_6_6_n3), .B2(
        npu_inst_int_data_x_6__7__0_), .ZN(npu_inst_pe_1_6_6_n61) );
  INV_X1 npu_inst_pe_1_6_6_U30 ( .A(npu_inst_pe_1_6_6_int_data_0_), .ZN(
        npu_inst_pe_1_6_6_n13) );
  INV_X1 npu_inst_pe_1_6_6_U29 ( .A(npu_inst_n67), .ZN(npu_inst_pe_1_6_6_n5)
         );
  OR3_X1 npu_inst_pe_1_6_6_U28 ( .A1(npu_inst_pe_1_6_6_n6), .A2(
        npu_inst_pe_1_6_6_n8), .A3(npu_inst_pe_1_6_6_n5), .ZN(
        npu_inst_pe_1_6_6_n56) );
  OR3_X1 npu_inst_pe_1_6_6_U27 ( .A1(npu_inst_pe_1_6_6_n5), .A2(
        npu_inst_pe_1_6_6_n8), .A3(npu_inst_pe_1_6_6_n7), .ZN(
        npu_inst_pe_1_6_6_n48) );
  INV_X1 npu_inst_pe_1_6_6_U26 ( .A(npu_inst_pe_1_6_6_n5), .ZN(
        npu_inst_pe_1_6_6_n4) );
  OR3_X1 npu_inst_pe_1_6_6_U25 ( .A1(npu_inst_pe_1_6_6_n4), .A2(
        npu_inst_pe_1_6_6_n8), .A3(npu_inst_pe_1_6_6_n7), .ZN(
        npu_inst_pe_1_6_6_n52) );
  OR3_X1 npu_inst_pe_1_6_6_U24 ( .A1(npu_inst_pe_1_6_6_n6), .A2(
        npu_inst_pe_1_6_6_n8), .A3(npu_inst_pe_1_6_6_n4), .ZN(
        npu_inst_pe_1_6_6_n60) );
  NOR2_X1 npu_inst_pe_1_6_6_U23 ( .A1(npu_inst_pe_1_6_6_n60), .A2(
        npu_inst_pe_1_6_6_n3), .ZN(npu_inst_pe_1_6_6_n58) );
  NOR2_X1 npu_inst_pe_1_6_6_U22 ( .A1(npu_inst_pe_1_6_6_n56), .A2(
        npu_inst_pe_1_6_6_n3), .ZN(npu_inst_pe_1_6_6_n54) );
  NOR2_X1 npu_inst_pe_1_6_6_U21 ( .A1(npu_inst_pe_1_6_6_n52), .A2(
        npu_inst_pe_1_6_6_n3), .ZN(npu_inst_pe_1_6_6_n50) );
  NOR2_X1 npu_inst_pe_1_6_6_U20 ( .A1(npu_inst_pe_1_6_6_n48), .A2(
        npu_inst_pe_1_6_6_n3), .ZN(npu_inst_pe_1_6_6_n46) );
  NOR2_X1 npu_inst_pe_1_6_6_U19 ( .A1(npu_inst_pe_1_6_6_n40), .A2(
        npu_inst_pe_1_6_6_n3), .ZN(npu_inst_pe_1_6_6_n38) );
  NOR2_X1 npu_inst_pe_1_6_6_U18 ( .A1(npu_inst_pe_1_6_6_n44), .A2(
        npu_inst_pe_1_6_6_n3), .ZN(npu_inst_pe_1_6_6_n42) );
  BUF_X1 npu_inst_pe_1_6_6_U17 ( .A(npu_inst_n94), .Z(npu_inst_pe_1_6_6_n8) );
  INV_X1 npu_inst_pe_1_6_6_U16 ( .A(npu_inst_n122), .ZN(npu_inst_pe_1_6_6_n12)
         );
  INV_X1 npu_inst_pe_1_6_6_U15 ( .A(npu_inst_pe_1_6_6_n38), .ZN(
        npu_inst_pe_1_6_6_n114) );
  INV_X1 npu_inst_pe_1_6_6_U14 ( .A(npu_inst_pe_1_6_6_n58), .ZN(
        npu_inst_pe_1_6_6_n119) );
  INV_X1 npu_inst_pe_1_6_6_U13 ( .A(npu_inst_pe_1_6_6_n54), .ZN(
        npu_inst_pe_1_6_6_n118) );
  INV_X1 npu_inst_pe_1_6_6_U12 ( .A(npu_inst_pe_1_6_6_n50), .ZN(
        npu_inst_pe_1_6_6_n117) );
  INV_X1 npu_inst_pe_1_6_6_U11 ( .A(npu_inst_pe_1_6_6_n46), .ZN(
        npu_inst_pe_1_6_6_n116) );
  INV_X1 npu_inst_pe_1_6_6_U10 ( .A(npu_inst_pe_1_6_6_n42), .ZN(
        npu_inst_pe_1_6_6_n115) );
  BUF_X1 npu_inst_pe_1_6_6_U9 ( .A(npu_inst_n11), .Z(npu_inst_pe_1_6_6_n2) );
  BUF_X1 npu_inst_pe_1_6_6_U8 ( .A(npu_inst_n11), .Z(npu_inst_pe_1_6_6_n1) );
  BUF_X1 npu_inst_pe_1_6_6_U7 ( .A(npu_inst_pe_1_6_6_n12), .Z(
        npu_inst_pe_1_6_6_n11) );
  BUF_X1 npu_inst_pe_1_6_6_U6 ( .A(npu_inst_pe_1_6_6_n12), .Z(
        npu_inst_pe_1_6_6_n10) );
  BUF_X1 npu_inst_pe_1_6_6_U5 ( .A(npu_inst_pe_1_6_6_n12), .Z(
        npu_inst_pe_1_6_6_n9) );
  NOR2_X1 npu_inst_pe_1_6_6_U4 ( .A1(npu_inst_pe_1_6_6_int_q_weight_0_), .A2(
        npu_inst_pe_1_6_6_n1), .ZN(npu_inst_pe_1_6_6_n76) );
  NOR2_X1 npu_inst_pe_1_6_6_U3 ( .A1(npu_inst_pe_1_6_6_n27), .A2(
        npu_inst_pe_1_6_6_n1), .ZN(npu_inst_pe_1_6_6_n77) );
  FA_X1 npu_inst_pe_1_6_6_sub_67_U2_1 ( .A(npu_inst_pe_1_6_6_int_q_acc_1_), 
        .B(npu_inst_pe_1_6_6_n14), .CI(npu_inst_pe_1_6_6_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_6_6_sub_67_carry_2_), .S(npu_inst_pe_1_6_6_N66) );
  FA_X1 npu_inst_pe_1_6_6_add_69_U1_1 ( .A(npu_inst_pe_1_6_6_int_q_acc_1_), 
        .B(npu_inst_pe_1_6_6_int_data_1_), .CI(
        npu_inst_pe_1_6_6_add_69_carry_1_), .CO(
        npu_inst_pe_1_6_6_add_69_carry_2_), .S(npu_inst_pe_1_6_6_N74) );
  NAND3_X1 npu_inst_pe_1_6_6_U109 ( .A1(npu_inst_pe_1_6_6_n5), .A2(
        npu_inst_pe_1_6_6_n7), .A3(npu_inst_pe_1_6_6_n8), .ZN(
        npu_inst_pe_1_6_6_n44) );
  NAND3_X1 npu_inst_pe_1_6_6_U108 ( .A1(npu_inst_pe_1_6_6_n4), .A2(
        npu_inst_pe_1_6_6_n7), .A3(npu_inst_pe_1_6_6_n8), .ZN(
        npu_inst_pe_1_6_6_n40) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_6_6_n34), .CK(
        npu_inst_pe_1_6_6_net3320), .RN(npu_inst_pe_1_6_6_n9), .Q(
        npu_inst_pe_1_6_6_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_6_6_n35), .CK(
        npu_inst_pe_1_6_6_net3320), .RN(npu_inst_pe_1_6_6_n9), .Q(
        npu_inst_pe_1_6_6_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_6_6_n36), .CK(
        npu_inst_pe_1_6_6_net3320), .RN(npu_inst_pe_1_6_6_n9), .Q(
        npu_inst_pe_1_6_6_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_6_6_n98), .CK(
        npu_inst_pe_1_6_6_net3320), .RN(npu_inst_pe_1_6_6_n9), .Q(
        npu_inst_pe_1_6_6_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_6_6_n99), .CK(
        npu_inst_pe_1_6_6_net3320), .RN(npu_inst_pe_1_6_6_n9), .Q(
        npu_inst_pe_1_6_6_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_6_6_n100), 
        .CK(npu_inst_pe_1_6_6_net3320), .RN(npu_inst_pe_1_6_6_n9), .Q(
        npu_inst_pe_1_6_6_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_6_6_n33), .CK(
        npu_inst_pe_1_6_6_net3320), .RN(npu_inst_pe_1_6_6_n9), .Q(
        npu_inst_pe_1_6_6_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_6_6_n101), 
        .CK(npu_inst_pe_1_6_6_net3320), .RN(npu_inst_pe_1_6_6_n9), .Q(
        npu_inst_pe_1_6_6_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_weight_reg_0_ ( .D(npu_inst_n108), .CK(
        npu_inst_pe_1_6_6_net3326), .RN(npu_inst_pe_1_6_6_n9), .Q(
        npu_inst_pe_1_6_6_int_q_weight_0_), .QN(npu_inst_pe_1_6_6_n27) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_weight_reg_1_ ( .D(npu_inst_n114), .CK(
        npu_inst_pe_1_6_6_net3326), .RN(npu_inst_pe_1_6_6_n9), .Q(
        npu_inst_pe_1_6_6_int_q_weight_1_), .QN(npu_inst_pe_1_6_6_n26) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_6_6_n113), 
        .CK(npu_inst_pe_1_6_6_net3326), .RN(npu_inst_pe_1_6_6_n9), .Q(
        npu_inst_pe_1_6_6_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_6_6_n107), 
        .CK(npu_inst_pe_1_6_6_net3326), .RN(npu_inst_pe_1_6_6_n9), .Q(
        npu_inst_pe_1_6_6_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_6_6_n112), 
        .CK(npu_inst_pe_1_6_6_net3326), .RN(npu_inst_pe_1_6_6_n10), .Q(
        npu_inst_pe_1_6_6_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_6_6_n106), 
        .CK(npu_inst_pe_1_6_6_net3326), .RN(npu_inst_pe_1_6_6_n10), .Q(
        npu_inst_pe_1_6_6_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_6_6_n111), 
        .CK(npu_inst_pe_1_6_6_net3326), .RN(npu_inst_pe_1_6_6_n10), .Q(
        npu_inst_pe_1_6_6_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_6_6_n105), 
        .CK(npu_inst_pe_1_6_6_net3326), .RN(npu_inst_pe_1_6_6_n10), .Q(
        npu_inst_pe_1_6_6_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_6_6_n110), 
        .CK(npu_inst_pe_1_6_6_net3326), .RN(npu_inst_pe_1_6_6_n10), .Q(
        npu_inst_pe_1_6_6_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_6_6_n104), 
        .CK(npu_inst_pe_1_6_6_net3326), .RN(npu_inst_pe_1_6_6_n10), .Q(
        npu_inst_pe_1_6_6_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_6_6_n109), 
        .CK(npu_inst_pe_1_6_6_net3326), .RN(npu_inst_pe_1_6_6_n10), .Q(
        npu_inst_pe_1_6_6_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_6_6_n103), 
        .CK(npu_inst_pe_1_6_6_net3326), .RN(npu_inst_pe_1_6_6_n10), .Q(
        npu_inst_pe_1_6_6_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_6_6_n108), 
        .CK(npu_inst_pe_1_6_6_net3326), .RN(npu_inst_pe_1_6_6_n10), .Q(
        npu_inst_pe_1_6_6_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_6_6_n102), 
        .CK(npu_inst_pe_1_6_6_net3326), .RN(npu_inst_pe_1_6_6_n10), .Q(
        npu_inst_pe_1_6_6_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_6_6_n86), 
        .CK(npu_inst_pe_1_6_6_net3326), .RN(npu_inst_pe_1_6_6_n10), .Q(
        npu_inst_pe_1_6_6_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_6_6_n87), 
        .CK(npu_inst_pe_1_6_6_net3326), .RN(npu_inst_pe_1_6_6_n10), .Q(
        npu_inst_pe_1_6_6_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_6_6_n88), 
        .CK(npu_inst_pe_1_6_6_net3326), .RN(npu_inst_pe_1_6_6_n11), .Q(
        npu_inst_pe_1_6_6_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_6_6_n89), 
        .CK(npu_inst_pe_1_6_6_net3326), .RN(npu_inst_pe_1_6_6_n11), .Q(
        npu_inst_pe_1_6_6_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_6_6_n90), 
        .CK(npu_inst_pe_1_6_6_net3326), .RN(npu_inst_pe_1_6_6_n11), .Q(
        npu_inst_pe_1_6_6_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_6_6_n91), 
        .CK(npu_inst_pe_1_6_6_net3326), .RN(npu_inst_pe_1_6_6_n11), .Q(
        npu_inst_pe_1_6_6_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_6_6_n92), 
        .CK(npu_inst_pe_1_6_6_net3326), .RN(npu_inst_pe_1_6_6_n11), .Q(
        npu_inst_pe_1_6_6_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_6_6_n93), 
        .CK(npu_inst_pe_1_6_6_net3326), .RN(npu_inst_pe_1_6_6_n11), .Q(
        npu_inst_pe_1_6_6_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_6_6_n94), 
        .CK(npu_inst_pe_1_6_6_net3326), .RN(npu_inst_pe_1_6_6_n11), .Q(
        npu_inst_pe_1_6_6_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_6_6_n95), 
        .CK(npu_inst_pe_1_6_6_net3326), .RN(npu_inst_pe_1_6_6_n11), .Q(
        npu_inst_pe_1_6_6_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_6_6_n96), 
        .CK(npu_inst_pe_1_6_6_net3326), .RN(npu_inst_pe_1_6_6_n11), .Q(
        npu_inst_pe_1_6_6_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_6_6_n97), 
        .CK(npu_inst_pe_1_6_6_net3326), .RN(npu_inst_pe_1_6_6_n11), .Q(
        npu_inst_pe_1_6_6_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_6_6_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_6_6_N84), .SE(1'b0), .GCK(npu_inst_pe_1_6_6_net3320) );
  CLKGATETST_X1 npu_inst_pe_1_6_6_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n61), .SE(1'b0), .GCK(npu_inst_pe_1_6_6_net3326) );
  MUX2_X1 npu_inst_pe_1_6_7_U162 ( .A(npu_inst_pe_1_6_7_n32), .B(
        npu_inst_pe_1_6_7_n29), .S(npu_inst_pe_1_6_7_n8), .Z(
        npu_inst_pe_1_6_7_N93) );
  MUX2_X1 npu_inst_pe_1_6_7_U161 ( .A(npu_inst_pe_1_6_7_n31), .B(
        npu_inst_pe_1_6_7_n30), .S(npu_inst_pe_1_6_7_n6), .Z(
        npu_inst_pe_1_6_7_n32) );
  MUX2_X1 npu_inst_pe_1_6_7_U160 ( .A(npu_inst_pe_1_6_7_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_6_7_int_q_reg_v_1__0_), .S(npu_inst_pe_1_6_7_n4), .Z(
        npu_inst_pe_1_6_7_n31) );
  MUX2_X1 npu_inst_pe_1_6_7_U159 ( .A(npu_inst_pe_1_6_7_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_6_7_int_q_reg_v_3__0_), .S(npu_inst_pe_1_6_7_n4), .Z(
        npu_inst_pe_1_6_7_n30) );
  MUX2_X1 npu_inst_pe_1_6_7_U158 ( .A(npu_inst_pe_1_6_7_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_6_7_int_q_reg_v_5__0_), .S(npu_inst_pe_1_6_7_n4), .Z(
        npu_inst_pe_1_6_7_n29) );
  MUX2_X1 npu_inst_pe_1_6_7_U157 ( .A(npu_inst_pe_1_6_7_n28), .B(
        npu_inst_pe_1_6_7_n23), .S(npu_inst_pe_1_6_7_n8), .Z(
        npu_inst_pe_1_6_7_N94) );
  MUX2_X1 npu_inst_pe_1_6_7_U156 ( .A(npu_inst_pe_1_6_7_n25), .B(
        npu_inst_pe_1_6_7_n24), .S(npu_inst_pe_1_6_7_n6), .Z(
        npu_inst_pe_1_6_7_n28) );
  MUX2_X1 npu_inst_pe_1_6_7_U155 ( .A(npu_inst_pe_1_6_7_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_6_7_int_q_reg_v_1__1_), .S(npu_inst_pe_1_6_7_n4), .Z(
        npu_inst_pe_1_6_7_n25) );
  MUX2_X1 npu_inst_pe_1_6_7_U154 ( .A(npu_inst_pe_1_6_7_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_6_7_int_q_reg_v_3__1_), .S(npu_inst_pe_1_6_7_n4), .Z(
        npu_inst_pe_1_6_7_n24) );
  MUX2_X1 npu_inst_pe_1_6_7_U153 ( .A(npu_inst_pe_1_6_7_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_6_7_int_q_reg_v_5__1_), .S(npu_inst_pe_1_6_7_n4), .Z(
        npu_inst_pe_1_6_7_n23) );
  MUX2_X1 npu_inst_pe_1_6_7_U152 ( .A(npu_inst_pe_1_6_7_n22), .B(
        npu_inst_pe_1_6_7_n19), .S(npu_inst_pe_1_6_7_n8), .Z(
        npu_inst_int_data_x_6__7__1_) );
  MUX2_X1 npu_inst_pe_1_6_7_U151 ( .A(npu_inst_pe_1_6_7_n21), .B(
        npu_inst_pe_1_6_7_n20), .S(npu_inst_pe_1_6_7_n6), .Z(
        npu_inst_pe_1_6_7_n22) );
  MUX2_X1 npu_inst_pe_1_6_7_U150 ( .A(npu_inst_pe_1_6_7_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_6_7_int_q_reg_h_1__1_), .S(npu_inst_pe_1_6_7_n4), .Z(
        npu_inst_pe_1_6_7_n21) );
  MUX2_X1 npu_inst_pe_1_6_7_U149 ( .A(npu_inst_pe_1_6_7_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_6_7_int_q_reg_h_3__1_), .S(npu_inst_pe_1_6_7_n4), .Z(
        npu_inst_pe_1_6_7_n20) );
  MUX2_X1 npu_inst_pe_1_6_7_U148 ( .A(npu_inst_pe_1_6_7_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_6_7_int_q_reg_h_5__1_), .S(npu_inst_pe_1_6_7_n4), .Z(
        npu_inst_pe_1_6_7_n19) );
  MUX2_X1 npu_inst_pe_1_6_7_U147 ( .A(npu_inst_pe_1_6_7_n18), .B(
        npu_inst_pe_1_6_7_n15), .S(npu_inst_pe_1_6_7_n8), .Z(
        npu_inst_int_data_x_6__7__0_) );
  MUX2_X1 npu_inst_pe_1_6_7_U146 ( .A(npu_inst_pe_1_6_7_n17), .B(
        npu_inst_pe_1_6_7_n16), .S(npu_inst_pe_1_6_7_n6), .Z(
        npu_inst_pe_1_6_7_n18) );
  MUX2_X1 npu_inst_pe_1_6_7_U145 ( .A(npu_inst_pe_1_6_7_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_6_7_int_q_reg_h_1__0_), .S(npu_inst_pe_1_6_7_n4), .Z(
        npu_inst_pe_1_6_7_n17) );
  MUX2_X1 npu_inst_pe_1_6_7_U144 ( .A(npu_inst_pe_1_6_7_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_6_7_int_q_reg_h_3__0_), .S(npu_inst_pe_1_6_7_n4), .Z(
        npu_inst_pe_1_6_7_n16) );
  MUX2_X1 npu_inst_pe_1_6_7_U143 ( .A(npu_inst_pe_1_6_7_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_6_7_int_q_reg_h_5__0_), .S(npu_inst_pe_1_6_7_n4), .Z(
        npu_inst_pe_1_6_7_n15) );
  XOR2_X1 npu_inst_pe_1_6_7_U142 ( .A(npu_inst_pe_1_6_7_int_data_0_), .B(
        npu_inst_pe_1_6_7_int_q_acc_0_), .Z(npu_inst_pe_1_6_7_N73) );
  AND2_X1 npu_inst_pe_1_6_7_U141 ( .A1(npu_inst_pe_1_6_7_int_q_acc_0_), .A2(
        npu_inst_pe_1_6_7_int_data_0_), .ZN(npu_inst_pe_1_6_7_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_6_7_U140 ( .A(npu_inst_pe_1_6_7_int_q_acc_0_), .B(
        npu_inst_pe_1_6_7_n13), .ZN(npu_inst_pe_1_6_7_N65) );
  OR2_X1 npu_inst_pe_1_6_7_U139 ( .A1(npu_inst_pe_1_6_7_n13), .A2(
        npu_inst_pe_1_6_7_int_q_acc_0_), .ZN(npu_inst_pe_1_6_7_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_6_7_U138 ( .A(npu_inst_pe_1_6_7_int_q_acc_2_), .B(
        npu_inst_pe_1_6_7_add_69_carry_2_), .Z(npu_inst_pe_1_6_7_N75) );
  AND2_X1 npu_inst_pe_1_6_7_U137 ( .A1(npu_inst_pe_1_6_7_add_69_carry_2_), 
        .A2(npu_inst_pe_1_6_7_int_q_acc_2_), .ZN(
        npu_inst_pe_1_6_7_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_6_7_U136 ( .A(npu_inst_pe_1_6_7_int_q_acc_3_), .B(
        npu_inst_pe_1_6_7_add_69_carry_3_), .Z(npu_inst_pe_1_6_7_N76) );
  AND2_X1 npu_inst_pe_1_6_7_U135 ( .A1(npu_inst_pe_1_6_7_add_69_carry_3_), 
        .A2(npu_inst_pe_1_6_7_int_q_acc_3_), .ZN(
        npu_inst_pe_1_6_7_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_6_7_U134 ( .A(npu_inst_pe_1_6_7_int_q_acc_4_), .B(
        npu_inst_pe_1_6_7_add_69_carry_4_), .Z(npu_inst_pe_1_6_7_N77) );
  AND2_X1 npu_inst_pe_1_6_7_U133 ( .A1(npu_inst_pe_1_6_7_add_69_carry_4_), 
        .A2(npu_inst_pe_1_6_7_int_q_acc_4_), .ZN(
        npu_inst_pe_1_6_7_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_6_7_U132 ( .A(npu_inst_pe_1_6_7_int_q_acc_5_), .B(
        npu_inst_pe_1_6_7_add_69_carry_5_), .Z(npu_inst_pe_1_6_7_N78) );
  AND2_X1 npu_inst_pe_1_6_7_U131 ( .A1(npu_inst_pe_1_6_7_add_69_carry_5_), 
        .A2(npu_inst_pe_1_6_7_int_q_acc_5_), .ZN(
        npu_inst_pe_1_6_7_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_6_7_U130 ( .A(npu_inst_pe_1_6_7_int_q_acc_6_), .B(
        npu_inst_pe_1_6_7_add_69_carry_6_), .Z(npu_inst_pe_1_6_7_N79) );
  AND2_X1 npu_inst_pe_1_6_7_U129 ( .A1(npu_inst_pe_1_6_7_add_69_carry_6_), 
        .A2(npu_inst_pe_1_6_7_int_q_acc_6_), .ZN(
        npu_inst_pe_1_6_7_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_6_7_U128 ( .A(npu_inst_pe_1_6_7_int_q_acc_7_), .B(
        npu_inst_pe_1_6_7_add_69_carry_7_), .Z(npu_inst_pe_1_6_7_N80) );
  XNOR2_X1 npu_inst_pe_1_6_7_U127 ( .A(npu_inst_pe_1_6_7_sub_67_carry_2_), .B(
        npu_inst_pe_1_6_7_int_q_acc_2_), .ZN(npu_inst_pe_1_6_7_N67) );
  OR2_X1 npu_inst_pe_1_6_7_U126 ( .A1(npu_inst_pe_1_6_7_int_q_acc_2_), .A2(
        npu_inst_pe_1_6_7_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_6_7_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_6_7_U125 ( .A(npu_inst_pe_1_6_7_sub_67_carry_3_), .B(
        npu_inst_pe_1_6_7_int_q_acc_3_), .ZN(npu_inst_pe_1_6_7_N68) );
  OR2_X1 npu_inst_pe_1_6_7_U124 ( .A1(npu_inst_pe_1_6_7_int_q_acc_3_), .A2(
        npu_inst_pe_1_6_7_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_6_7_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_6_7_U123 ( .A(npu_inst_pe_1_6_7_sub_67_carry_4_), .B(
        npu_inst_pe_1_6_7_int_q_acc_4_), .ZN(npu_inst_pe_1_6_7_N69) );
  OR2_X1 npu_inst_pe_1_6_7_U122 ( .A1(npu_inst_pe_1_6_7_int_q_acc_4_), .A2(
        npu_inst_pe_1_6_7_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_6_7_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_6_7_U121 ( .A(npu_inst_pe_1_6_7_sub_67_carry_5_), .B(
        npu_inst_pe_1_6_7_int_q_acc_5_), .ZN(npu_inst_pe_1_6_7_N70) );
  OR2_X1 npu_inst_pe_1_6_7_U120 ( .A1(npu_inst_pe_1_6_7_int_q_acc_5_), .A2(
        npu_inst_pe_1_6_7_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_6_7_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_6_7_U119 ( .A(npu_inst_pe_1_6_7_sub_67_carry_6_), .B(
        npu_inst_pe_1_6_7_int_q_acc_6_), .ZN(npu_inst_pe_1_6_7_N71) );
  OR2_X1 npu_inst_pe_1_6_7_U118 ( .A1(npu_inst_pe_1_6_7_int_q_acc_6_), .A2(
        npu_inst_pe_1_6_7_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_6_7_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_6_7_U117 ( .A(npu_inst_pe_1_6_7_int_q_acc_7_), .B(
        npu_inst_pe_1_6_7_sub_67_carry_7_), .ZN(npu_inst_pe_1_6_7_N72) );
  INV_X1 npu_inst_pe_1_6_7_U116 ( .A(npu_inst_n75), .ZN(npu_inst_pe_1_6_7_n7)
         );
  INV_X1 npu_inst_pe_1_6_7_U115 ( .A(npu_inst_pe_1_6_7_n7), .ZN(
        npu_inst_pe_1_6_7_n6) );
  INV_X1 npu_inst_pe_1_6_7_U114 ( .A(npu_inst_n53), .ZN(npu_inst_pe_1_6_7_n3)
         );
  AOI22_X1 npu_inst_pe_1_6_7_U113 ( .A1(npu_inst_int_data_y_7__7__0_), .A2(
        npu_inst_pe_1_6_7_n58), .B1(npu_inst_pe_1_6_7_n119), .B2(
        npu_inst_pe_1_6_7_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_6_7_n57) );
  INV_X1 npu_inst_pe_1_6_7_U112 ( .A(npu_inst_pe_1_6_7_n57), .ZN(
        npu_inst_pe_1_6_7_n108) );
  AOI22_X1 npu_inst_pe_1_6_7_U111 ( .A1(npu_inst_int_data_y_7__7__0_), .A2(
        npu_inst_pe_1_6_7_n54), .B1(npu_inst_pe_1_6_7_n118), .B2(
        npu_inst_pe_1_6_7_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_6_7_n53) );
  INV_X1 npu_inst_pe_1_6_7_U110 ( .A(npu_inst_pe_1_6_7_n53), .ZN(
        npu_inst_pe_1_6_7_n109) );
  AOI22_X1 npu_inst_pe_1_6_7_U107 ( .A1(npu_inst_int_data_y_7__7__0_), .A2(
        npu_inst_pe_1_6_7_n50), .B1(npu_inst_pe_1_6_7_n117), .B2(
        npu_inst_pe_1_6_7_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_6_7_n49) );
  INV_X1 npu_inst_pe_1_6_7_U106 ( .A(npu_inst_pe_1_6_7_n49), .ZN(
        npu_inst_pe_1_6_7_n110) );
  AOI22_X1 npu_inst_pe_1_6_7_U105 ( .A1(npu_inst_int_data_y_7__7__0_), .A2(
        npu_inst_pe_1_6_7_n46), .B1(npu_inst_pe_1_6_7_n116), .B2(
        npu_inst_pe_1_6_7_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_6_7_n45) );
  INV_X1 npu_inst_pe_1_6_7_U104 ( .A(npu_inst_pe_1_6_7_n45), .ZN(
        npu_inst_pe_1_6_7_n111) );
  AOI22_X1 npu_inst_pe_1_6_7_U103 ( .A1(npu_inst_int_data_y_7__7__0_), .A2(
        npu_inst_pe_1_6_7_n42), .B1(npu_inst_pe_1_6_7_n115), .B2(
        npu_inst_pe_1_6_7_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_6_7_n41) );
  INV_X1 npu_inst_pe_1_6_7_U102 ( .A(npu_inst_pe_1_6_7_n41), .ZN(
        npu_inst_pe_1_6_7_n112) );
  AOI22_X1 npu_inst_pe_1_6_7_U101 ( .A1(npu_inst_int_data_y_7__7__1_), .A2(
        npu_inst_pe_1_6_7_n58), .B1(npu_inst_pe_1_6_7_n119), .B2(
        npu_inst_pe_1_6_7_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_6_7_n59) );
  INV_X1 npu_inst_pe_1_6_7_U100 ( .A(npu_inst_pe_1_6_7_n59), .ZN(
        npu_inst_pe_1_6_7_n102) );
  AOI22_X1 npu_inst_pe_1_6_7_U99 ( .A1(npu_inst_int_data_y_7__7__1_), .A2(
        npu_inst_pe_1_6_7_n54), .B1(npu_inst_pe_1_6_7_n118), .B2(
        npu_inst_pe_1_6_7_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_6_7_n55) );
  INV_X1 npu_inst_pe_1_6_7_U98 ( .A(npu_inst_pe_1_6_7_n55), .ZN(
        npu_inst_pe_1_6_7_n103) );
  AOI22_X1 npu_inst_pe_1_6_7_U97 ( .A1(npu_inst_int_data_y_7__7__1_), .A2(
        npu_inst_pe_1_6_7_n50), .B1(npu_inst_pe_1_6_7_n117), .B2(
        npu_inst_pe_1_6_7_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_6_7_n51) );
  INV_X1 npu_inst_pe_1_6_7_U96 ( .A(npu_inst_pe_1_6_7_n51), .ZN(
        npu_inst_pe_1_6_7_n104) );
  AOI22_X1 npu_inst_pe_1_6_7_U95 ( .A1(npu_inst_int_data_y_7__7__1_), .A2(
        npu_inst_pe_1_6_7_n46), .B1(npu_inst_pe_1_6_7_n116), .B2(
        npu_inst_pe_1_6_7_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_6_7_n47) );
  INV_X1 npu_inst_pe_1_6_7_U94 ( .A(npu_inst_pe_1_6_7_n47), .ZN(
        npu_inst_pe_1_6_7_n105) );
  AOI22_X1 npu_inst_pe_1_6_7_U93 ( .A1(npu_inst_int_data_y_7__7__1_), .A2(
        npu_inst_pe_1_6_7_n42), .B1(npu_inst_pe_1_6_7_n115), .B2(
        npu_inst_pe_1_6_7_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_6_7_n43) );
  INV_X1 npu_inst_pe_1_6_7_U92 ( .A(npu_inst_pe_1_6_7_n43), .ZN(
        npu_inst_pe_1_6_7_n106) );
  AOI22_X1 npu_inst_pe_1_6_7_U91 ( .A1(npu_inst_pe_1_6_7_n38), .A2(
        npu_inst_int_data_y_7__7__1_), .B1(npu_inst_pe_1_6_7_n114), .B2(
        npu_inst_pe_1_6_7_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_6_7_n39) );
  INV_X1 npu_inst_pe_1_6_7_U90 ( .A(npu_inst_pe_1_6_7_n39), .ZN(
        npu_inst_pe_1_6_7_n107) );
  AOI22_X1 npu_inst_pe_1_6_7_U89 ( .A1(npu_inst_pe_1_6_7_n38), .A2(
        npu_inst_int_data_y_7__7__0_), .B1(npu_inst_pe_1_6_7_n114), .B2(
        npu_inst_pe_1_6_7_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_6_7_n37) );
  INV_X1 npu_inst_pe_1_6_7_U88 ( .A(npu_inst_pe_1_6_7_n37), .ZN(
        npu_inst_pe_1_6_7_n113) );
  AND2_X1 npu_inst_pe_1_6_7_U87 ( .A1(npu_inst_pe_1_6_7_N93), .A2(npu_inst_n53), .ZN(npu_inst_int_data_y_6__7__0_) );
  AND2_X1 npu_inst_pe_1_6_7_U86 ( .A1(npu_inst_n53), .A2(npu_inst_pe_1_6_7_N94), .ZN(npu_inst_int_data_y_6__7__1_) );
  NOR3_X1 npu_inst_pe_1_6_7_U85 ( .A1(npu_inst_pe_1_6_7_n26), .A2(npu_inst_n53), .A3(npu_inst_int_ckg[8]), .ZN(npu_inst_pe_1_6_7_n85) );
  OR2_X1 npu_inst_pe_1_6_7_U84 ( .A1(npu_inst_pe_1_6_7_n85), .A2(
        npu_inst_pe_1_6_7_n2), .ZN(npu_inst_pe_1_6_7_N84) );
  AND2_X1 npu_inst_pe_1_6_7_U83 ( .A1(npu_inst_pe_1_6_7_int_q_acc_0_), .A2(
        npu_inst_pe_1_6_7_n1), .ZN(npu_inst_int_data_res_6__7__0_) );
  AND2_X1 npu_inst_pe_1_6_7_U82 ( .A1(npu_inst_pe_1_6_7_n2), .A2(
        npu_inst_pe_1_6_7_int_q_acc_7_), .ZN(npu_inst_int_data_res_6__7__7_)
         );
  AND2_X1 npu_inst_pe_1_6_7_U81 ( .A1(npu_inst_pe_1_6_7_int_q_acc_1_), .A2(
        npu_inst_pe_1_6_7_n1), .ZN(npu_inst_int_data_res_6__7__1_) );
  AND2_X1 npu_inst_pe_1_6_7_U80 ( .A1(npu_inst_pe_1_6_7_int_q_acc_2_), .A2(
        npu_inst_pe_1_6_7_n1), .ZN(npu_inst_int_data_res_6__7__2_) );
  AND2_X1 npu_inst_pe_1_6_7_U79 ( .A1(npu_inst_pe_1_6_7_int_q_acc_3_), .A2(
        npu_inst_pe_1_6_7_n2), .ZN(npu_inst_int_data_res_6__7__3_) );
  AND2_X1 npu_inst_pe_1_6_7_U78 ( .A1(npu_inst_pe_1_6_7_int_q_acc_4_), .A2(
        npu_inst_pe_1_6_7_n2), .ZN(npu_inst_int_data_res_6__7__4_) );
  AND2_X1 npu_inst_pe_1_6_7_U77 ( .A1(npu_inst_pe_1_6_7_int_q_acc_5_), .A2(
        npu_inst_pe_1_6_7_n2), .ZN(npu_inst_int_data_res_6__7__5_) );
  AND2_X1 npu_inst_pe_1_6_7_U76 ( .A1(npu_inst_pe_1_6_7_int_q_acc_6_), .A2(
        npu_inst_pe_1_6_7_n2), .ZN(npu_inst_int_data_res_6__7__6_) );
  AOI222_X1 npu_inst_pe_1_6_7_U75 ( .A1(npu_inst_int_data_res_7__7__0_), .A2(
        npu_inst_pe_1_6_7_n1), .B1(npu_inst_pe_1_6_7_N73), .B2(
        npu_inst_pe_1_6_7_n76), .C1(npu_inst_pe_1_6_7_N65), .C2(
        npu_inst_pe_1_6_7_n77), .ZN(npu_inst_pe_1_6_7_n84) );
  INV_X1 npu_inst_pe_1_6_7_U74 ( .A(npu_inst_pe_1_6_7_n84), .ZN(
        npu_inst_pe_1_6_7_n101) );
  AOI222_X1 npu_inst_pe_1_6_7_U73 ( .A1(npu_inst_int_data_res_7__7__7_), .A2(
        npu_inst_pe_1_6_7_n1), .B1(npu_inst_pe_1_6_7_N80), .B2(
        npu_inst_pe_1_6_7_n76), .C1(npu_inst_pe_1_6_7_N72), .C2(
        npu_inst_pe_1_6_7_n77), .ZN(npu_inst_pe_1_6_7_n75) );
  INV_X1 npu_inst_pe_1_6_7_U72 ( .A(npu_inst_pe_1_6_7_n75), .ZN(
        npu_inst_pe_1_6_7_n33) );
  AOI222_X1 npu_inst_pe_1_6_7_U71 ( .A1(npu_inst_int_data_res_7__7__1_), .A2(
        npu_inst_pe_1_6_7_n1), .B1(npu_inst_pe_1_6_7_N74), .B2(
        npu_inst_pe_1_6_7_n76), .C1(npu_inst_pe_1_6_7_N66), .C2(
        npu_inst_pe_1_6_7_n77), .ZN(npu_inst_pe_1_6_7_n83) );
  INV_X1 npu_inst_pe_1_6_7_U70 ( .A(npu_inst_pe_1_6_7_n83), .ZN(
        npu_inst_pe_1_6_7_n100) );
  AOI222_X1 npu_inst_pe_1_6_7_U69 ( .A1(npu_inst_int_data_res_7__7__2_), .A2(
        npu_inst_pe_1_6_7_n1), .B1(npu_inst_pe_1_6_7_N75), .B2(
        npu_inst_pe_1_6_7_n76), .C1(npu_inst_pe_1_6_7_N67), .C2(
        npu_inst_pe_1_6_7_n77), .ZN(npu_inst_pe_1_6_7_n82) );
  INV_X1 npu_inst_pe_1_6_7_U68 ( .A(npu_inst_pe_1_6_7_n82), .ZN(
        npu_inst_pe_1_6_7_n99) );
  AOI222_X1 npu_inst_pe_1_6_7_U67 ( .A1(npu_inst_int_data_res_7__7__3_), .A2(
        npu_inst_pe_1_6_7_n1), .B1(npu_inst_pe_1_6_7_N76), .B2(
        npu_inst_pe_1_6_7_n76), .C1(npu_inst_pe_1_6_7_N68), .C2(
        npu_inst_pe_1_6_7_n77), .ZN(npu_inst_pe_1_6_7_n81) );
  INV_X1 npu_inst_pe_1_6_7_U66 ( .A(npu_inst_pe_1_6_7_n81), .ZN(
        npu_inst_pe_1_6_7_n98) );
  AOI222_X1 npu_inst_pe_1_6_7_U65 ( .A1(npu_inst_int_data_res_7__7__4_), .A2(
        npu_inst_pe_1_6_7_n1), .B1(npu_inst_pe_1_6_7_N77), .B2(
        npu_inst_pe_1_6_7_n76), .C1(npu_inst_pe_1_6_7_N69), .C2(
        npu_inst_pe_1_6_7_n77), .ZN(npu_inst_pe_1_6_7_n80) );
  INV_X1 npu_inst_pe_1_6_7_U64 ( .A(npu_inst_pe_1_6_7_n80), .ZN(
        npu_inst_pe_1_6_7_n36) );
  AOI222_X1 npu_inst_pe_1_6_7_U63 ( .A1(npu_inst_int_data_res_7__7__5_), .A2(
        npu_inst_pe_1_6_7_n1), .B1(npu_inst_pe_1_6_7_N78), .B2(
        npu_inst_pe_1_6_7_n76), .C1(npu_inst_pe_1_6_7_N70), .C2(
        npu_inst_pe_1_6_7_n77), .ZN(npu_inst_pe_1_6_7_n79) );
  INV_X1 npu_inst_pe_1_6_7_U62 ( .A(npu_inst_pe_1_6_7_n79), .ZN(
        npu_inst_pe_1_6_7_n35) );
  AOI222_X1 npu_inst_pe_1_6_7_U61 ( .A1(npu_inst_int_data_res_7__7__6_), .A2(
        npu_inst_pe_1_6_7_n1), .B1(npu_inst_pe_1_6_7_N79), .B2(
        npu_inst_pe_1_6_7_n76), .C1(npu_inst_pe_1_6_7_N71), .C2(
        npu_inst_pe_1_6_7_n77), .ZN(npu_inst_pe_1_6_7_n78) );
  INV_X1 npu_inst_pe_1_6_7_U60 ( .A(npu_inst_pe_1_6_7_n78), .ZN(
        npu_inst_pe_1_6_7_n34) );
  INV_X1 npu_inst_pe_1_6_7_U59 ( .A(npu_inst_pe_1_6_7_int_data_1_), .ZN(
        npu_inst_pe_1_6_7_n14) );
  AND2_X1 npu_inst_pe_1_6_7_U58 ( .A1(npu_inst_int_data_x_6__7__1_), .A2(
        npu_inst_pe_1_6_7_int_q_weight_1_), .ZN(npu_inst_pe_1_6_7_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_6_7_U57 ( .A1(npu_inst_int_data_x_6__7__0_), .A2(
        npu_inst_pe_1_6_7_int_q_weight_1_), .ZN(npu_inst_pe_1_6_7_int_data_0_)
         );
  NAND2_X1 npu_inst_pe_1_6_7_U56 ( .A1(npu_inst_pe_1_6_7_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_6_7_n60), .ZN(npu_inst_pe_1_6_7_n74) );
  OAI21_X1 npu_inst_pe_1_6_7_U55 ( .B1(npu_inst_pe_1_6_7_n63), .B2(
        npu_inst_pe_1_6_7_n60), .A(npu_inst_pe_1_6_7_n74), .ZN(
        npu_inst_pe_1_6_7_n97) );
  NAND2_X1 npu_inst_pe_1_6_7_U54 ( .A1(npu_inst_pe_1_6_7_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_6_7_n60), .ZN(npu_inst_pe_1_6_7_n73) );
  OAI21_X1 npu_inst_pe_1_6_7_U53 ( .B1(npu_inst_pe_1_6_7_n61), .B2(
        npu_inst_pe_1_6_7_n60), .A(npu_inst_pe_1_6_7_n73), .ZN(
        npu_inst_pe_1_6_7_n96) );
  NAND2_X1 npu_inst_pe_1_6_7_U52 ( .A1(npu_inst_pe_1_6_7_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_6_7_n56), .ZN(npu_inst_pe_1_6_7_n72) );
  OAI21_X1 npu_inst_pe_1_6_7_U51 ( .B1(npu_inst_pe_1_6_7_n63), .B2(
        npu_inst_pe_1_6_7_n56), .A(npu_inst_pe_1_6_7_n72), .ZN(
        npu_inst_pe_1_6_7_n95) );
  NAND2_X1 npu_inst_pe_1_6_7_U50 ( .A1(npu_inst_pe_1_6_7_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_6_7_n56), .ZN(npu_inst_pe_1_6_7_n71) );
  OAI21_X1 npu_inst_pe_1_6_7_U49 ( .B1(npu_inst_pe_1_6_7_n61), .B2(
        npu_inst_pe_1_6_7_n56), .A(npu_inst_pe_1_6_7_n71), .ZN(
        npu_inst_pe_1_6_7_n94) );
  NAND2_X1 npu_inst_pe_1_6_7_U48 ( .A1(npu_inst_pe_1_6_7_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_6_7_n52), .ZN(npu_inst_pe_1_6_7_n70) );
  OAI21_X1 npu_inst_pe_1_6_7_U47 ( .B1(npu_inst_pe_1_6_7_n63), .B2(
        npu_inst_pe_1_6_7_n52), .A(npu_inst_pe_1_6_7_n70), .ZN(
        npu_inst_pe_1_6_7_n93) );
  NAND2_X1 npu_inst_pe_1_6_7_U46 ( .A1(npu_inst_pe_1_6_7_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_6_7_n52), .ZN(npu_inst_pe_1_6_7_n69) );
  OAI21_X1 npu_inst_pe_1_6_7_U45 ( .B1(npu_inst_pe_1_6_7_n61), .B2(
        npu_inst_pe_1_6_7_n52), .A(npu_inst_pe_1_6_7_n69), .ZN(
        npu_inst_pe_1_6_7_n92) );
  NAND2_X1 npu_inst_pe_1_6_7_U44 ( .A1(npu_inst_pe_1_6_7_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_6_7_n48), .ZN(npu_inst_pe_1_6_7_n68) );
  OAI21_X1 npu_inst_pe_1_6_7_U43 ( .B1(npu_inst_pe_1_6_7_n63), .B2(
        npu_inst_pe_1_6_7_n48), .A(npu_inst_pe_1_6_7_n68), .ZN(
        npu_inst_pe_1_6_7_n91) );
  NAND2_X1 npu_inst_pe_1_6_7_U42 ( .A1(npu_inst_pe_1_6_7_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_6_7_n48), .ZN(npu_inst_pe_1_6_7_n67) );
  OAI21_X1 npu_inst_pe_1_6_7_U41 ( .B1(npu_inst_pe_1_6_7_n61), .B2(
        npu_inst_pe_1_6_7_n48), .A(npu_inst_pe_1_6_7_n67), .ZN(
        npu_inst_pe_1_6_7_n90) );
  NAND2_X1 npu_inst_pe_1_6_7_U40 ( .A1(npu_inst_pe_1_6_7_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_6_7_n44), .ZN(npu_inst_pe_1_6_7_n66) );
  OAI21_X1 npu_inst_pe_1_6_7_U39 ( .B1(npu_inst_pe_1_6_7_n63), .B2(
        npu_inst_pe_1_6_7_n44), .A(npu_inst_pe_1_6_7_n66), .ZN(
        npu_inst_pe_1_6_7_n89) );
  NAND2_X1 npu_inst_pe_1_6_7_U38 ( .A1(npu_inst_pe_1_6_7_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_6_7_n44), .ZN(npu_inst_pe_1_6_7_n65) );
  OAI21_X1 npu_inst_pe_1_6_7_U37 ( .B1(npu_inst_pe_1_6_7_n61), .B2(
        npu_inst_pe_1_6_7_n44), .A(npu_inst_pe_1_6_7_n65), .ZN(
        npu_inst_pe_1_6_7_n88) );
  NAND2_X1 npu_inst_pe_1_6_7_U36 ( .A1(npu_inst_pe_1_6_7_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_6_7_n40), .ZN(npu_inst_pe_1_6_7_n64) );
  OAI21_X1 npu_inst_pe_1_6_7_U35 ( .B1(npu_inst_pe_1_6_7_n63), .B2(
        npu_inst_pe_1_6_7_n40), .A(npu_inst_pe_1_6_7_n64), .ZN(
        npu_inst_pe_1_6_7_n87) );
  NAND2_X1 npu_inst_pe_1_6_7_U34 ( .A1(npu_inst_pe_1_6_7_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_6_7_n40), .ZN(npu_inst_pe_1_6_7_n62) );
  OAI21_X1 npu_inst_pe_1_6_7_U33 ( .B1(npu_inst_pe_1_6_7_n61), .B2(
        npu_inst_pe_1_6_7_n40), .A(npu_inst_pe_1_6_7_n62), .ZN(
        npu_inst_pe_1_6_7_n86) );
  INV_X1 npu_inst_pe_1_6_7_U32 ( .A(npu_inst_pe_1_6_7_int_data_0_), .ZN(
        npu_inst_pe_1_6_7_n13) );
  INV_X1 npu_inst_pe_1_6_7_U31 ( .A(npu_inst_n67), .ZN(npu_inst_pe_1_6_7_n5)
         );
  AOI22_X1 npu_inst_pe_1_6_7_U30 ( .A1(npu_inst_n53), .A2(
        npu_inst_int_data_y_7__7__1_), .B1(npu_inst_pe_1_6_7_n3), .B2(
        int_i_data_h_npu[3]), .ZN(npu_inst_pe_1_6_7_n63) );
  AOI22_X1 npu_inst_pe_1_6_7_U29 ( .A1(npu_inst_n53), .A2(
        npu_inst_int_data_y_7__7__0_), .B1(npu_inst_pe_1_6_7_n3), .B2(
        int_i_data_h_npu[2]), .ZN(npu_inst_pe_1_6_7_n61) );
  OR3_X1 npu_inst_pe_1_6_7_U28 ( .A1(npu_inst_pe_1_6_7_n6), .A2(
        npu_inst_pe_1_6_7_n8), .A3(npu_inst_pe_1_6_7_n5), .ZN(
        npu_inst_pe_1_6_7_n56) );
  OR3_X1 npu_inst_pe_1_6_7_U27 ( .A1(npu_inst_pe_1_6_7_n5), .A2(
        npu_inst_pe_1_6_7_n8), .A3(npu_inst_pe_1_6_7_n7), .ZN(
        npu_inst_pe_1_6_7_n48) );
  INV_X1 npu_inst_pe_1_6_7_U26 ( .A(npu_inst_pe_1_6_7_n5), .ZN(
        npu_inst_pe_1_6_7_n4) );
  OR3_X1 npu_inst_pe_1_6_7_U25 ( .A1(npu_inst_pe_1_6_7_n4), .A2(
        npu_inst_pe_1_6_7_n8), .A3(npu_inst_pe_1_6_7_n7), .ZN(
        npu_inst_pe_1_6_7_n52) );
  OR3_X1 npu_inst_pe_1_6_7_U24 ( .A1(npu_inst_pe_1_6_7_n6), .A2(
        npu_inst_pe_1_6_7_n8), .A3(npu_inst_pe_1_6_7_n4), .ZN(
        npu_inst_pe_1_6_7_n60) );
  NOR2_X1 npu_inst_pe_1_6_7_U23 ( .A1(npu_inst_pe_1_6_7_n60), .A2(
        npu_inst_pe_1_6_7_n3), .ZN(npu_inst_pe_1_6_7_n58) );
  NOR2_X1 npu_inst_pe_1_6_7_U22 ( .A1(npu_inst_pe_1_6_7_n56), .A2(
        npu_inst_pe_1_6_7_n3), .ZN(npu_inst_pe_1_6_7_n54) );
  NOR2_X1 npu_inst_pe_1_6_7_U21 ( .A1(npu_inst_pe_1_6_7_n52), .A2(
        npu_inst_pe_1_6_7_n3), .ZN(npu_inst_pe_1_6_7_n50) );
  NOR2_X1 npu_inst_pe_1_6_7_U20 ( .A1(npu_inst_pe_1_6_7_n48), .A2(
        npu_inst_pe_1_6_7_n3), .ZN(npu_inst_pe_1_6_7_n46) );
  NOR2_X1 npu_inst_pe_1_6_7_U19 ( .A1(npu_inst_pe_1_6_7_n40), .A2(
        npu_inst_pe_1_6_7_n3), .ZN(npu_inst_pe_1_6_7_n38) );
  NOR2_X1 npu_inst_pe_1_6_7_U18 ( .A1(npu_inst_pe_1_6_7_n44), .A2(
        npu_inst_pe_1_6_7_n3), .ZN(npu_inst_pe_1_6_7_n42) );
  BUF_X1 npu_inst_pe_1_6_7_U17 ( .A(npu_inst_n94), .Z(npu_inst_pe_1_6_7_n8) );
  INV_X1 npu_inst_pe_1_6_7_U16 ( .A(npu_inst_n122), .ZN(npu_inst_pe_1_6_7_n12)
         );
  INV_X1 npu_inst_pe_1_6_7_U15 ( .A(npu_inst_pe_1_6_7_n38), .ZN(
        npu_inst_pe_1_6_7_n114) );
  INV_X1 npu_inst_pe_1_6_7_U14 ( .A(npu_inst_pe_1_6_7_n58), .ZN(
        npu_inst_pe_1_6_7_n119) );
  INV_X1 npu_inst_pe_1_6_7_U13 ( .A(npu_inst_pe_1_6_7_n54), .ZN(
        npu_inst_pe_1_6_7_n118) );
  INV_X1 npu_inst_pe_1_6_7_U12 ( .A(npu_inst_pe_1_6_7_n50), .ZN(
        npu_inst_pe_1_6_7_n117) );
  INV_X1 npu_inst_pe_1_6_7_U11 ( .A(npu_inst_pe_1_6_7_n46), .ZN(
        npu_inst_pe_1_6_7_n116) );
  INV_X1 npu_inst_pe_1_6_7_U10 ( .A(npu_inst_pe_1_6_7_n42), .ZN(
        npu_inst_pe_1_6_7_n115) );
  BUF_X1 npu_inst_pe_1_6_7_U9 ( .A(npu_inst_n11), .Z(npu_inst_pe_1_6_7_n2) );
  BUF_X1 npu_inst_pe_1_6_7_U8 ( .A(npu_inst_n11), .Z(npu_inst_pe_1_6_7_n1) );
  BUF_X1 npu_inst_pe_1_6_7_U7 ( .A(npu_inst_pe_1_6_7_n12), .Z(
        npu_inst_pe_1_6_7_n11) );
  BUF_X1 npu_inst_pe_1_6_7_U6 ( .A(npu_inst_pe_1_6_7_n12), .Z(
        npu_inst_pe_1_6_7_n10) );
  BUF_X1 npu_inst_pe_1_6_7_U5 ( .A(npu_inst_pe_1_6_7_n12), .Z(
        npu_inst_pe_1_6_7_n9) );
  NOR2_X1 npu_inst_pe_1_6_7_U4 ( .A1(npu_inst_pe_1_6_7_int_q_weight_0_), .A2(
        npu_inst_pe_1_6_7_n1), .ZN(npu_inst_pe_1_6_7_n76) );
  NOR2_X1 npu_inst_pe_1_6_7_U3 ( .A1(npu_inst_pe_1_6_7_n27), .A2(
        npu_inst_pe_1_6_7_n1), .ZN(npu_inst_pe_1_6_7_n77) );
  FA_X1 npu_inst_pe_1_6_7_sub_67_U2_1 ( .A(npu_inst_pe_1_6_7_int_q_acc_1_), 
        .B(npu_inst_pe_1_6_7_n14), .CI(npu_inst_pe_1_6_7_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_6_7_sub_67_carry_2_), .S(npu_inst_pe_1_6_7_N66) );
  FA_X1 npu_inst_pe_1_6_7_add_69_U1_1 ( .A(npu_inst_pe_1_6_7_int_q_acc_1_), 
        .B(npu_inst_pe_1_6_7_int_data_1_), .CI(
        npu_inst_pe_1_6_7_add_69_carry_1_), .CO(
        npu_inst_pe_1_6_7_add_69_carry_2_), .S(npu_inst_pe_1_6_7_N74) );
  NAND3_X1 npu_inst_pe_1_6_7_U109 ( .A1(npu_inst_pe_1_6_7_n5), .A2(
        npu_inst_pe_1_6_7_n7), .A3(npu_inst_pe_1_6_7_n8), .ZN(
        npu_inst_pe_1_6_7_n44) );
  NAND3_X1 npu_inst_pe_1_6_7_U108 ( .A1(npu_inst_pe_1_6_7_n4), .A2(
        npu_inst_pe_1_6_7_n7), .A3(npu_inst_pe_1_6_7_n8), .ZN(
        npu_inst_pe_1_6_7_n40) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_6_7_n34), .CK(
        npu_inst_pe_1_6_7_net3297), .RN(npu_inst_pe_1_6_7_n9), .Q(
        npu_inst_pe_1_6_7_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_6_7_n35), .CK(
        npu_inst_pe_1_6_7_net3297), .RN(npu_inst_pe_1_6_7_n9), .Q(
        npu_inst_pe_1_6_7_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_6_7_n36), .CK(
        npu_inst_pe_1_6_7_net3297), .RN(npu_inst_pe_1_6_7_n9), .Q(
        npu_inst_pe_1_6_7_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_6_7_n98), .CK(
        npu_inst_pe_1_6_7_net3297), .RN(npu_inst_pe_1_6_7_n9), .Q(
        npu_inst_pe_1_6_7_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_6_7_n99), .CK(
        npu_inst_pe_1_6_7_net3297), .RN(npu_inst_pe_1_6_7_n9), .Q(
        npu_inst_pe_1_6_7_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_6_7_n100), 
        .CK(npu_inst_pe_1_6_7_net3297), .RN(npu_inst_pe_1_6_7_n9), .Q(
        npu_inst_pe_1_6_7_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_6_7_n33), .CK(
        npu_inst_pe_1_6_7_net3297), .RN(npu_inst_pe_1_6_7_n9), .Q(
        npu_inst_pe_1_6_7_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_6_7_n101), 
        .CK(npu_inst_pe_1_6_7_net3297), .RN(npu_inst_pe_1_6_7_n9), .Q(
        npu_inst_pe_1_6_7_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_weight_reg_0_ ( .D(npu_inst_n108), .CK(
        npu_inst_pe_1_6_7_net3303), .RN(npu_inst_pe_1_6_7_n9), .Q(
        npu_inst_pe_1_6_7_int_q_weight_0_), .QN(npu_inst_pe_1_6_7_n27) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_weight_reg_1_ ( .D(npu_inst_n114), .CK(
        npu_inst_pe_1_6_7_net3303), .RN(npu_inst_pe_1_6_7_n9), .Q(
        npu_inst_pe_1_6_7_int_q_weight_1_), .QN(npu_inst_pe_1_6_7_n26) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_6_7_n113), 
        .CK(npu_inst_pe_1_6_7_net3303), .RN(npu_inst_pe_1_6_7_n9), .Q(
        npu_inst_pe_1_6_7_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_6_7_n107), 
        .CK(npu_inst_pe_1_6_7_net3303), .RN(npu_inst_pe_1_6_7_n9), .Q(
        npu_inst_pe_1_6_7_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_6_7_n112), 
        .CK(npu_inst_pe_1_6_7_net3303), .RN(npu_inst_pe_1_6_7_n10), .Q(
        npu_inst_pe_1_6_7_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_6_7_n106), 
        .CK(npu_inst_pe_1_6_7_net3303), .RN(npu_inst_pe_1_6_7_n10), .Q(
        npu_inst_pe_1_6_7_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_6_7_n111), 
        .CK(npu_inst_pe_1_6_7_net3303), .RN(npu_inst_pe_1_6_7_n10), .Q(
        npu_inst_pe_1_6_7_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_6_7_n105), 
        .CK(npu_inst_pe_1_6_7_net3303), .RN(npu_inst_pe_1_6_7_n10), .Q(
        npu_inst_pe_1_6_7_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_6_7_n110), 
        .CK(npu_inst_pe_1_6_7_net3303), .RN(npu_inst_pe_1_6_7_n10), .Q(
        npu_inst_pe_1_6_7_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_6_7_n104), 
        .CK(npu_inst_pe_1_6_7_net3303), .RN(npu_inst_pe_1_6_7_n10), .Q(
        npu_inst_pe_1_6_7_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_6_7_n109), 
        .CK(npu_inst_pe_1_6_7_net3303), .RN(npu_inst_pe_1_6_7_n10), .Q(
        npu_inst_pe_1_6_7_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_6_7_n103), 
        .CK(npu_inst_pe_1_6_7_net3303), .RN(npu_inst_pe_1_6_7_n10), .Q(
        npu_inst_pe_1_6_7_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_6_7_n108), 
        .CK(npu_inst_pe_1_6_7_net3303), .RN(npu_inst_pe_1_6_7_n10), .Q(
        npu_inst_pe_1_6_7_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_6_7_n102), 
        .CK(npu_inst_pe_1_6_7_net3303), .RN(npu_inst_pe_1_6_7_n10), .Q(
        npu_inst_pe_1_6_7_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_6_7_n86), 
        .CK(npu_inst_pe_1_6_7_net3303), .RN(npu_inst_pe_1_6_7_n10), .Q(
        npu_inst_pe_1_6_7_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_6_7_n87), 
        .CK(npu_inst_pe_1_6_7_net3303), .RN(npu_inst_pe_1_6_7_n10), .Q(
        npu_inst_pe_1_6_7_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_6_7_n88), 
        .CK(npu_inst_pe_1_6_7_net3303), .RN(npu_inst_pe_1_6_7_n11), .Q(
        npu_inst_pe_1_6_7_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_6_7_n89), 
        .CK(npu_inst_pe_1_6_7_net3303), .RN(npu_inst_pe_1_6_7_n11), .Q(
        npu_inst_pe_1_6_7_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_6_7_n90), 
        .CK(npu_inst_pe_1_6_7_net3303), .RN(npu_inst_pe_1_6_7_n11), .Q(
        npu_inst_pe_1_6_7_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_6_7_n91), 
        .CK(npu_inst_pe_1_6_7_net3303), .RN(npu_inst_pe_1_6_7_n11), .Q(
        npu_inst_pe_1_6_7_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_6_7_n92), 
        .CK(npu_inst_pe_1_6_7_net3303), .RN(npu_inst_pe_1_6_7_n11), .Q(
        npu_inst_pe_1_6_7_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_6_7_n93), 
        .CK(npu_inst_pe_1_6_7_net3303), .RN(npu_inst_pe_1_6_7_n11), .Q(
        npu_inst_pe_1_6_7_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_6_7_n94), 
        .CK(npu_inst_pe_1_6_7_net3303), .RN(npu_inst_pe_1_6_7_n11), .Q(
        npu_inst_pe_1_6_7_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_6_7_n95), 
        .CK(npu_inst_pe_1_6_7_net3303), .RN(npu_inst_pe_1_6_7_n11), .Q(
        npu_inst_pe_1_6_7_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_6_7_n96), 
        .CK(npu_inst_pe_1_6_7_net3303), .RN(npu_inst_pe_1_6_7_n11), .Q(
        npu_inst_pe_1_6_7_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_6_7_n97), 
        .CK(npu_inst_pe_1_6_7_net3303), .RN(npu_inst_pe_1_6_7_n11), .Q(
        npu_inst_pe_1_6_7_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_6_7_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_6_7_N84), .SE(1'b0), .GCK(npu_inst_pe_1_6_7_net3297) );
  CLKGATETST_X1 npu_inst_pe_1_6_7_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n61), .SE(1'b0), .GCK(npu_inst_pe_1_6_7_net3303) );
  MUX2_X1 npu_inst_pe_1_7_0_U162 ( .A(npu_inst_pe_1_7_0_n32), .B(
        npu_inst_pe_1_7_0_n29), .S(npu_inst_pe_1_7_0_n8), .Z(
        npu_inst_pe_1_7_0_N93) );
  MUX2_X1 npu_inst_pe_1_7_0_U161 ( .A(npu_inst_pe_1_7_0_n31), .B(
        npu_inst_pe_1_7_0_n30), .S(npu_inst_pe_1_7_0_n6), .Z(
        npu_inst_pe_1_7_0_n32) );
  MUX2_X1 npu_inst_pe_1_7_0_U160 ( .A(npu_inst_pe_1_7_0_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_7_0_int_q_reg_v_1__0_), .S(npu_inst_pe_1_7_0_n4), .Z(
        npu_inst_pe_1_7_0_n31) );
  MUX2_X1 npu_inst_pe_1_7_0_U159 ( .A(npu_inst_pe_1_7_0_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_7_0_int_q_reg_v_3__0_), .S(npu_inst_pe_1_7_0_n4), .Z(
        npu_inst_pe_1_7_0_n30) );
  MUX2_X1 npu_inst_pe_1_7_0_U158 ( .A(npu_inst_pe_1_7_0_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_7_0_int_q_reg_v_5__0_), .S(npu_inst_pe_1_7_0_n4), .Z(
        npu_inst_pe_1_7_0_n29) );
  MUX2_X1 npu_inst_pe_1_7_0_U157 ( .A(npu_inst_pe_1_7_0_n28), .B(
        npu_inst_pe_1_7_0_n23), .S(npu_inst_pe_1_7_0_n8), .Z(
        npu_inst_pe_1_7_0_N94) );
  MUX2_X1 npu_inst_pe_1_7_0_U156 ( .A(npu_inst_pe_1_7_0_n25), .B(
        npu_inst_pe_1_7_0_n24), .S(npu_inst_pe_1_7_0_n6), .Z(
        npu_inst_pe_1_7_0_n28) );
  MUX2_X1 npu_inst_pe_1_7_0_U155 ( .A(npu_inst_pe_1_7_0_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_7_0_int_q_reg_v_1__1_), .S(npu_inst_pe_1_7_0_n4), .Z(
        npu_inst_pe_1_7_0_n25) );
  MUX2_X1 npu_inst_pe_1_7_0_U154 ( .A(npu_inst_pe_1_7_0_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_7_0_int_q_reg_v_3__1_), .S(npu_inst_pe_1_7_0_n4), .Z(
        npu_inst_pe_1_7_0_n24) );
  MUX2_X1 npu_inst_pe_1_7_0_U153 ( .A(npu_inst_pe_1_7_0_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_7_0_int_q_reg_v_5__1_), .S(npu_inst_pe_1_7_0_n4), .Z(
        npu_inst_pe_1_7_0_n23) );
  MUX2_X1 npu_inst_pe_1_7_0_U152 ( .A(npu_inst_pe_1_7_0_n22), .B(
        npu_inst_pe_1_7_0_n19), .S(npu_inst_pe_1_7_0_n8), .Z(
        npu_inst_pe_1_7_0_o_data_h_1_) );
  MUX2_X1 npu_inst_pe_1_7_0_U151 ( .A(npu_inst_pe_1_7_0_n21), .B(
        npu_inst_pe_1_7_0_n20), .S(npu_inst_pe_1_7_0_n6), .Z(
        npu_inst_pe_1_7_0_n22) );
  MUX2_X1 npu_inst_pe_1_7_0_U150 ( .A(npu_inst_pe_1_7_0_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_7_0_int_q_reg_h_1__1_), .S(npu_inst_pe_1_7_0_n4), .Z(
        npu_inst_pe_1_7_0_n21) );
  MUX2_X1 npu_inst_pe_1_7_0_U149 ( .A(npu_inst_pe_1_7_0_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_7_0_int_q_reg_h_3__1_), .S(npu_inst_pe_1_7_0_n4), .Z(
        npu_inst_pe_1_7_0_n20) );
  MUX2_X1 npu_inst_pe_1_7_0_U148 ( .A(npu_inst_pe_1_7_0_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_7_0_int_q_reg_h_5__1_), .S(npu_inst_pe_1_7_0_n4), .Z(
        npu_inst_pe_1_7_0_n19) );
  MUX2_X1 npu_inst_pe_1_7_0_U147 ( .A(npu_inst_pe_1_7_0_n18), .B(
        npu_inst_pe_1_7_0_n15), .S(npu_inst_pe_1_7_0_n8), .Z(
        npu_inst_pe_1_7_0_o_data_h_0_) );
  MUX2_X1 npu_inst_pe_1_7_0_U146 ( .A(npu_inst_pe_1_7_0_n17), .B(
        npu_inst_pe_1_7_0_n16), .S(npu_inst_pe_1_7_0_n6), .Z(
        npu_inst_pe_1_7_0_n18) );
  MUX2_X1 npu_inst_pe_1_7_0_U145 ( .A(npu_inst_pe_1_7_0_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_7_0_int_q_reg_h_1__0_), .S(npu_inst_pe_1_7_0_n4), .Z(
        npu_inst_pe_1_7_0_n17) );
  MUX2_X1 npu_inst_pe_1_7_0_U144 ( .A(npu_inst_pe_1_7_0_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_7_0_int_q_reg_h_3__0_), .S(npu_inst_pe_1_7_0_n4), .Z(
        npu_inst_pe_1_7_0_n16) );
  MUX2_X1 npu_inst_pe_1_7_0_U143 ( .A(npu_inst_pe_1_7_0_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_7_0_int_q_reg_h_5__0_), .S(npu_inst_pe_1_7_0_n4), .Z(
        npu_inst_pe_1_7_0_n15) );
  XOR2_X1 npu_inst_pe_1_7_0_U142 ( .A(npu_inst_pe_1_7_0_int_data_0_), .B(
        npu_inst_pe_1_7_0_int_q_acc_0_), .Z(npu_inst_pe_1_7_0_N73) );
  AND2_X1 npu_inst_pe_1_7_0_U141 ( .A1(npu_inst_pe_1_7_0_int_q_acc_0_), .A2(
        npu_inst_pe_1_7_0_int_data_0_), .ZN(npu_inst_pe_1_7_0_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_7_0_U140 ( .A(npu_inst_pe_1_7_0_int_q_acc_0_), .B(
        npu_inst_pe_1_7_0_n13), .ZN(npu_inst_pe_1_7_0_N65) );
  OR2_X1 npu_inst_pe_1_7_0_U139 ( .A1(npu_inst_pe_1_7_0_n13), .A2(
        npu_inst_pe_1_7_0_int_q_acc_0_), .ZN(npu_inst_pe_1_7_0_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_7_0_U138 ( .A(npu_inst_pe_1_7_0_int_q_acc_2_), .B(
        npu_inst_pe_1_7_0_add_69_carry_2_), .Z(npu_inst_pe_1_7_0_N75) );
  AND2_X1 npu_inst_pe_1_7_0_U137 ( .A1(npu_inst_pe_1_7_0_add_69_carry_2_), 
        .A2(npu_inst_pe_1_7_0_int_q_acc_2_), .ZN(
        npu_inst_pe_1_7_0_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_7_0_U136 ( .A(npu_inst_pe_1_7_0_int_q_acc_3_), .B(
        npu_inst_pe_1_7_0_add_69_carry_3_), .Z(npu_inst_pe_1_7_0_N76) );
  AND2_X1 npu_inst_pe_1_7_0_U135 ( .A1(npu_inst_pe_1_7_0_add_69_carry_3_), 
        .A2(npu_inst_pe_1_7_0_int_q_acc_3_), .ZN(
        npu_inst_pe_1_7_0_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_7_0_U134 ( .A(npu_inst_pe_1_7_0_int_q_acc_4_), .B(
        npu_inst_pe_1_7_0_add_69_carry_4_), .Z(npu_inst_pe_1_7_0_N77) );
  AND2_X1 npu_inst_pe_1_7_0_U133 ( .A1(npu_inst_pe_1_7_0_add_69_carry_4_), 
        .A2(npu_inst_pe_1_7_0_int_q_acc_4_), .ZN(
        npu_inst_pe_1_7_0_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_7_0_U132 ( .A(npu_inst_pe_1_7_0_int_q_acc_5_), .B(
        npu_inst_pe_1_7_0_add_69_carry_5_), .Z(npu_inst_pe_1_7_0_N78) );
  AND2_X1 npu_inst_pe_1_7_0_U131 ( .A1(npu_inst_pe_1_7_0_add_69_carry_5_), 
        .A2(npu_inst_pe_1_7_0_int_q_acc_5_), .ZN(
        npu_inst_pe_1_7_0_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_7_0_U130 ( .A(npu_inst_pe_1_7_0_int_q_acc_6_), .B(
        npu_inst_pe_1_7_0_add_69_carry_6_), .Z(npu_inst_pe_1_7_0_N79) );
  AND2_X1 npu_inst_pe_1_7_0_U129 ( .A1(npu_inst_pe_1_7_0_add_69_carry_6_), 
        .A2(npu_inst_pe_1_7_0_int_q_acc_6_), .ZN(
        npu_inst_pe_1_7_0_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_7_0_U128 ( .A(npu_inst_pe_1_7_0_int_q_acc_7_), .B(
        npu_inst_pe_1_7_0_add_69_carry_7_), .Z(npu_inst_pe_1_7_0_N80) );
  XNOR2_X1 npu_inst_pe_1_7_0_U127 ( .A(npu_inst_pe_1_7_0_sub_67_carry_2_), .B(
        npu_inst_pe_1_7_0_int_q_acc_2_), .ZN(npu_inst_pe_1_7_0_N67) );
  OR2_X1 npu_inst_pe_1_7_0_U126 ( .A1(npu_inst_pe_1_7_0_int_q_acc_2_), .A2(
        npu_inst_pe_1_7_0_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_7_0_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_7_0_U125 ( .A(npu_inst_pe_1_7_0_sub_67_carry_3_), .B(
        npu_inst_pe_1_7_0_int_q_acc_3_), .ZN(npu_inst_pe_1_7_0_N68) );
  OR2_X1 npu_inst_pe_1_7_0_U124 ( .A1(npu_inst_pe_1_7_0_int_q_acc_3_), .A2(
        npu_inst_pe_1_7_0_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_7_0_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_7_0_U123 ( .A(npu_inst_pe_1_7_0_sub_67_carry_4_), .B(
        npu_inst_pe_1_7_0_int_q_acc_4_), .ZN(npu_inst_pe_1_7_0_N69) );
  OR2_X1 npu_inst_pe_1_7_0_U122 ( .A1(npu_inst_pe_1_7_0_int_q_acc_4_), .A2(
        npu_inst_pe_1_7_0_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_7_0_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_7_0_U121 ( .A(npu_inst_pe_1_7_0_sub_67_carry_5_), .B(
        npu_inst_pe_1_7_0_int_q_acc_5_), .ZN(npu_inst_pe_1_7_0_N70) );
  OR2_X1 npu_inst_pe_1_7_0_U120 ( .A1(npu_inst_pe_1_7_0_int_q_acc_5_), .A2(
        npu_inst_pe_1_7_0_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_7_0_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_7_0_U119 ( .A(npu_inst_pe_1_7_0_sub_67_carry_6_), .B(
        npu_inst_pe_1_7_0_int_q_acc_6_), .ZN(npu_inst_pe_1_7_0_N71) );
  OR2_X1 npu_inst_pe_1_7_0_U118 ( .A1(npu_inst_pe_1_7_0_int_q_acc_6_), .A2(
        npu_inst_pe_1_7_0_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_7_0_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_7_0_U117 ( .A(npu_inst_pe_1_7_0_int_q_acc_7_), .B(
        npu_inst_pe_1_7_0_sub_67_carry_7_), .ZN(npu_inst_pe_1_7_0_N72) );
  INV_X1 npu_inst_pe_1_7_0_U116 ( .A(npu_inst_n75), .ZN(npu_inst_pe_1_7_0_n7)
         );
  INV_X1 npu_inst_pe_1_7_0_U115 ( .A(npu_inst_pe_1_7_0_n7), .ZN(
        npu_inst_pe_1_7_0_n6) );
  INV_X1 npu_inst_pe_1_7_0_U114 ( .A(npu_inst_n53), .ZN(npu_inst_pe_1_7_0_n3)
         );
  AOI22_X1 npu_inst_pe_1_7_0_U113 ( .A1(npu_inst_pe_1_7_0_n38), .A2(
        int_i_data_v_npu[15]), .B1(npu_inst_pe_1_7_0_n114), .B2(
        npu_inst_pe_1_7_0_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_7_0_n39) );
  INV_X1 npu_inst_pe_1_7_0_U112 ( .A(npu_inst_pe_1_7_0_n39), .ZN(
        npu_inst_pe_1_7_0_n112) );
  AOI22_X1 npu_inst_pe_1_7_0_U111 ( .A1(npu_inst_pe_1_7_0_n38), .A2(
        int_i_data_v_npu[14]), .B1(npu_inst_pe_1_7_0_n114), .B2(
        npu_inst_pe_1_7_0_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_7_0_n37) );
  INV_X1 npu_inst_pe_1_7_0_U110 ( .A(npu_inst_pe_1_7_0_n37), .ZN(
        npu_inst_pe_1_7_0_n113) );
  AOI22_X1 npu_inst_pe_1_7_0_U107 ( .A1(int_i_data_v_npu[15]), .A2(
        npu_inst_pe_1_7_0_n58), .B1(npu_inst_pe_1_7_0_n119), .B2(
        npu_inst_pe_1_7_0_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_7_0_n59) );
  INV_X1 npu_inst_pe_1_7_0_U106 ( .A(npu_inst_pe_1_7_0_n59), .ZN(
        npu_inst_pe_1_7_0_n102) );
  AOI22_X1 npu_inst_pe_1_7_0_U105 ( .A1(int_i_data_v_npu[14]), .A2(
        npu_inst_pe_1_7_0_n58), .B1(npu_inst_pe_1_7_0_n119), .B2(
        npu_inst_pe_1_7_0_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_7_0_n57) );
  INV_X1 npu_inst_pe_1_7_0_U104 ( .A(npu_inst_pe_1_7_0_n57), .ZN(
        npu_inst_pe_1_7_0_n103) );
  AOI22_X1 npu_inst_pe_1_7_0_U103 ( .A1(int_i_data_v_npu[15]), .A2(
        npu_inst_pe_1_7_0_n54), .B1(npu_inst_pe_1_7_0_n118), .B2(
        npu_inst_pe_1_7_0_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_7_0_n55) );
  INV_X1 npu_inst_pe_1_7_0_U102 ( .A(npu_inst_pe_1_7_0_n55), .ZN(
        npu_inst_pe_1_7_0_n104) );
  AOI22_X1 npu_inst_pe_1_7_0_U101 ( .A1(int_i_data_v_npu[14]), .A2(
        npu_inst_pe_1_7_0_n54), .B1(npu_inst_pe_1_7_0_n118), .B2(
        npu_inst_pe_1_7_0_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_7_0_n53) );
  INV_X1 npu_inst_pe_1_7_0_U100 ( .A(npu_inst_pe_1_7_0_n53), .ZN(
        npu_inst_pe_1_7_0_n105) );
  AOI22_X1 npu_inst_pe_1_7_0_U99 ( .A1(int_i_data_v_npu[15]), .A2(
        npu_inst_pe_1_7_0_n50), .B1(npu_inst_pe_1_7_0_n117), .B2(
        npu_inst_pe_1_7_0_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_7_0_n51) );
  INV_X1 npu_inst_pe_1_7_0_U98 ( .A(npu_inst_pe_1_7_0_n51), .ZN(
        npu_inst_pe_1_7_0_n106) );
  AOI22_X1 npu_inst_pe_1_7_0_U97 ( .A1(int_i_data_v_npu[14]), .A2(
        npu_inst_pe_1_7_0_n50), .B1(npu_inst_pe_1_7_0_n117), .B2(
        npu_inst_pe_1_7_0_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_7_0_n49) );
  INV_X1 npu_inst_pe_1_7_0_U96 ( .A(npu_inst_pe_1_7_0_n49), .ZN(
        npu_inst_pe_1_7_0_n107) );
  AOI22_X1 npu_inst_pe_1_7_0_U95 ( .A1(int_i_data_v_npu[15]), .A2(
        npu_inst_pe_1_7_0_n46), .B1(npu_inst_pe_1_7_0_n116), .B2(
        npu_inst_pe_1_7_0_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_7_0_n47) );
  INV_X1 npu_inst_pe_1_7_0_U94 ( .A(npu_inst_pe_1_7_0_n47), .ZN(
        npu_inst_pe_1_7_0_n108) );
  AOI22_X1 npu_inst_pe_1_7_0_U93 ( .A1(int_i_data_v_npu[14]), .A2(
        npu_inst_pe_1_7_0_n46), .B1(npu_inst_pe_1_7_0_n116), .B2(
        npu_inst_pe_1_7_0_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_7_0_n45) );
  INV_X1 npu_inst_pe_1_7_0_U92 ( .A(npu_inst_pe_1_7_0_n45), .ZN(
        npu_inst_pe_1_7_0_n109) );
  AOI22_X1 npu_inst_pe_1_7_0_U91 ( .A1(int_i_data_v_npu[15]), .A2(
        npu_inst_pe_1_7_0_n42), .B1(npu_inst_pe_1_7_0_n115), .B2(
        npu_inst_pe_1_7_0_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_7_0_n43) );
  INV_X1 npu_inst_pe_1_7_0_U90 ( .A(npu_inst_pe_1_7_0_n43), .ZN(
        npu_inst_pe_1_7_0_n110) );
  AOI22_X1 npu_inst_pe_1_7_0_U89 ( .A1(int_i_data_v_npu[14]), .A2(
        npu_inst_pe_1_7_0_n42), .B1(npu_inst_pe_1_7_0_n115), .B2(
        npu_inst_pe_1_7_0_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_7_0_n41) );
  INV_X1 npu_inst_pe_1_7_0_U88 ( .A(npu_inst_pe_1_7_0_n41), .ZN(
        npu_inst_pe_1_7_0_n111) );
  NAND2_X1 npu_inst_pe_1_7_0_U87 ( .A1(npu_inst_pe_1_7_0_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_7_0_n60), .ZN(npu_inst_pe_1_7_0_n74) );
  OAI21_X1 npu_inst_pe_1_7_0_U86 ( .B1(npu_inst_pe_1_7_0_n63), .B2(
        npu_inst_pe_1_7_0_n60), .A(npu_inst_pe_1_7_0_n74), .ZN(
        npu_inst_pe_1_7_0_n97) );
  NAND2_X1 npu_inst_pe_1_7_0_U85 ( .A1(npu_inst_pe_1_7_0_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_7_0_n60), .ZN(npu_inst_pe_1_7_0_n73) );
  OAI21_X1 npu_inst_pe_1_7_0_U84 ( .B1(npu_inst_pe_1_7_0_n61), .B2(
        npu_inst_pe_1_7_0_n60), .A(npu_inst_pe_1_7_0_n73), .ZN(
        npu_inst_pe_1_7_0_n96) );
  NAND2_X1 npu_inst_pe_1_7_0_U83 ( .A1(npu_inst_pe_1_7_0_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_7_0_n56), .ZN(npu_inst_pe_1_7_0_n72) );
  OAI21_X1 npu_inst_pe_1_7_0_U82 ( .B1(npu_inst_pe_1_7_0_n63), .B2(
        npu_inst_pe_1_7_0_n56), .A(npu_inst_pe_1_7_0_n72), .ZN(
        npu_inst_pe_1_7_0_n95) );
  NAND2_X1 npu_inst_pe_1_7_0_U81 ( .A1(npu_inst_pe_1_7_0_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_7_0_n56), .ZN(npu_inst_pe_1_7_0_n71) );
  OAI21_X1 npu_inst_pe_1_7_0_U80 ( .B1(npu_inst_pe_1_7_0_n61), .B2(
        npu_inst_pe_1_7_0_n56), .A(npu_inst_pe_1_7_0_n71), .ZN(
        npu_inst_pe_1_7_0_n94) );
  NAND2_X1 npu_inst_pe_1_7_0_U79 ( .A1(npu_inst_pe_1_7_0_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_7_0_n52), .ZN(npu_inst_pe_1_7_0_n70) );
  OAI21_X1 npu_inst_pe_1_7_0_U78 ( .B1(npu_inst_pe_1_7_0_n63), .B2(
        npu_inst_pe_1_7_0_n52), .A(npu_inst_pe_1_7_0_n70), .ZN(
        npu_inst_pe_1_7_0_n93) );
  NAND2_X1 npu_inst_pe_1_7_0_U77 ( .A1(npu_inst_pe_1_7_0_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_7_0_n52), .ZN(npu_inst_pe_1_7_0_n69) );
  OAI21_X1 npu_inst_pe_1_7_0_U76 ( .B1(npu_inst_pe_1_7_0_n61), .B2(
        npu_inst_pe_1_7_0_n52), .A(npu_inst_pe_1_7_0_n69), .ZN(
        npu_inst_pe_1_7_0_n92) );
  NAND2_X1 npu_inst_pe_1_7_0_U75 ( .A1(npu_inst_pe_1_7_0_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_7_0_n48), .ZN(npu_inst_pe_1_7_0_n68) );
  OAI21_X1 npu_inst_pe_1_7_0_U74 ( .B1(npu_inst_pe_1_7_0_n63), .B2(
        npu_inst_pe_1_7_0_n48), .A(npu_inst_pe_1_7_0_n68), .ZN(
        npu_inst_pe_1_7_0_n91) );
  NAND2_X1 npu_inst_pe_1_7_0_U73 ( .A1(npu_inst_pe_1_7_0_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_7_0_n48), .ZN(npu_inst_pe_1_7_0_n67) );
  OAI21_X1 npu_inst_pe_1_7_0_U72 ( .B1(npu_inst_pe_1_7_0_n61), .B2(
        npu_inst_pe_1_7_0_n48), .A(npu_inst_pe_1_7_0_n67), .ZN(
        npu_inst_pe_1_7_0_n90) );
  NAND2_X1 npu_inst_pe_1_7_0_U71 ( .A1(npu_inst_pe_1_7_0_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_7_0_n44), .ZN(npu_inst_pe_1_7_0_n66) );
  OAI21_X1 npu_inst_pe_1_7_0_U70 ( .B1(npu_inst_pe_1_7_0_n63), .B2(
        npu_inst_pe_1_7_0_n44), .A(npu_inst_pe_1_7_0_n66), .ZN(
        npu_inst_pe_1_7_0_n89) );
  NAND2_X1 npu_inst_pe_1_7_0_U69 ( .A1(npu_inst_pe_1_7_0_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_7_0_n44), .ZN(npu_inst_pe_1_7_0_n65) );
  OAI21_X1 npu_inst_pe_1_7_0_U68 ( .B1(npu_inst_pe_1_7_0_n61), .B2(
        npu_inst_pe_1_7_0_n44), .A(npu_inst_pe_1_7_0_n65), .ZN(
        npu_inst_pe_1_7_0_n88) );
  NAND2_X1 npu_inst_pe_1_7_0_U67 ( .A1(npu_inst_pe_1_7_0_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_7_0_n40), .ZN(npu_inst_pe_1_7_0_n64) );
  OAI21_X1 npu_inst_pe_1_7_0_U66 ( .B1(npu_inst_pe_1_7_0_n63), .B2(
        npu_inst_pe_1_7_0_n40), .A(npu_inst_pe_1_7_0_n64), .ZN(
        npu_inst_pe_1_7_0_n87) );
  NAND2_X1 npu_inst_pe_1_7_0_U65 ( .A1(npu_inst_pe_1_7_0_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_7_0_n40), .ZN(npu_inst_pe_1_7_0_n62) );
  OAI21_X1 npu_inst_pe_1_7_0_U64 ( .B1(npu_inst_pe_1_7_0_n61), .B2(
        npu_inst_pe_1_7_0_n40), .A(npu_inst_pe_1_7_0_n62), .ZN(
        npu_inst_pe_1_7_0_n86) );
  AND2_X1 npu_inst_pe_1_7_0_U63 ( .A1(npu_inst_pe_1_7_0_N93), .A2(npu_inst_n53), .ZN(npu_inst_int_data_y_7__0__0_) );
  AND2_X1 npu_inst_pe_1_7_0_U62 ( .A1(npu_inst_n53), .A2(npu_inst_pe_1_7_0_N94), .ZN(npu_inst_int_data_y_7__0__1_) );
  AOI22_X1 npu_inst_pe_1_7_0_U61 ( .A1(npu_inst_n53), .A2(int_i_data_v_npu[15]), .B1(npu_inst_pe_1_7_0_n3), .B2(npu_inst_int_data_x_7__1__1_), .ZN(
        npu_inst_pe_1_7_0_n63) );
  AOI22_X1 npu_inst_pe_1_7_0_U60 ( .A1(npu_inst_n53), .A2(int_i_data_v_npu[14]), .B1(npu_inst_pe_1_7_0_n3), .B2(npu_inst_int_data_x_7__1__0_), .ZN(
        npu_inst_pe_1_7_0_n61) );
  AOI222_X1 npu_inst_pe_1_7_0_U59 ( .A1(1'b0), .A2(npu_inst_pe_1_7_0_n1), .B1(
        npu_inst_pe_1_7_0_N73), .B2(npu_inst_pe_1_7_0_n76), .C1(
        npu_inst_pe_1_7_0_N65), .C2(npu_inst_pe_1_7_0_n77), .ZN(
        npu_inst_pe_1_7_0_n84) );
  INV_X1 npu_inst_pe_1_7_0_U58 ( .A(npu_inst_pe_1_7_0_n84), .ZN(
        npu_inst_pe_1_7_0_n101) );
  AOI222_X1 npu_inst_pe_1_7_0_U57 ( .A1(1'b0), .A2(npu_inst_pe_1_7_0_n1), .B1(
        npu_inst_pe_1_7_0_N80), .B2(npu_inst_pe_1_7_0_n76), .C1(
        npu_inst_pe_1_7_0_N72), .C2(npu_inst_pe_1_7_0_n77), .ZN(
        npu_inst_pe_1_7_0_n75) );
  INV_X1 npu_inst_pe_1_7_0_U56 ( .A(npu_inst_pe_1_7_0_n75), .ZN(
        npu_inst_pe_1_7_0_n33) );
  AOI222_X1 npu_inst_pe_1_7_0_U55 ( .A1(1'b0), .A2(npu_inst_pe_1_7_0_n1), .B1(
        npu_inst_pe_1_7_0_N74), .B2(npu_inst_pe_1_7_0_n76), .C1(
        npu_inst_pe_1_7_0_N66), .C2(npu_inst_pe_1_7_0_n77), .ZN(
        npu_inst_pe_1_7_0_n83) );
  INV_X1 npu_inst_pe_1_7_0_U54 ( .A(npu_inst_pe_1_7_0_n83), .ZN(
        npu_inst_pe_1_7_0_n100) );
  AOI222_X1 npu_inst_pe_1_7_0_U53 ( .A1(1'b0), .A2(npu_inst_pe_1_7_0_n1), .B1(
        npu_inst_pe_1_7_0_N75), .B2(npu_inst_pe_1_7_0_n76), .C1(
        npu_inst_pe_1_7_0_N67), .C2(npu_inst_pe_1_7_0_n77), .ZN(
        npu_inst_pe_1_7_0_n82) );
  INV_X1 npu_inst_pe_1_7_0_U52 ( .A(npu_inst_pe_1_7_0_n82), .ZN(
        npu_inst_pe_1_7_0_n99) );
  AOI222_X1 npu_inst_pe_1_7_0_U51 ( .A1(1'b0), .A2(npu_inst_pe_1_7_0_n1), .B1(
        npu_inst_pe_1_7_0_N76), .B2(npu_inst_pe_1_7_0_n76), .C1(
        npu_inst_pe_1_7_0_N68), .C2(npu_inst_pe_1_7_0_n77), .ZN(
        npu_inst_pe_1_7_0_n81) );
  INV_X1 npu_inst_pe_1_7_0_U50 ( .A(npu_inst_pe_1_7_0_n81), .ZN(
        npu_inst_pe_1_7_0_n98) );
  AOI222_X1 npu_inst_pe_1_7_0_U49 ( .A1(1'b0), .A2(npu_inst_pe_1_7_0_n1), .B1(
        npu_inst_pe_1_7_0_N77), .B2(npu_inst_pe_1_7_0_n76), .C1(
        npu_inst_pe_1_7_0_N69), .C2(npu_inst_pe_1_7_0_n77), .ZN(
        npu_inst_pe_1_7_0_n80) );
  INV_X1 npu_inst_pe_1_7_0_U48 ( .A(npu_inst_pe_1_7_0_n80), .ZN(
        npu_inst_pe_1_7_0_n36) );
  AOI222_X1 npu_inst_pe_1_7_0_U47 ( .A1(1'b0), .A2(npu_inst_pe_1_7_0_n1), .B1(
        npu_inst_pe_1_7_0_N78), .B2(npu_inst_pe_1_7_0_n76), .C1(
        npu_inst_pe_1_7_0_N70), .C2(npu_inst_pe_1_7_0_n77), .ZN(
        npu_inst_pe_1_7_0_n79) );
  INV_X1 npu_inst_pe_1_7_0_U46 ( .A(npu_inst_pe_1_7_0_n79), .ZN(
        npu_inst_pe_1_7_0_n35) );
  AOI222_X1 npu_inst_pe_1_7_0_U45 ( .A1(1'b0), .A2(npu_inst_pe_1_7_0_n1), .B1(
        npu_inst_pe_1_7_0_N79), .B2(npu_inst_pe_1_7_0_n76), .C1(
        npu_inst_pe_1_7_0_N71), .C2(npu_inst_pe_1_7_0_n77), .ZN(
        npu_inst_pe_1_7_0_n78) );
  INV_X1 npu_inst_pe_1_7_0_U44 ( .A(npu_inst_pe_1_7_0_n78), .ZN(
        npu_inst_pe_1_7_0_n34) );
  AND2_X1 npu_inst_pe_1_7_0_U43 ( .A1(npu_inst_pe_1_7_0_int_q_acc_0_), .A2(
        npu_inst_pe_1_7_0_n1), .ZN(npu_inst_int_data_res_7__0__0_) );
  AND2_X1 npu_inst_pe_1_7_0_U42 ( .A1(npu_inst_pe_1_7_0_n2), .A2(
        npu_inst_pe_1_7_0_int_q_acc_7_), .ZN(npu_inst_int_data_res_7__0__7_)
         );
  AND2_X1 npu_inst_pe_1_7_0_U41 ( .A1(npu_inst_pe_1_7_0_int_q_acc_1_), .A2(
        npu_inst_pe_1_7_0_n1), .ZN(npu_inst_int_data_res_7__0__1_) );
  AND2_X1 npu_inst_pe_1_7_0_U40 ( .A1(npu_inst_pe_1_7_0_int_q_acc_2_), .A2(
        npu_inst_pe_1_7_0_n1), .ZN(npu_inst_int_data_res_7__0__2_) );
  AND2_X1 npu_inst_pe_1_7_0_U39 ( .A1(npu_inst_pe_1_7_0_int_q_acc_3_), .A2(
        npu_inst_pe_1_7_0_n2), .ZN(npu_inst_int_data_res_7__0__3_) );
  AND2_X1 npu_inst_pe_1_7_0_U38 ( .A1(npu_inst_pe_1_7_0_int_q_acc_4_), .A2(
        npu_inst_pe_1_7_0_n2), .ZN(npu_inst_int_data_res_7__0__4_) );
  AND2_X1 npu_inst_pe_1_7_0_U37 ( .A1(npu_inst_pe_1_7_0_int_q_acc_5_), .A2(
        npu_inst_pe_1_7_0_n2), .ZN(npu_inst_int_data_res_7__0__5_) );
  AND2_X1 npu_inst_pe_1_7_0_U36 ( .A1(npu_inst_pe_1_7_0_int_q_acc_6_), .A2(
        npu_inst_pe_1_7_0_n2), .ZN(npu_inst_int_data_res_7__0__6_) );
  INV_X1 npu_inst_pe_1_7_0_U35 ( .A(npu_inst_pe_1_7_0_int_data_1_), .ZN(
        npu_inst_pe_1_7_0_n14) );
  NOR3_X1 npu_inst_pe_1_7_0_U34 ( .A1(npu_inst_pe_1_7_0_n26), .A2(npu_inst_n53), .A3(npu_inst_int_ckg[7]), .ZN(npu_inst_pe_1_7_0_n85) );
  OR2_X1 npu_inst_pe_1_7_0_U33 ( .A1(npu_inst_pe_1_7_0_n85), .A2(
        npu_inst_pe_1_7_0_n2), .ZN(npu_inst_pe_1_7_0_N84) );
  AND2_X1 npu_inst_pe_1_7_0_U32 ( .A1(npu_inst_pe_1_7_0_o_data_h_1_), .A2(
        npu_inst_pe_1_7_0_int_q_weight_1_), .ZN(npu_inst_pe_1_7_0_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_7_0_U31 ( .A1(npu_inst_pe_1_7_0_o_data_h_0_), .A2(
        npu_inst_pe_1_7_0_int_q_weight_1_), .ZN(npu_inst_pe_1_7_0_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_7_0_U30 ( .A(npu_inst_pe_1_7_0_int_data_0_), .ZN(
        npu_inst_pe_1_7_0_n13) );
  INV_X1 npu_inst_pe_1_7_0_U29 ( .A(npu_inst_n67), .ZN(npu_inst_pe_1_7_0_n5)
         );
  OR3_X1 npu_inst_pe_1_7_0_U28 ( .A1(npu_inst_pe_1_7_0_n6), .A2(
        npu_inst_pe_1_7_0_n8), .A3(npu_inst_pe_1_7_0_n5), .ZN(
        npu_inst_pe_1_7_0_n56) );
  OR3_X1 npu_inst_pe_1_7_0_U27 ( .A1(npu_inst_pe_1_7_0_n5), .A2(
        npu_inst_pe_1_7_0_n8), .A3(npu_inst_pe_1_7_0_n7), .ZN(
        npu_inst_pe_1_7_0_n48) );
  INV_X1 npu_inst_pe_1_7_0_U26 ( .A(npu_inst_pe_1_7_0_n5), .ZN(
        npu_inst_pe_1_7_0_n4) );
  OR3_X1 npu_inst_pe_1_7_0_U25 ( .A1(npu_inst_pe_1_7_0_n4), .A2(
        npu_inst_pe_1_7_0_n8), .A3(npu_inst_pe_1_7_0_n7), .ZN(
        npu_inst_pe_1_7_0_n52) );
  OR3_X1 npu_inst_pe_1_7_0_U24 ( .A1(npu_inst_pe_1_7_0_n6), .A2(
        npu_inst_pe_1_7_0_n8), .A3(npu_inst_pe_1_7_0_n4), .ZN(
        npu_inst_pe_1_7_0_n60) );
  NOR2_X1 npu_inst_pe_1_7_0_U23 ( .A1(npu_inst_pe_1_7_0_n60), .A2(
        npu_inst_pe_1_7_0_n3), .ZN(npu_inst_pe_1_7_0_n58) );
  NOR2_X1 npu_inst_pe_1_7_0_U22 ( .A1(npu_inst_pe_1_7_0_n56), .A2(
        npu_inst_pe_1_7_0_n3), .ZN(npu_inst_pe_1_7_0_n54) );
  NOR2_X1 npu_inst_pe_1_7_0_U21 ( .A1(npu_inst_pe_1_7_0_n52), .A2(
        npu_inst_pe_1_7_0_n3), .ZN(npu_inst_pe_1_7_0_n50) );
  NOR2_X1 npu_inst_pe_1_7_0_U20 ( .A1(npu_inst_pe_1_7_0_n48), .A2(
        npu_inst_pe_1_7_0_n3), .ZN(npu_inst_pe_1_7_0_n46) );
  NOR2_X1 npu_inst_pe_1_7_0_U19 ( .A1(npu_inst_pe_1_7_0_n40), .A2(
        npu_inst_pe_1_7_0_n3), .ZN(npu_inst_pe_1_7_0_n38) );
  NOR2_X1 npu_inst_pe_1_7_0_U18 ( .A1(npu_inst_pe_1_7_0_n44), .A2(
        npu_inst_pe_1_7_0_n3), .ZN(npu_inst_pe_1_7_0_n42) );
  BUF_X1 npu_inst_pe_1_7_0_U17 ( .A(npu_inst_n93), .Z(npu_inst_pe_1_7_0_n8) );
  INV_X1 npu_inst_pe_1_7_0_U16 ( .A(npu_inst_n122), .ZN(npu_inst_pe_1_7_0_n12)
         );
  INV_X1 npu_inst_pe_1_7_0_U15 ( .A(npu_inst_pe_1_7_0_n38), .ZN(
        npu_inst_pe_1_7_0_n114) );
  INV_X1 npu_inst_pe_1_7_0_U14 ( .A(npu_inst_pe_1_7_0_n58), .ZN(
        npu_inst_pe_1_7_0_n119) );
  INV_X1 npu_inst_pe_1_7_0_U13 ( .A(npu_inst_pe_1_7_0_n54), .ZN(
        npu_inst_pe_1_7_0_n118) );
  INV_X1 npu_inst_pe_1_7_0_U12 ( .A(npu_inst_pe_1_7_0_n50), .ZN(
        npu_inst_pe_1_7_0_n117) );
  INV_X1 npu_inst_pe_1_7_0_U11 ( .A(npu_inst_pe_1_7_0_n46), .ZN(
        npu_inst_pe_1_7_0_n116) );
  INV_X1 npu_inst_pe_1_7_0_U10 ( .A(npu_inst_pe_1_7_0_n42), .ZN(
        npu_inst_pe_1_7_0_n115) );
  BUF_X1 npu_inst_pe_1_7_0_U9 ( .A(npu_inst_n10), .Z(npu_inst_pe_1_7_0_n2) );
  BUF_X1 npu_inst_pe_1_7_0_U8 ( .A(npu_inst_n10), .Z(npu_inst_pe_1_7_0_n1) );
  BUF_X1 npu_inst_pe_1_7_0_U7 ( .A(npu_inst_pe_1_7_0_n12), .Z(
        npu_inst_pe_1_7_0_n11) );
  BUF_X1 npu_inst_pe_1_7_0_U6 ( .A(npu_inst_pe_1_7_0_n12), .Z(
        npu_inst_pe_1_7_0_n10) );
  BUF_X1 npu_inst_pe_1_7_0_U5 ( .A(npu_inst_pe_1_7_0_n12), .Z(
        npu_inst_pe_1_7_0_n9) );
  NOR2_X1 npu_inst_pe_1_7_0_U4 ( .A1(npu_inst_pe_1_7_0_int_q_weight_0_), .A2(
        npu_inst_pe_1_7_0_n1), .ZN(npu_inst_pe_1_7_0_n76) );
  NOR2_X1 npu_inst_pe_1_7_0_U3 ( .A1(npu_inst_pe_1_7_0_n27), .A2(
        npu_inst_pe_1_7_0_n1), .ZN(npu_inst_pe_1_7_0_n77) );
  FA_X1 npu_inst_pe_1_7_0_sub_67_U2_1 ( .A(npu_inst_pe_1_7_0_int_q_acc_1_), 
        .B(npu_inst_pe_1_7_0_n14), .CI(npu_inst_pe_1_7_0_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_7_0_sub_67_carry_2_), .S(npu_inst_pe_1_7_0_N66) );
  FA_X1 npu_inst_pe_1_7_0_add_69_U1_1 ( .A(npu_inst_pe_1_7_0_int_q_acc_1_), 
        .B(npu_inst_pe_1_7_0_int_data_1_), .CI(
        npu_inst_pe_1_7_0_add_69_carry_1_), .CO(
        npu_inst_pe_1_7_0_add_69_carry_2_), .S(npu_inst_pe_1_7_0_N74) );
  NAND3_X1 npu_inst_pe_1_7_0_U109 ( .A1(npu_inst_pe_1_7_0_n5), .A2(
        npu_inst_pe_1_7_0_n7), .A3(npu_inst_pe_1_7_0_n8), .ZN(
        npu_inst_pe_1_7_0_n44) );
  NAND3_X1 npu_inst_pe_1_7_0_U108 ( .A1(npu_inst_pe_1_7_0_n4), .A2(
        npu_inst_pe_1_7_0_n7), .A3(npu_inst_pe_1_7_0_n8), .ZN(
        npu_inst_pe_1_7_0_n40) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_7_0_n34), .CK(
        npu_inst_pe_1_7_0_net3274), .RN(npu_inst_pe_1_7_0_n9), .Q(
        npu_inst_pe_1_7_0_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_7_0_n35), .CK(
        npu_inst_pe_1_7_0_net3274), .RN(npu_inst_pe_1_7_0_n9), .Q(
        npu_inst_pe_1_7_0_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_7_0_n36), .CK(
        npu_inst_pe_1_7_0_net3274), .RN(npu_inst_pe_1_7_0_n9), .Q(
        npu_inst_pe_1_7_0_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_7_0_n98), .CK(
        npu_inst_pe_1_7_0_net3274), .RN(npu_inst_pe_1_7_0_n9), .Q(
        npu_inst_pe_1_7_0_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_7_0_n99), .CK(
        npu_inst_pe_1_7_0_net3274), .RN(npu_inst_pe_1_7_0_n9), .Q(
        npu_inst_pe_1_7_0_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_7_0_n100), 
        .CK(npu_inst_pe_1_7_0_net3274), .RN(npu_inst_pe_1_7_0_n9), .Q(
        npu_inst_pe_1_7_0_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_7_0_n33), .CK(
        npu_inst_pe_1_7_0_net3274), .RN(npu_inst_pe_1_7_0_n9), .Q(
        npu_inst_pe_1_7_0_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_7_0_n101), 
        .CK(npu_inst_pe_1_7_0_net3274), .RN(npu_inst_pe_1_7_0_n9), .Q(
        npu_inst_pe_1_7_0_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_weight_reg_0_ ( .D(npu_inst_n108), .CK(
        npu_inst_pe_1_7_0_net3280), .RN(npu_inst_pe_1_7_0_n9), .Q(
        npu_inst_pe_1_7_0_int_q_weight_0_), .QN(npu_inst_pe_1_7_0_n27) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_weight_reg_1_ ( .D(npu_inst_n114), .CK(
        npu_inst_pe_1_7_0_net3280), .RN(npu_inst_pe_1_7_0_n9), .Q(
        npu_inst_pe_1_7_0_int_q_weight_1_), .QN(npu_inst_pe_1_7_0_n26) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_7_0_n113), 
        .CK(npu_inst_pe_1_7_0_net3280), .RN(npu_inst_pe_1_7_0_n9), .Q(
        npu_inst_pe_1_7_0_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_7_0_n112), 
        .CK(npu_inst_pe_1_7_0_net3280), .RN(npu_inst_pe_1_7_0_n9), .Q(
        npu_inst_pe_1_7_0_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_7_0_n111), 
        .CK(npu_inst_pe_1_7_0_net3280), .RN(npu_inst_pe_1_7_0_n10), .Q(
        npu_inst_pe_1_7_0_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_7_0_n110), 
        .CK(npu_inst_pe_1_7_0_net3280), .RN(npu_inst_pe_1_7_0_n10), .Q(
        npu_inst_pe_1_7_0_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_7_0_n109), 
        .CK(npu_inst_pe_1_7_0_net3280), .RN(npu_inst_pe_1_7_0_n10), .Q(
        npu_inst_pe_1_7_0_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_7_0_n108), 
        .CK(npu_inst_pe_1_7_0_net3280), .RN(npu_inst_pe_1_7_0_n10), .Q(
        npu_inst_pe_1_7_0_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_7_0_n107), 
        .CK(npu_inst_pe_1_7_0_net3280), .RN(npu_inst_pe_1_7_0_n10), .Q(
        npu_inst_pe_1_7_0_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_7_0_n106), 
        .CK(npu_inst_pe_1_7_0_net3280), .RN(npu_inst_pe_1_7_0_n10), .Q(
        npu_inst_pe_1_7_0_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_7_0_n105), 
        .CK(npu_inst_pe_1_7_0_net3280), .RN(npu_inst_pe_1_7_0_n10), .Q(
        npu_inst_pe_1_7_0_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_7_0_n104), 
        .CK(npu_inst_pe_1_7_0_net3280), .RN(npu_inst_pe_1_7_0_n10), .Q(
        npu_inst_pe_1_7_0_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_7_0_n103), 
        .CK(npu_inst_pe_1_7_0_net3280), .RN(npu_inst_pe_1_7_0_n10), .Q(
        npu_inst_pe_1_7_0_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_7_0_n102), 
        .CK(npu_inst_pe_1_7_0_net3280), .RN(npu_inst_pe_1_7_0_n10), .Q(
        npu_inst_pe_1_7_0_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_7_0_n86), 
        .CK(npu_inst_pe_1_7_0_net3280), .RN(npu_inst_pe_1_7_0_n10), .Q(
        npu_inst_pe_1_7_0_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_7_0_n87), 
        .CK(npu_inst_pe_1_7_0_net3280), .RN(npu_inst_pe_1_7_0_n10), .Q(
        npu_inst_pe_1_7_0_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_7_0_n88), 
        .CK(npu_inst_pe_1_7_0_net3280), .RN(npu_inst_pe_1_7_0_n11), .Q(
        npu_inst_pe_1_7_0_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_7_0_n89), 
        .CK(npu_inst_pe_1_7_0_net3280), .RN(npu_inst_pe_1_7_0_n11), .Q(
        npu_inst_pe_1_7_0_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_7_0_n90), 
        .CK(npu_inst_pe_1_7_0_net3280), .RN(npu_inst_pe_1_7_0_n11), .Q(
        npu_inst_pe_1_7_0_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_7_0_n91), 
        .CK(npu_inst_pe_1_7_0_net3280), .RN(npu_inst_pe_1_7_0_n11), .Q(
        npu_inst_pe_1_7_0_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_7_0_n92), 
        .CK(npu_inst_pe_1_7_0_net3280), .RN(npu_inst_pe_1_7_0_n11), .Q(
        npu_inst_pe_1_7_0_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_7_0_n93), 
        .CK(npu_inst_pe_1_7_0_net3280), .RN(npu_inst_pe_1_7_0_n11), .Q(
        npu_inst_pe_1_7_0_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_7_0_n94), 
        .CK(npu_inst_pe_1_7_0_net3280), .RN(npu_inst_pe_1_7_0_n11), .Q(
        npu_inst_pe_1_7_0_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_7_0_n95), 
        .CK(npu_inst_pe_1_7_0_net3280), .RN(npu_inst_pe_1_7_0_n11), .Q(
        npu_inst_pe_1_7_0_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_7_0_n96), 
        .CK(npu_inst_pe_1_7_0_net3280), .RN(npu_inst_pe_1_7_0_n11), .Q(
        npu_inst_pe_1_7_0_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_7_0_n97), 
        .CK(npu_inst_pe_1_7_0_net3280), .RN(npu_inst_pe_1_7_0_n11), .Q(
        npu_inst_pe_1_7_0_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_7_0_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_7_0_N84), .SE(1'b0), .GCK(npu_inst_pe_1_7_0_net3274) );
  CLKGATETST_X1 npu_inst_pe_1_7_0_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n61), .SE(1'b0), .GCK(npu_inst_pe_1_7_0_net3280) );
  MUX2_X1 npu_inst_pe_1_7_1_U162 ( .A(npu_inst_pe_1_7_1_n32), .B(
        npu_inst_pe_1_7_1_n29), .S(npu_inst_pe_1_7_1_n8), .Z(
        npu_inst_pe_1_7_1_N93) );
  MUX2_X1 npu_inst_pe_1_7_1_U161 ( .A(npu_inst_pe_1_7_1_n31), .B(
        npu_inst_pe_1_7_1_n30), .S(npu_inst_pe_1_7_1_n6), .Z(
        npu_inst_pe_1_7_1_n32) );
  MUX2_X1 npu_inst_pe_1_7_1_U160 ( .A(npu_inst_pe_1_7_1_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_7_1_int_q_reg_v_1__0_), .S(npu_inst_pe_1_7_1_n4), .Z(
        npu_inst_pe_1_7_1_n31) );
  MUX2_X1 npu_inst_pe_1_7_1_U159 ( .A(npu_inst_pe_1_7_1_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_7_1_int_q_reg_v_3__0_), .S(npu_inst_pe_1_7_1_n4), .Z(
        npu_inst_pe_1_7_1_n30) );
  MUX2_X1 npu_inst_pe_1_7_1_U158 ( .A(npu_inst_pe_1_7_1_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_7_1_int_q_reg_v_5__0_), .S(npu_inst_pe_1_7_1_n4), .Z(
        npu_inst_pe_1_7_1_n29) );
  MUX2_X1 npu_inst_pe_1_7_1_U157 ( .A(npu_inst_pe_1_7_1_n28), .B(
        npu_inst_pe_1_7_1_n23), .S(npu_inst_pe_1_7_1_n8), .Z(
        npu_inst_pe_1_7_1_N94) );
  MUX2_X1 npu_inst_pe_1_7_1_U156 ( .A(npu_inst_pe_1_7_1_n25), .B(
        npu_inst_pe_1_7_1_n24), .S(npu_inst_pe_1_7_1_n6), .Z(
        npu_inst_pe_1_7_1_n28) );
  MUX2_X1 npu_inst_pe_1_7_1_U155 ( .A(npu_inst_pe_1_7_1_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_7_1_int_q_reg_v_1__1_), .S(npu_inst_pe_1_7_1_n4), .Z(
        npu_inst_pe_1_7_1_n25) );
  MUX2_X1 npu_inst_pe_1_7_1_U154 ( .A(npu_inst_pe_1_7_1_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_7_1_int_q_reg_v_3__1_), .S(npu_inst_pe_1_7_1_n4), .Z(
        npu_inst_pe_1_7_1_n24) );
  MUX2_X1 npu_inst_pe_1_7_1_U153 ( .A(npu_inst_pe_1_7_1_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_7_1_int_q_reg_v_5__1_), .S(npu_inst_pe_1_7_1_n4), .Z(
        npu_inst_pe_1_7_1_n23) );
  MUX2_X1 npu_inst_pe_1_7_1_U152 ( .A(npu_inst_pe_1_7_1_n22), .B(
        npu_inst_pe_1_7_1_n19), .S(npu_inst_pe_1_7_1_n8), .Z(
        npu_inst_int_data_x_7__1__1_) );
  MUX2_X1 npu_inst_pe_1_7_1_U151 ( .A(npu_inst_pe_1_7_1_n21), .B(
        npu_inst_pe_1_7_1_n20), .S(npu_inst_pe_1_7_1_n6), .Z(
        npu_inst_pe_1_7_1_n22) );
  MUX2_X1 npu_inst_pe_1_7_1_U150 ( .A(npu_inst_pe_1_7_1_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_7_1_int_q_reg_h_1__1_), .S(npu_inst_pe_1_7_1_n4), .Z(
        npu_inst_pe_1_7_1_n21) );
  MUX2_X1 npu_inst_pe_1_7_1_U149 ( .A(npu_inst_pe_1_7_1_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_7_1_int_q_reg_h_3__1_), .S(npu_inst_pe_1_7_1_n4), .Z(
        npu_inst_pe_1_7_1_n20) );
  MUX2_X1 npu_inst_pe_1_7_1_U148 ( .A(npu_inst_pe_1_7_1_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_7_1_int_q_reg_h_5__1_), .S(npu_inst_pe_1_7_1_n4), .Z(
        npu_inst_pe_1_7_1_n19) );
  MUX2_X1 npu_inst_pe_1_7_1_U147 ( .A(npu_inst_pe_1_7_1_n18), .B(
        npu_inst_pe_1_7_1_n15), .S(npu_inst_pe_1_7_1_n8), .Z(
        npu_inst_int_data_x_7__1__0_) );
  MUX2_X1 npu_inst_pe_1_7_1_U146 ( .A(npu_inst_pe_1_7_1_n17), .B(
        npu_inst_pe_1_7_1_n16), .S(npu_inst_pe_1_7_1_n6), .Z(
        npu_inst_pe_1_7_1_n18) );
  MUX2_X1 npu_inst_pe_1_7_1_U145 ( .A(npu_inst_pe_1_7_1_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_7_1_int_q_reg_h_1__0_), .S(npu_inst_pe_1_7_1_n4), .Z(
        npu_inst_pe_1_7_1_n17) );
  MUX2_X1 npu_inst_pe_1_7_1_U144 ( .A(npu_inst_pe_1_7_1_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_7_1_int_q_reg_h_3__0_), .S(npu_inst_pe_1_7_1_n4), .Z(
        npu_inst_pe_1_7_1_n16) );
  MUX2_X1 npu_inst_pe_1_7_1_U143 ( .A(npu_inst_pe_1_7_1_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_7_1_int_q_reg_h_5__0_), .S(npu_inst_pe_1_7_1_n4), .Z(
        npu_inst_pe_1_7_1_n15) );
  XOR2_X1 npu_inst_pe_1_7_1_U142 ( .A(npu_inst_pe_1_7_1_int_data_0_), .B(
        npu_inst_pe_1_7_1_int_q_acc_0_), .Z(npu_inst_pe_1_7_1_N73) );
  AND2_X1 npu_inst_pe_1_7_1_U141 ( .A1(npu_inst_pe_1_7_1_int_q_acc_0_), .A2(
        npu_inst_pe_1_7_1_int_data_0_), .ZN(npu_inst_pe_1_7_1_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_7_1_U140 ( .A(npu_inst_pe_1_7_1_int_q_acc_0_), .B(
        npu_inst_pe_1_7_1_n13), .ZN(npu_inst_pe_1_7_1_N65) );
  OR2_X1 npu_inst_pe_1_7_1_U139 ( .A1(npu_inst_pe_1_7_1_n13), .A2(
        npu_inst_pe_1_7_1_int_q_acc_0_), .ZN(npu_inst_pe_1_7_1_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_7_1_U138 ( .A(npu_inst_pe_1_7_1_int_q_acc_2_), .B(
        npu_inst_pe_1_7_1_add_69_carry_2_), .Z(npu_inst_pe_1_7_1_N75) );
  AND2_X1 npu_inst_pe_1_7_1_U137 ( .A1(npu_inst_pe_1_7_1_add_69_carry_2_), 
        .A2(npu_inst_pe_1_7_1_int_q_acc_2_), .ZN(
        npu_inst_pe_1_7_1_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_7_1_U136 ( .A(npu_inst_pe_1_7_1_int_q_acc_3_), .B(
        npu_inst_pe_1_7_1_add_69_carry_3_), .Z(npu_inst_pe_1_7_1_N76) );
  AND2_X1 npu_inst_pe_1_7_1_U135 ( .A1(npu_inst_pe_1_7_1_add_69_carry_3_), 
        .A2(npu_inst_pe_1_7_1_int_q_acc_3_), .ZN(
        npu_inst_pe_1_7_1_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_7_1_U134 ( .A(npu_inst_pe_1_7_1_int_q_acc_4_), .B(
        npu_inst_pe_1_7_1_add_69_carry_4_), .Z(npu_inst_pe_1_7_1_N77) );
  AND2_X1 npu_inst_pe_1_7_1_U133 ( .A1(npu_inst_pe_1_7_1_add_69_carry_4_), 
        .A2(npu_inst_pe_1_7_1_int_q_acc_4_), .ZN(
        npu_inst_pe_1_7_1_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_7_1_U132 ( .A(npu_inst_pe_1_7_1_int_q_acc_5_), .B(
        npu_inst_pe_1_7_1_add_69_carry_5_), .Z(npu_inst_pe_1_7_1_N78) );
  AND2_X1 npu_inst_pe_1_7_1_U131 ( .A1(npu_inst_pe_1_7_1_add_69_carry_5_), 
        .A2(npu_inst_pe_1_7_1_int_q_acc_5_), .ZN(
        npu_inst_pe_1_7_1_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_7_1_U130 ( .A(npu_inst_pe_1_7_1_int_q_acc_6_), .B(
        npu_inst_pe_1_7_1_add_69_carry_6_), .Z(npu_inst_pe_1_7_1_N79) );
  AND2_X1 npu_inst_pe_1_7_1_U129 ( .A1(npu_inst_pe_1_7_1_add_69_carry_6_), 
        .A2(npu_inst_pe_1_7_1_int_q_acc_6_), .ZN(
        npu_inst_pe_1_7_1_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_7_1_U128 ( .A(npu_inst_pe_1_7_1_int_q_acc_7_), .B(
        npu_inst_pe_1_7_1_add_69_carry_7_), .Z(npu_inst_pe_1_7_1_N80) );
  XNOR2_X1 npu_inst_pe_1_7_1_U127 ( .A(npu_inst_pe_1_7_1_sub_67_carry_2_), .B(
        npu_inst_pe_1_7_1_int_q_acc_2_), .ZN(npu_inst_pe_1_7_1_N67) );
  OR2_X1 npu_inst_pe_1_7_1_U126 ( .A1(npu_inst_pe_1_7_1_int_q_acc_2_), .A2(
        npu_inst_pe_1_7_1_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_7_1_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_7_1_U125 ( .A(npu_inst_pe_1_7_1_sub_67_carry_3_), .B(
        npu_inst_pe_1_7_1_int_q_acc_3_), .ZN(npu_inst_pe_1_7_1_N68) );
  OR2_X1 npu_inst_pe_1_7_1_U124 ( .A1(npu_inst_pe_1_7_1_int_q_acc_3_), .A2(
        npu_inst_pe_1_7_1_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_7_1_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_7_1_U123 ( .A(npu_inst_pe_1_7_1_sub_67_carry_4_), .B(
        npu_inst_pe_1_7_1_int_q_acc_4_), .ZN(npu_inst_pe_1_7_1_N69) );
  OR2_X1 npu_inst_pe_1_7_1_U122 ( .A1(npu_inst_pe_1_7_1_int_q_acc_4_), .A2(
        npu_inst_pe_1_7_1_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_7_1_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_7_1_U121 ( .A(npu_inst_pe_1_7_1_sub_67_carry_5_), .B(
        npu_inst_pe_1_7_1_int_q_acc_5_), .ZN(npu_inst_pe_1_7_1_N70) );
  OR2_X1 npu_inst_pe_1_7_1_U120 ( .A1(npu_inst_pe_1_7_1_int_q_acc_5_), .A2(
        npu_inst_pe_1_7_1_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_7_1_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_7_1_U119 ( .A(npu_inst_pe_1_7_1_sub_67_carry_6_), .B(
        npu_inst_pe_1_7_1_int_q_acc_6_), .ZN(npu_inst_pe_1_7_1_N71) );
  OR2_X1 npu_inst_pe_1_7_1_U118 ( .A1(npu_inst_pe_1_7_1_int_q_acc_6_), .A2(
        npu_inst_pe_1_7_1_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_7_1_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_7_1_U117 ( .A(npu_inst_pe_1_7_1_int_q_acc_7_), .B(
        npu_inst_pe_1_7_1_sub_67_carry_7_), .ZN(npu_inst_pe_1_7_1_N72) );
  INV_X1 npu_inst_pe_1_7_1_U116 ( .A(npu_inst_n75), .ZN(npu_inst_pe_1_7_1_n7)
         );
  INV_X1 npu_inst_pe_1_7_1_U115 ( .A(npu_inst_pe_1_7_1_n7), .ZN(
        npu_inst_pe_1_7_1_n6) );
  INV_X1 npu_inst_pe_1_7_1_U114 ( .A(npu_inst_n52), .ZN(npu_inst_pe_1_7_1_n3)
         );
  AOI22_X1 npu_inst_pe_1_7_1_U113 ( .A1(npu_inst_pe_1_7_1_n38), .A2(
        int_i_data_v_npu[13]), .B1(npu_inst_pe_1_7_1_n114), .B2(
        npu_inst_pe_1_7_1_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_7_1_n39) );
  INV_X1 npu_inst_pe_1_7_1_U112 ( .A(npu_inst_pe_1_7_1_n39), .ZN(
        npu_inst_pe_1_7_1_n112) );
  AOI22_X1 npu_inst_pe_1_7_1_U111 ( .A1(npu_inst_pe_1_7_1_n38), .A2(
        int_i_data_v_npu[12]), .B1(npu_inst_pe_1_7_1_n114), .B2(
        npu_inst_pe_1_7_1_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_7_1_n37) );
  INV_X1 npu_inst_pe_1_7_1_U110 ( .A(npu_inst_pe_1_7_1_n37), .ZN(
        npu_inst_pe_1_7_1_n113) );
  AOI22_X1 npu_inst_pe_1_7_1_U107 ( .A1(int_i_data_v_npu[13]), .A2(
        npu_inst_pe_1_7_1_n58), .B1(npu_inst_pe_1_7_1_n119), .B2(
        npu_inst_pe_1_7_1_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_7_1_n59) );
  INV_X1 npu_inst_pe_1_7_1_U106 ( .A(npu_inst_pe_1_7_1_n59), .ZN(
        npu_inst_pe_1_7_1_n102) );
  AOI22_X1 npu_inst_pe_1_7_1_U105 ( .A1(int_i_data_v_npu[12]), .A2(
        npu_inst_pe_1_7_1_n58), .B1(npu_inst_pe_1_7_1_n119), .B2(
        npu_inst_pe_1_7_1_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_7_1_n57) );
  INV_X1 npu_inst_pe_1_7_1_U104 ( .A(npu_inst_pe_1_7_1_n57), .ZN(
        npu_inst_pe_1_7_1_n103) );
  AOI22_X1 npu_inst_pe_1_7_1_U103 ( .A1(int_i_data_v_npu[13]), .A2(
        npu_inst_pe_1_7_1_n54), .B1(npu_inst_pe_1_7_1_n118), .B2(
        npu_inst_pe_1_7_1_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_7_1_n55) );
  INV_X1 npu_inst_pe_1_7_1_U102 ( .A(npu_inst_pe_1_7_1_n55), .ZN(
        npu_inst_pe_1_7_1_n104) );
  AOI22_X1 npu_inst_pe_1_7_1_U101 ( .A1(int_i_data_v_npu[12]), .A2(
        npu_inst_pe_1_7_1_n54), .B1(npu_inst_pe_1_7_1_n118), .B2(
        npu_inst_pe_1_7_1_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_7_1_n53) );
  INV_X1 npu_inst_pe_1_7_1_U100 ( .A(npu_inst_pe_1_7_1_n53), .ZN(
        npu_inst_pe_1_7_1_n105) );
  AOI22_X1 npu_inst_pe_1_7_1_U99 ( .A1(int_i_data_v_npu[13]), .A2(
        npu_inst_pe_1_7_1_n50), .B1(npu_inst_pe_1_7_1_n117), .B2(
        npu_inst_pe_1_7_1_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_7_1_n51) );
  INV_X1 npu_inst_pe_1_7_1_U98 ( .A(npu_inst_pe_1_7_1_n51), .ZN(
        npu_inst_pe_1_7_1_n106) );
  AOI22_X1 npu_inst_pe_1_7_1_U97 ( .A1(int_i_data_v_npu[12]), .A2(
        npu_inst_pe_1_7_1_n50), .B1(npu_inst_pe_1_7_1_n117), .B2(
        npu_inst_pe_1_7_1_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_7_1_n49) );
  INV_X1 npu_inst_pe_1_7_1_U96 ( .A(npu_inst_pe_1_7_1_n49), .ZN(
        npu_inst_pe_1_7_1_n107) );
  AOI22_X1 npu_inst_pe_1_7_1_U95 ( .A1(int_i_data_v_npu[13]), .A2(
        npu_inst_pe_1_7_1_n46), .B1(npu_inst_pe_1_7_1_n116), .B2(
        npu_inst_pe_1_7_1_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_7_1_n47) );
  INV_X1 npu_inst_pe_1_7_1_U94 ( .A(npu_inst_pe_1_7_1_n47), .ZN(
        npu_inst_pe_1_7_1_n108) );
  AOI22_X1 npu_inst_pe_1_7_1_U93 ( .A1(int_i_data_v_npu[12]), .A2(
        npu_inst_pe_1_7_1_n46), .B1(npu_inst_pe_1_7_1_n116), .B2(
        npu_inst_pe_1_7_1_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_7_1_n45) );
  INV_X1 npu_inst_pe_1_7_1_U92 ( .A(npu_inst_pe_1_7_1_n45), .ZN(
        npu_inst_pe_1_7_1_n109) );
  AOI22_X1 npu_inst_pe_1_7_1_U91 ( .A1(int_i_data_v_npu[13]), .A2(
        npu_inst_pe_1_7_1_n42), .B1(npu_inst_pe_1_7_1_n115), .B2(
        npu_inst_pe_1_7_1_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_7_1_n43) );
  INV_X1 npu_inst_pe_1_7_1_U90 ( .A(npu_inst_pe_1_7_1_n43), .ZN(
        npu_inst_pe_1_7_1_n110) );
  AOI22_X1 npu_inst_pe_1_7_1_U89 ( .A1(int_i_data_v_npu[12]), .A2(
        npu_inst_pe_1_7_1_n42), .B1(npu_inst_pe_1_7_1_n115), .B2(
        npu_inst_pe_1_7_1_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_7_1_n41) );
  INV_X1 npu_inst_pe_1_7_1_U88 ( .A(npu_inst_pe_1_7_1_n41), .ZN(
        npu_inst_pe_1_7_1_n111) );
  NAND2_X1 npu_inst_pe_1_7_1_U87 ( .A1(npu_inst_pe_1_7_1_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_7_1_n60), .ZN(npu_inst_pe_1_7_1_n74) );
  OAI21_X1 npu_inst_pe_1_7_1_U86 ( .B1(npu_inst_pe_1_7_1_n63), .B2(
        npu_inst_pe_1_7_1_n60), .A(npu_inst_pe_1_7_1_n74), .ZN(
        npu_inst_pe_1_7_1_n97) );
  NAND2_X1 npu_inst_pe_1_7_1_U85 ( .A1(npu_inst_pe_1_7_1_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_7_1_n60), .ZN(npu_inst_pe_1_7_1_n73) );
  OAI21_X1 npu_inst_pe_1_7_1_U84 ( .B1(npu_inst_pe_1_7_1_n61), .B2(
        npu_inst_pe_1_7_1_n60), .A(npu_inst_pe_1_7_1_n73), .ZN(
        npu_inst_pe_1_7_1_n96) );
  NAND2_X1 npu_inst_pe_1_7_1_U83 ( .A1(npu_inst_pe_1_7_1_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_7_1_n56), .ZN(npu_inst_pe_1_7_1_n72) );
  OAI21_X1 npu_inst_pe_1_7_1_U82 ( .B1(npu_inst_pe_1_7_1_n63), .B2(
        npu_inst_pe_1_7_1_n56), .A(npu_inst_pe_1_7_1_n72), .ZN(
        npu_inst_pe_1_7_1_n95) );
  NAND2_X1 npu_inst_pe_1_7_1_U81 ( .A1(npu_inst_pe_1_7_1_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_7_1_n56), .ZN(npu_inst_pe_1_7_1_n71) );
  OAI21_X1 npu_inst_pe_1_7_1_U80 ( .B1(npu_inst_pe_1_7_1_n61), .B2(
        npu_inst_pe_1_7_1_n56), .A(npu_inst_pe_1_7_1_n71), .ZN(
        npu_inst_pe_1_7_1_n94) );
  NAND2_X1 npu_inst_pe_1_7_1_U79 ( .A1(npu_inst_pe_1_7_1_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_7_1_n52), .ZN(npu_inst_pe_1_7_1_n70) );
  OAI21_X1 npu_inst_pe_1_7_1_U78 ( .B1(npu_inst_pe_1_7_1_n63), .B2(
        npu_inst_pe_1_7_1_n52), .A(npu_inst_pe_1_7_1_n70), .ZN(
        npu_inst_pe_1_7_1_n93) );
  NAND2_X1 npu_inst_pe_1_7_1_U77 ( .A1(npu_inst_pe_1_7_1_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_7_1_n52), .ZN(npu_inst_pe_1_7_1_n69) );
  OAI21_X1 npu_inst_pe_1_7_1_U76 ( .B1(npu_inst_pe_1_7_1_n61), .B2(
        npu_inst_pe_1_7_1_n52), .A(npu_inst_pe_1_7_1_n69), .ZN(
        npu_inst_pe_1_7_1_n92) );
  NAND2_X1 npu_inst_pe_1_7_1_U75 ( .A1(npu_inst_pe_1_7_1_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_7_1_n48), .ZN(npu_inst_pe_1_7_1_n68) );
  OAI21_X1 npu_inst_pe_1_7_1_U74 ( .B1(npu_inst_pe_1_7_1_n63), .B2(
        npu_inst_pe_1_7_1_n48), .A(npu_inst_pe_1_7_1_n68), .ZN(
        npu_inst_pe_1_7_1_n91) );
  NAND2_X1 npu_inst_pe_1_7_1_U73 ( .A1(npu_inst_pe_1_7_1_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_7_1_n48), .ZN(npu_inst_pe_1_7_1_n67) );
  OAI21_X1 npu_inst_pe_1_7_1_U72 ( .B1(npu_inst_pe_1_7_1_n61), .B2(
        npu_inst_pe_1_7_1_n48), .A(npu_inst_pe_1_7_1_n67), .ZN(
        npu_inst_pe_1_7_1_n90) );
  NAND2_X1 npu_inst_pe_1_7_1_U71 ( .A1(npu_inst_pe_1_7_1_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_7_1_n44), .ZN(npu_inst_pe_1_7_1_n66) );
  OAI21_X1 npu_inst_pe_1_7_1_U70 ( .B1(npu_inst_pe_1_7_1_n63), .B2(
        npu_inst_pe_1_7_1_n44), .A(npu_inst_pe_1_7_1_n66), .ZN(
        npu_inst_pe_1_7_1_n89) );
  NAND2_X1 npu_inst_pe_1_7_1_U69 ( .A1(npu_inst_pe_1_7_1_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_7_1_n44), .ZN(npu_inst_pe_1_7_1_n65) );
  OAI21_X1 npu_inst_pe_1_7_1_U68 ( .B1(npu_inst_pe_1_7_1_n61), .B2(
        npu_inst_pe_1_7_1_n44), .A(npu_inst_pe_1_7_1_n65), .ZN(
        npu_inst_pe_1_7_1_n88) );
  NAND2_X1 npu_inst_pe_1_7_1_U67 ( .A1(npu_inst_pe_1_7_1_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_7_1_n40), .ZN(npu_inst_pe_1_7_1_n64) );
  OAI21_X1 npu_inst_pe_1_7_1_U66 ( .B1(npu_inst_pe_1_7_1_n63), .B2(
        npu_inst_pe_1_7_1_n40), .A(npu_inst_pe_1_7_1_n64), .ZN(
        npu_inst_pe_1_7_1_n87) );
  NAND2_X1 npu_inst_pe_1_7_1_U65 ( .A1(npu_inst_pe_1_7_1_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_7_1_n40), .ZN(npu_inst_pe_1_7_1_n62) );
  OAI21_X1 npu_inst_pe_1_7_1_U64 ( .B1(npu_inst_pe_1_7_1_n61), .B2(
        npu_inst_pe_1_7_1_n40), .A(npu_inst_pe_1_7_1_n62), .ZN(
        npu_inst_pe_1_7_1_n86) );
  AND2_X1 npu_inst_pe_1_7_1_U63 ( .A1(npu_inst_pe_1_7_1_N93), .A2(npu_inst_n52), .ZN(npu_inst_int_data_y_7__1__0_) );
  AND2_X1 npu_inst_pe_1_7_1_U62 ( .A1(npu_inst_n52), .A2(npu_inst_pe_1_7_1_N94), .ZN(npu_inst_int_data_y_7__1__1_) );
  AOI22_X1 npu_inst_pe_1_7_1_U61 ( .A1(npu_inst_n52), .A2(int_i_data_v_npu[13]), .B1(npu_inst_pe_1_7_1_n3), .B2(npu_inst_int_data_x_7__2__1_), .ZN(
        npu_inst_pe_1_7_1_n63) );
  AOI22_X1 npu_inst_pe_1_7_1_U60 ( .A1(npu_inst_n52), .A2(int_i_data_v_npu[12]), .B1(npu_inst_pe_1_7_1_n3), .B2(npu_inst_int_data_x_7__2__0_), .ZN(
        npu_inst_pe_1_7_1_n61) );
  AOI222_X1 npu_inst_pe_1_7_1_U59 ( .A1(1'b0), .A2(npu_inst_pe_1_7_1_n1), .B1(
        npu_inst_pe_1_7_1_N73), .B2(npu_inst_pe_1_7_1_n76), .C1(
        npu_inst_pe_1_7_1_N65), .C2(npu_inst_pe_1_7_1_n77), .ZN(
        npu_inst_pe_1_7_1_n84) );
  INV_X1 npu_inst_pe_1_7_1_U58 ( .A(npu_inst_pe_1_7_1_n84), .ZN(
        npu_inst_pe_1_7_1_n101) );
  AOI222_X1 npu_inst_pe_1_7_1_U57 ( .A1(1'b0), .A2(npu_inst_pe_1_7_1_n1), .B1(
        npu_inst_pe_1_7_1_N80), .B2(npu_inst_pe_1_7_1_n76), .C1(
        npu_inst_pe_1_7_1_N72), .C2(npu_inst_pe_1_7_1_n77), .ZN(
        npu_inst_pe_1_7_1_n75) );
  INV_X1 npu_inst_pe_1_7_1_U56 ( .A(npu_inst_pe_1_7_1_n75), .ZN(
        npu_inst_pe_1_7_1_n33) );
  AOI222_X1 npu_inst_pe_1_7_1_U55 ( .A1(1'b0), .A2(npu_inst_pe_1_7_1_n1), .B1(
        npu_inst_pe_1_7_1_N74), .B2(npu_inst_pe_1_7_1_n76), .C1(
        npu_inst_pe_1_7_1_N66), .C2(npu_inst_pe_1_7_1_n77), .ZN(
        npu_inst_pe_1_7_1_n83) );
  INV_X1 npu_inst_pe_1_7_1_U54 ( .A(npu_inst_pe_1_7_1_n83), .ZN(
        npu_inst_pe_1_7_1_n100) );
  AOI222_X1 npu_inst_pe_1_7_1_U53 ( .A1(1'b0), .A2(npu_inst_pe_1_7_1_n1), .B1(
        npu_inst_pe_1_7_1_N75), .B2(npu_inst_pe_1_7_1_n76), .C1(
        npu_inst_pe_1_7_1_N67), .C2(npu_inst_pe_1_7_1_n77), .ZN(
        npu_inst_pe_1_7_1_n82) );
  INV_X1 npu_inst_pe_1_7_1_U52 ( .A(npu_inst_pe_1_7_1_n82), .ZN(
        npu_inst_pe_1_7_1_n99) );
  AOI222_X1 npu_inst_pe_1_7_1_U51 ( .A1(1'b0), .A2(npu_inst_pe_1_7_1_n1), .B1(
        npu_inst_pe_1_7_1_N76), .B2(npu_inst_pe_1_7_1_n76), .C1(
        npu_inst_pe_1_7_1_N68), .C2(npu_inst_pe_1_7_1_n77), .ZN(
        npu_inst_pe_1_7_1_n81) );
  INV_X1 npu_inst_pe_1_7_1_U50 ( .A(npu_inst_pe_1_7_1_n81), .ZN(
        npu_inst_pe_1_7_1_n98) );
  AOI222_X1 npu_inst_pe_1_7_1_U49 ( .A1(1'b0), .A2(npu_inst_pe_1_7_1_n1), .B1(
        npu_inst_pe_1_7_1_N77), .B2(npu_inst_pe_1_7_1_n76), .C1(
        npu_inst_pe_1_7_1_N69), .C2(npu_inst_pe_1_7_1_n77), .ZN(
        npu_inst_pe_1_7_1_n80) );
  INV_X1 npu_inst_pe_1_7_1_U48 ( .A(npu_inst_pe_1_7_1_n80), .ZN(
        npu_inst_pe_1_7_1_n36) );
  AOI222_X1 npu_inst_pe_1_7_1_U47 ( .A1(1'b0), .A2(npu_inst_pe_1_7_1_n1), .B1(
        npu_inst_pe_1_7_1_N78), .B2(npu_inst_pe_1_7_1_n76), .C1(
        npu_inst_pe_1_7_1_N70), .C2(npu_inst_pe_1_7_1_n77), .ZN(
        npu_inst_pe_1_7_1_n79) );
  INV_X1 npu_inst_pe_1_7_1_U46 ( .A(npu_inst_pe_1_7_1_n79), .ZN(
        npu_inst_pe_1_7_1_n35) );
  AOI222_X1 npu_inst_pe_1_7_1_U45 ( .A1(1'b0), .A2(npu_inst_pe_1_7_1_n1), .B1(
        npu_inst_pe_1_7_1_N79), .B2(npu_inst_pe_1_7_1_n76), .C1(
        npu_inst_pe_1_7_1_N71), .C2(npu_inst_pe_1_7_1_n77), .ZN(
        npu_inst_pe_1_7_1_n78) );
  INV_X1 npu_inst_pe_1_7_1_U44 ( .A(npu_inst_pe_1_7_1_n78), .ZN(
        npu_inst_pe_1_7_1_n34) );
  AND2_X1 npu_inst_pe_1_7_1_U43 ( .A1(npu_inst_pe_1_7_1_int_q_acc_0_), .A2(
        npu_inst_pe_1_7_1_n1), .ZN(npu_inst_int_data_res_7__1__0_) );
  AND2_X1 npu_inst_pe_1_7_1_U42 ( .A1(npu_inst_pe_1_7_1_n2), .A2(
        npu_inst_pe_1_7_1_int_q_acc_7_), .ZN(npu_inst_int_data_res_7__1__7_)
         );
  AND2_X1 npu_inst_pe_1_7_1_U41 ( .A1(npu_inst_pe_1_7_1_int_q_acc_1_), .A2(
        npu_inst_pe_1_7_1_n1), .ZN(npu_inst_int_data_res_7__1__1_) );
  AND2_X1 npu_inst_pe_1_7_1_U40 ( .A1(npu_inst_pe_1_7_1_int_q_acc_2_), .A2(
        npu_inst_pe_1_7_1_n1), .ZN(npu_inst_int_data_res_7__1__2_) );
  AND2_X1 npu_inst_pe_1_7_1_U39 ( .A1(npu_inst_pe_1_7_1_int_q_acc_3_), .A2(
        npu_inst_pe_1_7_1_n2), .ZN(npu_inst_int_data_res_7__1__3_) );
  AND2_X1 npu_inst_pe_1_7_1_U38 ( .A1(npu_inst_pe_1_7_1_int_q_acc_4_), .A2(
        npu_inst_pe_1_7_1_n2), .ZN(npu_inst_int_data_res_7__1__4_) );
  AND2_X1 npu_inst_pe_1_7_1_U37 ( .A1(npu_inst_pe_1_7_1_int_q_acc_5_), .A2(
        npu_inst_pe_1_7_1_n2), .ZN(npu_inst_int_data_res_7__1__5_) );
  AND2_X1 npu_inst_pe_1_7_1_U36 ( .A1(npu_inst_pe_1_7_1_int_q_acc_6_), .A2(
        npu_inst_pe_1_7_1_n2), .ZN(npu_inst_int_data_res_7__1__6_) );
  INV_X1 npu_inst_pe_1_7_1_U35 ( .A(npu_inst_pe_1_7_1_int_data_1_), .ZN(
        npu_inst_pe_1_7_1_n14) );
  NOR3_X1 npu_inst_pe_1_7_1_U34 ( .A1(npu_inst_pe_1_7_1_n26), .A2(npu_inst_n52), .A3(npu_inst_int_ckg[6]), .ZN(npu_inst_pe_1_7_1_n85) );
  OR2_X1 npu_inst_pe_1_7_1_U33 ( .A1(npu_inst_pe_1_7_1_n85), .A2(
        npu_inst_pe_1_7_1_n2), .ZN(npu_inst_pe_1_7_1_N84) );
  AND2_X1 npu_inst_pe_1_7_1_U32 ( .A1(npu_inst_int_data_x_7__1__1_), .A2(
        npu_inst_pe_1_7_1_int_q_weight_1_), .ZN(npu_inst_pe_1_7_1_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_7_1_U31 ( .A1(npu_inst_int_data_x_7__1__0_), .A2(
        npu_inst_pe_1_7_1_int_q_weight_1_), .ZN(npu_inst_pe_1_7_1_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_7_1_U30 ( .A(npu_inst_pe_1_7_1_int_data_0_), .ZN(
        npu_inst_pe_1_7_1_n13) );
  INV_X1 npu_inst_pe_1_7_1_U29 ( .A(npu_inst_n67), .ZN(npu_inst_pe_1_7_1_n5)
         );
  OR3_X1 npu_inst_pe_1_7_1_U28 ( .A1(npu_inst_pe_1_7_1_n6), .A2(
        npu_inst_pe_1_7_1_n8), .A3(npu_inst_pe_1_7_1_n5), .ZN(
        npu_inst_pe_1_7_1_n56) );
  OR3_X1 npu_inst_pe_1_7_1_U27 ( .A1(npu_inst_pe_1_7_1_n5), .A2(
        npu_inst_pe_1_7_1_n8), .A3(npu_inst_pe_1_7_1_n7), .ZN(
        npu_inst_pe_1_7_1_n48) );
  INV_X1 npu_inst_pe_1_7_1_U26 ( .A(npu_inst_pe_1_7_1_n5), .ZN(
        npu_inst_pe_1_7_1_n4) );
  OR3_X1 npu_inst_pe_1_7_1_U25 ( .A1(npu_inst_pe_1_7_1_n4), .A2(
        npu_inst_pe_1_7_1_n8), .A3(npu_inst_pe_1_7_1_n7), .ZN(
        npu_inst_pe_1_7_1_n52) );
  OR3_X1 npu_inst_pe_1_7_1_U24 ( .A1(npu_inst_pe_1_7_1_n6), .A2(
        npu_inst_pe_1_7_1_n8), .A3(npu_inst_pe_1_7_1_n4), .ZN(
        npu_inst_pe_1_7_1_n60) );
  NOR2_X1 npu_inst_pe_1_7_1_U23 ( .A1(npu_inst_pe_1_7_1_n60), .A2(
        npu_inst_pe_1_7_1_n3), .ZN(npu_inst_pe_1_7_1_n58) );
  NOR2_X1 npu_inst_pe_1_7_1_U22 ( .A1(npu_inst_pe_1_7_1_n56), .A2(
        npu_inst_pe_1_7_1_n3), .ZN(npu_inst_pe_1_7_1_n54) );
  NOR2_X1 npu_inst_pe_1_7_1_U21 ( .A1(npu_inst_pe_1_7_1_n52), .A2(
        npu_inst_pe_1_7_1_n3), .ZN(npu_inst_pe_1_7_1_n50) );
  NOR2_X1 npu_inst_pe_1_7_1_U20 ( .A1(npu_inst_pe_1_7_1_n48), .A2(
        npu_inst_pe_1_7_1_n3), .ZN(npu_inst_pe_1_7_1_n46) );
  NOR2_X1 npu_inst_pe_1_7_1_U19 ( .A1(npu_inst_pe_1_7_1_n40), .A2(
        npu_inst_pe_1_7_1_n3), .ZN(npu_inst_pe_1_7_1_n38) );
  NOR2_X1 npu_inst_pe_1_7_1_U18 ( .A1(npu_inst_pe_1_7_1_n44), .A2(
        npu_inst_pe_1_7_1_n3), .ZN(npu_inst_pe_1_7_1_n42) );
  BUF_X1 npu_inst_pe_1_7_1_U17 ( .A(npu_inst_n93), .Z(npu_inst_pe_1_7_1_n8) );
  INV_X1 npu_inst_pe_1_7_1_U16 ( .A(npu_inst_n122), .ZN(npu_inst_pe_1_7_1_n12)
         );
  INV_X1 npu_inst_pe_1_7_1_U15 ( .A(npu_inst_pe_1_7_1_n38), .ZN(
        npu_inst_pe_1_7_1_n114) );
  INV_X1 npu_inst_pe_1_7_1_U14 ( .A(npu_inst_pe_1_7_1_n58), .ZN(
        npu_inst_pe_1_7_1_n119) );
  INV_X1 npu_inst_pe_1_7_1_U13 ( .A(npu_inst_pe_1_7_1_n54), .ZN(
        npu_inst_pe_1_7_1_n118) );
  INV_X1 npu_inst_pe_1_7_1_U12 ( .A(npu_inst_pe_1_7_1_n50), .ZN(
        npu_inst_pe_1_7_1_n117) );
  INV_X1 npu_inst_pe_1_7_1_U11 ( .A(npu_inst_pe_1_7_1_n46), .ZN(
        npu_inst_pe_1_7_1_n116) );
  INV_X1 npu_inst_pe_1_7_1_U10 ( .A(npu_inst_pe_1_7_1_n42), .ZN(
        npu_inst_pe_1_7_1_n115) );
  BUF_X1 npu_inst_pe_1_7_1_U9 ( .A(npu_inst_n10), .Z(npu_inst_pe_1_7_1_n2) );
  BUF_X1 npu_inst_pe_1_7_1_U8 ( .A(npu_inst_n10), .Z(npu_inst_pe_1_7_1_n1) );
  BUF_X1 npu_inst_pe_1_7_1_U7 ( .A(npu_inst_pe_1_7_1_n12), .Z(
        npu_inst_pe_1_7_1_n11) );
  BUF_X1 npu_inst_pe_1_7_1_U6 ( .A(npu_inst_pe_1_7_1_n12), .Z(
        npu_inst_pe_1_7_1_n10) );
  BUF_X1 npu_inst_pe_1_7_1_U5 ( .A(npu_inst_pe_1_7_1_n12), .Z(
        npu_inst_pe_1_7_1_n9) );
  NOR2_X1 npu_inst_pe_1_7_1_U4 ( .A1(npu_inst_pe_1_7_1_int_q_weight_0_), .A2(
        npu_inst_pe_1_7_1_n1), .ZN(npu_inst_pe_1_7_1_n76) );
  NOR2_X1 npu_inst_pe_1_7_1_U3 ( .A1(npu_inst_pe_1_7_1_n27), .A2(
        npu_inst_pe_1_7_1_n1), .ZN(npu_inst_pe_1_7_1_n77) );
  FA_X1 npu_inst_pe_1_7_1_sub_67_U2_1 ( .A(npu_inst_pe_1_7_1_int_q_acc_1_), 
        .B(npu_inst_pe_1_7_1_n14), .CI(npu_inst_pe_1_7_1_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_7_1_sub_67_carry_2_), .S(npu_inst_pe_1_7_1_N66) );
  FA_X1 npu_inst_pe_1_7_1_add_69_U1_1 ( .A(npu_inst_pe_1_7_1_int_q_acc_1_), 
        .B(npu_inst_pe_1_7_1_int_data_1_), .CI(
        npu_inst_pe_1_7_1_add_69_carry_1_), .CO(
        npu_inst_pe_1_7_1_add_69_carry_2_), .S(npu_inst_pe_1_7_1_N74) );
  NAND3_X1 npu_inst_pe_1_7_1_U109 ( .A1(npu_inst_pe_1_7_1_n5), .A2(
        npu_inst_pe_1_7_1_n7), .A3(npu_inst_pe_1_7_1_n8), .ZN(
        npu_inst_pe_1_7_1_n44) );
  NAND3_X1 npu_inst_pe_1_7_1_U108 ( .A1(npu_inst_pe_1_7_1_n4), .A2(
        npu_inst_pe_1_7_1_n7), .A3(npu_inst_pe_1_7_1_n8), .ZN(
        npu_inst_pe_1_7_1_n40) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_7_1_n34), .CK(
        npu_inst_pe_1_7_1_net3251), .RN(npu_inst_pe_1_7_1_n9), .Q(
        npu_inst_pe_1_7_1_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_7_1_n35), .CK(
        npu_inst_pe_1_7_1_net3251), .RN(npu_inst_pe_1_7_1_n9), .Q(
        npu_inst_pe_1_7_1_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_7_1_n36), .CK(
        npu_inst_pe_1_7_1_net3251), .RN(npu_inst_pe_1_7_1_n9), .Q(
        npu_inst_pe_1_7_1_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_7_1_n98), .CK(
        npu_inst_pe_1_7_1_net3251), .RN(npu_inst_pe_1_7_1_n9), .Q(
        npu_inst_pe_1_7_1_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_7_1_n99), .CK(
        npu_inst_pe_1_7_1_net3251), .RN(npu_inst_pe_1_7_1_n9), .Q(
        npu_inst_pe_1_7_1_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_7_1_n100), 
        .CK(npu_inst_pe_1_7_1_net3251), .RN(npu_inst_pe_1_7_1_n9), .Q(
        npu_inst_pe_1_7_1_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_7_1_n33), .CK(
        npu_inst_pe_1_7_1_net3251), .RN(npu_inst_pe_1_7_1_n9), .Q(
        npu_inst_pe_1_7_1_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_7_1_n101), 
        .CK(npu_inst_pe_1_7_1_net3251), .RN(npu_inst_pe_1_7_1_n9), .Q(
        npu_inst_pe_1_7_1_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_weight_reg_0_ ( .D(npu_inst_n108), .CK(
        npu_inst_pe_1_7_1_net3257), .RN(npu_inst_pe_1_7_1_n9), .Q(
        npu_inst_pe_1_7_1_int_q_weight_0_), .QN(npu_inst_pe_1_7_1_n27) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_weight_reg_1_ ( .D(npu_inst_n114), .CK(
        npu_inst_pe_1_7_1_net3257), .RN(npu_inst_pe_1_7_1_n9), .Q(
        npu_inst_pe_1_7_1_int_q_weight_1_), .QN(npu_inst_pe_1_7_1_n26) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_7_1_n113), 
        .CK(npu_inst_pe_1_7_1_net3257), .RN(npu_inst_pe_1_7_1_n9), .Q(
        npu_inst_pe_1_7_1_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_7_1_n112), 
        .CK(npu_inst_pe_1_7_1_net3257), .RN(npu_inst_pe_1_7_1_n9), .Q(
        npu_inst_pe_1_7_1_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_7_1_n111), 
        .CK(npu_inst_pe_1_7_1_net3257), .RN(npu_inst_pe_1_7_1_n10), .Q(
        npu_inst_pe_1_7_1_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_7_1_n110), 
        .CK(npu_inst_pe_1_7_1_net3257), .RN(npu_inst_pe_1_7_1_n10), .Q(
        npu_inst_pe_1_7_1_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_7_1_n109), 
        .CK(npu_inst_pe_1_7_1_net3257), .RN(npu_inst_pe_1_7_1_n10), .Q(
        npu_inst_pe_1_7_1_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_7_1_n108), 
        .CK(npu_inst_pe_1_7_1_net3257), .RN(npu_inst_pe_1_7_1_n10), .Q(
        npu_inst_pe_1_7_1_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_7_1_n107), 
        .CK(npu_inst_pe_1_7_1_net3257), .RN(npu_inst_pe_1_7_1_n10), .Q(
        npu_inst_pe_1_7_1_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_7_1_n106), 
        .CK(npu_inst_pe_1_7_1_net3257), .RN(npu_inst_pe_1_7_1_n10), .Q(
        npu_inst_pe_1_7_1_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_7_1_n105), 
        .CK(npu_inst_pe_1_7_1_net3257), .RN(npu_inst_pe_1_7_1_n10), .Q(
        npu_inst_pe_1_7_1_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_7_1_n104), 
        .CK(npu_inst_pe_1_7_1_net3257), .RN(npu_inst_pe_1_7_1_n10), .Q(
        npu_inst_pe_1_7_1_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_7_1_n103), 
        .CK(npu_inst_pe_1_7_1_net3257), .RN(npu_inst_pe_1_7_1_n10), .Q(
        npu_inst_pe_1_7_1_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_7_1_n102), 
        .CK(npu_inst_pe_1_7_1_net3257), .RN(npu_inst_pe_1_7_1_n10), .Q(
        npu_inst_pe_1_7_1_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_7_1_n86), 
        .CK(npu_inst_pe_1_7_1_net3257), .RN(npu_inst_pe_1_7_1_n10), .Q(
        npu_inst_pe_1_7_1_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_7_1_n87), 
        .CK(npu_inst_pe_1_7_1_net3257), .RN(npu_inst_pe_1_7_1_n10), .Q(
        npu_inst_pe_1_7_1_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_7_1_n88), 
        .CK(npu_inst_pe_1_7_1_net3257), .RN(npu_inst_pe_1_7_1_n11), .Q(
        npu_inst_pe_1_7_1_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_7_1_n89), 
        .CK(npu_inst_pe_1_7_1_net3257), .RN(npu_inst_pe_1_7_1_n11), .Q(
        npu_inst_pe_1_7_1_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_7_1_n90), 
        .CK(npu_inst_pe_1_7_1_net3257), .RN(npu_inst_pe_1_7_1_n11), .Q(
        npu_inst_pe_1_7_1_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_7_1_n91), 
        .CK(npu_inst_pe_1_7_1_net3257), .RN(npu_inst_pe_1_7_1_n11), .Q(
        npu_inst_pe_1_7_1_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_7_1_n92), 
        .CK(npu_inst_pe_1_7_1_net3257), .RN(npu_inst_pe_1_7_1_n11), .Q(
        npu_inst_pe_1_7_1_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_7_1_n93), 
        .CK(npu_inst_pe_1_7_1_net3257), .RN(npu_inst_pe_1_7_1_n11), .Q(
        npu_inst_pe_1_7_1_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_7_1_n94), 
        .CK(npu_inst_pe_1_7_1_net3257), .RN(npu_inst_pe_1_7_1_n11), .Q(
        npu_inst_pe_1_7_1_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_7_1_n95), 
        .CK(npu_inst_pe_1_7_1_net3257), .RN(npu_inst_pe_1_7_1_n11), .Q(
        npu_inst_pe_1_7_1_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_7_1_n96), 
        .CK(npu_inst_pe_1_7_1_net3257), .RN(npu_inst_pe_1_7_1_n11), .Q(
        npu_inst_pe_1_7_1_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_7_1_n97), 
        .CK(npu_inst_pe_1_7_1_net3257), .RN(npu_inst_pe_1_7_1_n11), .Q(
        npu_inst_pe_1_7_1_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_7_1_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_7_1_N84), .SE(1'b0), .GCK(npu_inst_pe_1_7_1_net3251) );
  CLKGATETST_X1 npu_inst_pe_1_7_1_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n61), .SE(1'b0), .GCK(npu_inst_pe_1_7_1_net3257) );
  MUX2_X1 npu_inst_pe_1_7_2_U162 ( .A(npu_inst_pe_1_7_2_n32), .B(
        npu_inst_pe_1_7_2_n29), .S(npu_inst_pe_1_7_2_n8), .Z(
        npu_inst_pe_1_7_2_N93) );
  MUX2_X1 npu_inst_pe_1_7_2_U161 ( .A(npu_inst_pe_1_7_2_n31), .B(
        npu_inst_pe_1_7_2_n30), .S(npu_inst_pe_1_7_2_n6), .Z(
        npu_inst_pe_1_7_2_n32) );
  MUX2_X1 npu_inst_pe_1_7_2_U160 ( .A(npu_inst_pe_1_7_2_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_7_2_int_q_reg_v_1__0_), .S(npu_inst_pe_1_7_2_n4), .Z(
        npu_inst_pe_1_7_2_n31) );
  MUX2_X1 npu_inst_pe_1_7_2_U159 ( .A(npu_inst_pe_1_7_2_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_7_2_int_q_reg_v_3__0_), .S(npu_inst_pe_1_7_2_n4), .Z(
        npu_inst_pe_1_7_2_n30) );
  MUX2_X1 npu_inst_pe_1_7_2_U158 ( .A(npu_inst_pe_1_7_2_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_7_2_int_q_reg_v_5__0_), .S(npu_inst_pe_1_7_2_n4), .Z(
        npu_inst_pe_1_7_2_n29) );
  MUX2_X1 npu_inst_pe_1_7_2_U157 ( .A(npu_inst_pe_1_7_2_n28), .B(
        npu_inst_pe_1_7_2_n23), .S(npu_inst_pe_1_7_2_n8), .Z(
        npu_inst_pe_1_7_2_N94) );
  MUX2_X1 npu_inst_pe_1_7_2_U156 ( .A(npu_inst_pe_1_7_2_n25), .B(
        npu_inst_pe_1_7_2_n24), .S(npu_inst_pe_1_7_2_n6), .Z(
        npu_inst_pe_1_7_2_n28) );
  MUX2_X1 npu_inst_pe_1_7_2_U155 ( .A(npu_inst_pe_1_7_2_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_7_2_int_q_reg_v_1__1_), .S(npu_inst_pe_1_7_2_n4), .Z(
        npu_inst_pe_1_7_2_n25) );
  MUX2_X1 npu_inst_pe_1_7_2_U154 ( .A(npu_inst_pe_1_7_2_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_7_2_int_q_reg_v_3__1_), .S(npu_inst_pe_1_7_2_n4), .Z(
        npu_inst_pe_1_7_2_n24) );
  MUX2_X1 npu_inst_pe_1_7_2_U153 ( .A(npu_inst_pe_1_7_2_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_7_2_int_q_reg_v_5__1_), .S(npu_inst_pe_1_7_2_n4), .Z(
        npu_inst_pe_1_7_2_n23) );
  MUX2_X1 npu_inst_pe_1_7_2_U152 ( .A(npu_inst_pe_1_7_2_n22), .B(
        npu_inst_pe_1_7_2_n19), .S(npu_inst_pe_1_7_2_n8), .Z(
        npu_inst_int_data_x_7__2__1_) );
  MUX2_X1 npu_inst_pe_1_7_2_U151 ( .A(npu_inst_pe_1_7_2_n21), .B(
        npu_inst_pe_1_7_2_n20), .S(npu_inst_pe_1_7_2_n6), .Z(
        npu_inst_pe_1_7_2_n22) );
  MUX2_X1 npu_inst_pe_1_7_2_U150 ( .A(npu_inst_pe_1_7_2_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_7_2_int_q_reg_h_1__1_), .S(npu_inst_pe_1_7_2_n4), .Z(
        npu_inst_pe_1_7_2_n21) );
  MUX2_X1 npu_inst_pe_1_7_2_U149 ( .A(npu_inst_pe_1_7_2_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_7_2_int_q_reg_h_3__1_), .S(npu_inst_pe_1_7_2_n4), .Z(
        npu_inst_pe_1_7_2_n20) );
  MUX2_X1 npu_inst_pe_1_7_2_U148 ( .A(npu_inst_pe_1_7_2_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_7_2_int_q_reg_h_5__1_), .S(npu_inst_pe_1_7_2_n4), .Z(
        npu_inst_pe_1_7_2_n19) );
  MUX2_X1 npu_inst_pe_1_7_2_U147 ( .A(npu_inst_pe_1_7_2_n18), .B(
        npu_inst_pe_1_7_2_n15), .S(npu_inst_pe_1_7_2_n8), .Z(
        npu_inst_int_data_x_7__2__0_) );
  MUX2_X1 npu_inst_pe_1_7_2_U146 ( .A(npu_inst_pe_1_7_2_n17), .B(
        npu_inst_pe_1_7_2_n16), .S(npu_inst_pe_1_7_2_n6), .Z(
        npu_inst_pe_1_7_2_n18) );
  MUX2_X1 npu_inst_pe_1_7_2_U145 ( .A(npu_inst_pe_1_7_2_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_7_2_int_q_reg_h_1__0_), .S(npu_inst_pe_1_7_2_n4), .Z(
        npu_inst_pe_1_7_2_n17) );
  MUX2_X1 npu_inst_pe_1_7_2_U144 ( .A(npu_inst_pe_1_7_2_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_7_2_int_q_reg_h_3__0_), .S(npu_inst_pe_1_7_2_n4), .Z(
        npu_inst_pe_1_7_2_n16) );
  MUX2_X1 npu_inst_pe_1_7_2_U143 ( .A(npu_inst_pe_1_7_2_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_7_2_int_q_reg_h_5__0_), .S(npu_inst_pe_1_7_2_n4), .Z(
        npu_inst_pe_1_7_2_n15) );
  XOR2_X1 npu_inst_pe_1_7_2_U142 ( .A(npu_inst_pe_1_7_2_int_data_0_), .B(
        npu_inst_pe_1_7_2_int_q_acc_0_), .Z(npu_inst_pe_1_7_2_N73) );
  AND2_X1 npu_inst_pe_1_7_2_U141 ( .A1(npu_inst_pe_1_7_2_int_q_acc_0_), .A2(
        npu_inst_pe_1_7_2_int_data_0_), .ZN(npu_inst_pe_1_7_2_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_7_2_U140 ( .A(npu_inst_pe_1_7_2_int_q_acc_0_), .B(
        npu_inst_pe_1_7_2_n13), .ZN(npu_inst_pe_1_7_2_N65) );
  OR2_X1 npu_inst_pe_1_7_2_U139 ( .A1(npu_inst_pe_1_7_2_n13), .A2(
        npu_inst_pe_1_7_2_int_q_acc_0_), .ZN(npu_inst_pe_1_7_2_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_7_2_U138 ( .A(npu_inst_pe_1_7_2_int_q_acc_2_), .B(
        npu_inst_pe_1_7_2_add_69_carry_2_), .Z(npu_inst_pe_1_7_2_N75) );
  AND2_X1 npu_inst_pe_1_7_2_U137 ( .A1(npu_inst_pe_1_7_2_add_69_carry_2_), 
        .A2(npu_inst_pe_1_7_2_int_q_acc_2_), .ZN(
        npu_inst_pe_1_7_2_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_7_2_U136 ( .A(npu_inst_pe_1_7_2_int_q_acc_3_), .B(
        npu_inst_pe_1_7_2_add_69_carry_3_), .Z(npu_inst_pe_1_7_2_N76) );
  AND2_X1 npu_inst_pe_1_7_2_U135 ( .A1(npu_inst_pe_1_7_2_add_69_carry_3_), 
        .A2(npu_inst_pe_1_7_2_int_q_acc_3_), .ZN(
        npu_inst_pe_1_7_2_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_7_2_U134 ( .A(npu_inst_pe_1_7_2_int_q_acc_4_), .B(
        npu_inst_pe_1_7_2_add_69_carry_4_), .Z(npu_inst_pe_1_7_2_N77) );
  AND2_X1 npu_inst_pe_1_7_2_U133 ( .A1(npu_inst_pe_1_7_2_add_69_carry_4_), 
        .A2(npu_inst_pe_1_7_2_int_q_acc_4_), .ZN(
        npu_inst_pe_1_7_2_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_7_2_U132 ( .A(npu_inst_pe_1_7_2_int_q_acc_5_), .B(
        npu_inst_pe_1_7_2_add_69_carry_5_), .Z(npu_inst_pe_1_7_2_N78) );
  AND2_X1 npu_inst_pe_1_7_2_U131 ( .A1(npu_inst_pe_1_7_2_add_69_carry_5_), 
        .A2(npu_inst_pe_1_7_2_int_q_acc_5_), .ZN(
        npu_inst_pe_1_7_2_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_7_2_U130 ( .A(npu_inst_pe_1_7_2_int_q_acc_6_), .B(
        npu_inst_pe_1_7_2_add_69_carry_6_), .Z(npu_inst_pe_1_7_2_N79) );
  AND2_X1 npu_inst_pe_1_7_2_U129 ( .A1(npu_inst_pe_1_7_2_add_69_carry_6_), 
        .A2(npu_inst_pe_1_7_2_int_q_acc_6_), .ZN(
        npu_inst_pe_1_7_2_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_7_2_U128 ( .A(npu_inst_pe_1_7_2_int_q_acc_7_), .B(
        npu_inst_pe_1_7_2_add_69_carry_7_), .Z(npu_inst_pe_1_7_2_N80) );
  XNOR2_X1 npu_inst_pe_1_7_2_U127 ( .A(npu_inst_pe_1_7_2_sub_67_carry_2_), .B(
        npu_inst_pe_1_7_2_int_q_acc_2_), .ZN(npu_inst_pe_1_7_2_N67) );
  OR2_X1 npu_inst_pe_1_7_2_U126 ( .A1(npu_inst_pe_1_7_2_int_q_acc_2_), .A2(
        npu_inst_pe_1_7_2_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_7_2_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_7_2_U125 ( .A(npu_inst_pe_1_7_2_sub_67_carry_3_), .B(
        npu_inst_pe_1_7_2_int_q_acc_3_), .ZN(npu_inst_pe_1_7_2_N68) );
  OR2_X1 npu_inst_pe_1_7_2_U124 ( .A1(npu_inst_pe_1_7_2_int_q_acc_3_), .A2(
        npu_inst_pe_1_7_2_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_7_2_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_7_2_U123 ( .A(npu_inst_pe_1_7_2_sub_67_carry_4_), .B(
        npu_inst_pe_1_7_2_int_q_acc_4_), .ZN(npu_inst_pe_1_7_2_N69) );
  OR2_X1 npu_inst_pe_1_7_2_U122 ( .A1(npu_inst_pe_1_7_2_int_q_acc_4_), .A2(
        npu_inst_pe_1_7_2_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_7_2_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_7_2_U121 ( .A(npu_inst_pe_1_7_2_sub_67_carry_5_), .B(
        npu_inst_pe_1_7_2_int_q_acc_5_), .ZN(npu_inst_pe_1_7_2_N70) );
  OR2_X1 npu_inst_pe_1_7_2_U120 ( .A1(npu_inst_pe_1_7_2_int_q_acc_5_), .A2(
        npu_inst_pe_1_7_2_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_7_2_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_7_2_U119 ( .A(npu_inst_pe_1_7_2_sub_67_carry_6_), .B(
        npu_inst_pe_1_7_2_int_q_acc_6_), .ZN(npu_inst_pe_1_7_2_N71) );
  OR2_X1 npu_inst_pe_1_7_2_U118 ( .A1(npu_inst_pe_1_7_2_int_q_acc_6_), .A2(
        npu_inst_pe_1_7_2_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_7_2_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_7_2_U117 ( .A(npu_inst_pe_1_7_2_int_q_acc_7_), .B(
        npu_inst_pe_1_7_2_sub_67_carry_7_), .ZN(npu_inst_pe_1_7_2_N72) );
  INV_X1 npu_inst_pe_1_7_2_U116 ( .A(npu_inst_n75), .ZN(npu_inst_pe_1_7_2_n7)
         );
  INV_X1 npu_inst_pe_1_7_2_U115 ( .A(npu_inst_pe_1_7_2_n7), .ZN(
        npu_inst_pe_1_7_2_n6) );
  INV_X1 npu_inst_pe_1_7_2_U114 ( .A(npu_inst_n52), .ZN(npu_inst_pe_1_7_2_n3)
         );
  AOI22_X1 npu_inst_pe_1_7_2_U113 ( .A1(npu_inst_pe_1_7_2_n38), .A2(
        int_i_data_v_npu[11]), .B1(npu_inst_pe_1_7_2_n114), .B2(
        npu_inst_pe_1_7_2_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_7_2_n39) );
  INV_X1 npu_inst_pe_1_7_2_U112 ( .A(npu_inst_pe_1_7_2_n39), .ZN(
        npu_inst_pe_1_7_2_n112) );
  AOI22_X1 npu_inst_pe_1_7_2_U111 ( .A1(npu_inst_pe_1_7_2_n38), .A2(
        int_i_data_v_npu[10]), .B1(npu_inst_pe_1_7_2_n114), .B2(
        npu_inst_pe_1_7_2_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_7_2_n37) );
  INV_X1 npu_inst_pe_1_7_2_U110 ( .A(npu_inst_pe_1_7_2_n37), .ZN(
        npu_inst_pe_1_7_2_n113) );
  AOI22_X1 npu_inst_pe_1_7_2_U107 ( .A1(int_i_data_v_npu[11]), .A2(
        npu_inst_pe_1_7_2_n58), .B1(npu_inst_pe_1_7_2_n119), .B2(
        npu_inst_pe_1_7_2_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_7_2_n59) );
  INV_X1 npu_inst_pe_1_7_2_U106 ( .A(npu_inst_pe_1_7_2_n59), .ZN(
        npu_inst_pe_1_7_2_n102) );
  AOI22_X1 npu_inst_pe_1_7_2_U105 ( .A1(int_i_data_v_npu[10]), .A2(
        npu_inst_pe_1_7_2_n58), .B1(npu_inst_pe_1_7_2_n119), .B2(
        npu_inst_pe_1_7_2_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_7_2_n57) );
  INV_X1 npu_inst_pe_1_7_2_U104 ( .A(npu_inst_pe_1_7_2_n57), .ZN(
        npu_inst_pe_1_7_2_n103) );
  AOI22_X1 npu_inst_pe_1_7_2_U103 ( .A1(int_i_data_v_npu[11]), .A2(
        npu_inst_pe_1_7_2_n54), .B1(npu_inst_pe_1_7_2_n118), .B2(
        npu_inst_pe_1_7_2_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_7_2_n55) );
  INV_X1 npu_inst_pe_1_7_2_U102 ( .A(npu_inst_pe_1_7_2_n55), .ZN(
        npu_inst_pe_1_7_2_n104) );
  AOI22_X1 npu_inst_pe_1_7_2_U101 ( .A1(int_i_data_v_npu[10]), .A2(
        npu_inst_pe_1_7_2_n54), .B1(npu_inst_pe_1_7_2_n118), .B2(
        npu_inst_pe_1_7_2_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_7_2_n53) );
  INV_X1 npu_inst_pe_1_7_2_U100 ( .A(npu_inst_pe_1_7_2_n53), .ZN(
        npu_inst_pe_1_7_2_n105) );
  AOI22_X1 npu_inst_pe_1_7_2_U99 ( .A1(int_i_data_v_npu[11]), .A2(
        npu_inst_pe_1_7_2_n50), .B1(npu_inst_pe_1_7_2_n117), .B2(
        npu_inst_pe_1_7_2_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_7_2_n51) );
  INV_X1 npu_inst_pe_1_7_2_U98 ( .A(npu_inst_pe_1_7_2_n51), .ZN(
        npu_inst_pe_1_7_2_n106) );
  AOI22_X1 npu_inst_pe_1_7_2_U97 ( .A1(int_i_data_v_npu[10]), .A2(
        npu_inst_pe_1_7_2_n50), .B1(npu_inst_pe_1_7_2_n117), .B2(
        npu_inst_pe_1_7_2_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_7_2_n49) );
  INV_X1 npu_inst_pe_1_7_2_U96 ( .A(npu_inst_pe_1_7_2_n49), .ZN(
        npu_inst_pe_1_7_2_n107) );
  AOI22_X1 npu_inst_pe_1_7_2_U95 ( .A1(int_i_data_v_npu[11]), .A2(
        npu_inst_pe_1_7_2_n46), .B1(npu_inst_pe_1_7_2_n116), .B2(
        npu_inst_pe_1_7_2_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_7_2_n47) );
  INV_X1 npu_inst_pe_1_7_2_U94 ( .A(npu_inst_pe_1_7_2_n47), .ZN(
        npu_inst_pe_1_7_2_n108) );
  AOI22_X1 npu_inst_pe_1_7_2_U93 ( .A1(int_i_data_v_npu[10]), .A2(
        npu_inst_pe_1_7_2_n46), .B1(npu_inst_pe_1_7_2_n116), .B2(
        npu_inst_pe_1_7_2_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_7_2_n45) );
  INV_X1 npu_inst_pe_1_7_2_U92 ( .A(npu_inst_pe_1_7_2_n45), .ZN(
        npu_inst_pe_1_7_2_n109) );
  AOI22_X1 npu_inst_pe_1_7_2_U91 ( .A1(int_i_data_v_npu[11]), .A2(
        npu_inst_pe_1_7_2_n42), .B1(npu_inst_pe_1_7_2_n115), .B2(
        npu_inst_pe_1_7_2_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_7_2_n43) );
  INV_X1 npu_inst_pe_1_7_2_U90 ( .A(npu_inst_pe_1_7_2_n43), .ZN(
        npu_inst_pe_1_7_2_n110) );
  AOI22_X1 npu_inst_pe_1_7_2_U89 ( .A1(int_i_data_v_npu[10]), .A2(
        npu_inst_pe_1_7_2_n42), .B1(npu_inst_pe_1_7_2_n115), .B2(
        npu_inst_pe_1_7_2_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_7_2_n41) );
  INV_X1 npu_inst_pe_1_7_2_U88 ( .A(npu_inst_pe_1_7_2_n41), .ZN(
        npu_inst_pe_1_7_2_n111) );
  NAND2_X1 npu_inst_pe_1_7_2_U87 ( .A1(npu_inst_pe_1_7_2_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_7_2_n60), .ZN(npu_inst_pe_1_7_2_n74) );
  OAI21_X1 npu_inst_pe_1_7_2_U86 ( .B1(npu_inst_pe_1_7_2_n63), .B2(
        npu_inst_pe_1_7_2_n60), .A(npu_inst_pe_1_7_2_n74), .ZN(
        npu_inst_pe_1_7_2_n97) );
  NAND2_X1 npu_inst_pe_1_7_2_U85 ( .A1(npu_inst_pe_1_7_2_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_7_2_n60), .ZN(npu_inst_pe_1_7_2_n73) );
  OAI21_X1 npu_inst_pe_1_7_2_U84 ( .B1(npu_inst_pe_1_7_2_n61), .B2(
        npu_inst_pe_1_7_2_n60), .A(npu_inst_pe_1_7_2_n73), .ZN(
        npu_inst_pe_1_7_2_n96) );
  NAND2_X1 npu_inst_pe_1_7_2_U83 ( .A1(npu_inst_pe_1_7_2_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_7_2_n56), .ZN(npu_inst_pe_1_7_2_n72) );
  OAI21_X1 npu_inst_pe_1_7_2_U82 ( .B1(npu_inst_pe_1_7_2_n63), .B2(
        npu_inst_pe_1_7_2_n56), .A(npu_inst_pe_1_7_2_n72), .ZN(
        npu_inst_pe_1_7_2_n95) );
  NAND2_X1 npu_inst_pe_1_7_2_U81 ( .A1(npu_inst_pe_1_7_2_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_7_2_n56), .ZN(npu_inst_pe_1_7_2_n71) );
  OAI21_X1 npu_inst_pe_1_7_2_U80 ( .B1(npu_inst_pe_1_7_2_n61), .B2(
        npu_inst_pe_1_7_2_n56), .A(npu_inst_pe_1_7_2_n71), .ZN(
        npu_inst_pe_1_7_2_n94) );
  NAND2_X1 npu_inst_pe_1_7_2_U79 ( .A1(npu_inst_pe_1_7_2_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_7_2_n52), .ZN(npu_inst_pe_1_7_2_n70) );
  OAI21_X1 npu_inst_pe_1_7_2_U78 ( .B1(npu_inst_pe_1_7_2_n63), .B2(
        npu_inst_pe_1_7_2_n52), .A(npu_inst_pe_1_7_2_n70), .ZN(
        npu_inst_pe_1_7_2_n93) );
  NAND2_X1 npu_inst_pe_1_7_2_U77 ( .A1(npu_inst_pe_1_7_2_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_7_2_n52), .ZN(npu_inst_pe_1_7_2_n69) );
  OAI21_X1 npu_inst_pe_1_7_2_U76 ( .B1(npu_inst_pe_1_7_2_n61), .B2(
        npu_inst_pe_1_7_2_n52), .A(npu_inst_pe_1_7_2_n69), .ZN(
        npu_inst_pe_1_7_2_n92) );
  NAND2_X1 npu_inst_pe_1_7_2_U75 ( .A1(npu_inst_pe_1_7_2_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_7_2_n48), .ZN(npu_inst_pe_1_7_2_n68) );
  OAI21_X1 npu_inst_pe_1_7_2_U74 ( .B1(npu_inst_pe_1_7_2_n63), .B2(
        npu_inst_pe_1_7_2_n48), .A(npu_inst_pe_1_7_2_n68), .ZN(
        npu_inst_pe_1_7_2_n91) );
  NAND2_X1 npu_inst_pe_1_7_2_U73 ( .A1(npu_inst_pe_1_7_2_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_7_2_n48), .ZN(npu_inst_pe_1_7_2_n67) );
  OAI21_X1 npu_inst_pe_1_7_2_U72 ( .B1(npu_inst_pe_1_7_2_n61), .B2(
        npu_inst_pe_1_7_2_n48), .A(npu_inst_pe_1_7_2_n67), .ZN(
        npu_inst_pe_1_7_2_n90) );
  NAND2_X1 npu_inst_pe_1_7_2_U71 ( .A1(npu_inst_pe_1_7_2_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_7_2_n44), .ZN(npu_inst_pe_1_7_2_n66) );
  OAI21_X1 npu_inst_pe_1_7_2_U70 ( .B1(npu_inst_pe_1_7_2_n63), .B2(
        npu_inst_pe_1_7_2_n44), .A(npu_inst_pe_1_7_2_n66), .ZN(
        npu_inst_pe_1_7_2_n89) );
  NAND2_X1 npu_inst_pe_1_7_2_U69 ( .A1(npu_inst_pe_1_7_2_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_7_2_n44), .ZN(npu_inst_pe_1_7_2_n65) );
  OAI21_X1 npu_inst_pe_1_7_2_U68 ( .B1(npu_inst_pe_1_7_2_n61), .B2(
        npu_inst_pe_1_7_2_n44), .A(npu_inst_pe_1_7_2_n65), .ZN(
        npu_inst_pe_1_7_2_n88) );
  NAND2_X1 npu_inst_pe_1_7_2_U67 ( .A1(npu_inst_pe_1_7_2_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_7_2_n40), .ZN(npu_inst_pe_1_7_2_n64) );
  OAI21_X1 npu_inst_pe_1_7_2_U66 ( .B1(npu_inst_pe_1_7_2_n63), .B2(
        npu_inst_pe_1_7_2_n40), .A(npu_inst_pe_1_7_2_n64), .ZN(
        npu_inst_pe_1_7_2_n87) );
  NAND2_X1 npu_inst_pe_1_7_2_U65 ( .A1(npu_inst_pe_1_7_2_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_7_2_n40), .ZN(npu_inst_pe_1_7_2_n62) );
  OAI21_X1 npu_inst_pe_1_7_2_U64 ( .B1(npu_inst_pe_1_7_2_n61), .B2(
        npu_inst_pe_1_7_2_n40), .A(npu_inst_pe_1_7_2_n62), .ZN(
        npu_inst_pe_1_7_2_n86) );
  AND2_X1 npu_inst_pe_1_7_2_U63 ( .A1(npu_inst_pe_1_7_2_N93), .A2(npu_inst_n52), .ZN(npu_inst_int_data_y_7__2__0_) );
  AND2_X1 npu_inst_pe_1_7_2_U62 ( .A1(npu_inst_n52), .A2(npu_inst_pe_1_7_2_N94), .ZN(npu_inst_int_data_y_7__2__1_) );
  AOI22_X1 npu_inst_pe_1_7_2_U61 ( .A1(npu_inst_n52), .A2(int_i_data_v_npu[11]), .B1(npu_inst_pe_1_7_2_n3), .B2(npu_inst_int_data_x_7__3__1_), .ZN(
        npu_inst_pe_1_7_2_n63) );
  AOI22_X1 npu_inst_pe_1_7_2_U60 ( .A1(npu_inst_n52), .A2(int_i_data_v_npu[10]), .B1(npu_inst_pe_1_7_2_n3), .B2(npu_inst_int_data_x_7__3__0_), .ZN(
        npu_inst_pe_1_7_2_n61) );
  AOI222_X1 npu_inst_pe_1_7_2_U59 ( .A1(1'b0), .A2(npu_inst_pe_1_7_2_n1), .B1(
        npu_inst_pe_1_7_2_N73), .B2(npu_inst_pe_1_7_2_n76), .C1(
        npu_inst_pe_1_7_2_N65), .C2(npu_inst_pe_1_7_2_n77), .ZN(
        npu_inst_pe_1_7_2_n84) );
  INV_X1 npu_inst_pe_1_7_2_U58 ( .A(npu_inst_pe_1_7_2_n84), .ZN(
        npu_inst_pe_1_7_2_n101) );
  AOI222_X1 npu_inst_pe_1_7_2_U57 ( .A1(1'b0), .A2(npu_inst_pe_1_7_2_n1), .B1(
        npu_inst_pe_1_7_2_N80), .B2(npu_inst_pe_1_7_2_n76), .C1(
        npu_inst_pe_1_7_2_N72), .C2(npu_inst_pe_1_7_2_n77), .ZN(
        npu_inst_pe_1_7_2_n75) );
  INV_X1 npu_inst_pe_1_7_2_U56 ( .A(npu_inst_pe_1_7_2_n75), .ZN(
        npu_inst_pe_1_7_2_n33) );
  AOI222_X1 npu_inst_pe_1_7_2_U55 ( .A1(1'b0), .A2(npu_inst_pe_1_7_2_n1), .B1(
        npu_inst_pe_1_7_2_N74), .B2(npu_inst_pe_1_7_2_n76), .C1(
        npu_inst_pe_1_7_2_N66), .C2(npu_inst_pe_1_7_2_n77), .ZN(
        npu_inst_pe_1_7_2_n83) );
  INV_X1 npu_inst_pe_1_7_2_U54 ( .A(npu_inst_pe_1_7_2_n83), .ZN(
        npu_inst_pe_1_7_2_n100) );
  AOI222_X1 npu_inst_pe_1_7_2_U53 ( .A1(1'b0), .A2(npu_inst_pe_1_7_2_n1), .B1(
        npu_inst_pe_1_7_2_N75), .B2(npu_inst_pe_1_7_2_n76), .C1(
        npu_inst_pe_1_7_2_N67), .C2(npu_inst_pe_1_7_2_n77), .ZN(
        npu_inst_pe_1_7_2_n82) );
  INV_X1 npu_inst_pe_1_7_2_U52 ( .A(npu_inst_pe_1_7_2_n82), .ZN(
        npu_inst_pe_1_7_2_n99) );
  AOI222_X1 npu_inst_pe_1_7_2_U51 ( .A1(1'b0), .A2(npu_inst_pe_1_7_2_n1), .B1(
        npu_inst_pe_1_7_2_N76), .B2(npu_inst_pe_1_7_2_n76), .C1(
        npu_inst_pe_1_7_2_N68), .C2(npu_inst_pe_1_7_2_n77), .ZN(
        npu_inst_pe_1_7_2_n81) );
  INV_X1 npu_inst_pe_1_7_2_U50 ( .A(npu_inst_pe_1_7_2_n81), .ZN(
        npu_inst_pe_1_7_2_n98) );
  AOI222_X1 npu_inst_pe_1_7_2_U49 ( .A1(1'b0), .A2(npu_inst_pe_1_7_2_n1), .B1(
        npu_inst_pe_1_7_2_N77), .B2(npu_inst_pe_1_7_2_n76), .C1(
        npu_inst_pe_1_7_2_N69), .C2(npu_inst_pe_1_7_2_n77), .ZN(
        npu_inst_pe_1_7_2_n80) );
  INV_X1 npu_inst_pe_1_7_2_U48 ( .A(npu_inst_pe_1_7_2_n80), .ZN(
        npu_inst_pe_1_7_2_n36) );
  AOI222_X1 npu_inst_pe_1_7_2_U47 ( .A1(1'b0), .A2(npu_inst_pe_1_7_2_n1), .B1(
        npu_inst_pe_1_7_2_N78), .B2(npu_inst_pe_1_7_2_n76), .C1(
        npu_inst_pe_1_7_2_N70), .C2(npu_inst_pe_1_7_2_n77), .ZN(
        npu_inst_pe_1_7_2_n79) );
  INV_X1 npu_inst_pe_1_7_2_U46 ( .A(npu_inst_pe_1_7_2_n79), .ZN(
        npu_inst_pe_1_7_2_n35) );
  AOI222_X1 npu_inst_pe_1_7_2_U45 ( .A1(1'b0), .A2(npu_inst_pe_1_7_2_n1), .B1(
        npu_inst_pe_1_7_2_N79), .B2(npu_inst_pe_1_7_2_n76), .C1(
        npu_inst_pe_1_7_2_N71), .C2(npu_inst_pe_1_7_2_n77), .ZN(
        npu_inst_pe_1_7_2_n78) );
  INV_X1 npu_inst_pe_1_7_2_U44 ( .A(npu_inst_pe_1_7_2_n78), .ZN(
        npu_inst_pe_1_7_2_n34) );
  AND2_X1 npu_inst_pe_1_7_2_U43 ( .A1(npu_inst_pe_1_7_2_int_q_acc_0_), .A2(
        npu_inst_pe_1_7_2_n1), .ZN(npu_inst_int_data_res_7__2__0_) );
  AND2_X1 npu_inst_pe_1_7_2_U42 ( .A1(npu_inst_pe_1_7_2_n2), .A2(
        npu_inst_pe_1_7_2_int_q_acc_7_), .ZN(npu_inst_int_data_res_7__2__7_)
         );
  AND2_X1 npu_inst_pe_1_7_2_U41 ( .A1(npu_inst_pe_1_7_2_int_q_acc_1_), .A2(
        npu_inst_pe_1_7_2_n1), .ZN(npu_inst_int_data_res_7__2__1_) );
  AND2_X1 npu_inst_pe_1_7_2_U40 ( .A1(npu_inst_pe_1_7_2_int_q_acc_2_), .A2(
        npu_inst_pe_1_7_2_n1), .ZN(npu_inst_int_data_res_7__2__2_) );
  AND2_X1 npu_inst_pe_1_7_2_U39 ( .A1(npu_inst_pe_1_7_2_int_q_acc_3_), .A2(
        npu_inst_pe_1_7_2_n2), .ZN(npu_inst_int_data_res_7__2__3_) );
  AND2_X1 npu_inst_pe_1_7_2_U38 ( .A1(npu_inst_pe_1_7_2_int_q_acc_4_), .A2(
        npu_inst_pe_1_7_2_n2), .ZN(npu_inst_int_data_res_7__2__4_) );
  AND2_X1 npu_inst_pe_1_7_2_U37 ( .A1(npu_inst_pe_1_7_2_int_q_acc_5_), .A2(
        npu_inst_pe_1_7_2_n2), .ZN(npu_inst_int_data_res_7__2__5_) );
  AND2_X1 npu_inst_pe_1_7_2_U36 ( .A1(npu_inst_pe_1_7_2_int_q_acc_6_), .A2(
        npu_inst_pe_1_7_2_n2), .ZN(npu_inst_int_data_res_7__2__6_) );
  INV_X1 npu_inst_pe_1_7_2_U35 ( .A(npu_inst_pe_1_7_2_int_data_1_), .ZN(
        npu_inst_pe_1_7_2_n14) );
  NOR3_X1 npu_inst_pe_1_7_2_U34 ( .A1(npu_inst_pe_1_7_2_n26), .A2(npu_inst_n52), .A3(npu_inst_int_ckg[5]), .ZN(npu_inst_pe_1_7_2_n85) );
  OR2_X1 npu_inst_pe_1_7_2_U33 ( .A1(npu_inst_pe_1_7_2_n85), .A2(
        npu_inst_pe_1_7_2_n2), .ZN(npu_inst_pe_1_7_2_N84) );
  AND2_X1 npu_inst_pe_1_7_2_U32 ( .A1(npu_inst_int_data_x_7__2__1_), .A2(
        npu_inst_pe_1_7_2_int_q_weight_1_), .ZN(npu_inst_pe_1_7_2_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_7_2_U31 ( .A1(npu_inst_int_data_x_7__2__0_), .A2(
        npu_inst_pe_1_7_2_int_q_weight_1_), .ZN(npu_inst_pe_1_7_2_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_7_2_U30 ( .A(npu_inst_pe_1_7_2_int_data_0_), .ZN(
        npu_inst_pe_1_7_2_n13) );
  INV_X1 npu_inst_pe_1_7_2_U29 ( .A(npu_inst_n67), .ZN(npu_inst_pe_1_7_2_n5)
         );
  OR3_X1 npu_inst_pe_1_7_2_U28 ( .A1(npu_inst_pe_1_7_2_n6), .A2(
        npu_inst_pe_1_7_2_n8), .A3(npu_inst_pe_1_7_2_n5), .ZN(
        npu_inst_pe_1_7_2_n56) );
  OR3_X1 npu_inst_pe_1_7_2_U27 ( .A1(npu_inst_pe_1_7_2_n5), .A2(
        npu_inst_pe_1_7_2_n8), .A3(npu_inst_pe_1_7_2_n7), .ZN(
        npu_inst_pe_1_7_2_n48) );
  INV_X1 npu_inst_pe_1_7_2_U26 ( .A(npu_inst_pe_1_7_2_n5), .ZN(
        npu_inst_pe_1_7_2_n4) );
  OR3_X1 npu_inst_pe_1_7_2_U25 ( .A1(npu_inst_pe_1_7_2_n4), .A2(
        npu_inst_pe_1_7_2_n8), .A3(npu_inst_pe_1_7_2_n7), .ZN(
        npu_inst_pe_1_7_2_n52) );
  OR3_X1 npu_inst_pe_1_7_2_U24 ( .A1(npu_inst_pe_1_7_2_n6), .A2(
        npu_inst_pe_1_7_2_n8), .A3(npu_inst_pe_1_7_2_n4), .ZN(
        npu_inst_pe_1_7_2_n60) );
  NOR2_X1 npu_inst_pe_1_7_2_U23 ( .A1(npu_inst_pe_1_7_2_n60), .A2(
        npu_inst_pe_1_7_2_n3), .ZN(npu_inst_pe_1_7_2_n58) );
  NOR2_X1 npu_inst_pe_1_7_2_U22 ( .A1(npu_inst_pe_1_7_2_n56), .A2(
        npu_inst_pe_1_7_2_n3), .ZN(npu_inst_pe_1_7_2_n54) );
  NOR2_X1 npu_inst_pe_1_7_2_U21 ( .A1(npu_inst_pe_1_7_2_n52), .A2(
        npu_inst_pe_1_7_2_n3), .ZN(npu_inst_pe_1_7_2_n50) );
  NOR2_X1 npu_inst_pe_1_7_2_U20 ( .A1(npu_inst_pe_1_7_2_n48), .A2(
        npu_inst_pe_1_7_2_n3), .ZN(npu_inst_pe_1_7_2_n46) );
  NOR2_X1 npu_inst_pe_1_7_2_U19 ( .A1(npu_inst_pe_1_7_2_n40), .A2(
        npu_inst_pe_1_7_2_n3), .ZN(npu_inst_pe_1_7_2_n38) );
  NOR2_X1 npu_inst_pe_1_7_2_U18 ( .A1(npu_inst_pe_1_7_2_n44), .A2(
        npu_inst_pe_1_7_2_n3), .ZN(npu_inst_pe_1_7_2_n42) );
  BUF_X1 npu_inst_pe_1_7_2_U17 ( .A(npu_inst_n93), .Z(npu_inst_pe_1_7_2_n8) );
  INV_X1 npu_inst_pe_1_7_2_U16 ( .A(npu_inst_n122), .ZN(npu_inst_pe_1_7_2_n12)
         );
  INV_X1 npu_inst_pe_1_7_2_U15 ( .A(npu_inst_pe_1_7_2_n38), .ZN(
        npu_inst_pe_1_7_2_n114) );
  INV_X1 npu_inst_pe_1_7_2_U14 ( .A(npu_inst_pe_1_7_2_n58), .ZN(
        npu_inst_pe_1_7_2_n119) );
  INV_X1 npu_inst_pe_1_7_2_U13 ( .A(npu_inst_pe_1_7_2_n54), .ZN(
        npu_inst_pe_1_7_2_n118) );
  INV_X1 npu_inst_pe_1_7_2_U12 ( .A(npu_inst_pe_1_7_2_n50), .ZN(
        npu_inst_pe_1_7_2_n117) );
  INV_X1 npu_inst_pe_1_7_2_U11 ( .A(npu_inst_pe_1_7_2_n46), .ZN(
        npu_inst_pe_1_7_2_n116) );
  INV_X1 npu_inst_pe_1_7_2_U10 ( .A(npu_inst_pe_1_7_2_n42), .ZN(
        npu_inst_pe_1_7_2_n115) );
  BUF_X1 npu_inst_pe_1_7_2_U9 ( .A(npu_inst_n9), .Z(npu_inst_pe_1_7_2_n2) );
  BUF_X1 npu_inst_pe_1_7_2_U8 ( .A(npu_inst_n9), .Z(npu_inst_pe_1_7_2_n1) );
  BUF_X1 npu_inst_pe_1_7_2_U7 ( .A(npu_inst_pe_1_7_2_n12), .Z(
        npu_inst_pe_1_7_2_n11) );
  BUF_X1 npu_inst_pe_1_7_2_U6 ( .A(npu_inst_pe_1_7_2_n12), .Z(
        npu_inst_pe_1_7_2_n10) );
  BUF_X1 npu_inst_pe_1_7_2_U5 ( .A(npu_inst_pe_1_7_2_n12), .Z(
        npu_inst_pe_1_7_2_n9) );
  NOR2_X1 npu_inst_pe_1_7_2_U4 ( .A1(npu_inst_pe_1_7_2_int_q_weight_0_), .A2(
        npu_inst_pe_1_7_2_n1), .ZN(npu_inst_pe_1_7_2_n76) );
  NOR2_X1 npu_inst_pe_1_7_2_U3 ( .A1(npu_inst_pe_1_7_2_n27), .A2(
        npu_inst_pe_1_7_2_n1), .ZN(npu_inst_pe_1_7_2_n77) );
  FA_X1 npu_inst_pe_1_7_2_sub_67_U2_1 ( .A(npu_inst_pe_1_7_2_int_q_acc_1_), 
        .B(npu_inst_pe_1_7_2_n14), .CI(npu_inst_pe_1_7_2_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_7_2_sub_67_carry_2_), .S(npu_inst_pe_1_7_2_N66) );
  FA_X1 npu_inst_pe_1_7_2_add_69_U1_1 ( .A(npu_inst_pe_1_7_2_int_q_acc_1_), 
        .B(npu_inst_pe_1_7_2_int_data_1_), .CI(
        npu_inst_pe_1_7_2_add_69_carry_1_), .CO(
        npu_inst_pe_1_7_2_add_69_carry_2_), .S(npu_inst_pe_1_7_2_N74) );
  NAND3_X1 npu_inst_pe_1_7_2_U109 ( .A1(npu_inst_pe_1_7_2_n5), .A2(
        npu_inst_pe_1_7_2_n7), .A3(npu_inst_pe_1_7_2_n8), .ZN(
        npu_inst_pe_1_7_2_n44) );
  NAND3_X1 npu_inst_pe_1_7_2_U108 ( .A1(npu_inst_pe_1_7_2_n4), .A2(
        npu_inst_pe_1_7_2_n7), .A3(npu_inst_pe_1_7_2_n8), .ZN(
        npu_inst_pe_1_7_2_n40) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_7_2_n34), .CK(
        npu_inst_pe_1_7_2_net3228), .RN(npu_inst_pe_1_7_2_n9), .Q(
        npu_inst_pe_1_7_2_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_7_2_n35), .CK(
        npu_inst_pe_1_7_2_net3228), .RN(npu_inst_pe_1_7_2_n9), .Q(
        npu_inst_pe_1_7_2_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_7_2_n36), .CK(
        npu_inst_pe_1_7_2_net3228), .RN(npu_inst_pe_1_7_2_n9), .Q(
        npu_inst_pe_1_7_2_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_7_2_n98), .CK(
        npu_inst_pe_1_7_2_net3228), .RN(npu_inst_pe_1_7_2_n9), .Q(
        npu_inst_pe_1_7_2_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_7_2_n99), .CK(
        npu_inst_pe_1_7_2_net3228), .RN(npu_inst_pe_1_7_2_n9), .Q(
        npu_inst_pe_1_7_2_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_7_2_n100), 
        .CK(npu_inst_pe_1_7_2_net3228), .RN(npu_inst_pe_1_7_2_n9), .Q(
        npu_inst_pe_1_7_2_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_7_2_n33), .CK(
        npu_inst_pe_1_7_2_net3228), .RN(npu_inst_pe_1_7_2_n9), .Q(
        npu_inst_pe_1_7_2_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_7_2_n101), 
        .CK(npu_inst_pe_1_7_2_net3228), .RN(npu_inst_pe_1_7_2_n9), .Q(
        npu_inst_pe_1_7_2_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_weight_reg_0_ ( .D(npu_inst_n108), .CK(
        npu_inst_pe_1_7_2_net3234), .RN(npu_inst_pe_1_7_2_n9), .Q(
        npu_inst_pe_1_7_2_int_q_weight_0_), .QN(npu_inst_pe_1_7_2_n27) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_weight_reg_1_ ( .D(npu_inst_n114), .CK(
        npu_inst_pe_1_7_2_net3234), .RN(npu_inst_pe_1_7_2_n9), .Q(
        npu_inst_pe_1_7_2_int_q_weight_1_), .QN(npu_inst_pe_1_7_2_n26) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_7_2_n113), 
        .CK(npu_inst_pe_1_7_2_net3234), .RN(npu_inst_pe_1_7_2_n9), .Q(
        npu_inst_pe_1_7_2_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_7_2_n112), 
        .CK(npu_inst_pe_1_7_2_net3234), .RN(npu_inst_pe_1_7_2_n9), .Q(
        npu_inst_pe_1_7_2_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_7_2_n111), 
        .CK(npu_inst_pe_1_7_2_net3234), .RN(npu_inst_pe_1_7_2_n10), .Q(
        npu_inst_pe_1_7_2_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_7_2_n110), 
        .CK(npu_inst_pe_1_7_2_net3234), .RN(npu_inst_pe_1_7_2_n10), .Q(
        npu_inst_pe_1_7_2_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_7_2_n109), 
        .CK(npu_inst_pe_1_7_2_net3234), .RN(npu_inst_pe_1_7_2_n10), .Q(
        npu_inst_pe_1_7_2_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_7_2_n108), 
        .CK(npu_inst_pe_1_7_2_net3234), .RN(npu_inst_pe_1_7_2_n10), .Q(
        npu_inst_pe_1_7_2_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_7_2_n107), 
        .CK(npu_inst_pe_1_7_2_net3234), .RN(npu_inst_pe_1_7_2_n10), .Q(
        npu_inst_pe_1_7_2_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_7_2_n106), 
        .CK(npu_inst_pe_1_7_2_net3234), .RN(npu_inst_pe_1_7_2_n10), .Q(
        npu_inst_pe_1_7_2_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_7_2_n105), 
        .CK(npu_inst_pe_1_7_2_net3234), .RN(npu_inst_pe_1_7_2_n10), .Q(
        npu_inst_pe_1_7_2_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_7_2_n104), 
        .CK(npu_inst_pe_1_7_2_net3234), .RN(npu_inst_pe_1_7_2_n10), .Q(
        npu_inst_pe_1_7_2_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_7_2_n103), 
        .CK(npu_inst_pe_1_7_2_net3234), .RN(npu_inst_pe_1_7_2_n10), .Q(
        npu_inst_pe_1_7_2_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_7_2_n102), 
        .CK(npu_inst_pe_1_7_2_net3234), .RN(npu_inst_pe_1_7_2_n10), .Q(
        npu_inst_pe_1_7_2_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_7_2_n86), 
        .CK(npu_inst_pe_1_7_2_net3234), .RN(npu_inst_pe_1_7_2_n10), .Q(
        npu_inst_pe_1_7_2_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_7_2_n87), 
        .CK(npu_inst_pe_1_7_2_net3234), .RN(npu_inst_pe_1_7_2_n10), .Q(
        npu_inst_pe_1_7_2_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_7_2_n88), 
        .CK(npu_inst_pe_1_7_2_net3234), .RN(npu_inst_pe_1_7_2_n11), .Q(
        npu_inst_pe_1_7_2_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_7_2_n89), 
        .CK(npu_inst_pe_1_7_2_net3234), .RN(npu_inst_pe_1_7_2_n11), .Q(
        npu_inst_pe_1_7_2_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_7_2_n90), 
        .CK(npu_inst_pe_1_7_2_net3234), .RN(npu_inst_pe_1_7_2_n11), .Q(
        npu_inst_pe_1_7_2_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_7_2_n91), 
        .CK(npu_inst_pe_1_7_2_net3234), .RN(npu_inst_pe_1_7_2_n11), .Q(
        npu_inst_pe_1_7_2_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_7_2_n92), 
        .CK(npu_inst_pe_1_7_2_net3234), .RN(npu_inst_pe_1_7_2_n11), .Q(
        npu_inst_pe_1_7_2_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_7_2_n93), 
        .CK(npu_inst_pe_1_7_2_net3234), .RN(npu_inst_pe_1_7_2_n11), .Q(
        npu_inst_pe_1_7_2_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_7_2_n94), 
        .CK(npu_inst_pe_1_7_2_net3234), .RN(npu_inst_pe_1_7_2_n11), .Q(
        npu_inst_pe_1_7_2_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_7_2_n95), 
        .CK(npu_inst_pe_1_7_2_net3234), .RN(npu_inst_pe_1_7_2_n11), .Q(
        npu_inst_pe_1_7_2_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_7_2_n96), 
        .CK(npu_inst_pe_1_7_2_net3234), .RN(npu_inst_pe_1_7_2_n11), .Q(
        npu_inst_pe_1_7_2_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_7_2_n97), 
        .CK(npu_inst_pe_1_7_2_net3234), .RN(npu_inst_pe_1_7_2_n11), .Q(
        npu_inst_pe_1_7_2_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_7_2_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_7_2_N84), .SE(1'b0), .GCK(npu_inst_pe_1_7_2_net3228) );
  CLKGATETST_X1 npu_inst_pe_1_7_2_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n61), .SE(1'b0), .GCK(npu_inst_pe_1_7_2_net3234) );
  MUX2_X1 npu_inst_pe_1_7_3_U162 ( .A(npu_inst_pe_1_7_3_n32), .B(
        npu_inst_pe_1_7_3_n29), .S(npu_inst_pe_1_7_3_n8), .Z(
        npu_inst_pe_1_7_3_N93) );
  MUX2_X1 npu_inst_pe_1_7_3_U161 ( .A(npu_inst_pe_1_7_3_n31), .B(
        npu_inst_pe_1_7_3_n30), .S(npu_inst_pe_1_7_3_n6), .Z(
        npu_inst_pe_1_7_3_n32) );
  MUX2_X1 npu_inst_pe_1_7_3_U160 ( .A(npu_inst_pe_1_7_3_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_7_3_int_q_reg_v_1__0_), .S(npu_inst_pe_1_7_3_n4), .Z(
        npu_inst_pe_1_7_3_n31) );
  MUX2_X1 npu_inst_pe_1_7_3_U159 ( .A(npu_inst_pe_1_7_3_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_7_3_int_q_reg_v_3__0_), .S(npu_inst_pe_1_7_3_n4), .Z(
        npu_inst_pe_1_7_3_n30) );
  MUX2_X1 npu_inst_pe_1_7_3_U158 ( .A(npu_inst_pe_1_7_3_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_7_3_int_q_reg_v_5__0_), .S(npu_inst_pe_1_7_3_n4), .Z(
        npu_inst_pe_1_7_3_n29) );
  MUX2_X1 npu_inst_pe_1_7_3_U157 ( .A(npu_inst_pe_1_7_3_n28), .B(
        npu_inst_pe_1_7_3_n23), .S(npu_inst_pe_1_7_3_n8), .Z(
        npu_inst_pe_1_7_3_N94) );
  MUX2_X1 npu_inst_pe_1_7_3_U156 ( .A(npu_inst_pe_1_7_3_n25), .B(
        npu_inst_pe_1_7_3_n24), .S(npu_inst_pe_1_7_3_n6), .Z(
        npu_inst_pe_1_7_3_n28) );
  MUX2_X1 npu_inst_pe_1_7_3_U155 ( .A(npu_inst_pe_1_7_3_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_7_3_int_q_reg_v_1__1_), .S(npu_inst_pe_1_7_3_n4), .Z(
        npu_inst_pe_1_7_3_n25) );
  MUX2_X1 npu_inst_pe_1_7_3_U154 ( .A(npu_inst_pe_1_7_3_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_7_3_int_q_reg_v_3__1_), .S(npu_inst_pe_1_7_3_n4), .Z(
        npu_inst_pe_1_7_3_n24) );
  MUX2_X1 npu_inst_pe_1_7_3_U153 ( .A(npu_inst_pe_1_7_3_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_7_3_int_q_reg_v_5__1_), .S(npu_inst_pe_1_7_3_n4), .Z(
        npu_inst_pe_1_7_3_n23) );
  MUX2_X1 npu_inst_pe_1_7_3_U152 ( .A(npu_inst_pe_1_7_3_n22), .B(
        npu_inst_pe_1_7_3_n19), .S(npu_inst_pe_1_7_3_n8), .Z(
        npu_inst_int_data_x_7__3__1_) );
  MUX2_X1 npu_inst_pe_1_7_3_U151 ( .A(npu_inst_pe_1_7_3_n21), .B(
        npu_inst_pe_1_7_3_n20), .S(npu_inst_pe_1_7_3_n6), .Z(
        npu_inst_pe_1_7_3_n22) );
  MUX2_X1 npu_inst_pe_1_7_3_U150 ( .A(npu_inst_pe_1_7_3_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_7_3_int_q_reg_h_1__1_), .S(npu_inst_pe_1_7_3_n4), .Z(
        npu_inst_pe_1_7_3_n21) );
  MUX2_X1 npu_inst_pe_1_7_3_U149 ( .A(npu_inst_pe_1_7_3_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_7_3_int_q_reg_h_3__1_), .S(npu_inst_pe_1_7_3_n4), .Z(
        npu_inst_pe_1_7_3_n20) );
  MUX2_X1 npu_inst_pe_1_7_3_U148 ( .A(npu_inst_pe_1_7_3_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_7_3_int_q_reg_h_5__1_), .S(npu_inst_pe_1_7_3_n4), .Z(
        npu_inst_pe_1_7_3_n19) );
  MUX2_X1 npu_inst_pe_1_7_3_U147 ( .A(npu_inst_pe_1_7_3_n18), .B(
        npu_inst_pe_1_7_3_n15), .S(npu_inst_pe_1_7_3_n8), .Z(
        npu_inst_int_data_x_7__3__0_) );
  MUX2_X1 npu_inst_pe_1_7_3_U146 ( .A(npu_inst_pe_1_7_3_n17), .B(
        npu_inst_pe_1_7_3_n16), .S(npu_inst_pe_1_7_3_n6), .Z(
        npu_inst_pe_1_7_3_n18) );
  MUX2_X1 npu_inst_pe_1_7_3_U145 ( .A(npu_inst_pe_1_7_3_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_7_3_int_q_reg_h_1__0_), .S(npu_inst_pe_1_7_3_n4), .Z(
        npu_inst_pe_1_7_3_n17) );
  MUX2_X1 npu_inst_pe_1_7_3_U144 ( .A(npu_inst_pe_1_7_3_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_7_3_int_q_reg_h_3__0_), .S(npu_inst_pe_1_7_3_n4), .Z(
        npu_inst_pe_1_7_3_n16) );
  MUX2_X1 npu_inst_pe_1_7_3_U143 ( .A(npu_inst_pe_1_7_3_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_7_3_int_q_reg_h_5__0_), .S(npu_inst_pe_1_7_3_n4), .Z(
        npu_inst_pe_1_7_3_n15) );
  XOR2_X1 npu_inst_pe_1_7_3_U142 ( .A(npu_inst_pe_1_7_3_int_data_0_), .B(
        npu_inst_pe_1_7_3_int_q_acc_0_), .Z(npu_inst_pe_1_7_3_N73) );
  AND2_X1 npu_inst_pe_1_7_3_U141 ( .A1(npu_inst_pe_1_7_3_int_q_acc_0_), .A2(
        npu_inst_pe_1_7_3_int_data_0_), .ZN(npu_inst_pe_1_7_3_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_7_3_U140 ( .A(npu_inst_pe_1_7_3_int_q_acc_0_), .B(
        npu_inst_pe_1_7_3_n13), .ZN(npu_inst_pe_1_7_3_N65) );
  OR2_X1 npu_inst_pe_1_7_3_U139 ( .A1(npu_inst_pe_1_7_3_n13), .A2(
        npu_inst_pe_1_7_3_int_q_acc_0_), .ZN(npu_inst_pe_1_7_3_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_7_3_U138 ( .A(npu_inst_pe_1_7_3_int_q_acc_2_), .B(
        npu_inst_pe_1_7_3_add_69_carry_2_), .Z(npu_inst_pe_1_7_3_N75) );
  AND2_X1 npu_inst_pe_1_7_3_U137 ( .A1(npu_inst_pe_1_7_3_add_69_carry_2_), 
        .A2(npu_inst_pe_1_7_3_int_q_acc_2_), .ZN(
        npu_inst_pe_1_7_3_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_7_3_U136 ( .A(npu_inst_pe_1_7_3_int_q_acc_3_), .B(
        npu_inst_pe_1_7_3_add_69_carry_3_), .Z(npu_inst_pe_1_7_3_N76) );
  AND2_X1 npu_inst_pe_1_7_3_U135 ( .A1(npu_inst_pe_1_7_3_add_69_carry_3_), 
        .A2(npu_inst_pe_1_7_3_int_q_acc_3_), .ZN(
        npu_inst_pe_1_7_3_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_7_3_U134 ( .A(npu_inst_pe_1_7_3_int_q_acc_4_), .B(
        npu_inst_pe_1_7_3_add_69_carry_4_), .Z(npu_inst_pe_1_7_3_N77) );
  AND2_X1 npu_inst_pe_1_7_3_U133 ( .A1(npu_inst_pe_1_7_3_add_69_carry_4_), 
        .A2(npu_inst_pe_1_7_3_int_q_acc_4_), .ZN(
        npu_inst_pe_1_7_3_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_7_3_U132 ( .A(npu_inst_pe_1_7_3_int_q_acc_5_), .B(
        npu_inst_pe_1_7_3_add_69_carry_5_), .Z(npu_inst_pe_1_7_3_N78) );
  AND2_X1 npu_inst_pe_1_7_3_U131 ( .A1(npu_inst_pe_1_7_3_add_69_carry_5_), 
        .A2(npu_inst_pe_1_7_3_int_q_acc_5_), .ZN(
        npu_inst_pe_1_7_3_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_7_3_U130 ( .A(npu_inst_pe_1_7_3_int_q_acc_6_), .B(
        npu_inst_pe_1_7_3_add_69_carry_6_), .Z(npu_inst_pe_1_7_3_N79) );
  AND2_X1 npu_inst_pe_1_7_3_U129 ( .A1(npu_inst_pe_1_7_3_add_69_carry_6_), 
        .A2(npu_inst_pe_1_7_3_int_q_acc_6_), .ZN(
        npu_inst_pe_1_7_3_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_7_3_U128 ( .A(npu_inst_pe_1_7_3_int_q_acc_7_), .B(
        npu_inst_pe_1_7_3_add_69_carry_7_), .Z(npu_inst_pe_1_7_3_N80) );
  XNOR2_X1 npu_inst_pe_1_7_3_U127 ( .A(npu_inst_pe_1_7_3_sub_67_carry_2_), .B(
        npu_inst_pe_1_7_3_int_q_acc_2_), .ZN(npu_inst_pe_1_7_3_N67) );
  OR2_X1 npu_inst_pe_1_7_3_U126 ( .A1(npu_inst_pe_1_7_3_int_q_acc_2_), .A2(
        npu_inst_pe_1_7_3_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_7_3_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_7_3_U125 ( .A(npu_inst_pe_1_7_3_sub_67_carry_3_), .B(
        npu_inst_pe_1_7_3_int_q_acc_3_), .ZN(npu_inst_pe_1_7_3_N68) );
  OR2_X1 npu_inst_pe_1_7_3_U124 ( .A1(npu_inst_pe_1_7_3_int_q_acc_3_), .A2(
        npu_inst_pe_1_7_3_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_7_3_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_7_3_U123 ( .A(npu_inst_pe_1_7_3_sub_67_carry_4_), .B(
        npu_inst_pe_1_7_3_int_q_acc_4_), .ZN(npu_inst_pe_1_7_3_N69) );
  OR2_X1 npu_inst_pe_1_7_3_U122 ( .A1(npu_inst_pe_1_7_3_int_q_acc_4_), .A2(
        npu_inst_pe_1_7_3_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_7_3_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_7_3_U121 ( .A(npu_inst_pe_1_7_3_sub_67_carry_5_), .B(
        npu_inst_pe_1_7_3_int_q_acc_5_), .ZN(npu_inst_pe_1_7_3_N70) );
  OR2_X1 npu_inst_pe_1_7_3_U120 ( .A1(npu_inst_pe_1_7_3_int_q_acc_5_), .A2(
        npu_inst_pe_1_7_3_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_7_3_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_7_3_U119 ( .A(npu_inst_pe_1_7_3_sub_67_carry_6_), .B(
        npu_inst_pe_1_7_3_int_q_acc_6_), .ZN(npu_inst_pe_1_7_3_N71) );
  OR2_X1 npu_inst_pe_1_7_3_U118 ( .A1(npu_inst_pe_1_7_3_int_q_acc_6_), .A2(
        npu_inst_pe_1_7_3_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_7_3_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_7_3_U117 ( .A(npu_inst_pe_1_7_3_int_q_acc_7_), .B(
        npu_inst_pe_1_7_3_sub_67_carry_7_), .ZN(npu_inst_pe_1_7_3_N72) );
  INV_X1 npu_inst_pe_1_7_3_U116 ( .A(npu_inst_n75), .ZN(npu_inst_pe_1_7_3_n7)
         );
  INV_X1 npu_inst_pe_1_7_3_U115 ( .A(npu_inst_pe_1_7_3_n7), .ZN(
        npu_inst_pe_1_7_3_n6) );
  INV_X1 npu_inst_pe_1_7_3_U114 ( .A(npu_inst_n52), .ZN(npu_inst_pe_1_7_3_n3)
         );
  AOI22_X1 npu_inst_pe_1_7_3_U113 ( .A1(npu_inst_pe_1_7_3_n38), .A2(
        int_i_data_v_npu[9]), .B1(npu_inst_pe_1_7_3_n114), .B2(
        npu_inst_pe_1_7_3_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_7_3_n39) );
  INV_X1 npu_inst_pe_1_7_3_U112 ( .A(npu_inst_pe_1_7_3_n39), .ZN(
        npu_inst_pe_1_7_3_n112) );
  AOI22_X1 npu_inst_pe_1_7_3_U111 ( .A1(npu_inst_pe_1_7_3_n38), .A2(
        int_i_data_v_npu[8]), .B1(npu_inst_pe_1_7_3_n114), .B2(
        npu_inst_pe_1_7_3_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_7_3_n37) );
  INV_X1 npu_inst_pe_1_7_3_U110 ( .A(npu_inst_pe_1_7_3_n37), .ZN(
        npu_inst_pe_1_7_3_n113) );
  AOI22_X1 npu_inst_pe_1_7_3_U107 ( .A1(int_i_data_v_npu[9]), .A2(
        npu_inst_pe_1_7_3_n58), .B1(npu_inst_pe_1_7_3_n119), .B2(
        npu_inst_pe_1_7_3_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_7_3_n59) );
  INV_X1 npu_inst_pe_1_7_3_U106 ( .A(npu_inst_pe_1_7_3_n59), .ZN(
        npu_inst_pe_1_7_3_n102) );
  AOI22_X1 npu_inst_pe_1_7_3_U105 ( .A1(int_i_data_v_npu[8]), .A2(
        npu_inst_pe_1_7_3_n58), .B1(npu_inst_pe_1_7_3_n119), .B2(
        npu_inst_pe_1_7_3_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_7_3_n57) );
  INV_X1 npu_inst_pe_1_7_3_U104 ( .A(npu_inst_pe_1_7_3_n57), .ZN(
        npu_inst_pe_1_7_3_n103) );
  AOI22_X1 npu_inst_pe_1_7_3_U103 ( .A1(int_i_data_v_npu[9]), .A2(
        npu_inst_pe_1_7_3_n54), .B1(npu_inst_pe_1_7_3_n118), .B2(
        npu_inst_pe_1_7_3_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_7_3_n55) );
  INV_X1 npu_inst_pe_1_7_3_U102 ( .A(npu_inst_pe_1_7_3_n55), .ZN(
        npu_inst_pe_1_7_3_n104) );
  AOI22_X1 npu_inst_pe_1_7_3_U101 ( .A1(int_i_data_v_npu[8]), .A2(
        npu_inst_pe_1_7_3_n54), .B1(npu_inst_pe_1_7_3_n118), .B2(
        npu_inst_pe_1_7_3_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_7_3_n53) );
  INV_X1 npu_inst_pe_1_7_3_U100 ( .A(npu_inst_pe_1_7_3_n53), .ZN(
        npu_inst_pe_1_7_3_n105) );
  AOI22_X1 npu_inst_pe_1_7_3_U99 ( .A1(int_i_data_v_npu[9]), .A2(
        npu_inst_pe_1_7_3_n50), .B1(npu_inst_pe_1_7_3_n117), .B2(
        npu_inst_pe_1_7_3_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_7_3_n51) );
  INV_X1 npu_inst_pe_1_7_3_U98 ( .A(npu_inst_pe_1_7_3_n51), .ZN(
        npu_inst_pe_1_7_3_n106) );
  AOI22_X1 npu_inst_pe_1_7_3_U97 ( .A1(int_i_data_v_npu[8]), .A2(
        npu_inst_pe_1_7_3_n50), .B1(npu_inst_pe_1_7_3_n117), .B2(
        npu_inst_pe_1_7_3_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_7_3_n49) );
  INV_X1 npu_inst_pe_1_7_3_U96 ( .A(npu_inst_pe_1_7_3_n49), .ZN(
        npu_inst_pe_1_7_3_n107) );
  AOI22_X1 npu_inst_pe_1_7_3_U95 ( .A1(int_i_data_v_npu[9]), .A2(
        npu_inst_pe_1_7_3_n46), .B1(npu_inst_pe_1_7_3_n116), .B2(
        npu_inst_pe_1_7_3_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_7_3_n47) );
  INV_X1 npu_inst_pe_1_7_3_U94 ( .A(npu_inst_pe_1_7_3_n47), .ZN(
        npu_inst_pe_1_7_3_n108) );
  AOI22_X1 npu_inst_pe_1_7_3_U93 ( .A1(int_i_data_v_npu[8]), .A2(
        npu_inst_pe_1_7_3_n46), .B1(npu_inst_pe_1_7_3_n116), .B2(
        npu_inst_pe_1_7_3_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_7_3_n45) );
  INV_X1 npu_inst_pe_1_7_3_U92 ( .A(npu_inst_pe_1_7_3_n45), .ZN(
        npu_inst_pe_1_7_3_n109) );
  AOI22_X1 npu_inst_pe_1_7_3_U91 ( .A1(int_i_data_v_npu[9]), .A2(
        npu_inst_pe_1_7_3_n42), .B1(npu_inst_pe_1_7_3_n115), .B2(
        npu_inst_pe_1_7_3_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_7_3_n43) );
  INV_X1 npu_inst_pe_1_7_3_U90 ( .A(npu_inst_pe_1_7_3_n43), .ZN(
        npu_inst_pe_1_7_3_n110) );
  AOI22_X1 npu_inst_pe_1_7_3_U89 ( .A1(int_i_data_v_npu[8]), .A2(
        npu_inst_pe_1_7_3_n42), .B1(npu_inst_pe_1_7_3_n115), .B2(
        npu_inst_pe_1_7_3_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_7_3_n41) );
  INV_X1 npu_inst_pe_1_7_3_U88 ( .A(npu_inst_pe_1_7_3_n41), .ZN(
        npu_inst_pe_1_7_3_n111) );
  NAND2_X1 npu_inst_pe_1_7_3_U87 ( .A1(npu_inst_pe_1_7_3_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_7_3_n60), .ZN(npu_inst_pe_1_7_3_n74) );
  OAI21_X1 npu_inst_pe_1_7_3_U86 ( .B1(npu_inst_pe_1_7_3_n63), .B2(
        npu_inst_pe_1_7_3_n60), .A(npu_inst_pe_1_7_3_n74), .ZN(
        npu_inst_pe_1_7_3_n97) );
  NAND2_X1 npu_inst_pe_1_7_3_U85 ( .A1(npu_inst_pe_1_7_3_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_7_3_n60), .ZN(npu_inst_pe_1_7_3_n73) );
  OAI21_X1 npu_inst_pe_1_7_3_U84 ( .B1(npu_inst_pe_1_7_3_n61), .B2(
        npu_inst_pe_1_7_3_n60), .A(npu_inst_pe_1_7_3_n73), .ZN(
        npu_inst_pe_1_7_3_n96) );
  NAND2_X1 npu_inst_pe_1_7_3_U83 ( .A1(npu_inst_pe_1_7_3_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_7_3_n56), .ZN(npu_inst_pe_1_7_3_n72) );
  OAI21_X1 npu_inst_pe_1_7_3_U82 ( .B1(npu_inst_pe_1_7_3_n63), .B2(
        npu_inst_pe_1_7_3_n56), .A(npu_inst_pe_1_7_3_n72), .ZN(
        npu_inst_pe_1_7_3_n95) );
  NAND2_X1 npu_inst_pe_1_7_3_U81 ( .A1(npu_inst_pe_1_7_3_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_7_3_n56), .ZN(npu_inst_pe_1_7_3_n71) );
  OAI21_X1 npu_inst_pe_1_7_3_U80 ( .B1(npu_inst_pe_1_7_3_n61), .B2(
        npu_inst_pe_1_7_3_n56), .A(npu_inst_pe_1_7_3_n71), .ZN(
        npu_inst_pe_1_7_3_n94) );
  NAND2_X1 npu_inst_pe_1_7_3_U79 ( .A1(npu_inst_pe_1_7_3_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_7_3_n52), .ZN(npu_inst_pe_1_7_3_n70) );
  OAI21_X1 npu_inst_pe_1_7_3_U78 ( .B1(npu_inst_pe_1_7_3_n63), .B2(
        npu_inst_pe_1_7_3_n52), .A(npu_inst_pe_1_7_3_n70), .ZN(
        npu_inst_pe_1_7_3_n93) );
  NAND2_X1 npu_inst_pe_1_7_3_U77 ( .A1(npu_inst_pe_1_7_3_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_7_3_n52), .ZN(npu_inst_pe_1_7_3_n69) );
  OAI21_X1 npu_inst_pe_1_7_3_U76 ( .B1(npu_inst_pe_1_7_3_n61), .B2(
        npu_inst_pe_1_7_3_n52), .A(npu_inst_pe_1_7_3_n69), .ZN(
        npu_inst_pe_1_7_3_n92) );
  NAND2_X1 npu_inst_pe_1_7_3_U75 ( .A1(npu_inst_pe_1_7_3_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_7_3_n48), .ZN(npu_inst_pe_1_7_3_n68) );
  OAI21_X1 npu_inst_pe_1_7_3_U74 ( .B1(npu_inst_pe_1_7_3_n63), .B2(
        npu_inst_pe_1_7_3_n48), .A(npu_inst_pe_1_7_3_n68), .ZN(
        npu_inst_pe_1_7_3_n91) );
  NAND2_X1 npu_inst_pe_1_7_3_U73 ( .A1(npu_inst_pe_1_7_3_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_7_3_n48), .ZN(npu_inst_pe_1_7_3_n67) );
  OAI21_X1 npu_inst_pe_1_7_3_U72 ( .B1(npu_inst_pe_1_7_3_n61), .B2(
        npu_inst_pe_1_7_3_n48), .A(npu_inst_pe_1_7_3_n67), .ZN(
        npu_inst_pe_1_7_3_n90) );
  NAND2_X1 npu_inst_pe_1_7_3_U71 ( .A1(npu_inst_pe_1_7_3_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_7_3_n44), .ZN(npu_inst_pe_1_7_3_n66) );
  OAI21_X1 npu_inst_pe_1_7_3_U70 ( .B1(npu_inst_pe_1_7_3_n63), .B2(
        npu_inst_pe_1_7_3_n44), .A(npu_inst_pe_1_7_3_n66), .ZN(
        npu_inst_pe_1_7_3_n89) );
  NAND2_X1 npu_inst_pe_1_7_3_U69 ( .A1(npu_inst_pe_1_7_3_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_7_3_n44), .ZN(npu_inst_pe_1_7_3_n65) );
  OAI21_X1 npu_inst_pe_1_7_3_U68 ( .B1(npu_inst_pe_1_7_3_n61), .B2(
        npu_inst_pe_1_7_3_n44), .A(npu_inst_pe_1_7_3_n65), .ZN(
        npu_inst_pe_1_7_3_n88) );
  NAND2_X1 npu_inst_pe_1_7_3_U67 ( .A1(npu_inst_pe_1_7_3_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_7_3_n40), .ZN(npu_inst_pe_1_7_3_n64) );
  OAI21_X1 npu_inst_pe_1_7_3_U66 ( .B1(npu_inst_pe_1_7_3_n63), .B2(
        npu_inst_pe_1_7_3_n40), .A(npu_inst_pe_1_7_3_n64), .ZN(
        npu_inst_pe_1_7_3_n87) );
  NAND2_X1 npu_inst_pe_1_7_3_U65 ( .A1(npu_inst_pe_1_7_3_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_7_3_n40), .ZN(npu_inst_pe_1_7_3_n62) );
  OAI21_X1 npu_inst_pe_1_7_3_U64 ( .B1(npu_inst_pe_1_7_3_n61), .B2(
        npu_inst_pe_1_7_3_n40), .A(npu_inst_pe_1_7_3_n62), .ZN(
        npu_inst_pe_1_7_3_n86) );
  AND2_X1 npu_inst_pe_1_7_3_U63 ( .A1(npu_inst_pe_1_7_3_N93), .A2(npu_inst_n52), .ZN(npu_inst_int_data_y_7__3__0_) );
  AND2_X1 npu_inst_pe_1_7_3_U62 ( .A1(npu_inst_n52), .A2(npu_inst_pe_1_7_3_N94), .ZN(npu_inst_int_data_y_7__3__1_) );
  AOI22_X1 npu_inst_pe_1_7_3_U61 ( .A1(npu_inst_n52), .A2(int_i_data_v_npu[9]), 
        .B1(npu_inst_pe_1_7_3_n3), .B2(npu_inst_int_data_x_7__4__1_), .ZN(
        npu_inst_pe_1_7_3_n63) );
  AOI22_X1 npu_inst_pe_1_7_3_U60 ( .A1(npu_inst_n52), .A2(int_i_data_v_npu[8]), 
        .B1(npu_inst_pe_1_7_3_n3), .B2(npu_inst_int_data_x_7__4__0_), .ZN(
        npu_inst_pe_1_7_3_n61) );
  AOI222_X1 npu_inst_pe_1_7_3_U59 ( .A1(1'b0), .A2(npu_inst_pe_1_7_3_n1), .B1(
        npu_inst_pe_1_7_3_N73), .B2(npu_inst_pe_1_7_3_n76), .C1(
        npu_inst_pe_1_7_3_N65), .C2(npu_inst_pe_1_7_3_n77), .ZN(
        npu_inst_pe_1_7_3_n84) );
  INV_X1 npu_inst_pe_1_7_3_U58 ( .A(npu_inst_pe_1_7_3_n84), .ZN(
        npu_inst_pe_1_7_3_n101) );
  AOI222_X1 npu_inst_pe_1_7_3_U57 ( .A1(1'b0), .A2(npu_inst_pe_1_7_3_n1), .B1(
        npu_inst_pe_1_7_3_N80), .B2(npu_inst_pe_1_7_3_n76), .C1(
        npu_inst_pe_1_7_3_N72), .C2(npu_inst_pe_1_7_3_n77), .ZN(
        npu_inst_pe_1_7_3_n75) );
  INV_X1 npu_inst_pe_1_7_3_U56 ( .A(npu_inst_pe_1_7_3_n75), .ZN(
        npu_inst_pe_1_7_3_n33) );
  AOI222_X1 npu_inst_pe_1_7_3_U55 ( .A1(1'b0), .A2(npu_inst_pe_1_7_3_n1), .B1(
        npu_inst_pe_1_7_3_N74), .B2(npu_inst_pe_1_7_3_n76), .C1(
        npu_inst_pe_1_7_3_N66), .C2(npu_inst_pe_1_7_3_n77), .ZN(
        npu_inst_pe_1_7_3_n83) );
  INV_X1 npu_inst_pe_1_7_3_U54 ( .A(npu_inst_pe_1_7_3_n83), .ZN(
        npu_inst_pe_1_7_3_n100) );
  AOI222_X1 npu_inst_pe_1_7_3_U53 ( .A1(1'b0), .A2(npu_inst_pe_1_7_3_n1), .B1(
        npu_inst_pe_1_7_3_N75), .B2(npu_inst_pe_1_7_3_n76), .C1(
        npu_inst_pe_1_7_3_N67), .C2(npu_inst_pe_1_7_3_n77), .ZN(
        npu_inst_pe_1_7_3_n82) );
  INV_X1 npu_inst_pe_1_7_3_U52 ( .A(npu_inst_pe_1_7_3_n82), .ZN(
        npu_inst_pe_1_7_3_n99) );
  AOI222_X1 npu_inst_pe_1_7_3_U51 ( .A1(1'b0), .A2(npu_inst_pe_1_7_3_n1), .B1(
        npu_inst_pe_1_7_3_N76), .B2(npu_inst_pe_1_7_3_n76), .C1(
        npu_inst_pe_1_7_3_N68), .C2(npu_inst_pe_1_7_3_n77), .ZN(
        npu_inst_pe_1_7_3_n81) );
  INV_X1 npu_inst_pe_1_7_3_U50 ( .A(npu_inst_pe_1_7_3_n81), .ZN(
        npu_inst_pe_1_7_3_n98) );
  AOI222_X1 npu_inst_pe_1_7_3_U49 ( .A1(1'b0), .A2(npu_inst_pe_1_7_3_n1), .B1(
        npu_inst_pe_1_7_3_N77), .B2(npu_inst_pe_1_7_3_n76), .C1(
        npu_inst_pe_1_7_3_N69), .C2(npu_inst_pe_1_7_3_n77), .ZN(
        npu_inst_pe_1_7_3_n80) );
  INV_X1 npu_inst_pe_1_7_3_U48 ( .A(npu_inst_pe_1_7_3_n80), .ZN(
        npu_inst_pe_1_7_3_n36) );
  AOI222_X1 npu_inst_pe_1_7_3_U47 ( .A1(1'b0), .A2(npu_inst_pe_1_7_3_n1), .B1(
        npu_inst_pe_1_7_3_N78), .B2(npu_inst_pe_1_7_3_n76), .C1(
        npu_inst_pe_1_7_3_N70), .C2(npu_inst_pe_1_7_3_n77), .ZN(
        npu_inst_pe_1_7_3_n79) );
  INV_X1 npu_inst_pe_1_7_3_U46 ( .A(npu_inst_pe_1_7_3_n79), .ZN(
        npu_inst_pe_1_7_3_n35) );
  AOI222_X1 npu_inst_pe_1_7_3_U45 ( .A1(1'b0), .A2(npu_inst_pe_1_7_3_n1), .B1(
        npu_inst_pe_1_7_3_N79), .B2(npu_inst_pe_1_7_3_n76), .C1(
        npu_inst_pe_1_7_3_N71), .C2(npu_inst_pe_1_7_3_n77), .ZN(
        npu_inst_pe_1_7_3_n78) );
  INV_X1 npu_inst_pe_1_7_3_U44 ( .A(npu_inst_pe_1_7_3_n78), .ZN(
        npu_inst_pe_1_7_3_n34) );
  AND2_X1 npu_inst_pe_1_7_3_U43 ( .A1(npu_inst_pe_1_7_3_int_q_acc_0_), .A2(
        npu_inst_pe_1_7_3_n1), .ZN(npu_inst_int_data_res_7__3__0_) );
  AND2_X1 npu_inst_pe_1_7_3_U42 ( .A1(npu_inst_pe_1_7_3_n2), .A2(
        npu_inst_pe_1_7_3_int_q_acc_7_), .ZN(npu_inst_int_data_res_7__3__7_)
         );
  AND2_X1 npu_inst_pe_1_7_3_U41 ( .A1(npu_inst_pe_1_7_3_int_q_acc_1_), .A2(
        npu_inst_pe_1_7_3_n1), .ZN(npu_inst_int_data_res_7__3__1_) );
  AND2_X1 npu_inst_pe_1_7_3_U40 ( .A1(npu_inst_pe_1_7_3_int_q_acc_2_), .A2(
        npu_inst_pe_1_7_3_n1), .ZN(npu_inst_int_data_res_7__3__2_) );
  AND2_X1 npu_inst_pe_1_7_3_U39 ( .A1(npu_inst_pe_1_7_3_int_q_acc_3_), .A2(
        npu_inst_pe_1_7_3_n2), .ZN(npu_inst_int_data_res_7__3__3_) );
  AND2_X1 npu_inst_pe_1_7_3_U38 ( .A1(npu_inst_pe_1_7_3_int_q_acc_4_), .A2(
        npu_inst_pe_1_7_3_n2), .ZN(npu_inst_int_data_res_7__3__4_) );
  AND2_X1 npu_inst_pe_1_7_3_U37 ( .A1(npu_inst_pe_1_7_3_int_q_acc_5_), .A2(
        npu_inst_pe_1_7_3_n2), .ZN(npu_inst_int_data_res_7__3__5_) );
  AND2_X1 npu_inst_pe_1_7_3_U36 ( .A1(npu_inst_pe_1_7_3_int_q_acc_6_), .A2(
        npu_inst_pe_1_7_3_n2), .ZN(npu_inst_int_data_res_7__3__6_) );
  INV_X1 npu_inst_pe_1_7_3_U35 ( .A(npu_inst_pe_1_7_3_int_data_1_), .ZN(
        npu_inst_pe_1_7_3_n14) );
  NOR3_X1 npu_inst_pe_1_7_3_U34 ( .A1(npu_inst_pe_1_7_3_n26), .A2(npu_inst_n52), .A3(npu_inst_int_ckg[4]), .ZN(npu_inst_pe_1_7_3_n85) );
  OR2_X1 npu_inst_pe_1_7_3_U33 ( .A1(npu_inst_pe_1_7_3_n85), .A2(
        npu_inst_pe_1_7_3_n2), .ZN(npu_inst_pe_1_7_3_N84) );
  AND2_X1 npu_inst_pe_1_7_3_U32 ( .A1(npu_inst_int_data_x_7__3__1_), .A2(
        npu_inst_pe_1_7_3_int_q_weight_1_), .ZN(npu_inst_pe_1_7_3_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_7_3_U31 ( .A1(npu_inst_int_data_x_7__3__0_), .A2(
        npu_inst_pe_1_7_3_int_q_weight_1_), .ZN(npu_inst_pe_1_7_3_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_7_3_U30 ( .A(npu_inst_pe_1_7_3_int_data_0_), .ZN(
        npu_inst_pe_1_7_3_n13) );
  INV_X1 npu_inst_pe_1_7_3_U29 ( .A(npu_inst_n67), .ZN(npu_inst_pe_1_7_3_n5)
         );
  OR3_X1 npu_inst_pe_1_7_3_U28 ( .A1(npu_inst_pe_1_7_3_n6), .A2(
        npu_inst_pe_1_7_3_n8), .A3(npu_inst_pe_1_7_3_n5), .ZN(
        npu_inst_pe_1_7_3_n56) );
  OR3_X1 npu_inst_pe_1_7_3_U27 ( .A1(npu_inst_pe_1_7_3_n5), .A2(
        npu_inst_pe_1_7_3_n8), .A3(npu_inst_pe_1_7_3_n7), .ZN(
        npu_inst_pe_1_7_3_n48) );
  INV_X1 npu_inst_pe_1_7_3_U26 ( .A(npu_inst_pe_1_7_3_n5), .ZN(
        npu_inst_pe_1_7_3_n4) );
  OR3_X1 npu_inst_pe_1_7_3_U25 ( .A1(npu_inst_pe_1_7_3_n4), .A2(
        npu_inst_pe_1_7_3_n8), .A3(npu_inst_pe_1_7_3_n7), .ZN(
        npu_inst_pe_1_7_3_n52) );
  OR3_X1 npu_inst_pe_1_7_3_U24 ( .A1(npu_inst_pe_1_7_3_n6), .A2(
        npu_inst_pe_1_7_3_n8), .A3(npu_inst_pe_1_7_3_n4), .ZN(
        npu_inst_pe_1_7_3_n60) );
  NOR2_X1 npu_inst_pe_1_7_3_U23 ( .A1(npu_inst_pe_1_7_3_n60), .A2(
        npu_inst_pe_1_7_3_n3), .ZN(npu_inst_pe_1_7_3_n58) );
  NOR2_X1 npu_inst_pe_1_7_3_U22 ( .A1(npu_inst_pe_1_7_3_n56), .A2(
        npu_inst_pe_1_7_3_n3), .ZN(npu_inst_pe_1_7_3_n54) );
  NOR2_X1 npu_inst_pe_1_7_3_U21 ( .A1(npu_inst_pe_1_7_3_n52), .A2(
        npu_inst_pe_1_7_3_n3), .ZN(npu_inst_pe_1_7_3_n50) );
  NOR2_X1 npu_inst_pe_1_7_3_U20 ( .A1(npu_inst_pe_1_7_3_n48), .A2(
        npu_inst_pe_1_7_3_n3), .ZN(npu_inst_pe_1_7_3_n46) );
  NOR2_X1 npu_inst_pe_1_7_3_U19 ( .A1(npu_inst_pe_1_7_3_n40), .A2(
        npu_inst_pe_1_7_3_n3), .ZN(npu_inst_pe_1_7_3_n38) );
  NOR2_X1 npu_inst_pe_1_7_3_U18 ( .A1(npu_inst_pe_1_7_3_n44), .A2(
        npu_inst_pe_1_7_3_n3), .ZN(npu_inst_pe_1_7_3_n42) );
  BUF_X1 npu_inst_pe_1_7_3_U17 ( .A(npu_inst_n93), .Z(npu_inst_pe_1_7_3_n8) );
  INV_X1 npu_inst_pe_1_7_3_U16 ( .A(npu_inst_n122), .ZN(npu_inst_pe_1_7_3_n12)
         );
  INV_X1 npu_inst_pe_1_7_3_U15 ( .A(npu_inst_pe_1_7_3_n38), .ZN(
        npu_inst_pe_1_7_3_n114) );
  INV_X1 npu_inst_pe_1_7_3_U14 ( .A(npu_inst_pe_1_7_3_n58), .ZN(
        npu_inst_pe_1_7_3_n119) );
  INV_X1 npu_inst_pe_1_7_3_U13 ( .A(npu_inst_pe_1_7_3_n54), .ZN(
        npu_inst_pe_1_7_3_n118) );
  INV_X1 npu_inst_pe_1_7_3_U12 ( .A(npu_inst_pe_1_7_3_n50), .ZN(
        npu_inst_pe_1_7_3_n117) );
  INV_X1 npu_inst_pe_1_7_3_U11 ( .A(npu_inst_pe_1_7_3_n46), .ZN(
        npu_inst_pe_1_7_3_n116) );
  INV_X1 npu_inst_pe_1_7_3_U10 ( .A(npu_inst_pe_1_7_3_n42), .ZN(
        npu_inst_pe_1_7_3_n115) );
  BUF_X1 npu_inst_pe_1_7_3_U9 ( .A(npu_inst_n9), .Z(npu_inst_pe_1_7_3_n2) );
  BUF_X1 npu_inst_pe_1_7_3_U8 ( .A(npu_inst_n9), .Z(npu_inst_pe_1_7_3_n1) );
  BUF_X1 npu_inst_pe_1_7_3_U7 ( .A(npu_inst_pe_1_7_3_n12), .Z(
        npu_inst_pe_1_7_3_n11) );
  BUF_X1 npu_inst_pe_1_7_3_U6 ( .A(npu_inst_pe_1_7_3_n12), .Z(
        npu_inst_pe_1_7_3_n10) );
  BUF_X1 npu_inst_pe_1_7_3_U5 ( .A(npu_inst_pe_1_7_3_n12), .Z(
        npu_inst_pe_1_7_3_n9) );
  NOR2_X1 npu_inst_pe_1_7_3_U4 ( .A1(npu_inst_pe_1_7_3_int_q_weight_0_), .A2(
        npu_inst_pe_1_7_3_n1), .ZN(npu_inst_pe_1_7_3_n76) );
  NOR2_X1 npu_inst_pe_1_7_3_U3 ( .A1(npu_inst_pe_1_7_3_n27), .A2(
        npu_inst_pe_1_7_3_n1), .ZN(npu_inst_pe_1_7_3_n77) );
  FA_X1 npu_inst_pe_1_7_3_sub_67_U2_1 ( .A(npu_inst_pe_1_7_3_int_q_acc_1_), 
        .B(npu_inst_pe_1_7_3_n14), .CI(npu_inst_pe_1_7_3_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_7_3_sub_67_carry_2_), .S(npu_inst_pe_1_7_3_N66) );
  FA_X1 npu_inst_pe_1_7_3_add_69_U1_1 ( .A(npu_inst_pe_1_7_3_int_q_acc_1_), 
        .B(npu_inst_pe_1_7_3_int_data_1_), .CI(
        npu_inst_pe_1_7_3_add_69_carry_1_), .CO(
        npu_inst_pe_1_7_3_add_69_carry_2_), .S(npu_inst_pe_1_7_3_N74) );
  NAND3_X1 npu_inst_pe_1_7_3_U109 ( .A1(npu_inst_pe_1_7_3_n5), .A2(
        npu_inst_pe_1_7_3_n7), .A3(npu_inst_pe_1_7_3_n8), .ZN(
        npu_inst_pe_1_7_3_n44) );
  NAND3_X1 npu_inst_pe_1_7_3_U108 ( .A1(npu_inst_pe_1_7_3_n4), .A2(
        npu_inst_pe_1_7_3_n7), .A3(npu_inst_pe_1_7_3_n8), .ZN(
        npu_inst_pe_1_7_3_n40) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_7_3_n34), .CK(
        npu_inst_pe_1_7_3_net3205), .RN(npu_inst_pe_1_7_3_n9), .Q(
        npu_inst_pe_1_7_3_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_7_3_n35), .CK(
        npu_inst_pe_1_7_3_net3205), .RN(npu_inst_pe_1_7_3_n9), .Q(
        npu_inst_pe_1_7_3_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_7_3_n36), .CK(
        npu_inst_pe_1_7_3_net3205), .RN(npu_inst_pe_1_7_3_n9), .Q(
        npu_inst_pe_1_7_3_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_7_3_n98), .CK(
        npu_inst_pe_1_7_3_net3205), .RN(npu_inst_pe_1_7_3_n9), .Q(
        npu_inst_pe_1_7_3_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_7_3_n99), .CK(
        npu_inst_pe_1_7_3_net3205), .RN(npu_inst_pe_1_7_3_n9), .Q(
        npu_inst_pe_1_7_3_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_7_3_n100), 
        .CK(npu_inst_pe_1_7_3_net3205), .RN(npu_inst_pe_1_7_3_n9), .Q(
        npu_inst_pe_1_7_3_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_7_3_n33), .CK(
        npu_inst_pe_1_7_3_net3205), .RN(npu_inst_pe_1_7_3_n9), .Q(
        npu_inst_pe_1_7_3_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_7_3_n101), 
        .CK(npu_inst_pe_1_7_3_net3205), .RN(npu_inst_pe_1_7_3_n9), .Q(
        npu_inst_pe_1_7_3_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_weight_reg_0_ ( .D(npu_inst_n108), .CK(
        npu_inst_pe_1_7_3_net3211), .RN(npu_inst_pe_1_7_3_n9), .Q(
        npu_inst_pe_1_7_3_int_q_weight_0_), .QN(npu_inst_pe_1_7_3_n27) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_weight_reg_1_ ( .D(npu_inst_n114), .CK(
        npu_inst_pe_1_7_3_net3211), .RN(npu_inst_pe_1_7_3_n9), .Q(
        npu_inst_pe_1_7_3_int_q_weight_1_), .QN(npu_inst_pe_1_7_3_n26) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_7_3_n113), 
        .CK(npu_inst_pe_1_7_3_net3211), .RN(npu_inst_pe_1_7_3_n9), .Q(
        npu_inst_pe_1_7_3_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_7_3_n112), 
        .CK(npu_inst_pe_1_7_3_net3211), .RN(npu_inst_pe_1_7_3_n9), .Q(
        npu_inst_pe_1_7_3_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_7_3_n111), 
        .CK(npu_inst_pe_1_7_3_net3211), .RN(npu_inst_pe_1_7_3_n10), .Q(
        npu_inst_pe_1_7_3_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_7_3_n110), 
        .CK(npu_inst_pe_1_7_3_net3211), .RN(npu_inst_pe_1_7_3_n10), .Q(
        npu_inst_pe_1_7_3_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_7_3_n109), 
        .CK(npu_inst_pe_1_7_3_net3211), .RN(npu_inst_pe_1_7_3_n10), .Q(
        npu_inst_pe_1_7_3_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_7_3_n108), 
        .CK(npu_inst_pe_1_7_3_net3211), .RN(npu_inst_pe_1_7_3_n10), .Q(
        npu_inst_pe_1_7_3_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_7_3_n107), 
        .CK(npu_inst_pe_1_7_3_net3211), .RN(npu_inst_pe_1_7_3_n10), .Q(
        npu_inst_pe_1_7_3_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_7_3_n106), 
        .CK(npu_inst_pe_1_7_3_net3211), .RN(npu_inst_pe_1_7_3_n10), .Q(
        npu_inst_pe_1_7_3_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_7_3_n105), 
        .CK(npu_inst_pe_1_7_3_net3211), .RN(npu_inst_pe_1_7_3_n10), .Q(
        npu_inst_pe_1_7_3_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_7_3_n104), 
        .CK(npu_inst_pe_1_7_3_net3211), .RN(npu_inst_pe_1_7_3_n10), .Q(
        npu_inst_pe_1_7_3_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_7_3_n103), 
        .CK(npu_inst_pe_1_7_3_net3211), .RN(npu_inst_pe_1_7_3_n10), .Q(
        npu_inst_pe_1_7_3_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_7_3_n102), 
        .CK(npu_inst_pe_1_7_3_net3211), .RN(npu_inst_pe_1_7_3_n10), .Q(
        npu_inst_pe_1_7_3_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_7_3_n86), 
        .CK(npu_inst_pe_1_7_3_net3211), .RN(npu_inst_pe_1_7_3_n10), .Q(
        npu_inst_pe_1_7_3_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_7_3_n87), 
        .CK(npu_inst_pe_1_7_3_net3211), .RN(npu_inst_pe_1_7_3_n10), .Q(
        npu_inst_pe_1_7_3_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_7_3_n88), 
        .CK(npu_inst_pe_1_7_3_net3211), .RN(npu_inst_pe_1_7_3_n11), .Q(
        npu_inst_pe_1_7_3_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_7_3_n89), 
        .CK(npu_inst_pe_1_7_3_net3211), .RN(npu_inst_pe_1_7_3_n11), .Q(
        npu_inst_pe_1_7_3_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_7_3_n90), 
        .CK(npu_inst_pe_1_7_3_net3211), .RN(npu_inst_pe_1_7_3_n11), .Q(
        npu_inst_pe_1_7_3_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_7_3_n91), 
        .CK(npu_inst_pe_1_7_3_net3211), .RN(npu_inst_pe_1_7_3_n11), .Q(
        npu_inst_pe_1_7_3_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_7_3_n92), 
        .CK(npu_inst_pe_1_7_3_net3211), .RN(npu_inst_pe_1_7_3_n11), .Q(
        npu_inst_pe_1_7_3_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_7_3_n93), 
        .CK(npu_inst_pe_1_7_3_net3211), .RN(npu_inst_pe_1_7_3_n11), .Q(
        npu_inst_pe_1_7_3_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_7_3_n94), 
        .CK(npu_inst_pe_1_7_3_net3211), .RN(npu_inst_pe_1_7_3_n11), .Q(
        npu_inst_pe_1_7_3_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_7_3_n95), 
        .CK(npu_inst_pe_1_7_3_net3211), .RN(npu_inst_pe_1_7_3_n11), .Q(
        npu_inst_pe_1_7_3_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_7_3_n96), 
        .CK(npu_inst_pe_1_7_3_net3211), .RN(npu_inst_pe_1_7_3_n11), .Q(
        npu_inst_pe_1_7_3_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_7_3_n97), 
        .CK(npu_inst_pe_1_7_3_net3211), .RN(npu_inst_pe_1_7_3_n11), .Q(
        npu_inst_pe_1_7_3_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_7_3_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_7_3_N84), .SE(1'b0), .GCK(npu_inst_pe_1_7_3_net3205) );
  CLKGATETST_X1 npu_inst_pe_1_7_3_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n61), .SE(1'b0), .GCK(npu_inst_pe_1_7_3_net3211) );
  MUX2_X1 npu_inst_pe_1_7_4_U162 ( .A(npu_inst_pe_1_7_4_n32), .B(
        npu_inst_pe_1_7_4_n29), .S(npu_inst_pe_1_7_4_n8), .Z(
        npu_inst_pe_1_7_4_N93) );
  MUX2_X1 npu_inst_pe_1_7_4_U161 ( .A(npu_inst_pe_1_7_4_n31), .B(
        npu_inst_pe_1_7_4_n30), .S(npu_inst_pe_1_7_4_n6), .Z(
        npu_inst_pe_1_7_4_n32) );
  MUX2_X1 npu_inst_pe_1_7_4_U160 ( .A(npu_inst_pe_1_7_4_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_7_4_int_q_reg_v_1__0_), .S(npu_inst_pe_1_7_4_n4), .Z(
        npu_inst_pe_1_7_4_n31) );
  MUX2_X1 npu_inst_pe_1_7_4_U159 ( .A(npu_inst_pe_1_7_4_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_7_4_int_q_reg_v_3__0_), .S(npu_inst_pe_1_7_4_n4), .Z(
        npu_inst_pe_1_7_4_n30) );
  MUX2_X1 npu_inst_pe_1_7_4_U158 ( .A(npu_inst_pe_1_7_4_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_7_4_int_q_reg_v_5__0_), .S(npu_inst_pe_1_7_4_n4), .Z(
        npu_inst_pe_1_7_4_n29) );
  MUX2_X1 npu_inst_pe_1_7_4_U157 ( .A(npu_inst_pe_1_7_4_n28), .B(
        npu_inst_pe_1_7_4_n23), .S(npu_inst_pe_1_7_4_n8), .Z(
        npu_inst_pe_1_7_4_N94) );
  MUX2_X1 npu_inst_pe_1_7_4_U156 ( .A(npu_inst_pe_1_7_4_n25), .B(
        npu_inst_pe_1_7_4_n24), .S(npu_inst_pe_1_7_4_n6), .Z(
        npu_inst_pe_1_7_4_n28) );
  MUX2_X1 npu_inst_pe_1_7_4_U155 ( .A(npu_inst_pe_1_7_4_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_7_4_int_q_reg_v_1__1_), .S(npu_inst_pe_1_7_4_n4), .Z(
        npu_inst_pe_1_7_4_n25) );
  MUX2_X1 npu_inst_pe_1_7_4_U154 ( .A(npu_inst_pe_1_7_4_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_7_4_int_q_reg_v_3__1_), .S(npu_inst_pe_1_7_4_n4), .Z(
        npu_inst_pe_1_7_4_n24) );
  MUX2_X1 npu_inst_pe_1_7_4_U153 ( .A(npu_inst_pe_1_7_4_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_7_4_int_q_reg_v_5__1_), .S(npu_inst_pe_1_7_4_n4), .Z(
        npu_inst_pe_1_7_4_n23) );
  MUX2_X1 npu_inst_pe_1_7_4_U152 ( .A(npu_inst_pe_1_7_4_n22), .B(
        npu_inst_pe_1_7_4_n19), .S(npu_inst_pe_1_7_4_n8), .Z(
        npu_inst_int_data_x_7__4__1_) );
  MUX2_X1 npu_inst_pe_1_7_4_U151 ( .A(npu_inst_pe_1_7_4_n21), .B(
        npu_inst_pe_1_7_4_n20), .S(npu_inst_pe_1_7_4_n6), .Z(
        npu_inst_pe_1_7_4_n22) );
  MUX2_X1 npu_inst_pe_1_7_4_U150 ( .A(npu_inst_pe_1_7_4_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_7_4_int_q_reg_h_1__1_), .S(npu_inst_pe_1_7_4_n4), .Z(
        npu_inst_pe_1_7_4_n21) );
  MUX2_X1 npu_inst_pe_1_7_4_U149 ( .A(npu_inst_pe_1_7_4_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_7_4_int_q_reg_h_3__1_), .S(npu_inst_pe_1_7_4_n4), .Z(
        npu_inst_pe_1_7_4_n20) );
  MUX2_X1 npu_inst_pe_1_7_4_U148 ( .A(npu_inst_pe_1_7_4_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_7_4_int_q_reg_h_5__1_), .S(npu_inst_pe_1_7_4_n4), .Z(
        npu_inst_pe_1_7_4_n19) );
  MUX2_X1 npu_inst_pe_1_7_4_U147 ( .A(npu_inst_pe_1_7_4_n18), .B(
        npu_inst_pe_1_7_4_n15), .S(npu_inst_pe_1_7_4_n8), .Z(
        npu_inst_int_data_x_7__4__0_) );
  MUX2_X1 npu_inst_pe_1_7_4_U146 ( .A(npu_inst_pe_1_7_4_n17), .B(
        npu_inst_pe_1_7_4_n16), .S(npu_inst_pe_1_7_4_n6), .Z(
        npu_inst_pe_1_7_4_n18) );
  MUX2_X1 npu_inst_pe_1_7_4_U145 ( .A(npu_inst_pe_1_7_4_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_7_4_int_q_reg_h_1__0_), .S(npu_inst_pe_1_7_4_n4), .Z(
        npu_inst_pe_1_7_4_n17) );
  MUX2_X1 npu_inst_pe_1_7_4_U144 ( .A(npu_inst_pe_1_7_4_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_7_4_int_q_reg_h_3__0_), .S(npu_inst_pe_1_7_4_n4), .Z(
        npu_inst_pe_1_7_4_n16) );
  MUX2_X1 npu_inst_pe_1_7_4_U143 ( .A(npu_inst_pe_1_7_4_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_7_4_int_q_reg_h_5__0_), .S(npu_inst_pe_1_7_4_n4), .Z(
        npu_inst_pe_1_7_4_n15) );
  XOR2_X1 npu_inst_pe_1_7_4_U142 ( .A(npu_inst_pe_1_7_4_int_data_0_), .B(
        npu_inst_pe_1_7_4_int_q_acc_0_), .Z(npu_inst_pe_1_7_4_N73) );
  AND2_X1 npu_inst_pe_1_7_4_U141 ( .A1(npu_inst_pe_1_7_4_int_q_acc_0_), .A2(
        npu_inst_pe_1_7_4_int_data_0_), .ZN(npu_inst_pe_1_7_4_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_7_4_U140 ( .A(npu_inst_pe_1_7_4_int_q_acc_0_), .B(
        npu_inst_pe_1_7_4_n13), .ZN(npu_inst_pe_1_7_4_N65) );
  OR2_X1 npu_inst_pe_1_7_4_U139 ( .A1(npu_inst_pe_1_7_4_n13), .A2(
        npu_inst_pe_1_7_4_int_q_acc_0_), .ZN(npu_inst_pe_1_7_4_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_7_4_U138 ( .A(npu_inst_pe_1_7_4_int_q_acc_2_), .B(
        npu_inst_pe_1_7_4_add_69_carry_2_), .Z(npu_inst_pe_1_7_4_N75) );
  AND2_X1 npu_inst_pe_1_7_4_U137 ( .A1(npu_inst_pe_1_7_4_add_69_carry_2_), 
        .A2(npu_inst_pe_1_7_4_int_q_acc_2_), .ZN(
        npu_inst_pe_1_7_4_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_7_4_U136 ( .A(npu_inst_pe_1_7_4_int_q_acc_3_), .B(
        npu_inst_pe_1_7_4_add_69_carry_3_), .Z(npu_inst_pe_1_7_4_N76) );
  AND2_X1 npu_inst_pe_1_7_4_U135 ( .A1(npu_inst_pe_1_7_4_add_69_carry_3_), 
        .A2(npu_inst_pe_1_7_4_int_q_acc_3_), .ZN(
        npu_inst_pe_1_7_4_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_7_4_U134 ( .A(npu_inst_pe_1_7_4_int_q_acc_4_), .B(
        npu_inst_pe_1_7_4_add_69_carry_4_), .Z(npu_inst_pe_1_7_4_N77) );
  AND2_X1 npu_inst_pe_1_7_4_U133 ( .A1(npu_inst_pe_1_7_4_add_69_carry_4_), 
        .A2(npu_inst_pe_1_7_4_int_q_acc_4_), .ZN(
        npu_inst_pe_1_7_4_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_7_4_U132 ( .A(npu_inst_pe_1_7_4_int_q_acc_5_), .B(
        npu_inst_pe_1_7_4_add_69_carry_5_), .Z(npu_inst_pe_1_7_4_N78) );
  AND2_X1 npu_inst_pe_1_7_4_U131 ( .A1(npu_inst_pe_1_7_4_add_69_carry_5_), 
        .A2(npu_inst_pe_1_7_4_int_q_acc_5_), .ZN(
        npu_inst_pe_1_7_4_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_7_4_U130 ( .A(npu_inst_pe_1_7_4_int_q_acc_6_), .B(
        npu_inst_pe_1_7_4_add_69_carry_6_), .Z(npu_inst_pe_1_7_4_N79) );
  AND2_X1 npu_inst_pe_1_7_4_U129 ( .A1(npu_inst_pe_1_7_4_add_69_carry_6_), 
        .A2(npu_inst_pe_1_7_4_int_q_acc_6_), .ZN(
        npu_inst_pe_1_7_4_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_7_4_U128 ( .A(npu_inst_pe_1_7_4_int_q_acc_7_), .B(
        npu_inst_pe_1_7_4_add_69_carry_7_), .Z(npu_inst_pe_1_7_4_N80) );
  XNOR2_X1 npu_inst_pe_1_7_4_U127 ( .A(npu_inst_pe_1_7_4_sub_67_carry_2_), .B(
        npu_inst_pe_1_7_4_int_q_acc_2_), .ZN(npu_inst_pe_1_7_4_N67) );
  OR2_X1 npu_inst_pe_1_7_4_U126 ( .A1(npu_inst_pe_1_7_4_int_q_acc_2_), .A2(
        npu_inst_pe_1_7_4_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_7_4_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_7_4_U125 ( .A(npu_inst_pe_1_7_4_sub_67_carry_3_), .B(
        npu_inst_pe_1_7_4_int_q_acc_3_), .ZN(npu_inst_pe_1_7_4_N68) );
  OR2_X1 npu_inst_pe_1_7_4_U124 ( .A1(npu_inst_pe_1_7_4_int_q_acc_3_), .A2(
        npu_inst_pe_1_7_4_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_7_4_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_7_4_U123 ( .A(npu_inst_pe_1_7_4_sub_67_carry_4_), .B(
        npu_inst_pe_1_7_4_int_q_acc_4_), .ZN(npu_inst_pe_1_7_4_N69) );
  OR2_X1 npu_inst_pe_1_7_4_U122 ( .A1(npu_inst_pe_1_7_4_int_q_acc_4_), .A2(
        npu_inst_pe_1_7_4_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_7_4_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_7_4_U121 ( .A(npu_inst_pe_1_7_4_sub_67_carry_5_), .B(
        npu_inst_pe_1_7_4_int_q_acc_5_), .ZN(npu_inst_pe_1_7_4_N70) );
  OR2_X1 npu_inst_pe_1_7_4_U120 ( .A1(npu_inst_pe_1_7_4_int_q_acc_5_), .A2(
        npu_inst_pe_1_7_4_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_7_4_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_7_4_U119 ( .A(npu_inst_pe_1_7_4_sub_67_carry_6_), .B(
        npu_inst_pe_1_7_4_int_q_acc_6_), .ZN(npu_inst_pe_1_7_4_N71) );
  OR2_X1 npu_inst_pe_1_7_4_U118 ( .A1(npu_inst_pe_1_7_4_int_q_acc_6_), .A2(
        npu_inst_pe_1_7_4_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_7_4_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_7_4_U117 ( .A(npu_inst_pe_1_7_4_int_q_acc_7_), .B(
        npu_inst_pe_1_7_4_sub_67_carry_7_), .ZN(npu_inst_pe_1_7_4_N72) );
  INV_X1 npu_inst_pe_1_7_4_U116 ( .A(npu_inst_n75), .ZN(npu_inst_pe_1_7_4_n7)
         );
  INV_X1 npu_inst_pe_1_7_4_U115 ( .A(npu_inst_pe_1_7_4_n7), .ZN(
        npu_inst_pe_1_7_4_n6) );
  INV_X1 npu_inst_pe_1_7_4_U114 ( .A(npu_inst_n52), .ZN(npu_inst_pe_1_7_4_n3)
         );
  AOI22_X1 npu_inst_pe_1_7_4_U113 ( .A1(npu_inst_pe_1_7_4_n38), .A2(
        int_i_data_v_npu[7]), .B1(npu_inst_pe_1_7_4_n114), .B2(
        npu_inst_pe_1_7_4_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_7_4_n39) );
  INV_X1 npu_inst_pe_1_7_4_U112 ( .A(npu_inst_pe_1_7_4_n39), .ZN(
        npu_inst_pe_1_7_4_n112) );
  AOI22_X1 npu_inst_pe_1_7_4_U111 ( .A1(npu_inst_pe_1_7_4_n38), .A2(
        int_i_data_v_npu[6]), .B1(npu_inst_pe_1_7_4_n114), .B2(
        npu_inst_pe_1_7_4_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_7_4_n37) );
  INV_X1 npu_inst_pe_1_7_4_U110 ( .A(npu_inst_pe_1_7_4_n37), .ZN(
        npu_inst_pe_1_7_4_n113) );
  AOI22_X1 npu_inst_pe_1_7_4_U107 ( .A1(int_i_data_v_npu[7]), .A2(
        npu_inst_pe_1_7_4_n58), .B1(npu_inst_pe_1_7_4_n119), .B2(
        npu_inst_pe_1_7_4_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_7_4_n59) );
  INV_X1 npu_inst_pe_1_7_4_U106 ( .A(npu_inst_pe_1_7_4_n59), .ZN(
        npu_inst_pe_1_7_4_n102) );
  AOI22_X1 npu_inst_pe_1_7_4_U105 ( .A1(int_i_data_v_npu[6]), .A2(
        npu_inst_pe_1_7_4_n58), .B1(npu_inst_pe_1_7_4_n119), .B2(
        npu_inst_pe_1_7_4_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_7_4_n57) );
  INV_X1 npu_inst_pe_1_7_4_U104 ( .A(npu_inst_pe_1_7_4_n57), .ZN(
        npu_inst_pe_1_7_4_n103) );
  AOI22_X1 npu_inst_pe_1_7_4_U103 ( .A1(int_i_data_v_npu[7]), .A2(
        npu_inst_pe_1_7_4_n54), .B1(npu_inst_pe_1_7_4_n118), .B2(
        npu_inst_pe_1_7_4_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_7_4_n55) );
  INV_X1 npu_inst_pe_1_7_4_U102 ( .A(npu_inst_pe_1_7_4_n55), .ZN(
        npu_inst_pe_1_7_4_n104) );
  AOI22_X1 npu_inst_pe_1_7_4_U101 ( .A1(int_i_data_v_npu[6]), .A2(
        npu_inst_pe_1_7_4_n54), .B1(npu_inst_pe_1_7_4_n118), .B2(
        npu_inst_pe_1_7_4_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_7_4_n53) );
  INV_X1 npu_inst_pe_1_7_4_U100 ( .A(npu_inst_pe_1_7_4_n53), .ZN(
        npu_inst_pe_1_7_4_n105) );
  AOI22_X1 npu_inst_pe_1_7_4_U99 ( .A1(int_i_data_v_npu[7]), .A2(
        npu_inst_pe_1_7_4_n50), .B1(npu_inst_pe_1_7_4_n117), .B2(
        npu_inst_pe_1_7_4_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_7_4_n51) );
  INV_X1 npu_inst_pe_1_7_4_U98 ( .A(npu_inst_pe_1_7_4_n51), .ZN(
        npu_inst_pe_1_7_4_n106) );
  AOI22_X1 npu_inst_pe_1_7_4_U97 ( .A1(int_i_data_v_npu[6]), .A2(
        npu_inst_pe_1_7_4_n50), .B1(npu_inst_pe_1_7_4_n117), .B2(
        npu_inst_pe_1_7_4_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_7_4_n49) );
  INV_X1 npu_inst_pe_1_7_4_U96 ( .A(npu_inst_pe_1_7_4_n49), .ZN(
        npu_inst_pe_1_7_4_n107) );
  AOI22_X1 npu_inst_pe_1_7_4_U95 ( .A1(int_i_data_v_npu[7]), .A2(
        npu_inst_pe_1_7_4_n46), .B1(npu_inst_pe_1_7_4_n116), .B2(
        npu_inst_pe_1_7_4_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_7_4_n47) );
  INV_X1 npu_inst_pe_1_7_4_U94 ( .A(npu_inst_pe_1_7_4_n47), .ZN(
        npu_inst_pe_1_7_4_n108) );
  AOI22_X1 npu_inst_pe_1_7_4_U93 ( .A1(int_i_data_v_npu[6]), .A2(
        npu_inst_pe_1_7_4_n46), .B1(npu_inst_pe_1_7_4_n116), .B2(
        npu_inst_pe_1_7_4_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_7_4_n45) );
  INV_X1 npu_inst_pe_1_7_4_U92 ( .A(npu_inst_pe_1_7_4_n45), .ZN(
        npu_inst_pe_1_7_4_n109) );
  AOI22_X1 npu_inst_pe_1_7_4_U91 ( .A1(int_i_data_v_npu[7]), .A2(
        npu_inst_pe_1_7_4_n42), .B1(npu_inst_pe_1_7_4_n115), .B2(
        npu_inst_pe_1_7_4_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_7_4_n43) );
  INV_X1 npu_inst_pe_1_7_4_U90 ( .A(npu_inst_pe_1_7_4_n43), .ZN(
        npu_inst_pe_1_7_4_n110) );
  AOI22_X1 npu_inst_pe_1_7_4_U89 ( .A1(int_i_data_v_npu[6]), .A2(
        npu_inst_pe_1_7_4_n42), .B1(npu_inst_pe_1_7_4_n115), .B2(
        npu_inst_pe_1_7_4_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_7_4_n41) );
  INV_X1 npu_inst_pe_1_7_4_U88 ( .A(npu_inst_pe_1_7_4_n41), .ZN(
        npu_inst_pe_1_7_4_n111) );
  NAND2_X1 npu_inst_pe_1_7_4_U87 ( .A1(npu_inst_pe_1_7_4_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_7_4_n60), .ZN(npu_inst_pe_1_7_4_n74) );
  OAI21_X1 npu_inst_pe_1_7_4_U86 ( .B1(npu_inst_pe_1_7_4_n63), .B2(
        npu_inst_pe_1_7_4_n60), .A(npu_inst_pe_1_7_4_n74), .ZN(
        npu_inst_pe_1_7_4_n97) );
  NAND2_X1 npu_inst_pe_1_7_4_U85 ( .A1(npu_inst_pe_1_7_4_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_7_4_n60), .ZN(npu_inst_pe_1_7_4_n73) );
  OAI21_X1 npu_inst_pe_1_7_4_U84 ( .B1(npu_inst_pe_1_7_4_n61), .B2(
        npu_inst_pe_1_7_4_n60), .A(npu_inst_pe_1_7_4_n73), .ZN(
        npu_inst_pe_1_7_4_n96) );
  NAND2_X1 npu_inst_pe_1_7_4_U83 ( .A1(npu_inst_pe_1_7_4_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_7_4_n56), .ZN(npu_inst_pe_1_7_4_n72) );
  OAI21_X1 npu_inst_pe_1_7_4_U82 ( .B1(npu_inst_pe_1_7_4_n63), .B2(
        npu_inst_pe_1_7_4_n56), .A(npu_inst_pe_1_7_4_n72), .ZN(
        npu_inst_pe_1_7_4_n95) );
  NAND2_X1 npu_inst_pe_1_7_4_U81 ( .A1(npu_inst_pe_1_7_4_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_7_4_n56), .ZN(npu_inst_pe_1_7_4_n71) );
  OAI21_X1 npu_inst_pe_1_7_4_U80 ( .B1(npu_inst_pe_1_7_4_n61), .B2(
        npu_inst_pe_1_7_4_n56), .A(npu_inst_pe_1_7_4_n71), .ZN(
        npu_inst_pe_1_7_4_n94) );
  NAND2_X1 npu_inst_pe_1_7_4_U79 ( .A1(npu_inst_pe_1_7_4_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_7_4_n52), .ZN(npu_inst_pe_1_7_4_n70) );
  OAI21_X1 npu_inst_pe_1_7_4_U78 ( .B1(npu_inst_pe_1_7_4_n63), .B2(
        npu_inst_pe_1_7_4_n52), .A(npu_inst_pe_1_7_4_n70), .ZN(
        npu_inst_pe_1_7_4_n93) );
  NAND2_X1 npu_inst_pe_1_7_4_U77 ( .A1(npu_inst_pe_1_7_4_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_7_4_n52), .ZN(npu_inst_pe_1_7_4_n69) );
  OAI21_X1 npu_inst_pe_1_7_4_U76 ( .B1(npu_inst_pe_1_7_4_n61), .B2(
        npu_inst_pe_1_7_4_n52), .A(npu_inst_pe_1_7_4_n69), .ZN(
        npu_inst_pe_1_7_4_n92) );
  NAND2_X1 npu_inst_pe_1_7_4_U75 ( .A1(npu_inst_pe_1_7_4_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_7_4_n48), .ZN(npu_inst_pe_1_7_4_n68) );
  OAI21_X1 npu_inst_pe_1_7_4_U74 ( .B1(npu_inst_pe_1_7_4_n63), .B2(
        npu_inst_pe_1_7_4_n48), .A(npu_inst_pe_1_7_4_n68), .ZN(
        npu_inst_pe_1_7_4_n91) );
  NAND2_X1 npu_inst_pe_1_7_4_U73 ( .A1(npu_inst_pe_1_7_4_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_7_4_n48), .ZN(npu_inst_pe_1_7_4_n67) );
  OAI21_X1 npu_inst_pe_1_7_4_U72 ( .B1(npu_inst_pe_1_7_4_n61), .B2(
        npu_inst_pe_1_7_4_n48), .A(npu_inst_pe_1_7_4_n67), .ZN(
        npu_inst_pe_1_7_4_n90) );
  NAND2_X1 npu_inst_pe_1_7_4_U71 ( .A1(npu_inst_pe_1_7_4_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_7_4_n44), .ZN(npu_inst_pe_1_7_4_n66) );
  OAI21_X1 npu_inst_pe_1_7_4_U70 ( .B1(npu_inst_pe_1_7_4_n63), .B2(
        npu_inst_pe_1_7_4_n44), .A(npu_inst_pe_1_7_4_n66), .ZN(
        npu_inst_pe_1_7_4_n89) );
  NAND2_X1 npu_inst_pe_1_7_4_U69 ( .A1(npu_inst_pe_1_7_4_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_7_4_n44), .ZN(npu_inst_pe_1_7_4_n65) );
  OAI21_X1 npu_inst_pe_1_7_4_U68 ( .B1(npu_inst_pe_1_7_4_n61), .B2(
        npu_inst_pe_1_7_4_n44), .A(npu_inst_pe_1_7_4_n65), .ZN(
        npu_inst_pe_1_7_4_n88) );
  NAND2_X1 npu_inst_pe_1_7_4_U67 ( .A1(npu_inst_pe_1_7_4_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_7_4_n40), .ZN(npu_inst_pe_1_7_4_n64) );
  OAI21_X1 npu_inst_pe_1_7_4_U66 ( .B1(npu_inst_pe_1_7_4_n63), .B2(
        npu_inst_pe_1_7_4_n40), .A(npu_inst_pe_1_7_4_n64), .ZN(
        npu_inst_pe_1_7_4_n87) );
  NAND2_X1 npu_inst_pe_1_7_4_U65 ( .A1(npu_inst_pe_1_7_4_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_7_4_n40), .ZN(npu_inst_pe_1_7_4_n62) );
  OAI21_X1 npu_inst_pe_1_7_4_U64 ( .B1(npu_inst_pe_1_7_4_n61), .B2(
        npu_inst_pe_1_7_4_n40), .A(npu_inst_pe_1_7_4_n62), .ZN(
        npu_inst_pe_1_7_4_n86) );
  AND2_X1 npu_inst_pe_1_7_4_U63 ( .A1(npu_inst_pe_1_7_4_N93), .A2(npu_inst_n52), .ZN(npu_inst_int_data_y_7__4__0_) );
  AND2_X1 npu_inst_pe_1_7_4_U62 ( .A1(npu_inst_n52), .A2(npu_inst_pe_1_7_4_N94), .ZN(npu_inst_int_data_y_7__4__1_) );
  AOI22_X1 npu_inst_pe_1_7_4_U61 ( .A1(npu_inst_n52), .A2(int_i_data_v_npu[7]), 
        .B1(npu_inst_pe_1_7_4_n3), .B2(npu_inst_int_data_x_7__5__1_), .ZN(
        npu_inst_pe_1_7_4_n63) );
  AOI22_X1 npu_inst_pe_1_7_4_U60 ( .A1(npu_inst_n52), .A2(int_i_data_v_npu[6]), 
        .B1(npu_inst_pe_1_7_4_n3), .B2(npu_inst_int_data_x_7__5__0_), .ZN(
        npu_inst_pe_1_7_4_n61) );
  AOI222_X1 npu_inst_pe_1_7_4_U59 ( .A1(1'b0), .A2(npu_inst_pe_1_7_4_n1), .B1(
        npu_inst_pe_1_7_4_N73), .B2(npu_inst_pe_1_7_4_n76), .C1(
        npu_inst_pe_1_7_4_N65), .C2(npu_inst_pe_1_7_4_n77), .ZN(
        npu_inst_pe_1_7_4_n84) );
  INV_X1 npu_inst_pe_1_7_4_U58 ( .A(npu_inst_pe_1_7_4_n84), .ZN(
        npu_inst_pe_1_7_4_n101) );
  AOI222_X1 npu_inst_pe_1_7_4_U57 ( .A1(1'b0), .A2(npu_inst_pe_1_7_4_n1), .B1(
        npu_inst_pe_1_7_4_N80), .B2(npu_inst_pe_1_7_4_n76), .C1(
        npu_inst_pe_1_7_4_N72), .C2(npu_inst_pe_1_7_4_n77), .ZN(
        npu_inst_pe_1_7_4_n75) );
  INV_X1 npu_inst_pe_1_7_4_U56 ( .A(npu_inst_pe_1_7_4_n75), .ZN(
        npu_inst_pe_1_7_4_n33) );
  AOI222_X1 npu_inst_pe_1_7_4_U55 ( .A1(1'b0), .A2(npu_inst_pe_1_7_4_n1), .B1(
        npu_inst_pe_1_7_4_N74), .B2(npu_inst_pe_1_7_4_n76), .C1(
        npu_inst_pe_1_7_4_N66), .C2(npu_inst_pe_1_7_4_n77), .ZN(
        npu_inst_pe_1_7_4_n83) );
  INV_X1 npu_inst_pe_1_7_4_U54 ( .A(npu_inst_pe_1_7_4_n83), .ZN(
        npu_inst_pe_1_7_4_n100) );
  AOI222_X1 npu_inst_pe_1_7_4_U53 ( .A1(1'b0), .A2(npu_inst_pe_1_7_4_n1), .B1(
        npu_inst_pe_1_7_4_N75), .B2(npu_inst_pe_1_7_4_n76), .C1(
        npu_inst_pe_1_7_4_N67), .C2(npu_inst_pe_1_7_4_n77), .ZN(
        npu_inst_pe_1_7_4_n82) );
  INV_X1 npu_inst_pe_1_7_4_U52 ( .A(npu_inst_pe_1_7_4_n82), .ZN(
        npu_inst_pe_1_7_4_n99) );
  AOI222_X1 npu_inst_pe_1_7_4_U51 ( .A1(1'b0), .A2(npu_inst_pe_1_7_4_n1), .B1(
        npu_inst_pe_1_7_4_N76), .B2(npu_inst_pe_1_7_4_n76), .C1(
        npu_inst_pe_1_7_4_N68), .C2(npu_inst_pe_1_7_4_n77), .ZN(
        npu_inst_pe_1_7_4_n81) );
  INV_X1 npu_inst_pe_1_7_4_U50 ( .A(npu_inst_pe_1_7_4_n81), .ZN(
        npu_inst_pe_1_7_4_n98) );
  AOI222_X1 npu_inst_pe_1_7_4_U49 ( .A1(1'b0), .A2(npu_inst_pe_1_7_4_n1), .B1(
        npu_inst_pe_1_7_4_N77), .B2(npu_inst_pe_1_7_4_n76), .C1(
        npu_inst_pe_1_7_4_N69), .C2(npu_inst_pe_1_7_4_n77), .ZN(
        npu_inst_pe_1_7_4_n80) );
  INV_X1 npu_inst_pe_1_7_4_U48 ( .A(npu_inst_pe_1_7_4_n80), .ZN(
        npu_inst_pe_1_7_4_n36) );
  AOI222_X1 npu_inst_pe_1_7_4_U47 ( .A1(1'b0), .A2(npu_inst_pe_1_7_4_n1), .B1(
        npu_inst_pe_1_7_4_N78), .B2(npu_inst_pe_1_7_4_n76), .C1(
        npu_inst_pe_1_7_4_N70), .C2(npu_inst_pe_1_7_4_n77), .ZN(
        npu_inst_pe_1_7_4_n79) );
  INV_X1 npu_inst_pe_1_7_4_U46 ( .A(npu_inst_pe_1_7_4_n79), .ZN(
        npu_inst_pe_1_7_4_n35) );
  AOI222_X1 npu_inst_pe_1_7_4_U45 ( .A1(1'b0), .A2(npu_inst_pe_1_7_4_n1), .B1(
        npu_inst_pe_1_7_4_N79), .B2(npu_inst_pe_1_7_4_n76), .C1(
        npu_inst_pe_1_7_4_N71), .C2(npu_inst_pe_1_7_4_n77), .ZN(
        npu_inst_pe_1_7_4_n78) );
  INV_X1 npu_inst_pe_1_7_4_U44 ( .A(npu_inst_pe_1_7_4_n78), .ZN(
        npu_inst_pe_1_7_4_n34) );
  AND2_X1 npu_inst_pe_1_7_4_U43 ( .A1(npu_inst_pe_1_7_4_int_q_acc_0_), .A2(
        npu_inst_pe_1_7_4_n1), .ZN(npu_inst_int_data_res_7__4__0_) );
  AND2_X1 npu_inst_pe_1_7_4_U42 ( .A1(npu_inst_pe_1_7_4_n2), .A2(
        npu_inst_pe_1_7_4_int_q_acc_7_), .ZN(npu_inst_int_data_res_7__4__7_)
         );
  AND2_X1 npu_inst_pe_1_7_4_U41 ( .A1(npu_inst_pe_1_7_4_int_q_acc_1_), .A2(
        npu_inst_pe_1_7_4_n1), .ZN(npu_inst_int_data_res_7__4__1_) );
  AND2_X1 npu_inst_pe_1_7_4_U40 ( .A1(npu_inst_pe_1_7_4_int_q_acc_2_), .A2(
        npu_inst_pe_1_7_4_n1), .ZN(npu_inst_int_data_res_7__4__2_) );
  AND2_X1 npu_inst_pe_1_7_4_U39 ( .A1(npu_inst_pe_1_7_4_int_q_acc_3_), .A2(
        npu_inst_pe_1_7_4_n2), .ZN(npu_inst_int_data_res_7__4__3_) );
  AND2_X1 npu_inst_pe_1_7_4_U38 ( .A1(npu_inst_pe_1_7_4_int_q_acc_4_), .A2(
        npu_inst_pe_1_7_4_n2), .ZN(npu_inst_int_data_res_7__4__4_) );
  AND2_X1 npu_inst_pe_1_7_4_U37 ( .A1(npu_inst_pe_1_7_4_int_q_acc_5_), .A2(
        npu_inst_pe_1_7_4_n2), .ZN(npu_inst_int_data_res_7__4__5_) );
  AND2_X1 npu_inst_pe_1_7_4_U36 ( .A1(npu_inst_pe_1_7_4_int_q_acc_6_), .A2(
        npu_inst_pe_1_7_4_n2), .ZN(npu_inst_int_data_res_7__4__6_) );
  INV_X1 npu_inst_pe_1_7_4_U35 ( .A(npu_inst_pe_1_7_4_int_data_1_), .ZN(
        npu_inst_pe_1_7_4_n14) );
  NOR3_X1 npu_inst_pe_1_7_4_U34 ( .A1(npu_inst_pe_1_7_4_n26), .A2(npu_inst_n52), .A3(npu_inst_int_ckg[3]), .ZN(npu_inst_pe_1_7_4_n85) );
  OR2_X1 npu_inst_pe_1_7_4_U33 ( .A1(npu_inst_pe_1_7_4_n85), .A2(
        npu_inst_pe_1_7_4_n2), .ZN(npu_inst_pe_1_7_4_N84) );
  AND2_X1 npu_inst_pe_1_7_4_U32 ( .A1(npu_inst_int_data_x_7__4__1_), .A2(
        npu_inst_pe_1_7_4_int_q_weight_1_), .ZN(npu_inst_pe_1_7_4_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_7_4_U31 ( .A1(npu_inst_int_data_x_7__4__0_), .A2(
        npu_inst_pe_1_7_4_int_q_weight_1_), .ZN(npu_inst_pe_1_7_4_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_7_4_U30 ( .A(npu_inst_pe_1_7_4_int_data_0_), .ZN(
        npu_inst_pe_1_7_4_n13) );
  INV_X1 npu_inst_pe_1_7_4_U29 ( .A(npu_inst_n67), .ZN(npu_inst_pe_1_7_4_n5)
         );
  OR3_X1 npu_inst_pe_1_7_4_U28 ( .A1(npu_inst_pe_1_7_4_n6), .A2(
        npu_inst_pe_1_7_4_n8), .A3(npu_inst_pe_1_7_4_n5), .ZN(
        npu_inst_pe_1_7_4_n56) );
  OR3_X1 npu_inst_pe_1_7_4_U27 ( .A1(npu_inst_pe_1_7_4_n5), .A2(
        npu_inst_pe_1_7_4_n8), .A3(npu_inst_pe_1_7_4_n7), .ZN(
        npu_inst_pe_1_7_4_n48) );
  INV_X1 npu_inst_pe_1_7_4_U26 ( .A(npu_inst_pe_1_7_4_n5), .ZN(
        npu_inst_pe_1_7_4_n4) );
  OR3_X1 npu_inst_pe_1_7_4_U25 ( .A1(npu_inst_pe_1_7_4_n4), .A2(
        npu_inst_pe_1_7_4_n8), .A3(npu_inst_pe_1_7_4_n7), .ZN(
        npu_inst_pe_1_7_4_n52) );
  OR3_X1 npu_inst_pe_1_7_4_U24 ( .A1(npu_inst_pe_1_7_4_n6), .A2(
        npu_inst_pe_1_7_4_n8), .A3(npu_inst_pe_1_7_4_n4), .ZN(
        npu_inst_pe_1_7_4_n60) );
  NOR2_X1 npu_inst_pe_1_7_4_U23 ( .A1(npu_inst_pe_1_7_4_n60), .A2(
        npu_inst_pe_1_7_4_n3), .ZN(npu_inst_pe_1_7_4_n58) );
  NOR2_X1 npu_inst_pe_1_7_4_U22 ( .A1(npu_inst_pe_1_7_4_n56), .A2(
        npu_inst_pe_1_7_4_n3), .ZN(npu_inst_pe_1_7_4_n54) );
  NOR2_X1 npu_inst_pe_1_7_4_U21 ( .A1(npu_inst_pe_1_7_4_n52), .A2(
        npu_inst_pe_1_7_4_n3), .ZN(npu_inst_pe_1_7_4_n50) );
  NOR2_X1 npu_inst_pe_1_7_4_U20 ( .A1(npu_inst_pe_1_7_4_n48), .A2(
        npu_inst_pe_1_7_4_n3), .ZN(npu_inst_pe_1_7_4_n46) );
  NOR2_X1 npu_inst_pe_1_7_4_U19 ( .A1(npu_inst_pe_1_7_4_n40), .A2(
        npu_inst_pe_1_7_4_n3), .ZN(npu_inst_pe_1_7_4_n38) );
  NOR2_X1 npu_inst_pe_1_7_4_U18 ( .A1(npu_inst_pe_1_7_4_n44), .A2(
        npu_inst_pe_1_7_4_n3), .ZN(npu_inst_pe_1_7_4_n42) );
  BUF_X1 npu_inst_pe_1_7_4_U17 ( .A(npu_inst_n92), .Z(npu_inst_pe_1_7_4_n8) );
  INV_X1 npu_inst_pe_1_7_4_U16 ( .A(npu_inst_n122), .ZN(npu_inst_pe_1_7_4_n12)
         );
  INV_X1 npu_inst_pe_1_7_4_U15 ( .A(npu_inst_pe_1_7_4_n38), .ZN(
        npu_inst_pe_1_7_4_n114) );
  INV_X1 npu_inst_pe_1_7_4_U14 ( .A(npu_inst_pe_1_7_4_n58), .ZN(
        npu_inst_pe_1_7_4_n119) );
  INV_X1 npu_inst_pe_1_7_4_U13 ( .A(npu_inst_pe_1_7_4_n54), .ZN(
        npu_inst_pe_1_7_4_n118) );
  INV_X1 npu_inst_pe_1_7_4_U12 ( .A(npu_inst_pe_1_7_4_n50), .ZN(
        npu_inst_pe_1_7_4_n117) );
  INV_X1 npu_inst_pe_1_7_4_U11 ( .A(npu_inst_pe_1_7_4_n46), .ZN(
        npu_inst_pe_1_7_4_n116) );
  INV_X1 npu_inst_pe_1_7_4_U10 ( .A(npu_inst_pe_1_7_4_n42), .ZN(
        npu_inst_pe_1_7_4_n115) );
  BUF_X1 npu_inst_pe_1_7_4_U9 ( .A(npu_inst_n8), .Z(npu_inst_pe_1_7_4_n2) );
  BUF_X1 npu_inst_pe_1_7_4_U8 ( .A(npu_inst_n8), .Z(npu_inst_pe_1_7_4_n1) );
  BUF_X1 npu_inst_pe_1_7_4_U7 ( .A(npu_inst_pe_1_7_4_n12), .Z(
        npu_inst_pe_1_7_4_n11) );
  BUF_X1 npu_inst_pe_1_7_4_U6 ( .A(npu_inst_pe_1_7_4_n12), .Z(
        npu_inst_pe_1_7_4_n10) );
  BUF_X1 npu_inst_pe_1_7_4_U5 ( .A(npu_inst_pe_1_7_4_n12), .Z(
        npu_inst_pe_1_7_4_n9) );
  NOR2_X1 npu_inst_pe_1_7_4_U4 ( .A1(npu_inst_pe_1_7_4_int_q_weight_0_), .A2(
        npu_inst_pe_1_7_4_n1), .ZN(npu_inst_pe_1_7_4_n76) );
  NOR2_X1 npu_inst_pe_1_7_4_U3 ( .A1(npu_inst_pe_1_7_4_n27), .A2(
        npu_inst_pe_1_7_4_n1), .ZN(npu_inst_pe_1_7_4_n77) );
  FA_X1 npu_inst_pe_1_7_4_sub_67_U2_1 ( .A(npu_inst_pe_1_7_4_int_q_acc_1_), 
        .B(npu_inst_pe_1_7_4_n14), .CI(npu_inst_pe_1_7_4_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_7_4_sub_67_carry_2_), .S(npu_inst_pe_1_7_4_N66) );
  FA_X1 npu_inst_pe_1_7_4_add_69_U1_1 ( .A(npu_inst_pe_1_7_4_int_q_acc_1_), 
        .B(npu_inst_pe_1_7_4_int_data_1_), .CI(
        npu_inst_pe_1_7_4_add_69_carry_1_), .CO(
        npu_inst_pe_1_7_4_add_69_carry_2_), .S(npu_inst_pe_1_7_4_N74) );
  NAND3_X1 npu_inst_pe_1_7_4_U109 ( .A1(npu_inst_pe_1_7_4_n5), .A2(
        npu_inst_pe_1_7_4_n7), .A3(npu_inst_pe_1_7_4_n8), .ZN(
        npu_inst_pe_1_7_4_n44) );
  NAND3_X1 npu_inst_pe_1_7_4_U108 ( .A1(npu_inst_pe_1_7_4_n4), .A2(
        npu_inst_pe_1_7_4_n7), .A3(npu_inst_pe_1_7_4_n8), .ZN(
        npu_inst_pe_1_7_4_n40) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_7_4_n34), .CK(
        npu_inst_pe_1_7_4_net3182), .RN(npu_inst_pe_1_7_4_n9), .Q(
        npu_inst_pe_1_7_4_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_7_4_n35), .CK(
        npu_inst_pe_1_7_4_net3182), .RN(npu_inst_pe_1_7_4_n9), .Q(
        npu_inst_pe_1_7_4_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_7_4_n36), .CK(
        npu_inst_pe_1_7_4_net3182), .RN(npu_inst_pe_1_7_4_n9), .Q(
        npu_inst_pe_1_7_4_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_7_4_n98), .CK(
        npu_inst_pe_1_7_4_net3182), .RN(npu_inst_pe_1_7_4_n9), .Q(
        npu_inst_pe_1_7_4_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_7_4_n99), .CK(
        npu_inst_pe_1_7_4_net3182), .RN(npu_inst_pe_1_7_4_n9), .Q(
        npu_inst_pe_1_7_4_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_7_4_n100), 
        .CK(npu_inst_pe_1_7_4_net3182), .RN(npu_inst_pe_1_7_4_n9), .Q(
        npu_inst_pe_1_7_4_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_7_4_n33), .CK(
        npu_inst_pe_1_7_4_net3182), .RN(npu_inst_pe_1_7_4_n9), .Q(
        npu_inst_pe_1_7_4_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_7_4_n101), 
        .CK(npu_inst_pe_1_7_4_net3182), .RN(npu_inst_pe_1_7_4_n9), .Q(
        npu_inst_pe_1_7_4_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_weight_reg_0_ ( .D(npu_inst_n108), .CK(
        npu_inst_pe_1_7_4_net3188), .RN(npu_inst_pe_1_7_4_n9), .Q(
        npu_inst_pe_1_7_4_int_q_weight_0_), .QN(npu_inst_pe_1_7_4_n27) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_weight_reg_1_ ( .D(npu_inst_n114), .CK(
        npu_inst_pe_1_7_4_net3188), .RN(npu_inst_pe_1_7_4_n9), .Q(
        npu_inst_pe_1_7_4_int_q_weight_1_), .QN(npu_inst_pe_1_7_4_n26) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_7_4_n113), 
        .CK(npu_inst_pe_1_7_4_net3188), .RN(npu_inst_pe_1_7_4_n9), .Q(
        npu_inst_pe_1_7_4_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_7_4_n112), 
        .CK(npu_inst_pe_1_7_4_net3188), .RN(npu_inst_pe_1_7_4_n9), .Q(
        npu_inst_pe_1_7_4_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_7_4_n111), 
        .CK(npu_inst_pe_1_7_4_net3188), .RN(npu_inst_pe_1_7_4_n10), .Q(
        npu_inst_pe_1_7_4_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_7_4_n110), 
        .CK(npu_inst_pe_1_7_4_net3188), .RN(npu_inst_pe_1_7_4_n10), .Q(
        npu_inst_pe_1_7_4_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_7_4_n109), 
        .CK(npu_inst_pe_1_7_4_net3188), .RN(npu_inst_pe_1_7_4_n10), .Q(
        npu_inst_pe_1_7_4_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_7_4_n108), 
        .CK(npu_inst_pe_1_7_4_net3188), .RN(npu_inst_pe_1_7_4_n10), .Q(
        npu_inst_pe_1_7_4_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_7_4_n107), 
        .CK(npu_inst_pe_1_7_4_net3188), .RN(npu_inst_pe_1_7_4_n10), .Q(
        npu_inst_pe_1_7_4_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_7_4_n106), 
        .CK(npu_inst_pe_1_7_4_net3188), .RN(npu_inst_pe_1_7_4_n10), .Q(
        npu_inst_pe_1_7_4_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_7_4_n105), 
        .CK(npu_inst_pe_1_7_4_net3188), .RN(npu_inst_pe_1_7_4_n10), .Q(
        npu_inst_pe_1_7_4_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_7_4_n104), 
        .CK(npu_inst_pe_1_7_4_net3188), .RN(npu_inst_pe_1_7_4_n10), .Q(
        npu_inst_pe_1_7_4_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_7_4_n103), 
        .CK(npu_inst_pe_1_7_4_net3188), .RN(npu_inst_pe_1_7_4_n10), .Q(
        npu_inst_pe_1_7_4_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_7_4_n102), 
        .CK(npu_inst_pe_1_7_4_net3188), .RN(npu_inst_pe_1_7_4_n10), .Q(
        npu_inst_pe_1_7_4_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_7_4_n86), 
        .CK(npu_inst_pe_1_7_4_net3188), .RN(npu_inst_pe_1_7_4_n10), .Q(
        npu_inst_pe_1_7_4_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_7_4_n87), 
        .CK(npu_inst_pe_1_7_4_net3188), .RN(npu_inst_pe_1_7_4_n10), .Q(
        npu_inst_pe_1_7_4_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_7_4_n88), 
        .CK(npu_inst_pe_1_7_4_net3188), .RN(npu_inst_pe_1_7_4_n11), .Q(
        npu_inst_pe_1_7_4_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_7_4_n89), 
        .CK(npu_inst_pe_1_7_4_net3188), .RN(npu_inst_pe_1_7_4_n11), .Q(
        npu_inst_pe_1_7_4_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_7_4_n90), 
        .CK(npu_inst_pe_1_7_4_net3188), .RN(npu_inst_pe_1_7_4_n11), .Q(
        npu_inst_pe_1_7_4_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_7_4_n91), 
        .CK(npu_inst_pe_1_7_4_net3188), .RN(npu_inst_pe_1_7_4_n11), .Q(
        npu_inst_pe_1_7_4_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_7_4_n92), 
        .CK(npu_inst_pe_1_7_4_net3188), .RN(npu_inst_pe_1_7_4_n11), .Q(
        npu_inst_pe_1_7_4_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_7_4_n93), 
        .CK(npu_inst_pe_1_7_4_net3188), .RN(npu_inst_pe_1_7_4_n11), .Q(
        npu_inst_pe_1_7_4_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_7_4_n94), 
        .CK(npu_inst_pe_1_7_4_net3188), .RN(npu_inst_pe_1_7_4_n11), .Q(
        npu_inst_pe_1_7_4_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_7_4_n95), 
        .CK(npu_inst_pe_1_7_4_net3188), .RN(npu_inst_pe_1_7_4_n11), .Q(
        npu_inst_pe_1_7_4_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_7_4_n96), 
        .CK(npu_inst_pe_1_7_4_net3188), .RN(npu_inst_pe_1_7_4_n11), .Q(
        npu_inst_pe_1_7_4_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_7_4_n97), 
        .CK(npu_inst_pe_1_7_4_net3188), .RN(npu_inst_pe_1_7_4_n11), .Q(
        npu_inst_pe_1_7_4_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_7_4_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_7_4_N84), .SE(1'b0), .GCK(npu_inst_pe_1_7_4_net3182) );
  CLKGATETST_X1 npu_inst_pe_1_7_4_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n61), .SE(1'b0), .GCK(npu_inst_pe_1_7_4_net3188) );
  MUX2_X1 npu_inst_pe_1_7_5_U162 ( .A(npu_inst_pe_1_7_5_n32), .B(
        npu_inst_pe_1_7_5_n29), .S(npu_inst_pe_1_7_5_n8), .Z(
        npu_inst_pe_1_7_5_N93) );
  MUX2_X1 npu_inst_pe_1_7_5_U161 ( .A(npu_inst_pe_1_7_5_n31), .B(
        npu_inst_pe_1_7_5_n30), .S(npu_inst_pe_1_7_5_n6), .Z(
        npu_inst_pe_1_7_5_n32) );
  MUX2_X1 npu_inst_pe_1_7_5_U160 ( .A(npu_inst_pe_1_7_5_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_7_5_int_q_reg_v_1__0_), .S(npu_inst_pe_1_7_5_n4), .Z(
        npu_inst_pe_1_7_5_n31) );
  MUX2_X1 npu_inst_pe_1_7_5_U159 ( .A(npu_inst_pe_1_7_5_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_7_5_int_q_reg_v_3__0_), .S(npu_inst_pe_1_7_5_n4), .Z(
        npu_inst_pe_1_7_5_n30) );
  MUX2_X1 npu_inst_pe_1_7_5_U158 ( .A(npu_inst_pe_1_7_5_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_7_5_int_q_reg_v_5__0_), .S(npu_inst_pe_1_7_5_n4), .Z(
        npu_inst_pe_1_7_5_n29) );
  MUX2_X1 npu_inst_pe_1_7_5_U157 ( .A(npu_inst_pe_1_7_5_n28), .B(
        npu_inst_pe_1_7_5_n23), .S(npu_inst_pe_1_7_5_n8), .Z(
        npu_inst_pe_1_7_5_N94) );
  MUX2_X1 npu_inst_pe_1_7_5_U156 ( .A(npu_inst_pe_1_7_5_n25), .B(
        npu_inst_pe_1_7_5_n24), .S(npu_inst_pe_1_7_5_n6), .Z(
        npu_inst_pe_1_7_5_n28) );
  MUX2_X1 npu_inst_pe_1_7_5_U155 ( .A(npu_inst_pe_1_7_5_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_7_5_int_q_reg_v_1__1_), .S(npu_inst_pe_1_7_5_n4), .Z(
        npu_inst_pe_1_7_5_n25) );
  MUX2_X1 npu_inst_pe_1_7_5_U154 ( .A(npu_inst_pe_1_7_5_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_7_5_int_q_reg_v_3__1_), .S(npu_inst_pe_1_7_5_n4), .Z(
        npu_inst_pe_1_7_5_n24) );
  MUX2_X1 npu_inst_pe_1_7_5_U153 ( .A(npu_inst_pe_1_7_5_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_7_5_int_q_reg_v_5__1_), .S(npu_inst_pe_1_7_5_n4), .Z(
        npu_inst_pe_1_7_5_n23) );
  MUX2_X1 npu_inst_pe_1_7_5_U152 ( .A(npu_inst_pe_1_7_5_n22), .B(
        npu_inst_pe_1_7_5_n19), .S(npu_inst_pe_1_7_5_n8), .Z(
        npu_inst_int_data_x_7__5__1_) );
  MUX2_X1 npu_inst_pe_1_7_5_U151 ( .A(npu_inst_pe_1_7_5_n21), .B(
        npu_inst_pe_1_7_5_n20), .S(npu_inst_pe_1_7_5_n6), .Z(
        npu_inst_pe_1_7_5_n22) );
  MUX2_X1 npu_inst_pe_1_7_5_U150 ( .A(npu_inst_pe_1_7_5_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_7_5_int_q_reg_h_1__1_), .S(npu_inst_pe_1_7_5_n4), .Z(
        npu_inst_pe_1_7_5_n21) );
  MUX2_X1 npu_inst_pe_1_7_5_U149 ( .A(npu_inst_pe_1_7_5_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_7_5_int_q_reg_h_3__1_), .S(npu_inst_pe_1_7_5_n4), .Z(
        npu_inst_pe_1_7_5_n20) );
  MUX2_X1 npu_inst_pe_1_7_5_U148 ( .A(npu_inst_pe_1_7_5_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_7_5_int_q_reg_h_5__1_), .S(npu_inst_pe_1_7_5_n4), .Z(
        npu_inst_pe_1_7_5_n19) );
  MUX2_X1 npu_inst_pe_1_7_5_U147 ( .A(npu_inst_pe_1_7_5_n18), .B(
        npu_inst_pe_1_7_5_n15), .S(npu_inst_pe_1_7_5_n8), .Z(
        npu_inst_int_data_x_7__5__0_) );
  MUX2_X1 npu_inst_pe_1_7_5_U146 ( .A(npu_inst_pe_1_7_5_n17), .B(
        npu_inst_pe_1_7_5_n16), .S(npu_inst_pe_1_7_5_n6), .Z(
        npu_inst_pe_1_7_5_n18) );
  MUX2_X1 npu_inst_pe_1_7_5_U145 ( .A(npu_inst_pe_1_7_5_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_7_5_int_q_reg_h_1__0_), .S(npu_inst_pe_1_7_5_n4), .Z(
        npu_inst_pe_1_7_5_n17) );
  MUX2_X1 npu_inst_pe_1_7_5_U144 ( .A(npu_inst_pe_1_7_5_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_7_5_int_q_reg_h_3__0_), .S(npu_inst_pe_1_7_5_n4), .Z(
        npu_inst_pe_1_7_5_n16) );
  MUX2_X1 npu_inst_pe_1_7_5_U143 ( .A(npu_inst_pe_1_7_5_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_7_5_int_q_reg_h_5__0_), .S(npu_inst_pe_1_7_5_n4), .Z(
        npu_inst_pe_1_7_5_n15) );
  XOR2_X1 npu_inst_pe_1_7_5_U142 ( .A(npu_inst_pe_1_7_5_int_data_0_), .B(
        npu_inst_pe_1_7_5_int_q_acc_0_), .Z(npu_inst_pe_1_7_5_N73) );
  AND2_X1 npu_inst_pe_1_7_5_U141 ( .A1(npu_inst_pe_1_7_5_int_q_acc_0_), .A2(
        npu_inst_pe_1_7_5_int_data_0_), .ZN(npu_inst_pe_1_7_5_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_7_5_U140 ( .A(npu_inst_pe_1_7_5_int_q_acc_0_), .B(
        npu_inst_pe_1_7_5_n13), .ZN(npu_inst_pe_1_7_5_N65) );
  OR2_X1 npu_inst_pe_1_7_5_U139 ( .A1(npu_inst_pe_1_7_5_n13), .A2(
        npu_inst_pe_1_7_5_int_q_acc_0_), .ZN(npu_inst_pe_1_7_5_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_7_5_U138 ( .A(npu_inst_pe_1_7_5_int_q_acc_2_), .B(
        npu_inst_pe_1_7_5_add_69_carry_2_), .Z(npu_inst_pe_1_7_5_N75) );
  AND2_X1 npu_inst_pe_1_7_5_U137 ( .A1(npu_inst_pe_1_7_5_add_69_carry_2_), 
        .A2(npu_inst_pe_1_7_5_int_q_acc_2_), .ZN(
        npu_inst_pe_1_7_5_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_7_5_U136 ( .A(npu_inst_pe_1_7_5_int_q_acc_3_), .B(
        npu_inst_pe_1_7_5_add_69_carry_3_), .Z(npu_inst_pe_1_7_5_N76) );
  AND2_X1 npu_inst_pe_1_7_5_U135 ( .A1(npu_inst_pe_1_7_5_add_69_carry_3_), 
        .A2(npu_inst_pe_1_7_5_int_q_acc_3_), .ZN(
        npu_inst_pe_1_7_5_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_7_5_U134 ( .A(npu_inst_pe_1_7_5_int_q_acc_4_), .B(
        npu_inst_pe_1_7_5_add_69_carry_4_), .Z(npu_inst_pe_1_7_5_N77) );
  AND2_X1 npu_inst_pe_1_7_5_U133 ( .A1(npu_inst_pe_1_7_5_add_69_carry_4_), 
        .A2(npu_inst_pe_1_7_5_int_q_acc_4_), .ZN(
        npu_inst_pe_1_7_5_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_7_5_U132 ( .A(npu_inst_pe_1_7_5_int_q_acc_5_), .B(
        npu_inst_pe_1_7_5_add_69_carry_5_), .Z(npu_inst_pe_1_7_5_N78) );
  AND2_X1 npu_inst_pe_1_7_5_U131 ( .A1(npu_inst_pe_1_7_5_add_69_carry_5_), 
        .A2(npu_inst_pe_1_7_5_int_q_acc_5_), .ZN(
        npu_inst_pe_1_7_5_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_7_5_U130 ( .A(npu_inst_pe_1_7_5_int_q_acc_6_), .B(
        npu_inst_pe_1_7_5_add_69_carry_6_), .Z(npu_inst_pe_1_7_5_N79) );
  AND2_X1 npu_inst_pe_1_7_5_U129 ( .A1(npu_inst_pe_1_7_5_add_69_carry_6_), 
        .A2(npu_inst_pe_1_7_5_int_q_acc_6_), .ZN(
        npu_inst_pe_1_7_5_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_7_5_U128 ( .A(npu_inst_pe_1_7_5_int_q_acc_7_), .B(
        npu_inst_pe_1_7_5_add_69_carry_7_), .Z(npu_inst_pe_1_7_5_N80) );
  XNOR2_X1 npu_inst_pe_1_7_5_U127 ( .A(npu_inst_pe_1_7_5_sub_67_carry_2_), .B(
        npu_inst_pe_1_7_5_int_q_acc_2_), .ZN(npu_inst_pe_1_7_5_N67) );
  OR2_X1 npu_inst_pe_1_7_5_U126 ( .A1(npu_inst_pe_1_7_5_int_q_acc_2_), .A2(
        npu_inst_pe_1_7_5_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_7_5_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_7_5_U125 ( .A(npu_inst_pe_1_7_5_sub_67_carry_3_), .B(
        npu_inst_pe_1_7_5_int_q_acc_3_), .ZN(npu_inst_pe_1_7_5_N68) );
  OR2_X1 npu_inst_pe_1_7_5_U124 ( .A1(npu_inst_pe_1_7_5_int_q_acc_3_), .A2(
        npu_inst_pe_1_7_5_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_7_5_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_7_5_U123 ( .A(npu_inst_pe_1_7_5_sub_67_carry_4_), .B(
        npu_inst_pe_1_7_5_int_q_acc_4_), .ZN(npu_inst_pe_1_7_5_N69) );
  OR2_X1 npu_inst_pe_1_7_5_U122 ( .A1(npu_inst_pe_1_7_5_int_q_acc_4_), .A2(
        npu_inst_pe_1_7_5_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_7_5_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_7_5_U121 ( .A(npu_inst_pe_1_7_5_sub_67_carry_5_), .B(
        npu_inst_pe_1_7_5_int_q_acc_5_), .ZN(npu_inst_pe_1_7_5_N70) );
  OR2_X1 npu_inst_pe_1_7_5_U120 ( .A1(npu_inst_pe_1_7_5_int_q_acc_5_), .A2(
        npu_inst_pe_1_7_5_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_7_5_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_7_5_U119 ( .A(npu_inst_pe_1_7_5_sub_67_carry_6_), .B(
        npu_inst_pe_1_7_5_int_q_acc_6_), .ZN(npu_inst_pe_1_7_5_N71) );
  OR2_X1 npu_inst_pe_1_7_5_U118 ( .A1(npu_inst_pe_1_7_5_int_q_acc_6_), .A2(
        npu_inst_pe_1_7_5_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_7_5_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_7_5_U117 ( .A(npu_inst_pe_1_7_5_int_q_acc_7_), .B(
        npu_inst_pe_1_7_5_sub_67_carry_7_), .ZN(npu_inst_pe_1_7_5_N72) );
  INV_X1 npu_inst_pe_1_7_5_U116 ( .A(npu_inst_n75), .ZN(npu_inst_pe_1_7_5_n7)
         );
  INV_X1 npu_inst_pe_1_7_5_U115 ( .A(npu_inst_pe_1_7_5_n7), .ZN(
        npu_inst_pe_1_7_5_n6) );
  INV_X1 npu_inst_pe_1_7_5_U114 ( .A(npu_inst_n52), .ZN(npu_inst_pe_1_7_5_n3)
         );
  AOI22_X1 npu_inst_pe_1_7_5_U113 ( .A1(npu_inst_pe_1_7_5_n38), .A2(
        int_i_data_v_npu[5]), .B1(npu_inst_pe_1_7_5_n114), .B2(
        npu_inst_pe_1_7_5_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_7_5_n39) );
  INV_X1 npu_inst_pe_1_7_5_U112 ( .A(npu_inst_pe_1_7_5_n39), .ZN(
        npu_inst_pe_1_7_5_n112) );
  AOI22_X1 npu_inst_pe_1_7_5_U111 ( .A1(npu_inst_pe_1_7_5_n38), .A2(
        int_i_data_v_npu[4]), .B1(npu_inst_pe_1_7_5_n114), .B2(
        npu_inst_pe_1_7_5_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_7_5_n37) );
  INV_X1 npu_inst_pe_1_7_5_U110 ( .A(npu_inst_pe_1_7_5_n37), .ZN(
        npu_inst_pe_1_7_5_n113) );
  AOI22_X1 npu_inst_pe_1_7_5_U107 ( .A1(int_i_data_v_npu[5]), .A2(
        npu_inst_pe_1_7_5_n58), .B1(npu_inst_pe_1_7_5_n119), .B2(
        npu_inst_pe_1_7_5_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_7_5_n59) );
  INV_X1 npu_inst_pe_1_7_5_U106 ( .A(npu_inst_pe_1_7_5_n59), .ZN(
        npu_inst_pe_1_7_5_n102) );
  AOI22_X1 npu_inst_pe_1_7_5_U105 ( .A1(int_i_data_v_npu[4]), .A2(
        npu_inst_pe_1_7_5_n58), .B1(npu_inst_pe_1_7_5_n119), .B2(
        npu_inst_pe_1_7_5_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_7_5_n57) );
  INV_X1 npu_inst_pe_1_7_5_U104 ( .A(npu_inst_pe_1_7_5_n57), .ZN(
        npu_inst_pe_1_7_5_n103) );
  AOI22_X1 npu_inst_pe_1_7_5_U103 ( .A1(int_i_data_v_npu[5]), .A2(
        npu_inst_pe_1_7_5_n54), .B1(npu_inst_pe_1_7_5_n118), .B2(
        npu_inst_pe_1_7_5_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_7_5_n55) );
  INV_X1 npu_inst_pe_1_7_5_U102 ( .A(npu_inst_pe_1_7_5_n55), .ZN(
        npu_inst_pe_1_7_5_n104) );
  AOI22_X1 npu_inst_pe_1_7_5_U101 ( .A1(int_i_data_v_npu[4]), .A2(
        npu_inst_pe_1_7_5_n54), .B1(npu_inst_pe_1_7_5_n118), .B2(
        npu_inst_pe_1_7_5_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_7_5_n53) );
  INV_X1 npu_inst_pe_1_7_5_U100 ( .A(npu_inst_pe_1_7_5_n53), .ZN(
        npu_inst_pe_1_7_5_n105) );
  AOI22_X1 npu_inst_pe_1_7_5_U99 ( .A1(int_i_data_v_npu[5]), .A2(
        npu_inst_pe_1_7_5_n50), .B1(npu_inst_pe_1_7_5_n117), .B2(
        npu_inst_pe_1_7_5_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_7_5_n51) );
  INV_X1 npu_inst_pe_1_7_5_U98 ( .A(npu_inst_pe_1_7_5_n51), .ZN(
        npu_inst_pe_1_7_5_n106) );
  AOI22_X1 npu_inst_pe_1_7_5_U97 ( .A1(int_i_data_v_npu[4]), .A2(
        npu_inst_pe_1_7_5_n50), .B1(npu_inst_pe_1_7_5_n117), .B2(
        npu_inst_pe_1_7_5_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_7_5_n49) );
  INV_X1 npu_inst_pe_1_7_5_U96 ( .A(npu_inst_pe_1_7_5_n49), .ZN(
        npu_inst_pe_1_7_5_n107) );
  AOI22_X1 npu_inst_pe_1_7_5_U95 ( .A1(int_i_data_v_npu[5]), .A2(
        npu_inst_pe_1_7_5_n46), .B1(npu_inst_pe_1_7_5_n116), .B2(
        npu_inst_pe_1_7_5_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_7_5_n47) );
  INV_X1 npu_inst_pe_1_7_5_U94 ( .A(npu_inst_pe_1_7_5_n47), .ZN(
        npu_inst_pe_1_7_5_n108) );
  AOI22_X1 npu_inst_pe_1_7_5_U93 ( .A1(int_i_data_v_npu[4]), .A2(
        npu_inst_pe_1_7_5_n46), .B1(npu_inst_pe_1_7_5_n116), .B2(
        npu_inst_pe_1_7_5_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_7_5_n45) );
  INV_X1 npu_inst_pe_1_7_5_U92 ( .A(npu_inst_pe_1_7_5_n45), .ZN(
        npu_inst_pe_1_7_5_n109) );
  AOI22_X1 npu_inst_pe_1_7_5_U91 ( .A1(int_i_data_v_npu[5]), .A2(
        npu_inst_pe_1_7_5_n42), .B1(npu_inst_pe_1_7_5_n115), .B2(
        npu_inst_pe_1_7_5_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_7_5_n43) );
  INV_X1 npu_inst_pe_1_7_5_U90 ( .A(npu_inst_pe_1_7_5_n43), .ZN(
        npu_inst_pe_1_7_5_n110) );
  AOI22_X1 npu_inst_pe_1_7_5_U89 ( .A1(int_i_data_v_npu[4]), .A2(
        npu_inst_pe_1_7_5_n42), .B1(npu_inst_pe_1_7_5_n115), .B2(
        npu_inst_pe_1_7_5_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_7_5_n41) );
  INV_X1 npu_inst_pe_1_7_5_U88 ( .A(npu_inst_pe_1_7_5_n41), .ZN(
        npu_inst_pe_1_7_5_n111) );
  NAND2_X1 npu_inst_pe_1_7_5_U87 ( .A1(npu_inst_pe_1_7_5_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_7_5_n60), .ZN(npu_inst_pe_1_7_5_n74) );
  OAI21_X1 npu_inst_pe_1_7_5_U86 ( .B1(npu_inst_pe_1_7_5_n63), .B2(
        npu_inst_pe_1_7_5_n60), .A(npu_inst_pe_1_7_5_n74), .ZN(
        npu_inst_pe_1_7_5_n97) );
  NAND2_X1 npu_inst_pe_1_7_5_U85 ( .A1(npu_inst_pe_1_7_5_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_7_5_n60), .ZN(npu_inst_pe_1_7_5_n73) );
  OAI21_X1 npu_inst_pe_1_7_5_U84 ( .B1(npu_inst_pe_1_7_5_n61), .B2(
        npu_inst_pe_1_7_5_n60), .A(npu_inst_pe_1_7_5_n73), .ZN(
        npu_inst_pe_1_7_5_n96) );
  NAND2_X1 npu_inst_pe_1_7_5_U83 ( .A1(npu_inst_pe_1_7_5_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_7_5_n56), .ZN(npu_inst_pe_1_7_5_n72) );
  OAI21_X1 npu_inst_pe_1_7_5_U82 ( .B1(npu_inst_pe_1_7_5_n63), .B2(
        npu_inst_pe_1_7_5_n56), .A(npu_inst_pe_1_7_5_n72), .ZN(
        npu_inst_pe_1_7_5_n95) );
  NAND2_X1 npu_inst_pe_1_7_5_U81 ( .A1(npu_inst_pe_1_7_5_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_7_5_n56), .ZN(npu_inst_pe_1_7_5_n71) );
  OAI21_X1 npu_inst_pe_1_7_5_U80 ( .B1(npu_inst_pe_1_7_5_n61), .B2(
        npu_inst_pe_1_7_5_n56), .A(npu_inst_pe_1_7_5_n71), .ZN(
        npu_inst_pe_1_7_5_n94) );
  NAND2_X1 npu_inst_pe_1_7_5_U79 ( .A1(npu_inst_pe_1_7_5_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_7_5_n52), .ZN(npu_inst_pe_1_7_5_n70) );
  OAI21_X1 npu_inst_pe_1_7_5_U78 ( .B1(npu_inst_pe_1_7_5_n63), .B2(
        npu_inst_pe_1_7_5_n52), .A(npu_inst_pe_1_7_5_n70), .ZN(
        npu_inst_pe_1_7_5_n93) );
  NAND2_X1 npu_inst_pe_1_7_5_U77 ( .A1(npu_inst_pe_1_7_5_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_7_5_n52), .ZN(npu_inst_pe_1_7_5_n69) );
  OAI21_X1 npu_inst_pe_1_7_5_U76 ( .B1(npu_inst_pe_1_7_5_n61), .B2(
        npu_inst_pe_1_7_5_n52), .A(npu_inst_pe_1_7_5_n69), .ZN(
        npu_inst_pe_1_7_5_n92) );
  NAND2_X1 npu_inst_pe_1_7_5_U75 ( .A1(npu_inst_pe_1_7_5_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_7_5_n48), .ZN(npu_inst_pe_1_7_5_n68) );
  OAI21_X1 npu_inst_pe_1_7_5_U74 ( .B1(npu_inst_pe_1_7_5_n63), .B2(
        npu_inst_pe_1_7_5_n48), .A(npu_inst_pe_1_7_5_n68), .ZN(
        npu_inst_pe_1_7_5_n91) );
  NAND2_X1 npu_inst_pe_1_7_5_U73 ( .A1(npu_inst_pe_1_7_5_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_7_5_n48), .ZN(npu_inst_pe_1_7_5_n67) );
  OAI21_X1 npu_inst_pe_1_7_5_U72 ( .B1(npu_inst_pe_1_7_5_n61), .B2(
        npu_inst_pe_1_7_5_n48), .A(npu_inst_pe_1_7_5_n67), .ZN(
        npu_inst_pe_1_7_5_n90) );
  NAND2_X1 npu_inst_pe_1_7_5_U71 ( .A1(npu_inst_pe_1_7_5_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_7_5_n44), .ZN(npu_inst_pe_1_7_5_n66) );
  OAI21_X1 npu_inst_pe_1_7_5_U70 ( .B1(npu_inst_pe_1_7_5_n63), .B2(
        npu_inst_pe_1_7_5_n44), .A(npu_inst_pe_1_7_5_n66), .ZN(
        npu_inst_pe_1_7_5_n89) );
  NAND2_X1 npu_inst_pe_1_7_5_U69 ( .A1(npu_inst_pe_1_7_5_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_7_5_n44), .ZN(npu_inst_pe_1_7_5_n65) );
  OAI21_X1 npu_inst_pe_1_7_5_U68 ( .B1(npu_inst_pe_1_7_5_n61), .B2(
        npu_inst_pe_1_7_5_n44), .A(npu_inst_pe_1_7_5_n65), .ZN(
        npu_inst_pe_1_7_5_n88) );
  NAND2_X1 npu_inst_pe_1_7_5_U67 ( .A1(npu_inst_pe_1_7_5_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_7_5_n40), .ZN(npu_inst_pe_1_7_5_n64) );
  OAI21_X1 npu_inst_pe_1_7_5_U66 ( .B1(npu_inst_pe_1_7_5_n63), .B2(
        npu_inst_pe_1_7_5_n40), .A(npu_inst_pe_1_7_5_n64), .ZN(
        npu_inst_pe_1_7_5_n87) );
  NAND2_X1 npu_inst_pe_1_7_5_U65 ( .A1(npu_inst_pe_1_7_5_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_7_5_n40), .ZN(npu_inst_pe_1_7_5_n62) );
  OAI21_X1 npu_inst_pe_1_7_5_U64 ( .B1(npu_inst_pe_1_7_5_n61), .B2(
        npu_inst_pe_1_7_5_n40), .A(npu_inst_pe_1_7_5_n62), .ZN(
        npu_inst_pe_1_7_5_n86) );
  AND2_X1 npu_inst_pe_1_7_5_U63 ( .A1(npu_inst_pe_1_7_5_N93), .A2(npu_inst_n52), .ZN(npu_inst_int_data_y_7__5__0_) );
  AND2_X1 npu_inst_pe_1_7_5_U62 ( .A1(npu_inst_n52), .A2(npu_inst_pe_1_7_5_N94), .ZN(npu_inst_int_data_y_7__5__1_) );
  AOI22_X1 npu_inst_pe_1_7_5_U61 ( .A1(npu_inst_n52), .A2(int_i_data_v_npu[5]), 
        .B1(npu_inst_pe_1_7_5_n3), .B2(npu_inst_int_data_x_7__6__1_), .ZN(
        npu_inst_pe_1_7_5_n63) );
  AOI22_X1 npu_inst_pe_1_7_5_U60 ( .A1(npu_inst_n52), .A2(int_i_data_v_npu[4]), 
        .B1(npu_inst_pe_1_7_5_n3), .B2(npu_inst_int_data_x_7__6__0_), .ZN(
        npu_inst_pe_1_7_5_n61) );
  AOI222_X1 npu_inst_pe_1_7_5_U59 ( .A1(1'b0), .A2(npu_inst_pe_1_7_5_n1), .B1(
        npu_inst_pe_1_7_5_N73), .B2(npu_inst_pe_1_7_5_n76), .C1(
        npu_inst_pe_1_7_5_N65), .C2(npu_inst_pe_1_7_5_n77), .ZN(
        npu_inst_pe_1_7_5_n84) );
  INV_X1 npu_inst_pe_1_7_5_U58 ( .A(npu_inst_pe_1_7_5_n84), .ZN(
        npu_inst_pe_1_7_5_n101) );
  AOI222_X1 npu_inst_pe_1_7_5_U57 ( .A1(1'b0), .A2(npu_inst_pe_1_7_5_n1), .B1(
        npu_inst_pe_1_7_5_N80), .B2(npu_inst_pe_1_7_5_n76), .C1(
        npu_inst_pe_1_7_5_N72), .C2(npu_inst_pe_1_7_5_n77), .ZN(
        npu_inst_pe_1_7_5_n75) );
  INV_X1 npu_inst_pe_1_7_5_U56 ( .A(npu_inst_pe_1_7_5_n75), .ZN(
        npu_inst_pe_1_7_5_n33) );
  AOI222_X1 npu_inst_pe_1_7_5_U55 ( .A1(1'b0), .A2(npu_inst_pe_1_7_5_n1), .B1(
        npu_inst_pe_1_7_5_N74), .B2(npu_inst_pe_1_7_5_n76), .C1(
        npu_inst_pe_1_7_5_N66), .C2(npu_inst_pe_1_7_5_n77), .ZN(
        npu_inst_pe_1_7_5_n83) );
  INV_X1 npu_inst_pe_1_7_5_U54 ( .A(npu_inst_pe_1_7_5_n83), .ZN(
        npu_inst_pe_1_7_5_n100) );
  AOI222_X1 npu_inst_pe_1_7_5_U53 ( .A1(1'b0), .A2(npu_inst_pe_1_7_5_n1), .B1(
        npu_inst_pe_1_7_5_N75), .B2(npu_inst_pe_1_7_5_n76), .C1(
        npu_inst_pe_1_7_5_N67), .C2(npu_inst_pe_1_7_5_n77), .ZN(
        npu_inst_pe_1_7_5_n82) );
  INV_X1 npu_inst_pe_1_7_5_U52 ( .A(npu_inst_pe_1_7_5_n82), .ZN(
        npu_inst_pe_1_7_5_n99) );
  AOI222_X1 npu_inst_pe_1_7_5_U51 ( .A1(1'b0), .A2(npu_inst_pe_1_7_5_n1), .B1(
        npu_inst_pe_1_7_5_N76), .B2(npu_inst_pe_1_7_5_n76), .C1(
        npu_inst_pe_1_7_5_N68), .C2(npu_inst_pe_1_7_5_n77), .ZN(
        npu_inst_pe_1_7_5_n81) );
  INV_X1 npu_inst_pe_1_7_5_U50 ( .A(npu_inst_pe_1_7_5_n81), .ZN(
        npu_inst_pe_1_7_5_n98) );
  AOI222_X1 npu_inst_pe_1_7_5_U49 ( .A1(1'b0), .A2(npu_inst_pe_1_7_5_n1), .B1(
        npu_inst_pe_1_7_5_N77), .B2(npu_inst_pe_1_7_5_n76), .C1(
        npu_inst_pe_1_7_5_N69), .C2(npu_inst_pe_1_7_5_n77), .ZN(
        npu_inst_pe_1_7_5_n80) );
  INV_X1 npu_inst_pe_1_7_5_U48 ( .A(npu_inst_pe_1_7_5_n80), .ZN(
        npu_inst_pe_1_7_5_n36) );
  AOI222_X1 npu_inst_pe_1_7_5_U47 ( .A1(1'b0), .A2(npu_inst_pe_1_7_5_n1), .B1(
        npu_inst_pe_1_7_5_N78), .B2(npu_inst_pe_1_7_5_n76), .C1(
        npu_inst_pe_1_7_5_N70), .C2(npu_inst_pe_1_7_5_n77), .ZN(
        npu_inst_pe_1_7_5_n79) );
  INV_X1 npu_inst_pe_1_7_5_U46 ( .A(npu_inst_pe_1_7_5_n79), .ZN(
        npu_inst_pe_1_7_5_n35) );
  AOI222_X1 npu_inst_pe_1_7_5_U45 ( .A1(1'b0), .A2(npu_inst_pe_1_7_5_n1), .B1(
        npu_inst_pe_1_7_5_N79), .B2(npu_inst_pe_1_7_5_n76), .C1(
        npu_inst_pe_1_7_5_N71), .C2(npu_inst_pe_1_7_5_n77), .ZN(
        npu_inst_pe_1_7_5_n78) );
  INV_X1 npu_inst_pe_1_7_5_U44 ( .A(npu_inst_pe_1_7_5_n78), .ZN(
        npu_inst_pe_1_7_5_n34) );
  AND2_X1 npu_inst_pe_1_7_5_U43 ( .A1(npu_inst_pe_1_7_5_int_q_acc_0_), .A2(
        npu_inst_pe_1_7_5_n1), .ZN(npu_inst_int_data_res_7__5__0_) );
  AND2_X1 npu_inst_pe_1_7_5_U42 ( .A1(npu_inst_pe_1_7_5_n2), .A2(
        npu_inst_pe_1_7_5_int_q_acc_7_), .ZN(npu_inst_int_data_res_7__5__7_)
         );
  AND2_X1 npu_inst_pe_1_7_5_U41 ( .A1(npu_inst_pe_1_7_5_int_q_acc_1_), .A2(
        npu_inst_pe_1_7_5_n1), .ZN(npu_inst_int_data_res_7__5__1_) );
  AND2_X1 npu_inst_pe_1_7_5_U40 ( .A1(npu_inst_pe_1_7_5_int_q_acc_2_), .A2(
        npu_inst_pe_1_7_5_n1), .ZN(npu_inst_int_data_res_7__5__2_) );
  AND2_X1 npu_inst_pe_1_7_5_U39 ( .A1(npu_inst_pe_1_7_5_int_q_acc_3_), .A2(
        npu_inst_pe_1_7_5_n2), .ZN(npu_inst_int_data_res_7__5__3_) );
  AND2_X1 npu_inst_pe_1_7_5_U38 ( .A1(npu_inst_pe_1_7_5_int_q_acc_4_), .A2(
        npu_inst_pe_1_7_5_n2), .ZN(npu_inst_int_data_res_7__5__4_) );
  AND2_X1 npu_inst_pe_1_7_5_U37 ( .A1(npu_inst_pe_1_7_5_int_q_acc_5_), .A2(
        npu_inst_pe_1_7_5_n2), .ZN(npu_inst_int_data_res_7__5__5_) );
  AND2_X1 npu_inst_pe_1_7_5_U36 ( .A1(npu_inst_pe_1_7_5_int_q_acc_6_), .A2(
        npu_inst_pe_1_7_5_n2), .ZN(npu_inst_int_data_res_7__5__6_) );
  INV_X1 npu_inst_pe_1_7_5_U35 ( .A(npu_inst_pe_1_7_5_int_data_1_), .ZN(
        npu_inst_pe_1_7_5_n14) );
  NOR3_X1 npu_inst_pe_1_7_5_U34 ( .A1(npu_inst_pe_1_7_5_n26), .A2(npu_inst_n52), .A3(npu_inst_int_ckg[2]), .ZN(npu_inst_pe_1_7_5_n85) );
  OR2_X1 npu_inst_pe_1_7_5_U33 ( .A1(npu_inst_pe_1_7_5_n85), .A2(
        npu_inst_pe_1_7_5_n2), .ZN(npu_inst_pe_1_7_5_N84) );
  AND2_X1 npu_inst_pe_1_7_5_U32 ( .A1(npu_inst_int_data_x_7__5__1_), .A2(
        npu_inst_pe_1_7_5_int_q_weight_1_), .ZN(npu_inst_pe_1_7_5_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_7_5_U31 ( .A1(npu_inst_int_data_x_7__5__0_), .A2(
        npu_inst_pe_1_7_5_int_q_weight_1_), .ZN(npu_inst_pe_1_7_5_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_7_5_U30 ( .A(npu_inst_pe_1_7_5_int_data_0_), .ZN(
        npu_inst_pe_1_7_5_n13) );
  INV_X1 npu_inst_pe_1_7_5_U29 ( .A(npu_inst_n67), .ZN(npu_inst_pe_1_7_5_n5)
         );
  OR3_X1 npu_inst_pe_1_7_5_U28 ( .A1(npu_inst_pe_1_7_5_n6), .A2(
        npu_inst_pe_1_7_5_n8), .A3(npu_inst_pe_1_7_5_n5), .ZN(
        npu_inst_pe_1_7_5_n56) );
  OR3_X1 npu_inst_pe_1_7_5_U27 ( .A1(npu_inst_pe_1_7_5_n5), .A2(
        npu_inst_pe_1_7_5_n8), .A3(npu_inst_pe_1_7_5_n7), .ZN(
        npu_inst_pe_1_7_5_n48) );
  INV_X1 npu_inst_pe_1_7_5_U26 ( .A(npu_inst_pe_1_7_5_n5), .ZN(
        npu_inst_pe_1_7_5_n4) );
  OR3_X1 npu_inst_pe_1_7_5_U25 ( .A1(npu_inst_pe_1_7_5_n4), .A2(
        npu_inst_pe_1_7_5_n8), .A3(npu_inst_pe_1_7_5_n7), .ZN(
        npu_inst_pe_1_7_5_n52) );
  OR3_X1 npu_inst_pe_1_7_5_U24 ( .A1(npu_inst_pe_1_7_5_n6), .A2(
        npu_inst_pe_1_7_5_n8), .A3(npu_inst_pe_1_7_5_n4), .ZN(
        npu_inst_pe_1_7_5_n60) );
  NOR2_X1 npu_inst_pe_1_7_5_U23 ( .A1(npu_inst_pe_1_7_5_n60), .A2(
        npu_inst_pe_1_7_5_n3), .ZN(npu_inst_pe_1_7_5_n58) );
  NOR2_X1 npu_inst_pe_1_7_5_U22 ( .A1(npu_inst_pe_1_7_5_n56), .A2(
        npu_inst_pe_1_7_5_n3), .ZN(npu_inst_pe_1_7_5_n54) );
  NOR2_X1 npu_inst_pe_1_7_5_U21 ( .A1(npu_inst_pe_1_7_5_n52), .A2(
        npu_inst_pe_1_7_5_n3), .ZN(npu_inst_pe_1_7_5_n50) );
  NOR2_X1 npu_inst_pe_1_7_5_U20 ( .A1(npu_inst_pe_1_7_5_n48), .A2(
        npu_inst_pe_1_7_5_n3), .ZN(npu_inst_pe_1_7_5_n46) );
  NOR2_X1 npu_inst_pe_1_7_5_U19 ( .A1(npu_inst_pe_1_7_5_n40), .A2(
        npu_inst_pe_1_7_5_n3), .ZN(npu_inst_pe_1_7_5_n38) );
  NOR2_X1 npu_inst_pe_1_7_5_U18 ( .A1(npu_inst_pe_1_7_5_n44), .A2(
        npu_inst_pe_1_7_5_n3), .ZN(npu_inst_pe_1_7_5_n42) );
  BUF_X1 npu_inst_pe_1_7_5_U17 ( .A(npu_inst_n92), .Z(npu_inst_pe_1_7_5_n8) );
  INV_X1 npu_inst_pe_1_7_5_U16 ( .A(npu_inst_n122), .ZN(npu_inst_pe_1_7_5_n12)
         );
  INV_X1 npu_inst_pe_1_7_5_U15 ( .A(npu_inst_pe_1_7_5_n38), .ZN(
        npu_inst_pe_1_7_5_n114) );
  INV_X1 npu_inst_pe_1_7_5_U14 ( .A(npu_inst_pe_1_7_5_n58), .ZN(
        npu_inst_pe_1_7_5_n119) );
  INV_X1 npu_inst_pe_1_7_5_U13 ( .A(npu_inst_pe_1_7_5_n54), .ZN(
        npu_inst_pe_1_7_5_n118) );
  INV_X1 npu_inst_pe_1_7_5_U12 ( .A(npu_inst_pe_1_7_5_n50), .ZN(
        npu_inst_pe_1_7_5_n117) );
  INV_X1 npu_inst_pe_1_7_5_U11 ( .A(npu_inst_pe_1_7_5_n46), .ZN(
        npu_inst_pe_1_7_5_n116) );
  INV_X1 npu_inst_pe_1_7_5_U10 ( .A(npu_inst_pe_1_7_5_n42), .ZN(
        npu_inst_pe_1_7_5_n115) );
  BUF_X1 npu_inst_pe_1_7_5_U9 ( .A(npu_inst_n8), .Z(npu_inst_pe_1_7_5_n2) );
  BUF_X1 npu_inst_pe_1_7_5_U8 ( .A(npu_inst_n8), .Z(npu_inst_pe_1_7_5_n1) );
  BUF_X1 npu_inst_pe_1_7_5_U7 ( .A(npu_inst_pe_1_7_5_n12), .Z(
        npu_inst_pe_1_7_5_n11) );
  BUF_X1 npu_inst_pe_1_7_5_U6 ( .A(npu_inst_pe_1_7_5_n12), .Z(
        npu_inst_pe_1_7_5_n10) );
  BUF_X1 npu_inst_pe_1_7_5_U5 ( .A(npu_inst_pe_1_7_5_n12), .Z(
        npu_inst_pe_1_7_5_n9) );
  NOR2_X1 npu_inst_pe_1_7_5_U4 ( .A1(npu_inst_pe_1_7_5_int_q_weight_0_), .A2(
        npu_inst_pe_1_7_5_n1), .ZN(npu_inst_pe_1_7_5_n76) );
  NOR2_X1 npu_inst_pe_1_7_5_U3 ( .A1(npu_inst_pe_1_7_5_n27), .A2(
        npu_inst_pe_1_7_5_n1), .ZN(npu_inst_pe_1_7_5_n77) );
  FA_X1 npu_inst_pe_1_7_5_sub_67_U2_1 ( .A(npu_inst_pe_1_7_5_int_q_acc_1_), 
        .B(npu_inst_pe_1_7_5_n14), .CI(npu_inst_pe_1_7_5_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_7_5_sub_67_carry_2_), .S(npu_inst_pe_1_7_5_N66) );
  FA_X1 npu_inst_pe_1_7_5_add_69_U1_1 ( .A(npu_inst_pe_1_7_5_int_q_acc_1_), 
        .B(npu_inst_pe_1_7_5_int_data_1_), .CI(
        npu_inst_pe_1_7_5_add_69_carry_1_), .CO(
        npu_inst_pe_1_7_5_add_69_carry_2_), .S(npu_inst_pe_1_7_5_N74) );
  NAND3_X1 npu_inst_pe_1_7_5_U109 ( .A1(npu_inst_pe_1_7_5_n5), .A2(
        npu_inst_pe_1_7_5_n7), .A3(npu_inst_pe_1_7_5_n8), .ZN(
        npu_inst_pe_1_7_5_n44) );
  NAND3_X1 npu_inst_pe_1_7_5_U108 ( .A1(npu_inst_pe_1_7_5_n4), .A2(
        npu_inst_pe_1_7_5_n7), .A3(npu_inst_pe_1_7_5_n8), .ZN(
        npu_inst_pe_1_7_5_n40) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_7_5_n34), .CK(
        npu_inst_pe_1_7_5_net3159), .RN(npu_inst_pe_1_7_5_n9), .Q(
        npu_inst_pe_1_7_5_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_7_5_n35), .CK(
        npu_inst_pe_1_7_5_net3159), .RN(npu_inst_pe_1_7_5_n9), .Q(
        npu_inst_pe_1_7_5_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_7_5_n36), .CK(
        npu_inst_pe_1_7_5_net3159), .RN(npu_inst_pe_1_7_5_n9), .Q(
        npu_inst_pe_1_7_5_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_7_5_n98), .CK(
        npu_inst_pe_1_7_5_net3159), .RN(npu_inst_pe_1_7_5_n9), .Q(
        npu_inst_pe_1_7_5_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_7_5_n99), .CK(
        npu_inst_pe_1_7_5_net3159), .RN(npu_inst_pe_1_7_5_n9), .Q(
        npu_inst_pe_1_7_5_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_7_5_n100), 
        .CK(npu_inst_pe_1_7_5_net3159), .RN(npu_inst_pe_1_7_5_n9), .Q(
        npu_inst_pe_1_7_5_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_7_5_n33), .CK(
        npu_inst_pe_1_7_5_net3159), .RN(npu_inst_pe_1_7_5_n9), .Q(
        npu_inst_pe_1_7_5_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_7_5_n101), 
        .CK(npu_inst_pe_1_7_5_net3159), .RN(npu_inst_pe_1_7_5_n9), .Q(
        npu_inst_pe_1_7_5_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_weight_reg_0_ ( .D(npu_inst_n108), .CK(
        npu_inst_pe_1_7_5_net3165), .RN(npu_inst_pe_1_7_5_n9), .Q(
        npu_inst_pe_1_7_5_int_q_weight_0_), .QN(npu_inst_pe_1_7_5_n27) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_weight_reg_1_ ( .D(npu_inst_n114), .CK(
        npu_inst_pe_1_7_5_net3165), .RN(npu_inst_pe_1_7_5_n9), .Q(
        npu_inst_pe_1_7_5_int_q_weight_1_), .QN(npu_inst_pe_1_7_5_n26) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_7_5_n113), 
        .CK(npu_inst_pe_1_7_5_net3165), .RN(npu_inst_pe_1_7_5_n9), .Q(
        npu_inst_pe_1_7_5_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_7_5_n112), 
        .CK(npu_inst_pe_1_7_5_net3165), .RN(npu_inst_pe_1_7_5_n9), .Q(
        npu_inst_pe_1_7_5_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_7_5_n111), 
        .CK(npu_inst_pe_1_7_5_net3165), .RN(npu_inst_pe_1_7_5_n10), .Q(
        npu_inst_pe_1_7_5_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_7_5_n110), 
        .CK(npu_inst_pe_1_7_5_net3165), .RN(npu_inst_pe_1_7_5_n10), .Q(
        npu_inst_pe_1_7_5_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_7_5_n109), 
        .CK(npu_inst_pe_1_7_5_net3165), .RN(npu_inst_pe_1_7_5_n10), .Q(
        npu_inst_pe_1_7_5_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_7_5_n108), 
        .CK(npu_inst_pe_1_7_5_net3165), .RN(npu_inst_pe_1_7_5_n10), .Q(
        npu_inst_pe_1_7_5_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_7_5_n107), 
        .CK(npu_inst_pe_1_7_5_net3165), .RN(npu_inst_pe_1_7_5_n10), .Q(
        npu_inst_pe_1_7_5_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_7_5_n106), 
        .CK(npu_inst_pe_1_7_5_net3165), .RN(npu_inst_pe_1_7_5_n10), .Q(
        npu_inst_pe_1_7_5_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_7_5_n105), 
        .CK(npu_inst_pe_1_7_5_net3165), .RN(npu_inst_pe_1_7_5_n10), .Q(
        npu_inst_pe_1_7_5_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_7_5_n104), 
        .CK(npu_inst_pe_1_7_5_net3165), .RN(npu_inst_pe_1_7_5_n10), .Q(
        npu_inst_pe_1_7_5_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_7_5_n103), 
        .CK(npu_inst_pe_1_7_5_net3165), .RN(npu_inst_pe_1_7_5_n10), .Q(
        npu_inst_pe_1_7_5_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_7_5_n102), 
        .CK(npu_inst_pe_1_7_5_net3165), .RN(npu_inst_pe_1_7_5_n10), .Q(
        npu_inst_pe_1_7_5_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_7_5_n86), 
        .CK(npu_inst_pe_1_7_5_net3165), .RN(npu_inst_pe_1_7_5_n10), .Q(
        npu_inst_pe_1_7_5_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_7_5_n87), 
        .CK(npu_inst_pe_1_7_5_net3165), .RN(npu_inst_pe_1_7_5_n10), .Q(
        npu_inst_pe_1_7_5_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_7_5_n88), 
        .CK(npu_inst_pe_1_7_5_net3165), .RN(npu_inst_pe_1_7_5_n11), .Q(
        npu_inst_pe_1_7_5_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_7_5_n89), 
        .CK(npu_inst_pe_1_7_5_net3165), .RN(npu_inst_pe_1_7_5_n11), .Q(
        npu_inst_pe_1_7_5_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_7_5_n90), 
        .CK(npu_inst_pe_1_7_5_net3165), .RN(npu_inst_pe_1_7_5_n11), .Q(
        npu_inst_pe_1_7_5_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_7_5_n91), 
        .CK(npu_inst_pe_1_7_5_net3165), .RN(npu_inst_pe_1_7_5_n11), .Q(
        npu_inst_pe_1_7_5_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_7_5_n92), 
        .CK(npu_inst_pe_1_7_5_net3165), .RN(npu_inst_pe_1_7_5_n11), .Q(
        npu_inst_pe_1_7_5_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_7_5_n93), 
        .CK(npu_inst_pe_1_7_5_net3165), .RN(npu_inst_pe_1_7_5_n11), .Q(
        npu_inst_pe_1_7_5_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_7_5_n94), 
        .CK(npu_inst_pe_1_7_5_net3165), .RN(npu_inst_pe_1_7_5_n11), .Q(
        npu_inst_pe_1_7_5_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_7_5_n95), 
        .CK(npu_inst_pe_1_7_5_net3165), .RN(npu_inst_pe_1_7_5_n11), .Q(
        npu_inst_pe_1_7_5_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_7_5_n96), 
        .CK(npu_inst_pe_1_7_5_net3165), .RN(npu_inst_pe_1_7_5_n11), .Q(
        npu_inst_pe_1_7_5_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_7_5_n97), 
        .CK(npu_inst_pe_1_7_5_net3165), .RN(npu_inst_pe_1_7_5_n11), .Q(
        npu_inst_pe_1_7_5_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_7_5_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_7_5_N84), .SE(1'b0), .GCK(npu_inst_pe_1_7_5_net3159) );
  CLKGATETST_X1 npu_inst_pe_1_7_5_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n61), .SE(1'b0), .GCK(npu_inst_pe_1_7_5_net3165) );
  MUX2_X1 npu_inst_pe_1_7_6_U162 ( .A(npu_inst_pe_1_7_6_n32), .B(
        npu_inst_pe_1_7_6_n29), .S(npu_inst_pe_1_7_6_n8), .Z(
        npu_inst_pe_1_7_6_N93) );
  MUX2_X1 npu_inst_pe_1_7_6_U161 ( .A(npu_inst_pe_1_7_6_n31), .B(
        npu_inst_pe_1_7_6_n30), .S(npu_inst_pe_1_7_6_n6), .Z(
        npu_inst_pe_1_7_6_n32) );
  MUX2_X1 npu_inst_pe_1_7_6_U160 ( .A(npu_inst_pe_1_7_6_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_7_6_int_q_reg_v_1__0_), .S(npu_inst_pe_1_7_6_n4), .Z(
        npu_inst_pe_1_7_6_n31) );
  MUX2_X1 npu_inst_pe_1_7_6_U159 ( .A(npu_inst_pe_1_7_6_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_7_6_int_q_reg_v_3__0_), .S(npu_inst_pe_1_7_6_n4), .Z(
        npu_inst_pe_1_7_6_n30) );
  MUX2_X1 npu_inst_pe_1_7_6_U158 ( .A(npu_inst_pe_1_7_6_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_7_6_int_q_reg_v_5__0_), .S(npu_inst_pe_1_7_6_n4), .Z(
        npu_inst_pe_1_7_6_n29) );
  MUX2_X1 npu_inst_pe_1_7_6_U157 ( .A(npu_inst_pe_1_7_6_n28), .B(
        npu_inst_pe_1_7_6_n23), .S(npu_inst_pe_1_7_6_n8), .Z(
        npu_inst_pe_1_7_6_N94) );
  MUX2_X1 npu_inst_pe_1_7_6_U156 ( .A(npu_inst_pe_1_7_6_n25), .B(
        npu_inst_pe_1_7_6_n24), .S(npu_inst_pe_1_7_6_n6), .Z(
        npu_inst_pe_1_7_6_n28) );
  MUX2_X1 npu_inst_pe_1_7_6_U155 ( .A(npu_inst_pe_1_7_6_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_7_6_int_q_reg_v_1__1_), .S(npu_inst_pe_1_7_6_n4), .Z(
        npu_inst_pe_1_7_6_n25) );
  MUX2_X1 npu_inst_pe_1_7_6_U154 ( .A(npu_inst_pe_1_7_6_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_7_6_int_q_reg_v_3__1_), .S(npu_inst_pe_1_7_6_n4), .Z(
        npu_inst_pe_1_7_6_n24) );
  MUX2_X1 npu_inst_pe_1_7_6_U153 ( .A(npu_inst_pe_1_7_6_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_7_6_int_q_reg_v_5__1_), .S(npu_inst_pe_1_7_6_n4), .Z(
        npu_inst_pe_1_7_6_n23) );
  MUX2_X1 npu_inst_pe_1_7_6_U152 ( .A(npu_inst_pe_1_7_6_n22), .B(
        npu_inst_pe_1_7_6_n19), .S(npu_inst_pe_1_7_6_n8), .Z(
        npu_inst_int_data_x_7__6__1_) );
  MUX2_X1 npu_inst_pe_1_7_6_U151 ( .A(npu_inst_pe_1_7_6_n21), .B(
        npu_inst_pe_1_7_6_n20), .S(npu_inst_pe_1_7_6_n6), .Z(
        npu_inst_pe_1_7_6_n22) );
  MUX2_X1 npu_inst_pe_1_7_6_U150 ( .A(npu_inst_pe_1_7_6_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_7_6_int_q_reg_h_1__1_), .S(npu_inst_pe_1_7_6_n4), .Z(
        npu_inst_pe_1_7_6_n21) );
  MUX2_X1 npu_inst_pe_1_7_6_U149 ( .A(npu_inst_pe_1_7_6_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_7_6_int_q_reg_h_3__1_), .S(npu_inst_pe_1_7_6_n4), .Z(
        npu_inst_pe_1_7_6_n20) );
  MUX2_X1 npu_inst_pe_1_7_6_U148 ( .A(npu_inst_pe_1_7_6_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_7_6_int_q_reg_h_5__1_), .S(npu_inst_pe_1_7_6_n4), .Z(
        npu_inst_pe_1_7_6_n19) );
  MUX2_X1 npu_inst_pe_1_7_6_U147 ( .A(npu_inst_pe_1_7_6_n18), .B(
        npu_inst_pe_1_7_6_n15), .S(npu_inst_pe_1_7_6_n8), .Z(
        npu_inst_int_data_x_7__6__0_) );
  MUX2_X1 npu_inst_pe_1_7_6_U146 ( .A(npu_inst_pe_1_7_6_n17), .B(
        npu_inst_pe_1_7_6_n16), .S(npu_inst_pe_1_7_6_n6), .Z(
        npu_inst_pe_1_7_6_n18) );
  MUX2_X1 npu_inst_pe_1_7_6_U145 ( .A(npu_inst_pe_1_7_6_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_7_6_int_q_reg_h_1__0_), .S(npu_inst_pe_1_7_6_n4), .Z(
        npu_inst_pe_1_7_6_n17) );
  MUX2_X1 npu_inst_pe_1_7_6_U144 ( .A(npu_inst_pe_1_7_6_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_7_6_int_q_reg_h_3__0_), .S(npu_inst_pe_1_7_6_n4), .Z(
        npu_inst_pe_1_7_6_n16) );
  MUX2_X1 npu_inst_pe_1_7_6_U143 ( .A(npu_inst_pe_1_7_6_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_7_6_int_q_reg_h_5__0_), .S(npu_inst_pe_1_7_6_n4), .Z(
        npu_inst_pe_1_7_6_n15) );
  XOR2_X1 npu_inst_pe_1_7_6_U142 ( .A(npu_inst_pe_1_7_6_int_data_0_), .B(
        npu_inst_pe_1_7_6_int_q_acc_0_), .Z(npu_inst_pe_1_7_6_N73) );
  AND2_X1 npu_inst_pe_1_7_6_U141 ( .A1(npu_inst_pe_1_7_6_int_q_acc_0_), .A2(
        npu_inst_pe_1_7_6_int_data_0_), .ZN(npu_inst_pe_1_7_6_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_7_6_U140 ( .A(npu_inst_pe_1_7_6_int_q_acc_0_), .B(
        npu_inst_pe_1_7_6_n13), .ZN(npu_inst_pe_1_7_6_N65) );
  OR2_X1 npu_inst_pe_1_7_6_U139 ( .A1(npu_inst_pe_1_7_6_n13), .A2(
        npu_inst_pe_1_7_6_int_q_acc_0_), .ZN(npu_inst_pe_1_7_6_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_7_6_U138 ( .A(npu_inst_pe_1_7_6_int_q_acc_2_), .B(
        npu_inst_pe_1_7_6_add_69_carry_2_), .Z(npu_inst_pe_1_7_6_N75) );
  AND2_X1 npu_inst_pe_1_7_6_U137 ( .A1(npu_inst_pe_1_7_6_add_69_carry_2_), 
        .A2(npu_inst_pe_1_7_6_int_q_acc_2_), .ZN(
        npu_inst_pe_1_7_6_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_7_6_U136 ( .A(npu_inst_pe_1_7_6_int_q_acc_3_), .B(
        npu_inst_pe_1_7_6_add_69_carry_3_), .Z(npu_inst_pe_1_7_6_N76) );
  AND2_X1 npu_inst_pe_1_7_6_U135 ( .A1(npu_inst_pe_1_7_6_add_69_carry_3_), 
        .A2(npu_inst_pe_1_7_6_int_q_acc_3_), .ZN(
        npu_inst_pe_1_7_6_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_7_6_U134 ( .A(npu_inst_pe_1_7_6_int_q_acc_4_), .B(
        npu_inst_pe_1_7_6_add_69_carry_4_), .Z(npu_inst_pe_1_7_6_N77) );
  AND2_X1 npu_inst_pe_1_7_6_U133 ( .A1(npu_inst_pe_1_7_6_add_69_carry_4_), 
        .A2(npu_inst_pe_1_7_6_int_q_acc_4_), .ZN(
        npu_inst_pe_1_7_6_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_7_6_U132 ( .A(npu_inst_pe_1_7_6_int_q_acc_5_), .B(
        npu_inst_pe_1_7_6_add_69_carry_5_), .Z(npu_inst_pe_1_7_6_N78) );
  AND2_X1 npu_inst_pe_1_7_6_U131 ( .A1(npu_inst_pe_1_7_6_add_69_carry_5_), 
        .A2(npu_inst_pe_1_7_6_int_q_acc_5_), .ZN(
        npu_inst_pe_1_7_6_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_7_6_U130 ( .A(npu_inst_pe_1_7_6_int_q_acc_6_), .B(
        npu_inst_pe_1_7_6_add_69_carry_6_), .Z(npu_inst_pe_1_7_6_N79) );
  AND2_X1 npu_inst_pe_1_7_6_U129 ( .A1(npu_inst_pe_1_7_6_add_69_carry_6_), 
        .A2(npu_inst_pe_1_7_6_int_q_acc_6_), .ZN(
        npu_inst_pe_1_7_6_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_7_6_U128 ( .A(npu_inst_pe_1_7_6_int_q_acc_7_), .B(
        npu_inst_pe_1_7_6_add_69_carry_7_), .Z(npu_inst_pe_1_7_6_N80) );
  XNOR2_X1 npu_inst_pe_1_7_6_U127 ( .A(npu_inst_pe_1_7_6_sub_67_carry_2_), .B(
        npu_inst_pe_1_7_6_int_q_acc_2_), .ZN(npu_inst_pe_1_7_6_N67) );
  OR2_X1 npu_inst_pe_1_7_6_U126 ( .A1(npu_inst_pe_1_7_6_int_q_acc_2_), .A2(
        npu_inst_pe_1_7_6_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_7_6_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_7_6_U125 ( .A(npu_inst_pe_1_7_6_sub_67_carry_3_), .B(
        npu_inst_pe_1_7_6_int_q_acc_3_), .ZN(npu_inst_pe_1_7_6_N68) );
  OR2_X1 npu_inst_pe_1_7_6_U124 ( .A1(npu_inst_pe_1_7_6_int_q_acc_3_), .A2(
        npu_inst_pe_1_7_6_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_7_6_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_7_6_U123 ( .A(npu_inst_pe_1_7_6_sub_67_carry_4_), .B(
        npu_inst_pe_1_7_6_int_q_acc_4_), .ZN(npu_inst_pe_1_7_6_N69) );
  OR2_X1 npu_inst_pe_1_7_6_U122 ( .A1(npu_inst_pe_1_7_6_int_q_acc_4_), .A2(
        npu_inst_pe_1_7_6_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_7_6_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_7_6_U121 ( .A(npu_inst_pe_1_7_6_sub_67_carry_5_), .B(
        npu_inst_pe_1_7_6_int_q_acc_5_), .ZN(npu_inst_pe_1_7_6_N70) );
  OR2_X1 npu_inst_pe_1_7_6_U120 ( .A1(npu_inst_pe_1_7_6_int_q_acc_5_), .A2(
        npu_inst_pe_1_7_6_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_7_6_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_7_6_U119 ( .A(npu_inst_pe_1_7_6_sub_67_carry_6_), .B(
        npu_inst_pe_1_7_6_int_q_acc_6_), .ZN(npu_inst_pe_1_7_6_N71) );
  OR2_X1 npu_inst_pe_1_7_6_U118 ( .A1(npu_inst_pe_1_7_6_int_q_acc_6_), .A2(
        npu_inst_pe_1_7_6_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_7_6_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_7_6_U117 ( .A(npu_inst_pe_1_7_6_int_q_acc_7_), .B(
        npu_inst_pe_1_7_6_sub_67_carry_7_), .ZN(npu_inst_pe_1_7_6_N72) );
  INV_X1 npu_inst_pe_1_7_6_U116 ( .A(npu_inst_n75), .ZN(npu_inst_pe_1_7_6_n7)
         );
  INV_X1 npu_inst_pe_1_7_6_U115 ( .A(npu_inst_pe_1_7_6_n7), .ZN(
        npu_inst_pe_1_7_6_n6) );
  INV_X1 npu_inst_pe_1_7_6_U114 ( .A(npu_inst_n52), .ZN(npu_inst_pe_1_7_6_n3)
         );
  AOI22_X1 npu_inst_pe_1_7_6_U113 ( .A1(npu_inst_pe_1_7_6_n38), .A2(
        int_i_data_v_npu[3]), .B1(npu_inst_pe_1_7_6_n114), .B2(
        npu_inst_pe_1_7_6_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_7_6_n39) );
  INV_X1 npu_inst_pe_1_7_6_U112 ( .A(npu_inst_pe_1_7_6_n39), .ZN(
        npu_inst_pe_1_7_6_n112) );
  AOI22_X1 npu_inst_pe_1_7_6_U111 ( .A1(npu_inst_pe_1_7_6_n38), .A2(
        int_i_data_v_npu[2]), .B1(npu_inst_pe_1_7_6_n114), .B2(
        npu_inst_pe_1_7_6_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_7_6_n37) );
  INV_X1 npu_inst_pe_1_7_6_U110 ( .A(npu_inst_pe_1_7_6_n37), .ZN(
        npu_inst_pe_1_7_6_n113) );
  AOI22_X1 npu_inst_pe_1_7_6_U107 ( .A1(int_i_data_v_npu[3]), .A2(
        npu_inst_pe_1_7_6_n58), .B1(npu_inst_pe_1_7_6_n119), .B2(
        npu_inst_pe_1_7_6_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_7_6_n59) );
  INV_X1 npu_inst_pe_1_7_6_U106 ( .A(npu_inst_pe_1_7_6_n59), .ZN(
        npu_inst_pe_1_7_6_n102) );
  AOI22_X1 npu_inst_pe_1_7_6_U105 ( .A1(int_i_data_v_npu[2]), .A2(
        npu_inst_pe_1_7_6_n58), .B1(npu_inst_pe_1_7_6_n119), .B2(
        npu_inst_pe_1_7_6_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_7_6_n57) );
  INV_X1 npu_inst_pe_1_7_6_U104 ( .A(npu_inst_pe_1_7_6_n57), .ZN(
        npu_inst_pe_1_7_6_n103) );
  AOI22_X1 npu_inst_pe_1_7_6_U103 ( .A1(int_i_data_v_npu[3]), .A2(
        npu_inst_pe_1_7_6_n54), .B1(npu_inst_pe_1_7_6_n118), .B2(
        npu_inst_pe_1_7_6_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_7_6_n55) );
  INV_X1 npu_inst_pe_1_7_6_U102 ( .A(npu_inst_pe_1_7_6_n55), .ZN(
        npu_inst_pe_1_7_6_n104) );
  AOI22_X1 npu_inst_pe_1_7_6_U101 ( .A1(int_i_data_v_npu[2]), .A2(
        npu_inst_pe_1_7_6_n54), .B1(npu_inst_pe_1_7_6_n118), .B2(
        npu_inst_pe_1_7_6_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_7_6_n53) );
  INV_X1 npu_inst_pe_1_7_6_U100 ( .A(npu_inst_pe_1_7_6_n53), .ZN(
        npu_inst_pe_1_7_6_n105) );
  AOI22_X1 npu_inst_pe_1_7_6_U99 ( .A1(int_i_data_v_npu[3]), .A2(
        npu_inst_pe_1_7_6_n50), .B1(npu_inst_pe_1_7_6_n117), .B2(
        npu_inst_pe_1_7_6_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_7_6_n51) );
  INV_X1 npu_inst_pe_1_7_6_U98 ( .A(npu_inst_pe_1_7_6_n51), .ZN(
        npu_inst_pe_1_7_6_n106) );
  AOI22_X1 npu_inst_pe_1_7_6_U97 ( .A1(int_i_data_v_npu[2]), .A2(
        npu_inst_pe_1_7_6_n50), .B1(npu_inst_pe_1_7_6_n117), .B2(
        npu_inst_pe_1_7_6_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_7_6_n49) );
  INV_X1 npu_inst_pe_1_7_6_U96 ( .A(npu_inst_pe_1_7_6_n49), .ZN(
        npu_inst_pe_1_7_6_n107) );
  AOI22_X1 npu_inst_pe_1_7_6_U95 ( .A1(int_i_data_v_npu[3]), .A2(
        npu_inst_pe_1_7_6_n46), .B1(npu_inst_pe_1_7_6_n116), .B2(
        npu_inst_pe_1_7_6_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_7_6_n47) );
  INV_X1 npu_inst_pe_1_7_6_U94 ( .A(npu_inst_pe_1_7_6_n47), .ZN(
        npu_inst_pe_1_7_6_n108) );
  AOI22_X1 npu_inst_pe_1_7_6_U93 ( .A1(int_i_data_v_npu[2]), .A2(
        npu_inst_pe_1_7_6_n46), .B1(npu_inst_pe_1_7_6_n116), .B2(
        npu_inst_pe_1_7_6_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_7_6_n45) );
  INV_X1 npu_inst_pe_1_7_6_U92 ( .A(npu_inst_pe_1_7_6_n45), .ZN(
        npu_inst_pe_1_7_6_n109) );
  AOI22_X1 npu_inst_pe_1_7_6_U91 ( .A1(int_i_data_v_npu[3]), .A2(
        npu_inst_pe_1_7_6_n42), .B1(npu_inst_pe_1_7_6_n115), .B2(
        npu_inst_pe_1_7_6_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_7_6_n43) );
  INV_X1 npu_inst_pe_1_7_6_U90 ( .A(npu_inst_pe_1_7_6_n43), .ZN(
        npu_inst_pe_1_7_6_n110) );
  AOI22_X1 npu_inst_pe_1_7_6_U89 ( .A1(int_i_data_v_npu[2]), .A2(
        npu_inst_pe_1_7_6_n42), .B1(npu_inst_pe_1_7_6_n115), .B2(
        npu_inst_pe_1_7_6_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_7_6_n41) );
  INV_X1 npu_inst_pe_1_7_6_U88 ( .A(npu_inst_pe_1_7_6_n41), .ZN(
        npu_inst_pe_1_7_6_n111) );
  NAND2_X1 npu_inst_pe_1_7_6_U87 ( .A1(npu_inst_pe_1_7_6_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_7_6_n60), .ZN(npu_inst_pe_1_7_6_n74) );
  OAI21_X1 npu_inst_pe_1_7_6_U86 ( .B1(npu_inst_pe_1_7_6_n63), .B2(
        npu_inst_pe_1_7_6_n60), .A(npu_inst_pe_1_7_6_n74), .ZN(
        npu_inst_pe_1_7_6_n97) );
  NAND2_X1 npu_inst_pe_1_7_6_U85 ( .A1(npu_inst_pe_1_7_6_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_7_6_n60), .ZN(npu_inst_pe_1_7_6_n73) );
  OAI21_X1 npu_inst_pe_1_7_6_U84 ( .B1(npu_inst_pe_1_7_6_n61), .B2(
        npu_inst_pe_1_7_6_n60), .A(npu_inst_pe_1_7_6_n73), .ZN(
        npu_inst_pe_1_7_6_n96) );
  NAND2_X1 npu_inst_pe_1_7_6_U83 ( .A1(npu_inst_pe_1_7_6_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_7_6_n56), .ZN(npu_inst_pe_1_7_6_n72) );
  OAI21_X1 npu_inst_pe_1_7_6_U82 ( .B1(npu_inst_pe_1_7_6_n63), .B2(
        npu_inst_pe_1_7_6_n56), .A(npu_inst_pe_1_7_6_n72), .ZN(
        npu_inst_pe_1_7_6_n95) );
  NAND2_X1 npu_inst_pe_1_7_6_U81 ( .A1(npu_inst_pe_1_7_6_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_7_6_n56), .ZN(npu_inst_pe_1_7_6_n71) );
  OAI21_X1 npu_inst_pe_1_7_6_U80 ( .B1(npu_inst_pe_1_7_6_n61), .B2(
        npu_inst_pe_1_7_6_n56), .A(npu_inst_pe_1_7_6_n71), .ZN(
        npu_inst_pe_1_7_6_n94) );
  NAND2_X1 npu_inst_pe_1_7_6_U79 ( .A1(npu_inst_pe_1_7_6_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_7_6_n52), .ZN(npu_inst_pe_1_7_6_n70) );
  OAI21_X1 npu_inst_pe_1_7_6_U78 ( .B1(npu_inst_pe_1_7_6_n63), .B2(
        npu_inst_pe_1_7_6_n52), .A(npu_inst_pe_1_7_6_n70), .ZN(
        npu_inst_pe_1_7_6_n93) );
  NAND2_X1 npu_inst_pe_1_7_6_U77 ( .A1(npu_inst_pe_1_7_6_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_7_6_n52), .ZN(npu_inst_pe_1_7_6_n69) );
  OAI21_X1 npu_inst_pe_1_7_6_U76 ( .B1(npu_inst_pe_1_7_6_n61), .B2(
        npu_inst_pe_1_7_6_n52), .A(npu_inst_pe_1_7_6_n69), .ZN(
        npu_inst_pe_1_7_6_n92) );
  NAND2_X1 npu_inst_pe_1_7_6_U75 ( .A1(npu_inst_pe_1_7_6_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_7_6_n48), .ZN(npu_inst_pe_1_7_6_n68) );
  OAI21_X1 npu_inst_pe_1_7_6_U74 ( .B1(npu_inst_pe_1_7_6_n63), .B2(
        npu_inst_pe_1_7_6_n48), .A(npu_inst_pe_1_7_6_n68), .ZN(
        npu_inst_pe_1_7_6_n91) );
  NAND2_X1 npu_inst_pe_1_7_6_U73 ( .A1(npu_inst_pe_1_7_6_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_7_6_n48), .ZN(npu_inst_pe_1_7_6_n67) );
  OAI21_X1 npu_inst_pe_1_7_6_U72 ( .B1(npu_inst_pe_1_7_6_n61), .B2(
        npu_inst_pe_1_7_6_n48), .A(npu_inst_pe_1_7_6_n67), .ZN(
        npu_inst_pe_1_7_6_n90) );
  NAND2_X1 npu_inst_pe_1_7_6_U71 ( .A1(npu_inst_pe_1_7_6_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_7_6_n44), .ZN(npu_inst_pe_1_7_6_n66) );
  OAI21_X1 npu_inst_pe_1_7_6_U70 ( .B1(npu_inst_pe_1_7_6_n63), .B2(
        npu_inst_pe_1_7_6_n44), .A(npu_inst_pe_1_7_6_n66), .ZN(
        npu_inst_pe_1_7_6_n89) );
  NAND2_X1 npu_inst_pe_1_7_6_U69 ( .A1(npu_inst_pe_1_7_6_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_7_6_n44), .ZN(npu_inst_pe_1_7_6_n65) );
  OAI21_X1 npu_inst_pe_1_7_6_U68 ( .B1(npu_inst_pe_1_7_6_n61), .B2(
        npu_inst_pe_1_7_6_n44), .A(npu_inst_pe_1_7_6_n65), .ZN(
        npu_inst_pe_1_7_6_n88) );
  NAND2_X1 npu_inst_pe_1_7_6_U67 ( .A1(npu_inst_pe_1_7_6_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_7_6_n40), .ZN(npu_inst_pe_1_7_6_n64) );
  OAI21_X1 npu_inst_pe_1_7_6_U66 ( .B1(npu_inst_pe_1_7_6_n63), .B2(
        npu_inst_pe_1_7_6_n40), .A(npu_inst_pe_1_7_6_n64), .ZN(
        npu_inst_pe_1_7_6_n87) );
  NAND2_X1 npu_inst_pe_1_7_6_U65 ( .A1(npu_inst_pe_1_7_6_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_7_6_n40), .ZN(npu_inst_pe_1_7_6_n62) );
  OAI21_X1 npu_inst_pe_1_7_6_U64 ( .B1(npu_inst_pe_1_7_6_n61), .B2(
        npu_inst_pe_1_7_6_n40), .A(npu_inst_pe_1_7_6_n62), .ZN(
        npu_inst_pe_1_7_6_n86) );
  AND2_X1 npu_inst_pe_1_7_6_U63 ( .A1(npu_inst_pe_1_7_6_N93), .A2(npu_inst_n52), .ZN(npu_inst_int_data_y_7__6__0_) );
  AND2_X1 npu_inst_pe_1_7_6_U62 ( .A1(npu_inst_n52), .A2(npu_inst_pe_1_7_6_N94), .ZN(npu_inst_int_data_y_7__6__1_) );
  AOI22_X1 npu_inst_pe_1_7_6_U61 ( .A1(npu_inst_n52), .A2(int_i_data_v_npu[3]), 
        .B1(npu_inst_pe_1_7_6_n3), .B2(npu_inst_int_data_x_7__7__1_), .ZN(
        npu_inst_pe_1_7_6_n63) );
  AOI22_X1 npu_inst_pe_1_7_6_U60 ( .A1(npu_inst_n52), .A2(int_i_data_v_npu[2]), 
        .B1(npu_inst_pe_1_7_6_n3), .B2(npu_inst_int_data_x_7__7__0_), .ZN(
        npu_inst_pe_1_7_6_n61) );
  AOI222_X1 npu_inst_pe_1_7_6_U59 ( .A1(1'b0), .A2(npu_inst_pe_1_7_6_n1), .B1(
        npu_inst_pe_1_7_6_N73), .B2(npu_inst_pe_1_7_6_n76), .C1(
        npu_inst_pe_1_7_6_N65), .C2(npu_inst_pe_1_7_6_n77), .ZN(
        npu_inst_pe_1_7_6_n84) );
  INV_X1 npu_inst_pe_1_7_6_U58 ( .A(npu_inst_pe_1_7_6_n84), .ZN(
        npu_inst_pe_1_7_6_n101) );
  AOI222_X1 npu_inst_pe_1_7_6_U57 ( .A1(1'b0), .A2(npu_inst_pe_1_7_6_n1), .B1(
        npu_inst_pe_1_7_6_N80), .B2(npu_inst_pe_1_7_6_n76), .C1(
        npu_inst_pe_1_7_6_N72), .C2(npu_inst_pe_1_7_6_n77), .ZN(
        npu_inst_pe_1_7_6_n75) );
  INV_X1 npu_inst_pe_1_7_6_U56 ( .A(npu_inst_pe_1_7_6_n75), .ZN(
        npu_inst_pe_1_7_6_n33) );
  AOI222_X1 npu_inst_pe_1_7_6_U55 ( .A1(1'b0), .A2(npu_inst_pe_1_7_6_n1), .B1(
        npu_inst_pe_1_7_6_N74), .B2(npu_inst_pe_1_7_6_n76), .C1(
        npu_inst_pe_1_7_6_N66), .C2(npu_inst_pe_1_7_6_n77), .ZN(
        npu_inst_pe_1_7_6_n83) );
  INV_X1 npu_inst_pe_1_7_6_U54 ( .A(npu_inst_pe_1_7_6_n83), .ZN(
        npu_inst_pe_1_7_6_n100) );
  AOI222_X1 npu_inst_pe_1_7_6_U53 ( .A1(1'b0), .A2(npu_inst_pe_1_7_6_n1), .B1(
        npu_inst_pe_1_7_6_N75), .B2(npu_inst_pe_1_7_6_n76), .C1(
        npu_inst_pe_1_7_6_N67), .C2(npu_inst_pe_1_7_6_n77), .ZN(
        npu_inst_pe_1_7_6_n82) );
  INV_X1 npu_inst_pe_1_7_6_U52 ( .A(npu_inst_pe_1_7_6_n82), .ZN(
        npu_inst_pe_1_7_6_n99) );
  AOI222_X1 npu_inst_pe_1_7_6_U51 ( .A1(1'b0), .A2(npu_inst_pe_1_7_6_n1), .B1(
        npu_inst_pe_1_7_6_N76), .B2(npu_inst_pe_1_7_6_n76), .C1(
        npu_inst_pe_1_7_6_N68), .C2(npu_inst_pe_1_7_6_n77), .ZN(
        npu_inst_pe_1_7_6_n81) );
  INV_X1 npu_inst_pe_1_7_6_U50 ( .A(npu_inst_pe_1_7_6_n81), .ZN(
        npu_inst_pe_1_7_6_n98) );
  AOI222_X1 npu_inst_pe_1_7_6_U49 ( .A1(1'b0), .A2(npu_inst_pe_1_7_6_n1), .B1(
        npu_inst_pe_1_7_6_N77), .B2(npu_inst_pe_1_7_6_n76), .C1(
        npu_inst_pe_1_7_6_N69), .C2(npu_inst_pe_1_7_6_n77), .ZN(
        npu_inst_pe_1_7_6_n80) );
  INV_X1 npu_inst_pe_1_7_6_U48 ( .A(npu_inst_pe_1_7_6_n80), .ZN(
        npu_inst_pe_1_7_6_n36) );
  AOI222_X1 npu_inst_pe_1_7_6_U47 ( .A1(1'b0), .A2(npu_inst_pe_1_7_6_n1), .B1(
        npu_inst_pe_1_7_6_N78), .B2(npu_inst_pe_1_7_6_n76), .C1(
        npu_inst_pe_1_7_6_N70), .C2(npu_inst_pe_1_7_6_n77), .ZN(
        npu_inst_pe_1_7_6_n79) );
  INV_X1 npu_inst_pe_1_7_6_U46 ( .A(npu_inst_pe_1_7_6_n79), .ZN(
        npu_inst_pe_1_7_6_n35) );
  AOI222_X1 npu_inst_pe_1_7_6_U45 ( .A1(1'b0), .A2(npu_inst_pe_1_7_6_n1), .B1(
        npu_inst_pe_1_7_6_N79), .B2(npu_inst_pe_1_7_6_n76), .C1(
        npu_inst_pe_1_7_6_N71), .C2(npu_inst_pe_1_7_6_n77), .ZN(
        npu_inst_pe_1_7_6_n78) );
  INV_X1 npu_inst_pe_1_7_6_U44 ( .A(npu_inst_pe_1_7_6_n78), .ZN(
        npu_inst_pe_1_7_6_n34) );
  AND2_X1 npu_inst_pe_1_7_6_U43 ( .A1(npu_inst_pe_1_7_6_int_q_acc_0_), .A2(
        npu_inst_pe_1_7_6_n1), .ZN(npu_inst_int_data_res_7__6__0_) );
  AND2_X1 npu_inst_pe_1_7_6_U42 ( .A1(npu_inst_pe_1_7_6_n2), .A2(
        npu_inst_pe_1_7_6_int_q_acc_7_), .ZN(npu_inst_int_data_res_7__6__7_)
         );
  AND2_X1 npu_inst_pe_1_7_6_U41 ( .A1(npu_inst_pe_1_7_6_int_q_acc_1_), .A2(
        npu_inst_pe_1_7_6_n1), .ZN(npu_inst_int_data_res_7__6__1_) );
  AND2_X1 npu_inst_pe_1_7_6_U40 ( .A1(npu_inst_pe_1_7_6_int_q_acc_2_), .A2(
        npu_inst_pe_1_7_6_n1), .ZN(npu_inst_int_data_res_7__6__2_) );
  AND2_X1 npu_inst_pe_1_7_6_U39 ( .A1(npu_inst_pe_1_7_6_int_q_acc_3_), .A2(
        npu_inst_pe_1_7_6_n2), .ZN(npu_inst_int_data_res_7__6__3_) );
  AND2_X1 npu_inst_pe_1_7_6_U38 ( .A1(npu_inst_pe_1_7_6_int_q_acc_4_), .A2(
        npu_inst_pe_1_7_6_n2), .ZN(npu_inst_int_data_res_7__6__4_) );
  AND2_X1 npu_inst_pe_1_7_6_U37 ( .A1(npu_inst_pe_1_7_6_int_q_acc_5_), .A2(
        npu_inst_pe_1_7_6_n2), .ZN(npu_inst_int_data_res_7__6__5_) );
  AND2_X1 npu_inst_pe_1_7_6_U36 ( .A1(npu_inst_pe_1_7_6_int_q_acc_6_), .A2(
        npu_inst_pe_1_7_6_n2), .ZN(npu_inst_int_data_res_7__6__6_) );
  INV_X1 npu_inst_pe_1_7_6_U35 ( .A(npu_inst_pe_1_7_6_int_data_1_), .ZN(
        npu_inst_pe_1_7_6_n14) );
  NOR3_X1 npu_inst_pe_1_7_6_U34 ( .A1(npu_inst_pe_1_7_6_n26), .A2(npu_inst_n52), .A3(npu_inst_int_ckg[1]), .ZN(npu_inst_pe_1_7_6_n85) );
  OR2_X1 npu_inst_pe_1_7_6_U33 ( .A1(npu_inst_pe_1_7_6_n85), .A2(
        npu_inst_pe_1_7_6_n2), .ZN(npu_inst_pe_1_7_6_N84) );
  AND2_X1 npu_inst_pe_1_7_6_U32 ( .A1(npu_inst_int_data_x_7__6__1_), .A2(
        npu_inst_pe_1_7_6_int_q_weight_1_), .ZN(npu_inst_pe_1_7_6_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_7_6_U31 ( .A1(npu_inst_int_data_x_7__6__0_), .A2(
        npu_inst_pe_1_7_6_int_q_weight_1_), .ZN(npu_inst_pe_1_7_6_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_7_6_U30 ( .A(npu_inst_pe_1_7_6_int_data_0_), .ZN(
        npu_inst_pe_1_7_6_n13) );
  INV_X1 npu_inst_pe_1_7_6_U29 ( .A(npu_inst_n67), .ZN(npu_inst_pe_1_7_6_n5)
         );
  OR3_X1 npu_inst_pe_1_7_6_U28 ( .A1(npu_inst_pe_1_7_6_n6), .A2(
        npu_inst_pe_1_7_6_n8), .A3(npu_inst_pe_1_7_6_n5), .ZN(
        npu_inst_pe_1_7_6_n56) );
  OR3_X1 npu_inst_pe_1_7_6_U27 ( .A1(npu_inst_pe_1_7_6_n5), .A2(
        npu_inst_pe_1_7_6_n8), .A3(npu_inst_pe_1_7_6_n7), .ZN(
        npu_inst_pe_1_7_6_n48) );
  INV_X1 npu_inst_pe_1_7_6_U26 ( .A(npu_inst_pe_1_7_6_n5), .ZN(
        npu_inst_pe_1_7_6_n4) );
  OR3_X1 npu_inst_pe_1_7_6_U25 ( .A1(npu_inst_pe_1_7_6_n4), .A2(
        npu_inst_pe_1_7_6_n8), .A3(npu_inst_pe_1_7_6_n7), .ZN(
        npu_inst_pe_1_7_6_n52) );
  OR3_X1 npu_inst_pe_1_7_6_U24 ( .A1(npu_inst_pe_1_7_6_n6), .A2(
        npu_inst_pe_1_7_6_n8), .A3(npu_inst_pe_1_7_6_n4), .ZN(
        npu_inst_pe_1_7_6_n60) );
  NOR2_X1 npu_inst_pe_1_7_6_U23 ( .A1(npu_inst_pe_1_7_6_n60), .A2(
        npu_inst_pe_1_7_6_n3), .ZN(npu_inst_pe_1_7_6_n58) );
  NOR2_X1 npu_inst_pe_1_7_6_U22 ( .A1(npu_inst_pe_1_7_6_n56), .A2(
        npu_inst_pe_1_7_6_n3), .ZN(npu_inst_pe_1_7_6_n54) );
  NOR2_X1 npu_inst_pe_1_7_6_U21 ( .A1(npu_inst_pe_1_7_6_n52), .A2(
        npu_inst_pe_1_7_6_n3), .ZN(npu_inst_pe_1_7_6_n50) );
  NOR2_X1 npu_inst_pe_1_7_6_U20 ( .A1(npu_inst_pe_1_7_6_n48), .A2(
        npu_inst_pe_1_7_6_n3), .ZN(npu_inst_pe_1_7_6_n46) );
  NOR2_X1 npu_inst_pe_1_7_6_U19 ( .A1(npu_inst_pe_1_7_6_n40), .A2(
        npu_inst_pe_1_7_6_n3), .ZN(npu_inst_pe_1_7_6_n38) );
  NOR2_X1 npu_inst_pe_1_7_6_U18 ( .A1(npu_inst_pe_1_7_6_n44), .A2(
        npu_inst_pe_1_7_6_n3), .ZN(npu_inst_pe_1_7_6_n42) );
  BUF_X1 npu_inst_pe_1_7_6_U17 ( .A(npu_inst_n92), .Z(npu_inst_pe_1_7_6_n8) );
  INV_X1 npu_inst_pe_1_7_6_U16 ( .A(npu_inst_n122), .ZN(npu_inst_pe_1_7_6_n12)
         );
  INV_X1 npu_inst_pe_1_7_6_U15 ( .A(npu_inst_pe_1_7_6_n38), .ZN(
        npu_inst_pe_1_7_6_n114) );
  INV_X1 npu_inst_pe_1_7_6_U14 ( .A(npu_inst_pe_1_7_6_n58), .ZN(
        npu_inst_pe_1_7_6_n119) );
  INV_X1 npu_inst_pe_1_7_6_U13 ( .A(npu_inst_pe_1_7_6_n54), .ZN(
        npu_inst_pe_1_7_6_n118) );
  INV_X1 npu_inst_pe_1_7_6_U12 ( .A(npu_inst_pe_1_7_6_n50), .ZN(
        npu_inst_pe_1_7_6_n117) );
  INV_X1 npu_inst_pe_1_7_6_U11 ( .A(npu_inst_pe_1_7_6_n46), .ZN(
        npu_inst_pe_1_7_6_n116) );
  INV_X1 npu_inst_pe_1_7_6_U10 ( .A(npu_inst_pe_1_7_6_n42), .ZN(
        npu_inst_pe_1_7_6_n115) );
  BUF_X1 npu_inst_pe_1_7_6_U9 ( .A(npu_inst_n7), .Z(npu_inst_pe_1_7_6_n2) );
  BUF_X1 npu_inst_pe_1_7_6_U8 ( .A(npu_inst_n7), .Z(npu_inst_pe_1_7_6_n1) );
  BUF_X1 npu_inst_pe_1_7_6_U7 ( .A(npu_inst_pe_1_7_6_n12), .Z(
        npu_inst_pe_1_7_6_n11) );
  BUF_X1 npu_inst_pe_1_7_6_U6 ( .A(npu_inst_pe_1_7_6_n12), .Z(
        npu_inst_pe_1_7_6_n10) );
  BUF_X1 npu_inst_pe_1_7_6_U5 ( .A(npu_inst_pe_1_7_6_n12), .Z(
        npu_inst_pe_1_7_6_n9) );
  NOR2_X1 npu_inst_pe_1_7_6_U4 ( .A1(npu_inst_pe_1_7_6_int_q_weight_0_), .A2(
        npu_inst_pe_1_7_6_n1), .ZN(npu_inst_pe_1_7_6_n76) );
  NOR2_X1 npu_inst_pe_1_7_6_U3 ( .A1(npu_inst_pe_1_7_6_n27), .A2(
        npu_inst_pe_1_7_6_n1), .ZN(npu_inst_pe_1_7_6_n77) );
  FA_X1 npu_inst_pe_1_7_6_sub_67_U2_1 ( .A(npu_inst_pe_1_7_6_int_q_acc_1_), 
        .B(npu_inst_pe_1_7_6_n14), .CI(npu_inst_pe_1_7_6_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_7_6_sub_67_carry_2_), .S(npu_inst_pe_1_7_6_N66) );
  FA_X1 npu_inst_pe_1_7_6_add_69_U1_1 ( .A(npu_inst_pe_1_7_6_int_q_acc_1_), 
        .B(npu_inst_pe_1_7_6_int_data_1_), .CI(
        npu_inst_pe_1_7_6_add_69_carry_1_), .CO(
        npu_inst_pe_1_7_6_add_69_carry_2_), .S(npu_inst_pe_1_7_6_N74) );
  NAND3_X1 npu_inst_pe_1_7_6_U109 ( .A1(npu_inst_pe_1_7_6_n5), .A2(
        npu_inst_pe_1_7_6_n7), .A3(npu_inst_pe_1_7_6_n8), .ZN(
        npu_inst_pe_1_7_6_n44) );
  NAND3_X1 npu_inst_pe_1_7_6_U108 ( .A1(npu_inst_pe_1_7_6_n4), .A2(
        npu_inst_pe_1_7_6_n7), .A3(npu_inst_pe_1_7_6_n8), .ZN(
        npu_inst_pe_1_7_6_n40) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_7_6_n34), .CK(
        npu_inst_pe_1_7_6_net3136), .RN(npu_inst_pe_1_7_6_n9), .Q(
        npu_inst_pe_1_7_6_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_7_6_n35), .CK(
        npu_inst_pe_1_7_6_net3136), .RN(npu_inst_pe_1_7_6_n9), .Q(
        npu_inst_pe_1_7_6_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_7_6_n36), .CK(
        npu_inst_pe_1_7_6_net3136), .RN(npu_inst_pe_1_7_6_n9), .Q(
        npu_inst_pe_1_7_6_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_7_6_n98), .CK(
        npu_inst_pe_1_7_6_net3136), .RN(npu_inst_pe_1_7_6_n9), .Q(
        npu_inst_pe_1_7_6_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_7_6_n99), .CK(
        npu_inst_pe_1_7_6_net3136), .RN(npu_inst_pe_1_7_6_n9), .Q(
        npu_inst_pe_1_7_6_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_7_6_n100), 
        .CK(npu_inst_pe_1_7_6_net3136), .RN(npu_inst_pe_1_7_6_n9), .Q(
        npu_inst_pe_1_7_6_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_7_6_n33), .CK(
        npu_inst_pe_1_7_6_net3136), .RN(npu_inst_pe_1_7_6_n9), .Q(
        npu_inst_pe_1_7_6_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_7_6_n101), 
        .CK(npu_inst_pe_1_7_6_net3136), .RN(npu_inst_pe_1_7_6_n9), .Q(
        npu_inst_pe_1_7_6_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_weight_reg_0_ ( .D(npu_inst_n108), .CK(
        npu_inst_pe_1_7_6_net3142), .RN(npu_inst_pe_1_7_6_n9), .Q(
        npu_inst_pe_1_7_6_int_q_weight_0_), .QN(npu_inst_pe_1_7_6_n27) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_weight_reg_1_ ( .D(npu_inst_n114), .CK(
        npu_inst_pe_1_7_6_net3142), .RN(npu_inst_pe_1_7_6_n9), .Q(
        npu_inst_pe_1_7_6_int_q_weight_1_), .QN(npu_inst_pe_1_7_6_n26) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_7_6_n113), 
        .CK(npu_inst_pe_1_7_6_net3142), .RN(npu_inst_pe_1_7_6_n9), .Q(
        npu_inst_pe_1_7_6_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_7_6_n112), 
        .CK(npu_inst_pe_1_7_6_net3142), .RN(npu_inst_pe_1_7_6_n9), .Q(
        npu_inst_pe_1_7_6_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_7_6_n111), 
        .CK(npu_inst_pe_1_7_6_net3142), .RN(npu_inst_pe_1_7_6_n10), .Q(
        npu_inst_pe_1_7_6_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_7_6_n110), 
        .CK(npu_inst_pe_1_7_6_net3142), .RN(npu_inst_pe_1_7_6_n10), .Q(
        npu_inst_pe_1_7_6_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_7_6_n109), 
        .CK(npu_inst_pe_1_7_6_net3142), .RN(npu_inst_pe_1_7_6_n10), .Q(
        npu_inst_pe_1_7_6_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_7_6_n108), 
        .CK(npu_inst_pe_1_7_6_net3142), .RN(npu_inst_pe_1_7_6_n10), .Q(
        npu_inst_pe_1_7_6_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_7_6_n107), 
        .CK(npu_inst_pe_1_7_6_net3142), .RN(npu_inst_pe_1_7_6_n10), .Q(
        npu_inst_pe_1_7_6_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_7_6_n106), 
        .CK(npu_inst_pe_1_7_6_net3142), .RN(npu_inst_pe_1_7_6_n10), .Q(
        npu_inst_pe_1_7_6_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_7_6_n105), 
        .CK(npu_inst_pe_1_7_6_net3142), .RN(npu_inst_pe_1_7_6_n10), .Q(
        npu_inst_pe_1_7_6_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_7_6_n104), 
        .CK(npu_inst_pe_1_7_6_net3142), .RN(npu_inst_pe_1_7_6_n10), .Q(
        npu_inst_pe_1_7_6_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_7_6_n103), 
        .CK(npu_inst_pe_1_7_6_net3142), .RN(npu_inst_pe_1_7_6_n10), .Q(
        npu_inst_pe_1_7_6_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_7_6_n102), 
        .CK(npu_inst_pe_1_7_6_net3142), .RN(npu_inst_pe_1_7_6_n10), .Q(
        npu_inst_pe_1_7_6_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_7_6_n86), 
        .CK(npu_inst_pe_1_7_6_net3142), .RN(npu_inst_pe_1_7_6_n10), .Q(
        npu_inst_pe_1_7_6_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_7_6_n87), 
        .CK(npu_inst_pe_1_7_6_net3142), .RN(npu_inst_pe_1_7_6_n10), .Q(
        npu_inst_pe_1_7_6_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_7_6_n88), 
        .CK(npu_inst_pe_1_7_6_net3142), .RN(npu_inst_pe_1_7_6_n11), .Q(
        npu_inst_pe_1_7_6_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_7_6_n89), 
        .CK(npu_inst_pe_1_7_6_net3142), .RN(npu_inst_pe_1_7_6_n11), .Q(
        npu_inst_pe_1_7_6_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_7_6_n90), 
        .CK(npu_inst_pe_1_7_6_net3142), .RN(npu_inst_pe_1_7_6_n11), .Q(
        npu_inst_pe_1_7_6_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_7_6_n91), 
        .CK(npu_inst_pe_1_7_6_net3142), .RN(npu_inst_pe_1_7_6_n11), .Q(
        npu_inst_pe_1_7_6_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_7_6_n92), 
        .CK(npu_inst_pe_1_7_6_net3142), .RN(npu_inst_pe_1_7_6_n11), .Q(
        npu_inst_pe_1_7_6_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_7_6_n93), 
        .CK(npu_inst_pe_1_7_6_net3142), .RN(npu_inst_pe_1_7_6_n11), .Q(
        npu_inst_pe_1_7_6_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_7_6_n94), 
        .CK(npu_inst_pe_1_7_6_net3142), .RN(npu_inst_pe_1_7_6_n11), .Q(
        npu_inst_pe_1_7_6_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_7_6_n95), 
        .CK(npu_inst_pe_1_7_6_net3142), .RN(npu_inst_pe_1_7_6_n11), .Q(
        npu_inst_pe_1_7_6_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_7_6_n96), 
        .CK(npu_inst_pe_1_7_6_net3142), .RN(npu_inst_pe_1_7_6_n11), .Q(
        npu_inst_pe_1_7_6_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_7_6_n97), 
        .CK(npu_inst_pe_1_7_6_net3142), .RN(npu_inst_pe_1_7_6_n11), .Q(
        npu_inst_pe_1_7_6_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_7_6_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_7_6_N84), .SE(1'b0), .GCK(npu_inst_pe_1_7_6_net3136) );
  CLKGATETST_X1 npu_inst_pe_1_7_6_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n61), .SE(1'b0), .GCK(npu_inst_pe_1_7_6_net3142) );
  MUX2_X1 npu_inst_pe_1_7_7_U162 ( .A(npu_inst_pe_1_7_7_n32), .B(
        npu_inst_pe_1_7_7_n29), .S(npu_inst_pe_1_7_7_n8), .Z(
        npu_inst_pe_1_7_7_N93) );
  MUX2_X1 npu_inst_pe_1_7_7_U161 ( .A(npu_inst_pe_1_7_7_n31), .B(
        npu_inst_pe_1_7_7_n30), .S(npu_inst_pe_1_7_7_n6), .Z(
        npu_inst_pe_1_7_7_n32) );
  MUX2_X1 npu_inst_pe_1_7_7_U160 ( .A(npu_inst_pe_1_7_7_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_7_7_int_q_reg_v_1__0_), .S(npu_inst_pe_1_7_7_n4), .Z(
        npu_inst_pe_1_7_7_n31) );
  MUX2_X1 npu_inst_pe_1_7_7_U159 ( .A(npu_inst_pe_1_7_7_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_7_7_int_q_reg_v_3__0_), .S(npu_inst_pe_1_7_7_n4), .Z(
        npu_inst_pe_1_7_7_n30) );
  MUX2_X1 npu_inst_pe_1_7_7_U158 ( .A(npu_inst_pe_1_7_7_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_7_7_int_q_reg_v_5__0_), .S(npu_inst_pe_1_7_7_n4), .Z(
        npu_inst_pe_1_7_7_n29) );
  MUX2_X1 npu_inst_pe_1_7_7_U157 ( .A(npu_inst_pe_1_7_7_n28), .B(
        npu_inst_pe_1_7_7_n23), .S(npu_inst_pe_1_7_7_n8), .Z(
        npu_inst_pe_1_7_7_N94) );
  MUX2_X1 npu_inst_pe_1_7_7_U156 ( .A(npu_inst_pe_1_7_7_n25), .B(
        npu_inst_pe_1_7_7_n24), .S(npu_inst_pe_1_7_7_n6), .Z(
        npu_inst_pe_1_7_7_n28) );
  MUX2_X1 npu_inst_pe_1_7_7_U155 ( .A(npu_inst_pe_1_7_7_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_7_7_int_q_reg_v_1__1_), .S(npu_inst_pe_1_7_7_n4), .Z(
        npu_inst_pe_1_7_7_n25) );
  MUX2_X1 npu_inst_pe_1_7_7_U154 ( .A(npu_inst_pe_1_7_7_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_7_7_int_q_reg_v_3__1_), .S(npu_inst_pe_1_7_7_n4), .Z(
        npu_inst_pe_1_7_7_n24) );
  MUX2_X1 npu_inst_pe_1_7_7_U153 ( .A(npu_inst_pe_1_7_7_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_7_7_int_q_reg_v_5__1_), .S(npu_inst_pe_1_7_7_n4), .Z(
        npu_inst_pe_1_7_7_n23) );
  MUX2_X1 npu_inst_pe_1_7_7_U152 ( .A(npu_inst_pe_1_7_7_n22), .B(
        npu_inst_pe_1_7_7_n19), .S(npu_inst_pe_1_7_7_n8), .Z(
        npu_inst_int_data_x_7__7__1_) );
  MUX2_X1 npu_inst_pe_1_7_7_U151 ( .A(npu_inst_pe_1_7_7_n21), .B(
        npu_inst_pe_1_7_7_n20), .S(npu_inst_pe_1_7_7_n6), .Z(
        npu_inst_pe_1_7_7_n22) );
  MUX2_X1 npu_inst_pe_1_7_7_U150 ( .A(npu_inst_pe_1_7_7_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_7_7_int_q_reg_h_1__1_), .S(npu_inst_pe_1_7_7_n4), .Z(
        npu_inst_pe_1_7_7_n21) );
  MUX2_X1 npu_inst_pe_1_7_7_U149 ( .A(npu_inst_pe_1_7_7_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_7_7_int_q_reg_h_3__1_), .S(npu_inst_pe_1_7_7_n4), .Z(
        npu_inst_pe_1_7_7_n20) );
  MUX2_X1 npu_inst_pe_1_7_7_U148 ( .A(npu_inst_pe_1_7_7_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_7_7_int_q_reg_h_5__1_), .S(npu_inst_pe_1_7_7_n4), .Z(
        npu_inst_pe_1_7_7_n19) );
  MUX2_X1 npu_inst_pe_1_7_7_U147 ( .A(npu_inst_pe_1_7_7_n18), .B(
        npu_inst_pe_1_7_7_n15), .S(npu_inst_pe_1_7_7_n8), .Z(
        npu_inst_int_data_x_7__7__0_) );
  MUX2_X1 npu_inst_pe_1_7_7_U146 ( .A(npu_inst_pe_1_7_7_n17), .B(
        npu_inst_pe_1_7_7_n16), .S(npu_inst_pe_1_7_7_n6), .Z(
        npu_inst_pe_1_7_7_n18) );
  MUX2_X1 npu_inst_pe_1_7_7_U145 ( .A(npu_inst_pe_1_7_7_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_7_7_int_q_reg_h_1__0_), .S(npu_inst_pe_1_7_7_n4), .Z(
        npu_inst_pe_1_7_7_n17) );
  MUX2_X1 npu_inst_pe_1_7_7_U144 ( .A(npu_inst_pe_1_7_7_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_7_7_int_q_reg_h_3__0_), .S(npu_inst_pe_1_7_7_n4), .Z(
        npu_inst_pe_1_7_7_n16) );
  MUX2_X1 npu_inst_pe_1_7_7_U143 ( .A(npu_inst_pe_1_7_7_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_7_7_int_q_reg_h_5__0_), .S(npu_inst_pe_1_7_7_n4), .Z(
        npu_inst_pe_1_7_7_n15) );
  XOR2_X1 npu_inst_pe_1_7_7_U142 ( .A(npu_inst_pe_1_7_7_int_data_0_), .B(
        npu_inst_pe_1_7_7_int_q_acc_0_), .Z(npu_inst_pe_1_7_7_N73) );
  AND2_X1 npu_inst_pe_1_7_7_U141 ( .A1(npu_inst_pe_1_7_7_int_q_acc_0_), .A2(
        npu_inst_pe_1_7_7_int_data_0_), .ZN(npu_inst_pe_1_7_7_add_69_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_7_7_U140 ( .A(npu_inst_pe_1_7_7_int_q_acc_0_), .B(
        npu_inst_pe_1_7_7_n13), .ZN(npu_inst_pe_1_7_7_N65) );
  OR2_X1 npu_inst_pe_1_7_7_U139 ( .A1(npu_inst_pe_1_7_7_n13), .A2(
        npu_inst_pe_1_7_7_int_q_acc_0_), .ZN(npu_inst_pe_1_7_7_sub_67_carry_1_) );
  XOR2_X1 npu_inst_pe_1_7_7_U138 ( .A(npu_inst_pe_1_7_7_int_q_acc_2_), .B(
        npu_inst_pe_1_7_7_add_69_carry_2_), .Z(npu_inst_pe_1_7_7_N75) );
  AND2_X1 npu_inst_pe_1_7_7_U137 ( .A1(npu_inst_pe_1_7_7_add_69_carry_2_), 
        .A2(npu_inst_pe_1_7_7_int_q_acc_2_), .ZN(
        npu_inst_pe_1_7_7_add_69_carry_3_) );
  XOR2_X1 npu_inst_pe_1_7_7_U136 ( .A(npu_inst_pe_1_7_7_int_q_acc_3_), .B(
        npu_inst_pe_1_7_7_add_69_carry_3_), .Z(npu_inst_pe_1_7_7_N76) );
  AND2_X1 npu_inst_pe_1_7_7_U135 ( .A1(npu_inst_pe_1_7_7_add_69_carry_3_), 
        .A2(npu_inst_pe_1_7_7_int_q_acc_3_), .ZN(
        npu_inst_pe_1_7_7_add_69_carry_4_) );
  XOR2_X1 npu_inst_pe_1_7_7_U134 ( .A(npu_inst_pe_1_7_7_int_q_acc_4_), .B(
        npu_inst_pe_1_7_7_add_69_carry_4_), .Z(npu_inst_pe_1_7_7_N77) );
  AND2_X1 npu_inst_pe_1_7_7_U133 ( .A1(npu_inst_pe_1_7_7_add_69_carry_4_), 
        .A2(npu_inst_pe_1_7_7_int_q_acc_4_), .ZN(
        npu_inst_pe_1_7_7_add_69_carry_5_) );
  XOR2_X1 npu_inst_pe_1_7_7_U132 ( .A(npu_inst_pe_1_7_7_int_q_acc_5_), .B(
        npu_inst_pe_1_7_7_add_69_carry_5_), .Z(npu_inst_pe_1_7_7_N78) );
  AND2_X1 npu_inst_pe_1_7_7_U131 ( .A1(npu_inst_pe_1_7_7_add_69_carry_5_), 
        .A2(npu_inst_pe_1_7_7_int_q_acc_5_), .ZN(
        npu_inst_pe_1_7_7_add_69_carry_6_) );
  XOR2_X1 npu_inst_pe_1_7_7_U130 ( .A(npu_inst_pe_1_7_7_int_q_acc_6_), .B(
        npu_inst_pe_1_7_7_add_69_carry_6_), .Z(npu_inst_pe_1_7_7_N79) );
  AND2_X1 npu_inst_pe_1_7_7_U129 ( .A1(npu_inst_pe_1_7_7_add_69_carry_6_), 
        .A2(npu_inst_pe_1_7_7_int_q_acc_6_), .ZN(
        npu_inst_pe_1_7_7_add_69_carry_7_) );
  XOR2_X1 npu_inst_pe_1_7_7_U128 ( .A(npu_inst_pe_1_7_7_int_q_acc_7_), .B(
        npu_inst_pe_1_7_7_add_69_carry_7_), .Z(npu_inst_pe_1_7_7_N80) );
  XNOR2_X1 npu_inst_pe_1_7_7_U127 ( .A(npu_inst_pe_1_7_7_sub_67_carry_2_), .B(
        npu_inst_pe_1_7_7_int_q_acc_2_), .ZN(npu_inst_pe_1_7_7_N67) );
  OR2_X1 npu_inst_pe_1_7_7_U126 ( .A1(npu_inst_pe_1_7_7_int_q_acc_2_), .A2(
        npu_inst_pe_1_7_7_sub_67_carry_2_), .ZN(
        npu_inst_pe_1_7_7_sub_67_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_7_7_U125 ( .A(npu_inst_pe_1_7_7_sub_67_carry_3_), .B(
        npu_inst_pe_1_7_7_int_q_acc_3_), .ZN(npu_inst_pe_1_7_7_N68) );
  OR2_X1 npu_inst_pe_1_7_7_U124 ( .A1(npu_inst_pe_1_7_7_int_q_acc_3_), .A2(
        npu_inst_pe_1_7_7_sub_67_carry_3_), .ZN(
        npu_inst_pe_1_7_7_sub_67_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_7_7_U123 ( .A(npu_inst_pe_1_7_7_sub_67_carry_4_), .B(
        npu_inst_pe_1_7_7_int_q_acc_4_), .ZN(npu_inst_pe_1_7_7_N69) );
  OR2_X1 npu_inst_pe_1_7_7_U122 ( .A1(npu_inst_pe_1_7_7_int_q_acc_4_), .A2(
        npu_inst_pe_1_7_7_sub_67_carry_4_), .ZN(
        npu_inst_pe_1_7_7_sub_67_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_7_7_U121 ( .A(npu_inst_pe_1_7_7_sub_67_carry_5_), .B(
        npu_inst_pe_1_7_7_int_q_acc_5_), .ZN(npu_inst_pe_1_7_7_N70) );
  OR2_X1 npu_inst_pe_1_7_7_U120 ( .A1(npu_inst_pe_1_7_7_int_q_acc_5_), .A2(
        npu_inst_pe_1_7_7_sub_67_carry_5_), .ZN(
        npu_inst_pe_1_7_7_sub_67_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_7_7_U119 ( .A(npu_inst_pe_1_7_7_sub_67_carry_6_), .B(
        npu_inst_pe_1_7_7_int_q_acc_6_), .ZN(npu_inst_pe_1_7_7_N71) );
  OR2_X1 npu_inst_pe_1_7_7_U118 ( .A1(npu_inst_pe_1_7_7_int_q_acc_6_), .A2(
        npu_inst_pe_1_7_7_sub_67_carry_6_), .ZN(
        npu_inst_pe_1_7_7_sub_67_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_7_7_U117 ( .A(npu_inst_pe_1_7_7_int_q_acc_7_), .B(
        npu_inst_pe_1_7_7_sub_67_carry_7_), .ZN(npu_inst_pe_1_7_7_N72) );
  INV_X1 npu_inst_pe_1_7_7_U116 ( .A(npu_inst_n75), .ZN(npu_inst_pe_1_7_7_n7)
         );
  INV_X1 npu_inst_pe_1_7_7_U115 ( .A(npu_inst_pe_1_7_7_n7), .ZN(
        npu_inst_pe_1_7_7_n6) );
  INV_X1 npu_inst_pe_1_7_7_U114 ( .A(npu_inst_n52), .ZN(npu_inst_pe_1_7_7_n3)
         );
  AOI22_X1 npu_inst_pe_1_7_7_U113 ( .A1(npu_inst_pe_1_7_7_n38), .A2(
        int_i_data_v_npu[1]), .B1(npu_inst_pe_1_7_7_n114), .B2(
        npu_inst_pe_1_7_7_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_7_7_n39) );
  INV_X1 npu_inst_pe_1_7_7_U112 ( .A(npu_inst_pe_1_7_7_n39), .ZN(
        npu_inst_pe_1_7_7_n112) );
  AOI22_X1 npu_inst_pe_1_7_7_U111 ( .A1(npu_inst_pe_1_7_7_n38), .A2(
        int_i_data_v_npu[0]), .B1(npu_inst_pe_1_7_7_n114), .B2(
        npu_inst_pe_1_7_7_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_7_7_n37) );
  INV_X1 npu_inst_pe_1_7_7_U110 ( .A(npu_inst_pe_1_7_7_n37), .ZN(
        npu_inst_pe_1_7_7_n113) );
  AOI22_X1 npu_inst_pe_1_7_7_U107 ( .A1(int_i_data_v_npu[1]), .A2(
        npu_inst_pe_1_7_7_n58), .B1(npu_inst_pe_1_7_7_n119), .B2(
        npu_inst_pe_1_7_7_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_7_7_n59) );
  INV_X1 npu_inst_pe_1_7_7_U106 ( .A(npu_inst_pe_1_7_7_n59), .ZN(
        npu_inst_pe_1_7_7_n102) );
  AOI22_X1 npu_inst_pe_1_7_7_U105 ( .A1(int_i_data_v_npu[0]), .A2(
        npu_inst_pe_1_7_7_n58), .B1(npu_inst_pe_1_7_7_n119), .B2(
        npu_inst_pe_1_7_7_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_7_7_n57) );
  INV_X1 npu_inst_pe_1_7_7_U104 ( .A(npu_inst_pe_1_7_7_n57), .ZN(
        npu_inst_pe_1_7_7_n103) );
  AOI22_X1 npu_inst_pe_1_7_7_U103 ( .A1(int_i_data_v_npu[1]), .A2(
        npu_inst_pe_1_7_7_n54), .B1(npu_inst_pe_1_7_7_n118), .B2(
        npu_inst_pe_1_7_7_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_7_7_n55) );
  INV_X1 npu_inst_pe_1_7_7_U102 ( .A(npu_inst_pe_1_7_7_n55), .ZN(
        npu_inst_pe_1_7_7_n104) );
  AOI22_X1 npu_inst_pe_1_7_7_U101 ( .A1(int_i_data_v_npu[0]), .A2(
        npu_inst_pe_1_7_7_n54), .B1(npu_inst_pe_1_7_7_n118), .B2(
        npu_inst_pe_1_7_7_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_7_7_n53) );
  INV_X1 npu_inst_pe_1_7_7_U100 ( .A(npu_inst_pe_1_7_7_n53), .ZN(
        npu_inst_pe_1_7_7_n105) );
  AOI22_X1 npu_inst_pe_1_7_7_U99 ( .A1(int_i_data_v_npu[1]), .A2(
        npu_inst_pe_1_7_7_n50), .B1(npu_inst_pe_1_7_7_n117), .B2(
        npu_inst_pe_1_7_7_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_7_7_n51) );
  INV_X1 npu_inst_pe_1_7_7_U98 ( .A(npu_inst_pe_1_7_7_n51), .ZN(
        npu_inst_pe_1_7_7_n106) );
  AOI22_X1 npu_inst_pe_1_7_7_U97 ( .A1(int_i_data_v_npu[0]), .A2(
        npu_inst_pe_1_7_7_n50), .B1(npu_inst_pe_1_7_7_n117), .B2(
        npu_inst_pe_1_7_7_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_7_7_n49) );
  INV_X1 npu_inst_pe_1_7_7_U96 ( .A(npu_inst_pe_1_7_7_n49), .ZN(
        npu_inst_pe_1_7_7_n107) );
  AOI22_X1 npu_inst_pe_1_7_7_U95 ( .A1(int_i_data_v_npu[1]), .A2(
        npu_inst_pe_1_7_7_n46), .B1(npu_inst_pe_1_7_7_n116), .B2(
        npu_inst_pe_1_7_7_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_7_7_n47) );
  INV_X1 npu_inst_pe_1_7_7_U94 ( .A(npu_inst_pe_1_7_7_n47), .ZN(
        npu_inst_pe_1_7_7_n108) );
  AOI22_X1 npu_inst_pe_1_7_7_U93 ( .A1(int_i_data_v_npu[0]), .A2(
        npu_inst_pe_1_7_7_n46), .B1(npu_inst_pe_1_7_7_n116), .B2(
        npu_inst_pe_1_7_7_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_7_7_n45) );
  INV_X1 npu_inst_pe_1_7_7_U92 ( .A(npu_inst_pe_1_7_7_n45), .ZN(
        npu_inst_pe_1_7_7_n109) );
  AOI22_X1 npu_inst_pe_1_7_7_U91 ( .A1(int_i_data_v_npu[1]), .A2(
        npu_inst_pe_1_7_7_n42), .B1(npu_inst_pe_1_7_7_n115), .B2(
        npu_inst_pe_1_7_7_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_7_7_n43) );
  INV_X1 npu_inst_pe_1_7_7_U90 ( .A(npu_inst_pe_1_7_7_n43), .ZN(
        npu_inst_pe_1_7_7_n110) );
  AOI22_X1 npu_inst_pe_1_7_7_U89 ( .A1(int_i_data_v_npu[0]), .A2(
        npu_inst_pe_1_7_7_n42), .B1(npu_inst_pe_1_7_7_n115), .B2(
        npu_inst_pe_1_7_7_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_7_7_n41) );
  INV_X1 npu_inst_pe_1_7_7_U88 ( .A(npu_inst_pe_1_7_7_n41), .ZN(
        npu_inst_pe_1_7_7_n111) );
  AND2_X1 npu_inst_pe_1_7_7_U87 ( .A1(npu_inst_pe_1_7_7_N93), .A2(npu_inst_n52), .ZN(npu_inst_int_data_y_7__7__0_) );
  AND2_X1 npu_inst_pe_1_7_7_U86 ( .A1(npu_inst_n52), .A2(npu_inst_pe_1_7_7_N94), .ZN(npu_inst_int_data_y_7__7__1_) );
  NOR3_X1 npu_inst_pe_1_7_7_U85 ( .A1(npu_inst_pe_1_7_7_n26), .A2(npu_inst_n52), .A3(npu_inst_int_ckg[0]), .ZN(npu_inst_pe_1_7_7_n85) );
  OR2_X1 npu_inst_pe_1_7_7_U84 ( .A1(npu_inst_pe_1_7_7_n85), .A2(
        npu_inst_pe_1_7_7_n2), .ZN(npu_inst_pe_1_7_7_N84) );
  AOI222_X1 npu_inst_pe_1_7_7_U83 ( .A1(1'b0), .A2(npu_inst_pe_1_7_7_n1), .B1(
        npu_inst_pe_1_7_7_N73), .B2(npu_inst_pe_1_7_7_n76), .C1(
        npu_inst_pe_1_7_7_N65), .C2(npu_inst_pe_1_7_7_n77), .ZN(
        npu_inst_pe_1_7_7_n84) );
  INV_X1 npu_inst_pe_1_7_7_U82 ( .A(npu_inst_pe_1_7_7_n84), .ZN(
        npu_inst_pe_1_7_7_n101) );
  AOI222_X1 npu_inst_pe_1_7_7_U81 ( .A1(1'b0), .A2(npu_inst_pe_1_7_7_n1), .B1(
        npu_inst_pe_1_7_7_N80), .B2(npu_inst_pe_1_7_7_n76), .C1(
        npu_inst_pe_1_7_7_N72), .C2(npu_inst_pe_1_7_7_n77), .ZN(
        npu_inst_pe_1_7_7_n75) );
  INV_X1 npu_inst_pe_1_7_7_U80 ( .A(npu_inst_pe_1_7_7_n75), .ZN(
        npu_inst_pe_1_7_7_n33) );
  AOI222_X1 npu_inst_pe_1_7_7_U79 ( .A1(1'b0), .A2(npu_inst_pe_1_7_7_n1), .B1(
        npu_inst_pe_1_7_7_N74), .B2(npu_inst_pe_1_7_7_n76), .C1(
        npu_inst_pe_1_7_7_N66), .C2(npu_inst_pe_1_7_7_n77), .ZN(
        npu_inst_pe_1_7_7_n83) );
  INV_X1 npu_inst_pe_1_7_7_U78 ( .A(npu_inst_pe_1_7_7_n83), .ZN(
        npu_inst_pe_1_7_7_n100) );
  AOI222_X1 npu_inst_pe_1_7_7_U77 ( .A1(1'b0), .A2(npu_inst_pe_1_7_7_n1), .B1(
        npu_inst_pe_1_7_7_N75), .B2(npu_inst_pe_1_7_7_n76), .C1(
        npu_inst_pe_1_7_7_N67), .C2(npu_inst_pe_1_7_7_n77), .ZN(
        npu_inst_pe_1_7_7_n82) );
  INV_X1 npu_inst_pe_1_7_7_U76 ( .A(npu_inst_pe_1_7_7_n82), .ZN(
        npu_inst_pe_1_7_7_n99) );
  AOI222_X1 npu_inst_pe_1_7_7_U75 ( .A1(1'b0), .A2(npu_inst_pe_1_7_7_n1), .B1(
        npu_inst_pe_1_7_7_N76), .B2(npu_inst_pe_1_7_7_n76), .C1(
        npu_inst_pe_1_7_7_N68), .C2(npu_inst_pe_1_7_7_n77), .ZN(
        npu_inst_pe_1_7_7_n81) );
  INV_X1 npu_inst_pe_1_7_7_U74 ( .A(npu_inst_pe_1_7_7_n81), .ZN(
        npu_inst_pe_1_7_7_n98) );
  AOI222_X1 npu_inst_pe_1_7_7_U73 ( .A1(1'b0), .A2(npu_inst_pe_1_7_7_n1), .B1(
        npu_inst_pe_1_7_7_N77), .B2(npu_inst_pe_1_7_7_n76), .C1(
        npu_inst_pe_1_7_7_N69), .C2(npu_inst_pe_1_7_7_n77), .ZN(
        npu_inst_pe_1_7_7_n80) );
  INV_X1 npu_inst_pe_1_7_7_U72 ( .A(npu_inst_pe_1_7_7_n80), .ZN(
        npu_inst_pe_1_7_7_n36) );
  AOI222_X1 npu_inst_pe_1_7_7_U71 ( .A1(1'b0), .A2(npu_inst_pe_1_7_7_n1), .B1(
        npu_inst_pe_1_7_7_N78), .B2(npu_inst_pe_1_7_7_n76), .C1(
        npu_inst_pe_1_7_7_N70), .C2(npu_inst_pe_1_7_7_n77), .ZN(
        npu_inst_pe_1_7_7_n79) );
  INV_X1 npu_inst_pe_1_7_7_U70 ( .A(npu_inst_pe_1_7_7_n79), .ZN(
        npu_inst_pe_1_7_7_n35) );
  AOI222_X1 npu_inst_pe_1_7_7_U69 ( .A1(1'b0), .A2(npu_inst_pe_1_7_7_n1), .B1(
        npu_inst_pe_1_7_7_N79), .B2(npu_inst_pe_1_7_7_n76), .C1(
        npu_inst_pe_1_7_7_N71), .C2(npu_inst_pe_1_7_7_n77), .ZN(
        npu_inst_pe_1_7_7_n78) );
  INV_X1 npu_inst_pe_1_7_7_U68 ( .A(npu_inst_pe_1_7_7_n78), .ZN(
        npu_inst_pe_1_7_7_n34) );
  AND2_X1 npu_inst_pe_1_7_7_U67 ( .A1(npu_inst_pe_1_7_7_int_q_acc_0_), .A2(
        npu_inst_pe_1_7_7_n1), .ZN(npu_inst_int_data_res_7__7__0_) );
  AND2_X1 npu_inst_pe_1_7_7_U66 ( .A1(npu_inst_pe_1_7_7_n2), .A2(
        npu_inst_pe_1_7_7_int_q_acc_7_), .ZN(npu_inst_int_data_res_7__7__7_)
         );
  AND2_X1 npu_inst_pe_1_7_7_U65 ( .A1(npu_inst_pe_1_7_7_int_q_acc_1_), .A2(
        npu_inst_pe_1_7_7_n1), .ZN(npu_inst_int_data_res_7__7__1_) );
  AND2_X1 npu_inst_pe_1_7_7_U64 ( .A1(npu_inst_pe_1_7_7_int_q_acc_2_), .A2(
        npu_inst_pe_1_7_7_n1), .ZN(npu_inst_int_data_res_7__7__2_) );
  AND2_X1 npu_inst_pe_1_7_7_U63 ( .A1(npu_inst_pe_1_7_7_int_q_acc_3_), .A2(
        npu_inst_pe_1_7_7_n2), .ZN(npu_inst_int_data_res_7__7__3_) );
  AND2_X1 npu_inst_pe_1_7_7_U62 ( .A1(npu_inst_pe_1_7_7_int_q_acc_4_), .A2(
        npu_inst_pe_1_7_7_n2), .ZN(npu_inst_int_data_res_7__7__4_) );
  AND2_X1 npu_inst_pe_1_7_7_U61 ( .A1(npu_inst_pe_1_7_7_int_q_acc_5_), .A2(
        npu_inst_pe_1_7_7_n2), .ZN(npu_inst_int_data_res_7__7__5_) );
  AND2_X1 npu_inst_pe_1_7_7_U60 ( .A1(npu_inst_pe_1_7_7_int_q_acc_6_), .A2(
        npu_inst_pe_1_7_7_n2), .ZN(npu_inst_int_data_res_7__7__6_) );
  INV_X1 npu_inst_pe_1_7_7_U59 ( .A(npu_inst_pe_1_7_7_int_data_1_), .ZN(
        npu_inst_pe_1_7_7_n14) );
  AND2_X1 npu_inst_pe_1_7_7_U58 ( .A1(npu_inst_int_data_x_7__7__1_), .A2(
        npu_inst_pe_1_7_7_int_q_weight_1_), .ZN(npu_inst_pe_1_7_7_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_7_7_U57 ( .A1(npu_inst_int_data_x_7__7__0_), .A2(
        npu_inst_pe_1_7_7_int_q_weight_1_), .ZN(npu_inst_pe_1_7_7_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_7_7_U56 ( .A1(npu_inst_n52), .A2(int_i_data_v_npu[0]), 
        .B1(npu_inst_pe_1_7_7_n3), .B2(int_i_data_h_npu[0]), .ZN(
        npu_inst_pe_1_7_7_n61) );
  NAND2_X1 npu_inst_pe_1_7_7_U55 ( .A1(npu_inst_pe_1_7_7_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_7_7_n60), .ZN(npu_inst_pe_1_7_7_n74) );
  OAI21_X1 npu_inst_pe_1_7_7_U54 ( .B1(npu_inst_pe_1_7_7_n63), .B2(
        npu_inst_pe_1_7_7_n60), .A(npu_inst_pe_1_7_7_n74), .ZN(
        npu_inst_pe_1_7_7_n97) );
  NAND2_X1 npu_inst_pe_1_7_7_U53 ( .A1(npu_inst_pe_1_7_7_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_7_7_n60), .ZN(npu_inst_pe_1_7_7_n73) );
  OAI21_X1 npu_inst_pe_1_7_7_U52 ( .B1(npu_inst_pe_1_7_7_n61), .B2(
        npu_inst_pe_1_7_7_n60), .A(npu_inst_pe_1_7_7_n73), .ZN(
        npu_inst_pe_1_7_7_n96) );
  NAND2_X1 npu_inst_pe_1_7_7_U51 ( .A1(npu_inst_pe_1_7_7_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_7_7_n56), .ZN(npu_inst_pe_1_7_7_n72) );
  OAI21_X1 npu_inst_pe_1_7_7_U50 ( .B1(npu_inst_pe_1_7_7_n63), .B2(
        npu_inst_pe_1_7_7_n56), .A(npu_inst_pe_1_7_7_n72), .ZN(
        npu_inst_pe_1_7_7_n95) );
  NAND2_X1 npu_inst_pe_1_7_7_U49 ( .A1(npu_inst_pe_1_7_7_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_7_7_n56), .ZN(npu_inst_pe_1_7_7_n71) );
  OAI21_X1 npu_inst_pe_1_7_7_U48 ( .B1(npu_inst_pe_1_7_7_n61), .B2(
        npu_inst_pe_1_7_7_n56), .A(npu_inst_pe_1_7_7_n71), .ZN(
        npu_inst_pe_1_7_7_n94) );
  NAND2_X1 npu_inst_pe_1_7_7_U47 ( .A1(npu_inst_pe_1_7_7_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_7_7_n52), .ZN(npu_inst_pe_1_7_7_n70) );
  OAI21_X1 npu_inst_pe_1_7_7_U46 ( .B1(npu_inst_pe_1_7_7_n63), .B2(
        npu_inst_pe_1_7_7_n52), .A(npu_inst_pe_1_7_7_n70), .ZN(
        npu_inst_pe_1_7_7_n93) );
  NAND2_X1 npu_inst_pe_1_7_7_U45 ( .A1(npu_inst_pe_1_7_7_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_7_7_n52), .ZN(npu_inst_pe_1_7_7_n69) );
  OAI21_X1 npu_inst_pe_1_7_7_U44 ( .B1(npu_inst_pe_1_7_7_n61), .B2(
        npu_inst_pe_1_7_7_n52), .A(npu_inst_pe_1_7_7_n69), .ZN(
        npu_inst_pe_1_7_7_n92) );
  NAND2_X1 npu_inst_pe_1_7_7_U43 ( .A1(npu_inst_pe_1_7_7_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_7_7_n48), .ZN(npu_inst_pe_1_7_7_n68) );
  OAI21_X1 npu_inst_pe_1_7_7_U42 ( .B1(npu_inst_pe_1_7_7_n63), .B2(
        npu_inst_pe_1_7_7_n48), .A(npu_inst_pe_1_7_7_n68), .ZN(
        npu_inst_pe_1_7_7_n91) );
  NAND2_X1 npu_inst_pe_1_7_7_U41 ( .A1(npu_inst_pe_1_7_7_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_7_7_n48), .ZN(npu_inst_pe_1_7_7_n67) );
  OAI21_X1 npu_inst_pe_1_7_7_U40 ( .B1(npu_inst_pe_1_7_7_n61), .B2(
        npu_inst_pe_1_7_7_n48), .A(npu_inst_pe_1_7_7_n67), .ZN(
        npu_inst_pe_1_7_7_n90) );
  NAND2_X1 npu_inst_pe_1_7_7_U39 ( .A1(npu_inst_pe_1_7_7_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_7_7_n44), .ZN(npu_inst_pe_1_7_7_n66) );
  OAI21_X1 npu_inst_pe_1_7_7_U38 ( .B1(npu_inst_pe_1_7_7_n63), .B2(
        npu_inst_pe_1_7_7_n44), .A(npu_inst_pe_1_7_7_n66), .ZN(
        npu_inst_pe_1_7_7_n89) );
  NAND2_X1 npu_inst_pe_1_7_7_U37 ( .A1(npu_inst_pe_1_7_7_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_7_7_n44), .ZN(npu_inst_pe_1_7_7_n65) );
  OAI21_X1 npu_inst_pe_1_7_7_U36 ( .B1(npu_inst_pe_1_7_7_n61), .B2(
        npu_inst_pe_1_7_7_n44), .A(npu_inst_pe_1_7_7_n65), .ZN(
        npu_inst_pe_1_7_7_n88) );
  NAND2_X1 npu_inst_pe_1_7_7_U35 ( .A1(npu_inst_pe_1_7_7_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_7_7_n40), .ZN(npu_inst_pe_1_7_7_n64) );
  OAI21_X1 npu_inst_pe_1_7_7_U34 ( .B1(npu_inst_pe_1_7_7_n63), .B2(
        npu_inst_pe_1_7_7_n40), .A(npu_inst_pe_1_7_7_n64), .ZN(
        npu_inst_pe_1_7_7_n87) );
  NAND2_X1 npu_inst_pe_1_7_7_U33 ( .A1(npu_inst_pe_1_7_7_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_7_7_n40), .ZN(npu_inst_pe_1_7_7_n62) );
  OAI21_X1 npu_inst_pe_1_7_7_U32 ( .B1(npu_inst_pe_1_7_7_n61), .B2(
        npu_inst_pe_1_7_7_n40), .A(npu_inst_pe_1_7_7_n62), .ZN(
        npu_inst_pe_1_7_7_n86) );
  AOI22_X1 npu_inst_pe_1_7_7_U31 ( .A1(npu_inst_n52), .A2(int_i_data_v_npu[1]), 
        .B1(npu_inst_pe_1_7_7_n3), .B2(int_i_data_h_npu[1]), .ZN(
        npu_inst_pe_1_7_7_n63) );
  INV_X1 npu_inst_pe_1_7_7_U30 ( .A(npu_inst_pe_1_7_7_int_data_0_), .ZN(
        npu_inst_pe_1_7_7_n13) );
  INV_X1 npu_inst_pe_1_7_7_U29 ( .A(npu_inst_n67), .ZN(npu_inst_pe_1_7_7_n5)
         );
  OR3_X1 npu_inst_pe_1_7_7_U28 ( .A1(npu_inst_pe_1_7_7_n6), .A2(
        npu_inst_pe_1_7_7_n8), .A3(npu_inst_pe_1_7_7_n5), .ZN(
        npu_inst_pe_1_7_7_n56) );
  OR3_X1 npu_inst_pe_1_7_7_U27 ( .A1(npu_inst_pe_1_7_7_n5), .A2(
        npu_inst_pe_1_7_7_n8), .A3(npu_inst_pe_1_7_7_n7), .ZN(
        npu_inst_pe_1_7_7_n48) );
  INV_X1 npu_inst_pe_1_7_7_U26 ( .A(npu_inst_pe_1_7_7_n5), .ZN(
        npu_inst_pe_1_7_7_n4) );
  OR3_X1 npu_inst_pe_1_7_7_U25 ( .A1(npu_inst_pe_1_7_7_n4), .A2(
        npu_inst_pe_1_7_7_n8), .A3(npu_inst_pe_1_7_7_n7), .ZN(
        npu_inst_pe_1_7_7_n52) );
  OR3_X1 npu_inst_pe_1_7_7_U24 ( .A1(npu_inst_pe_1_7_7_n6), .A2(
        npu_inst_pe_1_7_7_n8), .A3(npu_inst_pe_1_7_7_n4), .ZN(
        npu_inst_pe_1_7_7_n60) );
  NOR2_X1 npu_inst_pe_1_7_7_U23 ( .A1(npu_inst_pe_1_7_7_n60), .A2(
        npu_inst_pe_1_7_7_n3), .ZN(npu_inst_pe_1_7_7_n58) );
  NOR2_X1 npu_inst_pe_1_7_7_U22 ( .A1(npu_inst_pe_1_7_7_n56), .A2(
        npu_inst_pe_1_7_7_n3), .ZN(npu_inst_pe_1_7_7_n54) );
  NOR2_X1 npu_inst_pe_1_7_7_U21 ( .A1(npu_inst_pe_1_7_7_n52), .A2(
        npu_inst_pe_1_7_7_n3), .ZN(npu_inst_pe_1_7_7_n50) );
  NOR2_X1 npu_inst_pe_1_7_7_U20 ( .A1(npu_inst_pe_1_7_7_n48), .A2(
        npu_inst_pe_1_7_7_n3), .ZN(npu_inst_pe_1_7_7_n46) );
  NOR2_X1 npu_inst_pe_1_7_7_U19 ( .A1(npu_inst_pe_1_7_7_n40), .A2(
        npu_inst_pe_1_7_7_n3), .ZN(npu_inst_pe_1_7_7_n38) );
  NOR2_X1 npu_inst_pe_1_7_7_U18 ( .A1(npu_inst_pe_1_7_7_n44), .A2(
        npu_inst_pe_1_7_7_n3), .ZN(npu_inst_pe_1_7_7_n42) );
  BUF_X1 npu_inst_pe_1_7_7_U17 ( .A(npu_inst_n92), .Z(npu_inst_pe_1_7_7_n8) );
  INV_X1 npu_inst_pe_1_7_7_U16 ( .A(npu_inst_n122), .ZN(npu_inst_pe_1_7_7_n12)
         );
  INV_X1 npu_inst_pe_1_7_7_U15 ( .A(npu_inst_pe_1_7_7_n38), .ZN(
        npu_inst_pe_1_7_7_n114) );
  INV_X1 npu_inst_pe_1_7_7_U14 ( .A(npu_inst_pe_1_7_7_n58), .ZN(
        npu_inst_pe_1_7_7_n119) );
  INV_X1 npu_inst_pe_1_7_7_U13 ( .A(npu_inst_pe_1_7_7_n54), .ZN(
        npu_inst_pe_1_7_7_n118) );
  INV_X1 npu_inst_pe_1_7_7_U12 ( .A(npu_inst_pe_1_7_7_n50), .ZN(
        npu_inst_pe_1_7_7_n117) );
  INV_X1 npu_inst_pe_1_7_7_U11 ( .A(npu_inst_pe_1_7_7_n46), .ZN(
        npu_inst_pe_1_7_7_n116) );
  INV_X1 npu_inst_pe_1_7_7_U10 ( .A(npu_inst_pe_1_7_7_n42), .ZN(
        npu_inst_pe_1_7_7_n115) );
  BUF_X1 npu_inst_pe_1_7_7_U9 ( .A(npu_inst_n7), .Z(npu_inst_pe_1_7_7_n2) );
  BUF_X1 npu_inst_pe_1_7_7_U8 ( .A(npu_inst_n7), .Z(npu_inst_pe_1_7_7_n1) );
  BUF_X1 npu_inst_pe_1_7_7_U7 ( .A(npu_inst_pe_1_7_7_n12), .Z(
        npu_inst_pe_1_7_7_n11) );
  BUF_X1 npu_inst_pe_1_7_7_U6 ( .A(npu_inst_pe_1_7_7_n12), .Z(
        npu_inst_pe_1_7_7_n10) );
  BUF_X1 npu_inst_pe_1_7_7_U5 ( .A(npu_inst_pe_1_7_7_n12), .Z(
        npu_inst_pe_1_7_7_n9) );
  NOR2_X1 npu_inst_pe_1_7_7_U4 ( .A1(npu_inst_pe_1_7_7_int_q_weight_0_), .A2(
        npu_inst_pe_1_7_7_n1), .ZN(npu_inst_pe_1_7_7_n76) );
  NOR2_X1 npu_inst_pe_1_7_7_U3 ( .A1(npu_inst_pe_1_7_7_n27), .A2(
        npu_inst_pe_1_7_7_n1), .ZN(npu_inst_pe_1_7_7_n77) );
  FA_X1 npu_inst_pe_1_7_7_sub_67_U2_1 ( .A(npu_inst_pe_1_7_7_int_q_acc_1_), 
        .B(npu_inst_pe_1_7_7_n14), .CI(npu_inst_pe_1_7_7_sub_67_carry_1_), 
        .CO(npu_inst_pe_1_7_7_sub_67_carry_2_), .S(npu_inst_pe_1_7_7_N66) );
  FA_X1 npu_inst_pe_1_7_7_add_69_U1_1 ( .A(npu_inst_pe_1_7_7_int_q_acc_1_), 
        .B(npu_inst_pe_1_7_7_int_data_1_), .CI(
        npu_inst_pe_1_7_7_add_69_carry_1_), .CO(
        npu_inst_pe_1_7_7_add_69_carry_2_), .S(npu_inst_pe_1_7_7_N74) );
  NAND3_X1 npu_inst_pe_1_7_7_U109 ( .A1(npu_inst_pe_1_7_7_n5), .A2(
        npu_inst_pe_1_7_7_n7), .A3(npu_inst_pe_1_7_7_n8), .ZN(
        npu_inst_pe_1_7_7_n44) );
  NAND3_X1 npu_inst_pe_1_7_7_U108 ( .A1(npu_inst_pe_1_7_7_n4), .A2(
        npu_inst_pe_1_7_7_n7), .A3(npu_inst_pe_1_7_7_n8), .ZN(
        npu_inst_pe_1_7_7_n40) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_7_7_n34), .CK(
        npu_inst_pe_1_7_7_net3113), .RN(npu_inst_pe_1_7_7_n9), .Q(
        npu_inst_pe_1_7_7_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_7_7_n35), .CK(
        npu_inst_pe_1_7_7_net3113), .RN(npu_inst_pe_1_7_7_n9), .Q(
        npu_inst_pe_1_7_7_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_7_7_n36), .CK(
        npu_inst_pe_1_7_7_net3113), .RN(npu_inst_pe_1_7_7_n9), .Q(
        npu_inst_pe_1_7_7_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_7_7_n98), .CK(
        npu_inst_pe_1_7_7_net3113), .RN(npu_inst_pe_1_7_7_n9), .Q(
        npu_inst_pe_1_7_7_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_7_7_n99), .CK(
        npu_inst_pe_1_7_7_net3113), .RN(npu_inst_pe_1_7_7_n9), .Q(
        npu_inst_pe_1_7_7_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_7_7_n100), 
        .CK(npu_inst_pe_1_7_7_net3113), .RN(npu_inst_pe_1_7_7_n9), .Q(
        npu_inst_pe_1_7_7_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_7_7_n33), .CK(
        npu_inst_pe_1_7_7_net3113), .RN(npu_inst_pe_1_7_7_n9), .Q(
        npu_inst_pe_1_7_7_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_7_7_n101), 
        .CK(npu_inst_pe_1_7_7_net3113), .RN(npu_inst_pe_1_7_7_n9), .Q(
        npu_inst_pe_1_7_7_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_weight_reg_0_ ( .D(npu_inst_n108), .CK(
        npu_inst_pe_1_7_7_net3119), .RN(npu_inst_pe_1_7_7_n9), .Q(
        npu_inst_pe_1_7_7_int_q_weight_0_), .QN(npu_inst_pe_1_7_7_n27) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_weight_reg_1_ ( .D(npu_inst_n114), .CK(
        npu_inst_pe_1_7_7_net3119), .RN(npu_inst_pe_1_7_7_n9), .Q(
        npu_inst_pe_1_7_7_int_q_weight_1_), .QN(npu_inst_pe_1_7_7_n26) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_7_7_n113), 
        .CK(npu_inst_pe_1_7_7_net3119), .RN(npu_inst_pe_1_7_7_n9), .Q(
        npu_inst_pe_1_7_7_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_7_7_n112), 
        .CK(npu_inst_pe_1_7_7_net3119), .RN(npu_inst_pe_1_7_7_n9), .Q(
        npu_inst_pe_1_7_7_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_7_7_n111), 
        .CK(npu_inst_pe_1_7_7_net3119), .RN(npu_inst_pe_1_7_7_n10), .Q(
        npu_inst_pe_1_7_7_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_7_7_n110), 
        .CK(npu_inst_pe_1_7_7_net3119), .RN(npu_inst_pe_1_7_7_n10), .Q(
        npu_inst_pe_1_7_7_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_7_7_n109), 
        .CK(npu_inst_pe_1_7_7_net3119), .RN(npu_inst_pe_1_7_7_n10), .Q(
        npu_inst_pe_1_7_7_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_7_7_n108), 
        .CK(npu_inst_pe_1_7_7_net3119), .RN(npu_inst_pe_1_7_7_n10), .Q(
        npu_inst_pe_1_7_7_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_7_7_n107), 
        .CK(npu_inst_pe_1_7_7_net3119), .RN(npu_inst_pe_1_7_7_n10), .Q(
        npu_inst_pe_1_7_7_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_7_7_n106), 
        .CK(npu_inst_pe_1_7_7_net3119), .RN(npu_inst_pe_1_7_7_n10), .Q(
        npu_inst_pe_1_7_7_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_7_7_n105), 
        .CK(npu_inst_pe_1_7_7_net3119), .RN(npu_inst_pe_1_7_7_n10), .Q(
        npu_inst_pe_1_7_7_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_7_7_n104), 
        .CK(npu_inst_pe_1_7_7_net3119), .RN(npu_inst_pe_1_7_7_n10), .Q(
        npu_inst_pe_1_7_7_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_7_7_n103), 
        .CK(npu_inst_pe_1_7_7_net3119), .RN(npu_inst_pe_1_7_7_n10), .Q(
        npu_inst_pe_1_7_7_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_7_7_n102), 
        .CK(npu_inst_pe_1_7_7_net3119), .RN(npu_inst_pe_1_7_7_n10), .Q(
        npu_inst_pe_1_7_7_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_7_7_n86), 
        .CK(npu_inst_pe_1_7_7_net3119), .RN(npu_inst_pe_1_7_7_n10), .Q(
        npu_inst_pe_1_7_7_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_7_7_n87), 
        .CK(npu_inst_pe_1_7_7_net3119), .RN(npu_inst_pe_1_7_7_n10), .Q(
        npu_inst_pe_1_7_7_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_7_7_n88), 
        .CK(npu_inst_pe_1_7_7_net3119), .RN(npu_inst_pe_1_7_7_n11), .Q(
        npu_inst_pe_1_7_7_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_7_7_n89), 
        .CK(npu_inst_pe_1_7_7_net3119), .RN(npu_inst_pe_1_7_7_n11), .Q(
        npu_inst_pe_1_7_7_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_7_7_n90), 
        .CK(npu_inst_pe_1_7_7_net3119), .RN(npu_inst_pe_1_7_7_n11), .Q(
        npu_inst_pe_1_7_7_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_7_7_n91), 
        .CK(npu_inst_pe_1_7_7_net3119), .RN(npu_inst_pe_1_7_7_n11), .Q(
        npu_inst_pe_1_7_7_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_7_7_n92), 
        .CK(npu_inst_pe_1_7_7_net3119), .RN(npu_inst_pe_1_7_7_n11), .Q(
        npu_inst_pe_1_7_7_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_7_7_n93), 
        .CK(npu_inst_pe_1_7_7_net3119), .RN(npu_inst_pe_1_7_7_n11), .Q(
        npu_inst_pe_1_7_7_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_7_7_n94), 
        .CK(npu_inst_pe_1_7_7_net3119), .RN(npu_inst_pe_1_7_7_n11), .Q(
        npu_inst_pe_1_7_7_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_7_7_n95), 
        .CK(npu_inst_pe_1_7_7_net3119), .RN(npu_inst_pe_1_7_7_n11), .Q(
        npu_inst_pe_1_7_7_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_7_7_n96), 
        .CK(npu_inst_pe_1_7_7_net3119), .RN(npu_inst_pe_1_7_7_n11), .Q(
        npu_inst_pe_1_7_7_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_7_7_n97), 
        .CK(npu_inst_pe_1_7_7_net3119), .RN(npu_inst_pe_1_7_7_n11), .Q(
        npu_inst_pe_1_7_7_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_7_7_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_7_7_N84), .SE(1'b0), .GCK(npu_inst_pe_1_7_7_net3113) );
  CLKGATETST_X1 npu_inst_pe_1_7_7_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n61), .SE(1'b0), .GCK(npu_inst_pe_1_7_7_net3119) );
  INV_X1 qrelu_i_0_U8 ( .A(int_o_data_npu[57]), .ZN(qrelu_i_0_n3) );
  OAI21_X1 qrelu_i_0_U7 ( .B1(qrelu_i_0_n3), .B2(int_o_data_npu[63]), .A(
        qrelu_i_0_n4), .ZN(o_data_relu[15]) );
  INV_X1 qrelu_i_0_U6 ( .A(int_o_data_npu[56]), .ZN(qrelu_i_0_n1) );
  OAI21_X1 qrelu_i_0_U5 ( .B1(qrelu_i_0_n1), .B2(int_o_data_npu[63]), .A(
        qrelu_i_0_n4), .ZN(o_data_relu[14]) );
  OR3_X1 qrelu_i_0_U4 ( .A1(int_o_data_npu[62]), .A2(int_o_data_npu[61]), .A3(
        int_o_data_npu[60]), .ZN(qrelu_i_0_n5) );
  OR2_X1 qrelu_i_0_U3 ( .A1(int_o_data_npu[59]), .A2(int_o_data_npu[58]), .ZN(
        qrelu_i_0_n6) );
  INV_X1 qrelu_i_0_U2 ( .A(int_o_data_npu[63]), .ZN(qrelu_i_0_n2) );
  OAI21_X1 qrelu_i_0_U1 ( .B1(qrelu_i_0_n5), .B2(qrelu_i_0_n6), .A(
        qrelu_i_0_n2), .ZN(qrelu_i_0_n4) );
  INV_X1 qrelu_i_1_U8 ( .A(int_o_data_npu[49]), .ZN(qrelu_i_1_n3) );
  OAI21_X1 qrelu_i_1_U7 ( .B1(qrelu_i_1_n3), .B2(int_o_data_npu[55]), .A(
        qrelu_i_1_n9), .ZN(o_data_relu[13]) );
  INV_X1 qrelu_i_1_U6 ( .A(int_o_data_npu[48]), .ZN(qrelu_i_1_n1) );
  OAI21_X1 qrelu_i_1_U5 ( .B1(qrelu_i_1_n1), .B2(int_o_data_npu[55]), .A(
        qrelu_i_1_n9), .ZN(o_data_relu[12]) );
  OR3_X1 qrelu_i_1_U4 ( .A1(int_o_data_npu[54]), .A2(int_o_data_npu[53]), .A3(
        int_o_data_npu[52]), .ZN(qrelu_i_1_n8) );
  OR2_X1 qrelu_i_1_U3 ( .A1(int_o_data_npu[51]), .A2(int_o_data_npu[50]), .ZN(
        qrelu_i_1_n7) );
  INV_X1 qrelu_i_1_U2 ( .A(int_o_data_npu[55]), .ZN(qrelu_i_1_n2) );
  OAI21_X1 qrelu_i_1_U1 ( .B1(qrelu_i_1_n8), .B2(qrelu_i_1_n7), .A(
        qrelu_i_1_n2), .ZN(qrelu_i_1_n9) );
  INV_X1 qrelu_i_2_U8 ( .A(int_o_data_npu[41]), .ZN(qrelu_i_2_n3) );
  OAI21_X1 qrelu_i_2_U7 ( .B1(qrelu_i_2_n3), .B2(int_o_data_npu[47]), .A(
        qrelu_i_2_n9), .ZN(o_data_relu[11]) );
  INV_X1 qrelu_i_2_U6 ( .A(int_o_data_npu[40]), .ZN(qrelu_i_2_n1) );
  OAI21_X1 qrelu_i_2_U5 ( .B1(qrelu_i_2_n1), .B2(int_o_data_npu[47]), .A(
        qrelu_i_2_n9), .ZN(o_data_relu[10]) );
  OR3_X1 qrelu_i_2_U4 ( .A1(int_o_data_npu[46]), .A2(int_o_data_npu[45]), .A3(
        int_o_data_npu[44]), .ZN(qrelu_i_2_n8) );
  OR2_X1 qrelu_i_2_U3 ( .A1(int_o_data_npu[43]), .A2(int_o_data_npu[42]), .ZN(
        qrelu_i_2_n7) );
  INV_X1 qrelu_i_2_U2 ( .A(int_o_data_npu[47]), .ZN(qrelu_i_2_n2) );
  OAI21_X1 qrelu_i_2_U1 ( .B1(qrelu_i_2_n8), .B2(qrelu_i_2_n7), .A(
        qrelu_i_2_n2), .ZN(qrelu_i_2_n9) );
  INV_X1 qrelu_i_3_U8 ( .A(int_o_data_npu[33]), .ZN(qrelu_i_3_n3) );
  OAI21_X1 qrelu_i_3_U7 ( .B1(qrelu_i_3_n3), .B2(int_o_data_npu[39]), .A(
        qrelu_i_3_n9), .ZN(o_data_relu[9]) );
  INV_X1 qrelu_i_3_U6 ( .A(int_o_data_npu[32]), .ZN(qrelu_i_3_n1) );
  OAI21_X1 qrelu_i_3_U5 ( .B1(qrelu_i_3_n1), .B2(int_o_data_npu[39]), .A(
        qrelu_i_3_n9), .ZN(o_data_relu[8]) );
  OR3_X1 qrelu_i_3_U4 ( .A1(int_o_data_npu[38]), .A2(int_o_data_npu[37]), .A3(
        int_o_data_npu[36]), .ZN(qrelu_i_3_n8) );
  OR2_X1 qrelu_i_3_U3 ( .A1(int_o_data_npu[35]), .A2(int_o_data_npu[34]), .ZN(
        qrelu_i_3_n7) );
  INV_X1 qrelu_i_3_U2 ( .A(int_o_data_npu[39]), .ZN(qrelu_i_3_n2) );
  OAI21_X1 qrelu_i_3_U1 ( .B1(qrelu_i_3_n8), .B2(qrelu_i_3_n7), .A(
        qrelu_i_3_n2), .ZN(qrelu_i_3_n9) );
  INV_X1 qrelu_i_4_U8 ( .A(int_o_data_npu[25]), .ZN(qrelu_i_4_n3) );
  OAI21_X1 qrelu_i_4_U7 ( .B1(qrelu_i_4_n3), .B2(int_o_data_npu[31]), .A(
        qrelu_i_4_n9), .ZN(o_data_relu[7]) );
  INV_X1 qrelu_i_4_U6 ( .A(int_o_data_npu[24]), .ZN(qrelu_i_4_n1) );
  OAI21_X1 qrelu_i_4_U5 ( .B1(qrelu_i_4_n1), .B2(int_o_data_npu[31]), .A(
        qrelu_i_4_n9), .ZN(o_data_relu[6]) );
  OR3_X1 qrelu_i_4_U4 ( .A1(int_o_data_npu[30]), .A2(int_o_data_npu[29]), .A3(
        int_o_data_npu[28]), .ZN(qrelu_i_4_n8) );
  OR2_X1 qrelu_i_4_U3 ( .A1(int_o_data_npu[27]), .A2(int_o_data_npu[26]), .ZN(
        qrelu_i_4_n7) );
  INV_X1 qrelu_i_4_U2 ( .A(int_o_data_npu[31]), .ZN(qrelu_i_4_n2) );
  OAI21_X1 qrelu_i_4_U1 ( .B1(qrelu_i_4_n8), .B2(qrelu_i_4_n7), .A(
        qrelu_i_4_n2), .ZN(qrelu_i_4_n9) );
  INV_X1 qrelu_i_5_U8 ( .A(int_o_data_npu[17]), .ZN(qrelu_i_5_n3) );
  OAI21_X1 qrelu_i_5_U7 ( .B1(qrelu_i_5_n3), .B2(int_o_data_npu[23]), .A(
        qrelu_i_5_n9), .ZN(o_data_relu[5]) );
  INV_X1 qrelu_i_5_U6 ( .A(int_o_data_npu[16]), .ZN(qrelu_i_5_n1) );
  OAI21_X1 qrelu_i_5_U5 ( .B1(qrelu_i_5_n1), .B2(int_o_data_npu[23]), .A(
        qrelu_i_5_n9), .ZN(o_data_relu[4]) );
  OR3_X1 qrelu_i_5_U4 ( .A1(int_o_data_npu[22]), .A2(int_o_data_npu[21]), .A3(
        int_o_data_npu[20]), .ZN(qrelu_i_5_n8) );
  OR2_X1 qrelu_i_5_U3 ( .A1(int_o_data_npu[19]), .A2(int_o_data_npu[18]), .ZN(
        qrelu_i_5_n7) );
  INV_X1 qrelu_i_5_U2 ( .A(int_o_data_npu[23]), .ZN(qrelu_i_5_n2) );
  OAI21_X1 qrelu_i_5_U1 ( .B1(qrelu_i_5_n8), .B2(qrelu_i_5_n7), .A(
        qrelu_i_5_n2), .ZN(qrelu_i_5_n9) );
  INV_X1 qrelu_i_6_U8 ( .A(int_o_data_npu[9]), .ZN(qrelu_i_6_n3) );
  OAI21_X1 qrelu_i_6_U7 ( .B1(qrelu_i_6_n3), .B2(int_o_data_npu[15]), .A(
        qrelu_i_6_n9), .ZN(o_data_relu[3]) );
  INV_X1 qrelu_i_6_U6 ( .A(int_o_data_npu[8]), .ZN(qrelu_i_6_n1) );
  OAI21_X1 qrelu_i_6_U5 ( .B1(qrelu_i_6_n1), .B2(int_o_data_npu[15]), .A(
        qrelu_i_6_n9), .ZN(o_data_relu[2]) );
  OR3_X1 qrelu_i_6_U4 ( .A1(int_o_data_npu[14]), .A2(int_o_data_npu[13]), .A3(
        int_o_data_npu[12]), .ZN(qrelu_i_6_n8) );
  OR2_X1 qrelu_i_6_U3 ( .A1(int_o_data_npu[11]), .A2(int_o_data_npu[10]), .ZN(
        qrelu_i_6_n7) );
  INV_X1 qrelu_i_6_U2 ( .A(int_o_data_npu[15]), .ZN(qrelu_i_6_n2) );
  OAI21_X1 qrelu_i_6_U1 ( .B1(qrelu_i_6_n8), .B2(qrelu_i_6_n7), .A(
        qrelu_i_6_n2), .ZN(qrelu_i_6_n9) );
  INV_X1 qrelu_i_7_U8 ( .A(int_o_data_npu[1]), .ZN(qrelu_i_7_n3) );
  OAI21_X1 qrelu_i_7_U7 ( .B1(qrelu_i_7_n3), .B2(int_o_data_npu[7]), .A(
        qrelu_i_7_n9), .ZN(o_data_relu[1]) );
  INV_X1 qrelu_i_7_U6 ( .A(int_o_data_npu[0]), .ZN(qrelu_i_7_n1) );
  OAI21_X1 qrelu_i_7_U5 ( .B1(qrelu_i_7_n1), .B2(int_o_data_npu[7]), .A(
        qrelu_i_7_n9), .ZN(o_data_relu[0]) );
  OR3_X1 qrelu_i_7_U4 ( .A1(int_o_data_npu[6]), .A2(int_o_data_npu[5]), .A3(
        int_o_data_npu[4]), .ZN(qrelu_i_7_n8) );
  OR2_X1 qrelu_i_7_U3 ( .A1(int_o_data_npu[3]), .A2(int_o_data_npu[2]), .ZN(
        qrelu_i_7_n7) );
  INV_X1 qrelu_i_7_U2 ( .A(int_o_data_npu[7]), .ZN(qrelu_i_7_n2) );
  OAI21_X1 qrelu_i_7_U1 ( .B1(qrelu_i_7_n8), .B2(qrelu_i_7_n7), .A(
        qrelu_i_7_n2), .ZN(qrelu_i_7_n9) );
  INV_X1 p_unit_i_0_U18 ( .A(rst), .ZN(p_unit_i_0_n11) );
  INV_X1 p_unit_i_0_U17 ( .A(p_unit_i_0_n8), .ZN(p_unit_i_0_n16) );
  NOR2_X1 p_unit_i_0_U15 ( .A1(p_unit_i_0_int_ps0_2_), .A2(p_unit_i_0_n16), 
        .ZN(p_unit_i_0_n6) );
  OAI22_X1 p_unit_i_0_U14 ( .A1(p_unit_i_0_n8), .A2(p_unit_i_0_n5), .B1(
        p_unit_i_0_n6), .B2(p_unit_i_0_n7), .ZN(p_unit_i_0_n4) );
  OAI211_X1 p_unit_i_0_U13 ( .C1(p_unit_i_0_int_ps0_1_), .C2(
        p_unit_i_0_int_ps1_1_), .A(p_unit_i_0_int_ps0_0_), .B(
        p_unit_i_0_int_ps1_0_), .ZN(p_unit_i_0_n10) );
  INV_X1 p_unit_i_0_U12 ( .A(p_unit_i_0_n10), .ZN(p_unit_i_0_n17) );
  AOI21_X1 p_unit_i_0_U11 ( .B1(p_unit_i_0_int_ps0_1_), .B2(
        p_unit_i_0_int_ps1_1_), .A(p_unit_i_0_n17), .ZN(p_unit_i_0_n8) );
  XNOR2_X1 p_unit_i_0_U10 ( .A(p_unit_i_0_n8), .B(p_unit_i_0_n9), .ZN(
        p_unit_i_0_N7) );
  XNOR2_X1 p_unit_i_0_U9 ( .A(p_unit_i_0_int_ps1_1_), .B(p_unit_i_0_int_ps0_1_), .ZN(p_unit_i_0_n3) );
  NAND2_X1 p_unit_i_0_U8 ( .A1(p_unit_i_0_int_ps0_0_), .A2(
        p_unit_i_0_int_ps1_0_), .ZN(p_unit_i_0_n2) );
  XOR2_X1 p_unit_i_0_U7 ( .A(p_unit_i_0_n2), .B(p_unit_i_0_n3), .Z(
        p_unit_i_0_N6) );
  AND3_X1 p_unit_i_0_U6 ( .A1(o_data_relu[14]), .A2(p_unit_i_0_n15), .A3(
        o_data_relu[12]), .ZN(p_unit_i_0_n14) );
  AOI21_X1 p_unit_i_0_U5 ( .B1(o_data_relu[13]), .B2(o_data_relu[15]), .A(
        p_unit_i_0_n14), .ZN(p_unit_i_0_n13) );
  INV_X1 p_unit_i_0_U4 ( .A(p_unit_i_0_n13), .ZN(p_unit_i_0_n12) );
  NAND2_X1 p_unit_i_0_U3 ( .A1(o_data_relu[14]), .A2(o_data_relu[12]), .ZN(
        p_unit_i_0_n1) );
  XNOR2_X1 p_unit_i_0_U2 ( .A(p_unit_i_0_n1), .B(p_unit_i_0_n15), .ZN(
        p_unit_i_0_N3) );
  DFFR_X1 p_unit_i_0_o_data_reg_3_ ( .D(p_unit_i_0_n4), .CK(p_unit_i_0_net3095), .RN(p_unit_i_0_n11), .Q(int_o_data_p[15]) );
  DFFR_X1 p_unit_i_0_o_data_reg_2_ ( .D(p_unit_i_0_N7), .CK(p_unit_i_0_net3095), .RN(p_unit_i_0_n11), .Q(int_o_data_p[14]) );
  DFFR_X1 p_unit_i_0_o_data_reg_1_ ( .D(p_unit_i_0_N6), .CK(p_unit_i_0_net3095), .RN(p_unit_i_0_n11), .Q(int_o_data_p[13]) );
  DFFR_X1 p_unit_i_0_o_data_reg_0_ ( .D(p_unit_i_0_N5), .CK(p_unit_i_0_net3095), .RN(p_unit_i_0_n11), .Q(int_o_data_p[12]) );
  DFFR_X1 p_unit_i_0_int_ps1_reg_1_ ( .D(p_unit_i_0_int_ps0_1_), .CK(
        p_unit_i_0_net3095), .RN(p_unit_i_0_n11), .Q(p_unit_i_0_int_ps1_1_) );
  DFFR_X1 p_unit_i_0_int_ps1_reg_0_ ( .D(p_unit_i_0_int_ps0_0_), .CK(
        p_unit_i_0_net3095), .RN(p_unit_i_0_n11), .Q(p_unit_i_0_int_ps1_0_) );
  XOR2_X1 p_unit_i_0_U22 ( .A(o_data_relu[12]), .B(o_data_relu[14]), .Z(
        p_unit_i_0_N2) );
  XOR2_X1 p_unit_i_0_U21 ( .A(o_data_relu[15]), .B(o_data_relu[13]), .Z(
        p_unit_i_0_n15) );
  XOR2_X1 p_unit_i_0_U19 ( .A(p_unit_i_0_int_ps1_0_), .B(p_unit_i_0_int_ps0_0_), .Z(p_unit_i_0_N5) );
  XOR2_X1 p_unit_i_0_U16 ( .A(p_unit_i_0_int_ps1_2_), .B(p_unit_i_0_int_ps0_2_), .Z(p_unit_i_0_n9) );
  DFFR_X1 p_unit_i_0_int_ps1_reg_2_ ( .D(p_unit_i_0_int_ps0_2_), .CK(
        p_unit_i_0_net3095), .RN(p_unit_i_0_n11), .Q(p_unit_i_0_int_ps1_2_), 
        .QN(p_unit_i_0_n7) );
  DFFR_X1 p_unit_i_0_int_ps0_reg_0_ ( .D(p_unit_i_0_N2), .CK(
        p_unit_i_0_net3095), .RN(p_unit_i_0_n11), .Q(p_unit_i_0_int_ps0_0_) );
  DFFR_X1 p_unit_i_0_int_ps0_reg_1_ ( .D(p_unit_i_0_N3), .CK(
        p_unit_i_0_net3095), .RN(p_unit_i_0_n11), .Q(p_unit_i_0_int_ps0_1_) );
  DFFR_X1 p_unit_i_0_int_ps0_reg_2_ ( .D(p_unit_i_0_n12), .CK(
        p_unit_i_0_net3095), .RN(p_unit_i_0_n11), .Q(p_unit_i_0_int_ps0_2_), 
        .QN(p_unit_i_0_n5) );
  CLKGATETST_X1 p_unit_i_0_clk_gate_o_data_reg_latch ( .CK(ck), .E(
        ps_ctrl_en_p), .SE(1'b0), .GCK(p_unit_i_0_net3095) );
  INV_X1 p_unit_i_1_U18 ( .A(rst), .ZN(p_unit_i_1_n11) );
  INV_X1 p_unit_i_1_U17 ( .A(p_unit_i_1_n8), .ZN(p_unit_i_1_n16) );
  NOR2_X1 p_unit_i_1_U15 ( .A1(p_unit_i_1_int_ps0_2_), .A2(p_unit_i_1_n16), 
        .ZN(p_unit_i_1_n6) );
  OAI22_X1 p_unit_i_1_U14 ( .A1(p_unit_i_1_n8), .A2(p_unit_i_1_n5), .B1(
        p_unit_i_1_n6), .B2(p_unit_i_1_n7), .ZN(p_unit_i_1_n4) );
  OAI211_X1 p_unit_i_1_U13 ( .C1(p_unit_i_1_int_ps0_1_), .C2(
        p_unit_i_1_int_ps1_1_), .A(p_unit_i_1_int_ps0_0_), .B(
        p_unit_i_1_int_ps1_0_), .ZN(p_unit_i_1_n10) );
  INV_X1 p_unit_i_1_U12 ( .A(p_unit_i_1_n10), .ZN(p_unit_i_1_n17) );
  AOI21_X1 p_unit_i_1_U11 ( .B1(p_unit_i_1_int_ps0_1_), .B2(
        p_unit_i_1_int_ps1_1_), .A(p_unit_i_1_n17), .ZN(p_unit_i_1_n8) );
  XNOR2_X1 p_unit_i_1_U10 ( .A(p_unit_i_1_n8), .B(p_unit_i_1_n9), .ZN(
        p_unit_i_1_N7) );
  XNOR2_X1 p_unit_i_1_U9 ( .A(p_unit_i_1_int_ps1_1_), .B(p_unit_i_1_int_ps0_1_), .ZN(p_unit_i_1_n3) );
  NAND2_X1 p_unit_i_1_U8 ( .A1(p_unit_i_1_int_ps0_0_), .A2(
        p_unit_i_1_int_ps1_0_), .ZN(p_unit_i_1_n2) );
  XOR2_X1 p_unit_i_1_U7 ( .A(p_unit_i_1_n2), .B(p_unit_i_1_n3), .Z(
        p_unit_i_1_N6) );
  AND3_X1 p_unit_i_1_U6 ( .A1(o_data_relu[10]), .A2(p_unit_i_1_n15), .A3(
        o_data_relu[8]), .ZN(p_unit_i_1_n14) );
  AOI21_X1 p_unit_i_1_U5 ( .B1(o_data_relu[9]), .B2(o_data_relu[11]), .A(
        p_unit_i_1_n14), .ZN(p_unit_i_1_n13) );
  INV_X1 p_unit_i_1_U4 ( .A(p_unit_i_1_n13), .ZN(p_unit_i_1_n12) );
  NAND2_X1 p_unit_i_1_U3 ( .A1(o_data_relu[10]), .A2(o_data_relu[8]), .ZN(
        p_unit_i_1_n1) );
  XNOR2_X1 p_unit_i_1_U2 ( .A(p_unit_i_1_n1), .B(p_unit_i_1_n15), .ZN(
        p_unit_i_1_N3) );
  DFFR_X1 p_unit_i_1_o_data_reg_3_ ( .D(p_unit_i_1_n4), .CK(p_unit_i_1_net3077), .RN(p_unit_i_1_n11), .Q(int_o_data_p[11]) );
  DFFR_X1 p_unit_i_1_o_data_reg_2_ ( .D(p_unit_i_1_N7), .CK(p_unit_i_1_net3077), .RN(p_unit_i_1_n11), .Q(int_o_data_p[10]) );
  DFFR_X1 p_unit_i_1_o_data_reg_1_ ( .D(p_unit_i_1_N6), .CK(p_unit_i_1_net3077), .RN(p_unit_i_1_n11), .Q(int_o_data_p[9]) );
  DFFR_X1 p_unit_i_1_o_data_reg_0_ ( .D(p_unit_i_1_N5), .CK(p_unit_i_1_net3077), .RN(p_unit_i_1_n11), .Q(int_o_data_p[8]) );
  DFFR_X1 p_unit_i_1_int_ps1_reg_1_ ( .D(p_unit_i_1_int_ps0_1_), .CK(
        p_unit_i_1_net3077), .RN(p_unit_i_1_n11), .Q(p_unit_i_1_int_ps1_1_) );
  DFFR_X1 p_unit_i_1_int_ps1_reg_0_ ( .D(p_unit_i_1_int_ps0_0_), .CK(
        p_unit_i_1_net3077), .RN(p_unit_i_1_n11), .Q(p_unit_i_1_int_ps1_0_) );
  XOR2_X1 p_unit_i_1_U22 ( .A(o_data_relu[8]), .B(o_data_relu[10]), .Z(
        p_unit_i_1_N2) );
  XOR2_X1 p_unit_i_1_U21 ( .A(o_data_relu[11]), .B(o_data_relu[9]), .Z(
        p_unit_i_1_n15) );
  XOR2_X1 p_unit_i_1_U19 ( .A(p_unit_i_1_int_ps1_0_), .B(p_unit_i_1_int_ps0_0_), .Z(p_unit_i_1_N5) );
  XOR2_X1 p_unit_i_1_U16 ( .A(p_unit_i_1_int_ps1_2_), .B(p_unit_i_1_int_ps0_2_), .Z(p_unit_i_1_n9) );
  DFFR_X1 p_unit_i_1_int_ps1_reg_2_ ( .D(p_unit_i_1_int_ps0_2_), .CK(
        p_unit_i_1_net3077), .RN(p_unit_i_1_n11), .Q(p_unit_i_1_int_ps1_2_), 
        .QN(p_unit_i_1_n7) );
  DFFR_X1 p_unit_i_1_int_ps0_reg_0_ ( .D(p_unit_i_1_N2), .CK(
        p_unit_i_1_net3077), .RN(p_unit_i_1_n11), .Q(p_unit_i_1_int_ps0_0_) );
  DFFR_X1 p_unit_i_1_int_ps0_reg_1_ ( .D(p_unit_i_1_N3), .CK(
        p_unit_i_1_net3077), .RN(p_unit_i_1_n11), .Q(p_unit_i_1_int_ps0_1_) );
  DFFR_X1 p_unit_i_1_int_ps0_reg_2_ ( .D(p_unit_i_1_n12), .CK(
        p_unit_i_1_net3077), .RN(p_unit_i_1_n11), .Q(p_unit_i_1_int_ps0_2_), 
        .QN(p_unit_i_1_n5) );
  CLKGATETST_X1 p_unit_i_1_clk_gate_o_data_reg_latch ( .CK(ck), .E(
        ps_ctrl_en_p), .SE(1'b0), .GCK(p_unit_i_1_net3077) );
  INV_X1 p_unit_i_2_U18 ( .A(rst), .ZN(p_unit_i_2_n11) );
  INV_X1 p_unit_i_2_U17 ( .A(p_unit_i_2_n8), .ZN(p_unit_i_2_n16) );
  NOR2_X1 p_unit_i_2_U15 ( .A1(p_unit_i_2_int_ps0_2_), .A2(p_unit_i_2_n16), 
        .ZN(p_unit_i_2_n6) );
  OAI22_X1 p_unit_i_2_U14 ( .A1(p_unit_i_2_n8), .A2(p_unit_i_2_n5), .B1(
        p_unit_i_2_n6), .B2(p_unit_i_2_n7), .ZN(p_unit_i_2_n4) );
  OAI211_X1 p_unit_i_2_U13 ( .C1(p_unit_i_2_int_ps0_1_), .C2(
        p_unit_i_2_int_ps1_1_), .A(p_unit_i_2_int_ps0_0_), .B(
        p_unit_i_2_int_ps1_0_), .ZN(p_unit_i_2_n10) );
  INV_X1 p_unit_i_2_U12 ( .A(p_unit_i_2_n10), .ZN(p_unit_i_2_n17) );
  AOI21_X1 p_unit_i_2_U11 ( .B1(p_unit_i_2_int_ps0_1_), .B2(
        p_unit_i_2_int_ps1_1_), .A(p_unit_i_2_n17), .ZN(p_unit_i_2_n8) );
  XNOR2_X1 p_unit_i_2_U10 ( .A(p_unit_i_2_n8), .B(p_unit_i_2_n9), .ZN(
        p_unit_i_2_N7) );
  XNOR2_X1 p_unit_i_2_U9 ( .A(p_unit_i_2_int_ps1_1_), .B(p_unit_i_2_int_ps0_1_), .ZN(p_unit_i_2_n3) );
  NAND2_X1 p_unit_i_2_U8 ( .A1(p_unit_i_2_int_ps0_0_), .A2(
        p_unit_i_2_int_ps1_0_), .ZN(p_unit_i_2_n2) );
  XOR2_X1 p_unit_i_2_U7 ( .A(p_unit_i_2_n2), .B(p_unit_i_2_n3), .Z(
        p_unit_i_2_N6) );
  AND3_X1 p_unit_i_2_U6 ( .A1(o_data_relu[6]), .A2(p_unit_i_2_n15), .A3(
        o_data_relu[4]), .ZN(p_unit_i_2_n14) );
  AOI21_X1 p_unit_i_2_U5 ( .B1(o_data_relu[5]), .B2(o_data_relu[7]), .A(
        p_unit_i_2_n14), .ZN(p_unit_i_2_n13) );
  INV_X1 p_unit_i_2_U4 ( .A(p_unit_i_2_n13), .ZN(p_unit_i_2_n12) );
  NAND2_X1 p_unit_i_2_U3 ( .A1(o_data_relu[6]), .A2(o_data_relu[4]), .ZN(
        p_unit_i_2_n1) );
  XNOR2_X1 p_unit_i_2_U2 ( .A(p_unit_i_2_n1), .B(p_unit_i_2_n15), .ZN(
        p_unit_i_2_N3) );
  DFFR_X1 p_unit_i_2_o_data_reg_3_ ( .D(p_unit_i_2_n4), .CK(p_unit_i_2_net3059), .RN(p_unit_i_2_n11), .Q(int_o_data_p[7]) );
  DFFR_X1 p_unit_i_2_o_data_reg_2_ ( .D(p_unit_i_2_N7), .CK(p_unit_i_2_net3059), .RN(p_unit_i_2_n11), .Q(int_o_data_p[6]) );
  DFFR_X1 p_unit_i_2_o_data_reg_1_ ( .D(p_unit_i_2_N6), .CK(p_unit_i_2_net3059), .RN(p_unit_i_2_n11), .Q(int_o_data_p[5]) );
  DFFR_X1 p_unit_i_2_o_data_reg_0_ ( .D(p_unit_i_2_N5), .CK(p_unit_i_2_net3059), .RN(p_unit_i_2_n11), .Q(int_o_data_p[4]) );
  DFFR_X1 p_unit_i_2_int_ps1_reg_1_ ( .D(p_unit_i_2_int_ps0_1_), .CK(
        p_unit_i_2_net3059), .RN(p_unit_i_2_n11), .Q(p_unit_i_2_int_ps1_1_) );
  DFFR_X1 p_unit_i_2_int_ps1_reg_0_ ( .D(p_unit_i_2_int_ps0_0_), .CK(
        p_unit_i_2_net3059), .RN(p_unit_i_2_n11), .Q(p_unit_i_2_int_ps1_0_) );
  XOR2_X1 p_unit_i_2_U22 ( .A(o_data_relu[4]), .B(o_data_relu[6]), .Z(
        p_unit_i_2_N2) );
  XOR2_X1 p_unit_i_2_U21 ( .A(o_data_relu[7]), .B(o_data_relu[5]), .Z(
        p_unit_i_2_n15) );
  XOR2_X1 p_unit_i_2_U19 ( .A(p_unit_i_2_int_ps1_0_), .B(p_unit_i_2_int_ps0_0_), .Z(p_unit_i_2_N5) );
  XOR2_X1 p_unit_i_2_U16 ( .A(p_unit_i_2_int_ps1_2_), .B(p_unit_i_2_int_ps0_2_), .Z(p_unit_i_2_n9) );
  DFFR_X1 p_unit_i_2_int_ps1_reg_2_ ( .D(p_unit_i_2_int_ps0_2_), .CK(
        p_unit_i_2_net3059), .RN(p_unit_i_2_n11), .Q(p_unit_i_2_int_ps1_2_), 
        .QN(p_unit_i_2_n7) );
  DFFR_X1 p_unit_i_2_int_ps0_reg_0_ ( .D(p_unit_i_2_N2), .CK(
        p_unit_i_2_net3059), .RN(p_unit_i_2_n11), .Q(p_unit_i_2_int_ps0_0_) );
  DFFR_X1 p_unit_i_2_int_ps0_reg_1_ ( .D(p_unit_i_2_N3), .CK(
        p_unit_i_2_net3059), .RN(p_unit_i_2_n11), .Q(p_unit_i_2_int_ps0_1_) );
  DFFR_X1 p_unit_i_2_int_ps0_reg_2_ ( .D(p_unit_i_2_n12), .CK(
        p_unit_i_2_net3059), .RN(p_unit_i_2_n11), .Q(p_unit_i_2_int_ps0_2_), 
        .QN(p_unit_i_2_n5) );
  CLKGATETST_X1 p_unit_i_2_clk_gate_o_data_reg_latch ( .CK(ck), .E(
        ps_ctrl_en_p), .SE(1'b0), .GCK(p_unit_i_2_net3059) );
  INV_X1 p_unit_i_3_U18 ( .A(rst), .ZN(p_unit_i_3_n11) );
  INV_X1 p_unit_i_3_U17 ( .A(p_unit_i_3_n8), .ZN(p_unit_i_3_n16) );
  NOR2_X1 p_unit_i_3_U15 ( .A1(p_unit_i_3_int_ps0_2_), .A2(p_unit_i_3_n16), 
        .ZN(p_unit_i_3_n6) );
  OAI22_X1 p_unit_i_3_U14 ( .A1(p_unit_i_3_n8), .A2(p_unit_i_3_n5), .B1(
        p_unit_i_3_n6), .B2(p_unit_i_3_n7), .ZN(p_unit_i_3_n4) );
  OAI211_X1 p_unit_i_3_U13 ( .C1(p_unit_i_3_int_ps0_1_), .C2(
        p_unit_i_3_int_ps1_1_), .A(p_unit_i_3_int_ps0_0_), .B(
        p_unit_i_3_int_ps1_0_), .ZN(p_unit_i_3_n10) );
  INV_X1 p_unit_i_3_U12 ( .A(p_unit_i_3_n10), .ZN(p_unit_i_3_n17) );
  AOI21_X1 p_unit_i_3_U11 ( .B1(p_unit_i_3_int_ps0_1_), .B2(
        p_unit_i_3_int_ps1_1_), .A(p_unit_i_3_n17), .ZN(p_unit_i_3_n8) );
  XNOR2_X1 p_unit_i_3_U10 ( .A(p_unit_i_3_n8), .B(p_unit_i_3_n9), .ZN(
        p_unit_i_3_N7) );
  XNOR2_X1 p_unit_i_3_U9 ( .A(p_unit_i_3_int_ps1_1_), .B(p_unit_i_3_int_ps0_1_), .ZN(p_unit_i_3_n3) );
  NAND2_X1 p_unit_i_3_U8 ( .A1(p_unit_i_3_int_ps0_0_), .A2(
        p_unit_i_3_int_ps1_0_), .ZN(p_unit_i_3_n2) );
  XOR2_X1 p_unit_i_3_U7 ( .A(p_unit_i_3_n2), .B(p_unit_i_3_n3), .Z(
        p_unit_i_3_N6) );
  AND3_X1 p_unit_i_3_U6 ( .A1(o_data_relu[2]), .A2(p_unit_i_3_n15), .A3(
        o_data_relu[0]), .ZN(p_unit_i_3_n14) );
  AOI21_X1 p_unit_i_3_U5 ( .B1(o_data_relu[1]), .B2(o_data_relu[3]), .A(
        p_unit_i_3_n14), .ZN(p_unit_i_3_n13) );
  INV_X1 p_unit_i_3_U4 ( .A(p_unit_i_3_n13), .ZN(p_unit_i_3_n12) );
  NAND2_X1 p_unit_i_3_U3 ( .A1(o_data_relu[2]), .A2(o_data_relu[0]), .ZN(
        p_unit_i_3_n1) );
  XNOR2_X1 p_unit_i_3_U2 ( .A(p_unit_i_3_n1), .B(p_unit_i_3_n15), .ZN(
        p_unit_i_3_N3) );
  DFFR_X1 p_unit_i_3_o_data_reg_3_ ( .D(p_unit_i_3_n4), .CK(p_unit_i_3_net3041), .RN(p_unit_i_3_n11), .Q(int_o_data_p[3]) );
  DFFR_X1 p_unit_i_3_o_data_reg_2_ ( .D(p_unit_i_3_N7), .CK(p_unit_i_3_net3041), .RN(p_unit_i_3_n11), .Q(int_o_data_p[2]) );
  DFFR_X1 p_unit_i_3_o_data_reg_1_ ( .D(p_unit_i_3_N6), .CK(p_unit_i_3_net3041), .RN(p_unit_i_3_n11), .Q(int_o_data_p[1]) );
  DFFR_X1 p_unit_i_3_o_data_reg_0_ ( .D(p_unit_i_3_N5), .CK(p_unit_i_3_net3041), .RN(p_unit_i_3_n11), .Q(int_o_data_p[0]) );
  DFFR_X1 p_unit_i_3_int_ps1_reg_1_ ( .D(p_unit_i_3_int_ps0_1_), .CK(
        p_unit_i_3_net3041), .RN(p_unit_i_3_n11), .Q(p_unit_i_3_int_ps1_1_) );
  DFFR_X1 p_unit_i_3_int_ps1_reg_0_ ( .D(p_unit_i_3_int_ps0_0_), .CK(
        p_unit_i_3_net3041), .RN(p_unit_i_3_n11), .Q(p_unit_i_3_int_ps1_0_) );
  XOR2_X1 p_unit_i_3_U22 ( .A(o_data_relu[0]), .B(o_data_relu[2]), .Z(
        p_unit_i_3_N2) );
  XOR2_X1 p_unit_i_3_U21 ( .A(o_data_relu[3]), .B(o_data_relu[1]), .Z(
        p_unit_i_3_n15) );
  XOR2_X1 p_unit_i_3_U19 ( .A(p_unit_i_3_int_ps1_0_), .B(p_unit_i_3_int_ps0_0_), .Z(p_unit_i_3_N5) );
  XOR2_X1 p_unit_i_3_U16 ( .A(p_unit_i_3_int_ps1_2_), .B(p_unit_i_3_int_ps0_2_), .Z(p_unit_i_3_n9) );
  DFFR_X1 p_unit_i_3_int_ps1_reg_2_ ( .D(p_unit_i_3_int_ps0_2_), .CK(
        p_unit_i_3_net3041), .RN(p_unit_i_3_n11), .Q(p_unit_i_3_int_ps1_2_), 
        .QN(p_unit_i_3_n7) );
  DFFR_X1 p_unit_i_3_int_ps0_reg_0_ ( .D(p_unit_i_3_N2), .CK(
        p_unit_i_3_net3041), .RN(p_unit_i_3_n11), .Q(p_unit_i_3_int_ps0_0_) );
  DFFR_X1 p_unit_i_3_int_ps0_reg_1_ ( .D(p_unit_i_3_N3), .CK(
        p_unit_i_3_net3041), .RN(p_unit_i_3_n11), .Q(p_unit_i_3_int_ps0_1_) );
  DFFR_X1 p_unit_i_3_int_ps0_reg_2_ ( .D(p_unit_i_3_n12), .CK(
        p_unit_i_3_net3041), .RN(p_unit_i_3_n11), .Q(p_unit_i_3_int_ps0_2_), 
        .QN(p_unit_i_3_n5) );
  CLKGATETST_X1 p_unit_i_3_clk_gate_o_data_reg_latch ( .CK(ck), .E(
        ps_ctrl_en_p), .SE(1'b0), .GCK(p_unit_i_3_net3041) );
  INV_X1 round_i_0_U5 ( .A(int_o_data_p[14]), .ZN(round_i_0_n2) );
  OAI21_X1 round_i_0_U4 ( .B1(int_o_data_p[13]), .B2(round_i_0_n2), .A(
        round_i_0_n3), .ZN(o_data[6]) );
  NAND2_X1 round_i_0_U3 ( .A1(int_o_data_p[13]), .A2(int_o_data_p[14]), .ZN(
        round_i_0_n1) );
  XNOR2_X1 round_i_0_U2 ( .A(int_o_data_p[15]), .B(round_i_0_n1), .ZN(
        o_data[7]) );
  NAND3_X1 round_i_0_U6 ( .A1(int_o_data_p[13]), .A2(round_i_0_n2), .A3(
        int_o_data_p[12]), .ZN(round_i_0_n3) );
  INV_X1 round_i_1_U5 ( .A(int_o_data_p[10]), .ZN(round_i_1_n2) );
  OAI21_X1 round_i_1_U4 ( .B1(int_o_data_p[9]), .B2(round_i_1_n2), .A(
        round_i_1_n4), .ZN(o_data[4]) );
  NAND2_X1 round_i_1_U3 ( .A1(int_o_data_p[9]), .A2(int_o_data_p[10]), .ZN(
        round_i_1_n1) );
  XNOR2_X1 round_i_1_U2 ( .A(int_o_data_p[11]), .B(round_i_1_n1), .ZN(
        o_data[5]) );
  NAND3_X1 round_i_1_U6 ( .A1(int_o_data_p[9]), .A2(round_i_1_n2), .A3(
        int_o_data_p[8]), .ZN(round_i_1_n4) );
  INV_X1 round_i_2_U5 ( .A(int_o_data_p[6]), .ZN(round_i_2_n2) );
  OAI21_X1 round_i_2_U4 ( .B1(int_o_data_p[5]), .B2(round_i_2_n2), .A(
        round_i_2_n4), .ZN(o_data[2]) );
  NAND2_X1 round_i_2_U3 ( .A1(int_o_data_p[5]), .A2(int_o_data_p[6]), .ZN(
        round_i_2_n1) );
  XNOR2_X1 round_i_2_U2 ( .A(int_o_data_p[7]), .B(round_i_2_n1), .ZN(o_data[3]) );
  NAND3_X1 round_i_2_U6 ( .A1(int_o_data_p[5]), .A2(round_i_2_n2), .A3(
        int_o_data_p[4]), .ZN(round_i_2_n4) );
  INV_X1 round_i_3_U5 ( .A(int_o_data_p[2]), .ZN(round_i_3_n2) );
  OAI21_X1 round_i_3_U4 ( .B1(int_o_data_p[1]), .B2(round_i_3_n2), .A(
        round_i_3_n4), .ZN(o_data[0]) );
  NAND2_X1 round_i_3_U3 ( .A1(int_o_data_p[1]), .A2(int_o_data_p[2]), .ZN(
        round_i_3_n1) );
  XNOR2_X1 round_i_3_U2 ( .A(int_o_data_p[3]), .B(round_i_3_n1), .ZN(o_data[1]) );
  NAND3_X1 round_i_3_U6 ( .A1(int_o_data_p[1]), .A2(round_i_3_n2), .A3(
        int_o_data_p[0]), .ZN(round_i_3_n4) );
  INV_X1 hmode_cnt_inst_U14 ( .A(rst), .ZN(hmode_cnt_inst_n12) );
  AOI21_X1 hmode_cnt_inst_U13 ( .B1(hmode_cnt_inst_n10), .B2(hmode_cnt_inst_n7), .A(hmode_cnt_inst_N10), .ZN(hmode_cnt_inst_n8) );
  NAND4_X1 hmode_cnt_inst_U12 ( .A1(hmode_cnt_inst_n10), .A2(int_hmode_cnt[1]), 
        .A3(int_hmode_cnt[0]), .A4(hmode_cnt_inst_n5), .ZN(hmode_cnt_inst_n9)
         );
  OAI21_X1 hmode_cnt_inst_U11 ( .B1(hmode_cnt_inst_n8), .B2(hmode_cnt_inst_n5), 
        .A(hmode_cnt_inst_n9), .ZN(hmode_cnt_inst_N12) );
  XNOR2_X1 hmode_cnt_inst_U10 ( .A(int_hmode_cnt[0]), .B(int_hmode_cnt[1]), 
        .ZN(hmode_cnt_inst_n11) );
  AND2_X1 hmode_cnt_inst_U9 ( .A1(hmode_cnt_inst_n10), .A2(hmode_cnt_inst_n6), 
        .ZN(hmode_cnt_inst_N10) );
  NOR2_X1 hmode_cnt_inst_U8 ( .A1(s_tc_hmode), .A2(1'b0), .ZN(
        hmode_cnt_inst_n10) );
  XOR2_X1 hmode_cnt_inst_U7 ( .A(int_hmode_cnt[1]), .B(arv_KSI[1]), .Z(
        hmode_cnt_inst_n4) );
  XOR2_X1 hmode_cnt_inst_U6 ( .A(int_hmode_cnt[0]), .B(arv_KSI[0]), .Z(
        hmode_cnt_inst_n2) );
  XOR2_X1 hmode_cnt_inst_U5 ( .A(int_hmode_cnt[2]), .B(arv_KSI[2]), .Z(
        hmode_cnt_inst_n1) );
  NOR3_X1 hmode_cnt_inst_U4 ( .A1(hmode_cnt_inst_n1), .A2(hmode_cnt_inst_n2), 
        .A3(hmode_cnt_inst_n4), .ZN(s_tc_hmode) );
  DFFR_X1 hmode_cnt_inst_cnt_out_reg_2_ ( .D(hmode_cnt_inst_N12), .CK(
        hmode_cnt_inst_net3023), .RN(hmode_cnt_inst_n12), .Q(int_hmode_cnt[2]), 
        .QN(hmode_cnt_inst_n5) );
  SDFFR_X1 hmode_cnt_inst_cnt_out_reg_1_ ( .D(hmode_cnt_inst_n10), .SI(1'b0), 
        .SE(hmode_cnt_inst_n11), .CK(hmode_cnt_inst_net3023), .RN(
        hmode_cnt_inst_n12), .Q(int_hmode_cnt[1]), .QN(hmode_cnt_inst_n7) );
  DFFR_X1 hmode_cnt_inst_cnt_out_reg_0_ ( .D(hmode_cnt_inst_N10), .CK(
        hmode_cnt_inst_net3023), .RN(hmode_cnt_inst_n12), .Q(int_hmode_cnt[0]), 
        .QN(hmode_cnt_inst_n6) );
  CLKGATETST_X1 hmode_cnt_inst_clk_gate_cnt_out_reg_latch ( .CK(ck), .E(
        int_en_hmode), .SE(1'b0), .GCK(hmode_cnt_inst_net3023) );
  INV_X1 vmode_cnt_inst_U14 ( .A(rst), .ZN(vmode_cnt_inst_n12) );
  AOI21_X1 vmode_cnt_inst_U13 ( .B1(vmode_cnt_inst_n10), .B2(vmode_cnt_inst_n7), .A(vmode_cnt_inst_N10), .ZN(vmode_cnt_inst_n8) );
  NAND4_X1 vmode_cnt_inst_U12 ( .A1(vmode_cnt_inst_n10), .A2(
        vmode_cnt_inst_q_1_), .A3(vmode_cnt_inst_q_0_), .A4(vmode_cnt_inst_n5), 
        .ZN(vmode_cnt_inst_n9) );
  OAI21_X1 vmode_cnt_inst_U11 ( .B1(vmode_cnt_inst_n8), .B2(vmode_cnt_inst_n5), 
        .A(vmode_cnt_inst_n9), .ZN(vmode_cnt_inst_N12) );
  XNOR2_X1 vmode_cnt_inst_U10 ( .A(vmode_cnt_inst_q_0_), .B(
        vmode_cnt_inst_q_1_), .ZN(vmode_cnt_inst_n11) );
  AND2_X1 vmode_cnt_inst_U9 ( .A1(vmode_cnt_inst_n10), .A2(vmode_cnt_inst_n6), 
        .ZN(vmode_cnt_inst_N10) );
  NOR2_X1 vmode_cnt_inst_U8 ( .A1(s_tc_vmode), .A2(1'b0), .ZN(
        vmode_cnt_inst_n10) );
  XOR2_X1 vmode_cnt_inst_U7 ( .A(vmode_cnt_inst_q_1_), .B(arv_KSI[1]), .Z(
        vmode_cnt_inst_n4) );
  XOR2_X1 vmode_cnt_inst_U6 ( .A(vmode_cnt_inst_q_0_), .B(arv_KSI[0]), .Z(
        vmode_cnt_inst_n2) );
  XOR2_X1 vmode_cnt_inst_U5 ( .A(vmode_cnt_inst_q_2_), .B(arv_KSI[2]), .Z(
        vmode_cnt_inst_n1) );
  NOR3_X1 vmode_cnt_inst_U4 ( .A1(vmode_cnt_inst_n1), .A2(vmode_cnt_inst_n2), 
        .A3(vmode_cnt_inst_n4), .ZN(s_tc_vmode) );
  DFFR_X1 vmode_cnt_inst_cnt_out_reg_2_ ( .D(vmode_cnt_inst_N12), .CK(
        vmode_cnt_inst_net3005), .RN(vmode_cnt_inst_n12), .Q(
        vmode_cnt_inst_q_2_), .QN(vmode_cnt_inst_n5) );
  SDFFR_X1 vmode_cnt_inst_cnt_out_reg_1_ ( .D(vmode_cnt_inst_n10), .SI(1'b0), 
        .SE(vmode_cnt_inst_n11), .CK(vmode_cnt_inst_net3005), .RN(
        vmode_cnt_inst_n12), .Q(vmode_cnt_inst_q_1_), .QN(vmode_cnt_inst_n7)
         );
  DFFR_X1 vmode_cnt_inst_cnt_out_reg_0_ ( .D(vmode_cnt_inst_N10), .CK(
        vmode_cnt_inst_net3005), .RN(vmode_cnt_inst_n12), .Q(
        vmode_cnt_inst_q_0_), .QN(vmode_cnt_inst_n6) );
  CLKGATETST_X1 vmode_cnt_inst_clk_gate_cnt_out_reg_latch ( .CK(ck), .E(
        int_en_vmode), .SE(1'b0), .GCK(vmode_cnt_inst_net3005) );
  INV_X1 res_cnt_inst_U14 ( .A(rst), .ZN(res_cnt_inst_n2) );
  XNOR2_X1 res_cnt_inst_U13 ( .A(res_cnt_inst_q_0_), .B(res_cnt_inst_q_1_), 
        .ZN(res_cnt_inst_n11) );
  AND2_X1 res_cnt_inst_U12 ( .A1(res_cnt_inst_n10), .A2(res_cnt_inst_n1), .ZN(
        res_cnt_inst_N10) );
  AOI21_X1 res_cnt_inst_U11 ( .B1(res_cnt_inst_n10), .B2(res_cnt_inst_n7), .A(
        res_cnt_inst_N10), .ZN(res_cnt_inst_n8) );
  NAND4_X1 res_cnt_inst_U10 ( .A1(res_cnt_inst_n10), .A2(res_cnt_inst_q_1_), 
        .A3(res_cnt_inst_q_0_), .A4(res_cnt_inst_n5), .ZN(res_cnt_inst_n9) );
  OAI21_X1 res_cnt_inst_U9 ( .B1(res_cnt_inst_n8), .B2(res_cnt_inst_n5), .A(
        res_cnt_inst_n9), .ZN(res_cnt_inst_N12) );
  XNOR2_X1 res_cnt_inst_U8 ( .A(res_cnt_inst_q_1_), .B(int_arv_res[1]), .ZN(
        res_cnt_inst_n14) );
  XNOR2_X1 res_cnt_inst_U7 ( .A(res_cnt_inst_q_0_), .B(int_arv_res[0]), .ZN(
        res_cnt_inst_n13) );
  XNOR2_X1 res_cnt_inst_U6 ( .A(res_cnt_inst_q_2_), .B(int_arv_res[2]), .ZN(
        res_cnt_inst_n12) );
  AND3_X1 res_cnt_inst_U5 ( .A1(res_cnt_inst_n12), .A2(res_cnt_inst_n13), .A3(
        res_cnt_inst_n14), .ZN(s_tc_res) );
  NOR2_X1 res_cnt_inst_U4 ( .A1(s_tc_res), .A2(1'b0), .ZN(res_cnt_inst_n10) );
  DFFR_X1 res_cnt_inst_cnt_out_reg_2_ ( .D(res_cnt_inst_N12), .CK(
        res_cnt_inst_net2987), .RN(res_cnt_inst_n2), .Q(res_cnt_inst_q_2_), 
        .QN(res_cnt_inst_n5) );
  SDFFR_X1 res_cnt_inst_cnt_out_reg_1_ ( .D(res_cnt_inst_n10), .SI(1'b0), .SE(
        res_cnt_inst_n11), .CK(res_cnt_inst_net2987), .RN(res_cnt_inst_n2), 
        .Q(res_cnt_inst_q_1_), .QN(res_cnt_inst_n7) );
  DFFR_X1 res_cnt_inst_cnt_out_reg_0_ ( .D(res_cnt_inst_N10), .CK(
        res_cnt_inst_net2987), .RN(res_cnt_inst_n2), .Q(res_cnt_inst_q_0_), 
        .QN(res_cnt_inst_n1) );
  CLKGATETST_X1 res_cnt_inst_clk_gate_cnt_out_reg_latch ( .CK(ck), .E(
        ctrl_wr_pipe), .SE(1'b0), .GCK(res_cnt_inst_net2987) );
  INV_X1 i_data_npu_cnt_inst_U17 ( .A(rst), .ZN(i_data_npu_cnt_inst_n2) );
  XNOR2_X1 i_data_npu_cnt_inst_U16 ( .A(int_L1_ptr[0]), .B(int_L1_ptr[1]), 
        .ZN(i_data_npu_cnt_inst_n15) );
  XNOR2_X1 i_data_npu_cnt_inst_U15 ( .A(i_data_npu_cnt_inst_q_3_), .B(
        arv_L1[3]), .ZN(i_data_npu_cnt_inst_n18) );
  XNOR2_X1 i_data_npu_cnt_inst_U14 ( .A(int_L1_ptr[2]), .B(arv_L1[2]), .ZN(
        i_data_npu_cnt_inst_n17) );
  AND4_X1 i_data_npu_cnt_inst_U13 ( .A1(i_data_npu_cnt_inst_n16), .A2(
        i_data_npu_cnt_inst_n17), .A3(i_data_npu_cnt_inst_n18), .A4(
        i_data_npu_cnt_inst_n19), .ZN(s_tc_L1) );
  AND2_X1 i_data_npu_cnt_inst_U12 ( .A1(i_data_npu_cnt_inst_n13), .A2(
        i_data_npu_cnt_inst_n1), .ZN(i_data_npu_cnt_inst_N11) );
  INV_X1 i_data_npu_cnt_inst_U11 ( .A(i_data_npu_cnt_inst_n14), .ZN(
        i_data_npu_cnt_inst_n4) );
  AOI21_X1 i_data_npu_cnt_inst_U10 ( .B1(i_data_npu_cnt_inst_n13), .B2(
        i_data_npu_cnt_inst_n8), .A(i_data_npu_cnt_inst_n4), .ZN(
        i_data_npu_cnt_inst_n10) );
  OR3_X1 i_data_npu_cnt_inst_U9 ( .A1(i_data_npu_cnt_inst_n8), .A2(
        i_data_npu_cnt_inst_q_3_), .A3(i_data_npu_cnt_inst_n12), .ZN(
        i_data_npu_cnt_inst_n11) );
  OAI21_X1 i_data_npu_cnt_inst_U8 ( .B1(i_data_npu_cnt_inst_n10), .B2(
        i_data_npu_cnt_inst_n5), .A(i_data_npu_cnt_inst_n11), .ZN(
        i_data_npu_cnt_inst_N14) );
  XNOR2_X1 i_data_npu_cnt_inst_U7 ( .A(int_L1_ptr[0]), .B(arv_L1[0]), .ZN(
        i_data_npu_cnt_inst_n19) );
  OAI22_X1 i_data_npu_cnt_inst_U6 ( .A1(i_data_npu_cnt_inst_n14), .A2(
        i_data_npu_cnt_inst_n8), .B1(int_L1_ptr[2]), .B2(
        i_data_npu_cnt_inst_n12), .ZN(i_data_npu_cnt_inst_N13) );
  AOI21_X1 i_data_npu_cnt_inst_U5 ( .B1(i_data_npu_cnt_inst_n9), .B2(
        i_data_npu_cnt_inst_n13), .A(i_data_npu_cnt_inst_N11), .ZN(
        i_data_npu_cnt_inst_n14) );
  NOR2_X1 i_data_npu_cnt_inst_U4 ( .A1(s_tc_L1), .A2(1'b0), .ZN(
        i_data_npu_cnt_inst_n13) );
  XOR2_X1 i_data_npu_cnt_inst_U20 ( .A(i_data_npu_cnt_inst_n9), .B(arv_L1[1]), 
        .Z(i_data_npu_cnt_inst_n16) );
  NAND3_X1 i_data_npu_cnt_inst_U19 ( .A1(int_L1_ptr[1]), .A2(int_L1_ptr[0]), 
        .A3(i_data_npu_cnt_inst_n13), .ZN(i_data_npu_cnt_inst_n12) );
  DFFR_X1 i_data_npu_cnt_inst_cnt_out_reg_3_ ( .D(i_data_npu_cnt_inst_N14), 
        .CK(i_data_npu_cnt_inst_net2969), .RN(i_data_npu_cnt_inst_n2), .Q(
        i_data_npu_cnt_inst_q_3_), .QN(i_data_npu_cnt_inst_n5) );
  DFFR_X1 i_data_npu_cnt_inst_cnt_out_reg_2_ ( .D(i_data_npu_cnt_inst_N13), 
        .CK(i_data_npu_cnt_inst_net2969), .RN(i_data_npu_cnt_inst_n2), .Q(
        int_L1_ptr[2]), .QN(i_data_npu_cnt_inst_n8) );
  SDFFR_X1 i_data_npu_cnt_inst_cnt_out_reg_1_ ( .D(i_data_npu_cnt_inst_n13), 
        .SI(1'b0), .SE(i_data_npu_cnt_inst_n15), .CK(
        i_data_npu_cnt_inst_net2969), .RN(i_data_npu_cnt_inst_n2), .Q(
        int_L1_ptr[1]), .QN(i_data_npu_cnt_inst_n9) );
  DFFR_X1 i_data_npu_cnt_inst_cnt_out_reg_0_ ( .D(i_data_npu_cnt_inst_N11), 
        .CK(i_data_npu_cnt_inst_net2969), .RN(i_data_npu_cnt_inst_n2), .Q(
        int_L1_ptr[0]), .QN(i_data_npu_cnt_inst_n1) );
  CLKGATETST_X1 i_data_npu_cnt_inst_clk_gate_cnt_out_reg_latch ( .CK(ck), .E(
        int_en_L1_ptr), .SE(1'b0), .GCK(i_data_npu_cnt_inst_net2969) );
  INV_X1 i_data_L2_cnt_inst_U17 ( .A(rst), .ZN(i_data_L2_cnt_inst_n2) );
  XNOR2_X1 i_data_L2_cnt_inst_U16 ( .A(i_data_L2_cnt_inst_q_0_), .B(
        i_data_L2_cnt_inst_q_1_), .ZN(i_data_L2_cnt_inst_n15) );
  XNOR2_X1 i_data_L2_cnt_inst_U15 ( .A(i_data_L2_cnt_inst_q_3_), .B(arv_L2[3]), 
        .ZN(i_data_L2_cnt_inst_n18) );
  XNOR2_X1 i_data_L2_cnt_inst_U14 ( .A(i_data_L2_cnt_inst_q_2_), .B(arv_L2[2]), 
        .ZN(i_data_L2_cnt_inst_n17) );
  AND4_X1 i_data_L2_cnt_inst_U13 ( .A1(i_data_L2_cnt_inst_n16), .A2(
        i_data_L2_cnt_inst_n17), .A3(i_data_L2_cnt_inst_n18), .A4(
        i_data_L2_cnt_inst_n19), .ZN(int_d_tc[2]) );
  INV_X1 i_data_L2_cnt_inst_U12 ( .A(i_data_L2_cnt_inst_n14), .ZN(
        i_data_L2_cnt_inst_n4) );
  AOI21_X1 i_data_L2_cnt_inst_U11 ( .B1(i_data_L2_cnt_inst_n13), .B2(
        i_data_L2_cnt_inst_n8), .A(i_data_L2_cnt_inst_n4), .ZN(
        i_data_L2_cnt_inst_n10) );
  OR3_X1 i_data_L2_cnt_inst_U10 ( .A1(i_data_L2_cnt_inst_n8), .A2(
        i_data_L2_cnt_inst_q_3_), .A3(i_data_L2_cnt_inst_n12), .ZN(
        i_data_L2_cnt_inst_n11) );
  OAI21_X1 i_data_L2_cnt_inst_U9 ( .B1(i_data_L2_cnt_inst_n10), .B2(
        i_data_L2_cnt_inst_n5), .A(i_data_L2_cnt_inst_n11), .ZN(
        i_data_L2_cnt_inst_N14) );
  AND2_X1 i_data_L2_cnt_inst_U8 ( .A1(i_data_L2_cnt_inst_n13), .A2(
        i_data_L2_cnt_inst_n1), .ZN(i_data_L2_cnt_inst_N11) );
  XNOR2_X1 i_data_L2_cnt_inst_U7 ( .A(i_data_L2_cnt_inst_q_0_), .B(arv_L2[0]), 
        .ZN(i_data_L2_cnt_inst_n19) );
  OAI22_X1 i_data_L2_cnt_inst_U6 ( .A1(i_data_L2_cnt_inst_n14), .A2(
        i_data_L2_cnt_inst_n8), .B1(i_data_L2_cnt_inst_q_2_), .B2(
        i_data_L2_cnt_inst_n12), .ZN(i_data_L2_cnt_inst_N13) );
  AOI21_X1 i_data_L2_cnt_inst_U5 ( .B1(i_data_L2_cnt_inst_n9), .B2(
        i_data_L2_cnt_inst_n13), .A(i_data_L2_cnt_inst_N11), .ZN(
        i_data_L2_cnt_inst_n14) );
  NOR2_X1 i_data_L2_cnt_inst_U4 ( .A1(int_d_tc[2]), .A2(1'b0), .ZN(
        i_data_L2_cnt_inst_n13) );
  XOR2_X1 i_data_L2_cnt_inst_U20 ( .A(i_data_L2_cnt_inst_n9), .B(arv_L2[1]), 
        .Z(i_data_L2_cnt_inst_n16) );
  NAND3_X1 i_data_L2_cnt_inst_U19 ( .A1(i_data_L2_cnt_inst_q_1_), .A2(
        i_data_L2_cnt_inst_q_0_), .A3(i_data_L2_cnt_inst_n13), .ZN(
        i_data_L2_cnt_inst_n12) );
  DFFR_X1 i_data_L2_cnt_inst_cnt_out_reg_3_ ( .D(i_data_L2_cnt_inst_N14), .CK(
        i_data_L2_cnt_inst_net2951), .RN(i_data_L2_cnt_inst_n2), .Q(
        i_data_L2_cnt_inst_q_3_), .QN(i_data_L2_cnt_inst_n5) );
  DFFR_X1 i_data_L2_cnt_inst_cnt_out_reg_2_ ( .D(i_data_L2_cnt_inst_N13), .CK(
        i_data_L2_cnt_inst_net2951), .RN(i_data_L2_cnt_inst_n2), .Q(
        i_data_L2_cnt_inst_q_2_), .QN(i_data_L2_cnt_inst_n8) );
  SDFFR_X1 i_data_L2_cnt_inst_cnt_out_reg_1_ ( .D(i_data_L2_cnt_inst_n13), 
        .SI(1'b0), .SE(i_data_L2_cnt_inst_n15), .CK(i_data_L2_cnt_inst_net2951), .RN(i_data_L2_cnt_inst_n2), .Q(i_data_L2_cnt_inst_q_1_), .QN(
        i_data_L2_cnt_inst_n9) );
  DFFR_X1 i_data_L2_cnt_inst_cnt_out_reg_0_ ( .D(i_data_L2_cnt_inst_N11), .CK(
        i_data_L2_cnt_inst_net2951), .RN(i_data_L2_cnt_inst_n2), .Q(
        i_data_L2_cnt_inst_q_0_), .QN(i_data_L2_cnt_inst_n1) );
  CLKGATETST_X1 i_data_L2_cnt_inst_clk_gate_cnt_out_reg_latch ( .CK(ck), .E(
        int_en_L2_ptr), .SE(1'b0), .GCK(i_data_L2_cnt_inst_net2951) );
  INV_X1 i_data_L3_cnt_inst_U17 ( .A(rst), .ZN(i_data_L3_cnt_inst_n2) );
  XNOR2_X1 i_data_L3_cnt_inst_U16 ( .A(i_data_ev_odd_n), .B(int_L3_ptr_1_), 
        .ZN(i_data_L3_cnt_inst_n15) );
  XNOR2_X1 i_data_L3_cnt_inst_U15 ( .A(i_data_L3_cnt_inst_q_3_), .B(arv_L3[3]), 
        .ZN(i_data_L3_cnt_inst_n18) );
  XNOR2_X1 i_data_L3_cnt_inst_U14 ( .A(i_data_L3_cnt_inst_q_2_), .B(arv_L3[2]), 
        .ZN(i_data_L3_cnt_inst_n17) );
  AND4_X1 i_data_L3_cnt_inst_U13 ( .A1(i_data_L3_cnt_inst_n16), .A2(
        i_data_L3_cnt_inst_n17), .A3(i_data_L3_cnt_inst_n18), .A4(
        i_data_L3_cnt_inst_n19), .ZN(int_d_tc[1]) );
  AND2_X1 i_data_L3_cnt_inst_U12 ( .A1(i_data_L3_cnt_inst_n13), .A2(
        i_data_L3_cnt_inst_n1), .ZN(i_data_L3_cnt_inst_N11) );
  INV_X1 i_data_L3_cnt_inst_U11 ( .A(i_data_L3_cnt_inst_n14), .ZN(
        i_data_L3_cnt_inst_n4) );
  AOI21_X1 i_data_L3_cnt_inst_U10 ( .B1(i_data_L3_cnt_inst_n13), .B2(
        i_data_L3_cnt_inst_n8), .A(i_data_L3_cnt_inst_n4), .ZN(
        i_data_L3_cnt_inst_n10) );
  OR3_X1 i_data_L3_cnt_inst_U9 ( .A1(i_data_L3_cnt_inst_n8), .A2(
        i_data_L3_cnt_inst_q_3_), .A3(i_data_L3_cnt_inst_n12), .ZN(
        i_data_L3_cnt_inst_n11) );
  OAI21_X1 i_data_L3_cnt_inst_U8 ( .B1(i_data_L3_cnt_inst_n10), .B2(
        i_data_L3_cnt_inst_n5), .A(i_data_L3_cnt_inst_n11), .ZN(
        i_data_L3_cnt_inst_N14) );
  XNOR2_X1 i_data_L3_cnt_inst_U7 ( .A(i_data_ev_odd_n), .B(arv_L3[0]), .ZN(
        i_data_L3_cnt_inst_n19) );
  OAI22_X1 i_data_L3_cnt_inst_U6 ( .A1(i_data_L3_cnt_inst_n14), .A2(
        i_data_L3_cnt_inst_n8), .B1(i_data_L3_cnt_inst_q_2_), .B2(
        i_data_L3_cnt_inst_n12), .ZN(i_data_L3_cnt_inst_N13) );
  AOI21_X1 i_data_L3_cnt_inst_U5 ( .B1(i_data_L3_cnt_inst_n9), .B2(
        i_data_L3_cnt_inst_n13), .A(i_data_L3_cnt_inst_N11), .ZN(
        i_data_L3_cnt_inst_n14) );
  NOR2_X1 i_data_L3_cnt_inst_U4 ( .A1(int_d_tc[1]), .A2(1'b0), .ZN(
        i_data_L3_cnt_inst_n13) );
  XOR2_X1 i_data_L3_cnt_inst_U20 ( .A(i_data_L3_cnt_inst_n9), .B(arv_L3[1]), 
        .Z(i_data_L3_cnt_inst_n16) );
  NAND3_X1 i_data_L3_cnt_inst_U19 ( .A1(int_L3_ptr_1_), .A2(i_data_ev_odd_n), 
        .A3(i_data_L3_cnt_inst_n13), .ZN(i_data_L3_cnt_inst_n12) );
  DFFR_X1 i_data_L3_cnt_inst_cnt_out_reg_3_ ( .D(i_data_L3_cnt_inst_N14), .CK(
        i_data_L3_cnt_inst_net2933), .RN(i_data_L3_cnt_inst_n2), .Q(
        i_data_L3_cnt_inst_q_3_), .QN(i_data_L3_cnt_inst_n5) );
  DFFR_X1 i_data_L3_cnt_inst_cnt_out_reg_2_ ( .D(i_data_L3_cnt_inst_N13), .CK(
        i_data_L3_cnt_inst_net2933), .RN(i_data_L3_cnt_inst_n2), .Q(
        i_data_L3_cnt_inst_q_2_), .QN(i_data_L3_cnt_inst_n8) );
  SDFFR_X1 i_data_L3_cnt_inst_cnt_out_reg_1_ ( .D(i_data_L3_cnt_inst_n13), 
        .SI(1'b0), .SE(i_data_L3_cnt_inst_n15), .CK(i_data_L3_cnt_inst_net2933), .RN(i_data_L3_cnt_inst_n2), .Q(int_L3_ptr_1_), .QN(i_data_L3_cnt_inst_n9) );
  DFFR_X1 i_data_L3_cnt_inst_cnt_out_reg_0_ ( .D(i_data_L3_cnt_inst_N11), .CK(
        i_data_L3_cnt_inst_net2933), .RN(i_data_L3_cnt_inst_n2), .Q(
        i_data_ev_odd_n), .QN(i_data_L3_cnt_inst_n1) );
  CLKGATETST_X1 i_data_L3_cnt_inst_clk_gate_cnt_out_reg_latch ( .CK(ck), .E(
        n33), .SE(1'b0), .GCK(i_data_L3_cnt_inst_net2933) );
  INV_X1 L0_cnt_inst_U17 ( .A(rst), .ZN(L0_cnt_inst_n2) );
  XNOR2_X1 L0_cnt_inst_U16 ( .A(int_L0_ptr[0]), .B(int_L0_ptr[1]), .ZN(
        L0_cnt_inst_n15) );
  INV_X1 L0_cnt_inst_U15 ( .A(L0_cnt_inst_n14), .ZN(L0_cnt_inst_n4) );
  AOI21_X1 L0_cnt_inst_U14 ( .B1(L0_cnt_inst_n13), .B2(L0_cnt_inst_n8), .A(
        L0_cnt_inst_n4), .ZN(L0_cnt_inst_n10) );
  OR3_X1 L0_cnt_inst_U13 ( .A1(L0_cnt_inst_n8), .A2(L0_cnt_inst_q_3_), .A3(
        L0_cnt_inst_n12), .ZN(L0_cnt_inst_n11) );
  OAI21_X1 L0_cnt_inst_U12 ( .B1(L0_cnt_inst_n10), .B2(L0_cnt_inst_n5), .A(
        L0_cnt_inst_n11), .ZN(L0_cnt_inst_N14) );
  XNOR2_X1 L0_cnt_inst_U11 ( .A(L0_cnt_inst_q_3_), .B(arv_L0[3]), .ZN(
        L0_cnt_inst_n18) );
  XNOR2_X1 L0_cnt_inst_U10 ( .A(int_L0_ptr[2]), .B(arv_L0[2]), .ZN(
        L0_cnt_inst_n17) );
  AND4_X1 L0_cnt_inst_U9 ( .A1(L0_cnt_inst_n16), .A2(L0_cnt_inst_n17), .A3(
        L0_cnt_inst_n18), .A4(L0_cnt_inst_n19), .ZN(s_tc_L0) );
  AND2_X1 L0_cnt_inst_U8 ( .A1(L0_cnt_inst_n13), .A2(L0_cnt_inst_n1), .ZN(
        L0_cnt_inst_N11) );
  XNOR2_X1 L0_cnt_inst_U7 ( .A(int_L0_ptr[0]), .B(arv_L0[0]), .ZN(
        L0_cnt_inst_n19) );
  OAI22_X1 L0_cnt_inst_U6 ( .A1(L0_cnt_inst_n14), .A2(L0_cnt_inst_n8), .B1(
        int_L0_ptr[2]), .B2(L0_cnt_inst_n12), .ZN(L0_cnt_inst_N13) );
  AOI21_X1 L0_cnt_inst_U5 ( .B1(L0_cnt_inst_n9), .B2(L0_cnt_inst_n13), .A(
        L0_cnt_inst_N11), .ZN(L0_cnt_inst_n14) );
  NOR2_X1 L0_cnt_inst_U4 ( .A1(s_tc_L0), .A2(1'b0), .ZN(L0_cnt_inst_n13) );
  XOR2_X1 L0_cnt_inst_U20 ( .A(L0_cnt_inst_n9), .B(arv_L0[1]), .Z(
        L0_cnt_inst_n16) );
  NAND3_X1 L0_cnt_inst_U19 ( .A1(int_L0_ptr[1]), .A2(int_L0_ptr[0]), .A3(
        L0_cnt_inst_n13), .ZN(L0_cnt_inst_n12) );
  DFFR_X1 L0_cnt_inst_cnt_out_reg_3_ ( .D(L0_cnt_inst_N14), .CK(
        L0_cnt_inst_net2915), .RN(L0_cnt_inst_n2), .Q(L0_cnt_inst_q_3_), .QN(
        L0_cnt_inst_n5) );
  DFFR_X1 L0_cnt_inst_cnt_out_reg_2_ ( .D(L0_cnt_inst_N13), .CK(
        L0_cnt_inst_net2915), .RN(L0_cnt_inst_n2), .Q(int_L0_ptr[2]), .QN(
        L0_cnt_inst_n8) );
  SDFFR_X1 L0_cnt_inst_cnt_out_reg_1_ ( .D(L0_cnt_inst_n13), .SI(1'b0), .SE(
        L0_cnt_inst_n15), .CK(L0_cnt_inst_net2915), .RN(L0_cnt_inst_n2), .Q(
        int_L0_ptr[1]), .QN(L0_cnt_inst_n9) );
  DFFR_X1 L0_cnt_inst_cnt_out_reg_0_ ( .D(L0_cnt_inst_N11), .CK(
        L0_cnt_inst_net2915), .RN(L0_cnt_inst_n2), .Q(int_L0_ptr[0]), .QN(
        L0_cnt_inst_n1) );
  CLKGATETST_X1 L0_cnt_inst_clk_gate_cnt_out_reg_latch ( .CK(ck), .E(
        ctrl_en_npu), .SE(1'b0), .GCK(L0_cnt_inst_net2915) );
  INV_X1 L4_cnt_inst_U17 ( .A(rst), .ZN(L4_cnt_inst_n2) );
  XNOR2_X1 L4_cnt_inst_U16 ( .A(L4_cnt_inst_q_0_), .B(L4_cnt_inst_q_1_), .ZN(
        L4_cnt_inst_n15) );
  AND2_X1 L4_cnt_inst_U15 ( .A1(L4_cnt_inst_n13), .A2(L4_cnt_inst_n1), .ZN(
        L4_cnt_inst_N11) );
  XNOR2_X1 L4_cnt_inst_U14 ( .A(L4_cnt_inst_q_3_), .B(arv_L4[3]), .ZN(
        L4_cnt_inst_n18) );
  XNOR2_X1 L4_cnt_inst_U13 ( .A(L4_cnt_inst_q_2_), .B(arv_L4[2]), .ZN(
        L4_cnt_inst_n17) );
  AND4_X1 L4_cnt_inst_U12 ( .A1(L4_cnt_inst_n16), .A2(L4_cnt_inst_n17), .A3(
        L4_cnt_inst_n18), .A4(L4_cnt_inst_n19), .ZN(int_d_tc[0]) );
  INV_X1 L4_cnt_inst_U11 ( .A(L4_cnt_inst_n14), .ZN(L4_cnt_inst_n4) );
  AOI21_X1 L4_cnt_inst_U10 ( .B1(L4_cnt_inst_n13), .B2(L4_cnt_inst_n8), .A(
        L4_cnt_inst_n4), .ZN(L4_cnt_inst_n10) );
  OR3_X1 L4_cnt_inst_U9 ( .A1(L4_cnt_inst_n8), .A2(L4_cnt_inst_q_3_), .A3(
        L4_cnt_inst_n12), .ZN(L4_cnt_inst_n11) );
  OAI21_X1 L4_cnt_inst_U8 ( .B1(L4_cnt_inst_n10), .B2(L4_cnt_inst_n5), .A(
        L4_cnt_inst_n11), .ZN(L4_cnt_inst_N14) );
  XNOR2_X1 L4_cnt_inst_U7 ( .A(L4_cnt_inst_q_0_), .B(arv_L4[0]), .ZN(
        L4_cnt_inst_n19) );
  OAI22_X1 L4_cnt_inst_U6 ( .A1(L4_cnt_inst_n14), .A2(L4_cnt_inst_n8), .B1(
        L4_cnt_inst_q_2_), .B2(L4_cnt_inst_n12), .ZN(L4_cnt_inst_N13) );
  AOI21_X1 L4_cnt_inst_U5 ( .B1(L4_cnt_inst_n9), .B2(L4_cnt_inst_n13), .A(
        L4_cnt_inst_N11), .ZN(L4_cnt_inst_n14) );
  NOR2_X1 L4_cnt_inst_U4 ( .A1(int_d_tc[0]), .A2(1'b0), .ZN(L4_cnt_inst_n13)
         );
  XOR2_X1 L4_cnt_inst_U20 ( .A(L4_cnt_inst_n9), .B(arv_L4[1]), .Z(
        L4_cnt_inst_n16) );
  NAND3_X1 L4_cnt_inst_U19 ( .A1(L4_cnt_inst_q_1_), .A2(L4_cnt_inst_q_0_), 
        .A3(L4_cnt_inst_n13), .ZN(L4_cnt_inst_n12) );
  DFFR_X1 L4_cnt_inst_cnt_out_reg_3_ ( .D(L4_cnt_inst_N14), .CK(
        L4_cnt_inst_net2897), .RN(L4_cnt_inst_n2), .Q(L4_cnt_inst_q_3_), .QN(
        L4_cnt_inst_n5) );
  DFFR_X1 L4_cnt_inst_cnt_out_reg_2_ ( .D(L4_cnt_inst_N13), .CK(
        L4_cnt_inst_net2897), .RN(L4_cnt_inst_n2), .Q(L4_cnt_inst_q_2_), .QN(
        L4_cnt_inst_n8) );
  SDFFR_X1 L4_cnt_inst_cnt_out_reg_1_ ( .D(L4_cnt_inst_n13), .SI(1'b0), .SE(
        L4_cnt_inst_n15), .CK(L4_cnt_inst_net2897), .RN(L4_cnt_inst_n2), .Q(
        L4_cnt_inst_q_1_), .QN(L4_cnt_inst_n9) );
  DFFR_X1 L4_cnt_inst_cnt_out_reg_0_ ( .D(L4_cnt_inst_N11), .CK(
        L4_cnt_inst_net2897), .RN(L4_cnt_inst_n2), .Q(L4_cnt_inst_q_0_), .QN(
        L4_cnt_inst_n1) );
  CLKGATETST_X1 L4_cnt_inst_clk_gate_cnt_out_reg_latch ( .CK(ck), .E(
        int_en_L4_ptr), .SE(1'b0), .GCK(L4_cnt_inst_net2897) );
  INV_X1 i_weight_addr_gen_inst_U41 ( .A(rst), .ZN(i_weight_addr_gen_inst_n6)
         );
  INV_X1 i_weight_addr_gen_inst_U40 ( .A(rst), .ZN(i_weight_addr_gen_inst_n5)
         );
  OR2_X1 i_weight_addr_gen_inst_U39 ( .A1(ctrl_en_hmode), .A2(s_tc_res), .ZN(
        i_weight_addr_gen_inst_N60) );
  OR2_X1 i_weight_addr_gen_inst_U38 ( .A1(int_c_i_en_weight_addr), .A2(1'b0), 
        .ZN(i_weight_addr_gen_inst_N37) );
  AOI22_X1 i_weight_addr_gen_inst_U37 ( .A1(i_weight_addr_gen_inst_N27), .A2(
        i_weight_addr_gen_inst_n31), .B1(i_weight_addr_gen_inst_N18), .B2(
        i_weight_addr_gen_inst_n32), .ZN(i_weight_addr_gen_inst_n30) );
  INV_X1 i_weight_addr_gen_inst_U36 ( .A(i_weight_addr_gen_inst_n30), .ZN(
        i_weight_addr_gen_inst_n7) );
  INV_X1 i_weight_addr_gen_inst_U35 ( .A(int_c_i_en_weight_addr), .ZN(
        i_weight_addr_gen_inst_n26) );
  INV_X1 i_weight_addr_gen_inst_U34 ( .A(s_tc_res), .ZN(
        i_weight_addr_gen_inst_n25) );
  AOI22_X1 i_weight_addr_gen_inst_U33 ( .A1(i_weight_addr_gen_inst_N19), .A2(
        i_weight_addr_gen_inst_n31), .B1(i_weight_addr_gen_inst_N10), .B2(
        i_weight_addr_gen_inst_n32), .ZN(i_weight_addr_gen_inst_n40) );
  INV_X1 i_weight_addr_gen_inst_U32 ( .A(i_weight_addr_gen_inst_n40), .ZN(
        i_weight_addr_gen_inst_n24) );
  AOI22_X1 i_weight_addr_gen_inst_U31 ( .A1(i_weight_addr_gen_inst_N20), .A2(
        i_weight_addr_gen_inst_n31), .B1(i_weight_addr_gen_inst_N11), .B2(
        i_weight_addr_gen_inst_n32), .ZN(i_weight_addr_gen_inst_n39) );
  INV_X1 i_weight_addr_gen_inst_U30 ( .A(i_weight_addr_gen_inst_n39), .ZN(
        i_weight_addr_gen_inst_n23) );
  AOI22_X1 i_weight_addr_gen_inst_U29 ( .A1(i_weight_addr_gen_inst_N21), .A2(
        i_weight_addr_gen_inst_n31), .B1(i_weight_addr_gen_inst_N12), .B2(
        i_weight_addr_gen_inst_n32), .ZN(i_weight_addr_gen_inst_n38) );
  INV_X1 i_weight_addr_gen_inst_U28 ( .A(i_weight_addr_gen_inst_n38), .ZN(
        i_weight_addr_gen_inst_n22) );
  AOI22_X1 i_weight_addr_gen_inst_U27 ( .A1(i_weight_addr_gen_inst_N22), .A2(
        i_weight_addr_gen_inst_n31), .B1(i_weight_addr_gen_inst_N13), .B2(
        i_weight_addr_gen_inst_n32), .ZN(i_weight_addr_gen_inst_n37) );
  INV_X1 i_weight_addr_gen_inst_U26 ( .A(i_weight_addr_gen_inst_n37), .ZN(
        i_weight_addr_gen_inst_n21) );
  AOI22_X1 i_weight_addr_gen_inst_U25 ( .A1(i_weight_addr_gen_inst_N23), .A2(
        i_weight_addr_gen_inst_n31), .B1(i_weight_addr_gen_inst_N14), .B2(
        i_weight_addr_gen_inst_n32), .ZN(i_weight_addr_gen_inst_n36) );
  INV_X1 i_weight_addr_gen_inst_U24 ( .A(i_weight_addr_gen_inst_n36), .ZN(
        i_weight_addr_gen_inst_n20) );
  AOI22_X1 i_weight_addr_gen_inst_U23 ( .A1(i_weight_addr_gen_inst_N24), .A2(
        i_weight_addr_gen_inst_n31), .B1(i_weight_addr_gen_inst_N15), .B2(
        i_weight_addr_gen_inst_n32), .ZN(i_weight_addr_gen_inst_n35) );
  INV_X1 i_weight_addr_gen_inst_U22 ( .A(i_weight_addr_gen_inst_n35), .ZN(
        i_weight_addr_gen_inst_n19) );
  AOI22_X1 i_weight_addr_gen_inst_U21 ( .A1(i_weight_addr_gen_inst_N25), .A2(
        i_weight_addr_gen_inst_n31), .B1(i_weight_addr_gen_inst_N16), .B2(
        i_weight_addr_gen_inst_n32), .ZN(i_weight_addr_gen_inst_n34) );
  INV_X1 i_weight_addr_gen_inst_U20 ( .A(i_weight_addr_gen_inst_n34), .ZN(
        i_weight_addr_gen_inst_n17) );
  AOI22_X1 i_weight_addr_gen_inst_U19 ( .A1(i_weight_addr_gen_inst_N26), .A2(
        i_weight_addr_gen_inst_n31), .B1(i_weight_addr_gen_inst_N17), .B2(
        i_weight_addr_gen_inst_n32), .ZN(i_weight_addr_gen_inst_n33) );
  INV_X1 i_weight_addr_gen_inst_U18 ( .A(i_weight_addr_gen_inst_n33), .ZN(
        i_weight_addr_gen_inst_n8) );
  NOR2_X1 i_weight_addr_gen_inst_U17 ( .A1(i_weight_addr_gen_inst_n26), .A2(
        1'b0), .ZN(i_weight_addr_gen_inst_n32) );
  NOR2_X1 i_weight_addr_gen_inst_U15 ( .A1(int_c_i_en_weight_addr), .A2(1'b0), 
        .ZN(i_weight_addr_gen_inst_n31) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_7_ ( .D(
        i_weight_addr_gen_inst_n8), .CK(i_weight_addr_gen_inst_net2874), .RN(
        i_weight_addr_gen_inst_n5), .Q(i_weight_addr_gen_inst_int_base_addr_7_) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_6_ ( .D(
        i_weight_addr_gen_inst_n17), .CK(i_weight_addr_gen_inst_net2874), .RN(
        i_weight_addr_gen_inst_n5), .Q(i_weight_addr_gen_inst_int_base_addr_6_) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_5_ ( .D(
        i_weight_addr_gen_inst_n19), .CK(i_weight_addr_gen_inst_net2874), .RN(
        i_weight_addr_gen_inst_n5), .Q(i_weight_addr_gen_inst_int_base_addr_5_) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_4_ ( .D(
        i_weight_addr_gen_inst_n20), .CK(i_weight_addr_gen_inst_net2874), .RN(
        i_weight_addr_gen_inst_n5), .Q(i_weight_addr_gen_inst_int_base_addr_4_) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_3_ ( .D(
        i_weight_addr_gen_inst_n21), .CK(i_weight_addr_gen_inst_net2874), .RN(
        i_weight_addr_gen_inst_n5), .Q(i_weight_addr_gen_inst_int_base_addr_3_) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_2_ ( .D(
        i_weight_addr_gen_inst_n22), .CK(i_weight_addr_gen_inst_net2874), .RN(
        i_weight_addr_gen_inst_n5), .Q(i_weight_addr_gen_inst_int_base_addr_2_) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_1_ ( .D(
        i_weight_addr_gen_inst_n23), .CK(i_weight_addr_gen_inst_net2874), .RN(
        i_weight_addr_gen_inst_n5), .Q(i_weight_addr_gen_inst_int_base_addr_1_) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_0_ ( .D(
        i_weight_addr_gen_inst_n24), .CK(i_weight_addr_gen_inst_net2874), .RN(
        i_weight_addr_gen_inst_n5), .Q(i_weight_addr_gen_inst_int_base_addr_0_) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_8_ ( .D(
        i_weight_addr_gen_inst_n7), .CK(i_weight_addr_gen_inst_net2874), .RN(
        i_weight_addr_gen_inst_n5), .Q(i_weight_addr_gen_inst_int_base_addr_8_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_8_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n25), .SE(i_weight_addr_gen_inst_N59), .CK(
        i_weight_addr_gen_inst_net2880), .RN(i_weight_addr_gen_inst_n5), .Q(
        i_weight_addr_gen_inst_int_offs_addr_8_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_7_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n25), .SE(i_weight_addr_gen_inst_N58), .CK(
        i_weight_addr_gen_inst_net2880), .RN(i_weight_addr_gen_inst_n5), .Q(
        i_weight_addr_gen_inst_int_offs_addr_7_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_6_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n25), .SE(i_weight_addr_gen_inst_N57), .CK(
        i_weight_addr_gen_inst_net2880), .RN(i_weight_addr_gen_inst_n5), .Q(
        i_weight_addr_gen_inst_int_offs_addr_6_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_5_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n25), .SE(i_weight_addr_gen_inst_N56), .CK(
        i_weight_addr_gen_inst_net2880), .RN(i_weight_addr_gen_inst_n6), .Q(
        i_weight_addr_gen_inst_int_offs_addr_5_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_4_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n25), .SE(i_weight_addr_gen_inst_N55), .CK(
        i_weight_addr_gen_inst_net2880), .RN(i_weight_addr_gen_inst_n6), .Q(
        i_weight_addr_gen_inst_int_offs_addr_4_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_3_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n25), .SE(i_weight_addr_gen_inst_N54), .CK(
        i_weight_addr_gen_inst_net2880), .RN(i_weight_addr_gen_inst_n6), .Q(
        i_weight_addr_gen_inst_int_offs_addr_3_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_2_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n25), .SE(i_weight_addr_gen_inst_N53), .CK(
        i_weight_addr_gen_inst_net2880), .RN(i_weight_addr_gen_inst_n6), .Q(
        i_weight_addr_gen_inst_int_offs_addr_2_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_1_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n25), .SE(i_weight_addr_gen_inst_N52), .CK(
        i_weight_addr_gen_inst_net2880), .RN(i_weight_addr_gen_inst_n6), .Q(
        i_weight_addr_gen_inst_int_offs_addr_1_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_0_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n25), .SE(i_weight_addr_gen_inst_N51), .CK(
        i_weight_addr_gen_inst_net2880), .RN(i_weight_addr_gen_inst_n6), .Q(
        i_weight_addr_gen_inst_int_offs_addr_0_) );
  CLKGATETST_X1 i_weight_addr_gen_inst_clk_gate_int_base_addr_reg_latch ( .CK(
        ck), .E(i_weight_addr_gen_inst_N37), .SE(1'b0), .GCK(
        i_weight_addr_gen_inst_net2874) );
  CLKGATETST_X1 i_weight_addr_gen_inst_clk_gate_int_offs_addr_reg_latch ( .CK(
        ck), .E(i_weight_addr_gen_inst_N60), .SE(1'b0), .GCK(
        i_weight_addr_gen_inst_net2880) );
  XOR2_X1 i_weight_addr_gen_inst_add_60_U2 ( .A(1'b1), .B(
        i_weight_addr_gen_inst_int_offs_addr_0_), .Z(
        i_weight_addr_gen_inst_N51) );
  AND2_X1 i_weight_addr_gen_inst_add_60_U1 ( .A1(1'b1), .A2(
        i_weight_addr_gen_inst_int_offs_addr_0_), .ZN(
        i_weight_addr_gen_inst_add_60_n1) );
  FA_X1 i_weight_addr_gen_inst_add_60_U1_1 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_1_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_60_n1), .CO(
        i_weight_addr_gen_inst_add_60_carry[2]), .S(i_weight_addr_gen_inst_N52) );
  FA_X1 i_weight_addr_gen_inst_add_60_U1_2 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_2_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_60_carry[2]), .CO(
        i_weight_addr_gen_inst_add_60_carry[3]), .S(i_weight_addr_gen_inst_N53) );
  FA_X1 i_weight_addr_gen_inst_add_60_U1_3 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_3_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_60_carry[3]), .CO(
        i_weight_addr_gen_inst_add_60_carry[4]), .S(i_weight_addr_gen_inst_N54) );
  FA_X1 i_weight_addr_gen_inst_add_60_U1_4 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_4_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_60_carry[4]), .CO(
        i_weight_addr_gen_inst_add_60_carry[5]), .S(i_weight_addr_gen_inst_N55) );
  FA_X1 i_weight_addr_gen_inst_add_60_U1_5 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_5_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_60_carry[5]), .CO(
        i_weight_addr_gen_inst_add_60_carry[6]), .S(i_weight_addr_gen_inst_N56) );
  FA_X1 i_weight_addr_gen_inst_add_60_U1_6 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_6_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_60_carry[6]), .CO(
        i_weight_addr_gen_inst_add_60_carry[7]), .S(i_weight_addr_gen_inst_N57) );
  FA_X1 i_weight_addr_gen_inst_add_60_U1_7 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_7_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_60_carry[7]), .CO(
        i_weight_addr_gen_inst_add_60_carry[8]), .S(i_weight_addr_gen_inst_N58) );
  FA_X1 i_weight_addr_gen_inst_add_60_U1_8 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_8_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_60_carry[8]), .S(i_weight_addr_gen_inst_N59) );
  AND2_X1 i_weight_addr_gen_inst_add_45_U2 ( .A1(1'b0), .A2(
        i_weight_addr_gen_inst_int_base_addr_0_), .ZN(
        i_weight_addr_gen_inst_add_45_n2) );
  XOR2_X1 i_weight_addr_gen_inst_add_45_U1 ( .A(1'b0), .B(
        i_weight_addr_gen_inst_int_base_addr_0_), .Z(
        i_weight_addr_gen_inst_N19) );
  FA_X1 i_weight_addr_gen_inst_add_45_U1_1 ( .A(
        i_weight_addr_gen_inst_int_base_addr_1_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_45_n2), .CO(
        i_weight_addr_gen_inst_add_45_carry[2]), .S(i_weight_addr_gen_inst_N20) );
  FA_X1 i_weight_addr_gen_inst_add_45_U1_2 ( .A(
        i_weight_addr_gen_inst_int_base_addr_2_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_45_carry[2]), .CO(
        i_weight_addr_gen_inst_add_45_carry[3]), .S(i_weight_addr_gen_inst_N21) );
  FA_X1 i_weight_addr_gen_inst_add_45_U1_3 ( .A(
        i_weight_addr_gen_inst_int_base_addr_3_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_45_carry[3]), .CO(
        i_weight_addr_gen_inst_add_45_carry[4]), .S(i_weight_addr_gen_inst_N22) );
  FA_X1 i_weight_addr_gen_inst_add_45_U1_4 ( .A(
        i_weight_addr_gen_inst_int_base_addr_4_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_45_carry[4]), .CO(
        i_weight_addr_gen_inst_add_45_carry[5]), .S(i_weight_addr_gen_inst_N23) );
  FA_X1 i_weight_addr_gen_inst_add_45_U1_5 ( .A(
        i_weight_addr_gen_inst_int_base_addr_5_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_45_carry[5]), .CO(
        i_weight_addr_gen_inst_add_45_carry[6]), .S(i_weight_addr_gen_inst_N24) );
  FA_X1 i_weight_addr_gen_inst_add_45_U1_6 ( .A(
        i_weight_addr_gen_inst_int_base_addr_6_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_45_carry[6]), .CO(
        i_weight_addr_gen_inst_add_45_carry[7]), .S(i_weight_addr_gen_inst_N25) );
  FA_X1 i_weight_addr_gen_inst_add_45_U1_7 ( .A(
        i_weight_addr_gen_inst_int_base_addr_7_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_45_carry[7]), .CO(
        i_weight_addr_gen_inst_add_45_carry[8]), .S(i_weight_addr_gen_inst_N26) );
  FA_X1 i_weight_addr_gen_inst_add_45_U1_8 ( .A(
        i_weight_addr_gen_inst_int_base_addr_8_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_45_carry[8]), .S(i_weight_addr_gen_inst_N27) );
  AND2_X1 i_weight_addr_gen_inst_add_43_U2 ( .A1(1'b0), .A2(i_weight_addr[0]), 
        .ZN(i_weight_addr_gen_inst_add_43_n2) );
  XOR2_X1 i_weight_addr_gen_inst_add_43_U1 ( .A(1'b0), .B(i_weight_addr[0]), 
        .Z(i_weight_addr_gen_inst_N10) );
  FA_X1 i_weight_addr_gen_inst_add_43_U1_1 ( .A(i_weight_addr[1]), .B(1'b0), 
        .CI(i_weight_addr_gen_inst_add_43_n2), .CO(
        i_weight_addr_gen_inst_add_43_carry[2]), .S(i_weight_addr_gen_inst_N11) );
  FA_X1 i_weight_addr_gen_inst_add_43_U1_2 ( .A(i_weight_addr[2]), .B(1'b0), 
        .CI(i_weight_addr_gen_inst_add_43_carry[2]), .CO(
        i_weight_addr_gen_inst_add_43_carry[3]), .S(i_weight_addr_gen_inst_N12) );
  FA_X1 i_weight_addr_gen_inst_add_43_U1_3 ( .A(i_weight_addr[3]), .B(1'b0), 
        .CI(i_weight_addr_gen_inst_add_43_carry[3]), .CO(
        i_weight_addr_gen_inst_add_43_carry[4]), .S(i_weight_addr_gen_inst_N13) );
  FA_X1 i_weight_addr_gen_inst_add_43_U1_4 ( .A(i_weight_addr[4]), .B(1'b0), 
        .CI(i_weight_addr_gen_inst_add_43_carry[4]), .CO(
        i_weight_addr_gen_inst_add_43_carry[5]), .S(i_weight_addr_gen_inst_N14) );
  FA_X1 i_weight_addr_gen_inst_add_43_U1_5 ( .A(i_weight_addr[5]), .B(1'b0), 
        .CI(i_weight_addr_gen_inst_add_43_carry[5]), .CO(
        i_weight_addr_gen_inst_add_43_carry[6]), .S(i_weight_addr_gen_inst_N15) );
  FA_X1 i_weight_addr_gen_inst_add_43_U1_6 ( .A(i_weight_addr[6]), .B(1'b0), 
        .CI(i_weight_addr_gen_inst_add_43_carry[6]), .CO(
        i_weight_addr_gen_inst_add_43_carry[7]), .S(i_weight_addr_gen_inst_N16) );
  FA_X1 i_weight_addr_gen_inst_add_43_U1_7 ( .A(i_weight_addr[7]), .B(1'b0), 
        .CI(i_weight_addr_gen_inst_add_43_carry[7]), .CO(
        i_weight_addr_gen_inst_add_43_carry[8]), .S(i_weight_addr_gen_inst_N17) );
  FA_X1 i_weight_addr_gen_inst_add_43_U1_8 ( .A(i_weight_addr[8]), .B(1'b0), 
        .CI(i_weight_addr_gen_inst_add_43_carry[8]), .S(
        i_weight_addr_gen_inst_N18) );
  XOR2_X1 i_weight_addr_gen_inst_add_31_U2 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_0_), .B(
        i_weight_addr_gen_inst_int_base_addr_0_), .Z(i_weight_addr[0]) );
  AND2_X1 i_weight_addr_gen_inst_add_31_U1 ( .A1(
        i_weight_addr_gen_inst_int_offs_addr_0_), .A2(
        i_weight_addr_gen_inst_int_base_addr_0_), .ZN(
        i_weight_addr_gen_inst_add_31_n1) );
  FA_X1 i_weight_addr_gen_inst_add_31_U1_1 ( .A(
        i_weight_addr_gen_inst_int_base_addr_1_), .B(
        i_weight_addr_gen_inst_int_offs_addr_1_), .CI(
        i_weight_addr_gen_inst_add_31_n1), .CO(
        i_weight_addr_gen_inst_add_31_carry[2]), .S(i_weight_addr[1]) );
  FA_X1 i_weight_addr_gen_inst_add_31_U1_2 ( .A(
        i_weight_addr_gen_inst_int_base_addr_2_), .B(
        i_weight_addr_gen_inst_int_offs_addr_2_), .CI(
        i_weight_addr_gen_inst_add_31_carry[2]), .CO(
        i_weight_addr_gen_inst_add_31_carry[3]), .S(i_weight_addr[2]) );
  FA_X1 i_weight_addr_gen_inst_add_31_U1_3 ( .A(
        i_weight_addr_gen_inst_int_base_addr_3_), .B(
        i_weight_addr_gen_inst_int_offs_addr_3_), .CI(
        i_weight_addr_gen_inst_add_31_carry[3]), .CO(
        i_weight_addr_gen_inst_add_31_carry[4]), .S(i_weight_addr[3]) );
  FA_X1 i_weight_addr_gen_inst_add_31_U1_4 ( .A(
        i_weight_addr_gen_inst_int_base_addr_4_), .B(
        i_weight_addr_gen_inst_int_offs_addr_4_), .CI(
        i_weight_addr_gen_inst_add_31_carry[4]), .CO(
        i_weight_addr_gen_inst_add_31_carry[5]), .S(i_weight_addr[4]) );
  FA_X1 i_weight_addr_gen_inst_add_31_U1_5 ( .A(
        i_weight_addr_gen_inst_int_base_addr_5_), .B(
        i_weight_addr_gen_inst_int_offs_addr_5_), .CI(
        i_weight_addr_gen_inst_add_31_carry[5]), .CO(
        i_weight_addr_gen_inst_add_31_carry[6]), .S(i_weight_addr[5]) );
  FA_X1 i_weight_addr_gen_inst_add_31_U1_6 ( .A(
        i_weight_addr_gen_inst_int_base_addr_6_), .B(
        i_weight_addr_gen_inst_int_offs_addr_6_), .CI(
        i_weight_addr_gen_inst_add_31_carry[6]), .CO(
        i_weight_addr_gen_inst_add_31_carry[7]), .S(i_weight_addr[6]) );
  FA_X1 i_weight_addr_gen_inst_add_31_U1_7 ( .A(
        i_weight_addr_gen_inst_int_base_addr_7_), .B(
        i_weight_addr_gen_inst_int_offs_addr_7_), .CI(
        i_weight_addr_gen_inst_add_31_carry[7]), .CO(
        i_weight_addr_gen_inst_add_31_carry[8]), .S(i_weight_addr[7]) );
  FA_X1 i_weight_addr_gen_inst_add_31_U1_8 ( .A(
        i_weight_addr_gen_inst_int_base_addr_8_), .B(
        i_weight_addr_gen_inst_int_offs_addr_8_), .CI(
        i_weight_addr_gen_inst_add_31_carry[8]), .S(i_weight_addr[8]) );
  INV_X1 i_data_even_addr_gen_inst_U44 ( .A(rst), .ZN(
        i_data_even_addr_gen_inst_n6) );
  INV_X1 i_data_even_addr_gen_inst_U43 ( .A(rst), .ZN(
        i_data_even_addr_gen_inst_n5) );
  AOI22_X1 i_data_even_addr_gen_inst_U42 ( .A1(i_data_even_addr_gen_inst_N29), 
        .A2(i_data_even_addr_gen_inst_n33), .B1(i_data_even_addr_gen_inst_N19), 
        .B2(i_data_even_addr_gen_inst_n34), .ZN(i_data_even_addr_gen_inst_n32)
         );
  INV_X1 i_data_even_addr_gen_inst_U41 ( .A(i_data_even_addr_gen_inst_n32), 
        .ZN(i_data_even_addr_gen_inst_n7) );
  OR2_X1 i_data_even_addr_gen_inst_U40 ( .A1(n33), .A2(ctrl_ldh_v_n), .ZN(
        i_data_even_addr_gen_inst_N65) );
  AOI22_X1 i_data_even_addr_gen_inst_U39 ( .A1(i_data_even_addr_gen_inst_N20), 
        .A2(i_data_even_addr_gen_inst_n33), .B1(i_data_even_addr_gen_inst_N10), 
        .B2(i_data_even_addr_gen_inst_n34), .ZN(i_data_even_addr_gen_inst_n43)
         );
  INV_X1 i_data_even_addr_gen_inst_U38 ( .A(i_data_even_addr_gen_inst_n43), 
        .ZN(i_data_even_addr_gen_inst_n26) );
  AOI22_X1 i_data_even_addr_gen_inst_U37 ( .A1(i_data_even_addr_gen_inst_N21), 
        .A2(i_data_even_addr_gen_inst_n33), .B1(i_data_even_addr_gen_inst_N11), 
        .B2(i_data_even_addr_gen_inst_n34), .ZN(i_data_even_addr_gen_inst_n42)
         );
  INV_X1 i_data_even_addr_gen_inst_U36 ( .A(i_data_even_addr_gen_inst_n42), 
        .ZN(i_data_even_addr_gen_inst_n25) );
  AOI22_X1 i_data_even_addr_gen_inst_U35 ( .A1(i_data_even_addr_gen_inst_N22), 
        .A2(i_data_even_addr_gen_inst_n33), .B1(i_data_even_addr_gen_inst_N12), 
        .B2(i_data_even_addr_gen_inst_n34), .ZN(i_data_even_addr_gen_inst_n41)
         );
  INV_X1 i_data_even_addr_gen_inst_U34 ( .A(i_data_even_addr_gen_inst_n41), 
        .ZN(i_data_even_addr_gen_inst_n24) );
  AOI22_X1 i_data_even_addr_gen_inst_U33 ( .A1(i_data_even_addr_gen_inst_N23), 
        .A2(i_data_even_addr_gen_inst_n33), .B1(i_data_even_addr_gen_inst_N13), 
        .B2(i_data_even_addr_gen_inst_n34), .ZN(i_data_even_addr_gen_inst_n40)
         );
  INV_X1 i_data_even_addr_gen_inst_U32 ( .A(i_data_even_addr_gen_inst_n40), 
        .ZN(i_data_even_addr_gen_inst_n23) );
  AOI22_X1 i_data_even_addr_gen_inst_U31 ( .A1(i_data_even_addr_gen_inst_N24), 
        .A2(i_data_even_addr_gen_inst_n33), .B1(i_data_even_addr_gen_inst_N14), 
        .B2(i_data_even_addr_gen_inst_n34), .ZN(i_data_even_addr_gen_inst_n39)
         );
  INV_X1 i_data_even_addr_gen_inst_U30 ( .A(i_data_even_addr_gen_inst_n39), 
        .ZN(i_data_even_addr_gen_inst_n22) );
  AOI22_X1 i_data_even_addr_gen_inst_U29 ( .A1(i_data_even_addr_gen_inst_N25), 
        .A2(i_data_even_addr_gen_inst_n33), .B1(i_data_even_addr_gen_inst_N15), 
        .B2(i_data_even_addr_gen_inst_n34), .ZN(i_data_even_addr_gen_inst_n38)
         );
  INV_X1 i_data_even_addr_gen_inst_U28 ( .A(i_data_even_addr_gen_inst_n38), 
        .ZN(i_data_even_addr_gen_inst_n21) );
  AOI22_X1 i_data_even_addr_gen_inst_U27 ( .A1(i_data_even_addr_gen_inst_N26), 
        .A2(i_data_even_addr_gen_inst_n33), .B1(i_data_even_addr_gen_inst_N16), 
        .B2(i_data_even_addr_gen_inst_n34), .ZN(i_data_even_addr_gen_inst_n37)
         );
  INV_X1 i_data_even_addr_gen_inst_U26 ( .A(i_data_even_addr_gen_inst_n37), 
        .ZN(i_data_even_addr_gen_inst_n20) );
  AOI22_X1 i_data_even_addr_gen_inst_U25 ( .A1(i_data_even_addr_gen_inst_N27), 
        .A2(i_data_even_addr_gen_inst_n33), .B1(i_data_even_addr_gen_inst_N17), 
        .B2(i_data_even_addr_gen_inst_n34), .ZN(i_data_even_addr_gen_inst_n36)
         );
  INV_X1 i_data_even_addr_gen_inst_U24 ( .A(i_data_even_addr_gen_inst_n36), 
        .ZN(i_data_even_addr_gen_inst_n18) );
  AOI22_X1 i_data_even_addr_gen_inst_U23 ( .A1(i_data_even_addr_gen_inst_N28), 
        .A2(i_data_even_addr_gen_inst_n33), .B1(i_data_even_addr_gen_inst_N18), 
        .B2(i_data_even_addr_gen_inst_n34), .ZN(i_data_even_addr_gen_inst_n35)
         );
  INV_X1 i_data_even_addr_gen_inst_U22 ( .A(i_data_even_addr_gen_inst_n35), 
        .ZN(i_data_even_addr_gen_inst_n8) );
  OR2_X1 i_data_even_addr_gen_inst_U21 ( .A1(int_c_i_en_even), .A2(
        int_en_L4_ptr), .ZN(i_data_even_addr_gen_inst_N40) );
  INV_X1 i_data_even_addr_gen_inst_U20 ( .A(int_c_i_en_even), .ZN(
        i_data_even_addr_gen_inst_n28) );
  NOR2_X1 i_data_even_addr_gen_inst_U19 ( .A1(i_data_even_addr_gen_inst_n28), 
        .A2(int_en_L4_ptr), .ZN(i_data_even_addr_gen_inst_n34) );
  NOR2_X1 i_data_even_addr_gen_inst_U18 ( .A1(int_c_i_en_even), .A2(
        int_en_L4_ptr), .ZN(i_data_even_addr_gen_inst_n33) );
  INV_X1 i_data_even_addr_gen_inst_U16 ( .A(n33), .ZN(
        i_data_even_addr_gen_inst_n27) );
  DFFR_X1 i_data_even_addr_gen_inst_int_base_addr_reg_8_ ( .D(
        i_data_even_addr_gen_inst_n8), .CK(i_data_even_addr_gen_inst_net2851), 
        .RN(i_data_even_addr_gen_inst_n5), .Q(
        i_data_even_addr_gen_inst_int_base_addr_8_) );
  DFFR_X1 i_data_even_addr_gen_inst_int_base_addr_reg_7_ ( .D(
        i_data_even_addr_gen_inst_n18), .CK(i_data_even_addr_gen_inst_net2851), 
        .RN(i_data_even_addr_gen_inst_n5), .Q(
        i_data_even_addr_gen_inst_int_base_addr_7_) );
  DFFR_X1 i_data_even_addr_gen_inst_int_base_addr_reg_6_ ( .D(
        i_data_even_addr_gen_inst_n20), .CK(i_data_even_addr_gen_inst_net2851), 
        .RN(i_data_even_addr_gen_inst_n5), .Q(
        i_data_even_addr_gen_inst_int_base_addr_6_) );
  DFFR_X1 i_data_even_addr_gen_inst_int_base_addr_reg_5_ ( .D(
        i_data_even_addr_gen_inst_n21), .CK(i_data_even_addr_gen_inst_net2851), 
        .RN(i_data_even_addr_gen_inst_n5), .Q(
        i_data_even_addr_gen_inst_int_base_addr_5_) );
  DFFR_X1 i_data_even_addr_gen_inst_int_base_addr_reg_4_ ( .D(
        i_data_even_addr_gen_inst_n22), .CK(i_data_even_addr_gen_inst_net2851), 
        .RN(i_data_even_addr_gen_inst_n5), .Q(
        i_data_even_addr_gen_inst_int_base_addr_4_) );
  DFFR_X1 i_data_even_addr_gen_inst_int_base_addr_reg_3_ ( .D(
        i_data_even_addr_gen_inst_n23), .CK(i_data_even_addr_gen_inst_net2851), 
        .RN(i_data_even_addr_gen_inst_n5), .Q(
        i_data_even_addr_gen_inst_int_base_addr_3_) );
  DFFR_X1 i_data_even_addr_gen_inst_int_base_addr_reg_2_ ( .D(
        i_data_even_addr_gen_inst_n24), .CK(i_data_even_addr_gen_inst_net2851), 
        .RN(i_data_even_addr_gen_inst_n5), .Q(
        i_data_even_addr_gen_inst_int_base_addr_2_) );
  DFFR_X1 i_data_even_addr_gen_inst_int_base_addr_reg_1_ ( .D(
        i_data_even_addr_gen_inst_n25), .CK(i_data_even_addr_gen_inst_net2851), 
        .RN(i_data_even_addr_gen_inst_n5), .Q(
        i_data_even_addr_gen_inst_int_base_addr_1_) );
  DFFR_X1 i_data_even_addr_gen_inst_int_base_addr_reg_0_ ( .D(
        i_data_even_addr_gen_inst_n26), .CK(i_data_even_addr_gen_inst_net2851), 
        .RN(i_data_even_addr_gen_inst_n5), .Q(
        i_data_even_addr_gen_inst_int_base_addr_0_) );
  DFFR_X1 i_data_even_addr_gen_inst_int_base_addr_reg_9_ ( .D(
        i_data_even_addr_gen_inst_n7), .CK(i_data_even_addr_gen_inst_net2851), 
        .RN(i_data_even_addr_gen_inst_n5), .Q(
        i_data_even_addr_gen_inst_int_base_addr_9_) );
  SDFFR_X1 i_data_even_addr_gen_inst_int_offs_addr_reg_9_ ( .D(1'b0), .SI(
        i_data_even_addr_gen_inst_n27), .SE(i_data_even_addr_gen_inst_N64), 
        .CK(i_data_even_addr_gen_inst_net2857), .RN(
        i_data_even_addr_gen_inst_n5), .Q(
        i_data_even_addr_gen_inst_int_offs_addr_9_) );
  SDFFR_X1 i_data_even_addr_gen_inst_int_offs_addr_reg_8_ ( .D(1'b0), .SI(
        i_data_even_addr_gen_inst_n27), .SE(i_data_even_addr_gen_inst_N63), 
        .CK(i_data_even_addr_gen_inst_net2857), .RN(
        i_data_even_addr_gen_inst_n5), .Q(
        i_data_even_addr_gen_inst_int_offs_addr_8_) );
  SDFFR_X1 i_data_even_addr_gen_inst_int_offs_addr_reg_7_ ( .D(1'b0), .SI(
        i_data_even_addr_gen_inst_n27), .SE(i_data_even_addr_gen_inst_N62), 
        .CK(i_data_even_addr_gen_inst_net2857), .RN(
        i_data_even_addr_gen_inst_n6), .Q(
        i_data_even_addr_gen_inst_int_offs_addr_7_) );
  SDFFR_X1 i_data_even_addr_gen_inst_int_offs_addr_reg_6_ ( .D(1'b0), .SI(
        i_data_even_addr_gen_inst_n27), .SE(i_data_even_addr_gen_inst_N61), 
        .CK(i_data_even_addr_gen_inst_net2857), .RN(
        i_data_even_addr_gen_inst_n6), .Q(
        i_data_even_addr_gen_inst_int_offs_addr_6_) );
  SDFFR_X1 i_data_even_addr_gen_inst_int_offs_addr_reg_5_ ( .D(1'b0), .SI(
        i_data_even_addr_gen_inst_n27), .SE(i_data_even_addr_gen_inst_N60), 
        .CK(i_data_even_addr_gen_inst_net2857), .RN(
        i_data_even_addr_gen_inst_n6), .Q(
        i_data_even_addr_gen_inst_int_offs_addr_5_) );
  SDFFR_X1 i_data_even_addr_gen_inst_int_offs_addr_reg_4_ ( .D(1'b0), .SI(
        i_data_even_addr_gen_inst_n27), .SE(i_data_even_addr_gen_inst_N59), 
        .CK(i_data_even_addr_gen_inst_net2857), .RN(
        i_data_even_addr_gen_inst_n6), .Q(
        i_data_even_addr_gen_inst_int_offs_addr_4_) );
  SDFFR_X1 i_data_even_addr_gen_inst_int_offs_addr_reg_3_ ( .D(1'b0), .SI(
        i_data_even_addr_gen_inst_n27), .SE(i_data_even_addr_gen_inst_N58), 
        .CK(i_data_even_addr_gen_inst_net2857), .RN(
        i_data_even_addr_gen_inst_n6), .Q(
        i_data_even_addr_gen_inst_int_offs_addr_3_) );
  SDFFR_X1 i_data_even_addr_gen_inst_int_offs_addr_reg_2_ ( .D(1'b0), .SI(
        i_data_even_addr_gen_inst_n27), .SE(i_data_even_addr_gen_inst_N57), 
        .CK(i_data_even_addr_gen_inst_net2857), .RN(
        i_data_even_addr_gen_inst_n6), .Q(
        i_data_even_addr_gen_inst_int_offs_addr_2_) );
  SDFFR_X1 i_data_even_addr_gen_inst_int_offs_addr_reg_1_ ( .D(1'b0), .SI(
        i_data_even_addr_gen_inst_n27), .SE(i_data_even_addr_gen_inst_N56), 
        .CK(i_data_even_addr_gen_inst_net2857), .RN(
        i_data_even_addr_gen_inst_n6), .Q(
        i_data_even_addr_gen_inst_int_offs_addr_1_) );
  SDFFR_X1 i_data_even_addr_gen_inst_int_offs_addr_reg_0_ ( .D(1'b0), .SI(
        i_data_even_addr_gen_inst_n27), .SE(i_data_even_addr_gen_inst_N55), 
        .CK(i_data_even_addr_gen_inst_net2857), .RN(
        i_data_even_addr_gen_inst_n6), .Q(
        i_data_even_addr_gen_inst_int_offs_addr_0_) );
  CLKGATETST_X1 i_data_even_addr_gen_inst_clk_gate_int_base_addr_reg_latch ( 
        .CK(ck), .E(i_data_even_addr_gen_inst_N40), .SE(1'b0), .GCK(
        i_data_even_addr_gen_inst_net2851) );
  CLKGATETST_X1 i_data_even_addr_gen_inst_clk_gate_int_offs_addr_reg_latch ( 
        .CK(ck), .E(i_data_even_addr_gen_inst_N65), .SE(1'b0), .GCK(
        i_data_even_addr_gen_inst_net2857) );
  XOR2_X1 i_data_even_addr_gen_inst_add_60_U2 ( .A(1'b1), .B(
        i_data_even_addr_gen_inst_int_offs_addr_0_), .Z(
        i_data_even_addr_gen_inst_N55) );
  AND2_X1 i_data_even_addr_gen_inst_add_60_U1 ( .A1(1'b1), .A2(
        i_data_even_addr_gen_inst_int_offs_addr_0_), .ZN(
        i_data_even_addr_gen_inst_add_60_n1) );
  FA_X1 i_data_even_addr_gen_inst_add_60_U1_1 ( .A(
        i_data_even_addr_gen_inst_int_offs_addr_1_), .B(1'b0), .CI(
        i_data_even_addr_gen_inst_add_60_n1), .CO(
        i_data_even_addr_gen_inst_add_60_carry[2]), .S(
        i_data_even_addr_gen_inst_N56) );
  FA_X1 i_data_even_addr_gen_inst_add_60_U1_2 ( .A(
        i_data_even_addr_gen_inst_int_offs_addr_2_), .B(1'b0), .CI(
        i_data_even_addr_gen_inst_add_60_carry[2]), .CO(
        i_data_even_addr_gen_inst_add_60_carry[3]), .S(
        i_data_even_addr_gen_inst_N57) );
  FA_X1 i_data_even_addr_gen_inst_add_60_U1_3 ( .A(
        i_data_even_addr_gen_inst_int_offs_addr_3_), .B(1'b0), .CI(
        i_data_even_addr_gen_inst_add_60_carry[3]), .CO(
        i_data_even_addr_gen_inst_add_60_carry[4]), .S(
        i_data_even_addr_gen_inst_N58) );
  FA_X1 i_data_even_addr_gen_inst_add_60_U1_4 ( .A(
        i_data_even_addr_gen_inst_int_offs_addr_4_), .B(1'b0), .CI(
        i_data_even_addr_gen_inst_add_60_carry[4]), .CO(
        i_data_even_addr_gen_inst_add_60_carry[5]), .S(
        i_data_even_addr_gen_inst_N59) );
  FA_X1 i_data_even_addr_gen_inst_add_60_U1_5 ( .A(
        i_data_even_addr_gen_inst_int_offs_addr_5_), .B(1'b0), .CI(
        i_data_even_addr_gen_inst_add_60_carry[5]), .CO(
        i_data_even_addr_gen_inst_add_60_carry[6]), .S(
        i_data_even_addr_gen_inst_N60) );
  FA_X1 i_data_even_addr_gen_inst_add_60_U1_6 ( .A(
        i_data_even_addr_gen_inst_int_offs_addr_6_), .B(1'b0), .CI(
        i_data_even_addr_gen_inst_add_60_carry[6]), .CO(
        i_data_even_addr_gen_inst_add_60_carry[7]), .S(
        i_data_even_addr_gen_inst_N61) );
  FA_X1 i_data_even_addr_gen_inst_add_60_U1_7 ( .A(
        i_data_even_addr_gen_inst_int_offs_addr_7_), .B(1'b0), .CI(
        i_data_even_addr_gen_inst_add_60_carry[7]), .CO(
        i_data_even_addr_gen_inst_add_60_carry[8]), .S(
        i_data_even_addr_gen_inst_N62) );
  FA_X1 i_data_even_addr_gen_inst_add_60_U1_8 ( .A(
        i_data_even_addr_gen_inst_int_offs_addr_8_), .B(1'b0), .CI(
        i_data_even_addr_gen_inst_add_60_carry[8]), .CO(
        i_data_even_addr_gen_inst_add_60_carry[9]), .S(
        i_data_even_addr_gen_inst_N63) );
  FA_X1 i_data_even_addr_gen_inst_add_60_U1_9 ( .A(
        i_data_even_addr_gen_inst_int_offs_addr_9_), .B(1'b0), .CI(
        i_data_even_addr_gen_inst_add_60_carry[9]), .S(
        i_data_even_addr_gen_inst_N64) );
  AND2_X1 i_data_even_addr_gen_inst_add_45_U2 ( .A1(1'b1), .A2(
        i_data_even_addr_gen_inst_int_base_addr_0_), .ZN(
        i_data_even_addr_gen_inst_add_45_n2) );
  XOR2_X1 i_data_even_addr_gen_inst_add_45_U1 ( .A(1'b1), .B(
        i_data_even_addr_gen_inst_int_base_addr_0_), .Z(
        i_data_even_addr_gen_inst_N20) );
  FA_X1 i_data_even_addr_gen_inst_add_45_U1_1 ( .A(
        i_data_even_addr_gen_inst_int_base_addr_1_), .B(1'b0), .CI(
        i_data_even_addr_gen_inst_add_45_n2), .CO(
        i_data_even_addr_gen_inst_add_45_carry[2]), .S(
        i_data_even_addr_gen_inst_N21) );
  FA_X1 i_data_even_addr_gen_inst_add_45_U1_2 ( .A(
        i_data_even_addr_gen_inst_int_base_addr_2_), .B(1'b0), .CI(
        i_data_even_addr_gen_inst_add_45_carry[2]), .CO(
        i_data_even_addr_gen_inst_add_45_carry[3]), .S(
        i_data_even_addr_gen_inst_N22) );
  FA_X1 i_data_even_addr_gen_inst_add_45_U1_3 ( .A(
        i_data_even_addr_gen_inst_int_base_addr_3_), .B(1'b0), .CI(
        i_data_even_addr_gen_inst_add_45_carry[3]), .CO(
        i_data_even_addr_gen_inst_add_45_carry[4]), .S(
        i_data_even_addr_gen_inst_N23) );
  FA_X1 i_data_even_addr_gen_inst_add_45_U1_4 ( .A(
        i_data_even_addr_gen_inst_int_base_addr_4_), .B(1'b0), .CI(
        i_data_even_addr_gen_inst_add_45_carry[4]), .CO(
        i_data_even_addr_gen_inst_add_45_carry[5]), .S(
        i_data_even_addr_gen_inst_N24) );
  FA_X1 i_data_even_addr_gen_inst_add_45_U1_5 ( .A(
        i_data_even_addr_gen_inst_int_base_addr_5_), .B(1'b0), .CI(
        i_data_even_addr_gen_inst_add_45_carry[5]), .CO(
        i_data_even_addr_gen_inst_add_45_carry[6]), .S(
        i_data_even_addr_gen_inst_N25) );
  FA_X1 i_data_even_addr_gen_inst_add_45_U1_6 ( .A(
        i_data_even_addr_gen_inst_int_base_addr_6_), .B(1'b0), .CI(
        i_data_even_addr_gen_inst_add_45_carry[6]), .CO(
        i_data_even_addr_gen_inst_add_45_carry[7]), .S(
        i_data_even_addr_gen_inst_N26) );
  FA_X1 i_data_even_addr_gen_inst_add_45_U1_7 ( .A(
        i_data_even_addr_gen_inst_int_base_addr_7_), .B(1'b0), .CI(
        i_data_even_addr_gen_inst_add_45_carry[7]), .CO(
        i_data_even_addr_gen_inst_add_45_carry[8]), .S(
        i_data_even_addr_gen_inst_N27) );
  FA_X1 i_data_even_addr_gen_inst_add_45_U1_8 ( .A(
        i_data_even_addr_gen_inst_int_base_addr_8_), .B(1'b0), .CI(
        i_data_even_addr_gen_inst_add_45_carry[8]), .CO(
        i_data_even_addr_gen_inst_add_45_carry[9]), .S(
        i_data_even_addr_gen_inst_N28) );
  FA_X1 i_data_even_addr_gen_inst_add_45_U1_9 ( .A(
        i_data_even_addr_gen_inst_int_base_addr_9_), .B(1'b0), .CI(
        i_data_even_addr_gen_inst_add_45_carry[9]), .S(
        i_data_even_addr_gen_inst_N29) );
  AND2_X1 i_data_even_addr_gen_inst_add_43_U2 ( .A1(1'b1), .A2(
        i_data_even_addr[0]), .ZN(i_data_even_addr_gen_inst_add_43_n2) );
  XOR2_X1 i_data_even_addr_gen_inst_add_43_U1 ( .A(1'b1), .B(
        i_data_even_addr[0]), .Z(i_data_even_addr_gen_inst_N10) );
  FA_X1 i_data_even_addr_gen_inst_add_43_U1_1 ( .A(i_data_even_addr[1]), .B(
        1'b0), .CI(i_data_even_addr_gen_inst_add_43_n2), .CO(
        i_data_even_addr_gen_inst_add_43_carry[2]), .S(
        i_data_even_addr_gen_inst_N11) );
  FA_X1 i_data_even_addr_gen_inst_add_43_U1_2 ( .A(i_data_even_addr[2]), .B(
        1'b0), .CI(i_data_even_addr_gen_inst_add_43_carry[2]), .CO(
        i_data_even_addr_gen_inst_add_43_carry[3]), .S(
        i_data_even_addr_gen_inst_N12) );
  FA_X1 i_data_even_addr_gen_inst_add_43_U1_3 ( .A(i_data_even_addr[3]), .B(
        1'b0), .CI(i_data_even_addr_gen_inst_add_43_carry[3]), .CO(
        i_data_even_addr_gen_inst_add_43_carry[4]), .S(
        i_data_even_addr_gen_inst_N13) );
  FA_X1 i_data_even_addr_gen_inst_add_43_U1_4 ( .A(i_data_even_addr[4]), .B(
        1'b0), .CI(i_data_even_addr_gen_inst_add_43_carry[4]), .CO(
        i_data_even_addr_gen_inst_add_43_carry[5]), .S(
        i_data_even_addr_gen_inst_N14) );
  FA_X1 i_data_even_addr_gen_inst_add_43_U1_5 ( .A(i_data_even_addr[5]), .B(
        1'b0), .CI(i_data_even_addr_gen_inst_add_43_carry[5]), .CO(
        i_data_even_addr_gen_inst_add_43_carry[6]), .S(
        i_data_even_addr_gen_inst_N15) );
  FA_X1 i_data_even_addr_gen_inst_add_43_U1_6 ( .A(i_data_even_addr[6]), .B(
        1'b0), .CI(i_data_even_addr_gen_inst_add_43_carry[6]), .CO(
        i_data_even_addr_gen_inst_add_43_carry[7]), .S(
        i_data_even_addr_gen_inst_N16) );
  FA_X1 i_data_even_addr_gen_inst_add_43_U1_7 ( .A(i_data_even_addr[7]), .B(
        1'b0), .CI(i_data_even_addr_gen_inst_add_43_carry[7]), .CO(
        i_data_even_addr_gen_inst_add_43_carry[8]), .S(
        i_data_even_addr_gen_inst_N17) );
  FA_X1 i_data_even_addr_gen_inst_add_43_U1_8 ( .A(i_data_even_addr[8]), .B(
        1'b0), .CI(i_data_even_addr_gen_inst_add_43_carry[8]), .CO(
        i_data_even_addr_gen_inst_add_43_carry[9]), .S(
        i_data_even_addr_gen_inst_N18) );
  FA_X1 i_data_even_addr_gen_inst_add_43_U1_9 ( .A(i_data_even_addr[9]), .B(
        1'b0), .CI(i_data_even_addr_gen_inst_add_43_carry[9]), .S(
        i_data_even_addr_gen_inst_N19) );
  AND2_X1 i_data_even_addr_gen_inst_add_31_U2 ( .A1(
        i_data_even_addr_gen_inst_int_offs_addr_0_), .A2(
        i_data_even_addr_gen_inst_int_base_addr_0_), .ZN(
        i_data_even_addr_gen_inst_add_31_n2) );
  XOR2_X1 i_data_even_addr_gen_inst_add_31_U1 ( .A(
        i_data_even_addr_gen_inst_int_offs_addr_0_), .B(
        i_data_even_addr_gen_inst_int_base_addr_0_), .Z(i_data_even_addr[0])
         );
  FA_X1 i_data_even_addr_gen_inst_add_31_U1_1 ( .A(
        i_data_even_addr_gen_inst_int_base_addr_1_), .B(
        i_data_even_addr_gen_inst_int_offs_addr_1_), .CI(
        i_data_even_addr_gen_inst_add_31_n2), .CO(
        i_data_even_addr_gen_inst_add_31_carry[2]), .S(i_data_even_addr[1]) );
  FA_X1 i_data_even_addr_gen_inst_add_31_U1_2 ( .A(
        i_data_even_addr_gen_inst_int_base_addr_2_), .B(
        i_data_even_addr_gen_inst_int_offs_addr_2_), .CI(
        i_data_even_addr_gen_inst_add_31_carry[2]), .CO(
        i_data_even_addr_gen_inst_add_31_carry[3]), .S(i_data_even_addr[2]) );
  FA_X1 i_data_even_addr_gen_inst_add_31_U1_3 ( .A(
        i_data_even_addr_gen_inst_int_base_addr_3_), .B(
        i_data_even_addr_gen_inst_int_offs_addr_3_), .CI(
        i_data_even_addr_gen_inst_add_31_carry[3]), .CO(
        i_data_even_addr_gen_inst_add_31_carry[4]), .S(i_data_even_addr[3]) );
  FA_X1 i_data_even_addr_gen_inst_add_31_U1_4 ( .A(
        i_data_even_addr_gen_inst_int_base_addr_4_), .B(
        i_data_even_addr_gen_inst_int_offs_addr_4_), .CI(
        i_data_even_addr_gen_inst_add_31_carry[4]), .CO(
        i_data_even_addr_gen_inst_add_31_carry[5]), .S(i_data_even_addr[4]) );
  FA_X1 i_data_even_addr_gen_inst_add_31_U1_5 ( .A(
        i_data_even_addr_gen_inst_int_base_addr_5_), .B(
        i_data_even_addr_gen_inst_int_offs_addr_5_), .CI(
        i_data_even_addr_gen_inst_add_31_carry[5]), .CO(
        i_data_even_addr_gen_inst_add_31_carry[6]), .S(i_data_even_addr[5]) );
  FA_X1 i_data_even_addr_gen_inst_add_31_U1_6 ( .A(
        i_data_even_addr_gen_inst_int_base_addr_6_), .B(
        i_data_even_addr_gen_inst_int_offs_addr_6_), .CI(
        i_data_even_addr_gen_inst_add_31_carry[6]), .CO(
        i_data_even_addr_gen_inst_add_31_carry[7]), .S(i_data_even_addr[6]) );
  FA_X1 i_data_even_addr_gen_inst_add_31_U1_7 ( .A(
        i_data_even_addr_gen_inst_int_base_addr_7_), .B(
        i_data_even_addr_gen_inst_int_offs_addr_7_), .CI(
        i_data_even_addr_gen_inst_add_31_carry[7]), .CO(
        i_data_even_addr_gen_inst_add_31_carry[8]), .S(i_data_even_addr[7]) );
  FA_X1 i_data_even_addr_gen_inst_add_31_U1_8 ( .A(
        i_data_even_addr_gen_inst_int_base_addr_8_), .B(
        i_data_even_addr_gen_inst_int_offs_addr_8_), .CI(
        i_data_even_addr_gen_inst_add_31_carry[8]), .CO(
        i_data_even_addr_gen_inst_add_31_carry[9]), .S(i_data_even_addr[8]) );
  FA_X1 i_data_even_addr_gen_inst_add_31_U1_9 ( .A(
        i_data_even_addr_gen_inst_int_base_addr_9_), .B(
        i_data_even_addr_gen_inst_int_offs_addr_9_), .CI(
        i_data_even_addr_gen_inst_add_31_carry[9]), .S(i_data_even_addr[9]) );
  INV_X1 i_data_odd_addr_gen_inst_U44 ( .A(rst), .ZN(
        i_data_odd_addr_gen_inst_n6) );
  INV_X1 i_data_odd_addr_gen_inst_U43 ( .A(rst), .ZN(
        i_data_odd_addr_gen_inst_n5) );
  AOI22_X1 i_data_odd_addr_gen_inst_U42 ( .A1(i_data_odd_addr_gen_inst_N29), 
        .A2(i_data_odd_addr_gen_inst_n33), .B1(i_data_odd_addr_gen_inst_N19), 
        .B2(i_data_odd_addr_gen_inst_n34), .ZN(i_data_odd_addr_gen_inst_n32)
         );
  INV_X1 i_data_odd_addr_gen_inst_U41 ( .A(i_data_odd_addr_gen_inst_n32), .ZN(
        i_data_odd_addr_gen_inst_n7) );
  OR2_X1 i_data_odd_addr_gen_inst_U40 ( .A1(n33), .A2(ctrl_ldh_v_n), .ZN(
        i_data_odd_addr_gen_inst_N65) );
  AOI22_X1 i_data_odd_addr_gen_inst_U39 ( .A1(i_data_odd_addr_gen_inst_N20), 
        .A2(i_data_odd_addr_gen_inst_n33), .B1(i_data_odd_addr_gen_inst_N10), 
        .B2(i_data_odd_addr_gen_inst_n34), .ZN(i_data_odd_addr_gen_inst_n43)
         );
  INV_X1 i_data_odd_addr_gen_inst_U38 ( .A(i_data_odd_addr_gen_inst_n43), .ZN(
        i_data_odd_addr_gen_inst_n26) );
  AOI22_X1 i_data_odd_addr_gen_inst_U37 ( .A1(i_data_odd_addr_gen_inst_N21), 
        .A2(i_data_odd_addr_gen_inst_n33), .B1(i_data_odd_addr_gen_inst_N11), 
        .B2(i_data_odd_addr_gen_inst_n34), .ZN(i_data_odd_addr_gen_inst_n42)
         );
  INV_X1 i_data_odd_addr_gen_inst_U36 ( .A(i_data_odd_addr_gen_inst_n42), .ZN(
        i_data_odd_addr_gen_inst_n25) );
  AOI22_X1 i_data_odd_addr_gen_inst_U35 ( .A1(i_data_odd_addr_gen_inst_N22), 
        .A2(i_data_odd_addr_gen_inst_n33), .B1(i_data_odd_addr_gen_inst_N12), 
        .B2(i_data_odd_addr_gen_inst_n34), .ZN(i_data_odd_addr_gen_inst_n41)
         );
  INV_X1 i_data_odd_addr_gen_inst_U34 ( .A(i_data_odd_addr_gen_inst_n41), .ZN(
        i_data_odd_addr_gen_inst_n24) );
  AOI22_X1 i_data_odd_addr_gen_inst_U33 ( .A1(i_data_odd_addr_gen_inst_N23), 
        .A2(i_data_odd_addr_gen_inst_n33), .B1(i_data_odd_addr_gen_inst_N13), 
        .B2(i_data_odd_addr_gen_inst_n34), .ZN(i_data_odd_addr_gen_inst_n40)
         );
  INV_X1 i_data_odd_addr_gen_inst_U32 ( .A(i_data_odd_addr_gen_inst_n40), .ZN(
        i_data_odd_addr_gen_inst_n23) );
  AOI22_X1 i_data_odd_addr_gen_inst_U31 ( .A1(i_data_odd_addr_gen_inst_N24), 
        .A2(i_data_odd_addr_gen_inst_n33), .B1(i_data_odd_addr_gen_inst_N14), 
        .B2(i_data_odd_addr_gen_inst_n34), .ZN(i_data_odd_addr_gen_inst_n39)
         );
  INV_X1 i_data_odd_addr_gen_inst_U30 ( .A(i_data_odd_addr_gen_inst_n39), .ZN(
        i_data_odd_addr_gen_inst_n22) );
  AOI22_X1 i_data_odd_addr_gen_inst_U29 ( .A1(i_data_odd_addr_gen_inst_N25), 
        .A2(i_data_odd_addr_gen_inst_n33), .B1(i_data_odd_addr_gen_inst_N15), 
        .B2(i_data_odd_addr_gen_inst_n34), .ZN(i_data_odd_addr_gen_inst_n38)
         );
  INV_X1 i_data_odd_addr_gen_inst_U28 ( .A(i_data_odd_addr_gen_inst_n38), .ZN(
        i_data_odd_addr_gen_inst_n21) );
  AOI22_X1 i_data_odd_addr_gen_inst_U27 ( .A1(i_data_odd_addr_gen_inst_N26), 
        .A2(i_data_odd_addr_gen_inst_n33), .B1(i_data_odd_addr_gen_inst_N16), 
        .B2(i_data_odd_addr_gen_inst_n34), .ZN(i_data_odd_addr_gen_inst_n37)
         );
  INV_X1 i_data_odd_addr_gen_inst_U26 ( .A(i_data_odd_addr_gen_inst_n37), .ZN(
        i_data_odd_addr_gen_inst_n20) );
  AOI22_X1 i_data_odd_addr_gen_inst_U25 ( .A1(i_data_odd_addr_gen_inst_N27), 
        .A2(i_data_odd_addr_gen_inst_n33), .B1(i_data_odd_addr_gen_inst_N17), 
        .B2(i_data_odd_addr_gen_inst_n34), .ZN(i_data_odd_addr_gen_inst_n36)
         );
  INV_X1 i_data_odd_addr_gen_inst_U24 ( .A(i_data_odd_addr_gen_inst_n36), .ZN(
        i_data_odd_addr_gen_inst_n18) );
  AOI22_X1 i_data_odd_addr_gen_inst_U23 ( .A1(i_data_odd_addr_gen_inst_N28), 
        .A2(i_data_odd_addr_gen_inst_n33), .B1(i_data_odd_addr_gen_inst_N18), 
        .B2(i_data_odd_addr_gen_inst_n34), .ZN(i_data_odd_addr_gen_inst_n35)
         );
  INV_X1 i_data_odd_addr_gen_inst_U22 ( .A(i_data_odd_addr_gen_inst_n35), .ZN(
        i_data_odd_addr_gen_inst_n8) );
  OR2_X1 i_data_odd_addr_gen_inst_U21 ( .A1(int_c_i_en_odd), .A2(int_en_L4_ptr), .ZN(i_data_odd_addr_gen_inst_N40) );
  INV_X1 i_data_odd_addr_gen_inst_U20 ( .A(int_c_i_en_odd), .ZN(
        i_data_odd_addr_gen_inst_n28) );
  NOR2_X1 i_data_odd_addr_gen_inst_U19 ( .A1(i_data_odd_addr_gen_inst_n28), 
        .A2(int_en_L4_ptr), .ZN(i_data_odd_addr_gen_inst_n34) );
  NOR2_X1 i_data_odd_addr_gen_inst_U18 ( .A1(int_c_i_en_odd), .A2(
        int_en_L4_ptr), .ZN(i_data_odd_addr_gen_inst_n33) );
  INV_X1 i_data_odd_addr_gen_inst_U16 ( .A(n33), .ZN(
        i_data_odd_addr_gen_inst_n27) );
  DFFR_X1 i_data_odd_addr_gen_inst_int_base_addr_reg_8_ ( .D(
        i_data_odd_addr_gen_inst_n8), .CK(i_data_odd_addr_gen_inst_net2828), 
        .RN(i_data_odd_addr_gen_inst_n5), .Q(
        i_data_odd_addr_gen_inst_int_base_addr_8_) );
  DFFR_X1 i_data_odd_addr_gen_inst_int_base_addr_reg_7_ ( .D(
        i_data_odd_addr_gen_inst_n18), .CK(i_data_odd_addr_gen_inst_net2828), 
        .RN(i_data_odd_addr_gen_inst_n5), .Q(
        i_data_odd_addr_gen_inst_int_base_addr_7_) );
  DFFR_X1 i_data_odd_addr_gen_inst_int_base_addr_reg_6_ ( .D(
        i_data_odd_addr_gen_inst_n20), .CK(i_data_odd_addr_gen_inst_net2828), 
        .RN(i_data_odd_addr_gen_inst_n5), .Q(
        i_data_odd_addr_gen_inst_int_base_addr_6_) );
  DFFR_X1 i_data_odd_addr_gen_inst_int_base_addr_reg_5_ ( .D(
        i_data_odd_addr_gen_inst_n21), .CK(i_data_odd_addr_gen_inst_net2828), 
        .RN(i_data_odd_addr_gen_inst_n5), .Q(
        i_data_odd_addr_gen_inst_int_base_addr_5_) );
  DFFR_X1 i_data_odd_addr_gen_inst_int_base_addr_reg_4_ ( .D(
        i_data_odd_addr_gen_inst_n22), .CK(i_data_odd_addr_gen_inst_net2828), 
        .RN(i_data_odd_addr_gen_inst_n5), .Q(
        i_data_odd_addr_gen_inst_int_base_addr_4_) );
  DFFR_X1 i_data_odd_addr_gen_inst_int_base_addr_reg_3_ ( .D(
        i_data_odd_addr_gen_inst_n23), .CK(i_data_odd_addr_gen_inst_net2828), 
        .RN(i_data_odd_addr_gen_inst_n5), .Q(
        i_data_odd_addr_gen_inst_int_base_addr_3_) );
  DFFR_X1 i_data_odd_addr_gen_inst_int_base_addr_reg_2_ ( .D(
        i_data_odd_addr_gen_inst_n24), .CK(i_data_odd_addr_gen_inst_net2828), 
        .RN(i_data_odd_addr_gen_inst_n5), .Q(
        i_data_odd_addr_gen_inst_int_base_addr_2_) );
  DFFR_X1 i_data_odd_addr_gen_inst_int_base_addr_reg_1_ ( .D(
        i_data_odd_addr_gen_inst_n25), .CK(i_data_odd_addr_gen_inst_net2828), 
        .RN(i_data_odd_addr_gen_inst_n5), .Q(
        i_data_odd_addr_gen_inst_int_base_addr_1_) );
  DFFR_X1 i_data_odd_addr_gen_inst_int_base_addr_reg_0_ ( .D(
        i_data_odd_addr_gen_inst_n26), .CK(i_data_odd_addr_gen_inst_net2828), 
        .RN(i_data_odd_addr_gen_inst_n5), .Q(
        i_data_odd_addr_gen_inst_int_base_addr_0_) );
  DFFR_X1 i_data_odd_addr_gen_inst_int_base_addr_reg_9_ ( .D(
        i_data_odd_addr_gen_inst_n7), .CK(i_data_odd_addr_gen_inst_net2828), 
        .RN(i_data_odd_addr_gen_inst_n5), .Q(
        i_data_odd_addr_gen_inst_int_base_addr_9_) );
  SDFFR_X1 i_data_odd_addr_gen_inst_int_offs_addr_reg_9_ ( .D(1'b0), .SI(
        i_data_odd_addr_gen_inst_n27), .SE(i_data_odd_addr_gen_inst_N64), .CK(
        i_data_odd_addr_gen_inst_net2834), .RN(i_data_odd_addr_gen_inst_n5), 
        .Q(i_data_odd_addr_gen_inst_int_offs_addr_9_) );
  SDFFR_X1 i_data_odd_addr_gen_inst_int_offs_addr_reg_8_ ( .D(1'b0), .SI(
        i_data_odd_addr_gen_inst_n27), .SE(i_data_odd_addr_gen_inst_N63), .CK(
        i_data_odd_addr_gen_inst_net2834), .RN(i_data_odd_addr_gen_inst_n5), 
        .Q(i_data_odd_addr_gen_inst_int_offs_addr_8_) );
  SDFFR_X1 i_data_odd_addr_gen_inst_int_offs_addr_reg_7_ ( .D(1'b0), .SI(
        i_data_odd_addr_gen_inst_n27), .SE(i_data_odd_addr_gen_inst_N62), .CK(
        i_data_odd_addr_gen_inst_net2834), .RN(i_data_odd_addr_gen_inst_n6), 
        .Q(i_data_odd_addr_gen_inst_int_offs_addr_7_) );
  SDFFR_X1 i_data_odd_addr_gen_inst_int_offs_addr_reg_6_ ( .D(1'b0), .SI(
        i_data_odd_addr_gen_inst_n27), .SE(i_data_odd_addr_gen_inst_N61), .CK(
        i_data_odd_addr_gen_inst_net2834), .RN(i_data_odd_addr_gen_inst_n6), 
        .Q(i_data_odd_addr_gen_inst_int_offs_addr_6_) );
  SDFFR_X1 i_data_odd_addr_gen_inst_int_offs_addr_reg_5_ ( .D(1'b0), .SI(
        i_data_odd_addr_gen_inst_n27), .SE(i_data_odd_addr_gen_inst_N60), .CK(
        i_data_odd_addr_gen_inst_net2834), .RN(i_data_odd_addr_gen_inst_n6), 
        .Q(i_data_odd_addr_gen_inst_int_offs_addr_5_) );
  SDFFR_X1 i_data_odd_addr_gen_inst_int_offs_addr_reg_4_ ( .D(1'b0), .SI(
        i_data_odd_addr_gen_inst_n27), .SE(i_data_odd_addr_gen_inst_N59), .CK(
        i_data_odd_addr_gen_inst_net2834), .RN(i_data_odd_addr_gen_inst_n6), 
        .Q(i_data_odd_addr_gen_inst_int_offs_addr_4_) );
  SDFFR_X1 i_data_odd_addr_gen_inst_int_offs_addr_reg_3_ ( .D(1'b0), .SI(
        i_data_odd_addr_gen_inst_n27), .SE(i_data_odd_addr_gen_inst_N58), .CK(
        i_data_odd_addr_gen_inst_net2834), .RN(i_data_odd_addr_gen_inst_n6), 
        .Q(i_data_odd_addr_gen_inst_int_offs_addr_3_) );
  SDFFR_X1 i_data_odd_addr_gen_inst_int_offs_addr_reg_2_ ( .D(1'b0), .SI(
        i_data_odd_addr_gen_inst_n27), .SE(i_data_odd_addr_gen_inst_N57), .CK(
        i_data_odd_addr_gen_inst_net2834), .RN(i_data_odd_addr_gen_inst_n6), 
        .Q(i_data_odd_addr_gen_inst_int_offs_addr_2_) );
  SDFFR_X1 i_data_odd_addr_gen_inst_int_offs_addr_reg_1_ ( .D(1'b0), .SI(
        i_data_odd_addr_gen_inst_n27), .SE(i_data_odd_addr_gen_inst_N56), .CK(
        i_data_odd_addr_gen_inst_net2834), .RN(i_data_odd_addr_gen_inst_n6), 
        .Q(i_data_odd_addr_gen_inst_int_offs_addr_1_) );
  SDFFR_X1 i_data_odd_addr_gen_inst_int_offs_addr_reg_0_ ( .D(1'b0), .SI(
        i_data_odd_addr_gen_inst_n27), .SE(i_data_odd_addr_gen_inst_N55), .CK(
        i_data_odd_addr_gen_inst_net2834), .RN(i_data_odd_addr_gen_inst_n6), 
        .Q(i_data_odd_addr_gen_inst_int_offs_addr_0_) );
  CLKGATETST_X1 i_data_odd_addr_gen_inst_clk_gate_int_base_addr_reg_latch ( 
        .CK(ck), .E(i_data_odd_addr_gen_inst_N40), .SE(1'b0), .GCK(
        i_data_odd_addr_gen_inst_net2828) );
  CLKGATETST_X1 i_data_odd_addr_gen_inst_clk_gate_int_offs_addr_reg_latch ( 
        .CK(ck), .E(i_data_odd_addr_gen_inst_N65), .SE(1'b0), .GCK(
        i_data_odd_addr_gen_inst_net2834) );
  XOR2_X1 i_data_odd_addr_gen_inst_add_60_U2 ( .A(1'b1), .B(
        i_data_odd_addr_gen_inst_int_offs_addr_0_), .Z(
        i_data_odd_addr_gen_inst_N55) );
  AND2_X1 i_data_odd_addr_gen_inst_add_60_U1 ( .A1(1'b1), .A2(
        i_data_odd_addr_gen_inst_int_offs_addr_0_), .ZN(
        i_data_odd_addr_gen_inst_add_60_n1) );
  FA_X1 i_data_odd_addr_gen_inst_add_60_U1_1 ( .A(
        i_data_odd_addr_gen_inst_int_offs_addr_1_), .B(1'b0), .CI(
        i_data_odd_addr_gen_inst_add_60_n1), .CO(
        i_data_odd_addr_gen_inst_add_60_carry[2]), .S(
        i_data_odd_addr_gen_inst_N56) );
  FA_X1 i_data_odd_addr_gen_inst_add_60_U1_2 ( .A(
        i_data_odd_addr_gen_inst_int_offs_addr_2_), .B(1'b0), .CI(
        i_data_odd_addr_gen_inst_add_60_carry[2]), .CO(
        i_data_odd_addr_gen_inst_add_60_carry[3]), .S(
        i_data_odd_addr_gen_inst_N57) );
  FA_X1 i_data_odd_addr_gen_inst_add_60_U1_3 ( .A(
        i_data_odd_addr_gen_inst_int_offs_addr_3_), .B(1'b0), .CI(
        i_data_odd_addr_gen_inst_add_60_carry[3]), .CO(
        i_data_odd_addr_gen_inst_add_60_carry[4]), .S(
        i_data_odd_addr_gen_inst_N58) );
  FA_X1 i_data_odd_addr_gen_inst_add_60_U1_4 ( .A(
        i_data_odd_addr_gen_inst_int_offs_addr_4_), .B(1'b0), .CI(
        i_data_odd_addr_gen_inst_add_60_carry[4]), .CO(
        i_data_odd_addr_gen_inst_add_60_carry[5]), .S(
        i_data_odd_addr_gen_inst_N59) );
  FA_X1 i_data_odd_addr_gen_inst_add_60_U1_5 ( .A(
        i_data_odd_addr_gen_inst_int_offs_addr_5_), .B(1'b0), .CI(
        i_data_odd_addr_gen_inst_add_60_carry[5]), .CO(
        i_data_odd_addr_gen_inst_add_60_carry[6]), .S(
        i_data_odd_addr_gen_inst_N60) );
  FA_X1 i_data_odd_addr_gen_inst_add_60_U1_6 ( .A(
        i_data_odd_addr_gen_inst_int_offs_addr_6_), .B(1'b0), .CI(
        i_data_odd_addr_gen_inst_add_60_carry[6]), .CO(
        i_data_odd_addr_gen_inst_add_60_carry[7]), .S(
        i_data_odd_addr_gen_inst_N61) );
  FA_X1 i_data_odd_addr_gen_inst_add_60_U1_7 ( .A(
        i_data_odd_addr_gen_inst_int_offs_addr_7_), .B(1'b0), .CI(
        i_data_odd_addr_gen_inst_add_60_carry[7]), .CO(
        i_data_odd_addr_gen_inst_add_60_carry[8]), .S(
        i_data_odd_addr_gen_inst_N62) );
  FA_X1 i_data_odd_addr_gen_inst_add_60_U1_8 ( .A(
        i_data_odd_addr_gen_inst_int_offs_addr_8_), .B(1'b0), .CI(
        i_data_odd_addr_gen_inst_add_60_carry[8]), .CO(
        i_data_odd_addr_gen_inst_add_60_carry[9]), .S(
        i_data_odd_addr_gen_inst_N63) );
  FA_X1 i_data_odd_addr_gen_inst_add_60_U1_9 ( .A(
        i_data_odd_addr_gen_inst_int_offs_addr_9_), .B(1'b0), .CI(
        i_data_odd_addr_gen_inst_add_60_carry[9]), .S(
        i_data_odd_addr_gen_inst_N64) );
  AND2_X1 i_data_odd_addr_gen_inst_add_45_U2 ( .A1(1'b1), .A2(
        i_data_odd_addr_gen_inst_int_base_addr_0_), .ZN(
        i_data_odd_addr_gen_inst_add_45_n2) );
  XOR2_X1 i_data_odd_addr_gen_inst_add_45_U1 ( .A(1'b1), .B(
        i_data_odd_addr_gen_inst_int_base_addr_0_), .Z(
        i_data_odd_addr_gen_inst_N20) );
  FA_X1 i_data_odd_addr_gen_inst_add_45_U1_1 ( .A(
        i_data_odd_addr_gen_inst_int_base_addr_1_), .B(1'b0), .CI(
        i_data_odd_addr_gen_inst_add_45_n2), .CO(
        i_data_odd_addr_gen_inst_add_45_carry[2]), .S(
        i_data_odd_addr_gen_inst_N21) );
  FA_X1 i_data_odd_addr_gen_inst_add_45_U1_2 ( .A(
        i_data_odd_addr_gen_inst_int_base_addr_2_), .B(1'b0), .CI(
        i_data_odd_addr_gen_inst_add_45_carry[2]), .CO(
        i_data_odd_addr_gen_inst_add_45_carry[3]), .S(
        i_data_odd_addr_gen_inst_N22) );
  FA_X1 i_data_odd_addr_gen_inst_add_45_U1_3 ( .A(
        i_data_odd_addr_gen_inst_int_base_addr_3_), .B(1'b0), .CI(
        i_data_odd_addr_gen_inst_add_45_carry[3]), .CO(
        i_data_odd_addr_gen_inst_add_45_carry[4]), .S(
        i_data_odd_addr_gen_inst_N23) );
  FA_X1 i_data_odd_addr_gen_inst_add_45_U1_4 ( .A(
        i_data_odd_addr_gen_inst_int_base_addr_4_), .B(1'b0), .CI(
        i_data_odd_addr_gen_inst_add_45_carry[4]), .CO(
        i_data_odd_addr_gen_inst_add_45_carry[5]), .S(
        i_data_odd_addr_gen_inst_N24) );
  FA_X1 i_data_odd_addr_gen_inst_add_45_U1_5 ( .A(
        i_data_odd_addr_gen_inst_int_base_addr_5_), .B(1'b0), .CI(
        i_data_odd_addr_gen_inst_add_45_carry[5]), .CO(
        i_data_odd_addr_gen_inst_add_45_carry[6]), .S(
        i_data_odd_addr_gen_inst_N25) );
  FA_X1 i_data_odd_addr_gen_inst_add_45_U1_6 ( .A(
        i_data_odd_addr_gen_inst_int_base_addr_6_), .B(1'b0), .CI(
        i_data_odd_addr_gen_inst_add_45_carry[6]), .CO(
        i_data_odd_addr_gen_inst_add_45_carry[7]), .S(
        i_data_odd_addr_gen_inst_N26) );
  FA_X1 i_data_odd_addr_gen_inst_add_45_U1_7 ( .A(
        i_data_odd_addr_gen_inst_int_base_addr_7_), .B(1'b0), .CI(
        i_data_odd_addr_gen_inst_add_45_carry[7]), .CO(
        i_data_odd_addr_gen_inst_add_45_carry[8]), .S(
        i_data_odd_addr_gen_inst_N27) );
  FA_X1 i_data_odd_addr_gen_inst_add_45_U1_8 ( .A(
        i_data_odd_addr_gen_inst_int_base_addr_8_), .B(1'b0), .CI(
        i_data_odd_addr_gen_inst_add_45_carry[8]), .CO(
        i_data_odd_addr_gen_inst_add_45_carry[9]), .S(
        i_data_odd_addr_gen_inst_N28) );
  FA_X1 i_data_odd_addr_gen_inst_add_45_U1_9 ( .A(
        i_data_odd_addr_gen_inst_int_base_addr_9_), .B(1'b0), .CI(
        i_data_odd_addr_gen_inst_add_45_carry[9]), .S(
        i_data_odd_addr_gen_inst_N29) );
  AND2_X1 i_data_odd_addr_gen_inst_add_43_U2 ( .A1(1'b1), .A2(
        i_data_odd_addr[0]), .ZN(i_data_odd_addr_gen_inst_add_43_n2) );
  XOR2_X1 i_data_odd_addr_gen_inst_add_43_U1 ( .A(1'b1), .B(i_data_odd_addr[0]), .Z(i_data_odd_addr_gen_inst_N10) );
  FA_X1 i_data_odd_addr_gen_inst_add_43_U1_1 ( .A(i_data_odd_addr[1]), .B(1'b0), .CI(i_data_odd_addr_gen_inst_add_43_n2), .CO(
        i_data_odd_addr_gen_inst_add_43_carry[2]), .S(
        i_data_odd_addr_gen_inst_N11) );
  FA_X1 i_data_odd_addr_gen_inst_add_43_U1_2 ( .A(i_data_odd_addr[2]), .B(1'b0), .CI(i_data_odd_addr_gen_inst_add_43_carry[2]), .CO(
        i_data_odd_addr_gen_inst_add_43_carry[3]), .S(
        i_data_odd_addr_gen_inst_N12) );
  FA_X1 i_data_odd_addr_gen_inst_add_43_U1_3 ( .A(i_data_odd_addr[3]), .B(1'b0), .CI(i_data_odd_addr_gen_inst_add_43_carry[3]), .CO(
        i_data_odd_addr_gen_inst_add_43_carry[4]), .S(
        i_data_odd_addr_gen_inst_N13) );
  FA_X1 i_data_odd_addr_gen_inst_add_43_U1_4 ( .A(i_data_odd_addr[4]), .B(1'b0), .CI(i_data_odd_addr_gen_inst_add_43_carry[4]), .CO(
        i_data_odd_addr_gen_inst_add_43_carry[5]), .S(
        i_data_odd_addr_gen_inst_N14) );
  FA_X1 i_data_odd_addr_gen_inst_add_43_U1_5 ( .A(i_data_odd_addr[5]), .B(1'b0), .CI(i_data_odd_addr_gen_inst_add_43_carry[5]), .CO(
        i_data_odd_addr_gen_inst_add_43_carry[6]), .S(
        i_data_odd_addr_gen_inst_N15) );
  FA_X1 i_data_odd_addr_gen_inst_add_43_U1_6 ( .A(i_data_odd_addr[6]), .B(1'b0), .CI(i_data_odd_addr_gen_inst_add_43_carry[6]), .CO(
        i_data_odd_addr_gen_inst_add_43_carry[7]), .S(
        i_data_odd_addr_gen_inst_N16) );
  FA_X1 i_data_odd_addr_gen_inst_add_43_U1_7 ( .A(i_data_odd_addr[7]), .B(1'b0), .CI(i_data_odd_addr_gen_inst_add_43_carry[7]), .CO(
        i_data_odd_addr_gen_inst_add_43_carry[8]), .S(
        i_data_odd_addr_gen_inst_N17) );
  FA_X1 i_data_odd_addr_gen_inst_add_43_U1_8 ( .A(i_data_odd_addr[8]), .B(1'b0), .CI(i_data_odd_addr_gen_inst_add_43_carry[8]), .CO(
        i_data_odd_addr_gen_inst_add_43_carry[9]), .S(
        i_data_odd_addr_gen_inst_N18) );
  FA_X1 i_data_odd_addr_gen_inst_add_43_U1_9 ( .A(i_data_odd_addr[9]), .B(1'b0), .CI(i_data_odd_addr_gen_inst_add_43_carry[9]), .S(
        i_data_odd_addr_gen_inst_N19) );
  AND2_X1 i_data_odd_addr_gen_inst_add_31_U2 ( .A1(
        i_data_odd_addr_gen_inst_int_offs_addr_0_), .A2(
        i_data_odd_addr_gen_inst_int_base_addr_0_), .ZN(
        i_data_odd_addr_gen_inst_add_31_n2) );
  XOR2_X1 i_data_odd_addr_gen_inst_add_31_U1 ( .A(
        i_data_odd_addr_gen_inst_int_offs_addr_0_), .B(
        i_data_odd_addr_gen_inst_int_base_addr_0_), .Z(i_data_odd_addr[0]) );
  FA_X1 i_data_odd_addr_gen_inst_add_31_U1_1 ( .A(
        i_data_odd_addr_gen_inst_int_base_addr_1_), .B(
        i_data_odd_addr_gen_inst_int_offs_addr_1_), .CI(
        i_data_odd_addr_gen_inst_add_31_n2), .CO(
        i_data_odd_addr_gen_inst_add_31_carry[2]), .S(i_data_odd_addr[1]) );
  FA_X1 i_data_odd_addr_gen_inst_add_31_U1_2 ( .A(
        i_data_odd_addr_gen_inst_int_base_addr_2_), .B(
        i_data_odd_addr_gen_inst_int_offs_addr_2_), .CI(
        i_data_odd_addr_gen_inst_add_31_carry[2]), .CO(
        i_data_odd_addr_gen_inst_add_31_carry[3]), .S(i_data_odd_addr[2]) );
  FA_X1 i_data_odd_addr_gen_inst_add_31_U1_3 ( .A(
        i_data_odd_addr_gen_inst_int_base_addr_3_), .B(
        i_data_odd_addr_gen_inst_int_offs_addr_3_), .CI(
        i_data_odd_addr_gen_inst_add_31_carry[3]), .CO(
        i_data_odd_addr_gen_inst_add_31_carry[4]), .S(i_data_odd_addr[3]) );
  FA_X1 i_data_odd_addr_gen_inst_add_31_U1_4 ( .A(
        i_data_odd_addr_gen_inst_int_base_addr_4_), .B(
        i_data_odd_addr_gen_inst_int_offs_addr_4_), .CI(
        i_data_odd_addr_gen_inst_add_31_carry[4]), .CO(
        i_data_odd_addr_gen_inst_add_31_carry[5]), .S(i_data_odd_addr[4]) );
  FA_X1 i_data_odd_addr_gen_inst_add_31_U1_5 ( .A(
        i_data_odd_addr_gen_inst_int_base_addr_5_), .B(
        i_data_odd_addr_gen_inst_int_offs_addr_5_), .CI(
        i_data_odd_addr_gen_inst_add_31_carry[5]), .CO(
        i_data_odd_addr_gen_inst_add_31_carry[6]), .S(i_data_odd_addr[5]) );
  FA_X1 i_data_odd_addr_gen_inst_add_31_U1_6 ( .A(
        i_data_odd_addr_gen_inst_int_base_addr_6_), .B(
        i_data_odd_addr_gen_inst_int_offs_addr_6_), .CI(
        i_data_odd_addr_gen_inst_add_31_carry[6]), .CO(
        i_data_odd_addr_gen_inst_add_31_carry[7]), .S(i_data_odd_addr[6]) );
  FA_X1 i_data_odd_addr_gen_inst_add_31_U1_7 ( .A(
        i_data_odd_addr_gen_inst_int_base_addr_7_), .B(
        i_data_odd_addr_gen_inst_int_offs_addr_7_), .CI(
        i_data_odd_addr_gen_inst_add_31_carry[7]), .CO(
        i_data_odd_addr_gen_inst_add_31_carry[8]), .S(i_data_odd_addr[7]) );
  FA_X1 i_data_odd_addr_gen_inst_add_31_U1_8 ( .A(
        i_data_odd_addr_gen_inst_int_base_addr_8_), .B(
        i_data_odd_addr_gen_inst_int_offs_addr_8_), .CI(
        i_data_odd_addr_gen_inst_add_31_carry[8]), .CO(
        i_data_odd_addr_gen_inst_add_31_carry[9]), .S(i_data_odd_addr[8]) );
  FA_X1 i_data_odd_addr_gen_inst_add_31_U1_9 ( .A(
        i_data_odd_addr_gen_inst_int_base_addr_9_), .B(
        i_data_odd_addr_gen_inst_int_offs_addr_9_), .CI(
        i_data_odd_addr_gen_inst_add_31_carry[9]), .S(i_data_odd_addr[9]) );
  INV_X1 o_data_even_addr_gen_inst_U44 ( .A(rst), .ZN(
        o_data_even_addr_gen_inst_n6) );
  INV_X1 o_data_even_addr_gen_inst_U43 ( .A(rst), .ZN(
        o_data_even_addr_gen_inst_n5) );
  INV_X1 o_data_even_addr_gen_inst_U42 ( .A(1'b0), .ZN(
        o_data_even_addr_gen_inst_n27) );
  OR2_X1 o_data_even_addr_gen_inst_U41 ( .A1(int_c_o_en_base_odd), .A2(1'b0), 
        .ZN(o_data_even_addr_gen_inst_N40) );
  OR2_X1 o_data_even_addr_gen_inst_U40 ( .A1(int_c_o_en_base_odd), .A2(
        int_c_o_en_offs_even), .ZN(o_data_even_addr_gen_inst_N65) );
  AOI22_X1 o_data_even_addr_gen_inst_U39 ( .A1(o_data_even_addr_gen_inst_N29), 
        .A2(o_data_even_addr_gen_inst_n33), .B1(o_data_even_addr_gen_inst_N19), 
        .B2(o_data_even_addr_gen_inst_n34), .ZN(o_data_even_addr_gen_inst_n32)
         );
  INV_X1 o_data_even_addr_gen_inst_U38 ( .A(o_data_even_addr_gen_inst_n32), 
        .ZN(o_data_even_addr_gen_inst_n7) );
  AOI22_X1 o_data_even_addr_gen_inst_U37 ( .A1(o_data_even_addr_gen_inst_N21), 
        .A2(o_data_even_addr_gen_inst_n33), .B1(o_data_even_addr_gen_inst_N11), 
        .B2(o_data_even_addr_gen_inst_n34), .ZN(o_data_even_addr_gen_inst_n42)
         );
  INV_X1 o_data_even_addr_gen_inst_U36 ( .A(o_data_even_addr_gen_inst_n42), 
        .ZN(o_data_even_addr_gen_inst_n25) );
  AOI22_X1 o_data_even_addr_gen_inst_U35 ( .A1(o_data_even_addr_gen_inst_N22), 
        .A2(o_data_even_addr_gen_inst_n33), .B1(o_data_even_addr_gen_inst_N12), 
        .B2(o_data_even_addr_gen_inst_n34), .ZN(o_data_even_addr_gen_inst_n41)
         );
  INV_X1 o_data_even_addr_gen_inst_U34 ( .A(o_data_even_addr_gen_inst_n41), 
        .ZN(o_data_even_addr_gen_inst_n24) );
  AOI22_X1 o_data_even_addr_gen_inst_U33 ( .A1(o_data_even_addr_gen_inst_N23), 
        .A2(o_data_even_addr_gen_inst_n33), .B1(o_data_even_addr_gen_inst_N13), 
        .B2(o_data_even_addr_gen_inst_n34), .ZN(o_data_even_addr_gen_inst_n40)
         );
  INV_X1 o_data_even_addr_gen_inst_U32 ( .A(o_data_even_addr_gen_inst_n40), 
        .ZN(o_data_even_addr_gen_inst_n23) );
  AOI22_X1 o_data_even_addr_gen_inst_U31 ( .A1(o_data_even_addr_gen_inst_N24), 
        .A2(o_data_even_addr_gen_inst_n33), .B1(o_data_even_addr_gen_inst_N14), 
        .B2(o_data_even_addr_gen_inst_n34), .ZN(o_data_even_addr_gen_inst_n39)
         );
  INV_X1 o_data_even_addr_gen_inst_U30 ( .A(o_data_even_addr_gen_inst_n39), 
        .ZN(o_data_even_addr_gen_inst_n22) );
  AOI22_X1 o_data_even_addr_gen_inst_U29 ( .A1(o_data_even_addr_gen_inst_N25), 
        .A2(o_data_even_addr_gen_inst_n33), .B1(o_data_even_addr_gen_inst_N15), 
        .B2(o_data_even_addr_gen_inst_n34), .ZN(o_data_even_addr_gen_inst_n38)
         );
  INV_X1 o_data_even_addr_gen_inst_U28 ( .A(o_data_even_addr_gen_inst_n38), 
        .ZN(o_data_even_addr_gen_inst_n21) );
  AOI22_X1 o_data_even_addr_gen_inst_U27 ( .A1(o_data_even_addr_gen_inst_N26), 
        .A2(o_data_even_addr_gen_inst_n33), .B1(o_data_even_addr_gen_inst_N16), 
        .B2(o_data_even_addr_gen_inst_n34), .ZN(o_data_even_addr_gen_inst_n37)
         );
  INV_X1 o_data_even_addr_gen_inst_U26 ( .A(o_data_even_addr_gen_inst_n37), 
        .ZN(o_data_even_addr_gen_inst_n20) );
  AOI22_X1 o_data_even_addr_gen_inst_U25 ( .A1(o_data_even_addr_gen_inst_N20), 
        .A2(o_data_even_addr_gen_inst_n33), .B1(o_data_even_addr_gen_inst_N10), 
        .B2(o_data_even_addr_gen_inst_n34), .ZN(o_data_even_addr_gen_inst_n43)
         );
  INV_X1 o_data_even_addr_gen_inst_U24 ( .A(o_data_even_addr_gen_inst_n43), 
        .ZN(o_data_even_addr_gen_inst_n26) );
  INV_X1 o_data_even_addr_gen_inst_U23 ( .A(int_c_o_en_base_odd), .ZN(
        o_data_even_addr_gen_inst_n28) );
  AOI22_X1 o_data_even_addr_gen_inst_U22 ( .A1(o_data_even_addr_gen_inst_N27), 
        .A2(o_data_even_addr_gen_inst_n33), .B1(o_data_even_addr_gen_inst_N17), 
        .B2(o_data_even_addr_gen_inst_n34), .ZN(o_data_even_addr_gen_inst_n36)
         );
  INV_X1 o_data_even_addr_gen_inst_U21 ( .A(o_data_even_addr_gen_inst_n36), 
        .ZN(o_data_even_addr_gen_inst_n18) );
  AOI22_X1 o_data_even_addr_gen_inst_U20 ( .A1(o_data_even_addr_gen_inst_N28), 
        .A2(o_data_even_addr_gen_inst_n33), .B1(o_data_even_addr_gen_inst_N18), 
        .B2(o_data_even_addr_gen_inst_n34), .ZN(o_data_even_addr_gen_inst_n35)
         );
  INV_X1 o_data_even_addr_gen_inst_U19 ( .A(o_data_even_addr_gen_inst_n35), 
        .ZN(o_data_even_addr_gen_inst_n8) );
  NOR2_X1 o_data_even_addr_gen_inst_U18 ( .A1(o_data_even_addr_gen_inst_n27), 
        .A2(1'b0), .ZN(o_data_even_addr_gen_inst_n34) );
  NOR2_X1 o_data_even_addr_gen_inst_U16 ( .A1(1'b0), .A2(1'b0), .ZN(
        o_data_even_addr_gen_inst_n33) );
  DFFR_X1 o_data_even_addr_gen_inst_int_base_addr_reg_4_ ( .D(
        o_data_even_addr_gen_inst_n22), .CK(o_data_even_addr_gen_inst_net2805), 
        .RN(o_data_even_addr_gen_inst_n6), .Q(
        o_data_even_addr_gen_inst_int_base_addr_4_) );
  DFFR_X1 o_data_even_addr_gen_inst_int_base_addr_reg_3_ ( .D(
        o_data_even_addr_gen_inst_n23), .CK(o_data_even_addr_gen_inst_net2805), 
        .RN(o_data_even_addr_gen_inst_n6), .Q(
        o_data_even_addr_gen_inst_int_base_addr_3_) );
  DFFR_X1 o_data_even_addr_gen_inst_int_base_addr_reg_2_ ( .D(
        o_data_even_addr_gen_inst_n24), .CK(o_data_even_addr_gen_inst_net2805), 
        .RN(o_data_even_addr_gen_inst_n6), .Q(
        o_data_even_addr_gen_inst_int_base_addr_2_) );
  DFFR_X1 o_data_even_addr_gen_inst_int_base_addr_reg_1_ ( .D(
        o_data_even_addr_gen_inst_n25), .CK(o_data_even_addr_gen_inst_net2805), 
        .RN(o_data_even_addr_gen_inst_n6), .Q(
        o_data_even_addr_gen_inst_int_base_addr_1_) );
  DFFR_X1 o_data_even_addr_gen_inst_int_base_addr_reg_0_ ( .D(
        o_data_even_addr_gen_inst_n26), .CK(o_data_even_addr_gen_inst_net2805), 
        .RN(o_data_even_addr_gen_inst_n6), .Q(
        o_data_even_addr_gen_inst_int_base_addr_0_) );
  DFFR_X1 o_data_even_addr_gen_inst_int_base_addr_reg_8_ ( .D(
        o_data_even_addr_gen_inst_n8), .CK(o_data_even_addr_gen_inst_net2805), 
        .RN(o_data_even_addr_gen_inst_n5), .Q(
        o_data_even_addr_gen_inst_int_base_addr_8_) );
  DFFR_X1 o_data_even_addr_gen_inst_int_base_addr_reg_7_ ( .D(
        o_data_even_addr_gen_inst_n18), .CK(o_data_even_addr_gen_inst_net2805), 
        .RN(o_data_even_addr_gen_inst_n5), .Q(
        o_data_even_addr_gen_inst_int_base_addr_7_) );
  DFFR_X1 o_data_even_addr_gen_inst_int_base_addr_reg_6_ ( .D(
        o_data_even_addr_gen_inst_n20), .CK(o_data_even_addr_gen_inst_net2805), 
        .RN(o_data_even_addr_gen_inst_n5), .Q(
        o_data_even_addr_gen_inst_int_base_addr_6_) );
  DFFR_X1 o_data_even_addr_gen_inst_int_base_addr_reg_5_ ( .D(
        o_data_even_addr_gen_inst_n21), .CK(o_data_even_addr_gen_inst_net2805), 
        .RN(o_data_even_addr_gen_inst_n5), .Q(
        o_data_even_addr_gen_inst_int_base_addr_5_) );
  DFFR_X1 o_data_even_addr_gen_inst_int_base_addr_reg_9_ ( .D(
        o_data_even_addr_gen_inst_n7), .CK(o_data_even_addr_gen_inst_net2805), 
        .RN(o_data_even_addr_gen_inst_n5), .Q(
        o_data_even_addr_gen_inst_int_base_addr_9_) );
  SDFFR_X1 o_data_even_addr_gen_inst_int_offs_addr_reg_9_ ( .D(1'b0), .SI(
        o_data_even_addr_gen_inst_n28), .SE(o_data_even_addr_gen_inst_N64), 
        .CK(o_data_even_addr_gen_inst_net2811), .RN(
        o_data_even_addr_gen_inst_n5), .Q(
        o_data_even_addr_gen_inst_int_offs_addr_9_) );
  SDFFR_X1 o_data_even_addr_gen_inst_int_offs_addr_reg_8_ ( .D(1'b0), .SI(
        o_data_even_addr_gen_inst_n28), .SE(o_data_even_addr_gen_inst_N63), 
        .CK(o_data_even_addr_gen_inst_net2811), .RN(
        o_data_even_addr_gen_inst_n5), .Q(
        o_data_even_addr_gen_inst_int_offs_addr_8_) );
  SDFFR_X1 o_data_even_addr_gen_inst_int_offs_addr_reg_7_ ( .D(1'b0), .SI(
        o_data_even_addr_gen_inst_n28), .SE(o_data_even_addr_gen_inst_N62), 
        .CK(o_data_even_addr_gen_inst_net2811), .RN(
        o_data_even_addr_gen_inst_n6), .Q(
        o_data_even_addr_gen_inst_int_offs_addr_7_) );
  SDFFR_X1 o_data_even_addr_gen_inst_int_offs_addr_reg_6_ ( .D(1'b0), .SI(
        o_data_even_addr_gen_inst_n28), .SE(o_data_even_addr_gen_inst_N61), 
        .CK(o_data_even_addr_gen_inst_net2811), .RN(
        o_data_even_addr_gen_inst_n6), .Q(
        o_data_even_addr_gen_inst_int_offs_addr_6_) );
  SDFFR_X1 o_data_even_addr_gen_inst_int_offs_addr_reg_5_ ( .D(1'b0), .SI(
        o_data_even_addr_gen_inst_n28), .SE(o_data_even_addr_gen_inst_N60), 
        .CK(o_data_even_addr_gen_inst_net2811), .RN(
        o_data_even_addr_gen_inst_n6), .Q(
        o_data_even_addr_gen_inst_int_offs_addr_5_) );
  SDFFR_X1 o_data_even_addr_gen_inst_int_offs_addr_reg_4_ ( .D(1'b0), .SI(
        o_data_even_addr_gen_inst_n28), .SE(o_data_even_addr_gen_inst_N59), 
        .CK(o_data_even_addr_gen_inst_net2811), .RN(
        o_data_even_addr_gen_inst_n6), .Q(
        o_data_even_addr_gen_inst_int_offs_addr_4_) );
  SDFFR_X1 o_data_even_addr_gen_inst_int_offs_addr_reg_3_ ( .D(1'b0), .SI(
        o_data_even_addr_gen_inst_n28), .SE(o_data_even_addr_gen_inst_N58), 
        .CK(o_data_even_addr_gen_inst_net2811), .RN(
        o_data_even_addr_gen_inst_n6), .Q(
        o_data_even_addr_gen_inst_int_offs_addr_3_) );
  SDFFR_X1 o_data_even_addr_gen_inst_int_offs_addr_reg_2_ ( .D(1'b0), .SI(
        o_data_even_addr_gen_inst_n28), .SE(o_data_even_addr_gen_inst_N57), 
        .CK(o_data_even_addr_gen_inst_net2811), .RN(
        o_data_even_addr_gen_inst_n6), .Q(
        o_data_even_addr_gen_inst_int_offs_addr_2_) );
  SDFFR_X1 o_data_even_addr_gen_inst_int_offs_addr_reg_1_ ( .D(1'b0), .SI(
        o_data_even_addr_gen_inst_n28), .SE(o_data_even_addr_gen_inst_N56), 
        .CK(o_data_even_addr_gen_inst_net2811), .RN(
        o_data_even_addr_gen_inst_n6), .Q(
        o_data_even_addr_gen_inst_int_offs_addr_1_) );
  SDFFR_X1 o_data_even_addr_gen_inst_int_offs_addr_reg_0_ ( .D(1'b0), .SI(
        o_data_even_addr_gen_inst_n28), .SE(o_data_even_addr_gen_inst_N55), 
        .CK(o_data_even_addr_gen_inst_net2811), .RN(
        o_data_even_addr_gen_inst_n6), .Q(
        o_data_even_addr_gen_inst_int_offs_addr_0_) );
  CLKGATETST_X1 o_data_even_addr_gen_inst_clk_gate_int_base_addr_reg_latch ( 
        .CK(ck), .E(o_data_even_addr_gen_inst_N40), .SE(1'b0), .GCK(
        o_data_even_addr_gen_inst_net2805) );
  CLKGATETST_X1 o_data_even_addr_gen_inst_clk_gate_int_offs_addr_reg_latch ( 
        .CK(ck), .E(o_data_even_addr_gen_inst_N65), .SE(1'b0), .GCK(
        o_data_even_addr_gen_inst_net2811) );
  XOR2_X1 o_data_even_addr_gen_inst_add_60_U2 ( .A(int_c_o_inc_value_offs[0]), 
        .B(o_data_even_addr_gen_inst_int_offs_addr_0_), .Z(
        o_data_even_addr_gen_inst_N55) );
  AND2_X1 o_data_even_addr_gen_inst_add_60_U1 ( .A1(int_c_o_inc_value_offs[0]), 
        .A2(o_data_even_addr_gen_inst_int_offs_addr_0_), .ZN(
        o_data_even_addr_gen_inst_add_60_n1) );
  FA_X1 o_data_even_addr_gen_inst_add_60_U1_1 ( .A(
        o_data_even_addr_gen_inst_int_offs_addr_1_), .B(
        int_c_o_inc_value_offs[1]), .CI(o_data_even_addr_gen_inst_add_60_n1), 
        .CO(o_data_even_addr_gen_inst_add_60_carry[2]), .S(
        o_data_even_addr_gen_inst_N56) );
  FA_X1 o_data_even_addr_gen_inst_add_60_U1_2 ( .A(
        o_data_even_addr_gen_inst_int_offs_addr_2_), .B(
        int_c_o_inc_value_offs[2]), .CI(
        o_data_even_addr_gen_inst_add_60_carry[2]), .CO(
        o_data_even_addr_gen_inst_add_60_carry[3]), .S(
        o_data_even_addr_gen_inst_N57) );
  FA_X1 o_data_even_addr_gen_inst_add_60_U1_3 ( .A(
        o_data_even_addr_gen_inst_int_offs_addr_3_), .B(
        int_c_o_inc_value_offs[3]), .CI(
        o_data_even_addr_gen_inst_add_60_carry[3]), .CO(
        o_data_even_addr_gen_inst_add_60_carry[4]), .S(
        o_data_even_addr_gen_inst_N58) );
  FA_X1 o_data_even_addr_gen_inst_add_60_U1_4 ( .A(
        o_data_even_addr_gen_inst_int_offs_addr_4_), .B(
        int_c_o_inc_value_offs[4]), .CI(
        o_data_even_addr_gen_inst_add_60_carry[4]), .CO(
        o_data_even_addr_gen_inst_add_60_carry[5]), .S(
        o_data_even_addr_gen_inst_N59) );
  FA_X1 o_data_even_addr_gen_inst_add_60_U1_5 ( .A(
        o_data_even_addr_gen_inst_int_offs_addr_5_), .B(1'b0), .CI(
        o_data_even_addr_gen_inst_add_60_carry[5]), .CO(
        o_data_even_addr_gen_inst_add_60_carry[6]), .S(
        o_data_even_addr_gen_inst_N60) );
  FA_X1 o_data_even_addr_gen_inst_add_60_U1_6 ( .A(
        o_data_even_addr_gen_inst_int_offs_addr_6_), .B(1'b0), .CI(
        o_data_even_addr_gen_inst_add_60_carry[6]), .CO(
        o_data_even_addr_gen_inst_add_60_carry[7]), .S(
        o_data_even_addr_gen_inst_N61) );
  FA_X1 o_data_even_addr_gen_inst_add_60_U1_7 ( .A(
        o_data_even_addr_gen_inst_int_offs_addr_7_), .B(1'b0), .CI(
        o_data_even_addr_gen_inst_add_60_carry[7]), .CO(
        o_data_even_addr_gen_inst_add_60_carry[8]), .S(
        o_data_even_addr_gen_inst_N62) );
  FA_X1 o_data_even_addr_gen_inst_add_60_U1_8 ( .A(
        o_data_even_addr_gen_inst_int_offs_addr_8_), .B(1'b0), .CI(
        o_data_even_addr_gen_inst_add_60_carry[8]), .CO(
        o_data_even_addr_gen_inst_add_60_carry[9]), .S(
        o_data_even_addr_gen_inst_N63) );
  FA_X1 o_data_even_addr_gen_inst_add_60_U1_9 ( .A(
        o_data_even_addr_gen_inst_int_offs_addr_9_), .B(1'b0), .CI(
        o_data_even_addr_gen_inst_add_60_carry[9]), .S(
        o_data_even_addr_gen_inst_N64) );
  AND2_X1 o_data_even_addr_gen_inst_add_45_U2 ( .A1(1'b1), .A2(
        o_data_even_addr_gen_inst_int_base_addr_0_), .ZN(
        o_data_even_addr_gen_inst_add_45_n2) );
  XOR2_X1 o_data_even_addr_gen_inst_add_45_U1 ( .A(1'b1), .B(
        o_data_even_addr_gen_inst_int_base_addr_0_), .Z(
        o_data_even_addr_gen_inst_N20) );
  FA_X1 o_data_even_addr_gen_inst_add_45_U1_1 ( .A(
        o_data_even_addr_gen_inst_int_base_addr_1_), .B(1'b0), .CI(
        o_data_even_addr_gen_inst_add_45_n2), .CO(
        o_data_even_addr_gen_inst_add_45_carry[2]), .S(
        o_data_even_addr_gen_inst_N21) );
  FA_X1 o_data_even_addr_gen_inst_add_45_U1_2 ( .A(
        o_data_even_addr_gen_inst_int_base_addr_2_), .B(1'b0), .CI(
        o_data_even_addr_gen_inst_add_45_carry[2]), .CO(
        o_data_even_addr_gen_inst_add_45_carry[3]), .S(
        o_data_even_addr_gen_inst_N22) );
  FA_X1 o_data_even_addr_gen_inst_add_45_U1_3 ( .A(
        o_data_even_addr_gen_inst_int_base_addr_3_), .B(1'b0), .CI(
        o_data_even_addr_gen_inst_add_45_carry[3]), .CO(
        o_data_even_addr_gen_inst_add_45_carry[4]), .S(
        o_data_even_addr_gen_inst_N23) );
  FA_X1 o_data_even_addr_gen_inst_add_45_U1_4 ( .A(
        o_data_even_addr_gen_inst_int_base_addr_4_), .B(1'b0), .CI(
        o_data_even_addr_gen_inst_add_45_carry[4]), .CO(
        o_data_even_addr_gen_inst_add_45_carry[5]), .S(
        o_data_even_addr_gen_inst_N24) );
  FA_X1 o_data_even_addr_gen_inst_add_45_U1_5 ( .A(
        o_data_even_addr_gen_inst_int_base_addr_5_), .B(1'b0), .CI(
        o_data_even_addr_gen_inst_add_45_carry[5]), .CO(
        o_data_even_addr_gen_inst_add_45_carry[6]), .S(
        o_data_even_addr_gen_inst_N25) );
  FA_X1 o_data_even_addr_gen_inst_add_45_U1_6 ( .A(
        o_data_even_addr_gen_inst_int_base_addr_6_), .B(1'b0), .CI(
        o_data_even_addr_gen_inst_add_45_carry[6]), .CO(
        o_data_even_addr_gen_inst_add_45_carry[7]), .S(
        o_data_even_addr_gen_inst_N26) );
  FA_X1 o_data_even_addr_gen_inst_add_45_U1_7 ( .A(
        o_data_even_addr_gen_inst_int_base_addr_7_), .B(1'b0), .CI(
        o_data_even_addr_gen_inst_add_45_carry[7]), .CO(
        o_data_even_addr_gen_inst_add_45_carry[8]), .S(
        o_data_even_addr_gen_inst_N27) );
  FA_X1 o_data_even_addr_gen_inst_add_45_U1_8 ( .A(
        o_data_even_addr_gen_inst_int_base_addr_8_), .B(1'b0), .CI(
        o_data_even_addr_gen_inst_add_45_carry[8]), .CO(
        o_data_even_addr_gen_inst_add_45_carry[9]), .S(
        o_data_even_addr_gen_inst_N28) );
  FA_X1 o_data_even_addr_gen_inst_add_45_U1_9 ( .A(
        o_data_even_addr_gen_inst_int_base_addr_9_), .B(1'b0), .CI(
        o_data_even_addr_gen_inst_add_45_carry[9]), .S(
        o_data_even_addr_gen_inst_N29) );
  AND2_X1 o_data_even_addr_gen_inst_add_43_U2 ( .A1(1'b1), .A2(
        o_data_even_addr[0]), .ZN(o_data_even_addr_gen_inst_add_43_n2) );
  XOR2_X1 o_data_even_addr_gen_inst_add_43_U1 ( .A(1'b1), .B(
        o_data_even_addr[0]), .Z(o_data_even_addr_gen_inst_N10) );
  FA_X1 o_data_even_addr_gen_inst_add_43_U1_1 ( .A(o_data_even_addr[1]), .B(
        1'b0), .CI(o_data_even_addr_gen_inst_add_43_n2), .CO(
        o_data_even_addr_gen_inst_add_43_carry[2]), .S(
        o_data_even_addr_gen_inst_N11) );
  FA_X1 o_data_even_addr_gen_inst_add_43_U1_2 ( .A(o_data_even_addr[2]), .B(
        1'b0), .CI(o_data_even_addr_gen_inst_add_43_carry[2]), .CO(
        o_data_even_addr_gen_inst_add_43_carry[3]), .S(
        o_data_even_addr_gen_inst_N12) );
  FA_X1 o_data_even_addr_gen_inst_add_43_U1_3 ( .A(o_data_even_addr[3]), .B(
        1'b0), .CI(o_data_even_addr_gen_inst_add_43_carry[3]), .CO(
        o_data_even_addr_gen_inst_add_43_carry[4]), .S(
        o_data_even_addr_gen_inst_N13) );
  FA_X1 o_data_even_addr_gen_inst_add_43_U1_4 ( .A(o_data_even_addr[4]), .B(
        1'b0), .CI(o_data_even_addr_gen_inst_add_43_carry[4]), .CO(
        o_data_even_addr_gen_inst_add_43_carry[5]), .S(
        o_data_even_addr_gen_inst_N14) );
  FA_X1 o_data_even_addr_gen_inst_add_43_U1_5 ( .A(o_data_even_addr[5]), .B(
        1'b0), .CI(o_data_even_addr_gen_inst_add_43_carry[5]), .CO(
        o_data_even_addr_gen_inst_add_43_carry[6]), .S(
        o_data_even_addr_gen_inst_N15) );
  FA_X1 o_data_even_addr_gen_inst_add_43_U1_6 ( .A(o_data_even_addr[6]), .B(
        1'b0), .CI(o_data_even_addr_gen_inst_add_43_carry[6]), .CO(
        o_data_even_addr_gen_inst_add_43_carry[7]), .S(
        o_data_even_addr_gen_inst_N16) );
  FA_X1 o_data_even_addr_gen_inst_add_43_U1_7 ( .A(o_data_even_addr[7]), .B(
        1'b0), .CI(o_data_even_addr_gen_inst_add_43_carry[7]), .CO(
        o_data_even_addr_gen_inst_add_43_carry[8]), .S(
        o_data_even_addr_gen_inst_N17) );
  FA_X1 o_data_even_addr_gen_inst_add_43_U1_8 ( .A(o_data_even_addr[8]), .B(
        1'b0), .CI(o_data_even_addr_gen_inst_add_43_carry[8]), .CO(
        o_data_even_addr_gen_inst_add_43_carry[9]), .S(
        o_data_even_addr_gen_inst_N18) );
  FA_X1 o_data_even_addr_gen_inst_add_43_U1_9 ( .A(o_data_even_addr[9]), .B(
        1'b0), .CI(o_data_even_addr_gen_inst_add_43_carry[9]), .S(
        o_data_even_addr_gen_inst_N19) );
  XOR2_X1 o_data_even_addr_gen_inst_add_31_U2 ( .A(
        o_data_even_addr_gen_inst_int_offs_addr_0_), .B(
        o_data_even_addr_gen_inst_int_base_addr_0_), .Z(o_data_even_addr[0])
         );
  AND2_X1 o_data_even_addr_gen_inst_add_31_U1 ( .A1(
        o_data_even_addr_gen_inst_int_offs_addr_0_), .A2(
        o_data_even_addr_gen_inst_int_base_addr_0_), .ZN(
        o_data_even_addr_gen_inst_add_31_n1) );
  FA_X1 o_data_even_addr_gen_inst_add_31_U1_1 ( .A(
        o_data_even_addr_gen_inst_int_base_addr_1_), .B(
        o_data_even_addr_gen_inst_int_offs_addr_1_), .CI(
        o_data_even_addr_gen_inst_add_31_n1), .CO(
        o_data_even_addr_gen_inst_add_31_carry[2]), .S(o_data_even_addr[1]) );
  FA_X1 o_data_even_addr_gen_inst_add_31_U1_2 ( .A(
        o_data_even_addr_gen_inst_int_base_addr_2_), .B(
        o_data_even_addr_gen_inst_int_offs_addr_2_), .CI(
        o_data_even_addr_gen_inst_add_31_carry[2]), .CO(
        o_data_even_addr_gen_inst_add_31_carry[3]), .S(o_data_even_addr[2]) );
  FA_X1 o_data_even_addr_gen_inst_add_31_U1_3 ( .A(
        o_data_even_addr_gen_inst_int_base_addr_3_), .B(
        o_data_even_addr_gen_inst_int_offs_addr_3_), .CI(
        o_data_even_addr_gen_inst_add_31_carry[3]), .CO(
        o_data_even_addr_gen_inst_add_31_carry[4]), .S(o_data_even_addr[3]) );
  FA_X1 o_data_even_addr_gen_inst_add_31_U1_4 ( .A(
        o_data_even_addr_gen_inst_int_base_addr_4_), .B(
        o_data_even_addr_gen_inst_int_offs_addr_4_), .CI(
        o_data_even_addr_gen_inst_add_31_carry[4]), .CO(
        o_data_even_addr_gen_inst_add_31_carry[5]), .S(o_data_even_addr[4]) );
  FA_X1 o_data_even_addr_gen_inst_add_31_U1_5 ( .A(
        o_data_even_addr_gen_inst_int_base_addr_5_), .B(
        o_data_even_addr_gen_inst_int_offs_addr_5_), .CI(
        o_data_even_addr_gen_inst_add_31_carry[5]), .CO(
        o_data_even_addr_gen_inst_add_31_carry[6]), .S(o_data_even_addr[5]) );
  FA_X1 o_data_even_addr_gen_inst_add_31_U1_6 ( .A(
        o_data_even_addr_gen_inst_int_base_addr_6_), .B(
        o_data_even_addr_gen_inst_int_offs_addr_6_), .CI(
        o_data_even_addr_gen_inst_add_31_carry[6]), .CO(
        o_data_even_addr_gen_inst_add_31_carry[7]), .S(o_data_even_addr[6]) );
  FA_X1 o_data_even_addr_gen_inst_add_31_U1_7 ( .A(
        o_data_even_addr_gen_inst_int_base_addr_7_), .B(
        o_data_even_addr_gen_inst_int_offs_addr_7_), .CI(
        o_data_even_addr_gen_inst_add_31_carry[7]), .CO(
        o_data_even_addr_gen_inst_add_31_carry[8]), .S(o_data_even_addr[7]) );
  FA_X1 o_data_even_addr_gen_inst_add_31_U1_8 ( .A(
        o_data_even_addr_gen_inst_int_base_addr_8_), .B(
        o_data_even_addr_gen_inst_int_offs_addr_8_), .CI(
        o_data_even_addr_gen_inst_add_31_carry[8]), .CO(
        o_data_even_addr_gen_inst_add_31_carry[9]), .S(o_data_even_addr[8]) );
  FA_X1 o_data_even_addr_gen_inst_add_31_U1_9 ( .A(
        o_data_even_addr_gen_inst_int_base_addr_9_), .B(
        o_data_even_addr_gen_inst_int_offs_addr_9_), .CI(
        o_data_even_addr_gen_inst_add_31_carry[9]), .S(o_data_even_addr[9]) );
  INV_X1 o_data_odd_addr_gen_inst_U44 ( .A(rst), .ZN(
        o_data_odd_addr_gen_inst_n6) );
  INV_X1 o_data_odd_addr_gen_inst_U43 ( .A(rst), .ZN(
        o_data_odd_addr_gen_inst_n5) );
  INV_X1 o_data_odd_addr_gen_inst_U42 ( .A(1'b0), .ZN(
        o_data_odd_addr_gen_inst_n27) );
  OR2_X1 o_data_odd_addr_gen_inst_U41 ( .A1(int_c_o_en_base_odd), .A2(1'b0), 
        .ZN(o_data_odd_addr_gen_inst_N40) );
  OR2_X1 o_data_odd_addr_gen_inst_U40 ( .A1(int_c_o_en_base_odd), .A2(
        int_c_o_en_offs_odd), .ZN(o_data_odd_addr_gen_inst_N65) );
  AOI22_X1 o_data_odd_addr_gen_inst_U39 ( .A1(o_data_odd_addr_gen_inst_N29), 
        .A2(o_data_odd_addr_gen_inst_n33), .B1(o_data_odd_addr_gen_inst_N19), 
        .B2(o_data_odd_addr_gen_inst_n34), .ZN(o_data_odd_addr_gen_inst_n32)
         );
  INV_X1 o_data_odd_addr_gen_inst_U38 ( .A(o_data_odd_addr_gen_inst_n32), .ZN(
        o_data_odd_addr_gen_inst_n7) );
  AOI22_X1 o_data_odd_addr_gen_inst_U37 ( .A1(o_data_odd_addr_gen_inst_N21), 
        .A2(o_data_odd_addr_gen_inst_n33), .B1(o_data_odd_addr_gen_inst_N11), 
        .B2(o_data_odd_addr_gen_inst_n34), .ZN(o_data_odd_addr_gen_inst_n42)
         );
  INV_X1 o_data_odd_addr_gen_inst_U36 ( .A(o_data_odd_addr_gen_inst_n42), .ZN(
        o_data_odd_addr_gen_inst_n25) );
  AOI22_X1 o_data_odd_addr_gen_inst_U35 ( .A1(o_data_odd_addr_gen_inst_N22), 
        .A2(o_data_odd_addr_gen_inst_n33), .B1(o_data_odd_addr_gen_inst_N12), 
        .B2(o_data_odd_addr_gen_inst_n34), .ZN(o_data_odd_addr_gen_inst_n41)
         );
  INV_X1 o_data_odd_addr_gen_inst_U34 ( .A(o_data_odd_addr_gen_inst_n41), .ZN(
        o_data_odd_addr_gen_inst_n24) );
  AOI22_X1 o_data_odd_addr_gen_inst_U33 ( .A1(o_data_odd_addr_gen_inst_N23), 
        .A2(o_data_odd_addr_gen_inst_n33), .B1(o_data_odd_addr_gen_inst_N13), 
        .B2(o_data_odd_addr_gen_inst_n34), .ZN(o_data_odd_addr_gen_inst_n40)
         );
  INV_X1 o_data_odd_addr_gen_inst_U32 ( .A(o_data_odd_addr_gen_inst_n40), .ZN(
        o_data_odd_addr_gen_inst_n23) );
  AOI22_X1 o_data_odd_addr_gen_inst_U31 ( .A1(o_data_odd_addr_gen_inst_N24), 
        .A2(o_data_odd_addr_gen_inst_n33), .B1(o_data_odd_addr_gen_inst_N14), 
        .B2(o_data_odd_addr_gen_inst_n34), .ZN(o_data_odd_addr_gen_inst_n39)
         );
  INV_X1 o_data_odd_addr_gen_inst_U30 ( .A(o_data_odd_addr_gen_inst_n39), .ZN(
        o_data_odd_addr_gen_inst_n22) );
  AOI22_X1 o_data_odd_addr_gen_inst_U29 ( .A1(o_data_odd_addr_gen_inst_N25), 
        .A2(o_data_odd_addr_gen_inst_n33), .B1(o_data_odd_addr_gen_inst_N15), 
        .B2(o_data_odd_addr_gen_inst_n34), .ZN(o_data_odd_addr_gen_inst_n38)
         );
  INV_X1 o_data_odd_addr_gen_inst_U28 ( .A(o_data_odd_addr_gen_inst_n38), .ZN(
        o_data_odd_addr_gen_inst_n21) );
  AOI22_X1 o_data_odd_addr_gen_inst_U27 ( .A1(o_data_odd_addr_gen_inst_N26), 
        .A2(o_data_odd_addr_gen_inst_n33), .B1(o_data_odd_addr_gen_inst_N16), 
        .B2(o_data_odd_addr_gen_inst_n34), .ZN(o_data_odd_addr_gen_inst_n37)
         );
  INV_X1 o_data_odd_addr_gen_inst_U26 ( .A(o_data_odd_addr_gen_inst_n37), .ZN(
        o_data_odd_addr_gen_inst_n20) );
  AOI22_X1 o_data_odd_addr_gen_inst_U25 ( .A1(o_data_odd_addr_gen_inst_N20), 
        .A2(o_data_odd_addr_gen_inst_n33), .B1(o_data_odd_addr_gen_inst_N10), 
        .B2(o_data_odd_addr_gen_inst_n34), .ZN(o_data_odd_addr_gen_inst_n43)
         );
  INV_X1 o_data_odd_addr_gen_inst_U24 ( .A(o_data_odd_addr_gen_inst_n43), .ZN(
        o_data_odd_addr_gen_inst_n26) );
  INV_X1 o_data_odd_addr_gen_inst_U23 ( .A(int_c_o_en_base_odd), .ZN(
        o_data_odd_addr_gen_inst_n28) );
  AOI22_X1 o_data_odd_addr_gen_inst_U22 ( .A1(o_data_odd_addr_gen_inst_N27), 
        .A2(o_data_odd_addr_gen_inst_n33), .B1(o_data_odd_addr_gen_inst_N17), 
        .B2(o_data_odd_addr_gen_inst_n34), .ZN(o_data_odd_addr_gen_inst_n36)
         );
  INV_X1 o_data_odd_addr_gen_inst_U21 ( .A(o_data_odd_addr_gen_inst_n36), .ZN(
        o_data_odd_addr_gen_inst_n18) );
  AOI22_X1 o_data_odd_addr_gen_inst_U20 ( .A1(o_data_odd_addr_gen_inst_N28), 
        .A2(o_data_odd_addr_gen_inst_n33), .B1(o_data_odd_addr_gen_inst_N18), 
        .B2(o_data_odd_addr_gen_inst_n34), .ZN(o_data_odd_addr_gen_inst_n35)
         );
  INV_X1 o_data_odd_addr_gen_inst_U19 ( .A(o_data_odd_addr_gen_inst_n35), .ZN(
        o_data_odd_addr_gen_inst_n8) );
  NOR2_X1 o_data_odd_addr_gen_inst_U18 ( .A1(o_data_odd_addr_gen_inst_n27), 
        .A2(1'b0), .ZN(o_data_odd_addr_gen_inst_n34) );
  NOR2_X1 o_data_odd_addr_gen_inst_U16 ( .A1(1'b0), .A2(1'b0), .ZN(
        o_data_odd_addr_gen_inst_n33) );
  DFFR_X1 o_data_odd_addr_gen_inst_int_base_addr_reg_4_ ( .D(
        o_data_odd_addr_gen_inst_n22), .CK(o_data_odd_addr_gen_inst_net2782), 
        .RN(o_data_odd_addr_gen_inst_n6), .Q(
        o_data_odd_addr_gen_inst_int_base_addr_4_) );
  DFFR_X1 o_data_odd_addr_gen_inst_int_base_addr_reg_3_ ( .D(
        o_data_odd_addr_gen_inst_n23), .CK(o_data_odd_addr_gen_inst_net2782), 
        .RN(o_data_odd_addr_gen_inst_n6), .Q(
        o_data_odd_addr_gen_inst_int_base_addr_3_) );
  DFFR_X1 o_data_odd_addr_gen_inst_int_base_addr_reg_2_ ( .D(
        o_data_odd_addr_gen_inst_n24), .CK(o_data_odd_addr_gen_inst_net2782), 
        .RN(o_data_odd_addr_gen_inst_n6), .Q(
        o_data_odd_addr_gen_inst_int_base_addr_2_) );
  DFFR_X1 o_data_odd_addr_gen_inst_int_base_addr_reg_1_ ( .D(
        o_data_odd_addr_gen_inst_n25), .CK(o_data_odd_addr_gen_inst_net2782), 
        .RN(o_data_odd_addr_gen_inst_n6), .Q(
        o_data_odd_addr_gen_inst_int_base_addr_1_) );
  DFFR_X1 o_data_odd_addr_gen_inst_int_base_addr_reg_0_ ( .D(
        o_data_odd_addr_gen_inst_n26), .CK(o_data_odd_addr_gen_inst_net2782), 
        .RN(o_data_odd_addr_gen_inst_n6), .Q(
        o_data_odd_addr_gen_inst_int_base_addr_0_) );
  DFFR_X1 o_data_odd_addr_gen_inst_int_base_addr_reg_8_ ( .D(
        o_data_odd_addr_gen_inst_n8), .CK(o_data_odd_addr_gen_inst_net2782), 
        .RN(o_data_odd_addr_gen_inst_n5), .Q(
        o_data_odd_addr_gen_inst_int_base_addr_8_) );
  DFFR_X1 o_data_odd_addr_gen_inst_int_base_addr_reg_7_ ( .D(
        o_data_odd_addr_gen_inst_n18), .CK(o_data_odd_addr_gen_inst_net2782), 
        .RN(o_data_odd_addr_gen_inst_n5), .Q(
        o_data_odd_addr_gen_inst_int_base_addr_7_) );
  DFFR_X1 o_data_odd_addr_gen_inst_int_base_addr_reg_6_ ( .D(
        o_data_odd_addr_gen_inst_n20), .CK(o_data_odd_addr_gen_inst_net2782), 
        .RN(o_data_odd_addr_gen_inst_n5), .Q(
        o_data_odd_addr_gen_inst_int_base_addr_6_) );
  DFFR_X1 o_data_odd_addr_gen_inst_int_base_addr_reg_5_ ( .D(
        o_data_odd_addr_gen_inst_n21), .CK(o_data_odd_addr_gen_inst_net2782), 
        .RN(o_data_odd_addr_gen_inst_n5), .Q(
        o_data_odd_addr_gen_inst_int_base_addr_5_) );
  DFFR_X1 o_data_odd_addr_gen_inst_int_base_addr_reg_9_ ( .D(
        o_data_odd_addr_gen_inst_n7), .CK(o_data_odd_addr_gen_inst_net2782), 
        .RN(o_data_odd_addr_gen_inst_n5), .Q(
        o_data_odd_addr_gen_inst_int_base_addr_9_) );
  SDFFR_X1 o_data_odd_addr_gen_inst_int_offs_addr_reg_9_ ( .D(1'b0), .SI(
        o_data_odd_addr_gen_inst_n28), .SE(o_data_odd_addr_gen_inst_N64), .CK(
        o_data_odd_addr_gen_inst_net2788), .RN(o_data_odd_addr_gen_inst_n5), 
        .Q(o_data_odd_addr_gen_inst_int_offs_addr_9_) );
  SDFFR_X1 o_data_odd_addr_gen_inst_int_offs_addr_reg_8_ ( .D(1'b0), .SI(
        o_data_odd_addr_gen_inst_n28), .SE(o_data_odd_addr_gen_inst_N63), .CK(
        o_data_odd_addr_gen_inst_net2788), .RN(o_data_odd_addr_gen_inst_n5), 
        .Q(o_data_odd_addr_gen_inst_int_offs_addr_8_) );
  SDFFR_X1 o_data_odd_addr_gen_inst_int_offs_addr_reg_7_ ( .D(1'b0), .SI(
        o_data_odd_addr_gen_inst_n28), .SE(o_data_odd_addr_gen_inst_N62), .CK(
        o_data_odd_addr_gen_inst_net2788), .RN(o_data_odd_addr_gen_inst_n6), 
        .Q(o_data_odd_addr_gen_inst_int_offs_addr_7_) );
  SDFFR_X1 o_data_odd_addr_gen_inst_int_offs_addr_reg_6_ ( .D(1'b0), .SI(
        o_data_odd_addr_gen_inst_n28), .SE(o_data_odd_addr_gen_inst_N61), .CK(
        o_data_odd_addr_gen_inst_net2788), .RN(o_data_odd_addr_gen_inst_n6), 
        .Q(o_data_odd_addr_gen_inst_int_offs_addr_6_) );
  SDFFR_X1 o_data_odd_addr_gen_inst_int_offs_addr_reg_5_ ( .D(1'b0), .SI(
        o_data_odd_addr_gen_inst_n28), .SE(o_data_odd_addr_gen_inst_N60), .CK(
        o_data_odd_addr_gen_inst_net2788), .RN(o_data_odd_addr_gen_inst_n6), 
        .Q(o_data_odd_addr_gen_inst_int_offs_addr_5_) );
  SDFFR_X1 o_data_odd_addr_gen_inst_int_offs_addr_reg_4_ ( .D(1'b0), .SI(
        o_data_odd_addr_gen_inst_n28), .SE(o_data_odd_addr_gen_inst_N59), .CK(
        o_data_odd_addr_gen_inst_net2788), .RN(o_data_odd_addr_gen_inst_n6), 
        .Q(o_data_odd_addr_gen_inst_int_offs_addr_4_) );
  SDFFR_X1 o_data_odd_addr_gen_inst_int_offs_addr_reg_3_ ( .D(1'b0), .SI(
        o_data_odd_addr_gen_inst_n28), .SE(o_data_odd_addr_gen_inst_N58), .CK(
        o_data_odd_addr_gen_inst_net2788), .RN(o_data_odd_addr_gen_inst_n6), 
        .Q(o_data_odd_addr_gen_inst_int_offs_addr_3_) );
  SDFFR_X1 o_data_odd_addr_gen_inst_int_offs_addr_reg_2_ ( .D(1'b0), .SI(
        o_data_odd_addr_gen_inst_n28), .SE(o_data_odd_addr_gen_inst_N57), .CK(
        o_data_odd_addr_gen_inst_net2788), .RN(o_data_odd_addr_gen_inst_n6), 
        .Q(o_data_odd_addr_gen_inst_int_offs_addr_2_) );
  SDFFR_X1 o_data_odd_addr_gen_inst_int_offs_addr_reg_1_ ( .D(1'b0), .SI(
        o_data_odd_addr_gen_inst_n28), .SE(o_data_odd_addr_gen_inst_N56), .CK(
        o_data_odd_addr_gen_inst_net2788), .RN(o_data_odd_addr_gen_inst_n6), 
        .Q(o_data_odd_addr_gen_inst_int_offs_addr_1_) );
  SDFFR_X1 o_data_odd_addr_gen_inst_int_offs_addr_reg_0_ ( .D(1'b0), .SI(
        o_data_odd_addr_gen_inst_n28), .SE(o_data_odd_addr_gen_inst_N55), .CK(
        o_data_odd_addr_gen_inst_net2788), .RN(o_data_odd_addr_gen_inst_n6), 
        .Q(o_data_odd_addr_gen_inst_int_offs_addr_0_) );
  CLKGATETST_X1 o_data_odd_addr_gen_inst_clk_gate_int_base_addr_reg_latch ( 
        .CK(ck), .E(o_data_odd_addr_gen_inst_N40), .SE(1'b0), .GCK(
        o_data_odd_addr_gen_inst_net2782) );
  CLKGATETST_X1 o_data_odd_addr_gen_inst_clk_gate_int_offs_addr_reg_latch ( 
        .CK(ck), .E(o_data_odd_addr_gen_inst_N65), .SE(1'b0), .GCK(
        o_data_odd_addr_gen_inst_net2788) );
  XOR2_X1 o_data_odd_addr_gen_inst_add_60_U2 ( .A(int_c_o_inc_value_offs[0]), 
        .B(o_data_odd_addr_gen_inst_int_offs_addr_0_), .Z(
        o_data_odd_addr_gen_inst_N55) );
  AND2_X1 o_data_odd_addr_gen_inst_add_60_U1 ( .A1(int_c_o_inc_value_offs[0]), 
        .A2(o_data_odd_addr_gen_inst_int_offs_addr_0_), .ZN(
        o_data_odd_addr_gen_inst_add_60_n1) );
  FA_X1 o_data_odd_addr_gen_inst_add_60_U1_1 ( .A(
        o_data_odd_addr_gen_inst_int_offs_addr_1_), .B(
        int_c_o_inc_value_offs[1]), .CI(o_data_odd_addr_gen_inst_add_60_n1), 
        .CO(o_data_odd_addr_gen_inst_add_60_carry[2]), .S(
        o_data_odd_addr_gen_inst_N56) );
  FA_X1 o_data_odd_addr_gen_inst_add_60_U1_2 ( .A(
        o_data_odd_addr_gen_inst_int_offs_addr_2_), .B(
        int_c_o_inc_value_offs[2]), .CI(
        o_data_odd_addr_gen_inst_add_60_carry[2]), .CO(
        o_data_odd_addr_gen_inst_add_60_carry[3]), .S(
        o_data_odd_addr_gen_inst_N57) );
  FA_X1 o_data_odd_addr_gen_inst_add_60_U1_3 ( .A(
        o_data_odd_addr_gen_inst_int_offs_addr_3_), .B(
        int_c_o_inc_value_offs[3]), .CI(
        o_data_odd_addr_gen_inst_add_60_carry[3]), .CO(
        o_data_odd_addr_gen_inst_add_60_carry[4]), .S(
        o_data_odd_addr_gen_inst_N58) );
  FA_X1 o_data_odd_addr_gen_inst_add_60_U1_4 ( .A(
        o_data_odd_addr_gen_inst_int_offs_addr_4_), .B(
        int_c_o_inc_value_offs[4]), .CI(
        o_data_odd_addr_gen_inst_add_60_carry[4]), .CO(
        o_data_odd_addr_gen_inst_add_60_carry[5]), .S(
        o_data_odd_addr_gen_inst_N59) );
  FA_X1 o_data_odd_addr_gen_inst_add_60_U1_5 ( .A(
        o_data_odd_addr_gen_inst_int_offs_addr_5_), .B(1'b0), .CI(
        o_data_odd_addr_gen_inst_add_60_carry[5]), .CO(
        o_data_odd_addr_gen_inst_add_60_carry[6]), .S(
        o_data_odd_addr_gen_inst_N60) );
  FA_X1 o_data_odd_addr_gen_inst_add_60_U1_6 ( .A(
        o_data_odd_addr_gen_inst_int_offs_addr_6_), .B(1'b0), .CI(
        o_data_odd_addr_gen_inst_add_60_carry[6]), .CO(
        o_data_odd_addr_gen_inst_add_60_carry[7]), .S(
        o_data_odd_addr_gen_inst_N61) );
  FA_X1 o_data_odd_addr_gen_inst_add_60_U1_7 ( .A(
        o_data_odd_addr_gen_inst_int_offs_addr_7_), .B(1'b0), .CI(
        o_data_odd_addr_gen_inst_add_60_carry[7]), .CO(
        o_data_odd_addr_gen_inst_add_60_carry[8]), .S(
        o_data_odd_addr_gen_inst_N62) );
  FA_X1 o_data_odd_addr_gen_inst_add_60_U1_8 ( .A(
        o_data_odd_addr_gen_inst_int_offs_addr_8_), .B(1'b0), .CI(
        o_data_odd_addr_gen_inst_add_60_carry[8]), .CO(
        o_data_odd_addr_gen_inst_add_60_carry[9]), .S(
        o_data_odd_addr_gen_inst_N63) );
  FA_X1 o_data_odd_addr_gen_inst_add_60_U1_9 ( .A(
        o_data_odd_addr_gen_inst_int_offs_addr_9_), .B(1'b0), .CI(
        o_data_odd_addr_gen_inst_add_60_carry[9]), .S(
        o_data_odd_addr_gen_inst_N64) );
  AND2_X1 o_data_odd_addr_gen_inst_add_45_U2 ( .A1(1'b1), .A2(
        o_data_odd_addr_gen_inst_int_base_addr_0_), .ZN(
        o_data_odd_addr_gen_inst_add_45_n2) );
  XOR2_X1 o_data_odd_addr_gen_inst_add_45_U1 ( .A(1'b1), .B(
        o_data_odd_addr_gen_inst_int_base_addr_0_), .Z(
        o_data_odd_addr_gen_inst_N20) );
  FA_X1 o_data_odd_addr_gen_inst_add_45_U1_1 ( .A(
        o_data_odd_addr_gen_inst_int_base_addr_1_), .B(1'b0), .CI(
        o_data_odd_addr_gen_inst_add_45_n2), .CO(
        o_data_odd_addr_gen_inst_add_45_carry[2]), .S(
        o_data_odd_addr_gen_inst_N21) );
  FA_X1 o_data_odd_addr_gen_inst_add_45_U1_2 ( .A(
        o_data_odd_addr_gen_inst_int_base_addr_2_), .B(1'b0), .CI(
        o_data_odd_addr_gen_inst_add_45_carry[2]), .CO(
        o_data_odd_addr_gen_inst_add_45_carry[3]), .S(
        o_data_odd_addr_gen_inst_N22) );
  FA_X1 o_data_odd_addr_gen_inst_add_45_U1_3 ( .A(
        o_data_odd_addr_gen_inst_int_base_addr_3_), .B(1'b0), .CI(
        o_data_odd_addr_gen_inst_add_45_carry[3]), .CO(
        o_data_odd_addr_gen_inst_add_45_carry[4]), .S(
        o_data_odd_addr_gen_inst_N23) );
  FA_X1 o_data_odd_addr_gen_inst_add_45_U1_4 ( .A(
        o_data_odd_addr_gen_inst_int_base_addr_4_), .B(1'b0), .CI(
        o_data_odd_addr_gen_inst_add_45_carry[4]), .CO(
        o_data_odd_addr_gen_inst_add_45_carry[5]), .S(
        o_data_odd_addr_gen_inst_N24) );
  FA_X1 o_data_odd_addr_gen_inst_add_45_U1_5 ( .A(
        o_data_odd_addr_gen_inst_int_base_addr_5_), .B(1'b0), .CI(
        o_data_odd_addr_gen_inst_add_45_carry[5]), .CO(
        o_data_odd_addr_gen_inst_add_45_carry[6]), .S(
        o_data_odd_addr_gen_inst_N25) );
  FA_X1 o_data_odd_addr_gen_inst_add_45_U1_6 ( .A(
        o_data_odd_addr_gen_inst_int_base_addr_6_), .B(1'b0), .CI(
        o_data_odd_addr_gen_inst_add_45_carry[6]), .CO(
        o_data_odd_addr_gen_inst_add_45_carry[7]), .S(
        o_data_odd_addr_gen_inst_N26) );
  FA_X1 o_data_odd_addr_gen_inst_add_45_U1_7 ( .A(
        o_data_odd_addr_gen_inst_int_base_addr_7_), .B(1'b0), .CI(
        o_data_odd_addr_gen_inst_add_45_carry[7]), .CO(
        o_data_odd_addr_gen_inst_add_45_carry[8]), .S(
        o_data_odd_addr_gen_inst_N27) );
  FA_X1 o_data_odd_addr_gen_inst_add_45_U1_8 ( .A(
        o_data_odd_addr_gen_inst_int_base_addr_8_), .B(1'b0), .CI(
        o_data_odd_addr_gen_inst_add_45_carry[8]), .CO(
        o_data_odd_addr_gen_inst_add_45_carry[9]), .S(
        o_data_odd_addr_gen_inst_N28) );
  FA_X1 o_data_odd_addr_gen_inst_add_45_U1_9 ( .A(
        o_data_odd_addr_gen_inst_int_base_addr_9_), .B(1'b0), .CI(
        o_data_odd_addr_gen_inst_add_45_carry[9]), .S(
        o_data_odd_addr_gen_inst_N29) );
  AND2_X1 o_data_odd_addr_gen_inst_add_43_U2 ( .A1(1'b1), .A2(
        o_data_odd_addr[0]), .ZN(o_data_odd_addr_gen_inst_add_43_n2) );
  XOR2_X1 o_data_odd_addr_gen_inst_add_43_U1 ( .A(1'b1), .B(o_data_odd_addr[0]), .Z(o_data_odd_addr_gen_inst_N10) );
  FA_X1 o_data_odd_addr_gen_inst_add_43_U1_1 ( .A(o_data_odd_addr[1]), .B(1'b0), .CI(o_data_odd_addr_gen_inst_add_43_n2), .CO(
        o_data_odd_addr_gen_inst_add_43_carry[2]), .S(
        o_data_odd_addr_gen_inst_N11) );
  FA_X1 o_data_odd_addr_gen_inst_add_43_U1_2 ( .A(o_data_odd_addr[2]), .B(1'b0), .CI(o_data_odd_addr_gen_inst_add_43_carry[2]), .CO(
        o_data_odd_addr_gen_inst_add_43_carry[3]), .S(
        o_data_odd_addr_gen_inst_N12) );
  FA_X1 o_data_odd_addr_gen_inst_add_43_U1_3 ( .A(o_data_odd_addr[3]), .B(1'b0), .CI(o_data_odd_addr_gen_inst_add_43_carry[3]), .CO(
        o_data_odd_addr_gen_inst_add_43_carry[4]), .S(
        o_data_odd_addr_gen_inst_N13) );
  FA_X1 o_data_odd_addr_gen_inst_add_43_U1_4 ( .A(o_data_odd_addr[4]), .B(1'b0), .CI(o_data_odd_addr_gen_inst_add_43_carry[4]), .CO(
        o_data_odd_addr_gen_inst_add_43_carry[5]), .S(
        o_data_odd_addr_gen_inst_N14) );
  FA_X1 o_data_odd_addr_gen_inst_add_43_U1_5 ( .A(o_data_odd_addr[5]), .B(1'b0), .CI(o_data_odd_addr_gen_inst_add_43_carry[5]), .CO(
        o_data_odd_addr_gen_inst_add_43_carry[6]), .S(
        o_data_odd_addr_gen_inst_N15) );
  FA_X1 o_data_odd_addr_gen_inst_add_43_U1_6 ( .A(o_data_odd_addr[6]), .B(1'b0), .CI(o_data_odd_addr_gen_inst_add_43_carry[6]), .CO(
        o_data_odd_addr_gen_inst_add_43_carry[7]), .S(
        o_data_odd_addr_gen_inst_N16) );
  FA_X1 o_data_odd_addr_gen_inst_add_43_U1_7 ( .A(o_data_odd_addr[7]), .B(1'b0), .CI(o_data_odd_addr_gen_inst_add_43_carry[7]), .CO(
        o_data_odd_addr_gen_inst_add_43_carry[8]), .S(
        o_data_odd_addr_gen_inst_N17) );
  FA_X1 o_data_odd_addr_gen_inst_add_43_U1_8 ( .A(o_data_odd_addr[8]), .B(1'b0), .CI(o_data_odd_addr_gen_inst_add_43_carry[8]), .CO(
        o_data_odd_addr_gen_inst_add_43_carry[9]), .S(
        o_data_odd_addr_gen_inst_N18) );
  FA_X1 o_data_odd_addr_gen_inst_add_43_U1_9 ( .A(o_data_odd_addr[9]), .B(1'b0), .CI(o_data_odd_addr_gen_inst_add_43_carry[9]), .S(
        o_data_odd_addr_gen_inst_N19) );
  XOR2_X1 o_data_odd_addr_gen_inst_add_31_U2 ( .A(
        o_data_odd_addr_gen_inst_int_offs_addr_0_), .B(
        o_data_odd_addr_gen_inst_int_base_addr_0_), .Z(o_data_odd_addr[0]) );
  AND2_X1 o_data_odd_addr_gen_inst_add_31_U1 ( .A1(
        o_data_odd_addr_gen_inst_int_offs_addr_0_), .A2(
        o_data_odd_addr_gen_inst_int_base_addr_0_), .ZN(
        o_data_odd_addr_gen_inst_add_31_n1) );
  FA_X1 o_data_odd_addr_gen_inst_add_31_U1_1 ( .A(
        o_data_odd_addr_gen_inst_int_base_addr_1_), .B(
        o_data_odd_addr_gen_inst_int_offs_addr_1_), .CI(
        o_data_odd_addr_gen_inst_add_31_n1), .CO(
        o_data_odd_addr_gen_inst_add_31_carry[2]), .S(o_data_odd_addr[1]) );
  FA_X1 o_data_odd_addr_gen_inst_add_31_U1_2 ( .A(
        o_data_odd_addr_gen_inst_int_base_addr_2_), .B(
        o_data_odd_addr_gen_inst_int_offs_addr_2_), .CI(
        o_data_odd_addr_gen_inst_add_31_carry[2]), .CO(
        o_data_odd_addr_gen_inst_add_31_carry[3]), .S(o_data_odd_addr[2]) );
  FA_X1 o_data_odd_addr_gen_inst_add_31_U1_3 ( .A(
        o_data_odd_addr_gen_inst_int_base_addr_3_), .B(
        o_data_odd_addr_gen_inst_int_offs_addr_3_), .CI(
        o_data_odd_addr_gen_inst_add_31_carry[3]), .CO(
        o_data_odd_addr_gen_inst_add_31_carry[4]), .S(o_data_odd_addr[3]) );
  FA_X1 o_data_odd_addr_gen_inst_add_31_U1_4 ( .A(
        o_data_odd_addr_gen_inst_int_base_addr_4_), .B(
        o_data_odd_addr_gen_inst_int_offs_addr_4_), .CI(
        o_data_odd_addr_gen_inst_add_31_carry[4]), .CO(
        o_data_odd_addr_gen_inst_add_31_carry[5]), .S(o_data_odd_addr[4]) );
  FA_X1 o_data_odd_addr_gen_inst_add_31_U1_5 ( .A(
        o_data_odd_addr_gen_inst_int_base_addr_5_), .B(
        o_data_odd_addr_gen_inst_int_offs_addr_5_), .CI(
        o_data_odd_addr_gen_inst_add_31_carry[5]), .CO(
        o_data_odd_addr_gen_inst_add_31_carry[6]), .S(o_data_odd_addr[5]) );
  FA_X1 o_data_odd_addr_gen_inst_add_31_U1_6 ( .A(
        o_data_odd_addr_gen_inst_int_base_addr_6_), .B(
        o_data_odd_addr_gen_inst_int_offs_addr_6_), .CI(
        o_data_odd_addr_gen_inst_add_31_carry[6]), .CO(
        o_data_odd_addr_gen_inst_add_31_carry[7]), .S(o_data_odd_addr[6]) );
  FA_X1 o_data_odd_addr_gen_inst_add_31_U1_7 ( .A(
        o_data_odd_addr_gen_inst_int_base_addr_7_), .B(
        o_data_odd_addr_gen_inst_int_offs_addr_7_), .CI(
        o_data_odd_addr_gen_inst_add_31_carry[7]), .CO(
        o_data_odd_addr_gen_inst_add_31_carry[8]), .S(o_data_odd_addr[7]) );
  FA_X1 o_data_odd_addr_gen_inst_add_31_U1_8 ( .A(
        o_data_odd_addr_gen_inst_int_base_addr_8_), .B(
        o_data_odd_addr_gen_inst_int_offs_addr_8_), .CI(
        o_data_odd_addr_gen_inst_add_31_carry[8]), .CO(
        o_data_odd_addr_gen_inst_add_31_carry[9]), .S(o_data_odd_addr[8]) );
  FA_X1 o_data_odd_addr_gen_inst_add_31_U1_9 ( .A(
        o_data_odd_addr_gen_inst_int_base_addr_9_), .B(
        o_data_odd_addr_gen_inst_int_offs_addr_9_), .CI(
        o_data_odd_addr_gen_inst_add_31_carry[9]), .S(o_data_odd_addr[9]) );
  CLKGATETST_X1 clk_gate_int_q_tc_reg_latch ( .CK(ck), .E(s_tc_res), .SE(1'b0), 
        .GCK(net2764) );
endmodule

