
module npu ( ck, rst, en, ldh_v_n, wr_pipe, ckg_rmask, ckg_cmask, i_ifmap_ptr, 
        i_weight, i_data_conv_h, i_data_conv_v, i_data_acc, o_data );
  input [0:7] ckg_rmask;
  input [0:7] ckg_cmask;
  input [2:0] i_ifmap_ptr;
  input [1:0] i_weight;
  input [31:0] i_data_conv_h;
  input [31:0] i_data_conv_v;
  input [63:0] i_data_acc;
  output [63:0] o_data;
  input ck, rst, en, ldh_v_n, wr_pipe;
  wire   int_data_x_0__1__3_, int_data_x_0__1__2_, int_data_x_0__1__1_,
         int_data_x_0__1__0_, int_data_x_0__2__3_, int_data_x_0__2__2_,
         int_data_x_0__2__1_, int_data_x_0__2__0_, int_data_x_0__3__3_,
         int_data_x_0__3__2_, int_data_x_0__3__1_, int_data_x_0__3__0_,
         int_data_x_0__4__3_, int_data_x_0__4__2_, int_data_x_0__4__1_,
         int_data_x_0__4__0_, int_data_x_0__5__3_, int_data_x_0__5__2_,
         int_data_x_0__5__1_, int_data_x_0__5__0_, int_data_x_0__6__3_,
         int_data_x_0__6__2_, int_data_x_0__6__1_, int_data_x_0__6__0_,
         int_data_x_0__7__3_, int_data_x_0__7__2_, int_data_x_0__7__1_,
         int_data_x_0__7__0_, int_data_x_1__1__3_, int_data_x_1__1__2_,
         int_data_x_1__1__1_, int_data_x_1__1__0_, int_data_x_1__2__3_,
         int_data_x_1__2__2_, int_data_x_1__2__1_, int_data_x_1__2__0_,
         int_data_x_1__3__3_, int_data_x_1__3__2_, int_data_x_1__3__1_,
         int_data_x_1__3__0_, int_data_x_1__4__3_, int_data_x_1__4__2_,
         int_data_x_1__4__1_, int_data_x_1__4__0_, int_data_x_1__5__3_,
         int_data_x_1__5__2_, int_data_x_1__5__1_, int_data_x_1__5__0_,
         int_data_x_1__6__3_, int_data_x_1__6__2_, int_data_x_1__6__1_,
         int_data_x_1__6__0_, int_data_x_1__7__3_, int_data_x_1__7__2_,
         int_data_x_1__7__1_, int_data_x_1__7__0_, int_data_x_2__1__3_,
         int_data_x_2__1__2_, int_data_x_2__1__1_, int_data_x_2__1__0_,
         int_data_x_2__2__3_, int_data_x_2__2__2_, int_data_x_2__2__1_,
         int_data_x_2__2__0_, int_data_x_2__3__3_, int_data_x_2__3__2_,
         int_data_x_2__3__1_, int_data_x_2__3__0_, int_data_x_2__4__3_,
         int_data_x_2__4__2_, int_data_x_2__4__1_, int_data_x_2__4__0_,
         int_data_x_2__5__3_, int_data_x_2__5__2_, int_data_x_2__5__1_,
         int_data_x_2__5__0_, int_data_x_2__6__3_, int_data_x_2__6__2_,
         int_data_x_2__6__1_, int_data_x_2__6__0_, int_data_x_2__7__3_,
         int_data_x_2__7__2_, int_data_x_2__7__1_, int_data_x_2__7__0_,
         int_data_x_3__1__3_, int_data_x_3__1__2_, int_data_x_3__1__1_,
         int_data_x_3__1__0_, int_data_x_3__2__3_, int_data_x_3__2__2_,
         int_data_x_3__2__1_, int_data_x_3__2__0_, int_data_x_3__3__3_,
         int_data_x_3__3__2_, int_data_x_3__3__1_, int_data_x_3__3__0_,
         int_data_x_3__4__3_, int_data_x_3__4__2_, int_data_x_3__4__1_,
         int_data_x_3__4__0_, int_data_x_3__5__3_, int_data_x_3__5__2_,
         int_data_x_3__5__1_, int_data_x_3__5__0_, int_data_x_3__6__3_,
         int_data_x_3__6__2_, int_data_x_3__6__1_, int_data_x_3__6__0_,
         int_data_x_3__7__3_, int_data_x_3__7__2_, int_data_x_3__7__1_,
         int_data_x_3__7__0_, int_data_x_4__1__3_, int_data_x_4__1__2_,
         int_data_x_4__1__1_, int_data_x_4__1__0_, int_data_x_4__2__3_,
         int_data_x_4__2__2_, int_data_x_4__2__1_, int_data_x_4__2__0_,
         int_data_x_4__3__3_, int_data_x_4__3__2_, int_data_x_4__3__1_,
         int_data_x_4__3__0_, int_data_x_4__4__3_, int_data_x_4__4__2_,
         int_data_x_4__4__1_, int_data_x_4__4__0_, int_data_x_4__5__3_,
         int_data_x_4__5__2_, int_data_x_4__5__1_, int_data_x_4__5__0_,
         int_data_x_4__6__3_, int_data_x_4__6__2_, int_data_x_4__6__1_,
         int_data_x_4__6__0_, int_data_x_4__7__3_, int_data_x_4__7__2_,
         int_data_x_4__7__1_, int_data_x_4__7__0_, int_data_x_5__1__3_,
         int_data_x_5__1__2_, int_data_x_5__1__1_, int_data_x_5__1__0_,
         int_data_x_5__2__3_, int_data_x_5__2__2_, int_data_x_5__2__1_,
         int_data_x_5__2__0_, int_data_x_5__3__3_, int_data_x_5__3__2_,
         int_data_x_5__3__1_, int_data_x_5__3__0_, int_data_x_5__4__3_,
         int_data_x_5__4__2_, int_data_x_5__4__1_, int_data_x_5__4__0_,
         int_data_x_5__5__3_, int_data_x_5__5__2_, int_data_x_5__5__1_,
         int_data_x_5__5__0_, int_data_x_5__6__3_, int_data_x_5__6__2_,
         int_data_x_5__6__1_, int_data_x_5__6__0_, int_data_x_5__7__3_,
         int_data_x_5__7__2_, int_data_x_5__7__1_, int_data_x_5__7__0_,
         int_data_x_6__1__3_, int_data_x_6__1__2_, int_data_x_6__1__1_,
         int_data_x_6__1__0_, int_data_x_6__2__3_, int_data_x_6__2__2_,
         int_data_x_6__2__1_, int_data_x_6__2__0_, int_data_x_6__3__3_,
         int_data_x_6__3__2_, int_data_x_6__3__1_, int_data_x_6__3__0_,
         int_data_x_6__4__3_, int_data_x_6__4__2_, int_data_x_6__4__1_,
         int_data_x_6__4__0_, int_data_x_6__5__3_, int_data_x_6__5__2_,
         int_data_x_6__5__1_, int_data_x_6__5__0_, int_data_x_6__6__3_,
         int_data_x_6__6__2_, int_data_x_6__6__1_, int_data_x_6__6__0_,
         int_data_x_6__7__3_, int_data_x_6__7__2_, int_data_x_6__7__1_,
         int_data_x_6__7__0_, int_data_x_7__1__3_, int_data_x_7__1__2_,
         int_data_x_7__1__1_, int_data_x_7__1__0_, int_data_x_7__2__3_,
         int_data_x_7__2__2_, int_data_x_7__2__1_, int_data_x_7__2__0_,
         int_data_x_7__3__3_, int_data_x_7__3__2_, int_data_x_7__3__1_,
         int_data_x_7__3__0_, int_data_x_7__4__3_, int_data_x_7__4__2_,
         int_data_x_7__4__1_, int_data_x_7__4__0_, int_data_x_7__5__3_,
         int_data_x_7__5__2_, int_data_x_7__5__1_, int_data_x_7__5__0_,
         int_data_x_7__6__3_, int_data_x_7__6__2_, int_data_x_7__6__1_,
         int_data_x_7__6__0_, int_data_x_7__7__3_, int_data_x_7__7__2_,
         int_data_x_7__7__1_, int_data_x_7__7__0_, int_data_y_1__0__3_,
         int_data_y_1__0__2_, int_data_y_1__0__1_, int_data_y_1__0__0_,
         int_data_y_1__1__3_, int_data_y_1__1__2_, int_data_y_1__1__1_,
         int_data_y_1__1__0_, int_data_y_1__2__3_, int_data_y_1__2__2_,
         int_data_y_1__2__1_, int_data_y_1__2__0_, int_data_y_1__3__3_,
         int_data_y_1__3__2_, int_data_y_1__3__1_, int_data_y_1__3__0_,
         int_data_y_1__4__3_, int_data_y_1__4__2_, int_data_y_1__4__1_,
         int_data_y_1__4__0_, int_data_y_1__5__3_, int_data_y_1__5__2_,
         int_data_y_1__5__1_, int_data_y_1__5__0_, int_data_y_1__6__3_,
         int_data_y_1__6__2_, int_data_y_1__6__1_, int_data_y_1__6__0_,
         int_data_y_1__7__3_, int_data_y_1__7__2_, int_data_y_1__7__1_,
         int_data_y_1__7__0_, int_data_y_2__0__3_, int_data_y_2__0__2_,
         int_data_y_2__0__1_, int_data_y_2__0__0_, int_data_y_2__1__3_,
         int_data_y_2__1__2_, int_data_y_2__1__1_, int_data_y_2__1__0_,
         int_data_y_2__2__3_, int_data_y_2__2__2_, int_data_y_2__2__1_,
         int_data_y_2__2__0_, int_data_y_2__3__3_, int_data_y_2__3__2_,
         int_data_y_2__3__1_, int_data_y_2__3__0_, int_data_y_2__4__3_,
         int_data_y_2__4__2_, int_data_y_2__4__1_, int_data_y_2__4__0_,
         int_data_y_2__5__3_, int_data_y_2__5__2_, int_data_y_2__5__1_,
         int_data_y_2__5__0_, int_data_y_2__6__3_, int_data_y_2__6__2_,
         int_data_y_2__6__1_, int_data_y_2__6__0_, int_data_y_2__7__3_,
         int_data_y_2__7__2_, int_data_y_2__7__1_, int_data_y_2__7__0_,
         int_data_y_3__0__3_, int_data_y_3__0__2_, int_data_y_3__0__1_,
         int_data_y_3__0__0_, int_data_y_3__1__3_, int_data_y_3__1__2_,
         int_data_y_3__1__1_, int_data_y_3__1__0_, int_data_y_3__2__3_,
         int_data_y_3__2__2_, int_data_y_3__2__1_, int_data_y_3__2__0_,
         int_data_y_3__3__3_, int_data_y_3__3__2_, int_data_y_3__3__1_,
         int_data_y_3__3__0_, int_data_y_3__4__3_, int_data_y_3__4__2_,
         int_data_y_3__4__1_, int_data_y_3__4__0_, int_data_y_3__5__3_,
         int_data_y_3__5__2_, int_data_y_3__5__1_, int_data_y_3__5__0_,
         int_data_y_3__6__3_, int_data_y_3__6__2_, int_data_y_3__6__1_,
         int_data_y_3__6__0_, int_data_y_3__7__3_, int_data_y_3__7__2_,
         int_data_y_3__7__1_, int_data_y_3__7__0_, int_data_y_4__0__3_,
         int_data_y_4__0__2_, int_data_y_4__0__1_, int_data_y_4__0__0_,
         int_data_y_4__1__3_, int_data_y_4__1__2_, int_data_y_4__1__1_,
         int_data_y_4__1__0_, int_data_y_4__2__3_, int_data_y_4__2__2_,
         int_data_y_4__2__1_, int_data_y_4__2__0_, int_data_y_4__3__3_,
         int_data_y_4__3__2_, int_data_y_4__3__1_, int_data_y_4__3__0_,
         int_data_y_4__4__3_, int_data_y_4__4__2_, int_data_y_4__4__1_,
         int_data_y_4__4__0_, int_data_y_4__5__3_, int_data_y_4__5__2_,
         int_data_y_4__5__1_, int_data_y_4__5__0_, int_data_y_4__6__3_,
         int_data_y_4__6__2_, int_data_y_4__6__1_, int_data_y_4__6__0_,
         int_data_y_4__7__3_, int_data_y_4__7__2_, int_data_y_4__7__1_,
         int_data_y_4__7__0_, int_data_y_5__0__3_, int_data_y_5__0__2_,
         int_data_y_5__0__1_, int_data_y_5__0__0_, int_data_y_5__1__3_,
         int_data_y_5__1__2_, int_data_y_5__1__1_, int_data_y_5__1__0_,
         int_data_y_5__2__3_, int_data_y_5__2__2_, int_data_y_5__2__1_,
         int_data_y_5__2__0_, int_data_y_5__3__3_, int_data_y_5__3__2_,
         int_data_y_5__3__1_, int_data_y_5__3__0_, int_data_y_5__4__3_,
         int_data_y_5__4__2_, int_data_y_5__4__1_, int_data_y_5__4__0_,
         int_data_y_5__5__3_, int_data_y_5__5__2_, int_data_y_5__5__1_,
         int_data_y_5__5__0_, int_data_y_5__6__3_, int_data_y_5__6__2_,
         int_data_y_5__6__1_, int_data_y_5__6__0_, int_data_y_5__7__3_,
         int_data_y_5__7__2_, int_data_y_5__7__1_, int_data_y_5__7__0_,
         int_data_y_6__0__3_, int_data_y_6__0__2_, int_data_y_6__0__1_,
         int_data_y_6__0__0_, int_data_y_6__1__3_, int_data_y_6__1__2_,
         int_data_y_6__1__1_, int_data_y_6__1__0_, int_data_y_6__2__3_,
         int_data_y_6__2__2_, int_data_y_6__2__1_, int_data_y_6__2__0_,
         int_data_y_6__3__3_, int_data_y_6__3__2_, int_data_y_6__3__1_,
         int_data_y_6__3__0_, int_data_y_6__4__3_, int_data_y_6__4__2_,
         int_data_y_6__4__1_, int_data_y_6__4__0_, int_data_y_6__5__3_,
         int_data_y_6__5__2_, int_data_y_6__5__1_, int_data_y_6__5__0_,
         int_data_y_6__6__3_, int_data_y_6__6__2_, int_data_y_6__6__1_,
         int_data_y_6__6__0_, int_data_y_6__7__3_, int_data_y_6__7__2_,
         int_data_y_6__7__1_, int_data_y_6__7__0_, int_data_y_7__0__3_,
         int_data_y_7__0__2_, int_data_y_7__0__1_, int_data_y_7__0__0_,
         int_data_y_7__1__3_, int_data_y_7__1__2_, int_data_y_7__1__1_,
         int_data_y_7__1__0_, int_data_y_7__2__3_, int_data_y_7__2__2_,
         int_data_y_7__2__1_, int_data_y_7__2__0_, int_data_y_7__3__3_,
         int_data_y_7__3__2_, int_data_y_7__3__1_, int_data_y_7__3__0_,
         int_data_y_7__4__3_, int_data_y_7__4__2_, int_data_y_7__4__1_,
         int_data_y_7__4__0_, int_data_y_7__5__3_, int_data_y_7__5__2_,
         int_data_y_7__5__1_, int_data_y_7__5__0_, int_data_y_7__6__3_,
         int_data_y_7__6__2_, int_data_y_7__6__1_, int_data_y_7__6__0_,
         int_data_y_7__7__3_, int_data_y_7__7__2_, int_data_y_7__7__1_,
         int_data_y_7__7__0_, int_data_res_1__0__7_, int_data_res_1__0__6_,
         int_data_res_1__0__5_, int_data_res_1__0__4_, int_data_res_1__0__3_,
         int_data_res_1__0__2_, int_data_res_1__0__1_, int_data_res_1__0__0_,
         int_data_res_1__1__7_, int_data_res_1__1__6_, int_data_res_1__1__5_,
         int_data_res_1__1__4_, int_data_res_1__1__3_, int_data_res_1__1__2_,
         int_data_res_1__1__1_, int_data_res_1__1__0_, int_data_res_1__2__7_,
         int_data_res_1__2__6_, int_data_res_1__2__5_, int_data_res_1__2__4_,
         int_data_res_1__2__3_, int_data_res_1__2__2_, int_data_res_1__2__1_,
         int_data_res_1__2__0_, int_data_res_1__3__7_, int_data_res_1__3__6_,
         int_data_res_1__3__5_, int_data_res_1__3__4_, int_data_res_1__3__3_,
         int_data_res_1__3__2_, int_data_res_1__3__1_, int_data_res_1__3__0_,
         int_data_res_1__4__7_, int_data_res_1__4__6_, int_data_res_1__4__5_,
         int_data_res_1__4__4_, int_data_res_1__4__3_, int_data_res_1__4__2_,
         int_data_res_1__4__1_, int_data_res_1__4__0_, int_data_res_1__5__7_,
         int_data_res_1__5__6_, int_data_res_1__5__5_, int_data_res_1__5__4_,
         int_data_res_1__5__3_, int_data_res_1__5__2_, int_data_res_1__5__1_,
         int_data_res_1__5__0_, int_data_res_1__6__7_, int_data_res_1__6__6_,
         int_data_res_1__6__5_, int_data_res_1__6__4_, int_data_res_1__6__3_,
         int_data_res_1__6__2_, int_data_res_1__6__1_, int_data_res_1__6__0_,
         int_data_res_1__7__7_, int_data_res_1__7__6_, int_data_res_1__7__5_,
         int_data_res_1__7__4_, int_data_res_1__7__3_, int_data_res_1__7__2_,
         int_data_res_1__7__1_, int_data_res_1__7__0_, int_data_res_2__0__7_,
         int_data_res_2__0__6_, int_data_res_2__0__5_, int_data_res_2__0__4_,
         int_data_res_2__0__3_, int_data_res_2__0__2_, int_data_res_2__0__1_,
         int_data_res_2__0__0_, int_data_res_2__1__7_, int_data_res_2__1__6_,
         int_data_res_2__1__5_, int_data_res_2__1__4_, int_data_res_2__1__3_,
         int_data_res_2__1__2_, int_data_res_2__1__1_, int_data_res_2__1__0_,
         int_data_res_2__2__7_, int_data_res_2__2__6_, int_data_res_2__2__5_,
         int_data_res_2__2__4_, int_data_res_2__2__3_, int_data_res_2__2__2_,
         int_data_res_2__2__1_, int_data_res_2__2__0_, int_data_res_2__3__7_,
         int_data_res_2__3__6_, int_data_res_2__3__5_, int_data_res_2__3__4_,
         int_data_res_2__3__3_, int_data_res_2__3__2_, int_data_res_2__3__1_,
         int_data_res_2__3__0_, int_data_res_2__4__7_, int_data_res_2__4__6_,
         int_data_res_2__4__5_, int_data_res_2__4__4_, int_data_res_2__4__3_,
         int_data_res_2__4__2_, int_data_res_2__4__1_, int_data_res_2__4__0_,
         int_data_res_2__5__7_, int_data_res_2__5__6_, int_data_res_2__5__5_,
         int_data_res_2__5__4_, int_data_res_2__5__3_, int_data_res_2__5__2_,
         int_data_res_2__5__1_, int_data_res_2__5__0_, int_data_res_2__6__7_,
         int_data_res_2__6__6_, int_data_res_2__6__5_, int_data_res_2__6__4_,
         int_data_res_2__6__3_, int_data_res_2__6__2_, int_data_res_2__6__1_,
         int_data_res_2__6__0_, int_data_res_2__7__7_, int_data_res_2__7__6_,
         int_data_res_2__7__5_, int_data_res_2__7__4_, int_data_res_2__7__3_,
         int_data_res_2__7__2_, int_data_res_2__7__1_, int_data_res_2__7__0_,
         int_data_res_3__0__7_, int_data_res_3__0__6_, int_data_res_3__0__5_,
         int_data_res_3__0__4_, int_data_res_3__0__3_, int_data_res_3__0__2_,
         int_data_res_3__0__1_, int_data_res_3__0__0_, int_data_res_3__1__7_,
         int_data_res_3__1__6_, int_data_res_3__1__5_, int_data_res_3__1__4_,
         int_data_res_3__1__3_, int_data_res_3__1__2_, int_data_res_3__1__1_,
         int_data_res_3__1__0_, int_data_res_3__2__7_, int_data_res_3__2__6_,
         int_data_res_3__2__5_, int_data_res_3__2__4_, int_data_res_3__2__3_,
         int_data_res_3__2__2_, int_data_res_3__2__1_, int_data_res_3__2__0_,
         int_data_res_3__3__7_, int_data_res_3__3__6_, int_data_res_3__3__5_,
         int_data_res_3__3__4_, int_data_res_3__3__3_, int_data_res_3__3__2_,
         int_data_res_3__3__1_, int_data_res_3__3__0_, int_data_res_3__4__7_,
         int_data_res_3__4__6_, int_data_res_3__4__5_, int_data_res_3__4__4_,
         int_data_res_3__4__3_, int_data_res_3__4__2_, int_data_res_3__4__1_,
         int_data_res_3__4__0_, int_data_res_3__5__7_, int_data_res_3__5__6_,
         int_data_res_3__5__5_, int_data_res_3__5__4_, int_data_res_3__5__3_,
         int_data_res_3__5__2_, int_data_res_3__5__1_, int_data_res_3__5__0_,
         int_data_res_3__6__7_, int_data_res_3__6__6_, int_data_res_3__6__5_,
         int_data_res_3__6__4_, int_data_res_3__6__3_, int_data_res_3__6__2_,
         int_data_res_3__6__1_, int_data_res_3__6__0_, int_data_res_3__7__7_,
         int_data_res_3__7__6_, int_data_res_3__7__5_, int_data_res_3__7__4_,
         int_data_res_3__7__3_, int_data_res_3__7__2_, int_data_res_3__7__1_,
         int_data_res_3__7__0_, int_data_res_4__0__7_, int_data_res_4__0__6_,
         int_data_res_4__0__5_, int_data_res_4__0__4_, int_data_res_4__0__3_,
         int_data_res_4__0__2_, int_data_res_4__0__1_, int_data_res_4__0__0_,
         int_data_res_4__1__7_, int_data_res_4__1__6_, int_data_res_4__1__5_,
         int_data_res_4__1__4_, int_data_res_4__1__3_, int_data_res_4__1__2_,
         int_data_res_4__1__1_, int_data_res_4__1__0_, int_data_res_4__2__7_,
         int_data_res_4__2__6_, int_data_res_4__2__5_, int_data_res_4__2__4_,
         int_data_res_4__2__3_, int_data_res_4__2__2_, int_data_res_4__2__1_,
         int_data_res_4__2__0_, int_data_res_4__3__7_, int_data_res_4__3__6_,
         int_data_res_4__3__5_, int_data_res_4__3__4_, int_data_res_4__3__3_,
         int_data_res_4__3__2_, int_data_res_4__3__1_, int_data_res_4__3__0_,
         int_data_res_4__4__7_, int_data_res_4__4__6_, int_data_res_4__4__5_,
         int_data_res_4__4__4_, int_data_res_4__4__3_, int_data_res_4__4__2_,
         int_data_res_4__4__1_, int_data_res_4__4__0_, int_data_res_4__5__7_,
         int_data_res_4__5__6_, int_data_res_4__5__5_, int_data_res_4__5__4_,
         int_data_res_4__5__3_, int_data_res_4__5__2_, int_data_res_4__5__1_,
         int_data_res_4__5__0_, int_data_res_4__6__7_, int_data_res_4__6__6_,
         int_data_res_4__6__5_, int_data_res_4__6__4_, int_data_res_4__6__3_,
         int_data_res_4__6__2_, int_data_res_4__6__1_, int_data_res_4__6__0_,
         int_data_res_4__7__7_, int_data_res_4__7__6_, int_data_res_4__7__5_,
         int_data_res_4__7__4_, int_data_res_4__7__3_, int_data_res_4__7__2_,
         int_data_res_4__7__1_, int_data_res_4__7__0_, int_data_res_5__0__7_,
         int_data_res_5__0__6_, int_data_res_5__0__5_, int_data_res_5__0__4_,
         int_data_res_5__0__3_, int_data_res_5__0__2_, int_data_res_5__0__1_,
         int_data_res_5__0__0_, int_data_res_5__1__7_, int_data_res_5__1__6_,
         int_data_res_5__1__5_, int_data_res_5__1__4_, int_data_res_5__1__3_,
         int_data_res_5__1__2_, int_data_res_5__1__1_, int_data_res_5__1__0_,
         int_data_res_5__2__7_, int_data_res_5__2__6_, int_data_res_5__2__5_,
         int_data_res_5__2__4_, int_data_res_5__2__3_, int_data_res_5__2__2_,
         int_data_res_5__2__1_, int_data_res_5__2__0_, int_data_res_5__3__7_,
         int_data_res_5__3__6_, int_data_res_5__3__5_, int_data_res_5__3__4_,
         int_data_res_5__3__3_, int_data_res_5__3__2_, int_data_res_5__3__1_,
         int_data_res_5__3__0_, int_data_res_5__4__7_, int_data_res_5__4__6_,
         int_data_res_5__4__5_, int_data_res_5__4__4_, int_data_res_5__4__3_,
         int_data_res_5__4__2_, int_data_res_5__4__1_, int_data_res_5__4__0_,
         int_data_res_5__5__7_, int_data_res_5__5__6_, int_data_res_5__5__5_,
         int_data_res_5__5__4_, int_data_res_5__5__3_, int_data_res_5__5__2_,
         int_data_res_5__5__1_, int_data_res_5__5__0_, int_data_res_5__6__7_,
         int_data_res_5__6__6_, int_data_res_5__6__5_, int_data_res_5__6__4_,
         int_data_res_5__6__3_, int_data_res_5__6__2_, int_data_res_5__6__1_,
         int_data_res_5__6__0_, int_data_res_5__7__7_, int_data_res_5__7__6_,
         int_data_res_5__7__5_, int_data_res_5__7__4_, int_data_res_5__7__3_,
         int_data_res_5__7__2_, int_data_res_5__7__1_, int_data_res_5__7__0_,
         int_data_res_6__0__7_, int_data_res_6__0__6_, int_data_res_6__0__5_,
         int_data_res_6__0__4_, int_data_res_6__0__3_, int_data_res_6__0__2_,
         int_data_res_6__0__1_, int_data_res_6__0__0_, int_data_res_6__1__7_,
         int_data_res_6__1__6_, int_data_res_6__1__5_, int_data_res_6__1__4_,
         int_data_res_6__1__3_, int_data_res_6__1__2_, int_data_res_6__1__1_,
         int_data_res_6__1__0_, int_data_res_6__2__7_, int_data_res_6__2__6_,
         int_data_res_6__2__5_, int_data_res_6__2__4_, int_data_res_6__2__3_,
         int_data_res_6__2__2_, int_data_res_6__2__1_, int_data_res_6__2__0_,
         int_data_res_6__3__7_, int_data_res_6__3__6_, int_data_res_6__3__5_,
         int_data_res_6__3__4_, int_data_res_6__3__3_, int_data_res_6__3__2_,
         int_data_res_6__3__1_, int_data_res_6__3__0_, int_data_res_6__4__7_,
         int_data_res_6__4__6_, int_data_res_6__4__5_, int_data_res_6__4__4_,
         int_data_res_6__4__3_, int_data_res_6__4__2_, int_data_res_6__4__1_,
         int_data_res_6__4__0_, int_data_res_6__5__7_, int_data_res_6__5__6_,
         int_data_res_6__5__5_, int_data_res_6__5__4_, int_data_res_6__5__3_,
         int_data_res_6__5__2_, int_data_res_6__5__1_, int_data_res_6__5__0_,
         int_data_res_6__6__7_, int_data_res_6__6__6_, int_data_res_6__6__5_,
         int_data_res_6__6__4_, int_data_res_6__6__3_, int_data_res_6__6__2_,
         int_data_res_6__6__1_, int_data_res_6__6__0_, int_data_res_6__7__7_,
         int_data_res_6__7__6_, int_data_res_6__7__5_, int_data_res_6__7__4_,
         int_data_res_6__7__3_, int_data_res_6__7__2_, int_data_res_6__7__1_,
         int_data_res_6__7__0_, int_data_res_7__0__7_, int_data_res_7__0__6_,
         int_data_res_7__0__5_, int_data_res_7__0__4_, int_data_res_7__0__3_,
         int_data_res_7__0__2_, int_data_res_7__0__1_, int_data_res_7__0__0_,
         int_data_res_7__1__7_, int_data_res_7__1__6_, int_data_res_7__1__5_,
         int_data_res_7__1__4_, int_data_res_7__1__3_, int_data_res_7__1__2_,
         int_data_res_7__1__1_, int_data_res_7__1__0_, int_data_res_7__2__7_,
         int_data_res_7__2__6_, int_data_res_7__2__5_, int_data_res_7__2__4_,
         int_data_res_7__2__3_, int_data_res_7__2__2_, int_data_res_7__2__1_,
         int_data_res_7__2__0_, int_data_res_7__3__7_, int_data_res_7__3__6_,
         int_data_res_7__3__5_, int_data_res_7__3__4_, int_data_res_7__3__3_,
         int_data_res_7__3__2_, int_data_res_7__3__1_, int_data_res_7__3__0_,
         int_data_res_7__4__7_, int_data_res_7__4__6_, int_data_res_7__4__5_,
         int_data_res_7__4__4_, int_data_res_7__4__3_, int_data_res_7__4__2_,
         int_data_res_7__4__1_, int_data_res_7__4__0_, int_data_res_7__5__7_,
         int_data_res_7__5__6_, int_data_res_7__5__5_, int_data_res_7__5__4_,
         int_data_res_7__5__3_, int_data_res_7__5__2_, int_data_res_7__5__1_,
         int_data_res_7__5__0_, int_data_res_7__6__7_, int_data_res_7__6__6_,
         int_data_res_7__6__5_, int_data_res_7__6__4_, int_data_res_7__6__3_,
         int_data_res_7__6__2_, int_data_res_7__6__1_, int_data_res_7__6__0_,
         int_data_res_7__7__7_, int_data_res_7__7__6_, int_data_res_7__7__5_,
         int_data_res_7__7__4_, int_data_res_7__7__3_, int_data_res_7__7__2_,
         int_data_res_7__7__1_, int_data_res_7__7__0_, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         pe_1_0_0_n87, pe_1_0_0_n86, pe_1_0_0_n85, pe_1_0_0_n84, pe_1_0_0_n83,
         pe_1_0_0_n82, pe_1_0_0_n81, pe_1_0_0_n80, pe_1_0_0_n79, pe_1_0_0_n78,
         pe_1_0_0_n77, pe_1_0_0_n76, pe_1_0_0_n75, pe_1_0_0_n74, pe_1_0_0_n73,
         pe_1_0_0_n72, pe_1_0_0_n71, pe_1_0_0_n70, pe_1_0_0_n69, pe_1_0_0_n68,
         pe_1_0_0_n67, pe_1_0_0_n66, pe_1_0_0_n65, pe_1_0_0_n64, pe_1_0_0_n63,
         pe_1_0_0_n62, pe_1_0_0_n61, pe_1_0_0_n60, pe_1_0_0_n59, pe_1_0_0_n58,
         pe_1_0_0_n57, pe_1_0_0_n56, pe_1_0_0_n55, pe_1_0_0_n54, pe_1_0_0_n53,
         pe_1_0_0_n52, pe_1_0_0_n51, pe_1_0_0_n50, pe_1_0_0_n49, pe_1_0_0_n48,
         pe_1_0_0_n47, pe_1_0_0_n46, pe_1_0_0_n45, pe_1_0_0_n25, pe_1_0_0_n24,
         pe_1_0_0_n23, pe_1_0_0_n22, pe_1_0_0_n21, pe_1_0_0_n20, pe_1_0_0_n19,
         pe_1_0_0_n18, pe_1_0_0_n17, pe_1_0_0_n16, pe_1_0_0_n15, pe_1_0_0_n14,
         pe_1_0_0_n13, pe_1_0_0_n12, pe_1_0_0_n11, pe_1_0_0_n10, pe_1_0_0_n9,
         pe_1_0_0_n8, pe_1_0_0_n7, pe_1_0_0_n6, pe_1_0_0_n5, pe_1_0_0_n4,
         pe_1_0_0_n3, pe_1_0_0_n2, pe_1_0_0_n1, pe_1_0_0_n44, pe_1_0_0_n43,
         pe_1_0_0_n42, pe_1_0_0_n41, pe_1_0_0_n40, pe_1_0_0_n39, pe_1_0_0_n38,
         pe_1_0_0_n37, pe_1_0_0_n36, pe_1_0_0_n35, pe_1_0_0_n34, pe_1_0_0_n33,
         pe_1_0_0_n32, pe_1_0_0_n31, pe_1_0_0_n30, pe_1_0_0_n29, pe_1_0_0_n28,
         pe_1_0_0_n27, pe_1_0_0_n26, pe_1_0_0_net7552, pe_1_0_0_net7547,
         pe_1_0_0_net7542, pe_1_0_0_net7537, pe_1_0_0_net7532,
         pe_1_0_0_net7527, pe_1_0_0_net7522, pe_1_0_0_net7517,
         pe_1_0_0_net7512, pe_1_0_0_net7507, pe_1_0_0_net7502,
         pe_1_0_0_net7497, pe_1_0_0_net7491, pe_1_0_0_N90, pe_1_0_0_N85,
         pe_1_0_0_N84, pe_1_0_0_N83, pe_1_0_0_N82, pe_1_0_0_N81, pe_1_0_0_N80,
         pe_1_0_0_N79, pe_1_0_0_N77, pe_1_0_0_N76, pe_1_0_0_N75, pe_1_0_0_N74,
         pe_1_0_0_N73, pe_1_0_0_N72, pe_1_0_0_N71, pe_1_0_0_N70,
         pe_1_0_0_int_data_0_, pe_1_0_0_int_data_1_, pe_1_0_0_int_data_2_,
         pe_1_0_0_int_data_3_, pe_1_0_0_N64, pe_1_0_0_N63, pe_1_0_0_N62,
         pe_1_0_0_N61, pe_1_0_0_N60, pe_1_0_0_N59, pe_1_0_0_o_data_v_0_,
         pe_1_0_0_o_data_v_1_, pe_1_0_0_o_data_v_2_, pe_1_0_0_o_data_v_3_,
         pe_1_0_0_o_data_h_0_, pe_1_0_0_o_data_h_1_, pe_1_0_0_o_data_h_2_,
         pe_1_0_0_o_data_h_3_, pe_1_0_1_n86, pe_1_0_1_n85, pe_1_0_1_n84,
         pe_1_0_1_n83, pe_1_0_1_n82, pe_1_0_1_n81, pe_1_0_1_n80, pe_1_0_1_n79,
         pe_1_0_1_n78, pe_1_0_1_n77, pe_1_0_1_n76, pe_1_0_1_n75, pe_1_0_1_n74,
         pe_1_0_1_n73, pe_1_0_1_n72, pe_1_0_1_n71, pe_1_0_1_n70, pe_1_0_1_n69,
         pe_1_0_1_n68, pe_1_0_1_n67, pe_1_0_1_n66, pe_1_0_1_n65, pe_1_0_1_n64,
         pe_1_0_1_n63, pe_1_0_1_n62, pe_1_0_1_n61, pe_1_0_1_n60, pe_1_0_1_n59,
         pe_1_0_1_n58, pe_1_0_1_n57, pe_1_0_1_n56, pe_1_0_1_n55, pe_1_0_1_n54,
         pe_1_0_1_n53, pe_1_0_1_n52, pe_1_0_1_n51, pe_1_0_1_n50, pe_1_0_1_n49,
         pe_1_0_1_n48, pe_1_0_1_n47, pe_1_0_1_n46, pe_1_0_1_n45, pe_1_0_1_n25,
         pe_1_0_1_n24, pe_1_0_1_n23, pe_1_0_1_n22, pe_1_0_1_n21, pe_1_0_1_n20,
         pe_1_0_1_n19, pe_1_0_1_n18, pe_1_0_1_n17, pe_1_0_1_n16, pe_1_0_1_n15,
         pe_1_0_1_n14, pe_1_0_1_n13, pe_1_0_1_n12, pe_1_0_1_n11, pe_1_0_1_n10,
         pe_1_0_1_n9, pe_1_0_1_n8, pe_1_0_1_n7, pe_1_0_1_n6, pe_1_0_1_n5,
         pe_1_0_1_n4, pe_1_0_1_n3, pe_1_0_1_n2, pe_1_0_1_n1, pe_1_0_1_n44,
         pe_1_0_1_n43, pe_1_0_1_n42, pe_1_0_1_n41, pe_1_0_1_n40, pe_1_0_1_n39,
         pe_1_0_1_n38, pe_1_0_1_n37, pe_1_0_1_n36, pe_1_0_1_n35, pe_1_0_1_n34,
         pe_1_0_1_n33, pe_1_0_1_n32, pe_1_0_1_n31, pe_1_0_1_n30, pe_1_0_1_n29,
         pe_1_0_1_n28, pe_1_0_1_n27, pe_1_0_1_n26, pe_1_0_1_net7474,
         pe_1_0_1_net7469, pe_1_0_1_net7464, pe_1_0_1_net7459,
         pe_1_0_1_net7454, pe_1_0_1_net7449, pe_1_0_1_net7444,
         pe_1_0_1_net7439, pe_1_0_1_net7434, pe_1_0_1_net7429,
         pe_1_0_1_net7424, pe_1_0_1_net7419, pe_1_0_1_net7413, pe_1_0_1_N90,
         pe_1_0_1_N85, pe_1_0_1_N84, pe_1_0_1_N83, pe_1_0_1_N82, pe_1_0_1_N81,
         pe_1_0_1_N80, pe_1_0_1_N79, pe_1_0_1_N77, pe_1_0_1_N76, pe_1_0_1_N75,
         pe_1_0_1_N74, pe_1_0_1_N73, pe_1_0_1_N72, pe_1_0_1_N71, pe_1_0_1_N70,
         pe_1_0_1_int_data_0_, pe_1_0_1_int_data_1_, pe_1_0_1_int_data_2_,
         pe_1_0_1_int_data_3_, pe_1_0_1_N64, pe_1_0_1_N63, pe_1_0_1_N62,
         pe_1_0_1_N61, pe_1_0_1_N60, pe_1_0_1_N59, pe_1_0_1_o_data_v_0_,
         pe_1_0_1_o_data_v_1_, pe_1_0_1_o_data_v_2_, pe_1_0_1_o_data_v_3_,
         pe_1_0_2_n87, pe_1_0_2_n86, pe_1_0_2_n85, pe_1_0_2_n84, pe_1_0_2_n83,
         pe_1_0_2_n82, pe_1_0_2_n81, pe_1_0_2_n80, pe_1_0_2_n79, pe_1_0_2_n78,
         pe_1_0_2_n77, pe_1_0_2_n76, pe_1_0_2_n75, pe_1_0_2_n74, pe_1_0_2_n73,
         pe_1_0_2_n72, pe_1_0_2_n71, pe_1_0_2_n70, pe_1_0_2_n69, pe_1_0_2_n68,
         pe_1_0_2_n67, pe_1_0_2_n66, pe_1_0_2_n65, pe_1_0_2_n64, pe_1_0_2_n63,
         pe_1_0_2_n62, pe_1_0_2_n61, pe_1_0_2_n60, pe_1_0_2_n59, pe_1_0_2_n58,
         pe_1_0_2_n57, pe_1_0_2_n56, pe_1_0_2_n55, pe_1_0_2_n54, pe_1_0_2_n53,
         pe_1_0_2_n52, pe_1_0_2_n51, pe_1_0_2_n50, pe_1_0_2_n49, pe_1_0_2_n48,
         pe_1_0_2_n47, pe_1_0_2_n46, pe_1_0_2_n45, pe_1_0_2_n25, pe_1_0_2_n24,
         pe_1_0_2_n23, pe_1_0_2_n22, pe_1_0_2_n21, pe_1_0_2_n20, pe_1_0_2_n19,
         pe_1_0_2_n18, pe_1_0_2_n17, pe_1_0_2_n16, pe_1_0_2_n15, pe_1_0_2_n14,
         pe_1_0_2_n13, pe_1_0_2_n12, pe_1_0_2_n11, pe_1_0_2_n10, pe_1_0_2_n9,
         pe_1_0_2_n8, pe_1_0_2_n7, pe_1_0_2_n6, pe_1_0_2_n5, pe_1_0_2_n4,
         pe_1_0_2_n3, pe_1_0_2_n2, pe_1_0_2_n1, pe_1_0_2_n44, pe_1_0_2_n43,
         pe_1_0_2_n42, pe_1_0_2_n41, pe_1_0_2_n40, pe_1_0_2_n39, pe_1_0_2_n38,
         pe_1_0_2_n37, pe_1_0_2_n36, pe_1_0_2_n35, pe_1_0_2_n34, pe_1_0_2_n33,
         pe_1_0_2_n32, pe_1_0_2_n31, pe_1_0_2_n30, pe_1_0_2_n29, pe_1_0_2_n28,
         pe_1_0_2_n27, pe_1_0_2_n26, pe_1_0_2_net7396, pe_1_0_2_net7391,
         pe_1_0_2_net7386, pe_1_0_2_net7381, pe_1_0_2_net7376,
         pe_1_0_2_net7371, pe_1_0_2_net7366, pe_1_0_2_net7361,
         pe_1_0_2_net7356, pe_1_0_2_net7351, pe_1_0_2_net7346,
         pe_1_0_2_net7341, pe_1_0_2_net7335, pe_1_0_2_N90, pe_1_0_2_N85,
         pe_1_0_2_N84, pe_1_0_2_N83, pe_1_0_2_N82, pe_1_0_2_N81, pe_1_0_2_N80,
         pe_1_0_2_N79, pe_1_0_2_N77, pe_1_0_2_N76, pe_1_0_2_N75, pe_1_0_2_N74,
         pe_1_0_2_N73, pe_1_0_2_N72, pe_1_0_2_N71, pe_1_0_2_N70,
         pe_1_0_2_int_data_0_, pe_1_0_2_int_data_1_, pe_1_0_2_int_data_2_,
         pe_1_0_2_int_data_3_, pe_1_0_2_N64, pe_1_0_2_N63, pe_1_0_2_N62,
         pe_1_0_2_N61, pe_1_0_2_N60, pe_1_0_2_N59, pe_1_0_2_o_data_v_0_,
         pe_1_0_2_o_data_v_1_, pe_1_0_2_o_data_v_2_, pe_1_0_2_o_data_v_3_,
         pe_1_0_3_n88, pe_1_0_3_n87, pe_1_0_3_n86, pe_1_0_3_n85, pe_1_0_3_n84,
         pe_1_0_3_n83, pe_1_0_3_n82, pe_1_0_3_n81, pe_1_0_3_n80, pe_1_0_3_n79,
         pe_1_0_3_n78, pe_1_0_3_n77, pe_1_0_3_n76, pe_1_0_3_n75, pe_1_0_3_n74,
         pe_1_0_3_n73, pe_1_0_3_n72, pe_1_0_3_n71, pe_1_0_3_n70, pe_1_0_3_n69,
         pe_1_0_3_n68, pe_1_0_3_n67, pe_1_0_3_n66, pe_1_0_3_n65, pe_1_0_3_n64,
         pe_1_0_3_n63, pe_1_0_3_n62, pe_1_0_3_n61, pe_1_0_3_n60, pe_1_0_3_n59,
         pe_1_0_3_n58, pe_1_0_3_n57, pe_1_0_3_n56, pe_1_0_3_n55, pe_1_0_3_n54,
         pe_1_0_3_n53, pe_1_0_3_n52, pe_1_0_3_n51, pe_1_0_3_n50, pe_1_0_3_n49,
         pe_1_0_3_n48, pe_1_0_3_n47, pe_1_0_3_n46, pe_1_0_3_n45, pe_1_0_3_n25,
         pe_1_0_3_n24, pe_1_0_3_n23, pe_1_0_3_n22, pe_1_0_3_n21, pe_1_0_3_n20,
         pe_1_0_3_n19, pe_1_0_3_n18, pe_1_0_3_n17, pe_1_0_3_n16, pe_1_0_3_n15,
         pe_1_0_3_n14, pe_1_0_3_n13, pe_1_0_3_n12, pe_1_0_3_n11, pe_1_0_3_n10,
         pe_1_0_3_n9, pe_1_0_3_n8, pe_1_0_3_n7, pe_1_0_3_n6, pe_1_0_3_n5,
         pe_1_0_3_n4, pe_1_0_3_n3, pe_1_0_3_n2, pe_1_0_3_n1, pe_1_0_3_n44,
         pe_1_0_3_n43, pe_1_0_3_n42, pe_1_0_3_n41, pe_1_0_3_n40, pe_1_0_3_n39,
         pe_1_0_3_n38, pe_1_0_3_n37, pe_1_0_3_n36, pe_1_0_3_n35, pe_1_0_3_n34,
         pe_1_0_3_n33, pe_1_0_3_n32, pe_1_0_3_n31, pe_1_0_3_n30, pe_1_0_3_n29,
         pe_1_0_3_n28, pe_1_0_3_n27, pe_1_0_3_n26, pe_1_0_3_net7318,
         pe_1_0_3_net7313, pe_1_0_3_net7308, pe_1_0_3_net7303,
         pe_1_0_3_net7298, pe_1_0_3_net7293, pe_1_0_3_net7288,
         pe_1_0_3_net7283, pe_1_0_3_net7278, pe_1_0_3_net7273,
         pe_1_0_3_net7268, pe_1_0_3_net7263, pe_1_0_3_net7257, pe_1_0_3_N90,
         pe_1_0_3_N85, pe_1_0_3_N84, pe_1_0_3_N83, pe_1_0_3_N82, pe_1_0_3_N81,
         pe_1_0_3_N80, pe_1_0_3_N79, pe_1_0_3_N77, pe_1_0_3_N76, pe_1_0_3_N75,
         pe_1_0_3_N74, pe_1_0_3_N73, pe_1_0_3_N72, pe_1_0_3_N71, pe_1_0_3_N70,
         pe_1_0_3_int_data_0_, pe_1_0_3_int_data_1_, pe_1_0_3_int_data_2_,
         pe_1_0_3_int_data_3_, pe_1_0_3_N64, pe_1_0_3_N63, pe_1_0_3_N62,
         pe_1_0_3_N61, pe_1_0_3_N60, pe_1_0_3_N59, pe_1_0_3_o_data_v_0_,
         pe_1_0_3_o_data_v_1_, pe_1_0_3_o_data_v_2_, pe_1_0_3_o_data_v_3_,
         pe_1_0_4_n90, pe_1_0_4_n89, pe_1_0_4_n88, pe_1_0_4_n87, pe_1_0_4_n86,
         pe_1_0_4_n85, pe_1_0_4_n84, pe_1_0_4_n83, pe_1_0_4_n82, pe_1_0_4_n81,
         pe_1_0_4_n80, pe_1_0_4_n79, pe_1_0_4_n78, pe_1_0_4_n77, pe_1_0_4_n76,
         pe_1_0_4_n75, pe_1_0_4_n74, pe_1_0_4_n73, pe_1_0_4_n72, pe_1_0_4_n71,
         pe_1_0_4_n70, pe_1_0_4_n69, pe_1_0_4_n68, pe_1_0_4_n67, pe_1_0_4_n66,
         pe_1_0_4_n65, pe_1_0_4_n64, pe_1_0_4_n63, pe_1_0_4_n62, pe_1_0_4_n61,
         pe_1_0_4_n60, pe_1_0_4_n59, pe_1_0_4_n58, pe_1_0_4_n57, pe_1_0_4_n56,
         pe_1_0_4_n55, pe_1_0_4_n54, pe_1_0_4_n53, pe_1_0_4_n52, pe_1_0_4_n51,
         pe_1_0_4_n50, pe_1_0_4_n49, pe_1_0_4_n48, pe_1_0_4_n47, pe_1_0_4_n46,
         pe_1_0_4_n45, pe_1_0_4_n25, pe_1_0_4_n24, pe_1_0_4_n23, pe_1_0_4_n22,
         pe_1_0_4_n21, pe_1_0_4_n20, pe_1_0_4_n19, pe_1_0_4_n18, pe_1_0_4_n17,
         pe_1_0_4_n16, pe_1_0_4_n15, pe_1_0_4_n14, pe_1_0_4_n13, pe_1_0_4_n12,
         pe_1_0_4_n11, pe_1_0_4_n10, pe_1_0_4_n9, pe_1_0_4_n8, pe_1_0_4_n7,
         pe_1_0_4_n6, pe_1_0_4_n5, pe_1_0_4_n4, pe_1_0_4_n3, pe_1_0_4_n2,
         pe_1_0_4_n1, pe_1_0_4_n44, pe_1_0_4_n43, pe_1_0_4_n42, pe_1_0_4_n41,
         pe_1_0_4_n40, pe_1_0_4_n39, pe_1_0_4_n38, pe_1_0_4_n37, pe_1_0_4_n36,
         pe_1_0_4_n35, pe_1_0_4_n34, pe_1_0_4_n33, pe_1_0_4_n32, pe_1_0_4_n31,
         pe_1_0_4_n30, pe_1_0_4_n29, pe_1_0_4_n28, pe_1_0_4_n27, pe_1_0_4_n26,
         pe_1_0_4_net7240, pe_1_0_4_net7235, pe_1_0_4_net7230,
         pe_1_0_4_net7225, pe_1_0_4_net7220, pe_1_0_4_net7215,
         pe_1_0_4_net7210, pe_1_0_4_net7205, pe_1_0_4_net7200,
         pe_1_0_4_net7195, pe_1_0_4_net7190, pe_1_0_4_net7185,
         pe_1_0_4_net7179, pe_1_0_4_N90, pe_1_0_4_N85, pe_1_0_4_N84,
         pe_1_0_4_N83, pe_1_0_4_N82, pe_1_0_4_N81, pe_1_0_4_N80, pe_1_0_4_N79,
         pe_1_0_4_N77, pe_1_0_4_N76, pe_1_0_4_N75, pe_1_0_4_N74, pe_1_0_4_N73,
         pe_1_0_4_N72, pe_1_0_4_N71, pe_1_0_4_N70, pe_1_0_4_int_data_0_,
         pe_1_0_4_int_data_1_, pe_1_0_4_int_data_2_, pe_1_0_4_int_data_3_,
         pe_1_0_4_N64, pe_1_0_4_N63, pe_1_0_4_N62, pe_1_0_4_N61, pe_1_0_4_N60,
         pe_1_0_4_N59, pe_1_0_4_o_data_v_0_, pe_1_0_4_o_data_v_1_,
         pe_1_0_4_o_data_v_2_, pe_1_0_4_o_data_v_3_, pe_1_0_5_n90,
         pe_1_0_5_n89, pe_1_0_5_n88, pe_1_0_5_n87, pe_1_0_5_n86, pe_1_0_5_n85,
         pe_1_0_5_n84, pe_1_0_5_n83, pe_1_0_5_n82, pe_1_0_5_n81, pe_1_0_5_n80,
         pe_1_0_5_n79, pe_1_0_5_n78, pe_1_0_5_n77, pe_1_0_5_n76, pe_1_0_5_n75,
         pe_1_0_5_n74, pe_1_0_5_n73, pe_1_0_5_n72, pe_1_0_5_n71, pe_1_0_5_n70,
         pe_1_0_5_n69, pe_1_0_5_n68, pe_1_0_5_n67, pe_1_0_5_n66, pe_1_0_5_n65,
         pe_1_0_5_n64, pe_1_0_5_n63, pe_1_0_5_n62, pe_1_0_5_n61, pe_1_0_5_n60,
         pe_1_0_5_n59, pe_1_0_5_n58, pe_1_0_5_n57, pe_1_0_5_n56, pe_1_0_5_n55,
         pe_1_0_5_n54, pe_1_0_5_n53, pe_1_0_5_n52, pe_1_0_5_n51, pe_1_0_5_n50,
         pe_1_0_5_n49, pe_1_0_5_n48, pe_1_0_5_n47, pe_1_0_5_n46, pe_1_0_5_n45,
         pe_1_0_5_n25, pe_1_0_5_n24, pe_1_0_5_n23, pe_1_0_5_n22, pe_1_0_5_n21,
         pe_1_0_5_n20, pe_1_0_5_n19, pe_1_0_5_n18, pe_1_0_5_n17, pe_1_0_5_n16,
         pe_1_0_5_n15, pe_1_0_5_n14, pe_1_0_5_n13, pe_1_0_5_n12, pe_1_0_5_n11,
         pe_1_0_5_n10, pe_1_0_5_n9, pe_1_0_5_n8, pe_1_0_5_n7, pe_1_0_5_n6,
         pe_1_0_5_n5, pe_1_0_5_n4, pe_1_0_5_n3, pe_1_0_5_n2, pe_1_0_5_n1,
         pe_1_0_5_n44, pe_1_0_5_n43, pe_1_0_5_n42, pe_1_0_5_n41, pe_1_0_5_n40,
         pe_1_0_5_n39, pe_1_0_5_n38, pe_1_0_5_n37, pe_1_0_5_n36, pe_1_0_5_n35,
         pe_1_0_5_n34, pe_1_0_5_n33, pe_1_0_5_n32, pe_1_0_5_n31, pe_1_0_5_n30,
         pe_1_0_5_n29, pe_1_0_5_n28, pe_1_0_5_n27, pe_1_0_5_n26,
         pe_1_0_5_net7162, pe_1_0_5_net7157, pe_1_0_5_net7152,
         pe_1_0_5_net7147, pe_1_0_5_net7142, pe_1_0_5_net7137,
         pe_1_0_5_net7132, pe_1_0_5_net7127, pe_1_0_5_net7122,
         pe_1_0_5_net7117, pe_1_0_5_net7112, pe_1_0_5_net7107,
         pe_1_0_5_net7101, pe_1_0_5_N90, pe_1_0_5_N85, pe_1_0_5_N84,
         pe_1_0_5_N83, pe_1_0_5_N82, pe_1_0_5_N81, pe_1_0_5_N80, pe_1_0_5_N79,
         pe_1_0_5_N77, pe_1_0_5_N76, pe_1_0_5_N75, pe_1_0_5_N74, pe_1_0_5_N73,
         pe_1_0_5_N72, pe_1_0_5_N71, pe_1_0_5_N70, pe_1_0_5_int_data_0_,
         pe_1_0_5_int_data_1_, pe_1_0_5_int_data_2_, pe_1_0_5_int_data_3_,
         pe_1_0_5_N64, pe_1_0_5_N63, pe_1_0_5_N62, pe_1_0_5_N61, pe_1_0_5_N60,
         pe_1_0_5_N59, pe_1_0_5_o_data_v_0_, pe_1_0_5_o_data_v_1_,
         pe_1_0_5_o_data_v_2_, pe_1_0_5_o_data_v_3_, pe_1_0_6_n90,
         pe_1_0_6_n89, pe_1_0_6_n88, pe_1_0_6_n87, pe_1_0_6_n86, pe_1_0_6_n85,
         pe_1_0_6_n84, pe_1_0_6_n83, pe_1_0_6_n82, pe_1_0_6_n81, pe_1_0_6_n80,
         pe_1_0_6_n79, pe_1_0_6_n78, pe_1_0_6_n77, pe_1_0_6_n76, pe_1_0_6_n75,
         pe_1_0_6_n74, pe_1_0_6_n73, pe_1_0_6_n72, pe_1_0_6_n71, pe_1_0_6_n70,
         pe_1_0_6_n69, pe_1_0_6_n68, pe_1_0_6_n67, pe_1_0_6_n66, pe_1_0_6_n65,
         pe_1_0_6_n64, pe_1_0_6_n63, pe_1_0_6_n62, pe_1_0_6_n61, pe_1_0_6_n60,
         pe_1_0_6_n59, pe_1_0_6_n58, pe_1_0_6_n57, pe_1_0_6_n56, pe_1_0_6_n55,
         pe_1_0_6_n54, pe_1_0_6_n53, pe_1_0_6_n52, pe_1_0_6_n51, pe_1_0_6_n50,
         pe_1_0_6_n49, pe_1_0_6_n48, pe_1_0_6_n47, pe_1_0_6_n46, pe_1_0_6_n45,
         pe_1_0_6_n25, pe_1_0_6_n24, pe_1_0_6_n23, pe_1_0_6_n22, pe_1_0_6_n21,
         pe_1_0_6_n20, pe_1_0_6_n19, pe_1_0_6_n18, pe_1_0_6_n17, pe_1_0_6_n16,
         pe_1_0_6_n15, pe_1_0_6_n14, pe_1_0_6_n13, pe_1_0_6_n12, pe_1_0_6_n11,
         pe_1_0_6_n10, pe_1_0_6_n9, pe_1_0_6_n8, pe_1_0_6_n7, pe_1_0_6_n6,
         pe_1_0_6_n5, pe_1_0_6_n4, pe_1_0_6_n3, pe_1_0_6_n2, pe_1_0_6_n1,
         pe_1_0_6_n44, pe_1_0_6_n43, pe_1_0_6_n42, pe_1_0_6_n41, pe_1_0_6_n40,
         pe_1_0_6_n39, pe_1_0_6_n38, pe_1_0_6_n37, pe_1_0_6_n36, pe_1_0_6_n35,
         pe_1_0_6_n34, pe_1_0_6_n33, pe_1_0_6_n32, pe_1_0_6_n31, pe_1_0_6_n30,
         pe_1_0_6_n29, pe_1_0_6_n28, pe_1_0_6_n27, pe_1_0_6_n26,
         pe_1_0_6_net7084, pe_1_0_6_net7079, pe_1_0_6_net7074,
         pe_1_0_6_net7069, pe_1_0_6_net7064, pe_1_0_6_net7059,
         pe_1_0_6_net7054, pe_1_0_6_net7049, pe_1_0_6_net7044,
         pe_1_0_6_net7039, pe_1_0_6_net7034, pe_1_0_6_net7029,
         pe_1_0_6_net7023, pe_1_0_6_N90, pe_1_0_6_N85, pe_1_0_6_N84,
         pe_1_0_6_N83, pe_1_0_6_N82, pe_1_0_6_N81, pe_1_0_6_N80, pe_1_0_6_N79,
         pe_1_0_6_N77, pe_1_0_6_N76, pe_1_0_6_N75, pe_1_0_6_N74, pe_1_0_6_N73,
         pe_1_0_6_N72, pe_1_0_6_N71, pe_1_0_6_N70, pe_1_0_6_int_data_0_,
         pe_1_0_6_int_data_1_, pe_1_0_6_int_data_2_, pe_1_0_6_int_data_3_,
         pe_1_0_6_N64, pe_1_0_6_N63, pe_1_0_6_N62, pe_1_0_6_N61, pe_1_0_6_N60,
         pe_1_0_6_N59, pe_1_0_6_o_data_v_0_, pe_1_0_6_o_data_v_1_,
         pe_1_0_6_o_data_v_2_, pe_1_0_6_o_data_v_3_, pe_1_0_7_n90,
         pe_1_0_7_n89, pe_1_0_7_n88, pe_1_0_7_n87, pe_1_0_7_n86, pe_1_0_7_n85,
         pe_1_0_7_n84, pe_1_0_7_n83, pe_1_0_7_n82, pe_1_0_7_n81, pe_1_0_7_n80,
         pe_1_0_7_n79, pe_1_0_7_n78, pe_1_0_7_n77, pe_1_0_7_n76, pe_1_0_7_n75,
         pe_1_0_7_n74, pe_1_0_7_n73, pe_1_0_7_n72, pe_1_0_7_n71, pe_1_0_7_n70,
         pe_1_0_7_n69, pe_1_0_7_n68, pe_1_0_7_n67, pe_1_0_7_n66, pe_1_0_7_n65,
         pe_1_0_7_n64, pe_1_0_7_n63, pe_1_0_7_n62, pe_1_0_7_n61, pe_1_0_7_n60,
         pe_1_0_7_n59, pe_1_0_7_n58, pe_1_0_7_n57, pe_1_0_7_n56, pe_1_0_7_n55,
         pe_1_0_7_n54, pe_1_0_7_n53, pe_1_0_7_n52, pe_1_0_7_n51, pe_1_0_7_n50,
         pe_1_0_7_n49, pe_1_0_7_n48, pe_1_0_7_n47, pe_1_0_7_n46, pe_1_0_7_n45,
         pe_1_0_7_n25, pe_1_0_7_n24, pe_1_0_7_n23, pe_1_0_7_n22, pe_1_0_7_n21,
         pe_1_0_7_n20, pe_1_0_7_n19, pe_1_0_7_n18, pe_1_0_7_n17, pe_1_0_7_n16,
         pe_1_0_7_n15, pe_1_0_7_n14, pe_1_0_7_n13, pe_1_0_7_n12, pe_1_0_7_n11,
         pe_1_0_7_n10, pe_1_0_7_n9, pe_1_0_7_n8, pe_1_0_7_n7, pe_1_0_7_n6,
         pe_1_0_7_n5, pe_1_0_7_n4, pe_1_0_7_n3, pe_1_0_7_n2, pe_1_0_7_n1,
         pe_1_0_7_n44, pe_1_0_7_n43, pe_1_0_7_n42, pe_1_0_7_n41, pe_1_0_7_n40,
         pe_1_0_7_n39, pe_1_0_7_n38, pe_1_0_7_n37, pe_1_0_7_n36, pe_1_0_7_n35,
         pe_1_0_7_n34, pe_1_0_7_n33, pe_1_0_7_n32, pe_1_0_7_n31, pe_1_0_7_n30,
         pe_1_0_7_n29, pe_1_0_7_n28, pe_1_0_7_n27, pe_1_0_7_n26,
         pe_1_0_7_net7006, pe_1_0_7_net7001, pe_1_0_7_net6996,
         pe_1_0_7_net6991, pe_1_0_7_net6986, pe_1_0_7_net6981,
         pe_1_0_7_net6976, pe_1_0_7_net6971, pe_1_0_7_net6966,
         pe_1_0_7_net6961, pe_1_0_7_net6956, pe_1_0_7_net6951,
         pe_1_0_7_net6945, pe_1_0_7_N90, pe_1_0_7_N85, pe_1_0_7_N84,
         pe_1_0_7_N83, pe_1_0_7_N82, pe_1_0_7_N81, pe_1_0_7_N80, pe_1_0_7_N79,
         pe_1_0_7_N77, pe_1_0_7_N76, pe_1_0_7_N75, pe_1_0_7_N74, pe_1_0_7_N73,
         pe_1_0_7_N72, pe_1_0_7_N71, pe_1_0_7_N70, pe_1_0_7_int_data_0_,
         pe_1_0_7_int_data_1_, pe_1_0_7_int_data_2_, pe_1_0_7_int_data_3_,
         pe_1_0_7_N64, pe_1_0_7_N63, pe_1_0_7_N62, pe_1_0_7_N61, pe_1_0_7_N60,
         pe_1_0_7_N59, pe_1_0_7_o_data_v_0_, pe_1_0_7_o_data_v_1_,
         pe_1_0_7_o_data_v_2_, pe_1_0_7_o_data_v_3_, pe_1_1_0_n90,
         pe_1_1_0_n89, pe_1_1_0_n88, pe_1_1_0_n87, pe_1_1_0_n86, pe_1_1_0_n85,
         pe_1_1_0_n84, pe_1_1_0_n83, pe_1_1_0_n82, pe_1_1_0_n81, pe_1_1_0_n80,
         pe_1_1_0_n79, pe_1_1_0_n78, pe_1_1_0_n77, pe_1_1_0_n76, pe_1_1_0_n75,
         pe_1_1_0_n74, pe_1_1_0_n73, pe_1_1_0_n72, pe_1_1_0_n71, pe_1_1_0_n70,
         pe_1_1_0_n69, pe_1_1_0_n68, pe_1_1_0_n67, pe_1_1_0_n66, pe_1_1_0_n65,
         pe_1_1_0_n64, pe_1_1_0_n63, pe_1_1_0_n62, pe_1_1_0_n61, pe_1_1_0_n60,
         pe_1_1_0_n59, pe_1_1_0_n58, pe_1_1_0_n57, pe_1_1_0_n56, pe_1_1_0_n55,
         pe_1_1_0_n54, pe_1_1_0_n53, pe_1_1_0_n52, pe_1_1_0_n51, pe_1_1_0_n50,
         pe_1_1_0_n49, pe_1_1_0_n48, pe_1_1_0_n47, pe_1_1_0_n46, pe_1_1_0_n45,
         pe_1_1_0_n25, pe_1_1_0_n24, pe_1_1_0_n23, pe_1_1_0_n22, pe_1_1_0_n21,
         pe_1_1_0_n20, pe_1_1_0_n19, pe_1_1_0_n18, pe_1_1_0_n17, pe_1_1_0_n16,
         pe_1_1_0_n15, pe_1_1_0_n14, pe_1_1_0_n13, pe_1_1_0_n12, pe_1_1_0_n11,
         pe_1_1_0_n10, pe_1_1_0_n9, pe_1_1_0_n8, pe_1_1_0_n7, pe_1_1_0_n6,
         pe_1_1_0_n5, pe_1_1_0_n4, pe_1_1_0_n3, pe_1_1_0_n2, pe_1_1_0_n1,
         pe_1_1_0_n44, pe_1_1_0_n43, pe_1_1_0_n42, pe_1_1_0_n41, pe_1_1_0_n40,
         pe_1_1_0_n39, pe_1_1_0_n38, pe_1_1_0_n37, pe_1_1_0_n36, pe_1_1_0_n35,
         pe_1_1_0_n34, pe_1_1_0_n33, pe_1_1_0_n32, pe_1_1_0_n31, pe_1_1_0_n30,
         pe_1_1_0_n29, pe_1_1_0_n28, pe_1_1_0_n27, pe_1_1_0_n26,
         pe_1_1_0_net6928, pe_1_1_0_net6923, pe_1_1_0_net6918,
         pe_1_1_0_net6913, pe_1_1_0_net6908, pe_1_1_0_net6903,
         pe_1_1_0_net6898, pe_1_1_0_net6893, pe_1_1_0_net6888,
         pe_1_1_0_net6883, pe_1_1_0_net6878, pe_1_1_0_net6873,
         pe_1_1_0_net6867, pe_1_1_0_N90, pe_1_1_0_N85, pe_1_1_0_N84,
         pe_1_1_0_N83, pe_1_1_0_N82, pe_1_1_0_N81, pe_1_1_0_N80, pe_1_1_0_N79,
         pe_1_1_0_N77, pe_1_1_0_N76, pe_1_1_0_N75, pe_1_1_0_N74, pe_1_1_0_N73,
         pe_1_1_0_N72, pe_1_1_0_N71, pe_1_1_0_N70, pe_1_1_0_int_data_0_,
         pe_1_1_0_int_data_1_, pe_1_1_0_int_data_2_, pe_1_1_0_int_data_3_,
         pe_1_1_0_N64, pe_1_1_0_N63, pe_1_1_0_N62, pe_1_1_0_N61, pe_1_1_0_N60,
         pe_1_1_0_N59, pe_1_1_0_o_data_h_0_, pe_1_1_0_o_data_h_1_,
         pe_1_1_0_o_data_h_2_, pe_1_1_0_o_data_h_3_, pe_1_1_1_n90,
         pe_1_1_1_n89, pe_1_1_1_n88, pe_1_1_1_n87, pe_1_1_1_n86, pe_1_1_1_n85,
         pe_1_1_1_n84, pe_1_1_1_n83, pe_1_1_1_n82, pe_1_1_1_n81, pe_1_1_1_n80,
         pe_1_1_1_n79, pe_1_1_1_n78, pe_1_1_1_n77, pe_1_1_1_n76, pe_1_1_1_n75,
         pe_1_1_1_n74, pe_1_1_1_n73, pe_1_1_1_n72, pe_1_1_1_n71, pe_1_1_1_n70,
         pe_1_1_1_n69, pe_1_1_1_n68, pe_1_1_1_n67, pe_1_1_1_n66, pe_1_1_1_n65,
         pe_1_1_1_n64, pe_1_1_1_n63, pe_1_1_1_n62, pe_1_1_1_n61, pe_1_1_1_n60,
         pe_1_1_1_n59, pe_1_1_1_n58, pe_1_1_1_n57, pe_1_1_1_n56, pe_1_1_1_n55,
         pe_1_1_1_n54, pe_1_1_1_n53, pe_1_1_1_n52, pe_1_1_1_n51, pe_1_1_1_n50,
         pe_1_1_1_n49, pe_1_1_1_n48, pe_1_1_1_n47, pe_1_1_1_n46, pe_1_1_1_n45,
         pe_1_1_1_n25, pe_1_1_1_n24, pe_1_1_1_n23, pe_1_1_1_n22, pe_1_1_1_n21,
         pe_1_1_1_n20, pe_1_1_1_n19, pe_1_1_1_n18, pe_1_1_1_n17, pe_1_1_1_n16,
         pe_1_1_1_n15, pe_1_1_1_n14, pe_1_1_1_n13, pe_1_1_1_n12, pe_1_1_1_n11,
         pe_1_1_1_n10, pe_1_1_1_n9, pe_1_1_1_n8, pe_1_1_1_n7, pe_1_1_1_n6,
         pe_1_1_1_n5, pe_1_1_1_n4, pe_1_1_1_n3, pe_1_1_1_n2, pe_1_1_1_n1,
         pe_1_1_1_n44, pe_1_1_1_n43, pe_1_1_1_n42, pe_1_1_1_n41, pe_1_1_1_n40,
         pe_1_1_1_n39, pe_1_1_1_n38, pe_1_1_1_n37, pe_1_1_1_n36, pe_1_1_1_n35,
         pe_1_1_1_n34, pe_1_1_1_n33, pe_1_1_1_n32, pe_1_1_1_n31, pe_1_1_1_n30,
         pe_1_1_1_n29, pe_1_1_1_n28, pe_1_1_1_n27, pe_1_1_1_n26,
         pe_1_1_1_net6850, pe_1_1_1_net6845, pe_1_1_1_net6840,
         pe_1_1_1_net6835, pe_1_1_1_net6830, pe_1_1_1_net6825,
         pe_1_1_1_net6820, pe_1_1_1_net6815, pe_1_1_1_net6810,
         pe_1_1_1_net6805, pe_1_1_1_net6800, pe_1_1_1_net6795,
         pe_1_1_1_net6789, pe_1_1_1_N90, pe_1_1_1_N85, pe_1_1_1_N84,
         pe_1_1_1_N83, pe_1_1_1_N82, pe_1_1_1_N81, pe_1_1_1_N80, pe_1_1_1_N79,
         pe_1_1_1_N77, pe_1_1_1_N76, pe_1_1_1_N75, pe_1_1_1_N74, pe_1_1_1_N73,
         pe_1_1_1_N72, pe_1_1_1_N71, pe_1_1_1_N70, pe_1_1_1_int_data_0_,
         pe_1_1_1_int_data_1_, pe_1_1_1_int_data_2_, pe_1_1_1_int_data_3_,
         pe_1_1_1_N64, pe_1_1_1_N63, pe_1_1_1_N62, pe_1_1_1_N61, pe_1_1_1_N60,
         pe_1_1_1_N59, pe_1_1_2_n90, pe_1_1_2_n89, pe_1_1_2_n88, pe_1_1_2_n87,
         pe_1_1_2_n86, pe_1_1_2_n85, pe_1_1_2_n84, pe_1_1_2_n83, pe_1_1_2_n82,
         pe_1_1_2_n81, pe_1_1_2_n80, pe_1_1_2_n79, pe_1_1_2_n78, pe_1_1_2_n77,
         pe_1_1_2_n76, pe_1_1_2_n75, pe_1_1_2_n74, pe_1_1_2_n73, pe_1_1_2_n72,
         pe_1_1_2_n71, pe_1_1_2_n70, pe_1_1_2_n69, pe_1_1_2_n68, pe_1_1_2_n67,
         pe_1_1_2_n66, pe_1_1_2_n65, pe_1_1_2_n64, pe_1_1_2_n63, pe_1_1_2_n62,
         pe_1_1_2_n61, pe_1_1_2_n60, pe_1_1_2_n59, pe_1_1_2_n58, pe_1_1_2_n57,
         pe_1_1_2_n56, pe_1_1_2_n55, pe_1_1_2_n54, pe_1_1_2_n53, pe_1_1_2_n52,
         pe_1_1_2_n51, pe_1_1_2_n50, pe_1_1_2_n49, pe_1_1_2_n48, pe_1_1_2_n47,
         pe_1_1_2_n46, pe_1_1_2_n45, pe_1_1_2_n25, pe_1_1_2_n24, pe_1_1_2_n23,
         pe_1_1_2_n22, pe_1_1_2_n21, pe_1_1_2_n20, pe_1_1_2_n19, pe_1_1_2_n18,
         pe_1_1_2_n17, pe_1_1_2_n16, pe_1_1_2_n15, pe_1_1_2_n14, pe_1_1_2_n13,
         pe_1_1_2_n12, pe_1_1_2_n11, pe_1_1_2_n10, pe_1_1_2_n9, pe_1_1_2_n8,
         pe_1_1_2_n7, pe_1_1_2_n6, pe_1_1_2_n5, pe_1_1_2_n4, pe_1_1_2_n3,
         pe_1_1_2_n2, pe_1_1_2_n1, pe_1_1_2_n44, pe_1_1_2_n43, pe_1_1_2_n42,
         pe_1_1_2_n41, pe_1_1_2_n40, pe_1_1_2_n39, pe_1_1_2_n38, pe_1_1_2_n37,
         pe_1_1_2_n36, pe_1_1_2_n35, pe_1_1_2_n34, pe_1_1_2_n33, pe_1_1_2_n32,
         pe_1_1_2_n31, pe_1_1_2_n30, pe_1_1_2_n29, pe_1_1_2_n28, pe_1_1_2_n27,
         pe_1_1_2_n26, pe_1_1_2_net6772, pe_1_1_2_net6767, pe_1_1_2_net6762,
         pe_1_1_2_net6757, pe_1_1_2_net6752, pe_1_1_2_net6747,
         pe_1_1_2_net6742, pe_1_1_2_net6737, pe_1_1_2_net6732,
         pe_1_1_2_net6727, pe_1_1_2_net6722, pe_1_1_2_net6717,
         pe_1_1_2_net6711, pe_1_1_2_N90, pe_1_1_2_N85, pe_1_1_2_N84,
         pe_1_1_2_N83, pe_1_1_2_N82, pe_1_1_2_N81, pe_1_1_2_N80, pe_1_1_2_N79,
         pe_1_1_2_N77, pe_1_1_2_N76, pe_1_1_2_N75, pe_1_1_2_N74, pe_1_1_2_N73,
         pe_1_1_2_N72, pe_1_1_2_N71, pe_1_1_2_N70, pe_1_1_2_int_data_0_,
         pe_1_1_2_int_data_1_, pe_1_1_2_int_data_2_, pe_1_1_2_int_data_3_,
         pe_1_1_2_N64, pe_1_1_2_N63, pe_1_1_2_N62, pe_1_1_2_N61, pe_1_1_2_N60,
         pe_1_1_2_N59, pe_1_1_3_n90, pe_1_1_3_n89, pe_1_1_3_n88, pe_1_1_3_n87,
         pe_1_1_3_n86, pe_1_1_3_n85, pe_1_1_3_n84, pe_1_1_3_n83, pe_1_1_3_n82,
         pe_1_1_3_n81, pe_1_1_3_n80, pe_1_1_3_n79, pe_1_1_3_n78, pe_1_1_3_n77,
         pe_1_1_3_n76, pe_1_1_3_n75, pe_1_1_3_n74, pe_1_1_3_n73, pe_1_1_3_n72,
         pe_1_1_3_n71, pe_1_1_3_n70, pe_1_1_3_n69, pe_1_1_3_n68, pe_1_1_3_n67,
         pe_1_1_3_n66, pe_1_1_3_n65, pe_1_1_3_n64, pe_1_1_3_n63, pe_1_1_3_n62,
         pe_1_1_3_n61, pe_1_1_3_n60, pe_1_1_3_n59, pe_1_1_3_n58, pe_1_1_3_n57,
         pe_1_1_3_n56, pe_1_1_3_n55, pe_1_1_3_n54, pe_1_1_3_n53, pe_1_1_3_n52,
         pe_1_1_3_n51, pe_1_1_3_n50, pe_1_1_3_n49, pe_1_1_3_n48, pe_1_1_3_n47,
         pe_1_1_3_n46, pe_1_1_3_n45, pe_1_1_3_n25, pe_1_1_3_n24, pe_1_1_3_n23,
         pe_1_1_3_n22, pe_1_1_3_n21, pe_1_1_3_n20, pe_1_1_3_n19, pe_1_1_3_n18,
         pe_1_1_3_n17, pe_1_1_3_n16, pe_1_1_3_n15, pe_1_1_3_n14, pe_1_1_3_n13,
         pe_1_1_3_n12, pe_1_1_3_n11, pe_1_1_3_n10, pe_1_1_3_n9, pe_1_1_3_n8,
         pe_1_1_3_n7, pe_1_1_3_n6, pe_1_1_3_n5, pe_1_1_3_n4, pe_1_1_3_n3,
         pe_1_1_3_n2, pe_1_1_3_n1, pe_1_1_3_n44, pe_1_1_3_n43, pe_1_1_3_n42,
         pe_1_1_3_n41, pe_1_1_3_n40, pe_1_1_3_n39, pe_1_1_3_n38, pe_1_1_3_n37,
         pe_1_1_3_n36, pe_1_1_3_n35, pe_1_1_3_n34, pe_1_1_3_n33, pe_1_1_3_n32,
         pe_1_1_3_n31, pe_1_1_3_n30, pe_1_1_3_n29, pe_1_1_3_n28, pe_1_1_3_n27,
         pe_1_1_3_n26, pe_1_1_3_net6694, pe_1_1_3_net6689, pe_1_1_3_net6684,
         pe_1_1_3_net6679, pe_1_1_3_net6674, pe_1_1_3_net6669,
         pe_1_1_3_net6664, pe_1_1_3_net6659, pe_1_1_3_net6654,
         pe_1_1_3_net6649, pe_1_1_3_net6644, pe_1_1_3_net6639,
         pe_1_1_3_net6633, pe_1_1_3_N90, pe_1_1_3_N85, pe_1_1_3_N84,
         pe_1_1_3_N83, pe_1_1_3_N82, pe_1_1_3_N81, pe_1_1_3_N80, pe_1_1_3_N79,
         pe_1_1_3_N77, pe_1_1_3_N76, pe_1_1_3_N75, pe_1_1_3_N74, pe_1_1_3_N73,
         pe_1_1_3_N72, pe_1_1_3_N71, pe_1_1_3_N70, pe_1_1_3_int_data_0_,
         pe_1_1_3_int_data_1_, pe_1_1_3_int_data_2_, pe_1_1_3_int_data_3_,
         pe_1_1_3_N64, pe_1_1_3_N63, pe_1_1_3_N62, pe_1_1_3_N61, pe_1_1_3_N60,
         pe_1_1_3_N59, pe_1_1_4_n86, pe_1_1_4_n85, pe_1_1_4_n84, pe_1_1_4_n83,
         pe_1_1_4_n82, pe_1_1_4_n81, pe_1_1_4_n80, pe_1_1_4_n79, pe_1_1_4_n78,
         pe_1_1_4_n77, pe_1_1_4_n76, pe_1_1_4_n75, pe_1_1_4_n74, pe_1_1_4_n73,
         pe_1_1_4_n72, pe_1_1_4_n71, pe_1_1_4_n70, pe_1_1_4_n69, pe_1_1_4_n68,
         pe_1_1_4_n67, pe_1_1_4_n66, pe_1_1_4_n65, pe_1_1_4_n64, pe_1_1_4_n63,
         pe_1_1_4_n62, pe_1_1_4_n61, pe_1_1_4_n60, pe_1_1_4_n59, pe_1_1_4_n58,
         pe_1_1_4_n57, pe_1_1_4_n56, pe_1_1_4_n55, pe_1_1_4_n54, pe_1_1_4_n53,
         pe_1_1_4_n52, pe_1_1_4_n51, pe_1_1_4_n50, pe_1_1_4_n49, pe_1_1_4_n48,
         pe_1_1_4_n47, pe_1_1_4_n46, pe_1_1_4_n45, pe_1_1_4_n25, pe_1_1_4_n24,
         pe_1_1_4_n23, pe_1_1_4_n22, pe_1_1_4_n21, pe_1_1_4_n20, pe_1_1_4_n19,
         pe_1_1_4_n18, pe_1_1_4_n17, pe_1_1_4_n16, pe_1_1_4_n15, pe_1_1_4_n14,
         pe_1_1_4_n13, pe_1_1_4_n12, pe_1_1_4_n11, pe_1_1_4_n10, pe_1_1_4_n9,
         pe_1_1_4_n8, pe_1_1_4_n7, pe_1_1_4_n6, pe_1_1_4_n5, pe_1_1_4_n4,
         pe_1_1_4_n3, pe_1_1_4_n2, pe_1_1_4_n1, pe_1_1_4_n44, pe_1_1_4_n43,
         pe_1_1_4_n42, pe_1_1_4_n41, pe_1_1_4_n40, pe_1_1_4_n39, pe_1_1_4_n38,
         pe_1_1_4_n37, pe_1_1_4_n36, pe_1_1_4_n35, pe_1_1_4_n34, pe_1_1_4_n33,
         pe_1_1_4_n32, pe_1_1_4_n31, pe_1_1_4_n30, pe_1_1_4_n29, pe_1_1_4_n28,
         pe_1_1_4_n27, pe_1_1_4_n26, pe_1_1_4_net6616, pe_1_1_4_net6611,
         pe_1_1_4_net6606, pe_1_1_4_net6601, pe_1_1_4_net6596,
         pe_1_1_4_net6591, pe_1_1_4_net6586, pe_1_1_4_net6581,
         pe_1_1_4_net6576, pe_1_1_4_net6571, pe_1_1_4_net6566,
         pe_1_1_4_net6561, pe_1_1_4_net6555, pe_1_1_4_N90, pe_1_1_4_N85,
         pe_1_1_4_N84, pe_1_1_4_N83, pe_1_1_4_N82, pe_1_1_4_N81, pe_1_1_4_N80,
         pe_1_1_4_N79, pe_1_1_4_N77, pe_1_1_4_N76, pe_1_1_4_N75, pe_1_1_4_N74,
         pe_1_1_4_N73, pe_1_1_4_N72, pe_1_1_4_N71, pe_1_1_4_N70,
         pe_1_1_4_int_data_0_, pe_1_1_4_int_data_1_, pe_1_1_4_int_data_2_,
         pe_1_1_4_int_data_3_, pe_1_1_4_N64, pe_1_1_4_N63, pe_1_1_4_N62,
         pe_1_1_4_N61, pe_1_1_4_N60, pe_1_1_4_N59, pe_1_1_5_n87, pe_1_1_5_n86,
         pe_1_1_5_n85, pe_1_1_5_n84, pe_1_1_5_n83, pe_1_1_5_n82, pe_1_1_5_n81,
         pe_1_1_5_n80, pe_1_1_5_n79, pe_1_1_5_n78, pe_1_1_5_n77, pe_1_1_5_n76,
         pe_1_1_5_n75, pe_1_1_5_n74, pe_1_1_5_n73, pe_1_1_5_n72, pe_1_1_5_n71,
         pe_1_1_5_n70, pe_1_1_5_n69, pe_1_1_5_n68, pe_1_1_5_n67, pe_1_1_5_n66,
         pe_1_1_5_n65, pe_1_1_5_n64, pe_1_1_5_n63, pe_1_1_5_n62, pe_1_1_5_n61,
         pe_1_1_5_n60, pe_1_1_5_n59, pe_1_1_5_n58, pe_1_1_5_n57, pe_1_1_5_n56,
         pe_1_1_5_n55, pe_1_1_5_n54, pe_1_1_5_n53, pe_1_1_5_n52, pe_1_1_5_n51,
         pe_1_1_5_n50, pe_1_1_5_n49, pe_1_1_5_n48, pe_1_1_5_n47, pe_1_1_5_n46,
         pe_1_1_5_n45, pe_1_1_5_n25, pe_1_1_5_n24, pe_1_1_5_n23, pe_1_1_5_n22,
         pe_1_1_5_n21, pe_1_1_5_n20, pe_1_1_5_n19, pe_1_1_5_n18, pe_1_1_5_n17,
         pe_1_1_5_n16, pe_1_1_5_n15, pe_1_1_5_n14, pe_1_1_5_n13, pe_1_1_5_n12,
         pe_1_1_5_n11, pe_1_1_5_n10, pe_1_1_5_n9, pe_1_1_5_n8, pe_1_1_5_n7,
         pe_1_1_5_n6, pe_1_1_5_n5, pe_1_1_5_n4, pe_1_1_5_n3, pe_1_1_5_n2,
         pe_1_1_5_n1, pe_1_1_5_n44, pe_1_1_5_n43, pe_1_1_5_n42, pe_1_1_5_n41,
         pe_1_1_5_n40, pe_1_1_5_n39, pe_1_1_5_n38, pe_1_1_5_n37, pe_1_1_5_n36,
         pe_1_1_5_n35, pe_1_1_5_n34, pe_1_1_5_n33, pe_1_1_5_n32, pe_1_1_5_n31,
         pe_1_1_5_n30, pe_1_1_5_n29, pe_1_1_5_n28, pe_1_1_5_n27, pe_1_1_5_n26,
         pe_1_1_5_net6538, pe_1_1_5_net6533, pe_1_1_5_net6528,
         pe_1_1_5_net6523, pe_1_1_5_net6518, pe_1_1_5_net6513,
         pe_1_1_5_net6508, pe_1_1_5_net6503, pe_1_1_5_net6498,
         pe_1_1_5_net6493, pe_1_1_5_net6488, pe_1_1_5_net6483,
         pe_1_1_5_net6477, pe_1_1_5_N90, pe_1_1_5_N85, pe_1_1_5_N84,
         pe_1_1_5_N83, pe_1_1_5_N82, pe_1_1_5_N81, pe_1_1_5_N80, pe_1_1_5_N79,
         pe_1_1_5_N77, pe_1_1_5_N76, pe_1_1_5_N75, pe_1_1_5_N74, pe_1_1_5_N73,
         pe_1_1_5_N72, pe_1_1_5_N71, pe_1_1_5_N70, pe_1_1_5_int_data_0_,
         pe_1_1_5_int_data_1_, pe_1_1_5_int_data_2_, pe_1_1_5_int_data_3_,
         pe_1_1_5_N64, pe_1_1_5_N63, pe_1_1_5_N62, pe_1_1_5_N61, pe_1_1_5_N60,
         pe_1_1_5_N59, pe_1_1_6_n88, pe_1_1_6_n87, pe_1_1_6_n86, pe_1_1_6_n85,
         pe_1_1_6_n84, pe_1_1_6_n83, pe_1_1_6_n82, pe_1_1_6_n81, pe_1_1_6_n80,
         pe_1_1_6_n79, pe_1_1_6_n78, pe_1_1_6_n77, pe_1_1_6_n76, pe_1_1_6_n75,
         pe_1_1_6_n74, pe_1_1_6_n73, pe_1_1_6_n72, pe_1_1_6_n71, pe_1_1_6_n70,
         pe_1_1_6_n69, pe_1_1_6_n68, pe_1_1_6_n67, pe_1_1_6_n66, pe_1_1_6_n65,
         pe_1_1_6_n64, pe_1_1_6_n63, pe_1_1_6_n62, pe_1_1_6_n61, pe_1_1_6_n60,
         pe_1_1_6_n59, pe_1_1_6_n58, pe_1_1_6_n57, pe_1_1_6_n56, pe_1_1_6_n55,
         pe_1_1_6_n54, pe_1_1_6_n53, pe_1_1_6_n52, pe_1_1_6_n51, pe_1_1_6_n50,
         pe_1_1_6_n49, pe_1_1_6_n48, pe_1_1_6_n47, pe_1_1_6_n46, pe_1_1_6_n45,
         pe_1_1_6_n25, pe_1_1_6_n24, pe_1_1_6_n23, pe_1_1_6_n22, pe_1_1_6_n21,
         pe_1_1_6_n20, pe_1_1_6_n19, pe_1_1_6_n18, pe_1_1_6_n17, pe_1_1_6_n16,
         pe_1_1_6_n15, pe_1_1_6_n14, pe_1_1_6_n13, pe_1_1_6_n12, pe_1_1_6_n11,
         pe_1_1_6_n10, pe_1_1_6_n9, pe_1_1_6_n8, pe_1_1_6_n7, pe_1_1_6_n6,
         pe_1_1_6_n5, pe_1_1_6_n4, pe_1_1_6_n3, pe_1_1_6_n2, pe_1_1_6_n1,
         pe_1_1_6_n44, pe_1_1_6_n43, pe_1_1_6_n42, pe_1_1_6_n41, pe_1_1_6_n40,
         pe_1_1_6_n39, pe_1_1_6_n38, pe_1_1_6_n37, pe_1_1_6_n36, pe_1_1_6_n35,
         pe_1_1_6_n34, pe_1_1_6_n33, pe_1_1_6_n32, pe_1_1_6_n31, pe_1_1_6_n30,
         pe_1_1_6_n29, pe_1_1_6_n28, pe_1_1_6_n27, pe_1_1_6_n26,
         pe_1_1_6_net6460, pe_1_1_6_net6455, pe_1_1_6_net6450,
         pe_1_1_6_net6445, pe_1_1_6_net6440, pe_1_1_6_net6435,
         pe_1_1_6_net6430, pe_1_1_6_net6425, pe_1_1_6_net6420,
         pe_1_1_6_net6415, pe_1_1_6_net6410, pe_1_1_6_net6405,
         pe_1_1_6_net6399, pe_1_1_6_N90, pe_1_1_6_N85, pe_1_1_6_N84,
         pe_1_1_6_N83, pe_1_1_6_N82, pe_1_1_6_N81, pe_1_1_6_N80, pe_1_1_6_N79,
         pe_1_1_6_N77, pe_1_1_6_N76, pe_1_1_6_N75, pe_1_1_6_N74, pe_1_1_6_N73,
         pe_1_1_6_N72, pe_1_1_6_N71, pe_1_1_6_N70, pe_1_1_6_int_data_0_,
         pe_1_1_6_int_data_1_, pe_1_1_6_int_data_2_, pe_1_1_6_int_data_3_,
         pe_1_1_6_N64, pe_1_1_6_N63, pe_1_1_6_N62, pe_1_1_6_N61, pe_1_1_6_N60,
         pe_1_1_6_N59, pe_1_1_7_n88, pe_1_1_7_n87, pe_1_1_7_n86, pe_1_1_7_n85,
         pe_1_1_7_n84, pe_1_1_7_n83, pe_1_1_7_n82, pe_1_1_7_n81, pe_1_1_7_n80,
         pe_1_1_7_n79, pe_1_1_7_n78, pe_1_1_7_n77, pe_1_1_7_n76, pe_1_1_7_n75,
         pe_1_1_7_n74, pe_1_1_7_n73, pe_1_1_7_n72, pe_1_1_7_n71, pe_1_1_7_n70,
         pe_1_1_7_n69, pe_1_1_7_n68, pe_1_1_7_n67, pe_1_1_7_n66, pe_1_1_7_n65,
         pe_1_1_7_n64, pe_1_1_7_n63, pe_1_1_7_n62, pe_1_1_7_n61, pe_1_1_7_n60,
         pe_1_1_7_n59, pe_1_1_7_n58, pe_1_1_7_n57, pe_1_1_7_n56, pe_1_1_7_n55,
         pe_1_1_7_n54, pe_1_1_7_n53, pe_1_1_7_n52, pe_1_1_7_n51, pe_1_1_7_n50,
         pe_1_1_7_n49, pe_1_1_7_n48, pe_1_1_7_n47, pe_1_1_7_n46, pe_1_1_7_n45,
         pe_1_1_7_n25, pe_1_1_7_n24, pe_1_1_7_n23, pe_1_1_7_n22, pe_1_1_7_n21,
         pe_1_1_7_n20, pe_1_1_7_n19, pe_1_1_7_n18, pe_1_1_7_n17, pe_1_1_7_n16,
         pe_1_1_7_n15, pe_1_1_7_n14, pe_1_1_7_n13, pe_1_1_7_n12, pe_1_1_7_n11,
         pe_1_1_7_n10, pe_1_1_7_n9, pe_1_1_7_n8, pe_1_1_7_n7, pe_1_1_7_n6,
         pe_1_1_7_n5, pe_1_1_7_n4, pe_1_1_7_n3, pe_1_1_7_n2, pe_1_1_7_n1,
         pe_1_1_7_n44, pe_1_1_7_n43, pe_1_1_7_n42, pe_1_1_7_n41, pe_1_1_7_n40,
         pe_1_1_7_n39, pe_1_1_7_n38, pe_1_1_7_n37, pe_1_1_7_n36, pe_1_1_7_n35,
         pe_1_1_7_n34, pe_1_1_7_n33, pe_1_1_7_n32, pe_1_1_7_n31, pe_1_1_7_n30,
         pe_1_1_7_n29, pe_1_1_7_n28, pe_1_1_7_n27, pe_1_1_7_n26,
         pe_1_1_7_net6382, pe_1_1_7_net6377, pe_1_1_7_net6372,
         pe_1_1_7_net6367, pe_1_1_7_net6362, pe_1_1_7_net6357,
         pe_1_1_7_net6352, pe_1_1_7_net6347, pe_1_1_7_net6342,
         pe_1_1_7_net6337, pe_1_1_7_net6332, pe_1_1_7_net6327,
         pe_1_1_7_net6321, pe_1_1_7_N90, pe_1_1_7_N85, pe_1_1_7_N84,
         pe_1_1_7_N83, pe_1_1_7_N82, pe_1_1_7_N81, pe_1_1_7_N80, pe_1_1_7_N79,
         pe_1_1_7_N77, pe_1_1_7_N76, pe_1_1_7_N75, pe_1_1_7_N74, pe_1_1_7_N73,
         pe_1_1_7_N72, pe_1_1_7_N71, pe_1_1_7_N70, pe_1_1_7_int_data_0_,
         pe_1_1_7_int_data_1_, pe_1_1_7_int_data_2_, pe_1_1_7_int_data_3_,
         pe_1_1_7_N64, pe_1_1_7_N63, pe_1_1_7_N62, pe_1_1_7_N61, pe_1_1_7_N60,
         pe_1_1_7_N59, pe_1_2_0_n89, pe_1_2_0_n88, pe_1_2_0_n87, pe_1_2_0_n86,
         pe_1_2_0_n85, pe_1_2_0_n84, pe_1_2_0_n83, pe_1_2_0_n82, pe_1_2_0_n81,
         pe_1_2_0_n80, pe_1_2_0_n79, pe_1_2_0_n78, pe_1_2_0_n77, pe_1_2_0_n76,
         pe_1_2_0_n75, pe_1_2_0_n74, pe_1_2_0_n73, pe_1_2_0_n72, pe_1_2_0_n71,
         pe_1_2_0_n70, pe_1_2_0_n69, pe_1_2_0_n68, pe_1_2_0_n67, pe_1_2_0_n66,
         pe_1_2_0_n65, pe_1_2_0_n64, pe_1_2_0_n63, pe_1_2_0_n62, pe_1_2_0_n61,
         pe_1_2_0_n60, pe_1_2_0_n59, pe_1_2_0_n58, pe_1_2_0_n57, pe_1_2_0_n56,
         pe_1_2_0_n55, pe_1_2_0_n54, pe_1_2_0_n53, pe_1_2_0_n52, pe_1_2_0_n51,
         pe_1_2_0_n50, pe_1_2_0_n49, pe_1_2_0_n48, pe_1_2_0_n47, pe_1_2_0_n46,
         pe_1_2_0_n45, pe_1_2_0_n25, pe_1_2_0_n24, pe_1_2_0_n23, pe_1_2_0_n22,
         pe_1_2_0_n21, pe_1_2_0_n20, pe_1_2_0_n19, pe_1_2_0_n18, pe_1_2_0_n17,
         pe_1_2_0_n16, pe_1_2_0_n15, pe_1_2_0_n14, pe_1_2_0_n13, pe_1_2_0_n12,
         pe_1_2_0_n11, pe_1_2_0_n10, pe_1_2_0_n9, pe_1_2_0_n8, pe_1_2_0_n7,
         pe_1_2_0_n6, pe_1_2_0_n5, pe_1_2_0_n4, pe_1_2_0_n3, pe_1_2_0_n2,
         pe_1_2_0_n1, pe_1_2_0_n44, pe_1_2_0_n43, pe_1_2_0_n42, pe_1_2_0_n41,
         pe_1_2_0_n40, pe_1_2_0_n39, pe_1_2_0_n38, pe_1_2_0_n37, pe_1_2_0_n36,
         pe_1_2_0_n35, pe_1_2_0_n34, pe_1_2_0_n33, pe_1_2_0_n32, pe_1_2_0_n31,
         pe_1_2_0_n30, pe_1_2_0_n29, pe_1_2_0_n28, pe_1_2_0_n27, pe_1_2_0_n26,
         pe_1_2_0_net6304, pe_1_2_0_net6299, pe_1_2_0_net6294,
         pe_1_2_0_net6289, pe_1_2_0_net6284, pe_1_2_0_net6279,
         pe_1_2_0_net6274, pe_1_2_0_net6269, pe_1_2_0_net6264,
         pe_1_2_0_net6259, pe_1_2_0_net6254, pe_1_2_0_net6249,
         pe_1_2_0_net6243, pe_1_2_0_N90, pe_1_2_0_N85, pe_1_2_0_N84,
         pe_1_2_0_N83, pe_1_2_0_N82, pe_1_2_0_N81, pe_1_2_0_N80, pe_1_2_0_N79,
         pe_1_2_0_N77, pe_1_2_0_N76, pe_1_2_0_N75, pe_1_2_0_N74, pe_1_2_0_N73,
         pe_1_2_0_N72, pe_1_2_0_N71, pe_1_2_0_N70, pe_1_2_0_int_data_0_,
         pe_1_2_0_int_data_1_, pe_1_2_0_int_data_2_, pe_1_2_0_int_data_3_,
         pe_1_2_0_N64, pe_1_2_0_N63, pe_1_2_0_N62, pe_1_2_0_N61, pe_1_2_0_N60,
         pe_1_2_0_N59, pe_1_2_0_o_data_h_0_, pe_1_2_0_o_data_h_1_,
         pe_1_2_0_o_data_h_2_, pe_1_2_0_o_data_h_3_, pe_1_2_1_n90,
         pe_1_2_1_n89, pe_1_2_1_n88, pe_1_2_1_n87, pe_1_2_1_n86, pe_1_2_1_n85,
         pe_1_2_1_n84, pe_1_2_1_n83, pe_1_2_1_n82, pe_1_2_1_n81, pe_1_2_1_n80,
         pe_1_2_1_n79, pe_1_2_1_n78, pe_1_2_1_n77, pe_1_2_1_n76, pe_1_2_1_n75,
         pe_1_2_1_n74, pe_1_2_1_n73, pe_1_2_1_n72, pe_1_2_1_n71, pe_1_2_1_n70,
         pe_1_2_1_n69, pe_1_2_1_n68, pe_1_2_1_n67, pe_1_2_1_n66, pe_1_2_1_n65,
         pe_1_2_1_n64, pe_1_2_1_n63, pe_1_2_1_n62, pe_1_2_1_n61, pe_1_2_1_n60,
         pe_1_2_1_n59, pe_1_2_1_n58, pe_1_2_1_n57, pe_1_2_1_n56, pe_1_2_1_n55,
         pe_1_2_1_n54, pe_1_2_1_n53, pe_1_2_1_n52, pe_1_2_1_n51, pe_1_2_1_n50,
         pe_1_2_1_n49, pe_1_2_1_n48, pe_1_2_1_n47, pe_1_2_1_n46, pe_1_2_1_n45,
         pe_1_2_1_n25, pe_1_2_1_n24, pe_1_2_1_n23, pe_1_2_1_n22, pe_1_2_1_n21,
         pe_1_2_1_n20, pe_1_2_1_n19, pe_1_2_1_n18, pe_1_2_1_n17, pe_1_2_1_n16,
         pe_1_2_1_n15, pe_1_2_1_n14, pe_1_2_1_n13, pe_1_2_1_n12, pe_1_2_1_n11,
         pe_1_2_1_n10, pe_1_2_1_n9, pe_1_2_1_n8, pe_1_2_1_n7, pe_1_2_1_n6,
         pe_1_2_1_n5, pe_1_2_1_n4, pe_1_2_1_n3, pe_1_2_1_n2, pe_1_2_1_n1,
         pe_1_2_1_n44, pe_1_2_1_n43, pe_1_2_1_n42, pe_1_2_1_n41, pe_1_2_1_n40,
         pe_1_2_1_n39, pe_1_2_1_n38, pe_1_2_1_n37, pe_1_2_1_n36, pe_1_2_1_n35,
         pe_1_2_1_n34, pe_1_2_1_n33, pe_1_2_1_n32, pe_1_2_1_n31, pe_1_2_1_n30,
         pe_1_2_1_n29, pe_1_2_1_n28, pe_1_2_1_n27, pe_1_2_1_n26,
         pe_1_2_1_net6226, pe_1_2_1_net6221, pe_1_2_1_net6216,
         pe_1_2_1_net6211, pe_1_2_1_net6206, pe_1_2_1_net6201,
         pe_1_2_1_net6196, pe_1_2_1_net6191, pe_1_2_1_net6186,
         pe_1_2_1_net6181, pe_1_2_1_net6176, pe_1_2_1_net6171,
         pe_1_2_1_net6165, pe_1_2_1_N90, pe_1_2_1_N85, pe_1_2_1_N84,
         pe_1_2_1_N83, pe_1_2_1_N82, pe_1_2_1_N81, pe_1_2_1_N80, pe_1_2_1_N79,
         pe_1_2_1_N77, pe_1_2_1_N76, pe_1_2_1_N75, pe_1_2_1_N74, pe_1_2_1_N73,
         pe_1_2_1_N72, pe_1_2_1_N71, pe_1_2_1_N70, pe_1_2_1_int_data_0_,
         pe_1_2_1_int_data_1_, pe_1_2_1_int_data_2_, pe_1_2_1_int_data_3_,
         pe_1_2_1_N64, pe_1_2_1_N63, pe_1_2_1_N62, pe_1_2_1_N61, pe_1_2_1_N60,
         pe_1_2_1_N59, pe_1_2_2_n90, pe_1_2_2_n89, pe_1_2_2_n88, pe_1_2_2_n87,
         pe_1_2_2_n86, pe_1_2_2_n85, pe_1_2_2_n84, pe_1_2_2_n83, pe_1_2_2_n82,
         pe_1_2_2_n81, pe_1_2_2_n80, pe_1_2_2_n79, pe_1_2_2_n78, pe_1_2_2_n77,
         pe_1_2_2_n76, pe_1_2_2_n75, pe_1_2_2_n74, pe_1_2_2_n73, pe_1_2_2_n72,
         pe_1_2_2_n71, pe_1_2_2_n70, pe_1_2_2_n69, pe_1_2_2_n68, pe_1_2_2_n67,
         pe_1_2_2_n66, pe_1_2_2_n65, pe_1_2_2_n64, pe_1_2_2_n63, pe_1_2_2_n62,
         pe_1_2_2_n61, pe_1_2_2_n60, pe_1_2_2_n59, pe_1_2_2_n58, pe_1_2_2_n57,
         pe_1_2_2_n56, pe_1_2_2_n55, pe_1_2_2_n54, pe_1_2_2_n53, pe_1_2_2_n52,
         pe_1_2_2_n51, pe_1_2_2_n50, pe_1_2_2_n49, pe_1_2_2_n48, pe_1_2_2_n47,
         pe_1_2_2_n46, pe_1_2_2_n45, pe_1_2_2_n25, pe_1_2_2_n24, pe_1_2_2_n23,
         pe_1_2_2_n22, pe_1_2_2_n21, pe_1_2_2_n20, pe_1_2_2_n19, pe_1_2_2_n18,
         pe_1_2_2_n17, pe_1_2_2_n16, pe_1_2_2_n15, pe_1_2_2_n14, pe_1_2_2_n13,
         pe_1_2_2_n12, pe_1_2_2_n11, pe_1_2_2_n10, pe_1_2_2_n9, pe_1_2_2_n8,
         pe_1_2_2_n7, pe_1_2_2_n6, pe_1_2_2_n5, pe_1_2_2_n4, pe_1_2_2_n3,
         pe_1_2_2_n2, pe_1_2_2_n1, pe_1_2_2_n44, pe_1_2_2_n43, pe_1_2_2_n42,
         pe_1_2_2_n41, pe_1_2_2_n40, pe_1_2_2_n39, pe_1_2_2_n38, pe_1_2_2_n37,
         pe_1_2_2_n36, pe_1_2_2_n35, pe_1_2_2_n34, pe_1_2_2_n33, pe_1_2_2_n32,
         pe_1_2_2_n31, pe_1_2_2_n30, pe_1_2_2_n29, pe_1_2_2_n28, pe_1_2_2_n27,
         pe_1_2_2_n26, pe_1_2_2_net6148, pe_1_2_2_net6143, pe_1_2_2_net6138,
         pe_1_2_2_net6133, pe_1_2_2_net6128, pe_1_2_2_net6123,
         pe_1_2_2_net6118, pe_1_2_2_net6113, pe_1_2_2_net6108,
         pe_1_2_2_net6103, pe_1_2_2_net6098, pe_1_2_2_net6093,
         pe_1_2_2_net6087, pe_1_2_2_N90, pe_1_2_2_N85, pe_1_2_2_N84,
         pe_1_2_2_N83, pe_1_2_2_N82, pe_1_2_2_N81, pe_1_2_2_N80, pe_1_2_2_N79,
         pe_1_2_2_N77, pe_1_2_2_N76, pe_1_2_2_N75, pe_1_2_2_N74, pe_1_2_2_N73,
         pe_1_2_2_N72, pe_1_2_2_N71, pe_1_2_2_N70, pe_1_2_2_int_data_0_,
         pe_1_2_2_int_data_1_, pe_1_2_2_int_data_2_, pe_1_2_2_int_data_3_,
         pe_1_2_2_N64, pe_1_2_2_N63, pe_1_2_2_N62, pe_1_2_2_N61, pe_1_2_2_N60,
         pe_1_2_2_N59, pe_1_2_3_n90, pe_1_2_3_n89, pe_1_2_3_n88, pe_1_2_3_n87,
         pe_1_2_3_n86, pe_1_2_3_n85, pe_1_2_3_n84, pe_1_2_3_n83, pe_1_2_3_n82,
         pe_1_2_3_n81, pe_1_2_3_n80, pe_1_2_3_n79, pe_1_2_3_n78, pe_1_2_3_n77,
         pe_1_2_3_n76, pe_1_2_3_n75, pe_1_2_3_n74, pe_1_2_3_n73, pe_1_2_3_n72,
         pe_1_2_3_n71, pe_1_2_3_n70, pe_1_2_3_n69, pe_1_2_3_n68, pe_1_2_3_n67,
         pe_1_2_3_n66, pe_1_2_3_n65, pe_1_2_3_n64, pe_1_2_3_n63, pe_1_2_3_n62,
         pe_1_2_3_n61, pe_1_2_3_n60, pe_1_2_3_n59, pe_1_2_3_n58, pe_1_2_3_n57,
         pe_1_2_3_n56, pe_1_2_3_n55, pe_1_2_3_n54, pe_1_2_3_n53, pe_1_2_3_n52,
         pe_1_2_3_n51, pe_1_2_3_n50, pe_1_2_3_n49, pe_1_2_3_n48, pe_1_2_3_n47,
         pe_1_2_3_n46, pe_1_2_3_n45, pe_1_2_3_n25, pe_1_2_3_n24, pe_1_2_3_n23,
         pe_1_2_3_n22, pe_1_2_3_n21, pe_1_2_3_n20, pe_1_2_3_n19, pe_1_2_3_n18,
         pe_1_2_3_n17, pe_1_2_3_n16, pe_1_2_3_n15, pe_1_2_3_n14, pe_1_2_3_n13,
         pe_1_2_3_n12, pe_1_2_3_n11, pe_1_2_3_n10, pe_1_2_3_n9, pe_1_2_3_n8,
         pe_1_2_3_n7, pe_1_2_3_n6, pe_1_2_3_n5, pe_1_2_3_n4, pe_1_2_3_n3,
         pe_1_2_3_n2, pe_1_2_3_n1, pe_1_2_3_n44, pe_1_2_3_n43, pe_1_2_3_n42,
         pe_1_2_3_n41, pe_1_2_3_n40, pe_1_2_3_n39, pe_1_2_3_n38, pe_1_2_3_n37,
         pe_1_2_3_n36, pe_1_2_3_n35, pe_1_2_3_n34, pe_1_2_3_n33, pe_1_2_3_n32,
         pe_1_2_3_n31, pe_1_2_3_n30, pe_1_2_3_n29, pe_1_2_3_n28, pe_1_2_3_n27,
         pe_1_2_3_n26, pe_1_2_3_net6070, pe_1_2_3_net6065, pe_1_2_3_net6060,
         pe_1_2_3_net6055, pe_1_2_3_net6050, pe_1_2_3_net6045,
         pe_1_2_3_net6040, pe_1_2_3_net6035, pe_1_2_3_net6030,
         pe_1_2_3_net6025, pe_1_2_3_net6020, pe_1_2_3_net6015,
         pe_1_2_3_net6009, pe_1_2_3_N90, pe_1_2_3_N85, pe_1_2_3_N84,
         pe_1_2_3_N83, pe_1_2_3_N82, pe_1_2_3_N81, pe_1_2_3_N80, pe_1_2_3_N79,
         pe_1_2_3_N77, pe_1_2_3_N76, pe_1_2_3_N75, pe_1_2_3_N74, pe_1_2_3_N73,
         pe_1_2_3_N72, pe_1_2_3_N71, pe_1_2_3_N70, pe_1_2_3_int_data_0_,
         pe_1_2_3_int_data_1_, pe_1_2_3_int_data_2_, pe_1_2_3_int_data_3_,
         pe_1_2_3_N64, pe_1_2_3_N63, pe_1_2_3_N62, pe_1_2_3_N61, pe_1_2_3_N60,
         pe_1_2_3_N59, pe_1_2_4_n90, pe_1_2_4_n89, pe_1_2_4_n88, pe_1_2_4_n87,
         pe_1_2_4_n86, pe_1_2_4_n85, pe_1_2_4_n84, pe_1_2_4_n83, pe_1_2_4_n82,
         pe_1_2_4_n81, pe_1_2_4_n80, pe_1_2_4_n79, pe_1_2_4_n78, pe_1_2_4_n77,
         pe_1_2_4_n76, pe_1_2_4_n75, pe_1_2_4_n74, pe_1_2_4_n73, pe_1_2_4_n72,
         pe_1_2_4_n71, pe_1_2_4_n70, pe_1_2_4_n69, pe_1_2_4_n68, pe_1_2_4_n67,
         pe_1_2_4_n66, pe_1_2_4_n65, pe_1_2_4_n64, pe_1_2_4_n63, pe_1_2_4_n62,
         pe_1_2_4_n61, pe_1_2_4_n60, pe_1_2_4_n59, pe_1_2_4_n58, pe_1_2_4_n57,
         pe_1_2_4_n56, pe_1_2_4_n55, pe_1_2_4_n54, pe_1_2_4_n53, pe_1_2_4_n52,
         pe_1_2_4_n51, pe_1_2_4_n50, pe_1_2_4_n49, pe_1_2_4_n48, pe_1_2_4_n47,
         pe_1_2_4_n46, pe_1_2_4_n45, pe_1_2_4_n25, pe_1_2_4_n24, pe_1_2_4_n23,
         pe_1_2_4_n22, pe_1_2_4_n21, pe_1_2_4_n20, pe_1_2_4_n19, pe_1_2_4_n18,
         pe_1_2_4_n17, pe_1_2_4_n16, pe_1_2_4_n15, pe_1_2_4_n14, pe_1_2_4_n13,
         pe_1_2_4_n12, pe_1_2_4_n11, pe_1_2_4_n10, pe_1_2_4_n9, pe_1_2_4_n8,
         pe_1_2_4_n7, pe_1_2_4_n6, pe_1_2_4_n5, pe_1_2_4_n4, pe_1_2_4_n3,
         pe_1_2_4_n2, pe_1_2_4_n1, pe_1_2_4_n44, pe_1_2_4_n43, pe_1_2_4_n42,
         pe_1_2_4_n41, pe_1_2_4_n40, pe_1_2_4_n39, pe_1_2_4_n38, pe_1_2_4_n37,
         pe_1_2_4_n36, pe_1_2_4_n35, pe_1_2_4_n34, pe_1_2_4_n33, pe_1_2_4_n32,
         pe_1_2_4_n31, pe_1_2_4_n30, pe_1_2_4_n29, pe_1_2_4_n28, pe_1_2_4_n27,
         pe_1_2_4_n26, pe_1_2_4_net5992, pe_1_2_4_net5987, pe_1_2_4_net5982,
         pe_1_2_4_net5977, pe_1_2_4_net5972, pe_1_2_4_net5967,
         pe_1_2_4_net5962, pe_1_2_4_net5957, pe_1_2_4_net5952,
         pe_1_2_4_net5947, pe_1_2_4_net5942, pe_1_2_4_net5937,
         pe_1_2_4_net5931, pe_1_2_4_N90, pe_1_2_4_N85, pe_1_2_4_N84,
         pe_1_2_4_N83, pe_1_2_4_N82, pe_1_2_4_N81, pe_1_2_4_N80, pe_1_2_4_N79,
         pe_1_2_4_N77, pe_1_2_4_N76, pe_1_2_4_N75, pe_1_2_4_N74, pe_1_2_4_N73,
         pe_1_2_4_N72, pe_1_2_4_N71, pe_1_2_4_N70, pe_1_2_4_int_data_0_,
         pe_1_2_4_int_data_1_, pe_1_2_4_int_data_2_, pe_1_2_4_int_data_3_,
         pe_1_2_4_N64, pe_1_2_4_N63, pe_1_2_4_N62, pe_1_2_4_N61, pe_1_2_4_N60,
         pe_1_2_4_N59, pe_1_2_5_n90, pe_1_2_5_n89, pe_1_2_5_n88, pe_1_2_5_n87,
         pe_1_2_5_n86, pe_1_2_5_n85, pe_1_2_5_n84, pe_1_2_5_n83, pe_1_2_5_n82,
         pe_1_2_5_n81, pe_1_2_5_n80, pe_1_2_5_n79, pe_1_2_5_n78, pe_1_2_5_n77,
         pe_1_2_5_n76, pe_1_2_5_n75, pe_1_2_5_n74, pe_1_2_5_n73, pe_1_2_5_n72,
         pe_1_2_5_n71, pe_1_2_5_n70, pe_1_2_5_n69, pe_1_2_5_n68, pe_1_2_5_n67,
         pe_1_2_5_n66, pe_1_2_5_n65, pe_1_2_5_n64, pe_1_2_5_n63, pe_1_2_5_n62,
         pe_1_2_5_n61, pe_1_2_5_n60, pe_1_2_5_n59, pe_1_2_5_n58, pe_1_2_5_n57,
         pe_1_2_5_n56, pe_1_2_5_n55, pe_1_2_5_n54, pe_1_2_5_n53, pe_1_2_5_n52,
         pe_1_2_5_n51, pe_1_2_5_n50, pe_1_2_5_n49, pe_1_2_5_n48, pe_1_2_5_n47,
         pe_1_2_5_n46, pe_1_2_5_n45, pe_1_2_5_n25, pe_1_2_5_n24, pe_1_2_5_n23,
         pe_1_2_5_n22, pe_1_2_5_n21, pe_1_2_5_n20, pe_1_2_5_n19, pe_1_2_5_n18,
         pe_1_2_5_n17, pe_1_2_5_n16, pe_1_2_5_n15, pe_1_2_5_n14, pe_1_2_5_n13,
         pe_1_2_5_n12, pe_1_2_5_n11, pe_1_2_5_n10, pe_1_2_5_n9, pe_1_2_5_n8,
         pe_1_2_5_n7, pe_1_2_5_n6, pe_1_2_5_n5, pe_1_2_5_n4, pe_1_2_5_n3,
         pe_1_2_5_n2, pe_1_2_5_n1, pe_1_2_5_n44, pe_1_2_5_n43, pe_1_2_5_n42,
         pe_1_2_5_n41, pe_1_2_5_n40, pe_1_2_5_n39, pe_1_2_5_n38, pe_1_2_5_n37,
         pe_1_2_5_n36, pe_1_2_5_n35, pe_1_2_5_n34, pe_1_2_5_n33, pe_1_2_5_n32,
         pe_1_2_5_n31, pe_1_2_5_n30, pe_1_2_5_n29, pe_1_2_5_n28, pe_1_2_5_n27,
         pe_1_2_5_n26, pe_1_2_5_net5914, pe_1_2_5_net5909, pe_1_2_5_net5904,
         pe_1_2_5_net5899, pe_1_2_5_net5894, pe_1_2_5_net5889,
         pe_1_2_5_net5884, pe_1_2_5_net5879, pe_1_2_5_net5874,
         pe_1_2_5_net5869, pe_1_2_5_net5864, pe_1_2_5_net5859,
         pe_1_2_5_net5853, pe_1_2_5_N90, pe_1_2_5_N85, pe_1_2_5_N84,
         pe_1_2_5_N83, pe_1_2_5_N82, pe_1_2_5_N81, pe_1_2_5_N80, pe_1_2_5_N79,
         pe_1_2_5_N77, pe_1_2_5_N76, pe_1_2_5_N75, pe_1_2_5_N74, pe_1_2_5_N73,
         pe_1_2_5_N72, pe_1_2_5_N71, pe_1_2_5_N70, pe_1_2_5_int_data_0_,
         pe_1_2_5_int_data_1_, pe_1_2_5_int_data_2_, pe_1_2_5_int_data_3_,
         pe_1_2_5_N64, pe_1_2_5_N63, pe_1_2_5_N62, pe_1_2_5_N61, pe_1_2_5_N60,
         pe_1_2_5_N59, pe_1_2_6_n90, pe_1_2_6_n89, pe_1_2_6_n88, pe_1_2_6_n87,
         pe_1_2_6_n86, pe_1_2_6_n85, pe_1_2_6_n84, pe_1_2_6_n83, pe_1_2_6_n82,
         pe_1_2_6_n81, pe_1_2_6_n80, pe_1_2_6_n79, pe_1_2_6_n78, pe_1_2_6_n77,
         pe_1_2_6_n76, pe_1_2_6_n75, pe_1_2_6_n74, pe_1_2_6_n73, pe_1_2_6_n72,
         pe_1_2_6_n71, pe_1_2_6_n70, pe_1_2_6_n69, pe_1_2_6_n68, pe_1_2_6_n67,
         pe_1_2_6_n66, pe_1_2_6_n65, pe_1_2_6_n64, pe_1_2_6_n63, pe_1_2_6_n62,
         pe_1_2_6_n61, pe_1_2_6_n60, pe_1_2_6_n59, pe_1_2_6_n58, pe_1_2_6_n57,
         pe_1_2_6_n56, pe_1_2_6_n55, pe_1_2_6_n54, pe_1_2_6_n53, pe_1_2_6_n52,
         pe_1_2_6_n51, pe_1_2_6_n50, pe_1_2_6_n49, pe_1_2_6_n48, pe_1_2_6_n47,
         pe_1_2_6_n46, pe_1_2_6_n45, pe_1_2_6_n25, pe_1_2_6_n24, pe_1_2_6_n23,
         pe_1_2_6_n22, pe_1_2_6_n21, pe_1_2_6_n20, pe_1_2_6_n19, pe_1_2_6_n18,
         pe_1_2_6_n17, pe_1_2_6_n16, pe_1_2_6_n15, pe_1_2_6_n14, pe_1_2_6_n13,
         pe_1_2_6_n12, pe_1_2_6_n11, pe_1_2_6_n10, pe_1_2_6_n9, pe_1_2_6_n8,
         pe_1_2_6_n7, pe_1_2_6_n6, pe_1_2_6_n5, pe_1_2_6_n4, pe_1_2_6_n3,
         pe_1_2_6_n2, pe_1_2_6_n1, pe_1_2_6_n44, pe_1_2_6_n43, pe_1_2_6_n42,
         pe_1_2_6_n41, pe_1_2_6_n40, pe_1_2_6_n39, pe_1_2_6_n38, pe_1_2_6_n37,
         pe_1_2_6_n36, pe_1_2_6_n35, pe_1_2_6_n34, pe_1_2_6_n33, pe_1_2_6_n32,
         pe_1_2_6_n31, pe_1_2_6_n30, pe_1_2_6_n29, pe_1_2_6_n28, pe_1_2_6_n27,
         pe_1_2_6_n26, pe_1_2_6_net5836, pe_1_2_6_net5831, pe_1_2_6_net5826,
         pe_1_2_6_net5821, pe_1_2_6_net5816, pe_1_2_6_net5811,
         pe_1_2_6_net5806, pe_1_2_6_net5801, pe_1_2_6_net5796,
         pe_1_2_6_net5791, pe_1_2_6_net5786, pe_1_2_6_net5781,
         pe_1_2_6_net5775, pe_1_2_6_N90, pe_1_2_6_N85, pe_1_2_6_N84,
         pe_1_2_6_N83, pe_1_2_6_N82, pe_1_2_6_N81, pe_1_2_6_N80, pe_1_2_6_N79,
         pe_1_2_6_N77, pe_1_2_6_N76, pe_1_2_6_N75, pe_1_2_6_N74, pe_1_2_6_N73,
         pe_1_2_6_N72, pe_1_2_6_N71, pe_1_2_6_N70, pe_1_2_6_int_data_0_,
         pe_1_2_6_int_data_1_, pe_1_2_6_int_data_2_, pe_1_2_6_int_data_3_,
         pe_1_2_6_N64, pe_1_2_6_N63, pe_1_2_6_N62, pe_1_2_6_N61, pe_1_2_6_N60,
         pe_1_2_6_N59, pe_1_2_7_n90, pe_1_2_7_n89, pe_1_2_7_n88, pe_1_2_7_n87,
         pe_1_2_7_n86, pe_1_2_7_n85, pe_1_2_7_n84, pe_1_2_7_n83, pe_1_2_7_n82,
         pe_1_2_7_n81, pe_1_2_7_n80, pe_1_2_7_n79, pe_1_2_7_n78, pe_1_2_7_n77,
         pe_1_2_7_n76, pe_1_2_7_n75, pe_1_2_7_n74, pe_1_2_7_n73, pe_1_2_7_n72,
         pe_1_2_7_n71, pe_1_2_7_n70, pe_1_2_7_n69, pe_1_2_7_n68, pe_1_2_7_n67,
         pe_1_2_7_n66, pe_1_2_7_n65, pe_1_2_7_n64, pe_1_2_7_n63, pe_1_2_7_n62,
         pe_1_2_7_n61, pe_1_2_7_n60, pe_1_2_7_n59, pe_1_2_7_n58, pe_1_2_7_n57,
         pe_1_2_7_n56, pe_1_2_7_n55, pe_1_2_7_n54, pe_1_2_7_n53, pe_1_2_7_n52,
         pe_1_2_7_n51, pe_1_2_7_n50, pe_1_2_7_n49, pe_1_2_7_n48, pe_1_2_7_n47,
         pe_1_2_7_n46, pe_1_2_7_n45, pe_1_2_7_n25, pe_1_2_7_n24, pe_1_2_7_n23,
         pe_1_2_7_n22, pe_1_2_7_n21, pe_1_2_7_n20, pe_1_2_7_n19, pe_1_2_7_n18,
         pe_1_2_7_n17, pe_1_2_7_n16, pe_1_2_7_n15, pe_1_2_7_n14, pe_1_2_7_n13,
         pe_1_2_7_n12, pe_1_2_7_n11, pe_1_2_7_n10, pe_1_2_7_n9, pe_1_2_7_n8,
         pe_1_2_7_n7, pe_1_2_7_n6, pe_1_2_7_n5, pe_1_2_7_n4, pe_1_2_7_n3,
         pe_1_2_7_n2, pe_1_2_7_n1, pe_1_2_7_n44, pe_1_2_7_n43, pe_1_2_7_n42,
         pe_1_2_7_n41, pe_1_2_7_n40, pe_1_2_7_n39, pe_1_2_7_n38, pe_1_2_7_n37,
         pe_1_2_7_n36, pe_1_2_7_n35, pe_1_2_7_n34, pe_1_2_7_n33, pe_1_2_7_n32,
         pe_1_2_7_n31, pe_1_2_7_n30, pe_1_2_7_n29, pe_1_2_7_n28, pe_1_2_7_n27,
         pe_1_2_7_n26, pe_1_2_7_net5758, pe_1_2_7_net5753, pe_1_2_7_net5748,
         pe_1_2_7_net5743, pe_1_2_7_net5738, pe_1_2_7_net5733,
         pe_1_2_7_net5728, pe_1_2_7_net5723, pe_1_2_7_net5718,
         pe_1_2_7_net5713, pe_1_2_7_net5708, pe_1_2_7_net5703,
         pe_1_2_7_net5697, pe_1_2_7_N90, pe_1_2_7_N85, pe_1_2_7_N84,
         pe_1_2_7_N83, pe_1_2_7_N82, pe_1_2_7_N81, pe_1_2_7_N80, pe_1_2_7_N79,
         pe_1_2_7_N77, pe_1_2_7_N76, pe_1_2_7_N75, pe_1_2_7_N74, pe_1_2_7_N73,
         pe_1_2_7_N72, pe_1_2_7_N71, pe_1_2_7_N70, pe_1_2_7_int_data_0_,
         pe_1_2_7_int_data_1_, pe_1_2_7_int_data_2_, pe_1_2_7_int_data_3_,
         pe_1_2_7_N64, pe_1_2_7_N63, pe_1_2_7_N62, pe_1_2_7_N61, pe_1_2_7_N60,
         pe_1_2_7_N59, pe_1_3_0_n87, pe_1_3_0_n86, pe_1_3_0_n85, pe_1_3_0_n84,
         pe_1_3_0_n83, pe_1_3_0_n82, pe_1_3_0_n81, pe_1_3_0_n80, pe_1_3_0_n79,
         pe_1_3_0_n78, pe_1_3_0_n77, pe_1_3_0_n76, pe_1_3_0_n75, pe_1_3_0_n74,
         pe_1_3_0_n73, pe_1_3_0_n72, pe_1_3_0_n71, pe_1_3_0_n70, pe_1_3_0_n69,
         pe_1_3_0_n68, pe_1_3_0_n67, pe_1_3_0_n66, pe_1_3_0_n65, pe_1_3_0_n64,
         pe_1_3_0_n63, pe_1_3_0_n62, pe_1_3_0_n61, pe_1_3_0_n60, pe_1_3_0_n59,
         pe_1_3_0_n58, pe_1_3_0_n57, pe_1_3_0_n56, pe_1_3_0_n55, pe_1_3_0_n54,
         pe_1_3_0_n53, pe_1_3_0_n52, pe_1_3_0_n51, pe_1_3_0_n50, pe_1_3_0_n49,
         pe_1_3_0_n48, pe_1_3_0_n47, pe_1_3_0_n46, pe_1_3_0_n45, pe_1_3_0_n25,
         pe_1_3_0_n24, pe_1_3_0_n23, pe_1_3_0_n22, pe_1_3_0_n21, pe_1_3_0_n20,
         pe_1_3_0_n19, pe_1_3_0_n18, pe_1_3_0_n17, pe_1_3_0_n16, pe_1_3_0_n15,
         pe_1_3_0_n14, pe_1_3_0_n13, pe_1_3_0_n12, pe_1_3_0_n11, pe_1_3_0_n10,
         pe_1_3_0_n9, pe_1_3_0_n8, pe_1_3_0_n7, pe_1_3_0_n6, pe_1_3_0_n5,
         pe_1_3_0_n4, pe_1_3_0_n3, pe_1_3_0_n2, pe_1_3_0_n1, pe_1_3_0_n44,
         pe_1_3_0_n43, pe_1_3_0_n42, pe_1_3_0_n41, pe_1_3_0_n40, pe_1_3_0_n39,
         pe_1_3_0_n38, pe_1_3_0_n37, pe_1_3_0_n36, pe_1_3_0_n35, pe_1_3_0_n34,
         pe_1_3_0_n33, pe_1_3_0_n32, pe_1_3_0_n31, pe_1_3_0_n30, pe_1_3_0_n29,
         pe_1_3_0_n28, pe_1_3_0_n27, pe_1_3_0_n26, pe_1_3_0_net5680,
         pe_1_3_0_net5675, pe_1_3_0_net5670, pe_1_3_0_net5665,
         pe_1_3_0_net5660, pe_1_3_0_net5655, pe_1_3_0_net5650,
         pe_1_3_0_net5645, pe_1_3_0_net5640, pe_1_3_0_net5635,
         pe_1_3_0_net5630, pe_1_3_0_net5625, pe_1_3_0_net5619, pe_1_3_0_N90,
         pe_1_3_0_N85, pe_1_3_0_N84, pe_1_3_0_N83, pe_1_3_0_N82, pe_1_3_0_N81,
         pe_1_3_0_N80, pe_1_3_0_N79, pe_1_3_0_N77, pe_1_3_0_N76, pe_1_3_0_N75,
         pe_1_3_0_N74, pe_1_3_0_N73, pe_1_3_0_N72, pe_1_3_0_N71, pe_1_3_0_N70,
         pe_1_3_0_int_data_0_, pe_1_3_0_int_data_1_, pe_1_3_0_int_data_2_,
         pe_1_3_0_int_data_3_, pe_1_3_0_N64, pe_1_3_0_N63, pe_1_3_0_N62,
         pe_1_3_0_N61, pe_1_3_0_N60, pe_1_3_0_N59, pe_1_3_0_o_data_h_0_,
         pe_1_3_0_o_data_h_1_, pe_1_3_0_o_data_h_2_, pe_1_3_0_o_data_h_3_,
         pe_1_3_1_n86, pe_1_3_1_n85, pe_1_3_1_n84, pe_1_3_1_n83, pe_1_3_1_n82,
         pe_1_3_1_n81, pe_1_3_1_n80, pe_1_3_1_n79, pe_1_3_1_n78, pe_1_3_1_n77,
         pe_1_3_1_n76, pe_1_3_1_n75, pe_1_3_1_n74, pe_1_3_1_n73, pe_1_3_1_n72,
         pe_1_3_1_n71, pe_1_3_1_n70, pe_1_3_1_n69, pe_1_3_1_n68, pe_1_3_1_n67,
         pe_1_3_1_n66, pe_1_3_1_n65, pe_1_3_1_n64, pe_1_3_1_n63, pe_1_3_1_n62,
         pe_1_3_1_n61, pe_1_3_1_n60, pe_1_3_1_n59, pe_1_3_1_n58, pe_1_3_1_n57,
         pe_1_3_1_n56, pe_1_3_1_n55, pe_1_3_1_n54, pe_1_3_1_n53, pe_1_3_1_n52,
         pe_1_3_1_n51, pe_1_3_1_n50, pe_1_3_1_n49, pe_1_3_1_n48, pe_1_3_1_n47,
         pe_1_3_1_n46, pe_1_3_1_n45, pe_1_3_1_n25, pe_1_3_1_n24, pe_1_3_1_n23,
         pe_1_3_1_n22, pe_1_3_1_n21, pe_1_3_1_n20, pe_1_3_1_n19, pe_1_3_1_n18,
         pe_1_3_1_n17, pe_1_3_1_n16, pe_1_3_1_n15, pe_1_3_1_n14, pe_1_3_1_n13,
         pe_1_3_1_n12, pe_1_3_1_n11, pe_1_3_1_n10, pe_1_3_1_n9, pe_1_3_1_n8,
         pe_1_3_1_n7, pe_1_3_1_n6, pe_1_3_1_n5, pe_1_3_1_n4, pe_1_3_1_n3,
         pe_1_3_1_n2, pe_1_3_1_n1, pe_1_3_1_n44, pe_1_3_1_n43, pe_1_3_1_n42,
         pe_1_3_1_n41, pe_1_3_1_n40, pe_1_3_1_n39, pe_1_3_1_n38, pe_1_3_1_n37,
         pe_1_3_1_n36, pe_1_3_1_n35, pe_1_3_1_n34, pe_1_3_1_n33, pe_1_3_1_n32,
         pe_1_3_1_n31, pe_1_3_1_n30, pe_1_3_1_n29, pe_1_3_1_n28, pe_1_3_1_n27,
         pe_1_3_1_n26, pe_1_3_1_net5602, pe_1_3_1_net5597, pe_1_3_1_net5592,
         pe_1_3_1_net5587, pe_1_3_1_net5582, pe_1_3_1_net5577,
         pe_1_3_1_net5572, pe_1_3_1_net5567, pe_1_3_1_net5562,
         pe_1_3_1_net5557, pe_1_3_1_net5552, pe_1_3_1_net5547,
         pe_1_3_1_net5541, pe_1_3_1_N90, pe_1_3_1_N85, pe_1_3_1_N84,
         pe_1_3_1_N83, pe_1_3_1_N82, pe_1_3_1_N81, pe_1_3_1_N80, pe_1_3_1_N79,
         pe_1_3_1_N77, pe_1_3_1_N76, pe_1_3_1_N75, pe_1_3_1_N74, pe_1_3_1_N73,
         pe_1_3_1_N72, pe_1_3_1_N71, pe_1_3_1_N70, pe_1_3_1_int_data_0_,
         pe_1_3_1_int_data_1_, pe_1_3_1_int_data_2_, pe_1_3_1_int_data_3_,
         pe_1_3_1_N64, pe_1_3_1_N63, pe_1_3_1_N62, pe_1_3_1_N61, pe_1_3_1_N60,
         pe_1_3_1_N59, pe_1_3_2_n87, pe_1_3_2_n86, pe_1_3_2_n85, pe_1_3_2_n84,
         pe_1_3_2_n83, pe_1_3_2_n82, pe_1_3_2_n81, pe_1_3_2_n80, pe_1_3_2_n79,
         pe_1_3_2_n78, pe_1_3_2_n77, pe_1_3_2_n76, pe_1_3_2_n75, pe_1_3_2_n74,
         pe_1_3_2_n73, pe_1_3_2_n72, pe_1_3_2_n71, pe_1_3_2_n70, pe_1_3_2_n69,
         pe_1_3_2_n68, pe_1_3_2_n67, pe_1_3_2_n66, pe_1_3_2_n65, pe_1_3_2_n64,
         pe_1_3_2_n63, pe_1_3_2_n62, pe_1_3_2_n61, pe_1_3_2_n60, pe_1_3_2_n59,
         pe_1_3_2_n58, pe_1_3_2_n57, pe_1_3_2_n56, pe_1_3_2_n55, pe_1_3_2_n54,
         pe_1_3_2_n53, pe_1_3_2_n52, pe_1_3_2_n51, pe_1_3_2_n50, pe_1_3_2_n49,
         pe_1_3_2_n48, pe_1_3_2_n47, pe_1_3_2_n46, pe_1_3_2_n45, pe_1_3_2_n25,
         pe_1_3_2_n24, pe_1_3_2_n23, pe_1_3_2_n22, pe_1_3_2_n21, pe_1_3_2_n20,
         pe_1_3_2_n19, pe_1_3_2_n18, pe_1_3_2_n17, pe_1_3_2_n16, pe_1_3_2_n15,
         pe_1_3_2_n14, pe_1_3_2_n13, pe_1_3_2_n12, pe_1_3_2_n11, pe_1_3_2_n10,
         pe_1_3_2_n9, pe_1_3_2_n8, pe_1_3_2_n7, pe_1_3_2_n6, pe_1_3_2_n5,
         pe_1_3_2_n4, pe_1_3_2_n3, pe_1_3_2_n2, pe_1_3_2_n1, pe_1_3_2_n44,
         pe_1_3_2_n43, pe_1_3_2_n42, pe_1_3_2_n41, pe_1_3_2_n40, pe_1_3_2_n39,
         pe_1_3_2_n38, pe_1_3_2_n37, pe_1_3_2_n36, pe_1_3_2_n35, pe_1_3_2_n34,
         pe_1_3_2_n33, pe_1_3_2_n32, pe_1_3_2_n31, pe_1_3_2_n30, pe_1_3_2_n29,
         pe_1_3_2_n28, pe_1_3_2_n27, pe_1_3_2_n26, pe_1_3_2_net5524,
         pe_1_3_2_net5519, pe_1_3_2_net5514, pe_1_3_2_net5509,
         pe_1_3_2_net5504, pe_1_3_2_net5499, pe_1_3_2_net5494,
         pe_1_3_2_net5489, pe_1_3_2_net5484, pe_1_3_2_net5479,
         pe_1_3_2_net5474, pe_1_3_2_net5469, pe_1_3_2_net5463, pe_1_3_2_N90,
         pe_1_3_2_N85, pe_1_3_2_N84, pe_1_3_2_N83, pe_1_3_2_N82, pe_1_3_2_N81,
         pe_1_3_2_N80, pe_1_3_2_N79, pe_1_3_2_N77, pe_1_3_2_N76, pe_1_3_2_N75,
         pe_1_3_2_N74, pe_1_3_2_N73, pe_1_3_2_N72, pe_1_3_2_N71, pe_1_3_2_N70,
         pe_1_3_2_int_data_0_, pe_1_3_2_int_data_1_, pe_1_3_2_int_data_2_,
         pe_1_3_2_int_data_3_, pe_1_3_2_N64, pe_1_3_2_N63, pe_1_3_2_N62,
         pe_1_3_2_N61, pe_1_3_2_N60, pe_1_3_2_N59, pe_1_3_3_n88, pe_1_3_3_n87,
         pe_1_3_3_n86, pe_1_3_3_n85, pe_1_3_3_n84, pe_1_3_3_n83, pe_1_3_3_n82,
         pe_1_3_3_n81, pe_1_3_3_n80, pe_1_3_3_n79, pe_1_3_3_n78, pe_1_3_3_n77,
         pe_1_3_3_n76, pe_1_3_3_n75, pe_1_3_3_n74, pe_1_3_3_n73, pe_1_3_3_n72,
         pe_1_3_3_n71, pe_1_3_3_n70, pe_1_3_3_n69, pe_1_3_3_n68, pe_1_3_3_n67,
         pe_1_3_3_n66, pe_1_3_3_n65, pe_1_3_3_n64, pe_1_3_3_n63, pe_1_3_3_n62,
         pe_1_3_3_n61, pe_1_3_3_n60, pe_1_3_3_n59, pe_1_3_3_n58, pe_1_3_3_n57,
         pe_1_3_3_n56, pe_1_3_3_n55, pe_1_3_3_n54, pe_1_3_3_n53, pe_1_3_3_n52,
         pe_1_3_3_n51, pe_1_3_3_n50, pe_1_3_3_n49, pe_1_3_3_n48, pe_1_3_3_n47,
         pe_1_3_3_n46, pe_1_3_3_n45, pe_1_3_3_n25, pe_1_3_3_n24, pe_1_3_3_n23,
         pe_1_3_3_n22, pe_1_3_3_n21, pe_1_3_3_n20, pe_1_3_3_n19, pe_1_3_3_n18,
         pe_1_3_3_n17, pe_1_3_3_n16, pe_1_3_3_n15, pe_1_3_3_n14, pe_1_3_3_n13,
         pe_1_3_3_n12, pe_1_3_3_n11, pe_1_3_3_n10, pe_1_3_3_n9, pe_1_3_3_n8,
         pe_1_3_3_n7, pe_1_3_3_n6, pe_1_3_3_n5, pe_1_3_3_n4, pe_1_3_3_n3,
         pe_1_3_3_n2, pe_1_3_3_n1, pe_1_3_3_n44, pe_1_3_3_n43, pe_1_3_3_n42,
         pe_1_3_3_n41, pe_1_3_3_n40, pe_1_3_3_n39, pe_1_3_3_n38, pe_1_3_3_n37,
         pe_1_3_3_n36, pe_1_3_3_n35, pe_1_3_3_n34, pe_1_3_3_n33, pe_1_3_3_n32,
         pe_1_3_3_n31, pe_1_3_3_n30, pe_1_3_3_n29, pe_1_3_3_n28, pe_1_3_3_n27,
         pe_1_3_3_n26, pe_1_3_3_net5446, pe_1_3_3_net5441, pe_1_3_3_net5436,
         pe_1_3_3_net5431, pe_1_3_3_net5426, pe_1_3_3_net5421,
         pe_1_3_3_net5416, pe_1_3_3_net5411, pe_1_3_3_net5406,
         pe_1_3_3_net5401, pe_1_3_3_net5396, pe_1_3_3_net5391,
         pe_1_3_3_net5385, pe_1_3_3_N90, pe_1_3_3_N85, pe_1_3_3_N84,
         pe_1_3_3_N83, pe_1_3_3_N82, pe_1_3_3_N81, pe_1_3_3_N80, pe_1_3_3_N79,
         pe_1_3_3_N77, pe_1_3_3_N76, pe_1_3_3_N75, pe_1_3_3_N74, pe_1_3_3_N73,
         pe_1_3_3_N72, pe_1_3_3_N71, pe_1_3_3_N70, pe_1_3_3_int_data_0_,
         pe_1_3_3_int_data_1_, pe_1_3_3_int_data_2_, pe_1_3_3_int_data_3_,
         pe_1_3_3_N64, pe_1_3_3_N63, pe_1_3_3_N62, pe_1_3_3_N61, pe_1_3_3_N60,
         pe_1_3_3_N59, pe_1_3_4_n90, pe_1_3_4_n89, pe_1_3_4_n88, pe_1_3_4_n87,
         pe_1_3_4_n86, pe_1_3_4_n85, pe_1_3_4_n84, pe_1_3_4_n83, pe_1_3_4_n82,
         pe_1_3_4_n81, pe_1_3_4_n80, pe_1_3_4_n79, pe_1_3_4_n78, pe_1_3_4_n77,
         pe_1_3_4_n76, pe_1_3_4_n75, pe_1_3_4_n74, pe_1_3_4_n73, pe_1_3_4_n72,
         pe_1_3_4_n71, pe_1_3_4_n70, pe_1_3_4_n69, pe_1_3_4_n68, pe_1_3_4_n67,
         pe_1_3_4_n66, pe_1_3_4_n65, pe_1_3_4_n64, pe_1_3_4_n63, pe_1_3_4_n62,
         pe_1_3_4_n61, pe_1_3_4_n60, pe_1_3_4_n59, pe_1_3_4_n58, pe_1_3_4_n57,
         pe_1_3_4_n56, pe_1_3_4_n55, pe_1_3_4_n54, pe_1_3_4_n53, pe_1_3_4_n52,
         pe_1_3_4_n51, pe_1_3_4_n50, pe_1_3_4_n49, pe_1_3_4_n48, pe_1_3_4_n47,
         pe_1_3_4_n46, pe_1_3_4_n45, pe_1_3_4_n25, pe_1_3_4_n24, pe_1_3_4_n23,
         pe_1_3_4_n22, pe_1_3_4_n21, pe_1_3_4_n20, pe_1_3_4_n19, pe_1_3_4_n18,
         pe_1_3_4_n17, pe_1_3_4_n16, pe_1_3_4_n15, pe_1_3_4_n14, pe_1_3_4_n13,
         pe_1_3_4_n12, pe_1_3_4_n11, pe_1_3_4_n10, pe_1_3_4_n9, pe_1_3_4_n8,
         pe_1_3_4_n7, pe_1_3_4_n6, pe_1_3_4_n5, pe_1_3_4_n4, pe_1_3_4_n3,
         pe_1_3_4_n2, pe_1_3_4_n1, pe_1_3_4_n44, pe_1_3_4_n43, pe_1_3_4_n42,
         pe_1_3_4_n41, pe_1_3_4_n40, pe_1_3_4_n39, pe_1_3_4_n38, pe_1_3_4_n37,
         pe_1_3_4_n36, pe_1_3_4_n35, pe_1_3_4_n34, pe_1_3_4_n33, pe_1_3_4_n32,
         pe_1_3_4_n31, pe_1_3_4_n30, pe_1_3_4_n29, pe_1_3_4_n28, pe_1_3_4_n27,
         pe_1_3_4_n26, pe_1_3_4_net5368, pe_1_3_4_net5363, pe_1_3_4_net5358,
         pe_1_3_4_net5353, pe_1_3_4_net5348, pe_1_3_4_net5343,
         pe_1_3_4_net5338, pe_1_3_4_net5333, pe_1_3_4_net5328,
         pe_1_3_4_net5323, pe_1_3_4_net5318, pe_1_3_4_net5313,
         pe_1_3_4_net5307, pe_1_3_4_N90, pe_1_3_4_N85, pe_1_3_4_N84,
         pe_1_3_4_N83, pe_1_3_4_N82, pe_1_3_4_N81, pe_1_3_4_N80, pe_1_3_4_N79,
         pe_1_3_4_N77, pe_1_3_4_N76, pe_1_3_4_N75, pe_1_3_4_N74, pe_1_3_4_N73,
         pe_1_3_4_N72, pe_1_3_4_N71, pe_1_3_4_N70, pe_1_3_4_int_data_0_,
         pe_1_3_4_int_data_1_, pe_1_3_4_int_data_2_, pe_1_3_4_int_data_3_,
         pe_1_3_4_N64, pe_1_3_4_N63, pe_1_3_4_N62, pe_1_3_4_N61, pe_1_3_4_N60,
         pe_1_3_4_N59, pe_1_3_5_n90, pe_1_3_5_n89, pe_1_3_5_n88, pe_1_3_5_n87,
         pe_1_3_5_n86, pe_1_3_5_n85, pe_1_3_5_n84, pe_1_3_5_n83, pe_1_3_5_n82,
         pe_1_3_5_n81, pe_1_3_5_n80, pe_1_3_5_n79, pe_1_3_5_n78, pe_1_3_5_n77,
         pe_1_3_5_n76, pe_1_3_5_n75, pe_1_3_5_n74, pe_1_3_5_n73, pe_1_3_5_n72,
         pe_1_3_5_n71, pe_1_3_5_n70, pe_1_3_5_n69, pe_1_3_5_n68, pe_1_3_5_n67,
         pe_1_3_5_n66, pe_1_3_5_n65, pe_1_3_5_n64, pe_1_3_5_n63, pe_1_3_5_n62,
         pe_1_3_5_n61, pe_1_3_5_n60, pe_1_3_5_n59, pe_1_3_5_n58, pe_1_3_5_n57,
         pe_1_3_5_n56, pe_1_3_5_n55, pe_1_3_5_n54, pe_1_3_5_n53, pe_1_3_5_n52,
         pe_1_3_5_n51, pe_1_3_5_n50, pe_1_3_5_n49, pe_1_3_5_n48, pe_1_3_5_n47,
         pe_1_3_5_n46, pe_1_3_5_n45, pe_1_3_5_n25, pe_1_3_5_n24, pe_1_3_5_n23,
         pe_1_3_5_n22, pe_1_3_5_n21, pe_1_3_5_n20, pe_1_3_5_n19, pe_1_3_5_n18,
         pe_1_3_5_n17, pe_1_3_5_n16, pe_1_3_5_n15, pe_1_3_5_n14, pe_1_3_5_n13,
         pe_1_3_5_n12, pe_1_3_5_n11, pe_1_3_5_n10, pe_1_3_5_n9, pe_1_3_5_n8,
         pe_1_3_5_n7, pe_1_3_5_n6, pe_1_3_5_n5, pe_1_3_5_n4, pe_1_3_5_n3,
         pe_1_3_5_n2, pe_1_3_5_n1, pe_1_3_5_n44, pe_1_3_5_n43, pe_1_3_5_n42,
         pe_1_3_5_n41, pe_1_3_5_n40, pe_1_3_5_n39, pe_1_3_5_n38, pe_1_3_5_n37,
         pe_1_3_5_n36, pe_1_3_5_n35, pe_1_3_5_n34, pe_1_3_5_n33, pe_1_3_5_n32,
         pe_1_3_5_n31, pe_1_3_5_n30, pe_1_3_5_n29, pe_1_3_5_n28, pe_1_3_5_n27,
         pe_1_3_5_n26, pe_1_3_5_net5290, pe_1_3_5_net5285, pe_1_3_5_net5280,
         pe_1_3_5_net5275, pe_1_3_5_net5270, pe_1_3_5_net5265,
         pe_1_3_5_net5260, pe_1_3_5_net5255, pe_1_3_5_net5250,
         pe_1_3_5_net5245, pe_1_3_5_net5240, pe_1_3_5_net5235,
         pe_1_3_5_net5229, pe_1_3_5_N90, pe_1_3_5_N85, pe_1_3_5_N84,
         pe_1_3_5_N83, pe_1_3_5_N82, pe_1_3_5_N81, pe_1_3_5_N80, pe_1_3_5_N79,
         pe_1_3_5_N77, pe_1_3_5_N76, pe_1_3_5_N75, pe_1_3_5_N74, pe_1_3_5_N73,
         pe_1_3_5_N72, pe_1_3_5_N71, pe_1_3_5_N70, pe_1_3_5_int_data_0_,
         pe_1_3_5_int_data_1_, pe_1_3_5_int_data_2_, pe_1_3_5_int_data_3_,
         pe_1_3_5_N64, pe_1_3_5_N63, pe_1_3_5_N62, pe_1_3_5_N61, pe_1_3_5_N60,
         pe_1_3_5_N59, pe_1_3_6_n90, pe_1_3_6_n89, pe_1_3_6_n88, pe_1_3_6_n87,
         pe_1_3_6_n86, pe_1_3_6_n85, pe_1_3_6_n84, pe_1_3_6_n83, pe_1_3_6_n82,
         pe_1_3_6_n81, pe_1_3_6_n80, pe_1_3_6_n79, pe_1_3_6_n78, pe_1_3_6_n77,
         pe_1_3_6_n76, pe_1_3_6_n75, pe_1_3_6_n74, pe_1_3_6_n73, pe_1_3_6_n72,
         pe_1_3_6_n71, pe_1_3_6_n70, pe_1_3_6_n69, pe_1_3_6_n68, pe_1_3_6_n67,
         pe_1_3_6_n66, pe_1_3_6_n65, pe_1_3_6_n64, pe_1_3_6_n63, pe_1_3_6_n62,
         pe_1_3_6_n61, pe_1_3_6_n60, pe_1_3_6_n59, pe_1_3_6_n58, pe_1_3_6_n57,
         pe_1_3_6_n56, pe_1_3_6_n55, pe_1_3_6_n54, pe_1_3_6_n53, pe_1_3_6_n52,
         pe_1_3_6_n51, pe_1_3_6_n50, pe_1_3_6_n49, pe_1_3_6_n48, pe_1_3_6_n47,
         pe_1_3_6_n46, pe_1_3_6_n45, pe_1_3_6_n25, pe_1_3_6_n24, pe_1_3_6_n23,
         pe_1_3_6_n22, pe_1_3_6_n21, pe_1_3_6_n20, pe_1_3_6_n19, pe_1_3_6_n18,
         pe_1_3_6_n17, pe_1_3_6_n16, pe_1_3_6_n15, pe_1_3_6_n14, pe_1_3_6_n13,
         pe_1_3_6_n12, pe_1_3_6_n11, pe_1_3_6_n10, pe_1_3_6_n9, pe_1_3_6_n8,
         pe_1_3_6_n7, pe_1_3_6_n6, pe_1_3_6_n5, pe_1_3_6_n4, pe_1_3_6_n3,
         pe_1_3_6_n2, pe_1_3_6_n1, pe_1_3_6_n44, pe_1_3_6_n43, pe_1_3_6_n42,
         pe_1_3_6_n41, pe_1_3_6_n40, pe_1_3_6_n39, pe_1_3_6_n38, pe_1_3_6_n37,
         pe_1_3_6_n36, pe_1_3_6_n35, pe_1_3_6_n34, pe_1_3_6_n33, pe_1_3_6_n32,
         pe_1_3_6_n31, pe_1_3_6_n30, pe_1_3_6_n29, pe_1_3_6_n28, pe_1_3_6_n27,
         pe_1_3_6_n26, pe_1_3_6_net5212, pe_1_3_6_net5207, pe_1_3_6_net5202,
         pe_1_3_6_net5197, pe_1_3_6_net5192, pe_1_3_6_net5187,
         pe_1_3_6_net5182, pe_1_3_6_net5177, pe_1_3_6_net5172,
         pe_1_3_6_net5167, pe_1_3_6_net5162, pe_1_3_6_net5157,
         pe_1_3_6_net5151, pe_1_3_6_N90, pe_1_3_6_N85, pe_1_3_6_N84,
         pe_1_3_6_N83, pe_1_3_6_N82, pe_1_3_6_N81, pe_1_3_6_N80, pe_1_3_6_N79,
         pe_1_3_6_N77, pe_1_3_6_N76, pe_1_3_6_N75, pe_1_3_6_N74, pe_1_3_6_N73,
         pe_1_3_6_N72, pe_1_3_6_N71, pe_1_3_6_N70, pe_1_3_6_int_data_0_,
         pe_1_3_6_int_data_1_, pe_1_3_6_int_data_2_, pe_1_3_6_int_data_3_,
         pe_1_3_6_N64, pe_1_3_6_N63, pe_1_3_6_N62, pe_1_3_6_N61, pe_1_3_6_N60,
         pe_1_3_6_N59, pe_1_3_7_n90, pe_1_3_7_n89, pe_1_3_7_n88, pe_1_3_7_n87,
         pe_1_3_7_n86, pe_1_3_7_n85, pe_1_3_7_n84, pe_1_3_7_n83, pe_1_3_7_n82,
         pe_1_3_7_n81, pe_1_3_7_n80, pe_1_3_7_n79, pe_1_3_7_n78, pe_1_3_7_n77,
         pe_1_3_7_n76, pe_1_3_7_n75, pe_1_3_7_n74, pe_1_3_7_n73, pe_1_3_7_n72,
         pe_1_3_7_n71, pe_1_3_7_n70, pe_1_3_7_n69, pe_1_3_7_n68, pe_1_3_7_n67,
         pe_1_3_7_n66, pe_1_3_7_n65, pe_1_3_7_n64, pe_1_3_7_n63, pe_1_3_7_n62,
         pe_1_3_7_n61, pe_1_3_7_n60, pe_1_3_7_n59, pe_1_3_7_n58, pe_1_3_7_n57,
         pe_1_3_7_n56, pe_1_3_7_n55, pe_1_3_7_n54, pe_1_3_7_n53, pe_1_3_7_n52,
         pe_1_3_7_n51, pe_1_3_7_n50, pe_1_3_7_n49, pe_1_3_7_n48, pe_1_3_7_n47,
         pe_1_3_7_n46, pe_1_3_7_n45, pe_1_3_7_n25, pe_1_3_7_n24, pe_1_3_7_n23,
         pe_1_3_7_n22, pe_1_3_7_n21, pe_1_3_7_n20, pe_1_3_7_n19, pe_1_3_7_n18,
         pe_1_3_7_n17, pe_1_3_7_n16, pe_1_3_7_n15, pe_1_3_7_n14, pe_1_3_7_n13,
         pe_1_3_7_n12, pe_1_3_7_n11, pe_1_3_7_n10, pe_1_3_7_n9, pe_1_3_7_n8,
         pe_1_3_7_n7, pe_1_3_7_n6, pe_1_3_7_n5, pe_1_3_7_n4, pe_1_3_7_n3,
         pe_1_3_7_n2, pe_1_3_7_n1, pe_1_3_7_n44, pe_1_3_7_n43, pe_1_3_7_n42,
         pe_1_3_7_n41, pe_1_3_7_n40, pe_1_3_7_n39, pe_1_3_7_n38, pe_1_3_7_n37,
         pe_1_3_7_n36, pe_1_3_7_n35, pe_1_3_7_n34, pe_1_3_7_n33, pe_1_3_7_n32,
         pe_1_3_7_n31, pe_1_3_7_n30, pe_1_3_7_n29, pe_1_3_7_n28, pe_1_3_7_n27,
         pe_1_3_7_n26, pe_1_3_7_net5134, pe_1_3_7_net5129, pe_1_3_7_net5124,
         pe_1_3_7_net5119, pe_1_3_7_net5114, pe_1_3_7_net5109,
         pe_1_3_7_net5104, pe_1_3_7_net5099, pe_1_3_7_net5094,
         pe_1_3_7_net5089, pe_1_3_7_net5084, pe_1_3_7_net5079,
         pe_1_3_7_net5073, pe_1_3_7_N90, pe_1_3_7_N85, pe_1_3_7_N84,
         pe_1_3_7_N83, pe_1_3_7_N82, pe_1_3_7_N81, pe_1_3_7_N80, pe_1_3_7_N79,
         pe_1_3_7_N77, pe_1_3_7_N76, pe_1_3_7_N75, pe_1_3_7_N74, pe_1_3_7_N73,
         pe_1_3_7_N72, pe_1_3_7_N71, pe_1_3_7_N70, pe_1_3_7_int_data_0_,
         pe_1_3_7_int_data_1_, pe_1_3_7_int_data_2_, pe_1_3_7_int_data_3_,
         pe_1_3_7_N64, pe_1_3_7_N63, pe_1_3_7_N62, pe_1_3_7_N61, pe_1_3_7_N60,
         pe_1_3_7_N59, pe_1_4_0_n90, pe_1_4_0_n89, pe_1_4_0_n88, pe_1_4_0_n87,
         pe_1_4_0_n86, pe_1_4_0_n85, pe_1_4_0_n84, pe_1_4_0_n83, pe_1_4_0_n82,
         pe_1_4_0_n81, pe_1_4_0_n80, pe_1_4_0_n79, pe_1_4_0_n78, pe_1_4_0_n77,
         pe_1_4_0_n76, pe_1_4_0_n75, pe_1_4_0_n74, pe_1_4_0_n73, pe_1_4_0_n72,
         pe_1_4_0_n71, pe_1_4_0_n70, pe_1_4_0_n69, pe_1_4_0_n68, pe_1_4_0_n67,
         pe_1_4_0_n66, pe_1_4_0_n65, pe_1_4_0_n64, pe_1_4_0_n63, pe_1_4_0_n62,
         pe_1_4_0_n61, pe_1_4_0_n60, pe_1_4_0_n59, pe_1_4_0_n58, pe_1_4_0_n57,
         pe_1_4_0_n56, pe_1_4_0_n55, pe_1_4_0_n54, pe_1_4_0_n53, pe_1_4_0_n52,
         pe_1_4_0_n51, pe_1_4_0_n50, pe_1_4_0_n49, pe_1_4_0_n48, pe_1_4_0_n47,
         pe_1_4_0_n46, pe_1_4_0_n45, pe_1_4_0_n25, pe_1_4_0_n24, pe_1_4_0_n23,
         pe_1_4_0_n22, pe_1_4_0_n21, pe_1_4_0_n20, pe_1_4_0_n19, pe_1_4_0_n18,
         pe_1_4_0_n17, pe_1_4_0_n16, pe_1_4_0_n15, pe_1_4_0_n14, pe_1_4_0_n13,
         pe_1_4_0_n12, pe_1_4_0_n11, pe_1_4_0_n10, pe_1_4_0_n9, pe_1_4_0_n8,
         pe_1_4_0_n7, pe_1_4_0_n6, pe_1_4_0_n5, pe_1_4_0_n4, pe_1_4_0_n3,
         pe_1_4_0_n2, pe_1_4_0_n1, pe_1_4_0_n44, pe_1_4_0_n43, pe_1_4_0_n42,
         pe_1_4_0_n41, pe_1_4_0_n40, pe_1_4_0_n39, pe_1_4_0_n38, pe_1_4_0_n37,
         pe_1_4_0_n36, pe_1_4_0_n35, pe_1_4_0_n34, pe_1_4_0_n33, pe_1_4_0_n32,
         pe_1_4_0_n31, pe_1_4_0_n30, pe_1_4_0_n29, pe_1_4_0_n28, pe_1_4_0_n27,
         pe_1_4_0_n26, pe_1_4_0_net5056, pe_1_4_0_net5051, pe_1_4_0_net5046,
         pe_1_4_0_net5041, pe_1_4_0_net5036, pe_1_4_0_net5031,
         pe_1_4_0_net5026, pe_1_4_0_net5021, pe_1_4_0_net5016,
         pe_1_4_0_net5011, pe_1_4_0_net5006, pe_1_4_0_net5001,
         pe_1_4_0_net4995, pe_1_4_0_N90, pe_1_4_0_N85, pe_1_4_0_N84,
         pe_1_4_0_N83, pe_1_4_0_N82, pe_1_4_0_N81, pe_1_4_0_N80, pe_1_4_0_N79,
         pe_1_4_0_N77, pe_1_4_0_N76, pe_1_4_0_N75, pe_1_4_0_N74, pe_1_4_0_N73,
         pe_1_4_0_N72, pe_1_4_0_N71, pe_1_4_0_N70, pe_1_4_0_int_data_0_,
         pe_1_4_0_int_data_1_, pe_1_4_0_int_data_2_, pe_1_4_0_int_data_3_,
         pe_1_4_0_N64, pe_1_4_0_N63, pe_1_4_0_N62, pe_1_4_0_N61, pe_1_4_0_N60,
         pe_1_4_0_N59, pe_1_4_0_o_data_h_0_, pe_1_4_0_o_data_h_1_,
         pe_1_4_0_o_data_h_2_, pe_1_4_0_o_data_h_3_, pe_1_4_1_n90,
         pe_1_4_1_n89, pe_1_4_1_n88, pe_1_4_1_n87, pe_1_4_1_n86, pe_1_4_1_n85,
         pe_1_4_1_n84, pe_1_4_1_n83, pe_1_4_1_n82, pe_1_4_1_n81, pe_1_4_1_n80,
         pe_1_4_1_n79, pe_1_4_1_n78, pe_1_4_1_n77, pe_1_4_1_n76, pe_1_4_1_n75,
         pe_1_4_1_n74, pe_1_4_1_n73, pe_1_4_1_n72, pe_1_4_1_n71, pe_1_4_1_n70,
         pe_1_4_1_n69, pe_1_4_1_n68, pe_1_4_1_n67, pe_1_4_1_n66, pe_1_4_1_n65,
         pe_1_4_1_n64, pe_1_4_1_n63, pe_1_4_1_n62, pe_1_4_1_n61, pe_1_4_1_n60,
         pe_1_4_1_n59, pe_1_4_1_n58, pe_1_4_1_n57, pe_1_4_1_n56, pe_1_4_1_n55,
         pe_1_4_1_n54, pe_1_4_1_n53, pe_1_4_1_n52, pe_1_4_1_n51, pe_1_4_1_n50,
         pe_1_4_1_n49, pe_1_4_1_n48, pe_1_4_1_n47, pe_1_4_1_n46, pe_1_4_1_n45,
         pe_1_4_1_n25, pe_1_4_1_n24, pe_1_4_1_n23, pe_1_4_1_n22, pe_1_4_1_n21,
         pe_1_4_1_n20, pe_1_4_1_n19, pe_1_4_1_n18, pe_1_4_1_n17, pe_1_4_1_n16,
         pe_1_4_1_n15, pe_1_4_1_n14, pe_1_4_1_n13, pe_1_4_1_n12, pe_1_4_1_n11,
         pe_1_4_1_n10, pe_1_4_1_n9, pe_1_4_1_n8, pe_1_4_1_n7, pe_1_4_1_n6,
         pe_1_4_1_n5, pe_1_4_1_n4, pe_1_4_1_n3, pe_1_4_1_n2, pe_1_4_1_n1,
         pe_1_4_1_n44, pe_1_4_1_n43, pe_1_4_1_n42, pe_1_4_1_n41, pe_1_4_1_n40,
         pe_1_4_1_n39, pe_1_4_1_n38, pe_1_4_1_n37, pe_1_4_1_n36, pe_1_4_1_n35,
         pe_1_4_1_n34, pe_1_4_1_n33, pe_1_4_1_n32, pe_1_4_1_n31, pe_1_4_1_n30,
         pe_1_4_1_n29, pe_1_4_1_n28, pe_1_4_1_n27, pe_1_4_1_n26,
         pe_1_4_1_net4978, pe_1_4_1_net4973, pe_1_4_1_net4968,
         pe_1_4_1_net4963, pe_1_4_1_net4958, pe_1_4_1_net4953,
         pe_1_4_1_net4948, pe_1_4_1_net4943, pe_1_4_1_net4938,
         pe_1_4_1_net4933, pe_1_4_1_net4928, pe_1_4_1_net4923,
         pe_1_4_1_net4917, pe_1_4_1_N90, pe_1_4_1_N85, pe_1_4_1_N84,
         pe_1_4_1_N83, pe_1_4_1_N82, pe_1_4_1_N81, pe_1_4_1_N80, pe_1_4_1_N79,
         pe_1_4_1_N77, pe_1_4_1_N76, pe_1_4_1_N75, pe_1_4_1_N74, pe_1_4_1_N73,
         pe_1_4_1_N72, pe_1_4_1_N71, pe_1_4_1_N70, pe_1_4_1_int_data_0_,
         pe_1_4_1_int_data_1_, pe_1_4_1_int_data_2_, pe_1_4_1_int_data_3_,
         pe_1_4_1_N64, pe_1_4_1_N63, pe_1_4_1_N62, pe_1_4_1_N61, pe_1_4_1_N60,
         pe_1_4_1_N59, pe_1_4_2_n90, pe_1_4_2_n89, pe_1_4_2_n88, pe_1_4_2_n87,
         pe_1_4_2_n86, pe_1_4_2_n85, pe_1_4_2_n84, pe_1_4_2_n83, pe_1_4_2_n82,
         pe_1_4_2_n81, pe_1_4_2_n80, pe_1_4_2_n79, pe_1_4_2_n78, pe_1_4_2_n77,
         pe_1_4_2_n76, pe_1_4_2_n75, pe_1_4_2_n74, pe_1_4_2_n73, pe_1_4_2_n72,
         pe_1_4_2_n71, pe_1_4_2_n70, pe_1_4_2_n69, pe_1_4_2_n68, pe_1_4_2_n67,
         pe_1_4_2_n66, pe_1_4_2_n65, pe_1_4_2_n64, pe_1_4_2_n63, pe_1_4_2_n62,
         pe_1_4_2_n61, pe_1_4_2_n60, pe_1_4_2_n59, pe_1_4_2_n58, pe_1_4_2_n57,
         pe_1_4_2_n56, pe_1_4_2_n55, pe_1_4_2_n54, pe_1_4_2_n53, pe_1_4_2_n52,
         pe_1_4_2_n51, pe_1_4_2_n50, pe_1_4_2_n49, pe_1_4_2_n48, pe_1_4_2_n47,
         pe_1_4_2_n46, pe_1_4_2_n45, pe_1_4_2_n25, pe_1_4_2_n24, pe_1_4_2_n23,
         pe_1_4_2_n22, pe_1_4_2_n21, pe_1_4_2_n20, pe_1_4_2_n19, pe_1_4_2_n18,
         pe_1_4_2_n17, pe_1_4_2_n16, pe_1_4_2_n15, pe_1_4_2_n14, pe_1_4_2_n13,
         pe_1_4_2_n12, pe_1_4_2_n11, pe_1_4_2_n10, pe_1_4_2_n9, pe_1_4_2_n8,
         pe_1_4_2_n7, pe_1_4_2_n6, pe_1_4_2_n5, pe_1_4_2_n4, pe_1_4_2_n3,
         pe_1_4_2_n2, pe_1_4_2_n1, pe_1_4_2_n44, pe_1_4_2_n43, pe_1_4_2_n42,
         pe_1_4_2_n41, pe_1_4_2_n40, pe_1_4_2_n39, pe_1_4_2_n38, pe_1_4_2_n37,
         pe_1_4_2_n36, pe_1_4_2_n35, pe_1_4_2_n34, pe_1_4_2_n33, pe_1_4_2_n32,
         pe_1_4_2_n31, pe_1_4_2_n30, pe_1_4_2_n29, pe_1_4_2_n28, pe_1_4_2_n27,
         pe_1_4_2_n26, pe_1_4_2_net4900, pe_1_4_2_net4895, pe_1_4_2_net4890,
         pe_1_4_2_net4885, pe_1_4_2_net4880, pe_1_4_2_net4875,
         pe_1_4_2_net4870, pe_1_4_2_net4865, pe_1_4_2_net4860,
         pe_1_4_2_net4855, pe_1_4_2_net4850, pe_1_4_2_net4845,
         pe_1_4_2_net4839, pe_1_4_2_N90, pe_1_4_2_N85, pe_1_4_2_N84,
         pe_1_4_2_N83, pe_1_4_2_N82, pe_1_4_2_N81, pe_1_4_2_N80, pe_1_4_2_N79,
         pe_1_4_2_N77, pe_1_4_2_N76, pe_1_4_2_N75, pe_1_4_2_N74, pe_1_4_2_N73,
         pe_1_4_2_N72, pe_1_4_2_N71, pe_1_4_2_N70, pe_1_4_2_int_data_0_,
         pe_1_4_2_int_data_1_, pe_1_4_2_int_data_2_, pe_1_4_2_int_data_3_,
         pe_1_4_2_N64, pe_1_4_2_N63, pe_1_4_2_N62, pe_1_4_2_N61, pe_1_4_2_N60,
         pe_1_4_2_N59, pe_1_4_3_n90, pe_1_4_3_n89, pe_1_4_3_n88, pe_1_4_3_n87,
         pe_1_4_3_n86, pe_1_4_3_n85, pe_1_4_3_n84, pe_1_4_3_n83, pe_1_4_3_n82,
         pe_1_4_3_n81, pe_1_4_3_n80, pe_1_4_3_n79, pe_1_4_3_n78, pe_1_4_3_n77,
         pe_1_4_3_n76, pe_1_4_3_n75, pe_1_4_3_n74, pe_1_4_3_n73, pe_1_4_3_n72,
         pe_1_4_3_n71, pe_1_4_3_n70, pe_1_4_3_n69, pe_1_4_3_n68, pe_1_4_3_n67,
         pe_1_4_3_n66, pe_1_4_3_n65, pe_1_4_3_n64, pe_1_4_3_n63, pe_1_4_3_n62,
         pe_1_4_3_n61, pe_1_4_3_n60, pe_1_4_3_n59, pe_1_4_3_n58, pe_1_4_3_n57,
         pe_1_4_3_n56, pe_1_4_3_n55, pe_1_4_3_n54, pe_1_4_3_n53, pe_1_4_3_n52,
         pe_1_4_3_n51, pe_1_4_3_n50, pe_1_4_3_n49, pe_1_4_3_n48, pe_1_4_3_n47,
         pe_1_4_3_n46, pe_1_4_3_n45, pe_1_4_3_n25, pe_1_4_3_n24, pe_1_4_3_n23,
         pe_1_4_3_n22, pe_1_4_3_n21, pe_1_4_3_n20, pe_1_4_3_n19, pe_1_4_3_n18,
         pe_1_4_3_n17, pe_1_4_3_n16, pe_1_4_3_n15, pe_1_4_3_n14, pe_1_4_3_n13,
         pe_1_4_3_n12, pe_1_4_3_n11, pe_1_4_3_n10, pe_1_4_3_n9, pe_1_4_3_n8,
         pe_1_4_3_n7, pe_1_4_3_n6, pe_1_4_3_n5, pe_1_4_3_n4, pe_1_4_3_n3,
         pe_1_4_3_n2, pe_1_4_3_n1, pe_1_4_3_n44, pe_1_4_3_n43, pe_1_4_3_n42,
         pe_1_4_3_n41, pe_1_4_3_n40, pe_1_4_3_n39, pe_1_4_3_n38, pe_1_4_3_n37,
         pe_1_4_3_n36, pe_1_4_3_n35, pe_1_4_3_n34, pe_1_4_3_n33, pe_1_4_3_n32,
         pe_1_4_3_n31, pe_1_4_3_n30, pe_1_4_3_n29, pe_1_4_3_n28, pe_1_4_3_n27,
         pe_1_4_3_n26, pe_1_4_3_net4822, pe_1_4_3_net4817, pe_1_4_3_net4812,
         pe_1_4_3_net4807, pe_1_4_3_net4802, pe_1_4_3_net4797,
         pe_1_4_3_net4792, pe_1_4_3_net4787, pe_1_4_3_net4782,
         pe_1_4_3_net4777, pe_1_4_3_net4772, pe_1_4_3_net4767,
         pe_1_4_3_net4761, pe_1_4_3_N90, pe_1_4_3_N85, pe_1_4_3_N84,
         pe_1_4_3_N83, pe_1_4_3_N82, pe_1_4_3_N81, pe_1_4_3_N80, pe_1_4_3_N79,
         pe_1_4_3_N77, pe_1_4_3_N76, pe_1_4_3_N75, pe_1_4_3_N74, pe_1_4_3_N73,
         pe_1_4_3_N72, pe_1_4_3_N71, pe_1_4_3_N70, pe_1_4_3_int_data_0_,
         pe_1_4_3_int_data_1_, pe_1_4_3_int_data_2_, pe_1_4_3_int_data_3_,
         pe_1_4_3_N64, pe_1_4_3_N63, pe_1_4_3_N62, pe_1_4_3_N61, pe_1_4_3_N60,
         pe_1_4_3_N59, pe_1_4_4_n86, pe_1_4_4_n85, pe_1_4_4_n84, pe_1_4_4_n83,
         pe_1_4_4_n82, pe_1_4_4_n81, pe_1_4_4_n80, pe_1_4_4_n79, pe_1_4_4_n78,
         pe_1_4_4_n77, pe_1_4_4_n76, pe_1_4_4_n75, pe_1_4_4_n74, pe_1_4_4_n73,
         pe_1_4_4_n72, pe_1_4_4_n71, pe_1_4_4_n70, pe_1_4_4_n69, pe_1_4_4_n68,
         pe_1_4_4_n67, pe_1_4_4_n66, pe_1_4_4_n65, pe_1_4_4_n64, pe_1_4_4_n63,
         pe_1_4_4_n62, pe_1_4_4_n61, pe_1_4_4_n60, pe_1_4_4_n59, pe_1_4_4_n58,
         pe_1_4_4_n57, pe_1_4_4_n56, pe_1_4_4_n55, pe_1_4_4_n54, pe_1_4_4_n53,
         pe_1_4_4_n52, pe_1_4_4_n51, pe_1_4_4_n50, pe_1_4_4_n49, pe_1_4_4_n48,
         pe_1_4_4_n47, pe_1_4_4_n46, pe_1_4_4_n45, pe_1_4_4_n25, pe_1_4_4_n24,
         pe_1_4_4_n23, pe_1_4_4_n22, pe_1_4_4_n21, pe_1_4_4_n20, pe_1_4_4_n19,
         pe_1_4_4_n18, pe_1_4_4_n17, pe_1_4_4_n16, pe_1_4_4_n15, pe_1_4_4_n14,
         pe_1_4_4_n13, pe_1_4_4_n12, pe_1_4_4_n11, pe_1_4_4_n10, pe_1_4_4_n9,
         pe_1_4_4_n8, pe_1_4_4_n7, pe_1_4_4_n6, pe_1_4_4_n5, pe_1_4_4_n4,
         pe_1_4_4_n3, pe_1_4_4_n2, pe_1_4_4_n1, pe_1_4_4_n44, pe_1_4_4_n43,
         pe_1_4_4_n42, pe_1_4_4_n41, pe_1_4_4_n40, pe_1_4_4_n39, pe_1_4_4_n38,
         pe_1_4_4_n37, pe_1_4_4_n36, pe_1_4_4_n35, pe_1_4_4_n34, pe_1_4_4_n33,
         pe_1_4_4_n32, pe_1_4_4_n31, pe_1_4_4_n30, pe_1_4_4_n29, pe_1_4_4_n28,
         pe_1_4_4_n27, pe_1_4_4_n26, pe_1_4_4_net4744, pe_1_4_4_net4739,
         pe_1_4_4_net4734, pe_1_4_4_net4729, pe_1_4_4_net4724,
         pe_1_4_4_net4719, pe_1_4_4_net4714, pe_1_4_4_net4709,
         pe_1_4_4_net4704, pe_1_4_4_net4699, pe_1_4_4_net4694,
         pe_1_4_4_net4689, pe_1_4_4_net4683, pe_1_4_4_N90, pe_1_4_4_N85,
         pe_1_4_4_N84, pe_1_4_4_N83, pe_1_4_4_N82, pe_1_4_4_N81, pe_1_4_4_N80,
         pe_1_4_4_N79, pe_1_4_4_N77, pe_1_4_4_N76, pe_1_4_4_N75, pe_1_4_4_N74,
         pe_1_4_4_N73, pe_1_4_4_N72, pe_1_4_4_N71, pe_1_4_4_N70,
         pe_1_4_4_int_data_0_, pe_1_4_4_int_data_1_, pe_1_4_4_int_data_2_,
         pe_1_4_4_int_data_3_, pe_1_4_4_N64, pe_1_4_4_N63, pe_1_4_4_N62,
         pe_1_4_4_N61, pe_1_4_4_N60, pe_1_4_4_N59, pe_1_4_5_n87, pe_1_4_5_n86,
         pe_1_4_5_n85, pe_1_4_5_n84, pe_1_4_5_n83, pe_1_4_5_n82, pe_1_4_5_n81,
         pe_1_4_5_n80, pe_1_4_5_n79, pe_1_4_5_n78, pe_1_4_5_n77, pe_1_4_5_n76,
         pe_1_4_5_n75, pe_1_4_5_n74, pe_1_4_5_n73, pe_1_4_5_n72, pe_1_4_5_n71,
         pe_1_4_5_n70, pe_1_4_5_n69, pe_1_4_5_n68, pe_1_4_5_n67, pe_1_4_5_n66,
         pe_1_4_5_n65, pe_1_4_5_n64, pe_1_4_5_n63, pe_1_4_5_n62, pe_1_4_5_n61,
         pe_1_4_5_n60, pe_1_4_5_n59, pe_1_4_5_n58, pe_1_4_5_n57, pe_1_4_5_n56,
         pe_1_4_5_n55, pe_1_4_5_n54, pe_1_4_5_n53, pe_1_4_5_n52, pe_1_4_5_n51,
         pe_1_4_5_n50, pe_1_4_5_n49, pe_1_4_5_n48, pe_1_4_5_n47, pe_1_4_5_n46,
         pe_1_4_5_n45, pe_1_4_5_n25, pe_1_4_5_n24, pe_1_4_5_n23, pe_1_4_5_n22,
         pe_1_4_5_n21, pe_1_4_5_n20, pe_1_4_5_n19, pe_1_4_5_n18, pe_1_4_5_n17,
         pe_1_4_5_n16, pe_1_4_5_n15, pe_1_4_5_n14, pe_1_4_5_n13, pe_1_4_5_n12,
         pe_1_4_5_n11, pe_1_4_5_n10, pe_1_4_5_n9, pe_1_4_5_n8, pe_1_4_5_n7,
         pe_1_4_5_n6, pe_1_4_5_n5, pe_1_4_5_n4, pe_1_4_5_n3, pe_1_4_5_n2,
         pe_1_4_5_n1, pe_1_4_5_n44, pe_1_4_5_n43, pe_1_4_5_n42, pe_1_4_5_n41,
         pe_1_4_5_n40, pe_1_4_5_n39, pe_1_4_5_n38, pe_1_4_5_n37, pe_1_4_5_n36,
         pe_1_4_5_n35, pe_1_4_5_n34, pe_1_4_5_n33, pe_1_4_5_n32, pe_1_4_5_n31,
         pe_1_4_5_n30, pe_1_4_5_n29, pe_1_4_5_n28, pe_1_4_5_n27, pe_1_4_5_n26,
         pe_1_4_5_net4666, pe_1_4_5_net4661, pe_1_4_5_net4656,
         pe_1_4_5_net4651, pe_1_4_5_net4646, pe_1_4_5_net4641,
         pe_1_4_5_net4636, pe_1_4_5_net4631, pe_1_4_5_net4626,
         pe_1_4_5_net4621, pe_1_4_5_net4616, pe_1_4_5_net4611,
         pe_1_4_5_net4605, pe_1_4_5_N90, pe_1_4_5_N85, pe_1_4_5_N84,
         pe_1_4_5_N83, pe_1_4_5_N82, pe_1_4_5_N81, pe_1_4_5_N80, pe_1_4_5_N79,
         pe_1_4_5_N77, pe_1_4_5_N76, pe_1_4_5_N75, pe_1_4_5_N74, pe_1_4_5_N73,
         pe_1_4_5_N72, pe_1_4_5_N71, pe_1_4_5_N70, pe_1_4_5_int_data_0_,
         pe_1_4_5_int_data_1_, pe_1_4_5_int_data_2_, pe_1_4_5_int_data_3_,
         pe_1_4_5_N64, pe_1_4_5_N63, pe_1_4_5_N62, pe_1_4_5_N61, pe_1_4_5_N60,
         pe_1_4_5_N59, pe_1_4_6_n88, pe_1_4_6_n87, pe_1_4_6_n86, pe_1_4_6_n85,
         pe_1_4_6_n84, pe_1_4_6_n83, pe_1_4_6_n82, pe_1_4_6_n81, pe_1_4_6_n80,
         pe_1_4_6_n79, pe_1_4_6_n78, pe_1_4_6_n77, pe_1_4_6_n76, pe_1_4_6_n75,
         pe_1_4_6_n74, pe_1_4_6_n73, pe_1_4_6_n72, pe_1_4_6_n71, pe_1_4_6_n70,
         pe_1_4_6_n69, pe_1_4_6_n68, pe_1_4_6_n67, pe_1_4_6_n66, pe_1_4_6_n65,
         pe_1_4_6_n64, pe_1_4_6_n63, pe_1_4_6_n62, pe_1_4_6_n61, pe_1_4_6_n60,
         pe_1_4_6_n59, pe_1_4_6_n58, pe_1_4_6_n57, pe_1_4_6_n56, pe_1_4_6_n55,
         pe_1_4_6_n54, pe_1_4_6_n53, pe_1_4_6_n52, pe_1_4_6_n51, pe_1_4_6_n50,
         pe_1_4_6_n49, pe_1_4_6_n48, pe_1_4_6_n47, pe_1_4_6_n46, pe_1_4_6_n45,
         pe_1_4_6_n25, pe_1_4_6_n24, pe_1_4_6_n23, pe_1_4_6_n22, pe_1_4_6_n21,
         pe_1_4_6_n20, pe_1_4_6_n19, pe_1_4_6_n18, pe_1_4_6_n17, pe_1_4_6_n16,
         pe_1_4_6_n15, pe_1_4_6_n14, pe_1_4_6_n13, pe_1_4_6_n12, pe_1_4_6_n11,
         pe_1_4_6_n10, pe_1_4_6_n9, pe_1_4_6_n8, pe_1_4_6_n7, pe_1_4_6_n6,
         pe_1_4_6_n5, pe_1_4_6_n4, pe_1_4_6_n3, pe_1_4_6_n2, pe_1_4_6_n1,
         pe_1_4_6_n44, pe_1_4_6_n43, pe_1_4_6_n42, pe_1_4_6_n41, pe_1_4_6_n40,
         pe_1_4_6_n39, pe_1_4_6_n38, pe_1_4_6_n37, pe_1_4_6_n36, pe_1_4_6_n35,
         pe_1_4_6_n34, pe_1_4_6_n33, pe_1_4_6_n32, pe_1_4_6_n31, pe_1_4_6_n30,
         pe_1_4_6_n29, pe_1_4_6_n28, pe_1_4_6_n27, pe_1_4_6_n26,
         pe_1_4_6_net4588, pe_1_4_6_net4583, pe_1_4_6_net4578,
         pe_1_4_6_net4573, pe_1_4_6_net4568, pe_1_4_6_net4563,
         pe_1_4_6_net4558, pe_1_4_6_net4553, pe_1_4_6_net4548,
         pe_1_4_6_net4543, pe_1_4_6_net4538, pe_1_4_6_net4533,
         pe_1_4_6_net4527, pe_1_4_6_N90, pe_1_4_6_N85, pe_1_4_6_N84,
         pe_1_4_6_N83, pe_1_4_6_N82, pe_1_4_6_N81, pe_1_4_6_N80, pe_1_4_6_N79,
         pe_1_4_6_N77, pe_1_4_6_N76, pe_1_4_6_N75, pe_1_4_6_N74, pe_1_4_6_N73,
         pe_1_4_6_N72, pe_1_4_6_N71, pe_1_4_6_N70, pe_1_4_6_int_data_0_,
         pe_1_4_6_int_data_1_, pe_1_4_6_int_data_2_, pe_1_4_6_int_data_3_,
         pe_1_4_6_N64, pe_1_4_6_N63, pe_1_4_6_N62, pe_1_4_6_N61, pe_1_4_6_N60,
         pe_1_4_6_N59, pe_1_4_7_n88, pe_1_4_7_n87, pe_1_4_7_n86, pe_1_4_7_n85,
         pe_1_4_7_n84, pe_1_4_7_n83, pe_1_4_7_n82, pe_1_4_7_n81, pe_1_4_7_n80,
         pe_1_4_7_n79, pe_1_4_7_n78, pe_1_4_7_n77, pe_1_4_7_n76, pe_1_4_7_n75,
         pe_1_4_7_n74, pe_1_4_7_n73, pe_1_4_7_n72, pe_1_4_7_n71, pe_1_4_7_n70,
         pe_1_4_7_n69, pe_1_4_7_n68, pe_1_4_7_n67, pe_1_4_7_n66, pe_1_4_7_n65,
         pe_1_4_7_n64, pe_1_4_7_n63, pe_1_4_7_n62, pe_1_4_7_n61, pe_1_4_7_n60,
         pe_1_4_7_n59, pe_1_4_7_n58, pe_1_4_7_n57, pe_1_4_7_n56, pe_1_4_7_n55,
         pe_1_4_7_n54, pe_1_4_7_n53, pe_1_4_7_n52, pe_1_4_7_n51, pe_1_4_7_n50,
         pe_1_4_7_n49, pe_1_4_7_n48, pe_1_4_7_n47, pe_1_4_7_n46, pe_1_4_7_n45,
         pe_1_4_7_n25, pe_1_4_7_n24, pe_1_4_7_n23, pe_1_4_7_n22, pe_1_4_7_n21,
         pe_1_4_7_n20, pe_1_4_7_n19, pe_1_4_7_n18, pe_1_4_7_n17, pe_1_4_7_n16,
         pe_1_4_7_n15, pe_1_4_7_n14, pe_1_4_7_n13, pe_1_4_7_n12, pe_1_4_7_n11,
         pe_1_4_7_n10, pe_1_4_7_n9, pe_1_4_7_n8, pe_1_4_7_n7, pe_1_4_7_n6,
         pe_1_4_7_n5, pe_1_4_7_n4, pe_1_4_7_n3, pe_1_4_7_n2, pe_1_4_7_n1,
         pe_1_4_7_n44, pe_1_4_7_n43, pe_1_4_7_n42, pe_1_4_7_n41, pe_1_4_7_n40,
         pe_1_4_7_n39, pe_1_4_7_n38, pe_1_4_7_n37, pe_1_4_7_n36, pe_1_4_7_n35,
         pe_1_4_7_n34, pe_1_4_7_n33, pe_1_4_7_n32, pe_1_4_7_n31, pe_1_4_7_n30,
         pe_1_4_7_n29, pe_1_4_7_n28, pe_1_4_7_n27, pe_1_4_7_n26,
         pe_1_4_7_net4510, pe_1_4_7_net4505, pe_1_4_7_net4500,
         pe_1_4_7_net4495, pe_1_4_7_net4490, pe_1_4_7_net4485,
         pe_1_4_7_net4480, pe_1_4_7_net4475, pe_1_4_7_net4470,
         pe_1_4_7_net4465, pe_1_4_7_net4460, pe_1_4_7_net4455,
         pe_1_4_7_net4449, pe_1_4_7_N90, pe_1_4_7_N85, pe_1_4_7_N84,
         pe_1_4_7_N83, pe_1_4_7_N82, pe_1_4_7_N81, pe_1_4_7_N80, pe_1_4_7_N79,
         pe_1_4_7_N77, pe_1_4_7_N76, pe_1_4_7_N75, pe_1_4_7_N74, pe_1_4_7_N73,
         pe_1_4_7_N72, pe_1_4_7_N71, pe_1_4_7_N70, pe_1_4_7_int_data_0_,
         pe_1_4_7_int_data_1_, pe_1_4_7_int_data_2_, pe_1_4_7_int_data_3_,
         pe_1_4_7_N64, pe_1_4_7_N63, pe_1_4_7_N62, pe_1_4_7_N61, pe_1_4_7_N60,
         pe_1_4_7_N59, pe_1_5_0_n89, pe_1_5_0_n88, pe_1_5_0_n87, pe_1_5_0_n86,
         pe_1_5_0_n85, pe_1_5_0_n84, pe_1_5_0_n83, pe_1_5_0_n82, pe_1_5_0_n81,
         pe_1_5_0_n80, pe_1_5_0_n79, pe_1_5_0_n78, pe_1_5_0_n77, pe_1_5_0_n76,
         pe_1_5_0_n75, pe_1_5_0_n74, pe_1_5_0_n73, pe_1_5_0_n72, pe_1_5_0_n71,
         pe_1_5_0_n70, pe_1_5_0_n69, pe_1_5_0_n68, pe_1_5_0_n67, pe_1_5_0_n66,
         pe_1_5_0_n65, pe_1_5_0_n64, pe_1_5_0_n63, pe_1_5_0_n62, pe_1_5_0_n61,
         pe_1_5_0_n60, pe_1_5_0_n59, pe_1_5_0_n58, pe_1_5_0_n57, pe_1_5_0_n56,
         pe_1_5_0_n55, pe_1_5_0_n54, pe_1_5_0_n53, pe_1_5_0_n52, pe_1_5_0_n51,
         pe_1_5_0_n50, pe_1_5_0_n49, pe_1_5_0_n48, pe_1_5_0_n47, pe_1_5_0_n46,
         pe_1_5_0_n45, pe_1_5_0_n25, pe_1_5_0_n24, pe_1_5_0_n23, pe_1_5_0_n22,
         pe_1_5_0_n21, pe_1_5_0_n20, pe_1_5_0_n19, pe_1_5_0_n18, pe_1_5_0_n17,
         pe_1_5_0_n16, pe_1_5_0_n15, pe_1_5_0_n14, pe_1_5_0_n13, pe_1_5_0_n12,
         pe_1_5_0_n11, pe_1_5_0_n10, pe_1_5_0_n9, pe_1_5_0_n8, pe_1_5_0_n7,
         pe_1_5_0_n6, pe_1_5_0_n5, pe_1_5_0_n4, pe_1_5_0_n3, pe_1_5_0_n2,
         pe_1_5_0_n1, pe_1_5_0_n44, pe_1_5_0_n43, pe_1_5_0_n42, pe_1_5_0_n41,
         pe_1_5_0_n40, pe_1_5_0_n39, pe_1_5_0_n38, pe_1_5_0_n37, pe_1_5_0_n36,
         pe_1_5_0_n35, pe_1_5_0_n34, pe_1_5_0_n33, pe_1_5_0_n32, pe_1_5_0_n31,
         pe_1_5_0_n30, pe_1_5_0_n29, pe_1_5_0_n28, pe_1_5_0_n27, pe_1_5_0_n26,
         pe_1_5_0_net4432, pe_1_5_0_net4427, pe_1_5_0_net4422,
         pe_1_5_0_net4417, pe_1_5_0_net4412, pe_1_5_0_net4407,
         pe_1_5_0_net4402, pe_1_5_0_net4397, pe_1_5_0_net4392,
         pe_1_5_0_net4387, pe_1_5_0_net4382, pe_1_5_0_net4377,
         pe_1_5_0_net4371, pe_1_5_0_N90, pe_1_5_0_N85, pe_1_5_0_N84,
         pe_1_5_0_N83, pe_1_5_0_N82, pe_1_5_0_N81, pe_1_5_0_N80, pe_1_5_0_N79,
         pe_1_5_0_N77, pe_1_5_0_N76, pe_1_5_0_N75, pe_1_5_0_N74, pe_1_5_0_N73,
         pe_1_5_0_N72, pe_1_5_0_N71, pe_1_5_0_N70, pe_1_5_0_int_data_0_,
         pe_1_5_0_int_data_1_, pe_1_5_0_int_data_2_, pe_1_5_0_int_data_3_,
         pe_1_5_0_N64, pe_1_5_0_N63, pe_1_5_0_N62, pe_1_5_0_N61, pe_1_5_0_N60,
         pe_1_5_0_N59, pe_1_5_0_o_data_h_0_, pe_1_5_0_o_data_h_1_,
         pe_1_5_0_o_data_h_2_, pe_1_5_0_o_data_h_3_, pe_1_5_1_n90,
         pe_1_5_1_n89, pe_1_5_1_n88, pe_1_5_1_n87, pe_1_5_1_n86, pe_1_5_1_n85,
         pe_1_5_1_n84, pe_1_5_1_n83, pe_1_5_1_n82, pe_1_5_1_n81, pe_1_5_1_n80,
         pe_1_5_1_n79, pe_1_5_1_n78, pe_1_5_1_n77, pe_1_5_1_n76, pe_1_5_1_n75,
         pe_1_5_1_n74, pe_1_5_1_n73, pe_1_5_1_n72, pe_1_5_1_n71, pe_1_5_1_n70,
         pe_1_5_1_n69, pe_1_5_1_n68, pe_1_5_1_n67, pe_1_5_1_n66, pe_1_5_1_n65,
         pe_1_5_1_n64, pe_1_5_1_n63, pe_1_5_1_n62, pe_1_5_1_n61, pe_1_5_1_n60,
         pe_1_5_1_n59, pe_1_5_1_n58, pe_1_5_1_n57, pe_1_5_1_n56, pe_1_5_1_n55,
         pe_1_5_1_n54, pe_1_5_1_n53, pe_1_5_1_n52, pe_1_5_1_n51, pe_1_5_1_n50,
         pe_1_5_1_n49, pe_1_5_1_n48, pe_1_5_1_n47, pe_1_5_1_n46, pe_1_5_1_n45,
         pe_1_5_1_n25, pe_1_5_1_n24, pe_1_5_1_n23, pe_1_5_1_n22, pe_1_5_1_n21,
         pe_1_5_1_n20, pe_1_5_1_n19, pe_1_5_1_n18, pe_1_5_1_n17, pe_1_5_1_n16,
         pe_1_5_1_n15, pe_1_5_1_n14, pe_1_5_1_n13, pe_1_5_1_n12, pe_1_5_1_n11,
         pe_1_5_1_n10, pe_1_5_1_n9, pe_1_5_1_n8, pe_1_5_1_n7, pe_1_5_1_n6,
         pe_1_5_1_n5, pe_1_5_1_n4, pe_1_5_1_n3, pe_1_5_1_n2, pe_1_5_1_n1,
         pe_1_5_1_n44, pe_1_5_1_n43, pe_1_5_1_n42, pe_1_5_1_n41, pe_1_5_1_n40,
         pe_1_5_1_n39, pe_1_5_1_n38, pe_1_5_1_n37, pe_1_5_1_n36, pe_1_5_1_n35,
         pe_1_5_1_n34, pe_1_5_1_n33, pe_1_5_1_n32, pe_1_5_1_n31, pe_1_5_1_n30,
         pe_1_5_1_n29, pe_1_5_1_n28, pe_1_5_1_n27, pe_1_5_1_n26,
         pe_1_5_1_net4354, pe_1_5_1_net4349, pe_1_5_1_net4344,
         pe_1_5_1_net4339, pe_1_5_1_net4334, pe_1_5_1_net4329,
         pe_1_5_1_net4324, pe_1_5_1_net4319, pe_1_5_1_net4314,
         pe_1_5_1_net4309, pe_1_5_1_net4304, pe_1_5_1_net4299,
         pe_1_5_1_net4293, pe_1_5_1_N90, pe_1_5_1_N85, pe_1_5_1_N84,
         pe_1_5_1_N83, pe_1_5_1_N82, pe_1_5_1_N81, pe_1_5_1_N80, pe_1_5_1_N79,
         pe_1_5_1_N77, pe_1_5_1_N76, pe_1_5_1_N75, pe_1_5_1_N74, pe_1_5_1_N73,
         pe_1_5_1_N72, pe_1_5_1_N71, pe_1_5_1_N70, pe_1_5_1_int_data_0_,
         pe_1_5_1_int_data_1_, pe_1_5_1_int_data_2_, pe_1_5_1_int_data_3_,
         pe_1_5_1_N64, pe_1_5_1_N63, pe_1_5_1_N62, pe_1_5_1_N61, pe_1_5_1_N60,
         pe_1_5_1_N59, pe_1_5_2_n90, pe_1_5_2_n89, pe_1_5_2_n88, pe_1_5_2_n87,
         pe_1_5_2_n86, pe_1_5_2_n85, pe_1_5_2_n84, pe_1_5_2_n83, pe_1_5_2_n82,
         pe_1_5_2_n81, pe_1_5_2_n80, pe_1_5_2_n79, pe_1_5_2_n78, pe_1_5_2_n77,
         pe_1_5_2_n76, pe_1_5_2_n75, pe_1_5_2_n74, pe_1_5_2_n73, pe_1_5_2_n72,
         pe_1_5_2_n71, pe_1_5_2_n70, pe_1_5_2_n69, pe_1_5_2_n68, pe_1_5_2_n67,
         pe_1_5_2_n66, pe_1_5_2_n65, pe_1_5_2_n64, pe_1_5_2_n63, pe_1_5_2_n62,
         pe_1_5_2_n61, pe_1_5_2_n60, pe_1_5_2_n59, pe_1_5_2_n58, pe_1_5_2_n57,
         pe_1_5_2_n56, pe_1_5_2_n55, pe_1_5_2_n54, pe_1_5_2_n53, pe_1_5_2_n52,
         pe_1_5_2_n51, pe_1_5_2_n50, pe_1_5_2_n49, pe_1_5_2_n48, pe_1_5_2_n47,
         pe_1_5_2_n46, pe_1_5_2_n45, pe_1_5_2_n25, pe_1_5_2_n24, pe_1_5_2_n23,
         pe_1_5_2_n22, pe_1_5_2_n21, pe_1_5_2_n20, pe_1_5_2_n19, pe_1_5_2_n18,
         pe_1_5_2_n17, pe_1_5_2_n16, pe_1_5_2_n15, pe_1_5_2_n14, pe_1_5_2_n13,
         pe_1_5_2_n12, pe_1_5_2_n11, pe_1_5_2_n10, pe_1_5_2_n9, pe_1_5_2_n8,
         pe_1_5_2_n7, pe_1_5_2_n6, pe_1_5_2_n5, pe_1_5_2_n4, pe_1_5_2_n3,
         pe_1_5_2_n2, pe_1_5_2_n1, pe_1_5_2_n44, pe_1_5_2_n43, pe_1_5_2_n42,
         pe_1_5_2_n41, pe_1_5_2_n40, pe_1_5_2_n39, pe_1_5_2_n38, pe_1_5_2_n37,
         pe_1_5_2_n36, pe_1_5_2_n35, pe_1_5_2_n34, pe_1_5_2_n33, pe_1_5_2_n32,
         pe_1_5_2_n31, pe_1_5_2_n30, pe_1_5_2_n29, pe_1_5_2_n28, pe_1_5_2_n27,
         pe_1_5_2_n26, pe_1_5_2_net4276, pe_1_5_2_net4271, pe_1_5_2_net4266,
         pe_1_5_2_net4261, pe_1_5_2_net4256, pe_1_5_2_net4251,
         pe_1_5_2_net4246, pe_1_5_2_net4241, pe_1_5_2_net4236,
         pe_1_5_2_net4231, pe_1_5_2_net4226, pe_1_5_2_net4221,
         pe_1_5_2_net4215, pe_1_5_2_N90, pe_1_5_2_N85, pe_1_5_2_N84,
         pe_1_5_2_N83, pe_1_5_2_N82, pe_1_5_2_N81, pe_1_5_2_N80, pe_1_5_2_N79,
         pe_1_5_2_N77, pe_1_5_2_N76, pe_1_5_2_N75, pe_1_5_2_N74, pe_1_5_2_N73,
         pe_1_5_2_N72, pe_1_5_2_N71, pe_1_5_2_N70, pe_1_5_2_int_data_0_,
         pe_1_5_2_int_data_1_, pe_1_5_2_int_data_2_, pe_1_5_2_int_data_3_,
         pe_1_5_2_N64, pe_1_5_2_N63, pe_1_5_2_N62, pe_1_5_2_N61, pe_1_5_2_N60,
         pe_1_5_2_N59, pe_1_5_3_n90, pe_1_5_3_n89, pe_1_5_3_n88, pe_1_5_3_n87,
         pe_1_5_3_n86, pe_1_5_3_n85, pe_1_5_3_n84, pe_1_5_3_n83, pe_1_5_3_n82,
         pe_1_5_3_n81, pe_1_5_3_n80, pe_1_5_3_n79, pe_1_5_3_n78, pe_1_5_3_n77,
         pe_1_5_3_n76, pe_1_5_3_n75, pe_1_5_3_n74, pe_1_5_3_n73, pe_1_5_3_n72,
         pe_1_5_3_n71, pe_1_5_3_n70, pe_1_5_3_n69, pe_1_5_3_n68, pe_1_5_3_n67,
         pe_1_5_3_n66, pe_1_5_3_n65, pe_1_5_3_n64, pe_1_5_3_n63, pe_1_5_3_n62,
         pe_1_5_3_n61, pe_1_5_3_n60, pe_1_5_3_n59, pe_1_5_3_n58, pe_1_5_3_n57,
         pe_1_5_3_n56, pe_1_5_3_n55, pe_1_5_3_n54, pe_1_5_3_n53, pe_1_5_3_n52,
         pe_1_5_3_n51, pe_1_5_3_n50, pe_1_5_3_n49, pe_1_5_3_n48, pe_1_5_3_n47,
         pe_1_5_3_n46, pe_1_5_3_n45, pe_1_5_3_n25, pe_1_5_3_n24, pe_1_5_3_n23,
         pe_1_5_3_n22, pe_1_5_3_n21, pe_1_5_3_n20, pe_1_5_3_n19, pe_1_5_3_n18,
         pe_1_5_3_n17, pe_1_5_3_n16, pe_1_5_3_n15, pe_1_5_3_n14, pe_1_5_3_n13,
         pe_1_5_3_n12, pe_1_5_3_n11, pe_1_5_3_n10, pe_1_5_3_n9, pe_1_5_3_n8,
         pe_1_5_3_n7, pe_1_5_3_n6, pe_1_5_3_n5, pe_1_5_3_n4, pe_1_5_3_n3,
         pe_1_5_3_n2, pe_1_5_3_n1, pe_1_5_3_n44, pe_1_5_3_n43, pe_1_5_3_n42,
         pe_1_5_3_n41, pe_1_5_3_n40, pe_1_5_3_n39, pe_1_5_3_n38, pe_1_5_3_n37,
         pe_1_5_3_n36, pe_1_5_3_n35, pe_1_5_3_n34, pe_1_5_3_n33, pe_1_5_3_n32,
         pe_1_5_3_n31, pe_1_5_3_n30, pe_1_5_3_n29, pe_1_5_3_n28, pe_1_5_3_n27,
         pe_1_5_3_n26, pe_1_5_3_net4198, pe_1_5_3_net4193, pe_1_5_3_net4188,
         pe_1_5_3_net4183, pe_1_5_3_net4178, pe_1_5_3_net4173,
         pe_1_5_3_net4168, pe_1_5_3_net4163, pe_1_5_3_net4158,
         pe_1_5_3_net4153, pe_1_5_3_net4148, pe_1_5_3_net4143,
         pe_1_5_3_net4137, pe_1_5_3_N90, pe_1_5_3_N85, pe_1_5_3_N84,
         pe_1_5_3_N83, pe_1_5_3_N82, pe_1_5_3_N81, pe_1_5_3_N80, pe_1_5_3_N79,
         pe_1_5_3_N77, pe_1_5_3_N76, pe_1_5_3_N75, pe_1_5_3_N74, pe_1_5_3_N73,
         pe_1_5_3_N72, pe_1_5_3_N71, pe_1_5_3_N70, pe_1_5_3_int_data_0_,
         pe_1_5_3_int_data_1_, pe_1_5_3_int_data_2_, pe_1_5_3_int_data_3_,
         pe_1_5_3_N64, pe_1_5_3_N63, pe_1_5_3_N62, pe_1_5_3_N61, pe_1_5_3_N60,
         pe_1_5_3_N59, pe_1_5_4_n90, pe_1_5_4_n89, pe_1_5_4_n88, pe_1_5_4_n87,
         pe_1_5_4_n86, pe_1_5_4_n85, pe_1_5_4_n84, pe_1_5_4_n83, pe_1_5_4_n82,
         pe_1_5_4_n81, pe_1_5_4_n80, pe_1_5_4_n79, pe_1_5_4_n78, pe_1_5_4_n77,
         pe_1_5_4_n76, pe_1_5_4_n75, pe_1_5_4_n74, pe_1_5_4_n73, pe_1_5_4_n72,
         pe_1_5_4_n71, pe_1_5_4_n70, pe_1_5_4_n69, pe_1_5_4_n68, pe_1_5_4_n67,
         pe_1_5_4_n66, pe_1_5_4_n65, pe_1_5_4_n64, pe_1_5_4_n63, pe_1_5_4_n62,
         pe_1_5_4_n61, pe_1_5_4_n60, pe_1_5_4_n59, pe_1_5_4_n58, pe_1_5_4_n57,
         pe_1_5_4_n56, pe_1_5_4_n55, pe_1_5_4_n54, pe_1_5_4_n53, pe_1_5_4_n52,
         pe_1_5_4_n51, pe_1_5_4_n50, pe_1_5_4_n49, pe_1_5_4_n48, pe_1_5_4_n47,
         pe_1_5_4_n46, pe_1_5_4_n45, pe_1_5_4_n25, pe_1_5_4_n24, pe_1_5_4_n23,
         pe_1_5_4_n22, pe_1_5_4_n21, pe_1_5_4_n20, pe_1_5_4_n19, pe_1_5_4_n18,
         pe_1_5_4_n17, pe_1_5_4_n16, pe_1_5_4_n15, pe_1_5_4_n14, pe_1_5_4_n13,
         pe_1_5_4_n12, pe_1_5_4_n11, pe_1_5_4_n10, pe_1_5_4_n9, pe_1_5_4_n8,
         pe_1_5_4_n7, pe_1_5_4_n6, pe_1_5_4_n5, pe_1_5_4_n4, pe_1_5_4_n3,
         pe_1_5_4_n2, pe_1_5_4_n1, pe_1_5_4_n44, pe_1_5_4_n43, pe_1_5_4_n42,
         pe_1_5_4_n41, pe_1_5_4_n40, pe_1_5_4_n39, pe_1_5_4_n38, pe_1_5_4_n37,
         pe_1_5_4_n36, pe_1_5_4_n35, pe_1_5_4_n34, pe_1_5_4_n33, pe_1_5_4_n32,
         pe_1_5_4_n31, pe_1_5_4_n30, pe_1_5_4_n29, pe_1_5_4_n28, pe_1_5_4_n27,
         pe_1_5_4_n26, pe_1_5_4_net4120, pe_1_5_4_net4115, pe_1_5_4_net4110,
         pe_1_5_4_net4105, pe_1_5_4_net4100, pe_1_5_4_net4095,
         pe_1_5_4_net4090, pe_1_5_4_net4085, pe_1_5_4_net4080,
         pe_1_5_4_net4075, pe_1_5_4_net4070, pe_1_5_4_net4065,
         pe_1_5_4_net4059, pe_1_5_4_N90, pe_1_5_4_N85, pe_1_5_4_N84,
         pe_1_5_4_N83, pe_1_5_4_N82, pe_1_5_4_N81, pe_1_5_4_N80, pe_1_5_4_N79,
         pe_1_5_4_N77, pe_1_5_4_N76, pe_1_5_4_N75, pe_1_5_4_N74, pe_1_5_4_N73,
         pe_1_5_4_N72, pe_1_5_4_N71, pe_1_5_4_N70, pe_1_5_4_int_data_0_,
         pe_1_5_4_int_data_1_, pe_1_5_4_int_data_2_, pe_1_5_4_int_data_3_,
         pe_1_5_4_N64, pe_1_5_4_N63, pe_1_5_4_N62, pe_1_5_4_N61, pe_1_5_4_N60,
         pe_1_5_4_N59, pe_1_5_5_n90, pe_1_5_5_n89, pe_1_5_5_n88, pe_1_5_5_n87,
         pe_1_5_5_n86, pe_1_5_5_n85, pe_1_5_5_n84, pe_1_5_5_n83, pe_1_5_5_n82,
         pe_1_5_5_n81, pe_1_5_5_n80, pe_1_5_5_n79, pe_1_5_5_n78, pe_1_5_5_n77,
         pe_1_5_5_n76, pe_1_5_5_n75, pe_1_5_5_n74, pe_1_5_5_n73, pe_1_5_5_n72,
         pe_1_5_5_n71, pe_1_5_5_n70, pe_1_5_5_n69, pe_1_5_5_n68, pe_1_5_5_n67,
         pe_1_5_5_n66, pe_1_5_5_n65, pe_1_5_5_n64, pe_1_5_5_n63, pe_1_5_5_n62,
         pe_1_5_5_n61, pe_1_5_5_n60, pe_1_5_5_n59, pe_1_5_5_n58, pe_1_5_5_n57,
         pe_1_5_5_n56, pe_1_5_5_n55, pe_1_5_5_n54, pe_1_5_5_n53, pe_1_5_5_n52,
         pe_1_5_5_n51, pe_1_5_5_n50, pe_1_5_5_n49, pe_1_5_5_n48, pe_1_5_5_n47,
         pe_1_5_5_n46, pe_1_5_5_n45, pe_1_5_5_n25, pe_1_5_5_n24, pe_1_5_5_n23,
         pe_1_5_5_n22, pe_1_5_5_n21, pe_1_5_5_n20, pe_1_5_5_n19, pe_1_5_5_n18,
         pe_1_5_5_n17, pe_1_5_5_n16, pe_1_5_5_n15, pe_1_5_5_n14, pe_1_5_5_n13,
         pe_1_5_5_n12, pe_1_5_5_n11, pe_1_5_5_n10, pe_1_5_5_n9, pe_1_5_5_n8,
         pe_1_5_5_n7, pe_1_5_5_n6, pe_1_5_5_n5, pe_1_5_5_n4, pe_1_5_5_n3,
         pe_1_5_5_n2, pe_1_5_5_n1, pe_1_5_5_n44, pe_1_5_5_n43, pe_1_5_5_n42,
         pe_1_5_5_n41, pe_1_5_5_n40, pe_1_5_5_n39, pe_1_5_5_n38, pe_1_5_5_n37,
         pe_1_5_5_n36, pe_1_5_5_n35, pe_1_5_5_n34, pe_1_5_5_n33, pe_1_5_5_n32,
         pe_1_5_5_n31, pe_1_5_5_n30, pe_1_5_5_n29, pe_1_5_5_n28, pe_1_5_5_n27,
         pe_1_5_5_n26, pe_1_5_5_net4042, pe_1_5_5_net4037, pe_1_5_5_net4032,
         pe_1_5_5_net4027, pe_1_5_5_net4022, pe_1_5_5_net4017,
         pe_1_5_5_net4012, pe_1_5_5_net4007, pe_1_5_5_net4002,
         pe_1_5_5_net3997, pe_1_5_5_net3992, pe_1_5_5_net3987,
         pe_1_5_5_net3981, pe_1_5_5_N90, pe_1_5_5_N85, pe_1_5_5_N84,
         pe_1_5_5_N83, pe_1_5_5_N82, pe_1_5_5_N81, pe_1_5_5_N80, pe_1_5_5_N79,
         pe_1_5_5_N77, pe_1_5_5_N76, pe_1_5_5_N75, pe_1_5_5_N74, pe_1_5_5_N73,
         pe_1_5_5_N72, pe_1_5_5_N71, pe_1_5_5_N70, pe_1_5_5_int_data_0_,
         pe_1_5_5_int_data_1_, pe_1_5_5_int_data_2_, pe_1_5_5_int_data_3_,
         pe_1_5_5_N64, pe_1_5_5_N63, pe_1_5_5_N62, pe_1_5_5_N61, pe_1_5_5_N60,
         pe_1_5_5_N59, pe_1_5_6_n90, pe_1_5_6_n89, pe_1_5_6_n88, pe_1_5_6_n87,
         pe_1_5_6_n86, pe_1_5_6_n85, pe_1_5_6_n84, pe_1_5_6_n83, pe_1_5_6_n82,
         pe_1_5_6_n81, pe_1_5_6_n80, pe_1_5_6_n79, pe_1_5_6_n78, pe_1_5_6_n77,
         pe_1_5_6_n76, pe_1_5_6_n75, pe_1_5_6_n74, pe_1_5_6_n73, pe_1_5_6_n72,
         pe_1_5_6_n71, pe_1_5_6_n70, pe_1_5_6_n69, pe_1_5_6_n68, pe_1_5_6_n67,
         pe_1_5_6_n66, pe_1_5_6_n65, pe_1_5_6_n64, pe_1_5_6_n63, pe_1_5_6_n62,
         pe_1_5_6_n61, pe_1_5_6_n60, pe_1_5_6_n59, pe_1_5_6_n58, pe_1_5_6_n57,
         pe_1_5_6_n56, pe_1_5_6_n55, pe_1_5_6_n54, pe_1_5_6_n53, pe_1_5_6_n52,
         pe_1_5_6_n51, pe_1_5_6_n50, pe_1_5_6_n49, pe_1_5_6_n48, pe_1_5_6_n47,
         pe_1_5_6_n46, pe_1_5_6_n45, pe_1_5_6_n25, pe_1_5_6_n24, pe_1_5_6_n23,
         pe_1_5_6_n22, pe_1_5_6_n21, pe_1_5_6_n20, pe_1_5_6_n19, pe_1_5_6_n18,
         pe_1_5_6_n17, pe_1_5_6_n16, pe_1_5_6_n15, pe_1_5_6_n14, pe_1_5_6_n13,
         pe_1_5_6_n12, pe_1_5_6_n11, pe_1_5_6_n10, pe_1_5_6_n9, pe_1_5_6_n8,
         pe_1_5_6_n7, pe_1_5_6_n6, pe_1_5_6_n5, pe_1_5_6_n4, pe_1_5_6_n3,
         pe_1_5_6_n2, pe_1_5_6_n1, pe_1_5_6_n44, pe_1_5_6_n43, pe_1_5_6_n42,
         pe_1_5_6_n41, pe_1_5_6_n40, pe_1_5_6_n39, pe_1_5_6_n38, pe_1_5_6_n37,
         pe_1_5_6_n36, pe_1_5_6_n35, pe_1_5_6_n34, pe_1_5_6_n33, pe_1_5_6_n32,
         pe_1_5_6_n31, pe_1_5_6_n30, pe_1_5_6_n29, pe_1_5_6_n28, pe_1_5_6_n27,
         pe_1_5_6_n26, pe_1_5_6_net3964, pe_1_5_6_net3959, pe_1_5_6_net3954,
         pe_1_5_6_net3949, pe_1_5_6_net3944, pe_1_5_6_net3939,
         pe_1_5_6_net3934, pe_1_5_6_net3929, pe_1_5_6_net3924,
         pe_1_5_6_net3919, pe_1_5_6_net3914, pe_1_5_6_net3909,
         pe_1_5_6_net3903, pe_1_5_6_N90, pe_1_5_6_N85, pe_1_5_6_N84,
         pe_1_5_6_N83, pe_1_5_6_N82, pe_1_5_6_N81, pe_1_5_6_N80, pe_1_5_6_N79,
         pe_1_5_6_N77, pe_1_5_6_N76, pe_1_5_6_N75, pe_1_5_6_N74, pe_1_5_6_N73,
         pe_1_5_6_N72, pe_1_5_6_N71, pe_1_5_6_N70, pe_1_5_6_int_data_0_,
         pe_1_5_6_int_data_1_, pe_1_5_6_int_data_2_, pe_1_5_6_int_data_3_,
         pe_1_5_6_N64, pe_1_5_6_N63, pe_1_5_6_N62, pe_1_5_6_N61, pe_1_5_6_N60,
         pe_1_5_6_N59, pe_1_5_7_n90, pe_1_5_7_n89, pe_1_5_7_n88, pe_1_5_7_n87,
         pe_1_5_7_n86, pe_1_5_7_n85, pe_1_5_7_n84, pe_1_5_7_n83, pe_1_5_7_n82,
         pe_1_5_7_n81, pe_1_5_7_n80, pe_1_5_7_n79, pe_1_5_7_n78, pe_1_5_7_n77,
         pe_1_5_7_n76, pe_1_5_7_n75, pe_1_5_7_n74, pe_1_5_7_n73, pe_1_5_7_n72,
         pe_1_5_7_n71, pe_1_5_7_n70, pe_1_5_7_n69, pe_1_5_7_n68, pe_1_5_7_n67,
         pe_1_5_7_n66, pe_1_5_7_n65, pe_1_5_7_n64, pe_1_5_7_n63, pe_1_5_7_n62,
         pe_1_5_7_n61, pe_1_5_7_n60, pe_1_5_7_n59, pe_1_5_7_n58, pe_1_5_7_n57,
         pe_1_5_7_n56, pe_1_5_7_n55, pe_1_5_7_n54, pe_1_5_7_n53, pe_1_5_7_n52,
         pe_1_5_7_n51, pe_1_5_7_n50, pe_1_5_7_n49, pe_1_5_7_n48, pe_1_5_7_n47,
         pe_1_5_7_n46, pe_1_5_7_n45, pe_1_5_7_n25, pe_1_5_7_n24, pe_1_5_7_n23,
         pe_1_5_7_n22, pe_1_5_7_n21, pe_1_5_7_n20, pe_1_5_7_n19, pe_1_5_7_n18,
         pe_1_5_7_n17, pe_1_5_7_n16, pe_1_5_7_n15, pe_1_5_7_n14, pe_1_5_7_n13,
         pe_1_5_7_n12, pe_1_5_7_n11, pe_1_5_7_n10, pe_1_5_7_n9, pe_1_5_7_n8,
         pe_1_5_7_n7, pe_1_5_7_n6, pe_1_5_7_n5, pe_1_5_7_n4, pe_1_5_7_n3,
         pe_1_5_7_n2, pe_1_5_7_n1, pe_1_5_7_n44, pe_1_5_7_n43, pe_1_5_7_n42,
         pe_1_5_7_n41, pe_1_5_7_n40, pe_1_5_7_n39, pe_1_5_7_n38, pe_1_5_7_n37,
         pe_1_5_7_n36, pe_1_5_7_n35, pe_1_5_7_n34, pe_1_5_7_n33, pe_1_5_7_n32,
         pe_1_5_7_n31, pe_1_5_7_n30, pe_1_5_7_n29, pe_1_5_7_n28, pe_1_5_7_n27,
         pe_1_5_7_n26, pe_1_5_7_net3886, pe_1_5_7_net3881, pe_1_5_7_net3876,
         pe_1_5_7_net3871, pe_1_5_7_net3866, pe_1_5_7_net3861,
         pe_1_5_7_net3856, pe_1_5_7_net3851, pe_1_5_7_net3846,
         pe_1_5_7_net3841, pe_1_5_7_net3836, pe_1_5_7_net3831,
         pe_1_5_7_net3825, pe_1_5_7_N90, pe_1_5_7_N85, pe_1_5_7_N84,
         pe_1_5_7_N83, pe_1_5_7_N82, pe_1_5_7_N81, pe_1_5_7_N80, pe_1_5_7_N79,
         pe_1_5_7_N77, pe_1_5_7_N76, pe_1_5_7_N75, pe_1_5_7_N74, pe_1_5_7_N73,
         pe_1_5_7_N72, pe_1_5_7_N71, pe_1_5_7_N70, pe_1_5_7_int_data_0_,
         pe_1_5_7_int_data_1_, pe_1_5_7_int_data_2_, pe_1_5_7_int_data_3_,
         pe_1_5_7_N64, pe_1_5_7_N63, pe_1_5_7_N62, pe_1_5_7_N61, pe_1_5_7_N60,
         pe_1_5_7_N59, pe_1_6_0_n87, pe_1_6_0_n86, pe_1_6_0_n85, pe_1_6_0_n84,
         pe_1_6_0_n83, pe_1_6_0_n82, pe_1_6_0_n81, pe_1_6_0_n80, pe_1_6_0_n79,
         pe_1_6_0_n78, pe_1_6_0_n77, pe_1_6_0_n76, pe_1_6_0_n75, pe_1_6_0_n74,
         pe_1_6_0_n73, pe_1_6_0_n72, pe_1_6_0_n71, pe_1_6_0_n70, pe_1_6_0_n69,
         pe_1_6_0_n68, pe_1_6_0_n67, pe_1_6_0_n66, pe_1_6_0_n65, pe_1_6_0_n64,
         pe_1_6_0_n63, pe_1_6_0_n62, pe_1_6_0_n61, pe_1_6_0_n60, pe_1_6_0_n59,
         pe_1_6_0_n58, pe_1_6_0_n57, pe_1_6_0_n56, pe_1_6_0_n55, pe_1_6_0_n54,
         pe_1_6_0_n53, pe_1_6_0_n52, pe_1_6_0_n51, pe_1_6_0_n50, pe_1_6_0_n49,
         pe_1_6_0_n48, pe_1_6_0_n47, pe_1_6_0_n46, pe_1_6_0_n45, pe_1_6_0_n25,
         pe_1_6_0_n24, pe_1_6_0_n23, pe_1_6_0_n22, pe_1_6_0_n21, pe_1_6_0_n20,
         pe_1_6_0_n19, pe_1_6_0_n18, pe_1_6_0_n17, pe_1_6_0_n16, pe_1_6_0_n15,
         pe_1_6_0_n14, pe_1_6_0_n13, pe_1_6_0_n12, pe_1_6_0_n11, pe_1_6_0_n10,
         pe_1_6_0_n9, pe_1_6_0_n8, pe_1_6_0_n7, pe_1_6_0_n6, pe_1_6_0_n5,
         pe_1_6_0_n4, pe_1_6_0_n3, pe_1_6_0_n2, pe_1_6_0_n1, pe_1_6_0_n44,
         pe_1_6_0_n43, pe_1_6_0_n42, pe_1_6_0_n41, pe_1_6_0_n40, pe_1_6_0_n39,
         pe_1_6_0_n38, pe_1_6_0_n37, pe_1_6_0_n36, pe_1_6_0_n35, pe_1_6_0_n34,
         pe_1_6_0_n33, pe_1_6_0_n32, pe_1_6_0_n31, pe_1_6_0_n30, pe_1_6_0_n29,
         pe_1_6_0_n28, pe_1_6_0_n27, pe_1_6_0_n26, pe_1_6_0_net3808,
         pe_1_6_0_net3803, pe_1_6_0_net3798, pe_1_6_0_net3793,
         pe_1_6_0_net3788, pe_1_6_0_net3783, pe_1_6_0_net3778,
         pe_1_6_0_net3773, pe_1_6_0_net3768, pe_1_6_0_net3763,
         pe_1_6_0_net3758, pe_1_6_0_net3753, pe_1_6_0_net3747, pe_1_6_0_N90,
         pe_1_6_0_N85, pe_1_6_0_N84, pe_1_6_0_N83, pe_1_6_0_N82, pe_1_6_0_N81,
         pe_1_6_0_N80, pe_1_6_0_N79, pe_1_6_0_N77, pe_1_6_0_N76, pe_1_6_0_N75,
         pe_1_6_0_N74, pe_1_6_0_N73, pe_1_6_0_N72, pe_1_6_0_N71, pe_1_6_0_N70,
         pe_1_6_0_int_data_0_, pe_1_6_0_int_data_1_, pe_1_6_0_int_data_2_,
         pe_1_6_0_int_data_3_, pe_1_6_0_N64, pe_1_6_0_N63, pe_1_6_0_N62,
         pe_1_6_0_N61, pe_1_6_0_N60, pe_1_6_0_N59, pe_1_6_0_o_data_h_0_,
         pe_1_6_0_o_data_h_1_, pe_1_6_0_o_data_h_2_, pe_1_6_0_o_data_h_3_,
         pe_1_6_1_n86, pe_1_6_1_n85, pe_1_6_1_n84, pe_1_6_1_n83, pe_1_6_1_n82,
         pe_1_6_1_n81, pe_1_6_1_n80, pe_1_6_1_n79, pe_1_6_1_n78, pe_1_6_1_n77,
         pe_1_6_1_n76, pe_1_6_1_n75, pe_1_6_1_n74, pe_1_6_1_n73, pe_1_6_1_n72,
         pe_1_6_1_n71, pe_1_6_1_n70, pe_1_6_1_n69, pe_1_6_1_n68, pe_1_6_1_n67,
         pe_1_6_1_n66, pe_1_6_1_n65, pe_1_6_1_n64, pe_1_6_1_n63, pe_1_6_1_n62,
         pe_1_6_1_n61, pe_1_6_1_n60, pe_1_6_1_n59, pe_1_6_1_n58, pe_1_6_1_n57,
         pe_1_6_1_n56, pe_1_6_1_n55, pe_1_6_1_n54, pe_1_6_1_n53, pe_1_6_1_n52,
         pe_1_6_1_n51, pe_1_6_1_n50, pe_1_6_1_n49, pe_1_6_1_n48, pe_1_6_1_n47,
         pe_1_6_1_n46, pe_1_6_1_n45, pe_1_6_1_n25, pe_1_6_1_n24, pe_1_6_1_n23,
         pe_1_6_1_n22, pe_1_6_1_n21, pe_1_6_1_n20, pe_1_6_1_n19, pe_1_6_1_n18,
         pe_1_6_1_n17, pe_1_6_1_n16, pe_1_6_1_n15, pe_1_6_1_n14, pe_1_6_1_n13,
         pe_1_6_1_n12, pe_1_6_1_n11, pe_1_6_1_n10, pe_1_6_1_n9, pe_1_6_1_n8,
         pe_1_6_1_n7, pe_1_6_1_n6, pe_1_6_1_n5, pe_1_6_1_n4, pe_1_6_1_n3,
         pe_1_6_1_n2, pe_1_6_1_n1, pe_1_6_1_n44, pe_1_6_1_n43, pe_1_6_1_n42,
         pe_1_6_1_n41, pe_1_6_1_n40, pe_1_6_1_n39, pe_1_6_1_n38, pe_1_6_1_n37,
         pe_1_6_1_n36, pe_1_6_1_n35, pe_1_6_1_n34, pe_1_6_1_n33, pe_1_6_1_n32,
         pe_1_6_1_n31, pe_1_6_1_n30, pe_1_6_1_n29, pe_1_6_1_n28, pe_1_6_1_n27,
         pe_1_6_1_n26, pe_1_6_1_net3730, pe_1_6_1_net3725, pe_1_6_1_net3720,
         pe_1_6_1_net3715, pe_1_6_1_net3710, pe_1_6_1_net3705,
         pe_1_6_1_net3700, pe_1_6_1_net3695, pe_1_6_1_net3690,
         pe_1_6_1_net3685, pe_1_6_1_net3680, pe_1_6_1_net3675,
         pe_1_6_1_net3669, pe_1_6_1_N90, pe_1_6_1_N85, pe_1_6_1_N84,
         pe_1_6_1_N83, pe_1_6_1_N82, pe_1_6_1_N81, pe_1_6_1_N80, pe_1_6_1_N79,
         pe_1_6_1_N77, pe_1_6_1_N76, pe_1_6_1_N75, pe_1_6_1_N74, pe_1_6_1_N73,
         pe_1_6_1_N72, pe_1_6_1_N71, pe_1_6_1_N70, pe_1_6_1_int_data_0_,
         pe_1_6_1_int_data_1_, pe_1_6_1_int_data_2_, pe_1_6_1_int_data_3_,
         pe_1_6_1_N64, pe_1_6_1_N63, pe_1_6_1_N62, pe_1_6_1_N61, pe_1_6_1_N60,
         pe_1_6_1_N59, pe_1_6_2_n87, pe_1_6_2_n86, pe_1_6_2_n85, pe_1_6_2_n84,
         pe_1_6_2_n83, pe_1_6_2_n82, pe_1_6_2_n81, pe_1_6_2_n80, pe_1_6_2_n79,
         pe_1_6_2_n78, pe_1_6_2_n77, pe_1_6_2_n76, pe_1_6_2_n75, pe_1_6_2_n74,
         pe_1_6_2_n73, pe_1_6_2_n72, pe_1_6_2_n71, pe_1_6_2_n70, pe_1_6_2_n69,
         pe_1_6_2_n68, pe_1_6_2_n67, pe_1_6_2_n66, pe_1_6_2_n65, pe_1_6_2_n64,
         pe_1_6_2_n63, pe_1_6_2_n62, pe_1_6_2_n61, pe_1_6_2_n60, pe_1_6_2_n59,
         pe_1_6_2_n58, pe_1_6_2_n57, pe_1_6_2_n56, pe_1_6_2_n55, pe_1_6_2_n54,
         pe_1_6_2_n53, pe_1_6_2_n52, pe_1_6_2_n51, pe_1_6_2_n50, pe_1_6_2_n49,
         pe_1_6_2_n48, pe_1_6_2_n47, pe_1_6_2_n46, pe_1_6_2_n45, pe_1_6_2_n25,
         pe_1_6_2_n24, pe_1_6_2_n23, pe_1_6_2_n22, pe_1_6_2_n21, pe_1_6_2_n20,
         pe_1_6_2_n19, pe_1_6_2_n18, pe_1_6_2_n17, pe_1_6_2_n16, pe_1_6_2_n15,
         pe_1_6_2_n14, pe_1_6_2_n13, pe_1_6_2_n12, pe_1_6_2_n11, pe_1_6_2_n10,
         pe_1_6_2_n9, pe_1_6_2_n8, pe_1_6_2_n7, pe_1_6_2_n6, pe_1_6_2_n5,
         pe_1_6_2_n4, pe_1_6_2_n3, pe_1_6_2_n2, pe_1_6_2_n1, pe_1_6_2_n44,
         pe_1_6_2_n43, pe_1_6_2_n42, pe_1_6_2_n41, pe_1_6_2_n40, pe_1_6_2_n39,
         pe_1_6_2_n38, pe_1_6_2_n37, pe_1_6_2_n36, pe_1_6_2_n35, pe_1_6_2_n34,
         pe_1_6_2_n33, pe_1_6_2_n32, pe_1_6_2_n31, pe_1_6_2_n30, pe_1_6_2_n29,
         pe_1_6_2_n28, pe_1_6_2_n27, pe_1_6_2_n26, pe_1_6_2_net3652,
         pe_1_6_2_net3647, pe_1_6_2_net3642, pe_1_6_2_net3637,
         pe_1_6_2_net3632, pe_1_6_2_net3627, pe_1_6_2_net3622,
         pe_1_6_2_net3617, pe_1_6_2_net3612, pe_1_6_2_net3607,
         pe_1_6_2_net3602, pe_1_6_2_net3597, pe_1_6_2_net3591, pe_1_6_2_N90,
         pe_1_6_2_N85, pe_1_6_2_N84, pe_1_6_2_N83, pe_1_6_2_N82, pe_1_6_2_N81,
         pe_1_6_2_N80, pe_1_6_2_N79, pe_1_6_2_N77, pe_1_6_2_N76, pe_1_6_2_N75,
         pe_1_6_2_N74, pe_1_6_2_N73, pe_1_6_2_N72, pe_1_6_2_N71, pe_1_6_2_N70,
         pe_1_6_2_int_data_0_, pe_1_6_2_int_data_1_, pe_1_6_2_int_data_2_,
         pe_1_6_2_int_data_3_, pe_1_6_2_N64, pe_1_6_2_N63, pe_1_6_2_N62,
         pe_1_6_2_N61, pe_1_6_2_N60, pe_1_6_2_N59, pe_1_6_3_n88, pe_1_6_3_n87,
         pe_1_6_3_n86, pe_1_6_3_n85, pe_1_6_3_n84, pe_1_6_3_n83, pe_1_6_3_n82,
         pe_1_6_3_n81, pe_1_6_3_n80, pe_1_6_3_n79, pe_1_6_3_n78, pe_1_6_3_n77,
         pe_1_6_3_n76, pe_1_6_3_n75, pe_1_6_3_n74, pe_1_6_3_n73, pe_1_6_3_n72,
         pe_1_6_3_n71, pe_1_6_3_n70, pe_1_6_3_n69, pe_1_6_3_n68, pe_1_6_3_n67,
         pe_1_6_3_n66, pe_1_6_3_n65, pe_1_6_3_n64, pe_1_6_3_n63, pe_1_6_3_n62,
         pe_1_6_3_n61, pe_1_6_3_n60, pe_1_6_3_n59, pe_1_6_3_n58, pe_1_6_3_n57,
         pe_1_6_3_n56, pe_1_6_3_n55, pe_1_6_3_n54, pe_1_6_3_n53, pe_1_6_3_n52,
         pe_1_6_3_n51, pe_1_6_3_n50, pe_1_6_3_n49, pe_1_6_3_n48, pe_1_6_3_n47,
         pe_1_6_3_n46, pe_1_6_3_n45, pe_1_6_3_n25, pe_1_6_3_n24, pe_1_6_3_n23,
         pe_1_6_3_n22, pe_1_6_3_n21, pe_1_6_3_n20, pe_1_6_3_n19, pe_1_6_3_n18,
         pe_1_6_3_n17, pe_1_6_3_n16, pe_1_6_3_n15, pe_1_6_3_n14, pe_1_6_3_n13,
         pe_1_6_3_n12, pe_1_6_3_n11, pe_1_6_3_n10, pe_1_6_3_n9, pe_1_6_3_n8,
         pe_1_6_3_n7, pe_1_6_3_n6, pe_1_6_3_n5, pe_1_6_3_n4, pe_1_6_3_n3,
         pe_1_6_3_n2, pe_1_6_3_n1, pe_1_6_3_n44, pe_1_6_3_n43, pe_1_6_3_n42,
         pe_1_6_3_n41, pe_1_6_3_n40, pe_1_6_3_n39, pe_1_6_3_n38, pe_1_6_3_n37,
         pe_1_6_3_n36, pe_1_6_3_n35, pe_1_6_3_n34, pe_1_6_3_n33, pe_1_6_3_n32,
         pe_1_6_3_n31, pe_1_6_3_n30, pe_1_6_3_n29, pe_1_6_3_n28, pe_1_6_3_n27,
         pe_1_6_3_n26, pe_1_6_3_net3574, pe_1_6_3_net3569, pe_1_6_3_net3564,
         pe_1_6_3_net3559, pe_1_6_3_net3554, pe_1_6_3_net3549,
         pe_1_6_3_net3544, pe_1_6_3_net3539, pe_1_6_3_net3534,
         pe_1_6_3_net3529, pe_1_6_3_net3524, pe_1_6_3_net3519,
         pe_1_6_3_net3513, pe_1_6_3_N90, pe_1_6_3_N85, pe_1_6_3_N84,
         pe_1_6_3_N83, pe_1_6_3_N82, pe_1_6_3_N81, pe_1_6_3_N80, pe_1_6_3_N79,
         pe_1_6_3_N77, pe_1_6_3_N76, pe_1_6_3_N75, pe_1_6_3_N74, pe_1_6_3_N73,
         pe_1_6_3_N72, pe_1_6_3_N71, pe_1_6_3_N70, pe_1_6_3_int_data_0_,
         pe_1_6_3_int_data_1_, pe_1_6_3_int_data_2_, pe_1_6_3_int_data_3_,
         pe_1_6_3_N64, pe_1_6_3_N63, pe_1_6_3_N62, pe_1_6_3_N61, pe_1_6_3_N60,
         pe_1_6_3_N59, pe_1_6_4_n90, pe_1_6_4_n89, pe_1_6_4_n88, pe_1_6_4_n87,
         pe_1_6_4_n86, pe_1_6_4_n85, pe_1_6_4_n84, pe_1_6_4_n83, pe_1_6_4_n82,
         pe_1_6_4_n81, pe_1_6_4_n80, pe_1_6_4_n79, pe_1_6_4_n78, pe_1_6_4_n77,
         pe_1_6_4_n76, pe_1_6_4_n75, pe_1_6_4_n74, pe_1_6_4_n73, pe_1_6_4_n72,
         pe_1_6_4_n71, pe_1_6_4_n70, pe_1_6_4_n69, pe_1_6_4_n68, pe_1_6_4_n67,
         pe_1_6_4_n66, pe_1_6_4_n65, pe_1_6_4_n64, pe_1_6_4_n63, pe_1_6_4_n62,
         pe_1_6_4_n61, pe_1_6_4_n60, pe_1_6_4_n59, pe_1_6_4_n58, pe_1_6_4_n57,
         pe_1_6_4_n56, pe_1_6_4_n55, pe_1_6_4_n54, pe_1_6_4_n53, pe_1_6_4_n52,
         pe_1_6_4_n51, pe_1_6_4_n50, pe_1_6_4_n49, pe_1_6_4_n48, pe_1_6_4_n47,
         pe_1_6_4_n46, pe_1_6_4_n45, pe_1_6_4_n25, pe_1_6_4_n24, pe_1_6_4_n23,
         pe_1_6_4_n22, pe_1_6_4_n21, pe_1_6_4_n20, pe_1_6_4_n19, pe_1_6_4_n18,
         pe_1_6_4_n17, pe_1_6_4_n16, pe_1_6_4_n15, pe_1_6_4_n14, pe_1_6_4_n13,
         pe_1_6_4_n12, pe_1_6_4_n11, pe_1_6_4_n10, pe_1_6_4_n9, pe_1_6_4_n8,
         pe_1_6_4_n7, pe_1_6_4_n6, pe_1_6_4_n5, pe_1_6_4_n4, pe_1_6_4_n3,
         pe_1_6_4_n2, pe_1_6_4_n1, pe_1_6_4_n44, pe_1_6_4_n43, pe_1_6_4_n42,
         pe_1_6_4_n41, pe_1_6_4_n40, pe_1_6_4_n39, pe_1_6_4_n38, pe_1_6_4_n37,
         pe_1_6_4_n36, pe_1_6_4_n35, pe_1_6_4_n34, pe_1_6_4_n33, pe_1_6_4_n32,
         pe_1_6_4_n31, pe_1_6_4_n30, pe_1_6_4_n29, pe_1_6_4_n28, pe_1_6_4_n27,
         pe_1_6_4_n26, pe_1_6_4_net3496, pe_1_6_4_net3491, pe_1_6_4_net3486,
         pe_1_6_4_net3481, pe_1_6_4_net3476, pe_1_6_4_net3471,
         pe_1_6_4_net3466, pe_1_6_4_net3461, pe_1_6_4_net3456,
         pe_1_6_4_net3451, pe_1_6_4_net3446, pe_1_6_4_net3441,
         pe_1_6_4_net3435, pe_1_6_4_N90, pe_1_6_4_N85, pe_1_6_4_N84,
         pe_1_6_4_N83, pe_1_6_4_N82, pe_1_6_4_N81, pe_1_6_4_N80, pe_1_6_4_N79,
         pe_1_6_4_N77, pe_1_6_4_N76, pe_1_6_4_N75, pe_1_6_4_N74, pe_1_6_4_N73,
         pe_1_6_4_N72, pe_1_6_4_N71, pe_1_6_4_N70, pe_1_6_4_int_data_0_,
         pe_1_6_4_int_data_1_, pe_1_6_4_int_data_2_, pe_1_6_4_int_data_3_,
         pe_1_6_4_N64, pe_1_6_4_N63, pe_1_6_4_N62, pe_1_6_4_N61, pe_1_6_4_N60,
         pe_1_6_4_N59, pe_1_6_5_n90, pe_1_6_5_n89, pe_1_6_5_n88, pe_1_6_5_n87,
         pe_1_6_5_n86, pe_1_6_5_n85, pe_1_6_5_n84, pe_1_6_5_n83, pe_1_6_5_n82,
         pe_1_6_5_n81, pe_1_6_5_n80, pe_1_6_5_n79, pe_1_6_5_n78, pe_1_6_5_n77,
         pe_1_6_5_n76, pe_1_6_5_n75, pe_1_6_5_n74, pe_1_6_5_n73, pe_1_6_5_n72,
         pe_1_6_5_n71, pe_1_6_5_n70, pe_1_6_5_n69, pe_1_6_5_n68, pe_1_6_5_n67,
         pe_1_6_5_n66, pe_1_6_5_n65, pe_1_6_5_n64, pe_1_6_5_n63, pe_1_6_5_n62,
         pe_1_6_5_n61, pe_1_6_5_n60, pe_1_6_5_n59, pe_1_6_5_n58, pe_1_6_5_n57,
         pe_1_6_5_n56, pe_1_6_5_n55, pe_1_6_5_n54, pe_1_6_5_n53, pe_1_6_5_n52,
         pe_1_6_5_n51, pe_1_6_5_n50, pe_1_6_5_n49, pe_1_6_5_n48, pe_1_6_5_n47,
         pe_1_6_5_n46, pe_1_6_5_n45, pe_1_6_5_n25, pe_1_6_5_n24, pe_1_6_5_n23,
         pe_1_6_5_n22, pe_1_6_5_n21, pe_1_6_5_n20, pe_1_6_5_n19, pe_1_6_5_n18,
         pe_1_6_5_n17, pe_1_6_5_n16, pe_1_6_5_n15, pe_1_6_5_n14, pe_1_6_5_n13,
         pe_1_6_5_n12, pe_1_6_5_n11, pe_1_6_5_n10, pe_1_6_5_n9, pe_1_6_5_n8,
         pe_1_6_5_n7, pe_1_6_5_n6, pe_1_6_5_n5, pe_1_6_5_n4, pe_1_6_5_n3,
         pe_1_6_5_n2, pe_1_6_5_n1, pe_1_6_5_n44, pe_1_6_5_n43, pe_1_6_5_n42,
         pe_1_6_5_n41, pe_1_6_5_n40, pe_1_6_5_n39, pe_1_6_5_n38, pe_1_6_5_n37,
         pe_1_6_5_n36, pe_1_6_5_n35, pe_1_6_5_n34, pe_1_6_5_n33, pe_1_6_5_n32,
         pe_1_6_5_n31, pe_1_6_5_n30, pe_1_6_5_n29, pe_1_6_5_n28, pe_1_6_5_n27,
         pe_1_6_5_n26, pe_1_6_5_net3418, pe_1_6_5_net3413, pe_1_6_5_net3408,
         pe_1_6_5_net3403, pe_1_6_5_net3398, pe_1_6_5_net3393,
         pe_1_6_5_net3388, pe_1_6_5_net3383, pe_1_6_5_net3378,
         pe_1_6_5_net3373, pe_1_6_5_net3368, pe_1_6_5_net3363,
         pe_1_6_5_net3357, pe_1_6_5_N90, pe_1_6_5_N85, pe_1_6_5_N84,
         pe_1_6_5_N83, pe_1_6_5_N82, pe_1_6_5_N81, pe_1_6_5_N80, pe_1_6_5_N79,
         pe_1_6_5_N77, pe_1_6_5_N76, pe_1_6_5_N75, pe_1_6_5_N74, pe_1_6_5_N73,
         pe_1_6_5_N72, pe_1_6_5_N71, pe_1_6_5_N70, pe_1_6_5_int_data_0_,
         pe_1_6_5_int_data_1_, pe_1_6_5_int_data_2_, pe_1_6_5_int_data_3_,
         pe_1_6_5_N64, pe_1_6_5_N63, pe_1_6_5_N62, pe_1_6_5_N61, pe_1_6_5_N60,
         pe_1_6_5_N59, pe_1_6_6_n90, pe_1_6_6_n89, pe_1_6_6_n88, pe_1_6_6_n87,
         pe_1_6_6_n86, pe_1_6_6_n85, pe_1_6_6_n84, pe_1_6_6_n83, pe_1_6_6_n82,
         pe_1_6_6_n81, pe_1_6_6_n80, pe_1_6_6_n79, pe_1_6_6_n78, pe_1_6_6_n77,
         pe_1_6_6_n76, pe_1_6_6_n75, pe_1_6_6_n74, pe_1_6_6_n73, pe_1_6_6_n72,
         pe_1_6_6_n71, pe_1_6_6_n70, pe_1_6_6_n69, pe_1_6_6_n68, pe_1_6_6_n67,
         pe_1_6_6_n66, pe_1_6_6_n65, pe_1_6_6_n64, pe_1_6_6_n63, pe_1_6_6_n62,
         pe_1_6_6_n61, pe_1_6_6_n60, pe_1_6_6_n59, pe_1_6_6_n58, pe_1_6_6_n57,
         pe_1_6_6_n56, pe_1_6_6_n55, pe_1_6_6_n54, pe_1_6_6_n53, pe_1_6_6_n52,
         pe_1_6_6_n51, pe_1_6_6_n50, pe_1_6_6_n49, pe_1_6_6_n48, pe_1_6_6_n47,
         pe_1_6_6_n46, pe_1_6_6_n45, pe_1_6_6_n25, pe_1_6_6_n24, pe_1_6_6_n23,
         pe_1_6_6_n22, pe_1_6_6_n21, pe_1_6_6_n20, pe_1_6_6_n19, pe_1_6_6_n18,
         pe_1_6_6_n17, pe_1_6_6_n16, pe_1_6_6_n15, pe_1_6_6_n14, pe_1_6_6_n13,
         pe_1_6_6_n12, pe_1_6_6_n11, pe_1_6_6_n10, pe_1_6_6_n9, pe_1_6_6_n8,
         pe_1_6_6_n7, pe_1_6_6_n6, pe_1_6_6_n5, pe_1_6_6_n4, pe_1_6_6_n3,
         pe_1_6_6_n2, pe_1_6_6_n1, pe_1_6_6_n44, pe_1_6_6_n43, pe_1_6_6_n42,
         pe_1_6_6_n41, pe_1_6_6_n40, pe_1_6_6_n39, pe_1_6_6_n38, pe_1_6_6_n37,
         pe_1_6_6_n36, pe_1_6_6_n35, pe_1_6_6_n34, pe_1_6_6_n33, pe_1_6_6_n32,
         pe_1_6_6_n31, pe_1_6_6_n30, pe_1_6_6_n29, pe_1_6_6_n28, pe_1_6_6_n27,
         pe_1_6_6_n26, pe_1_6_6_net3340, pe_1_6_6_net3335, pe_1_6_6_net3330,
         pe_1_6_6_net3325, pe_1_6_6_net3320, pe_1_6_6_net3315,
         pe_1_6_6_net3310, pe_1_6_6_net3305, pe_1_6_6_net3300,
         pe_1_6_6_net3295, pe_1_6_6_net3290, pe_1_6_6_net3285,
         pe_1_6_6_net3279, pe_1_6_6_N90, pe_1_6_6_N85, pe_1_6_6_N84,
         pe_1_6_6_N83, pe_1_6_6_N82, pe_1_6_6_N81, pe_1_6_6_N80, pe_1_6_6_N79,
         pe_1_6_6_N77, pe_1_6_6_N76, pe_1_6_6_N75, pe_1_6_6_N74, pe_1_6_6_N73,
         pe_1_6_6_N72, pe_1_6_6_N71, pe_1_6_6_N70, pe_1_6_6_int_data_0_,
         pe_1_6_6_int_data_1_, pe_1_6_6_int_data_2_, pe_1_6_6_int_data_3_,
         pe_1_6_6_N64, pe_1_6_6_N63, pe_1_6_6_N62, pe_1_6_6_N61, pe_1_6_6_N60,
         pe_1_6_6_N59, pe_1_6_7_n90, pe_1_6_7_n89, pe_1_6_7_n88, pe_1_6_7_n87,
         pe_1_6_7_n86, pe_1_6_7_n85, pe_1_6_7_n84, pe_1_6_7_n83, pe_1_6_7_n82,
         pe_1_6_7_n81, pe_1_6_7_n80, pe_1_6_7_n79, pe_1_6_7_n78, pe_1_6_7_n77,
         pe_1_6_7_n76, pe_1_6_7_n75, pe_1_6_7_n74, pe_1_6_7_n73, pe_1_6_7_n72,
         pe_1_6_7_n71, pe_1_6_7_n70, pe_1_6_7_n69, pe_1_6_7_n68, pe_1_6_7_n67,
         pe_1_6_7_n66, pe_1_6_7_n65, pe_1_6_7_n64, pe_1_6_7_n63, pe_1_6_7_n62,
         pe_1_6_7_n61, pe_1_6_7_n60, pe_1_6_7_n59, pe_1_6_7_n58, pe_1_6_7_n57,
         pe_1_6_7_n56, pe_1_6_7_n55, pe_1_6_7_n54, pe_1_6_7_n53, pe_1_6_7_n52,
         pe_1_6_7_n51, pe_1_6_7_n50, pe_1_6_7_n49, pe_1_6_7_n48, pe_1_6_7_n47,
         pe_1_6_7_n46, pe_1_6_7_n45, pe_1_6_7_n25, pe_1_6_7_n24, pe_1_6_7_n23,
         pe_1_6_7_n22, pe_1_6_7_n21, pe_1_6_7_n20, pe_1_6_7_n19, pe_1_6_7_n18,
         pe_1_6_7_n17, pe_1_6_7_n16, pe_1_6_7_n15, pe_1_6_7_n14, pe_1_6_7_n13,
         pe_1_6_7_n12, pe_1_6_7_n11, pe_1_6_7_n10, pe_1_6_7_n9, pe_1_6_7_n8,
         pe_1_6_7_n7, pe_1_6_7_n6, pe_1_6_7_n5, pe_1_6_7_n4, pe_1_6_7_n3,
         pe_1_6_7_n2, pe_1_6_7_n1, pe_1_6_7_n44, pe_1_6_7_n43, pe_1_6_7_n42,
         pe_1_6_7_n41, pe_1_6_7_n40, pe_1_6_7_n39, pe_1_6_7_n38, pe_1_6_7_n37,
         pe_1_6_7_n36, pe_1_6_7_n35, pe_1_6_7_n34, pe_1_6_7_n33, pe_1_6_7_n32,
         pe_1_6_7_n31, pe_1_6_7_n30, pe_1_6_7_n29, pe_1_6_7_n28, pe_1_6_7_n27,
         pe_1_6_7_n26, pe_1_6_7_net3262, pe_1_6_7_net3257, pe_1_6_7_net3252,
         pe_1_6_7_net3247, pe_1_6_7_net3242, pe_1_6_7_net3237,
         pe_1_6_7_net3232, pe_1_6_7_net3227, pe_1_6_7_net3222,
         pe_1_6_7_net3217, pe_1_6_7_net3212, pe_1_6_7_net3207,
         pe_1_6_7_net3201, pe_1_6_7_N90, pe_1_6_7_N85, pe_1_6_7_N84,
         pe_1_6_7_N83, pe_1_6_7_N82, pe_1_6_7_N81, pe_1_6_7_N80, pe_1_6_7_N79,
         pe_1_6_7_N77, pe_1_6_7_N76, pe_1_6_7_N75, pe_1_6_7_N74, pe_1_6_7_N73,
         pe_1_6_7_N72, pe_1_6_7_N71, pe_1_6_7_N70, pe_1_6_7_int_data_0_,
         pe_1_6_7_int_data_1_, pe_1_6_7_int_data_2_, pe_1_6_7_int_data_3_,
         pe_1_6_7_N64, pe_1_6_7_N63, pe_1_6_7_N62, pe_1_6_7_N61, pe_1_6_7_N60,
         pe_1_6_7_N59, pe_1_7_0_n90, pe_1_7_0_n89, pe_1_7_0_n88, pe_1_7_0_n87,
         pe_1_7_0_n86, pe_1_7_0_n85, pe_1_7_0_n84, pe_1_7_0_n83, pe_1_7_0_n82,
         pe_1_7_0_n81, pe_1_7_0_n80, pe_1_7_0_n79, pe_1_7_0_n78, pe_1_7_0_n77,
         pe_1_7_0_n76, pe_1_7_0_n75, pe_1_7_0_n74, pe_1_7_0_n73, pe_1_7_0_n72,
         pe_1_7_0_n71, pe_1_7_0_n70, pe_1_7_0_n69, pe_1_7_0_n68, pe_1_7_0_n67,
         pe_1_7_0_n66, pe_1_7_0_n65, pe_1_7_0_n64, pe_1_7_0_n63, pe_1_7_0_n62,
         pe_1_7_0_n61, pe_1_7_0_n60, pe_1_7_0_n59, pe_1_7_0_n58, pe_1_7_0_n57,
         pe_1_7_0_n56, pe_1_7_0_n55, pe_1_7_0_n54, pe_1_7_0_n53, pe_1_7_0_n52,
         pe_1_7_0_n51, pe_1_7_0_n50, pe_1_7_0_n49, pe_1_7_0_n48, pe_1_7_0_n47,
         pe_1_7_0_n46, pe_1_7_0_n45, pe_1_7_0_n25, pe_1_7_0_n24, pe_1_7_0_n23,
         pe_1_7_0_n22, pe_1_7_0_n21, pe_1_7_0_n20, pe_1_7_0_n19, pe_1_7_0_n18,
         pe_1_7_0_n17, pe_1_7_0_n16, pe_1_7_0_n15, pe_1_7_0_n14, pe_1_7_0_n13,
         pe_1_7_0_n12, pe_1_7_0_n11, pe_1_7_0_n10, pe_1_7_0_n9, pe_1_7_0_n8,
         pe_1_7_0_n7, pe_1_7_0_n6, pe_1_7_0_n5, pe_1_7_0_n4, pe_1_7_0_n3,
         pe_1_7_0_n2, pe_1_7_0_n1, pe_1_7_0_n44, pe_1_7_0_n43, pe_1_7_0_n42,
         pe_1_7_0_n41, pe_1_7_0_n40, pe_1_7_0_n39, pe_1_7_0_n38, pe_1_7_0_n37,
         pe_1_7_0_n36, pe_1_7_0_n35, pe_1_7_0_n34, pe_1_7_0_n33, pe_1_7_0_n32,
         pe_1_7_0_n31, pe_1_7_0_n30, pe_1_7_0_n29, pe_1_7_0_n28, pe_1_7_0_n27,
         pe_1_7_0_n26, pe_1_7_0_net3184, pe_1_7_0_net3179, pe_1_7_0_net3174,
         pe_1_7_0_net3169, pe_1_7_0_net3164, pe_1_7_0_net3159,
         pe_1_7_0_net3154, pe_1_7_0_net3149, pe_1_7_0_net3144,
         pe_1_7_0_net3139, pe_1_7_0_net3134, pe_1_7_0_net3129,
         pe_1_7_0_net3123, pe_1_7_0_N90, pe_1_7_0_N85, pe_1_7_0_N84,
         pe_1_7_0_N83, pe_1_7_0_N82, pe_1_7_0_N81, pe_1_7_0_N80, pe_1_7_0_N79,
         pe_1_7_0_N77, pe_1_7_0_N76, pe_1_7_0_N75, pe_1_7_0_N74, pe_1_7_0_N73,
         pe_1_7_0_N72, pe_1_7_0_N71, pe_1_7_0_N70, pe_1_7_0_int_data_0_,
         pe_1_7_0_int_data_1_, pe_1_7_0_int_data_2_, pe_1_7_0_int_data_3_,
         pe_1_7_0_N64, pe_1_7_0_N63, pe_1_7_0_N62, pe_1_7_0_N61, pe_1_7_0_N60,
         pe_1_7_0_N59, pe_1_7_0_o_data_h_0_, pe_1_7_0_o_data_h_1_,
         pe_1_7_0_o_data_h_2_, pe_1_7_0_o_data_h_3_, pe_1_7_1_n90,
         pe_1_7_1_n89, pe_1_7_1_n88, pe_1_7_1_n87, pe_1_7_1_n86, pe_1_7_1_n85,
         pe_1_7_1_n84, pe_1_7_1_n83, pe_1_7_1_n82, pe_1_7_1_n81, pe_1_7_1_n80,
         pe_1_7_1_n79, pe_1_7_1_n78, pe_1_7_1_n77, pe_1_7_1_n76, pe_1_7_1_n75,
         pe_1_7_1_n74, pe_1_7_1_n73, pe_1_7_1_n72, pe_1_7_1_n71, pe_1_7_1_n70,
         pe_1_7_1_n69, pe_1_7_1_n68, pe_1_7_1_n67, pe_1_7_1_n66, pe_1_7_1_n65,
         pe_1_7_1_n64, pe_1_7_1_n63, pe_1_7_1_n62, pe_1_7_1_n61, pe_1_7_1_n60,
         pe_1_7_1_n59, pe_1_7_1_n58, pe_1_7_1_n57, pe_1_7_1_n56, pe_1_7_1_n55,
         pe_1_7_1_n54, pe_1_7_1_n53, pe_1_7_1_n52, pe_1_7_1_n51, pe_1_7_1_n50,
         pe_1_7_1_n49, pe_1_7_1_n48, pe_1_7_1_n47, pe_1_7_1_n46, pe_1_7_1_n45,
         pe_1_7_1_n25, pe_1_7_1_n24, pe_1_7_1_n23, pe_1_7_1_n22, pe_1_7_1_n21,
         pe_1_7_1_n20, pe_1_7_1_n19, pe_1_7_1_n18, pe_1_7_1_n17, pe_1_7_1_n16,
         pe_1_7_1_n15, pe_1_7_1_n14, pe_1_7_1_n13, pe_1_7_1_n12, pe_1_7_1_n11,
         pe_1_7_1_n10, pe_1_7_1_n9, pe_1_7_1_n8, pe_1_7_1_n7, pe_1_7_1_n6,
         pe_1_7_1_n5, pe_1_7_1_n4, pe_1_7_1_n3, pe_1_7_1_n2, pe_1_7_1_n1,
         pe_1_7_1_n44, pe_1_7_1_n43, pe_1_7_1_n42, pe_1_7_1_n41, pe_1_7_1_n40,
         pe_1_7_1_n39, pe_1_7_1_n38, pe_1_7_1_n37, pe_1_7_1_n36, pe_1_7_1_n35,
         pe_1_7_1_n34, pe_1_7_1_n33, pe_1_7_1_n32, pe_1_7_1_n31, pe_1_7_1_n30,
         pe_1_7_1_n29, pe_1_7_1_n28, pe_1_7_1_n27, pe_1_7_1_n26,
         pe_1_7_1_net3106, pe_1_7_1_net3101, pe_1_7_1_net3096,
         pe_1_7_1_net3091, pe_1_7_1_net3086, pe_1_7_1_net3081,
         pe_1_7_1_net3076, pe_1_7_1_net3071, pe_1_7_1_net3066,
         pe_1_7_1_net3061, pe_1_7_1_net3056, pe_1_7_1_net3051,
         pe_1_7_1_net3045, pe_1_7_1_N90, pe_1_7_1_N85, pe_1_7_1_N84,
         pe_1_7_1_N83, pe_1_7_1_N82, pe_1_7_1_N81, pe_1_7_1_N80, pe_1_7_1_N79,
         pe_1_7_1_N77, pe_1_7_1_N76, pe_1_7_1_N75, pe_1_7_1_N74, pe_1_7_1_N73,
         pe_1_7_1_N72, pe_1_7_1_N71, pe_1_7_1_N70, pe_1_7_1_int_data_0_,
         pe_1_7_1_int_data_1_, pe_1_7_1_int_data_2_, pe_1_7_1_int_data_3_,
         pe_1_7_1_N64, pe_1_7_1_N63, pe_1_7_1_N62, pe_1_7_1_N61, pe_1_7_1_N60,
         pe_1_7_1_N59, pe_1_7_2_n90, pe_1_7_2_n89, pe_1_7_2_n88, pe_1_7_2_n87,
         pe_1_7_2_n86, pe_1_7_2_n85, pe_1_7_2_n84, pe_1_7_2_n83, pe_1_7_2_n82,
         pe_1_7_2_n81, pe_1_7_2_n80, pe_1_7_2_n79, pe_1_7_2_n78, pe_1_7_2_n77,
         pe_1_7_2_n76, pe_1_7_2_n75, pe_1_7_2_n74, pe_1_7_2_n73, pe_1_7_2_n72,
         pe_1_7_2_n71, pe_1_7_2_n70, pe_1_7_2_n69, pe_1_7_2_n68, pe_1_7_2_n67,
         pe_1_7_2_n66, pe_1_7_2_n65, pe_1_7_2_n64, pe_1_7_2_n63, pe_1_7_2_n62,
         pe_1_7_2_n61, pe_1_7_2_n60, pe_1_7_2_n59, pe_1_7_2_n58, pe_1_7_2_n57,
         pe_1_7_2_n56, pe_1_7_2_n55, pe_1_7_2_n54, pe_1_7_2_n53, pe_1_7_2_n52,
         pe_1_7_2_n51, pe_1_7_2_n50, pe_1_7_2_n49, pe_1_7_2_n48, pe_1_7_2_n47,
         pe_1_7_2_n46, pe_1_7_2_n45, pe_1_7_2_n25, pe_1_7_2_n24, pe_1_7_2_n23,
         pe_1_7_2_n22, pe_1_7_2_n21, pe_1_7_2_n20, pe_1_7_2_n19, pe_1_7_2_n18,
         pe_1_7_2_n17, pe_1_7_2_n16, pe_1_7_2_n15, pe_1_7_2_n14, pe_1_7_2_n13,
         pe_1_7_2_n12, pe_1_7_2_n11, pe_1_7_2_n10, pe_1_7_2_n9, pe_1_7_2_n8,
         pe_1_7_2_n7, pe_1_7_2_n6, pe_1_7_2_n5, pe_1_7_2_n4, pe_1_7_2_n3,
         pe_1_7_2_n2, pe_1_7_2_n1, pe_1_7_2_n44, pe_1_7_2_n43, pe_1_7_2_n42,
         pe_1_7_2_n41, pe_1_7_2_n40, pe_1_7_2_n39, pe_1_7_2_n38, pe_1_7_2_n37,
         pe_1_7_2_n36, pe_1_7_2_n35, pe_1_7_2_n34, pe_1_7_2_n33, pe_1_7_2_n32,
         pe_1_7_2_n31, pe_1_7_2_n30, pe_1_7_2_n29, pe_1_7_2_n28, pe_1_7_2_n27,
         pe_1_7_2_n26, pe_1_7_2_net3028, pe_1_7_2_net3023, pe_1_7_2_net3018,
         pe_1_7_2_net3013, pe_1_7_2_net3008, pe_1_7_2_net3003,
         pe_1_7_2_net2998, pe_1_7_2_net2993, pe_1_7_2_net2988,
         pe_1_7_2_net2983, pe_1_7_2_net2978, pe_1_7_2_net2973,
         pe_1_7_2_net2967, pe_1_7_2_N90, pe_1_7_2_N85, pe_1_7_2_N84,
         pe_1_7_2_N83, pe_1_7_2_N82, pe_1_7_2_N81, pe_1_7_2_N80, pe_1_7_2_N79,
         pe_1_7_2_N77, pe_1_7_2_N76, pe_1_7_2_N75, pe_1_7_2_N74, pe_1_7_2_N73,
         pe_1_7_2_N72, pe_1_7_2_N71, pe_1_7_2_N70, pe_1_7_2_int_data_0_,
         pe_1_7_2_int_data_1_, pe_1_7_2_int_data_2_, pe_1_7_2_int_data_3_,
         pe_1_7_2_N64, pe_1_7_2_N63, pe_1_7_2_N62, pe_1_7_2_N61, pe_1_7_2_N60,
         pe_1_7_2_N59, pe_1_7_3_n90, pe_1_7_3_n89, pe_1_7_3_n88, pe_1_7_3_n87,
         pe_1_7_3_n86, pe_1_7_3_n85, pe_1_7_3_n84, pe_1_7_3_n83, pe_1_7_3_n82,
         pe_1_7_3_n81, pe_1_7_3_n80, pe_1_7_3_n79, pe_1_7_3_n78, pe_1_7_3_n77,
         pe_1_7_3_n76, pe_1_7_3_n75, pe_1_7_3_n74, pe_1_7_3_n73, pe_1_7_3_n72,
         pe_1_7_3_n71, pe_1_7_3_n70, pe_1_7_3_n69, pe_1_7_3_n68, pe_1_7_3_n67,
         pe_1_7_3_n66, pe_1_7_3_n65, pe_1_7_3_n64, pe_1_7_3_n63, pe_1_7_3_n62,
         pe_1_7_3_n61, pe_1_7_3_n60, pe_1_7_3_n59, pe_1_7_3_n58, pe_1_7_3_n57,
         pe_1_7_3_n56, pe_1_7_3_n55, pe_1_7_3_n54, pe_1_7_3_n53, pe_1_7_3_n52,
         pe_1_7_3_n51, pe_1_7_3_n50, pe_1_7_3_n49, pe_1_7_3_n48, pe_1_7_3_n47,
         pe_1_7_3_n46, pe_1_7_3_n45, pe_1_7_3_n25, pe_1_7_3_n24, pe_1_7_3_n23,
         pe_1_7_3_n22, pe_1_7_3_n21, pe_1_7_3_n20, pe_1_7_3_n19, pe_1_7_3_n18,
         pe_1_7_3_n17, pe_1_7_3_n16, pe_1_7_3_n15, pe_1_7_3_n14, pe_1_7_3_n13,
         pe_1_7_3_n12, pe_1_7_3_n11, pe_1_7_3_n10, pe_1_7_3_n9, pe_1_7_3_n8,
         pe_1_7_3_n7, pe_1_7_3_n6, pe_1_7_3_n5, pe_1_7_3_n4, pe_1_7_3_n3,
         pe_1_7_3_n2, pe_1_7_3_n1, pe_1_7_3_n44, pe_1_7_3_n43, pe_1_7_3_n42,
         pe_1_7_3_n41, pe_1_7_3_n40, pe_1_7_3_n39, pe_1_7_3_n38, pe_1_7_3_n37,
         pe_1_7_3_n36, pe_1_7_3_n35, pe_1_7_3_n34, pe_1_7_3_n33, pe_1_7_3_n32,
         pe_1_7_3_n31, pe_1_7_3_n30, pe_1_7_3_n29, pe_1_7_3_n28, pe_1_7_3_n27,
         pe_1_7_3_n26, pe_1_7_3_net2950, pe_1_7_3_net2945, pe_1_7_3_net2940,
         pe_1_7_3_net2935, pe_1_7_3_net2930, pe_1_7_3_net2925,
         pe_1_7_3_net2920, pe_1_7_3_net2915, pe_1_7_3_net2910,
         pe_1_7_3_net2905, pe_1_7_3_net2900, pe_1_7_3_net2895,
         pe_1_7_3_net2889, pe_1_7_3_N90, pe_1_7_3_N85, pe_1_7_3_N84,
         pe_1_7_3_N83, pe_1_7_3_N82, pe_1_7_3_N81, pe_1_7_3_N80, pe_1_7_3_N79,
         pe_1_7_3_N77, pe_1_7_3_N76, pe_1_7_3_N75, pe_1_7_3_N74, pe_1_7_3_N73,
         pe_1_7_3_N72, pe_1_7_3_N71, pe_1_7_3_N70, pe_1_7_3_int_data_0_,
         pe_1_7_3_int_data_1_, pe_1_7_3_int_data_2_, pe_1_7_3_int_data_3_,
         pe_1_7_3_N64, pe_1_7_3_N63, pe_1_7_3_N62, pe_1_7_3_N61, pe_1_7_3_N60,
         pe_1_7_3_N59, pe_1_7_4_n84, pe_1_7_4_n83, pe_1_7_4_n82, pe_1_7_4_n81,
         pe_1_7_4_n80, pe_1_7_4_n79, pe_1_7_4_n78, pe_1_7_4_n77, pe_1_7_4_n76,
         pe_1_7_4_n75, pe_1_7_4_n74, pe_1_7_4_n73, pe_1_7_4_n72, pe_1_7_4_n71,
         pe_1_7_4_n70, pe_1_7_4_n69, pe_1_7_4_n68, pe_1_7_4_n67, pe_1_7_4_n66,
         pe_1_7_4_n65, pe_1_7_4_n64, pe_1_7_4_n63, pe_1_7_4_n62, pe_1_7_4_n61,
         pe_1_7_4_n60, pe_1_7_4_n59, pe_1_7_4_n58, pe_1_7_4_n57, pe_1_7_4_n56,
         pe_1_7_4_n55, pe_1_7_4_n54, pe_1_7_4_n53, pe_1_7_4_n52, pe_1_7_4_n51,
         pe_1_7_4_n50, pe_1_7_4_n49, pe_1_7_4_n48, pe_1_7_4_n47, pe_1_7_4_n46,
         pe_1_7_4_n45, pe_1_7_4_n25, pe_1_7_4_n24, pe_1_7_4_n23, pe_1_7_4_n22,
         pe_1_7_4_n21, pe_1_7_4_n20, pe_1_7_4_n19, pe_1_7_4_n18, pe_1_7_4_n17,
         pe_1_7_4_n16, pe_1_7_4_n15, pe_1_7_4_n14, pe_1_7_4_n13, pe_1_7_4_n12,
         pe_1_7_4_n11, pe_1_7_4_n10, pe_1_7_4_n9, pe_1_7_4_n8, pe_1_7_4_n7,
         pe_1_7_4_n6, pe_1_7_4_n5, pe_1_7_4_n4, pe_1_7_4_n3, pe_1_7_4_n2,
         pe_1_7_4_n1, pe_1_7_4_n44, pe_1_7_4_n43, pe_1_7_4_n42, pe_1_7_4_n41,
         pe_1_7_4_n40, pe_1_7_4_n39, pe_1_7_4_n38, pe_1_7_4_n37, pe_1_7_4_n36,
         pe_1_7_4_n35, pe_1_7_4_n34, pe_1_7_4_n33, pe_1_7_4_n32, pe_1_7_4_n31,
         pe_1_7_4_n30, pe_1_7_4_n29, pe_1_7_4_n28, pe_1_7_4_n27, pe_1_7_4_n26,
         pe_1_7_4_net2872, pe_1_7_4_net2867, pe_1_7_4_net2862,
         pe_1_7_4_net2857, pe_1_7_4_net2852, pe_1_7_4_net2847,
         pe_1_7_4_net2842, pe_1_7_4_net2837, pe_1_7_4_net2832,
         pe_1_7_4_net2827, pe_1_7_4_net2822, pe_1_7_4_net2817,
         pe_1_7_4_net2811, pe_1_7_4_N90, pe_1_7_4_N85, pe_1_7_4_N84,
         pe_1_7_4_N83, pe_1_7_4_N82, pe_1_7_4_N81, pe_1_7_4_N80, pe_1_7_4_N79,
         pe_1_7_4_N77, pe_1_7_4_N76, pe_1_7_4_N75, pe_1_7_4_N74, pe_1_7_4_N73,
         pe_1_7_4_N72, pe_1_7_4_N71, pe_1_7_4_N70, pe_1_7_4_int_data_0_,
         pe_1_7_4_int_data_1_, pe_1_7_4_int_data_2_, pe_1_7_4_int_data_3_,
         pe_1_7_4_N64, pe_1_7_4_N63, pe_1_7_4_N62, pe_1_7_4_N61, pe_1_7_4_N60,
         pe_1_7_4_N59, pe_1_7_5_n84, pe_1_7_5_n83, pe_1_7_5_n82, pe_1_7_5_n81,
         pe_1_7_5_n80, pe_1_7_5_n79, pe_1_7_5_n78, pe_1_7_5_n77, pe_1_7_5_n76,
         pe_1_7_5_n75, pe_1_7_5_n74, pe_1_7_5_n73, pe_1_7_5_n72, pe_1_7_5_n71,
         pe_1_7_5_n70, pe_1_7_5_n69, pe_1_7_5_n68, pe_1_7_5_n67, pe_1_7_5_n66,
         pe_1_7_5_n65, pe_1_7_5_n64, pe_1_7_5_n63, pe_1_7_5_n62, pe_1_7_5_n61,
         pe_1_7_5_n60, pe_1_7_5_n59, pe_1_7_5_n58, pe_1_7_5_n57, pe_1_7_5_n56,
         pe_1_7_5_n55, pe_1_7_5_n54, pe_1_7_5_n53, pe_1_7_5_n52, pe_1_7_5_n51,
         pe_1_7_5_n50, pe_1_7_5_n49, pe_1_7_5_n48, pe_1_7_5_n47, pe_1_7_5_n46,
         pe_1_7_5_n45, pe_1_7_5_n25, pe_1_7_5_n24, pe_1_7_5_n23, pe_1_7_5_n22,
         pe_1_7_5_n21, pe_1_7_5_n20, pe_1_7_5_n19, pe_1_7_5_n18, pe_1_7_5_n17,
         pe_1_7_5_n16, pe_1_7_5_n15, pe_1_7_5_n14, pe_1_7_5_n13, pe_1_7_5_n12,
         pe_1_7_5_n11, pe_1_7_5_n10, pe_1_7_5_n9, pe_1_7_5_n8, pe_1_7_5_n7,
         pe_1_7_5_n6, pe_1_7_5_n5, pe_1_7_5_n4, pe_1_7_5_n3, pe_1_7_5_n2,
         pe_1_7_5_n1, pe_1_7_5_n44, pe_1_7_5_n43, pe_1_7_5_n42, pe_1_7_5_n41,
         pe_1_7_5_n40, pe_1_7_5_n39, pe_1_7_5_n38, pe_1_7_5_n37, pe_1_7_5_n36,
         pe_1_7_5_n35, pe_1_7_5_n34, pe_1_7_5_n33, pe_1_7_5_n32, pe_1_7_5_n31,
         pe_1_7_5_n30, pe_1_7_5_n29, pe_1_7_5_n28, pe_1_7_5_n27, pe_1_7_5_n26,
         pe_1_7_5_net2794, pe_1_7_5_net2789, pe_1_7_5_net2784,
         pe_1_7_5_net2779, pe_1_7_5_net2774, pe_1_7_5_net2769,
         pe_1_7_5_net2764, pe_1_7_5_net2759, pe_1_7_5_net2754,
         pe_1_7_5_net2749, pe_1_7_5_net2744, pe_1_7_5_net2739,
         pe_1_7_5_net2733, pe_1_7_5_N90, pe_1_7_5_N85, pe_1_7_5_N84,
         pe_1_7_5_N83, pe_1_7_5_N82, pe_1_7_5_N81, pe_1_7_5_N80, pe_1_7_5_N79,
         pe_1_7_5_N77, pe_1_7_5_N76, pe_1_7_5_N75, pe_1_7_5_N74, pe_1_7_5_N73,
         pe_1_7_5_N72, pe_1_7_5_N71, pe_1_7_5_N70, pe_1_7_5_int_data_0_,
         pe_1_7_5_int_data_1_, pe_1_7_5_int_data_2_, pe_1_7_5_int_data_3_,
         pe_1_7_5_N64, pe_1_7_5_N63, pe_1_7_5_N62, pe_1_7_5_N61, pe_1_7_5_N60,
         pe_1_7_5_N59, pe_1_7_6_n85, pe_1_7_6_n84, pe_1_7_6_n83, pe_1_7_6_n82,
         pe_1_7_6_n81, pe_1_7_6_n80, pe_1_7_6_n79, pe_1_7_6_n78, pe_1_7_6_n77,
         pe_1_7_6_n76, pe_1_7_6_n75, pe_1_7_6_n74, pe_1_7_6_n73, pe_1_7_6_n72,
         pe_1_7_6_n71, pe_1_7_6_n70, pe_1_7_6_n69, pe_1_7_6_n68, pe_1_7_6_n67,
         pe_1_7_6_n66, pe_1_7_6_n65, pe_1_7_6_n64, pe_1_7_6_n63, pe_1_7_6_n62,
         pe_1_7_6_n61, pe_1_7_6_n60, pe_1_7_6_n59, pe_1_7_6_n58, pe_1_7_6_n57,
         pe_1_7_6_n56, pe_1_7_6_n55, pe_1_7_6_n54, pe_1_7_6_n53, pe_1_7_6_n52,
         pe_1_7_6_n51, pe_1_7_6_n50, pe_1_7_6_n49, pe_1_7_6_n48, pe_1_7_6_n47,
         pe_1_7_6_n46, pe_1_7_6_n45, pe_1_7_6_n25, pe_1_7_6_n24, pe_1_7_6_n23,
         pe_1_7_6_n22, pe_1_7_6_n21, pe_1_7_6_n20, pe_1_7_6_n19, pe_1_7_6_n18,
         pe_1_7_6_n17, pe_1_7_6_n16, pe_1_7_6_n15, pe_1_7_6_n14, pe_1_7_6_n13,
         pe_1_7_6_n12, pe_1_7_6_n11, pe_1_7_6_n10, pe_1_7_6_n9, pe_1_7_6_n8,
         pe_1_7_6_n7, pe_1_7_6_n6, pe_1_7_6_n5, pe_1_7_6_n4, pe_1_7_6_n3,
         pe_1_7_6_n2, pe_1_7_6_n1, pe_1_7_6_n44, pe_1_7_6_n43, pe_1_7_6_n42,
         pe_1_7_6_n41, pe_1_7_6_n40, pe_1_7_6_n39, pe_1_7_6_n38, pe_1_7_6_n37,
         pe_1_7_6_n36, pe_1_7_6_n35, pe_1_7_6_n34, pe_1_7_6_n33, pe_1_7_6_n32,
         pe_1_7_6_n31, pe_1_7_6_n30, pe_1_7_6_n29, pe_1_7_6_n28, pe_1_7_6_n27,
         pe_1_7_6_n26, pe_1_7_6_net2716, pe_1_7_6_net2711, pe_1_7_6_net2706,
         pe_1_7_6_net2701, pe_1_7_6_net2696, pe_1_7_6_net2691,
         pe_1_7_6_net2686, pe_1_7_6_net2681, pe_1_7_6_net2676,
         pe_1_7_6_net2671, pe_1_7_6_net2666, pe_1_7_6_net2661,
         pe_1_7_6_net2655, pe_1_7_6_N90, pe_1_7_6_N85, pe_1_7_6_N84,
         pe_1_7_6_N83, pe_1_7_6_N82, pe_1_7_6_N81, pe_1_7_6_N80, pe_1_7_6_N79,
         pe_1_7_6_N77, pe_1_7_6_N76, pe_1_7_6_N75, pe_1_7_6_N74, pe_1_7_6_N73,
         pe_1_7_6_N72, pe_1_7_6_N71, pe_1_7_6_N70, pe_1_7_6_int_data_0_,
         pe_1_7_6_int_data_1_, pe_1_7_6_int_data_2_, pe_1_7_6_int_data_3_,
         pe_1_7_6_N64, pe_1_7_6_N63, pe_1_7_6_N62, pe_1_7_6_N61, pe_1_7_6_N60,
         pe_1_7_6_N59, pe_1_7_7_n86, pe_1_7_7_n85, pe_1_7_7_n84, pe_1_7_7_n83,
         pe_1_7_7_n82, pe_1_7_7_n81, pe_1_7_7_n80, pe_1_7_7_n79, pe_1_7_7_n78,
         pe_1_7_7_n77, pe_1_7_7_n76, pe_1_7_7_n75, pe_1_7_7_n74, pe_1_7_7_n73,
         pe_1_7_7_n72, pe_1_7_7_n71, pe_1_7_7_n70, pe_1_7_7_n69, pe_1_7_7_n68,
         pe_1_7_7_n67, pe_1_7_7_n66, pe_1_7_7_n65, pe_1_7_7_n64, pe_1_7_7_n63,
         pe_1_7_7_n62, pe_1_7_7_n61, pe_1_7_7_n60, pe_1_7_7_n59, pe_1_7_7_n58,
         pe_1_7_7_n57, pe_1_7_7_n56, pe_1_7_7_n55, pe_1_7_7_n54, pe_1_7_7_n53,
         pe_1_7_7_n52, pe_1_7_7_n51, pe_1_7_7_n50, pe_1_7_7_n49, pe_1_7_7_n48,
         pe_1_7_7_n47, pe_1_7_7_n46, pe_1_7_7_n45, pe_1_7_7_n25, pe_1_7_7_n24,
         pe_1_7_7_n23, pe_1_7_7_n22, pe_1_7_7_n21, pe_1_7_7_n20, pe_1_7_7_n19,
         pe_1_7_7_n18, pe_1_7_7_n17, pe_1_7_7_n16, pe_1_7_7_n15, pe_1_7_7_n14,
         pe_1_7_7_n13, pe_1_7_7_n12, pe_1_7_7_n11, pe_1_7_7_n10, pe_1_7_7_n9,
         pe_1_7_7_n8, pe_1_7_7_n7, pe_1_7_7_n6, pe_1_7_7_n5, pe_1_7_7_n4,
         pe_1_7_7_n3, pe_1_7_7_n2, pe_1_7_7_n1, pe_1_7_7_n44, pe_1_7_7_n43,
         pe_1_7_7_n42, pe_1_7_7_n41, pe_1_7_7_n40, pe_1_7_7_n39, pe_1_7_7_n38,
         pe_1_7_7_n37, pe_1_7_7_n36, pe_1_7_7_n35, pe_1_7_7_n34, pe_1_7_7_n33,
         pe_1_7_7_n32, pe_1_7_7_n31, pe_1_7_7_n30, pe_1_7_7_n29, pe_1_7_7_n28,
         pe_1_7_7_n27, pe_1_7_7_n26, pe_1_7_7_net2638, pe_1_7_7_net2633,
         pe_1_7_7_net2628, pe_1_7_7_net2623, pe_1_7_7_net2618,
         pe_1_7_7_net2613, pe_1_7_7_net2608, pe_1_7_7_net2603,
         pe_1_7_7_net2598, pe_1_7_7_net2593, pe_1_7_7_net2588,
         pe_1_7_7_net2583, pe_1_7_7_net2577, pe_1_7_7_N90, pe_1_7_7_N85,
         pe_1_7_7_N84, pe_1_7_7_N83, pe_1_7_7_N82, pe_1_7_7_N81, pe_1_7_7_N80,
         pe_1_7_7_N79, pe_1_7_7_N77, pe_1_7_7_N76, pe_1_7_7_N75, pe_1_7_7_N74,
         pe_1_7_7_N73, pe_1_7_7_N72, pe_1_7_7_N71, pe_1_7_7_N70,
         pe_1_7_7_int_data_0_, pe_1_7_7_int_data_1_, pe_1_7_7_int_data_2_,
         pe_1_7_7_int_data_3_, pe_1_7_7_N64, pe_1_7_7_N63, pe_1_7_7_N62,
         pe_1_7_7_N61, pe_1_7_7_N60, pe_1_7_7_N59;
  wire   [63:0] int_ckg;
  wire   [1:7] pe_1_0_0_sub_81_carry;
  wire   [2:7] pe_1_0_0_add_83_carry;
  wire   [23:0] pe_1_0_0_int_q_reg_v;
  wire   [23:0] pe_1_0_0_int_q_reg_h;
  wire   [1:7] pe_1_0_1_sub_81_carry;
  wire   [2:7] pe_1_0_1_add_83_carry;
  wire   [23:0] pe_1_0_1_int_q_reg_v;
  wire   [23:0] pe_1_0_1_int_q_reg_h;
  wire   [1:7] pe_1_0_2_sub_81_carry;
  wire   [2:7] pe_1_0_2_add_83_carry;
  wire   [23:0] pe_1_0_2_int_q_reg_v;
  wire   [23:0] pe_1_0_2_int_q_reg_h;
  wire   [1:7] pe_1_0_3_sub_81_carry;
  wire   [2:7] pe_1_0_3_add_83_carry;
  wire   [23:0] pe_1_0_3_int_q_reg_v;
  wire   [23:0] pe_1_0_3_int_q_reg_h;
  wire   [1:7] pe_1_0_4_sub_81_carry;
  wire   [2:7] pe_1_0_4_add_83_carry;
  wire   [23:0] pe_1_0_4_int_q_reg_v;
  wire   [23:0] pe_1_0_4_int_q_reg_h;
  wire   [1:7] pe_1_0_5_sub_81_carry;
  wire   [2:7] pe_1_0_5_add_83_carry;
  wire   [23:0] pe_1_0_5_int_q_reg_v;
  wire   [23:0] pe_1_0_5_int_q_reg_h;
  wire   [1:7] pe_1_0_6_sub_81_carry;
  wire   [2:7] pe_1_0_6_add_83_carry;
  wire   [23:0] pe_1_0_6_int_q_reg_v;
  wire   [23:0] pe_1_0_6_int_q_reg_h;
  wire   [1:7] pe_1_0_7_sub_81_carry;
  wire   [2:7] pe_1_0_7_add_83_carry;
  wire   [23:0] pe_1_0_7_int_q_reg_v;
  wire   [23:0] pe_1_0_7_int_q_reg_h;
  wire   [1:7] pe_1_1_0_sub_81_carry;
  wire   [2:7] pe_1_1_0_add_83_carry;
  wire   [23:0] pe_1_1_0_int_q_reg_v;
  wire   [23:0] pe_1_1_0_int_q_reg_h;
  wire   [1:7] pe_1_1_1_sub_81_carry;
  wire   [2:7] pe_1_1_1_add_83_carry;
  wire   [23:0] pe_1_1_1_int_q_reg_v;
  wire   [23:0] pe_1_1_1_int_q_reg_h;
  wire   [1:7] pe_1_1_2_sub_81_carry;
  wire   [2:7] pe_1_1_2_add_83_carry;
  wire   [23:0] pe_1_1_2_int_q_reg_v;
  wire   [23:0] pe_1_1_2_int_q_reg_h;
  wire   [1:7] pe_1_1_3_sub_81_carry;
  wire   [2:7] pe_1_1_3_add_83_carry;
  wire   [23:0] pe_1_1_3_int_q_reg_v;
  wire   [23:0] pe_1_1_3_int_q_reg_h;
  wire   [1:7] pe_1_1_4_sub_81_carry;
  wire   [2:7] pe_1_1_4_add_83_carry;
  wire   [23:0] pe_1_1_4_int_q_reg_v;
  wire   [23:0] pe_1_1_4_int_q_reg_h;
  wire   [1:7] pe_1_1_5_sub_81_carry;
  wire   [2:7] pe_1_1_5_add_83_carry;
  wire   [23:0] pe_1_1_5_int_q_reg_v;
  wire   [23:0] pe_1_1_5_int_q_reg_h;
  wire   [1:7] pe_1_1_6_sub_81_carry;
  wire   [2:7] pe_1_1_6_add_83_carry;
  wire   [23:0] pe_1_1_6_int_q_reg_v;
  wire   [23:0] pe_1_1_6_int_q_reg_h;
  wire   [1:7] pe_1_1_7_sub_81_carry;
  wire   [2:7] pe_1_1_7_add_83_carry;
  wire   [23:0] pe_1_1_7_int_q_reg_v;
  wire   [23:0] pe_1_1_7_int_q_reg_h;
  wire   [1:7] pe_1_2_0_sub_81_carry;
  wire   [2:7] pe_1_2_0_add_83_carry;
  wire   [23:0] pe_1_2_0_int_q_reg_v;
  wire   [23:0] pe_1_2_0_int_q_reg_h;
  wire   [1:7] pe_1_2_1_sub_81_carry;
  wire   [2:7] pe_1_2_1_add_83_carry;
  wire   [23:0] pe_1_2_1_int_q_reg_v;
  wire   [23:0] pe_1_2_1_int_q_reg_h;
  wire   [1:7] pe_1_2_2_sub_81_carry;
  wire   [2:7] pe_1_2_2_add_83_carry;
  wire   [23:0] pe_1_2_2_int_q_reg_v;
  wire   [23:0] pe_1_2_2_int_q_reg_h;
  wire   [1:7] pe_1_2_3_sub_81_carry;
  wire   [2:7] pe_1_2_3_add_83_carry;
  wire   [23:0] pe_1_2_3_int_q_reg_v;
  wire   [23:0] pe_1_2_3_int_q_reg_h;
  wire   [1:7] pe_1_2_4_sub_81_carry;
  wire   [2:7] pe_1_2_4_add_83_carry;
  wire   [23:0] pe_1_2_4_int_q_reg_v;
  wire   [23:0] pe_1_2_4_int_q_reg_h;
  wire   [1:7] pe_1_2_5_sub_81_carry;
  wire   [2:7] pe_1_2_5_add_83_carry;
  wire   [23:0] pe_1_2_5_int_q_reg_v;
  wire   [23:0] pe_1_2_5_int_q_reg_h;
  wire   [1:7] pe_1_2_6_sub_81_carry;
  wire   [2:7] pe_1_2_6_add_83_carry;
  wire   [23:0] pe_1_2_6_int_q_reg_v;
  wire   [23:0] pe_1_2_6_int_q_reg_h;
  wire   [1:7] pe_1_2_7_sub_81_carry;
  wire   [2:7] pe_1_2_7_add_83_carry;
  wire   [23:0] pe_1_2_7_int_q_reg_v;
  wire   [23:0] pe_1_2_7_int_q_reg_h;
  wire   [1:7] pe_1_3_0_sub_81_carry;
  wire   [2:7] pe_1_3_0_add_83_carry;
  wire   [23:0] pe_1_3_0_int_q_reg_v;
  wire   [23:0] pe_1_3_0_int_q_reg_h;
  wire   [1:7] pe_1_3_1_sub_81_carry;
  wire   [2:7] pe_1_3_1_add_83_carry;
  wire   [23:0] pe_1_3_1_int_q_reg_v;
  wire   [23:0] pe_1_3_1_int_q_reg_h;
  wire   [1:7] pe_1_3_2_sub_81_carry;
  wire   [2:7] pe_1_3_2_add_83_carry;
  wire   [23:0] pe_1_3_2_int_q_reg_v;
  wire   [23:0] pe_1_3_2_int_q_reg_h;
  wire   [1:7] pe_1_3_3_sub_81_carry;
  wire   [2:7] pe_1_3_3_add_83_carry;
  wire   [23:0] pe_1_3_3_int_q_reg_v;
  wire   [23:0] pe_1_3_3_int_q_reg_h;
  wire   [1:7] pe_1_3_4_sub_81_carry;
  wire   [2:7] pe_1_3_4_add_83_carry;
  wire   [23:0] pe_1_3_4_int_q_reg_v;
  wire   [23:0] pe_1_3_4_int_q_reg_h;
  wire   [1:7] pe_1_3_5_sub_81_carry;
  wire   [2:7] pe_1_3_5_add_83_carry;
  wire   [23:0] pe_1_3_5_int_q_reg_v;
  wire   [23:0] pe_1_3_5_int_q_reg_h;
  wire   [1:7] pe_1_3_6_sub_81_carry;
  wire   [2:7] pe_1_3_6_add_83_carry;
  wire   [23:0] pe_1_3_6_int_q_reg_v;
  wire   [23:0] pe_1_3_6_int_q_reg_h;
  wire   [1:7] pe_1_3_7_sub_81_carry;
  wire   [2:7] pe_1_3_7_add_83_carry;
  wire   [23:0] pe_1_3_7_int_q_reg_v;
  wire   [23:0] pe_1_3_7_int_q_reg_h;
  wire   [1:7] pe_1_4_0_sub_81_carry;
  wire   [2:7] pe_1_4_0_add_83_carry;
  wire   [23:0] pe_1_4_0_int_q_reg_v;
  wire   [23:0] pe_1_4_0_int_q_reg_h;
  wire   [1:7] pe_1_4_1_sub_81_carry;
  wire   [2:7] pe_1_4_1_add_83_carry;
  wire   [23:0] pe_1_4_1_int_q_reg_v;
  wire   [23:0] pe_1_4_1_int_q_reg_h;
  wire   [1:7] pe_1_4_2_sub_81_carry;
  wire   [2:7] pe_1_4_2_add_83_carry;
  wire   [23:0] pe_1_4_2_int_q_reg_v;
  wire   [23:0] pe_1_4_2_int_q_reg_h;
  wire   [1:7] pe_1_4_3_sub_81_carry;
  wire   [2:7] pe_1_4_3_add_83_carry;
  wire   [23:0] pe_1_4_3_int_q_reg_v;
  wire   [23:0] pe_1_4_3_int_q_reg_h;
  wire   [1:7] pe_1_4_4_sub_81_carry;
  wire   [2:7] pe_1_4_4_add_83_carry;
  wire   [23:0] pe_1_4_4_int_q_reg_v;
  wire   [23:0] pe_1_4_4_int_q_reg_h;
  wire   [1:7] pe_1_4_5_sub_81_carry;
  wire   [2:7] pe_1_4_5_add_83_carry;
  wire   [23:0] pe_1_4_5_int_q_reg_v;
  wire   [23:0] pe_1_4_5_int_q_reg_h;
  wire   [1:7] pe_1_4_6_sub_81_carry;
  wire   [2:7] pe_1_4_6_add_83_carry;
  wire   [23:0] pe_1_4_6_int_q_reg_v;
  wire   [23:0] pe_1_4_6_int_q_reg_h;
  wire   [1:7] pe_1_4_7_sub_81_carry;
  wire   [2:7] pe_1_4_7_add_83_carry;
  wire   [23:0] pe_1_4_7_int_q_reg_v;
  wire   [23:0] pe_1_4_7_int_q_reg_h;
  wire   [1:7] pe_1_5_0_sub_81_carry;
  wire   [2:7] pe_1_5_0_add_83_carry;
  wire   [23:0] pe_1_5_0_int_q_reg_v;
  wire   [23:0] pe_1_5_0_int_q_reg_h;
  wire   [1:7] pe_1_5_1_sub_81_carry;
  wire   [2:7] pe_1_5_1_add_83_carry;
  wire   [23:0] pe_1_5_1_int_q_reg_v;
  wire   [23:0] pe_1_5_1_int_q_reg_h;
  wire   [1:7] pe_1_5_2_sub_81_carry;
  wire   [2:7] pe_1_5_2_add_83_carry;
  wire   [23:0] pe_1_5_2_int_q_reg_v;
  wire   [23:0] pe_1_5_2_int_q_reg_h;
  wire   [1:7] pe_1_5_3_sub_81_carry;
  wire   [2:7] pe_1_5_3_add_83_carry;
  wire   [23:0] pe_1_5_3_int_q_reg_v;
  wire   [23:0] pe_1_5_3_int_q_reg_h;
  wire   [1:7] pe_1_5_4_sub_81_carry;
  wire   [2:7] pe_1_5_4_add_83_carry;
  wire   [23:0] pe_1_5_4_int_q_reg_v;
  wire   [23:0] pe_1_5_4_int_q_reg_h;
  wire   [1:7] pe_1_5_5_sub_81_carry;
  wire   [2:7] pe_1_5_5_add_83_carry;
  wire   [23:0] pe_1_5_5_int_q_reg_v;
  wire   [23:0] pe_1_5_5_int_q_reg_h;
  wire   [1:7] pe_1_5_6_sub_81_carry;
  wire   [2:7] pe_1_5_6_add_83_carry;
  wire   [23:0] pe_1_5_6_int_q_reg_v;
  wire   [23:0] pe_1_5_6_int_q_reg_h;
  wire   [1:7] pe_1_5_7_sub_81_carry;
  wire   [2:7] pe_1_5_7_add_83_carry;
  wire   [23:0] pe_1_5_7_int_q_reg_v;
  wire   [23:0] pe_1_5_7_int_q_reg_h;
  wire   [1:7] pe_1_6_0_sub_81_carry;
  wire   [2:7] pe_1_6_0_add_83_carry;
  wire   [23:0] pe_1_6_0_int_q_reg_v;
  wire   [23:0] pe_1_6_0_int_q_reg_h;
  wire   [1:7] pe_1_6_1_sub_81_carry;
  wire   [2:7] pe_1_6_1_add_83_carry;
  wire   [23:0] pe_1_6_1_int_q_reg_v;
  wire   [23:0] pe_1_6_1_int_q_reg_h;
  wire   [1:7] pe_1_6_2_sub_81_carry;
  wire   [2:7] pe_1_6_2_add_83_carry;
  wire   [23:0] pe_1_6_2_int_q_reg_v;
  wire   [23:0] pe_1_6_2_int_q_reg_h;
  wire   [1:7] pe_1_6_3_sub_81_carry;
  wire   [2:7] pe_1_6_3_add_83_carry;
  wire   [23:0] pe_1_6_3_int_q_reg_v;
  wire   [23:0] pe_1_6_3_int_q_reg_h;
  wire   [1:7] pe_1_6_4_sub_81_carry;
  wire   [2:7] pe_1_6_4_add_83_carry;
  wire   [23:0] pe_1_6_4_int_q_reg_v;
  wire   [23:0] pe_1_6_4_int_q_reg_h;
  wire   [1:7] pe_1_6_5_sub_81_carry;
  wire   [2:7] pe_1_6_5_add_83_carry;
  wire   [23:0] pe_1_6_5_int_q_reg_v;
  wire   [23:0] pe_1_6_5_int_q_reg_h;
  wire   [1:7] pe_1_6_6_sub_81_carry;
  wire   [2:7] pe_1_6_6_add_83_carry;
  wire   [23:0] pe_1_6_6_int_q_reg_v;
  wire   [23:0] pe_1_6_6_int_q_reg_h;
  wire   [1:7] pe_1_6_7_sub_81_carry;
  wire   [2:7] pe_1_6_7_add_83_carry;
  wire   [23:0] pe_1_6_7_int_q_reg_v;
  wire   [23:0] pe_1_6_7_int_q_reg_h;
  wire   [1:7] pe_1_7_0_sub_81_carry;
  wire   [2:7] pe_1_7_0_add_83_carry;
  wire   [23:0] pe_1_7_0_int_q_reg_v;
  wire   [23:0] pe_1_7_0_int_q_reg_h;
  wire   [1:7] pe_1_7_1_sub_81_carry;
  wire   [2:7] pe_1_7_1_add_83_carry;
  wire   [23:0] pe_1_7_1_int_q_reg_v;
  wire   [23:0] pe_1_7_1_int_q_reg_h;
  wire   [1:7] pe_1_7_2_sub_81_carry;
  wire   [2:7] pe_1_7_2_add_83_carry;
  wire   [23:0] pe_1_7_2_int_q_reg_v;
  wire   [23:0] pe_1_7_2_int_q_reg_h;
  wire   [1:7] pe_1_7_3_sub_81_carry;
  wire   [2:7] pe_1_7_3_add_83_carry;
  wire   [23:0] pe_1_7_3_int_q_reg_v;
  wire   [23:0] pe_1_7_3_int_q_reg_h;
  wire   [1:7] pe_1_7_4_sub_81_carry;
  wire   [2:7] pe_1_7_4_add_83_carry;
  wire   [23:0] pe_1_7_4_int_q_reg_v;
  wire   [23:0] pe_1_7_4_int_q_reg_h;
  wire   [1:7] pe_1_7_5_sub_81_carry;
  wire   [2:7] pe_1_7_5_add_83_carry;
  wire   [23:0] pe_1_7_5_int_q_reg_v;
  wire   [23:0] pe_1_7_5_int_q_reg_h;
  wire   [1:7] pe_1_7_6_sub_81_carry;
  wire   [2:7] pe_1_7_6_add_83_carry;
  wire   [23:0] pe_1_7_6_int_q_reg_v;
  wire   [23:0] pe_1_7_6_int_q_reg_h;
  wire   [1:7] pe_1_7_7_sub_81_carry;
  wire   [2:7] pe_1_7_7_add_83_carry;
  wire   [23:0] pe_1_7_7_int_q_reg_v;
  wire   [23:0] pe_1_7_7_int_q_reg_h;

  CLKBUF_X1 U81 ( .A(rst), .Z(n81) );
  BUF_X1 U82 ( .A(n24), .Z(n19) );
  BUF_X1 U83 ( .A(n24), .Z(n18) );
  BUF_X1 U84 ( .A(n24), .Z(n17) );
  BUF_X1 U85 ( .A(n23), .Z(n21) );
  BUF_X1 U86 ( .A(n23), .Z(n20) );
  BUF_X2 U87 ( .A(n56), .Z(n55) );
  BUF_X2 U88 ( .A(n72), .Z(n67) );
  BUF_X2 U89 ( .A(n72), .Z(n66) );
  BUF_X2 U90 ( .A(n72), .Z(n65) );
  BUF_X2 U91 ( .A(n71), .Z(n69) );
  BUF_X2 U92 ( .A(n71), .Z(n68) );
  BUF_X1 U93 ( .A(n80), .Z(n73) );
  BUF_X1 U94 ( .A(n80), .Z(n74) );
  BUF_X1 U95 ( .A(n80), .Z(n75) );
  BUF_X1 U96 ( .A(n79), .Z(n76) );
  BUF_X1 U97 ( .A(n79), .Z(n77) );
  BUF_X1 U98 ( .A(n71), .Z(n70) );
  NAND2_X1 U99 ( .A1(n87), .A2(n95), .ZN(int_ckg[63]) );
  NAND2_X1 U100 ( .A1(n87), .A2(n96), .ZN(int_ckg[62]) );
  NAND2_X1 U101 ( .A1(n87), .A2(n97), .ZN(int_ckg[61]) );
  NAND2_X1 U102 ( .A1(n87), .A2(n98), .ZN(int_ckg[60]) );
  NAND2_X1 U103 ( .A1(n87), .A2(n99), .ZN(int_ckg[59]) );
  NAND2_X1 U104 ( .A1(n87), .A2(n100), .ZN(int_ckg[58]) );
  NAND2_X1 U105 ( .A1(n87), .A2(n101), .ZN(int_ckg[57]) );
  NAND2_X1 U106 ( .A1(n87), .A2(n102), .ZN(int_ckg[56]) );
  NAND2_X1 U107 ( .A1(n88), .A2(n95), .ZN(int_ckg[55]) );
  NAND2_X1 U108 ( .A1(n88), .A2(n96), .ZN(int_ckg[54]) );
  NAND2_X1 U109 ( .A1(n88), .A2(n97), .ZN(int_ckg[53]) );
  NAND2_X1 U110 ( .A1(n88), .A2(n98), .ZN(int_ckg[52]) );
  NAND2_X1 U111 ( .A1(n88), .A2(n99), .ZN(int_ckg[51]) );
  NAND2_X1 U112 ( .A1(n88), .A2(n100), .ZN(int_ckg[50]) );
  NAND2_X1 U113 ( .A1(n88), .A2(n101), .ZN(int_ckg[49]) );
  NAND2_X1 U114 ( .A1(n88), .A2(n102), .ZN(int_ckg[48]) );
  NAND2_X1 U115 ( .A1(n89), .A2(n95), .ZN(int_ckg[47]) );
  NAND2_X1 U116 ( .A1(n89), .A2(n96), .ZN(int_ckg[46]) );
  NAND2_X1 U117 ( .A1(n89), .A2(n97), .ZN(int_ckg[45]) );
  NAND2_X1 U118 ( .A1(n89), .A2(n98), .ZN(int_ckg[44]) );
  NAND2_X1 U119 ( .A1(n89), .A2(n99), .ZN(int_ckg[43]) );
  NAND2_X1 U120 ( .A1(n89), .A2(n100), .ZN(int_ckg[42]) );
  NAND2_X1 U121 ( .A1(n89), .A2(n101), .ZN(int_ckg[41]) );
  NAND2_X1 U122 ( .A1(n89), .A2(n102), .ZN(int_ckg[40]) );
  NAND2_X1 U123 ( .A1(n90), .A2(n95), .ZN(int_ckg[39]) );
  NAND2_X1 U124 ( .A1(n90), .A2(n96), .ZN(int_ckg[38]) );
  NAND2_X1 U125 ( .A1(n90), .A2(n97), .ZN(int_ckg[37]) );
  NAND2_X1 U126 ( .A1(n90), .A2(n98), .ZN(int_ckg[36]) );
  NAND2_X1 U127 ( .A1(n90), .A2(n99), .ZN(int_ckg[35]) );
  NAND2_X1 U128 ( .A1(n90), .A2(n100), .ZN(int_ckg[34]) );
  NAND2_X1 U129 ( .A1(n90), .A2(n101), .ZN(int_ckg[33]) );
  NAND2_X1 U130 ( .A1(n90), .A2(n102), .ZN(int_ckg[32]) );
  NAND2_X1 U131 ( .A1(n91), .A2(n95), .ZN(int_ckg[31]) );
  NAND2_X1 U132 ( .A1(n91), .A2(n96), .ZN(int_ckg[30]) );
  NAND2_X1 U133 ( .A1(n91), .A2(n97), .ZN(int_ckg[29]) );
  NAND2_X1 U134 ( .A1(n91), .A2(n98), .ZN(int_ckg[28]) );
  NAND2_X1 U135 ( .A1(n91), .A2(n99), .ZN(int_ckg[27]) );
  NAND2_X1 U136 ( .A1(n91), .A2(n100), .ZN(int_ckg[26]) );
  NAND2_X1 U137 ( .A1(n91), .A2(n101), .ZN(int_ckg[25]) );
  NAND2_X1 U138 ( .A1(n91), .A2(n102), .ZN(int_ckg[24]) );
  NAND2_X1 U139 ( .A1(n92), .A2(n95), .ZN(int_ckg[23]) );
  NAND2_X1 U140 ( .A1(n92), .A2(n96), .ZN(int_ckg[22]) );
  NAND2_X1 U141 ( .A1(n92), .A2(n97), .ZN(int_ckg[21]) );
  NAND2_X1 U142 ( .A1(n92), .A2(n98), .ZN(int_ckg[20]) );
  NAND2_X1 U143 ( .A1(n92), .A2(n99), .ZN(int_ckg[19]) );
  NAND2_X1 U144 ( .A1(n92), .A2(n100), .ZN(int_ckg[18]) );
  NAND2_X1 U145 ( .A1(n92), .A2(n101), .ZN(int_ckg[17]) );
  NAND2_X1 U146 ( .A1(n92), .A2(n102), .ZN(int_ckg[16]) );
  NAND2_X1 U147 ( .A1(n93), .A2(n95), .ZN(int_ckg[15]) );
  NAND2_X1 U148 ( .A1(n93), .A2(n96), .ZN(int_ckg[14]) );
  NAND2_X1 U149 ( .A1(n93), .A2(n97), .ZN(int_ckg[13]) );
  NAND2_X1 U150 ( .A1(n93), .A2(n98), .ZN(int_ckg[12]) );
  NAND2_X1 U151 ( .A1(n93), .A2(n99), .ZN(int_ckg[11]) );
  NAND2_X1 U152 ( .A1(n93), .A2(n100), .ZN(int_ckg[10]) );
  NAND2_X1 U153 ( .A1(n93), .A2(n101), .ZN(int_ckg[9]) );
  NAND2_X1 U154 ( .A1(n93), .A2(n102), .ZN(int_ckg[8]) );
  NAND2_X1 U155 ( .A1(n94), .A2(n95), .ZN(int_ckg[7]) );
  NAND2_X1 U156 ( .A1(n94), .A2(n96), .ZN(int_ckg[6]) );
  NAND2_X1 U157 ( .A1(n94), .A2(n97), .ZN(int_ckg[5]) );
  NAND2_X1 U158 ( .A1(n94), .A2(n98), .ZN(int_ckg[4]) );
  NAND2_X1 U159 ( .A1(n94), .A2(n99), .ZN(int_ckg[3]) );
  NAND2_X1 U160 ( .A1(n94), .A2(n100), .ZN(int_ckg[2]) );
  NAND2_X1 U161 ( .A1(n94), .A2(n101), .ZN(int_ckg[1]) );
  NAND2_X1 U162 ( .A1(n94), .A2(n102), .ZN(int_ckg[0]) );
  BUF_X1 U163 ( .A(n23), .Z(n22) );
  BUF_X1 U164 ( .A(n79), .Z(n78) );
  BUF_X1 U165 ( .A(i_ifmap_ptr[0]), .Z(n35) );
  BUF_X1 U166 ( .A(i_ifmap_ptr[0]), .Z(n34) );
  BUF_X1 U167 ( .A(i_ifmap_ptr[0]), .Z(n33) );
  BUF_X1 U168 ( .A(i_ifmap_ptr[0]), .Z(n32) );
  BUF_X1 U169 ( .A(i_ifmap_ptr[0]), .Z(n31) );
  BUF_X1 U170 ( .A(wr_pipe), .Z(n59) );
  BUF_X1 U171 ( .A(wr_pipe), .Z(n60) );
  BUF_X1 U172 ( .A(wr_pipe), .Z(n61) );
  BUF_X1 U173 ( .A(wr_pipe), .Z(n62) );
  BUF_X1 U174 ( .A(wr_pipe), .Z(n63) );
  BUF_X1 U175 ( .A(i_ifmap_ptr[1]), .Z(n41) );
  BUF_X1 U176 ( .A(i_ifmap_ptr[1]), .Z(n40) );
  BUF_X1 U177 ( .A(i_ifmap_ptr[1]), .Z(n39) );
  BUF_X1 U178 ( .A(i_ifmap_ptr[1]), .Z(n38) );
  BUF_X1 U179 ( .A(i_ifmap_ptr[1]), .Z(n37) );
  BUF_X1 U180 ( .A(ldh_v_n), .Z(n72) );
  BUF_X1 U181 ( .A(i_weight[1]), .Z(n29) );
  BUF_X1 U182 ( .A(i_weight[1]), .Z(n28) );
  BUF_X1 U183 ( .A(i_weight[1]), .Z(n27) );
  BUF_X1 U184 ( .A(i_weight[1]), .Z(n26) );
  BUF_X1 U185 ( .A(i_weight[1]), .Z(n25) );
  BUF_X1 U186 ( .A(ldh_v_n), .Z(n71) );
  BUF_X1 U187 ( .A(i_weight[0]), .Z(n24) );
  BUF_X1 U188 ( .A(en), .Z(n80) );
  BUF_X1 U189 ( .A(i_weight[0]), .Z(n23) );
  BUF_X1 U190 ( .A(en), .Z(n79) );
  BUF_X1 U191 ( .A(i_ifmap_ptr[2]), .Z(n56) );
  BUF_X1 U192 ( .A(i_ifmap_ptr[2]), .Z(n57) );
  BUF_X1 U193 ( .A(i_ifmap_ptr[2]), .Z(n58) );
  INV_X1 U194 ( .A(ckg_cmask[0]), .ZN(n95) );
  INV_X1 U195 ( .A(ckg_cmask[1]), .ZN(n96) );
  INV_X1 U196 ( .A(ckg_cmask[2]), .ZN(n97) );
  INV_X1 U197 ( .A(ckg_cmask[3]), .ZN(n98) );
  INV_X1 U198 ( .A(ckg_cmask[4]), .ZN(n99) );
  INV_X1 U199 ( .A(ckg_cmask[5]), .ZN(n100) );
  INV_X1 U200 ( .A(ckg_cmask[6]), .ZN(n101) );
  INV_X1 U201 ( .A(ckg_cmask[7]), .ZN(n102) );
  INV_X1 U202 ( .A(ckg_rmask[0]), .ZN(n87) );
  INV_X1 U203 ( .A(ckg_rmask[1]), .ZN(n88) );
  INV_X1 U204 ( .A(ckg_rmask[2]), .ZN(n89) );
  INV_X1 U205 ( .A(ckg_rmask[3]), .ZN(n90) );
  INV_X1 U206 ( .A(ckg_rmask[4]), .ZN(n91) );
  INV_X1 U207 ( .A(ckg_rmask[5]), .ZN(n92) );
  INV_X1 U208 ( .A(ckg_rmask[6]), .ZN(n93) );
  INV_X1 U209 ( .A(ckg_rmask[7]), .ZN(n94) );
  BUF_X1 U210 ( .A(rst), .Z(n85) );
  BUF_X1 U211 ( .A(rst), .Z(n84) );
  BUF_X1 U212 ( .A(rst), .Z(n83) );
  BUF_X1 U213 ( .A(rst), .Z(n82) );
  CLKBUF_X1 U214 ( .A(i_weight[1]), .Z(n30) );
  CLKBUF_X1 U215 ( .A(i_ifmap_ptr[0]), .Z(n36) );
  CLKBUF_X1 U216 ( .A(i_ifmap_ptr[1]), .Z(n42) );
  CLKBUF_X3 U217 ( .A(n58), .Z(n43) );
  CLKBUF_X3 U218 ( .A(n58), .Z(n44) );
  CLKBUF_X3 U219 ( .A(n58), .Z(n45) );
  CLKBUF_X3 U220 ( .A(n57), .Z(n46) );
  CLKBUF_X3 U221 ( .A(n57), .Z(n47) );
  CLKBUF_X3 U222 ( .A(n57), .Z(n48) );
  CLKBUF_X3 U223 ( .A(n57), .Z(n49) );
  CLKBUF_X3 U224 ( .A(n57), .Z(n50) );
  CLKBUF_X3 U225 ( .A(n56), .Z(n51) );
  CLKBUF_X3 U226 ( .A(n56), .Z(n52) );
  CLKBUF_X3 U227 ( .A(n56), .Z(n53) );
  CLKBUF_X3 U228 ( .A(n56), .Z(n54) );
  CLKBUF_X1 U229 ( .A(wr_pipe), .Z(n64) );
  CLKBUF_X1 U230 ( .A(rst), .Z(n86) );
  CLKBUF_X1 pe_1_0_0_U109 ( .A(pe_1_0_0_n69), .Z(pe_1_0_0_n68) );
  INV_X1 pe_1_0_0_U108 ( .A(n73), .ZN(pe_1_0_0_n67) );
  INV_X1 pe_1_0_0_U107 ( .A(n65), .ZN(pe_1_0_0_n66) );
  INV_X1 pe_1_0_0_U106 ( .A(n65), .ZN(pe_1_0_0_n65) );
  INV_X1 pe_1_0_0_U105 ( .A(pe_1_0_0_n66), .ZN(pe_1_0_0_n64) );
  INV_X1 pe_1_0_0_U104 ( .A(pe_1_0_0_n61), .ZN(pe_1_0_0_n60) );
  INV_X1 pe_1_0_0_U103 ( .A(n25), .ZN(pe_1_0_0_n58) );
  INV_X1 pe_1_0_0_U102 ( .A(n17), .ZN(pe_1_0_0_n57) );
  MUX2_X1 pe_1_0_0_U101 ( .A(pe_1_0_0_n54), .B(pe_1_0_0_n51), .S(n43), .Z(
        pe_1_0_0_o_data_h_3_) );
  MUX2_X1 pe_1_0_0_U100 ( .A(pe_1_0_0_n53), .B(pe_1_0_0_n52), .S(pe_1_0_0_n60), 
        .Z(pe_1_0_0_n54) );
  MUX2_X1 pe_1_0_0_U99 ( .A(pe_1_0_0_int_q_reg_h[23]), .B(
        pe_1_0_0_int_q_reg_h[19]), .S(pe_1_0_0_n56), .Z(pe_1_0_0_n53) );
  MUX2_X1 pe_1_0_0_U98 ( .A(pe_1_0_0_int_q_reg_h[15]), .B(
        pe_1_0_0_int_q_reg_h[11]), .S(pe_1_0_0_n56), .Z(pe_1_0_0_n52) );
  MUX2_X1 pe_1_0_0_U97 ( .A(pe_1_0_0_int_q_reg_h[7]), .B(
        pe_1_0_0_int_q_reg_h[3]), .S(pe_1_0_0_n56), .Z(pe_1_0_0_n51) );
  MUX2_X1 pe_1_0_0_U96 ( .A(pe_1_0_0_n50), .B(pe_1_0_0_n47), .S(n43), .Z(
        pe_1_0_0_o_data_h_2_) );
  MUX2_X1 pe_1_0_0_U95 ( .A(pe_1_0_0_n49), .B(pe_1_0_0_n48), .S(pe_1_0_0_n60), 
        .Z(pe_1_0_0_n50) );
  MUX2_X1 pe_1_0_0_U94 ( .A(pe_1_0_0_int_q_reg_h[22]), .B(
        pe_1_0_0_int_q_reg_h[18]), .S(pe_1_0_0_n56), .Z(pe_1_0_0_n49) );
  MUX2_X1 pe_1_0_0_U93 ( .A(pe_1_0_0_int_q_reg_h[14]), .B(
        pe_1_0_0_int_q_reg_h[10]), .S(pe_1_0_0_n56), .Z(pe_1_0_0_n48) );
  MUX2_X1 pe_1_0_0_U92 ( .A(pe_1_0_0_int_q_reg_h[6]), .B(
        pe_1_0_0_int_q_reg_h[2]), .S(pe_1_0_0_n56), .Z(pe_1_0_0_n47) );
  MUX2_X1 pe_1_0_0_U91 ( .A(pe_1_0_0_n46), .B(pe_1_0_0_n24), .S(n43), .Z(
        pe_1_0_0_o_data_h_1_) );
  MUX2_X1 pe_1_0_0_U90 ( .A(pe_1_0_0_n45), .B(pe_1_0_0_n25), .S(pe_1_0_0_n60), 
        .Z(pe_1_0_0_n46) );
  MUX2_X1 pe_1_0_0_U89 ( .A(pe_1_0_0_int_q_reg_h[21]), .B(
        pe_1_0_0_int_q_reg_h[17]), .S(pe_1_0_0_n56), .Z(pe_1_0_0_n45) );
  MUX2_X1 pe_1_0_0_U88 ( .A(pe_1_0_0_int_q_reg_h[13]), .B(
        pe_1_0_0_int_q_reg_h[9]), .S(pe_1_0_0_n56), .Z(pe_1_0_0_n25) );
  MUX2_X1 pe_1_0_0_U87 ( .A(pe_1_0_0_int_q_reg_h[5]), .B(
        pe_1_0_0_int_q_reg_h[1]), .S(pe_1_0_0_n56), .Z(pe_1_0_0_n24) );
  MUX2_X1 pe_1_0_0_U86 ( .A(pe_1_0_0_n23), .B(pe_1_0_0_n20), .S(n43), .Z(
        pe_1_0_0_o_data_h_0_) );
  MUX2_X1 pe_1_0_0_U85 ( .A(pe_1_0_0_n22), .B(pe_1_0_0_n21), .S(pe_1_0_0_n60), 
        .Z(pe_1_0_0_n23) );
  MUX2_X1 pe_1_0_0_U84 ( .A(pe_1_0_0_int_q_reg_h[20]), .B(
        pe_1_0_0_int_q_reg_h[16]), .S(pe_1_0_0_n56), .Z(pe_1_0_0_n22) );
  MUX2_X1 pe_1_0_0_U83 ( .A(pe_1_0_0_int_q_reg_h[12]), .B(
        pe_1_0_0_int_q_reg_h[8]), .S(pe_1_0_0_n56), .Z(pe_1_0_0_n21) );
  MUX2_X1 pe_1_0_0_U82 ( .A(pe_1_0_0_int_q_reg_h[4]), .B(
        pe_1_0_0_int_q_reg_h[0]), .S(pe_1_0_0_n56), .Z(pe_1_0_0_n20) );
  MUX2_X1 pe_1_0_0_U81 ( .A(pe_1_0_0_n19), .B(pe_1_0_0_n16), .S(n43), .Z(
        pe_1_0_0_o_data_v_3_) );
  MUX2_X1 pe_1_0_0_U80 ( .A(pe_1_0_0_n18), .B(pe_1_0_0_n17), .S(pe_1_0_0_n60), 
        .Z(pe_1_0_0_n19) );
  MUX2_X1 pe_1_0_0_U79 ( .A(pe_1_0_0_int_q_reg_v[23]), .B(
        pe_1_0_0_int_q_reg_v[19]), .S(pe_1_0_0_n55), .Z(pe_1_0_0_n18) );
  MUX2_X1 pe_1_0_0_U78 ( .A(pe_1_0_0_int_q_reg_v[15]), .B(
        pe_1_0_0_int_q_reg_v[11]), .S(pe_1_0_0_n55), .Z(pe_1_0_0_n17) );
  MUX2_X1 pe_1_0_0_U77 ( .A(pe_1_0_0_int_q_reg_v[7]), .B(
        pe_1_0_0_int_q_reg_v[3]), .S(pe_1_0_0_n55), .Z(pe_1_0_0_n16) );
  MUX2_X1 pe_1_0_0_U76 ( .A(pe_1_0_0_n15), .B(pe_1_0_0_n12), .S(n43), .Z(
        pe_1_0_0_o_data_v_2_) );
  MUX2_X1 pe_1_0_0_U75 ( .A(pe_1_0_0_n14), .B(pe_1_0_0_n13), .S(pe_1_0_0_n60), 
        .Z(pe_1_0_0_n15) );
  MUX2_X1 pe_1_0_0_U74 ( .A(pe_1_0_0_int_q_reg_v[22]), .B(
        pe_1_0_0_int_q_reg_v[18]), .S(pe_1_0_0_n55), .Z(pe_1_0_0_n14) );
  MUX2_X1 pe_1_0_0_U73 ( .A(pe_1_0_0_int_q_reg_v[14]), .B(
        pe_1_0_0_int_q_reg_v[10]), .S(pe_1_0_0_n55), .Z(pe_1_0_0_n13) );
  MUX2_X1 pe_1_0_0_U72 ( .A(pe_1_0_0_int_q_reg_v[6]), .B(
        pe_1_0_0_int_q_reg_v[2]), .S(pe_1_0_0_n55), .Z(pe_1_0_0_n12) );
  MUX2_X1 pe_1_0_0_U71 ( .A(pe_1_0_0_n11), .B(pe_1_0_0_n8), .S(n43), .Z(
        pe_1_0_0_o_data_v_1_) );
  MUX2_X1 pe_1_0_0_U70 ( .A(pe_1_0_0_n10), .B(pe_1_0_0_n9), .S(pe_1_0_0_n60), 
        .Z(pe_1_0_0_n11) );
  MUX2_X1 pe_1_0_0_U69 ( .A(pe_1_0_0_int_q_reg_v[21]), .B(
        pe_1_0_0_int_q_reg_v[17]), .S(pe_1_0_0_n55), .Z(pe_1_0_0_n10) );
  MUX2_X1 pe_1_0_0_U68 ( .A(pe_1_0_0_int_q_reg_v[13]), .B(
        pe_1_0_0_int_q_reg_v[9]), .S(pe_1_0_0_n55), .Z(pe_1_0_0_n9) );
  MUX2_X1 pe_1_0_0_U67 ( .A(pe_1_0_0_int_q_reg_v[5]), .B(
        pe_1_0_0_int_q_reg_v[1]), .S(pe_1_0_0_n55), .Z(pe_1_0_0_n8) );
  MUX2_X1 pe_1_0_0_U66 ( .A(pe_1_0_0_n7), .B(pe_1_0_0_n4), .S(n43), .Z(
        pe_1_0_0_o_data_v_0_) );
  MUX2_X1 pe_1_0_0_U65 ( .A(pe_1_0_0_n6), .B(pe_1_0_0_n5), .S(pe_1_0_0_n60), 
        .Z(pe_1_0_0_n7) );
  MUX2_X1 pe_1_0_0_U64 ( .A(pe_1_0_0_int_q_reg_v[20]), .B(
        pe_1_0_0_int_q_reg_v[16]), .S(pe_1_0_0_n55), .Z(pe_1_0_0_n6) );
  MUX2_X1 pe_1_0_0_U63 ( .A(pe_1_0_0_int_q_reg_v[12]), .B(
        pe_1_0_0_int_q_reg_v[8]), .S(pe_1_0_0_n55), .Z(pe_1_0_0_n5) );
  MUX2_X1 pe_1_0_0_U62 ( .A(pe_1_0_0_int_q_reg_v[4]), .B(
        pe_1_0_0_int_q_reg_v[0]), .S(pe_1_0_0_n55), .Z(pe_1_0_0_n4) );
  AND2_X1 pe_1_0_0_U61 ( .A1(pe_1_0_0_o_data_h_3_), .A2(n25), .ZN(
        pe_1_0_0_int_data_3_) );
  AOI222_X1 pe_1_0_0_U60 ( .A1(pe_1_0_0_n62), .A2(int_data_res_1__0__7_), .B1(
        pe_1_0_0_N85), .B2(pe_1_0_0_n27), .C1(pe_1_0_0_N77), .C2(pe_1_0_0_n28), 
        .ZN(pe_1_0_0_n26) );
  INV_X1 pe_1_0_0_U59 ( .A(pe_1_0_0_n26), .ZN(pe_1_0_0_n74) );
  AOI222_X1 pe_1_0_0_U58 ( .A1(int_data_res_1__0__2_), .A2(pe_1_0_0_n62), .B1(
        pe_1_0_0_N80), .B2(pe_1_0_0_n27), .C1(pe_1_0_0_N72), .C2(pe_1_0_0_n28), 
        .ZN(pe_1_0_0_n33) );
  INV_X1 pe_1_0_0_U57 ( .A(pe_1_0_0_n33), .ZN(pe_1_0_0_n79) );
  AOI222_X1 pe_1_0_0_U52 ( .A1(int_data_res_1__0__3_), .A2(pe_1_0_0_n62), .B1(
        pe_1_0_0_N81), .B2(pe_1_0_0_n27), .C1(pe_1_0_0_N73), .C2(pe_1_0_0_n28), 
        .ZN(pe_1_0_0_n32) );
  INV_X1 pe_1_0_0_U51 ( .A(pe_1_0_0_n32), .ZN(pe_1_0_0_n78) );
  AOI222_X1 pe_1_0_0_U50 ( .A1(int_data_res_1__0__6_), .A2(pe_1_0_0_n62), .B1(
        pe_1_0_0_N84), .B2(pe_1_0_0_n27), .C1(pe_1_0_0_N76), .C2(pe_1_0_0_n28), 
        .ZN(pe_1_0_0_n29) );
  INV_X1 pe_1_0_0_U49 ( .A(pe_1_0_0_n29), .ZN(pe_1_0_0_n75) );
  AND2_X1 pe_1_0_0_U48 ( .A1(pe_1_0_0_o_data_h_2_), .A2(n25), .ZN(
        pe_1_0_0_int_data_2_) );
  AND2_X1 pe_1_0_0_U47 ( .A1(pe_1_0_0_o_data_h_1_), .A2(n25), .ZN(
        pe_1_0_0_int_data_1_) );
  INV_X1 pe_1_0_0_U46 ( .A(pe_1_0_0_int_data_2_), .ZN(pe_1_0_0_n72) );
  NAND2_X1 pe_1_0_0_U45 ( .A1(pe_1_0_0_int_data_0_), .A2(pe_1_0_0_n3), .ZN(
        pe_1_0_0_sub_81_carry[1]) );
  INV_X1 pe_1_0_0_U44 ( .A(pe_1_0_0_int_data_1_), .ZN(pe_1_0_0_n71) );
  AND2_X1 pe_1_0_0_U43 ( .A1(pe_1_0_0_int_data_0_), .A2(o_data[56]), .ZN(
        pe_1_0_0_n2) );
  AND2_X1 pe_1_0_0_U42 ( .A1(pe_1_0_0_o_data_h_0_), .A2(n25), .ZN(
        pe_1_0_0_int_data_0_) );
  XNOR2_X1 pe_1_0_0_U41 ( .A(pe_1_0_0_n70), .B(o_data[56]), .ZN(pe_1_0_0_N70)
         );
  AOI222_X1 pe_1_0_0_U40 ( .A1(int_data_res_1__0__0_), .A2(pe_1_0_0_n62), .B1(
        pe_1_0_0_n1), .B2(pe_1_0_0_n27), .C1(pe_1_0_0_N70), .C2(pe_1_0_0_n28), 
        .ZN(pe_1_0_0_n35) );
  INV_X1 pe_1_0_0_U39 ( .A(pe_1_0_0_n35), .ZN(pe_1_0_0_n81) );
  AOI222_X1 pe_1_0_0_U38 ( .A1(int_data_res_1__0__1_), .A2(pe_1_0_0_n62), .B1(
        pe_1_0_0_N79), .B2(pe_1_0_0_n27), .C1(pe_1_0_0_N71), .C2(pe_1_0_0_n28), 
        .ZN(pe_1_0_0_n34) );
  INV_X1 pe_1_0_0_U37 ( .A(pe_1_0_0_n34), .ZN(pe_1_0_0_n80) );
  AOI222_X1 pe_1_0_0_U36 ( .A1(int_data_res_1__0__4_), .A2(pe_1_0_0_n62), .B1(
        pe_1_0_0_N82), .B2(pe_1_0_0_n27), .C1(pe_1_0_0_N74), .C2(pe_1_0_0_n28), 
        .ZN(pe_1_0_0_n31) );
  INV_X1 pe_1_0_0_U35 ( .A(pe_1_0_0_n31), .ZN(pe_1_0_0_n77) );
  AOI222_X1 pe_1_0_0_U34 ( .A1(int_data_res_1__0__5_), .A2(pe_1_0_0_n62), .B1(
        pe_1_0_0_N83), .B2(pe_1_0_0_n27), .C1(pe_1_0_0_N75), .C2(pe_1_0_0_n28), 
        .ZN(pe_1_0_0_n30) );
  INV_X1 pe_1_0_0_U33 ( .A(pe_1_0_0_n30), .ZN(pe_1_0_0_n76) );
  NOR3_X1 pe_1_0_0_U32 ( .A1(pe_1_0_0_n58), .A2(pe_1_0_0_n63), .A3(int_ckg[63]), .ZN(pe_1_0_0_n36) );
  OR2_X1 pe_1_0_0_U31 ( .A1(pe_1_0_0_n36), .A2(pe_1_0_0_n62), .ZN(pe_1_0_0_N90) );
  INV_X1 pe_1_0_0_U30 ( .A(pe_1_0_0_int_data_0_), .ZN(pe_1_0_0_n70) );
  INV_X1 pe_1_0_0_U29 ( .A(n37), .ZN(pe_1_0_0_n61) );
  INV_X1 pe_1_0_0_U28 ( .A(n31), .ZN(pe_1_0_0_n59) );
  INV_X1 pe_1_0_0_U27 ( .A(pe_1_0_0_int_data_3_), .ZN(pe_1_0_0_n73) );
  BUF_X1 pe_1_0_0_U26 ( .A(n59), .Z(pe_1_0_0_n62) );
  NAND2_X1 pe_1_0_0_U25 ( .A1(pe_1_0_0_n44), .A2(pe_1_0_0_n59), .ZN(
        pe_1_0_0_n41) );
  AND3_X1 pe_1_0_0_U24 ( .A1(n73), .A2(pe_1_0_0_n61), .A3(n43), .ZN(
        pe_1_0_0_n44) );
  NOR2_X1 pe_1_0_0_U23 ( .A1(pe_1_0_0_n67), .A2(n43), .ZN(pe_1_0_0_n43) );
  NOR2_X1 pe_1_0_0_U22 ( .A1(pe_1_0_0_n57), .A2(pe_1_0_0_n62), .ZN(
        pe_1_0_0_n28) );
  NOR2_X1 pe_1_0_0_U21 ( .A1(n17), .A2(pe_1_0_0_n62), .ZN(pe_1_0_0_n27) );
  BUF_X1 pe_1_0_0_U20 ( .A(n31), .Z(pe_1_0_0_n55) );
  INV_X1 pe_1_0_0_U19 ( .A(pe_1_0_0_n41), .ZN(pe_1_0_0_n87) );
  INV_X1 pe_1_0_0_U18 ( .A(pe_1_0_0_n37), .ZN(pe_1_0_0_n85) );
  INV_X1 pe_1_0_0_U17 ( .A(pe_1_0_0_n38), .ZN(pe_1_0_0_n84) );
  INV_X1 pe_1_0_0_U16 ( .A(pe_1_0_0_n39), .ZN(pe_1_0_0_n83) );
  NOR2_X1 pe_1_0_0_U15 ( .A1(pe_1_0_0_n65), .A2(pe_1_0_0_n42), .ZN(
        pe_1_0_0_N59) );
  NOR2_X1 pe_1_0_0_U14 ( .A1(pe_1_0_0_n65), .A2(pe_1_0_0_n41), .ZN(
        pe_1_0_0_N60) );
  NOR2_X1 pe_1_0_0_U13 ( .A1(pe_1_0_0_n65), .A2(pe_1_0_0_n38), .ZN(
        pe_1_0_0_N63) );
  NOR2_X1 pe_1_0_0_U12 ( .A1(pe_1_0_0_n65), .A2(pe_1_0_0_n40), .ZN(
        pe_1_0_0_N61) );
  NOR2_X1 pe_1_0_0_U11 ( .A1(pe_1_0_0_n65), .A2(pe_1_0_0_n39), .ZN(
        pe_1_0_0_N62) );
  NOR2_X1 pe_1_0_0_U10 ( .A1(pe_1_0_0_n37), .A2(pe_1_0_0_n65), .ZN(
        pe_1_0_0_N64) );
  NAND2_X1 pe_1_0_0_U9 ( .A1(pe_1_0_0_n44), .A2(n31), .ZN(pe_1_0_0_n42) );
  BUF_X1 pe_1_0_0_U8 ( .A(n31), .Z(pe_1_0_0_n56) );
  INV_X1 pe_1_0_0_U7 ( .A(pe_1_0_0_n66), .ZN(pe_1_0_0_n63) );
  INV_X1 pe_1_0_0_U6 ( .A(pe_1_0_0_n42), .ZN(pe_1_0_0_n86) );
  INV_X1 pe_1_0_0_U5 ( .A(pe_1_0_0_n40), .ZN(pe_1_0_0_n82) );
  INV_X2 pe_1_0_0_U4 ( .A(n81), .ZN(pe_1_0_0_n69) );
  XOR2_X1 pe_1_0_0_U3 ( .A(pe_1_0_0_int_data_0_), .B(o_data[56]), .Z(
        pe_1_0_0_n1) );
  DFFR_X1 pe_1_0_0_int_q_acc_reg_0_ ( .D(pe_1_0_0_n81), .CK(pe_1_0_0_net7552), 
        .RN(pe_1_0_0_n69), .Q(o_data[56]), .QN(pe_1_0_0_n3) );
  DFFR_X1 pe_1_0_0_int_q_reg_v_reg_0__0_ ( .D(int_data_y_1__0__0_), .CK(
        pe_1_0_0_net7522), .RN(pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_v[20]) );
  DFFR_X1 pe_1_0_0_int_q_reg_v_reg_0__1_ ( .D(int_data_y_1__0__1_), .CK(
        pe_1_0_0_net7522), .RN(pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_v[21]) );
  DFFR_X1 pe_1_0_0_int_q_reg_v_reg_0__2_ ( .D(int_data_y_1__0__2_), .CK(
        pe_1_0_0_net7522), .RN(pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_v[22]) );
  DFFR_X1 pe_1_0_0_int_q_reg_v_reg_0__3_ ( .D(int_data_y_1__0__3_), .CK(
        pe_1_0_0_net7522), .RN(pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_v[23]) );
  DFFR_X1 pe_1_0_0_int_q_reg_v_reg_1__0_ ( .D(int_data_y_1__0__0_), .CK(
        pe_1_0_0_net7527), .RN(pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_v[16]) );
  DFFR_X1 pe_1_0_0_int_q_reg_v_reg_1__1_ ( .D(int_data_y_1__0__1_), .CK(
        pe_1_0_0_net7527), .RN(pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_v[17]) );
  DFFR_X1 pe_1_0_0_int_q_reg_v_reg_1__2_ ( .D(int_data_y_1__0__2_), .CK(
        pe_1_0_0_net7527), .RN(pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_v[18]) );
  DFFR_X1 pe_1_0_0_int_q_reg_v_reg_1__3_ ( .D(int_data_y_1__0__3_), .CK(
        pe_1_0_0_net7527), .RN(pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_v[19]) );
  DFFR_X1 pe_1_0_0_int_q_reg_v_reg_2__0_ ( .D(int_data_y_1__0__0_), .CK(
        pe_1_0_0_net7532), .RN(pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_v[12]) );
  DFFR_X1 pe_1_0_0_int_q_reg_v_reg_2__1_ ( .D(int_data_y_1__0__1_), .CK(
        pe_1_0_0_net7532), .RN(pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_v[13]) );
  DFFR_X1 pe_1_0_0_int_q_reg_v_reg_2__2_ ( .D(int_data_y_1__0__2_), .CK(
        pe_1_0_0_net7532), .RN(pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_v[14]) );
  DFFR_X1 pe_1_0_0_int_q_reg_v_reg_2__3_ ( .D(int_data_y_1__0__3_), .CK(
        pe_1_0_0_net7532), .RN(pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_v[15]) );
  DFFR_X1 pe_1_0_0_int_q_reg_v_reg_3__0_ ( .D(int_data_y_1__0__0_), .CK(
        pe_1_0_0_net7537), .RN(pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_v[8]) );
  DFFR_X1 pe_1_0_0_int_q_reg_v_reg_3__1_ ( .D(int_data_y_1__0__1_), .CK(
        pe_1_0_0_net7537), .RN(pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_v[9]) );
  DFFR_X1 pe_1_0_0_int_q_reg_v_reg_3__2_ ( .D(int_data_y_1__0__2_), .CK(
        pe_1_0_0_net7537), .RN(pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_v[10]) );
  DFFR_X1 pe_1_0_0_int_q_reg_v_reg_3__3_ ( .D(int_data_y_1__0__3_), .CK(
        pe_1_0_0_net7537), .RN(pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_v[11]) );
  DFFR_X1 pe_1_0_0_int_q_reg_v_reg_4__0_ ( .D(int_data_y_1__0__0_), .CK(
        pe_1_0_0_net7542), .RN(pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_v[4]) );
  DFFR_X1 pe_1_0_0_int_q_reg_v_reg_4__1_ ( .D(int_data_y_1__0__1_), .CK(
        pe_1_0_0_net7542), .RN(pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_v[5]) );
  DFFR_X1 pe_1_0_0_int_q_reg_v_reg_4__2_ ( .D(int_data_y_1__0__2_), .CK(
        pe_1_0_0_net7542), .RN(pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_v[6]) );
  DFFR_X1 pe_1_0_0_int_q_reg_v_reg_4__3_ ( .D(int_data_y_1__0__3_), .CK(
        pe_1_0_0_net7542), .RN(pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_v[7]) );
  DFFR_X1 pe_1_0_0_int_q_reg_v_reg_5__0_ ( .D(int_data_y_1__0__0_), .CK(
        pe_1_0_0_net7547), .RN(pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_v[0]) );
  DFFR_X1 pe_1_0_0_int_q_reg_v_reg_5__1_ ( .D(int_data_y_1__0__1_), .CK(
        pe_1_0_0_net7547), .RN(pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_v[1]) );
  DFFR_X1 pe_1_0_0_int_q_reg_v_reg_5__2_ ( .D(int_data_y_1__0__2_), .CK(
        pe_1_0_0_net7547), .RN(pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_v[2]) );
  DFFR_X1 pe_1_0_0_int_q_reg_v_reg_5__3_ ( .D(int_data_y_1__0__3_), .CK(
        pe_1_0_0_net7547), .RN(pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_0_0_int_q_reg_h_reg_0__0_ ( .D(int_data_x_0__1__0_), .SI(
        int_data_y_1__0__0_), .SE(pe_1_0_0_n63), .CK(pe_1_0_0_net7491), .RN(
        pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_0_0_int_q_reg_h_reg_0__1_ ( .D(int_data_x_0__1__1_), .SI(
        int_data_y_1__0__1_), .SE(pe_1_0_0_n63), .CK(pe_1_0_0_net7491), .RN(
        pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_0_0_int_q_reg_h_reg_0__2_ ( .D(int_data_x_0__1__2_), .SI(
        int_data_y_1__0__2_), .SE(pe_1_0_0_n63), .CK(pe_1_0_0_net7491), .RN(
        pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_0_0_int_q_reg_h_reg_0__3_ ( .D(int_data_x_0__1__3_), .SI(
        int_data_y_1__0__3_), .SE(pe_1_0_0_n63), .CK(pe_1_0_0_net7491), .RN(
        pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_0_0_int_q_reg_h_reg_1__0_ ( .D(int_data_x_0__1__0_), .SI(
        int_data_y_1__0__0_), .SE(pe_1_0_0_n63), .CK(pe_1_0_0_net7497), .RN(
        pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_0_0_int_q_reg_h_reg_1__1_ ( .D(int_data_x_0__1__1_), .SI(
        int_data_y_1__0__1_), .SE(pe_1_0_0_n63), .CK(pe_1_0_0_net7497), .RN(
        pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_0_0_int_q_reg_h_reg_1__2_ ( .D(int_data_x_0__1__2_), .SI(
        int_data_y_1__0__2_), .SE(pe_1_0_0_n63), .CK(pe_1_0_0_net7497), .RN(
        pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_0_0_int_q_reg_h_reg_1__3_ ( .D(int_data_x_0__1__3_), .SI(
        int_data_y_1__0__3_), .SE(pe_1_0_0_n63), .CK(pe_1_0_0_net7497), .RN(
        pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_0_0_int_q_reg_h_reg_2__0_ ( .D(int_data_x_0__1__0_), .SI(
        int_data_y_1__0__0_), .SE(pe_1_0_0_n63), .CK(pe_1_0_0_net7502), .RN(
        pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_0_0_int_q_reg_h_reg_2__1_ ( .D(int_data_x_0__1__1_), .SI(
        int_data_y_1__0__1_), .SE(pe_1_0_0_n63), .CK(pe_1_0_0_net7502), .RN(
        pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_0_0_int_q_reg_h_reg_2__2_ ( .D(int_data_x_0__1__2_), .SI(
        int_data_y_1__0__2_), .SE(pe_1_0_0_n63), .CK(pe_1_0_0_net7502), .RN(
        pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_0_0_int_q_reg_h_reg_2__3_ ( .D(int_data_x_0__1__3_), .SI(
        int_data_y_1__0__3_), .SE(pe_1_0_0_n63), .CK(pe_1_0_0_net7502), .RN(
        pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_0_0_int_q_reg_h_reg_3__0_ ( .D(int_data_x_0__1__0_), .SI(
        int_data_y_1__0__0_), .SE(pe_1_0_0_n63), .CK(pe_1_0_0_net7507), .RN(
        pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_0_0_int_q_reg_h_reg_3__1_ ( .D(int_data_x_0__1__1_), .SI(
        int_data_y_1__0__1_), .SE(pe_1_0_0_n63), .CK(pe_1_0_0_net7507), .RN(
        pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_0_0_int_q_reg_h_reg_3__2_ ( .D(int_data_x_0__1__2_), .SI(
        int_data_y_1__0__2_), .SE(pe_1_0_0_n63), .CK(pe_1_0_0_net7507), .RN(
        pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_0_0_int_q_reg_h_reg_3__3_ ( .D(int_data_x_0__1__3_), .SI(
        int_data_y_1__0__3_), .SE(pe_1_0_0_n63), .CK(pe_1_0_0_net7507), .RN(
        pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_0_0_int_q_reg_h_reg_4__0_ ( .D(int_data_x_0__1__0_), .SI(
        int_data_y_1__0__0_), .SE(pe_1_0_0_n64), .CK(pe_1_0_0_net7512), .RN(
        pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_0_0_int_q_reg_h_reg_4__1_ ( .D(int_data_x_0__1__1_), .SI(
        int_data_y_1__0__1_), .SE(pe_1_0_0_n64), .CK(pe_1_0_0_net7512), .RN(
        pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_0_0_int_q_reg_h_reg_4__2_ ( .D(int_data_x_0__1__2_), .SI(
        int_data_y_1__0__2_), .SE(pe_1_0_0_n64), .CK(pe_1_0_0_net7512), .RN(
        pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_0_0_int_q_reg_h_reg_4__3_ ( .D(int_data_x_0__1__3_), .SI(
        int_data_y_1__0__3_), .SE(pe_1_0_0_n64), .CK(pe_1_0_0_net7512), .RN(
        pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_0_0_int_q_reg_h_reg_5__0_ ( .D(int_data_x_0__1__0_), .SI(
        int_data_y_1__0__0_), .SE(pe_1_0_0_n64), .CK(pe_1_0_0_net7517), .RN(
        pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_0_0_int_q_reg_h_reg_5__1_ ( .D(int_data_x_0__1__1_), .SI(
        int_data_y_1__0__1_), .SE(pe_1_0_0_n64), .CK(pe_1_0_0_net7517), .RN(
        pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_0_0_int_q_reg_h_reg_5__2_ ( .D(int_data_x_0__1__2_), .SI(
        int_data_y_1__0__2_), .SE(pe_1_0_0_n64), .CK(pe_1_0_0_net7517), .RN(
        pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_0_0_int_q_reg_h_reg_5__3_ ( .D(int_data_x_0__1__3_), .SI(
        int_data_y_1__0__3_), .SE(pe_1_0_0_n64), .CK(pe_1_0_0_net7517), .RN(
        pe_1_0_0_n69), .Q(pe_1_0_0_int_q_reg_h[3]) );
  FA_X1 pe_1_0_0_sub_81_U2_7 ( .A(o_data[63]), .B(pe_1_0_0_n73), .CI(
        pe_1_0_0_sub_81_carry[7]), .S(pe_1_0_0_N77) );
  FA_X1 pe_1_0_0_sub_81_U2_6 ( .A(o_data[62]), .B(pe_1_0_0_n73), .CI(
        pe_1_0_0_sub_81_carry[6]), .CO(pe_1_0_0_sub_81_carry[7]), .S(
        pe_1_0_0_N76) );
  FA_X1 pe_1_0_0_sub_81_U2_5 ( .A(o_data[61]), .B(pe_1_0_0_n73), .CI(
        pe_1_0_0_sub_81_carry[5]), .CO(pe_1_0_0_sub_81_carry[6]), .S(
        pe_1_0_0_N75) );
  FA_X1 pe_1_0_0_sub_81_U2_4 ( .A(o_data[60]), .B(pe_1_0_0_n73), .CI(
        pe_1_0_0_sub_81_carry[4]), .CO(pe_1_0_0_sub_81_carry[5]), .S(
        pe_1_0_0_N74) );
  FA_X1 pe_1_0_0_sub_81_U2_3 ( .A(o_data[59]), .B(pe_1_0_0_n73), .CI(
        pe_1_0_0_sub_81_carry[3]), .CO(pe_1_0_0_sub_81_carry[4]), .S(
        pe_1_0_0_N73) );
  FA_X1 pe_1_0_0_sub_81_U2_2 ( .A(o_data[58]), .B(pe_1_0_0_n72), .CI(
        pe_1_0_0_sub_81_carry[2]), .CO(pe_1_0_0_sub_81_carry[3]), .S(
        pe_1_0_0_N72) );
  FA_X1 pe_1_0_0_sub_81_U2_1 ( .A(o_data[57]), .B(pe_1_0_0_n71), .CI(
        pe_1_0_0_sub_81_carry[1]), .CO(pe_1_0_0_sub_81_carry[2]), .S(
        pe_1_0_0_N71) );
  FA_X1 pe_1_0_0_add_83_U1_7 ( .A(o_data[63]), .B(pe_1_0_0_int_data_3_), .CI(
        pe_1_0_0_add_83_carry[7]), .S(pe_1_0_0_N85) );
  FA_X1 pe_1_0_0_add_83_U1_6 ( .A(o_data[62]), .B(pe_1_0_0_int_data_3_), .CI(
        pe_1_0_0_add_83_carry[6]), .CO(pe_1_0_0_add_83_carry[7]), .S(
        pe_1_0_0_N84) );
  FA_X1 pe_1_0_0_add_83_U1_5 ( .A(o_data[61]), .B(pe_1_0_0_int_data_3_), .CI(
        pe_1_0_0_add_83_carry[5]), .CO(pe_1_0_0_add_83_carry[6]), .S(
        pe_1_0_0_N83) );
  FA_X1 pe_1_0_0_add_83_U1_4 ( .A(o_data[60]), .B(pe_1_0_0_int_data_3_), .CI(
        pe_1_0_0_add_83_carry[4]), .CO(pe_1_0_0_add_83_carry[5]), .S(
        pe_1_0_0_N82) );
  FA_X1 pe_1_0_0_add_83_U1_3 ( .A(o_data[59]), .B(pe_1_0_0_int_data_3_), .CI(
        pe_1_0_0_add_83_carry[3]), .CO(pe_1_0_0_add_83_carry[4]), .S(
        pe_1_0_0_N81) );
  FA_X1 pe_1_0_0_add_83_U1_2 ( .A(o_data[58]), .B(pe_1_0_0_int_data_2_), .CI(
        pe_1_0_0_add_83_carry[2]), .CO(pe_1_0_0_add_83_carry[3]), .S(
        pe_1_0_0_N80) );
  FA_X1 pe_1_0_0_add_83_U1_1 ( .A(o_data[57]), .B(pe_1_0_0_int_data_1_), .CI(
        pe_1_0_0_n2), .CO(pe_1_0_0_add_83_carry[2]), .S(pe_1_0_0_N79) );
  NAND3_X1 pe_1_0_0_U56 ( .A1(n31), .A2(pe_1_0_0_n43), .A3(pe_1_0_0_n60), .ZN(
        pe_1_0_0_n40) );
  NAND3_X1 pe_1_0_0_U55 ( .A1(pe_1_0_0_n43), .A2(pe_1_0_0_n59), .A3(
        pe_1_0_0_n60), .ZN(pe_1_0_0_n39) );
  NAND3_X1 pe_1_0_0_U54 ( .A1(pe_1_0_0_n43), .A2(pe_1_0_0_n61), .A3(n31), .ZN(
        pe_1_0_0_n38) );
  NAND3_X1 pe_1_0_0_U53 ( .A1(pe_1_0_0_n59), .A2(pe_1_0_0_n61), .A3(
        pe_1_0_0_n43), .ZN(pe_1_0_0_n37) );
  DFFR_X1 pe_1_0_0_int_q_acc_reg_6_ ( .D(pe_1_0_0_n75), .CK(pe_1_0_0_net7552), 
        .RN(pe_1_0_0_n68), .Q(o_data[62]) );
  DFFR_X1 pe_1_0_0_int_q_acc_reg_5_ ( .D(pe_1_0_0_n76), .CK(pe_1_0_0_net7552), 
        .RN(pe_1_0_0_n68), .Q(o_data[61]) );
  DFFR_X1 pe_1_0_0_int_q_acc_reg_4_ ( .D(pe_1_0_0_n77), .CK(pe_1_0_0_net7552), 
        .RN(pe_1_0_0_n68), .Q(o_data[60]) );
  DFFR_X1 pe_1_0_0_int_q_acc_reg_3_ ( .D(pe_1_0_0_n78), .CK(pe_1_0_0_net7552), 
        .RN(pe_1_0_0_n68), .Q(o_data[59]) );
  DFFR_X1 pe_1_0_0_int_q_acc_reg_2_ ( .D(pe_1_0_0_n79), .CK(pe_1_0_0_net7552), 
        .RN(pe_1_0_0_n68), .Q(o_data[58]) );
  DFFR_X1 pe_1_0_0_int_q_acc_reg_1_ ( .D(pe_1_0_0_n80), .CK(pe_1_0_0_net7552), 
        .RN(pe_1_0_0_n68), .Q(o_data[57]) );
  DFFR_X1 pe_1_0_0_int_q_acc_reg_7_ ( .D(pe_1_0_0_n74), .CK(pe_1_0_0_net7552), 
        .RN(pe_1_0_0_n68), .Q(o_data[63]) );
  CLKGATETST_X1 pe_1_0_0_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_0_0_n85), .SE(1'b0), .GCK(pe_1_0_0_net7491) );
  CLKGATETST_X1 pe_1_0_0_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_0_0_n84), .SE(1'b0), .GCK(pe_1_0_0_net7497) );
  CLKGATETST_X1 pe_1_0_0_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_0_0_n83), .SE(1'b0), .GCK(pe_1_0_0_net7502) );
  CLKGATETST_X1 pe_1_0_0_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_0_0_n82), .SE(1'b0), .GCK(pe_1_0_0_net7507) );
  CLKGATETST_X1 pe_1_0_0_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_0_0_n87), .SE(1'b0), .GCK(pe_1_0_0_net7512) );
  CLKGATETST_X1 pe_1_0_0_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_0_0_n86), .SE(1'b0), .GCK(pe_1_0_0_net7517) );
  CLKGATETST_X1 pe_1_0_0_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_0_0_N64), .SE(1'b0), .GCK(pe_1_0_0_net7522) );
  CLKGATETST_X1 pe_1_0_0_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_0_0_N63), .SE(1'b0), .GCK(pe_1_0_0_net7527) );
  CLKGATETST_X1 pe_1_0_0_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_0_0_N62), .SE(1'b0), .GCK(pe_1_0_0_net7532) );
  CLKGATETST_X1 pe_1_0_0_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_0_0_N61), .SE(1'b0), .GCK(pe_1_0_0_net7537) );
  CLKGATETST_X1 pe_1_0_0_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_0_0_N60), .SE(1'b0), .GCK(pe_1_0_0_net7542) );
  CLKGATETST_X1 pe_1_0_0_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_0_0_N59), .SE(1'b0), .GCK(pe_1_0_0_net7547) );
  CLKGATETST_X1 pe_1_0_0_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_0_0_N90), .SE(1'b0), .GCK(pe_1_0_0_net7552) );
  CLKBUF_X1 pe_1_0_1_U108 ( .A(pe_1_0_1_n68), .Z(pe_1_0_1_n67) );
  INV_X1 pe_1_0_1_U107 ( .A(n73), .ZN(pe_1_0_1_n66) );
  INV_X1 pe_1_0_1_U106 ( .A(n65), .ZN(pe_1_0_1_n65) );
  INV_X1 pe_1_0_1_U105 ( .A(n65), .ZN(pe_1_0_1_n64) );
  INV_X1 pe_1_0_1_U104 ( .A(pe_1_0_1_n65), .ZN(pe_1_0_1_n63) );
  INV_X1 pe_1_0_1_U103 ( .A(n25), .ZN(pe_1_0_1_n58) );
  INV_X1 pe_1_0_1_U102 ( .A(n17), .ZN(pe_1_0_1_n57) );
  MUX2_X1 pe_1_0_1_U101 ( .A(pe_1_0_1_n54), .B(pe_1_0_1_n51), .S(n43), .Z(
        int_data_x_0__1__3_) );
  MUX2_X1 pe_1_0_1_U100 ( .A(pe_1_0_1_n53), .B(pe_1_0_1_n52), .S(n37), .Z(
        pe_1_0_1_n54) );
  MUX2_X1 pe_1_0_1_U99 ( .A(pe_1_0_1_int_q_reg_h[23]), .B(
        pe_1_0_1_int_q_reg_h[19]), .S(pe_1_0_1_n56), .Z(pe_1_0_1_n53) );
  MUX2_X1 pe_1_0_1_U98 ( .A(pe_1_0_1_int_q_reg_h[15]), .B(
        pe_1_0_1_int_q_reg_h[11]), .S(pe_1_0_1_n56), .Z(pe_1_0_1_n52) );
  MUX2_X1 pe_1_0_1_U97 ( .A(pe_1_0_1_int_q_reg_h[7]), .B(
        pe_1_0_1_int_q_reg_h[3]), .S(pe_1_0_1_n56), .Z(pe_1_0_1_n51) );
  MUX2_X1 pe_1_0_1_U96 ( .A(pe_1_0_1_n50), .B(pe_1_0_1_n47), .S(n43), .Z(
        int_data_x_0__1__2_) );
  MUX2_X1 pe_1_0_1_U95 ( .A(pe_1_0_1_n49), .B(pe_1_0_1_n48), .S(n37), .Z(
        pe_1_0_1_n50) );
  MUX2_X1 pe_1_0_1_U94 ( .A(pe_1_0_1_int_q_reg_h[22]), .B(
        pe_1_0_1_int_q_reg_h[18]), .S(pe_1_0_1_n56), .Z(pe_1_0_1_n49) );
  MUX2_X1 pe_1_0_1_U93 ( .A(pe_1_0_1_int_q_reg_h[14]), .B(
        pe_1_0_1_int_q_reg_h[10]), .S(pe_1_0_1_n56), .Z(pe_1_0_1_n48) );
  MUX2_X1 pe_1_0_1_U92 ( .A(pe_1_0_1_int_q_reg_h[6]), .B(
        pe_1_0_1_int_q_reg_h[2]), .S(pe_1_0_1_n56), .Z(pe_1_0_1_n47) );
  MUX2_X1 pe_1_0_1_U91 ( .A(pe_1_0_1_n46), .B(pe_1_0_1_n24), .S(n43), .Z(
        int_data_x_0__1__1_) );
  MUX2_X1 pe_1_0_1_U90 ( .A(pe_1_0_1_n45), .B(pe_1_0_1_n25), .S(n37), .Z(
        pe_1_0_1_n46) );
  MUX2_X1 pe_1_0_1_U89 ( .A(pe_1_0_1_int_q_reg_h[21]), .B(
        pe_1_0_1_int_q_reg_h[17]), .S(pe_1_0_1_n56), .Z(pe_1_0_1_n45) );
  MUX2_X1 pe_1_0_1_U88 ( .A(pe_1_0_1_int_q_reg_h[13]), .B(
        pe_1_0_1_int_q_reg_h[9]), .S(pe_1_0_1_n56), .Z(pe_1_0_1_n25) );
  MUX2_X1 pe_1_0_1_U87 ( .A(pe_1_0_1_int_q_reg_h[5]), .B(
        pe_1_0_1_int_q_reg_h[1]), .S(pe_1_0_1_n56), .Z(pe_1_0_1_n24) );
  MUX2_X1 pe_1_0_1_U86 ( .A(pe_1_0_1_n23), .B(pe_1_0_1_n20), .S(n43), .Z(
        int_data_x_0__1__0_) );
  MUX2_X1 pe_1_0_1_U85 ( .A(pe_1_0_1_n22), .B(pe_1_0_1_n21), .S(n37), .Z(
        pe_1_0_1_n23) );
  MUX2_X1 pe_1_0_1_U84 ( .A(pe_1_0_1_int_q_reg_h[20]), .B(
        pe_1_0_1_int_q_reg_h[16]), .S(pe_1_0_1_n56), .Z(pe_1_0_1_n22) );
  MUX2_X1 pe_1_0_1_U83 ( .A(pe_1_0_1_int_q_reg_h[12]), .B(
        pe_1_0_1_int_q_reg_h[8]), .S(pe_1_0_1_n56), .Z(pe_1_0_1_n21) );
  MUX2_X1 pe_1_0_1_U82 ( .A(pe_1_0_1_int_q_reg_h[4]), .B(
        pe_1_0_1_int_q_reg_h[0]), .S(pe_1_0_1_n56), .Z(pe_1_0_1_n20) );
  MUX2_X1 pe_1_0_1_U81 ( .A(pe_1_0_1_n19), .B(pe_1_0_1_n16), .S(n43), .Z(
        pe_1_0_1_o_data_v_3_) );
  MUX2_X1 pe_1_0_1_U80 ( .A(pe_1_0_1_n18), .B(pe_1_0_1_n17), .S(n37), .Z(
        pe_1_0_1_n19) );
  MUX2_X1 pe_1_0_1_U79 ( .A(pe_1_0_1_int_q_reg_v[23]), .B(
        pe_1_0_1_int_q_reg_v[19]), .S(pe_1_0_1_n55), .Z(pe_1_0_1_n18) );
  MUX2_X1 pe_1_0_1_U78 ( .A(pe_1_0_1_int_q_reg_v[15]), .B(
        pe_1_0_1_int_q_reg_v[11]), .S(pe_1_0_1_n55), .Z(pe_1_0_1_n17) );
  MUX2_X1 pe_1_0_1_U77 ( .A(pe_1_0_1_int_q_reg_v[7]), .B(
        pe_1_0_1_int_q_reg_v[3]), .S(pe_1_0_1_n55), .Z(pe_1_0_1_n16) );
  MUX2_X1 pe_1_0_1_U76 ( .A(pe_1_0_1_n15), .B(pe_1_0_1_n12), .S(n43), .Z(
        pe_1_0_1_o_data_v_2_) );
  MUX2_X1 pe_1_0_1_U75 ( .A(pe_1_0_1_n14), .B(pe_1_0_1_n13), .S(n37), .Z(
        pe_1_0_1_n15) );
  MUX2_X1 pe_1_0_1_U74 ( .A(pe_1_0_1_int_q_reg_v[22]), .B(
        pe_1_0_1_int_q_reg_v[18]), .S(pe_1_0_1_n55), .Z(pe_1_0_1_n14) );
  MUX2_X1 pe_1_0_1_U73 ( .A(pe_1_0_1_int_q_reg_v[14]), .B(
        pe_1_0_1_int_q_reg_v[10]), .S(pe_1_0_1_n55), .Z(pe_1_0_1_n13) );
  MUX2_X1 pe_1_0_1_U72 ( .A(pe_1_0_1_int_q_reg_v[6]), .B(
        pe_1_0_1_int_q_reg_v[2]), .S(pe_1_0_1_n55), .Z(pe_1_0_1_n12) );
  MUX2_X1 pe_1_0_1_U71 ( .A(pe_1_0_1_n11), .B(pe_1_0_1_n8), .S(n43), .Z(
        pe_1_0_1_o_data_v_1_) );
  MUX2_X1 pe_1_0_1_U70 ( .A(pe_1_0_1_n10), .B(pe_1_0_1_n9), .S(n37), .Z(
        pe_1_0_1_n11) );
  MUX2_X1 pe_1_0_1_U69 ( .A(pe_1_0_1_int_q_reg_v[21]), .B(
        pe_1_0_1_int_q_reg_v[17]), .S(pe_1_0_1_n55), .Z(pe_1_0_1_n10) );
  MUX2_X1 pe_1_0_1_U68 ( .A(pe_1_0_1_int_q_reg_v[13]), .B(
        pe_1_0_1_int_q_reg_v[9]), .S(pe_1_0_1_n55), .Z(pe_1_0_1_n9) );
  MUX2_X1 pe_1_0_1_U67 ( .A(pe_1_0_1_int_q_reg_v[5]), .B(
        pe_1_0_1_int_q_reg_v[1]), .S(pe_1_0_1_n55), .Z(pe_1_0_1_n8) );
  MUX2_X1 pe_1_0_1_U66 ( .A(pe_1_0_1_n7), .B(pe_1_0_1_n4), .S(n43), .Z(
        pe_1_0_1_o_data_v_0_) );
  MUX2_X1 pe_1_0_1_U65 ( .A(pe_1_0_1_n6), .B(pe_1_0_1_n5), .S(n37), .Z(
        pe_1_0_1_n7) );
  MUX2_X1 pe_1_0_1_U64 ( .A(pe_1_0_1_int_q_reg_v[20]), .B(
        pe_1_0_1_int_q_reg_v[16]), .S(pe_1_0_1_n55), .Z(pe_1_0_1_n6) );
  MUX2_X1 pe_1_0_1_U63 ( .A(pe_1_0_1_int_q_reg_v[12]), .B(
        pe_1_0_1_int_q_reg_v[8]), .S(pe_1_0_1_n55), .Z(pe_1_0_1_n5) );
  MUX2_X1 pe_1_0_1_U62 ( .A(pe_1_0_1_int_q_reg_v[4]), .B(
        pe_1_0_1_int_q_reg_v[0]), .S(pe_1_0_1_n55), .Z(pe_1_0_1_n4) );
  XNOR2_X1 pe_1_0_1_U61 ( .A(pe_1_0_1_n69), .B(o_data[48]), .ZN(pe_1_0_1_N70)
         );
  AOI222_X1 pe_1_0_1_U60 ( .A1(int_data_res_1__1__0_), .A2(pe_1_0_1_n61), .B1(
        pe_1_0_1_n1), .B2(pe_1_0_1_n27), .C1(pe_1_0_1_N70), .C2(pe_1_0_1_n28), 
        .ZN(pe_1_0_1_n35) );
  INV_X1 pe_1_0_1_U59 ( .A(pe_1_0_1_n35), .ZN(pe_1_0_1_n80) );
  AOI222_X1 pe_1_0_1_U58 ( .A1(int_data_res_1__1__2_), .A2(pe_1_0_1_n61), .B1(
        pe_1_0_1_N80), .B2(pe_1_0_1_n27), .C1(pe_1_0_1_N72), .C2(pe_1_0_1_n28), 
        .ZN(pe_1_0_1_n33) );
  INV_X1 pe_1_0_1_U57 ( .A(pe_1_0_1_n33), .ZN(pe_1_0_1_n78) );
  AOI222_X1 pe_1_0_1_U52 ( .A1(int_data_res_1__1__6_), .A2(pe_1_0_1_n61), .B1(
        pe_1_0_1_N84), .B2(pe_1_0_1_n27), .C1(pe_1_0_1_N76), .C2(pe_1_0_1_n28), 
        .ZN(pe_1_0_1_n29) );
  INV_X1 pe_1_0_1_U51 ( .A(pe_1_0_1_n29), .ZN(pe_1_0_1_n74) );
  AOI222_X1 pe_1_0_1_U50 ( .A1(int_data_res_1__1__1_), .A2(pe_1_0_1_n61), .B1(
        pe_1_0_1_N79), .B2(pe_1_0_1_n27), .C1(pe_1_0_1_N71), .C2(pe_1_0_1_n28), 
        .ZN(pe_1_0_1_n34) );
  INV_X1 pe_1_0_1_U49 ( .A(pe_1_0_1_n34), .ZN(pe_1_0_1_n79) );
  AOI222_X1 pe_1_0_1_U48 ( .A1(int_data_res_1__1__3_), .A2(pe_1_0_1_n61), .B1(
        pe_1_0_1_N81), .B2(pe_1_0_1_n27), .C1(pe_1_0_1_N73), .C2(pe_1_0_1_n28), 
        .ZN(pe_1_0_1_n32) );
  INV_X1 pe_1_0_1_U47 ( .A(pe_1_0_1_n32), .ZN(pe_1_0_1_n77) );
  AOI222_X1 pe_1_0_1_U46 ( .A1(int_data_res_1__1__4_), .A2(pe_1_0_1_n61), .B1(
        pe_1_0_1_N82), .B2(pe_1_0_1_n27), .C1(pe_1_0_1_N74), .C2(pe_1_0_1_n28), 
        .ZN(pe_1_0_1_n31) );
  INV_X1 pe_1_0_1_U45 ( .A(pe_1_0_1_n31), .ZN(pe_1_0_1_n76) );
  AOI222_X1 pe_1_0_1_U44 ( .A1(int_data_res_1__1__5_), .A2(pe_1_0_1_n61), .B1(
        pe_1_0_1_N83), .B2(pe_1_0_1_n27), .C1(pe_1_0_1_N75), .C2(pe_1_0_1_n28), 
        .ZN(pe_1_0_1_n30) );
  INV_X1 pe_1_0_1_U43 ( .A(pe_1_0_1_n30), .ZN(pe_1_0_1_n75) );
  INV_X1 pe_1_0_1_U42 ( .A(pe_1_0_1_int_data_2_), .ZN(pe_1_0_1_n71) );
  NAND2_X1 pe_1_0_1_U41 ( .A1(pe_1_0_1_int_data_0_), .A2(pe_1_0_1_n3), .ZN(
        pe_1_0_1_sub_81_carry[1]) );
  INV_X1 pe_1_0_1_U40 ( .A(pe_1_0_1_int_data_1_), .ZN(pe_1_0_1_n70) );
  AND2_X1 pe_1_0_1_U39 ( .A1(pe_1_0_1_int_data_0_), .A2(o_data[48]), .ZN(
        pe_1_0_1_n2) );
  AOI222_X1 pe_1_0_1_U38 ( .A1(pe_1_0_1_n61), .A2(int_data_res_1__1__7_), .B1(
        pe_1_0_1_N85), .B2(pe_1_0_1_n27), .C1(pe_1_0_1_N77), .C2(pe_1_0_1_n28), 
        .ZN(pe_1_0_1_n26) );
  INV_X1 pe_1_0_1_U37 ( .A(pe_1_0_1_n26), .ZN(pe_1_0_1_n73) );
  NOR3_X1 pe_1_0_1_U36 ( .A1(pe_1_0_1_n58), .A2(pe_1_0_1_n62), .A3(int_ckg[62]), .ZN(pe_1_0_1_n36) );
  OR2_X1 pe_1_0_1_U35 ( .A1(pe_1_0_1_n36), .A2(pe_1_0_1_n61), .ZN(pe_1_0_1_N90) );
  INV_X1 pe_1_0_1_U34 ( .A(n37), .ZN(pe_1_0_1_n60) );
  AND2_X1 pe_1_0_1_U33 ( .A1(int_data_x_0__1__2_), .A2(n25), .ZN(
        pe_1_0_1_int_data_2_) );
  AND2_X1 pe_1_0_1_U32 ( .A1(int_data_x_0__1__1_), .A2(n25), .ZN(
        pe_1_0_1_int_data_1_) );
  AND2_X1 pe_1_0_1_U31 ( .A1(int_data_x_0__1__3_), .A2(n25), .ZN(
        pe_1_0_1_int_data_3_) );
  BUF_X1 pe_1_0_1_U30 ( .A(n59), .Z(pe_1_0_1_n61) );
  INV_X1 pe_1_0_1_U29 ( .A(n31), .ZN(pe_1_0_1_n59) );
  AND2_X1 pe_1_0_1_U28 ( .A1(int_data_x_0__1__0_), .A2(n25), .ZN(
        pe_1_0_1_int_data_0_) );
  NAND2_X1 pe_1_0_1_U27 ( .A1(pe_1_0_1_n44), .A2(pe_1_0_1_n59), .ZN(
        pe_1_0_1_n41) );
  AND3_X1 pe_1_0_1_U26 ( .A1(n73), .A2(pe_1_0_1_n60), .A3(n43), .ZN(
        pe_1_0_1_n44) );
  INV_X1 pe_1_0_1_U25 ( .A(pe_1_0_1_int_data_3_), .ZN(pe_1_0_1_n72) );
  NOR2_X1 pe_1_0_1_U24 ( .A1(pe_1_0_1_n66), .A2(n43), .ZN(pe_1_0_1_n43) );
  NOR2_X1 pe_1_0_1_U23 ( .A1(pe_1_0_1_n57), .A2(pe_1_0_1_n61), .ZN(
        pe_1_0_1_n28) );
  NOR2_X1 pe_1_0_1_U22 ( .A1(n17), .A2(pe_1_0_1_n61), .ZN(pe_1_0_1_n27) );
  INV_X1 pe_1_0_1_U21 ( .A(pe_1_0_1_int_data_0_), .ZN(pe_1_0_1_n69) );
  BUF_X1 pe_1_0_1_U20 ( .A(n31), .Z(pe_1_0_1_n55) );
  INV_X1 pe_1_0_1_U19 ( .A(pe_1_0_1_n41), .ZN(pe_1_0_1_n86) );
  INV_X1 pe_1_0_1_U18 ( .A(pe_1_0_1_n37), .ZN(pe_1_0_1_n84) );
  INV_X1 pe_1_0_1_U17 ( .A(pe_1_0_1_n38), .ZN(pe_1_0_1_n83) );
  INV_X1 pe_1_0_1_U16 ( .A(pe_1_0_1_n39), .ZN(pe_1_0_1_n82) );
  NOR2_X1 pe_1_0_1_U15 ( .A1(pe_1_0_1_n64), .A2(pe_1_0_1_n42), .ZN(
        pe_1_0_1_N59) );
  NOR2_X1 pe_1_0_1_U14 ( .A1(pe_1_0_1_n64), .A2(pe_1_0_1_n41), .ZN(
        pe_1_0_1_N60) );
  NOR2_X1 pe_1_0_1_U13 ( .A1(pe_1_0_1_n64), .A2(pe_1_0_1_n38), .ZN(
        pe_1_0_1_N63) );
  NOR2_X1 pe_1_0_1_U12 ( .A1(pe_1_0_1_n64), .A2(pe_1_0_1_n40), .ZN(
        pe_1_0_1_N61) );
  NOR2_X1 pe_1_0_1_U11 ( .A1(pe_1_0_1_n64), .A2(pe_1_0_1_n39), .ZN(
        pe_1_0_1_N62) );
  NOR2_X1 pe_1_0_1_U10 ( .A1(pe_1_0_1_n37), .A2(pe_1_0_1_n64), .ZN(
        pe_1_0_1_N64) );
  NAND2_X1 pe_1_0_1_U9 ( .A1(pe_1_0_1_n44), .A2(n31), .ZN(pe_1_0_1_n42) );
  INV_X1 pe_1_0_1_U8 ( .A(pe_1_0_1_n65), .ZN(pe_1_0_1_n62) );
  BUF_X1 pe_1_0_1_U7 ( .A(n31), .Z(pe_1_0_1_n56) );
  INV_X1 pe_1_0_1_U6 ( .A(pe_1_0_1_n42), .ZN(pe_1_0_1_n85) );
  INV_X1 pe_1_0_1_U5 ( .A(pe_1_0_1_n40), .ZN(pe_1_0_1_n81) );
  INV_X2 pe_1_0_1_U4 ( .A(n81), .ZN(pe_1_0_1_n68) );
  XOR2_X1 pe_1_0_1_U3 ( .A(pe_1_0_1_int_data_0_), .B(o_data[48]), .Z(
        pe_1_0_1_n1) );
  DFFR_X1 pe_1_0_1_int_q_acc_reg_0_ ( .D(pe_1_0_1_n80), .CK(pe_1_0_1_net7474), 
        .RN(pe_1_0_1_n68), .Q(o_data[48]), .QN(pe_1_0_1_n3) );
  DFFR_X1 pe_1_0_1_int_q_reg_v_reg_0__0_ ( .D(int_data_y_1__1__0_), .CK(
        pe_1_0_1_net7444), .RN(pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_v[20]) );
  DFFR_X1 pe_1_0_1_int_q_reg_v_reg_0__1_ ( .D(int_data_y_1__1__1_), .CK(
        pe_1_0_1_net7444), .RN(pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_v[21]) );
  DFFR_X1 pe_1_0_1_int_q_reg_v_reg_0__2_ ( .D(int_data_y_1__1__2_), .CK(
        pe_1_0_1_net7444), .RN(pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_v[22]) );
  DFFR_X1 pe_1_0_1_int_q_reg_v_reg_0__3_ ( .D(int_data_y_1__1__3_), .CK(
        pe_1_0_1_net7444), .RN(pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_v[23]) );
  DFFR_X1 pe_1_0_1_int_q_reg_v_reg_1__0_ ( .D(int_data_y_1__1__0_), .CK(
        pe_1_0_1_net7449), .RN(pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_v[16]) );
  DFFR_X1 pe_1_0_1_int_q_reg_v_reg_1__1_ ( .D(int_data_y_1__1__1_), .CK(
        pe_1_0_1_net7449), .RN(pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_v[17]) );
  DFFR_X1 pe_1_0_1_int_q_reg_v_reg_1__2_ ( .D(int_data_y_1__1__2_), .CK(
        pe_1_0_1_net7449), .RN(pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_v[18]) );
  DFFR_X1 pe_1_0_1_int_q_reg_v_reg_1__3_ ( .D(int_data_y_1__1__3_), .CK(
        pe_1_0_1_net7449), .RN(pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_v[19]) );
  DFFR_X1 pe_1_0_1_int_q_reg_v_reg_2__0_ ( .D(int_data_y_1__1__0_), .CK(
        pe_1_0_1_net7454), .RN(pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_v[12]) );
  DFFR_X1 pe_1_0_1_int_q_reg_v_reg_2__1_ ( .D(int_data_y_1__1__1_), .CK(
        pe_1_0_1_net7454), .RN(pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_v[13]) );
  DFFR_X1 pe_1_0_1_int_q_reg_v_reg_2__2_ ( .D(int_data_y_1__1__2_), .CK(
        pe_1_0_1_net7454), .RN(pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_v[14]) );
  DFFR_X1 pe_1_0_1_int_q_reg_v_reg_2__3_ ( .D(int_data_y_1__1__3_), .CK(
        pe_1_0_1_net7454), .RN(pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_v[15]) );
  DFFR_X1 pe_1_0_1_int_q_reg_v_reg_3__0_ ( .D(int_data_y_1__1__0_), .CK(
        pe_1_0_1_net7459), .RN(pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_v[8]) );
  DFFR_X1 pe_1_0_1_int_q_reg_v_reg_3__1_ ( .D(int_data_y_1__1__1_), .CK(
        pe_1_0_1_net7459), .RN(pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_v[9]) );
  DFFR_X1 pe_1_0_1_int_q_reg_v_reg_3__2_ ( .D(int_data_y_1__1__2_), .CK(
        pe_1_0_1_net7459), .RN(pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_v[10]) );
  DFFR_X1 pe_1_0_1_int_q_reg_v_reg_3__3_ ( .D(int_data_y_1__1__3_), .CK(
        pe_1_0_1_net7459), .RN(pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_v[11]) );
  DFFR_X1 pe_1_0_1_int_q_reg_v_reg_4__0_ ( .D(int_data_y_1__1__0_), .CK(
        pe_1_0_1_net7464), .RN(pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_v[4]) );
  DFFR_X1 pe_1_0_1_int_q_reg_v_reg_4__1_ ( .D(int_data_y_1__1__1_), .CK(
        pe_1_0_1_net7464), .RN(pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_v[5]) );
  DFFR_X1 pe_1_0_1_int_q_reg_v_reg_4__2_ ( .D(int_data_y_1__1__2_), .CK(
        pe_1_0_1_net7464), .RN(pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_v[6]) );
  DFFR_X1 pe_1_0_1_int_q_reg_v_reg_4__3_ ( .D(int_data_y_1__1__3_), .CK(
        pe_1_0_1_net7464), .RN(pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_v[7]) );
  DFFR_X1 pe_1_0_1_int_q_reg_v_reg_5__0_ ( .D(int_data_y_1__1__0_), .CK(
        pe_1_0_1_net7469), .RN(pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_v[0]) );
  DFFR_X1 pe_1_0_1_int_q_reg_v_reg_5__1_ ( .D(int_data_y_1__1__1_), .CK(
        pe_1_0_1_net7469), .RN(pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_v[1]) );
  DFFR_X1 pe_1_0_1_int_q_reg_v_reg_5__2_ ( .D(int_data_y_1__1__2_), .CK(
        pe_1_0_1_net7469), .RN(pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_v[2]) );
  DFFR_X1 pe_1_0_1_int_q_reg_v_reg_5__3_ ( .D(int_data_y_1__1__3_), .CK(
        pe_1_0_1_net7469), .RN(pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_0_1_int_q_reg_h_reg_0__0_ ( .D(int_data_x_0__2__0_), .SI(
        int_data_y_1__1__0_), .SE(pe_1_0_1_n62), .CK(pe_1_0_1_net7413), .RN(
        pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_0_1_int_q_reg_h_reg_0__1_ ( .D(int_data_x_0__2__1_), .SI(
        int_data_y_1__1__1_), .SE(pe_1_0_1_n62), .CK(pe_1_0_1_net7413), .RN(
        pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_0_1_int_q_reg_h_reg_0__2_ ( .D(int_data_x_0__2__2_), .SI(
        int_data_y_1__1__2_), .SE(pe_1_0_1_n62), .CK(pe_1_0_1_net7413), .RN(
        pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_0_1_int_q_reg_h_reg_0__3_ ( .D(int_data_x_0__2__3_), .SI(
        int_data_y_1__1__3_), .SE(pe_1_0_1_n62), .CK(pe_1_0_1_net7413), .RN(
        pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_0_1_int_q_reg_h_reg_1__0_ ( .D(int_data_x_0__2__0_), .SI(
        int_data_y_1__1__0_), .SE(pe_1_0_1_n62), .CK(pe_1_0_1_net7419), .RN(
        pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_0_1_int_q_reg_h_reg_1__1_ ( .D(int_data_x_0__2__1_), .SI(
        int_data_y_1__1__1_), .SE(pe_1_0_1_n62), .CK(pe_1_0_1_net7419), .RN(
        pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_0_1_int_q_reg_h_reg_1__2_ ( .D(int_data_x_0__2__2_), .SI(
        int_data_y_1__1__2_), .SE(pe_1_0_1_n62), .CK(pe_1_0_1_net7419), .RN(
        pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_0_1_int_q_reg_h_reg_1__3_ ( .D(int_data_x_0__2__3_), .SI(
        int_data_y_1__1__3_), .SE(pe_1_0_1_n62), .CK(pe_1_0_1_net7419), .RN(
        pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_0_1_int_q_reg_h_reg_2__0_ ( .D(int_data_x_0__2__0_), .SI(
        int_data_y_1__1__0_), .SE(pe_1_0_1_n62), .CK(pe_1_0_1_net7424), .RN(
        pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_0_1_int_q_reg_h_reg_2__1_ ( .D(int_data_x_0__2__1_), .SI(
        int_data_y_1__1__1_), .SE(pe_1_0_1_n62), .CK(pe_1_0_1_net7424), .RN(
        pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_0_1_int_q_reg_h_reg_2__2_ ( .D(int_data_x_0__2__2_), .SI(
        int_data_y_1__1__2_), .SE(pe_1_0_1_n62), .CK(pe_1_0_1_net7424), .RN(
        pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_0_1_int_q_reg_h_reg_2__3_ ( .D(int_data_x_0__2__3_), .SI(
        int_data_y_1__1__3_), .SE(pe_1_0_1_n62), .CK(pe_1_0_1_net7424), .RN(
        pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_0_1_int_q_reg_h_reg_3__0_ ( .D(int_data_x_0__2__0_), .SI(
        int_data_y_1__1__0_), .SE(pe_1_0_1_n62), .CK(pe_1_0_1_net7429), .RN(
        pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_0_1_int_q_reg_h_reg_3__1_ ( .D(int_data_x_0__2__1_), .SI(
        int_data_y_1__1__1_), .SE(pe_1_0_1_n62), .CK(pe_1_0_1_net7429), .RN(
        pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_0_1_int_q_reg_h_reg_3__2_ ( .D(int_data_x_0__2__2_), .SI(
        int_data_y_1__1__2_), .SE(pe_1_0_1_n62), .CK(pe_1_0_1_net7429), .RN(
        pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_0_1_int_q_reg_h_reg_3__3_ ( .D(int_data_x_0__2__3_), .SI(
        int_data_y_1__1__3_), .SE(pe_1_0_1_n62), .CK(pe_1_0_1_net7429), .RN(
        pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_0_1_int_q_reg_h_reg_4__0_ ( .D(int_data_x_0__2__0_), .SI(
        int_data_y_1__1__0_), .SE(pe_1_0_1_n63), .CK(pe_1_0_1_net7434), .RN(
        pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_0_1_int_q_reg_h_reg_4__1_ ( .D(int_data_x_0__2__1_), .SI(
        int_data_y_1__1__1_), .SE(pe_1_0_1_n63), .CK(pe_1_0_1_net7434), .RN(
        pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_0_1_int_q_reg_h_reg_4__2_ ( .D(int_data_x_0__2__2_), .SI(
        int_data_y_1__1__2_), .SE(pe_1_0_1_n63), .CK(pe_1_0_1_net7434), .RN(
        pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_0_1_int_q_reg_h_reg_4__3_ ( .D(int_data_x_0__2__3_), .SI(
        int_data_y_1__1__3_), .SE(pe_1_0_1_n63), .CK(pe_1_0_1_net7434), .RN(
        pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_0_1_int_q_reg_h_reg_5__0_ ( .D(int_data_x_0__2__0_), .SI(
        int_data_y_1__1__0_), .SE(pe_1_0_1_n63), .CK(pe_1_0_1_net7439), .RN(
        pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_0_1_int_q_reg_h_reg_5__1_ ( .D(int_data_x_0__2__1_), .SI(
        int_data_y_1__1__1_), .SE(pe_1_0_1_n63), .CK(pe_1_0_1_net7439), .RN(
        pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_0_1_int_q_reg_h_reg_5__2_ ( .D(int_data_x_0__2__2_), .SI(
        int_data_y_1__1__2_), .SE(pe_1_0_1_n63), .CK(pe_1_0_1_net7439), .RN(
        pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_0_1_int_q_reg_h_reg_5__3_ ( .D(int_data_x_0__2__3_), .SI(
        int_data_y_1__1__3_), .SE(pe_1_0_1_n63), .CK(pe_1_0_1_net7439), .RN(
        pe_1_0_1_n68), .Q(pe_1_0_1_int_q_reg_h[3]) );
  FA_X1 pe_1_0_1_sub_81_U2_7 ( .A(o_data[55]), .B(pe_1_0_1_n72), .CI(
        pe_1_0_1_sub_81_carry[7]), .S(pe_1_0_1_N77) );
  FA_X1 pe_1_0_1_sub_81_U2_6 ( .A(o_data[54]), .B(pe_1_0_1_n72), .CI(
        pe_1_0_1_sub_81_carry[6]), .CO(pe_1_0_1_sub_81_carry[7]), .S(
        pe_1_0_1_N76) );
  FA_X1 pe_1_0_1_sub_81_U2_5 ( .A(o_data[53]), .B(pe_1_0_1_n72), .CI(
        pe_1_0_1_sub_81_carry[5]), .CO(pe_1_0_1_sub_81_carry[6]), .S(
        pe_1_0_1_N75) );
  FA_X1 pe_1_0_1_sub_81_U2_4 ( .A(o_data[52]), .B(pe_1_0_1_n72), .CI(
        pe_1_0_1_sub_81_carry[4]), .CO(pe_1_0_1_sub_81_carry[5]), .S(
        pe_1_0_1_N74) );
  FA_X1 pe_1_0_1_sub_81_U2_3 ( .A(o_data[51]), .B(pe_1_0_1_n72), .CI(
        pe_1_0_1_sub_81_carry[3]), .CO(pe_1_0_1_sub_81_carry[4]), .S(
        pe_1_0_1_N73) );
  FA_X1 pe_1_0_1_sub_81_U2_2 ( .A(o_data[50]), .B(pe_1_0_1_n71), .CI(
        pe_1_0_1_sub_81_carry[2]), .CO(pe_1_0_1_sub_81_carry[3]), .S(
        pe_1_0_1_N72) );
  FA_X1 pe_1_0_1_sub_81_U2_1 ( .A(o_data[49]), .B(pe_1_0_1_n70), .CI(
        pe_1_0_1_sub_81_carry[1]), .CO(pe_1_0_1_sub_81_carry[2]), .S(
        pe_1_0_1_N71) );
  FA_X1 pe_1_0_1_add_83_U1_7 ( .A(o_data[55]), .B(pe_1_0_1_int_data_3_), .CI(
        pe_1_0_1_add_83_carry[7]), .S(pe_1_0_1_N85) );
  FA_X1 pe_1_0_1_add_83_U1_6 ( .A(o_data[54]), .B(pe_1_0_1_int_data_3_), .CI(
        pe_1_0_1_add_83_carry[6]), .CO(pe_1_0_1_add_83_carry[7]), .S(
        pe_1_0_1_N84) );
  FA_X1 pe_1_0_1_add_83_U1_5 ( .A(o_data[53]), .B(pe_1_0_1_int_data_3_), .CI(
        pe_1_0_1_add_83_carry[5]), .CO(pe_1_0_1_add_83_carry[6]), .S(
        pe_1_0_1_N83) );
  FA_X1 pe_1_0_1_add_83_U1_4 ( .A(o_data[52]), .B(pe_1_0_1_int_data_3_), .CI(
        pe_1_0_1_add_83_carry[4]), .CO(pe_1_0_1_add_83_carry[5]), .S(
        pe_1_0_1_N82) );
  FA_X1 pe_1_0_1_add_83_U1_3 ( .A(o_data[51]), .B(pe_1_0_1_int_data_3_), .CI(
        pe_1_0_1_add_83_carry[3]), .CO(pe_1_0_1_add_83_carry[4]), .S(
        pe_1_0_1_N81) );
  FA_X1 pe_1_0_1_add_83_U1_2 ( .A(o_data[50]), .B(pe_1_0_1_int_data_2_), .CI(
        pe_1_0_1_add_83_carry[2]), .CO(pe_1_0_1_add_83_carry[3]), .S(
        pe_1_0_1_N80) );
  FA_X1 pe_1_0_1_add_83_U1_1 ( .A(o_data[49]), .B(pe_1_0_1_int_data_1_), .CI(
        pe_1_0_1_n2), .CO(pe_1_0_1_add_83_carry[2]), .S(pe_1_0_1_N79) );
  NAND3_X1 pe_1_0_1_U56 ( .A1(n31), .A2(pe_1_0_1_n43), .A3(n37), .ZN(
        pe_1_0_1_n40) );
  NAND3_X1 pe_1_0_1_U55 ( .A1(pe_1_0_1_n43), .A2(pe_1_0_1_n59), .A3(n37), .ZN(
        pe_1_0_1_n39) );
  NAND3_X1 pe_1_0_1_U54 ( .A1(pe_1_0_1_n43), .A2(pe_1_0_1_n60), .A3(n31), .ZN(
        pe_1_0_1_n38) );
  NAND3_X1 pe_1_0_1_U53 ( .A1(pe_1_0_1_n59), .A2(pe_1_0_1_n60), .A3(
        pe_1_0_1_n43), .ZN(pe_1_0_1_n37) );
  DFFR_X1 pe_1_0_1_int_q_acc_reg_6_ ( .D(pe_1_0_1_n74), .CK(pe_1_0_1_net7474), 
        .RN(pe_1_0_1_n67), .Q(o_data[54]) );
  DFFR_X1 pe_1_0_1_int_q_acc_reg_5_ ( .D(pe_1_0_1_n75), .CK(pe_1_0_1_net7474), 
        .RN(pe_1_0_1_n67), .Q(o_data[53]) );
  DFFR_X1 pe_1_0_1_int_q_acc_reg_4_ ( .D(pe_1_0_1_n76), .CK(pe_1_0_1_net7474), 
        .RN(pe_1_0_1_n67), .Q(o_data[52]) );
  DFFR_X1 pe_1_0_1_int_q_acc_reg_3_ ( .D(pe_1_0_1_n77), .CK(pe_1_0_1_net7474), 
        .RN(pe_1_0_1_n67), .Q(o_data[51]) );
  DFFR_X1 pe_1_0_1_int_q_acc_reg_2_ ( .D(pe_1_0_1_n78), .CK(pe_1_0_1_net7474), 
        .RN(pe_1_0_1_n67), .Q(o_data[50]) );
  DFFR_X1 pe_1_0_1_int_q_acc_reg_1_ ( .D(pe_1_0_1_n79), .CK(pe_1_0_1_net7474), 
        .RN(pe_1_0_1_n67), .Q(o_data[49]) );
  DFFR_X1 pe_1_0_1_int_q_acc_reg_7_ ( .D(pe_1_0_1_n73), .CK(pe_1_0_1_net7474), 
        .RN(pe_1_0_1_n67), .Q(o_data[55]) );
  CLKGATETST_X1 pe_1_0_1_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_0_1_n84), .SE(1'b0), .GCK(pe_1_0_1_net7413) );
  CLKGATETST_X1 pe_1_0_1_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_0_1_n83), .SE(1'b0), .GCK(pe_1_0_1_net7419) );
  CLKGATETST_X1 pe_1_0_1_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_0_1_n82), .SE(1'b0), .GCK(pe_1_0_1_net7424) );
  CLKGATETST_X1 pe_1_0_1_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_0_1_n81), .SE(1'b0), .GCK(pe_1_0_1_net7429) );
  CLKGATETST_X1 pe_1_0_1_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_0_1_n86), .SE(1'b0), .GCK(pe_1_0_1_net7434) );
  CLKGATETST_X1 pe_1_0_1_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_0_1_n85), .SE(1'b0), .GCK(pe_1_0_1_net7439) );
  CLKGATETST_X1 pe_1_0_1_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_0_1_N64), .SE(1'b0), .GCK(pe_1_0_1_net7444) );
  CLKGATETST_X1 pe_1_0_1_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_0_1_N63), .SE(1'b0), .GCK(pe_1_0_1_net7449) );
  CLKGATETST_X1 pe_1_0_1_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_0_1_N62), .SE(1'b0), .GCK(pe_1_0_1_net7454) );
  CLKGATETST_X1 pe_1_0_1_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_0_1_N61), .SE(1'b0), .GCK(pe_1_0_1_net7459) );
  CLKGATETST_X1 pe_1_0_1_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_0_1_N60), .SE(1'b0), .GCK(pe_1_0_1_net7464) );
  CLKGATETST_X1 pe_1_0_1_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_0_1_N59), .SE(1'b0), .GCK(pe_1_0_1_net7469) );
  CLKGATETST_X1 pe_1_0_1_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_0_1_N90), .SE(1'b0), .GCK(pe_1_0_1_net7474) );
  CLKBUF_X1 pe_1_0_2_U109 ( .A(pe_1_0_2_n69), .Z(pe_1_0_2_n68) );
  INV_X1 pe_1_0_2_U108 ( .A(n73), .ZN(pe_1_0_2_n67) );
  INV_X1 pe_1_0_2_U107 ( .A(n65), .ZN(pe_1_0_2_n66) );
  INV_X1 pe_1_0_2_U106 ( .A(n65), .ZN(pe_1_0_2_n65) );
  INV_X1 pe_1_0_2_U105 ( .A(pe_1_0_2_n66), .ZN(pe_1_0_2_n64) );
  INV_X1 pe_1_0_2_U104 ( .A(pe_1_0_2_n61), .ZN(pe_1_0_2_n60) );
  INV_X1 pe_1_0_2_U103 ( .A(n25), .ZN(pe_1_0_2_n58) );
  INV_X1 pe_1_0_2_U102 ( .A(n17), .ZN(pe_1_0_2_n57) );
  MUX2_X1 pe_1_0_2_U101 ( .A(pe_1_0_2_n54), .B(pe_1_0_2_n51), .S(n43), .Z(
        int_data_x_0__2__3_) );
  MUX2_X1 pe_1_0_2_U100 ( .A(pe_1_0_2_n53), .B(pe_1_0_2_n52), .S(pe_1_0_2_n60), 
        .Z(pe_1_0_2_n54) );
  MUX2_X1 pe_1_0_2_U99 ( .A(pe_1_0_2_int_q_reg_h[23]), .B(
        pe_1_0_2_int_q_reg_h[19]), .S(pe_1_0_2_n56), .Z(pe_1_0_2_n53) );
  MUX2_X1 pe_1_0_2_U98 ( .A(pe_1_0_2_int_q_reg_h[15]), .B(
        pe_1_0_2_int_q_reg_h[11]), .S(pe_1_0_2_n56), .Z(pe_1_0_2_n52) );
  MUX2_X1 pe_1_0_2_U97 ( .A(pe_1_0_2_int_q_reg_h[7]), .B(
        pe_1_0_2_int_q_reg_h[3]), .S(pe_1_0_2_n56), .Z(pe_1_0_2_n51) );
  MUX2_X1 pe_1_0_2_U96 ( .A(pe_1_0_2_n50), .B(pe_1_0_2_n47), .S(n43), .Z(
        int_data_x_0__2__2_) );
  MUX2_X1 pe_1_0_2_U95 ( .A(pe_1_0_2_n49), .B(pe_1_0_2_n48), .S(pe_1_0_2_n60), 
        .Z(pe_1_0_2_n50) );
  MUX2_X1 pe_1_0_2_U94 ( .A(pe_1_0_2_int_q_reg_h[22]), .B(
        pe_1_0_2_int_q_reg_h[18]), .S(pe_1_0_2_n56), .Z(pe_1_0_2_n49) );
  MUX2_X1 pe_1_0_2_U93 ( .A(pe_1_0_2_int_q_reg_h[14]), .B(
        pe_1_0_2_int_q_reg_h[10]), .S(pe_1_0_2_n56), .Z(pe_1_0_2_n48) );
  MUX2_X1 pe_1_0_2_U92 ( .A(pe_1_0_2_int_q_reg_h[6]), .B(
        pe_1_0_2_int_q_reg_h[2]), .S(pe_1_0_2_n56), .Z(pe_1_0_2_n47) );
  MUX2_X1 pe_1_0_2_U91 ( .A(pe_1_0_2_n46), .B(pe_1_0_2_n24), .S(n43), .Z(
        int_data_x_0__2__1_) );
  MUX2_X1 pe_1_0_2_U90 ( .A(pe_1_0_2_n45), .B(pe_1_0_2_n25), .S(pe_1_0_2_n60), 
        .Z(pe_1_0_2_n46) );
  MUX2_X1 pe_1_0_2_U89 ( .A(pe_1_0_2_int_q_reg_h[21]), .B(
        pe_1_0_2_int_q_reg_h[17]), .S(pe_1_0_2_n56), .Z(pe_1_0_2_n45) );
  MUX2_X1 pe_1_0_2_U88 ( .A(pe_1_0_2_int_q_reg_h[13]), .B(
        pe_1_0_2_int_q_reg_h[9]), .S(pe_1_0_2_n56), .Z(pe_1_0_2_n25) );
  MUX2_X1 pe_1_0_2_U87 ( .A(pe_1_0_2_int_q_reg_h[5]), .B(
        pe_1_0_2_int_q_reg_h[1]), .S(pe_1_0_2_n56), .Z(pe_1_0_2_n24) );
  MUX2_X1 pe_1_0_2_U86 ( .A(pe_1_0_2_n23), .B(pe_1_0_2_n20), .S(n43), .Z(
        int_data_x_0__2__0_) );
  MUX2_X1 pe_1_0_2_U85 ( .A(pe_1_0_2_n22), .B(pe_1_0_2_n21), .S(pe_1_0_2_n60), 
        .Z(pe_1_0_2_n23) );
  MUX2_X1 pe_1_0_2_U84 ( .A(pe_1_0_2_int_q_reg_h[20]), .B(
        pe_1_0_2_int_q_reg_h[16]), .S(pe_1_0_2_n56), .Z(pe_1_0_2_n22) );
  MUX2_X1 pe_1_0_2_U83 ( .A(pe_1_0_2_int_q_reg_h[12]), .B(
        pe_1_0_2_int_q_reg_h[8]), .S(pe_1_0_2_n56), .Z(pe_1_0_2_n21) );
  MUX2_X1 pe_1_0_2_U82 ( .A(pe_1_0_2_int_q_reg_h[4]), .B(
        pe_1_0_2_int_q_reg_h[0]), .S(pe_1_0_2_n56), .Z(pe_1_0_2_n20) );
  MUX2_X1 pe_1_0_2_U81 ( .A(pe_1_0_2_n19), .B(pe_1_0_2_n16), .S(n43), .Z(
        pe_1_0_2_o_data_v_3_) );
  MUX2_X1 pe_1_0_2_U80 ( .A(pe_1_0_2_n18), .B(pe_1_0_2_n17), .S(pe_1_0_2_n60), 
        .Z(pe_1_0_2_n19) );
  MUX2_X1 pe_1_0_2_U79 ( .A(pe_1_0_2_int_q_reg_v[23]), .B(
        pe_1_0_2_int_q_reg_v[19]), .S(pe_1_0_2_n55), .Z(pe_1_0_2_n18) );
  MUX2_X1 pe_1_0_2_U78 ( .A(pe_1_0_2_int_q_reg_v[15]), .B(
        pe_1_0_2_int_q_reg_v[11]), .S(pe_1_0_2_n55), .Z(pe_1_0_2_n17) );
  MUX2_X1 pe_1_0_2_U77 ( .A(pe_1_0_2_int_q_reg_v[7]), .B(
        pe_1_0_2_int_q_reg_v[3]), .S(pe_1_0_2_n55), .Z(pe_1_0_2_n16) );
  MUX2_X1 pe_1_0_2_U76 ( .A(pe_1_0_2_n15), .B(pe_1_0_2_n12), .S(n43), .Z(
        pe_1_0_2_o_data_v_2_) );
  MUX2_X1 pe_1_0_2_U75 ( .A(pe_1_0_2_n14), .B(pe_1_0_2_n13), .S(pe_1_0_2_n60), 
        .Z(pe_1_0_2_n15) );
  MUX2_X1 pe_1_0_2_U74 ( .A(pe_1_0_2_int_q_reg_v[22]), .B(
        pe_1_0_2_int_q_reg_v[18]), .S(pe_1_0_2_n55), .Z(pe_1_0_2_n14) );
  MUX2_X1 pe_1_0_2_U73 ( .A(pe_1_0_2_int_q_reg_v[14]), .B(
        pe_1_0_2_int_q_reg_v[10]), .S(pe_1_0_2_n55), .Z(pe_1_0_2_n13) );
  MUX2_X1 pe_1_0_2_U72 ( .A(pe_1_0_2_int_q_reg_v[6]), .B(
        pe_1_0_2_int_q_reg_v[2]), .S(pe_1_0_2_n55), .Z(pe_1_0_2_n12) );
  MUX2_X1 pe_1_0_2_U71 ( .A(pe_1_0_2_n11), .B(pe_1_0_2_n8), .S(n43), .Z(
        pe_1_0_2_o_data_v_1_) );
  MUX2_X1 pe_1_0_2_U70 ( .A(pe_1_0_2_n10), .B(pe_1_0_2_n9), .S(pe_1_0_2_n60), 
        .Z(pe_1_0_2_n11) );
  MUX2_X1 pe_1_0_2_U69 ( .A(pe_1_0_2_int_q_reg_v[21]), .B(
        pe_1_0_2_int_q_reg_v[17]), .S(pe_1_0_2_n55), .Z(pe_1_0_2_n10) );
  MUX2_X1 pe_1_0_2_U68 ( .A(pe_1_0_2_int_q_reg_v[13]), .B(
        pe_1_0_2_int_q_reg_v[9]), .S(pe_1_0_2_n55), .Z(pe_1_0_2_n9) );
  MUX2_X1 pe_1_0_2_U67 ( .A(pe_1_0_2_int_q_reg_v[5]), .B(
        pe_1_0_2_int_q_reg_v[1]), .S(pe_1_0_2_n55), .Z(pe_1_0_2_n8) );
  MUX2_X1 pe_1_0_2_U66 ( .A(pe_1_0_2_n7), .B(pe_1_0_2_n4), .S(n43), .Z(
        pe_1_0_2_o_data_v_0_) );
  MUX2_X1 pe_1_0_2_U65 ( .A(pe_1_0_2_n6), .B(pe_1_0_2_n5), .S(pe_1_0_2_n60), 
        .Z(pe_1_0_2_n7) );
  MUX2_X1 pe_1_0_2_U64 ( .A(pe_1_0_2_int_q_reg_v[20]), .B(
        pe_1_0_2_int_q_reg_v[16]), .S(pe_1_0_2_n55), .Z(pe_1_0_2_n6) );
  MUX2_X1 pe_1_0_2_U63 ( .A(pe_1_0_2_int_q_reg_v[12]), .B(
        pe_1_0_2_int_q_reg_v[8]), .S(pe_1_0_2_n55), .Z(pe_1_0_2_n5) );
  MUX2_X1 pe_1_0_2_U62 ( .A(pe_1_0_2_int_q_reg_v[4]), .B(
        pe_1_0_2_int_q_reg_v[0]), .S(pe_1_0_2_n55), .Z(pe_1_0_2_n4) );
  XNOR2_X1 pe_1_0_2_U61 ( .A(pe_1_0_2_n70), .B(o_data[40]), .ZN(pe_1_0_2_N70)
         );
  AOI222_X1 pe_1_0_2_U60 ( .A1(int_data_res_1__2__0_), .A2(pe_1_0_2_n62), .B1(
        pe_1_0_2_n1), .B2(pe_1_0_2_n27), .C1(pe_1_0_2_N70), .C2(pe_1_0_2_n28), 
        .ZN(pe_1_0_2_n35) );
  INV_X1 pe_1_0_2_U59 ( .A(pe_1_0_2_n35), .ZN(pe_1_0_2_n81) );
  AOI222_X1 pe_1_0_2_U58 ( .A1(int_data_res_1__2__2_), .A2(pe_1_0_2_n62), .B1(
        pe_1_0_2_N80), .B2(pe_1_0_2_n27), .C1(pe_1_0_2_N72), .C2(pe_1_0_2_n28), 
        .ZN(pe_1_0_2_n33) );
  INV_X1 pe_1_0_2_U57 ( .A(pe_1_0_2_n33), .ZN(pe_1_0_2_n79) );
  AOI222_X1 pe_1_0_2_U52 ( .A1(int_data_res_1__2__6_), .A2(pe_1_0_2_n62), .B1(
        pe_1_0_2_N84), .B2(pe_1_0_2_n27), .C1(pe_1_0_2_N76), .C2(pe_1_0_2_n28), 
        .ZN(pe_1_0_2_n29) );
  INV_X1 pe_1_0_2_U51 ( .A(pe_1_0_2_n29), .ZN(pe_1_0_2_n75) );
  AOI222_X1 pe_1_0_2_U50 ( .A1(int_data_res_1__2__1_), .A2(pe_1_0_2_n62), .B1(
        pe_1_0_2_N79), .B2(pe_1_0_2_n27), .C1(pe_1_0_2_N71), .C2(pe_1_0_2_n28), 
        .ZN(pe_1_0_2_n34) );
  INV_X1 pe_1_0_2_U49 ( .A(pe_1_0_2_n34), .ZN(pe_1_0_2_n80) );
  AOI222_X1 pe_1_0_2_U48 ( .A1(int_data_res_1__2__3_), .A2(pe_1_0_2_n62), .B1(
        pe_1_0_2_N81), .B2(pe_1_0_2_n27), .C1(pe_1_0_2_N73), .C2(pe_1_0_2_n28), 
        .ZN(pe_1_0_2_n32) );
  INV_X1 pe_1_0_2_U47 ( .A(pe_1_0_2_n32), .ZN(pe_1_0_2_n78) );
  AOI222_X1 pe_1_0_2_U46 ( .A1(int_data_res_1__2__4_), .A2(pe_1_0_2_n62), .B1(
        pe_1_0_2_N82), .B2(pe_1_0_2_n27), .C1(pe_1_0_2_N74), .C2(pe_1_0_2_n28), 
        .ZN(pe_1_0_2_n31) );
  INV_X1 pe_1_0_2_U45 ( .A(pe_1_0_2_n31), .ZN(pe_1_0_2_n77) );
  AOI222_X1 pe_1_0_2_U44 ( .A1(int_data_res_1__2__5_), .A2(pe_1_0_2_n62), .B1(
        pe_1_0_2_N83), .B2(pe_1_0_2_n27), .C1(pe_1_0_2_N75), .C2(pe_1_0_2_n28), 
        .ZN(pe_1_0_2_n30) );
  INV_X1 pe_1_0_2_U43 ( .A(pe_1_0_2_n30), .ZN(pe_1_0_2_n76) );
  INV_X1 pe_1_0_2_U42 ( .A(pe_1_0_2_int_data_2_), .ZN(pe_1_0_2_n72) );
  NAND2_X1 pe_1_0_2_U41 ( .A1(pe_1_0_2_int_data_0_), .A2(pe_1_0_2_n3), .ZN(
        pe_1_0_2_sub_81_carry[1]) );
  INV_X1 pe_1_0_2_U40 ( .A(pe_1_0_2_int_data_1_), .ZN(pe_1_0_2_n71) );
  AND2_X1 pe_1_0_2_U39 ( .A1(pe_1_0_2_int_data_0_), .A2(o_data[40]), .ZN(
        pe_1_0_2_n2) );
  AOI222_X1 pe_1_0_2_U38 ( .A1(pe_1_0_2_n62), .A2(int_data_res_1__2__7_), .B1(
        pe_1_0_2_N85), .B2(pe_1_0_2_n27), .C1(pe_1_0_2_N77), .C2(pe_1_0_2_n28), 
        .ZN(pe_1_0_2_n26) );
  INV_X1 pe_1_0_2_U37 ( .A(pe_1_0_2_n26), .ZN(pe_1_0_2_n74) );
  NOR3_X1 pe_1_0_2_U36 ( .A1(pe_1_0_2_n58), .A2(pe_1_0_2_n63), .A3(int_ckg[61]), .ZN(pe_1_0_2_n36) );
  OR2_X1 pe_1_0_2_U35 ( .A1(pe_1_0_2_n36), .A2(pe_1_0_2_n62), .ZN(pe_1_0_2_N90) );
  INV_X1 pe_1_0_2_U34 ( .A(n37), .ZN(pe_1_0_2_n61) );
  AND2_X1 pe_1_0_2_U33 ( .A1(int_data_x_0__2__2_), .A2(n25), .ZN(
        pe_1_0_2_int_data_2_) );
  AND2_X1 pe_1_0_2_U32 ( .A1(int_data_x_0__2__1_), .A2(n25), .ZN(
        pe_1_0_2_int_data_1_) );
  AND2_X1 pe_1_0_2_U31 ( .A1(int_data_x_0__2__3_), .A2(n25), .ZN(
        pe_1_0_2_int_data_3_) );
  BUF_X1 pe_1_0_2_U30 ( .A(n59), .Z(pe_1_0_2_n62) );
  INV_X1 pe_1_0_2_U29 ( .A(n31), .ZN(pe_1_0_2_n59) );
  AND2_X1 pe_1_0_2_U28 ( .A1(int_data_x_0__2__0_), .A2(n25), .ZN(
        pe_1_0_2_int_data_0_) );
  NAND2_X1 pe_1_0_2_U27 ( .A1(pe_1_0_2_n44), .A2(pe_1_0_2_n59), .ZN(
        pe_1_0_2_n41) );
  AND3_X1 pe_1_0_2_U26 ( .A1(n73), .A2(pe_1_0_2_n61), .A3(n43), .ZN(
        pe_1_0_2_n44) );
  INV_X1 pe_1_0_2_U25 ( .A(pe_1_0_2_int_data_3_), .ZN(pe_1_0_2_n73) );
  NOR2_X1 pe_1_0_2_U24 ( .A1(pe_1_0_2_n67), .A2(n43), .ZN(pe_1_0_2_n43) );
  NOR2_X1 pe_1_0_2_U23 ( .A1(pe_1_0_2_n57), .A2(pe_1_0_2_n62), .ZN(
        pe_1_0_2_n28) );
  NOR2_X1 pe_1_0_2_U22 ( .A1(n17), .A2(pe_1_0_2_n62), .ZN(pe_1_0_2_n27) );
  INV_X1 pe_1_0_2_U21 ( .A(pe_1_0_2_int_data_0_), .ZN(pe_1_0_2_n70) );
  BUF_X1 pe_1_0_2_U20 ( .A(n31), .Z(pe_1_0_2_n55) );
  INV_X1 pe_1_0_2_U19 ( .A(pe_1_0_2_n41), .ZN(pe_1_0_2_n87) );
  INV_X1 pe_1_0_2_U18 ( .A(pe_1_0_2_n37), .ZN(pe_1_0_2_n85) );
  INV_X1 pe_1_0_2_U17 ( .A(pe_1_0_2_n38), .ZN(pe_1_0_2_n84) );
  INV_X1 pe_1_0_2_U16 ( .A(pe_1_0_2_n39), .ZN(pe_1_0_2_n83) );
  NOR2_X1 pe_1_0_2_U15 ( .A1(pe_1_0_2_n65), .A2(pe_1_0_2_n42), .ZN(
        pe_1_0_2_N59) );
  NOR2_X1 pe_1_0_2_U14 ( .A1(pe_1_0_2_n65), .A2(pe_1_0_2_n41), .ZN(
        pe_1_0_2_N60) );
  NOR2_X1 pe_1_0_2_U13 ( .A1(pe_1_0_2_n65), .A2(pe_1_0_2_n38), .ZN(
        pe_1_0_2_N63) );
  NOR2_X1 pe_1_0_2_U12 ( .A1(pe_1_0_2_n65), .A2(pe_1_0_2_n40), .ZN(
        pe_1_0_2_N61) );
  NOR2_X1 pe_1_0_2_U11 ( .A1(pe_1_0_2_n65), .A2(pe_1_0_2_n39), .ZN(
        pe_1_0_2_N62) );
  NOR2_X1 pe_1_0_2_U10 ( .A1(pe_1_0_2_n37), .A2(pe_1_0_2_n65), .ZN(
        pe_1_0_2_N64) );
  NAND2_X1 pe_1_0_2_U9 ( .A1(pe_1_0_2_n44), .A2(n31), .ZN(pe_1_0_2_n42) );
  INV_X1 pe_1_0_2_U8 ( .A(pe_1_0_2_n66), .ZN(pe_1_0_2_n63) );
  BUF_X1 pe_1_0_2_U7 ( .A(n31), .Z(pe_1_0_2_n56) );
  INV_X1 pe_1_0_2_U6 ( .A(pe_1_0_2_n42), .ZN(pe_1_0_2_n86) );
  INV_X1 pe_1_0_2_U5 ( .A(pe_1_0_2_n40), .ZN(pe_1_0_2_n82) );
  INV_X2 pe_1_0_2_U4 ( .A(n81), .ZN(pe_1_0_2_n69) );
  XOR2_X1 pe_1_0_2_U3 ( .A(pe_1_0_2_int_data_0_), .B(o_data[40]), .Z(
        pe_1_0_2_n1) );
  DFFR_X1 pe_1_0_2_int_q_acc_reg_0_ ( .D(pe_1_0_2_n81), .CK(pe_1_0_2_net7396), 
        .RN(pe_1_0_2_n69), .Q(o_data[40]), .QN(pe_1_0_2_n3) );
  DFFR_X1 pe_1_0_2_int_q_reg_v_reg_0__0_ ( .D(int_data_y_1__2__0_), .CK(
        pe_1_0_2_net7366), .RN(pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_v[20]) );
  DFFR_X1 pe_1_0_2_int_q_reg_v_reg_0__1_ ( .D(int_data_y_1__2__1_), .CK(
        pe_1_0_2_net7366), .RN(pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_v[21]) );
  DFFR_X1 pe_1_0_2_int_q_reg_v_reg_0__2_ ( .D(int_data_y_1__2__2_), .CK(
        pe_1_0_2_net7366), .RN(pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_v[22]) );
  DFFR_X1 pe_1_0_2_int_q_reg_v_reg_0__3_ ( .D(int_data_y_1__2__3_), .CK(
        pe_1_0_2_net7366), .RN(pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_v[23]) );
  DFFR_X1 pe_1_0_2_int_q_reg_v_reg_1__0_ ( .D(int_data_y_1__2__0_), .CK(
        pe_1_0_2_net7371), .RN(pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_v[16]) );
  DFFR_X1 pe_1_0_2_int_q_reg_v_reg_1__1_ ( .D(int_data_y_1__2__1_), .CK(
        pe_1_0_2_net7371), .RN(pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_v[17]) );
  DFFR_X1 pe_1_0_2_int_q_reg_v_reg_1__2_ ( .D(int_data_y_1__2__2_), .CK(
        pe_1_0_2_net7371), .RN(pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_v[18]) );
  DFFR_X1 pe_1_0_2_int_q_reg_v_reg_1__3_ ( .D(int_data_y_1__2__3_), .CK(
        pe_1_0_2_net7371), .RN(pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_v[19]) );
  DFFR_X1 pe_1_0_2_int_q_reg_v_reg_2__0_ ( .D(int_data_y_1__2__0_), .CK(
        pe_1_0_2_net7376), .RN(pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_v[12]) );
  DFFR_X1 pe_1_0_2_int_q_reg_v_reg_2__1_ ( .D(int_data_y_1__2__1_), .CK(
        pe_1_0_2_net7376), .RN(pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_v[13]) );
  DFFR_X1 pe_1_0_2_int_q_reg_v_reg_2__2_ ( .D(int_data_y_1__2__2_), .CK(
        pe_1_0_2_net7376), .RN(pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_v[14]) );
  DFFR_X1 pe_1_0_2_int_q_reg_v_reg_2__3_ ( .D(int_data_y_1__2__3_), .CK(
        pe_1_0_2_net7376), .RN(pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_v[15]) );
  DFFR_X1 pe_1_0_2_int_q_reg_v_reg_3__0_ ( .D(int_data_y_1__2__0_), .CK(
        pe_1_0_2_net7381), .RN(pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_v[8]) );
  DFFR_X1 pe_1_0_2_int_q_reg_v_reg_3__1_ ( .D(int_data_y_1__2__1_), .CK(
        pe_1_0_2_net7381), .RN(pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_v[9]) );
  DFFR_X1 pe_1_0_2_int_q_reg_v_reg_3__2_ ( .D(int_data_y_1__2__2_), .CK(
        pe_1_0_2_net7381), .RN(pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_v[10]) );
  DFFR_X1 pe_1_0_2_int_q_reg_v_reg_3__3_ ( .D(int_data_y_1__2__3_), .CK(
        pe_1_0_2_net7381), .RN(pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_v[11]) );
  DFFR_X1 pe_1_0_2_int_q_reg_v_reg_4__0_ ( .D(int_data_y_1__2__0_), .CK(
        pe_1_0_2_net7386), .RN(pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_v[4]) );
  DFFR_X1 pe_1_0_2_int_q_reg_v_reg_4__1_ ( .D(int_data_y_1__2__1_), .CK(
        pe_1_0_2_net7386), .RN(pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_v[5]) );
  DFFR_X1 pe_1_0_2_int_q_reg_v_reg_4__2_ ( .D(int_data_y_1__2__2_), .CK(
        pe_1_0_2_net7386), .RN(pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_v[6]) );
  DFFR_X1 pe_1_0_2_int_q_reg_v_reg_4__3_ ( .D(int_data_y_1__2__3_), .CK(
        pe_1_0_2_net7386), .RN(pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_v[7]) );
  DFFR_X1 pe_1_0_2_int_q_reg_v_reg_5__0_ ( .D(int_data_y_1__2__0_), .CK(
        pe_1_0_2_net7391), .RN(pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_v[0]) );
  DFFR_X1 pe_1_0_2_int_q_reg_v_reg_5__1_ ( .D(int_data_y_1__2__1_), .CK(
        pe_1_0_2_net7391), .RN(pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_v[1]) );
  DFFR_X1 pe_1_0_2_int_q_reg_v_reg_5__2_ ( .D(int_data_y_1__2__2_), .CK(
        pe_1_0_2_net7391), .RN(pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_v[2]) );
  DFFR_X1 pe_1_0_2_int_q_reg_v_reg_5__3_ ( .D(int_data_y_1__2__3_), .CK(
        pe_1_0_2_net7391), .RN(pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_0_2_int_q_reg_h_reg_0__0_ ( .D(int_data_x_0__3__0_), .SI(
        int_data_y_1__2__0_), .SE(pe_1_0_2_n63), .CK(pe_1_0_2_net7335), .RN(
        pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_0_2_int_q_reg_h_reg_0__1_ ( .D(int_data_x_0__3__1_), .SI(
        int_data_y_1__2__1_), .SE(pe_1_0_2_n63), .CK(pe_1_0_2_net7335), .RN(
        pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_0_2_int_q_reg_h_reg_0__2_ ( .D(int_data_x_0__3__2_), .SI(
        int_data_y_1__2__2_), .SE(pe_1_0_2_n63), .CK(pe_1_0_2_net7335), .RN(
        pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_0_2_int_q_reg_h_reg_0__3_ ( .D(int_data_x_0__3__3_), .SI(
        int_data_y_1__2__3_), .SE(pe_1_0_2_n63), .CK(pe_1_0_2_net7335), .RN(
        pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_0_2_int_q_reg_h_reg_1__0_ ( .D(int_data_x_0__3__0_), .SI(
        int_data_y_1__2__0_), .SE(pe_1_0_2_n63), .CK(pe_1_0_2_net7341), .RN(
        pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_0_2_int_q_reg_h_reg_1__1_ ( .D(int_data_x_0__3__1_), .SI(
        int_data_y_1__2__1_), .SE(pe_1_0_2_n63), .CK(pe_1_0_2_net7341), .RN(
        pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_0_2_int_q_reg_h_reg_1__2_ ( .D(int_data_x_0__3__2_), .SI(
        int_data_y_1__2__2_), .SE(pe_1_0_2_n63), .CK(pe_1_0_2_net7341), .RN(
        pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_0_2_int_q_reg_h_reg_1__3_ ( .D(int_data_x_0__3__3_), .SI(
        int_data_y_1__2__3_), .SE(pe_1_0_2_n63), .CK(pe_1_0_2_net7341), .RN(
        pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_0_2_int_q_reg_h_reg_2__0_ ( .D(int_data_x_0__3__0_), .SI(
        int_data_y_1__2__0_), .SE(pe_1_0_2_n63), .CK(pe_1_0_2_net7346), .RN(
        pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_0_2_int_q_reg_h_reg_2__1_ ( .D(int_data_x_0__3__1_), .SI(
        int_data_y_1__2__1_), .SE(pe_1_0_2_n63), .CK(pe_1_0_2_net7346), .RN(
        pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_0_2_int_q_reg_h_reg_2__2_ ( .D(int_data_x_0__3__2_), .SI(
        int_data_y_1__2__2_), .SE(pe_1_0_2_n63), .CK(pe_1_0_2_net7346), .RN(
        pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_0_2_int_q_reg_h_reg_2__3_ ( .D(int_data_x_0__3__3_), .SI(
        int_data_y_1__2__3_), .SE(pe_1_0_2_n63), .CK(pe_1_0_2_net7346), .RN(
        pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_0_2_int_q_reg_h_reg_3__0_ ( .D(int_data_x_0__3__0_), .SI(
        int_data_y_1__2__0_), .SE(pe_1_0_2_n63), .CK(pe_1_0_2_net7351), .RN(
        pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_0_2_int_q_reg_h_reg_3__1_ ( .D(int_data_x_0__3__1_), .SI(
        int_data_y_1__2__1_), .SE(pe_1_0_2_n63), .CK(pe_1_0_2_net7351), .RN(
        pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_0_2_int_q_reg_h_reg_3__2_ ( .D(int_data_x_0__3__2_), .SI(
        int_data_y_1__2__2_), .SE(pe_1_0_2_n63), .CK(pe_1_0_2_net7351), .RN(
        pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_0_2_int_q_reg_h_reg_3__3_ ( .D(int_data_x_0__3__3_), .SI(
        int_data_y_1__2__3_), .SE(pe_1_0_2_n63), .CK(pe_1_0_2_net7351), .RN(
        pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_0_2_int_q_reg_h_reg_4__0_ ( .D(int_data_x_0__3__0_), .SI(
        int_data_y_1__2__0_), .SE(pe_1_0_2_n64), .CK(pe_1_0_2_net7356), .RN(
        pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_0_2_int_q_reg_h_reg_4__1_ ( .D(int_data_x_0__3__1_), .SI(
        int_data_y_1__2__1_), .SE(pe_1_0_2_n64), .CK(pe_1_0_2_net7356), .RN(
        pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_0_2_int_q_reg_h_reg_4__2_ ( .D(int_data_x_0__3__2_), .SI(
        int_data_y_1__2__2_), .SE(pe_1_0_2_n64), .CK(pe_1_0_2_net7356), .RN(
        pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_0_2_int_q_reg_h_reg_4__3_ ( .D(int_data_x_0__3__3_), .SI(
        int_data_y_1__2__3_), .SE(pe_1_0_2_n64), .CK(pe_1_0_2_net7356), .RN(
        pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_0_2_int_q_reg_h_reg_5__0_ ( .D(int_data_x_0__3__0_), .SI(
        int_data_y_1__2__0_), .SE(pe_1_0_2_n64), .CK(pe_1_0_2_net7361), .RN(
        pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_0_2_int_q_reg_h_reg_5__1_ ( .D(int_data_x_0__3__1_), .SI(
        int_data_y_1__2__1_), .SE(pe_1_0_2_n64), .CK(pe_1_0_2_net7361), .RN(
        pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_0_2_int_q_reg_h_reg_5__2_ ( .D(int_data_x_0__3__2_), .SI(
        int_data_y_1__2__2_), .SE(pe_1_0_2_n64), .CK(pe_1_0_2_net7361), .RN(
        pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_0_2_int_q_reg_h_reg_5__3_ ( .D(int_data_x_0__3__3_), .SI(
        int_data_y_1__2__3_), .SE(pe_1_0_2_n64), .CK(pe_1_0_2_net7361), .RN(
        pe_1_0_2_n69), .Q(pe_1_0_2_int_q_reg_h[3]) );
  FA_X1 pe_1_0_2_sub_81_U2_7 ( .A(o_data[47]), .B(pe_1_0_2_n73), .CI(
        pe_1_0_2_sub_81_carry[7]), .S(pe_1_0_2_N77) );
  FA_X1 pe_1_0_2_sub_81_U2_6 ( .A(o_data[46]), .B(pe_1_0_2_n73), .CI(
        pe_1_0_2_sub_81_carry[6]), .CO(pe_1_0_2_sub_81_carry[7]), .S(
        pe_1_0_2_N76) );
  FA_X1 pe_1_0_2_sub_81_U2_5 ( .A(o_data[45]), .B(pe_1_0_2_n73), .CI(
        pe_1_0_2_sub_81_carry[5]), .CO(pe_1_0_2_sub_81_carry[6]), .S(
        pe_1_0_2_N75) );
  FA_X1 pe_1_0_2_sub_81_U2_4 ( .A(o_data[44]), .B(pe_1_0_2_n73), .CI(
        pe_1_0_2_sub_81_carry[4]), .CO(pe_1_0_2_sub_81_carry[5]), .S(
        pe_1_0_2_N74) );
  FA_X1 pe_1_0_2_sub_81_U2_3 ( .A(o_data[43]), .B(pe_1_0_2_n73), .CI(
        pe_1_0_2_sub_81_carry[3]), .CO(pe_1_0_2_sub_81_carry[4]), .S(
        pe_1_0_2_N73) );
  FA_X1 pe_1_0_2_sub_81_U2_2 ( .A(o_data[42]), .B(pe_1_0_2_n72), .CI(
        pe_1_0_2_sub_81_carry[2]), .CO(pe_1_0_2_sub_81_carry[3]), .S(
        pe_1_0_2_N72) );
  FA_X1 pe_1_0_2_sub_81_U2_1 ( .A(o_data[41]), .B(pe_1_0_2_n71), .CI(
        pe_1_0_2_sub_81_carry[1]), .CO(pe_1_0_2_sub_81_carry[2]), .S(
        pe_1_0_2_N71) );
  FA_X1 pe_1_0_2_add_83_U1_7 ( .A(o_data[47]), .B(pe_1_0_2_int_data_3_), .CI(
        pe_1_0_2_add_83_carry[7]), .S(pe_1_0_2_N85) );
  FA_X1 pe_1_0_2_add_83_U1_6 ( .A(o_data[46]), .B(pe_1_0_2_int_data_3_), .CI(
        pe_1_0_2_add_83_carry[6]), .CO(pe_1_0_2_add_83_carry[7]), .S(
        pe_1_0_2_N84) );
  FA_X1 pe_1_0_2_add_83_U1_5 ( .A(o_data[45]), .B(pe_1_0_2_int_data_3_), .CI(
        pe_1_0_2_add_83_carry[5]), .CO(pe_1_0_2_add_83_carry[6]), .S(
        pe_1_0_2_N83) );
  FA_X1 pe_1_0_2_add_83_U1_4 ( .A(o_data[44]), .B(pe_1_0_2_int_data_3_), .CI(
        pe_1_0_2_add_83_carry[4]), .CO(pe_1_0_2_add_83_carry[5]), .S(
        pe_1_0_2_N82) );
  FA_X1 pe_1_0_2_add_83_U1_3 ( .A(o_data[43]), .B(pe_1_0_2_int_data_3_), .CI(
        pe_1_0_2_add_83_carry[3]), .CO(pe_1_0_2_add_83_carry[4]), .S(
        pe_1_0_2_N81) );
  FA_X1 pe_1_0_2_add_83_U1_2 ( .A(o_data[42]), .B(pe_1_0_2_int_data_2_), .CI(
        pe_1_0_2_add_83_carry[2]), .CO(pe_1_0_2_add_83_carry[3]), .S(
        pe_1_0_2_N80) );
  FA_X1 pe_1_0_2_add_83_U1_1 ( .A(o_data[41]), .B(pe_1_0_2_int_data_1_), .CI(
        pe_1_0_2_n2), .CO(pe_1_0_2_add_83_carry[2]), .S(pe_1_0_2_N79) );
  NAND3_X1 pe_1_0_2_U56 ( .A1(n31), .A2(pe_1_0_2_n43), .A3(pe_1_0_2_n60), .ZN(
        pe_1_0_2_n40) );
  NAND3_X1 pe_1_0_2_U55 ( .A1(pe_1_0_2_n43), .A2(pe_1_0_2_n59), .A3(
        pe_1_0_2_n60), .ZN(pe_1_0_2_n39) );
  NAND3_X1 pe_1_0_2_U54 ( .A1(pe_1_0_2_n43), .A2(pe_1_0_2_n61), .A3(n31), .ZN(
        pe_1_0_2_n38) );
  NAND3_X1 pe_1_0_2_U53 ( .A1(pe_1_0_2_n59), .A2(pe_1_0_2_n61), .A3(
        pe_1_0_2_n43), .ZN(pe_1_0_2_n37) );
  DFFR_X1 pe_1_0_2_int_q_acc_reg_6_ ( .D(pe_1_0_2_n75), .CK(pe_1_0_2_net7396), 
        .RN(pe_1_0_2_n68), .Q(o_data[46]) );
  DFFR_X1 pe_1_0_2_int_q_acc_reg_5_ ( .D(pe_1_0_2_n76), .CK(pe_1_0_2_net7396), 
        .RN(pe_1_0_2_n68), .Q(o_data[45]) );
  DFFR_X1 pe_1_0_2_int_q_acc_reg_4_ ( .D(pe_1_0_2_n77), .CK(pe_1_0_2_net7396), 
        .RN(pe_1_0_2_n68), .Q(o_data[44]) );
  DFFR_X1 pe_1_0_2_int_q_acc_reg_3_ ( .D(pe_1_0_2_n78), .CK(pe_1_0_2_net7396), 
        .RN(pe_1_0_2_n68), .Q(o_data[43]) );
  DFFR_X1 pe_1_0_2_int_q_acc_reg_2_ ( .D(pe_1_0_2_n79), .CK(pe_1_0_2_net7396), 
        .RN(pe_1_0_2_n68), .Q(o_data[42]) );
  DFFR_X1 pe_1_0_2_int_q_acc_reg_1_ ( .D(pe_1_0_2_n80), .CK(pe_1_0_2_net7396), 
        .RN(pe_1_0_2_n68), .Q(o_data[41]) );
  DFFR_X1 pe_1_0_2_int_q_acc_reg_7_ ( .D(pe_1_0_2_n74), .CK(pe_1_0_2_net7396), 
        .RN(pe_1_0_2_n68), .Q(o_data[47]) );
  CLKGATETST_X1 pe_1_0_2_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_0_2_n85), .SE(1'b0), .GCK(pe_1_0_2_net7335) );
  CLKGATETST_X1 pe_1_0_2_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_0_2_n84), .SE(1'b0), .GCK(pe_1_0_2_net7341) );
  CLKGATETST_X1 pe_1_0_2_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_0_2_n83), .SE(1'b0), .GCK(pe_1_0_2_net7346) );
  CLKGATETST_X1 pe_1_0_2_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_0_2_n82), .SE(1'b0), .GCK(pe_1_0_2_net7351) );
  CLKGATETST_X1 pe_1_0_2_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_0_2_n87), .SE(1'b0), .GCK(pe_1_0_2_net7356) );
  CLKGATETST_X1 pe_1_0_2_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_0_2_n86), .SE(1'b0), .GCK(pe_1_0_2_net7361) );
  CLKGATETST_X1 pe_1_0_2_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_0_2_N64), .SE(1'b0), .GCK(pe_1_0_2_net7366) );
  CLKGATETST_X1 pe_1_0_2_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_0_2_N63), .SE(1'b0), .GCK(pe_1_0_2_net7371) );
  CLKGATETST_X1 pe_1_0_2_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_0_2_N62), .SE(1'b0), .GCK(pe_1_0_2_net7376) );
  CLKGATETST_X1 pe_1_0_2_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_0_2_N61), .SE(1'b0), .GCK(pe_1_0_2_net7381) );
  CLKGATETST_X1 pe_1_0_2_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_0_2_N60), .SE(1'b0), .GCK(pe_1_0_2_net7386) );
  CLKGATETST_X1 pe_1_0_2_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_0_2_N59), .SE(1'b0), .GCK(pe_1_0_2_net7391) );
  CLKGATETST_X1 pe_1_0_2_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_0_2_N90), .SE(1'b0), .GCK(pe_1_0_2_net7396) );
  CLKBUF_X1 pe_1_0_3_U110 ( .A(pe_1_0_3_n70), .Z(pe_1_0_3_n69) );
  INV_X1 pe_1_0_3_U109 ( .A(n73), .ZN(pe_1_0_3_n68) );
  INV_X1 pe_1_0_3_U108 ( .A(n65), .ZN(pe_1_0_3_n67) );
  INV_X1 pe_1_0_3_U107 ( .A(n65), .ZN(pe_1_0_3_n66) );
  INV_X1 pe_1_0_3_U106 ( .A(pe_1_0_3_n67), .ZN(pe_1_0_3_n65) );
  INV_X1 pe_1_0_3_U105 ( .A(pe_1_0_3_n62), .ZN(pe_1_0_3_n61) );
  INV_X1 pe_1_0_3_U104 ( .A(pe_1_0_3_n60), .ZN(pe_1_0_3_n59) );
  INV_X1 pe_1_0_3_U103 ( .A(n25), .ZN(pe_1_0_3_n58) );
  INV_X1 pe_1_0_3_U102 ( .A(n17), .ZN(pe_1_0_3_n57) );
  MUX2_X1 pe_1_0_3_U101 ( .A(pe_1_0_3_n54), .B(pe_1_0_3_n51), .S(n43), .Z(
        int_data_x_0__3__3_) );
  MUX2_X1 pe_1_0_3_U100 ( .A(pe_1_0_3_n53), .B(pe_1_0_3_n52), .S(pe_1_0_3_n61), 
        .Z(pe_1_0_3_n54) );
  MUX2_X1 pe_1_0_3_U99 ( .A(pe_1_0_3_int_q_reg_h[23]), .B(
        pe_1_0_3_int_q_reg_h[19]), .S(pe_1_0_3_n56), .Z(pe_1_0_3_n53) );
  MUX2_X1 pe_1_0_3_U98 ( .A(pe_1_0_3_int_q_reg_h[15]), .B(
        pe_1_0_3_int_q_reg_h[11]), .S(pe_1_0_3_n56), .Z(pe_1_0_3_n52) );
  MUX2_X1 pe_1_0_3_U97 ( .A(pe_1_0_3_int_q_reg_h[7]), .B(
        pe_1_0_3_int_q_reg_h[3]), .S(pe_1_0_3_n56), .Z(pe_1_0_3_n51) );
  MUX2_X1 pe_1_0_3_U96 ( .A(pe_1_0_3_n50), .B(pe_1_0_3_n47), .S(n43), .Z(
        int_data_x_0__3__2_) );
  MUX2_X1 pe_1_0_3_U95 ( .A(pe_1_0_3_n49), .B(pe_1_0_3_n48), .S(pe_1_0_3_n61), 
        .Z(pe_1_0_3_n50) );
  MUX2_X1 pe_1_0_3_U94 ( .A(pe_1_0_3_int_q_reg_h[22]), .B(
        pe_1_0_3_int_q_reg_h[18]), .S(pe_1_0_3_n56), .Z(pe_1_0_3_n49) );
  MUX2_X1 pe_1_0_3_U93 ( .A(pe_1_0_3_int_q_reg_h[14]), .B(
        pe_1_0_3_int_q_reg_h[10]), .S(pe_1_0_3_n56), .Z(pe_1_0_3_n48) );
  MUX2_X1 pe_1_0_3_U92 ( .A(pe_1_0_3_int_q_reg_h[6]), .B(
        pe_1_0_3_int_q_reg_h[2]), .S(pe_1_0_3_n56), .Z(pe_1_0_3_n47) );
  MUX2_X1 pe_1_0_3_U91 ( .A(pe_1_0_3_n46), .B(pe_1_0_3_n24), .S(n43), .Z(
        int_data_x_0__3__1_) );
  MUX2_X1 pe_1_0_3_U90 ( .A(pe_1_0_3_n45), .B(pe_1_0_3_n25), .S(pe_1_0_3_n61), 
        .Z(pe_1_0_3_n46) );
  MUX2_X1 pe_1_0_3_U89 ( .A(pe_1_0_3_int_q_reg_h[21]), .B(
        pe_1_0_3_int_q_reg_h[17]), .S(pe_1_0_3_n56), .Z(pe_1_0_3_n45) );
  MUX2_X1 pe_1_0_3_U88 ( .A(pe_1_0_3_int_q_reg_h[13]), .B(
        pe_1_0_3_int_q_reg_h[9]), .S(pe_1_0_3_n56), .Z(pe_1_0_3_n25) );
  MUX2_X1 pe_1_0_3_U87 ( .A(pe_1_0_3_int_q_reg_h[5]), .B(
        pe_1_0_3_int_q_reg_h[1]), .S(pe_1_0_3_n56), .Z(pe_1_0_3_n24) );
  MUX2_X1 pe_1_0_3_U86 ( .A(pe_1_0_3_n23), .B(pe_1_0_3_n20), .S(n43), .Z(
        int_data_x_0__3__0_) );
  MUX2_X1 pe_1_0_3_U85 ( .A(pe_1_0_3_n22), .B(pe_1_0_3_n21), .S(pe_1_0_3_n61), 
        .Z(pe_1_0_3_n23) );
  MUX2_X1 pe_1_0_3_U84 ( .A(pe_1_0_3_int_q_reg_h[20]), .B(
        pe_1_0_3_int_q_reg_h[16]), .S(pe_1_0_3_n56), .Z(pe_1_0_3_n22) );
  MUX2_X1 pe_1_0_3_U83 ( .A(pe_1_0_3_int_q_reg_h[12]), .B(
        pe_1_0_3_int_q_reg_h[8]), .S(pe_1_0_3_n56), .Z(pe_1_0_3_n21) );
  MUX2_X1 pe_1_0_3_U82 ( .A(pe_1_0_3_int_q_reg_h[4]), .B(
        pe_1_0_3_int_q_reg_h[0]), .S(pe_1_0_3_n56), .Z(pe_1_0_3_n20) );
  MUX2_X1 pe_1_0_3_U81 ( .A(pe_1_0_3_n19), .B(pe_1_0_3_n16), .S(n43), .Z(
        pe_1_0_3_o_data_v_3_) );
  MUX2_X1 pe_1_0_3_U80 ( .A(pe_1_0_3_n18), .B(pe_1_0_3_n17), .S(pe_1_0_3_n61), 
        .Z(pe_1_0_3_n19) );
  MUX2_X1 pe_1_0_3_U79 ( .A(pe_1_0_3_int_q_reg_v[23]), .B(
        pe_1_0_3_int_q_reg_v[19]), .S(pe_1_0_3_n55), .Z(pe_1_0_3_n18) );
  MUX2_X1 pe_1_0_3_U78 ( .A(pe_1_0_3_int_q_reg_v[15]), .B(
        pe_1_0_3_int_q_reg_v[11]), .S(pe_1_0_3_n55), .Z(pe_1_0_3_n17) );
  MUX2_X1 pe_1_0_3_U77 ( .A(pe_1_0_3_int_q_reg_v[7]), .B(
        pe_1_0_3_int_q_reg_v[3]), .S(pe_1_0_3_n55), .Z(pe_1_0_3_n16) );
  MUX2_X1 pe_1_0_3_U76 ( .A(pe_1_0_3_n15), .B(pe_1_0_3_n12), .S(n43), .Z(
        pe_1_0_3_o_data_v_2_) );
  MUX2_X1 pe_1_0_3_U75 ( .A(pe_1_0_3_n14), .B(pe_1_0_3_n13), .S(pe_1_0_3_n61), 
        .Z(pe_1_0_3_n15) );
  MUX2_X1 pe_1_0_3_U74 ( .A(pe_1_0_3_int_q_reg_v[22]), .B(
        pe_1_0_3_int_q_reg_v[18]), .S(pe_1_0_3_n55), .Z(pe_1_0_3_n14) );
  MUX2_X1 pe_1_0_3_U73 ( .A(pe_1_0_3_int_q_reg_v[14]), .B(
        pe_1_0_3_int_q_reg_v[10]), .S(pe_1_0_3_n55), .Z(pe_1_0_3_n13) );
  MUX2_X1 pe_1_0_3_U72 ( .A(pe_1_0_3_int_q_reg_v[6]), .B(
        pe_1_0_3_int_q_reg_v[2]), .S(pe_1_0_3_n55), .Z(pe_1_0_3_n12) );
  MUX2_X1 pe_1_0_3_U71 ( .A(pe_1_0_3_n11), .B(pe_1_0_3_n8), .S(n43), .Z(
        pe_1_0_3_o_data_v_1_) );
  MUX2_X1 pe_1_0_3_U70 ( .A(pe_1_0_3_n10), .B(pe_1_0_3_n9), .S(pe_1_0_3_n61), 
        .Z(pe_1_0_3_n11) );
  MUX2_X1 pe_1_0_3_U69 ( .A(pe_1_0_3_int_q_reg_v[21]), .B(
        pe_1_0_3_int_q_reg_v[17]), .S(pe_1_0_3_n55), .Z(pe_1_0_3_n10) );
  MUX2_X1 pe_1_0_3_U68 ( .A(pe_1_0_3_int_q_reg_v[13]), .B(
        pe_1_0_3_int_q_reg_v[9]), .S(pe_1_0_3_n55), .Z(pe_1_0_3_n9) );
  MUX2_X1 pe_1_0_3_U67 ( .A(pe_1_0_3_int_q_reg_v[5]), .B(
        pe_1_0_3_int_q_reg_v[1]), .S(pe_1_0_3_n55), .Z(pe_1_0_3_n8) );
  MUX2_X1 pe_1_0_3_U66 ( .A(pe_1_0_3_n7), .B(pe_1_0_3_n4), .S(n43), .Z(
        pe_1_0_3_o_data_v_0_) );
  MUX2_X1 pe_1_0_3_U65 ( .A(pe_1_0_3_n6), .B(pe_1_0_3_n5), .S(pe_1_0_3_n61), 
        .Z(pe_1_0_3_n7) );
  MUX2_X1 pe_1_0_3_U64 ( .A(pe_1_0_3_int_q_reg_v[20]), .B(
        pe_1_0_3_int_q_reg_v[16]), .S(pe_1_0_3_n55), .Z(pe_1_0_3_n6) );
  MUX2_X1 pe_1_0_3_U63 ( .A(pe_1_0_3_int_q_reg_v[12]), .B(
        pe_1_0_3_int_q_reg_v[8]), .S(pe_1_0_3_n55), .Z(pe_1_0_3_n5) );
  MUX2_X1 pe_1_0_3_U62 ( .A(pe_1_0_3_int_q_reg_v[4]), .B(
        pe_1_0_3_int_q_reg_v[0]), .S(pe_1_0_3_n55), .Z(pe_1_0_3_n4) );
  XNOR2_X1 pe_1_0_3_U61 ( .A(pe_1_0_3_n71), .B(o_data[32]), .ZN(pe_1_0_3_N70)
         );
  AOI222_X1 pe_1_0_3_U60 ( .A1(int_data_res_1__3__0_), .A2(pe_1_0_3_n63), .B1(
        pe_1_0_3_n1), .B2(pe_1_0_3_n27), .C1(pe_1_0_3_N70), .C2(pe_1_0_3_n28), 
        .ZN(pe_1_0_3_n35) );
  INV_X1 pe_1_0_3_U59 ( .A(pe_1_0_3_n35), .ZN(pe_1_0_3_n82) );
  AOI222_X1 pe_1_0_3_U58 ( .A1(int_data_res_1__3__2_), .A2(pe_1_0_3_n63), .B1(
        pe_1_0_3_N80), .B2(pe_1_0_3_n27), .C1(pe_1_0_3_N72), .C2(pe_1_0_3_n28), 
        .ZN(pe_1_0_3_n33) );
  INV_X1 pe_1_0_3_U57 ( .A(pe_1_0_3_n33), .ZN(pe_1_0_3_n80) );
  AOI222_X1 pe_1_0_3_U52 ( .A1(int_data_res_1__3__6_), .A2(pe_1_0_3_n63), .B1(
        pe_1_0_3_N84), .B2(pe_1_0_3_n27), .C1(pe_1_0_3_N76), .C2(pe_1_0_3_n28), 
        .ZN(pe_1_0_3_n29) );
  INV_X1 pe_1_0_3_U51 ( .A(pe_1_0_3_n29), .ZN(pe_1_0_3_n76) );
  AOI222_X1 pe_1_0_3_U50 ( .A1(int_data_res_1__3__1_), .A2(pe_1_0_3_n63), .B1(
        pe_1_0_3_N79), .B2(pe_1_0_3_n27), .C1(pe_1_0_3_N71), .C2(pe_1_0_3_n28), 
        .ZN(pe_1_0_3_n34) );
  INV_X1 pe_1_0_3_U49 ( .A(pe_1_0_3_n34), .ZN(pe_1_0_3_n81) );
  AOI222_X1 pe_1_0_3_U48 ( .A1(int_data_res_1__3__3_), .A2(pe_1_0_3_n63), .B1(
        pe_1_0_3_N81), .B2(pe_1_0_3_n27), .C1(pe_1_0_3_N73), .C2(pe_1_0_3_n28), 
        .ZN(pe_1_0_3_n32) );
  INV_X1 pe_1_0_3_U47 ( .A(pe_1_0_3_n32), .ZN(pe_1_0_3_n79) );
  AOI222_X1 pe_1_0_3_U46 ( .A1(int_data_res_1__3__4_), .A2(pe_1_0_3_n63), .B1(
        pe_1_0_3_N82), .B2(pe_1_0_3_n27), .C1(pe_1_0_3_N74), .C2(pe_1_0_3_n28), 
        .ZN(pe_1_0_3_n31) );
  INV_X1 pe_1_0_3_U45 ( .A(pe_1_0_3_n31), .ZN(pe_1_0_3_n78) );
  AOI222_X1 pe_1_0_3_U44 ( .A1(int_data_res_1__3__5_), .A2(pe_1_0_3_n63), .B1(
        pe_1_0_3_N83), .B2(pe_1_0_3_n27), .C1(pe_1_0_3_N75), .C2(pe_1_0_3_n28), 
        .ZN(pe_1_0_3_n30) );
  INV_X1 pe_1_0_3_U43 ( .A(pe_1_0_3_n30), .ZN(pe_1_0_3_n77) );
  INV_X1 pe_1_0_3_U42 ( .A(pe_1_0_3_int_data_2_), .ZN(pe_1_0_3_n73) );
  NAND2_X1 pe_1_0_3_U41 ( .A1(pe_1_0_3_int_data_0_), .A2(pe_1_0_3_n3), .ZN(
        pe_1_0_3_sub_81_carry[1]) );
  INV_X1 pe_1_0_3_U40 ( .A(pe_1_0_3_int_data_1_), .ZN(pe_1_0_3_n72) );
  AND2_X1 pe_1_0_3_U39 ( .A1(pe_1_0_3_int_data_0_), .A2(o_data[32]), .ZN(
        pe_1_0_3_n2) );
  AOI222_X1 pe_1_0_3_U38 ( .A1(pe_1_0_3_n63), .A2(int_data_res_1__3__7_), .B1(
        pe_1_0_3_N85), .B2(pe_1_0_3_n27), .C1(pe_1_0_3_N77), .C2(pe_1_0_3_n28), 
        .ZN(pe_1_0_3_n26) );
  INV_X1 pe_1_0_3_U37 ( .A(pe_1_0_3_n26), .ZN(pe_1_0_3_n75) );
  NOR3_X1 pe_1_0_3_U36 ( .A1(pe_1_0_3_n58), .A2(pe_1_0_3_n64), .A3(int_ckg[60]), .ZN(pe_1_0_3_n36) );
  OR2_X1 pe_1_0_3_U35 ( .A1(pe_1_0_3_n36), .A2(pe_1_0_3_n63), .ZN(pe_1_0_3_N90) );
  INV_X1 pe_1_0_3_U34 ( .A(n37), .ZN(pe_1_0_3_n62) );
  AND2_X1 pe_1_0_3_U33 ( .A1(int_data_x_0__3__2_), .A2(n25), .ZN(
        pe_1_0_3_int_data_2_) );
  AND2_X1 pe_1_0_3_U32 ( .A1(int_data_x_0__3__1_), .A2(n25), .ZN(
        pe_1_0_3_int_data_1_) );
  AND2_X1 pe_1_0_3_U31 ( .A1(int_data_x_0__3__3_), .A2(n25), .ZN(
        pe_1_0_3_int_data_3_) );
  BUF_X1 pe_1_0_3_U30 ( .A(n59), .Z(pe_1_0_3_n63) );
  INV_X1 pe_1_0_3_U29 ( .A(n31), .ZN(pe_1_0_3_n60) );
  AND2_X1 pe_1_0_3_U28 ( .A1(int_data_x_0__3__0_), .A2(n25), .ZN(
        pe_1_0_3_int_data_0_) );
  NAND2_X1 pe_1_0_3_U27 ( .A1(pe_1_0_3_n44), .A2(pe_1_0_3_n60), .ZN(
        pe_1_0_3_n41) );
  AND3_X1 pe_1_0_3_U26 ( .A1(n73), .A2(pe_1_0_3_n62), .A3(n43), .ZN(
        pe_1_0_3_n44) );
  INV_X1 pe_1_0_3_U25 ( .A(pe_1_0_3_int_data_3_), .ZN(pe_1_0_3_n74) );
  NOR2_X1 pe_1_0_3_U24 ( .A1(pe_1_0_3_n68), .A2(n43), .ZN(pe_1_0_3_n43) );
  NOR2_X1 pe_1_0_3_U23 ( .A1(pe_1_0_3_n57), .A2(pe_1_0_3_n63), .ZN(
        pe_1_0_3_n28) );
  NOR2_X1 pe_1_0_3_U22 ( .A1(n17), .A2(pe_1_0_3_n63), .ZN(pe_1_0_3_n27) );
  INV_X1 pe_1_0_3_U21 ( .A(pe_1_0_3_int_data_0_), .ZN(pe_1_0_3_n71) );
  BUF_X1 pe_1_0_3_U20 ( .A(pe_1_0_3_n59), .Z(pe_1_0_3_n55) );
  INV_X1 pe_1_0_3_U19 ( .A(pe_1_0_3_n41), .ZN(pe_1_0_3_n88) );
  INV_X1 pe_1_0_3_U18 ( .A(pe_1_0_3_n37), .ZN(pe_1_0_3_n86) );
  INV_X1 pe_1_0_3_U17 ( .A(pe_1_0_3_n38), .ZN(pe_1_0_3_n85) );
  INV_X1 pe_1_0_3_U16 ( .A(pe_1_0_3_n39), .ZN(pe_1_0_3_n84) );
  NOR2_X1 pe_1_0_3_U15 ( .A1(pe_1_0_3_n66), .A2(pe_1_0_3_n42), .ZN(
        pe_1_0_3_N59) );
  NOR2_X1 pe_1_0_3_U14 ( .A1(pe_1_0_3_n66), .A2(pe_1_0_3_n41), .ZN(
        pe_1_0_3_N60) );
  NOR2_X1 pe_1_0_3_U13 ( .A1(pe_1_0_3_n66), .A2(pe_1_0_3_n38), .ZN(
        pe_1_0_3_N63) );
  NOR2_X1 pe_1_0_3_U12 ( .A1(pe_1_0_3_n66), .A2(pe_1_0_3_n40), .ZN(
        pe_1_0_3_N61) );
  NOR2_X1 pe_1_0_3_U11 ( .A1(pe_1_0_3_n66), .A2(pe_1_0_3_n39), .ZN(
        pe_1_0_3_N62) );
  NOR2_X1 pe_1_0_3_U10 ( .A1(pe_1_0_3_n37), .A2(pe_1_0_3_n66), .ZN(
        pe_1_0_3_N64) );
  NAND2_X1 pe_1_0_3_U9 ( .A1(pe_1_0_3_n44), .A2(pe_1_0_3_n59), .ZN(
        pe_1_0_3_n42) );
  INV_X1 pe_1_0_3_U8 ( .A(pe_1_0_3_n67), .ZN(pe_1_0_3_n64) );
  BUF_X1 pe_1_0_3_U7 ( .A(pe_1_0_3_n59), .Z(pe_1_0_3_n56) );
  INV_X1 pe_1_0_3_U6 ( .A(pe_1_0_3_n42), .ZN(pe_1_0_3_n87) );
  INV_X1 pe_1_0_3_U5 ( .A(pe_1_0_3_n40), .ZN(pe_1_0_3_n83) );
  INV_X2 pe_1_0_3_U4 ( .A(n81), .ZN(pe_1_0_3_n70) );
  XOR2_X1 pe_1_0_3_U3 ( .A(pe_1_0_3_int_data_0_), .B(o_data[32]), .Z(
        pe_1_0_3_n1) );
  DFFR_X1 pe_1_0_3_int_q_acc_reg_0_ ( .D(pe_1_0_3_n82), .CK(pe_1_0_3_net7318), 
        .RN(pe_1_0_3_n70), .Q(o_data[32]), .QN(pe_1_0_3_n3) );
  DFFR_X1 pe_1_0_3_int_q_reg_v_reg_0__0_ ( .D(int_data_y_1__3__0_), .CK(
        pe_1_0_3_net7288), .RN(pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_v[20]) );
  DFFR_X1 pe_1_0_3_int_q_reg_v_reg_0__1_ ( .D(int_data_y_1__3__1_), .CK(
        pe_1_0_3_net7288), .RN(pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_v[21]) );
  DFFR_X1 pe_1_0_3_int_q_reg_v_reg_0__2_ ( .D(int_data_y_1__3__2_), .CK(
        pe_1_0_3_net7288), .RN(pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_v[22]) );
  DFFR_X1 pe_1_0_3_int_q_reg_v_reg_0__3_ ( .D(int_data_y_1__3__3_), .CK(
        pe_1_0_3_net7288), .RN(pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_v[23]) );
  DFFR_X1 pe_1_0_3_int_q_reg_v_reg_1__0_ ( .D(int_data_y_1__3__0_), .CK(
        pe_1_0_3_net7293), .RN(pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_v[16]) );
  DFFR_X1 pe_1_0_3_int_q_reg_v_reg_1__1_ ( .D(int_data_y_1__3__1_), .CK(
        pe_1_0_3_net7293), .RN(pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_v[17]) );
  DFFR_X1 pe_1_0_3_int_q_reg_v_reg_1__2_ ( .D(int_data_y_1__3__2_), .CK(
        pe_1_0_3_net7293), .RN(pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_v[18]) );
  DFFR_X1 pe_1_0_3_int_q_reg_v_reg_1__3_ ( .D(int_data_y_1__3__3_), .CK(
        pe_1_0_3_net7293), .RN(pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_v[19]) );
  DFFR_X1 pe_1_0_3_int_q_reg_v_reg_2__0_ ( .D(int_data_y_1__3__0_), .CK(
        pe_1_0_3_net7298), .RN(pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_v[12]) );
  DFFR_X1 pe_1_0_3_int_q_reg_v_reg_2__1_ ( .D(int_data_y_1__3__1_), .CK(
        pe_1_0_3_net7298), .RN(pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_v[13]) );
  DFFR_X1 pe_1_0_3_int_q_reg_v_reg_2__2_ ( .D(int_data_y_1__3__2_), .CK(
        pe_1_0_3_net7298), .RN(pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_v[14]) );
  DFFR_X1 pe_1_0_3_int_q_reg_v_reg_2__3_ ( .D(int_data_y_1__3__3_), .CK(
        pe_1_0_3_net7298), .RN(pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_v[15]) );
  DFFR_X1 pe_1_0_3_int_q_reg_v_reg_3__0_ ( .D(int_data_y_1__3__0_), .CK(
        pe_1_0_3_net7303), .RN(pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_v[8]) );
  DFFR_X1 pe_1_0_3_int_q_reg_v_reg_3__1_ ( .D(int_data_y_1__3__1_), .CK(
        pe_1_0_3_net7303), .RN(pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_v[9]) );
  DFFR_X1 pe_1_0_3_int_q_reg_v_reg_3__2_ ( .D(int_data_y_1__3__2_), .CK(
        pe_1_0_3_net7303), .RN(pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_v[10]) );
  DFFR_X1 pe_1_0_3_int_q_reg_v_reg_3__3_ ( .D(int_data_y_1__3__3_), .CK(
        pe_1_0_3_net7303), .RN(pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_v[11]) );
  DFFR_X1 pe_1_0_3_int_q_reg_v_reg_4__0_ ( .D(int_data_y_1__3__0_), .CK(
        pe_1_0_3_net7308), .RN(pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_v[4]) );
  DFFR_X1 pe_1_0_3_int_q_reg_v_reg_4__1_ ( .D(int_data_y_1__3__1_), .CK(
        pe_1_0_3_net7308), .RN(pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_v[5]) );
  DFFR_X1 pe_1_0_3_int_q_reg_v_reg_4__2_ ( .D(int_data_y_1__3__2_), .CK(
        pe_1_0_3_net7308), .RN(pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_v[6]) );
  DFFR_X1 pe_1_0_3_int_q_reg_v_reg_4__3_ ( .D(int_data_y_1__3__3_), .CK(
        pe_1_0_3_net7308), .RN(pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_v[7]) );
  DFFR_X1 pe_1_0_3_int_q_reg_v_reg_5__0_ ( .D(int_data_y_1__3__0_), .CK(
        pe_1_0_3_net7313), .RN(pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_v[0]) );
  DFFR_X1 pe_1_0_3_int_q_reg_v_reg_5__1_ ( .D(int_data_y_1__3__1_), .CK(
        pe_1_0_3_net7313), .RN(pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_v[1]) );
  DFFR_X1 pe_1_0_3_int_q_reg_v_reg_5__2_ ( .D(int_data_y_1__3__2_), .CK(
        pe_1_0_3_net7313), .RN(pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_v[2]) );
  DFFR_X1 pe_1_0_3_int_q_reg_v_reg_5__3_ ( .D(int_data_y_1__3__3_), .CK(
        pe_1_0_3_net7313), .RN(pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_0_3_int_q_reg_h_reg_0__0_ ( .D(int_data_x_0__4__0_), .SI(
        int_data_y_1__3__0_), .SE(pe_1_0_3_n64), .CK(pe_1_0_3_net7257), .RN(
        pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_0_3_int_q_reg_h_reg_0__1_ ( .D(int_data_x_0__4__1_), .SI(
        int_data_y_1__3__1_), .SE(pe_1_0_3_n64), .CK(pe_1_0_3_net7257), .RN(
        pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_0_3_int_q_reg_h_reg_0__2_ ( .D(int_data_x_0__4__2_), .SI(
        int_data_y_1__3__2_), .SE(pe_1_0_3_n64), .CK(pe_1_0_3_net7257), .RN(
        pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_0_3_int_q_reg_h_reg_0__3_ ( .D(int_data_x_0__4__3_), .SI(
        int_data_y_1__3__3_), .SE(pe_1_0_3_n64), .CK(pe_1_0_3_net7257), .RN(
        pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_0_3_int_q_reg_h_reg_1__0_ ( .D(int_data_x_0__4__0_), .SI(
        int_data_y_1__3__0_), .SE(pe_1_0_3_n64), .CK(pe_1_0_3_net7263), .RN(
        pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_0_3_int_q_reg_h_reg_1__1_ ( .D(int_data_x_0__4__1_), .SI(
        int_data_y_1__3__1_), .SE(pe_1_0_3_n64), .CK(pe_1_0_3_net7263), .RN(
        pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_0_3_int_q_reg_h_reg_1__2_ ( .D(int_data_x_0__4__2_), .SI(
        int_data_y_1__3__2_), .SE(pe_1_0_3_n64), .CK(pe_1_0_3_net7263), .RN(
        pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_0_3_int_q_reg_h_reg_1__3_ ( .D(int_data_x_0__4__3_), .SI(
        int_data_y_1__3__3_), .SE(pe_1_0_3_n64), .CK(pe_1_0_3_net7263), .RN(
        pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_0_3_int_q_reg_h_reg_2__0_ ( .D(int_data_x_0__4__0_), .SI(
        int_data_y_1__3__0_), .SE(pe_1_0_3_n64), .CK(pe_1_0_3_net7268), .RN(
        pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_0_3_int_q_reg_h_reg_2__1_ ( .D(int_data_x_0__4__1_), .SI(
        int_data_y_1__3__1_), .SE(pe_1_0_3_n64), .CK(pe_1_0_3_net7268), .RN(
        pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_0_3_int_q_reg_h_reg_2__2_ ( .D(int_data_x_0__4__2_), .SI(
        int_data_y_1__3__2_), .SE(pe_1_0_3_n64), .CK(pe_1_0_3_net7268), .RN(
        pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_0_3_int_q_reg_h_reg_2__3_ ( .D(int_data_x_0__4__3_), .SI(
        int_data_y_1__3__3_), .SE(pe_1_0_3_n64), .CK(pe_1_0_3_net7268), .RN(
        pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_0_3_int_q_reg_h_reg_3__0_ ( .D(int_data_x_0__4__0_), .SI(
        int_data_y_1__3__0_), .SE(pe_1_0_3_n64), .CK(pe_1_0_3_net7273), .RN(
        pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_0_3_int_q_reg_h_reg_3__1_ ( .D(int_data_x_0__4__1_), .SI(
        int_data_y_1__3__1_), .SE(pe_1_0_3_n64), .CK(pe_1_0_3_net7273), .RN(
        pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_0_3_int_q_reg_h_reg_3__2_ ( .D(int_data_x_0__4__2_), .SI(
        int_data_y_1__3__2_), .SE(pe_1_0_3_n64), .CK(pe_1_0_3_net7273), .RN(
        pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_0_3_int_q_reg_h_reg_3__3_ ( .D(int_data_x_0__4__3_), .SI(
        int_data_y_1__3__3_), .SE(pe_1_0_3_n64), .CK(pe_1_0_3_net7273), .RN(
        pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_0_3_int_q_reg_h_reg_4__0_ ( .D(int_data_x_0__4__0_), .SI(
        int_data_y_1__3__0_), .SE(pe_1_0_3_n65), .CK(pe_1_0_3_net7278), .RN(
        pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_0_3_int_q_reg_h_reg_4__1_ ( .D(int_data_x_0__4__1_), .SI(
        int_data_y_1__3__1_), .SE(pe_1_0_3_n65), .CK(pe_1_0_3_net7278), .RN(
        pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_0_3_int_q_reg_h_reg_4__2_ ( .D(int_data_x_0__4__2_), .SI(
        int_data_y_1__3__2_), .SE(pe_1_0_3_n65), .CK(pe_1_0_3_net7278), .RN(
        pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_0_3_int_q_reg_h_reg_4__3_ ( .D(int_data_x_0__4__3_), .SI(
        int_data_y_1__3__3_), .SE(pe_1_0_3_n65), .CK(pe_1_0_3_net7278), .RN(
        pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_0_3_int_q_reg_h_reg_5__0_ ( .D(int_data_x_0__4__0_), .SI(
        int_data_y_1__3__0_), .SE(pe_1_0_3_n65), .CK(pe_1_0_3_net7283), .RN(
        pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_0_3_int_q_reg_h_reg_5__1_ ( .D(int_data_x_0__4__1_), .SI(
        int_data_y_1__3__1_), .SE(pe_1_0_3_n65), .CK(pe_1_0_3_net7283), .RN(
        pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_0_3_int_q_reg_h_reg_5__2_ ( .D(int_data_x_0__4__2_), .SI(
        int_data_y_1__3__2_), .SE(pe_1_0_3_n65), .CK(pe_1_0_3_net7283), .RN(
        pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_0_3_int_q_reg_h_reg_5__3_ ( .D(int_data_x_0__4__3_), .SI(
        int_data_y_1__3__3_), .SE(pe_1_0_3_n65), .CK(pe_1_0_3_net7283), .RN(
        pe_1_0_3_n70), .Q(pe_1_0_3_int_q_reg_h[3]) );
  FA_X1 pe_1_0_3_sub_81_U2_7 ( .A(o_data[39]), .B(pe_1_0_3_n74), .CI(
        pe_1_0_3_sub_81_carry[7]), .S(pe_1_0_3_N77) );
  FA_X1 pe_1_0_3_sub_81_U2_6 ( .A(o_data[38]), .B(pe_1_0_3_n74), .CI(
        pe_1_0_3_sub_81_carry[6]), .CO(pe_1_0_3_sub_81_carry[7]), .S(
        pe_1_0_3_N76) );
  FA_X1 pe_1_0_3_sub_81_U2_5 ( .A(o_data[37]), .B(pe_1_0_3_n74), .CI(
        pe_1_0_3_sub_81_carry[5]), .CO(pe_1_0_3_sub_81_carry[6]), .S(
        pe_1_0_3_N75) );
  FA_X1 pe_1_0_3_sub_81_U2_4 ( .A(o_data[36]), .B(pe_1_0_3_n74), .CI(
        pe_1_0_3_sub_81_carry[4]), .CO(pe_1_0_3_sub_81_carry[5]), .S(
        pe_1_0_3_N74) );
  FA_X1 pe_1_0_3_sub_81_U2_3 ( .A(o_data[35]), .B(pe_1_0_3_n74), .CI(
        pe_1_0_3_sub_81_carry[3]), .CO(pe_1_0_3_sub_81_carry[4]), .S(
        pe_1_0_3_N73) );
  FA_X1 pe_1_0_3_sub_81_U2_2 ( .A(o_data[34]), .B(pe_1_0_3_n73), .CI(
        pe_1_0_3_sub_81_carry[2]), .CO(pe_1_0_3_sub_81_carry[3]), .S(
        pe_1_0_3_N72) );
  FA_X1 pe_1_0_3_sub_81_U2_1 ( .A(o_data[33]), .B(pe_1_0_3_n72), .CI(
        pe_1_0_3_sub_81_carry[1]), .CO(pe_1_0_3_sub_81_carry[2]), .S(
        pe_1_0_3_N71) );
  FA_X1 pe_1_0_3_add_83_U1_7 ( .A(o_data[39]), .B(pe_1_0_3_int_data_3_), .CI(
        pe_1_0_3_add_83_carry[7]), .S(pe_1_0_3_N85) );
  FA_X1 pe_1_0_3_add_83_U1_6 ( .A(o_data[38]), .B(pe_1_0_3_int_data_3_), .CI(
        pe_1_0_3_add_83_carry[6]), .CO(pe_1_0_3_add_83_carry[7]), .S(
        pe_1_0_3_N84) );
  FA_X1 pe_1_0_3_add_83_U1_5 ( .A(o_data[37]), .B(pe_1_0_3_int_data_3_), .CI(
        pe_1_0_3_add_83_carry[5]), .CO(pe_1_0_3_add_83_carry[6]), .S(
        pe_1_0_3_N83) );
  FA_X1 pe_1_0_3_add_83_U1_4 ( .A(o_data[36]), .B(pe_1_0_3_int_data_3_), .CI(
        pe_1_0_3_add_83_carry[4]), .CO(pe_1_0_3_add_83_carry[5]), .S(
        pe_1_0_3_N82) );
  FA_X1 pe_1_0_3_add_83_U1_3 ( .A(o_data[35]), .B(pe_1_0_3_int_data_3_), .CI(
        pe_1_0_3_add_83_carry[3]), .CO(pe_1_0_3_add_83_carry[4]), .S(
        pe_1_0_3_N81) );
  FA_X1 pe_1_0_3_add_83_U1_2 ( .A(o_data[34]), .B(pe_1_0_3_int_data_2_), .CI(
        pe_1_0_3_add_83_carry[2]), .CO(pe_1_0_3_add_83_carry[3]), .S(
        pe_1_0_3_N80) );
  FA_X1 pe_1_0_3_add_83_U1_1 ( .A(o_data[33]), .B(pe_1_0_3_int_data_1_), .CI(
        pe_1_0_3_n2), .CO(pe_1_0_3_add_83_carry[2]), .S(pe_1_0_3_N79) );
  NAND3_X1 pe_1_0_3_U56 ( .A1(pe_1_0_3_n59), .A2(pe_1_0_3_n43), .A3(
        pe_1_0_3_n61), .ZN(pe_1_0_3_n40) );
  NAND3_X1 pe_1_0_3_U55 ( .A1(pe_1_0_3_n43), .A2(pe_1_0_3_n60), .A3(
        pe_1_0_3_n61), .ZN(pe_1_0_3_n39) );
  NAND3_X1 pe_1_0_3_U54 ( .A1(pe_1_0_3_n43), .A2(pe_1_0_3_n62), .A3(
        pe_1_0_3_n59), .ZN(pe_1_0_3_n38) );
  NAND3_X1 pe_1_0_3_U53 ( .A1(pe_1_0_3_n60), .A2(pe_1_0_3_n62), .A3(
        pe_1_0_3_n43), .ZN(pe_1_0_3_n37) );
  DFFR_X1 pe_1_0_3_int_q_acc_reg_6_ ( .D(pe_1_0_3_n76), .CK(pe_1_0_3_net7318), 
        .RN(pe_1_0_3_n69), .Q(o_data[38]) );
  DFFR_X1 pe_1_0_3_int_q_acc_reg_5_ ( .D(pe_1_0_3_n77), .CK(pe_1_0_3_net7318), 
        .RN(pe_1_0_3_n69), .Q(o_data[37]) );
  DFFR_X1 pe_1_0_3_int_q_acc_reg_4_ ( .D(pe_1_0_3_n78), .CK(pe_1_0_3_net7318), 
        .RN(pe_1_0_3_n69), .Q(o_data[36]) );
  DFFR_X1 pe_1_0_3_int_q_acc_reg_3_ ( .D(pe_1_0_3_n79), .CK(pe_1_0_3_net7318), 
        .RN(pe_1_0_3_n69), .Q(o_data[35]) );
  DFFR_X1 pe_1_0_3_int_q_acc_reg_2_ ( .D(pe_1_0_3_n80), .CK(pe_1_0_3_net7318), 
        .RN(pe_1_0_3_n69), .Q(o_data[34]) );
  DFFR_X1 pe_1_0_3_int_q_acc_reg_1_ ( .D(pe_1_0_3_n81), .CK(pe_1_0_3_net7318), 
        .RN(pe_1_0_3_n69), .Q(o_data[33]) );
  DFFR_X1 pe_1_0_3_int_q_acc_reg_7_ ( .D(pe_1_0_3_n75), .CK(pe_1_0_3_net7318), 
        .RN(pe_1_0_3_n69), .Q(o_data[39]) );
  CLKGATETST_X1 pe_1_0_3_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_0_3_n86), .SE(1'b0), .GCK(pe_1_0_3_net7257) );
  CLKGATETST_X1 pe_1_0_3_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_0_3_n85), .SE(1'b0), .GCK(pe_1_0_3_net7263) );
  CLKGATETST_X1 pe_1_0_3_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_0_3_n84), .SE(1'b0), .GCK(pe_1_0_3_net7268) );
  CLKGATETST_X1 pe_1_0_3_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_0_3_n83), .SE(1'b0), .GCK(pe_1_0_3_net7273) );
  CLKGATETST_X1 pe_1_0_3_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_0_3_n88), .SE(1'b0), .GCK(pe_1_0_3_net7278) );
  CLKGATETST_X1 pe_1_0_3_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_0_3_n87), .SE(1'b0), .GCK(pe_1_0_3_net7283) );
  CLKGATETST_X1 pe_1_0_3_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_0_3_N64), .SE(1'b0), .GCK(pe_1_0_3_net7288) );
  CLKGATETST_X1 pe_1_0_3_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_0_3_N63), .SE(1'b0), .GCK(pe_1_0_3_net7293) );
  CLKGATETST_X1 pe_1_0_3_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_0_3_N62), .SE(1'b0), .GCK(pe_1_0_3_net7298) );
  CLKGATETST_X1 pe_1_0_3_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_0_3_N61), .SE(1'b0), .GCK(pe_1_0_3_net7303) );
  CLKGATETST_X1 pe_1_0_3_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_0_3_N60), .SE(1'b0), .GCK(pe_1_0_3_net7308) );
  CLKGATETST_X1 pe_1_0_3_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_0_3_N59), .SE(1'b0), .GCK(pe_1_0_3_net7313) );
  CLKGATETST_X1 pe_1_0_3_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_0_3_N90), .SE(1'b0), .GCK(pe_1_0_3_net7318) );
  CLKBUF_X1 pe_1_0_4_U112 ( .A(pe_1_0_4_n72), .Z(pe_1_0_4_n71) );
  INV_X1 pe_1_0_4_U111 ( .A(n73), .ZN(pe_1_0_4_n70) );
  INV_X1 pe_1_0_4_U110 ( .A(n65), .ZN(pe_1_0_4_n69) );
  INV_X1 pe_1_0_4_U109 ( .A(n65), .ZN(pe_1_0_4_n68) );
  INV_X1 pe_1_0_4_U108 ( .A(n65), .ZN(pe_1_0_4_n67) );
  INV_X1 pe_1_0_4_U107 ( .A(pe_1_0_4_n69), .ZN(pe_1_0_4_n66) );
  INV_X1 pe_1_0_4_U106 ( .A(pe_1_0_4_n63), .ZN(pe_1_0_4_n62) );
  INV_X1 pe_1_0_4_U105 ( .A(pe_1_0_4_n61), .ZN(pe_1_0_4_n60) );
  INV_X1 pe_1_0_4_U104 ( .A(n25), .ZN(pe_1_0_4_n59) );
  INV_X1 pe_1_0_4_U103 ( .A(pe_1_0_4_n59), .ZN(pe_1_0_4_n58) );
  INV_X1 pe_1_0_4_U102 ( .A(n17), .ZN(pe_1_0_4_n57) );
  MUX2_X1 pe_1_0_4_U101 ( .A(pe_1_0_4_n54), .B(pe_1_0_4_n51), .S(n43), .Z(
        int_data_x_0__4__3_) );
  MUX2_X1 pe_1_0_4_U100 ( .A(pe_1_0_4_n53), .B(pe_1_0_4_n52), .S(pe_1_0_4_n62), 
        .Z(pe_1_0_4_n54) );
  MUX2_X1 pe_1_0_4_U99 ( .A(pe_1_0_4_int_q_reg_h[23]), .B(
        pe_1_0_4_int_q_reg_h[19]), .S(pe_1_0_4_n56), .Z(pe_1_0_4_n53) );
  MUX2_X1 pe_1_0_4_U98 ( .A(pe_1_0_4_int_q_reg_h[15]), .B(
        pe_1_0_4_int_q_reg_h[11]), .S(pe_1_0_4_n56), .Z(pe_1_0_4_n52) );
  MUX2_X1 pe_1_0_4_U97 ( .A(pe_1_0_4_int_q_reg_h[7]), .B(
        pe_1_0_4_int_q_reg_h[3]), .S(pe_1_0_4_n56), .Z(pe_1_0_4_n51) );
  MUX2_X1 pe_1_0_4_U96 ( .A(pe_1_0_4_n50), .B(pe_1_0_4_n47), .S(n43), .Z(
        int_data_x_0__4__2_) );
  MUX2_X1 pe_1_0_4_U95 ( .A(pe_1_0_4_n49), .B(pe_1_0_4_n48), .S(pe_1_0_4_n62), 
        .Z(pe_1_0_4_n50) );
  MUX2_X1 pe_1_0_4_U94 ( .A(pe_1_0_4_int_q_reg_h[22]), .B(
        pe_1_0_4_int_q_reg_h[18]), .S(pe_1_0_4_n56), .Z(pe_1_0_4_n49) );
  MUX2_X1 pe_1_0_4_U93 ( .A(pe_1_0_4_int_q_reg_h[14]), .B(
        pe_1_0_4_int_q_reg_h[10]), .S(pe_1_0_4_n56), .Z(pe_1_0_4_n48) );
  MUX2_X1 pe_1_0_4_U92 ( .A(pe_1_0_4_int_q_reg_h[6]), .B(
        pe_1_0_4_int_q_reg_h[2]), .S(pe_1_0_4_n56), .Z(pe_1_0_4_n47) );
  MUX2_X1 pe_1_0_4_U91 ( .A(pe_1_0_4_n46), .B(pe_1_0_4_n24), .S(n43), .Z(
        int_data_x_0__4__1_) );
  MUX2_X1 pe_1_0_4_U90 ( .A(pe_1_0_4_n45), .B(pe_1_0_4_n25), .S(pe_1_0_4_n62), 
        .Z(pe_1_0_4_n46) );
  MUX2_X1 pe_1_0_4_U89 ( .A(pe_1_0_4_int_q_reg_h[21]), .B(
        pe_1_0_4_int_q_reg_h[17]), .S(pe_1_0_4_n56), .Z(pe_1_0_4_n45) );
  MUX2_X1 pe_1_0_4_U88 ( .A(pe_1_0_4_int_q_reg_h[13]), .B(
        pe_1_0_4_int_q_reg_h[9]), .S(pe_1_0_4_n56), .Z(pe_1_0_4_n25) );
  MUX2_X1 pe_1_0_4_U87 ( .A(pe_1_0_4_int_q_reg_h[5]), .B(
        pe_1_0_4_int_q_reg_h[1]), .S(pe_1_0_4_n56), .Z(pe_1_0_4_n24) );
  MUX2_X1 pe_1_0_4_U86 ( .A(pe_1_0_4_n23), .B(pe_1_0_4_n20), .S(n43), .Z(
        int_data_x_0__4__0_) );
  MUX2_X1 pe_1_0_4_U85 ( .A(pe_1_0_4_n22), .B(pe_1_0_4_n21), .S(pe_1_0_4_n62), 
        .Z(pe_1_0_4_n23) );
  MUX2_X1 pe_1_0_4_U84 ( .A(pe_1_0_4_int_q_reg_h[20]), .B(
        pe_1_0_4_int_q_reg_h[16]), .S(pe_1_0_4_n56), .Z(pe_1_0_4_n22) );
  MUX2_X1 pe_1_0_4_U83 ( .A(pe_1_0_4_int_q_reg_h[12]), .B(
        pe_1_0_4_int_q_reg_h[8]), .S(pe_1_0_4_n56), .Z(pe_1_0_4_n21) );
  MUX2_X1 pe_1_0_4_U82 ( .A(pe_1_0_4_int_q_reg_h[4]), .B(
        pe_1_0_4_int_q_reg_h[0]), .S(pe_1_0_4_n56), .Z(pe_1_0_4_n20) );
  MUX2_X1 pe_1_0_4_U81 ( .A(pe_1_0_4_n19), .B(pe_1_0_4_n16), .S(n43), .Z(
        pe_1_0_4_o_data_v_3_) );
  MUX2_X1 pe_1_0_4_U80 ( .A(pe_1_0_4_n18), .B(pe_1_0_4_n17), .S(pe_1_0_4_n62), 
        .Z(pe_1_0_4_n19) );
  MUX2_X1 pe_1_0_4_U79 ( .A(pe_1_0_4_int_q_reg_v[23]), .B(
        pe_1_0_4_int_q_reg_v[19]), .S(pe_1_0_4_n55), .Z(pe_1_0_4_n18) );
  MUX2_X1 pe_1_0_4_U78 ( .A(pe_1_0_4_int_q_reg_v[15]), .B(
        pe_1_0_4_int_q_reg_v[11]), .S(pe_1_0_4_n55), .Z(pe_1_0_4_n17) );
  MUX2_X1 pe_1_0_4_U77 ( .A(pe_1_0_4_int_q_reg_v[7]), .B(
        pe_1_0_4_int_q_reg_v[3]), .S(pe_1_0_4_n55), .Z(pe_1_0_4_n16) );
  MUX2_X1 pe_1_0_4_U76 ( .A(pe_1_0_4_n15), .B(pe_1_0_4_n12), .S(n43), .Z(
        pe_1_0_4_o_data_v_2_) );
  MUX2_X1 pe_1_0_4_U75 ( .A(pe_1_0_4_n14), .B(pe_1_0_4_n13), .S(pe_1_0_4_n62), 
        .Z(pe_1_0_4_n15) );
  MUX2_X1 pe_1_0_4_U74 ( .A(pe_1_0_4_int_q_reg_v[22]), .B(
        pe_1_0_4_int_q_reg_v[18]), .S(pe_1_0_4_n55), .Z(pe_1_0_4_n14) );
  MUX2_X1 pe_1_0_4_U73 ( .A(pe_1_0_4_int_q_reg_v[14]), .B(
        pe_1_0_4_int_q_reg_v[10]), .S(pe_1_0_4_n55), .Z(pe_1_0_4_n13) );
  MUX2_X1 pe_1_0_4_U72 ( .A(pe_1_0_4_int_q_reg_v[6]), .B(
        pe_1_0_4_int_q_reg_v[2]), .S(pe_1_0_4_n55), .Z(pe_1_0_4_n12) );
  MUX2_X1 pe_1_0_4_U71 ( .A(pe_1_0_4_n11), .B(pe_1_0_4_n8), .S(n43), .Z(
        pe_1_0_4_o_data_v_1_) );
  MUX2_X1 pe_1_0_4_U70 ( .A(pe_1_0_4_n10), .B(pe_1_0_4_n9), .S(pe_1_0_4_n62), 
        .Z(pe_1_0_4_n11) );
  MUX2_X1 pe_1_0_4_U69 ( .A(pe_1_0_4_int_q_reg_v[21]), .B(
        pe_1_0_4_int_q_reg_v[17]), .S(pe_1_0_4_n55), .Z(pe_1_0_4_n10) );
  MUX2_X1 pe_1_0_4_U68 ( .A(pe_1_0_4_int_q_reg_v[13]), .B(
        pe_1_0_4_int_q_reg_v[9]), .S(pe_1_0_4_n55), .Z(pe_1_0_4_n9) );
  MUX2_X1 pe_1_0_4_U67 ( .A(pe_1_0_4_int_q_reg_v[5]), .B(
        pe_1_0_4_int_q_reg_v[1]), .S(pe_1_0_4_n55), .Z(pe_1_0_4_n8) );
  MUX2_X1 pe_1_0_4_U66 ( .A(pe_1_0_4_n7), .B(pe_1_0_4_n4), .S(n43), .Z(
        pe_1_0_4_o_data_v_0_) );
  MUX2_X1 pe_1_0_4_U65 ( .A(pe_1_0_4_n6), .B(pe_1_0_4_n5), .S(pe_1_0_4_n62), 
        .Z(pe_1_0_4_n7) );
  MUX2_X1 pe_1_0_4_U64 ( .A(pe_1_0_4_int_q_reg_v[20]), .B(
        pe_1_0_4_int_q_reg_v[16]), .S(pe_1_0_4_n55), .Z(pe_1_0_4_n6) );
  MUX2_X1 pe_1_0_4_U63 ( .A(pe_1_0_4_int_q_reg_v[12]), .B(
        pe_1_0_4_int_q_reg_v[8]), .S(pe_1_0_4_n55), .Z(pe_1_0_4_n5) );
  MUX2_X1 pe_1_0_4_U62 ( .A(pe_1_0_4_int_q_reg_v[4]), .B(
        pe_1_0_4_int_q_reg_v[0]), .S(pe_1_0_4_n55), .Z(pe_1_0_4_n4) );
  XNOR2_X1 pe_1_0_4_U61 ( .A(pe_1_0_4_n73), .B(o_data[24]), .ZN(pe_1_0_4_N70)
         );
  AOI222_X1 pe_1_0_4_U60 ( .A1(int_data_res_1__4__0_), .A2(pe_1_0_4_n64), .B1(
        pe_1_0_4_n1), .B2(pe_1_0_4_n27), .C1(pe_1_0_4_N70), .C2(pe_1_0_4_n28), 
        .ZN(pe_1_0_4_n35) );
  INV_X1 pe_1_0_4_U59 ( .A(pe_1_0_4_n35), .ZN(pe_1_0_4_n84) );
  AOI222_X1 pe_1_0_4_U58 ( .A1(int_data_res_1__4__2_), .A2(pe_1_0_4_n64), .B1(
        pe_1_0_4_N80), .B2(pe_1_0_4_n27), .C1(pe_1_0_4_N72), .C2(pe_1_0_4_n28), 
        .ZN(pe_1_0_4_n33) );
  INV_X1 pe_1_0_4_U57 ( .A(pe_1_0_4_n33), .ZN(pe_1_0_4_n82) );
  AOI222_X1 pe_1_0_4_U52 ( .A1(int_data_res_1__4__6_), .A2(pe_1_0_4_n64), .B1(
        pe_1_0_4_N84), .B2(pe_1_0_4_n27), .C1(pe_1_0_4_N76), .C2(pe_1_0_4_n28), 
        .ZN(pe_1_0_4_n29) );
  INV_X1 pe_1_0_4_U51 ( .A(pe_1_0_4_n29), .ZN(pe_1_0_4_n78) );
  AOI222_X1 pe_1_0_4_U50 ( .A1(int_data_res_1__4__1_), .A2(pe_1_0_4_n64), .B1(
        pe_1_0_4_N79), .B2(pe_1_0_4_n27), .C1(pe_1_0_4_N71), .C2(pe_1_0_4_n28), 
        .ZN(pe_1_0_4_n34) );
  INV_X1 pe_1_0_4_U49 ( .A(pe_1_0_4_n34), .ZN(pe_1_0_4_n83) );
  AOI222_X1 pe_1_0_4_U48 ( .A1(int_data_res_1__4__3_), .A2(pe_1_0_4_n64), .B1(
        pe_1_0_4_N81), .B2(pe_1_0_4_n27), .C1(pe_1_0_4_N73), .C2(pe_1_0_4_n28), 
        .ZN(pe_1_0_4_n32) );
  INV_X1 pe_1_0_4_U47 ( .A(pe_1_0_4_n32), .ZN(pe_1_0_4_n81) );
  AOI222_X1 pe_1_0_4_U46 ( .A1(int_data_res_1__4__4_), .A2(pe_1_0_4_n64), .B1(
        pe_1_0_4_N82), .B2(pe_1_0_4_n27), .C1(pe_1_0_4_N74), .C2(pe_1_0_4_n28), 
        .ZN(pe_1_0_4_n31) );
  INV_X1 pe_1_0_4_U45 ( .A(pe_1_0_4_n31), .ZN(pe_1_0_4_n80) );
  AOI222_X1 pe_1_0_4_U44 ( .A1(int_data_res_1__4__5_), .A2(pe_1_0_4_n64), .B1(
        pe_1_0_4_N83), .B2(pe_1_0_4_n27), .C1(pe_1_0_4_N75), .C2(pe_1_0_4_n28), 
        .ZN(pe_1_0_4_n30) );
  INV_X1 pe_1_0_4_U43 ( .A(pe_1_0_4_n30), .ZN(pe_1_0_4_n79) );
  INV_X1 pe_1_0_4_U42 ( .A(pe_1_0_4_int_data_2_), .ZN(pe_1_0_4_n75) );
  NAND2_X1 pe_1_0_4_U41 ( .A1(pe_1_0_4_int_data_0_), .A2(pe_1_0_4_n3), .ZN(
        pe_1_0_4_sub_81_carry[1]) );
  INV_X1 pe_1_0_4_U40 ( .A(pe_1_0_4_int_data_1_), .ZN(pe_1_0_4_n74) );
  AND2_X1 pe_1_0_4_U39 ( .A1(pe_1_0_4_int_data_0_), .A2(o_data[24]), .ZN(
        pe_1_0_4_n2) );
  AOI222_X1 pe_1_0_4_U38 ( .A1(pe_1_0_4_n64), .A2(int_data_res_1__4__7_), .B1(
        pe_1_0_4_N85), .B2(pe_1_0_4_n27), .C1(pe_1_0_4_N77), .C2(pe_1_0_4_n28), 
        .ZN(pe_1_0_4_n26) );
  INV_X1 pe_1_0_4_U37 ( .A(pe_1_0_4_n26), .ZN(pe_1_0_4_n77) );
  NOR3_X1 pe_1_0_4_U36 ( .A1(pe_1_0_4_n59), .A2(pe_1_0_4_n65), .A3(int_ckg[59]), .ZN(pe_1_0_4_n36) );
  OR2_X1 pe_1_0_4_U35 ( .A1(pe_1_0_4_n36), .A2(pe_1_0_4_n64), .ZN(pe_1_0_4_N90) );
  INV_X1 pe_1_0_4_U34 ( .A(n37), .ZN(pe_1_0_4_n63) );
  AND2_X1 pe_1_0_4_U33 ( .A1(int_data_x_0__4__2_), .A2(pe_1_0_4_n58), .ZN(
        pe_1_0_4_int_data_2_) );
  AND2_X1 pe_1_0_4_U32 ( .A1(int_data_x_0__4__1_), .A2(pe_1_0_4_n58), .ZN(
        pe_1_0_4_int_data_1_) );
  AND2_X1 pe_1_0_4_U31 ( .A1(int_data_x_0__4__3_), .A2(pe_1_0_4_n58), .ZN(
        pe_1_0_4_int_data_3_) );
  BUF_X1 pe_1_0_4_U30 ( .A(n59), .Z(pe_1_0_4_n64) );
  INV_X1 pe_1_0_4_U29 ( .A(n31), .ZN(pe_1_0_4_n61) );
  AND2_X1 pe_1_0_4_U28 ( .A1(int_data_x_0__4__0_), .A2(pe_1_0_4_n58), .ZN(
        pe_1_0_4_int_data_0_) );
  NAND2_X1 pe_1_0_4_U27 ( .A1(pe_1_0_4_n44), .A2(pe_1_0_4_n61), .ZN(
        pe_1_0_4_n41) );
  AND3_X1 pe_1_0_4_U26 ( .A1(n73), .A2(pe_1_0_4_n63), .A3(n43), .ZN(
        pe_1_0_4_n44) );
  INV_X1 pe_1_0_4_U25 ( .A(pe_1_0_4_int_data_3_), .ZN(pe_1_0_4_n76) );
  NOR2_X1 pe_1_0_4_U24 ( .A1(pe_1_0_4_n70), .A2(n43), .ZN(pe_1_0_4_n43) );
  NOR2_X1 pe_1_0_4_U23 ( .A1(pe_1_0_4_n57), .A2(pe_1_0_4_n64), .ZN(
        pe_1_0_4_n28) );
  NOR2_X1 pe_1_0_4_U22 ( .A1(n17), .A2(pe_1_0_4_n64), .ZN(pe_1_0_4_n27) );
  INV_X1 pe_1_0_4_U21 ( .A(pe_1_0_4_int_data_0_), .ZN(pe_1_0_4_n73) );
  BUF_X1 pe_1_0_4_U20 ( .A(pe_1_0_4_n60), .Z(pe_1_0_4_n55) );
  INV_X1 pe_1_0_4_U19 ( .A(pe_1_0_4_n41), .ZN(pe_1_0_4_n90) );
  INV_X1 pe_1_0_4_U18 ( .A(pe_1_0_4_n37), .ZN(pe_1_0_4_n88) );
  INV_X1 pe_1_0_4_U17 ( .A(pe_1_0_4_n38), .ZN(pe_1_0_4_n87) );
  INV_X1 pe_1_0_4_U16 ( .A(pe_1_0_4_n39), .ZN(pe_1_0_4_n86) );
  NOR2_X1 pe_1_0_4_U15 ( .A1(pe_1_0_4_n68), .A2(pe_1_0_4_n42), .ZN(
        pe_1_0_4_N59) );
  NOR2_X1 pe_1_0_4_U14 ( .A1(pe_1_0_4_n68), .A2(pe_1_0_4_n41), .ZN(
        pe_1_0_4_N60) );
  NOR2_X1 pe_1_0_4_U13 ( .A1(pe_1_0_4_n68), .A2(pe_1_0_4_n38), .ZN(
        pe_1_0_4_N63) );
  NOR2_X1 pe_1_0_4_U12 ( .A1(pe_1_0_4_n67), .A2(pe_1_0_4_n40), .ZN(
        pe_1_0_4_N61) );
  NOR2_X1 pe_1_0_4_U11 ( .A1(pe_1_0_4_n67), .A2(pe_1_0_4_n39), .ZN(
        pe_1_0_4_N62) );
  NOR2_X1 pe_1_0_4_U10 ( .A1(pe_1_0_4_n37), .A2(pe_1_0_4_n67), .ZN(
        pe_1_0_4_N64) );
  NAND2_X1 pe_1_0_4_U9 ( .A1(pe_1_0_4_n44), .A2(pe_1_0_4_n60), .ZN(
        pe_1_0_4_n42) );
  INV_X1 pe_1_0_4_U8 ( .A(pe_1_0_4_n69), .ZN(pe_1_0_4_n65) );
  BUF_X1 pe_1_0_4_U7 ( .A(pe_1_0_4_n60), .Z(pe_1_0_4_n56) );
  INV_X1 pe_1_0_4_U6 ( .A(pe_1_0_4_n42), .ZN(pe_1_0_4_n89) );
  INV_X1 pe_1_0_4_U5 ( .A(pe_1_0_4_n40), .ZN(pe_1_0_4_n85) );
  INV_X2 pe_1_0_4_U4 ( .A(n81), .ZN(pe_1_0_4_n72) );
  XOR2_X1 pe_1_0_4_U3 ( .A(pe_1_0_4_int_data_0_), .B(o_data[24]), .Z(
        pe_1_0_4_n1) );
  DFFR_X1 pe_1_0_4_int_q_acc_reg_0_ ( .D(pe_1_0_4_n84), .CK(pe_1_0_4_net7240), 
        .RN(pe_1_0_4_n72), .Q(o_data[24]), .QN(pe_1_0_4_n3) );
  DFFR_X1 pe_1_0_4_int_q_reg_v_reg_0__0_ ( .D(int_data_y_1__4__0_), .CK(
        pe_1_0_4_net7210), .RN(pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_v[20]) );
  DFFR_X1 pe_1_0_4_int_q_reg_v_reg_0__1_ ( .D(int_data_y_1__4__1_), .CK(
        pe_1_0_4_net7210), .RN(pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_v[21]) );
  DFFR_X1 pe_1_0_4_int_q_reg_v_reg_0__2_ ( .D(int_data_y_1__4__2_), .CK(
        pe_1_0_4_net7210), .RN(pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_v[22]) );
  DFFR_X1 pe_1_0_4_int_q_reg_v_reg_0__3_ ( .D(int_data_y_1__4__3_), .CK(
        pe_1_0_4_net7210), .RN(pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_v[23]) );
  DFFR_X1 pe_1_0_4_int_q_reg_v_reg_1__0_ ( .D(int_data_y_1__4__0_), .CK(
        pe_1_0_4_net7215), .RN(pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_v[16]) );
  DFFR_X1 pe_1_0_4_int_q_reg_v_reg_1__1_ ( .D(int_data_y_1__4__1_), .CK(
        pe_1_0_4_net7215), .RN(pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_v[17]) );
  DFFR_X1 pe_1_0_4_int_q_reg_v_reg_1__2_ ( .D(int_data_y_1__4__2_), .CK(
        pe_1_0_4_net7215), .RN(pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_v[18]) );
  DFFR_X1 pe_1_0_4_int_q_reg_v_reg_1__3_ ( .D(int_data_y_1__4__3_), .CK(
        pe_1_0_4_net7215), .RN(pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_v[19]) );
  DFFR_X1 pe_1_0_4_int_q_reg_v_reg_2__0_ ( .D(int_data_y_1__4__0_), .CK(
        pe_1_0_4_net7220), .RN(pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_v[12]) );
  DFFR_X1 pe_1_0_4_int_q_reg_v_reg_2__1_ ( .D(int_data_y_1__4__1_), .CK(
        pe_1_0_4_net7220), .RN(pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_v[13]) );
  DFFR_X1 pe_1_0_4_int_q_reg_v_reg_2__2_ ( .D(int_data_y_1__4__2_), .CK(
        pe_1_0_4_net7220), .RN(pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_v[14]) );
  DFFR_X1 pe_1_0_4_int_q_reg_v_reg_2__3_ ( .D(int_data_y_1__4__3_), .CK(
        pe_1_0_4_net7220), .RN(pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_v[15]) );
  DFFR_X1 pe_1_0_4_int_q_reg_v_reg_3__0_ ( .D(int_data_y_1__4__0_), .CK(
        pe_1_0_4_net7225), .RN(pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_v[8]) );
  DFFR_X1 pe_1_0_4_int_q_reg_v_reg_3__1_ ( .D(int_data_y_1__4__1_), .CK(
        pe_1_0_4_net7225), .RN(pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_v[9]) );
  DFFR_X1 pe_1_0_4_int_q_reg_v_reg_3__2_ ( .D(int_data_y_1__4__2_), .CK(
        pe_1_0_4_net7225), .RN(pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_v[10]) );
  DFFR_X1 pe_1_0_4_int_q_reg_v_reg_3__3_ ( .D(int_data_y_1__4__3_), .CK(
        pe_1_0_4_net7225), .RN(pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_v[11]) );
  DFFR_X1 pe_1_0_4_int_q_reg_v_reg_4__0_ ( .D(int_data_y_1__4__0_), .CK(
        pe_1_0_4_net7230), .RN(pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_v[4]) );
  DFFR_X1 pe_1_0_4_int_q_reg_v_reg_4__1_ ( .D(int_data_y_1__4__1_), .CK(
        pe_1_0_4_net7230), .RN(pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_v[5]) );
  DFFR_X1 pe_1_0_4_int_q_reg_v_reg_4__2_ ( .D(int_data_y_1__4__2_), .CK(
        pe_1_0_4_net7230), .RN(pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_v[6]) );
  DFFR_X1 pe_1_0_4_int_q_reg_v_reg_4__3_ ( .D(int_data_y_1__4__3_), .CK(
        pe_1_0_4_net7230), .RN(pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_v[7]) );
  DFFR_X1 pe_1_0_4_int_q_reg_v_reg_5__0_ ( .D(int_data_y_1__4__0_), .CK(
        pe_1_0_4_net7235), .RN(pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_v[0]) );
  DFFR_X1 pe_1_0_4_int_q_reg_v_reg_5__1_ ( .D(int_data_y_1__4__1_), .CK(
        pe_1_0_4_net7235), .RN(pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_v[1]) );
  DFFR_X1 pe_1_0_4_int_q_reg_v_reg_5__2_ ( .D(int_data_y_1__4__2_), .CK(
        pe_1_0_4_net7235), .RN(pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_v[2]) );
  DFFR_X1 pe_1_0_4_int_q_reg_v_reg_5__3_ ( .D(int_data_y_1__4__3_), .CK(
        pe_1_0_4_net7235), .RN(pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_0_4_int_q_reg_h_reg_0__0_ ( .D(int_data_x_0__5__0_), .SI(
        int_data_y_1__4__0_), .SE(pe_1_0_4_n65), .CK(pe_1_0_4_net7179), .RN(
        pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_0_4_int_q_reg_h_reg_0__1_ ( .D(int_data_x_0__5__1_), .SI(
        int_data_y_1__4__1_), .SE(pe_1_0_4_n65), .CK(pe_1_0_4_net7179), .RN(
        pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_0_4_int_q_reg_h_reg_0__2_ ( .D(int_data_x_0__5__2_), .SI(
        int_data_y_1__4__2_), .SE(pe_1_0_4_n65), .CK(pe_1_0_4_net7179), .RN(
        pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_0_4_int_q_reg_h_reg_0__3_ ( .D(int_data_x_0__5__3_), .SI(
        int_data_y_1__4__3_), .SE(pe_1_0_4_n65), .CK(pe_1_0_4_net7179), .RN(
        pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_0_4_int_q_reg_h_reg_1__0_ ( .D(int_data_x_0__5__0_), .SI(
        int_data_y_1__4__0_), .SE(pe_1_0_4_n65), .CK(pe_1_0_4_net7185), .RN(
        pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_0_4_int_q_reg_h_reg_1__1_ ( .D(int_data_x_0__5__1_), .SI(
        int_data_y_1__4__1_), .SE(pe_1_0_4_n65), .CK(pe_1_0_4_net7185), .RN(
        pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_0_4_int_q_reg_h_reg_1__2_ ( .D(int_data_x_0__5__2_), .SI(
        int_data_y_1__4__2_), .SE(pe_1_0_4_n65), .CK(pe_1_0_4_net7185), .RN(
        pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_0_4_int_q_reg_h_reg_1__3_ ( .D(int_data_x_0__5__3_), .SI(
        int_data_y_1__4__3_), .SE(pe_1_0_4_n65), .CK(pe_1_0_4_net7185), .RN(
        pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_0_4_int_q_reg_h_reg_2__0_ ( .D(int_data_x_0__5__0_), .SI(
        int_data_y_1__4__0_), .SE(pe_1_0_4_n65), .CK(pe_1_0_4_net7190), .RN(
        pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_0_4_int_q_reg_h_reg_2__1_ ( .D(int_data_x_0__5__1_), .SI(
        int_data_y_1__4__1_), .SE(pe_1_0_4_n65), .CK(pe_1_0_4_net7190), .RN(
        pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_0_4_int_q_reg_h_reg_2__2_ ( .D(int_data_x_0__5__2_), .SI(
        int_data_y_1__4__2_), .SE(pe_1_0_4_n65), .CK(pe_1_0_4_net7190), .RN(
        pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_0_4_int_q_reg_h_reg_2__3_ ( .D(int_data_x_0__5__3_), .SI(
        int_data_y_1__4__3_), .SE(pe_1_0_4_n65), .CK(pe_1_0_4_net7190), .RN(
        pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_0_4_int_q_reg_h_reg_3__0_ ( .D(int_data_x_0__5__0_), .SI(
        int_data_y_1__4__0_), .SE(pe_1_0_4_n65), .CK(pe_1_0_4_net7195), .RN(
        pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_0_4_int_q_reg_h_reg_3__1_ ( .D(int_data_x_0__5__1_), .SI(
        int_data_y_1__4__1_), .SE(pe_1_0_4_n65), .CK(pe_1_0_4_net7195), .RN(
        pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_0_4_int_q_reg_h_reg_3__2_ ( .D(int_data_x_0__5__2_), .SI(
        int_data_y_1__4__2_), .SE(pe_1_0_4_n65), .CK(pe_1_0_4_net7195), .RN(
        pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_0_4_int_q_reg_h_reg_3__3_ ( .D(int_data_x_0__5__3_), .SI(
        int_data_y_1__4__3_), .SE(pe_1_0_4_n65), .CK(pe_1_0_4_net7195), .RN(
        pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_0_4_int_q_reg_h_reg_4__0_ ( .D(int_data_x_0__5__0_), .SI(
        int_data_y_1__4__0_), .SE(pe_1_0_4_n66), .CK(pe_1_0_4_net7200), .RN(
        pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_0_4_int_q_reg_h_reg_4__1_ ( .D(int_data_x_0__5__1_), .SI(
        int_data_y_1__4__1_), .SE(pe_1_0_4_n66), .CK(pe_1_0_4_net7200), .RN(
        pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_0_4_int_q_reg_h_reg_4__2_ ( .D(int_data_x_0__5__2_), .SI(
        int_data_y_1__4__2_), .SE(pe_1_0_4_n66), .CK(pe_1_0_4_net7200), .RN(
        pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_0_4_int_q_reg_h_reg_4__3_ ( .D(int_data_x_0__5__3_), .SI(
        int_data_y_1__4__3_), .SE(pe_1_0_4_n66), .CK(pe_1_0_4_net7200), .RN(
        pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_0_4_int_q_reg_h_reg_5__0_ ( .D(int_data_x_0__5__0_), .SI(
        int_data_y_1__4__0_), .SE(pe_1_0_4_n66), .CK(pe_1_0_4_net7205), .RN(
        pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_0_4_int_q_reg_h_reg_5__1_ ( .D(int_data_x_0__5__1_), .SI(
        int_data_y_1__4__1_), .SE(pe_1_0_4_n66), .CK(pe_1_0_4_net7205), .RN(
        pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_0_4_int_q_reg_h_reg_5__2_ ( .D(int_data_x_0__5__2_), .SI(
        int_data_y_1__4__2_), .SE(pe_1_0_4_n66), .CK(pe_1_0_4_net7205), .RN(
        pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_0_4_int_q_reg_h_reg_5__3_ ( .D(int_data_x_0__5__3_), .SI(
        int_data_y_1__4__3_), .SE(pe_1_0_4_n66), .CK(pe_1_0_4_net7205), .RN(
        pe_1_0_4_n72), .Q(pe_1_0_4_int_q_reg_h[3]) );
  FA_X1 pe_1_0_4_sub_81_U2_7 ( .A(o_data[31]), .B(pe_1_0_4_n76), .CI(
        pe_1_0_4_sub_81_carry[7]), .S(pe_1_0_4_N77) );
  FA_X1 pe_1_0_4_sub_81_U2_6 ( .A(o_data[30]), .B(pe_1_0_4_n76), .CI(
        pe_1_0_4_sub_81_carry[6]), .CO(pe_1_0_4_sub_81_carry[7]), .S(
        pe_1_0_4_N76) );
  FA_X1 pe_1_0_4_sub_81_U2_5 ( .A(o_data[29]), .B(pe_1_0_4_n76), .CI(
        pe_1_0_4_sub_81_carry[5]), .CO(pe_1_0_4_sub_81_carry[6]), .S(
        pe_1_0_4_N75) );
  FA_X1 pe_1_0_4_sub_81_U2_4 ( .A(o_data[28]), .B(pe_1_0_4_n76), .CI(
        pe_1_0_4_sub_81_carry[4]), .CO(pe_1_0_4_sub_81_carry[5]), .S(
        pe_1_0_4_N74) );
  FA_X1 pe_1_0_4_sub_81_U2_3 ( .A(o_data[27]), .B(pe_1_0_4_n76), .CI(
        pe_1_0_4_sub_81_carry[3]), .CO(pe_1_0_4_sub_81_carry[4]), .S(
        pe_1_0_4_N73) );
  FA_X1 pe_1_0_4_sub_81_U2_2 ( .A(o_data[26]), .B(pe_1_0_4_n75), .CI(
        pe_1_0_4_sub_81_carry[2]), .CO(pe_1_0_4_sub_81_carry[3]), .S(
        pe_1_0_4_N72) );
  FA_X1 pe_1_0_4_sub_81_U2_1 ( .A(o_data[25]), .B(pe_1_0_4_n74), .CI(
        pe_1_0_4_sub_81_carry[1]), .CO(pe_1_0_4_sub_81_carry[2]), .S(
        pe_1_0_4_N71) );
  FA_X1 pe_1_0_4_add_83_U1_7 ( .A(o_data[31]), .B(pe_1_0_4_int_data_3_), .CI(
        pe_1_0_4_add_83_carry[7]), .S(pe_1_0_4_N85) );
  FA_X1 pe_1_0_4_add_83_U1_6 ( .A(o_data[30]), .B(pe_1_0_4_int_data_3_), .CI(
        pe_1_0_4_add_83_carry[6]), .CO(pe_1_0_4_add_83_carry[7]), .S(
        pe_1_0_4_N84) );
  FA_X1 pe_1_0_4_add_83_U1_5 ( .A(o_data[29]), .B(pe_1_0_4_int_data_3_), .CI(
        pe_1_0_4_add_83_carry[5]), .CO(pe_1_0_4_add_83_carry[6]), .S(
        pe_1_0_4_N83) );
  FA_X1 pe_1_0_4_add_83_U1_4 ( .A(o_data[28]), .B(pe_1_0_4_int_data_3_), .CI(
        pe_1_0_4_add_83_carry[4]), .CO(pe_1_0_4_add_83_carry[5]), .S(
        pe_1_0_4_N82) );
  FA_X1 pe_1_0_4_add_83_U1_3 ( .A(o_data[27]), .B(pe_1_0_4_int_data_3_), .CI(
        pe_1_0_4_add_83_carry[3]), .CO(pe_1_0_4_add_83_carry[4]), .S(
        pe_1_0_4_N81) );
  FA_X1 pe_1_0_4_add_83_U1_2 ( .A(o_data[26]), .B(pe_1_0_4_int_data_2_), .CI(
        pe_1_0_4_add_83_carry[2]), .CO(pe_1_0_4_add_83_carry[3]), .S(
        pe_1_0_4_N80) );
  FA_X1 pe_1_0_4_add_83_U1_1 ( .A(o_data[25]), .B(pe_1_0_4_int_data_1_), .CI(
        pe_1_0_4_n2), .CO(pe_1_0_4_add_83_carry[2]), .S(pe_1_0_4_N79) );
  NAND3_X1 pe_1_0_4_U56 ( .A1(pe_1_0_4_n60), .A2(pe_1_0_4_n43), .A3(
        pe_1_0_4_n62), .ZN(pe_1_0_4_n40) );
  NAND3_X1 pe_1_0_4_U55 ( .A1(pe_1_0_4_n43), .A2(pe_1_0_4_n61), .A3(
        pe_1_0_4_n62), .ZN(pe_1_0_4_n39) );
  NAND3_X1 pe_1_0_4_U54 ( .A1(pe_1_0_4_n43), .A2(pe_1_0_4_n63), .A3(
        pe_1_0_4_n60), .ZN(pe_1_0_4_n38) );
  NAND3_X1 pe_1_0_4_U53 ( .A1(pe_1_0_4_n61), .A2(pe_1_0_4_n63), .A3(
        pe_1_0_4_n43), .ZN(pe_1_0_4_n37) );
  DFFR_X1 pe_1_0_4_int_q_acc_reg_6_ ( .D(pe_1_0_4_n78), .CK(pe_1_0_4_net7240), 
        .RN(pe_1_0_4_n71), .Q(o_data[30]) );
  DFFR_X1 pe_1_0_4_int_q_acc_reg_5_ ( .D(pe_1_0_4_n79), .CK(pe_1_0_4_net7240), 
        .RN(pe_1_0_4_n71), .Q(o_data[29]) );
  DFFR_X1 pe_1_0_4_int_q_acc_reg_4_ ( .D(pe_1_0_4_n80), .CK(pe_1_0_4_net7240), 
        .RN(pe_1_0_4_n71), .Q(o_data[28]) );
  DFFR_X1 pe_1_0_4_int_q_acc_reg_3_ ( .D(pe_1_0_4_n81), .CK(pe_1_0_4_net7240), 
        .RN(pe_1_0_4_n71), .Q(o_data[27]) );
  DFFR_X1 pe_1_0_4_int_q_acc_reg_2_ ( .D(pe_1_0_4_n82), .CK(pe_1_0_4_net7240), 
        .RN(pe_1_0_4_n71), .Q(o_data[26]) );
  DFFR_X1 pe_1_0_4_int_q_acc_reg_1_ ( .D(pe_1_0_4_n83), .CK(pe_1_0_4_net7240), 
        .RN(pe_1_0_4_n71), .Q(o_data[25]) );
  DFFR_X1 pe_1_0_4_int_q_acc_reg_7_ ( .D(pe_1_0_4_n77), .CK(pe_1_0_4_net7240), 
        .RN(pe_1_0_4_n71), .Q(o_data[31]) );
  CLKGATETST_X1 pe_1_0_4_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_0_4_n88), .SE(1'b0), .GCK(pe_1_0_4_net7179) );
  CLKGATETST_X1 pe_1_0_4_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_0_4_n87), .SE(1'b0), .GCK(pe_1_0_4_net7185) );
  CLKGATETST_X1 pe_1_0_4_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_0_4_n86), .SE(1'b0), .GCK(pe_1_0_4_net7190) );
  CLKGATETST_X1 pe_1_0_4_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_0_4_n85), .SE(1'b0), .GCK(pe_1_0_4_net7195) );
  CLKGATETST_X1 pe_1_0_4_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_0_4_n90), .SE(1'b0), .GCK(pe_1_0_4_net7200) );
  CLKGATETST_X1 pe_1_0_4_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_0_4_n89), .SE(1'b0), .GCK(pe_1_0_4_net7205) );
  CLKGATETST_X1 pe_1_0_4_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_0_4_N64), .SE(1'b0), .GCK(pe_1_0_4_net7210) );
  CLKGATETST_X1 pe_1_0_4_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_0_4_N63), .SE(1'b0), .GCK(pe_1_0_4_net7215) );
  CLKGATETST_X1 pe_1_0_4_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_0_4_N62), .SE(1'b0), .GCK(pe_1_0_4_net7220) );
  CLKGATETST_X1 pe_1_0_4_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_0_4_N61), .SE(1'b0), .GCK(pe_1_0_4_net7225) );
  CLKGATETST_X1 pe_1_0_4_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_0_4_N60), .SE(1'b0), .GCK(pe_1_0_4_net7230) );
  CLKGATETST_X1 pe_1_0_4_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_0_4_N59), .SE(1'b0), .GCK(pe_1_0_4_net7235) );
  CLKGATETST_X1 pe_1_0_4_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_0_4_N90), .SE(1'b0), .GCK(pe_1_0_4_net7240) );
  CLKBUF_X1 pe_1_0_5_U112 ( .A(pe_1_0_5_n72), .Z(pe_1_0_5_n71) );
  INV_X1 pe_1_0_5_U111 ( .A(n73), .ZN(pe_1_0_5_n70) );
  INV_X1 pe_1_0_5_U110 ( .A(n65), .ZN(pe_1_0_5_n69) );
  INV_X1 pe_1_0_5_U109 ( .A(n65), .ZN(pe_1_0_5_n68) );
  INV_X1 pe_1_0_5_U108 ( .A(n65), .ZN(pe_1_0_5_n67) );
  INV_X1 pe_1_0_5_U107 ( .A(pe_1_0_5_n69), .ZN(pe_1_0_5_n66) );
  INV_X1 pe_1_0_5_U106 ( .A(pe_1_0_5_n63), .ZN(pe_1_0_5_n62) );
  INV_X1 pe_1_0_5_U105 ( .A(pe_1_0_5_n61), .ZN(pe_1_0_5_n60) );
  INV_X1 pe_1_0_5_U104 ( .A(n25), .ZN(pe_1_0_5_n59) );
  INV_X1 pe_1_0_5_U103 ( .A(pe_1_0_5_n59), .ZN(pe_1_0_5_n58) );
  INV_X1 pe_1_0_5_U102 ( .A(n17), .ZN(pe_1_0_5_n57) );
  MUX2_X1 pe_1_0_5_U101 ( .A(pe_1_0_5_n54), .B(pe_1_0_5_n51), .S(n44), .Z(
        int_data_x_0__5__3_) );
  MUX2_X1 pe_1_0_5_U100 ( .A(pe_1_0_5_n53), .B(pe_1_0_5_n52), .S(pe_1_0_5_n62), 
        .Z(pe_1_0_5_n54) );
  MUX2_X1 pe_1_0_5_U99 ( .A(pe_1_0_5_int_q_reg_h[23]), .B(
        pe_1_0_5_int_q_reg_h[19]), .S(pe_1_0_5_n56), .Z(pe_1_0_5_n53) );
  MUX2_X1 pe_1_0_5_U98 ( .A(pe_1_0_5_int_q_reg_h[15]), .B(
        pe_1_0_5_int_q_reg_h[11]), .S(pe_1_0_5_n56), .Z(pe_1_0_5_n52) );
  MUX2_X1 pe_1_0_5_U97 ( .A(pe_1_0_5_int_q_reg_h[7]), .B(
        pe_1_0_5_int_q_reg_h[3]), .S(pe_1_0_5_n56), .Z(pe_1_0_5_n51) );
  MUX2_X1 pe_1_0_5_U96 ( .A(pe_1_0_5_n50), .B(pe_1_0_5_n47), .S(n44), .Z(
        int_data_x_0__5__2_) );
  MUX2_X1 pe_1_0_5_U95 ( .A(pe_1_0_5_n49), .B(pe_1_0_5_n48), .S(pe_1_0_5_n62), 
        .Z(pe_1_0_5_n50) );
  MUX2_X1 pe_1_0_5_U94 ( .A(pe_1_0_5_int_q_reg_h[22]), .B(
        pe_1_0_5_int_q_reg_h[18]), .S(pe_1_0_5_n56), .Z(pe_1_0_5_n49) );
  MUX2_X1 pe_1_0_5_U93 ( .A(pe_1_0_5_int_q_reg_h[14]), .B(
        pe_1_0_5_int_q_reg_h[10]), .S(pe_1_0_5_n56), .Z(pe_1_0_5_n48) );
  MUX2_X1 pe_1_0_5_U92 ( .A(pe_1_0_5_int_q_reg_h[6]), .B(
        pe_1_0_5_int_q_reg_h[2]), .S(pe_1_0_5_n56), .Z(pe_1_0_5_n47) );
  MUX2_X1 pe_1_0_5_U91 ( .A(pe_1_0_5_n46), .B(pe_1_0_5_n24), .S(n44), .Z(
        int_data_x_0__5__1_) );
  MUX2_X1 pe_1_0_5_U90 ( .A(pe_1_0_5_n45), .B(pe_1_0_5_n25), .S(pe_1_0_5_n62), 
        .Z(pe_1_0_5_n46) );
  MUX2_X1 pe_1_0_5_U89 ( .A(pe_1_0_5_int_q_reg_h[21]), .B(
        pe_1_0_5_int_q_reg_h[17]), .S(pe_1_0_5_n56), .Z(pe_1_0_5_n45) );
  MUX2_X1 pe_1_0_5_U88 ( .A(pe_1_0_5_int_q_reg_h[13]), .B(
        pe_1_0_5_int_q_reg_h[9]), .S(pe_1_0_5_n56), .Z(pe_1_0_5_n25) );
  MUX2_X1 pe_1_0_5_U87 ( .A(pe_1_0_5_int_q_reg_h[5]), .B(
        pe_1_0_5_int_q_reg_h[1]), .S(pe_1_0_5_n56), .Z(pe_1_0_5_n24) );
  MUX2_X1 pe_1_0_5_U86 ( .A(pe_1_0_5_n23), .B(pe_1_0_5_n20), .S(n44), .Z(
        int_data_x_0__5__0_) );
  MUX2_X1 pe_1_0_5_U85 ( .A(pe_1_0_5_n22), .B(pe_1_0_5_n21), .S(pe_1_0_5_n62), 
        .Z(pe_1_0_5_n23) );
  MUX2_X1 pe_1_0_5_U84 ( .A(pe_1_0_5_int_q_reg_h[20]), .B(
        pe_1_0_5_int_q_reg_h[16]), .S(pe_1_0_5_n56), .Z(pe_1_0_5_n22) );
  MUX2_X1 pe_1_0_5_U83 ( .A(pe_1_0_5_int_q_reg_h[12]), .B(
        pe_1_0_5_int_q_reg_h[8]), .S(pe_1_0_5_n56), .Z(pe_1_0_5_n21) );
  MUX2_X1 pe_1_0_5_U82 ( .A(pe_1_0_5_int_q_reg_h[4]), .B(
        pe_1_0_5_int_q_reg_h[0]), .S(pe_1_0_5_n56), .Z(pe_1_0_5_n20) );
  MUX2_X1 pe_1_0_5_U81 ( .A(pe_1_0_5_n19), .B(pe_1_0_5_n16), .S(n44), .Z(
        pe_1_0_5_o_data_v_3_) );
  MUX2_X1 pe_1_0_5_U80 ( .A(pe_1_0_5_n18), .B(pe_1_0_5_n17), .S(pe_1_0_5_n62), 
        .Z(pe_1_0_5_n19) );
  MUX2_X1 pe_1_0_5_U79 ( .A(pe_1_0_5_int_q_reg_v[23]), .B(
        pe_1_0_5_int_q_reg_v[19]), .S(pe_1_0_5_n55), .Z(pe_1_0_5_n18) );
  MUX2_X1 pe_1_0_5_U78 ( .A(pe_1_0_5_int_q_reg_v[15]), .B(
        pe_1_0_5_int_q_reg_v[11]), .S(pe_1_0_5_n55), .Z(pe_1_0_5_n17) );
  MUX2_X1 pe_1_0_5_U77 ( .A(pe_1_0_5_int_q_reg_v[7]), .B(
        pe_1_0_5_int_q_reg_v[3]), .S(pe_1_0_5_n55), .Z(pe_1_0_5_n16) );
  MUX2_X1 pe_1_0_5_U76 ( .A(pe_1_0_5_n15), .B(pe_1_0_5_n12), .S(n44), .Z(
        pe_1_0_5_o_data_v_2_) );
  MUX2_X1 pe_1_0_5_U75 ( .A(pe_1_0_5_n14), .B(pe_1_0_5_n13), .S(pe_1_0_5_n62), 
        .Z(pe_1_0_5_n15) );
  MUX2_X1 pe_1_0_5_U74 ( .A(pe_1_0_5_int_q_reg_v[22]), .B(
        pe_1_0_5_int_q_reg_v[18]), .S(pe_1_0_5_n55), .Z(pe_1_0_5_n14) );
  MUX2_X1 pe_1_0_5_U73 ( .A(pe_1_0_5_int_q_reg_v[14]), .B(
        pe_1_0_5_int_q_reg_v[10]), .S(pe_1_0_5_n55), .Z(pe_1_0_5_n13) );
  MUX2_X1 pe_1_0_5_U72 ( .A(pe_1_0_5_int_q_reg_v[6]), .B(
        pe_1_0_5_int_q_reg_v[2]), .S(pe_1_0_5_n55), .Z(pe_1_0_5_n12) );
  MUX2_X1 pe_1_0_5_U71 ( .A(pe_1_0_5_n11), .B(pe_1_0_5_n8), .S(n44), .Z(
        pe_1_0_5_o_data_v_1_) );
  MUX2_X1 pe_1_0_5_U70 ( .A(pe_1_0_5_n10), .B(pe_1_0_5_n9), .S(pe_1_0_5_n62), 
        .Z(pe_1_0_5_n11) );
  MUX2_X1 pe_1_0_5_U69 ( .A(pe_1_0_5_int_q_reg_v[21]), .B(
        pe_1_0_5_int_q_reg_v[17]), .S(pe_1_0_5_n55), .Z(pe_1_0_5_n10) );
  MUX2_X1 pe_1_0_5_U68 ( .A(pe_1_0_5_int_q_reg_v[13]), .B(
        pe_1_0_5_int_q_reg_v[9]), .S(pe_1_0_5_n55), .Z(pe_1_0_5_n9) );
  MUX2_X1 pe_1_0_5_U67 ( .A(pe_1_0_5_int_q_reg_v[5]), .B(
        pe_1_0_5_int_q_reg_v[1]), .S(pe_1_0_5_n55), .Z(pe_1_0_5_n8) );
  MUX2_X1 pe_1_0_5_U66 ( .A(pe_1_0_5_n7), .B(pe_1_0_5_n4), .S(n44), .Z(
        pe_1_0_5_o_data_v_0_) );
  MUX2_X1 pe_1_0_5_U65 ( .A(pe_1_0_5_n6), .B(pe_1_0_5_n5), .S(pe_1_0_5_n62), 
        .Z(pe_1_0_5_n7) );
  MUX2_X1 pe_1_0_5_U64 ( .A(pe_1_0_5_int_q_reg_v[20]), .B(
        pe_1_0_5_int_q_reg_v[16]), .S(pe_1_0_5_n55), .Z(pe_1_0_5_n6) );
  MUX2_X1 pe_1_0_5_U63 ( .A(pe_1_0_5_int_q_reg_v[12]), .B(
        pe_1_0_5_int_q_reg_v[8]), .S(pe_1_0_5_n55), .Z(pe_1_0_5_n5) );
  MUX2_X1 pe_1_0_5_U62 ( .A(pe_1_0_5_int_q_reg_v[4]), .B(
        pe_1_0_5_int_q_reg_v[0]), .S(pe_1_0_5_n55), .Z(pe_1_0_5_n4) );
  XNOR2_X1 pe_1_0_5_U61 ( .A(pe_1_0_5_n73), .B(o_data[16]), .ZN(pe_1_0_5_N70)
         );
  AOI222_X1 pe_1_0_5_U60 ( .A1(int_data_res_1__5__0_), .A2(pe_1_0_5_n64), .B1(
        pe_1_0_5_n1), .B2(pe_1_0_5_n27), .C1(pe_1_0_5_N70), .C2(pe_1_0_5_n28), 
        .ZN(pe_1_0_5_n35) );
  INV_X1 pe_1_0_5_U59 ( .A(pe_1_0_5_n35), .ZN(pe_1_0_5_n84) );
  AOI222_X1 pe_1_0_5_U58 ( .A1(int_data_res_1__5__2_), .A2(pe_1_0_5_n64), .B1(
        pe_1_0_5_N80), .B2(pe_1_0_5_n27), .C1(pe_1_0_5_N72), .C2(pe_1_0_5_n28), 
        .ZN(pe_1_0_5_n33) );
  INV_X1 pe_1_0_5_U57 ( .A(pe_1_0_5_n33), .ZN(pe_1_0_5_n82) );
  AOI222_X1 pe_1_0_5_U52 ( .A1(int_data_res_1__5__6_), .A2(pe_1_0_5_n64), .B1(
        pe_1_0_5_N84), .B2(pe_1_0_5_n27), .C1(pe_1_0_5_N76), .C2(pe_1_0_5_n28), 
        .ZN(pe_1_0_5_n29) );
  INV_X1 pe_1_0_5_U51 ( .A(pe_1_0_5_n29), .ZN(pe_1_0_5_n78) );
  AOI222_X1 pe_1_0_5_U50 ( .A1(int_data_res_1__5__1_), .A2(pe_1_0_5_n64), .B1(
        pe_1_0_5_N79), .B2(pe_1_0_5_n27), .C1(pe_1_0_5_N71), .C2(pe_1_0_5_n28), 
        .ZN(pe_1_0_5_n34) );
  INV_X1 pe_1_0_5_U49 ( .A(pe_1_0_5_n34), .ZN(pe_1_0_5_n83) );
  AOI222_X1 pe_1_0_5_U48 ( .A1(int_data_res_1__5__3_), .A2(pe_1_0_5_n64), .B1(
        pe_1_0_5_N81), .B2(pe_1_0_5_n27), .C1(pe_1_0_5_N73), .C2(pe_1_0_5_n28), 
        .ZN(pe_1_0_5_n32) );
  INV_X1 pe_1_0_5_U47 ( .A(pe_1_0_5_n32), .ZN(pe_1_0_5_n81) );
  AOI222_X1 pe_1_0_5_U46 ( .A1(int_data_res_1__5__4_), .A2(pe_1_0_5_n64), .B1(
        pe_1_0_5_N82), .B2(pe_1_0_5_n27), .C1(pe_1_0_5_N74), .C2(pe_1_0_5_n28), 
        .ZN(pe_1_0_5_n31) );
  INV_X1 pe_1_0_5_U45 ( .A(pe_1_0_5_n31), .ZN(pe_1_0_5_n80) );
  AOI222_X1 pe_1_0_5_U44 ( .A1(int_data_res_1__5__5_), .A2(pe_1_0_5_n64), .B1(
        pe_1_0_5_N83), .B2(pe_1_0_5_n27), .C1(pe_1_0_5_N75), .C2(pe_1_0_5_n28), 
        .ZN(pe_1_0_5_n30) );
  INV_X1 pe_1_0_5_U43 ( .A(pe_1_0_5_n30), .ZN(pe_1_0_5_n79) );
  INV_X1 pe_1_0_5_U42 ( .A(pe_1_0_5_int_data_2_), .ZN(pe_1_0_5_n75) );
  NAND2_X1 pe_1_0_5_U41 ( .A1(pe_1_0_5_int_data_0_), .A2(pe_1_0_5_n3), .ZN(
        pe_1_0_5_sub_81_carry[1]) );
  INV_X1 pe_1_0_5_U40 ( .A(pe_1_0_5_int_data_1_), .ZN(pe_1_0_5_n74) );
  AND2_X1 pe_1_0_5_U39 ( .A1(pe_1_0_5_int_data_0_), .A2(o_data[16]), .ZN(
        pe_1_0_5_n2) );
  AOI222_X1 pe_1_0_5_U38 ( .A1(pe_1_0_5_n64), .A2(int_data_res_1__5__7_), .B1(
        pe_1_0_5_N85), .B2(pe_1_0_5_n27), .C1(pe_1_0_5_N77), .C2(pe_1_0_5_n28), 
        .ZN(pe_1_0_5_n26) );
  INV_X1 pe_1_0_5_U37 ( .A(pe_1_0_5_n26), .ZN(pe_1_0_5_n77) );
  NOR3_X1 pe_1_0_5_U36 ( .A1(pe_1_0_5_n59), .A2(pe_1_0_5_n65), .A3(int_ckg[58]), .ZN(pe_1_0_5_n36) );
  OR2_X1 pe_1_0_5_U35 ( .A1(pe_1_0_5_n36), .A2(pe_1_0_5_n64), .ZN(pe_1_0_5_N90) );
  INV_X1 pe_1_0_5_U34 ( .A(n37), .ZN(pe_1_0_5_n63) );
  AND2_X1 pe_1_0_5_U33 ( .A1(int_data_x_0__5__2_), .A2(pe_1_0_5_n58), .ZN(
        pe_1_0_5_int_data_2_) );
  AND2_X1 pe_1_0_5_U32 ( .A1(int_data_x_0__5__1_), .A2(pe_1_0_5_n58), .ZN(
        pe_1_0_5_int_data_1_) );
  AND2_X1 pe_1_0_5_U31 ( .A1(int_data_x_0__5__3_), .A2(pe_1_0_5_n58), .ZN(
        pe_1_0_5_int_data_3_) );
  BUF_X1 pe_1_0_5_U30 ( .A(n59), .Z(pe_1_0_5_n64) );
  INV_X1 pe_1_0_5_U29 ( .A(n31), .ZN(pe_1_0_5_n61) );
  AND2_X1 pe_1_0_5_U28 ( .A1(int_data_x_0__5__0_), .A2(pe_1_0_5_n58), .ZN(
        pe_1_0_5_int_data_0_) );
  NAND2_X1 pe_1_0_5_U27 ( .A1(pe_1_0_5_n44), .A2(pe_1_0_5_n61), .ZN(
        pe_1_0_5_n41) );
  AND3_X1 pe_1_0_5_U26 ( .A1(n73), .A2(pe_1_0_5_n63), .A3(n44), .ZN(
        pe_1_0_5_n44) );
  INV_X1 pe_1_0_5_U25 ( .A(pe_1_0_5_int_data_3_), .ZN(pe_1_0_5_n76) );
  NOR2_X1 pe_1_0_5_U24 ( .A1(pe_1_0_5_n70), .A2(n44), .ZN(pe_1_0_5_n43) );
  NOR2_X1 pe_1_0_5_U23 ( .A1(pe_1_0_5_n57), .A2(pe_1_0_5_n64), .ZN(
        pe_1_0_5_n28) );
  NOR2_X1 pe_1_0_5_U22 ( .A1(n17), .A2(pe_1_0_5_n64), .ZN(pe_1_0_5_n27) );
  INV_X1 pe_1_0_5_U21 ( .A(pe_1_0_5_int_data_0_), .ZN(pe_1_0_5_n73) );
  BUF_X1 pe_1_0_5_U20 ( .A(pe_1_0_5_n60), .Z(pe_1_0_5_n55) );
  INV_X1 pe_1_0_5_U19 ( .A(pe_1_0_5_n41), .ZN(pe_1_0_5_n90) );
  INV_X1 pe_1_0_5_U18 ( .A(pe_1_0_5_n37), .ZN(pe_1_0_5_n88) );
  INV_X1 pe_1_0_5_U17 ( .A(pe_1_0_5_n38), .ZN(pe_1_0_5_n87) );
  INV_X1 pe_1_0_5_U16 ( .A(pe_1_0_5_n39), .ZN(pe_1_0_5_n86) );
  NOR2_X1 pe_1_0_5_U15 ( .A1(pe_1_0_5_n68), .A2(pe_1_0_5_n42), .ZN(
        pe_1_0_5_N59) );
  NOR2_X1 pe_1_0_5_U14 ( .A1(pe_1_0_5_n68), .A2(pe_1_0_5_n41), .ZN(
        pe_1_0_5_N60) );
  NOR2_X1 pe_1_0_5_U13 ( .A1(pe_1_0_5_n68), .A2(pe_1_0_5_n38), .ZN(
        pe_1_0_5_N63) );
  NOR2_X1 pe_1_0_5_U12 ( .A1(pe_1_0_5_n67), .A2(pe_1_0_5_n40), .ZN(
        pe_1_0_5_N61) );
  NOR2_X1 pe_1_0_5_U11 ( .A1(pe_1_0_5_n67), .A2(pe_1_0_5_n39), .ZN(
        pe_1_0_5_N62) );
  NOR2_X1 pe_1_0_5_U10 ( .A1(pe_1_0_5_n37), .A2(pe_1_0_5_n67), .ZN(
        pe_1_0_5_N64) );
  NAND2_X1 pe_1_0_5_U9 ( .A1(pe_1_0_5_n44), .A2(pe_1_0_5_n60), .ZN(
        pe_1_0_5_n42) );
  INV_X1 pe_1_0_5_U8 ( .A(pe_1_0_5_n69), .ZN(pe_1_0_5_n65) );
  BUF_X1 pe_1_0_5_U7 ( .A(pe_1_0_5_n60), .Z(pe_1_0_5_n56) );
  INV_X1 pe_1_0_5_U6 ( .A(pe_1_0_5_n42), .ZN(pe_1_0_5_n89) );
  INV_X1 pe_1_0_5_U5 ( .A(pe_1_0_5_n40), .ZN(pe_1_0_5_n85) );
  INV_X2 pe_1_0_5_U4 ( .A(n81), .ZN(pe_1_0_5_n72) );
  XOR2_X1 pe_1_0_5_U3 ( .A(pe_1_0_5_int_data_0_), .B(o_data[16]), .Z(
        pe_1_0_5_n1) );
  DFFR_X1 pe_1_0_5_int_q_acc_reg_0_ ( .D(pe_1_0_5_n84), .CK(pe_1_0_5_net7162), 
        .RN(pe_1_0_5_n72), .Q(o_data[16]), .QN(pe_1_0_5_n3) );
  DFFR_X1 pe_1_0_5_int_q_reg_v_reg_0__0_ ( .D(int_data_y_1__5__0_), .CK(
        pe_1_0_5_net7132), .RN(pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_v[20]) );
  DFFR_X1 pe_1_0_5_int_q_reg_v_reg_0__1_ ( .D(int_data_y_1__5__1_), .CK(
        pe_1_0_5_net7132), .RN(pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_v[21]) );
  DFFR_X1 pe_1_0_5_int_q_reg_v_reg_0__2_ ( .D(int_data_y_1__5__2_), .CK(
        pe_1_0_5_net7132), .RN(pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_v[22]) );
  DFFR_X1 pe_1_0_5_int_q_reg_v_reg_0__3_ ( .D(int_data_y_1__5__3_), .CK(
        pe_1_0_5_net7132), .RN(pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_v[23]) );
  DFFR_X1 pe_1_0_5_int_q_reg_v_reg_1__0_ ( .D(int_data_y_1__5__0_), .CK(
        pe_1_0_5_net7137), .RN(pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_v[16]) );
  DFFR_X1 pe_1_0_5_int_q_reg_v_reg_1__1_ ( .D(int_data_y_1__5__1_), .CK(
        pe_1_0_5_net7137), .RN(pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_v[17]) );
  DFFR_X1 pe_1_0_5_int_q_reg_v_reg_1__2_ ( .D(int_data_y_1__5__2_), .CK(
        pe_1_0_5_net7137), .RN(pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_v[18]) );
  DFFR_X1 pe_1_0_5_int_q_reg_v_reg_1__3_ ( .D(int_data_y_1__5__3_), .CK(
        pe_1_0_5_net7137), .RN(pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_v[19]) );
  DFFR_X1 pe_1_0_5_int_q_reg_v_reg_2__0_ ( .D(int_data_y_1__5__0_), .CK(
        pe_1_0_5_net7142), .RN(pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_v[12]) );
  DFFR_X1 pe_1_0_5_int_q_reg_v_reg_2__1_ ( .D(int_data_y_1__5__1_), .CK(
        pe_1_0_5_net7142), .RN(pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_v[13]) );
  DFFR_X1 pe_1_0_5_int_q_reg_v_reg_2__2_ ( .D(int_data_y_1__5__2_), .CK(
        pe_1_0_5_net7142), .RN(pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_v[14]) );
  DFFR_X1 pe_1_0_5_int_q_reg_v_reg_2__3_ ( .D(int_data_y_1__5__3_), .CK(
        pe_1_0_5_net7142), .RN(pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_v[15]) );
  DFFR_X1 pe_1_0_5_int_q_reg_v_reg_3__0_ ( .D(int_data_y_1__5__0_), .CK(
        pe_1_0_5_net7147), .RN(pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_v[8]) );
  DFFR_X1 pe_1_0_5_int_q_reg_v_reg_3__1_ ( .D(int_data_y_1__5__1_), .CK(
        pe_1_0_5_net7147), .RN(pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_v[9]) );
  DFFR_X1 pe_1_0_5_int_q_reg_v_reg_3__2_ ( .D(int_data_y_1__5__2_), .CK(
        pe_1_0_5_net7147), .RN(pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_v[10]) );
  DFFR_X1 pe_1_0_5_int_q_reg_v_reg_3__3_ ( .D(int_data_y_1__5__3_), .CK(
        pe_1_0_5_net7147), .RN(pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_v[11]) );
  DFFR_X1 pe_1_0_5_int_q_reg_v_reg_4__0_ ( .D(int_data_y_1__5__0_), .CK(
        pe_1_0_5_net7152), .RN(pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_v[4]) );
  DFFR_X1 pe_1_0_5_int_q_reg_v_reg_4__1_ ( .D(int_data_y_1__5__1_), .CK(
        pe_1_0_5_net7152), .RN(pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_v[5]) );
  DFFR_X1 pe_1_0_5_int_q_reg_v_reg_4__2_ ( .D(int_data_y_1__5__2_), .CK(
        pe_1_0_5_net7152), .RN(pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_v[6]) );
  DFFR_X1 pe_1_0_5_int_q_reg_v_reg_4__3_ ( .D(int_data_y_1__5__3_), .CK(
        pe_1_0_5_net7152), .RN(pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_v[7]) );
  DFFR_X1 pe_1_0_5_int_q_reg_v_reg_5__0_ ( .D(int_data_y_1__5__0_), .CK(
        pe_1_0_5_net7157), .RN(pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_v[0]) );
  DFFR_X1 pe_1_0_5_int_q_reg_v_reg_5__1_ ( .D(int_data_y_1__5__1_), .CK(
        pe_1_0_5_net7157), .RN(pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_v[1]) );
  DFFR_X1 pe_1_0_5_int_q_reg_v_reg_5__2_ ( .D(int_data_y_1__5__2_), .CK(
        pe_1_0_5_net7157), .RN(pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_v[2]) );
  DFFR_X1 pe_1_0_5_int_q_reg_v_reg_5__3_ ( .D(int_data_y_1__5__3_), .CK(
        pe_1_0_5_net7157), .RN(pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_0_5_int_q_reg_h_reg_0__0_ ( .D(int_data_x_0__6__0_), .SI(
        int_data_y_1__5__0_), .SE(pe_1_0_5_n65), .CK(pe_1_0_5_net7101), .RN(
        pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_0_5_int_q_reg_h_reg_0__1_ ( .D(int_data_x_0__6__1_), .SI(
        int_data_y_1__5__1_), .SE(pe_1_0_5_n65), .CK(pe_1_0_5_net7101), .RN(
        pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_0_5_int_q_reg_h_reg_0__2_ ( .D(int_data_x_0__6__2_), .SI(
        int_data_y_1__5__2_), .SE(pe_1_0_5_n65), .CK(pe_1_0_5_net7101), .RN(
        pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_0_5_int_q_reg_h_reg_0__3_ ( .D(int_data_x_0__6__3_), .SI(
        int_data_y_1__5__3_), .SE(pe_1_0_5_n65), .CK(pe_1_0_5_net7101), .RN(
        pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_0_5_int_q_reg_h_reg_1__0_ ( .D(int_data_x_0__6__0_), .SI(
        int_data_y_1__5__0_), .SE(pe_1_0_5_n65), .CK(pe_1_0_5_net7107), .RN(
        pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_0_5_int_q_reg_h_reg_1__1_ ( .D(int_data_x_0__6__1_), .SI(
        int_data_y_1__5__1_), .SE(pe_1_0_5_n65), .CK(pe_1_0_5_net7107), .RN(
        pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_0_5_int_q_reg_h_reg_1__2_ ( .D(int_data_x_0__6__2_), .SI(
        int_data_y_1__5__2_), .SE(pe_1_0_5_n65), .CK(pe_1_0_5_net7107), .RN(
        pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_0_5_int_q_reg_h_reg_1__3_ ( .D(int_data_x_0__6__3_), .SI(
        int_data_y_1__5__3_), .SE(pe_1_0_5_n65), .CK(pe_1_0_5_net7107), .RN(
        pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_0_5_int_q_reg_h_reg_2__0_ ( .D(int_data_x_0__6__0_), .SI(
        int_data_y_1__5__0_), .SE(pe_1_0_5_n65), .CK(pe_1_0_5_net7112), .RN(
        pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_0_5_int_q_reg_h_reg_2__1_ ( .D(int_data_x_0__6__1_), .SI(
        int_data_y_1__5__1_), .SE(pe_1_0_5_n65), .CK(pe_1_0_5_net7112), .RN(
        pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_0_5_int_q_reg_h_reg_2__2_ ( .D(int_data_x_0__6__2_), .SI(
        int_data_y_1__5__2_), .SE(pe_1_0_5_n65), .CK(pe_1_0_5_net7112), .RN(
        pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_0_5_int_q_reg_h_reg_2__3_ ( .D(int_data_x_0__6__3_), .SI(
        int_data_y_1__5__3_), .SE(pe_1_0_5_n65), .CK(pe_1_0_5_net7112), .RN(
        pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_0_5_int_q_reg_h_reg_3__0_ ( .D(int_data_x_0__6__0_), .SI(
        int_data_y_1__5__0_), .SE(pe_1_0_5_n65), .CK(pe_1_0_5_net7117), .RN(
        pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_0_5_int_q_reg_h_reg_3__1_ ( .D(int_data_x_0__6__1_), .SI(
        int_data_y_1__5__1_), .SE(pe_1_0_5_n65), .CK(pe_1_0_5_net7117), .RN(
        pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_0_5_int_q_reg_h_reg_3__2_ ( .D(int_data_x_0__6__2_), .SI(
        int_data_y_1__5__2_), .SE(pe_1_0_5_n65), .CK(pe_1_0_5_net7117), .RN(
        pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_0_5_int_q_reg_h_reg_3__3_ ( .D(int_data_x_0__6__3_), .SI(
        int_data_y_1__5__3_), .SE(pe_1_0_5_n65), .CK(pe_1_0_5_net7117), .RN(
        pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_0_5_int_q_reg_h_reg_4__0_ ( .D(int_data_x_0__6__0_), .SI(
        int_data_y_1__5__0_), .SE(pe_1_0_5_n66), .CK(pe_1_0_5_net7122), .RN(
        pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_0_5_int_q_reg_h_reg_4__1_ ( .D(int_data_x_0__6__1_), .SI(
        int_data_y_1__5__1_), .SE(pe_1_0_5_n66), .CK(pe_1_0_5_net7122), .RN(
        pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_0_5_int_q_reg_h_reg_4__2_ ( .D(int_data_x_0__6__2_), .SI(
        int_data_y_1__5__2_), .SE(pe_1_0_5_n66), .CK(pe_1_0_5_net7122), .RN(
        pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_0_5_int_q_reg_h_reg_4__3_ ( .D(int_data_x_0__6__3_), .SI(
        int_data_y_1__5__3_), .SE(pe_1_0_5_n66), .CK(pe_1_0_5_net7122), .RN(
        pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_0_5_int_q_reg_h_reg_5__0_ ( .D(int_data_x_0__6__0_), .SI(
        int_data_y_1__5__0_), .SE(pe_1_0_5_n66), .CK(pe_1_0_5_net7127), .RN(
        pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_0_5_int_q_reg_h_reg_5__1_ ( .D(int_data_x_0__6__1_), .SI(
        int_data_y_1__5__1_), .SE(pe_1_0_5_n66), .CK(pe_1_0_5_net7127), .RN(
        pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_0_5_int_q_reg_h_reg_5__2_ ( .D(int_data_x_0__6__2_), .SI(
        int_data_y_1__5__2_), .SE(pe_1_0_5_n66), .CK(pe_1_0_5_net7127), .RN(
        pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_0_5_int_q_reg_h_reg_5__3_ ( .D(int_data_x_0__6__3_), .SI(
        int_data_y_1__5__3_), .SE(pe_1_0_5_n66), .CK(pe_1_0_5_net7127), .RN(
        pe_1_0_5_n72), .Q(pe_1_0_5_int_q_reg_h[3]) );
  FA_X1 pe_1_0_5_sub_81_U2_7 ( .A(o_data[23]), .B(pe_1_0_5_n76), .CI(
        pe_1_0_5_sub_81_carry[7]), .S(pe_1_0_5_N77) );
  FA_X1 pe_1_0_5_sub_81_U2_6 ( .A(o_data[22]), .B(pe_1_0_5_n76), .CI(
        pe_1_0_5_sub_81_carry[6]), .CO(pe_1_0_5_sub_81_carry[7]), .S(
        pe_1_0_5_N76) );
  FA_X1 pe_1_0_5_sub_81_U2_5 ( .A(o_data[21]), .B(pe_1_0_5_n76), .CI(
        pe_1_0_5_sub_81_carry[5]), .CO(pe_1_0_5_sub_81_carry[6]), .S(
        pe_1_0_5_N75) );
  FA_X1 pe_1_0_5_sub_81_U2_4 ( .A(o_data[20]), .B(pe_1_0_5_n76), .CI(
        pe_1_0_5_sub_81_carry[4]), .CO(pe_1_0_5_sub_81_carry[5]), .S(
        pe_1_0_5_N74) );
  FA_X1 pe_1_0_5_sub_81_U2_3 ( .A(o_data[19]), .B(pe_1_0_5_n76), .CI(
        pe_1_0_5_sub_81_carry[3]), .CO(pe_1_0_5_sub_81_carry[4]), .S(
        pe_1_0_5_N73) );
  FA_X1 pe_1_0_5_sub_81_U2_2 ( .A(o_data[18]), .B(pe_1_0_5_n75), .CI(
        pe_1_0_5_sub_81_carry[2]), .CO(pe_1_0_5_sub_81_carry[3]), .S(
        pe_1_0_5_N72) );
  FA_X1 pe_1_0_5_sub_81_U2_1 ( .A(o_data[17]), .B(pe_1_0_5_n74), .CI(
        pe_1_0_5_sub_81_carry[1]), .CO(pe_1_0_5_sub_81_carry[2]), .S(
        pe_1_0_5_N71) );
  FA_X1 pe_1_0_5_add_83_U1_7 ( .A(o_data[23]), .B(pe_1_0_5_int_data_3_), .CI(
        pe_1_0_5_add_83_carry[7]), .S(pe_1_0_5_N85) );
  FA_X1 pe_1_0_5_add_83_U1_6 ( .A(o_data[22]), .B(pe_1_0_5_int_data_3_), .CI(
        pe_1_0_5_add_83_carry[6]), .CO(pe_1_0_5_add_83_carry[7]), .S(
        pe_1_0_5_N84) );
  FA_X1 pe_1_0_5_add_83_U1_5 ( .A(o_data[21]), .B(pe_1_0_5_int_data_3_), .CI(
        pe_1_0_5_add_83_carry[5]), .CO(pe_1_0_5_add_83_carry[6]), .S(
        pe_1_0_5_N83) );
  FA_X1 pe_1_0_5_add_83_U1_4 ( .A(o_data[20]), .B(pe_1_0_5_int_data_3_), .CI(
        pe_1_0_5_add_83_carry[4]), .CO(pe_1_0_5_add_83_carry[5]), .S(
        pe_1_0_5_N82) );
  FA_X1 pe_1_0_5_add_83_U1_3 ( .A(o_data[19]), .B(pe_1_0_5_int_data_3_), .CI(
        pe_1_0_5_add_83_carry[3]), .CO(pe_1_0_5_add_83_carry[4]), .S(
        pe_1_0_5_N81) );
  FA_X1 pe_1_0_5_add_83_U1_2 ( .A(o_data[18]), .B(pe_1_0_5_int_data_2_), .CI(
        pe_1_0_5_add_83_carry[2]), .CO(pe_1_0_5_add_83_carry[3]), .S(
        pe_1_0_5_N80) );
  FA_X1 pe_1_0_5_add_83_U1_1 ( .A(o_data[17]), .B(pe_1_0_5_int_data_1_), .CI(
        pe_1_0_5_n2), .CO(pe_1_0_5_add_83_carry[2]), .S(pe_1_0_5_N79) );
  NAND3_X1 pe_1_0_5_U56 ( .A1(pe_1_0_5_n60), .A2(pe_1_0_5_n43), .A3(
        pe_1_0_5_n62), .ZN(pe_1_0_5_n40) );
  NAND3_X1 pe_1_0_5_U55 ( .A1(pe_1_0_5_n43), .A2(pe_1_0_5_n61), .A3(
        pe_1_0_5_n62), .ZN(pe_1_0_5_n39) );
  NAND3_X1 pe_1_0_5_U54 ( .A1(pe_1_0_5_n43), .A2(pe_1_0_5_n63), .A3(
        pe_1_0_5_n60), .ZN(pe_1_0_5_n38) );
  NAND3_X1 pe_1_0_5_U53 ( .A1(pe_1_0_5_n61), .A2(pe_1_0_5_n63), .A3(
        pe_1_0_5_n43), .ZN(pe_1_0_5_n37) );
  DFFR_X1 pe_1_0_5_int_q_acc_reg_6_ ( .D(pe_1_0_5_n78), .CK(pe_1_0_5_net7162), 
        .RN(pe_1_0_5_n71), .Q(o_data[22]) );
  DFFR_X1 pe_1_0_5_int_q_acc_reg_5_ ( .D(pe_1_0_5_n79), .CK(pe_1_0_5_net7162), 
        .RN(pe_1_0_5_n71), .Q(o_data[21]) );
  DFFR_X1 pe_1_0_5_int_q_acc_reg_4_ ( .D(pe_1_0_5_n80), .CK(pe_1_0_5_net7162), 
        .RN(pe_1_0_5_n71), .Q(o_data[20]) );
  DFFR_X1 pe_1_0_5_int_q_acc_reg_3_ ( .D(pe_1_0_5_n81), .CK(pe_1_0_5_net7162), 
        .RN(pe_1_0_5_n71), .Q(o_data[19]) );
  DFFR_X1 pe_1_0_5_int_q_acc_reg_2_ ( .D(pe_1_0_5_n82), .CK(pe_1_0_5_net7162), 
        .RN(pe_1_0_5_n71), .Q(o_data[18]) );
  DFFR_X1 pe_1_0_5_int_q_acc_reg_1_ ( .D(pe_1_0_5_n83), .CK(pe_1_0_5_net7162), 
        .RN(pe_1_0_5_n71), .Q(o_data[17]) );
  DFFR_X1 pe_1_0_5_int_q_acc_reg_7_ ( .D(pe_1_0_5_n77), .CK(pe_1_0_5_net7162), 
        .RN(pe_1_0_5_n71), .Q(o_data[23]) );
  CLKGATETST_X1 pe_1_0_5_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_0_5_n88), .SE(1'b0), .GCK(pe_1_0_5_net7101) );
  CLKGATETST_X1 pe_1_0_5_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_0_5_n87), .SE(1'b0), .GCK(pe_1_0_5_net7107) );
  CLKGATETST_X1 pe_1_0_5_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_0_5_n86), .SE(1'b0), .GCK(pe_1_0_5_net7112) );
  CLKGATETST_X1 pe_1_0_5_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_0_5_n85), .SE(1'b0), .GCK(pe_1_0_5_net7117) );
  CLKGATETST_X1 pe_1_0_5_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_0_5_n90), .SE(1'b0), .GCK(pe_1_0_5_net7122) );
  CLKGATETST_X1 pe_1_0_5_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_0_5_n89), .SE(1'b0), .GCK(pe_1_0_5_net7127) );
  CLKGATETST_X1 pe_1_0_5_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_0_5_N64), .SE(1'b0), .GCK(pe_1_0_5_net7132) );
  CLKGATETST_X1 pe_1_0_5_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_0_5_N63), .SE(1'b0), .GCK(pe_1_0_5_net7137) );
  CLKGATETST_X1 pe_1_0_5_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_0_5_N62), .SE(1'b0), .GCK(pe_1_0_5_net7142) );
  CLKGATETST_X1 pe_1_0_5_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_0_5_N61), .SE(1'b0), .GCK(pe_1_0_5_net7147) );
  CLKGATETST_X1 pe_1_0_5_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_0_5_N60), .SE(1'b0), .GCK(pe_1_0_5_net7152) );
  CLKGATETST_X1 pe_1_0_5_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_0_5_N59), .SE(1'b0), .GCK(pe_1_0_5_net7157) );
  CLKGATETST_X1 pe_1_0_5_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_0_5_N90), .SE(1'b0), .GCK(pe_1_0_5_net7162) );
  CLKBUF_X1 pe_1_0_6_U112 ( .A(pe_1_0_6_n72), .Z(pe_1_0_6_n71) );
  INV_X1 pe_1_0_6_U111 ( .A(n73), .ZN(pe_1_0_6_n70) );
  INV_X1 pe_1_0_6_U110 ( .A(n65), .ZN(pe_1_0_6_n69) );
  INV_X1 pe_1_0_6_U109 ( .A(n65), .ZN(pe_1_0_6_n68) );
  INV_X1 pe_1_0_6_U108 ( .A(n65), .ZN(pe_1_0_6_n67) );
  INV_X1 pe_1_0_6_U107 ( .A(pe_1_0_6_n69), .ZN(pe_1_0_6_n66) );
  INV_X1 pe_1_0_6_U106 ( .A(pe_1_0_6_n63), .ZN(pe_1_0_6_n62) );
  INV_X1 pe_1_0_6_U105 ( .A(pe_1_0_6_n61), .ZN(pe_1_0_6_n60) );
  INV_X1 pe_1_0_6_U104 ( .A(n25), .ZN(pe_1_0_6_n59) );
  INV_X1 pe_1_0_6_U103 ( .A(pe_1_0_6_n59), .ZN(pe_1_0_6_n58) );
  INV_X1 pe_1_0_6_U102 ( .A(n17), .ZN(pe_1_0_6_n57) );
  MUX2_X1 pe_1_0_6_U101 ( .A(pe_1_0_6_n54), .B(pe_1_0_6_n51), .S(n44), .Z(
        int_data_x_0__6__3_) );
  MUX2_X1 pe_1_0_6_U100 ( .A(pe_1_0_6_n53), .B(pe_1_0_6_n52), .S(pe_1_0_6_n62), 
        .Z(pe_1_0_6_n54) );
  MUX2_X1 pe_1_0_6_U99 ( .A(pe_1_0_6_int_q_reg_h[23]), .B(
        pe_1_0_6_int_q_reg_h[19]), .S(pe_1_0_6_n56), .Z(pe_1_0_6_n53) );
  MUX2_X1 pe_1_0_6_U98 ( .A(pe_1_0_6_int_q_reg_h[15]), .B(
        pe_1_0_6_int_q_reg_h[11]), .S(pe_1_0_6_n56), .Z(pe_1_0_6_n52) );
  MUX2_X1 pe_1_0_6_U97 ( .A(pe_1_0_6_int_q_reg_h[7]), .B(
        pe_1_0_6_int_q_reg_h[3]), .S(pe_1_0_6_n56), .Z(pe_1_0_6_n51) );
  MUX2_X1 pe_1_0_6_U96 ( .A(pe_1_0_6_n50), .B(pe_1_0_6_n47), .S(n44), .Z(
        int_data_x_0__6__2_) );
  MUX2_X1 pe_1_0_6_U95 ( .A(pe_1_0_6_n49), .B(pe_1_0_6_n48), .S(pe_1_0_6_n62), 
        .Z(pe_1_0_6_n50) );
  MUX2_X1 pe_1_0_6_U94 ( .A(pe_1_0_6_int_q_reg_h[22]), .B(
        pe_1_0_6_int_q_reg_h[18]), .S(pe_1_0_6_n56), .Z(pe_1_0_6_n49) );
  MUX2_X1 pe_1_0_6_U93 ( .A(pe_1_0_6_int_q_reg_h[14]), .B(
        pe_1_0_6_int_q_reg_h[10]), .S(pe_1_0_6_n56), .Z(pe_1_0_6_n48) );
  MUX2_X1 pe_1_0_6_U92 ( .A(pe_1_0_6_int_q_reg_h[6]), .B(
        pe_1_0_6_int_q_reg_h[2]), .S(pe_1_0_6_n56), .Z(pe_1_0_6_n47) );
  MUX2_X1 pe_1_0_6_U91 ( .A(pe_1_0_6_n46), .B(pe_1_0_6_n24), .S(n44), .Z(
        int_data_x_0__6__1_) );
  MUX2_X1 pe_1_0_6_U90 ( .A(pe_1_0_6_n45), .B(pe_1_0_6_n25), .S(pe_1_0_6_n62), 
        .Z(pe_1_0_6_n46) );
  MUX2_X1 pe_1_0_6_U89 ( .A(pe_1_0_6_int_q_reg_h[21]), .B(
        pe_1_0_6_int_q_reg_h[17]), .S(pe_1_0_6_n56), .Z(pe_1_0_6_n45) );
  MUX2_X1 pe_1_0_6_U88 ( .A(pe_1_0_6_int_q_reg_h[13]), .B(
        pe_1_0_6_int_q_reg_h[9]), .S(pe_1_0_6_n56), .Z(pe_1_0_6_n25) );
  MUX2_X1 pe_1_0_6_U87 ( .A(pe_1_0_6_int_q_reg_h[5]), .B(
        pe_1_0_6_int_q_reg_h[1]), .S(pe_1_0_6_n56), .Z(pe_1_0_6_n24) );
  MUX2_X1 pe_1_0_6_U86 ( .A(pe_1_0_6_n23), .B(pe_1_0_6_n20), .S(n44), .Z(
        int_data_x_0__6__0_) );
  MUX2_X1 pe_1_0_6_U85 ( .A(pe_1_0_6_n22), .B(pe_1_0_6_n21), .S(pe_1_0_6_n62), 
        .Z(pe_1_0_6_n23) );
  MUX2_X1 pe_1_0_6_U84 ( .A(pe_1_0_6_int_q_reg_h[20]), .B(
        pe_1_0_6_int_q_reg_h[16]), .S(pe_1_0_6_n56), .Z(pe_1_0_6_n22) );
  MUX2_X1 pe_1_0_6_U83 ( .A(pe_1_0_6_int_q_reg_h[12]), .B(
        pe_1_0_6_int_q_reg_h[8]), .S(pe_1_0_6_n56), .Z(pe_1_0_6_n21) );
  MUX2_X1 pe_1_0_6_U82 ( .A(pe_1_0_6_int_q_reg_h[4]), .B(
        pe_1_0_6_int_q_reg_h[0]), .S(pe_1_0_6_n56), .Z(pe_1_0_6_n20) );
  MUX2_X1 pe_1_0_6_U81 ( .A(pe_1_0_6_n19), .B(pe_1_0_6_n16), .S(n44), .Z(
        pe_1_0_6_o_data_v_3_) );
  MUX2_X1 pe_1_0_6_U80 ( .A(pe_1_0_6_n18), .B(pe_1_0_6_n17), .S(pe_1_0_6_n62), 
        .Z(pe_1_0_6_n19) );
  MUX2_X1 pe_1_0_6_U79 ( .A(pe_1_0_6_int_q_reg_v[23]), .B(
        pe_1_0_6_int_q_reg_v[19]), .S(pe_1_0_6_n55), .Z(pe_1_0_6_n18) );
  MUX2_X1 pe_1_0_6_U78 ( .A(pe_1_0_6_int_q_reg_v[15]), .B(
        pe_1_0_6_int_q_reg_v[11]), .S(pe_1_0_6_n55), .Z(pe_1_0_6_n17) );
  MUX2_X1 pe_1_0_6_U77 ( .A(pe_1_0_6_int_q_reg_v[7]), .B(
        pe_1_0_6_int_q_reg_v[3]), .S(pe_1_0_6_n55), .Z(pe_1_0_6_n16) );
  MUX2_X1 pe_1_0_6_U76 ( .A(pe_1_0_6_n15), .B(pe_1_0_6_n12), .S(n44), .Z(
        pe_1_0_6_o_data_v_2_) );
  MUX2_X1 pe_1_0_6_U75 ( .A(pe_1_0_6_n14), .B(pe_1_0_6_n13), .S(pe_1_0_6_n62), 
        .Z(pe_1_0_6_n15) );
  MUX2_X1 pe_1_0_6_U74 ( .A(pe_1_0_6_int_q_reg_v[22]), .B(
        pe_1_0_6_int_q_reg_v[18]), .S(pe_1_0_6_n55), .Z(pe_1_0_6_n14) );
  MUX2_X1 pe_1_0_6_U73 ( .A(pe_1_0_6_int_q_reg_v[14]), .B(
        pe_1_0_6_int_q_reg_v[10]), .S(pe_1_0_6_n55), .Z(pe_1_0_6_n13) );
  MUX2_X1 pe_1_0_6_U72 ( .A(pe_1_0_6_int_q_reg_v[6]), .B(
        pe_1_0_6_int_q_reg_v[2]), .S(pe_1_0_6_n55), .Z(pe_1_0_6_n12) );
  MUX2_X1 pe_1_0_6_U71 ( .A(pe_1_0_6_n11), .B(pe_1_0_6_n8), .S(n44), .Z(
        pe_1_0_6_o_data_v_1_) );
  MUX2_X1 pe_1_0_6_U70 ( .A(pe_1_0_6_n10), .B(pe_1_0_6_n9), .S(pe_1_0_6_n62), 
        .Z(pe_1_0_6_n11) );
  MUX2_X1 pe_1_0_6_U69 ( .A(pe_1_0_6_int_q_reg_v[21]), .B(
        pe_1_0_6_int_q_reg_v[17]), .S(pe_1_0_6_n55), .Z(pe_1_0_6_n10) );
  MUX2_X1 pe_1_0_6_U68 ( .A(pe_1_0_6_int_q_reg_v[13]), .B(
        pe_1_0_6_int_q_reg_v[9]), .S(pe_1_0_6_n55), .Z(pe_1_0_6_n9) );
  MUX2_X1 pe_1_0_6_U67 ( .A(pe_1_0_6_int_q_reg_v[5]), .B(
        pe_1_0_6_int_q_reg_v[1]), .S(pe_1_0_6_n55), .Z(pe_1_0_6_n8) );
  MUX2_X1 pe_1_0_6_U66 ( .A(pe_1_0_6_n7), .B(pe_1_0_6_n4), .S(n44), .Z(
        pe_1_0_6_o_data_v_0_) );
  MUX2_X1 pe_1_0_6_U65 ( .A(pe_1_0_6_n6), .B(pe_1_0_6_n5), .S(pe_1_0_6_n62), 
        .Z(pe_1_0_6_n7) );
  MUX2_X1 pe_1_0_6_U64 ( .A(pe_1_0_6_int_q_reg_v[20]), .B(
        pe_1_0_6_int_q_reg_v[16]), .S(pe_1_0_6_n55), .Z(pe_1_0_6_n6) );
  MUX2_X1 pe_1_0_6_U63 ( .A(pe_1_0_6_int_q_reg_v[12]), .B(
        pe_1_0_6_int_q_reg_v[8]), .S(pe_1_0_6_n55), .Z(pe_1_0_6_n5) );
  MUX2_X1 pe_1_0_6_U62 ( .A(pe_1_0_6_int_q_reg_v[4]), .B(
        pe_1_0_6_int_q_reg_v[0]), .S(pe_1_0_6_n55), .Z(pe_1_0_6_n4) );
  XNOR2_X1 pe_1_0_6_U61 ( .A(pe_1_0_6_n73), .B(o_data[8]), .ZN(pe_1_0_6_N70)
         );
  AOI222_X1 pe_1_0_6_U60 ( .A1(int_data_res_1__6__0_), .A2(pe_1_0_6_n64), .B1(
        pe_1_0_6_n1), .B2(pe_1_0_6_n27), .C1(pe_1_0_6_N70), .C2(pe_1_0_6_n28), 
        .ZN(pe_1_0_6_n35) );
  INV_X1 pe_1_0_6_U59 ( .A(pe_1_0_6_n35), .ZN(pe_1_0_6_n84) );
  AOI222_X1 pe_1_0_6_U58 ( .A1(int_data_res_1__6__2_), .A2(pe_1_0_6_n64), .B1(
        pe_1_0_6_N80), .B2(pe_1_0_6_n27), .C1(pe_1_0_6_N72), .C2(pe_1_0_6_n28), 
        .ZN(pe_1_0_6_n33) );
  INV_X1 pe_1_0_6_U57 ( .A(pe_1_0_6_n33), .ZN(pe_1_0_6_n82) );
  AOI222_X1 pe_1_0_6_U52 ( .A1(int_data_res_1__6__6_), .A2(pe_1_0_6_n64), .B1(
        pe_1_0_6_N84), .B2(pe_1_0_6_n27), .C1(pe_1_0_6_N76), .C2(pe_1_0_6_n28), 
        .ZN(pe_1_0_6_n29) );
  INV_X1 pe_1_0_6_U51 ( .A(pe_1_0_6_n29), .ZN(pe_1_0_6_n78) );
  AOI222_X1 pe_1_0_6_U50 ( .A1(int_data_res_1__6__1_), .A2(pe_1_0_6_n64), .B1(
        pe_1_0_6_N79), .B2(pe_1_0_6_n27), .C1(pe_1_0_6_N71), .C2(pe_1_0_6_n28), 
        .ZN(pe_1_0_6_n34) );
  INV_X1 pe_1_0_6_U49 ( .A(pe_1_0_6_n34), .ZN(pe_1_0_6_n83) );
  AOI222_X1 pe_1_0_6_U48 ( .A1(int_data_res_1__6__3_), .A2(pe_1_0_6_n64), .B1(
        pe_1_0_6_N81), .B2(pe_1_0_6_n27), .C1(pe_1_0_6_N73), .C2(pe_1_0_6_n28), 
        .ZN(pe_1_0_6_n32) );
  INV_X1 pe_1_0_6_U47 ( .A(pe_1_0_6_n32), .ZN(pe_1_0_6_n81) );
  AOI222_X1 pe_1_0_6_U46 ( .A1(int_data_res_1__6__4_), .A2(pe_1_0_6_n64), .B1(
        pe_1_0_6_N82), .B2(pe_1_0_6_n27), .C1(pe_1_0_6_N74), .C2(pe_1_0_6_n28), 
        .ZN(pe_1_0_6_n31) );
  INV_X1 pe_1_0_6_U45 ( .A(pe_1_0_6_n31), .ZN(pe_1_0_6_n80) );
  AOI222_X1 pe_1_0_6_U44 ( .A1(int_data_res_1__6__5_), .A2(pe_1_0_6_n64), .B1(
        pe_1_0_6_N83), .B2(pe_1_0_6_n27), .C1(pe_1_0_6_N75), .C2(pe_1_0_6_n28), 
        .ZN(pe_1_0_6_n30) );
  INV_X1 pe_1_0_6_U43 ( .A(pe_1_0_6_n30), .ZN(pe_1_0_6_n79) );
  INV_X1 pe_1_0_6_U42 ( .A(pe_1_0_6_int_data_2_), .ZN(pe_1_0_6_n75) );
  NAND2_X1 pe_1_0_6_U41 ( .A1(pe_1_0_6_int_data_0_), .A2(pe_1_0_6_n3), .ZN(
        pe_1_0_6_sub_81_carry[1]) );
  INV_X1 pe_1_0_6_U40 ( .A(pe_1_0_6_int_data_1_), .ZN(pe_1_0_6_n74) );
  AND2_X1 pe_1_0_6_U39 ( .A1(pe_1_0_6_int_data_0_), .A2(o_data[8]), .ZN(
        pe_1_0_6_n2) );
  AOI222_X1 pe_1_0_6_U38 ( .A1(pe_1_0_6_n64), .A2(int_data_res_1__6__7_), .B1(
        pe_1_0_6_N85), .B2(pe_1_0_6_n27), .C1(pe_1_0_6_N77), .C2(pe_1_0_6_n28), 
        .ZN(pe_1_0_6_n26) );
  INV_X1 pe_1_0_6_U37 ( .A(pe_1_0_6_n26), .ZN(pe_1_0_6_n77) );
  NOR3_X1 pe_1_0_6_U36 ( .A1(pe_1_0_6_n59), .A2(pe_1_0_6_n65), .A3(int_ckg[57]), .ZN(pe_1_0_6_n36) );
  OR2_X1 pe_1_0_6_U35 ( .A1(pe_1_0_6_n36), .A2(pe_1_0_6_n64), .ZN(pe_1_0_6_N90) );
  INV_X1 pe_1_0_6_U34 ( .A(n37), .ZN(pe_1_0_6_n63) );
  AND2_X1 pe_1_0_6_U33 ( .A1(int_data_x_0__6__2_), .A2(pe_1_0_6_n58), .ZN(
        pe_1_0_6_int_data_2_) );
  AND2_X1 pe_1_0_6_U32 ( .A1(int_data_x_0__6__1_), .A2(pe_1_0_6_n58), .ZN(
        pe_1_0_6_int_data_1_) );
  AND2_X1 pe_1_0_6_U31 ( .A1(int_data_x_0__6__3_), .A2(pe_1_0_6_n58), .ZN(
        pe_1_0_6_int_data_3_) );
  BUF_X1 pe_1_0_6_U30 ( .A(n59), .Z(pe_1_0_6_n64) );
  INV_X1 pe_1_0_6_U29 ( .A(n31), .ZN(pe_1_0_6_n61) );
  AND2_X1 pe_1_0_6_U28 ( .A1(int_data_x_0__6__0_), .A2(pe_1_0_6_n58), .ZN(
        pe_1_0_6_int_data_0_) );
  NAND2_X1 pe_1_0_6_U27 ( .A1(pe_1_0_6_n44), .A2(pe_1_0_6_n61), .ZN(
        pe_1_0_6_n41) );
  AND3_X1 pe_1_0_6_U26 ( .A1(n73), .A2(pe_1_0_6_n63), .A3(n44), .ZN(
        pe_1_0_6_n44) );
  INV_X1 pe_1_0_6_U25 ( .A(pe_1_0_6_int_data_3_), .ZN(pe_1_0_6_n76) );
  NOR2_X1 pe_1_0_6_U24 ( .A1(pe_1_0_6_n70), .A2(n44), .ZN(pe_1_0_6_n43) );
  NOR2_X1 pe_1_0_6_U23 ( .A1(pe_1_0_6_n57), .A2(pe_1_0_6_n64), .ZN(
        pe_1_0_6_n28) );
  NOR2_X1 pe_1_0_6_U22 ( .A1(n17), .A2(pe_1_0_6_n64), .ZN(pe_1_0_6_n27) );
  INV_X1 pe_1_0_6_U21 ( .A(pe_1_0_6_int_data_0_), .ZN(pe_1_0_6_n73) );
  BUF_X1 pe_1_0_6_U20 ( .A(pe_1_0_6_n60), .Z(pe_1_0_6_n55) );
  INV_X1 pe_1_0_6_U19 ( .A(pe_1_0_6_n41), .ZN(pe_1_0_6_n90) );
  INV_X1 pe_1_0_6_U18 ( .A(pe_1_0_6_n37), .ZN(pe_1_0_6_n88) );
  INV_X1 pe_1_0_6_U17 ( .A(pe_1_0_6_n38), .ZN(pe_1_0_6_n87) );
  INV_X1 pe_1_0_6_U16 ( .A(pe_1_0_6_n39), .ZN(pe_1_0_6_n86) );
  NOR2_X1 pe_1_0_6_U15 ( .A1(pe_1_0_6_n68), .A2(pe_1_0_6_n42), .ZN(
        pe_1_0_6_N59) );
  NOR2_X1 pe_1_0_6_U14 ( .A1(pe_1_0_6_n68), .A2(pe_1_0_6_n41), .ZN(
        pe_1_0_6_N60) );
  NOR2_X1 pe_1_0_6_U13 ( .A1(pe_1_0_6_n68), .A2(pe_1_0_6_n38), .ZN(
        pe_1_0_6_N63) );
  NOR2_X1 pe_1_0_6_U12 ( .A1(pe_1_0_6_n67), .A2(pe_1_0_6_n40), .ZN(
        pe_1_0_6_N61) );
  NOR2_X1 pe_1_0_6_U11 ( .A1(pe_1_0_6_n67), .A2(pe_1_0_6_n39), .ZN(
        pe_1_0_6_N62) );
  NOR2_X1 pe_1_0_6_U10 ( .A1(pe_1_0_6_n37), .A2(pe_1_0_6_n67), .ZN(
        pe_1_0_6_N64) );
  NAND2_X1 pe_1_0_6_U9 ( .A1(pe_1_0_6_n44), .A2(pe_1_0_6_n60), .ZN(
        pe_1_0_6_n42) );
  INV_X1 pe_1_0_6_U8 ( .A(pe_1_0_6_n69), .ZN(pe_1_0_6_n65) );
  BUF_X1 pe_1_0_6_U7 ( .A(pe_1_0_6_n60), .Z(pe_1_0_6_n56) );
  INV_X1 pe_1_0_6_U6 ( .A(pe_1_0_6_n42), .ZN(pe_1_0_6_n89) );
  INV_X1 pe_1_0_6_U5 ( .A(pe_1_0_6_n40), .ZN(pe_1_0_6_n85) );
  INV_X2 pe_1_0_6_U4 ( .A(n81), .ZN(pe_1_0_6_n72) );
  XOR2_X1 pe_1_0_6_U3 ( .A(pe_1_0_6_int_data_0_), .B(o_data[8]), .Z(
        pe_1_0_6_n1) );
  DFFR_X1 pe_1_0_6_int_q_acc_reg_0_ ( .D(pe_1_0_6_n84), .CK(pe_1_0_6_net7084), 
        .RN(pe_1_0_6_n72), .Q(o_data[8]), .QN(pe_1_0_6_n3) );
  DFFR_X1 pe_1_0_6_int_q_reg_v_reg_0__0_ ( .D(int_data_y_1__6__0_), .CK(
        pe_1_0_6_net7054), .RN(pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_v[20]) );
  DFFR_X1 pe_1_0_6_int_q_reg_v_reg_0__1_ ( .D(int_data_y_1__6__1_), .CK(
        pe_1_0_6_net7054), .RN(pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_v[21]) );
  DFFR_X1 pe_1_0_6_int_q_reg_v_reg_0__2_ ( .D(int_data_y_1__6__2_), .CK(
        pe_1_0_6_net7054), .RN(pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_v[22]) );
  DFFR_X1 pe_1_0_6_int_q_reg_v_reg_0__3_ ( .D(int_data_y_1__6__3_), .CK(
        pe_1_0_6_net7054), .RN(pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_v[23]) );
  DFFR_X1 pe_1_0_6_int_q_reg_v_reg_1__0_ ( .D(int_data_y_1__6__0_), .CK(
        pe_1_0_6_net7059), .RN(pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_v[16]) );
  DFFR_X1 pe_1_0_6_int_q_reg_v_reg_1__1_ ( .D(int_data_y_1__6__1_), .CK(
        pe_1_0_6_net7059), .RN(pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_v[17]) );
  DFFR_X1 pe_1_0_6_int_q_reg_v_reg_1__2_ ( .D(int_data_y_1__6__2_), .CK(
        pe_1_0_6_net7059), .RN(pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_v[18]) );
  DFFR_X1 pe_1_0_6_int_q_reg_v_reg_1__3_ ( .D(int_data_y_1__6__3_), .CK(
        pe_1_0_6_net7059), .RN(pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_v[19]) );
  DFFR_X1 pe_1_0_6_int_q_reg_v_reg_2__0_ ( .D(int_data_y_1__6__0_), .CK(
        pe_1_0_6_net7064), .RN(pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_v[12]) );
  DFFR_X1 pe_1_0_6_int_q_reg_v_reg_2__1_ ( .D(int_data_y_1__6__1_), .CK(
        pe_1_0_6_net7064), .RN(pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_v[13]) );
  DFFR_X1 pe_1_0_6_int_q_reg_v_reg_2__2_ ( .D(int_data_y_1__6__2_), .CK(
        pe_1_0_6_net7064), .RN(pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_v[14]) );
  DFFR_X1 pe_1_0_6_int_q_reg_v_reg_2__3_ ( .D(int_data_y_1__6__3_), .CK(
        pe_1_0_6_net7064), .RN(pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_v[15]) );
  DFFR_X1 pe_1_0_6_int_q_reg_v_reg_3__0_ ( .D(int_data_y_1__6__0_), .CK(
        pe_1_0_6_net7069), .RN(pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_v[8]) );
  DFFR_X1 pe_1_0_6_int_q_reg_v_reg_3__1_ ( .D(int_data_y_1__6__1_), .CK(
        pe_1_0_6_net7069), .RN(pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_v[9]) );
  DFFR_X1 pe_1_0_6_int_q_reg_v_reg_3__2_ ( .D(int_data_y_1__6__2_), .CK(
        pe_1_0_6_net7069), .RN(pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_v[10]) );
  DFFR_X1 pe_1_0_6_int_q_reg_v_reg_3__3_ ( .D(int_data_y_1__6__3_), .CK(
        pe_1_0_6_net7069), .RN(pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_v[11]) );
  DFFR_X1 pe_1_0_6_int_q_reg_v_reg_4__0_ ( .D(int_data_y_1__6__0_), .CK(
        pe_1_0_6_net7074), .RN(pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_v[4]) );
  DFFR_X1 pe_1_0_6_int_q_reg_v_reg_4__1_ ( .D(int_data_y_1__6__1_), .CK(
        pe_1_0_6_net7074), .RN(pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_v[5]) );
  DFFR_X1 pe_1_0_6_int_q_reg_v_reg_4__2_ ( .D(int_data_y_1__6__2_), .CK(
        pe_1_0_6_net7074), .RN(pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_v[6]) );
  DFFR_X1 pe_1_0_6_int_q_reg_v_reg_4__3_ ( .D(int_data_y_1__6__3_), .CK(
        pe_1_0_6_net7074), .RN(pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_v[7]) );
  DFFR_X1 pe_1_0_6_int_q_reg_v_reg_5__0_ ( .D(int_data_y_1__6__0_), .CK(
        pe_1_0_6_net7079), .RN(pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_v[0]) );
  DFFR_X1 pe_1_0_6_int_q_reg_v_reg_5__1_ ( .D(int_data_y_1__6__1_), .CK(
        pe_1_0_6_net7079), .RN(pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_v[1]) );
  DFFR_X1 pe_1_0_6_int_q_reg_v_reg_5__2_ ( .D(int_data_y_1__6__2_), .CK(
        pe_1_0_6_net7079), .RN(pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_v[2]) );
  DFFR_X1 pe_1_0_6_int_q_reg_v_reg_5__3_ ( .D(int_data_y_1__6__3_), .CK(
        pe_1_0_6_net7079), .RN(pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_0_6_int_q_reg_h_reg_0__0_ ( .D(int_data_x_0__7__0_), .SI(
        int_data_y_1__6__0_), .SE(pe_1_0_6_n65), .CK(pe_1_0_6_net7023), .RN(
        pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_0_6_int_q_reg_h_reg_0__1_ ( .D(int_data_x_0__7__1_), .SI(
        int_data_y_1__6__1_), .SE(pe_1_0_6_n65), .CK(pe_1_0_6_net7023), .RN(
        pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_0_6_int_q_reg_h_reg_0__2_ ( .D(int_data_x_0__7__2_), .SI(
        int_data_y_1__6__2_), .SE(pe_1_0_6_n65), .CK(pe_1_0_6_net7023), .RN(
        pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_0_6_int_q_reg_h_reg_0__3_ ( .D(int_data_x_0__7__3_), .SI(
        int_data_y_1__6__3_), .SE(pe_1_0_6_n65), .CK(pe_1_0_6_net7023), .RN(
        pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_0_6_int_q_reg_h_reg_1__0_ ( .D(int_data_x_0__7__0_), .SI(
        int_data_y_1__6__0_), .SE(pe_1_0_6_n65), .CK(pe_1_0_6_net7029), .RN(
        pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_0_6_int_q_reg_h_reg_1__1_ ( .D(int_data_x_0__7__1_), .SI(
        int_data_y_1__6__1_), .SE(pe_1_0_6_n65), .CK(pe_1_0_6_net7029), .RN(
        pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_0_6_int_q_reg_h_reg_1__2_ ( .D(int_data_x_0__7__2_), .SI(
        int_data_y_1__6__2_), .SE(pe_1_0_6_n65), .CK(pe_1_0_6_net7029), .RN(
        pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_0_6_int_q_reg_h_reg_1__3_ ( .D(int_data_x_0__7__3_), .SI(
        int_data_y_1__6__3_), .SE(pe_1_0_6_n65), .CK(pe_1_0_6_net7029), .RN(
        pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_0_6_int_q_reg_h_reg_2__0_ ( .D(int_data_x_0__7__0_), .SI(
        int_data_y_1__6__0_), .SE(pe_1_0_6_n65), .CK(pe_1_0_6_net7034), .RN(
        pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_0_6_int_q_reg_h_reg_2__1_ ( .D(int_data_x_0__7__1_), .SI(
        int_data_y_1__6__1_), .SE(pe_1_0_6_n65), .CK(pe_1_0_6_net7034), .RN(
        pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_0_6_int_q_reg_h_reg_2__2_ ( .D(int_data_x_0__7__2_), .SI(
        int_data_y_1__6__2_), .SE(pe_1_0_6_n65), .CK(pe_1_0_6_net7034), .RN(
        pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_0_6_int_q_reg_h_reg_2__3_ ( .D(int_data_x_0__7__3_), .SI(
        int_data_y_1__6__3_), .SE(pe_1_0_6_n65), .CK(pe_1_0_6_net7034), .RN(
        pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_0_6_int_q_reg_h_reg_3__0_ ( .D(int_data_x_0__7__0_), .SI(
        int_data_y_1__6__0_), .SE(pe_1_0_6_n65), .CK(pe_1_0_6_net7039), .RN(
        pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_0_6_int_q_reg_h_reg_3__1_ ( .D(int_data_x_0__7__1_), .SI(
        int_data_y_1__6__1_), .SE(pe_1_0_6_n65), .CK(pe_1_0_6_net7039), .RN(
        pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_0_6_int_q_reg_h_reg_3__2_ ( .D(int_data_x_0__7__2_), .SI(
        int_data_y_1__6__2_), .SE(pe_1_0_6_n65), .CK(pe_1_0_6_net7039), .RN(
        pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_0_6_int_q_reg_h_reg_3__3_ ( .D(int_data_x_0__7__3_), .SI(
        int_data_y_1__6__3_), .SE(pe_1_0_6_n65), .CK(pe_1_0_6_net7039), .RN(
        pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_0_6_int_q_reg_h_reg_4__0_ ( .D(int_data_x_0__7__0_), .SI(
        int_data_y_1__6__0_), .SE(pe_1_0_6_n66), .CK(pe_1_0_6_net7044), .RN(
        pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_0_6_int_q_reg_h_reg_4__1_ ( .D(int_data_x_0__7__1_), .SI(
        int_data_y_1__6__1_), .SE(pe_1_0_6_n66), .CK(pe_1_0_6_net7044), .RN(
        pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_0_6_int_q_reg_h_reg_4__2_ ( .D(int_data_x_0__7__2_), .SI(
        int_data_y_1__6__2_), .SE(pe_1_0_6_n66), .CK(pe_1_0_6_net7044), .RN(
        pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_0_6_int_q_reg_h_reg_4__3_ ( .D(int_data_x_0__7__3_), .SI(
        int_data_y_1__6__3_), .SE(pe_1_0_6_n66), .CK(pe_1_0_6_net7044), .RN(
        pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_0_6_int_q_reg_h_reg_5__0_ ( .D(int_data_x_0__7__0_), .SI(
        int_data_y_1__6__0_), .SE(pe_1_0_6_n66), .CK(pe_1_0_6_net7049), .RN(
        pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_0_6_int_q_reg_h_reg_5__1_ ( .D(int_data_x_0__7__1_), .SI(
        int_data_y_1__6__1_), .SE(pe_1_0_6_n66), .CK(pe_1_0_6_net7049), .RN(
        pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_0_6_int_q_reg_h_reg_5__2_ ( .D(int_data_x_0__7__2_), .SI(
        int_data_y_1__6__2_), .SE(pe_1_0_6_n66), .CK(pe_1_0_6_net7049), .RN(
        pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_0_6_int_q_reg_h_reg_5__3_ ( .D(int_data_x_0__7__3_), .SI(
        int_data_y_1__6__3_), .SE(pe_1_0_6_n66), .CK(pe_1_0_6_net7049), .RN(
        pe_1_0_6_n72), .Q(pe_1_0_6_int_q_reg_h[3]) );
  FA_X1 pe_1_0_6_sub_81_U2_7 ( .A(o_data[15]), .B(pe_1_0_6_n76), .CI(
        pe_1_0_6_sub_81_carry[7]), .S(pe_1_0_6_N77) );
  FA_X1 pe_1_0_6_sub_81_U2_6 ( .A(o_data[14]), .B(pe_1_0_6_n76), .CI(
        pe_1_0_6_sub_81_carry[6]), .CO(pe_1_0_6_sub_81_carry[7]), .S(
        pe_1_0_6_N76) );
  FA_X1 pe_1_0_6_sub_81_U2_5 ( .A(o_data[13]), .B(pe_1_0_6_n76), .CI(
        pe_1_0_6_sub_81_carry[5]), .CO(pe_1_0_6_sub_81_carry[6]), .S(
        pe_1_0_6_N75) );
  FA_X1 pe_1_0_6_sub_81_U2_4 ( .A(o_data[12]), .B(pe_1_0_6_n76), .CI(
        pe_1_0_6_sub_81_carry[4]), .CO(pe_1_0_6_sub_81_carry[5]), .S(
        pe_1_0_6_N74) );
  FA_X1 pe_1_0_6_sub_81_U2_3 ( .A(o_data[11]), .B(pe_1_0_6_n76), .CI(
        pe_1_0_6_sub_81_carry[3]), .CO(pe_1_0_6_sub_81_carry[4]), .S(
        pe_1_0_6_N73) );
  FA_X1 pe_1_0_6_sub_81_U2_2 ( .A(o_data[10]), .B(pe_1_0_6_n75), .CI(
        pe_1_0_6_sub_81_carry[2]), .CO(pe_1_0_6_sub_81_carry[3]), .S(
        pe_1_0_6_N72) );
  FA_X1 pe_1_0_6_sub_81_U2_1 ( .A(o_data[9]), .B(pe_1_0_6_n74), .CI(
        pe_1_0_6_sub_81_carry[1]), .CO(pe_1_0_6_sub_81_carry[2]), .S(
        pe_1_0_6_N71) );
  FA_X1 pe_1_0_6_add_83_U1_7 ( .A(o_data[15]), .B(pe_1_0_6_int_data_3_), .CI(
        pe_1_0_6_add_83_carry[7]), .S(pe_1_0_6_N85) );
  FA_X1 pe_1_0_6_add_83_U1_6 ( .A(o_data[14]), .B(pe_1_0_6_int_data_3_), .CI(
        pe_1_0_6_add_83_carry[6]), .CO(pe_1_0_6_add_83_carry[7]), .S(
        pe_1_0_6_N84) );
  FA_X1 pe_1_0_6_add_83_U1_5 ( .A(o_data[13]), .B(pe_1_0_6_int_data_3_), .CI(
        pe_1_0_6_add_83_carry[5]), .CO(pe_1_0_6_add_83_carry[6]), .S(
        pe_1_0_6_N83) );
  FA_X1 pe_1_0_6_add_83_U1_4 ( .A(o_data[12]), .B(pe_1_0_6_int_data_3_), .CI(
        pe_1_0_6_add_83_carry[4]), .CO(pe_1_0_6_add_83_carry[5]), .S(
        pe_1_0_6_N82) );
  FA_X1 pe_1_0_6_add_83_U1_3 ( .A(o_data[11]), .B(pe_1_0_6_int_data_3_), .CI(
        pe_1_0_6_add_83_carry[3]), .CO(pe_1_0_6_add_83_carry[4]), .S(
        pe_1_0_6_N81) );
  FA_X1 pe_1_0_6_add_83_U1_2 ( .A(o_data[10]), .B(pe_1_0_6_int_data_2_), .CI(
        pe_1_0_6_add_83_carry[2]), .CO(pe_1_0_6_add_83_carry[3]), .S(
        pe_1_0_6_N80) );
  FA_X1 pe_1_0_6_add_83_U1_1 ( .A(o_data[9]), .B(pe_1_0_6_int_data_1_), .CI(
        pe_1_0_6_n2), .CO(pe_1_0_6_add_83_carry[2]), .S(pe_1_0_6_N79) );
  NAND3_X1 pe_1_0_6_U56 ( .A1(pe_1_0_6_n60), .A2(pe_1_0_6_n43), .A3(
        pe_1_0_6_n62), .ZN(pe_1_0_6_n40) );
  NAND3_X1 pe_1_0_6_U55 ( .A1(pe_1_0_6_n43), .A2(pe_1_0_6_n61), .A3(
        pe_1_0_6_n62), .ZN(pe_1_0_6_n39) );
  NAND3_X1 pe_1_0_6_U54 ( .A1(pe_1_0_6_n43), .A2(pe_1_0_6_n63), .A3(
        pe_1_0_6_n60), .ZN(pe_1_0_6_n38) );
  NAND3_X1 pe_1_0_6_U53 ( .A1(pe_1_0_6_n61), .A2(pe_1_0_6_n63), .A3(
        pe_1_0_6_n43), .ZN(pe_1_0_6_n37) );
  DFFR_X1 pe_1_0_6_int_q_acc_reg_6_ ( .D(pe_1_0_6_n78), .CK(pe_1_0_6_net7084), 
        .RN(pe_1_0_6_n71), .Q(o_data[14]) );
  DFFR_X1 pe_1_0_6_int_q_acc_reg_5_ ( .D(pe_1_0_6_n79), .CK(pe_1_0_6_net7084), 
        .RN(pe_1_0_6_n71), .Q(o_data[13]) );
  DFFR_X1 pe_1_0_6_int_q_acc_reg_4_ ( .D(pe_1_0_6_n80), .CK(pe_1_0_6_net7084), 
        .RN(pe_1_0_6_n71), .Q(o_data[12]) );
  DFFR_X1 pe_1_0_6_int_q_acc_reg_3_ ( .D(pe_1_0_6_n81), .CK(pe_1_0_6_net7084), 
        .RN(pe_1_0_6_n71), .Q(o_data[11]) );
  DFFR_X1 pe_1_0_6_int_q_acc_reg_2_ ( .D(pe_1_0_6_n82), .CK(pe_1_0_6_net7084), 
        .RN(pe_1_0_6_n71), .Q(o_data[10]) );
  DFFR_X1 pe_1_0_6_int_q_acc_reg_1_ ( .D(pe_1_0_6_n83), .CK(pe_1_0_6_net7084), 
        .RN(pe_1_0_6_n71), .Q(o_data[9]) );
  DFFR_X1 pe_1_0_6_int_q_acc_reg_7_ ( .D(pe_1_0_6_n77), .CK(pe_1_0_6_net7084), 
        .RN(pe_1_0_6_n71), .Q(o_data[15]) );
  CLKGATETST_X1 pe_1_0_6_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_0_6_n88), .SE(1'b0), .GCK(pe_1_0_6_net7023) );
  CLKGATETST_X1 pe_1_0_6_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_0_6_n87), .SE(1'b0), .GCK(pe_1_0_6_net7029) );
  CLKGATETST_X1 pe_1_0_6_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_0_6_n86), .SE(1'b0), .GCK(pe_1_0_6_net7034) );
  CLKGATETST_X1 pe_1_0_6_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_0_6_n85), .SE(1'b0), .GCK(pe_1_0_6_net7039) );
  CLKGATETST_X1 pe_1_0_6_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_0_6_n90), .SE(1'b0), .GCK(pe_1_0_6_net7044) );
  CLKGATETST_X1 pe_1_0_6_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_0_6_n89), .SE(1'b0), .GCK(pe_1_0_6_net7049) );
  CLKGATETST_X1 pe_1_0_6_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_0_6_N64), .SE(1'b0), .GCK(pe_1_0_6_net7054) );
  CLKGATETST_X1 pe_1_0_6_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_0_6_N63), .SE(1'b0), .GCK(pe_1_0_6_net7059) );
  CLKGATETST_X1 pe_1_0_6_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_0_6_N62), .SE(1'b0), .GCK(pe_1_0_6_net7064) );
  CLKGATETST_X1 pe_1_0_6_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_0_6_N61), .SE(1'b0), .GCK(pe_1_0_6_net7069) );
  CLKGATETST_X1 pe_1_0_6_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_0_6_N60), .SE(1'b0), .GCK(pe_1_0_6_net7074) );
  CLKGATETST_X1 pe_1_0_6_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_0_6_N59), .SE(1'b0), .GCK(pe_1_0_6_net7079) );
  CLKGATETST_X1 pe_1_0_6_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_0_6_N90), .SE(1'b0), .GCK(pe_1_0_6_net7084) );
  CLKBUF_X1 pe_1_0_7_U112 ( .A(pe_1_0_7_n72), .Z(pe_1_0_7_n71) );
  INV_X1 pe_1_0_7_U111 ( .A(n73), .ZN(pe_1_0_7_n70) );
  INV_X1 pe_1_0_7_U110 ( .A(n65), .ZN(pe_1_0_7_n69) );
  INV_X1 pe_1_0_7_U109 ( .A(n65), .ZN(pe_1_0_7_n68) );
  INV_X1 pe_1_0_7_U108 ( .A(n65), .ZN(pe_1_0_7_n67) );
  INV_X1 pe_1_0_7_U107 ( .A(pe_1_0_7_n69), .ZN(pe_1_0_7_n66) );
  INV_X1 pe_1_0_7_U106 ( .A(pe_1_0_7_n63), .ZN(pe_1_0_7_n62) );
  INV_X1 pe_1_0_7_U105 ( .A(pe_1_0_7_n61), .ZN(pe_1_0_7_n60) );
  INV_X1 pe_1_0_7_U104 ( .A(n25), .ZN(pe_1_0_7_n59) );
  INV_X1 pe_1_0_7_U103 ( .A(pe_1_0_7_n59), .ZN(pe_1_0_7_n58) );
  INV_X1 pe_1_0_7_U102 ( .A(n17), .ZN(pe_1_0_7_n57) );
  MUX2_X1 pe_1_0_7_U101 ( .A(pe_1_0_7_n54), .B(pe_1_0_7_n51), .S(n44), .Z(
        int_data_x_0__7__3_) );
  MUX2_X1 pe_1_0_7_U100 ( .A(pe_1_0_7_n53), .B(pe_1_0_7_n52), .S(pe_1_0_7_n62), 
        .Z(pe_1_0_7_n54) );
  MUX2_X1 pe_1_0_7_U99 ( .A(pe_1_0_7_int_q_reg_h[23]), .B(
        pe_1_0_7_int_q_reg_h[19]), .S(pe_1_0_7_n56), .Z(pe_1_0_7_n53) );
  MUX2_X1 pe_1_0_7_U98 ( .A(pe_1_0_7_int_q_reg_h[15]), .B(
        pe_1_0_7_int_q_reg_h[11]), .S(pe_1_0_7_n56), .Z(pe_1_0_7_n52) );
  MUX2_X1 pe_1_0_7_U97 ( .A(pe_1_0_7_int_q_reg_h[7]), .B(
        pe_1_0_7_int_q_reg_h[3]), .S(pe_1_0_7_n56), .Z(pe_1_0_7_n51) );
  MUX2_X1 pe_1_0_7_U96 ( .A(pe_1_0_7_n50), .B(pe_1_0_7_n47), .S(n44), .Z(
        int_data_x_0__7__2_) );
  MUX2_X1 pe_1_0_7_U95 ( .A(pe_1_0_7_n49), .B(pe_1_0_7_n48), .S(pe_1_0_7_n62), 
        .Z(pe_1_0_7_n50) );
  MUX2_X1 pe_1_0_7_U94 ( .A(pe_1_0_7_int_q_reg_h[22]), .B(
        pe_1_0_7_int_q_reg_h[18]), .S(pe_1_0_7_n56), .Z(pe_1_0_7_n49) );
  MUX2_X1 pe_1_0_7_U93 ( .A(pe_1_0_7_int_q_reg_h[14]), .B(
        pe_1_0_7_int_q_reg_h[10]), .S(pe_1_0_7_n56), .Z(pe_1_0_7_n48) );
  MUX2_X1 pe_1_0_7_U92 ( .A(pe_1_0_7_int_q_reg_h[6]), .B(
        pe_1_0_7_int_q_reg_h[2]), .S(pe_1_0_7_n56), .Z(pe_1_0_7_n47) );
  MUX2_X1 pe_1_0_7_U91 ( .A(pe_1_0_7_n46), .B(pe_1_0_7_n24), .S(n44), .Z(
        int_data_x_0__7__1_) );
  MUX2_X1 pe_1_0_7_U90 ( .A(pe_1_0_7_n45), .B(pe_1_0_7_n25), .S(pe_1_0_7_n62), 
        .Z(pe_1_0_7_n46) );
  MUX2_X1 pe_1_0_7_U89 ( .A(pe_1_0_7_int_q_reg_h[21]), .B(
        pe_1_0_7_int_q_reg_h[17]), .S(pe_1_0_7_n56), .Z(pe_1_0_7_n45) );
  MUX2_X1 pe_1_0_7_U88 ( .A(pe_1_0_7_int_q_reg_h[13]), .B(
        pe_1_0_7_int_q_reg_h[9]), .S(pe_1_0_7_n56), .Z(pe_1_0_7_n25) );
  MUX2_X1 pe_1_0_7_U87 ( .A(pe_1_0_7_int_q_reg_h[5]), .B(
        pe_1_0_7_int_q_reg_h[1]), .S(pe_1_0_7_n56), .Z(pe_1_0_7_n24) );
  MUX2_X1 pe_1_0_7_U86 ( .A(pe_1_0_7_n23), .B(pe_1_0_7_n20), .S(n44), .Z(
        int_data_x_0__7__0_) );
  MUX2_X1 pe_1_0_7_U85 ( .A(pe_1_0_7_n22), .B(pe_1_0_7_n21), .S(pe_1_0_7_n62), 
        .Z(pe_1_0_7_n23) );
  MUX2_X1 pe_1_0_7_U84 ( .A(pe_1_0_7_int_q_reg_h[20]), .B(
        pe_1_0_7_int_q_reg_h[16]), .S(pe_1_0_7_n56), .Z(pe_1_0_7_n22) );
  MUX2_X1 pe_1_0_7_U83 ( .A(pe_1_0_7_int_q_reg_h[12]), .B(
        pe_1_0_7_int_q_reg_h[8]), .S(pe_1_0_7_n56), .Z(pe_1_0_7_n21) );
  MUX2_X1 pe_1_0_7_U82 ( .A(pe_1_0_7_int_q_reg_h[4]), .B(
        pe_1_0_7_int_q_reg_h[0]), .S(pe_1_0_7_n56), .Z(pe_1_0_7_n20) );
  MUX2_X1 pe_1_0_7_U81 ( .A(pe_1_0_7_n19), .B(pe_1_0_7_n16), .S(n44), .Z(
        pe_1_0_7_o_data_v_3_) );
  MUX2_X1 pe_1_0_7_U80 ( .A(pe_1_0_7_n18), .B(pe_1_0_7_n17), .S(pe_1_0_7_n62), 
        .Z(pe_1_0_7_n19) );
  MUX2_X1 pe_1_0_7_U79 ( .A(pe_1_0_7_int_q_reg_v[23]), .B(
        pe_1_0_7_int_q_reg_v[19]), .S(pe_1_0_7_n55), .Z(pe_1_0_7_n18) );
  MUX2_X1 pe_1_0_7_U78 ( .A(pe_1_0_7_int_q_reg_v[15]), .B(
        pe_1_0_7_int_q_reg_v[11]), .S(pe_1_0_7_n55), .Z(pe_1_0_7_n17) );
  MUX2_X1 pe_1_0_7_U77 ( .A(pe_1_0_7_int_q_reg_v[7]), .B(
        pe_1_0_7_int_q_reg_v[3]), .S(pe_1_0_7_n55), .Z(pe_1_0_7_n16) );
  MUX2_X1 pe_1_0_7_U76 ( .A(pe_1_0_7_n15), .B(pe_1_0_7_n12), .S(n44), .Z(
        pe_1_0_7_o_data_v_2_) );
  MUX2_X1 pe_1_0_7_U75 ( .A(pe_1_0_7_n14), .B(pe_1_0_7_n13), .S(pe_1_0_7_n62), 
        .Z(pe_1_0_7_n15) );
  MUX2_X1 pe_1_0_7_U74 ( .A(pe_1_0_7_int_q_reg_v[22]), .B(
        pe_1_0_7_int_q_reg_v[18]), .S(pe_1_0_7_n55), .Z(pe_1_0_7_n14) );
  MUX2_X1 pe_1_0_7_U73 ( .A(pe_1_0_7_int_q_reg_v[14]), .B(
        pe_1_0_7_int_q_reg_v[10]), .S(pe_1_0_7_n55), .Z(pe_1_0_7_n13) );
  MUX2_X1 pe_1_0_7_U72 ( .A(pe_1_0_7_int_q_reg_v[6]), .B(
        pe_1_0_7_int_q_reg_v[2]), .S(pe_1_0_7_n55), .Z(pe_1_0_7_n12) );
  MUX2_X1 pe_1_0_7_U71 ( .A(pe_1_0_7_n11), .B(pe_1_0_7_n8), .S(n44), .Z(
        pe_1_0_7_o_data_v_1_) );
  MUX2_X1 pe_1_0_7_U70 ( .A(pe_1_0_7_n10), .B(pe_1_0_7_n9), .S(pe_1_0_7_n62), 
        .Z(pe_1_0_7_n11) );
  MUX2_X1 pe_1_0_7_U69 ( .A(pe_1_0_7_int_q_reg_v[21]), .B(
        pe_1_0_7_int_q_reg_v[17]), .S(pe_1_0_7_n55), .Z(pe_1_0_7_n10) );
  MUX2_X1 pe_1_0_7_U68 ( .A(pe_1_0_7_int_q_reg_v[13]), .B(
        pe_1_0_7_int_q_reg_v[9]), .S(pe_1_0_7_n55), .Z(pe_1_0_7_n9) );
  MUX2_X1 pe_1_0_7_U67 ( .A(pe_1_0_7_int_q_reg_v[5]), .B(
        pe_1_0_7_int_q_reg_v[1]), .S(pe_1_0_7_n55), .Z(pe_1_0_7_n8) );
  MUX2_X1 pe_1_0_7_U66 ( .A(pe_1_0_7_n7), .B(pe_1_0_7_n4), .S(n44), .Z(
        pe_1_0_7_o_data_v_0_) );
  MUX2_X1 pe_1_0_7_U65 ( .A(pe_1_0_7_n6), .B(pe_1_0_7_n5), .S(pe_1_0_7_n62), 
        .Z(pe_1_0_7_n7) );
  MUX2_X1 pe_1_0_7_U64 ( .A(pe_1_0_7_int_q_reg_v[20]), .B(
        pe_1_0_7_int_q_reg_v[16]), .S(pe_1_0_7_n55), .Z(pe_1_0_7_n6) );
  MUX2_X1 pe_1_0_7_U63 ( .A(pe_1_0_7_int_q_reg_v[12]), .B(
        pe_1_0_7_int_q_reg_v[8]), .S(pe_1_0_7_n55), .Z(pe_1_0_7_n5) );
  MUX2_X1 pe_1_0_7_U62 ( .A(pe_1_0_7_int_q_reg_v[4]), .B(
        pe_1_0_7_int_q_reg_v[0]), .S(pe_1_0_7_n55), .Z(pe_1_0_7_n4) );
  XNOR2_X1 pe_1_0_7_U61 ( .A(pe_1_0_7_n73), .B(o_data[0]), .ZN(pe_1_0_7_N70)
         );
  AOI222_X1 pe_1_0_7_U60 ( .A1(int_data_res_1__7__0_), .A2(pe_1_0_7_n64), .B1(
        pe_1_0_7_n1), .B2(pe_1_0_7_n27), .C1(pe_1_0_7_N70), .C2(pe_1_0_7_n28), 
        .ZN(pe_1_0_7_n35) );
  INV_X1 pe_1_0_7_U59 ( .A(pe_1_0_7_n35), .ZN(pe_1_0_7_n84) );
  AOI222_X1 pe_1_0_7_U58 ( .A1(int_data_res_1__7__2_), .A2(pe_1_0_7_n64), .B1(
        pe_1_0_7_N80), .B2(pe_1_0_7_n27), .C1(pe_1_0_7_N72), .C2(pe_1_0_7_n28), 
        .ZN(pe_1_0_7_n33) );
  INV_X1 pe_1_0_7_U57 ( .A(pe_1_0_7_n33), .ZN(pe_1_0_7_n82) );
  AOI222_X1 pe_1_0_7_U52 ( .A1(int_data_res_1__7__6_), .A2(pe_1_0_7_n64), .B1(
        pe_1_0_7_N84), .B2(pe_1_0_7_n27), .C1(pe_1_0_7_N76), .C2(pe_1_0_7_n28), 
        .ZN(pe_1_0_7_n29) );
  INV_X1 pe_1_0_7_U51 ( .A(pe_1_0_7_n29), .ZN(pe_1_0_7_n78) );
  AOI222_X1 pe_1_0_7_U50 ( .A1(int_data_res_1__7__1_), .A2(pe_1_0_7_n64), .B1(
        pe_1_0_7_N79), .B2(pe_1_0_7_n27), .C1(pe_1_0_7_N71), .C2(pe_1_0_7_n28), 
        .ZN(pe_1_0_7_n34) );
  INV_X1 pe_1_0_7_U49 ( .A(pe_1_0_7_n34), .ZN(pe_1_0_7_n83) );
  AOI222_X1 pe_1_0_7_U48 ( .A1(int_data_res_1__7__3_), .A2(pe_1_0_7_n64), .B1(
        pe_1_0_7_N81), .B2(pe_1_0_7_n27), .C1(pe_1_0_7_N73), .C2(pe_1_0_7_n28), 
        .ZN(pe_1_0_7_n32) );
  INV_X1 pe_1_0_7_U47 ( .A(pe_1_0_7_n32), .ZN(pe_1_0_7_n81) );
  AOI222_X1 pe_1_0_7_U46 ( .A1(int_data_res_1__7__4_), .A2(pe_1_0_7_n64), .B1(
        pe_1_0_7_N82), .B2(pe_1_0_7_n27), .C1(pe_1_0_7_N74), .C2(pe_1_0_7_n28), 
        .ZN(pe_1_0_7_n31) );
  INV_X1 pe_1_0_7_U45 ( .A(pe_1_0_7_n31), .ZN(pe_1_0_7_n80) );
  AOI222_X1 pe_1_0_7_U44 ( .A1(int_data_res_1__7__5_), .A2(pe_1_0_7_n64), .B1(
        pe_1_0_7_N83), .B2(pe_1_0_7_n27), .C1(pe_1_0_7_N75), .C2(pe_1_0_7_n28), 
        .ZN(pe_1_0_7_n30) );
  INV_X1 pe_1_0_7_U43 ( .A(pe_1_0_7_n30), .ZN(pe_1_0_7_n79) );
  INV_X1 pe_1_0_7_U42 ( .A(pe_1_0_7_int_data_2_), .ZN(pe_1_0_7_n75) );
  NAND2_X1 pe_1_0_7_U41 ( .A1(pe_1_0_7_int_data_0_), .A2(pe_1_0_7_n3), .ZN(
        pe_1_0_7_sub_81_carry[1]) );
  INV_X1 pe_1_0_7_U40 ( .A(pe_1_0_7_int_data_1_), .ZN(pe_1_0_7_n74) );
  AND2_X1 pe_1_0_7_U39 ( .A1(pe_1_0_7_int_data_0_), .A2(o_data[0]), .ZN(
        pe_1_0_7_n2) );
  AOI222_X1 pe_1_0_7_U38 ( .A1(pe_1_0_7_n64), .A2(int_data_res_1__7__7_), .B1(
        pe_1_0_7_N85), .B2(pe_1_0_7_n27), .C1(pe_1_0_7_N77), .C2(pe_1_0_7_n28), 
        .ZN(pe_1_0_7_n26) );
  INV_X1 pe_1_0_7_U37 ( .A(pe_1_0_7_n26), .ZN(pe_1_0_7_n77) );
  NOR3_X1 pe_1_0_7_U36 ( .A1(pe_1_0_7_n59), .A2(pe_1_0_7_n65), .A3(int_ckg[56]), .ZN(pe_1_0_7_n36) );
  OR2_X1 pe_1_0_7_U35 ( .A1(pe_1_0_7_n36), .A2(pe_1_0_7_n64), .ZN(pe_1_0_7_N90) );
  INV_X1 pe_1_0_7_U34 ( .A(n37), .ZN(pe_1_0_7_n63) );
  AND2_X1 pe_1_0_7_U33 ( .A1(int_data_x_0__7__2_), .A2(pe_1_0_7_n58), .ZN(
        pe_1_0_7_int_data_2_) );
  AND2_X1 pe_1_0_7_U32 ( .A1(int_data_x_0__7__1_), .A2(pe_1_0_7_n58), .ZN(
        pe_1_0_7_int_data_1_) );
  AND2_X1 pe_1_0_7_U31 ( .A1(int_data_x_0__7__3_), .A2(pe_1_0_7_n58), .ZN(
        pe_1_0_7_int_data_3_) );
  BUF_X1 pe_1_0_7_U30 ( .A(n59), .Z(pe_1_0_7_n64) );
  INV_X1 pe_1_0_7_U29 ( .A(n31), .ZN(pe_1_0_7_n61) );
  AND2_X1 pe_1_0_7_U28 ( .A1(int_data_x_0__7__0_), .A2(pe_1_0_7_n58), .ZN(
        pe_1_0_7_int_data_0_) );
  NAND2_X1 pe_1_0_7_U27 ( .A1(pe_1_0_7_n44), .A2(pe_1_0_7_n61), .ZN(
        pe_1_0_7_n41) );
  AND3_X1 pe_1_0_7_U26 ( .A1(n73), .A2(pe_1_0_7_n63), .A3(n44), .ZN(
        pe_1_0_7_n44) );
  INV_X1 pe_1_0_7_U25 ( .A(pe_1_0_7_int_data_3_), .ZN(pe_1_0_7_n76) );
  NOR2_X1 pe_1_0_7_U24 ( .A1(pe_1_0_7_n70), .A2(n44), .ZN(pe_1_0_7_n43) );
  NOR2_X1 pe_1_0_7_U23 ( .A1(pe_1_0_7_n57), .A2(pe_1_0_7_n64), .ZN(
        pe_1_0_7_n28) );
  NOR2_X1 pe_1_0_7_U22 ( .A1(n17), .A2(pe_1_0_7_n64), .ZN(pe_1_0_7_n27) );
  INV_X1 pe_1_0_7_U21 ( .A(pe_1_0_7_int_data_0_), .ZN(pe_1_0_7_n73) );
  BUF_X1 pe_1_0_7_U20 ( .A(pe_1_0_7_n60), .Z(pe_1_0_7_n55) );
  INV_X1 pe_1_0_7_U19 ( .A(pe_1_0_7_n41), .ZN(pe_1_0_7_n90) );
  INV_X1 pe_1_0_7_U18 ( .A(pe_1_0_7_n37), .ZN(pe_1_0_7_n88) );
  INV_X1 pe_1_0_7_U17 ( .A(pe_1_0_7_n38), .ZN(pe_1_0_7_n87) );
  INV_X1 pe_1_0_7_U16 ( .A(pe_1_0_7_n39), .ZN(pe_1_0_7_n86) );
  NOR2_X1 pe_1_0_7_U15 ( .A1(pe_1_0_7_n68), .A2(pe_1_0_7_n42), .ZN(
        pe_1_0_7_N59) );
  NOR2_X1 pe_1_0_7_U14 ( .A1(pe_1_0_7_n68), .A2(pe_1_0_7_n41), .ZN(
        pe_1_0_7_N60) );
  NOR2_X1 pe_1_0_7_U13 ( .A1(pe_1_0_7_n68), .A2(pe_1_0_7_n38), .ZN(
        pe_1_0_7_N63) );
  NOR2_X1 pe_1_0_7_U12 ( .A1(pe_1_0_7_n67), .A2(pe_1_0_7_n40), .ZN(
        pe_1_0_7_N61) );
  NOR2_X1 pe_1_0_7_U11 ( .A1(pe_1_0_7_n67), .A2(pe_1_0_7_n39), .ZN(
        pe_1_0_7_N62) );
  NOR2_X1 pe_1_0_7_U10 ( .A1(pe_1_0_7_n37), .A2(pe_1_0_7_n67), .ZN(
        pe_1_0_7_N64) );
  NAND2_X1 pe_1_0_7_U9 ( .A1(pe_1_0_7_n44), .A2(pe_1_0_7_n60), .ZN(
        pe_1_0_7_n42) );
  INV_X1 pe_1_0_7_U8 ( .A(pe_1_0_7_n69), .ZN(pe_1_0_7_n65) );
  BUF_X1 pe_1_0_7_U7 ( .A(pe_1_0_7_n60), .Z(pe_1_0_7_n56) );
  INV_X1 pe_1_0_7_U6 ( .A(pe_1_0_7_n42), .ZN(pe_1_0_7_n89) );
  INV_X1 pe_1_0_7_U5 ( .A(pe_1_0_7_n40), .ZN(pe_1_0_7_n85) );
  INV_X2 pe_1_0_7_U4 ( .A(n81), .ZN(pe_1_0_7_n72) );
  XOR2_X1 pe_1_0_7_U3 ( .A(pe_1_0_7_int_data_0_), .B(o_data[0]), .Z(
        pe_1_0_7_n1) );
  DFFR_X1 pe_1_0_7_int_q_acc_reg_0_ ( .D(pe_1_0_7_n84), .CK(pe_1_0_7_net7006), 
        .RN(pe_1_0_7_n72), .Q(o_data[0]), .QN(pe_1_0_7_n3) );
  DFFR_X1 pe_1_0_7_int_q_reg_v_reg_0__0_ ( .D(int_data_y_1__7__0_), .CK(
        pe_1_0_7_net6976), .RN(pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_v[20]) );
  DFFR_X1 pe_1_0_7_int_q_reg_v_reg_0__1_ ( .D(int_data_y_1__7__1_), .CK(
        pe_1_0_7_net6976), .RN(pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_v[21]) );
  DFFR_X1 pe_1_0_7_int_q_reg_v_reg_0__2_ ( .D(int_data_y_1__7__2_), .CK(
        pe_1_0_7_net6976), .RN(pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_v[22]) );
  DFFR_X1 pe_1_0_7_int_q_reg_v_reg_0__3_ ( .D(int_data_y_1__7__3_), .CK(
        pe_1_0_7_net6976), .RN(pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_v[23]) );
  DFFR_X1 pe_1_0_7_int_q_reg_v_reg_1__0_ ( .D(int_data_y_1__7__0_), .CK(
        pe_1_0_7_net6981), .RN(pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_v[16]) );
  DFFR_X1 pe_1_0_7_int_q_reg_v_reg_1__1_ ( .D(int_data_y_1__7__1_), .CK(
        pe_1_0_7_net6981), .RN(pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_v[17]) );
  DFFR_X1 pe_1_0_7_int_q_reg_v_reg_1__2_ ( .D(int_data_y_1__7__2_), .CK(
        pe_1_0_7_net6981), .RN(pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_v[18]) );
  DFFR_X1 pe_1_0_7_int_q_reg_v_reg_1__3_ ( .D(int_data_y_1__7__3_), .CK(
        pe_1_0_7_net6981), .RN(pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_v[19]) );
  DFFR_X1 pe_1_0_7_int_q_reg_v_reg_2__0_ ( .D(int_data_y_1__7__0_), .CK(
        pe_1_0_7_net6986), .RN(pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_v[12]) );
  DFFR_X1 pe_1_0_7_int_q_reg_v_reg_2__1_ ( .D(int_data_y_1__7__1_), .CK(
        pe_1_0_7_net6986), .RN(pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_v[13]) );
  DFFR_X1 pe_1_0_7_int_q_reg_v_reg_2__2_ ( .D(int_data_y_1__7__2_), .CK(
        pe_1_0_7_net6986), .RN(pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_v[14]) );
  DFFR_X1 pe_1_0_7_int_q_reg_v_reg_2__3_ ( .D(int_data_y_1__7__3_), .CK(
        pe_1_0_7_net6986), .RN(pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_v[15]) );
  DFFR_X1 pe_1_0_7_int_q_reg_v_reg_3__0_ ( .D(int_data_y_1__7__0_), .CK(
        pe_1_0_7_net6991), .RN(pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_v[8]) );
  DFFR_X1 pe_1_0_7_int_q_reg_v_reg_3__1_ ( .D(int_data_y_1__7__1_), .CK(
        pe_1_0_7_net6991), .RN(pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_v[9]) );
  DFFR_X1 pe_1_0_7_int_q_reg_v_reg_3__2_ ( .D(int_data_y_1__7__2_), .CK(
        pe_1_0_7_net6991), .RN(pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_v[10]) );
  DFFR_X1 pe_1_0_7_int_q_reg_v_reg_3__3_ ( .D(int_data_y_1__7__3_), .CK(
        pe_1_0_7_net6991), .RN(pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_v[11]) );
  DFFR_X1 pe_1_0_7_int_q_reg_v_reg_4__0_ ( .D(int_data_y_1__7__0_), .CK(
        pe_1_0_7_net6996), .RN(pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_v[4]) );
  DFFR_X1 pe_1_0_7_int_q_reg_v_reg_4__1_ ( .D(int_data_y_1__7__1_), .CK(
        pe_1_0_7_net6996), .RN(pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_v[5]) );
  DFFR_X1 pe_1_0_7_int_q_reg_v_reg_4__2_ ( .D(int_data_y_1__7__2_), .CK(
        pe_1_0_7_net6996), .RN(pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_v[6]) );
  DFFR_X1 pe_1_0_7_int_q_reg_v_reg_4__3_ ( .D(int_data_y_1__7__3_), .CK(
        pe_1_0_7_net6996), .RN(pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_v[7]) );
  DFFR_X1 pe_1_0_7_int_q_reg_v_reg_5__0_ ( .D(int_data_y_1__7__0_), .CK(
        pe_1_0_7_net7001), .RN(pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_v[0]) );
  DFFR_X1 pe_1_0_7_int_q_reg_v_reg_5__1_ ( .D(int_data_y_1__7__1_), .CK(
        pe_1_0_7_net7001), .RN(pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_v[1]) );
  DFFR_X1 pe_1_0_7_int_q_reg_v_reg_5__2_ ( .D(int_data_y_1__7__2_), .CK(
        pe_1_0_7_net7001), .RN(pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_v[2]) );
  DFFR_X1 pe_1_0_7_int_q_reg_v_reg_5__3_ ( .D(int_data_y_1__7__3_), .CK(
        pe_1_0_7_net7001), .RN(pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_0_7_int_q_reg_h_reg_0__0_ ( .D(i_data_conv_h[28]), .SI(
        int_data_y_1__7__0_), .SE(pe_1_0_7_n65), .CK(pe_1_0_7_net6945), .RN(
        pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_0_7_int_q_reg_h_reg_0__1_ ( .D(i_data_conv_h[29]), .SI(
        int_data_y_1__7__1_), .SE(pe_1_0_7_n65), .CK(pe_1_0_7_net6945), .RN(
        pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_0_7_int_q_reg_h_reg_0__2_ ( .D(i_data_conv_h[30]), .SI(
        int_data_y_1__7__2_), .SE(pe_1_0_7_n65), .CK(pe_1_0_7_net6945), .RN(
        pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_0_7_int_q_reg_h_reg_0__3_ ( .D(i_data_conv_h[31]), .SI(
        int_data_y_1__7__3_), .SE(pe_1_0_7_n65), .CK(pe_1_0_7_net6945), .RN(
        pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_0_7_int_q_reg_h_reg_1__0_ ( .D(i_data_conv_h[28]), .SI(
        int_data_y_1__7__0_), .SE(pe_1_0_7_n65), .CK(pe_1_0_7_net6951), .RN(
        pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_0_7_int_q_reg_h_reg_1__1_ ( .D(i_data_conv_h[29]), .SI(
        int_data_y_1__7__1_), .SE(pe_1_0_7_n65), .CK(pe_1_0_7_net6951), .RN(
        pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_0_7_int_q_reg_h_reg_1__2_ ( .D(i_data_conv_h[30]), .SI(
        int_data_y_1__7__2_), .SE(pe_1_0_7_n65), .CK(pe_1_0_7_net6951), .RN(
        pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_0_7_int_q_reg_h_reg_1__3_ ( .D(i_data_conv_h[31]), .SI(
        int_data_y_1__7__3_), .SE(pe_1_0_7_n65), .CK(pe_1_0_7_net6951), .RN(
        pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_0_7_int_q_reg_h_reg_2__0_ ( .D(i_data_conv_h[28]), .SI(
        int_data_y_1__7__0_), .SE(pe_1_0_7_n65), .CK(pe_1_0_7_net6956), .RN(
        pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_0_7_int_q_reg_h_reg_2__1_ ( .D(i_data_conv_h[29]), .SI(
        int_data_y_1__7__1_), .SE(pe_1_0_7_n65), .CK(pe_1_0_7_net6956), .RN(
        pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_0_7_int_q_reg_h_reg_2__2_ ( .D(i_data_conv_h[30]), .SI(
        int_data_y_1__7__2_), .SE(pe_1_0_7_n65), .CK(pe_1_0_7_net6956), .RN(
        pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_0_7_int_q_reg_h_reg_2__3_ ( .D(i_data_conv_h[31]), .SI(
        int_data_y_1__7__3_), .SE(pe_1_0_7_n65), .CK(pe_1_0_7_net6956), .RN(
        pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_0_7_int_q_reg_h_reg_3__0_ ( .D(i_data_conv_h[28]), .SI(
        int_data_y_1__7__0_), .SE(pe_1_0_7_n65), .CK(pe_1_0_7_net6961), .RN(
        pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_0_7_int_q_reg_h_reg_3__1_ ( .D(i_data_conv_h[29]), .SI(
        int_data_y_1__7__1_), .SE(pe_1_0_7_n65), .CK(pe_1_0_7_net6961), .RN(
        pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_0_7_int_q_reg_h_reg_3__2_ ( .D(i_data_conv_h[30]), .SI(
        int_data_y_1__7__2_), .SE(pe_1_0_7_n65), .CK(pe_1_0_7_net6961), .RN(
        pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_0_7_int_q_reg_h_reg_3__3_ ( .D(i_data_conv_h[31]), .SI(
        int_data_y_1__7__3_), .SE(pe_1_0_7_n65), .CK(pe_1_0_7_net6961), .RN(
        pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_0_7_int_q_reg_h_reg_4__0_ ( .D(i_data_conv_h[28]), .SI(
        int_data_y_1__7__0_), .SE(pe_1_0_7_n66), .CK(pe_1_0_7_net6966), .RN(
        pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_0_7_int_q_reg_h_reg_4__1_ ( .D(i_data_conv_h[29]), .SI(
        int_data_y_1__7__1_), .SE(pe_1_0_7_n66), .CK(pe_1_0_7_net6966), .RN(
        pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_0_7_int_q_reg_h_reg_4__2_ ( .D(i_data_conv_h[30]), .SI(
        int_data_y_1__7__2_), .SE(pe_1_0_7_n66), .CK(pe_1_0_7_net6966), .RN(
        pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_0_7_int_q_reg_h_reg_4__3_ ( .D(i_data_conv_h[31]), .SI(
        int_data_y_1__7__3_), .SE(pe_1_0_7_n66), .CK(pe_1_0_7_net6966), .RN(
        pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_0_7_int_q_reg_h_reg_5__0_ ( .D(i_data_conv_h[28]), .SI(
        int_data_y_1__7__0_), .SE(pe_1_0_7_n66), .CK(pe_1_0_7_net6971), .RN(
        pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_0_7_int_q_reg_h_reg_5__1_ ( .D(i_data_conv_h[29]), .SI(
        int_data_y_1__7__1_), .SE(pe_1_0_7_n66), .CK(pe_1_0_7_net6971), .RN(
        pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_0_7_int_q_reg_h_reg_5__2_ ( .D(i_data_conv_h[30]), .SI(
        int_data_y_1__7__2_), .SE(pe_1_0_7_n66), .CK(pe_1_0_7_net6971), .RN(
        pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_0_7_int_q_reg_h_reg_5__3_ ( .D(i_data_conv_h[31]), .SI(
        int_data_y_1__7__3_), .SE(pe_1_0_7_n66), .CK(pe_1_0_7_net6971), .RN(
        pe_1_0_7_n72), .Q(pe_1_0_7_int_q_reg_h[3]) );
  FA_X1 pe_1_0_7_sub_81_U2_7 ( .A(o_data[7]), .B(pe_1_0_7_n76), .CI(
        pe_1_0_7_sub_81_carry[7]), .S(pe_1_0_7_N77) );
  FA_X1 pe_1_0_7_sub_81_U2_6 ( .A(o_data[6]), .B(pe_1_0_7_n76), .CI(
        pe_1_0_7_sub_81_carry[6]), .CO(pe_1_0_7_sub_81_carry[7]), .S(
        pe_1_0_7_N76) );
  FA_X1 pe_1_0_7_sub_81_U2_5 ( .A(o_data[5]), .B(pe_1_0_7_n76), .CI(
        pe_1_0_7_sub_81_carry[5]), .CO(pe_1_0_7_sub_81_carry[6]), .S(
        pe_1_0_7_N75) );
  FA_X1 pe_1_0_7_sub_81_U2_4 ( .A(o_data[4]), .B(pe_1_0_7_n76), .CI(
        pe_1_0_7_sub_81_carry[4]), .CO(pe_1_0_7_sub_81_carry[5]), .S(
        pe_1_0_7_N74) );
  FA_X1 pe_1_0_7_sub_81_U2_3 ( .A(o_data[3]), .B(pe_1_0_7_n76), .CI(
        pe_1_0_7_sub_81_carry[3]), .CO(pe_1_0_7_sub_81_carry[4]), .S(
        pe_1_0_7_N73) );
  FA_X1 pe_1_0_7_sub_81_U2_2 ( .A(o_data[2]), .B(pe_1_0_7_n75), .CI(
        pe_1_0_7_sub_81_carry[2]), .CO(pe_1_0_7_sub_81_carry[3]), .S(
        pe_1_0_7_N72) );
  FA_X1 pe_1_0_7_sub_81_U2_1 ( .A(o_data[1]), .B(pe_1_0_7_n74), .CI(
        pe_1_0_7_sub_81_carry[1]), .CO(pe_1_0_7_sub_81_carry[2]), .S(
        pe_1_0_7_N71) );
  FA_X1 pe_1_0_7_add_83_U1_7 ( .A(o_data[7]), .B(pe_1_0_7_int_data_3_), .CI(
        pe_1_0_7_add_83_carry[7]), .S(pe_1_0_7_N85) );
  FA_X1 pe_1_0_7_add_83_U1_6 ( .A(o_data[6]), .B(pe_1_0_7_int_data_3_), .CI(
        pe_1_0_7_add_83_carry[6]), .CO(pe_1_0_7_add_83_carry[7]), .S(
        pe_1_0_7_N84) );
  FA_X1 pe_1_0_7_add_83_U1_5 ( .A(o_data[5]), .B(pe_1_0_7_int_data_3_), .CI(
        pe_1_0_7_add_83_carry[5]), .CO(pe_1_0_7_add_83_carry[6]), .S(
        pe_1_0_7_N83) );
  FA_X1 pe_1_0_7_add_83_U1_4 ( .A(o_data[4]), .B(pe_1_0_7_int_data_3_), .CI(
        pe_1_0_7_add_83_carry[4]), .CO(pe_1_0_7_add_83_carry[5]), .S(
        pe_1_0_7_N82) );
  FA_X1 pe_1_0_7_add_83_U1_3 ( .A(o_data[3]), .B(pe_1_0_7_int_data_3_), .CI(
        pe_1_0_7_add_83_carry[3]), .CO(pe_1_0_7_add_83_carry[4]), .S(
        pe_1_0_7_N81) );
  FA_X1 pe_1_0_7_add_83_U1_2 ( .A(o_data[2]), .B(pe_1_0_7_int_data_2_), .CI(
        pe_1_0_7_add_83_carry[2]), .CO(pe_1_0_7_add_83_carry[3]), .S(
        pe_1_0_7_N80) );
  FA_X1 pe_1_0_7_add_83_U1_1 ( .A(o_data[1]), .B(pe_1_0_7_int_data_1_), .CI(
        pe_1_0_7_n2), .CO(pe_1_0_7_add_83_carry[2]), .S(pe_1_0_7_N79) );
  NAND3_X1 pe_1_0_7_U56 ( .A1(pe_1_0_7_n60), .A2(pe_1_0_7_n43), .A3(
        pe_1_0_7_n62), .ZN(pe_1_0_7_n40) );
  NAND3_X1 pe_1_0_7_U55 ( .A1(pe_1_0_7_n43), .A2(pe_1_0_7_n61), .A3(
        pe_1_0_7_n62), .ZN(pe_1_0_7_n39) );
  NAND3_X1 pe_1_0_7_U54 ( .A1(pe_1_0_7_n43), .A2(pe_1_0_7_n63), .A3(
        pe_1_0_7_n60), .ZN(pe_1_0_7_n38) );
  NAND3_X1 pe_1_0_7_U53 ( .A1(pe_1_0_7_n61), .A2(pe_1_0_7_n63), .A3(
        pe_1_0_7_n43), .ZN(pe_1_0_7_n37) );
  DFFR_X1 pe_1_0_7_int_q_acc_reg_6_ ( .D(pe_1_0_7_n78), .CK(pe_1_0_7_net7006), 
        .RN(pe_1_0_7_n71), .Q(o_data[6]) );
  DFFR_X1 pe_1_0_7_int_q_acc_reg_5_ ( .D(pe_1_0_7_n79), .CK(pe_1_0_7_net7006), 
        .RN(pe_1_0_7_n71), .Q(o_data[5]) );
  DFFR_X1 pe_1_0_7_int_q_acc_reg_4_ ( .D(pe_1_0_7_n80), .CK(pe_1_0_7_net7006), 
        .RN(pe_1_0_7_n71), .Q(o_data[4]) );
  DFFR_X1 pe_1_0_7_int_q_acc_reg_3_ ( .D(pe_1_0_7_n81), .CK(pe_1_0_7_net7006), 
        .RN(pe_1_0_7_n71), .Q(o_data[3]) );
  DFFR_X1 pe_1_0_7_int_q_acc_reg_2_ ( .D(pe_1_0_7_n82), .CK(pe_1_0_7_net7006), 
        .RN(pe_1_0_7_n71), .Q(o_data[2]) );
  DFFR_X1 pe_1_0_7_int_q_acc_reg_1_ ( .D(pe_1_0_7_n83), .CK(pe_1_0_7_net7006), 
        .RN(pe_1_0_7_n71), .Q(o_data[1]) );
  DFFR_X1 pe_1_0_7_int_q_acc_reg_7_ ( .D(pe_1_0_7_n77), .CK(pe_1_0_7_net7006), 
        .RN(pe_1_0_7_n71), .Q(o_data[7]) );
  CLKGATETST_X1 pe_1_0_7_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_0_7_n88), .SE(1'b0), .GCK(pe_1_0_7_net6945) );
  CLKGATETST_X1 pe_1_0_7_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_0_7_n87), .SE(1'b0), .GCK(pe_1_0_7_net6951) );
  CLKGATETST_X1 pe_1_0_7_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_0_7_n86), .SE(1'b0), .GCK(pe_1_0_7_net6956) );
  CLKGATETST_X1 pe_1_0_7_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_0_7_n85), .SE(1'b0), .GCK(pe_1_0_7_net6961) );
  CLKGATETST_X1 pe_1_0_7_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_0_7_n90), .SE(1'b0), .GCK(pe_1_0_7_net6966) );
  CLKGATETST_X1 pe_1_0_7_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_0_7_n89), .SE(1'b0), .GCK(pe_1_0_7_net6971) );
  CLKGATETST_X1 pe_1_0_7_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_0_7_N64), .SE(1'b0), .GCK(pe_1_0_7_net6976) );
  CLKGATETST_X1 pe_1_0_7_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_0_7_N63), .SE(1'b0), .GCK(pe_1_0_7_net6981) );
  CLKGATETST_X1 pe_1_0_7_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_0_7_N62), .SE(1'b0), .GCK(pe_1_0_7_net6986) );
  CLKGATETST_X1 pe_1_0_7_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_0_7_N61), .SE(1'b0), .GCK(pe_1_0_7_net6991) );
  CLKGATETST_X1 pe_1_0_7_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_0_7_N60), .SE(1'b0), .GCK(pe_1_0_7_net6996) );
  CLKGATETST_X1 pe_1_0_7_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_0_7_N59), .SE(1'b0), .GCK(pe_1_0_7_net7001) );
  CLKGATETST_X1 pe_1_0_7_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_0_7_N90), .SE(1'b0), .GCK(pe_1_0_7_net7006) );
  CLKBUF_X1 pe_1_1_0_U112 ( .A(pe_1_1_0_n72), .Z(pe_1_1_0_n71) );
  INV_X1 pe_1_1_0_U111 ( .A(n73), .ZN(pe_1_1_0_n70) );
  INV_X1 pe_1_1_0_U110 ( .A(n65), .ZN(pe_1_1_0_n69) );
  INV_X1 pe_1_1_0_U109 ( .A(n65), .ZN(pe_1_1_0_n68) );
  INV_X1 pe_1_1_0_U108 ( .A(n65), .ZN(pe_1_1_0_n67) );
  INV_X1 pe_1_1_0_U107 ( .A(pe_1_1_0_n69), .ZN(pe_1_1_0_n66) );
  INV_X1 pe_1_1_0_U106 ( .A(pe_1_1_0_n63), .ZN(pe_1_1_0_n62) );
  INV_X1 pe_1_1_0_U105 ( .A(pe_1_1_0_n61), .ZN(pe_1_1_0_n60) );
  INV_X1 pe_1_1_0_U104 ( .A(n25), .ZN(pe_1_1_0_n59) );
  INV_X1 pe_1_1_0_U103 ( .A(pe_1_1_0_n59), .ZN(pe_1_1_0_n58) );
  INV_X1 pe_1_1_0_U102 ( .A(n17), .ZN(pe_1_1_0_n57) );
  MUX2_X1 pe_1_1_0_U101 ( .A(pe_1_1_0_n54), .B(pe_1_1_0_n51), .S(n44), .Z(
        pe_1_1_0_o_data_h_3_) );
  MUX2_X1 pe_1_1_0_U100 ( .A(pe_1_1_0_n53), .B(pe_1_1_0_n52), .S(pe_1_1_0_n62), 
        .Z(pe_1_1_0_n54) );
  MUX2_X1 pe_1_1_0_U99 ( .A(pe_1_1_0_int_q_reg_h[23]), .B(
        pe_1_1_0_int_q_reg_h[19]), .S(pe_1_1_0_n56), .Z(pe_1_1_0_n53) );
  MUX2_X1 pe_1_1_0_U98 ( .A(pe_1_1_0_int_q_reg_h[15]), .B(
        pe_1_1_0_int_q_reg_h[11]), .S(pe_1_1_0_n56), .Z(pe_1_1_0_n52) );
  MUX2_X1 pe_1_1_0_U97 ( .A(pe_1_1_0_int_q_reg_h[7]), .B(
        pe_1_1_0_int_q_reg_h[3]), .S(pe_1_1_0_n56), .Z(pe_1_1_0_n51) );
  MUX2_X1 pe_1_1_0_U96 ( .A(pe_1_1_0_n50), .B(pe_1_1_0_n47), .S(n44), .Z(
        pe_1_1_0_o_data_h_2_) );
  MUX2_X1 pe_1_1_0_U95 ( .A(pe_1_1_0_n49), .B(pe_1_1_0_n48), .S(pe_1_1_0_n62), 
        .Z(pe_1_1_0_n50) );
  MUX2_X1 pe_1_1_0_U94 ( .A(pe_1_1_0_int_q_reg_h[22]), .B(
        pe_1_1_0_int_q_reg_h[18]), .S(pe_1_1_0_n56), .Z(pe_1_1_0_n49) );
  MUX2_X1 pe_1_1_0_U93 ( .A(pe_1_1_0_int_q_reg_h[14]), .B(
        pe_1_1_0_int_q_reg_h[10]), .S(pe_1_1_0_n56), .Z(pe_1_1_0_n48) );
  MUX2_X1 pe_1_1_0_U92 ( .A(pe_1_1_0_int_q_reg_h[6]), .B(
        pe_1_1_0_int_q_reg_h[2]), .S(pe_1_1_0_n56), .Z(pe_1_1_0_n47) );
  MUX2_X1 pe_1_1_0_U91 ( .A(pe_1_1_0_n46), .B(pe_1_1_0_n24), .S(n44), .Z(
        pe_1_1_0_o_data_h_1_) );
  MUX2_X1 pe_1_1_0_U90 ( .A(pe_1_1_0_n45), .B(pe_1_1_0_n25), .S(pe_1_1_0_n62), 
        .Z(pe_1_1_0_n46) );
  MUX2_X1 pe_1_1_0_U89 ( .A(pe_1_1_0_int_q_reg_h[21]), .B(
        pe_1_1_0_int_q_reg_h[17]), .S(pe_1_1_0_n56), .Z(pe_1_1_0_n45) );
  MUX2_X1 pe_1_1_0_U88 ( .A(pe_1_1_0_int_q_reg_h[13]), .B(
        pe_1_1_0_int_q_reg_h[9]), .S(pe_1_1_0_n56), .Z(pe_1_1_0_n25) );
  MUX2_X1 pe_1_1_0_U87 ( .A(pe_1_1_0_int_q_reg_h[5]), .B(
        pe_1_1_0_int_q_reg_h[1]), .S(pe_1_1_0_n56), .Z(pe_1_1_0_n24) );
  MUX2_X1 pe_1_1_0_U86 ( .A(pe_1_1_0_n23), .B(pe_1_1_0_n20), .S(n44), .Z(
        pe_1_1_0_o_data_h_0_) );
  MUX2_X1 pe_1_1_0_U85 ( .A(pe_1_1_0_n22), .B(pe_1_1_0_n21), .S(pe_1_1_0_n62), 
        .Z(pe_1_1_0_n23) );
  MUX2_X1 pe_1_1_0_U84 ( .A(pe_1_1_0_int_q_reg_h[20]), .B(
        pe_1_1_0_int_q_reg_h[16]), .S(pe_1_1_0_n56), .Z(pe_1_1_0_n22) );
  MUX2_X1 pe_1_1_0_U83 ( .A(pe_1_1_0_int_q_reg_h[12]), .B(
        pe_1_1_0_int_q_reg_h[8]), .S(pe_1_1_0_n56), .Z(pe_1_1_0_n21) );
  MUX2_X1 pe_1_1_0_U82 ( .A(pe_1_1_0_int_q_reg_h[4]), .B(
        pe_1_1_0_int_q_reg_h[0]), .S(pe_1_1_0_n56), .Z(pe_1_1_0_n20) );
  MUX2_X1 pe_1_1_0_U81 ( .A(pe_1_1_0_n19), .B(pe_1_1_0_n16), .S(n44), .Z(
        int_data_y_1__0__3_) );
  MUX2_X1 pe_1_1_0_U80 ( .A(pe_1_1_0_n18), .B(pe_1_1_0_n17), .S(pe_1_1_0_n62), 
        .Z(pe_1_1_0_n19) );
  MUX2_X1 pe_1_1_0_U79 ( .A(pe_1_1_0_int_q_reg_v[23]), .B(
        pe_1_1_0_int_q_reg_v[19]), .S(pe_1_1_0_n55), .Z(pe_1_1_0_n18) );
  MUX2_X1 pe_1_1_0_U78 ( .A(pe_1_1_0_int_q_reg_v[15]), .B(
        pe_1_1_0_int_q_reg_v[11]), .S(pe_1_1_0_n55), .Z(pe_1_1_0_n17) );
  MUX2_X1 pe_1_1_0_U77 ( .A(pe_1_1_0_int_q_reg_v[7]), .B(
        pe_1_1_0_int_q_reg_v[3]), .S(pe_1_1_0_n55), .Z(pe_1_1_0_n16) );
  MUX2_X1 pe_1_1_0_U76 ( .A(pe_1_1_0_n15), .B(pe_1_1_0_n12), .S(n44), .Z(
        int_data_y_1__0__2_) );
  MUX2_X1 pe_1_1_0_U75 ( .A(pe_1_1_0_n14), .B(pe_1_1_0_n13), .S(pe_1_1_0_n62), 
        .Z(pe_1_1_0_n15) );
  MUX2_X1 pe_1_1_0_U74 ( .A(pe_1_1_0_int_q_reg_v[22]), .B(
        pe_1_1_0_int_q_reg_v[18]), .S(pe_1_1_0_n55), .Z(pe_1_1_0_n14) );
  MUX2_X1 pe_1_1_0_U73 ( .A(pe_1_1_0_int_q_reg_v[14]), .B(
        pe_1_1_0_int_q_reg_v[10]), .S(pe_1_1_0_n55), .Z(pe_1_1_0_n13) );
  MUX2_X1 pe_1_1_0_U72 ( .A(pe_1_1_0_int_q_reg_v[6]), .B(
        pe_1_1_0_int_q_reg_v[2]), .S(pe_1_1_0_n55), .Z(pe_1_1_0_n12) );
  MUX2_X1 pe_1_1_0_U71 ( .A(pe_1_1_0_n11), .B(pe_1_1_0_n8), .S(n44), .Z(
        int_data_y_1__0__1_) );
  MUX2_X1 pe_1_1_0_U70 ( .A(pe_1_1_0_n10), .B(pe_1_1_0_n9), .S(pe_1_1_0_n62), 
        .Z(pe_1_1_0_n11) );
  MUX2_X1 pe_1_1_0_U69 ( .A(pe_1_1_0_int_q_reg_v[21]), .B(
        pe_1_1_0_int_q_reg_v[17]), .S(pe_1_1_0_n55), .Z(pe_1_1_0_n10) );
  MUX2_X1 pe_1_1_0_U68 ( .A(pe_1_1_0_int_q_reg_v[13]), .B(
        pe_1_1_0_int_q_reg_v[9]), .S(pe_1_1_0_n55), .Z(pe_1_1_0_n9) );
  MUX2_X1 pe_1_1_0_U67 ( .A(pe_1_1_0_int_q_reg_v[5]), .B(
        pe_1_1_0_int_q_reg_v[1]), .S(pe_1_1_0_n55), .Z(pe_1_1_0_n8) );
  MUX2_X1 pe_1_1_0_U66 ( .A(pe_1_1_0_n7), .B(pe_1_1_0_n4), .S(n44), .Z(
        int_data_y_1__0__0_) );
  MUX2_X1 pe_1_1_0_U65 ( .A(pe_1_1_0_n6), .B(pe_1_1_0_n5), .S(pe_1_1_0_n62), 
        .Z(pe_1_1_0_n7) );
  MUX2_X1 pe_1_1_0_U64 ( .A(pe_1_1_0_int_q_reg_v[20]), .B(
        pe_1_1_0_int_q_reg_v[16]), .S(pe_1_1_0_n55), .Z(pe_1_1_0_n6) );
  MUX2_X1 pe_1_1_0_U63 ( .A(pe_1_1_0_int_q_reg_v[12]), .B(
        pe_1_1_0_int_q_reg_v[8]), .S(pe_1_1_0_n55), .Z(pe_1_1_0_n5) );
  MUX2_X1 pe_1_1_0_U62 ( .A(pe_1_1_0_int_q_reg_v[4]), .B(
        pe_1_1_0_int_q_reg_v[0]), .S(pe_1_1_0_n55), .Z(pe_1_1_0_n4) );
  AND2_X1 pe_1_1_0_U61 ( .A1(pe_1_1_0_o_data_h_3_), .A2(pe_1_1_0_n58), .ZN(
        pe_1_1_0_int_data_3_) );
  NAND2_X1 pe_1_1_0_U60 ( .A1(pe_1_1_0_int_data_0_), .A2(pe_1_1_0_n3), .ZN(
        pe_1_1_0_sub_81_carry[1]) );
  INV_X1 pe_1_1_0_U59 ( .A(pe_1_1_0_int_data_1_), .ZN(pe_1_1_0_n74) );
  AOI222_X1 pe_1_1_0_U58 ( .A1(pe_1_1_0_n64), .A2(int_data_res_2__0__7_), .B1(
        pe_1_1_0_N85), .B2(pe_1_1_0_n27), .C1(pe_1_1_0_N77), .C2(pe_1_1_0_n28), 
        .ZN(pe_1_1_0_n26) );
  INV_X1 pe_1_1_0_U57 ( .A(pe_1_1_0_n26), .ZN(pe_1_1_0_n77) );
  AOI222_X1 pe_1_1_0_U52 ( .A1(int_data_res_2__0__1_), .A2(pe_1_1_0_n64), .B1(
        pe_1_1_0_N79), .B2(pe_1_1_0_n27), .C1(pe_1_1_0_N71), .C2(pe_1_1_0_n28), 
        .ZN(pe_1_1_0_n34) );
  INV_X1 pe_1_1_0_U51 ( .A(pe_1_1_0_n34), .ZN(pe_1_1_0_n83) );
  AOI222_X1 pe_1_1_0_U50 ( .A1(int_data_res_2__0__2_), .A2(pe_1_1_0_n64), .B1(
        pe_1_1_0_N80), .B2(pe_1_1_0_n27), .C1(pe_1_1_0_N72), .C2(pe_1_1_0_n28), 
        .ZN(pe_1_1_0_n33) );
  INV_X1 pe_1_1_0_U49 ( .A(pe_1_1_0_n33), .ZN(pe_1_1_0_n82) );
  AOI222_X1 pe_1_1_0_U48 ( .A1(int_data_res_2__0__6_), .A2(pe_1_1_0_n64), .B1(
        pe_1_1_0_N84), .B2(pe_1_1_0_n27), .C1(pe_1_1_0_N76), .C2(pe_1_1_0_n28), 
        .ZN(pe_1_1_0_n29) );
  INV_X1 pe_1_1_0_U47 ( .A(pe_1_1_0_n29), .ZN(pe_1_1_0_n78) );
  AND2_X1 pe_1_1_0_U46 ( .A1(pe_1_1_0_o_data_h_2_), .A2(pe_1_1_0_n58), .ZN(
        pe_1_1_0_int_data_2_) );
  AND2_X1 pe_1_1_0_U45 ( .A1(pe_1_1_0_o_data_h_1_), .A2(pe_1_1_0_n58), .ZN(
        pe_1_1_0_int_data_1_) );
  INV_X1 pe_1_1_0_U44 ( .A(pe_1_1_0_int_data_2_), .ZN(pe_1_1_0_n75) );
  AND2_X1 pe_1_1_0_U43 ( .A1(pe_1_1_0_int_data_0_), .A2(int_data_res_1__0__0_), 
        .ZN(pe_1_1_0_n2) );
  AND2_X1 pe_1_1_0_U42 ( .A1(pe_1_1_0_o_data_h_0_), .A2(pe_1_1_0_n58), .ZN(
        pe_1_1_0_int_data_0_) );
  XNOR2_X1 pe_1_1_0_U41 ( .A(pe_1_1_0_n73), .B(int_data_res_1__0__0_), .ZN(
        pe_1_1_0_N70) );
  AOI222_X1 pe_1_1_0_U40 ( .A1(int_data_res_2__0__0_), .A2(pe_1_1_0_n64), .B1(
        pe_1_1_0_n1), .B2(pe_1_1_0_n27), .C1(pe_1_1_0_N70), .C2(pe_1_1_0_n28), 
        .ZN(pe_1_1_0_n35) );
  INV_X1 pe_1_1_0_U39 ( .A(pe_1_1_0_n35), .ZN(pe_1_1_0_n84) );
  AOI222_X1 pe_1_1_0_U38 ( .A1(int_data_res_2__0__3_), .A2(pe_1_1_0_n64), .B1(
        pe_1_1_0_N81), .B2(pe_1_1_0_n27), .C1(pe_1_1_0_N73), .C2(pe_1_1_0_n28), 
        .ZN(pe_1_1_0_n32) );
  INV_X1 pe_1_1_0_U37 ( .A(pe_1_1_0_n32), .ZN(pe_1_1_0_n81) );
  AOI222_X1 pe_1_1_0_U36 ( .A1(int_data_res_2__0__4_), .A2(pe_1_1_0_n64), .B1(
        pe_1_1_0_N82), .B2(pe_1_1_0_n27), .C1(pe_1_1_0_N74), .C2(pe_1_1_0_n28), 
        .ZN(pe_1_1_0_n31) );
  INV_X1 pe_1_1_0_U35 ( .A(pe_1_1_0_n31), .ZN(pe_1_1_0_n80) );
  AOI222_X1 pe_1_1_0_U34 ( .A1(int_data_res_2__0__5_), .A2(pe_1_1_0_n64), .B1(
        pe_1_1_0_N83), .B2(pe_1_1_0_n27), .C1(pe_1_1_0_N75), .C2(pe_1_1_0_n28), 
        .ZN(pe_1_1_0_n30) );
  INV_X1 pe_1_1_0_U33 ( .A(pe_1_1_0_n30), .ZN(pe_1_1_0_n79) );
  NOR3_X1 pe_1_1_0_U32 ( .A1(pe_1_1_0_n59), .A2(pe_1_1_0_n65), .A3(int_ckg[55]), .ZN(pe_1_1_0_n36) );
  OR2_X1 pe_1_1_0_U31 ( .A1(pe_1_1_0_n36), .A2(pe_1_1_0_n64), .ZN(pe_1_1_0_N90) );
  INV_X1 pe_1_1_0_U30 ( .A(pe_1_1_0_int_data_0_), .ZN(pe_1_1_0_n73) );
  INV_X1 pe_1_1_0_U29 ( .A(n37), .ZN(pe_1_1_0_n63) );
  INV_X1 pe_1_1_0_U28 ( .A(n31), .ZN(pe_1_1_0_n61) );
  INV_X1 pe_1_1_0_U27 ( .A(pe_1_1_0_int_data_3_), .ZN(pe_1_1_0_n76) );
  BUF_X1 pe_1_1_0_U26 ( .A(n59), .Z(pe_1_1_0_n64) );
  NAND2_X1 pe_1_1_0_U25 ( .A1(pe_1_1_0_n44), .A2(pe_1_1_0_n61), .ZN(
        pe_1_1_0_n41) );
  AND3_X1 pe_1_1_0_U24 ( .A1(n73), .A2(pe_1_1_0_n63), .A3(n44), .ZN(
        pe_1_1_0_n44) );
  NOR2_X1 pe_1_1_0_U23 ( .A1(pe_1_1_0_n70), .A2(n44), .ZN(pe_1_1_0_n43) );
  NOR2_X1 pe_1_1_0_U22 ( .A1(pe_1_1_0_n57), .A2(pe_1_1_0_n64), .ZN(
        pe_1_1_0_n28) );
  NOR2_X1 pe_1_1_0_U21 ( .A1(n17), .A2(pe_1_1_0_n64), .ZN(pe_1_1_0_n27) );
  INV_X1 pe_1_1_0_U20 ( .A(pe_1_1_0_n41), .ZN(pe_1_1_0_n90) );
  INV_X1 pe_1_1_0_U19 ( .A(pe_1_1_0_n37), .ZN(pe_1_1_0_n88) );
  INV_X1 pe_1_1_0_U18 ( .A(pe_1_1_0_n38), .ZN(pe_1_1_0_n87) );
  INV_X1 pe_1_1_0_U17 ( .A(pe_1_1_0_n39), .ZN(pe_1_1_0_n86) );
  NOR2_X1 pe_1_1_0_U16 ( .A1(pe_1_1_0_n68), .A2(pe_1_1_0_n42), .ZN(
        pe_1_1_0_N59) );
  NOR2_X1 pe_1_1_0_U15 ( .A1(pe_1_1_0_n68), .A2(pe_1_1_0_n41), .ZN(
        pe_1_1_0_N60) );
  NOR2_X1 pe_1_1_0_U14 ( .A1(pe_1_1_0_n68), .A2(pe_1_1_0_n38), .ZN(
        pe_1_1_0_N63) );
  NOR2_X1 pe_1_1_0_U13 ( .A1(pe_1_1_0_n67), .A2(pe_1_1_0_n40), .ZN(
        pe_1_1_0_N61) );
  NOR2_X1 pe_1_1_0_U12 ( .A1(pe_1_1_0_n67), .A2(pe_1_1_0_n39), .ZN(
        pe_1_1_0_N62) );
  NOR2_X1 pe_1_1_0_U11 ( .A1(pe_1_1_0_n37), .A2(pe_1_1_0_n67), .ZN(
        pe_1_1_0_N64) );
  NAND2_X1 pe_1_1_0_U10 ( .A1(pe_1_1_0_n44), .A2(pe_1_1_0_n60), .ZN(
        pe_1_1_0_n42) );
  BUF_X1 pe_1_1_0_U9 ( .A(pe_1_1_0_n60), .Z(pe_1_1_0_n55) );
  BUF_X1 pe_1_1_0_U8 ( .A(pe_1_1_0_n60), .Z(pe_1_1_0_n56) );
  INV_X1 pe_1_1_0_U7 ( .A(pe_1_1_0_n69), .ZN(pe_1_1_0_n65) );
  INV_X1 pe_1_1_0_U6 ( .A(pe_1_1_0_n42), .ZN(pe_1_1_0_n89) );
  INV_X1 pe_1_1_0_U5 ( .A(pe_1_1_0_n40), .ZN(pe_1_1_0_n85) );
  INV_X2 pe_1_1_0_U4 ( .A(n81), .ZN(pe_1_1_0_n72) );
  XOR2_X1 pe_1_1_0_U3 ( .A(pe_1_1_0_int_data_0_), .B(int_data_res_1__0__0_), 
        .Z(pe_1_1_0_n1) );
  DFFR_X1 pe_1_1_0_int_q_acc_reg_0_ ( .D(pe_1_1_0_n84), .CK(pe_1_1_0_net6928), 
        .RN(pe_1_1_0_n72), .Q(int_data_res_1__0__0_), .QN(pe_1_1_0_n3) );
  DFFR_X1 pe_1_1_0_int_q_reg_v_reg_0__0_ ( .D(int_data_y_2__0__0_), .CK(
        pe_1_1_0_net6898), .RN(pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_v[20]) );
  DFFR_X1 pe_1_1_0_int_q_reg_v_reg_0__1_ ( .D(int_data_y_2__0__1_), .CK(
        pe_1_1_0_net6898), .RN(pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_v[21]) );
  DFFR_X1 pe_1_1_0_int_q_reg_v_reg_0__2_ ( .D(int_data_y_2__0__2_), .CK(
        pe_1_1_0_net6898), .RN(pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_v[22]) );
  DFFR_X1 pe_1_1_0_int_q_reg_v_reg_0__3_ ( .D(int_data_y_2__0__3_), .CK(
        pe_1_1_0_net6898), .RN(pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_v[23]) );
  DFFR_X1 pe_1_1_0_int_q_reg_v_reg_1__0_ ( .D(int_data_y_2__0__0_), .CK(
        pe_1_1_0_net6903), .RN(pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_v[16]) );
  DFFR_X1 pe_1_1_0_int_q_reg_v_reg_1__1_ ( .D(int_data_y_2__0__1_), .CK(
        pe_1_1_0_net6903), .RN(pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_v[17]) );
  DFFR_X1 pe_1_1_0_int_q_reg_v_reg_1__2_ ( .D(int_data_y_2__0__2_), .CK(
        pe_1_1_0_net6903), .RN(pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_v[18]) );
  DFFR_X1 pe_1_1_0_int_q_reg_v_reg_1__3_ ( .D(int_data_y_2__0__3_), .CK(
        pe_1_1_0_net6903), .RN(pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_v[19]) );
  DFFR_X1 pe_1_1_0_int_q_reg_v_reg_2__0_ ( .D(int_data_y_2__0__0_), .CK(
        pe_1_1_0_net6908), .RN(pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_v[12]) );
  DFFR_X1 pe_1_1_0_int_q_reg_v_reg_2__1_ ( .D(int_data_y_2__0__1_), .CK(
        pe_1_1_0_net6908), .RN(pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_v[13]) );
  DFFR_X1 pe_1_1_0_int_q_reg_v_reg_2__2_ ( .D(int_data_y_2__0__2_), .CK(
        pe_1_1_0_net6908), .RN(pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_v[14]) );
  DFFR_X1 pe_1_1_0_int_q_reg_v_reg_2__3_ ( .D(int_data_y_2__0__3_), .CK(
        pe_1_1_0_net6908), .RN(pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_v[15]) );
  DFFR_X1 pe_1_1_0_int_q_reg_v_reg_3__0_ ( .D(int_data_y_2__0__0_), .CK(
        pe_1_1_0_net6913), .RN(pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_v[8]) );
  DFFR_X1 pe_1_1_0_int_q_reg_v_reg_3__1_ ( .D(int_data_y_2__0__1_), .CK(
        pe_1_1_0_net6913), .RN(pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_v[9]) );
  DFFR_X1 pe_1_1_0_int_q_reg_v_reg_3__2_ ( .D(int_data_y_2__0__2_), .CK(
        pe_1_1_0_net6913), .RN(pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_v[10]) );
  DFFR_X1 pe_1_1_0_int_q_reg_v_reg_3__3_ ( .D(int_data_y_2__0__3_), .CK(
        pe_1_1_0_net6913), .RN(pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_v[11]) );
  DFFR_X1 pe_1_1_0_int_q_reg_v_reg_4__0_ ( .D(int_data_y_2__0__0_), .CK(
        pe_1_1_0_net6918), .RN(pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_v[4]) );
  DFFR_X1 pe_1_1_0_int_q_reg_v_reg_4__1_ ( .D(int_data_y_2__0__1_), .CK(
        pe_1_1_0_net6918), .RN(pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_v[5]) );
  DFFR_X1 pe_1_1_0_int_q_reg_v_reg_4__2_ ( .D(int_data_y_2__0__2_), .CK(
        pe_1_1_0_net6918), .RN(pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_v[6]) );
  DFFR_X1 pe_1_1_0_int_q_reg_v_reg_4__3_ ( .D(int_data_y_2__0__3_), .CK(
        pe_1_1_0_net6918), .RN(pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_v[7]) );
  DFFR_X1 pe_1_1_0_int_q_reg_v_reg_5__0_ ( .D(int_data_y_2__0__0_), .CK(
        pe_1_1_0_net6923), .RN(pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_v[0]) );
  DFFR_X1 pe_1_1_0_int_q_reg_v_reg_5__1_ ( .D(int_data_y_2__0__1_), .CK(
        pe_1_1_0_net6923), .RN(pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_v[1]) );
  DFFR_X1 pe_1_1_0_int_q_reg_v_reg_5__2_ ( .D(int_data_y_2__0__2_), .CK(
        pe_1_1_0_net6923), .RN(pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_v[2]) );
  DFFR_X1 pe_1_1_0_int_q_reg_v_reg_5__3_ ( .D(int_data_y_2__0__3_), .CK(
        pe_1_1_0_net6923), .RN(pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_1_0_int_q_reg_h_reg_0__0_ ( .D(int_data_x_1__1__0_), .SI(
        int_data_y_2__0__0_), .SE(pe_1_1_0_n65), .CK(pe_1_1_0_net6867), .RN(
        pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_1_0_int_q_reg_h_reg_0__1_ ( .D(int_data_x_1__1__1_), .SI(
        int_data_y_2__0__1_), .SE(pe_1_1_0_n65), .CK(pe_1_1_0_net6867), .RN(
        pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_1_0_int_q_reg_h_reg_0__2_ ( .D(int_data_x_1__1__2_), .SI(
        int_data_y_2__0__2_), .SE(pe_1_1_0_n65), .CK(pe_1_1_0_net6867), .RN(
        pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_1_0_int_q_reg_h_reg_0__3_ ( .D(int_data_x_1__1__3_), .SI(
        int_data_y_2__0__3_), .SE(pe_1_1_0_n65), .CK(pe_1_1_0_net6867), .RN(
        pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_1_0_int_q_reg_h_reg_1__0_ ( .D(int_data_x_1__1__0_), .SI(
        int_data_y_2__0__0_), .SE(pe_1_1_0_n65), .CK(pe_1_1_0_net6873), .RN(
        pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_1_0_int_q_reg_h_reg_1__1_ ( .D(int_data_x_1__1__1_), .SI(
        int_data_y_2__0__1_), .SE(pe_1_1_0_n65), .CK(pe_1_1_0_net6873), .RN(
        pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_1_0_int_q_reg_h_reg_1__2_ ( .D(int_data_x_1__1__2_), .SI(
        int_data_y_2__0__2_), .SE(pe_1_1_0_n65), .CK(pe_1_1_0_net6873), .RN(
        pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_1_0_int_q_reg_h_reg_1__3_ ( .D(int_data_x_1__1__3_), .SI(
        int_data_y_2__0__3_), .SE(pe_1_1_0_n65), .CK(pe_1_1_0_net6873), .RN(
        pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_1_0_int_q_reg_h_reg_2__0_ ( .D(int_data_x_1__1__0_), .SI(
        int_data_y_2__0__0_), .SE(pe_1_1_0_n65), .CK(pe_1_1_0_net6878), .RN(
        pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_1_0_int_q_reg_h_reg_2__1_ ( .D(int_data_x_1__1__1_), .SI(
        int_data_y_2__0__1_), .SE(pe_1_1_0_n65), .CK(pe_1_1_0_net6878), .RN(
        pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_1_0_int_q_reg_h_reg_2__2_ ( .D(int_data_x_1__1__2_), .SI(
        int_data_y_2__0__2_), .SE(pe_1_1_0_n65), .CK(pe_1_1_0_net6878), .RN(
        pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_1_0_int_q_reg_h_reg_2__3_ ( .D(int_data_x_1__1__3_), .SI(
        int_data_y_2__0__3_), .SE(pe_1_1_0_n65), .CK(pe_1_1_0_net6878), .RN(
        pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_1_0_int_q_reg_h_reg_3__0_ ( .D(int_data_x_1__1__0_), .SI(
        int_data_y_2__0__0_), .SE(pe_1_1_0_n65), .CK(pe_1_1_0_net6883), .RN(
        pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_1_0_int_q_reg_h_reg_3__1_ ( .D(int_data_x_1__1__1_), .SI(
        int_data_y_2__0__1_), .SE(pe_1_1_0_n65), .CK(pe_1_1_0_net6883), .RN(
        pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_1_0_int_q_reg_h_reg_3__2_ ( .D(int_data_x_1__1__2_), .SI(
        int_data_y_2__0__2_), .SE(pe_1_1_0_n65), .CK(pe_1_1_0_net6883), .RN(
        pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_1_0_int_q_reg_h_reg_3__3_ ( .D(int_data_x_1__1__3_), .SI(
        int_data_y_2__0__3_), .SE(pe_1_1_0_n65), .CK(pe_1_1_0_net6883), .RN(
        pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_1_0_int_q_reg_h_reg_4__0_ ( .D(int_data_x_1__1__0_), .SI(
        int_data_y_2__0__0_), .SE(pe_1_1_0_n66), .CK(pe_1_1_0_net6888), .RN(
        pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_1_0_int_q_reg_h_reg_4__1_ ( .D(int_data_x_1__1__1_), .SI(
        int_data_y_2__0__1_), .SE(pe_1_1_0_n66), .CK(pe_1_1_0_net6888), .RN(
        pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_1_0_int_q_reg_h_reg_4__2_ ( .D(int_data_x_1__1__2_), .SI(
        int_data_y_2__0__2_), .SE(pe_1_1_0_n66), .CK(pe_1_1_0_net6888), .RN(
        pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_1_0_int_q_reg_h_reg_4__3_ ( .D(int_data_x_1__1__3_), .SI(
        int_data_y_2__0__3_), .SE(pe_1_1_0_n66), .CK(pe_1_1_0_net6888), .RN(
        pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_1_0_int_q_reg_h_reg_5__0_ ( .D(int_data_x_1__1__0_), .SI(
        int_data_y_2__0__0_), .SE(pe_1_1_0_n66), .CK(pe_1_1_0_net6893), .RN(
        pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_1_0_int_q_reg_h_reg_5__1_ ( .D(int_data_x_1__1__1_), .SI(
        int_data_y_2__0__1_), .SE(pe_1_1_0_n66), .CK(pe_1_1_0_net6893), .RN(
        pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_1_0_int_q_reg_h_reg_5__2_ ( .D(int_data_x_1__1__2_), .SI(
        int_data_y_2__0__2_), .SE(pe_1_1_0_n66), .CK(pe_1_1_0_net6893), .RN(
        pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_1_0_int_q_reg_h_reg_5__3_ ( .D(int_data_x_1__1__3_), .SI(
        int_data_y_2__0__3_), .SE(pe_1_1_0_n66), .CK(pe_1_1_0_net6893), .RN(
        pe_1_1_0_n72), .Q(pe_1_1_0_int_q_reg_h[3]) );
  FA_X1 pe_1_1_0_sub_81_U2_7 ( .A(int_data_res_1__0__7_), .B(pe_1_1_0_n76), 
        .CI(pe_1_1_0_sub_81_carry[7]), .S(pe_1_1_0_N77) );
  FA_X1 pe_1_1_0_sub_81_U2_6 ( .A(int_data_res_1__0__6_), .B(pe_1_1_0_n76), 
        .CI(pe_1_1_0_sub_81_carry[6]), .CO(pe_1_1_0_sub_81_carry[7]), .S(
        pe_1_1_0_N76) );
  FA_X1 pe_1_1_0_sub_81_U2_5 ( .A(int_data_res_1__0__5_), .B(pe_1_1_0_n76), 
        .CI(pe_1_1_0_sub_81_carry[5]), .CO(pe_1_1_0_sub_81_carry[6]), .S(
        pe_1_1_0_N75) );
  FA_X1 pe_1_1_0_sub_81_U2_4 ( .A(int_data_res_1__0__4_), .B(pe_1_1_0_n76), 
        .CI(pe_1_1_0_sub_81_carry[4]), .CO(pe_1_1_0_sub_81_carry[5]), .S(
        pe_1_1_0_N74) );
  FA_X1 pe_1_1_0_sub_81_U2_3 ( .A(int_data_res_1__0__3_), .B(pe_1_1_0_n76), 
        .CI(pe_1_1_0_sub_81_carry[3]), .CO(pe_1_1_0_sub_81_carry[4]), .S(
        pe_1_1_0_N73) );
  FA_X1 pe_1_1_0_sub_81_U2_2 ( .A(int_data_res_1__0__2_), .B(pe_1_1_0_n75), 
        .CI(pe_1_1_0_sub_81_carry[2]), .CO(pe_1_1_0_sub_81_carry[3]), .S(
        pe_1_1_0_N72) );
  FA_X1 pe_1_1_0_sub_81_U2_1 ( .A(int_data_res_1__0__1_), .B(pe_1_1_0_n74), 
        .CI(pe_1_1_0_sub_81_carry[1]), .CO(pe_1_1_0_sub_81_carry[2]), .S(
        pe_1_1_0_N71) );
  FA_X1 pe_1_1_0_add_83_U1_7 ( .A(int_data_res_1__0__7_), .B(
        pe_1_1_0_int_data_3_), .CI(pe_1_1_0_add_83_carry[7]), .S(pe_1_1_0_N85)
         );
  FA_X1 pe_1_1_0_add_83_U1_6 ( .A(int_data_res_1__0__6_), .B(
        pe_1_1_0_int_data_3_), .CI(pe_1_1_0_add_83_carry[6]), .CO(
        pe_1_1_0_add_83_carry[7]), .S(pe_1_1_0_N84) );
  FA_X1 pe_1_1_0_add_83_U1_5 ( .A(int_data_res_1__0__5_), .B(
        pe_1_1_0_int_data_3_), .CI(pe_1_1_0_add_83_carry[5]), .CO(
        pe_1_1_0_add_83_carry[6]), .S(pe_1_1_0_N83) );
  FA_X1 pe_1_1_0_add_83_U1_4 ( .A(int_data_res_1__0__4_), .B(
        pe_1_1_0_int_data_3_), .CI(pe_1_1_0_add_83_carry[4]), .CO(
        pe_1_1_0_add_83_carry[5]), .S(pe_1_1_0_N82) );
  FA_X1 pe_1_1_0_add_83_U1_3 ( .A(int_data_res_1__0__3_), .B(
        pe_1_1_0_int_data_3_), .CI(pe_1_1_0_add_83_carry[3]), .CO(
        pe_1_1_0_add_83_carry[4]), .S(pe_1_1_0_N81) );
  FA_X1 pe_1_1_0_add_83_U1_2 ( .A(int_data_res_1__0__2_), .B(
        pe_1_1_0_int_data_2_), .CI(pe_1_1_0_add_83_carry[2]), .CO(
        pe_1_1_0_add_83_carry[3]), .S(pe_1_1_0_N80) );
  FA_X1 pe_1_1_0_add_83_U1_1 ( .A(int_data_res_1__0__1_), .B(
        pe_1_1_0_int_data_1_), .CI(pe_1_1_0_n2), .CO(pe_1_1_0_add_83_carry[2]), 
        .S(pe_1_1_0_N79) );
  NAND3_X1 pe_1_1_0_U56 ( .A1(pe_1_1_0_n60), .A2(pe_1_1_0_n43), .A3(
        pe_1_1_0_n62), .ZN(pe_1_1_0_n40) );
  NAND3_X1 pe_1_1_0_U55 ( .A1(pe_1_1_0_n43), .A2(pe_1_1_0_n61), .A3(
        pe_1_1_0_n62), .ZN(pe_1_1_0_n39) );
  NAND3_X1 pe_1_1_0_U54 ( .A1(pe_1_1_0_n43), .A2(pe_1_1_0_n63), .A3(
        pe_1_1_0_n60), .ZN(pe_1_1_0_n38) );
  NAND3_X1 pe_1_1_0_U53 ( .A1(pe_1_1_0_n61), .A2(pe_1_1_0_n63), .A3(
        pe_1_1_0_n43), .ZN(pe_1_1_0_n37) );
  DFFR_X1 pe_1_1_0_int_q_acc_reg_6_ ( .D(pe_1_1_0_n78), .CK(pe_1_1_0_net6928), 
        .RN(pe_1_1_0_n71), .Q(int_data_res_1__0__6_) );
  DFFR_X1 pe_1_1_0_int_q_acc_reg_5_ ( .D(pe_1_1_0_n79), .CK(pe_1_1_0_net6928), 
        .RN(pe_1_1_0_n71), .Q(int_data_res_1__0__5_) );
  DFFR_X1 pe_1_1_0_int_q_acc_reg_4_ ( .D(pe_1_1_0_n80), .CK(pe_1_1_0_net6928), 
        .RN(pe_1_1_0_n71), .Q(int_data_res_1__0__4_) );
  DFFR_X1 pe_1_1_0_int_q_acc_reg_3_ ( .D(pe_1_1_0_n81), .CK(pe_1_1_0_net6928), 
        .RN(pe_1_1_0_n71), .Q(int_data_res_1__0__3_) );
  DFFR_X1 pe_1_1_0_int_q_acc_reg_2_ ( .D(pe_1_1_0_n82), .CK(pe_1_1_0_net6928), 
        .RN(pe_1_1_0_n71), .Q(int_data_res_1__0__2_) );
  DFFR_X1 pe_1_1_0_int_q_acc_reg_1_ ( .D(pe_1_1_0_n83), .CK(pe_1_1_0_net6928), 
        .RN(pe_1_1_0_n71), .Q(int_data_res_1__0__1_) );
  DFFR_X1 pe_1_1_0_int_q_acc_reg_7_ ( .D(pe_1_1_0_n77), .CK(pe_1_1_0_net6928), 
        .RN(pe_1_1_0_n71), .Q(int_data_res_1__0__7_) );
  CLKGATETST_X1 pe_1_1_0_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_1_0_n88), .SE(1'b0), .GCK(pe_1_1_0_net6867) );
  CLKGATETST_X1 pe_1_1_0_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_1_0_n87), .SE(1'b0), .GCK(pe_1_1_0_net6873) );
  CLKGATETST_X1 pe_1_1_0_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_1_0_n86), .SE(1'b0), .GCK(pe_1_1_0_net6878) );
  CLKGATETST_X1 pe_1_1_0_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_1_0_n85), .SE(1'b0), .GCK(pe_1_1_0_net6883) );
  CLKGATETST_X1 pe_1_1_0_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_1_0_n90), .SE(1'b0), .GCK(pe_1_1_0_net6888) );
  CLKGATETST_X1 pe_1_1_0_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_1_0_n89), .SE(1'b0), .GCK(pe_1_1_0_net6893) );
  CLKGATETST_X1 pe_1_1_0_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_1_0_N64), .SE(1'b0), .GCK(pe_1_1_0_net6898) );
  CLKGATETST_X1 pe_1_1_0_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_1_0_N63), .SE(1'b0), .GCK(pe_1_1_0_net6903) );
  CLKGATETST_X1 pe_1_1_0_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_1_0_N62), .SE(1'b0), .GCK(pe_1_1_0_net6908) );
  CLKGATETST_X1 pe_1_1_0_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_1_0_N61), .SE(1'b0), .GCK(pe_1_1_0_net6913) );
  CLKGATETST_X1 pe_1_1_0_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_1_0_N60), .SE(1'b0), .GCK(pe_1_1_0_net6918) );
  CLKGATETST_X1 pe_1_1_0_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_1_0_N59), .SE(1'b0), .GCK(pe_1_1_0_net6923) );
  CLKGATETST_X1 pe_1_1_0_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_1_0_N90), .SE(1'b0), .GCK(pe_1_1_0_net6928) );
  CLKBUF_X1 pe_1_1_1_U112 ( .A(pe_1_1_1_n72), .Z(pe_1_1_1_n71) );
  INV_X1 pe_1_1_1_U111 ( .A(n73), .ZN(pe_1_1_1_n70) );
  INV_X1 pe_1_1_1_U110 ( .A(n65), .ZN(pe_1_1_1_n69) );
  INV_X1 pe_1_1_1_U109 ( .A(n65), .ZN(pe_1_1_1_n68) );
  INV_X1 pe_1_1_1_U108 ( .A(n65), .ZN(pe_1_1_1_n67) );
  INV_X1 pe_1_1_1_U107 ( .A(pe_1_1_1_n69), .ZN(pe_1_1_1_n66) );
  INV_X1 pe_1_1_1_U106 ( .A(pe_1_1_1_n63), .ZN(pe_1_1_1_n62) );
  INV_X1 pe_1_1_1_U105 ( .A(pe_1_1_1_n61), .ZN(pe_1_1_1_n60) );
  INV_X1 pe_1_1_1_U104 ( .A(n25), .ZN(pe_1_1_1_n59) );
  INV_X1 pe_1_1_1_U103 ( .A(pe_1_1_1_n59), .ZN(pe_1_1_1_n58) );
  INV_X1 pe_1_1_1_U102 ( .A(n17), .ZN(pe_1_1_1_n57) );
  MUX2_X1 pe_1_1_1_U101 ( .A(pe_1_1_1_n54), .B(pe_1_1_1_n51), .S(n44), .Z(
        int_data_x_1__1__3_) );
  MUX2_X1 pe_1_1_1_U100 ( .A(pe_1_1_1_n53), .B(pe_1_1_1_n52), .S(pe_1_1_1_n62), 
        .Z(pe_1_1_1_n54) );
  MUX2_X1 pe_1_1_1_U99 ( .A(pe_1_1_1_int_q_reg_h[23]), .B(
        pe_1_1_1_int_q_reg_h[19]), .S(pe_1_1_1_n56), .Z(pe_1_1_1_n53) );
  MUX2_X1 pe_1_1_1_U98 ( .A(pe_1_1_1_int_q_reg_h[15]), .B(
        pe_1_1_1_int_q_reg_h[11]), .S(pe_1_1_1_n56), .Z(pe_1_1_1_n52) );
  MUX2_X1 pe_1_1_1_U97 ( .A(pe_1_1_1_int_q_reg_h[7]), .B(
        pe_1_1_1_int_q_reg_h[3]), .S(pe_1_1_1_n56), .Z(pe_1_1_1_n51) );
  MUX2_X1 pe_1_1_1_U96 ( .A(pe_1_1_1_n50), .B(pe_1_1_1_n47), .S(n44), .Z(
        int_data_x_1__1__2_) );
  MUX2_X1 pe_1_1_1_U95 ( .A(pe_1_1_1_n49), .B(pe_1_1_1_n48), .S(pe_1_1_1_n62), 
        .Z(pe_1_1_1_n50) );
  MUX2_X1 pe_1_1_1_U94 ( .A(pe_1_1_1_int_q_reg_h[22]), .B(
        pe_1_1_1_int_q_reg_h[18]), .S(pe_1_1_1_n56), .Z(pe_1_1_1_n49) );
  MUX2_X1 pe_1_1_1_U93 ( .A(pe_1_1_1_int_q_reg_h[14]), .B(
        pe_1_1_1_int_q_reg_h[10]), .S(pe_1_1_1_n56), .Z(pe_1_1_1_n48) );
  MUX2_X1 pe_1_1_1_U92 ( .A(pe_1_1_1_int_q_reg_h[6]), .B(
        pe_1_1_1_int_q_reg_h[2]), .S(pe_1_1_1_n56), .Z(pe_1_1_1_n47) );
  MUX2_X1 pe_1_1_1_U91 ( .A(pe_1_1_1_n46), .B(pe_1_1_1_n24), .S(n44), .Z(
        int_data_x_1__1__1_) );
  MUX2_X1 pe_1_1_1_U90 ( .A(pe_1_1_1_n45), .B(pe_1_1_1_n25), .S(pe_1_1_1_n62), 
        .Z(pe_1_1_1_n46) );
  MUX2_X1 pe_1_1_1_U89 ( .A(pe_1_1_1_int_q_reg_h[21]), .B(
        pe_1_1_1_int_q_reg_h[17]), .S(pe_1_1_1_n56), .Z(pe_1_1_1_n45) );
  MUX2_X1 pe_1_1_1_U88 ( .A(pe_1_1_1_int_q_reg_h[13]), .B(
        pe_1_1_1_int_q_reg_h[9]), .S(pe_1_1_1_n56), .Z(pe_1_1_1_n25) );
  MUX2_X1 pe_1_1_1_U87 ( .A(pe_1_1_1_int_q_reg_h[5]), .B(
        pe_1_1_1_int_q_reg_h[1]), .S(pe_1_1_1_n56), .Z(pe_1_1_1_n24) );
  MUX2_X1 pe_1_1_1_U86 ( .A(pe_1_1_1_n23), .B(pe_1_1_1_n20), .S(n44), .Z(
        int_data_x_1__1__0_) );
  MUX2_X1 pe_1_1_1_U85 ( .A(pe_1_1_1_n22), .B(pe_1_1_1_n21), .S(pe_1_1_1_n62), 
        .Z(pe_1_1_1_n23) );
  MUX2_X1 pe_1_1_1_U84 ( .A(pe_1_1_1_int_q_reg_h[20]), .B(
        pe_1_1_1_int_q_reg_h[16]), .S(pe_1_1_1_n56), .Z(pe_1_1_1_n22) );
  MUX2_X1 pe_1_1_1_U83 ( .A(pe_1_1_1_int_q_reg_h[12]), .B(
        pe_1_1_1_int_q_reg_h[8]), .S(pe_1_1_1_n56), .Z(pe_1_1_1_n21) );
  MUX2_X1 pe_1_1_1_U82 ( .A(pe_1_1_1_int_q_reg_h[4]), .B(
        pe_1_1_1_int_q_reg_h[0]), .S(pe_1_1_1_n56), .Z(pe_1_1_1_n20) );
  MUX2_X1 pe_1_1_1_U81 ( .A(pe_1_1_1_n19), .B(pe_1_1_1_n16), .S(n44), .Z(
        int_data_y_1__1__3_) );
  MUX2_X1 pe_1_1_1_U80 ( .A(pe_1_1_1_n18), .B(pe_1_1_1_n17), .S(pe_1_1_1_n62), 
        .Z(pe_1_1_1_n19) );
  MUX2_X1 pe_1_1_1_U79 ( .A(pe_1_1_1_int_q_reg_v[23]), .B(
        pe_1_1_1_int_q_reg_v[19]), .S(pe_1_1_1_n55), .Z(pe_1_1_1_n18) );
  MUX2_X1 pe_1_1_1_U78 ( .A(pe_1_1_1_int_q_reg_v[15]), .B(
        pe_1_1_1_int_q_reg_v[11]), .S(pe_1_1_1_n55), .Z(pe_1_1_1_n17) );
  MUX2_X1 pe_1_1_1_U77 ( .A(pe_1_1_1_int_q_reg_v[7]), .B(
        pe_1_1_1_int_q_reg_v[3]), .S(pe_1_1_1_n55), .Z(pe_1_1_1_n16) );
  MUX2_X1 pe_1_1_1_U76 ( .A(pe_1_1_1_n15), .B(pe_1_1_1_n12), .S(n44), .Z(
        int_data_y_1__1__2_) );
  MUX2_X1 pe_1_1_1_U75 ( .A(pe_1_1_1_n14), .B(pe_1_1_1_n13), .S(pe_1_1_1_n62), 
        .Z(pe_1_1_1_n15) );
  MUX2_X1 pe_1_1_1_U74 ( .A(pe_1_1_1_int_q_reg_v[22]), .B(
        pe_1_1_1_int_q_reg_v[18]), .S(pe_1_1_1_n55), .Z(pe_1_1_1_n14) );
  MUX2_X1 pe_1_1_1_U73 ( .A(pe_1_1_1_int_q_reg_v[14]), .B(
        pe_1_1_1_int_q_reg_v[10]), .S(pe_1_1_1_n55), .Z(pe_1_1_1_n13) );
  MUX2_X1 pe_1_1_1_U72 ( .A(pe_1_1_1_int_q_reg_v[6]), .B(
        pe_1_1_1_int_q_reg_v[2]), .S(pe_1_1_1_n55), .Z(pe_1_1_1_n12) );
  MUX2_X1 pe_1_1_1_U71 ( .A(pe_1_1_1_n11), .B(pe_1_1_1_n8), .S(n44), .Z(
        int_data_y_1__1__1_) );
  MUX2_X1 pe_1_1_1_U70 ( .A(pe_1_1_1_n10), .B(pe_1_1_1_n9), .S(pe_1_1_1_n62), 
        .Z(pe_1_1_1_n11) );
  MUX2_X1 pe_1_1_1_U69 ( .A(pe_1_1_1_int_q_reg_v[21]), .B(
        pe_1_1_1_int_q_reg_v[17]), .S(pe_1_1_1_n55), .Z(pe_1_1_1_n10) );
  MUX2_X1 pe_1_1_1_U68 ( .A(pe_1_1_1_int_q_reg_v[13]), .B(
        pe_1_1_1_int_q_reg_v[9]), .S(pe_1_1_1_n55), .Z(pe_1_1_1_n9) );
  MUX2_X1 pe_1_1_1_U67 ( .A(pe_1_1_1_int_q_reg_v[5]), .B(
        pe_1_1_1_int_q_reg_v[1]), .S(pe_1_1_1_n55), .Z(pe_1_1_1_n8) );
  MUX2_X1 pe_1_1_1_U66 ( .A(pe_1_1_1_n7), .B(pe_1_1_1_n4), .S(n44), .Z(
        int_data_y_1__1__0_) );
  MUX2_X1 pe_1_1_1_U65 ( .A(pe_1_1_1_n6), .B(pe_1_1_1_n5), .S(pe_1_1_1_n62), 
        .Z(pe_1_1_1_n7) );
  MUX2_X1 pe_1_1_1_U64 ( .A(pe_1_1_1_int_q_reg_v[20]), .B(
        pe_1_1_1_int_q_reg_v[16]), .S(pe_1_1_1_n55), .Z(pe_1_1_1_n6) );
  MUX2_X1 pe_1_1_1_U63 ( .A(pe_1_1_1_int_q_reg_v[12]), .B(
        pe_1_1_1_int_q_reg_v[8]), .S(pe_1_1_1_n55), .Z(pe_1_1_1_n5) );
  MUX2_X1 pe_1_1_1_U62 ( .A(pe_1_1_1_int_q_reg_v[4]), .B(
        pe_1_1_1_int_q_reg_v[0]), .S(pe_1_1_1_n55), .Z(pe_1_1_1_n4) );
  AOI222_X1 pe_1_1_1_U61 ( .A1(int_data_res_2__1__2_), .A2(pe_1_1_1_n64), .B1(
        pe_1_1_1_N80), .B2(pe_1_1_1_n27), .C1(pe_1_1_1_N72), .C2(pe_1_1_1_n28), 
        .ZN(pe_1_1_1_n33) );
  INV_X1 pe_1_1_1_U60 ( .A(pe_1_1_1_n33), .ZN(pe_1_1_1_n82) );
  AOI222_X1 pe_1_1_1_U59 ( .A1(int_data_res_2__1__6_), .A2(pe_1_1_1_n64), .B1(
        pe_1_1_1_N84), .B2(pe_1_1_1_n27), .C1(pe_1_1_1_N76), .C2(pe_1_1_1_n28), 
        .ZN(pe_1_1_1_n29) );
  INV_X1 pe_1_1_1_U58 ( .A(pe_1_1_1_n29), .ZN(pe_1_1_1_n78) );
  XNOR2_X1 pe_1_1_1_U57 ( .A(pe_1_1_1_n73), .B(int_data_res_1__1__0_), .ZN(
        pe_1_1_1_N70) );
  AOI222_X1 pe_1_1_1_U52 ( .A1(int_data_res_2__1__0_), .A2(pe_1_1_1_n64), .B1(
        pe_1_1_1_n1), .B2(pe_1_1_1_n27), .C1(pe_1_1_1_N70), .C2(pe_1_1_1_n28), 
        .ZN(pe_1_1_1_n35) );
  INV_X1 pe_1_1_1_U51 ( .A(pe_1_1_1_n35), .ZN(pe_1_1_1_n84) );
  AOI222_X1 pe_1_1_1_U50 ( .A1(int_data_res_2__1__1_), .A2(pe_1_1_1_n64), .B1(
        pe_1_1_1_N79), .B2(pe_1_1_1_n27), .C1(pe_1_1_1_N71), .C2(pe_1_1_1_n28), 
        .ZN(pe_1_1_1_n34) );
  INV_X1 pe_1_1_1_U49 ( .A(pe_1_1_1_n34), .ZN(pe_1_1_1_n83) );
  AOI222_X1 pe_1_1_1_U48 ( .A1(int_data_res_2__1__3_), .A2(pe_1_1_1_n64), .B1(
        pe_1_1_1_N81), .B2(pe_1_1_1_n27), .C1(pe_1_1_1_N73), .C2(pe_1_1_1_n28), 
        .ZN(pe_1_1_1_n32) );
  INV_X1 pe_1_1_1_U47 ( .A(pe_1_1_1_n32), .ZN(pe_1_1_1_n81) );
  AOI222_X1 pe_1_1_1_U46 ( .A1(int_data_res_2__1__4_), .A2(pe_1_1_1_n64), .B1(
        pe_1_1_1_N82), .B2(pe_1_1_1_n27), .C1(pe_1_1_1_N74), .C2(pe_1_1_1_n28), 
        .ZN(pe_1_1_1_n31) );
  INV_X1 pe_1_1_1_U45 ( .A(pe_1_1_1_n31), .ZN(pe_1_1_1_n80) );
  AOI222_X1 pe_1_1_1_U44 ( .A1(int_data_res_2__1__5_), .A2(pe_1_1_1_n64), .B1(
        pe_1_1_1_N83), .B2(pe_1_1_1_n27), .C1(pe_1_1_1_N75), .C2(pe_1_1_1_n28), 
        .ZN(pe_1_1_1_n30) );
  INV_X1 pe_1_1_1_U43 ( .A(pe_1_1_1_n30), .ZN(pe_1_1_1_n79) );
  NAND2_X1 pe_1_1_1_U42 ( .A1(pe_1_1_1_int_data_0_), .A2(pe_1_1_1_n3), .ZN(
        pe_1_1_1_sub_81_carry[1]) );
  INV_X1 pe_1_1_1_U41 ( .A(pe_1_1_1_int_data_1_), .ZN(pe_1_1_1_n74) );
  INV_X1 pe_1_1_1_U40 ( .A(pe_1_1_1_int_data_2_), .ZN(pe_1_1_1_n75) );
  AND2_X1 pe_1_1_1_U39 ( .A1(pe_1_1_1_int_data_0_), .A2(int_data_res_1__1__0_), 
        .ZN(pe_1_1_1_n2) );
  AOI222_X1 pe_1_1_1_U38 ( .A1(pe_1_1_1_n64), .A2(int_data_res_2__1__7_), .B1(
        pe_1_1_1_N85), .B2(pe_1_1_1_n27), .C1(pe_1_1_1_N77), .C2(pe_1_1_1_n28), 
        .ZN(pe_1_1_1_n26) );
  INV_X1 pe_1_1_1_U37 ( .A(pe_1_1_1_n26), .ZN(pe_1_1_1_n77) );
  NOR3_X1 pe_1_1_1_U36 ( .A1(pe_1_1_1_n59), .A2(pe_1_1_1_n65), .A3(int_ckg[54]), .ZN(pe_1_1_1_n36) );
  OR2_X1 pe_1_1_1_U35 ( .A1(pe_1_1_1_n36), .A2(pe_1_1_1_n64), .ZN(pe_1_1_1_N90) );
  INV_X1 pe_1_1_1_U34 ( .A(n37), .ZN(pe_1_1_1_n63) );
  AND2_X1 pe_1_1_1_U33 ( .A1(int_data_x_1__1__2_), .A2(pe_1_1_1_n58), .ZN(
        pe_1_1_1_int_data_2_) );
  AND2_X1 pe_1_1_1_U32 ( .A1(int_data_x_1__1__1_), .A2(pe_1_1_1_n58), .ZN(
        pe_1_1_1_int_data_1_) );
  AND2_X1 pe_1_1_1_U31 ( .A1(int_data_x_1__1__3_), .A2(pe_1_1_1_n58), .ZN(
        pe_1_1_1_int_data_3_) );
  BUF_X1 pe_1_1_1_U30 ( .A(n59), .Z(pe_1_1_1_n64) );
  INV_X1 pe_1_1_1_U29 ( .A(n31), .ZN(pe_1_1_1_n61) );
  AND2_X1 pe_1_1_1_U28 ( .A1(int_data_x_1__1__0_), .A2(pe_1_1_1_n58), .ZN(
        pe_1_1_1_int_data_0_) );
  NAND2_X1 pe_1_1_1_U27 ( .A1(pe_1_1_1_n44), .A2(pe_1_1_1_n61), .ZN(
        pe_1_1_1_n41) );
  AND3_X1 pe_1_1_1_U26 ( .A1(n73), .A2(pe_1_1_1_n63), .A3(n44), .ZN(
        pe_1_1_1_n44) );
  INV_X1 pe_1_1_1_U25 ( .A(pe_1_1_1_int_data_3_), .ZN(pe_1_1_1_n76) );
  NOR2_X1 pe_1_1_1_U24 ( .A1(pe_1_1_1_n70), .A2(n44), .ZN(pe_1_1_1_n43) );
  NOR2_X1 pe_1_1_1_U23 ( .A1(pe_1_1_1_n57), .A2(pe_1_1_1_n64), .ZN(
        pe_1_1_1_n28) );
  NOR2_X1 pe_1_1_1_U22 ( .A1(n17), .A2(pe_1_1_1_n64), .ZN(pe_1_1_1_n27) );
  INV_X1 pe_1_1_1_U21 ( .A(pe_1_1_1_int_data_0_), .ZN(pe_1_1_1_n73) );
  INV_X1 pe_1_1_1_U20 ( .A(pe_1_1_1_n41), .ZN(pe_1_1_1_n90) );
  INV_X1 pe_1_1_1_U19 ( .A(pe_1_1_1_n37), .ZN(pe_1_1_1_n88) );
  INV_X1 pe_1_1_1_U18 ( .A(pe_1_1_1_n38), .ZN(pe_1_1_1_n87) );
  INV_X1 pe_1_1_1_U17 ( .A(pe_1_1_1_n39), .ZN(pe_1_1_1_n86) );
  NOR2_X1 pe_1_1_1_U16 ( .A1(pe_1_1_1_n68), .A2(pe_1_1_1_n42), .ZN(
        pe_1_1_1_N59) );
  NOR2_X1 pe_1_1_1_U15 ( .A1(pe_1_1_1_n68), .A2(pe_1_1_1_n41), .ZN(
        pe_1_1_1_N60) );
  NOR2_X1 pe_1_1_1_U14 ( .A1(pe_1_1_1_n68), .A2(pe_1_1_1_n38), .ZN(
        pe_1_1_1_N63) );
  NOR2_X1 pe_1_1_1_U13 ( .A1(pe_1_1_1_n67), .A2(pe_1_1_1_n40), .ZN(
        pe_1_1_1_N61) );
  NOR2_X1 pe_1_1_1_U12 ( .A1(pe_1_1_1_n67), .A2(pe_1_1_1_n39), .ZN(
        pe_1_1_1_N62) );
  NOR2_X1 pe_1_1_1_U11 ( .A1(pe_1_1_1_n37), .A2(pe_1_1_1_n67), .ZN(
        pe_1_1_1_N64) );
  NAND2_X1 pe_1_1_1_U10 ( .A1(pe_1_1_1_n44), .A2(pe_1_1_1_n60), .ZN(
        pe_1_1_1_n42) );
  BUF_X1 pe_1_1_1_U9 ( .A(pe_1_1_1_n60), .Z(pe_1_1_1_n55) );
  INV_X1 pe_1_1_1_U8 ( .A(pe_1_1_1_n69), .ZN(pe_1_1_1_n65) );
  BUF_X1 pe_1_1_1_U7 ( .A(pe_1_1_1_n60), .Z(pe_1_1_1_n56) );
  INV_X1 pe_1_1_1_U6 ( .A(pe_1_1_1_n42), .ZN(pe_1_1_1_n89) );
  INV_X1 pe_1_1_1_U5 ( .A(pe_1_1_1_n40), .ZN(pe_1_1_1_n85) );
  INV_X2 pe_1_1_1_U4 ( .A(n81), .ZN(pe_1_1_1_n72) );
  XOR2_X1 pe_1_1_1_U3 ( .A(pe_1_1_1_int_data_0_), .B(int_data_res_1__1__0_), 
        .Z(pe_1_1_1_n1) );
  DFFR_X1 pe_1_1_1_int_q_acc_reg_0_ ( .D(pe_1_1_1_n84), .CK(pe_1_1_1_net6850), 
        .RN(pe_1_1_1_n72), .Q(int_data_res_1__1__0_), .QN(pe_1_1_1_n3) );
  DFFR_X1 pe_1_1_1_int_q_reg_v_reg_0__0_ ( .D(int_data_y_2__1__0_), .CK(
        pe_1_1_1_net6820), .RN(pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_v[20]) );
  DFFR_X1 pe_1_1_1_int_q_reg_v_reg_0__1_ ( .D(int_data_y_2__1__1_), .CK(
        pe_1_1_1_net6820), .RN(pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_v[21]) );
  DFFR_X1 pe_1_1_1_int_q_reg_v_reg_0__2_ ( .D(int_data_y_2__1__2_), .CK(
        pe_1_1_1_net6820), .RN(pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_v[22]) );
  DFFR_X1 pe_1_1_1_int_q_reg_v_reg_0__3_ ( .D(int_data_y_2__1__3_), .CK(
        pe_1_1_1_net6820), .RN(pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_v[23]) );
  DFFR_X1 pe_1_1_1_int_q_reg_v_reg_1__0_ ( .D(int_data_y_2__1__0_), .CK(
        pe_1_1_1_net6825), .RN(pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_v[16]) );
  DFFR_X1 pe_1_1_1_int_q_reg_v_reg_1__1_ ( .D(int_data_y_2__1__1_), .CK(
        pe_1_1_1_net6825), .RN(pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_v[17]) );
  DFFR_X1 pe_1_1_1_int_q_reg_v_reg_1__2_ ( .D(int_data_y_2__1__2_), .CK(
        pe_1_1_1_net6825), .RN(pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_v[18]) );
  DFFR_X1 pe_1_1_1_int_q_reg_v_reg_1__3_ ( .D(int_data_y_2__1__3_), .CK(
        pe_1_1_1_net6825), .RN(pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_v[19]) );
  DFFR_X1 pe_1_1_1_int_q_reg_v_reg_2__0_ ( .D(int_data_y_2__1__0_), .CK(
        pe_1_1_1_net6830), .RN(pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_v[12]) );
  DFFR_X1 pe_1_1_1_int_q_reg_v_reg_2__1_ ( .D(int_data_y_2__1__1_), .CK(
        pe_1_1_1_net6830), .RN(pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_v[13]) );
  DFFR_X1 pe_1_1_1_int_q_reg_v_reg_2__2_ ( .D(int_data_y_2__1__2_), .CK(
        pe_1_1_1_net6830), .RN(pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_v[14]) );
  DFFR_X1 pe_1_1_1_int_q_reg_v_reg_2__3_ ( .D(int_data_y_2__1__3_), .CK(
        pe_1_1_1_net6830), .RN(pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_v[15]) );
  DFFR_X1 pe_1_1_1_int_q_reg_v_reg_3__0_ ( .D(int_data_y_2__1__0_), .CK(
        pe_1_1_1_net6835), .RN(pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_v[8]) );
  DFFR_X1 pe_1_1_1_int_q_reg_v_reg_3__1_ ( .D(int_data_y_2__1__1_), .CK(
        pe_1_1_1_net6835), .RN(pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_v[9]) );
  DFFR_X1 pe_1_1_1_int_q_reg_v_reg_3__2_ ( .D(int_data_y_2__1__2_), .CK(
        pe_1_1_1_net6835), .RN(pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_v[10]) );
  DFFR_X1 pe_1_1_1_int_q_reg_v_reg_3__3_ ( .D(int_data_y_2__1__3_), .CK(
        pe_1_1_1_net6835), .RN(pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_v[11]) );
  DFFR_X1 pe_1_1_1_int_q_reg_v_reg_4__0_ ( .D(int_data_y_2__1__0_), .CK(
        pe_1_1_1_net6840), .RN(pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_v[4]) );
  DFFR_X1 pe_1_1_1_int_q_reg_v_reg_4__1_ ( .D(int_data_y_2__1__1_), .CK(
        pe_1_1_1_net6840), .RN(pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_v[5]) );
  DFFR_X1 pe_1_1_1_int_q_reg_v_reg_4__2_ ( .D(int_data_y_2__1__2_), .CK(
        pe_1_1_1_net6840), .RN(pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_v[6]) );
  DFFR_X1 pe_1_1_1_int_q_reg_v_reg_4__3_ ( .D(int_data_y_2__1__3_), .CK(
        pe_1_1_1_net6840), .RN(pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_v[7]) );
  DFFR_X1 pe_1_1_1_int_q_reg_v_reg_5__0_ ( .D(int_data_y_2__1__0_), .CK(
        pe_1_1_1_net6845), .RN(pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_v[0]) );
  DFFR_X1 pe_1_1_1_int_q_reg_v_reg_5__1_ ( .D(int_data_y_2__1__1_), .CK(
        pe_1_1_1_net6845), .RN(pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_v[1]) );
  DFFR_X1 pe_1_1_1_int_q_reg_v_reg_5__2_ ( .D(int_data_y_2__1__2_), .CK(
        pe_1_1_1_net6845), .RN(pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_v[2]) );
  DFFR_X1 pe_1_1_1_int_q_reg_v_reg_5__3_ ( .D(int_data_y_2__1__3_), .CK(
        pe_1_1_1_net6845), .RN(pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_1_1_int_q_reg_h_reg_0__0_ ( .D(int_data_x_1__2__0_), .SI(
        int_data_y_2__1__0_), .SE(pe_1_1_1_n65), .CK(pe_1_1_1_net6789), .RN(
        pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_1_1_int_q_reg_h_reg_0__1_ ( .D(int_data_x_1__2__1_), .SI(
        int_data_y_2__1__1_), .SE(pe_1_1_1_n65), .CK(pe_1_1_1_net6789), .RN(
        pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_1_1_int_q_reg_h_reg_0__2_ ( .D(int_data_x_1__2__2_), .SI(
        int_data_y_2__1__2_), .SE(pe_1_1_1_n65), .CK(pe_1_1_1_net6789), .RN(
        pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_1_1_int_q_reg_h_reg_0__3_ ( .D(int_data_x_1__2__3_), .SI(
        int_data_y_2__1__3_), .SE(pe_1_1_1_n65), .CK(pe_1_1_1_net6789), .RN(
        pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_1_1_int_q_reg_h_reg_1__0_ ( .D(int_data_x_1__2__0_), .SI(
        int_data_y_2__1__0_), .SE(pe_1_1_1_n65), .CK(pe_1_1_1_net6795), .RN(
        pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_1_1_int_q_reg_h_reg_1__1_ ( .D(int_data_x_1__2__1_), .SI(
        int_data_y_2__1__1_), .SE(pe_1_1_1_n65), .CK(pe_1_1_1_net6795), .RN(
        pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_1_1_int_q_reg_h_reg_1__2_ ( .D(int_data_x_1__2__2_), .SI(
        int_data_y_2__1__2_), .SE(pe_1_1_1_n65), .CK(pe_1_1_1_net6795), .RN(
        pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_1_1_int_q_reg_h_reg_1__3_ ( .D(int_data_x_1__2__3_), .SI(
        int_data_y_2__1__3_), .SE(pe_1_1_1_n65), .CK(pe_1_1_1_net6795), .RN(
        pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_1_1_int_q_reg_h_reg_2__0_ ( .D(int_data_x_1__2__0_), .SI(
        int_data_y_2__1__0_), .SE(pe_1_1_1_n65), .CK(pe_1_1_1_net6800), .RN(
        pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_1_1_int_q_reg_h_reg_2__1_ ( .D(int_data_x_1__2__1_), .SI(
        int_data_y_2__1__1_), .SE(pe_1_1_1_n65), .CK(pe_1_1_1_net6800), .RN(
        pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_1_1_int_q_reg_h_reg_2__2_ ( .D(int_data_x_1__2__2_), .SI(
        int_data_y_2__1__2_), .SE(pe_1_1_1_n65), .CK(pe_1_1_1_net6800), .RN(
        pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_1_1_int_q_reg_h_reg_2__3_ ( .D(int_data_x_1__2__3_), .SI(
        int_data_y_2__1__3_), .SE(pe_1_1_1_n65), .CK(pe_1_1_1_net6800), .RN(
        pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_1_1_int_q_reg_h_reg_3__0_ ( .D(int_data_x_1__2__0_), .SI(
        int_data_y_2__1__0_), .SE(pe_1_1_1_n65), .CK(pe_1_1_1_net6805), .RN(
        pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_1_1_int_q_reg_h_reg_3__1_ ( .D(int_data_x_1__2__1_), .SI(
        int_data_y_2__1__1_), .SE(pe_1_1_1_n65), .CK(pe_1_1_1_net6805), .RN(
        pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_1_1_int_q_reg_h_reg_3__2_ ( .D(int_data_x_1__2__2_), .SI(
        int_data_y_2__1__2_), .SE(pe_1_1_1_n65), .CK(pe_1_1_1_net6805), .RN(
        pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_1_1_int_q_reg_h_reg_3__3_ ( .D(int_data_x_1__2__3_), .SI(
        int_data_y_2__1__3_), .SE(pe_1_1_1_n65), .CK(pe_1_1_1_net6805), .RN(
        pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_1_1_int_q_reg_h_reg_4__0_ ( .D(int_data_x_1__2__0_), .SI(
        int_data_y_2__1__0_), .SE(pe_1_1_1_n66), .CK(pe_1_1_1_net6810), .RN(
        pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_1_1_int_q_reg_h_reg_4__1_ ( .D(int_data_x_1__2__1_), .SI(
        int_data_y_2__1__1_), .SE(pe_1_1_1_n66), .CK(pe_1_1_1_net6810), .RN(
        pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_1_1_int_q_reg_h_reg_4__2_ ( .D(int_data_x_1__2__2_), .SI(
        int_data_y_2__1__2_), .SE(pe_1_1_1_n66), .CK(pe_1_1_1_net6810), .RN(
        pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_1_1_int_q_reg_h_reg_4__3_ ( .D(int_data_x_1__2__3_), .SI(
        int_data_y_2__1__3_), .SE(pe_1_1_1_n66), .CK(pe_1_1_1_net6810), .RN(
        pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_1_1_int_q_reg_h_reg_5__0_ ( .D(int_data_x_1__2__0_), .SI(
        int_data_y_2__1__0_), .SE(pe_1_1_1_n66), .CK(pe_1_1_1_net6815), .RN(
        pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_1_1_int_q_reg_h_reg_5__1_ ( .D(int_data_x_1__2__1_), .SI(
        int_data_y_2__1__1_), .SE(pe_1_1_1_n66), .CK(pe_1_1_1_net6815), .RN(
        pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_1_1_int_q_reg_h_reg_5__2_ ( .D(int_data_x_1__2__2_), .SI(
        int_data_y_2__1__2_), .SE(pe_1_1_1_n66), .CK(pe_1_1_1_net6815), .RN(
        pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_1_1_int_q_reg_h_reg_5__3_ ( .D(int_data_x_1__2__3_), .SI(
        int_data_y_2__1__3_), .SE(pe_1_1_1_n66), .CK(pe_1_1_1_net6815), .RN(
        pe_1_1_1_n72), .Q(pe_1_1_1_int_q_reg_h[3]) );
  FA_X1 pe_1_1_1_sub_81_U2_7 ( .A(int_data_res_1__1__7_), .B(pe_1_1_1_n76), 
        .CI(pe_1_1_1_sub_81_carry[7]), .S(pe_1_1_1_N77) );
  FA_X1 pe_1_1_1_sub_81_U2_6 ( .A(int_data_res_1__1__6_), .B(pe_1_1_1_n76), 
        .CI(pe_1_1_1_sub_81_carry[6]), .CO(pe_1_1_1_sub_81_carry[7]), .S(
        pe_1_1_1_N76) );
  FA_X1 pe_1_1_1_sub_81_U2_5 ( .A(int_data_res_1__1__5_), .B(pe_1_1_1_n76), 
        .CI(pe_1_1_1_sub_81_carry[5]), .CO(pe_1_1_1_sub_81_carry[6]), .S(
        pe_1_1_1_N75) );
  FA_X1 pe_1_1_1_sub_81_U2_4 ( .A(int_data_res_1__1__4_), .B(pe_1_1_1_n76), 
        .CI(pe_1_1_1_sub_81_carry[4]), .CO(pe_1_1_1_sub_81_carry[5]), .S(
        pe_1_1_1_N74) );
  FA_X1 pe_1_1_1_sub_81_U2_3 ( .A(int_data_res_1__1__3_), .B(pe_1_1_1_n76), 
        .CI(pe_1_1_1_sub_81_carry[3]), .CO(pe_1_1_1_sub_81_carry[4]), .S(
        pe_1_1_1_N73) );
  FA_X1 pe_1_1_1_sub_81_U2_2 ( .A(int_data_res_1__1__2_), .B(pe_1_1_1_n75), 
        .CI(pe_1_1_1_sub_81_carry[2]), .CO(pe_1_1_1_sub_81_carry[3]), .S(
        pe_1_1_1_N72) );
  FA_X1 pe_1_1_1_sub_81_U2_1 ( .A(int_data_res_1__1__1_), .B(pe_1_1_1_n74), 
        .CI(pe_1_1_1_sub_81_carry[1]), .CO(pe_1_1_1_sub_81_carry[2]), .S(
        pe_1_1_1_N71) );
  FA_X1 pe_1_1_1_add_83_U1_7 ( .A(int_data_res_1__1__7_), .B(
        pe_1_1_1_int_data_3_), .CI(pe_1_1_1_add_83_carry[7]), .S(pe_1_1_1_N85)
         );
  FA_X1 pe_1_1_1_add_83_U1_6 ( .A(int_data_res_1__1__6_), .B(
        pe_1_1_1_int_data_3_), .CI(pe_1_1_1_add_83_carry[6]), .CO(
        pe_1_1_1_add_83_carry[7]), .S(pe_1_1_1_N84) );
  FA_X1 pe_1_1_1_add_83_U1_5 ( .A(int_data_res_1__1__5_), .B(
        pe_1_1_1_int_data_3_), .CI(pe_1_1_1_add_83_carry[5]), .CO(
        pe_1_1_1_add_83_carry[6]), .S(pe_1_1_1_N83) );
  FA_X1 pe_1_1_1_add_83_U1_4 ( .A(int_data_res_1__1__4_), .B(
        pe_1_1_1_int_data_3_), .CI(pe_1_1_1_add_83_carry[4]), .CO(
        pe_1_1_1_add_83_carry[5]), .S(pe_1_1_1_N82) );
  FA_X1 pe_1_1_1_add_83_U1_3 ( .A(int_data_res_1__1__3_), .B(
        pe_1_1_1_int_data_3_), .CI(pe_1_1_1_add_83_carry[3]), .CO(
        pe_1_1_1_add_83_carry[4]), .S(pe_1_1_1_N81) );
  FA_X1 pe_1_1_1_add_83_U1_2 ( .A(int_data_res_1__1__2_), .B(
        pe_1_1_1_int_data_2_), .CI(pe_1_1_1_add_83_carry[2]), .CO(
        pe_1_1_1_add_83_carry[3]), .S(pe_1_1_1_N80) );
  FA_X1 pe_1_1_1_add_83_U1_1 ( .A(int_data_res_1__1__1_), .B(
        pe_1_1_1_int_data_1_), .CI(pe_1_1_1_n2), .CO(pe_1_1_1_add_83_carry[2]), 
        .S(pe_1_1_1_N79) );
  NAND3_X1 pe_1_1_1_U56 ( .A1(pe_1_1_1_n60), .A2(pe_1_1_1_n43), .A3(
        pe_1_1_1_n62), .ZN(pe_1_1_1_n40) );
  NAND3_X1 pe_1_1_1_U55 ( .A1(pe_1_1_1_n43), .A2(pe_1_1_1_n61), .A3(
        pe_1_1_1_n62), .ZN(pe_1_1_1_n39) );
  NAND3_X1 pe_1_1_1_U54 ( .A1(pe_1_1_1_n43), .A2(pe_1_1_1_n63), .A3(
        pe_1_1_1_n60), .ZN(pe_1_1_1_n38) );
  NAND3_X1 pe_1_1_1_U53 ( .A1(pe_1_1_1_n61), .A2(pe_1_1_1_n63), .A3(
        pe_1_1_1_n43), .ZN(pe_1_1_1_n37) );
  DFFR_X1 pe_1_1_1_int_q_acc_reg_6_ ( .D(pe_1_1_1_n78), .CK(pe_1_1_1_net6850), 
        .RN(pe_1_1_1_n71), .Q(int_data_res_1__1__6_) );
  DFFR_X1 pe_1_1_1_int_q_acc_reg_5_ ( .D(pe_1_1_1_n79), .CK(pe_1_1_1_net6850), 
        .RN(pe_1_1_1_n71), .Q(int_data_res_1__1__5_) );
  DFFR_X1 pe_1_1_1_int_q_acc_reg_4_ ( .D(pe_1_1_1_n80), .CK(pe_1_1_1_net6850), 
        .RN(pe_1_1_1_n71), .Q(int_data_res_1__1__4_) );
  DFFR_X1 pe_1_1_1_int_q_acc_reg_3_ ( .D(pe_1_1_1_n81), .CK(pe_1_1_1_net6850), 
        .RN(pe_1_1_1_n71), .Q(int_data_res_1__1__3_) );
  DFFR_X1 pe_1_1_1_int_q_acc_reg_2_ ( .D(pe_1_1_1_n82), .CK(pe_1_1_1_net6850), 
        .RN(pe_1_1_1_n71), .Q(int_data_res_1__1__2_) );
  DFFR_X1 pe_1_1_1_int_q_acc_reg_1_ ( .D(pe_1_1_1_n83), .CK(pe_1_1_1_net6850), 
        .RN(pe_1_1_1_n71), .Q(int_data_res_1__1__1_) );
  DFFR_X1 pe_1_1_1_int_q_acc_reg_7_ ( .D(pe_1_1_1_n77), .CK(pe_1_1_1_net6850), 
        .RN(pe_1_1_1_n71), .Q(int_data_res_1__1__7_) );
  CLKGATETST_X1 pe_1_1_1_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_1_1_n88), .SE(1'b0), .GCK(pe_1_1_1_net6789) );
  CLKGATETST_X1 pe_1_1_1_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_1_1_n87), .SE(1'b0), .GCK(pe_1_1_1_net6795) );
  CLKGATETST_X1 pe_1_1_1_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_1_1_n86), .SE(1'b0), .GCK(pe_1_1_1_net6800) );
  CLKGATETST_X1 pe_1_1_1_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_1_1_n85), .SE(1'b0), .GCK(pe_1_1_1_net6805) );
  CLKGATETST_X1 pe_1_1_1_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_1_1_n90), .SE(1'b0), .GCK(pe_1_1_1_net6810) );
  CLKGATETST_X1 pe_1_1_1_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_1_1_n89), .SE(1'b0), .GCK(pe_1_1_1_net6815) );
  CLKGATETST_X1 pe_1_1_1_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_1_1_N64), .SE(1'b0), .GCK(pe_1_1_1_net6820) );
  CLKGATETST_X1 pe_1_1_1_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_1_1_N63), .SE(1'b0), .GCK(pe_1_1_1_net6825) );
  CLKGATETST_X1 pe_1_1_1_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_1_1_N62), .SE(1'b0), .GCK(pe_1_1_1_net6830) );
  CLKGATETST_X1 pe_1_1_1_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_1_1_N61), .SE(1'b0), .GCK(pe_1_1_1_net6835) );
  CLKGATETST_X1 pe_1_1_1_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_1_1_N60), .SE(1'b0), .GCK(pe_1_1_1_net6840) );
  CLKGATETST_X1 pe_1_1_1_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_1_1_N59), .SE(1'b0), .GCK(pe_1_1_1_net6845) );
  CLKGATETST_X1 pe_1_1_1_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_1_1_N90), .SE(1'b0), .GCK(pe_1_1_1_net6850) );
  CLKBUF_X1 pe_1_1_2_U112 ( .A(pe_1_1_2_n72), .Z(pe_1_1_2_n71) );
  INV_X1 pe_1_1_2_U111 ( .A(n73), .ZN(pe_1_1_2_n70) );
  INV_X1 pe_1_1_2_U110 ( .A(n65), .ZN(pe_1_1_2_n69) );
  INV_X1 pe_1_1_2_U109 ( .A(n65), .ZN(pe_1_1_2_n68) );
  INV_X1 pe_1_1_2_U108 ( .A(n65), .ZN(pe_1_1_2_n67) );
  INV_X1 pe_1_1_2_U107 ( .A(pe_1_1_2_n69), .ZN(pe_1_1_2_n66) );
  INV_X1 pe_1_1_2_U106 ( .A(pe_1_1_2_n63), .ZN(pe_1_1_2_n62) );
  INV_X1 pe_1_1_2_U105 ( .A(pe_1_1_2_n61), .ZN(pe_1_1_2_n60) );
  INV_X1 pe_1_1_2_U104 ( .A(n25), .ZN(pe_1_1_2_n59) );
  INV_X1 pe_1_1_2_U103 ( .A(pe_1_1_2_n59), .ZN(pe_1_1_2_n58) );
  INV_X1 pe_1_1_2_U102 ( .A(n17), .ZN(pe_1_1_2_n57) );
  MUX2_X1 pe_1_1_2_U101 ( .A(pe_1_1_2_n54), .B(pe_1_1_2_n51), .S(n45), .Z(
        int_data_x_1__2__3_) );
  MUX2_X1 pe_1_1_2_U100 ( .A(pe_1_1_2_n53), .B(pe_1_1_2_n52), .S(pe_1_1_2_n62), 
        .Z(pe_1_1_2_n54) );
  MUX2_X1 pe_1_1_2_U99 ( .A(pe_1_1_2_int_q_reg_h[23]), .B(
        pe_1_1_2_int_q_reg_h[19]), .S(pe_1_1_2_n56), .Z(pe_1_1_2_n53) );
  MUX2_X1 pe_1_1_2_U98 ( .A(pe_1_1_2_int_q_reg_h[15]), .B(
        pe_1_1_2_int_q_reg_h[11]), .S(pe_1_1_2_n56), .Z(pe_1_1_2_n52) );
  MUX2_X1 pe_1_1_2_U97 ( .A(pe_1_1_2_int_q_reg_h[7]), .B(
        pe_1_1_2_int_q_reg_h[3]), .S(pe_1_1_2_n56), .Z(pe_1_1_2_n51) );
  MUX2_X1 pe_1_1_2_U96 ( .A(pe_1_1_2_n50), .B(pe_1_1_2_n47), .S(n45), .Z(
        int_data_x_1__2__2_) );
  MUX2_X1 pe_1_1_2_U95 ( .A(pe_1_1_2_n49), .B(pe_1_1_2_n48), .S(pe_1_1_2_n62), 
        .Z(pe_1_1_2_n50) );
  MUX2_X1 pe_1_1_2_U94 ( .A(pe_1_1_2_int_q_reg_h[22]), .B(
        pe_1_1_2_int_q_reg_h[18]), .S(pe_1_1_2_n56), .Z(pe_1_1_2_n49) );
  MUX2_X1 pe_1_1_2_U93 ( .A(pe_1_1_2_int_q_reg_h[14]), .B(
        pe_1_1_2_int_q_reg_h[10]), .S(pe_1_1_2_n56), .Z(pe_1_1_2_n48) );
  MUX2_X1 pe_1_1_2_U92 ( .A(pe_1_1_2_int_q_reg_h[6]), .B(
        pe_1_1_2_int_q_reg_h[2]), .S(pe_1_1_2_n56), .Z(pe_1_1_2_n47) );
  MUX2_X1 pe_1_1_2_U91 ( .A(pe_1_1_2_n46), .B(pe_1_1_2_n24), .S(n45), .Z(
        int_data_x_1__2__1_) );
  MUX2_X1 pe_1_1_2_U90 ( .A(pe_1_1_2_n45), .B(pe_1_1_2_n25), .S(pe_1_1_2_n62), 
        .Z(pe_1_1_2_n46) );
  MUX2_X1 pe_1_1_2_U89 ( .A(pe_1_1_2_int_q_reg_h[21]), .B(
        pe_1_1_2_int_q_reg_h[17]), .S(pe_1_1_2_n56), .Z(pe_1_1_2_n45) );
  MUX2_X1 pe_1_1_2_U88 ( .A(pe_1_1_2_int_q_reg_h[13]), .B(
        pe_1_1_2_int_q_reg_h[9]), .S(pe_1_1_2_n56), .Z(pe_1_1_2_n25) );
  MUX2_X1 pe_1_1_2_U87 ( .A(pe_1_1_2_int_q_reg_h[5]), .B(
        pe_1_1_2_int_q_reg_h[1]), .S(pe_1_1_2_n56), .Z(pe_1_1_2_n24) );
  MUX2_X1 pe_1_1_2_U86 ( .A(pe_1_1_2_n23), .B(pe_1_1_2_n20), .S(n45), .Z(
        int_data_x_1__2__0_) );
  MUX2_X1 pe_1_1_2_U85 ( .A(pe_1_1_2_n22), .B(pe_1_1_2_n21), .S(pe_1_1_2_n62), 
        .Z(pe_1_1_2_n23) );
  MUX2_X1 pe_1_1_2_U84 ( .A(pe_1_1_2_int_q_reg_h[20]), .B(
        pe_1_1_2_int_q_reg_h[16]), .S(pe_1_1_2_n56), .Z(pe_1_1_2_n22) );
  MUX2_X1 pe_1_1_2_U83 ( .A(pe_1_1_2_int_q_reg_h[12]), .B(
        pe_1_1_2_int_q_reg_h[8]), .S(pe_1_1_2_n56), .Z(pe_1_1_2_n21) );
  MUX2_X1 pe_1_1_2_U82 ( .A(pe_1_1_2_int_q_reg_h[4]), .B(
        pe_1_1_2_int_q_reg_h[0]), .S(pe_1_1_2_n56), .Z(pe_1_1_2_n20) );
  MUX2_X1 pe_1_1_2_U81 ( .A(pe_1_1_2_n19), .B(pe_1_1_2_n16), .S(n45), .Z(
        int_data_y_1__2__3_) );
  MUX2_X1 pe_1_1_2_U80 ( .A(pe_1_1_2_n18), .B(pe_1_1_2_n17), .S(pe_1_1_2_n62), 
        .Z(pe_1_1_2_n19) );
  MUX2_X1 pe_1_1_2_U79 ( .A(pe_1_1_2_int_q_reg_v[23]), .B(
        pe_1_1_2_int_q_reg_v[19]), .S(pe_1_1_2_n55), .Z(pe_1_1_2_n18) );
  MUX2_X1 pe_1_1_2_U78 ( .A(pe_1_1_2_int_q_reg_v[15]), .B(
        pe_1_1_2_int_q_reg_v[11]), .S(pe_1_1_2_n55), .Z(pe_1_1_2_n17) );
  MUX2_X1 pe_1_1_2_U77 ( .A(pe_1_1_2_int_q_reg_v[7]), .B(
        pe_1_1_2_int_q_reg_v[3]), .S(pe_1_1_2_n55), .Z(pe_1_1_2_n16) );
  MUX2_X1 pe_1_1_2_U76 ( .A(pe_1_1_2_n15), .B(pe_1_1_2_n12), .S(n45), .Z(
        int_data_y_1__2__2_) );
  MUX2_X1 pe_1_1_2_U75 ( .A(pe_1_1_2_n14), .B(pe_1_1_2_n13), .S(pe_1_1_2_n62), 
        .Z(pe_1_1_2_n15) );
  MUX2_X1 pe_1_1_2_U74 ( .A(pe_1_1_2_int_q_reg_v[22]), .B(
        pe_1_1_2_int_q_reg_v[18]), .S(pe_1_1_2_n55), .Z(pe_1_1_2_n14) );
  MUX2_X1 pe_1_1_2_U73 ( .A(pe_1_1_2_int_q_reg_v[14]), .B(
        pe_1_1_2_int_q_reg_v[10]), .S(pe_1_1_2_n55), .Z(pe_1_1_2_n13) );
  MUX2_X1 pe_1_1_2_U72 ( .A(pe_1_1_2_int_q_reg_v[6]), .B(
        pe_1_1_2_int_q_reg_v[2]), .S(pe_1_1_2_n55), .Z(pe_1_1_2_n12) );
  MUX2_X1 pe_1_1_2_U71 ( .A(pe_1_1_2_n11), .B(pe_1_1_2_n8), .S(n45), .Z(
        int_data_y_1__2__1_) );
  MUX2_X1 pe_1_1_2_U70 ( .A(pe_1_1_2_n10), .B(pe_1_1_2_n9), .S(pe_1_1_2_n62), 
        .Z(pe_1_1_2_n11) );
  MUX2_X1 pe_1_1_2_U69 ( .A(pe_1_1_2_int_q_reg_v[21]), .B(
        pe_1_1_2_int_q_reg_v[17]), .S(pe_1_1_2_n55), .Z(pe_1_1_2_n10) );
  MUX2_X1 pe_1_1_2_U68 ( .A(pe_1_1_2_int_q_reg_v[13]), .B(
        pe_1_1_2_int_q_reg_v[9]), .S(pe_1_1_2_n55), .Z(pe_1_1_2_n9) );
  MUX2_X1 pe_1_1_2_U67 ( .A(pe_1_1_2_int_q_reg_v[5]), .B(
        pe_1_1_2_int_q_reg_v[1]), .S(pe_1_1_2_n55), .Z(pe_1_1_2_n8) );
  MUX2_X1 pe_1_1_2_U66 ( .A(pe_1_1_2_n7), .B(pe_1_1_2_n4), .S(n45), .Z(
        int_data_y_1__2__0_) );
  MUX2_X1 pe_1_1_2_U65 ( .A(pe_1_1_2_n6), .B(pe_1_1_2_n5), .S(pe_1_1_2_n62), 
        .Z(pe_1_1_2_n7) );
  MUX2_X1 pe_1_1_2_U64 ( .A(pe_1_1_2_int_q_reg_v[20]), .B(
        pe_1_1_2_int_q_reg_v[16]), .S(pe_1_1_2_n55), .Z(pe_1_1_2_n6) );
  MUX2_X1 pe_1_1_2_U63 ( .A(pe_1_1_2_int_q_reg_v[12]), .B(
        pe_1_1_2_int_q_reg_v[8]), .S(pe_1_1_2_n55), .Z(pe_1_1_2_n5) );
  MUX2_X1 pe_1_1_2_U62 ( .A(pe_1_1_2_int_q_reg_v[4]), .B(
        pe_1_1_2_int_q_reg_v[0]), .S(pe_1_1_2_n55), .Z(pe_1_1_2_n4) );
  AOI222_X1 pe_1_1_2_U61 ( .A1(int_data_res_2__2__2_), .A2(pe_1_1_2_n64), .B1(
        pe_1_1_2_N80), .B2(pe_1_1_2_n27), .C1(pe_1_1_2_N72), .C2(pe_1_1_2_n28), 
        .ZN(pe_1_1_2_n33) );
  INV_X1 pe_1_1_2_U60 ( .A(pe_1_1_2_n33), .ZN(pe_1_1_2_n82) );
  AOI222_X1 pe_1_1_2_U59 ( .A1(int_data_res_2__2__6_), .A2(pe_1_1_2_n64), .B1(
        pe_1_1_2_N84), .B2(pe_1_1_2_n27), .C1(pe_1_1_2_N76), .C2(pe_1_1_2_n28), 
        .ZN(pe_1_1_2_n29) );
  INV_X1 pe_1_1_2_U58 ( .A(pe_1_1_2_n29), .ZN(pe_1_1_2_n78) );
  XNOR2_X1 pe_1_1_2_U57 ( .A(pe_1_1_2_n73), .B(int_data_res_1__2__0_), .ZN(
        pe_1_1_2_N70) );
  AOI222_X1 pe_1_1_2_U52 ( .A1(int_data_res_2__2__0_), .A2(pe_1_1_2_n64), .B1(
        pe_1_1_2_n1), .B2(pe_1_1_2_n27), .C1(pe_1_1_2_N70), .C2(pe_1_1_2_n28), 
        .ZN(pe_1_1_2_n35) );
  INV_X1 pe_1_1_2_U51 ( .A(pe_1_1_2_n35), .ZN(pe_1_1_2_n84) );
  AOI222_X1 pe_1_1_2_U50 ( .A1(int_data_res_2__2__1_), .A2(pe_1_1_2_n64), .B1(
        pe_1_1_2_N79), .B2(pe_1_1_2_n27), .C1(pe_1_1_2_N71), .C2(pe_1_1_2_n28), 
        .ZN(pe_1_1_2_n34) );
  INV_X1 pe_1_1_2_U49 ( .A(pe_1_1_2_n34), .ZN(pe_1_1_2_n83) );
  AOI222_X1 pe_1_1_2_U48 ( .A1(int_data_res_2__2__3_), .A2(pe_1_1_2_n64), .B1(
        pe_1_1_2_N81), .B2(pe_1_1_2_n27), .C1(pe_1_1_2_N73), .C2(pe_1_1_2_n28), 
        .ZN(pe_1_1_2_n32) );
  INV_X1 pe_1_1_2_U47 ( .A(pe_1_1_2_n32), .ZN(pe_1_1_2_n81) );
  AOI222_X1 pe_1_1_2_U46 ( .A1(int_data_res_2__2__4_), .A2(pe_1_1_2_n64), .B1(
        pe_1_1_2_N82), .B2(pe_1_1_2_n27), .C1(pe_1_1_2_N74), .C2(pe_1_1_2_n28), 
        .ZN(pe_1_1_2_n31) );
  INV_X1 pe_1_1_2_U45 ( .A(pe_1_1_2_n31), .ZN(pe_1_1_2_n80) );
  AOI222_X1 pe_1_1_2_U44 ( .A1(int_data_res_2__2__5_), .A2(pe_1_1_2_n64), .B1(
        pe_1_1_2_N83), .B2(pe_1_1_2_n27), .C1(pe_1_1_2_N75), .C2(pe_1_1_2_n28), 
        .ZN(pe_1_1_2_n30) );
  INV_X1 pe_1_1_2_U43 ( .A(pe_1_1_2_n30), .ZN(pe_1_1_2_n79) );
  NAND2_X1 pe_1_1_2_U42 ( .A1(pe_1_1_2_int_data_0_), .A2(pe_1_1_2_n3), .ZN(
        pe_1_1_2_sub_81_carry[1]) );
  INV_X1 pe_1_1_2_U41 ( .A(pe_1_1_2_int_data_1_), .ZN(pe_1_1_2_n74) );
  INV_X1 pe_1_1_2_U40 ( .A(pe_1_1_2_int_data_2_), .ZN(pe_1_1_2_n75) );
  AND2_X1 pe_1_1_2_U39 ( .A1(pe_1_1_2_int_data_0_), .A2(int_data_res_1__2__0_), 
        .ZN(pe_1_1_2_n2) );
  AOI222_X1 pe_1_1_2_U38 ( .A1(pe_1_1_2_n64), .A2(int_data_res_2__2__7_), .B1(
        pe_1_1_2_N85), .B2(pe_1_1_2_n27), .C1(pe_1_1_2_N77), .C2(pe_1_1_2_n28), 
        .ZN(pe_1_1_2_n26) );
  INV_X1 pe_1_1_2_U37 ( .A(pe_1_1_2_n26), .ZN(pe_1_1_2_n77) );
  NOR3_X1 pe_1_1_2_U36 ( .A1(pe_1_1_2_n59), .A2(pe_1_1_2_n65), .A3(int_ckg[53]), .ZN(pe_1_1_2_n36) );
  OR2_X1 pe_1_1_2_U35 ( .A1(pe_1_1_2_n36), .A2(pe_1_1_2_n64), .ZN(pe_1_1_2_N90) );
  INV_X1 pe_1_1_2_U34 ( .A(n37), .ZN(pe_1_1_2_n63) );
  AND2_X1 pe_1_1_2_U33 ( .A1(int_data_x_1__2__2_), .A2(pe_1_1_2_n58), .ZN(
        pe_1_1_2_int_data_2_) );
  AND2_X1 pe_1_1_2_U32 ( .A1(int_data_x_1__2__1_), .A2(pe_1_1_2_n58), .ZN(
        pe_1_1_2_int_data_1_) );
  AND2_X1 pe_1_1_2_U31 ( .A1(int_data_x_1__2__3_), .A2(pe_1_1_2_n58), .ZN(
        pe_1_1_2_int_data_3_) );
  BUF_X1 pe_1_1_2_U30 ( .A(n59), .Z(pe_1_1_2_n64) );
  INV_X1 pe_1_1_2_U29 ( .A(n31), .ZN(pe_1_1_2_n61) );
  AND2_X1 pe_1_1_2_U28 ( .A1(int_data_x_1__2__0_), .A2(pe_1_1_2_n58), .ZN(
        pe_1_1_2_int_data_0_) );
  NAND2_X1 pe_1_1_2_U27 ( .A1(pe_1_1_2_n44), .A2(pe_1_1_2_n61), .ZN(
        pe_1_1_2_n41) );
  AND3_X1 pe_1_1_2_U26 ( .A1(n73), .A2(pe_1_1_2_n63), .A3(n45), .ZN(
        pe_1_1_2_n44) );
  INV_X1 pe_1_1_2_U25 ( .A(pe_1_1_2_int_data_3_), .ZN(pe_1_1_2_n76) );
  NOR2_X1 pe_1_1_2_U24 ( .A1(pe_1_1_2_n70), .A2(n45), .ZN(pe_1_1_2_n43) );
  NOR2_X1 pe_1_1_2_U23 ( .A1(pe_1_1_2_n57), .A2(pe_1_1_2_n64), .ZN(
        pe_1_1_2_n28) );
  NOR2_X1 pe_1_1_2_U22 ( .A1(n17), .A2(pe_1_1_2_n64), .ZN(pe_1_1_2_n27) );
  INV_X1 pe_1_1_2_U21 ( .A(pe_1_1_2_int_data_0_), .ZN(pe_1_1_2_n73) );
  INV_X1 pe_1_1_2_U20 ( .A(pe_1_1_2_n41), .ZN(pe_1_1_2_n90) );
  INV_X1 pe_1_1_2_U19 ( .A(pe_1_1_2_n37), .ZN(pe_1_1_2_n88) );
  INV_X1 pe_1_1_2_U18 ( .A(pe_1_1_2_n38), .ZN(pe_1_1_2_n87) );
  INV_X1 pe_1_1_2_U17 ( .A(pe_1_1_2_n39), .ZN(pe_1_1_2_n86) );
  NOR2_X1 pe_1_1_2_U16 ( .A1(pe_1_1_2_n68), .A2(pe_1_1_2_n42), .ZN(
        pe_1_1_2_N59) );
  NOR2_X1 pe_1_1_2_U15 ( .A1(pe_1_1_2_n68), .A2(pe_1_1_2_n41), .ZN(
        pe_1_1_2_N60) );
  NOR2_X1 pe_1_1_2_U14 ( .A1(pe_1_1_2_n68), .A2(pe_1_1_2_n38), .ZN(
        pe_1_1_2_N63) );
  NOR2_X1 pe_1_1_2_U13 ( .A1(pe_1_1_2_n67), .A2(pe_1_1_2_n40), .ZN(
        pe_1_1_2_N61) );
  NOR2_X1 pe_1_1_2_U12 ( .A1(pe_1_1_2_n67), .A2(pe_1_1_2_n39), .ZN(
        pe_1_1_2_N62) );
  NOR2_X1 pe_1_1_2_U11 ( .A1(pe_1_1_2_n37), .A2(pe_1_1_2_n67), .ZN(
        pe_1_1_2_N64) );
  NAND2_X1 pe_1_1_2_U10 ( .A1(pe_1_1_2_n44), .A2(pe_1_1_2_n60), .ZN(
        pe_1_1_2_n42) );
  BUF_X1 pe_1_1_2_U9 ( .A(pe_1_1_2_n60), .Z(pe_1_1_2_n55) );
  INV_X1 pe_1_1_2_U8 ( .A(pe_1_1_2_n69), .ZN(pe_1_1_2_n65) );
  BUF_X1 pe_1_1_2_U7 ( .A(pe_1_1_2_n60), .Z(pe_1_1_2_n56) );
  INV_X1 pe_1_1_2_U6 ( .A(pe_1_1_2_n42), .ZN(pe_1_1_2_n89) );
  INV_X1 pe_1_1_2_U5 ( .A(pe_1_1_2_n40), .ZN(pe_1_1_2_n85) );
  INV_X2 pe_1_1_2_U4 ( .A(n81), .ZN(pe_1_1_2_n72) );
  XOR2_X1 pe_1_1_2_U3 ( .A(pe_1_1_2_int_data_0_), .B(int_data_res_1__2__0_), 
        .Z(pe_1_1_2_n1) );
  DFFR_X1 pe_1_1_2_int_q_acc_reg_0_ ( .D(pe_1_1_2_n84), .CK(pe_1_1_2_net6772), 
        .RN(pe_1_1_2_n72), .Q(int_data_res_1__2__0_), .QN(pe_1_1_2_n3) );
  DFFR_X1 pe_1_1_2_int_q_reg_v_reg_0__0_ ( .D(int_data_y_2__2__0_), .CK(
        pe_1_1_2_net6742), .RN(pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_v[20]) );
  DFFR_X1 pe_1_1_2_int_q_reg_v_reg_0__1_ ( .D(int_data_y_2__2__1_), .CK(
        pe_1_1_2_net6742), .RN(pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_v[21]) );
  DFFR_X1 pe_1_1_2_int_q_reg_v_reg_0__2_ ( .D(int_data_y_2__2__2_), .CK(
        pe_1_1_2_net6742), .RN(pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_v[22]) );
  DFFR_X1 pe_1_1_2_int_q_reg_v_reg_0__3_ ( .D(int_data_y_2__2__3_), .CK(
        pe_1_1_2_net6742), .RN(pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_v[23]) );
  DFFR_X1 pe_1_1_2_int_q_reg_v_reg_1__0_ ( .D(int_data_y_2__2__0_), .CK(
        pe_1_1_2_net6747), .RN(pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_v[16]) );
  DFFR_X1 pe_1_1_2_int_q_reg_v_reg_1__1_ ( .D(int_data_y_2__2__1_), .CK(
        pe_1_1_2_net6747), .RN(pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_v[17]) );
  DFFR_X1 pe_1_1_2_int_q_reg_v_reg_1__2_ ( .D(int_data_y_2__2__2_), .CK(
        pe_1_1_2_net6747), .RN(pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_v[18]) );
  DFFR_X1 pe_1_1_2_int_q_reg_v_reg_1__3_ ( .D(int_data_y_2__2__3_), .CK(
        pe_1_1_2_net6747), .RN(pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_v[19]) );
  DFFR_X1 pe_1_1_2_int_q_reg_v_reg_2__0_ ( .D(int_data_y_2__2__0_), .CK(
        pe_1_1_2_net6752), .RN(pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_v[12]) );
  DFFR_X1 pe_1_1_2_int_q_reg_v_reg_2__1_ ( .D(int_data_y_2__2__1_), .CK(
        pe_1_1_2_net6752), .RN(pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_v[13]) );
  DFFR_X1 pe_1_1_2_int_q_reg_v_reg_2__2_ ( .D(int_data_y_2__2__2_), .CK(
        pe_1_1_2_net6752), .RN(pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_v[14]) );
  DFFR_X1 pe_1_1_2_int_q_reg_v_reg_2__3_ ( .D(int_data_y_2__2__3_), .CK(
        pe_1_1_2_net6752), .RN(pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_v[15]) );
  DFFR_X1 pe_1_1_2_int_q_reg_v_reg_3__0_ ( .D(int_data_y_2__2__0_), .CK(
        pe_1_1_2_net6757), .RN(pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_v[8]) );
  DFFR_X1 pe_1_1_2_int_q_reg_v_reg_3__1_ ( .D(int_data_y_2__2__1_), .CK(
        pe_1_1_2_net6757), .RN(pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_v[9]) );
  DFFR_X1 pe_1_1_2_int_q_reg_v_reg_3__2_ ( .D(int_data_y_2__2__2_), .CK(
        pe_1_1_2_net6757), .RN(pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_v[10]) );
  DFFR_X1 pe_1_1_2_int_q_reg_v_reg_3__3_ ( .D(int_data_y_2__2__3_), .CK(
        pe_1_1_2_net6757), .RN(pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_v[11]) );
  DFFR_X1 pe_1_1_2_int_q_reg_v_reg_4__0_ ( .D(int_data_y_2__2__0_), .CK(
        pe_1_1_2_net6762), .RN(pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_v[4]) );
  DFFR_X1 pe_1_1_2_int_q_reg_v_reg_4__1_ ( .D(int_data_y_2__2__1_), .CK(
        pe_1_1_2_net6762), .RN(pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_v[5]) );
  DFFR_X1 pe_1_1_2_int_q_reg_v_reg_4__2_ ( .D(int_data_y_2__2__2_), .CK(
        pe_1_1_2_net6762), .RN(pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_v[6]) );
  DFFR_X1 pe_1_1_2_int_q_reg_v_reg_4__3_ ( .D(int_data_y_2__2__3_), .CK(
        pe_1_1_2_net6762), .RN(pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_v[7]) );
  DFFR_X1 pe_1_1_2_int_q_reg_v_reg_5__0_ ( .D(int_data_y_2__2__0_), .CK(
        pe_1_1_2_net6767), .RN(pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_v[0]) );
  DFFR_X1 pe_1_1_2_int_q_reg_v_reg_5__1_ ( .D(int_data_y_2__2__1_), .CK(
        pe_1_1_2_net6767), .RN(pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_v[1]) );
  DFFR_X1 pe_1_1_2_int_q_reg_v_reg_5__2_ ( .D(int_data_y_2__2__2_), .CK(
        pe_1_1_2_net6767), .RN(pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_v[2]) );
  DFFR_X1 pe_1_1_2_int_q_reg_v_reg_5__3_ ( .D(int_data_y_2__2__3_), .CK(
        pe_1_1_2_net6767), .RN(pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_1_2_int_q_reg_h_reg_0__0_ ( .D(int_data_x_1__3__0_), .SI(
        int_data_y_2__2__0_), .SE(pe_1_1_2_n65), .CK(pe_1_1_2_net6711), .RN(
        pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_1_2_int_q_reg_h_reg_0__1_ ( .D(int_data_x_1__3__1_), .SI(
        int_data_y_2__2__1_), .SE(pe_1_1_2_n65), .CK(pe_1_1_2_net6711), .RN(
        pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_1_2_int_q_reg_h_reg_0__2_ ( .D(int_data_x_1__3__2_), .SI(
        int_data_y_2__2__2_), .SE(pe_1_1_2_n65), .CK(pe_1_1_2_net6711), .RN(
        pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_1_2_int_q_reg_h_reg_0__3_ ( .D(int_data_x_1__3__3_), .SI(
        int_data_y_2__2__3_), .SE(pe_1_1_2_n65), .CK(pe_1_1_2_net6711), .RN(
        pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_1_2_int_q_reg_h_reg_1__0_ ( .D(int_data_x_1__3__0_), .SI(
        int_data_y_2__2__0_), .SE(pe_1_1_2_n65), .CK(pe_1_1_2_net6717), .RN(
        pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_1_2_int_q_reg_h_reg_1__1_ ( .D(int_data_x_1__3__1_), .SI(
        int_data_y_2__2__1_), .SE(pe_1_1_2_n65), .CK(pe_1_1_2_net6717), .RN(
        pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_1_2_int_q_reg_h_reg_1__2_ ( .D(int_data_x_1__3__2_), .SI(
        int_data_y_2__2__2_), .SE(pe_1_1_2_n65), .CK(pe_1_1_2_net6717), .RN(
        pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_1_2_int_q_reg_h_reg_1__3_ ( .D(int_data_x_1__3__3_), .SI(
        int_data_y_2__2__3_), .SE(pe_1_1_2_n65), .CK(pe_1_1_2_net6717), .RN(
        pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_1_2_int_q_reg_h_reg_2__0_ ( .D(int_data_x_1__3__0_), .SI(
        int_data_y_2__2__0_), .SE(pe_1_1_2_n65), .CK(pe_1_1_2_net6722), .RN(
        pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_1_2_int_q_reg_h_reg_2__1_ ( .D(int_data_x_1__3__1_), .SI(
        int_data_y_2__2__1_), .SE(pe_1_1_2_n65), .CK(pe_1_1_2_net6722), .RN(
        pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_1_2_int_q_reg_h_reg_2__2_ ( .D(int_data_x_1__3__2_), .SI(
        int_data_y_2__2__2_), .SE(pe_1_1_2_n65), .CK(pe_1_1_2_net6722), .RN(
        pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_1_2_int_q_reg_h_reg_2__3_ ( .D(int_data_x_1__3__3_), .SI(
        int_data_y_2__2__3_), .SE(pe_1_1_2_n65), .CK(pe_1_1_2_net6722), .RN(
        pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_1_2_int_q_reg_h_reg_3__0_ ( .D(int_data_x_1__3__0_), .SI(
        int_data_y_2__2__0_), .SE(pe_1_1_2_n65), .CK(pe_1_1_2_net6727), .RN(
        pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_1_2_int_q_reg_h_reg_3__1_ ( .D(int_data_x_1__3__1_), .SI(
        int_data_y_2__2__1_), .SE(pe_1_1_2_n65), .CK(pe_1_1_2_net6727), .RN(
        pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_1_2_int_q_reg_h_reg_3__2_ ( .D(int_data_x_1__3__2_), .SI(
        int_data_y_2__2__2_), .SE(pe_1_1_2_n65), .CK(pe_1_1_2_net6727), .RN(
        pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_1_2_int_q_reg_h_reg_3__3_ ( .D(int_data_x_1__3__3_), .SI(
        int_data_y_2__2__3_), .SE(pe_1_1_2_n65), .CK(pe_1_1_2_net6727), .RN(
        pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_1_2_int_q_reg_h_reg_4__0_ ( .D(int_data_x_1__3__0_), .SI(
        int_data_y_2__2__0_), .SE(pe_1_1_2_n66), .CK(pe_1_1_2_net6732), .RN(
        pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_1_2_int_q_reg_h_reg_4__1_ ( .D(int_data_x_1__3__1_), .SI(
        int_data_y_2__2__1_), .SE(pe_1_1_2_n66), .CK(pe_1_1_2_net6732), .RN(
        pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_1_2_int_q_reg_h_reg_4__2_ ( .D(int_data_x_1__3__2_), .SI(
        int_data_y_2__2__2_), .SE(pe_1_1_2_n66), .CK(pe_1_1_2_net6732), .RN(
        pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_1_2_int_q_reg_h_reg_4__3_ ( .D(int_data_x_1__3__3_), .SI(
        int_data_y_2__2__3_), .SE(pe_1_1_2_n66), .CK(pe_1_1_2_net6732), .RN(
        pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_1_2_int_q_reg_h_reg_5__0_ ( .D(int_data_x_1__3__0_), .SI(
        int_data_y_2__2__0_), .SE(pe_1_1_2_n66), .CK(pe_1_1_2_net6737), .RN(
        pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_1_2_int_q_reg_h_reg_5__1_ ( .D(int_data_x_1__3__1_), .SI(
        int_data_y_2__2__1_), .SE(pe_1_1_2_n66), .CK(pe_1_1_2_net6737), .RN(
        pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_1_2_int_q_reg_h_reg_5__2_ ( .D(int_data_x_1__3__2_), .SI(
        int_data_y_2__2__2_), .SE(pe_1_1_2_n66), .CK(pe_1_1_2_net6737), .RN(
        pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_1_2_int_q_reg_h_reg_5__3_ ( .D(int_data_x_1__3__3_), .SI(
        int_data_y_2__2__3_), .SE(pe_1_1_2_n66), .CK(pe_1_1_2_net6737), .RN(
        pe_1_1_2_n72), .Q(pe_1_1_2_int_q_reg_h[3]) );
  FA_X1 pe_1_1_2_sub_81_U2_7 ( .A(int_data_res_1__2__7_), .B(pe_1_1_2_n76), 
        .CI(pe_1_1_2_sub_81_carry[7]), .S(pe_1_1_2_N77) );
  FA_X1 pe_1_1_2_sub_81_U2_6 ( .A(int_data_res_1__2__6_), .B(pe_1_1_2_n76), 
        .CI(pe_1_1_2_sub_81_carry[6]), .CO(pe_1_1_2_sub_81_carry[7]), .S(
        pe_1_1_2_N76) );
  FA_X1 pe_1_1_2_sub_81_U2_5 ( .A(int_data_res_1__2__5_), .B(pe_1_1_2_n76), 
        .CI(pe_1_1_2_sub_81_carry[5]), .CO(pe_1_1_2_sub_81_carry[6]), .S(
        pe_1_1_2_N75) );
  FA_X1 pe_1_1_2_sub_81_U2_4 ( .A(int_data_res_1__2__4_), .B(pe_1_1_2_n76), 
        .CI(pe_1_1_2_sub_81_carry[4]), .CO(pe_1_1_2_sub_81_carry[5]), .S(
        pe_1_1_2_N74) );
  FA_X1 pe_1_1_2_sub_81_U2_3 ( .A(int_data_res_1__2__3_), .B(pe_1_1_2_n76), 
        .CI(pe_1_1_2_sub_81_carry[3]), .CO(pe_1_1_2_sub_81_carry[4]), .S(
        pe_1_1_2_N73) );
  FA_X1 pe_1_1_2_sub_81_U2_2 ( .A(int_data_res_1__2__2_), .B(pe_1_1_2_n75), 
        .CI(pe_1_1_2_sub_81_carry[2]), .CO(pe_1_1_2_sub_81_carry[3]), .S(
        pe_1_1_2_N72) );
  FA_X1 pe_1_1_2_sub_81_U2_1 ( .A(int_data_res_1__2__1_), .B(pe_1_1_2_n74), 
        .CI(pe_1_1_2_sub_81_carry[1]), .CO(pe_1_1_2_sub_81_carry[2]), .S(
        pe_1_1_2_N71) );
  FA_X1 pe_1_1_2_add_83_U1_7 ( .A(int_data_res_1__2__7_), .B(
        pe_1_1_2_int_data_3_), .CI(pe_1_1_2_add_83_carry[7]), .S(pe_1_1_2_N85)
         );
  FA_X1 pe_1_1_2_add_83_U1_6 ( .A(int_data_res_1__2__6_), .B(
        pe_1_1_2_int_data_3_), .CI(pe_1_1_2_add_83_carry[6]), .CO(
        pe_1_1_2_add_83_carry[7]), .S(pe_1_1_2_N84) );
  FA_X1 pe_1_1_2_add_83_U1_5 ( .A(int_data_res_1__2__5_), .B(
        pe_1_1_2_int_data_3_), .CI(pe_1_1_2_add_83_carry[5]), .CO(
        pe_1_1_2_add_83_carry[6]), .S(pe_1_1_2_N83) );
  FA_X1 pe_1_1_2_add_83_U1_4 ( .A(int_data_res_1__2__4_), .B(
        pe_1_1_2_int_data_3_), .CI(pe_1_1_2_add_83_carry[4]), .CO(
        pe_1_1_2_add_83_carry[5]), .S(pe_1_1_2_N82) );
  FA_X1 pe_1_1_2_add_83_U1_3 ( .A(int_data_res_1__2__3_), .B(
        pe_1_1_2_int_data_3_), .CI(pe_1_1_2_add_83_carry[3]), .CO(
        pe_1_1_2_add_83_carry[4]), .S(pe_1_1_2_N81) );
  FA_X1 pe_1_1_2_add_83_U1_2 ( .A(int_data_res_1__2__2_), .B(
        pe_1_1_2_int_data_2_), .CI(pe_1_1_2_add_83_carry[2]), .CO(
        pe_1_1_2_add_83_carry[3]), .S(pe_1_1_2_N80) );
  FA_X1 pe_1_1_2_add_83_U1_1 ( .A(int_data_res_1__2__1_), .B(
        pe_1_1_2_int_data_1_), .CI(pe_1_1_2_n2), .CO(pe_1_1_2_add_83_carry[2]), 
        .S(pe_1_1_2_N79) );
  NAND3_X1 pe_1_1_2_U56 ( .A1(pe_1_1_2_n60), .A2(pe_1_1_2_n43), .A3(
        pe_1_1_2_n62), .ZN(pe_1_1_2_n40) );
  NAND3_X1 pe_1_1_2_U55 ( .A1(pe_1_1_2_n43), .A2(pe_1_1_2_n61), .A3(
        pe_1_1_2_n62), .ZN(pe_1_1_2_n39) );
  NAND3_X1 pe_1_1_2_U54 ( .A1(pe_1_1_2_n43), .A2(pe_1_1_2_n63), .A3(
        pe_1_1_2_n60), .ZN(pe_1_1_2_n38) );
  NAND3_X1 pe_1_1_2_U53 ( .A1(pe_1_1_2_n61), .A2(pe_1_1_2_n63), .A3(
        pe_1_1_2_n43), .ZN(pe_1_1_2_n37) );
  DFFR_X1 pe_1_1_2_int_q_acc_reg_6_ ( .D(pe_1_1_2_n78), .CK(pe_1_1_2_net6772), 
        .RN(pe_1_1_2_n71), .Q(int_data_res_1__2__6_) );
  DFFR_X1 pe_1_1_2_int_q_acc_reg_5_ ( .D(pe_1_1_2_n79), .CK(pe_1_1_2_net6772), 
        .RN(pe_1_1_2_n71), .Q(int_data_res_1__2__5_) );
  DFFR_X1 pe_1_1_2_int_q_acc_reg_4_ ( .D(pe_1_1_2_n80), .CK(pe_1_1_2_net6772), 
        .RN(pe_1_1_2_n71), .Q(int_data_res_1__2__4_) );
  DFFR_X1 pe_1_1_2_int_q_acc_reg_3_ ( .D(pe_1_1_2_n81), .CK(pe_1_1_2_net6772), 
        .RN(pe_1_1_2_n71), .Q(int_data_res_1__2__3_) );
  DFFR_X1 pe_1_1_2_int_q_acc_reg_2_ ( .D(pe_1_1_2_n82), .CK(pe_1_1_2_net6772), 
        .RN(pe_1_1_2_n71), .Q(int_data_res_1__2__2_) );
  DFFR_X1 pe_1_1_2_int_q_acc_reg_1_ ( .D(pe_1_1_2_n83), .CK(pe_1_1_2_net6772), 
        .RN(pe_1_1_2_n71), .Q(int_data_res_1__2__1_) );
  DFFR_X1 pe_1_1_2_int_q_acc_reg_7_ ( .D(pe_1_1_2_n77), .CK(pe_1_1_2_net6772), 
        .RN(pe_1_1_2_n71), .Q(int_data_res_1__2__7_) );
  CLKGATETST_X1 pe_1_1_2_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_1_2_n88), .SE(1'b0), .GCK(pe_1_1_2_net6711) );
  CLKGATETST_X1 pe_1_1_2_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_1_2_n87), .SE(1'b0), .GCK(pe_1_1_2_net6717) );
  CLKGATETST_X1 pe_1_1_2_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_1_2_n86), .SE(1'b0), .GCK(pe_1_1_2_net6722) );
  CLKGATETST_X1 pe_1_1_2_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_1_2_n85), .SE(1'b0), .GCK(pe_1_1_2_net6727) );
  CLKGATETST_X1 pe_1_1_2_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_1_2_n90), .SE(1'b0), .GCK(pe_1_1_2_net6732) );
  CLKGATETST_X1 pe_1_1_2_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_1_2_n89), .SE(1'b0), .GCK(pe_1_1_2_net6737) );
  CLKGATETST_X1 pe_1_1_2_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_1_2_N64), .SE(1'b0), .GCK(pe_1_1_2_net6742) );
  CLKGATETST_X1 pe_1_1_2_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_1_2_N63), .SE(1'b0), .GCK(pe_1_1_2_net6747) );
  CLKGATETST_X1 pe_1_1_2_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_1_2_N62), .SE(1'b0), .GCK(pe_1_1_2_net6752) );
  CLKGATETST_X1 pe_1_1_2_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_1_2_N61), .SE(1'b0), .GCK(pe_1_1_2_net6757) );
  CLKGATETST_X1 pe_1_1_2_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_1_2_N60), .SE(1'b0), .GCK(pe_1_1_2_net6762) );
  CLKGATETST_X1 pe_1_1_2_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_1_2_N59), .SE(1'b0), .GCK(pe_1_1_2_net6767) );
  CLKGATETST_X1 pe_1_1_2_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_1_2_N90), .SE(1'b0), .GCK(pe_1_1_2_net6772) );
  CLKBUF_X1 pe_1_1_3_U112 ( .A(pe_1_1_3_n72), .Z(pe_1_1_3_n71) );
  INV_X1 pe_1_1_3_U111 ( .A(n73), .ZN(pe_1_1_3_n70) );
  INV_X1 pe_1_1_3_U110 ( .A(n65), .ZN(pe_1_1_3_n69) );
  INV_X1 pe_1_1_3_U109 ( .A(n65), .ZN(pe_1_1_3_n68) );
  INV_X1 pe_1_1_3_U108 ( .A(n65), .ZN(pe_1_1_3_n67) );
  INV_X1 pe_1_1_3_U107 ( .A(pe_1_1_3_n69), .ZN(pe_1_1_3_n66) );
  INV_X1 pe_1_1_3_U106 ( .A(pe_1_1_3_n63), .ZN(pe_1_1_3_n62) );
  INV_X1 pe_1_1_3_U105 ( .A(pe_1_1_3_n61), .ZN(pe_1_1_3_n60) );
  INV_X1 pe_1_1_3_U104 ( .A(n25), .ZN(pe_1_1_3_n59) );
  INV_X1 pe_1_1_3_U103 ( .A(pe_1_1_3_n59), .ZN(pe_1_1_3_n58) );
  INV_X1 pe_1_1_3_U102 ( .A(n17), .ZN(pe_1_1_3_n57) );
  MUX2_X1 pe_1_1_3_U101 ( .A(pe_1_1_3_n54), .B(pe_1_1_3_n51), .S(n45), .Z(
        int_data_x_1__3__3_) );
  MUX2_X1 pe_1_1_3_U100 ( .A(pe_1_1_3_n53), .B(pe_1_1_3_n52), .S(pe_1_1_3_n62), 
        .Z(pe_1_1_3_n54) );
  MUX2_X1 pe_1_1_3_U99 ( .A(pe_1_1_3_int_q_reg_h[23]), .B(
        pe_1_1_3_int_q_reg_h[19]), .S(pe_1_1_3_n56), .Z(pe_1_1_3_n53) );
  MUX2_X1 pe_1_1_3_U98 ( .A(pe_1_1_3_int_q_reg_h[15]), .B(
        pe_1_1_3_int_q_reg_h[11]), .S(pe_1_1_3_n56), .Z(pe_1_1_3_n52) );
  MUX2_X1 pe_1_1_3_U97 ( .A(pe_1_1_3_int_q_reg_h[7]), .B(
        pe_1_1_3_int_q_reg_h[3]), .S(pe_1_1_3_n56), .Z(pe_1_1_3_n51) );
  MUX2_X1 pe_1_1_3_U96 ( .A(pe_1_1_3_n50), .B(pe_1_1_3_n47), .S(n45), .Z(
        int_data_x_1__3__2_) );
  MUX2_X1 pe_1_1_3_U95 ( .A(pe_1_1_3_n49), .B(pe_1_1_3_n48), .S(pe_1_1_3_n62), 
        .Z(pe_1_1_3_n50) );
  MUX2_X1 pe_1_1_3_U94 ( .A(pe_1_1_3_int_q_reg_h[22]), .B(
        pe_1_1_3_int_q_reg_h[18]), .S(pe_1_1_3_n56), .Z(pe_1_1_3_n49) );
  MUX2_X1 pe_1_1_3_U93 ( .A(pe_1_1_3_int_q_reg_h[14]), .B(
        pe_1_1_3_int_q_reg_h[10]), .S(pe_1_1_3_n56), .Z(pe_1_1_3_n48) );
  MUX2_X1 pe_1_1_3_U92 ( .A(pe_1_1_3_int_q_reg_h[6]), .B(
        pe_1_1_3_int_q_reg_h[2]), .S(pe_1_1_3_n56), .Z(pe_1_1_3_n47) );
  MUX2_X1 pe_1_1_3_U91 ( .A(pe_1_1_3_n46), .B(pe_1_1_3_n24), .S(n45), .Z(
        int_data_x_1__3__1_) );
  MUX2_X1 pe_1_1_3_U90 ( .A(pe_1_1_3_n45), .B(pe_1_1_3_n25), .S(pe_1_1_3_n62), 
        .Z(pe_1_1_3_n46) );
  MUX2_X1 pe_1_1_3_U89 ( .A(pe_1_1_3_int_q_reg_h[21]), .B(
        pe_1_1_3_int_q_reg_h[17]), .S(pe_1_1_3_n56), .Z(pe_1_1_3_n45) );
  MUX2_X1 pe_1_1_3_U88 ( .A(pe_1_1_3_int_q_reg_h[13]), .B(
        pe_1_1_3_int_q_reg_h[9]), .S(pe_1_1_3_n56), .Z(pe_1_1_3_n25) );
  MUX2_X1 pe_1_1_3_U87 ( .A(pe_1_1_3_int_q_reg_h[5]), .B(
        pe_1_1_3_int_q_reg_h[1]), .S(pe_1_1_3_n56), .Z(pe_1_1_3_n24) );
  MUX2_X1 pe_1_1_3_U86 ( .A(pe_1_1_3_n23), .B(pe_1_1_3_n20), .S(n45), .Z(
        int_data_x_1__3__0_) );
  MUX2_X1 pe_1_1_3_U85 ( .A(pe_1_1_3_n22), .B(pe_1_1_3_n21), .S(pe_1_1_3_n62), 
        .Z(pe_1_1_3_n23) );
  MUX2_X1 pe_1_1_3_U84 ( .A(pe_1_1_3_int_q_reg_h[20]), .B(
        pe_1_1_3_int_q_reg_h[16]), .S(pe_1_1_3_n56), .Z(pe_1_1_3_n22) );
  MUX2_X1 pe_1_1_3_U83 ( .A(pe_1_1_3_int_q_reg_h[12]), .B(
        pe_1_1_3_int_q_reg_h[8]), .S(pe_1_1_3_n56), .Z(pe_1_1_3_n21) );
  MUX2_X1 pe_1_1_3_U82 ( .A(pe_1_1_3_int_q_reg_h[4]), .B(
        pe_1_1_3_int_q_reg_h[0]), .S(pe_1_1_3_n56), .Z(pe_1_1_3_n20) );
  MUX2_X1 pe_1_1_3_U81 ( .A(pe_1_1_3_n19), .B(pe_1_1_3_n16), .S(n45), .Z(
        int_data_y_1__3__3_) );
  MUX2_X1 pe_1_1_3_U80 ( .A(pe_1_1_3_n18), .B(pe_1_1_3_n17), .S(pe_1_1_3_n62), 
        .Z(pe_1_1_3_n19) );
  MUX2_X1 pe_1_1_3_U79 ( .A(pe_1_1_3_int_q_reg_v[23]), .B(
        pe_1_1_3_int_q_reg_v[19]), .S(pe_1_1_3_n55), .Z(pe_1_1_3_n18) );
  MUX2_X1 pe_1_1_3_U78 ( .A(pe_1_1_3_int_q_reg_v[15]), .B(
        pe_1_1_3_int_q_reg_v[11]), .S(pe_1_1_3_n55), .Z(pe_1_1_3_n17) );
  MUX2_X1 pe_1_1_3_U77 ( .A(pe_1_1_3_int_q_reg_v[7]), .B(
        pe_1_1_3_int_q_reg_v[3]), .S(pe_1_1_3_n55), .Z(pe_1_1_3_n16) );
  MUX2_X1 pe_1_1_3_U76 ( .A(pe_1_1_3_n15), .B(pe_1_1_3_n12), .S(n45), .Z(
        int_data_y_1__3__2_) );
  MUX2_X1 pe_1_1_3_U75 ( .A(pe_1_1_3_n14), .B(pe_1_1_3_n13), .S(pe_1_1_3_n62), 
        .Z(pe_1_1_3_n15) );
  MUX2_X1 pe_1_1_3_U74 ( .A(pe_1_1_3_int_q_reg_v[22]), .B(
        pe_1_1_3_int_q_reg_v[18]), .S(pe_1_1_3_n55), .Z(pe_1_1_3_n14) );
  MUX2_X1 pe_1_1_3_U73 ( .A(pe_1_1_3_int_q_reg_v[14]), .B(
        pe_1_1_3_int_q_reg_v[10]), .S(pe_1_1_3_n55), .Z(pe_1_1_3_n13) );
  MUX2_X1 pe_1_1_3_U72 ( .A(pe_1_1_3_int_q_reg_v[6]), .B(
        pe_1_1_3_int_q_reg_v[2]), .S(pe_1_1_3_n55), .Z(pe_1_1_3_n12) );
  MUX2_X1 pe_1_1_3_U71 ( .A(pe_1_1_3_n11), .B(pe_1_1_3_n8), .S(n45), .Z(
        int_data_y_1__3__1_) );
  MUX2_X1 pe_1_1_3_U70 ( .A(pe_1_1_3_n10), .B(pe_1_1_3_n9), .S(pe_1_1_3_n62), 
        .Z(pe_1_1_3_n11) );
  MUX2_X1 pe_1_1_3_U69 ( .A(pe_1_1_3_int_q_reg_v[21]), .B(
        pe_1_1_3_int_q_reg_v[17]), .S(pe_1_1_3_n55), .Z(pe_1_1_3_n10) );
  MUX2_X1 pe_1_1_3_U68 ( .A(pe_1_1_3_int_q_reg_v[13]), .B(
        pe_1_1_3_int_q_reg_v[9]), .S(pe_1_1_3_n55), .Z(pe_1_1_3_n9) );
  MUX2_X1 pe_1_1_3_U67 ( .A(pe_1_1_3_int_q_reg_v[5]), .B(
        pe_1_1_3_int_q_reg_v[1]), .S(pe_1_1_3_n55), .Z(pe_1_1_3_n8) );
  MUX2_X1 pe_1_1_3_U66 ( .A(pe_1_1_3_n7), .B(pe_1_1_3_n4), .S(n45), .Z(
        int_data_y_1__3__0_) );
  MUX2_X1 pe_1_1_3_U65 ( .A(pe_1_1_3_n6), .B(pe_1_1_3_n5), .S(pe_1_1_3_n62), 
        .Z(pe_1_1_3_n7) );
  MUX2_X1 pe_1_1_3_U64 ( .A(pe_1_1_3_int_q_reg_v[20]), .B(
        pe_1_1_3_int_q_reg_v[16]), .S(pe_1_1_3_n55), .Z(pe_1_1_3_n6) );
  MUX2_X1 pe_1_1_3_U63 ( .A(pe_1_1_3_int_q_reg_v[12]), .B(
        pe_1_1_3_int_q_reg_v[8]), .S(pe_1_1_3_n55), .Z(pe_1_1_3_n5) );
  MUX2_X1 pe_1_1_3_U62 ( .A(pe_1_1_3_int_q_reg_v[4]), .B(
        pe_1_1_3_int_q_reg_v[0]), .S(pe_1_1_3_n55), .Z(pe_1_1_3_n4) );
  AOI222_X1 pe_1_1_3_U61 ( .A1(int_data_res_2__3__2_), .A2(pe_1_1_3_n64), .B1(
        pe_1_1_3_N80), .B2(pe_1_1_3_n27), .C1(pe_1_1_3_N72), .C2(pe_1_1_3_n28), 
        .ZN(pe_1_1_3_n33) );
  INV_X1 pe_1_1_3_U60 ( .A(pe_1_1_3_n33), .ZN(pe_1_1_3_n82) );
  AOI222_X1 pe_1_1_3_U59 ( .A1(int_data_res_2__3__6_), .A2(pe_1_1_3_n64), .B1(
        pe_1_1_3_N84), .B2(pe_1_1_3_n27), .C1(pe_1_1_3_N76), .C2(pe_1_1_3_n28), 
        .ZN(pe_1_1_3_n29) );
  INV_X1 pe_1_1_3_U58 ( .A(pe_1_1_3_n29), .ZN(pe_1_1_3_n78) );
  XNOR2_X1 pe_1_1_3_U57 ( .A(pe_1_1_3_n73), .B(int_data_res_1__3__0_), .ZN(
        pe_1_1_3_N70) );
  AOI222_X1 pe_1_1_3_U52 ( .A1(int_data_res_2__3__0_), .A2(pe_1_1_3_n64), .B1(
        pe_1_1_3_n1), .B2(pe_1_1_3_n27), .C1(pe_1_1_3_N70), .C2(pe_1_1_3_n28), 
        .ZN(pe_1_1_3_n35) );
  INV_X1 pe_1_1_3_U51 ( .A(pe_1_1_3_n35), .ZN(pe_1_1_3_n84) );
  AOI222_X1 pe_1_1_3_U50 ( .A1(int_data_res_2__3__1_), .A2(pe_1_1_3_n64), .B1(
        pe_1_1_3_N79), .B2(pe_1_1_3_n27), .C1(pe_1_1_3_N71), .C2(pe_1_1_3_n28), 
        .ZN(pe_1_1_3_n34) );
  INV_X1 pe_1_1_3_U49 ( .A(pe_1_1_3_n34), .ZN(pe_1_1_3_n83) );
  AOI222_X1 pe_1_1_3_U48 ( .A1(int_data_res_2__3__3_), .A2(pe_1_1_3_n64), .B1(
        pe_1_1_3_N81), .B2(pe_1_1_3_n27), .C1(pe_1_1_3_N73), .C2(pe_1_1_3_n28), 
        .ZN(pe_1_1_3_n32) );
  INV_X1 pe_1_1_3_U47 ( .A(pe_1_1_3_n32), .ZN(pe_1_1_3_n81) );
  AOI222_X1 pe_1_1_3_U46 ( .A1(int_data_res_2__3__4_), .A2(pe_1_1_3_n64), .B1(
        pe_1_1_3_N82), .B2(pe_1_1_3_n27), .C1(pe_1_1_3_N74), .C2(pe_1_1_3_n28), 
        .ZN(pe_1_1_3_n31) );
  INV_X1 pe_1_1_3_U45 ( .A(pe_1_1_3_n31), .ZN(pe_1_1_3_n80) );
  AOI222_X1 pe_1_1_3_U44 ( .A1(int_data_res_2__3__5_), .A2(pe_1_1_3_n64), .B1(
        pe_1_1_3_N83), .B2(pe_1_1_3_n27), .C1(pe_1_1_3_N75), .C2(pe_1_1_3_n28), 
        .ZN(pe_1_1_3_n30) );
  INV_X1 pe_1_1_3_U43 ( .A(pe_1_1_3_n30), .ZN(pe_1_1_3_n79) );
  NAND2_X1 pe_1_1_3_U42 ( .A1(pe_1_1_3_int_data_0_), .A2(pe_1_1_3_n3), .ZN(
        pe_1_1_3_sub_81_carry[1]) );
  INV_X1 pe_1_1_3_U41 ( .A(pe_1_1_3_int_data_1_), .ZN(pe_1_1_3_n74) );
  INV_X1 pe_1_1_3_U40 ( .A(pe_1_1_3_int_data_2_), .ZN(pe_1_1_3_n75) );
  AND2_X1 pe_1_1_3_U39 ( .A1(pe_1_1_3_int_data_0_), .A2(int_data_res_1__3__0_), 
        .ZN(pe_1_1_3_n2) );
  AOI222_X1 pe_1_1_3_U38 ( .A1(pe_1_1_3_n64), .A2(int_data_res_2__3__7_), .B1(
        pe_1_1_3_N85), .B2(pe_1_1_3_n27), .C1(pe_1_1_3_N77), .C2(pe_1_1_3_n28), 
        .ZN(pe_1_1_3_n26) );
  INV_X1 pe_1_1_3_U37 ( .A(pe_1_1_3_n26), .ZN(pe_1_1_3_n77) );
  NOR3_X1 pe_1_1_3_U36 ( .A1(pe_1_1_3_n59), .A2(pe_1_1_3_n65), .A3(int_ckg[52]), .ZN(pe_1_1_3_n36) );
  OR2_X1 pe_1_1_3_U35 ( .A1(pe_1_1_3_n36), .A2(pe_1_1_3_n64), .ZN(pe_1_1_3_N90) );
  INV_X1 pe_1_1_3_U34 ( .A(n37), .ZN(pe_1_1_3_n63) );
  AND2_X1 pe_1_1_3_U33 ( .A1(int_data_x_1__3__2_), .A2(pe_1_1_3_n58), .ZN(
        pe_1_1_3_int_data_2_) );
  AND2_X1 pe_1_1_3_U32 ( .A1(int_data_x_1__3__1_), .A2(pe_1_1_3_n58), .ZN(
        pe_1_1_3_int_data_1_) );
  AND2_X1 pe_1_1_3_U31 ( .A1(int_data_x_1__3__3_), .A2(pe_1_1_3_n58), .ZN(
        pe_1_1_3_int_data_3_) );
  BUF_X1 pe_1_1_3_U30 ( .A(n59), .Z(pe_1_1_3_n64) );
  INV_X1 pe_1_1_3_U29 ( .A(n31), .ZN(pe_1_1_3_n61) );
  AND2_X1 pe_1_1_3_U28 ( .A1(int_data_x_1__3__0_), .A2(pe_1_1_3_n58), .ZN(
        pe_1_1_3_int_data_0_) );
  NAND2_X1 pe_1_1_3_U27 ( .A1(pe_1_1_3_n44), .A2(pe_1_1_3_n61), .ZN(
        pe_1_1_3_n41) );
  AND3_X1 pe_1_1_3_U26 ( .A1(n73), .A2(pe_1_1_3_n63), .A3(n45), .ZN(
        pe_1_1_3_n44) );
  INV_X1 pe_1_1_3_U25 ( .A(pe_1_1_3_int_data_3_), .ZN(pe_1_1_3_n76) );
  NOR2_X1 pe_1_1_3_U24 ( .A1(pe_1_1_3_n70), .A2(n45), .ZN(pe_1_1_3_n43) );
  NOR2_X1 pe_1_1_3_U23 ( .A1(pe_1_1_3_n57), .A2(pe_1_1_3_n64), .ZN(
        pe_1_1_3_n28) );
  NOR2_X1 pe_1_1_3_U22 ( .A1(n17), .A2(pe_1_1_3_n64), .ZN(pe_1_1_3_n27) );
  INV_X1 pe_1_1_3_U21 ( .A(pe_1_1_3_int_data_0_), .ZN(pe_1_1_3_n73) );
  INV_X1 pe_1_1_3_U20 ( .A(pe_1_1_3_n41), .ZN(pe_1_1_3_n90) );
  INV_X1 pe_1_1_3_U19 ( .A(pe_1_1_3_n37), .ZN(pe_1_1_3_n88) );
  INV_X1 pe_1_1_3_U18 ( .A(pe_1_1_3_n38), .ZN(pe_1_1_3_n87) );
  INV_X1 pe_1_1_3_U17 ( .A(pe_1_1_3_n39), .ZN(pe_1_1_3_n86) );
  NOR2_X1 pe_1_1_3_U16 ( .A1(pe_1_1_3_n68), .A2(pe_1_1_3_n42), .ZN(
        pe_1_1_3_N59) );
  NOR2_X1 pe_1_1_3_U15 ( .A1(pe_1_1_3_n68), .A2(pe_1_1_3_n41), .ZN(
        pe_1_1_3_N60) );
  NOR2_X1 pe_1_1_3_U14 ( .A1(pe_1_1_3_n68), .A2(pe_1_1_3_n38), .ZN(
        pe_1_1_3_N63) );
  NOR2_X1 pe_1_1_3_U13 ( .A1(pe_1_1_3_n67), .A2(pe_1_1_3_n40), .ZN(
        pe_1_1_3_N61) );
  NOR2_X1 pe_1_1_3_U12 ( .A1(pe_1_1_3_n67), .A2(pe_1_1_3_n39), .ZN(
        pe_1_1_3_N62) );
  NOR2_X1 pe_1_1_3_U11 ( .A1(pe_1_1_3_n37), .A2(pe_1_1_3_n67), .ZN(
        pe_1_1_3_N64) );
  NAND2_X1 pe_1_1_3_U10 ( .A1(pe_1_1_3_n44), .A2(pe_1_1_3_n60), .ZN(
        pe_1_1_3_n42) );
  BUF_X1 pe_1_1_3_U9 ( .A(pe_1_1_3_n60), .Z(pe_1_1_3_n55) );
  INV_X1 pe_1_1_3_U8 ( .A(pe_1_1_3_n69), .ZN(pe_1_1_3_n65) );
  BUF_X1 pe_1_1_3_U7 ( .A(pe_1_1_3_n60), .Z(pe_1_1_3_n56) );
  INV_X1 pe_1_1_3_U6 ( .A(pe_1_1_3_n42), .ZN(pe_1_1_3_n89) );
  INV_X1 pe_1_1_3_U5 ( .A(pe_1_1_3_n40), .ZN(pe_1_1_3_n85) );
  INV_X2 pe_1_1_3_U4 ( .A(n81), .ZN(pe_1_1_3_n72) );
  XOR2_X1 pe_1_1_3_U3 ( .A(pe_1_1_3_int_data_0_), .B(int_data_res_1__3__0_), 
        .Z(pe_1_1_3_n1) );
  DFFR_X1 pe_1_1_3_int_q_acc_reg_0_ ( .D(pe_1_1_3_n84), .CK(pe_1_1_3_net6694), 
        .RN(pe_1_1_3_n72), .Q(int_data_res_1__3__0_), .QN(pe_1_1_3_n3) );
  DFFR_X1 pe_1_1_3_int_q_reg_v_reg_0__0_ ( .D(int_data_y_2__3__0_), .CK(
        pe_1_1_3_net6664), .RN(pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_v[20]) );
  DFFR_X1 pe_1_1_3_int_q_reg_v_reg_0__1_ ( .D(int_data_y_2__3__1_), .CK(
        pe_1_1_3_net6664), .RN(pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_v[21]) );
  DFFR_X1 pe_1_1_3_int_q_reg_v_reg_0__2_ ( .D(int_data_y_2__3__2_), .CK(
        pe_1_1_3_net6664), .RN(pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_v[22]) );
  DFFR_X1 pe_1_1_3_int_q_reg_v_reg_0__3_ ( .D(int_data_y_2__3__3_), .CK(
        pe_1_1_3_net6664), .RN(pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_v[23]) );
  DFFR_X1 pe_1_1_3_int_q_reg_v_reg_1__0_ ( .D(int_data_y_2__3__0_), .CK(
        pe_1_1_3_net6669), .RN(pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_v[16]) );
  DFFR_X1 pe_1_1_3_int_q_reg_v_reg_1__1_ ( .D(int_data_y_2__3__1_), .CK(
        pe_1_1_3_net6669), .RN(pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_v[17]) );
  DFFR_X1 pe_1_1_3_int_q_reg_v_reg_1__2_ ( .D(int_data_y_2__3__2_), .CK(
        pe_1_1_3_net6669), .RN(pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_v[18]) );
  DFFR_X1 pe_1_1_3_int_q_reg_v_reg_1__3_ ( .D(int_data_y_2__3__3_), .CK(
        pe_1_1_3_net6669), .RN(pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_v[19]) );
  DFFR_X1 pe_1_1_3_int_q_reg_v_reg_2__0_ ( .D(int_data_y_2__3__0_), .CK(
        pe_1_1_3_net6674), .RN(pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_v[12]) );
  DFFR_X1 pe_1_1_3_int_q_reg_v_reg_2__1_ ( .D(int_data_y_2__3__1_), .CK(
        pe_1_1_3_net6674), .RN(pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_v[13]) );
  DFFR_X1 pe_1_1_3_int_q_reg_v_reg_2__2_ ( .D(int_data_y_2__3__2_), .CK(
        pe_1_1_3_net6674), .RN(pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_v[14]) );
  DFFR_X1 pe_1_1_3_int_q_reg_v_reg_2__3_ ( .D(int_data_y_2__3__3_), .CK(
        pe_1_1_3_net6674), .RN(pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_v[15]) );
  DFFR_X1 pe_1_1_3_int_q_reg_v_reg_3__0_ ( .D(int_data_y_2__3__0_), .CK(
        pe_1_1_3_net6679), .RN(pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_v[8]) );
  DFFR_X1 pe_1_1_3_int_q_reg_v_reg_3__1_ ( .D(int_data_y_2__3__1_), .CK(
        pe_1_1_3_net6679), .RN(pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_v[9]) );
  DFFR_X1 pe_1_1_3_int_q_reg_v_reg_3__2_ ( .D(int_data_y_2__3__2_), .CK(
        pe_1_1_3_net6679), .RN(pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_v[10]) );
  DFFR_X1 pe_1_1_3_int_q_reg_v_reg_3__3_ ( .D(int_data_y_2__3__3_), .CK(
        pe_1_1_3_net6679), .RN(pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_v[11]) );
  DFFR_X1 pe_1_1_3_int_q_reg_v_reg_4__0_ ( .D(int_data_y_2__3__0_), .CK(
        pe_1_1_3_net6684), .RN(pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_v[4]) );
  DFFR_X1 pe_1_1_3_int_q_reg_v_reg_4__1_ ( .D(int_data_y_2__3__1_), .CK(
        pe_1_1_3_net6684), .RN(pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_v[5]) );
  DFFR_X1 pe_1_1_3_int_q_reg_v_reg_4__2_ ( .D(int_data_y_2__3__2_), .CK(
        pe_1_1_3_net6684), .RN(pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_v[6]) );
  DFFR_X1 pe_1_1_3_int_q_reg_v_reg_4__3_ ( .D(int_data_y_2__3__3_), .CK(
        pe_1_1_3_net6684), .RN(pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_v[7]) );
  DFFR_X1 pe_1_1_3_int_q_reg_v_reg_5__0_ ( .D(int_data_y_2__3__0_), .CK(
        pe_1_1_3_net6689), .RN(pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_v[0]) );
  DFFR_X1 pe_1_1_3_int_q_reg_v_reg_5__1_ ( .D(int_data_y_2__3__1_), .CK(
        pe_1_1_3_net6689), .RN(pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_v[1]) );
  DFFR_X1 pe_1_1_3_int_q_reg_v_reg_5__2_ ( .D(int_data_y_2__3__2_), .CK(
        pe_1_1_3_net6689), .RN(pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_v[2]) );
  DFFR_X1 pe_1_1_3_int_q_reg_v_reg_5__3_ ( .D(int_data_y_2__3__3_), .CK(
        pe_1_1_3_net6689), .RN(pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_1_3_int_q_reg_h_reg_0__0_ ( .D(int_data_x_1__4__0_), .SI(
        int_data_y_2__3__0_), .SE(pe_1_1_3_n65), .CK(pe_1_1_3_net6633), .RN(
        pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_1_3_int_q_reg_h_reg_0__1_ ( .D(int_data_x_1__4__1_), .SI(
        int_data_y_2__3__1_), .SE(pe_1_1_3_n65), .CK(pe_1_1_3_net6633), .RN(
        pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_1_3_int_q_reg_h_reg_0__2_ ( .D(int_data_x_1__4__2_), .SI(
        int_data_y_2__3__2_), .SE(pe_1_1_3_n65), .CK(pe_1_1_3_net6633), .RN(
        pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_1_3_int_q_reg_h_reg_0__3_ ( .D(int_data_x_1__4__3_), .SI(
        int_data_y_2__3__3_), .SE(pe_1_1_3_n65), .CK(pe_1_1_3_net6633), .RN(
        pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_1_3_int_q_reg_h_reg_1__0_ ( .D(int_data_x_1__4__0_), .SI(
        int_data_y_2__3__0_), .SE(pe_1_1_3_n65), .CK(pe_1_1_3_net6639), .RN(
        pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_1_3_int_q_reg_h_reg_1__1_ ( .D(int_data_x_1__4__1_), .SI(
        int_data_y_2__3__1_), .SE(pe_1_1_3_n65), .CK(pe_1_1_3_net6639), .RN(
        pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_1_3_int_q_reg_h_reg_1__2_ ( .D(int_data_x_1__4__2_), .SI(
        int_data_y_2__3__2_), .SE(pe_1_1_3_n65), .CK(pe_1_1_3_net6639), .RN(
        pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_1_3_int_q_reg_h_reg_1__3_ ( .D(int_data_x_1__4__3_), .SI(
        int_data_y_2__3__3_), .SE(pe_1_1_3_n65), .CK(pe_1_1_3_net6639), .RN(
        pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_1_3_int_q_reg_h_reg_2__0_ ( .D(int_data_x_1__4__0_), .SI(
        int_data_y_2__3__0_), .SE(pe_1_1_3_n65), .CK(pe_1_1_3_net6644), .RN(
        pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_1_3_int_q_reg_h_reg_2__1_ ( .D(int_data_x_1__4__1_), .SI(
        int_data_y_2__3__1_), .SE(pe_1_1_3_n65), .CK(pe_1_1_3_net6644), .RN(
        pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_1_3_int_q_reg_h_reg_2__2_ ( .D(int_data_x_1__4__2_), .SI(
        int_data_y_2__3__2_), .SE(pe_1_1_3_n65), .CK(pe_1_1_3_net6644), .RN(
        pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_1_3_int_q_reg_h_reg_2__3_ ( .D(int_data_x_1__4__3_), .SI(
        int_data_y_2__3__3_), .SE(pe_1_1_3_n65), .CK(pe_1_1_3_net6644), .RN(
        pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_1_3_int_q_reg_h_reg_3__0_ ( .D(int_data_x_1__4__0_), .SI(
        int_data_y_2__3__0_), .SE(pe_1_1_3_n65), .CK(pe_1_1_3_net6649), .RN(
        pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_1_3_int_q_reg_h_reg_3__1_ ( .D(int_data_x_1__4__1_), .SI(
        int_data_y_2__3__1_), .SE(pe_1_1_3_n65), .CK(pe_1_1_3_net6649), .RN(
        pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_1_3_int_q_reg_h_reg_3__2_ ( .D(int_data_x_1__4__2_), .SI(
        int_data_y_2__3__2_), .SE(pe_1_1_3_n65), .CK(pe_1_1_3_net6649), .RN(
        pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_1_3_int_q_reg_h_reg_3__3_ ( .D(int_data_x_1__4__3_), .SI(
        int_data_y_2__3__3_), .SE(pe_1_1_3_n65), .CK(pe_1_1_3_net6649), .RN(
        pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_1_3_int_q_reg_h_reg_4__0_ ( .D(int_data_x_1__4__0_), .SI(
        int_data_y_2__3__0_), .SE(pe_1_1_3_n66), .CK(pe_1_1_3_net6654), .RN(
        pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_1_3_int_q_reg_h_reg_4__1_ ( .D(int_data_x_1__4__1_), .SI(
        int_data_y_2__3__1_), .SE(pe_1_1_3_n66), .CK(pe_1_1_3_net6654), .RN(
        pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_1_3_int_q_reg_h_reg_4__2_ ( .D(int_data_x_1__4__2_), .SI(
        int_data_y_2__3__2_), .SE(pe_1_1_3_n66), .CK(pe_1_1_3_net6654), .RN(
        pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_1_3_int_q_reg_h_reg_4__3_ ( .D(int_data_x_1__4__3_), .SI(
        int_data_y_2__3__3_), .SE(pe_1_1_3_n66), .CK(pe_1_1_3_net6654), .RN(
        pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_1_3_int_q_reg_h_reg_5__0_ ( .D(int_data_x_1__4__0_), .SI(
        int_data_y_2__3__0_), .SE(pe_1_1_3_n66), .CK(pe_1_1_3_net6659), .RN(
        pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_1_3_int_q_reg_h_reg_5__1_ ( .D(int_data_x_1__4__1_), .SI(
        int_data_y_2__3__1_), .SE(pe_1_1_3_n66), .CK(pe_1_1_3_net6659), .RN(
        pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_1_3_int_q_reg_h_reg_5__2_ ( .D(int_data_x_1__4__2_), .SI(
        int_data_y_2__3__2_), .SE(pe_1_1_3_n66), .CK(pe_1_1_3_net6659), .RN(
        pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_1_3_int_q_reg_h_reg_5__3_ ( .D(int_data_x_1__4__3_), .SI(
        int_data_y_2__3__3_), .SE(pe_1_1_3_n66), .CK(pe_1_1_3_net6659), .RN(
        pe_1_1_3_n72), .Q(pe_1_1_3_int_q_reg_h[3]) );
  FA_X1 pe_1_1_3_sub_81_U2_7 ( .A(int_data_res_1__3__7_), .B(pe_1_1_3_n76), 
        .CI(pe_1_1_3_sub_81_carry[7]), .S(pe_1_1_3_N77) );
  FA_X1 pe_1_1_3_sub_81_U2_6 ( .A(int_data_res_1__3__6_), .B(pe_1_1_3_n76), 
        .CI(pe_1_1_3_sub_81_carry[6]), .CO(pe_1_1_3_sub_81_carry[7]), .S(
        pe_1_1_3_N76) );
  FA_X1 pe_1_1_3_sub_81_U2_5 ( .A(int_data_res_1__3__5_), .B(pe_1_1_3_n76), 
        .CI(pe_1_1_3_sub_81_carry[5]), .CO(pe_1_1_3_sub_81_carry[6]), .S(
        pe_1_1_3_N75) );
  FA_X1 pe_1_1_3_sub_81_U2_4 ( .A(int_data_res_1__3__4_), .B(pe_1_1_3_n76), 
        .CI(pe_1_1_3_sub_81_carry[4]), .CO(pe_1_1_3_sub_81_carry[5]), .S(
        pe_1_1_3_N74) );
  FA_X1 pe_1_1_3_sub_81_U2_3 ( .A(int_data_res_1__3__3_), .B(pe_1_1_3_n76), 
        .CI(pe_1_1_3_sub_81_carry[3]), .CO(pe_1_1_3_sub_81_carry[4]), .S(
        pe_1_1_3_N73) );
  FA_X1 pe_1_1_3_sub_81_U2_2 ( .A(int_data_res_1__3__2_), .B(pe_1_1_3_n75), 
        .CI(pe_1_1_3_sub_81_carry[2]), .CO(pe_1_1_3_sub_81_carry[3]), .S(
        pe_1_1_3_N72) );
  FA_X1 pe_1_1_3_sub_81_U2_1 ( .A(int_data_res_1__3__1_), .B(pe_1_1_3_n74), 
        .CI(pe_1_1_3_sub_81_carry[1]), .CO(pe_1_1_3_sub_81_carry[2]), .S(
        pe_1_1_3_N71) );
  FA_X1 pe_1_1_3_add_83_U1_7 ( .A(int_data_res_1__3__7_), .B(
        pe_1_1_3_int_data_3_), .CI(pe_1_1_3_add_83_carry[7]), .S(pe_1_1_3_N85)
         );
  FA_X1 pe_1_1_3_add_83_U1_6 ( .A(int_data_res_1__3__6_), .B(
        pe_1_1_3_int_data_3_), .CI(pe_1_1_3_add_83_carry[6]), .CO(
        pe_1_1_3_add_83_carry[7]), .S(pe_1_1_3_N84) );
  FA_X1 pe_1_1_3_add_83_U1_5 ( .A(int_data_res_1__3__5_), .B(
        pe_1_1_3_int_data_3_), .CI(pe_1_1_3_add_83_carry[5]), .CO(
        pe_1_1_3_add_83_carry[6]), .S(pe_1_1_3_N83) );
  FA_X1 pe_1_1_3_add_83_U1_4 ( .A(int_data_res_1__3__4_), .B(
        pe_1_1_3_int_data_3_), .CI(pe_1_1_3_add_83_carry[4]), .CO(
        pe_1_1_3_add_83_carry[5]), .S(pe_1_1_3_N82) );
  FA_X1 pe_1_1_3_add_83_U1_3 ( .A(int_data_res_1__3__3_), .B(
        pe_1_1_3_int_data_3_), .CI(pe_1_1_3_add_83_carry[3]), .CO(
        pe_1_1_3_add_83_carry[4]), .S(pe_1_1_3_N81) );
  FA_X1 pe_1_1_3_add_83_U1_2 ( .A(int_data_res_1__3__2_), .B(
        pe_1_1_3_int_data_2_), .CI(pe_1_1_3_add_83_carry[2]), .CO(
        pe_1_1_3_add_83_carry[3]), .S(pe_1_1_3_N80) );
  FA_X1 pe_1_1_3_add_83_U1_1 ( .A(int_data_res_1__3__1_), .B(
        pe_1_1_3_int_data_1_), .CI(pe_1_1_3_n2), .CO(pe_1_1_3_add_83_carry[2]), 
        .S(pe_1_1_3_N79) );
  NAND3_X1 pe_1_1_3_U56 ( .A1(pe_1_1_3_n60), .A2(pe_1_1_3_n43), .A3(
        pe_1_1_3_n62), .ZN(pe_1_1_3_n40) );
  NAND3_X1 pe_1_1_3_U55 ( .A1(pe_1_1_3_n43), .A2(pe_1_1_3_n61), .A3(
        pe_1_1_3_n62), .ZN(pe_1_1_3_n39) );
  NAND3_X1 pe_1_1_3_U54 ( .A1(pe_1_1_3_n43), .A2(pe_1_1_3_n63), .A3(
        pe_1_1_3_n60), .ZN(pe_1_1_3_n38) );
  NAND3_X1 pe_1_1_3_U53 ( .A1(pe_1_1_3_n61), .A2(pe_1_1_3_n63), .A3(
        pe_1_1_3_n43), .ZN(pe_1_1_3_n37) );
  DFFR_X1 pe_1_1_3_int_q_acc_reg_6_ ( .D(pe_1_1_3_n78), .CK(pe_1_1_3_net6694), 
        .RN(pe_1_1_3_n71), .Q(int_data_res_1__3__6_) );
  DFFR_X1 pe_1_1_3_int_q_acc_reg_5_ ( .D(pe_1_1_3_n79), .CK(pe_1_1_3_net6694), 
        .RN(pe_1_1_3_n71), .Q(int_data_res_1__3__5_) );
  DFFR_X1 pe_1_1_3_int_q_acc_reg_4_ ( .D(pe_1_1_3_n80), .CK(pe_1_1_3_net6694), 
        .RN(pe_1_1_3_n71), .Q(int_data_res_1__3__4_) );
  DFFR_X1 pe_1_1_3_int_q_acc_reg_3_ ( .D(pe_1_1_3_n81), .CK(pe_1_1_3_net6694), 
        .RN(pe_1_1_3_n71), .Q(int_data_res_1__3__3_) );
  DFFR_X1 pe_1_1_3_int_q_acc_reg_2_ ( .D(pe_1_1_3_n82), .CK(pe_1_1_3_net6694), 
        .RN(pe_1_1_3_n71), .Q(int_data_res_1__3__2_) );
  DFFR_X1 pe_1_1_3_int_q_acc_reg_1_ ( .D(pe_1_1_3_n83), .CK(pe_1_1_3_net6694), 
        .RN(pe_1_1_3_n71), .Q(int_data_res_1__3__1_) );
  DFFR_X1 pe_1_1_3_int_q_acc_reg_7_ ( .D(pe_1_1_3_n77), .CK(pe_1_1_3_net6694), 
        .RN(pe_1_1_3_n71), .Q(int_data_res_1__3__7_) );
  CLKGATETST_X1 pe_1_1_3_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_1_3_n88), .SE(1'b0), .GCK(pe_1_1_3_net6633) );
  CLKGATETST_X1 pe_1_1_3_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_1_3_n87), .SE(1'b0), .GCK(pe_1_1_3_net6639) );
  CLKGATETST_X1 pe_1_1_3_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_1_3_n86), .SE(1'b0), .GCK(pe_1_1_3_net6644) );
  CLKGATETST_X1 pe_1_1_3_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_1_3_n85), .SE(1'b0), .GCK(pe_1_1_3_net6649) );
  CLKGATETST_X1 pe_1_1_3_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_1_3_n90), .SE(1'b0), .GCK(pe_1_1_3_net6654) );
  CLKGATETST_X1 pe_1_1_3_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_1_3_n89), .SE(1'b0), .GCK(pe_1_1_3_net6659) );
  CLKGATETST_X1 pe_1_1_3_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_1_3_N64), .SE(1'b0), .GCK(pe_1_1_3_net6664) );
  CLKGATETST_X1 pe_1_1_3_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_1_3_N63), .SE(1'b0), .GCK(pe_1_1_3_net6669) );
  CLKGATETST_X1 pe_1_1_3_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_1_3_N62), .SE(1'b0), .GCK(pe_1_1_3_net6674) );
  CLKGATETST_X1 pe_1_1_3_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_1_3_N61), .SE(1'b0), .GCK(pe_1_1_3_net6679) );
  CLKGATETST_X1 pe_1_1_3_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_1_3_N60), .SE(1'b0), .GCK(pe_1_1_3_net6684) );
  CLKGATETST_X1 pe_1_1_3_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_1_3_N59), .SE(1'b0), .GCK(pe_1_1_3_net6689) );
  CLKGATETST_X1 pe_1_1_3_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_1_3_N90), .SE(1'b0), .GCK(pe_1_1_3_net6694) );
  CLKBUF_X1 pe_1_1_4_U108 ( .A(pe_1_1_4_n68), .Z(pe_1_1_4_n67) );
  INV_X1 pe_1_1_4_U107 ( .A(n74), .ZN(pe_1_1_4_n66) );
  INV_X1 pe_1_1_4_U106 ( .A(n66), .ZN(pe_1_1_4_n65) );
  INV_X1 pe_1_1_4_U105 ( .A(n66), .ZN(pe_1_1_4_n64) );
  INV_X1 pe_1_1_4_U104 ( .A(pe_1_1_4_n65), .ZN(pe_1_1_4_n63) );
  INV_X1 pe_1_1_4_U103 ( .A(n26), .ZN(pe_1_1_4_n58) );
  INV_X1 pe_1_1_4_U102 ( .A(n18), .ZN(pe_1_1_4_n57) );
  MUX2_X1 pe_1_1_4_U101 ( .A(pe_1_1_4_n54), .B(pe_1_1_4_n51), .S(n45), .Z(
        int_data_x_1__4__3_) );
  MUX2_X1 pe_1_1_4_U100 ( .A(pe_1_1_4_n53), .B(pe_1_1_4_n52), .S(n38), .Z(
        pe_1_1_4_n54) );
  MUX2_X1 pe_1_1_4_U99 ( .A(pe_1_1_4_int_q_reg_h[23]), .B(
        pe_1_1_4_int_q_reg_h[19]), .S(pe_1_1_4_n56), .Z(pe_1_1_4_n53) );
  MUX2_X1 pe_1_1_4_U98 ( .A(pe_1_1_4_int_q_reg_h[15]), .B(
        pe_1_1_4_int_q_reg_h[11]), .S(pe_1_1_4_n56), .Z(pe_1_1_4_n52) );
  MUX2_X1 pe_1_1_4_U97 ( .A(pe_1_1_4_int_q_reg_h[7]), .B(
        pe_1_1_4_int_q_reg_h[3]), .S(pe_1_1_4_n56), .Z(pe_1_1_4_n51) );
  MUX2_X1 pe_1_1_4_U96 ( .A(pe_1_1_4_n50), .B(pe_1_1_4_n47), .S(n45), .Z(
        int_data_x_1__4__2_) );
  MUX2_X1 pe_1_1_4_U95 ( .A(pe_1_1_4_n49), .B(pe_1_1_4_n48), .S(n38), .Z(
        pe_1_1_4_n50) );
  MUX2_X1 pe_1_1_4_U94 ( .A(pe_1_1_4_int_q_reg_h[22]), .B(
        pe_1_1_4_int_q_reg_h[18]), .S(pe_1_1_4_n56), .Z(pe_1_1_4_n49) );
  MUX2_X1 pe_1_1_4_U93 ( .A(pe_1_1_4_int_q_reg_h[14]), .B(
        pe_1_1_4_int_q_reg_h[10]), .S(pe_1_1_4_n56), .Z(pe_1_1_4_n48) );
  MUX2_X1 pe_1_1_4_U92 ( .A(pe_1_1_4_int_q_reg_h[6]), .B(
        pe_1_1_4_int_q_reg_h[2]), .S(pe_1_1_4_n56), .Z(pe_1_1_4_n47) );
  MUX2_X1 pe_1_1_4_U91 ( .A(pe_1_1_4_n46), .B(pe_1_1_4_n24), .S(n45), .Z(
        int_data_x_1__4__1_) );
  MUX2_X1 pe_1_1_4_U90 ( .A(pe_1_1_4_n45), .B(pe_1_1_4_n25), .S(n38), .Z(
        pe_1_1_4_n46) );
  MUX2_X1 pe_1_1_4_U89 ( .A(pe_1_1_4_int_q_reg_h[21]), .B(
        pe_1_1_4_int_q_reg_h[17]), .S(pe_1_1_4_n56), .Z(pe_1_1_4_n45) );
  MUX2_X1 pe_1_1_4_U88 ( .A(pe_1_1_4_int_q_reg_h[13]), .B(
        pe_1_1_4_int_q_reg_h[9]), .S(pe_1_1_4_n56), .Z(pe_1_1_4_n25) );
  MUX2_X1 pe_1_1_4_U87 ( .A(pe_1_1_4_int_q_reg_h[5]), .B(
        pe_1_1_4_int_q_reg_h[1]), .S(pe_1_1_4_n56), .Z(pe_1_1_4_n24) );
  MUX2_X1 pe_1_1_4_U86 ( .A(pe_1_1_4_n23), .B(pe_1_1_4_n20), .S(n45), .Z(
        int_data_x_1__4__0_) );
  MUX2_X1 pe_1_1_4_U85 ( .A(pe_1_1_4_n22), .B(pe_1_1_4_n21), .S(n38), .Z(
        pe_1_1_4_n23) );
  MUX2_X1 pe_1_1_4_U84 ( .A(pe_1_1_4_int_q_reg_h[20]), .B(
        pe_1_1_4_int_q_reg_h[16]), .S(pe_1_1_4_n56), .Z(pe_1_1_4_n22) );
  MUX2_X1 pe_1_1_4_U83 ( .A(pe_1_1_4_int_q_reg_h[12]), .B(
        pe_1_1_4_int_q_reg_h[8]), .S(pe_1_1_4_n56), .Z(pe_1_1_4_n21) );
  MUX2_X1 pe_1_1_4_U82 ( .A(pe_1_1_4_int_q_reg_h[4]), .B(
        pe_1_1_4_int_q_reg_h[0]), .S(pe_1_1_4_n56), .Z(pe_1_1_4_n20) );
  MUX2_X1 pe_1_1_4_U81 ( .A(pe_1_1_4_n19), .B(pe_1_1_4_n16), .S(n45), .Z(
        int_data_y_1__4__3_) );
  MUX2_X1 pe_1_1_4_U80 ( .A(pe_1_1_4_n18), .B(pe_1_1_4_n17), .S(n38), .Z(
        pe_1_1_4_n19) );
  MUX2_X1 pe_1_1_4_U79 ( .A(pe_1_1_4_int_q_reg_v[23]), .B(
        pe_1_1_4_int_q_reg_v[19]), .S(pe_1_1_4_n55), .Z(pe_1_1_4_n18) );
  MUX2_X1 pe_1_1_4_U78 ( .A(pe_1_1_4_int_q_reg_v[15]), .B(
        pe_1_1_4_int_q_reg_v[11]), .S(pe_1_1_4_n55), .Z(pe_1_1_4_n17) );
  MUX2_X1 pe_1_1_4_U77 ( .A(pe_1_1_4_int_q_reg_v[7]), .B(
        pe_1_1_4_int_q_reg_v[3]), .S(pe_1_1_4_n55), .Z(pe_1_1_4_n16) );
  MUX2_X1 pe_1_1_4_U76 ( .A(pe_1_1_4_n15), .B(pe_1_1_4_n12), .S(n45), .Z(
        int_data_y_1__4__2_) );
  MUX2_X1 pe_1_1_4_U75 ( .A(pe_1_1_4_n14), .B(pe_1_1_4_n13), .S(n38), .Z(
        pe_1_1_4_n15) );
  MUX2_X1 pe_1_1_4_U74 ( .A(pe_1_1_4_int_q_reg_v[22]), .B(
        pe_1_1_4_int_q_reg_v[18]), .S(pe_1_1_4_n55), .Z(pe_1_1_4_n14) );
  MUX2_X1 pe_1_1_4_U73 ( .A(pe_1_1_4_int_q_reg_v[14]), .B(
        pe_1_1_4_int_q_reg_v[10]), .S(pe_1_1_4_n55), .Z(pe_1_1_4_n13) );
  MUX2_X1 pe_1_1_4_U72 ( .A(pe_1_1_4_int_q_reg_v[6]), .B(
        pe_1_1_4_int_q_reg_v[2]), .S(pe_1_1_4_n55), .Z(pe_1_1_4_n12) );
  MUX2_X1 pe_1_1_4_U71 ( .A(pe_1_1_4_n11), .B(pe_1_1_4_n8), .S(n45), .Z(
        int_data_y_1__4__1_) );
  MUX2_X1 pe_1_1_4_U70 ( .A(pe_1_1_4_n10), .B(pe_1_1_4_n9), .S(n38), .Z(
        pe_1_1_4_n11) );
  MUX2_X1 pe_1_1_4_U69 ( .A(pe_1_1_4_int_q_reg_v[21]), .B(
        pe_1_1_4_int_q_reg_v[17]), .S(pe_1_1_4_n55), .Z(pe_1_1_4_n10) );
  MUX2_X1 pe_1_1_4_U68 ( .A(pe_1_1_4_int_q_reg_v[13]), .B(
        pe_1_1_4_int_q_reg_v[9]), .S(pe_1_1_4_n55), .Z(pe_1_1_4_n9) );
  MUX2_X1 pe_1_1_4_U67 ( .A(pe_1_1_4_int_q_reg_v[5]), .B(
        pe_1_1_4_int_q_reg_v[1]), .S(pe_1_1_4_n55), .Z(pe_1_1_4_n8) );
  MUX2_X1 pe_1_1_4_U66 ( .A(pe_1_1_4_n7), .B(pe_1_1_4_n4), .S(n45), .Z(
        int_data_y_1__4__0_) );
  MUX2_X1 pe_1_1_4_U65 ( .A(pe_1_1_4_n6), .B(pe_1_1_4_n5), .S(n38), .Z(
        pe_1_1_4_n7) );
  MUX2_X1 pe_1_1_4_U64 ( .A(pe_1_1_4_int_q_reg_v[20]), .B(
        pe_1_1_4_int_q_reg_v[16]), .S(pe_1_1_4_n55), .Z(pe_1_1_4_n6) );
  MUX2_X1 pe_1_1_4_U63 ( .A(pe_1_1_4_int_q_reg_v[12]), .B(
        pe_1_1_4_int_q_reg_v[8]), .S(pe_1_1_4_n55), .Z(pe_1_1_4_n5) );
  MUX2_X1 pe_1_1_4_U62 ( .A(pe_1_1_4_int_q_reg_v[4]), .B(
        pe_1_1_4_int_q_reg_v[0]), .S(pe_1_1_4_n55), .Z(pe_1_1_4_n4) );
  AOI222_X1 pe_1_1_4_U61 ( .A1(int_data_res_2__4__2_), .A2(pe_1_1_4_n61), .B1(
        pe_1_1_4_N80), .B2(pe_1_1_4_n27), .C1(pe_1_1_4_N72), .C2(pe_1_1_4_n28), 
        .ZN(pe_1_1_4_n33) );
  INV_X1 pe_1_1_4_U60 ( .A(pe_1_1_4_n33), .ZN(pe_1_1_4_n78) );
  AOI222_X1 pe_1_1_4_U59 ( .A1(int_data_res_2__4__6_), .A2(pe_1_1_4_n61), .B1(
        pe_1_1_4_N84), .B2(pe_1_1_4_n27), .C1(pe_1_1_4_N76), .C2(pe_1_1_4_n28), 
        .ZN(pe_1_1_4_n29) );
  INV_X1 pe_1_1_4_U58 ( .A(pe_1_1_4_n29), .ZN(pe_1_1_4_n74) );
  XNOR2_X1 pe_1_1_4_U57 ( .A(pe_1_1_4_n69), .B(int_data_res_1__4__0_), .ZN(
        pe_1_1_4_N70) );
  AOI222_X1 pe_1_1_4_U52 ( .A1(int_data_res_2__4__0_), .A2(pe_1_1_4_n61), .B1(
        pe_1_1_4_n1), .B2(pe_1_1_4_n27), .C1(pe_1_1_4_N70), .C2(pe_1_1_4_n28), 
        .ZN(pe_1_1_4_n35) );
  INV_X1 pe_1_1_4_U51 ( .A(pe_1_1_4_n35), .ZN(pe_1_1_4_n80) );
  AOI222_X1 pe_1_1_4_U50 ( .A1(int_data_res_2__4__1_), .A2(pe_1_1_4_n61), .B1(
        pe_1_1_4_N79), .B2(pe_1_1_4_n27), .C1(pe_1_1_4_N71), .C2(pe_1_1_4_n28), 
        .ZN(pe_1_1_4_n34) );
  INV_X1 pe_1_1_4_U49 ( .A(pe_1_1_4_n34), .ZN(pe_1_1_4_n79) );
  AOI222_X1 pe_1_1_4_U48 ( .A1(int_data_res_2__4__3_), .A2(pe_1_1_4_n61), .B1(
        pe_1_1_4_N81), .B2(pe_1_1_4_n27), .C1(pe_1_1_4_N73), .C2(pe_1_1_4_n28), 
        .ZN(pe_1_1_4_n32) );
  INV_X1 pe_1_1_4_U47 ( .A(pe_1_1_4_n32), .ZN(pe_1_1_4_n77) );
  AOI222_X1 pe_1_1_4_U46 ( .A1(int_data_res_2__4__4_), .A2(pe_1_1_4_n61), .B1(
        pe_1_1_4_N82), .B2(pe_1_1_4_n27), .C1(pe_1_1_4_N74), .C2(pe_1_1_4_n28), 
        .ZN(pe_1_1_4_n31) );
  INV_X1 pe_1_1_4_U45 ( .A(pe_1_1_4_n31), .ZN(pe_1_1_4_n76) );
  AOI222_X1 pe_1_1_4_U44 ( .A1(int_data_res_2__4__5_), .A2(pe_1_1_4_n61), .B1(
        pe_1_1_4_N83), .B2(pe_1_1_4_n27), .C1(pe_1_1_4_N75), .C2(pe_1_1_4_n28), 
        .ZN(pe_1_1_4_n30) );
  INV_X1 pe_1_1_4_U43 ( .A(pe_1_1_4_n30), .ZN(pe_1_1_4_n75) );
  NAND2_X1 pe_1_1_4_U42 ( .A1(pe_1_1_4_int_data_0_), .A2(pe_1_1_4_n3), .ZN(
        pe_1_1_4_sub_81_carry[1]) );
  INV_X1 pe_1_1_4_U41 ( .A(pe_1_1_4_int_data_1_), .ZN(pe_1_1_4_n70) );
  INV_X1 pe_1_1_4_U40 ( .A(pe_1_1_4_int_data_2_), .ZN(pe_1_1_4_n71) );
  AND2_X1 pe_1_1_4_U39 ( .A1(pe_1_1_4_int_data_0_), .A2(int_data_res_1__4__0_), 
        .ZN(pe_1_1_4_n2) );
  AOI222_X1 pe_1_1_4_U38 ( .A1(pe_1_1_4_n61), .A2(int_data_res_2__4__7_), .B1(
        pe_1_1_4_N85), .B2(pe_1_1_4_n27), .C1(pe_1_1_4_N77), .C2(pe_1_1_4_n28), 
        .ZN(pe_1_1_4_n26) );
  INV_X1 pe_1_1_4_U37 ( .A(pe_1_1_4_n26), .ZN(pe_1_1_4_n73) );
  NOR3_X1 pe_1_1_4_U36 ( .A1(pe_1_1_4_n58), .A2(pe_1_1_4_n62), .A3(int_ckg[51]), .ZN(pe_1_1_4_n36) );
  OR2_X1 pe_1_1_4_U35 ( .A1(pe_1_1_4_n36), .A2(pe_1_1_4_n61), .ZN(pe_1_1_4_N90) );
  INV_X1 pe_1_1_4_U34 ( .A(n38), .ZN(pe_1_1_4_n60) );
  AND2_X1 pe_1_1_4_U33 ( .A1(int_data_x_1__4__2_), .A2(n26), .ZN(
        pe_1_1_4_int_data_2_) );
  AND2_X1 pe_1_1_4_U32 ( .A1(int_data_x_1__4__1_), .A2(n26), .ZN(
        pe_1_1_4_int_data_1_) );
  AND2_X1 pe_1_1_4_U31 ( .A1(int_data_x_1__4__3_), .A2(n26), .ZN(
        pe_1_1_4_int_data_3_) );
  BUF_X1 pe_1_1_4_U30 ( .A(n60), .Z(pe_1_1_4_n61) );
  INV_X1 pe_1_1_4_U29 ( .A(n32), .ZN(pe_1_1_4_n59) );
  AND2_X1 pe_1_1_4_U28 ( .A1(int_data_x_1__4__0_), .A2(n26), .ZN(
        pe_1_1_4_int_data_0_) );
  NAND2_X1 pe_1_1_4_U27 ( .A1(pe_1_1_4_n44), .A2(pe_1_1_4_n59), .ZN(
        pe_1_1_4_n41) );
  AND3_X1 pe_1_1_4_U26 ( .A1(n74), .A2(pe_1_1_4_n60), .A3(n45), .ZN(
        pe_1_1_4_n44) );
  INV_X1 pe_1_1_4_U25 ( .A(pe_1_1_4_int_data_3_), .ZN(pe_1_1_4_n72) );
  NOR2_X1 pe_1_1_4_U24 ( .A1(pe_1_1_4_n66), .A2(n45), .ZN(pe_1_1_4_n43) );
  NOR2_X1 pe_1_1_4_U23 ( .A1(pe_1_1_4_n57), .A2(pe_1_1_4_n61), .ZN(
        pe_1_1_4_n28) );
  NOR2_X1 pe_1_1_4_U22 ( .A1(n18), .A2(pe_1_1_4_n61), .ZN(pe_1_1_4_n27) );
  INV_X1 pe_1_1_4_U21 ( .A(pe_1_1_4_int_data_0_), .ZN(pe_1_1_4_n69) );
  INV_X1 pe_1_1_4_U20 ( .A(pe_1_1_4_n41), .ZN(pe_1_1_4_n86) );
  INV_X1 pe_1_1_4_U19 ( .A(pe_1_1_4_n37), .ZN(pe_1_1_4_n84) );
  INV_X1 pe_1_1_4_U18 ( .A(pe_1_1_4_n38), .ZN(pe_1_1_4_n83) );
  INV_X1 pe_1_1_4_U17 ( .A(pe_1_1_4_n39), .ZN(pe_1_1_4_n82) );
  NOR2_X1 pe_1_1_4_U16 ( .A1(pe_1_1_4_n64), .A2(pe_1_1_4_n42), .ZN(
        pe_1_1_4_N59) );
  NOR2_X1 pe_1_1_4_U15 ( .A1(pe_1_1_4_n64), .A2(pe_1_1_4_n41), .ZN(
        pe_1_1_4_N60) );
  NOR2_X1 pe_1_1_4_U14 ( .A1(pe_1_1_4_n64), .A2(pe_1_1_4_n38), .ZN(
        pe_1_1_4_N63) );
  NOR2_X1 pe_1_1_4_U13 ( .A1(pe_1_1_4_n64), .A2(pe_1_1_4_n40), .ZN(
        pe_1_1_4_N61) );
  NOR2_X1 pe_1_1_4_U12 ( .A1(pe_1_1_4_n64), .A2(pe_1_1_4_n39), .ZN(
        pe_1_1_4_N62) );
  NOR2_X1 pe_1_1_4_U11 ( .A1(pe_1_1_4_n37), .A2(pe_1_1_4_n64), .ZN(
        pe_1_1_4_N64) );
  NAND2_X1 pe_1_1_4_U10 ( .A1(pe_1_1_4_n44), .A2(n32), .ZN(pe_1_1_4_n42) );
  BUF_X1 pe_1_1_4_U9 ( .A(n32), .Z(pe_1_1_4_n55) );
  INV_X1 pe_1_1_4_U8 ( .A(pe_1_1_4_n65), .ZN(pe_1_1_4_n62) );
  BUF_X1 pe_1_1_4_U7 ( .A(n32), .Z(pe_1_1_4_n56) );
  INV_X1 pe_1_1_4_U6 ( .A(pe_1_1_4_n42), .ZN(pe_1_1_4_n85) );
  INV_X1 pe_1_1_4_U5 ( .A(pe_1_1_4_n40), .ZN(pe_1_1_4_n81) );
  INV_X2 pe_1_1_4_U4 ( .A(n82), .ZN(pe_1_1_4_n68) );
  XOR2_X1 pe_1_1_4_U3 ( .A(pe_1_1_4_int_data_0_), .B(int_data_res_1__4__0_), 
        .Z(pe_1_1_4_n1) );
  DFFR_X1 pe_1_1_4_int_q_acc_reg_0_ ( .D(pe_1_1_4_n80), .CK(pe_1_1_4_net6616), 
        .RN(pe_1_1_4_n68), .Q(int_data_res_1__4__0_), .QN(pe_1_1_4_n3) );
  DFFR_X1 pe_1_1_4_int_q_reg_v_reg_0__0_ ( .D(int_data_y_2__4__0_), .CK(
        pe_1_1_4_net6586), .RN(pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_v[20]) );
  DFFR_X1 pe_1_1_4_int_q_reg_v_reg_0__1_ ( .D(int_data_y_2__4__1_), .CK(
        pe_1_1_4_net6586), .RN(pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_v[21]) );
  DFFR_X1 pe_1_1_4_int_q_reg_v_reg_0__2_ ( .D(int_data_y_2__4__2_), .CK(
        pe_1_1_4_net6586), .RN(pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_v[22]) );
  DFFR_X1 pe_1_1_4_int_q_reg_v_reg_0__3_ ( .D(int_data_y_2__4__3_), .CK(
        pe_1_1_4_net6586), .RN(pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_v[23]) );
  DFFR_X1 pe_1_1_4_int_q_reg_v_reg_1__0_ ( .D(int_data_y_2__4__0_), .CK(
        pe_1_1_4_net6591), .RN(pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_v[16]) );
  DFFR_X1 pe_1_1_4_int_q_reg_v_reg_1__1_ ( .D(int_data_y_2__4__1_), .CK(
        pe_1_1_4_net6591), .RN(pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_v[17]) );
  DFFR_X1 pe_1_1_4_int_q_reg_v_reg_1__2_ ( .D(int_data_y_2__4__2_), .CK(
        pe_1_1_4_net6591), .RN(pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_v[18]) );
  DFFR_X1 pe_1_1_4_int_q_reg_v_reg_1__3_ ( .D(int_data_y_2__4__3_), .CK(
        pe_1_1_4_net6591), .RN(pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_v[19]) );
  DFFR_X1 pe_1_1_4_int_q_reg_v_reg_2__0_ ( .D(int_data_y_2__4__0_), .CK(
        pe_1_1_4_net6596), .RN(pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_v[12]) );
  DFFR_X1 pe_1_1_4_int_q_reg_v_reg_2__1_ ( .D(int_data_y_2__4__1_), .CK(
        pe_1_1_4_net6596), .RN(pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_v[13]) );
  DFFR_X1 pe_1_1_4_int_q_reg_v_reg_2__2_ ( .D(int_data_y_2__4__2_), .CK(
        pe_1_1_4_net6596), .RN(pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_v[14]) );
  DFFR_X1 pe_1_1_4_int_q_reg_v_reg_2__3_ ( .D(int_data_y_2__4__3_), .CK(
        pe_1_1_4_net6596), .RN(pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_v[15]) );
  DFFR_X1 pe_1_1_4_int_q_reg_v_reg_3__0_ ( .D(int_data_y_2__4__0_), .CK(
        pe_1_1_4_net6601), .RN(pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_v[8]) );
  DFFR_X1 pe_1_1_4_int_q_reg_v_reg_3__1_ ( .D(int_data_y_2__4__1_), .CK(
        pe_1_1_4_net6601), .RN(pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_v[9]) );
  DFFR_X1 pe_1_1_4_int_q_reg_v_reg_3__2_ ( .D(int_data_y_2__4__2_), .CK(
        pe_1_1_4_net6601), .RN(pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_v[10]) );
  DFFR_X1 pe_1_1_4_int_q_reg_v_reg_3__3_ ( .D(int_data_y_2__4__3_), .CK(
        pe_1_1_4_net6601), .RN(pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_v[11]) );
  DFFR_X1 pe_1_1_4_int_q_reg_v_reg_4__0_ ( .D(int_data_y_2__4__0_), .CK(
        pe_1_1_4_net6606), .RN(pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_v[4]) );
  DFFR_X1 pe_1_1_4_int_q_reg_v_reg_4__1_ ( .D(int_data_y_2__4__1_), .CK(
        pe_1_1_4_net6606), .RN(pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_v[5]) );
  DFFR_X1 pe_1_1_4_int_q_reg_v_reg_4__2_ ( .D(int_data_y_2__4__2_), .CK(
        pe_1_1_4_net6606), .RN(pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_v[6]) );
  DFFR_X1 pe_1_1_4_int_q_reg_v_reg_4__3_ ( .D(int_data_y_2__4__3_), .CK(
        pe_1_1_4_net6606), .RN(pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_v[7]) );
  DFFR_X1 pe_1_1_4_int_q_reg_v_reg_5__0_ ( .D(int_data_y_2__4__0_), .CK(
        pe_1_1_4_net6611), .RN(pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_v[0]) );
  DFFR_X1 pe_1_1_4_int_q_reg_v_reg_5__1_ ( .D(int_data_y_2__4__1_), .CK(
        pe_1_1_4_net6611), .RN(pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_v[1]) );
  DFFR_X1 pe_1_1_4_int_q_reg_v_reg_5__2_ ( .D(int_data_y_2__4__2_), .CK(
        pe_1_1_4_net6611), .RN(pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_v[2]) );
  DFFR_X1 pe_1_1_4_int_q_reg_v_reg_5__3_ ( .D(int_data_y_2__4__3_), .CK(
        pe_1_1_4_net6611), .RN(pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_1_4_int_q_reg_h_reg_0__0_ ( .D(int_data_x_1__5__0_), .SI(
        int_data_y_2__4__0_), .SE(pe_1_1_4_n62), .CK(pe_1_1_4_net6555), .RN(
        pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_1_4_int_q_reg_h_reg_0__1_ ( .D(int_data_x_1__5__1_), .SI(
        int_data_y_2__4__1_), .SE(pe_1_1_4_n62), .CK(pe_1_1_4_net6555), .RN(
        pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_1_4_int_q_reg_h_reg_0__2_ ( .D(int_data_x_1__5__2_), .SI(
        int_data_y_2__4__2_), .SE(pe_1_1_4_n62), .CK(pe_1_1_4_net6555), .RN(
        pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_1_4_int_q_reg_h_reg_0__3_ ( .D(int_data_x_1__5__3_), .SI(
        int_data_y_2__4__3_), .SE(pe_1_1_4_n62), .CK(pe_1_1_4_net6555), .RN(
        pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_1_4_int_q_reg_h_reg_1__0_ ( .D(int_data_x_1__5__0_), .SI(
        int_data_y_2__4__0_), .SE(pe_1_1_4_n62), .CK(pe_1_1_4_net6561), .RN(
        pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_1_4_int_q_reg_h_reg_1__1_ ( .D(int_data_x_1__5__1_), .SI(
        int_data_y_2__4__1_), .SE(pe_1_1_4_n62), .CK(pe_1_1_4_net6561), .RN(
        pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_1_4_int_q_reg_h_reg_1__2_ ( .D(int_data_x_1__5__2_), .SI(
        int_data_y_2__4__2_), .SE(pe_1_1_4_n62), .CK(pe_1_1_4_net6561), .RN(
        pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_1_4_int_q_reg_h_reg_1__3_ ( .D(int_data_x_1__5__3_), .SI(
        int_data_y_2__4__3_), .SE(pe_1_1_4_n62), .CK(pe_1_1_4_net6561), .RN(
        pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_1_4_int_q_reg_h_reg_2__0_ ( .D(int_data_x_1__5__0_), .SI(
        int_data_y_2__4__0_), .SE(pe_1_1_4_n62), .CK(pe_1_1_4_net6566), .RN(
        pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_1_4_int_q_reg_h_reg_2__1_ ( .D(int_data_x_1__5__1_), .SI(
        int_data_y_2__4__1_), .SE(pe_1_1_4_n62), .CK(pe_1_1_4_net6566), .RN(
        pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_1_4_int_q_reg_h_reg_2__2_ ( .D(int_data_x_1__5__2_), .SI(
        int_data_y_2__4__2_), .SE(pe_1_1_4_n62), .CK(pe_1_1_4_net6566), .RN(
        pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_1_4_int_q_reg_h_reg_2__3_ ( .D(int_data_x_1__5__3_), .SI(
        int_data_y_2__4__3_), .SE(pe_1_1_4_n62), .CK(pe_1_1_4_net6566), .RN(
        pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_1_4_int_q_reg_h_reg_3__0_ ( .D(int_data_x_1__5__0_), .SI(
        int_data_y_2__4__0_), .SE(pe_1_1_4_n62), .CK(pe_1_1_4_net6571), .RN(
        pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_1_4_int_q_reg_h_reg_3__1_ ( .D(int_data_x_1__5__1_), .SI(
        int_data_y_2__4__1_), .SE(pe_1_1_4_n62), .CK(pe_1_1_4_net6571), .RN(
        pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_1_4_int_q_reg_h_reg_3__2_ ( .D(int_data_x_1__5__2_), .SI(
        int_data_y_2__4__2_), .SE(pe_1_1_4_n62), .CK(pe_1_1_4_net6571), .RN(
        pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_1_4_int_q_reg_h_reg_3__3_ ( .D(int_data_x_1__5__3_), .SI(
        int_data_y_2__4__3_), .SE(pe_1_1_4_n62), .CK(pe_1_1_4_net6571), .RN(
        pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_1_4_int_q_reg_h_reg_4__0_ ( .D(int_data_x_1__5__0_), .SI(
        int_data_y_2__4__0_), .SE(pe_1_1_4_n63), .CK(pe_1_1_4_net6576), .RN(
        pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_1_4_int_q_reg_h_reg_4__1_ ( .D(int_data_x_1__5__1_), .SI(
        int_data_y_2__4__1_), .SE(pe_1_1_4_n63), .CK(pe_1_1_4_net6576), .RN(
        pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_1_4_int_q_reg_h_reg_4__2_ ( .D(int_data_x_1__5__2_), .SI(
        int_data_y_2__4__2_), .SE(pe_1_1_4_n63), .CK(pe_1_1_4_net6576), .RN(
        pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_1_4_int_q_reg_h_reg_4__3_ ( .D(int_data_x_1__5__3_), .SI(
        int_data_y_2__4__3_), .SE(pe_1_1_4_n63), .CK(pe_1_1_4_net6576), .RN(
        pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_1_4_int_q_reg_h_reg_5__0_ ( .D(int_data_x_1__5__0_), .SI(
        int_data_y_2__4__0_), .SE(pe_1_1_4_n63), .CK(pe_1_1_4_net6581), .RN(
        pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_1_4_int_q_reg_h_reg_5__1_ ( .D(int_data_x_1__5__1_), .SI(
        int_data_y_2__4__1_), .SE(pe_1_1_4_n63), .CK(pe_1_1_4_net6581), .RN(
        pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_1_4_int_q_reg_h_reg_5__2_ ( .D(int_data_x_1__5__2_), .SI(
        int_data_y_2__4__2_), .SE(pe_1_1_4_n63), .CK(pe_1_1_4_net6581), .RN(
        pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_1_4_int_q_reg_h_reg_5__3_ ( .D(int_data_x_1__5__3_), .SI(
        int_data_y_2__4__3_), .SE(pe_1_1_4_n63), .CK(pe_1_1_4_net6581), .RN(
        pe_1_1_4_n68), .Q(pe_1_1_4_int_q_reg_h[3]) );
  FA_X1 pe_1_1_4_sub_81_U2_7 ( .A(int_data_res_1__4__7_), .B(pe_1_1_4_n72), 
        .CI(pe_1_1_4_sub_81_carry[7]), .S(pe_1_1_4_N77) );
  FA_X1 pe_1_1_4_sub_81_U2_6 ( .A(int_data_res_1__4__6_), .B(pe_1_1_4_n72), 
        .CI(pe_1_1_4_sub_81_carry[6]), .CO(pe_1_1_4_sub_81_carry[7]), .S(
        pe_1_1_4_N76) );
  FA_X1 pe_1_1_4_sub_81_U2_5 ( .A(int_data_res_1__4__5_), .B(pe_1_1_4_n72), 
        .CI(pe_1_1_4_sub_81_carry[5]), .CO(pe_1_1_4_sub_81_carry[6]), .S(
        pe_1_1_4_N75) );
  FA_X1 pe_1_1_4_sub_81_U2_4 ( .A(int_data_res_1__4__4_), .B(pe_1_1_4_n72), 
        .CI(pe_1_1_4_sub_81_carry[4]), .CO(pe_1_1_4_sub_81_carry[5]), .S(
        pe_1_1_4_N74) );
  FA_X1 pe_1_1_4_sub_81_U2_3 ( .A(int_data_res_1__4__3_), .B(pe_1_1_4_n72), 
        .CI(pe_1_1_4_sub_81_carry[3]), .CO(pe_1_1_4_sub_81_carry[4]), .S(
        pe_1_1_4_N73) );
  FA_X1 pe_1_1_4_sub_81_U2_2 ( .A(int_data_res_1__4__2_), .B(pe_1_1_4_n71), 
        .CI(pe_1_1_4_sub_81_carry[2]), .CO(pe_1_1_4_sub_81_carry[3]), .S(
        pe_1_1_4_N72) );
  FA_X1 pe_1_1_4_sub_81_U2_1 ( .A(int_data_res_1__4__1_), .B(pe_1_1_4_n70), 
        .CI(pe_1_1_4_sub_81_carry[1]), .CO(pe_1_1_4_sub_81_carry[2]), .S(
        pe_1_1_4_N71) );
  FA_X1 pe_1_1_4_add_83_U1_7 ( .A(int_data_res_1__4__7_), .B(
        pe_1_1_4_int_data_3_), .CI(pe_1_1_4_add_83_carry[7]), .S(pe_1_1_4_N85)
         );
  FA_X1 pe_1_1_4_add_83_U1_6 ( .A(int_data_res_1__4__6_), .B(
        pe_1_1_4_int_data_3_), .CI(pe_1_1_4_add_83_carry[6]), .CO(
        pe_1_1_4_add_83_carry[7]), .S(pe_1_1_4_N84) );
  FA_X1 pe_1_1_4_add_83_U1_5 ( .A(int_data_res_1__4__5_), .B(
        pe_1_1_4_int_data_3_), .CI(pe_1_1_4_add_83_carry[5]), .CO(
        pe_1_1_4_add_83_carry[6]), .S(pe_1_1_4_N83) );
  FA_X1 pe_1_1_4_add_83_U1_4 ( .A(int_data_res_1__4__4_), .B(
        pe_1_1_4_int_data_3_), .CI(pe_1_1_4_add_83_carry[4]), .CO(
        pe_1_1_4_add_83_carry[5]), .S(pe_1_1_4_N82) );
  FA_X1 pe_1_1_4_add_83_U1_3 ( .A(int_data_res_1__4__3_), .B(
        pe_1_1_4_int_data_3_), .CI(pe_1_1_4_add_83_carry[3]), .CO(
        pe_1_1_4_add_83_carry[4]), .S(pe_1_1_4_N81) );
  FA_X1 pe_1_1_4_add_83_U1_2 ( .A(int_data_res_1__4__2_), .B(
        pe_1_1_4_int_data_2_), .CI(pe_1_1_4_add_83_carry[2]), .CO(
        pe_1_1_4_add_83_carry[3]), .S(pe_1_1_4_N80) );
  FA_X1 pe_1_1_4_add_83_U1_1 ( .A(int_data_res_1__4__1_), .B(
        pe_1_1_4_int_data_1_), .CI(pe_1_1_4_n2), .CO(pe_1_1_4_add_83_carry[2]), 
        .S(pe_1_1_4_N79) );
  NAND3_X1 pe_1_1_4_U56 ( .A1(n32), .A2(pe_1_1_4_n43), .A3(n38), .ZN(
        pe_1_1_4_n40) );
  NAND3_X1 pe_1_1_4_U55 ( .A1(pe_1_1_4_n43), .A2(pe_1_1_4_n59), .A3(n38), .ZN(
        pe_1_1_4_n39) );
  NAND3_X1 pe_1_1_4_U54 ( .A1(pe_1_1_4_n43), .A2(pe_1_1_4_n60), .A3(n32), .ZN(
        pe_1_1_4_n38) );
  NAND3_X1 pe_1_1_4_U53 ( .A1(pe_1_1_4_n59), .A2(pe_1_1_4_n60), .A3(
        pe_1_1_4_n43), .ZN(pe_1_1_4_n37) );
  DFFR_X1 pe_1_1_4_int_q_acc_reg_6_ ( .D(pe_1_1_4_n74), .CK(pe_1_1_4_net6616), 
        .RN(pe_1_1_4_n67), .Q(int_data_res_1__4__6_) );
  DFFR_X1 pe_1_1_4_int_q_acc_reg_5_ ( .D(pe_1_1_4_n75), .CK(pe_1_1_4_net6616), 
        .RN(pe_1_1_4_n67), .Q(int_data_res_1__4__5_) );
  DFFR_X1 pe_1_1_4_int_q_acc_reg_4_ ( .D(pe_1_1_4_n76), .CK(pe_1_1_4_net6616), 
        .RN(pe_1_1_4_n67), .Q(int_data_res_1__4__4_) );
  DFFR_X1 pe_1_1_4_int_q_acc_reg_3_ ( .D(pe_1_1_4_n77), .CK(pe_1_1_4_net6616), 
        .RN(pe_1_1_4_n67), .Q(int_data_res_1__4__3_) );
  DFFR_X1 pe_1_1_4_int_q_acc_reg_2_ ( .D(pe_1_1_4_n78), .CK(pe_1_1_4_net6616), 
        .RN(pe_1_1_4_n67), .Q(int_data_res_1__4__2_) );
  DFFR_X1 pe_1_1_4_int_q_acc_reg_1_ ( .D(pe_1_1_4_n79), .CK(pe_1_1_4_net6616), 
        .RN(pe_1_1_4_n67), .Q(int_data_res_1__4__1_) );
  DFFR_X1 pe_1_1_4_int_q_acc_reg_7_ ( .D(pe_1_1_4_n73), .CK(pe_1_1_4_net6616), 
        .RN(pe_1_1_4_n67), .Q(int_data_res_1__4__7_) );
  CLKGATETST_X1 pe_1_1_4_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_1_4_n84), .SE(1'b0), .GCK(pe_1_1_4_net6555) );
  CLKGATETST_X1 pe_1_1_4_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_1_4_n83), .SE(1'b0), .GCK(pe_1_1_4_net6561) );
  CLKGATETST_X1 pe_1_1_4_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_1_4_n82), .SE(1'b0), .GCK(pe_1_1_4_net6566) );
  CLKGATETST_X1 pe_1_1_4_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_1_4_n81), .SE(1'b0), .GCK(pe_1_1_4_net6571) );
  CLKGATETST_X1 pe_1_1_4_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_1_4_n86), .SE(1'b0), .GCK(pe_1_1_4_net6576) );
  CLKGATETST_X1 pe_1_1_4_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_1_4_n85), .SE(1'b0), .GCK(pe_1_1_4_net6581) );
  CLKGATETST_X1 pe_1_1_4_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_1_4_N64), .SE(1'b0), .GCK(pe_1_1_4_net6586) );
  CLKGATETST_X1 pe_1_1_4_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_1_4_N63), .SE(1'b0), .GCK(pe_1_1_4_net6591) );
  CLKGATETST_X1 pe_1_1_4_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_1_4_N62), .SE(1'b0), .GCK(pe_1_1_4_net6596) );
  CLKGATETST_X1 pe_1_1_4_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_1_4_N61), .SE(1'b0), .GCK(pe_1_1_4_net6601) );
  CLKGATETST_X1 pe_1_1_4_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_1_4_N60), .SE(1'b0), .GCK(pe_1_1_4_net6606) );
  CLKGATETST_X1 pe_1_1_4_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_1_4_N59), .SE(1'b0), .GCK(pe_1_1_4_net6611) );
  CLKGATETST_X1 pe_1_1_4_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_1_4_N90), .SE(1'b0), .GCK(pe_1_1_4_net6616) );
  CLKBUF_X1 pe_1_1_5_U109 ( .A(pe_1_1_5_n69), .Z(pe_1_1_5_n68) );
  INV_X1 pe_1_1_5_U108 ( .A(n74), .ZN(pe_1_1_5_n67) );
  INV_X1 pe_1_1_5_U107 ( .A(n66), .ZN(pe_1_1_5_n66) );
  INV_X1 pe_1_1_5_U106 ( .A(n66), .ZN(pe_1_1_5_n65) );
  INV_X1 pe_1_1_5_U105 ( .A(pe_1_1_5_n66), .ZN(pe_1_1_5_n64) );
  INV_X1 pe_1_1_5_U104 ( .A(pe_1_1_5_n61), .ZN(pe_1_1_5_n60) );
  INV_X1 pe_1_1_5_U103 ( .A(n26), .ZN(pe_1_1_5_n58) );
  INV_X1 pe_1_1_5_U102 ( .A(n18), .ZN(pe_1_1_5_n57) );
  MUX2_X1 pe_1_1_5_U101 ( .A(pe_1_1_5_n54), .B(pe_1_1_5_n51), .S(n45), .Z(
        int_data_x_1__5__3_) );
  MUX2_X1 pe_1_1_5_U100 ( .A(pe_1_1_5_n53), .B(pe_1_1_5_n52), .S(pe_1_1_5_n60), 
        .Z(pe_1_1_5_n54) );
  MUX2_X1 pe_1_1_5_U99 ( .A(pe_1_1_5_int_q_reg_h[23]), .B(
        pe_1_1_5_int_q_reg_h[19]), .S(pe_1_1_5_n56), .Z(pe_1_1_5_n53) );
  MUX2_X1 pe_1_1_5_U98 ( .A(pe_1_1_5_int_q_reg_h[15]), .B(
        pe_1_1_5_int_q_reg_h[11]), .S(pe_1_1_5_n56), .Z(pe_1_1_5_n52) );
  MUX2_X1 pe_1_1_5_U97 ( .A(pe_1_1_5_int_q_reg_h[7]), .B(
        pe_1_1_5_int_q_reg_h[3]), .S(pe_1_1_5_n56), .Z(pe_1_1_5_n51) );
  MUX2_X1 pe_1_1_5_U96 ( .A(pe_1_1_5_n50), .B(pe_1_1_5_n47), .S(n45), .Z(
        int_data_x_1__5__2_) );
  MUX2_X1 pe_1_1_5_U95 ( .A(pe_1_1_5_n49), .B(pe_1_1_5_n48), .S(pe_1_1_5_n60), 
        .Z(pe_1_1_5_n50) );
  MUX2_X1 pe_1_1_5_U94 ( .A(pe_1_1_5_int_q_reg_h[22]), .B(
        pe_1_1_5_int_q_reg_h[18]), .S(pe_1_1_5_n56), .Z(pe_1_1_5_n49) );
  MUX2_X1 pe_1_1_5_U93 ( .A(pe_1_1_5_int_q_reg_h[14]), .B(
        pe_1_1_5_int_q_reg_h[10]), .S(pe_1_1_5_n56), .Z(pe_1_1_5_n48) );
  MUX2_X1 pe_1_1_5_U92 ( .A(pe_1_1_5_int_q_reg_h[6]), .B(
        pe_1_1_5_int_q_reg_h[2]), .S(pe_1_1_5_n56), .Z(pe_1_1_5_n47) );
  MUX2_X1 pe_1_1_5_U91 ( .A(pe_1_1_5_n46), .B(pe_1_1_5_n24), .S(n45), .Z(
        int_data_x_1__5__1_) );
  MUX2_X1 pe_1_1_5_U90 ( .A(pe_1_1_5_n45), .B(pe_1_1_5_n25), .S(pe_1_1_5_n60), 
        .Z(pe_1_1_5_n46) );
  MUX2_X1 pe_1_1_5_U89 ( .A(pe_1_1_5_int_q_reg_h[21]), .B(
        pe_1_1_5_int_q_reg_h[17]), .S(pe_1_1_5_n56), .Z(pe_1_1_5_n45) );
  MUX2_X1 pe_1_1_5_U88 ( .A(pe_1_1_5_int_q_reg_h[13]), .B(
        pe_1_1_5_int_q_reg_h[9]), .S(pe_1_1_5_n56), .Z(pe_1_1_5_n25) );
  MUX2_X1 pe_1_1_5_U87 ( .A(pe_1_1_5_int_q_reg_h[5]), .B(
        pe_1_1_5_int_q_reg_h[1]), .S(pe_1_1_5_n56), .Z(pe_1_1_5_n24) );
  MUX2_X1 pe_1_1_5_U86 ( .A(pe_1_1_5_n23), .B(pe_1_1_5_n20), .S(n45), .Z(
        int_data_x_1__5__0_) );
  MUX2_X1 pe_1_1_5_U85 ( .A(pe_1_1_5_n22), .B(pe_1_1_5_n21), .S(pe_1_1_5_n60), 
        .Z(pe_1_1_5_n23) );
  MUX2_X1 pe_1_1_5_U84 ( .A(pe_1_1_5_int_q_reg_h[20]), .B(
        pe_1_1_5_int_q_reg_h[16]), .S(pe_1_1_5_n56), .Z(pe_1_1_5_n22) );
  MUX2_X1 pe_1_1_5_U83 ( .A(pe_1_1_5_int_q_reg_h[12]), .B(
        pe_1_1_5_int_q_reg_h[8]), .S(pe_1_1_5_n56), .Z(pe_1_1_5_n21) );
  MUX2_X1 pe_1_1_5_U82 ( .A(pe_1_1_5_int_q_reg_h[4]), .B(
        pe_1_1_5_int_q_reg_h[0]), .S(pe_1_1_5_n56), .Z(pe_1_1_5_n20) );
  MUX2_X1 pe_1_1_5_U81 ( .A(pe_1_1_5_n19), .B(pe_1_1_5_n16), .S(n45), .Z(
        int_data_y_1__5__3_) );
  MUX2_X1 pe_1_1_5_U80 ( .A(pe_1_1_5_n18), .B(pe_1_1_5_n17), .S(pe_1_1_5_n60), 
        .Z(pe_1_1_5_n19) );
  MUX2_X1 pe_1_1_5_U79 ( .A(pe_1_1_5_int_q_reg_v[23]), .B(
        pe_1_1_5_int_q_reg_v[19]), .S(pe_1_1_5_n55), .Z(pe_1_1_5_n18) );
  MUX2_X1 pe_1_1_5_U78 ( .A(pe_1_1_5_int_q_reg_v[15]), .B(
        pe_1_1_5_int_q_reg_v[11]), .S(pe_1_1_5_n55), .Z(pe_1_1_5_n17) );
  MUX2_X1 pe_1_1_5_U77 ( .A(pe_1_1_5_int_q_reg_v[7]), .B(
        pe_1_1_5_int_q_reg_v[3]), .S(pe_1_1_5_n55), .Z(pe_1_1_5_n16) );
  MUX2_X1 pe_1_1_5_U76 ( .A(pe_1_1_5_n15), .B(pe_1_1_5_n12), .S(n45), .Z(
        int_data_y_1__5__2_) );
  MUX2_X1 pe_1_1_5_U75 ( .A(pe_1_1_5_n14), .B(pe_1_1_5_n13), .S(pe_1_1_5_n60), 
        .Z(pe_1_1_5_n15) );
  MUX2_X1 pe_1_1_5_U74 ( .A(pe_1_1_5_int_q_reg_v[22]), .B(
        pe_1_1_5_int_q_reg_v[18]), .S(pe_1_1_5_n55), .Z(pe_1_1_5_n14) );
  MUX2_X1 pe_1_1_5_U73 ( .A(pe_1_1_5_int_q_reg_v[14]), .B(
        pe_1_1_5_int_q_reg_v[10]), .S(pe_1_1_5_n55), .Z(pe_1_1_5_n13) );
  MUX2_X1 pe_1_1_5_U72 ( .A(pe_1_1_5_int_q_reg_v[6]), .B(
        pe_1_1_5_int_q_reg_v[2]), .S(pe_1_1_5_n55), .Z(pe_1_1_5_n12) );
  MUX2_X1 pe_1_1_5_U71 ( .A(pe_1_1_5_n11), .B(pe_1_1_5_n8), .S(n45), .Z(
        int_data_y_1__5__1_) );
  MUX2_X1 pe_1_1_5_U70 ( .A(pe_1_1_5_n10), .B(pe_1_1_5_n9), .S(pe_1_1_5_n60), 
        .Z(pe_1_1_5_n11) );
  MUX2_X1 pe_1_1_5_U69 ( .A(pe_1_1_5_int_q_reg_v[21]), .B(
        pe_1_1_5_int_q_reg_v[17]), .S(pe_1_1_5_n55), .Z(pe_1_1_5_n10) );
  MUX2_X1 pe_1_1_5_U68 ( .A(pe_1_1_5_int_q_reg_v[13]), .B(
        pe_1_1_5_int_q_reg_v[9]), .S(pe_1_1_5_n55), .Z(pe_1_1_5_n9) );
  MUX2_X1 pe_1_1_5_U67 ( .A(pe_1_1_5_int_q_reg_v[5]), .B(
        pe_1_1_5_int_q_reg_v[1]), .S(pe_1_1_5_n55), .Z(pe_1_1_5_n8) );
  MUX2_X1 pe_1_1_5_U66 ( .A(pe_1_1_5_n7), .B(pe_1_1_5_n4), .S(n45), .Z(
        int_data_y_1__5__0_) );
  MUX2_X1 pe_1_1_5_U65 ( .A(pe_1_1_5_n6), .B(pe_1_1_5_n5), .S(pe_1_1_5_n60), 
        .Z(pe_1_1_5_n7) );
  MUX2_X1 pe_1_1_5_U64 ( .A(pe_1_1_5_int_q_reg_v[20]), .B(
        pe_1_1_5_int_q_reg_v[16]), .S(pe_1_1_5_n55), .Z(pe_1_1_5_n6) );
  MUX2_X1 pe_1_1_5_U63 ( .A(pe_1_1_5_int_q_reg_v[12]), .B(
        pe_1_1_5_int_q_reg_v[8]), .S(pe_1_1_5_n55), .Z(pe_1_1_5_n5) );
  MUX2_X1 pe_1_1_5_U62 ( .A(pe_1_1_5_int_q_reg_v[4]), .B(
        pe_1_1_5_int_q_reg_v[0]), .S(pe_1_1_5_n55), .Z(pe_1_1_5_n4) );
  AOI222_X1 pe_1_1_5_U61 ( .A1(int_data_res_2__5__2_), .A2(pe_1_1_5_n62), .B1(
        pe_1_1_5_N80), .B2(pe_1_1_5_n27), .C1(pe_1_1_5_N72), .C2(pe_1_1_5_n28), 
        .ZN(pe_1_1_5_n33) );
  INV_X1 pe_1_1_5_U60 ( .A(pe_1_1_5_n33), .ZN(pe_1_1_5_n79) );
  AOI222_X1 pe_1_1_5_U59 ( .A1(int_data_res_2__5__6_), .A2(pe_1_1_5_n62), .B1(
        pe_1_1_5_N84), .B2(pe_1_1_5_n27), .C1(pe_1_1_5_N76), .C2(pe_1_1_5_n28), 
        .ZN(pe_1_1_5_n29) );
  INV_X1 pe_1_1_5_U58 ( .A(pe_1_1_5_n29), .ZN(pe_1_1_5_n75) );
  XNOR2_X1 pe_1_1_5_U57 ( .A(pe_1_1_5_n70), .B(int_data_res_1__5__0_), .ZN(
        pe_1_1_5_N70) );
  AOI222_X1 pe_1_1_5_U52 ( .A1(int_data_res_2__5__0_), .A2(pe_1_1_5_n62), .B1(
        pe_1_1_5_n1), .B2(pe_1_1_5_n27), .C1(pe_1_1_5_N70), .C2(pe_1_1_5_n28), 
        .ZN(pe_1_1_5_n35) );
  INV_X1 pe_1_1_5_U51 ( .A(pe_1_1_5_n35), .ZN(pe_1_1_5_n81) );
  AOI222_X1 pe_1_1_5_U50 ( .A1(int_data_res_2__5__1_), .A2(pe_1_1_5_n62), .B1(
        pe_1_1_5_N79), .B2(pe_1_1_5_n27), .C1(pe_1_1_5_N71), .C2(pe_1_1_5_n28), 
        .ZN(pe_1_1_5_n34) );
  INV_X1 pe_1_1_5_U49 ( .A(pe_1_1_5_n34), .ZN(pe_1_1_5_n80) );
  AOI222_X1 pe_1_1_5_U48 ( .A1(int_data_res_2__5__3_), .A2(pe_1_1_5_n62), .B1(
        pe_1_1_5_N81), .B2(pe_1_1_5_n27), .C1(pe_1_1_5_N73), .C2(pe_1_1_5_n28), 
        .ZN(pe_1_1_5_n32) );
  INV_X1 pe_1_1_5_U47 ( .A(pe_1_1_5_n32), .ZN(pe_1_1_5_n78) );
  AOI222_X1 pe_1_1_5_U46 ( .A1(int_data_res_2__5__4_), .A2(pe_1_1_5_n62), .B1(
        pe_1_1_5_N82), .B2(pe_1_1_5_n27), .C1(pe_1_1_5_N74), .C2(pe_1_1_5_n28), 
        .ZN(pe_1_1_5_n31) );
  INV_X1 pe_1_1_5_U45 ( .A(pe_1_1_5_n31), .ZN(pe_1_1_5_n77) );
  AOI222_X1 pe_1_1_5_U44 ( .A1(int_data_res_2__5__5_), .A2(pe_1_1_5_n62), .B1(
        pe_1_1_5_N83), .B2(pe_1_1_5_n27), .C1(pe_1_1_5_N75), .C2(pe_1_1_5_n28), 
        .ZN(pe_1_1_5_n30) );
  INV_X1 pe_1_1_5_U43 ( .A(pe_1_1_5_n30), .ZN(pe_1_1_5_n76) );
  NAND2_X1 pe_1_1_5_U42 ( .A1(pe_1_1_5_int_data_0_), .A2(pe_1_1_5_n3), .ZN(
        pe_1_1_5_sub_81_carry[1]) );
  INV_X1 pe_1_1_5_U41 ( .A(pe_1_1_5_int_data_1_), .ZN(pe_1_1_5_n71) );
  INV_X1 pe_1_1_5_U40 ( .A(pe_1_1_5_int_data_2_), .ZN(pe_1_1_5_n72) );
  AND2_X1 pe_1_1_5_U39 ( .A1(pe_1_1_5_int_data_0_), .A2(int_data_res_1__5__0_), 
        .ZN(pe_1_1_5_n2) );
  AOI222_X1 pe_1_1_5_U38 ( .A1(pe_1_1_5_n62), .A2(int_data_res_2__5__7_), .B1(
        pe_1_1_5_N85), .B2(pe_1_1_5_n27), .C1(pe_1_1_5_N77), .C2(pe_1_1_5_n28), 
        .ZN(pe_1_1_5_n26) );
  INV_X1 pe_1_1_5_U37 ( .A(pe_1_1_5_n26), .ZN(pe_1_1_5_n74) );
  NOR3_X1 pe_1_1_5_U36 ( .A1(pe_1_1_5_n58), .A2(pe_1_1_5_n63), .A3(int_ckg[50]), .ZN(pe_1_1_5_n36) );
  OR2_X1 pe_1_1_5_U35 ( .A1(pe_1_1_5_n36), .A2(pe_1_1_5_n62), .ZN(pe_1_1_5_N90) );
  INV_X1 pe_1_1_5_U34 ( .A(n38), .ZN(pe_1_1_5_n61) );
  AND2_X1 pe_1_1_5_U33 ( .A1(int_data_x_1__5__2_), .A2(n26), .ZN(
        pe_1_1_5_int_data_2_) );
  AND2_X1 pe_1_1_5_U32 ( .A1(int_data_x_1__5__1_), .A2(n26), .ZN(
        pe_1_1_5_int_data_1_) );
  AND2_X1 pe_1_1_5_U31 ( .A1(int_data_x_1__5__3_), .A2(n26), .ZN(
        pe_1_1_5_int_data_3_) );
  BUF_X1 pe_1_1_5_U30 ( .A(n60), .Z(pe_1_1_5_n62) );
  INV_X1 pe_1_1_5_U29 ( .A(n32), .ZN(pe_1_1_5_n59) );
  AND2_X1 pe_1_1_5_U28 ( .A1(int_data_x_1__5__0_), .A2(n26), .ZN(
        pe_1_1_5_int_data_0_) );
  NAND2_X1 pe_1_1_5_U27 ( .A1(pe_1_1_5_n44), .A2(pe_1_1_5_n59), .ZN(
        pe_1_1_5_n41) );
  AND3_X1 pe_1_1_5_U26 ( .A1(n74), .A2(pe_1_1_5_n61), .A3(n45), .ZN(
        pe_1_1_5_n44) );
  INV_X1 pe_1_1_5_U25 ( .A(pe_1_1_5_int_data_3_), .ZN(pe_1_1_5_n73) );
  NOR2_X1 pe_1_1_5_U24 ( .A1(pe_1_1_5_n67), .A2(n45), .ZN(pe_1_1_5_n43) );
  NOR2_X1 pe_1_1_5_U23 ( .A1(pe_1_1_5_n57), .A2(pe_1_1_5_n62), .ZN(
        pe_1_1_5_n28) );
  NOR2_X1 pe_1_1_5_U22 ( .A1(n18), .A2(pe_1_1_5_n62), .ZN(pe_1_1_5_n27) );
  INV_X1 pe_1_1_5_U21 ( .A(pe_1_1_5_int_data_0_), .ZN(pe_1_1_5_n70) );
  INV_X1 pe_1_1_5_U20 ( .A(pe_1_1_5_n41), .ZN(pe_1_1_5_n87) );
  INV_X1 pe_1_1_5_U19 ( .A(pe_1_1_5_n37), .ZN(pe_1_1_5_n85) );
  INV_X1 pe_1_1_5_U18 ( .A(pe_1_1_5_n38), .ZN(pe_1_1_5_n84) );
  INV_X1 pe_1_1_5_U17 ( .A(pe_1_1_5_n39), .ZN(pe_1_1_5_n83) );
  NOR2_X1 pe_1_1_5_U16 ( .A1(pe_1_1_5_n65), .A2(pe_1_1_5_n42), .ZN(
        pe_1_1_5_N59) );
  NOR2_X1 pe_1_1_5_U15 ( .A1(pe_1_1_5_n65), .A2(pe_1_1_5_n41), .ZN(
        pe_1_1_5_N60) );
  NOR2_X1 pe_1_1_5_U14 ( .A1(pe_1_1_5_n65), .A2(pe_1_1_5_n38), .ZN(
        pe_1_1_5_N63) );
  NOR2_X1 pe_1_1_5_U13 ( .A1(pe_1_1_5_n65), .A2(pe_1_1_5_n40), .ZN(
        pe_1_1_5_N61) );
  NOR2_X1 pe_1_1_5_U12 ( .A1(pe_1_1_5_n65), .A2(pe_1_1_5_n39), .ZN(
        pe_1_1_5_N62) );
  NOR2_X1 pe_1_1_5_U11 ( .A1(pe_1_1_5_n37), .A2(pe_1_1_5_n65), .ZN(
        pe_1_1_5_N64) );
  NAND2_X1 pe_1_1_5_U10 ( .A1(pe_1_1_5_n44), .A2(n32), .ZN(pe_1_1_5_n42) );
  BUF_X1 pe_1_1_5_U9 ( .A(n32), .Z(pe_1_1_5_n55) );
  INV_X1 pe_1_1_5_U8 ( .A(pe_1_1_5_n66), .ZN(pe_1_1_5_n63) );
  BUF_X1 pe_1_1_5_U7 ( .A(n32), .Z(pe_1_1_5_n56) );
  INV_X1 pe_1_1_5_U6 ( .A(pe_1_1_5_n42), .ZN(pe_1_1_5_n86) );
  INV_X1 pe_1_1_5_U5 ( .A(pe_1_1_5_n40), .ZN(pe_1_1_5_n82) );
  INV_X2 pe_1_1_5_U4 ( .A(n82), .ZN(pe_1_1_5_n69) );
  XOR2_X1 pe_1_1_5_U3 ( .A(pe_1_1_5_int_data_0_), .B(int_data_res_1__5__0_), 
        .Z(pe_1_1_5_n1) );
  DFFR_X1 pe_1_1_5_int_q_acc_reg_0_ ( .D(pe_1_1_5_n81), .CK(pe_1_1_5_net6538), 
        .RN(pe_1_1_5_n69), .Q(int_data_res_1__5__0_), .QN(pe_1_1_5_n3) );
  DFFR_X1 pe_1_1_5_int_q_reg_v_reg_0__0_ ( .D(int_data_y_2__5__0_), .CK(
        pe_1_1_5_net6508), .RN(pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_v[20]) );
  DFFR_X1 pe_1_1_5_int_q_reg_v_reg_0__1_ ( .D(int_data_y_2__5__1_), .CK(
        pe_1_1_5_net6508), .RN(pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_v[21]) );
  DFFR_X1 pe_1_1_5_int_q_reg_v_reg_0__2_ ( .D(int_data_y_2__5__2_), .CK(
        pe_1_1_5_net6508), .RN(pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_v[22]) );
  DFFR_X1 pe_1_1_5_int_q_reg_v_reg_0__3_ ( .D(int_data_y_2__5__3_), .CK(
        pe_1_1_5_net6508), .RN(pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_v[23]) );
  DFFR_X1 pe_1_1_5_int_q_reg_v_reg_1__0_ ( .D(int_data_y_2__5__0_), .CK(
        pe_1_1_5_net6513), .RN(pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_v[16]) );
  DFFR_X1 pe_1_1_5_int_q_reg_v_reg_1__1_ ( .D(int_data_y_2__5__1_), .CK(
        pe_1_1_5_net6513), .RN(pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_v[17]) );
  DFFR_X1 pe_1_1_5_int_q_reg_v_reg_1__2_ ( .D(int_data_y_2__5__2_), .CK(
        pe_1_1_5_net6513), .RN(pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_v[18]) );
  DFFR_X1 pe_1_1_5_int_q_reg_v_reg_1__3_ ( .D(int_data_y_2__5__3_), .CK(
        pe_1_1_5_net6513), .RN(pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_v[19]) );
  DFFR_X1 pe_1_1_5_int_q_reg_v_reg_2__0_ ( .D(int_data_y_2__5__0_), .CK(
        pe_1_1_5_net6518), .RN(pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_v[12]) );
  DFFR_X1 pe_1_1_5_int_q_reg_v_reg_2__1_ ( .D(int_data_y_2__5__1_), .CK(
        pe_1_1_5_net6518), .RN(pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_v[13]) );
  DFFR_X1 pe_1_1_5_int_q_reg_v_reg_2__2_ ( .D(int_data_y_2__5__2_), .CK(
        pe_1_1_5_net6518), .RN(pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_v[14]) );
  DFFR_X1 pe_1_1_5_int_q_reg_v_reg_2__3_ ( .D(int_data_y_2__5__3_), .CK(
        pe_1_1_5_net6518), .RN(pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_v[15]) );
  DFFR_X1 pe_1_1_5_int_q_reg_v_reg_3__0_ ( .D(int_data_y_2__5__0_), .CK(
        pe_1_1_5_net6523), .RN(pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_v[8]) );
  DFFR_X1 pe_1_1_5_int_q_reg_v_reg_3__1_ ( .D(int_data_y_2__5__1_), .CK(
        pe_1_1_5_net6523), .RN(pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_v[9]) );
  DFFR_X1 pe_1_1_5_int_q_reg_v_reg_3__2_ ( .D(int_data_y_2__5__2_), .CK(
        pe_1_1_5_net6523), .RN(pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_v[10]) );
  DFFR_X1 pe_1_1_5_int_q_reg_v_reg_3__3_ ( .D(int_data_y_2__5__3_), .CK(
        pe_1_1_5_net6523), .RN(pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_v[11]) );
  DFFR_X1 pe_1_1_5_int_q_reg_v_reg_4__0_ ( .D(int_data_y_2__5__0_), .CK(
        pe_1_1_5_net6528), .RN(pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_v[4]) );
  DFFR_X1 pe_1_1_5_int_q_reg_v_reg_4__1_ ( .D(int_data_y_2__5__1_), .CK(
        pe_1_1_5_net6528), .RN(pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_v[5]) );
  DFFR_X1 pe_1_1_5_int_q_reg_v_reg_4__2_ ( .D(int_data_y_2__5__2_), .CK(
        pe_1_1_5_net6528), .RN(pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_v[6]) );
  DFFR_X1 pe_1_1_5_int_q_reg_v_reg_4__3_ ( .D(int_data_y_2__5__3_), .CK(
        pe_1_1_5_net6528), .RN(pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_v[7]) );
  DFFR_X1 pe_1_1_5_int_q_reg_v_reg_5__0_ ( .D(int_data_y_2__5__0_), .CK(
        pe_1_1_5_net6533), .RN(pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_v[0]) );
  DFFR_X1 pe_1_1_5_int_q_reg_v_reg_5__1_ ( .D(int_data_y_2__5__1_), .CK(
        pe_1_1_5_net6533), .RN(pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_v[1]) );
  DFFR_X1 pe_1_1_5_int_q_reg_v_reg_5__2_ ( .D(int_data_y_2__5__2_), .CK(
        pe_1_1_5_net6533), .RN(pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_v[2]) );
  DFFR_X1 pe_1_1_5_int_q_reg_v_reg_5__3_ ( .D(int_data_y_2__5__3_), .CK(
        pe_1_1_5_net6533), .RN(pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_1_5_int_q_reg_h_reg_0__0_ ( .D(int_data_x_1__6__0_), .SI(
        int_data_y_2__5__0_), .SE(pe_1_1_5_n63), .CK(pe_1_1_5_net6477), .RN(
        pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_1_5_int_q_reg_h_reg_0__1_ ( .D(int_data_x_1__6__1_), .SI(
        int_data_y_2__5__1_), .SE(pe_1_1_5_n63), .CK(pe_1_1_5_net6477), .RN(
        pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_1_5_int_q_reg_h_reg_0__2_ ( .D(int_data_x_1__6__2_), .SI(
        int_data_y_2__5__2_), .SE(pe_1_1_5_n63), .CK(pe_1_1_5_net6477), .RN(
        pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_1_5_int_q_reg_h_reg_0__3_ ( .D(int_data_x_1__6__3_), .SI(
        int_data_y_2__5__3_), .SE(pe_1_1_5_n63), .CK(pe_1_1_5_net6477), .RN(
        pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_1_5_int_q_reg_h_reg_1__0_ ( .D(int_data_x_1__6__0_), .SI(
        int_data_y_2__5__0_), .SE(pe_1_1_5_n63), .CK(pe_1_1_5_net6483), .RN(
        pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_1_5_int_q_reg_h_reg_1__1_ ( .D(int_data_x_1__6__1_), .SI(
        int_data_y_2__5__1_), .SE(pe_1_1_5_n63), .CK(pe_1_1_5_net6483), .RN(
        pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_1_5_int_q_reg_h_reg_1__2_ ( .D(int_data_x_1__6__2_), .SI(
        int_data_y_2__5__2_), .SE(pe_1_1_5_n63), .CK(pe_1_1_5_net6483), .RN(
        pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_1_5_int_q_reg_h_reg_1__3_ ( .D(int_data_x_1__6__3_), .SI(
        int_data_y_2__5__3_), .SE(pe_1_1_5_n63), .CK(pe_1_1_5_net6483), .RN(
        pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_1_5_int_q_reg_h_reg_2__0_ ( .D(int_data_x_1__6__0_), .SI(
        int_data_y_2__5__0_), .SE(pe_1_1_5_n63), .CK(pe_1_1_5_net6488), .RN(
        pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_1_5_int_q_reg_h_reg_2__1_ ( .D(int_data_x_1__6__1_), .SI(
        int_data_y_2__5__1_), .SE(pe_1_1_5_n63), .CK(pe_1_1_5_net6488), .RN(
        pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_1_5_int_q_reg_h_reg_2__2_ ( .D(int_data_x_1__6__2_), .SI(
        int_data_y_2__5__2_), .SE(pe_1_1_5_n63), .CK(pe_1_1_5_net6488), .RN(
        pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_1_5_int_q_reg_h_reg_2__3_ ( .D(int_data_x_1__6__3_), .SI(
        int_data_y_2__5__3_), .SE(pe_1_1_5_n63), .CK(pe_1_1_5_net6488), .RN(
        pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_1_5_int_q_reg_h_reg_3__0_ ( .D(int_data_x_1__6__0_), .SI(
        int_data_y_2__5__0_), .SE(pe_1_1_5_n63), .CK(pe_1_1_5_net6493), .RN(
        pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_1_5_int_q_reg_h_reg_3__1_ ( .D(int_data_x_1__6__1_), .SI(
        int_data_y_2__5__1_), .SE(pe_1_1_5_n63), .CK(pe_1_1_5_net6493), .RN(
        pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_1_5_int_q_reg_h_reg_3__2_ ( .D(int_data_x_1__6__2_), .SI(
        int_data_y_2__5__2_), .SE(pe_1_1_5_n63), .CK(pe_1_1_5_net6493), .RN(
        pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_1_5_int_q_reg_h_reg_3__3_ ( .D(int_data_x_1__6__3_), .SI(
        int_data_y_2__5__3_), .SE(pe_1_1_5_n63), .CK(pe_1_1_5_net6493), .RN(
        pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_1_5_int_q_reg_h_reg_4__0_ ( .D(int_data_x_1__6__0_), .SI(
        int_data_y_2__5__0_), .SE(pe_1_1_5_n64), .CK(pe_1_1_5_net6498), .RN(
        pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_1_5_int_q_reg_h_reg_4__1_ ( .D(int_data_x_1__6__1_), .SI(
        int_data_y_2__5__1_), .SE(pe_1_1_5_n64), .CK(pe_1_1_5_net6498), .RN(
        pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_1_5_int_q_reg_h_reg_4__2_ ( .D(int_data_x_1__6__2_), .SI(
        int_data_y_2__5__2_), .SE(pe_1_1_5_n64), .CK(pe_1_1_5_net6498), .RN(
        pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_1_5_int_q_reg_h_reg_4__3_ ( .D(int_data_x_1__6__3_), .SI(
        int_data_y_2__5__3_), .SE(pe_1_1_5_n64), .CK(pe_1_1_5_net6498), .RN(
        pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_1_5_int_q_reg_h_reg_5__0_ ( .D(int_data_x_1__6__0_), .SI(
        int_data_y_2__5__0_), .SE(pe_1_1_5_n64), .CK(pe_1_1_5_net6503), .RN(
        pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_1_5_int_q_reg_h_reg_5__1_ ( .D(int_data_x_1__6__1_), .SI(
        int_data_y_2__5__1_), .SE(pe_1_1_5_n64), .CK(pe_1_1_5_net6503), .RN(
        pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_1_5_int_q_reg_h_reg_5__2_ ( .D(int_data_x_1__6__2_), .SI(
        int_data_y_2__5__2_), .SE(pe_1_1_5_n64), .CK(pe_1_1_5_net6503), .RN(
        pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_1_5_int_q_reg_h_reg_5__3_ ( .D(int_data_x_1__6__3_), .SI(
        int_data_y_2__5__3_), .SE(pe_1_1_5_n64), .CK(pe_1_1_5_net6503), .RN(
        pe_1_1_5_n69), .Q(pe_1_1_5_int_q_reg_h[3]) );
  FA_X1 pe_1_1_5_sub_81_U2_7 ( .A(int_data_res_1__5__7_), .B(pe_1_1_5_n73), 
        .CI(pe_1_1_5_sub_81_carry[7]), .S(pe_1_1_5_N77) );
  FA_X1 pe_1_1_5_sub_81_U2_6 ( .A(int_data_res_1__5__6_), .B(pe_1_1_5_n73), 
        .CI(pe_1_1_5_sub_81_carry[6]), .CO(pe_1_1_5_sub_81_carry[7]), .S(
        pe_1_1_5_N76) );
  FA_X1 pe_1_1_5_sub_81_U2_5 ( .A(int_data_res_1__5__5_), .B(pe_1_1_5_n73), 
        .CI(pe_1_1_5_sub_81_carry[5]), .CO(pe_1_1_5_sub_81_carry[6]), .S(
        pe_1_1_5_N75) );
  FA_X1 pe_1_1_5_sub_81_U2_4 ( .A(int_data_res_1__5__4_), .B(pe_1_1_5_n73), 
        .CI(pe_1_1_5_sub_81_carry[4]), .CO(pe_1_1_5_sub_81_carry[5]), .S(
        pe_1_1_5_N74) );
  FA_X1 pe_1_1_5_sub_81_U2_3 ( .A(int_data_res_1__5__3_), .B(pe_1_1_5_n73), 
        .CI(pe_1_1_5_sub_81_carry[3]), .CO(pe_1_1_5_sub_81_carry[4]), .S(
        pe_1_1_5_N73) );
  FA_X1 pe_1_1_5_sub_81_U2_2 ( .A(int_data_res_1__5__2_), .B(pe_1_1_5_n72), 
        .CI(pe_1_1_5_sub_81_carry[2]), .CO(pe_1_1_5_sub_81_carry[3]), .S(
        pe_1_1_5_N72) );
  FA_X1 pe_1_1_5_sub_81_U2_1 ( .A(int_data_res_1__5__1_), .B(pe_1_1_5_n71), 
        .CI(pe_1_1_5_sub_81_carry[1]), .CO(pe_1_1_5_sub_81_carry[2]), .S(
        pe_1_1_5_N71) );
  FA_X1 pe_1_1_5_add_83_U1_7 ( .A(int_data_res_1__5__7_), .B(
        pe_1_1_5_int_data_3_), .CI(pe_1_1_5_add_83_carry[7]), .S(pe_1_1_5_N85)
         );
  FA_X1 pe_1_1_5_add_83_U1_6 ( .A(int_data_res_1__5__6_), .B(
        pe_1_1_5_int_data_3_), .CI(pe_1_1_5_add_83_carry[6]), .CO(
        pe_1_1_5_add_83_carry[7]), .S(pe_1_1_5_N84) );
  FA_X1 pe_1_1_5_add_83_U1_5 ( .A(int_data_res_1__5__5_), .B(
        pe_1_1_5_int_data_3_), .CI(pe_1_1_5_add_83_carry[5]), .CO(
        pe_1_1_5_add_83_carry[6]), .S(pe_1_1_5_N83) );
  FA_X1 pe_1_1_5_add_83_U1_4 ( .A(int_data_res_1__5__4_), .B(
        pe_1_1_5_int_data_3_), .CI(pe_1_1_5_add_83_carry[4]), .CO(
        pe_1_1_5_add_83_carry[5]), .S(pe_1_1_5_N82) );
  FA_X1 pe_1_1_5_add_83_U1_3 ( .A(int_data_res_1__5__3_), .B(
        pe_1_1_5_int_data_3_), .CI(pe_1_1_5_add_83_carry[3]), .CO(
        pe_1_1_5_add_83_carry[4]), .S(pe_1_1_5_N81) );
  FA_X1 pe_1_1_5_add_83_U1_2 ( .A(int_data_res_1__5__2_), .B(
        pe_1_1_5_int_data_2_), .CI(pe_1_1_5_add_83_carry[2]), .CO(
        pe_1_1_5_add_83_carry[3]), .S(pe_1_1_5_N80) );
  FA_X1 pe_1_1_5_add_83_U1_1 ( .A(int_data_res_1__5__1_), .B(
        pe_1_1_5_int_data_1_), .CI(pe_1_1_5_n2), .CO(pe_1_1_5_add_83_carry[2]), 
        .S(pe_1_1_5_N79) );
  NAND3_X1 pe_1_1_5_U56 ( .A1(n32), .A2(pe_1_1_5_n43), .A3(pe_1_1_5_n60), .ZN(
        pe_1_1_5_n40) );
  NAND3_X1 pe_1_1_5_U55 ( .A1(pe_1_1_5_n43), .A2(pe_1_1_5_n59), .A3(
        pe_1_1_5_n60), .ZN(pe_1_1_5_n39) );
  NAND3_X1 pe_1_1_5_U54 ( .A1(pe_1_1_5_n43), .A2(pe_1_1_5_n61), .A3(n32), .ZN(
        pe_1_1_5_n38) );
  NAND3_X1 pe_1_1_5_U53 ( .A1(pe_1_1_5_n59), .A2(pe_1_1_5_n61), .A3(
        pe_1_1_5_n43), .ZN(pe_1_1_5_n37) );
  DFFR_X1 pe_1_1_5_int_q_acc_reg_6_ ( .D(pe_1_1_5_n75), .CK(pe_1_1_5_net6538), 
        .RN(pe_1_1_5_n68), .Q(int_data_res_1__5__6_) );
  DFFR_X1 pe_1_1_5_int_q_acc_reg_5_ ( .D(pe_1_1_5_n76), .CK(pe_1_1_5_net6538), 
        .RN(pe_1_1_5_n68), .Q(int_data_res_1__5__5_) );
  DFFR_X1 pe_1_1_5_int_q_acc_reg_4_ ( .D(pe_1_1_5_n77), .CK(pe_1_1_5_net6538), 
        .RN(pe_1_1_5_n68), .Q(int_data_res_1__5__4_) );
  DFFR_X1 pe_1_1_5_int_q_acc_reg_3_ ( .D(pe_1_1_5_n78), .CK(pe_1_1_5_net6538), 
        .RN(pe_1_1_5_n68), .Q(int_data_res_1__5__3_) );
  DFFR_X1 pe_1_1_5_int_q_acc_reg_2_ ( .D(pe_1_1_5_n79), .CK(pe_1_1_5_net6538), 
        .RN(pe_1_1_5_n68), .Q(int_data_res_1__5__2_) );
  DFFR_X1 pe_1_1_5_int_q_acc_reg_1_ ( .D(pe_1_1_5_n80), .CK(pe_1_1_5_net6538), 
        .RN(pe_1_1_5_n68), .Q(int_data_res_1__5__1_) );
  DFFR_X1 pe_1_1_5_int_q_acc_reg_7_ ( .D(pe_1_1_5_n74), .CK(pe_1_1_5_net6538), 
        .RN(pe_1_1_5_n68), .Q(int_data_res_1__5__7_) );
  CLKGATETST_X1 pe_1_1_5_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_1_5_n85), .SE(1'b0), .GCK(pe_1_1_5_net6477) );
  CLKGATETST_X1 pe_1_1_5_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_1_5_n84), .SE(1'b0), .GCK(pe_1_1_5_net6483) );
  CLKGATETST_X1 pe_1_1_5_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_1_5_n83), .SE(1'b0), .GCK(pe_1_1_5_net6488) );
  CLKGATETST_X1 pe_1_1_5_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_1_5_n82), .SE(1'b0), .GCK(pe_1_1_5_net6493) );
  CLKGATETST_X1 pe_1_1_5_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_1_5_n87), .SE(1'b0), .GCK(pe_1_1_5_net6498) );
  CLKGATETST_X1 pe_1_1_5_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_1_5_n86), .SE(1'b0), .GCK(pe_1_1_5_net6503) );
  CLKGATETST_X1 pe_1_1_5_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_1_5_N64), .SE(1'b0), .GCK(pe_1_1_5_net6508) );
  CLKGATETST_X1 pe_1_1_5_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_1_5_N63), .SE(1'b0), .GCK(pe_1_1_5_net6513) );
  CLKGATETST_X1 pe_1_1_5_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_1_5_N62), .SE(1'b0), .GCK(pe_1_1_5_net6518) );
  CLKGATETST_X1 pe_1_1_5_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_1_5_N61), .SE(1'b0), .GCK(pe_1_1_5_net6523) );
  CLKGATETST_X1 pe_1_1_5_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_1_5_N60), .SE(1'b0), .GCK(pe_1_1_5_net6528) );
  CLKGATETST_X1 pe_1_1_5_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_1_5_N59), .SE(1'b0), .GCK(pe_1_1_5_net6533) );
  CLKGATETST_X1 pe_1_1_5_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_1_5_N90), .SE(1'b0), .GCK(pe_1_1_5_net6538) );
  CLKBUF_X1 pe_1_1_6_U110 ( .A(pe_1_1_6_n70), .Z(pe_1_1_6_n69) );
  INV_X1 pe_1_1_6_U109 ( .A(n74), .ZN(pe_1_1_6_n68) );
  INV_X1 pe_1_1_6_U108 ( .A(n66), .ZN(pe_1_1_6_n67) );
  INV_X1 pe_1_1_6_U107 ( .A(n66), .ZN(pe_1_1_6_n66) );
  INV_X1 pe_1_1_6_U106 ( .A(pe_1_1_6_n67), .ZN(pe_1_1_6_n65) );
  INV_X1 pe_1_1_6_U105 ( .A(pe_1_1_6_n62), .ZN(pe_1_1_6_n61) );
  INV_X1 pe_1_1_6_U104 ( .A(pe_1_1_6_n60), .ZN(pe_1_1_6_n59) );
  INV_X1 pe_1_1_6_U103 ( .A(n26), .ZN(pe_1_1_6_n58) );
  INV_X1 pe_1_1_6_U102 ( .A(n18), .ZN(pe_1_1_6_n57) );
  MUX2_X1 pe_1_1_6_U101 ( .A(pe_1_1_6_n54), .B(pe_1_1_6_n51), .S(n45), .Z(
        int_data_x_1__6__3_) );
  MUX2_X1 pe_1_1_6_U100 ( .A(pe_1_1_6_n53), .B(pe_1_1_6_n52), .S(pe_1_1_6_n61), 
        .Z(pe_1_1_6_n54) );
  MUX2_X1 pe_1_1_6_U99 ( .A(pe_1_1_6_int_q_reg_h[23]), .B(
        pe_1_1_6_int_q_reg_h[19]), .S(pe_1_1_6_n56), .Z(pe_1_1_6_n53) );
  MUX2_X1 pe_1_1_6_U98 ( .A(pe_1_1_6_int_q_reg_h[15]), .B(
        pe_1_1_6_int_q_reg_h[11]), .S(pe_1_1_6_n56), .Z(pe_1_1_6_n52) );
  MUX2_X1 pe_1_1_6_U97 ( .A(pe_1_1_6_int_q_reg_h[7]), .B(
        pe_1_1_6_int_q_reg_h[3]), .S(pe_1_1_6_n56), .Z(pe_1_1_6_n51) );
  MUX2_X1 pe_1_1_6_U96 ( .A(pe_1_1_6_n50), .B(pe_1_1_6_n47), .S(n45), .Z(
        int_data_x_1__6__2_) );
  MUX2_X1 pe_1_1_6_U95 ( .A(pe_1_1_6_n49), .B(pe_1_1_6_n48), .S(pe_1_1_6_n61), 
        .Z(pe_1_1_6_n50) );
  MUX2_X1 pe_1_1_6_U94 ( .A(pe_1_1_6_int_q_reg_h[22]), .B(
        pe_1_1_6_int_q_reg_h[18]), .S(pe_1_1_6_n56), .Z(pe_1_1_6_n49) );
  MUX2_X1 pe_1_1_6_U93 ( .A(pe_1_1_6_int_q_reg_h[14]), .B(
        pe_1_1_6_int_q_reg_h[10]), .S(pe_1_1_6_n56), .Z(pe_1_1_6_n48) );
  MUX2_X1 pe_1_1_6_U92 ( .A(pe_1_1_6_int_q_reg_h[6]), .B(
        pe_1_1_6_int_q_reg_h[2]), .S(pe_1_1_6_n56), .Z(pe_1_1_6_n47) );
  MUX2_X1 pe_1_1_6_U91 ( .A(pe_1_1_6_n46), .B(pe_1_1_6_n24), .S(n45), .Z(
        int_data_x_1__6__1_) );
  MUX2_X1 pe_1_1_6_U90 ( .A(pe_1_1_6_n45), .B(pe_1_1_6_n25), .S(pe_1_1_6_n61), 
        .Z(pe_1_1_6_n46) );
  MUX2_X1 pe_1_1_6_U89 ( .A(pe_1_1_6_int_q_reg_h[21]), .B(
        pe_1_1_6_int_q_reg_h[17]), .S(pe_1_1_6_n56), .Z(pe_1_1_6_n45) );
  MUX2_X1 pe_1_1_6_U88 ( .A(pe_1_1_6_int_q_reg_h[13]), .B(
        pe_1_1_6_int_q_reg_h[9]), .S(pe_1_1_6_n56), .Z(pe_1_1_6_n25) );
  MUX2_X1 pe_1_1_6_U87 ( .A(pe_1_1_6_int_q_reg_h[5]), .B(
        pe_1_1_6_int_q_reg_h[1]), .S(pe_1_1_6_n56), .Z(pe_1_1_6_n24) );
  MUX2_X1 pe_1_1_6_U86 ( .A(pe_1_1_6_n23), .B(pe_1_1_6_n20), .S(n45), .Z(
        int_data_x_1__6__0_) );
  MUX2_X1 pe_1_1_6_U85 ( .A(pe_1_1_6_n22), .B(pe_1_1_6_n21), .S(pe_1_1_6_n61), 
        .Z(pe_1_1_6_n23) );
  MUX2_X1 pe_1_1_6_U84 ( .A(pe_1_1_6_int_q_reg_h[20]), .B(
        pe_1_1_6_int_q_reg_h[16]), .S(pe_1_1_6_n56), .Z(pe_1_1_6_n22) );
  MUX2_X1 pe_1_1_6_U83 ( .A(pe_1_1_6_int_q_reg_h[12]), .B(
        pe_1_1_6_int_q_reg_h[8]), .S(pe_1_1_6_n56), .Z(pe_1_1_6_n21) );
  MUX2_X1 pe_1_1_6_U82 ( .A(pe_1_1_6_int_q_reg_h[4]), .B(
        pe_1_1_6_int_q_reg_h[0]), .S(pe_1_1_6_n56), .Z(pe_1_1_6_n20) );
  MUX2_X1 pe_1_1_6_U81 ( .A(pe_1_1_6_n19), .B(pe_1_1_6_n16), .S(n45), .Z(
        int_data_y_1__6__3_) );
  MUX2_X1 pe_1_1_6_U80 ( .A(pe_1_1_6_n18), .B(pe_1_1_6_n17), .S(pe_1_1_6_n61), 
        .Z(pe_1_1_6_n19) );
  MUX2_X1 pe_1_1_6_U79 ( .A(pe_1_1_6_int_q_reg_v[23]), .B(
        pe_1_1_6_int_q_reg_v[19]), .S(pe_1_1_6_n55), .Z(pe_1_1_6_n18) );
  MUX2_X1 pe_1_1_6_U78 ( .A(pe_1_1_6_int_q_reg_v[15]), .B(
        pe_1_1_6_int_q_reg_v[11]), .S(pe_1_1_6_n55), .Z(pe_1_1_6_n17) );
  MUX2_X1 pe_1_1_6_U77 ( .A(pe_1_1_6_int_q_reg_v[7]), .B(
        pe_1_1_6_int_q_reg_v[3]), .S(pe_1_1_6_n55), .Z(pe_1_1_6_n16) );
  MUX2_X1 pe_1_1_6_U76 ( .A(pe_1_1_6_n15), .B(pe_1_1_6_n12), .S(n45), .Z(
        int_data_y_1__6__2_) );
  MUX2_X1 pe_1_1_6_U75 ( .A(pe_1_1_6_n14), .B(pe_1_1_6_n13), .S(pe_1_1_6_n61), 
        .Z(pe_1_1_6_n15) );
  MUX2_X1 pe_1_1_6_U74 ( .A(pe_1_1_6_int_q_reg_v[22]), .B(
        pe_1_1_6_int_q_reg_v[18]), .S(pe_1_1_6_n55), .Z(pe_1_1_6_n14) );
  MUX2_X1 pe_1_1_6_U73 ( .A(pe_1_1_6_int_q_reg_v[14]), .B(
        pe_1_1_6_int_q_reg_v[10]), .S(pe_1_1_6_n55), .Z(pe_1_1_6_n13) );
  MUX2_X1 pe_1_1_6_U72 ( .A(pe_1_1_6_int_q_reg_v[6]), .B(
        pe_1_1_6_int_q_reg_v[2]), .S(pe_1_1_6_n55), .Z(pe_1_1_6_n12) );
  MUX2_X1 pe_1_1_6_U71 ( .A(pe_1_1_6_n11), .B(pe_1_1_6_n8), .S(n45), .Z(
        int_data_y_1__6__1_) );
  MUX2_X1 pe_1_1_6_U70 ( .A(pe_1_1_6_n10), .B(pe_1_1_6_n9), .S(pe_1_1_6_n61), 
        .Z(pe_1_1_6_n11) );
  MUX2_X1 pe_1_1_6_U69 ( .A(pe_1_1_6_int_q_reg_v[21]), .B(
        pe_1_1_6_int_q_reg_v[17]), .S(pe_1_1_6_n55), .Z(pe_1_1_6_n10) );
  MUX2_X1 pe_1_1_6_U68 ( .A(pe_1_1_6_int_q_reg_v[13]), .B(
        pe_1_1_6_int_q_reg_v[9]), .S(pe_1_1_6_n55), .Z(pe_1_1_6_n9) );
  MUX2_X1 pe_1_1_6_U67 ( .A(pe_1_1_6_int_q_reg_v[5]), .B(
        pe_1_1_6_int_q_reg_v[1]), .S(pe_1_1_6_n55), .Z(pe_1_1_6_n8) );
  MUX2_X1 pe_1_1_6_U66 ( .A(pe_1_1_6_n7), .B(pe_1_1_6_n4), .S(n45), .Z(
        int_data_y_1__6__0_) );
  MUX2_X1 pe_1_1_6_U65 ( .A(pe_1_1_6_n6), .B(pe_1_1_6_n5), .S(pe_1_1_6_n61), 
        .Z(pe_1_1_6_n7) );
  MUX2_X1 pe_1_1_6_U64 ( .A(pe_1_1_6_int_q_reg_v[20]), .B(
        pe_1_1_6_int_q_reg_v[16]), .S(pe_1_1_6_n55), .Z(pe_1_1_6_n6) );
  MUX2_X1 pe_1_1_6_U63 ( .A(pe_1_1_6_int_q_reg_v[12]), .B(
        pe_1_1_6_int_q_reg_v[8]), .S(pe_1_1_6_n55), .Z(pe_1_1_6_n5) );
  MUX2_X1 pe_1_1_6_U62 ( .A(pe_1_1_6_int_q_reg_v[4]), .B(
        pe_1_1_6_int_q_reg_v[0]), .S(pe_1_1_6_n55), .Z(pe_1_1_6_n4) );
  AOI222_X1 pe_1_1_6_U61 ( .A1(int_data_res_2__6__2_), .A2(pe_1_1_6_n63), .B1(
        pe_1_1_6_N80), .B2(pe_1_1_6_n27), .C1(pe_1_1_6_N72), .C2(pe_1_1_6_n28), 
        .ZN(pe_1_1_6_n33) );
  INV_X1 pe_1_1_6_U60 ( .A(pe_1_1_6_n33), .ZN(pe_1_1_6_n80) );
  AOI222_X1 pe_1_1_6_U59 ( .A1(int_data_res_2__6__6_), .A2(pe_1_1_6_n63), .B1(
        pe_1_1_6_N84), .B2(pe_1_1_6_n27), .C1(pe_1_1_6_N76), .C2(pe_1_1_6_n28), 
        .ZN(pe_1_1_6_n29) );
  INV_X1 pe_1_1_6_U58 ( .A(pe_1_1_6_n29), .ZN(pe_1_1_6_n76) );
  XNOR2_X1 pe_1_1_6_U57 ( .A(pe_1_1_6_n71), .B(int_data_res_1__6__0_), .ZN(
        pe_1_1_6_N70) );
  AOI222_X1 pe_1_1_6_U52 ( .A1(int_data_res_2__6__0_), .A2(pe_1_1_6_n63), .B1(
        pe_1_1_6_n1), .B2(pe_1_1_6_n27), .C1(pe_1_1_6_N70), .C2(pe_1_1_6_n28), 
        .ZN(pe_1_1_6_n35) );
  INV_X1 pe_1_1_6_U51 ( .A(pe_1_1_6_n35), .ZN(pe_1_1_6_n82) );
  AOI222_X1 pe_1_1_6_U50 ( .A1(int_data_res_2__6__1_), .A2(pe_1_1_6_n63), .B1(
        pe_1_1_6_N79), .B2(pe_1_1_6_n27), .C1(pe_1_1_6_N71), .C2(pe_1_1_6_n28), 
        .ZN(pe_1_1_6_n34) );
  INV_X1 pe_1_1_6_U49 ( .A(pe_1_1_6_n34), .ZN(pe_1_1_6_n81) );
  AOI222_X1 pe_1_1_6_U48 ( .A1(int_data_res_2__6__3_), .A2(pe_1_1_6_n63), .B1(
        pe_1_1_6_N81), .B2(pe_1_1_6_n27), .C1(pe_1_1_6_N73), .C2(pe_1_1_6_n28), 
        .ZN(pe_1_1_6_n32) );
  INV_X1 pe_1_1_6_U47 ( .A(pe_1_1_6_n32), .ZN(pe_1_1_6_n79) );
  AOI222_X1 pe_1_1_6_U46 ( .A1(int_data_res_2__6__4_), .A2(pe_1_1_6_n63), .B1(
        pe_1_1_6_N82), .B2(pe_1_1_6_n27), .C1(pe_1_1_6_N74), .C2(pe_1_1_6_n28), 
        .ZN(pe_1_1_6_n31) );
  INV_X1 pe_1_1_6_U45 ( .A(pe_1_1_6_n31), .ZN(pe_1_1_6_n78) );
  AOI222_X1 pe_1_1_6_U44 ( .A1(int_data_res_2__6__5_), .A2(pe_1_1_6_n63), .B1(
        pe_1_1_6_N83), .B2(pe_1_1_6_n27), .C1(pe_1_1_6_N75), .C2(pe_1_1_6_n28), 
        .ZN(pe_1_1_6_n30) );
  INV_X1 pe_1_1_6_U43 ( .A(pe_1_1_6_n30), .ZN(pe_1_1_6_n77) );
  NAND2_X1 pe_1_1_6_U42 ( .A1(pe_1_1_6_int_data_0_), .A2(pe_1_1_6_n3), .ZN(
        pe_1_1_6_sub_81_carry[1]) );
  INV_X1 pe_1_1_6_U41 ( .A(pe_1_1_6_int_data_1_), .ZN(pe_1_1_6_n72) );
  INV_X1 pe_1_1_6_U40 ( .A(pe_1_1_6_int_data_2_), .ZN(pe_1_1_6_n73) );
  AND2_X1 pe_1_1_6_U39 ( .A1(pe_1_1_6_int_data_0_), .A2(int_data_res_1__6__0_), 
        .ZN(pe_1_1_6_n2) );
  AOI222_X1 pe_1_1_6_U38 ( .A1(pe_1_1_6_n63), .A2(int_data_res_2__6__7_), .B1(
        pe_1_1_6_N85), .B2(pe_1_1_6_n27), .C1(pe_1_1_6_N77), .C2(pe_1_1_6_n28), 
        .ZN(pe_1_1_6_n26) );
  INV_X1 pe_1_1_6_U37 ( .A(pe_1_1_6_n26), .ZN(pe_1_1_6_n75) );
  NOR3_X1 pe_1_1_6_U36 ( .A1(pe_1_1_6_n58), .A2(pe_1_1_6_n64), .A3(int_ckg[49]), .ZN(pe_1_1_6_n36) );
  OR2_X1 pe_1_1_6_U35 ( .A1(pe_1_1_6_n36), .A2(pe_1_1_6_n63), .ZN(pe_1_1_6_N90) );
  INV_X1 pe_1_1_6_U34 ( .A(n38), .ZN(pe_1_1_6_n62) );
  AND2_X1 pe_1_1_6_U33 ( .A1(int_data_x_1__6__2_), .A2(n26), .ZN(
        pe_1_1_6_int_data_2_) );
  AND2_X1 pe_1_1_6_U32 ( .A1(int_data_x_1__6__1_), .A2(n26), .ZN(
        pe_1_1_6_int_data_1_) );
  AND2_X1 pe_1_1_6_U31 ( .A1(int_data_x_1__6__3_), .A2(n26), .ZN(
        pe_1_1_6_int_data_3_) );
  BUF_X1 pe_1_1_6_U30 ( .A(n60), .Z(pe_1_1_6_n63) );
  INV_X1 pe_1_1_6_U29 ( .A(n32), .ZN(pe_1_1_6_n60) );
  AND2_X1 pe_1_1_6_U28 ( .A1(int_data_x_1__6__0_), .A2(n26), .ZN(
        pe_1_1_6_int_data_0_) );
  NAND2_X1 pe_1_1_6_U27 ( .A1(pe_1_1_6_n44), .A2(pe_1_1_6_n60), .ZN(
        pe_1_1_6_n41) );
  AND3_X1 pe_1_1_6_U26 ( .A1(n74), .A2(pe_1_1_6_n62), .A3(n45), .ZN(
        pe_1_1_6_n44) );
  INV_X1 pe_1_1_6_U25 ( .A(pe_1_1_6_int_data_3_), .ZN(pe_1_1_6_n74) );
  NOR2_X1 pe_1_1_6_U24 ( .A1(pe_1_1_6_n68), .A2(n45), .ZN(pe_1_1_6_n43) );
  NOR2_X1 pe_1_1_6_U23 ( .A1(pe_1_1_6_n57), .A2(pe_1_1_6_n63), .ZN(
        pe_1_1_6_n28) );
  NOR2_X1 pe_1_1_6_U22 ( .A1(n18), .A2(pe_1_1_6_n63), .ZN(pe_1_1_6_n27) );
  INV_X1 pe_1_1_6_U21 ( .A(pe_1_1_6_int_data_0_), .ZN(pe_1_1_6_n71) );
  INV_X1 pe_1_1_6_U20 ( .A(pe_1_1_6_n41), .ZN(pe_1_1_6_n88) );
  INV_X1 pe_1_1_6_U19 ( .A(pe_1_1_6_n37), .ZN(pe_1_1_6_n86) );
  INV_X1 pe_1_1_6_U18 ( .A(pe_1_1_6_n38), .ZN(pe_1_1_6_n85) );
  INV_X1 pe_1_1_6_U17 ( .A(pe_1_1_6_n39), .ZN(pe_1_1_6_n84) );
  NOR2_X1 pe_1_1_6_U16 ( .A1(pe_1_1_6_n66), .A2(pe_1_1_6_n42), .ZN(
        pe_1_1_6_N59) );
  NOR2_X1 pe_1_1_6_U15 ( .A1(pe_1_1_6_n66), .A2(pe_1_1_6_n41), .ZN(
        pe_1_1_6_N60) );
  NOR2_X1 pe_1_1_6_U14 ( .A1(pe_1_1_6_n66), .A2(pe_1_1_6_n38), .ZN(
        pe_1_1_6_N63) );
  NOR2_X1 pe_1_1_6_U13 ( .A1(pe_1_1_6_n66), .A2(pe_1_1_6_n40), .ZN(
        pe_1_1_6_N61) );
  NOR2_X1 pe_1_1_6_U12 ( .A1(pe_1_1_6_n66), .A2(pe_1_1_6_n39), .ZN(
        pe_1_1_6_N62) );
  NOR2_X1 pe_1_1_6_U11 ( .A1(pe_1_1_6_n37), .A2(pe_1_1_6_n66), .ZN(
        pe_1_1_6_N64) );
  NAND2_X1 pe_1_1_6_U10 ( .A1(pe_1_1_6_n44), .A2(pe_1_1_6_n59), .ZN(
        pe_1_1_6_n42) );
  BUF_X1 pe_1_1_6_U9 ( .A(pe_1_1_6_n59), .Z(pe_1_1_6_n55) );
  INV_X1 pe_1_1_6_U8 ( .A(pe_1_1_6_n67), .ZN(pe_1_1_6_n64) );
  BUF_X1 pe_1_1_6_U7 ( .A(pe_1_1_6_n59), .Z(pe_1_1_6_n56) );
  INV_X1 pe_1_1_6_U6 ( .A(pe_1_1_6_n42), .ZN(pe_1_1_6_n87) );
  INV_X1 pe_1_1_6_U5 ( .A(pe_1_1_6_n40), .ZN(pe_1_1_6_n83) );
  INV_X2 pe_1_1_6_U4 ( .A(n82), .ZN(pe_1_1_6_n70) );
  XOR2_X1 pe_1_1_6_U3 ( .A(pe_1_1_6_int_data_0_), .B(int_data_res_1__6__0_), 
        .Z(pe_1_1_6_n1) );
  DFFR_X1 pe_1_1_6_int_q_acc_reg_0_ ( .D(pe_1_1_6_n82), .CK(pe_1_1_6_net6460), 
        .RN(pe_1_1_6_n70), .Q(int_data_res_1__6__0_), .QN(pe_1_1_6_n3) );
  DFFR_X1 pe_1_1_6_int_q_reg_v_reg_0__0_ ( .D(int_data_y_2__6__0_), .CK(
        pe_1_1_6_net6430), .RN(pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_v[20]) );
  DFFR_X1 pe_1_1_6_int_q_reg_v_reg_0__1_ ( .D(int_data_y_2__6__1_), .CK(
        pe_1_1_6_net6430), .RN(pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_v[21]) );
  DFFR_X1 pe_1_1_6_int_q_reg_v_reg_0__2_ ( .D(int_data_y_2__6__2_), .CK(
        pe_1_1_6_net6430), .RN(pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_v[22]) );
  DFFR_X1 pe_1_1_6_int_q_reg_v_reg_0__3_ ( .D(int_data_y_2__6__3_), .CK(
        pe_1_1_6_net6430), .RN(pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_v[23]) );
  DFFR_X1 pe_1_1_6_int_q_reg_v_reg_1__0_ ( .D(int_data_y_2__6__0_), .CK(
        pe_1_1_6_net6435), .RN(pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_v[16]) );
  DFFR_X1 pe_1_1_6_int_q_reg_v_reg_1__1_ ( .D(int_data_y_2__6__1_), .CK(
        pe_1_1_6_net6435), .RN(pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_v[17]) );
  DFFR_X1 pe_1_1_6_int_q_reg_v_reg_1__2_ ( .D(int_data_y_2__6__2_), .CK(
        pe_1_1_6_net6435), .RN(pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_v[18]) );
  DFFR_X1 pe_1_1_6_int_q_reg_v_reg_1__3_ ( .D(int_data_y_2__6__3_), .CK(
        pe_1_1_6_net6435), .RN(pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_v[19]) );
  DFFR_X1 pe_1_1_6_int_q_reg_v_reg_2__0_ ( .D(int_data_y_2__6__0_), .CK(
        pe_1_1_6_net6440), .RN(pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_v[12]) );
  DFFR_X1 pe_1_1_6_int_q_reg_v_reg_2__1_ ( .D(int_data_y_2__6__1_), .CK(
        pe_1_1_6_net6440), .RN(pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_v[13]) );
  DFFR_X1 pe_1_1_6_int_q_reg_v_reg_2__2_ ( .D(int_data_y_2__6__2_), .CK(
        pe_1_1_6_net6440), .RN(pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_v[14]) );
  DFFR_X1 pe_1_1_6_int_q_reg_v_reg_2__3_ ( .D(int_data_y_2__6__3_), .CK(
        pe_1_1_6_net6440), .RN(pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_v[15]) );
  DFFR_X1 pe_1_1_6_int_q_reg_v_reg_3__0_ ( .D(int_data_y_2__6__0_), .CK(
        pe_1_1_6_net6445), .RN(pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_v[8]) );
  DFFR_X1 pe_1_1_6_int_q_reg_v_reg_3__1_ ( .D(int_data_y_2__6__1_), .CK(
        pe_1_1_6_net6445), .RN(pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_v[9]) );
  DFFR_X1 pe_1_1_6_int_q_reg_v_reg_3__2_ ( .D(int_data_y_2__6__2_), .CK(
        pe_1_1_6_net6445), .RN(pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_v[10]) );
  DFFR_X1 pe_1_1_6_int_q_reg_v_reg_3__3_ ( .D(int_data_y_2__6__3_), .CK(
        pe_1_1_6_net6445), .RN(pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_v[11]) );
  DFFR_X1 pe_1_1_6_int_q_reg_v_reg_4__0_ ( .D(int_data_y_2__6__0_), .CK(
        pe_1_1_6_net6450), .RN(pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_v[4]) );
  DFFR_X1 pe_1_1_6_int_q_reg_v_reg_4__1_ ( .D(int_data_y_2__6__1_), .CK(
        pe_1_1_6_net6450), .RN(pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_v[5]) );
  DFFR_X1 pe_1_1_6_int_q_reg_v_reg_4__2_ ( .D(int_data_y_2__6__2_), .CK(
        pe_1_1_6_net6450), .RN(pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_v[6]) );
  DFFR_X1 pe_1_1_6_int_q_reg_v_reg_4__3_ ( .D(int_data_y_2__6__3_), .CK(
        pe_1_1_6_net6450), .RN(pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_v[7]) );
  DFFR_X1 pe_1_1_6_int_q_reg_v_reg_5__0_ ( .D(int_data_y_2__6__0_), .CK(
        pe_1_1_6_net6455), .RN(pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_v[0]) );
  DFFR_X1 pe_1_1_6_int_q_reg_v_reg_5__1_ ( .D(int_data_y_2__6__1_), .CK(
        pe_1_1_6_net6455), .RN(pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_v[1]) );
  DFFR_X1 pe_1_1_6_int_q_reg_v_reg_5__2_ ( .D(int_data_y_2__6__2_), .CK(
        pe_1_1_6_net6455), .RN(pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_v[2]) );
  DFFR_X1 pe_1_1_6_int_q_reg_v_reg_5__3_ ( .D(int_data_y_2__6__3_), .CK(
        pe_1_1_6_net6455), .RN(pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_1_6_int_q_reg_h_reg_0__0_ ( .D(int_data_x_1__7__0_), .SI(
        int_data_y_2__6__0_), .SE(pe_1_1_6_n64), .CK(pe_1_1_6_net6399), .RN(
        pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_1_6_int_q_reg_h_reg_0__1_ ( .D(int_data_x_1__7__1_), .SI(
        int_data_y_2__6__1_), .SE(pe_1_1_6_n64), .CK(pe_1_1_6_net6399), .RN(
        pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_1_6_int_q_reg_h_reg_0__2_ ( .D(int_data_x_1__7__2_), .SI(
        int_data_y_2__6__2_), .SE(pe_1_1_6_n64), .CK(pe_1_1_6_net6399), .RN(
        pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_1_6_int_q_reg_h_reg_0__3_ ( .D(int_data_x_1__7__3_), .SI(
        int_data_y_2__6__3_), .SE(pe_1_1_6_n64), .CK(pe_1_1_6_net6399), .RN(
        pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_1_6_int_q_reg_h_reg_1__0_ ( .D(int_data_x_1__7__0_), .SI(
        int_data_y_2__6__0_), .SE(pe_1_1_6_n64), .CK(pe_1_1_6_net6405), .RN(
        pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_1_6_int_q_reg_h_reg_1__1_ ( .D(int_data_x_1__7__1_), .SI(
        int_data_y_2__6__1_), .SE(pe_1_1_6_n64), .CK(pe_1_1_6_net6405), .RN(
        pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_1_6_int_q_reg_h_reg_1__2_ ( .D(int_data_x_1__7__2_), .SI(
        int_data_y_2__6__2_), .SE(pe_1_1_6_n64), .CK(pe_1_1_6_net6405), .RN(
        pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_1_6_int_q_reg_h_reg_1__3_ ( .D(int_data_x_1__7__3_), .SI(
        int_data_y_2__6__3_), .SE(pe_1_1_6_n64), .CK(pe_1_1_6_net6405), .RN(
        pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_1_6_int_q_reg_h_reg_2__0_ ( .D(int_data_x_1__7__0_), .SI(
        int_data_y_2__6__0_), .SE(pe_1_1_6_n64), .CK(pe_1_1_6_net6410), .RN(
        pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_1_6_int_q_reg_h_reg_2__1_ ( .D(int_data_x_1__7__1_), .SI(
        int_data_y_2__6__1_), .SE(pe_1_1_6_n64), .CK(pe_1_1_6_net6410), .RN(
        pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_1_6_int_q_reg_h_reg_2__2_ ( .D(int_data_x_1__7__2_), .SI(
        int_data_y_2__6__2_), .SE(pe_1_1_6_n64), .CK(pe_1_1_6_net6410), .RN(
        pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_1_6_int_q_reg_h_reg_2__3_ ( .D(int_data_x_1__7__3_), .SI(
        int_data_y_2__6__3_), .SE(pe_1_1_6_n64), .CK(pe_1_1_6_net6410), .RN(
        pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_1_6_int_q_reg_h_reg_3__0_ ( .D(int_data_x_1__7__0_), .SI(
        int_data_y_2__6__0_), .SE(pe_1_1_6_n64), .CK(pe_1_1_6_net6415), .RN(
        pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_1_6_int_q_reg_h_reg_3__1_ ( .D(int_data_x_1__7__1_), .SI(
        int_data_y_2__6__1_), .SE(pe_1_1_6_n64), .CK(pe_1_1_6_net6415), .RN(
        pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_1_6_int_q_reg_h_reg_3__2_ ( .D(int_data_x_1__7__2_), .SI(
        int_data_y_2__6__2_), .SE(pe_1_1_6_n64), .CK(pe_1_1_6_net6415), .RN(
        pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_1_6_int_q_reg_h_reg_3__3_ ( .D(int_data_x_1__7__3_), .SI(
        int_data_y_2__6__3_), .SE(pe_1_1_6_n64), .CK(pe_1_1_6_net6415), .RN(
        pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_1_6_int_q_reg_h_reg_4__0_ ( .D(int_data_x_1__7__0_), .SI(
        int_data_y_2__6__0_), .SE(pe_1_1_6_n65), .CK(pe_1_1_6_net6420), .RN(
        pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_1_6_int_q_reg_h_reg_4__1_ ( .D(int_data_x_1__7__1_), .SI(
        int_data_y_2__6__1_), .SE(pe_1_1_6_n65), .CK(pe_1_1_6_net6420), .RN(
        pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_1_6_int_q_reg_h_reg_4__2_ ( .D(int_data_x_1__7__2_), .SI(
        int_data_y_2__6__2_), .SE(pe_1_1_6_n65), .CK(pe_1_1_6_net6420), .RN(
        pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_1_6_int_q_reg_h_reg_4__3_ ( .D(int_data_x_1__7__3_), .SI(
        int_data_y_2__6__3_), .SE(pe_1_1_6_n65), .CK(pe_1_1_6_net6420), .RN(
        pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_1_6_int_q_reg_h_reg_5__0_ ( .D(int_data_x_1__7__0_), .SI(
        int_data_y_2__6__0_), .SE(pe_1_1_6_n65), .CK(pe_1_1_6_net6425), .RN(
        pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_1_6_int_q_reg_h_reg_5__1_ ( .D(int_data_x_1__7__1_), .SI(
        int_data_y_2__6__1_), .SE(pe_1_1_6_n65), .CK(pe_1_1_6_net6425), .RN(
        pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_1_6_int_q_reg_h_reg_5__2_ ( .D(int_data_x_1__7__2_), .SI(
        int_data_y_2__6__2_), .SE(pe_1_1_6_n65), .CK(pe_1_1_6_net6425), .RN(
        pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_1_6_int_q_reg_h_reg_5__3_ ( .D(int_data_x_1__7__3_), .SI(
        int_data_y_2__6__3_), .SE(pe_1_1_6_n65), .CK(pe_1_1_6_net6425), .RN(
        pe_1_1_6_n70), .Q(pe_1_1_6_int_q_reg_h[3]) );
  FA_X1 pe_1_1_6_sub_81_U2_7 ( .A(int_data_res_1__6__7_), .B(pe_1_1_6_n74), 
        .CI(pe_1_1_6_sub_81_carry[7]), .S(pe_1_1_6_N77) );
  FA_X1 pe_1_1_6_sub_81_U2_6 ( .A(int_data_res_1__6__6_), .B(pe_1_1_6_n74), 
        .CI(pe_1_1_6_sub_81_carry[6]), .CO(pe_1_1_6_sub_81_carry[7]), .S(
        pe_1_1_6_N76) );
  FA_X1 pe_1_1_6_sub_81_U2_5 ( .A(int_data_res_1__6__5_), .B(pe_1_1_6_n74), 
        .CI(pe_1_1_6_sub_81_carry[5]), .CO(pe_1_1_6_sub_81_carry[6]), .S(
        pe_1_1_6_N75) );
  FA_X1 pe_1_1_6_sub_81_U2_4 ( .A(int_data_res_1__6__4_), .B(pe_1_1_6_n74), 
        .CI(pe_1_1_6_sub_81_carry[4]), .CO(pe_1_1_6_sub_81_carry[5]), .S(
        pe_1_1_6_N74) );
  FA_X1 pe_1_1_6_sub_81_U2_3 ( .A(int_data_res_1__6__3_), .B(pe_1_1_6_n74), 
        .CI(pe_1_1_6_sub_81_carry[3]), .CO(pe_1_1_6_sub_81_carry[4]), .S(
        pe_1_1_6_N73) );
  FA_X1 pe_1_1_6_sub_81_U2_2 ( .A(int_data_res_1__6__2_), .B(pe_1_1_6_n73), 
        .CI(pe_1_1_6_sub_81_carry[2]), .CO(pe_1_1_6_sub_81_carry[3]), .S(
        pe_1_1_6_N72) );
  FA_X1 pe_1_1_6_sub_81_U2_1 ( .A(int_data_res_1__6__1_), .B(pe_1_1_6_n72), 
        .CI(pe_1_1_6_sub_81_carry[1]), .CO(pe_1_1_6_sub_81_carry[2]), .S(
        pe_1_1_6_N71) );
  FA_X1 pe_1_1_6_add_83_U1_7 ( .A(int_data_res_1__6__7_), .B(
        pe_1_1_6_int_data_3_), .CI(pe_1_1_6_add_83_carry[7]), .S(pe_1_1_6_N85)
         );
  FA_X1 pe_1_1_6_add_83_U1_6 ( .A(int_data_res_1__6__6_), .B(
        pe_1_1_6_int_data_3_), .CI(pe_1_1_6_add_83_carry[6]), .CO(
        pe_1_1_6_add_83_carry[7]), .S(pe_1_1_6_N84) );
  FA_X1 pe_1_1_6_add_83_U1_5 ( .A(int_data_res_1__6__5_), .B(
        pe_1_1_6_int_data_3_), .CI(pe_1_1_6_add_83_carry[5]), .CO(
        pe_1_1_6_add_83_carry[6]), .S(pe_1_1_6_N83) );
  FA_X1 pe_1_1_6_add_83_U1_4 ( .A(int_data_res_1__6__4_), .B(
        pe_1_1_6_int_data_3_), .CI(pe_1_1_6_add_83_carry[4]), .CO(
        pe_1_1_6_add_83_carry[5]), .S(pe_1_1_6_N82) );
  FA_X1 pe_1_1_6_add_83_U1_3 ( .A(int_data_res_1__6__3_), .B(
        pe_1_1_6_int_data_3_), .CI(pe_1_1_6_add_83_carry[3]), .CO(
        pe_1_1_6_add_83_carry[4]), .S(pe_1_1_6_N81) );
  FA_X1 pe_1_1_6_add_83_U1_2 ( .A(int_data_res_1__6__2_), .B(
        pe_1_1_6_int_data_2_), .CI(pe_1_1_6_add_83_carry[2]), .CO(
        pe_1_1_6_add_83_carry[3]), .S(pe_1_1_6_N80) );
  FA_X1 pe_1_1_6_add_83_U1_1 ( .A(int_data_res_1__6__1_), .B(
        pe_1_1_6_int_data_1_), .CI(pe_1_1_6_n2), .CO(pe_1_1_6_add_83_carry[2]), 
        .S(pe_1_1_6_N79) );
  NAND3_X1 pe_1_1_6_U56 ( .A1(pe_1_1_6_n59), .A2(pe_1_1_6_n43), .A3(
        pe_1_1_6_n61), .ZN(pe_1_1_6_n40) );
  NAND3_X1 pe_1_1_6_U55 ( .A1(pe_1_1_6_n43), .A2(pe_1_1_6_n60), .A3(
        pe_1_1_6_n61), .ZN(pe_1_1_6_n39) );
  NAND3_X1 pe_1_1_6_U54 ( .A1(pe_1_1_6_n43), .A2(pe_1_1_6_n62), .A3(
        pe_1_1_6_n59), .ZN(pe_1_1_6_n38) );
  NAND3_X1 pe_1_1_6_U53 ( .A1(pe_1_1_6_n60), .A2(pe_1_1_6_n62), .A3(
        pe_1_1_6_n43), .ZN(pe_1_1_6_n37) );
  DFFR_X1 pe_1_1_6_int_q_acc_reg_6_ ( .D(pe_1_1_6_n76), .CK(pe_1_1_6_net6460), 
        .RN(pe_1_1_6_n69), .Q(int_data_res_1__6__6_) );
  DFFR_X1 pe_1_1_6_int_q_acc_reg_5_ ( .D(pe_1_1_6_n77), .CK(pe_1_1_6_net6460), 
        .RN(pe_1_1_6_n69), .Q(int_data_res_1__6__5_) );
  DFFR_X1 pe_1_1_6_int_q_acc_reg_4_ ( .D(pe_1_1_6_n78), .CK(pe_1_1_6_net6460), 
        .RN(pe_1_1_6_n69), .Q(int_data_res_1__6__4_) );
  DFFR_X1 pe_1_1_6_int_q_acc_reg_3_ ( .D(pe_1_1_6_n79), .CK(pe_1_1_6_net6460), 
        .RN(pe_1_1_6_n69), .Q(int_data_res_1__6__3_) );
  DFFR_X1 pe_1_1_6_int_q_acc_reg_2_ ( .D(pe_1_1_6_n80), .CK(pe_1_1_6_net6460), 
        .RN(pe_1_1_6_n69), .Q(int_data_res_1__6__2_) );
  DFFR_X1 pe_1_1_6_int_q_acc_reg_1_ ( .D(pe_1_1_6_n81), .CK(pe_1_1_6_net6460), 
        .RN(pe_1_1_6_n69), .Q(int_data_res_1__6__1_) );
  DFFR_X1 pe_1_1_6_int_q_acc_reg_7_ ( .D(pe_1_1_6_n75), .CK(pe_1_1_6_net6460), 
        .RN(pe_1_1_6_n69), .Q(int_data_res_1__6__7_) );
  CLKGATETST_X1 pe_1_1_6_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_1_6_n86), .SE(1'b0), .GCK(pe_1_1_6_net6399) );
  CLKGATETST_X1 pe_1_1_6_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_1_6_n85), .SE(1'b0), .GCK(pe_1_1_6_net6405) );
  CLKGATETST_X1 pe_1_1_6_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_1_6_n84), .SE(1'b0), .GCK(pe_1_1_6_net6410) );
  CLKGATETST_X1 pe_1_1_6_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_1_6_n83), .SE(1'b0), .GCK(pe_1_1_6_net6415) );
  CLKGATETST_X1 pe_1_1_6_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_1_6_n88), .SE(1'b0), .GCK(pe_1_1_6_net6420) );
  CLKGATETST_X1 pe_1_1_6_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_1_6_n87), .SE(1'b0), .GCK(pe_1_1_6_net6425) );
  CLKGATETST_X1 pe_1_1_6_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_1_6_N64), .SE(1'b0), .GCK(pe_1_1_6_net6430) );
  CLKGATETST_X1 pe_1_1_6_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_1_6_N63), .SE(1'b0), .GCK(pe_1_1_6_net6435) );
  CLKGATETST_X1 pe_1_1_6_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_1_6_N62), .SE(1'b0), .GCK(pe_1_1_6_net6440) );
  CLKGATETST_X1 pe_1_1_6_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_1_6_N61), .SE(1'b0), .GCK(pe_1_1_6_net6445) );
  CLKGATETST_X1 pe_1_1_6_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_1_6_N60), .SE(1'b0), .GCK(pe_1_1_6_net6450) );
  CLKGATETST_X1 pe_1_1_6_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_1_6_N59), .SE(1'b0), .GCK(pe_1_1_6_net6455) );
  CLKGATETST_X1 pe_1_1_6_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_1_6_N90), .SE(1'b0), .GCK(pe_1_1_6_net6460) );
  CLKBUF_X1 pe_1_1_7_U110 ( .A(pe_1_1_7_n70), .Z(pe_1_1_7_n69) );
  INV_X1 pe_1_1_7_U109 ( .A(n74), .ZN(pe_1_1_7_n68) );
  INV_X1 pe_1_1_7_U108 ( .A(n66), .ZN(pe_1_1_7_n67) );
  INV_X1 pe_1_1_7_U107 ( .A(n66), .ZN(pe_1_1_7_n66) );
  INV_X1 pe_1_1_7_U106 ( .A(pe_1_1_7_n67), .ZN(pe_1_1_7_n65) );
  INV_X1 pe_1_1_7_U105 ( .A(pe_1_1_7_n62), .ZN(pe_1_1_7_n61) );
  INV_X1 pe_1_1_7_U104 ( .A(pe_1_1_7_n60), .ZN(pe_1_1_7_n59) );
  INV_X1 pe_1_1_7_U103 ( .A(n26), .ZN(pe_1_1_7_n58) );
  INV_X1 pe_1_1_7_U102 ( .A(n18), .ZN(pe_1_1_7_n57) );
  MUX2_X1 pe_1_1_7_U101 ( .A(pe_1_1_7_n54), .B(pe_1_1_7_n51), .S(n46), .Z(
        int_data_x_1__7__3_) );
  MUX2_X1 pe_1_1_7_U100 ( .A(pe_1_1_7_n53), .B(pe_1_1_7_n52), .S(pe_1_1_7_n61), 
        .Z(pe_1_1_7_n54) );
  MUX2_X1 pe_1_1_7_U99 ( .A(pe_1_1_7_int_q_reg_h[23]), .B(
        pe_1_1_7_int_q_reg_h[19]), .S(pe_1_1_7_n56), .Z(pe_1_1_7_n53) );
  MUX2_X1 pe_1_1_7_U98 ( .A(pe_1_1_7_int_q_reg_h[15]), .B(
        pe_1_1_7_int_q_reg_h[11]), .S(pe_1_1_7_n56), .Z(pe_1_1_7_n52) );
  MUX2_X1 pe_1_1_7_U97 ( .A(pe_1_1_7_int_q_reg_h[7]), .B(
        pe_1_1_7_int_q_reg_h[3]), .S(pe_1_1_7_n56), .Z(pe_1_1_7_n51) );
  MUX2_X1 pe_1_1_7_U96 ( .A(pe_1_1_7_n50), .B(pe_1_1_7_n47), .S(n46), .Z(
        int_data_x_1__7__2_) );
  MUX2_X1 pe_1_1_7_U95 ( .A(pe_1_1_7_n49), .B(pe_1_1_7_n48), .S(pe_1_1_7_n61), 
        .Z(pe_1_1_7_n50) );
  MUX2_X1 pe_1_1_7_U94 ( .A(pe_1_1_7_int_q_reg_h[22]), .B(
        pe_1_1_7_int_q_reg_h[18]), .S(pe_1_1_7_n56), .Z(pe_1_1_7_n49) );
  MUX2_X1 pe_1_1_7_U93 ( .A(pe_1_1_7_int_q_reg_h[14]), .B(
        pe_1_1_7_int_q_reg_h[10]), .S(pe_1_1_7_n56), .Z(pe_1_1_7_n48) );
  MUX2_X1 pe_1_1_7_U92 ( .A(pe_1_1_7_int_q_reg_h[6]), .B(
        pe_1_1_7_int_q_reg_h[2]), .S(pe_1_1_7_n56), .Z(pe_1_1_7_n47) );
  MUX2_X1 pe_1_1_7_U91 ( .A(pe_1_1_7_n46), .B(pe_1_1_7_n24), .S(n46), .Z(
        int_data_x_1__7__1_) );
  MUX2_X1 pe_1_1_7_U90 ( .A(pe_1_1_7_n45), .B(pe_1_1_7_n25), .S(pe_1_1_7_n61), 
        .Z(pe_1_1_7_n46) );
  MUX2_X1 pe_1_1_7_U89 ( .A(pe_1_1_7_int_q_reg_h[21]), .B(
        pe_1_1_7_int_q_reg_h[17]), .S(pe_1_1_7_n56), .Z(pe_1_1_7_n45) );
  MUX2_X1 pe_1_1_7_U88 ( .A(pe_1_1_7_int_q_reg_h[13]), .B(
        pe_1_1_7_int_q_reg_h[9]), .S(pe_1_1_7_n56), .Z(pe_1_1_7_n25) );
  MUX2_X1 pe_1_1_7_U87 ( .A(pe_1_1_7_int_q_reg_h[5]), .B(
        pe_1_1_7_int_q_reg_h[1]), .S(pe_1_1_7_n56), .Z(pe_1_1_7_n24) );
  MUX2_X1 pe_1_1_7_U86 ( .A(pe_1_1_7_n23), .B(pe_1_1_7_n20), .S(n46), .Z(
        int_data_x_1__7__0_) );
  MUX2_X1 pe_1_1_7_U85 ( .A(pe_1_1_7_n22), .B(pe_1_1_7_n21), .S(pe_1_1_7_n61), 
        .Z(pe_1_1_7_n23) );
  MUX2_X1 pe_1_1_7_U84 ( .A(pe_1_1_7_int_q_reg_h[20]), .B(
        pe_1_1_7_int_q_reg_h[16]), .S(pe_1_1_7_n56), .Z(pe_1_1_7_n22) );
  MUX2_X1 pe_1_1_7_U83 ( .A(pe_1_1_7_int_q_reg_h[12]), .B(
        pe_1_1_7_int_q_reg_h[8]), .S(pe_1_1_7_n56), .Z(pe_1_1_7_n21) );
  MUX2_X1 pe_1_1_7_U82 ( .A(pe_1_1_7_int_q_reg_h[4]), .B(
        pe_1_1_7_int_q_reg_h[0]), .S(pe_1_1_7_n56), .Z(pe_1_1_7_n20) );
  MUX2_X1 pe_1_1_7_U81 ( .A(pe_1_1_7_n19), .B(pe_1_1_7_n16), .S(n46), .Z(
        int_data_y_1__7__3_) );
  MUX2_X1 pe_1_1_7_U80 ( .A(pe_1_1_7_n18), .B(pe_1_1_7_n17), .S(pe_1_1_7_n61), 
        .Z(pe_1_1_7_n19) );
  MUX2_X1 pe_1_1_7_U79 ( .A(pe_1_1_7_int_q_reg_v[23]), .B(
        pe_1_1_7_int_q_reg_v[19]), .S(pe_1_1_7_n55), .Z(pe_1_1_7_n18) );
  MUX2_X1 pe_1_1_7_U78 ( .A(pe_1_1_7_int_q_reg_v[15]), .B(
        pe_1_1_7_int_q_reg_v[11]), .S(pe_1_1_7_n55), .Z(pe_1_1_7_n17) );
  MUX2_X1 pe_1_1_7_U77 ( .A(pe_1_1_7_int_q_reg_v[7]), .B(
        pe_1_1_7_int_q_reg_v[3]), .S(pe_1_1_7_n55), .Z(pe_1_1_7_n16) );
  MUX2_X1 pe_1_1_7_U76 ( .A(pe_1_1_7_n15), .B(pe_1_1_7_n12), .S(n46), .Z(
        int_data_y_1__7__2_) );
  MUX2_X1 pe_1_1_7_U75 ( .A(pe_1_1_7_n14), .B(pe_1_1_7_n13), .S(pe_1_1_7_n61), 
        .Z(pe_1_1_7_n15) );
  MUX2_X1 pe_1_1_7_U74 ( .A(pe_1_1_7_int_q_reg_v[22]), .B(
        pe_1_1_7_int_q_reg_v[18]), .S(pe_1_1_7_n55), .Z(pe_1_1_7_n14) );
  MUX2_X1 pe_1_1_7_U73 ( .A(pe_1_1_7_int_q_reg_v[14]), .B(
        pe_1_1_7_int_q_reg_v[10]), .S(pe_1_1_7_n55), .Z(pe_1_1_7_n13) );
  MUX2_X1 pe_1_1_7_U72 ( .A(pe_1_1_7_int_q_reg_v[6]), .B(
        pe_1_1_7_int_q_reg_v[2]), .S(pe_1_1_7_n55), .Z(pe_1_1_7_n12) );
  MUX2_X1 pe_1_1_7_U71 ( .A(pe_1_1_7_n11), .B(pe_1_1_7_n8), .S(n46), .Z(
        int_data_y_1__7__1_) );
  MUX2_X1 pe_1_1_7_U70 ( .A(pe_1_1_7_n10), .B(pe_1_1_7_n9), .S(pe_1_1_7_n61), 
        .Z(pe_1_1_7_n11) );
  MUX2_X1 pe_1_1_7_U69 ( .A(pe_1_1_7_int_q_reg_v[21]), .B(
        pe_1_1_7_int_q_reg_v[17]), .S(pe_1_1_7_n55), .Z(pe_1_1_7_n10) );
  MUX2_X1 pe_1_1_7_U68 ( .A(pe_1_1_7_int_q_reg_v[13]), .B(
        pe_1_1_7_int_q_reg_v[9]), .S(pe_1_1_7_n55), .Z(pe_1_1_7_n9) );
  MUX2_X1 pe_1_1_7_U67 ( .A(pe_1_1_7_int_q_reg_v[5]), .B(
        pe_1_1_7_int_q_reg_v[1]), .S(pe_1_1_7_n55), .Z(pe_1_1_7_n8) );
  MUX2_X1 pe_1_1_7_U66 ( .A(pe_1_1_7_n7), .B(pe_1_1_7_n4), .S(n46), .Z(
        int_data_y_1__7__0_) );
  MUX2_X1 pe_1_1_7_U65 ( .A(pe_1_1_7_n6), .B(pe_1_1_7_n5), .S(pe_1_1_7_n61), 
        .Z(pe_1_1_7_n7) );
  MUX2_X1 pe_1_1_7_U64 ( .A(pe_1_1_7_int_q_reg_v[20]), .B(
        pe_1_1_7_int_q_reg_v[16]), .S(pe_1_1_7_n55), .Z(pe_1_1_7_n6) );
  MUX2_X1 pe_1_1_7_U63 ( .A(pe_1_1_7_int_q_reg_v[12]), .B(
        pe_1_1_7_int_q_reg_v[8]), .S(pe_1_1_7_n55), .Z(pe_1_1_7_n5) );
  MUX2_X1 pe_1_1_7_U62 ( .A(pe_1_1_7_int_q_reg_v[4]), .B(
        pe_1_1_7_int_q_reg_v[0]), .S(pe_1_1_7_n55), .Z(pe_1_1_7_n4) );
  AOI222_X1 pe_1_1_7_U61 ( .A1(int_data_res_2__7__2_), .A2(pe_1_1_7_n63), .B1(
        pe_1_1_7_N80), .B2(pe_1_1_7_n27), .C1(pe_1_1_7_N72), .C2(pe_1_1_7_n28), 
        .ZN(pe_1_1_7_n33) );
  INV_X1 pe_1_1_7_U60 ( .A(pe_1_1_7_n33), .ZN(pe_1_1_7_n80) );
  AOI222_X1 pe_1_1_7_U59 ( .A1(int_data_res_2__7__6_), .A2(pe_1_1_7_n63), .B1(
        pe_1_1_7_N84), .B2(pe_1_1_7_n27), .C1(pe_1_1_7_N76), .C2(pe_1_1_7_n28), 
        .ZN(pe_1_1_7_n29) );
  INV_X1 pe_1_1_7_U58 ( .A(pe_1_1_7_n29), .ZN(pe_1_1_7_n76) );
  XNOR2_X1 pe_1_1_7_U57 ( .A(pe_1_1_7_n71), .B(int_data_res_1__7__0_), .ZN(
        pe_1_1_7_N70) );
  AOI222_X1 pe_1_1_7_U52 ( .A1(int_data_res_2__7__0_), .A2(pe_1_1_7_n63), .B1(
        pe_1_1_7_n1), .B2(pe_1_1_7_n27), .C1(pe_1_1_7_N70), .C2(pe_1_1_7_n28), 
        .ZN(pe_1_1_7_n35) );
  INV_X1 pe_1_1_7_U51 ( .A(pe_1_1_7_n35), .ZN(pe_1_1_7_n82) );
  AOI222_X1 pe_1_1_7_U50 ( .A1(int_data_res_2__7__1_), .A2(pe_1_1_7_n63), .B1(
        pe_1_1_7_N79), .B2(pe_1_1_7_n27), .C1(pe_1_1_7_N71), .C2(pe_1_1_7_n28), 
        .ZN(pe_1_1_7_n34) );
  INV_X1 pe_1_1_7_U49 ( .A(pe_1_1_7_n34), .ZN(pe_1_1_7_n81) );
  AOI222_X1 pe_1_1_7_U48 ( .A1(int_data_res_2__7__3_), .A2(pe_1_1_7_n63), .B1(
        pe_1_1_7_N81), .B2(pe_1_1_7_n27), .C1(pe_1_1_7_N73), .C2(pe_1_1_7_n28), 
        .ZN(pe_1_1_7_n32) );
  INV_X1 pe_1_1_7_U47 ( .A(pe_1_1_7_n32), .ZN(pe_1_1_7_n79) );
  AOI222_X1 pe_1_1_7_U46 ( .A1(int_data_res_2__7__4_), .A2(pe_1_1_7_n63), .B1(
        pe_1_1_7_N82), .B2(pe_1_1_7_n27), .C1(pe_1_1_7_N74), .C2(pe_1_1_7_n28), 
        .ZN(pe_1_1_7_n31) );
  INV_X1 pe_1_1_7_U45 ( .A(pe_1_1_7_n31), .ZN(pe_1_1_7_n78) );
  AOI222_X1 pe_1_1_7_U44 ( .A1(int_data_res_2__7__5_), .A2(pe_1_1_7_n63), .B1(
        pe_1_1_7_N83), .B2(pe_1_1_7_n27), .C1(pe_1_1_7_N75), .C2(pe_1_1_7_n28), 
        .ZN(pe_1_1_7_n30) );
  INV_X1 pe_1_1_7_U43 ( .A(pe_1_1_7_n30), .ZN(pe_1_1_7_n77) );
  NAND2_X1 pe_1_1_7_U42 ( .A1(pe_1_1_7_int_data_0_), .A2(pe_1_1_7_n3), .ZN(
        pe_1_1_7_sub_81_carry[1]) );
  INV_X1 pe_1_1_7_U41 ( .A(pe_1_1_7_int_data_1_), .ZN(pe_1_1_7_n72) );
  INV_X1 pe_1_1_7_U40 ( .A(pe_1_1_7_int_data_2_), .ZN(pe_1_1_7_n73) );
  AND2_X1 pe_1_1_7_U39 ( .A1(pe_1_1_7_int_data_0_), .A2(int_data_res_1__7__0_), 
        .ZN(pe_1_1_7_n2) );
  AOI222_X1 pe_1_1_7_U38 ( .A1(pe_1_1_7_n63), .A2(int_data_res_2__7__7_), .B1(
        pe_1_1_7_N85), .B2(pe_1_1_7_n27), .C1(pe_1_1_7_N77), .C2(pe_1_1_7_n28), 
        .ZN(pe_1_1_7_n26) );
  INV_X1 pe_1_1_7_U37 ( .A(pe_1_1_7_n26), .ZN(pe_1_1_7_n75) );
  NOR3_X1 pe_1_1_7_U36 ( .A1(pe_1_1_7_n58), .A2(pe_1_1_7_n64), .A3(int_ckg[48]), .ZN(pe_1_1_7_n36) );
  OR2_X1 pe_1_1_7_U35 ( .A1(pe_1_1_7_n36), .A2(pe_1_1_7_n63), .ZN(pe_1_1_7_N90) );
  INV_X1 pe_1_1_7_U34 ( .A(n38), .ZN(pe_1_1_7_n62) );
  AND2_X1 pe_1_1_7_U33 ( .A1(int_data_x_1__7__2_), .A2(n26), .ZN(
        pe_1_1_7_int_data_2_) );
  AND2_X1 pe_1_1_7_U32 ( .A1(int_data_x_1__7__1_), .A2(n26), .ZN(
        pe_1_1_7_int_data_1_) );
  AND2_X1 pe_1_1_7_U31 ( .A1(int_data_x_1__7__3_), .A2(n26), .ZN(
        pe_1_1_7_int_data_3_) );
  BUF_X1 pe_1_1_7_U30 ( .A(n60), .Z(pe_1_1_7_n63) );
  INV_X1 pe_1_1_7_U29 ( .A(n32), .ZN(pe_1_1_7_n60) );
  AND2_X1 pe_1_1_7_U28 ( .A1(int_data_x_1__7__0_), .A2(n26), .ZN(
        pe_1_1_7_int_data_0_) );
  NAND2_X1 pe_1_1_7_U27 ( .A1(pe_1_1_7_n44), .A2(pe_1_1_7_n60), .ZN(
        pe_1_1_7_n41) );
  AND3_X1 pe_1_1_7_U26 ( .A1(n74), .A2(pe_1_1_7_n62), .A3(n46), .ZN(
        pe_1_1_7_n44) );
  INV_X1 pe_1_1_7_U25 ( .A(pe_1_1_7_int_data_3_), .ZN(pe_1_1_7_n74) );
  NOR2_X1 pe_1_1_7_U24 ( .A1(pe_1_1_7_n68), .A2(n46), .ZN(pe_1_1_7_n43) );
  NOR2_X1 pe_1_1_7_U23 ( .A1(pe_1_1_7_n57), .A2(pe_1_1_7_n63), .ZN(
        pe_1_1_7_n28) );
  NOR2_X1 pe_1_1_7_U22 ( .A1(n18), .A2(pe_1_1_7_n63), .ZN(pe_1_1_7_n27) );
  INV_X1 pe_1_1_7_U21 ( .A(pe_1_1_7_int_data_0_), .ZN(pe_1_1_7_n71) );
  INV_X1 pe_1_1_7_U20 ( .A(pe_1_1_7_n41), .ZN(pe_1_1_7_n88) );
  INV_X1 pe_1_1_7_U19 ( .A(pe_1_1_7_n37), .ZN(pe_1_1_7_n86) );
  INV_X1 pe_1_1_7_U18 ( .A(pe_1_1_7_n38), .ZN(pe_1_1_7_n85) );
  INV_X1 pe_1_1_7_U17 ( .A(pe_1_1_7_n39), .ZN(pe_1_1_7_n84) );
  NOR2_X1 pe_1_1_7_U16 ( .A1(pe_1_1_7_n66), .A2(pe_1_1_7_n42), .ZN(
        pe_1_1_7_N59) );
  NOR2_X1 pe_1_1_7_U15 ( .A1(pe_1_1_7_n66), .A2(pe_1_1_7_n41), .ZN(
        pe_1_1_7_N60) );
  NOR2_X1 pe_1_1_7_U14 ( .A1(pe_1_1_7_n66), .A2(pe_1_1_7_n38), .ZN(
        pe_1_1_7_N63) );
  NOR2_X1 pe_1_1_7_U13 ( .A1(pe_1_1_7_n66), .A2(pe_1_1_7_n40), .ZN(
        pe_1_1_7_N61) );
  NOR2_X1 pe_1_1_7_U12 ( .A1(pe_1_1_7_n66), .A2(pe_1_1_7_n39), .ZN(
        pe_1_1_7_N62) );
  NOR2_X1 pe_1_1_7_U11 ( .A1(pe_1_1_7_n37), .A2(pe_1_1_7_n66), .ZN(
        pe_1_1_7_N64) );
  NAND2_X1 pe_1_1_7_U10 ( .A1(pe_1_1_7_n44), .A2(pe_1_1_7_n59), .ZN(
        pe_1_1_7_n42) );
  BUF_X1 pe_1_1_7_U9 ( .A(pe_1_1_7_n59), .Z(pe_1_1_7_n55) );
  INV_X1 pe_1_1_7_U8 ( .A(pe_1_1_7_n67), .ZN(pe_1_1_7_n64) );
  BUF_X1 pe_1_1_7_U7 ( .A(pe_1_1_7_n59), .Z(pe_1_1_7_n56) );
  INV_X1 pe_1_1_7_U6 ( .A(pe_1_1_7_n42), .ZN(pe_1_1_7_n87) );
  INV_X1 pe_1_1_7_U5 ( .A(pe_1_1_7_n40), .ZN(pe_1_1_7_n83) );
  INV_X2 pe_1_1_7_U4 ( .A(n82), .ZN(pe_1_1_7_n70) );
  XOR2_X1 pe_1_1_7_U3 ( .A(pe_1_1_7_int_data_0_), .B(int_data_res_1__7__0_), 
        .Z(pe_1_1_7_n1) );
  DFFR_X1 pe_1_1_7_int_q_acc_reg_0_ ( .D(pe_1_1_7_n82), .CK(pe_1_1_7_net6382), 
        .RN(pe_1_1_7_n70), .Q(int_data_res_1__7__0_), .QN(pe_1_1_7_n3) );
  DFFR_X1 pe_1_1_7_int_q_reg_v_reg_0__0_ ( .D(int_data_y_2__7__0_), .CK(
        pe_1_1_7_net6352), .RN(pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_v[20]) );
  DFFR_X1 pe_1_1_7_int_q_reg_v_reg_0__1_ ( .D(int_data_y_2__7__1_), .CK(
        pe_1_1_7_net6352), .RN(pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_v[21]) );
  DFFR_X1 pe_1_1_7_int_q_reg_v_reg_0__2_ ( .D(int_data_y_2__7__2_), .CK(
        pe_1_1_7_net6352), .RN(pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_v[22]) );
  DFFR_X1 pe_1_1_7_int_q_reg_v_reg_0__3_ ( .D(int_data_y_2__7__3_), .CK(
        pe_1_1_7_net6352), .RN(pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_v[23]) );
  DFFR_X1 pe_1_1_7_int_q_reg_v_reg_1__0_ ( .D(int_data_y_2__7__0_), .CK(
        pe_1_1_7_net6357), .RN(pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_v[16]) );
  DFFR_X1 pe_1_1_7_int_q_reg_v_reg_1__1_ ( .D(int_data_y_2__7__1_), .CK(
        pe_1_1_7_net6357), .RN(pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_v[17]) );
  DFFR_X1 pe_1_1_7_int_q_reg_v_reg_1__2_ ( .D(int_data_y_2__7__2_), .CK(
        pe_1_1_7_net6357), .RN(pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_v[18]) );
  DFFR_X1 pe_1_1_7_int_q_reg_v_reg_1__3_ ( .D(int_data_y_2__7__3_), .CK(
        pe_1_1_7_net6357), .RN(pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_v[19]) );
  DFFR_X1 pe_1_1_7_int_q_reg_v_reg_2__0_ ( .D(int_data_y_2__7__0_), .CK(
        pe_1_1_7_net6362), .RN(pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_v[12]) );
  DFFR_X1 pe_1_1_7_int_q_reg_v_reg_2__1_ ( .D(int_data_y_2__7__1_), .CK(
        pe_1_1_7_net6362), .RN(pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_v[13]) );
  DFFR_X1 pe_1_1_7_int_q_reg_v_reg_2__2_ ( .D(int_data_y_2__7__2_), .CK(
        pe_1_1_7_net6362), .RN(pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_v[14]) );
  DFFR_X1 pe_1_1_7_int_q_reg_v_reg_2__3_ ( .D(int_data_y_2__7__3_), .CK(
        pe_1_1_7_net6362), .RN(pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_v[15]) );
  DFFR_X1 pe_1_1_7_int_q_reg_v_reg_3__0_ ( .D(int_data_y_2__7__0_), .CK(
        pe_1_1_7_net6367), .RN(pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_v[8]) );
  DFFR_X1 pe_1_1_7_int_q_reg_v_reg_3__1_ ( .D(int_data_y_2__7__1_), .CK(
        pe_1_1_7_net6367), .RN(pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_v[9]) );
  DFFR_X1 pe_1_1_7_int_q_reg_v_reg_3__2_ ( .D(int_data_y_2__7__2_), .CK(
        pe_1_1_7_net6367), .RN(pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_v[10]) );
  DFFR_X1 pe_1_1_7_int_q_reg_v_reg_3__3_ ( .D(int_data_y_2__7__3_), .CK(
        pe_1_1_7_net6367), .RN(pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_v[11]) );
  DFFR_X1 pe_1_1_7_int_q_reg_v_reg_4__0_ ( .D(int_data_y_2__7__0_), .CK(
        pe_1_1_7_net6372), .RN(pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_v[4]) );
  DFFR_X1 pe_1_1_7_int_q_reg_v_reg_4__1_ ( .D(int_data_y_2__7__1_), .CK(
        pe_1_1_7_net6372), .RN(pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_v[5]) );
  DFFR_X1 pe_1_1_7_int_q_reg_v_reg_4__2_ ( .D(int_data_y_2__7__2_), .CK(
        pe_1_1_7_net6372), .RN(pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_v[6]) );
  DFFR_X1 pe_1_1_7_int_q_reg_v_reg_4__3_ ( .D(int_data_y_2__7__3_), .CK(
        pe_1_1_7_net6372), .RN(pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_v[7]) );
  DFFR_X1 pe_1_1_7_int_q_reg_v_reg_5__0_ ( .D(int_data_y_2__7__0_), .CK(
        pe_1_1_7_net6377), .RN(pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_v[0]) );
  DFFR_X1 pe_1_1_7_int_q_reg_v_reg_5__1_ ( .D(int_data_y_2__7__1_), .CK(
        pe_1_1_7_net6377), .RN(pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_v[1]) );
  DFFR_X1 pe_1_1_7_int_q_reg_v_reg_5__2_ ( .D(int_data_y_2__7__2_), .CK(
        pe_1_1_7_net6377), .RN(pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_v[2]) );
  DFFR_X1 pe_1_1_7_int_q_reg_v_reg_5__3_ ( .D(int_data_y_2__7__3_), .CK(
        pe_1_1_7_net6377), .RN(pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_1_7_int_q_reg_h_reg_0__0_ ( .D(i_data_conv_h[24]), .SI(
        int_data_y_2__7__0_), .SE(pe_1_1_7_n64), .CK(pe_1_1_7_net6321), .RN(
        pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_1_7_int_q_reg_h_reg_0__1_ ( .D(i_data_conv_h[25]), .SI(
        int_data_y_2__7__1_), .SE(pe_1_1_7_n64), .CK(pe_1_1_7_net6321), .RN(
        pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_1_7_int_q_reg_h_reg_0__2_ ( .D(i_data_conv_h[26]), .SI(
        int_data_y_2__7__2_), .SE(pe_1_1_7_n64), .CK(pe_1_1_7_net6321), .RN(
        pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_1_7_int_q_reg_h_reg_0__3_ ( .D(i_data_conv_h[27]), .SI(
        int_data_y_2__7__3_), .SE(pe_1_1_7_n64), .CK(pe_1_1_7_net6321), .RN(
        pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_1_7_int_q_reg_h_reg_1__0_ ( .D(i_data_conv_h[24]), .SI(
        int_data_y_2__7__0_), .SE(pe_1_1_7_n64), .CK(pe_1_1_7_net6327), .RN(
        pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_1_7_int_q_reg_h_reg_1__1_ ( .D(i_data_conv_h[25]), .SI(
        int_data_y_2__7__1_), .SE(pe_1_1_7_n64), .CK(pe_1_1_7_net6327), .RN(
        pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_1_7_int_q_reg_h_reg_1__2_ ( .D(i_data_conv_h[26]), .SI(
        int_data_y_2__7__2_), .SE(pe_1_1_7_n64), .CK(pe_1_1_7_net6327), .RN(
        pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_1_7_int_q_reg_h_reg_1__3_ ( .D(i_data_conv_h[27]), .SI(
        int_data_y_2__7__3_), .SE(pe_1_1_7_n64), .CK(pe_1_1_7_net6327), .RN(
        pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_1_7_int_q_reg_h_reg_2__0_ ( .D(i_data_conv_h[24]), .SI(
        int_data_y_2__7__0_), .SE(pe_1_1_7_n64), .CK(pe_1_1_7_net6332), .RN(
        pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_1_7_int_q_reg_h_reg_2__1_ ( .D(i_data_conv_h[25]), .SI(
        int_data_y_2__7__1_), .SE(pe_1_1_7_n64), .CK(pe_1_1_7_net6332), .RN(
        pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_1_7_int_q_reg_h_reg_2__2_ ( .D(i_data_conv_h[26]), .SI(
        int_data_y_2__7__2_), .SE(pe_1_1_7_n64), .CK(pe_1_1_7_net6332), .RN(
        pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_1_7_int_q_reg_h_reg_2__3_ ( .D(i_data_conv_h[27]), .SI(
        int_data_y_2__7__3_), .SE(pe_1_1_7_n64), .CK(pe_1_1_7_net6332), .RN(
        pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_1_7_int_q_reg_h_reg_3__0_ ( .D(i_data_conv_h[24]), .SI(
        int_data_y_2__7__0_), .SE(pe_1_1_7_n64), .CK(pe_1_1_7_net6337), .RN(
        pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_1_7_int_q_reg_h_reg_3__1_ ( .D(i_data_conv_h[25]), .SI(
        int_data_y_2__7__1_), .SE(pe_1_1_7_n64), .CK(pe_1_1_7_net6337), .RN(
        pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_1_7_int_q_reg_h_reg_3__2_ ( .D(i_data_conv_h[26]), .SI(
        int_data_y_2__7__2_), .SE(pe_1_1_7_n64), .CK(pe_1_1_7_net6337), .RN(
        pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_1_7_int_q_reg_h_reg_3__3_ ( .D(i_data_conv_h[27]), .SI(
        int_data_y_2__7__3_), .SE(pe_1_1_7_n64), .CK(pe_1_1_7_net6337), .RN(
        pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_1_7_int_q_reg_h_reg_4__0_ ( .D(i_data_conv_h[24]), .SI(
        int_data_y_2__7__0_), .SE(pe_1_1_7_n65), .CK(pe_1_1_7_net6342), .RN(
        pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_1_7_int_q_reg_h_reg_4__1_ ( .D(i_data_conv_h[25]), .SI(
        int_data_y_2__7__1_), .SE(pe_1_1_7_n65), .CK(pe_1_1_7_net6342), .RN(
        pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_1_7_int_q_reg_h_reg_4__2_ ( .D(i_data_conv_h[26]), .SI(
        int_data_y_2__7__2_), .SE(pe_1_1_7_n65), .CK(pe_1_1_7_net6342), .RN(
        pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_1_7_int_q_reg_h_reg_4__3_ ( .D(i_data_conv_h[27]), .SI(
        int_data_y_2__7__3_), .SE(pe_1_1_7_n65), .CK(pe_1_1_7_net6342), .RN(
        pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_1_7_int_q_reg_h_reg_5__0_ ( .D(i_data_conv_h[24]), .SI(
        int_data_y_2__7__0_), .SE(pe_1_1_7_n65), .CK(pe_1_1_7_net6347), .RN(
        pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_1_7_int_q_reg_h_reg_5__1_ ( .D(i_data_conv_h[25]), .SI(
        int_data_y_2__7__1_), .SE(pe_1_1_7_n65), .CK(pe_1_1_7_net6347), .RN(
        pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_1_7_int_q_reg_h_reg_5__2_ ( .D(i_data_conv_h[26]), .SI(
        int_data_y_2__7__2_), .SE(pe_1_1_7_n65), .CK(pe_1_1_7_net6347), .RN(
        pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_1_7_int_q_reg_h_reg_5__3_ ( .D(i_data_conv_h[27]), .SI(
        int_data_y_2__7__3_), .SE(pe_1_1_7_n65), .CK(pe_1_1_7_net6347), .RN(
        pe_1_1_7_n70), .Q(pe_1_1_7_int_q_reg_h[3]) );
  FA_X1 pe_1_1_7_sub_81_U2_7 ( .A(int_data_res_1__7__7_), .B(pe_1_1_7_n74), 
        .CI(pe_1_1_7_sub_81_carry[7]), .S(pe_1_1_7_N77) );
  FA_X1 pe_1_1_7_sub_81_U2_6 ( .A(int_data_res_1__7__6_), .B(pe_1_1_7_n74), 
        .CI(pe_1_1_7_sub_81_carry[6]), .CO(pe_1_1_7_sub_81_carry[7]), .S(
        pe_1_1_7_N76) );
  FA_X1 pe_1_1_7_sub_81_U2_5 ( .A(int_data_res_1__7__5_), .B(pe_1_1_7_n74), 
        .CI(pe_1_1_7_sub_81_carry[5]), .CO(pe_1_1_7_sub_81_carry[6]), .S(
        pe_1_1_7_N75) );
  FA_X1 pe_1_1_7_sub_81_U2_4 ( .A(int_data_res_1__7__4_), .B(pe_1_1_7_n74), 
        .CI(pe_1_1_7_sub_81_carry[4]), .CO(pe_1_1_7_sub_81_carry[5]), .S(
        pe_1_1_7_N74) );
  FA_X1 pe_1_1_7_sub_81_U2_3 ( .A(int_data_res_1__7__3_), .B(pe_1_1_7_n74), 
        .CI(pe_1_1_7_sub_81_carry[3]), .CO(pe_1_1_7_sub_81_carry[4]), .S(
        pe_1_1_7_N73) );
  FA_X1 pe_1_1_7_sub_81_U2_2 ( .A(int_data_res_1__7__2_), .B(pe_1_1_7_n73), 
        .CI(pe_1_1_7_sub_81_carry[2]), .CO(pe_1_1_7_sub_81_carry[3]), .S(
        pe_1_1_7_N72) );
  FA_X1 pe_1_1_7_sub_81_U2_1 ( .A(int_data_res_1__7__1_), .B(pe_1_1_7_n72), 
        .CI(pe_1_1_7_sub_81_carry[1]), .CO(pe_1_1_7_sub_81_carry[2]), .S(
        pe_1_1_7_N71) );
  FA_X1 pe_1_1_7_add_83_U1_7 ( .A(int_data_res_1__7__7_), .B(
        pe_1_1_7_int_data_3_), .CI(pe_1_1_7_add_83_carry[7]), .S(pe_1_1_7_N85)
         );
  FA_X1 pe_1_1_7_add_83_U1_6 ( .A(int_data_res_1__7__6_), .B(
        pe_1_1_7_int_data_3_), .CI(pe_1_1_7_add_83_carry[6]), .CO(
        pe_1_1_7_add_83_carry[7]), .S(pe_1_1_7_N84) );
  FA_X1 pe_1_1_7_add_83_U1_5 ( .A(int_data_res_1__7__5_), .B(
        pe_1_1_7_int_data_3_), .CI(pe_1_1_7_add_83_carry[5]), .CO(
        pe_1_1_7_add_83_carry[6]), .S(pe_1_1_7_N83) );
  FA_X1 pe_1_1_7_add_83_U1_4 ( .A(int_data_res_1__7__4_), .B(
        pe_1_1_7_int_data_3_), .CI(pe_1_1_7_add_83_carry[4]), .CO(
        pe_1_1_7_add_83_carry[5]), .S(pe_1_1_7_N82) );
  FA_X1 pe_1_1_7_add_83_U1_3 ( .A(int_data_res_1__7__3_), .B(
        pe_1_1_7_int_data_3_), .CI(pe_1_1_7_add_83_carry[3]), .CO(
        pe_1_1_7_add_83_carry[4]), .S(pe_1_1_7_N81) );
  FA_X1 pe_1_1_7_add_83_U1_2 ( .A(int_data_res_1__7__2_), .B(
        pe_1_1_7_int_data_2_), .CI(pe_1_1_7_add_83_carry[2]), .CO(
        pe_1_1_7_add_83_carry[3]), .S(pe_1_1_7_N80) );
  FA_X1 pe_1_1_7_add_83_U1_1 ( .A(int_data_res_1__7__1_), .B(
        pe_1_1_7_int_data_1_), .CI(pe_1_1_7_n2), .CO(pe_1_1_7_add_83_carry[2]), 
        .S(pe_1_1_7_N79) );
  NAND3_X1 pe_1_1_7_U56 ( .A1(pe_1_1_7_n59), .A2(pe_1_1_7_n43), .A3(
        pe_1_1_7_n61), .ZN(pe_1_1_7_n40) );
  NAND3_X1 pe_1_1_7_U55 ( .A1(pe_1_1_7_n43), .A2(pe_1_1_7_n60), .A3(
        pe_1_1_7_n61), .ZN(pe_1_1_7_n39) );
  NAND3_X1 pe_1_1_7_U54 ( .A1(pe_1_1_7_n43), .A2(pe_1_1_7_n62), .A3(
        pe_1_1_7_n59), .ZN(pe_1_1_7_n38) );
  NAND3_X1 pe_1_1_7_U53 ( .A1(pe_1_1_7_n60), .A2(pe_1_1_7_n62), .A3(
        pe_1_1_7_n43), .ZN(pe_1_1_7_n37) );
  DFFR_X1 pe_1_1_7_int_q_acc_reg_6_ ( .D(pe_1_1_7_n76), .CK(pe_1_1_7_net6382), 
        .RN(pe_1_1_7_n69), .Q(int_data_res_1__7__6_) );
  DFFR_X1 pe_1_1_7_int_q_acc_reg_5_ ( .D(pe_1_1_7_n77), .CK(pe_1_1_7_net6382), 
        .RN(pe_1_1_7_n69), .Q(int_data_res_1__7__5_) );
  DFFR_X1 pe_1_1_7_int_q_acc_reg_4_ ( .D(pe_1_1_7_n78), .CK(pe_1_1_7_net6382), 
        .RN(pe_1_1_7_n69), .Q(int_data_res_1__7__4_) );
  DFFR_X1 pe_1_1_7_int_q_acc_reg_3_ ( .D(pe_1_1_7_n79), .CK(pe_1_1_7_net6382), 
        .RN(pe_1_1_7_n69), .Q(int_data_res_1__7__3_) );
  DFFR_X1 pe_1_1_7_int_q_acc_reg_2_ ( .D(pe_1_1_7_n80), .CK(pe_1_1_7_net6382), 
        .RN(pe_1_1_7_n69), .Q(int_data_res_1__7__2_) );
  DFFR_X1 pe_1_1_7_int_q_acc_reg_1_ ( .D(pe_1_1_7_n81), .CK(pe_1_1_7_net6382), 
        .RN(pe_1_1_7_n69), .Q(int_data_res_1__7__1_) );
  DFFR_X1 pe_1_1_7_int_q_acc_reg_7_ ( .D(pe_1_1_7_n75), .CK(pe_1_1_7_net6382), 
        .RN(pe_1_1_7_n69), .Q(int_data_res_1__7__7_) );
  CLKGATETST_X1 pe_1_1_7_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_1_7_n86), .SE(1'b0), .GCK(pe_1_1_7_net6321) );
  CLKGATETST_X1 pe_1_1_7_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_1_7_n85), .SE(1'b0), .GCK(pe_1_1_7_net6327) );
  CLKGATETST_X1 pe_1_1_7_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_1_7_n84), .SE(1'b0), .GCK(pe_1_1_7_net6332) );
  CLKGATETST_X1 pe_1_1_7_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_1_7_n83), .SE(1'b0), .GCK(pe_1_1_7_net6337) );
  CLKGATETST_X1 pe_1_1_7_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_1_7_n88), .SE(1'b0), .GCK(pe_1_1_7_net6342) );
  CLKGATETST_X1 pe_1_1_7_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_1_7_n87), .SE(1'b0), .GCK(pe_1_1_7_net6347) );
  CLKGATETST_X1 pe_1_1_7_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_1_7_N64), .SE(1'b0), .GCK(pe_1_1_7_net6352) );
  CLKGATETST_X1 pe_1_1_7_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_1_7_N63), .SE(1'b0), .GCK(pe_1_1_7_net6357) );
  CLKGATETST_X1 pe_1_1_7_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_1_7_N62), .SE(1'b0), .GCK(pe_1_1_7_net6362) );
  CLKGATETST_X1 pe_1_1_7_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_1_7_N61), .SE(1'b0), .GCK(pe_1_1_7_net6367) );
  CLKGATETST_X1 pe_1_1_7_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_1_7_N60), .SE(1'b0), .GCK(pe_1_1_7_net6372) );
  CLKGATETST_X1 pe_1_1_7_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_1_7_N59), .SE(1'b0), .GCK(pe_1_1_7_net6377) );
  CLKGATETST_X1 pe_1_1_7_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_1_7_N90), .SE(1'b0), .GCK(pe_1_1_7_net6382) );
  CLKBUF_X1 pe_1_2_0_U111 ( .A(pe_1_2_0_n71), .Z(pe_1_2_0_n70) );
  INV_X1 pe_1_2_0_U110 ( .A(n74), .ZN(pe_1_2_0_n69) );
  INV_X1 pe_1_2_0_U109 ( .A(n66), .ZN(pe_1_2_0_n68) );
  INV_X1 pe_1_2_0_U108 ( .A(n66), .ZN(pe_1_2_0_n67) );
  INV_X1 pe_1_2_0_U107 ( .A(n66), .ZN(pe_1_2_0_n66) );
  INV_X1 pe_1_2_0_U106 ( .A(pe_1_2_0_n68), .ZN(pe_1_2_0_n65) );
  INV_X1 pe_1_2_0_U105 ( .A(pe_1_2_0_n62), .ZN(pe_1_2_0_n61) );
  INV_X1 pe_1_2_0_U104 ( .A(n26), .ZN(pe_1_2_0_n59) );
  INV_X1 pe_1_2_0_U103 ( .A(pe_1_2_0_n59), .ZN(pe_1_2_0_n58) );
  INV_X1 pe_1_2_0_U102 ( .A(n18), .ZN(pe_1_2_0_n57) );
  MUX2_X1 pe_1_2_0_U101 ( .A(pe_1_2_0_n54), .B(pe_1_2_0_n51), .S(n46), .Z(
        pe_1_2_0_o_data_h_3_) );
  MUX2_X1 pe_1_2_0_U100 ( .A(pe_1_2_0_n53), .B(pe_1_2_0_n52), .S(pe_1_2_0_n61), 
        .Z(pe_1_2_0_n54) );
  MUX2_X1 pe_1_2_0_U99 ( .A(pe_1_2_0_int_q_reg_h[23]), .B(
        pe_1_2_0_int_q_reg_h[19]), .S(pe_1_2_0_n56), .Z(pe_1_2_0_n53) );
  MUX2_X1 pe_1_2_0_U98 ( .A(pe_1_2_0_int_q_reg_h[15]), .B(
        pe_1_2_0_int_q_reg_h[11]), .S(pe_1_2_0_n56), .Z(pe_1_2_0_n52) );
  MUX2_X1 pe_1_2_0_U97 ( .A(pe_1_2_0_int_q_reg_h[7]), .B(
        pe_1_2_0_int_q_reg_h[3]), .S(pe_1_2_0_n56), .Z(pe_1_2_0_n51) );
  MUX2_X1 pe_1_2_0_U96 ( .A(pe_1_2_0_n50), .B(pe_1_2_0_n47), .S(n46), .Z(
        pe_1_2_0_o_data_h_2_) );
  MUX2_X1 pe_1_2_0_U95 ( .A(pe_1_2_0_n49), .B(pe_1_2_0_n48), .S(pe_1_2_0_n61), 
        .Z(pe_1_2_0_n50) );
  MUX2_X1 pe_1_2_0_U94 ( .A(pe_1_2_0_int_q_reg_h[22]), .B(
        pe_1_2_0_int_q_reg_h[18]), .S(pe_1_2_0_n56), .Z(pe_1_2_0_n49) );
  MUX2_X1 pe_1_2_0_U93 ( .A(pe_1_2_0_int_q_reg_h[14]), .B(
        pe_1_2_0_int_q_reg_h[10]), .S(pe_1_2_0_n56), .Z(pe_1_2_0_n48) );
  MUX2_X1 pe_1_2_0_U92 ( .A(pe_1_2_0_int_q_reg_h[6]), .B(
        pe_1_2_0_int_q_reg_h[2]), .S(pe_1_2_0_n56), .Z(pe_1_2_0_n47) );
  MUX2_X1 pe_1_2_0_U91 ( .A(pe_1_2_0_n46), .B(pe_1_2_0_n24), .S(n46), .Z(
        pe_1_2_0_o_data_h_1_) );
  MUX2_X1 pe_1_2_0_U90 ( .A(pe_1_2_0_n45), .B(pe_1_2_0_n25), .S(pe_1_2_0_n61), 
        .Z(pe_1_2_0_n46) );
  MUX2_X1 pe_1_2_0_U89 ( .A(pe_1_2_0_int_q_reg_h[21]), .B(
        pe_1_2_0_int_q_reg_h[17]), .S(pe_1_2_0_n56), .Z(pe_1_2_0_n45) );
  MUX2_X1 pe_1_2_0_U88 ( .A(pe_1_2_0_int_q_reg_h[13]), .B(
        pe_1_2_0_int_q_reg_h[9]), .S(pe_1_2_0_n56), .Z(pe_1_2_0_n25) );
  MUX2_X1 pe_1_2_0_U87 ( .A(pe_1_2_0_int_q_reg_h[5]), .B(
        pe_1_2_0_int_q_reg_h[1]), .S(pe_1_2_0_n56), .Z(pe_1_2_0_n24) );
  MUX2_X1 pe_1_2_0_U86 ( .A(pe_1_2_0_n23), .B(pe_1_2_0_n20), .S(n46), .Z(
        pe_1_2_0_o_data_h_0_) );
  MUX2_X1 pe_1_2_0_U85 ( .A(pe_1_2_0_n22), .B(pe_1_2_0_n21), .S(pe_1_2_0_n61), 
        .Z(pe_1_2_0_n23) );
  MUX2_X1 pe_1_2_0_U84 ( .A(pe_1_2_0_int_q_reg_h[20]), .B(
        pe_1_2_0_int_q_reg_h[16]), .S(pe_1_2_0_n56), .Z(pe_1_2_0_n22) );
  MUX2_X1 pe_1_2_0_U83 ( .A(pe_1_2_0_int_q_reg_h[12]), .B(
        pe_1_2_0_int_q_reg_h[8]), .S(pe_1_2_0_n56), .Z(pe_1_2_0_n21) );
  MUX2_X1 pe_1_2_0_U82 ( .A(pe_1_2_0_int_q_reg_h[4]), .B(
        pe_1_2_0_int_q_reg_h[0]), .S(pe_1_2_0_n56), .Z(pe_1_2_0_n20) );
  MUX2_X1 pe_1_2_0_U81 ( .A(pe_1_2_0_n19), .B(pe_1_2_0_n16), .S(n46), .Z(
        int_data_y_2__0__3_) );
  MUX2_X1 pe_1_2_0_U80 ( .A(pe_1_2_0_n18), .B(pe_1_2_0_n17), .S(pe_1_2_0_n61), 
        .Z(pe_1_2_0_n19) );
  MUX2_X1 pe_1_2_0_U79 ( .A(pe_1_2_0_int_q_reg_v[23]), .B(
        pe_1_2_0_int_q_reg_v[19]), .S(pe_1_2_0_n55), .Z(pe_1_2_0_n18) );
  MUX2_X1 pe_1_2_0_U78 ( .A(pe_1_2_0_int_q_reg_v[15]), .B(
        pe_1_2_0_int_q_reg_v[11]), .S(pe_1_2_0_n55), .Z(pe_1_2_0_n17) );
  MUX2_X1 pe_1_2_0_U77 ( .A(pe_1_2_0_int_q_reg_v[7]), .B(
        pe_1_2_0_int_q_reg_v[3]), .S(pe_1_2_0_n55), .Z(pe_1_2_0_n16) );
  MUX2_X1 pe_1_2_0_U76 ( .A(pe_1_2_0_n15), .B(pe_1_2_0_n12), .S(n46), .Z(
        int_data_y_2__0__2_) );
  MUX2_X1 pe_1_2_0_U75 ( .A(pe_1_2_0_n14), .B(pe_1_2_0_n13), .S(pe_1_2_0_n61), 
        .Z(pe_1_2_0_n15) );
  MUX2_X1 pe_1_2_0_U74 ( .A(pe_1_2_0_int_q_reg_v[22]), .B(
        pe_1_2_0_int_q_reg_v[18]), .S(pe_1_2_0_n55), .Z(pe_1_2_0_n14) );
  MUX2_X1 pe_1_2_0_U73 ( .A(pe_1_2_0_int_q_reg_v[14]), .B(
        pe_1_2_0_int_q_reg_v[10]), .S(pe_1_2_0_n55), .Z(pe_1_2_0_n13) );
  MUX2_X1 pe_1_2_0_U72 ( .A(pe_1_2_0_int_q_reg_v[6]), .B(
        pe_1_2_0_int_q_reg_v[2]), .S(pe_1_2_0_n55), .Z(pe_1_2_0_n12) );
  MUX2_X1 pe_1_2_0_U71 ( .A(pe_1_2_0_n11), .B(pe_1_2_0_n8), .S(n46), .Z(
        int_data_y_2__0__1_) );
  MUX2_X1 pe_1_2_0_U70 ( .A(pe_1_2_0_n10), .B(pe_1_2_0_n9), .S(pe_1_2_0_n61), 
        .Z(pe_1_2_0_n11) );
  MUX2_X1 pe_1_2_0_U69 ( .A(pe_1_2_0_int_q_reg_v[21]), .B(
        pe_1_2_0_int_q_reg_v[17]), .S(pe_1_2_0_n55), .Z(pe_1_2_0_n10) );
  MUX2_X1 pe_1_2_0_U68 ( .A(pe_1_2_0_int_q_reg_v[13]), .B(
        pe_1_2_0_int_q_reg_v[9]), .S(pe_1_2_0_n55), .Z(pe_1_2_0_n9) );
  MUX2_X1 pe_1_2_0_U67 ( .A(pe_1_2_0_int_q_reg_v[5]), .B(
        pe_1_2_0_int_q_reg_v[1]), .S(pe_1_2_0_n55), .Z(pe_1_2_0_n8) );
  MUX2_X1 pe_1_2_0_U66 ( .A(pe_1_2_0_n7), .B(pe_1_2_0_n4), .S(n46), .Z(
        int_data_y_2__0__0_) );
  MUX2_X1 pe_1_2_0_U65 ( .A(pe_1_2_0_n6), .B(pe_1_2_0_n5), .S(pe_1_2_0_n61), 
        .Z(pe_1_2_0_n7) );
  MUX2_X1 pe_1_2_0_U64 ( .A(pe_1_2_0_int_q_reg_v[20]), .B(
        pe_1_2_0_int_q_reg_v[16]), .S(pe_1_2_0_n55), .Z(pe_1_2_0_n6) );
  MUX2_X1 pe_1_2_0_U63 ( .A(pe_1_2_0_int_q_reg_v[12]), .B(
        pe_1_2_0_int_q_reg_v[8]), .S(pe_1_2_0_n55), .Z(pe_1_2_0_n5) );
  MUX2_X1 pe_1_2_0_U62 ( .A(pe_1_2_0_int_q_reg_v[4]), .B(
        pe_1_2_0_int_q_reg_v[0]), .S(pe_1_2_0_n55), .Z(pe_1_2_0_n4) );
  AND2_X1 pe_1_2_0_U61 ( .A1(pe_1_2_0_o_data_h_3_), .A2(pe_1_2_0_n58), .ZN(
        pe_1_2_0_int_data_3_) );
  NAND2_X1 pe_1_2_0_U60 ( .A1(pe_1_2_0_int_data_0_), .A2(pe_1_2_0_n3), .ZN(
        pe_1_2_0_sub_81_carry[1]) );
  INV_X1 pe_1_2_0_U59 ( .A(pe_1_2_0_int_data_1_), .ZN(pe_1_2_0_n73) );
  AOI222_X1 pe_1_2_0_U58 ( .A1(pe_1_2_0_n63), .A2(int_data_res_3__0__7_), .B1(
        pe_1_2_0_N85), .B2(pe_1_2_0_n27), .C1(pe_1_2_0_N77), .C2(pe_1_2_0_n28), 
        .ZN(pe_1_2_0_n26) );
  INV_X1 pe_1_2_0_U57 ( .A(pe_1_2_0_n26), .ZN(pe_1_2_0_n76) );
  AOI222_X1 pe_1_2_0_U52 ( .A1(int_data_res_3__0__1_), .A2(pe_1_2_0_n63), .B1(
        pe_1_2_0_N79), .B2(pe_1_2_0_n27), .C1(pe_1_2_0_N71), .C2(pe_1_2_0_n28), 
        .ZN(pe_1_2_0_n34) );
  INV_X1 pe_1_2_0_U51 ( .A(pe_1_2_0_n34), .ZN(pe_1_2_0_n82) );
  AOI222_X1 pe_1_2_0_U50 ( .A1(int_data_res_3__0__2_), .A2(pe_1_2_0_n63), .B1(
        pe_1_2_0_N80), .B2(pe_1_2_0_n27), .C1(pe_1_2_0_N72), .C2(pe_1_2_0_n28), 
        .ZN(pe_1_2_0_n33) );
  INV_X1 pe_1_2_0_U49 ( .A(pe_1_2_0_n33), .ZN(pe_1_2_0_n81) );
  AOI222_X1 pe_1_2_0_U48 ( .A1(int_data_res_3__0__6_), .A2(pe_1_2_0_n63), .B1(
        pe_1_2_0_N84), .B2(pe_1_2_0_n27), .C1(pe_1_2_0_N76), .C2(pe_1_2_0_n28), 
        .ZN(pe_1_2_0_n29) );
  INV_X1 pe_1_2_0_U47 ( .A(pe_1_2_0_n29), .ZN(pe_1_2_0_n77) );
  AND2_X1 pe_1_2_0_U46 ( .A1(pe_1_2_0_o_data_h_2_), .A2(pe_1_2_0_n58), .ZN(
        pe_1_2_0_int_data_2_) );
  AND2_X1 pe_1_2_0_U45 ( .A1(pe_1_2_0_o_data_h_1_), .A2(pe_1_2_0_n58), .ZN(
        pe_1_2_0_int_data_1_) );
  INV_X1 pe_1_2_0_U44 ( .A(pe_1_2_0_int_data_2_), .ZN(pe_1_2_0_n74) );
  AND2_X1 pe_1_2_0_U43 ( .A1(pe_1_2_0_int_data_0_), .A2(int_data_res_2__0__0_), 
        .ZN(pe_1_2_0_n2) );
  AND2_X1 pe_1_2_0_U42 ( .A1(pe_1_2_0_o_data_h_0_), .A2(pe_1_2_0_n58), .ZN(
        pe_1_2_0_int_data_0_) );
  XNOR2_X1 pe_1_2_0_U41 ( .A(pe_1_2_0_n72), .B(int_data_res_2__0__0_), .ZN(
        pe_1_2_0_N70) );
  AOI222_X1 pe_1_2_0_U40 ( .A1(int_data_res_3__0__0_), .A2(pe_1_2_0_n63), .B1(
        pe_1_2_0_n1), .B2(pe_1_2_0_n27), .C1(pe_1_2_0_N70), .C2(pe_1_2_0_n28), 
        .ZN(pe_1_2_0_n35) );
  INV_X1 pe_1_2_0_U39 ( .A(pe_1_2_0_n35), .ZN(pe_1_2_0_n83) );
  AOI222_X1 pe_1_2_0_U38 ( .A1(int_data_res_3__0__3_), .A2(pe_1_2_0_n63), .B1(
        pe_1_2_0_N81), .B2(pe_1_2_0_n27), .C1(pe_1_2_0_N73), .C2(pe_1_2_0_n28), 
        .ZN(pe_1_2_0_n32) );
  INV_X1 pe_1_2_0_U37 ( .A(pe_1_2_0_n32), .ZN(pe_1_2_0_n80) );
  AOI222_X1 pe_1_2_0_U36 ( .A1(int_data_res_3__0__4_), .A2(pe_1_2_0_n63), .B1(
        pe_1_2_0_N82), .B2(pe_1_2_0_n27), .C1(pe_1_2_0_N74), .C2(pe_1_2_0_n28), 
        .ZN(pe_1_2_0_n31) );
  INV_X1 pe_1_2_0_U35 ( .A(pe_1_2_0_n31), .ZN(pe_1_2_0_n79) );
  AOI222_X1 pe_1_2_0_U34 ( .A1(int_data_res_3__0__5_), .A2(pe_1_2_0_n63), .B1(
        pe_1_2_0_N83), .B2(pe_1_2_0_n27), .C1(pe_1_2_0_N75), .C2(pe_1_2_0_n28), 
        .ZN(pe_1_2_0_n30) );
  INV_X1 pe_1_2_0_U33 ( .A(pe_1_2_0_n30), .ZN(pe_1_2_0_n78) );
  NOR3_X1 pe_1_2_0_U32 ( .A1(pe_1_2_0_n59), .A2(pe_1_2_0_n64), .A3(int_ckg[47]), .ZN(pe_1_2_0_n36) );
  OR2_X1 pe_1_2_0_U31 ( .A1(pe_1_2_0_n36), .A2(pe_1_2_0_n63), .ZN(pe_1_2_0_N90) );
  INV_X1 pe_1_2_0_U30 ( .A(pe_1_2_0_int_data_0_), .ZN(pe_1_2_0_n72) );
  INV_X1 pe_1_2_0_U29 ( .A(n38), .ZN(pe_1_2_0_n62) );
  INV_X1 pe_1_2_0_U28 ( .A(n32), .ZN(pe_1_2_0_n60) );
  INV_X1 pe_1_2_0_U27 ( .A(pe_1_2_0_int_data_3_), .ZN(pe_1_2_0_n75) );
  BUF_X1 pe_1_2_0_U26 ( .A(n60), .Z(pe_1_2_0_n63) );
  NAND2_X1 pe_1_2_0_U25 ( .A1(pe_1_2_0_n44), .A2(pe_1_2_0_n60), .ZN(
        pe_1_2_0_n41) );
  AND3_X1 pe_1_2_0_U24 ( .A1(n74), .A2(pe_1_2_0_n62), .A3(n46), .ZN(
        pe_1_2_0_n44) );
  NOR2_X1 pe_1_2_0_U23 ( .A1(pe_1_2_0_n69), .A2(n46), .ZN(pe_1_2_0_n43) );
  NOR2_X1 pe_1_2_0_U22 ( .A1(pe_1_2_0_n57), .A2(pe_1_2_0_n63), .ZN(
        pe_1_2_0_n28) );
  NOR2_X1 pe_1_2_0_U21 ( .A1(n18), .A2(pe_1_2_0_n63), .ZN(pe_1_2_0_n27) );
  INV_X1 pe_1_2_0_U20 ( .A(pe_1_2_0_n41), .ZN(pe_1_2_0_n89) );
  INV_X1 pe_1_2_0_U19 ( .A(pe_1_2_0_n37), .ZN(pe_1_2_0_n87) );
  INV_X1 pe_1_2_0_U18 ( .A(pe_1_2_0_n38), .ZN(pe_1_2_0_n86) );
  INV_X1 pe_1_2_0_U17 ( .A(pe_1_2_0_n39), .ZN(pe_1_2_0_n85) );
  NOR2_X1 pe_1_2_0_U16 ( .A1(pe_1_2_0_n67), .A2(pe_1_2_0_n42), .ZN(
        pe_1_2_0_N59) );
  NOR2_X1 pe_1_2_0_U15 ( .A1(pe_1_2_0_n67), .A2(pe_1_2_0_n41), .ZN(
        pe_1_2_0_N60) );
  NOR2_X1 pe_1_2_0_U14 ( .A1(pe_1_2_0_n67), .A2(pe_1_2_0_n38), .ZN(
        pe_1_2_0_N63) );
  NOR2_X1 pe_1_2_0_U13 ( .A1(pe_1_2_0_n66), .A2(pe_1_2_0_n40), .ZN(
        pe_1_2_0_N61) );
  NOR2_X1 pe_1_2_0_U12 ( .A1(pe_1_2_0_n66), .A2(pe_1_2_0_n39), .ZN(
        pe_1_2_0_N62) );
  NOR2_X1 pe_1_2_0_U11 ( .A1(pe_1_2_0_n37), .A2(pe_1_2_0_n66), .ZN(
        pe_1_2_0_N64) );
  NAND2_X1 pe_1_2_0_U10 ( .A1(pe_1_2_0_n44), .A2(n32), .ZN(pe_1_2_0_n42) );
  BUF_X1 pe_1_2_0_U9 ( .A(n32), .Z(pe_1_2_0_n55) );
  BUF_X1 pe_1_2_0_U8 ( .A(n32), .Z(pe_1_2_0_n56) );
  INV_X1 pe_1_2_0_U7 ( .A(pe_1_2_0_n68), .ZN(pe_1_2_0_n64) );
  INV_X1 pe_1_2_0_U6 ( .A(pe_1_2_0_n42), .ZN(pe_1_2_0_n88) );
  INV_X1 pe_1_2_0_U5 ( .A(pe_1_2_0_n40), .ZN(pe_1_2_0_n84) );
  INV_X2 pe_1_2_0_U4 ( .A(n82), .ZN(pe_1_2_0_n71) );
  XOR2_X1 pe_1_2_0_U3 ( .A(pe_1_2_0_int_data_0_), .B(int_data_res_2__0__0_), 
        .Z(pe_1_2_0_n1) );
  DFFR_X1 pe_1_2_0_int_q_acc_reg_0_ ( .D(pe_1_2_0_n83), .CK(pe_1_2_0_net6304), 
        .RN(pe_1_2_0_n71), .Q(int_data_res_2__0__0_), .QN(pe_1_2_0_n3) );
  DFFR_X1 pe_1_2_0_int_q_reg_v_reg_0__0_ ( .D(int_data_y_3__0__0_), .CK(
        pe_1_2_0_net6274), .RN(pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_v[20]) );
  DFFR_X1 pe_1_2_0_int_q_reg_v_reg_0__1_ ( .D(int_data_y_3__0__1_), .CK(
        pe_1_2_0_net6274), .RN(pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_v[21]) );
  DFFR_X1 pe_1_2_0_int_q_reg_v_reg_0__2_ ( .D(int_data_y_3__0__2_), .CK(
        pe_1_2_0_net6274), .RN(pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_v[22]) );
  DFFR_X1 pe_1_2_0_int_q_reg_v_reg_0__3_ ( .D(int_data_y_3__0__3_), .CK(
        pe_1_2_0_net6274), .RN(pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_v[23]) );
  DFFR_X1 pe_1_2_0_int_q_reg_v_reg_1__0_ ( .D(int_data_y_3__0__0_), .CK(
        pe_1_2_0_net6279), .RN(pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_v[16]) );
  DFFR_X1 pe_1_2_0_int_q_reg_v_reg_1__1_ ( .D(int_data_y_3__0__1_), .CK(
        pe_1_2_0_net6279), .RN(pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_v[17]) );
  DFFR_X1 pe_1_2_0_int_q_reg_v_reg_1__2_ ( .D(int_data_y_3__0__2_), .CK(
        pe_1_2_0_net6279), .RN(pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_v[18]) );
  DFFR_X1 pe_1_2_0_int_q_reg_v_reg_1__3_ ( .D(int_data_y_3__0__3_), .CK(
        pe_1_2_0_net6279), .RN(pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_v[19]) );
  DFFR_X1 pe_1_2_0_int_q_reg_v_reg_2__0_ ( .D(int_data_y_3__0__0_), .CK(
        pe_1_2_0_net6284), .RN(pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_v[12]) );
  DFFR_X1 pe_1_2_0_int_q_reg_v_reg_2__1_ ( .D(int_data_y_3__0__1_), .CK(
        pe_1_2_0_net6284), .RN(pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_v[13]) );
  DFFR_X1 pe_1_2_0_int_q_reg_v_reg_2__2_ ( .D(int_data_y_3__0__2_), .CK(
        pe_1_2_0_net6284), .RN(pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_v[14]) );
  DFFR_X1 pe_1_2_0_int_q_reg_v_reg_2__3_ ( .D(int_data_y_3__0__3_), .CK(
        pe_1_2_0_net6284), .RN(pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_v[15]) );
  DFFR_X1 pe_1_2_0_int_q_reg_v_reg_3__0_ ( .D(int_data_y_3__0__0_), .CK(
        pe_1_2_0_net6289), .RN(pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_v[8]) );
  DFFR_X1 pe_1_2_0_int_q_reg_v_reg_3__1_ ( .D(int_data_y_3__0__1_), .CK(
        pe_1_2_0_net6289), .RN(pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_v[9]) );
  DFFR_X1 pe_1_2_0_int_q_reg_v_reg_3__2_ ( .D(int_data_y_3__0__2_), .CK(
        pe_1_2_0_net6289), .RN(pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_v[10]) );
  DFFR_X1 pe_1_2_0_int_q_reg_v_reg_3__3_ ( .D(int_data_y_3__0__3_), .CK(
        pe_1_2_0_net6289), .RN(pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_v[11]) );
  DFFR_X1 pe_1_2_0_int_q_reg_v_reg_4__0_ ( .D(int_data_y_3__0__0_), .CK(
        pe_1_2_0_net6294), .RN(pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_v[4]) );
  DFFR_X1 pe_1_2_0_int_q_reg_v_reg_4__1_ ( .D(int_data_y_3__0__1_), .CK(
        pe_1_2_0_net6294), .RN(pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_v[5]) );
  DFFR_X1 pe_1_2_0_int_q_reg_v_reg_4__2_ ( .D(int_data_y_3__0__2_), .CK(
        pe_1_2_0_net6294), .RN(pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_v[6]) );
  DFFR_X1 pe_1_2_0_int_q_reg_v_reg_4__3_ ( .D(int_data_y_3__0__3_), .CK(
        pe_1_2_0_net6294), .RN(pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_v[7]) );
  DFFR_X1 pe_1_2_0_int_q_reg_v_reg_5__0_ ( .D(int_data_y_3__0__0_), .CK(
        pe_1_2_0_net6299), .RN(pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_v[0]) );
  DFFR_X1 pe_1_2_0_int_q_reg_v_reg_5__1_ ( .D(int_data_y_3__0__1_), .CK(
        pe_1_2_0_net6299), .RN(pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_v[1]) );
  DFFR_X1 pe_1_2_0_int_q_reg_v_reg_5__2_ ( .D(int_data_y_3__0__2_), .CK(
        pe_1_2_0_net6299), .RN(pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_v[2]) );
  DFFR_X1 pe_1_2_0_int_q_reg_v_reg_5__3_ ( .D(int_data_y_3__0__3_), .CK(
        pe_1_2_0_net6299), .RN(pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_2_0_int_q_reg_h_reg_0__0_ ( .D(int_data_x_2__1__0_), .SI(
        int_data_y_3__0__0_), .SE(pe_1_2_0_n64), .CK(pe_1_2_0_net6243), .RN(
        pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_2_0_int_q_reg_h_reg_0__1_ ( .D(int_data_x_2__1__1_), .SI(
        int_data_y_3__0__1_), .SE(pe_1_2_0_n64), .CK(pe_1_2_0_net6243), .RN(
        pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_2_0_int_q_reg_h_reg_0__2_ ( .D(int_data_x_2__1__2_), .SI(
        int_data_y_3__0__2_), .SE(pe_1_2_0_n64), .CK(pe_1_2_0_net6243), .RN(
        pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_2_0_int_q_reg_h_reg_0__3_ ( .D(int_data_x_2__1__3_), .SI(
        int_data_y_3__0__3_), .SE(pe_1_2_0_n64), .CK(pe_1_2_0_net6243), .RN(
        pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_2_0_int_q_reg_h_reg_1__0_ ( .D(int_data_x_2__1__0_), .SI(
        int_data_y_3__0__0_), .SE(pe_1_2_0_n64), .CK(pe_1_2_0_net6249), .RN(
        pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_2_0_int_q_reg_h_reg_1__1_ ( .D(int_data_x_2__1__1_), .SI(
        int_data_y_3__0__1_), .SE(pe_1_2_0_n64), .CK(pe_1_2_0_net6249), .RN(
        pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_2_0_int_q_reg_h_reg_1__2_ ( .D(int_data_x_2__1__2_), .SI(
        int_data_y_3__0__2_), .SE(pe_1_2_0_n64), .CK(pe_1_2_0_net6249), .RN(
        pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_2_0_int_q_reg_h_reg_1__3_ ( .D(int_data_x_2__1__3_), .SI(
        int_data_y_3__0__3_), .SE(pe_1_2_0_n64), .CK(pe_1_2_0_net6249), .RN(
        pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_2_0_int_q_reg_h_reg_2__0_ ( .D(int_data_x_2__1__0_), .SI(
        int_data_y_3__0__0_), .SE(pe_1_2_0_n64), .CK(pe_1_2_0_net6254), .RN(
        pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_2_0_int_q_reg_h_reg_2__1_ ( .D(int_data_x_2__1__1_), .SI(
        int_data_y_3__0__1_), .SE(pe_1_2_0_n64), .CK(pe_1_2_0_net6254), .RN(
        pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_2_0_int_q_reg_h_reg_2__2_ ( .D(int_data_x_2__1__2_), .SI(
        int_data_y_3__0__2_), .SE(pe_1_2_0_n64), .CK(pe_1_2_0_net6254), .RN(
        pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_2_0_int_q_reg_h_reg_2__3_ ( .D(int_data_x_2__1__3_), .SI(
        int_data_y_3__0__3_), .SE(pe_1_2_0_n64), .CK(pe_1_2_0_net6254), .RN(
        pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_2_0_int_q_reg_h_reg_3__0_ ( .D(int_data_x_2__1__0_), .SI(
        int_data_y_3__0__0_), .SE(pe_1_2_0_n64), .CK(pe_1_2_0_net6259), .RN(
        pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_2_0_int_q_reg_h_reg_3__1_ ( .D(int_data_x_2__1__1_), .SI(
        int_data_y_3__0__1_), .SE(pe_1_2_0_n64), .CK(pe_1_2_0_net6259), .RN(
        pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_2_0_int_q_reg_h_reg_3__2_ ( .D(int_data_x_2__1__2_), .SI(
        int_data_y_3__0__2_), .SE(pe_1_2_0_n64), .CK(pe_1_2_0_net6259), .RN(
        pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_2_0_int_q_reg_h_reg_3__3_ ( .D(int_data_x_2__1__3_), .SI(
        int_data_y_3__0__3_), .SE(pe_1_2_0_n64), .CK(pe_1_2_0_net6259), .RN(
        pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_2_0_int_q_reg_h_reg_4__0_ ( .D(int_data_x_2__1__0_), .SI(
        int_data_y_3__0__0_), .SE(pe_1_2_0_n65), .CK(pe_1_2_0_net6264), .RN(
        pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_2_0_int_q_reg_h_reg_4__1_ ( .D(int_data_x_2__1__1_), .SI(
        int_data_y_3__0__1_), .SE(pe_1_2_0_n65), .CK(pe_1_2_0_net6264), .RN(
        pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_2_0_int_q_reg_h_reg_4__2_ ( .D(int_data_x_2__1__2_), .SI(
        int_data_y_3__0__2_), .SE(pe_1_2_0_n65), .CK(pe_1_2_0_net6264), .RN(
        pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_2_0_int_q_reg_h_reg_4__3_ ( .D(int_data_x_2__1__3_), .SI(
        int_data_y_3__0__3_), .SE(pe_1_2_0_n65), .CK(pe_1_2_0_net6264), .RN(
        pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_2_0_int_q_reg_h_reg_5__0_ ( .D(int_data_x_2__1__0_), .SI(
        int_data_y_3__0__0_), .SE(pe_1_2_0_n65), .CK(pe_1_2_0_net6269), .RN(
        pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_2_0_int_q_reg_h_reg_5__1_ ( .D(int_data_x_2__1__1_), .SI(
        int_data_y_3__0__1_), .SE(pe_1_2_0_n65), .CK(pe_1_2_0_net6269), .RN(
        pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_2_0_int_q_reg_h_reg_5__2_ ( .D(int_data_x_2__1__2_), .SI(
        int_data_y_3__0__2_), .SE(pe_1_2_0_n65), .CK(pe_1_2_0_net6269), .RN(
        pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_2_0_int_q_reg_h_reg_5__3_ ( .D(int_data_x_2__1__3_), .SI(
        int_data_y_3__0__3_), .SE(pe_1_2_0_n65), .CK(pe_1_2_0_net6269), .RN(
        pe_1_2_0_n71), .Q(pe_1_2_0_int_q_reg_h[3]) );
  FA_X1 pe_1_2_0_sub_81_U2_7 ( .A(int_data_res_2__0__7_), .B(pe_1_2_0_n75), 
        .CI(pe_1_2_0_sub_81_carry[7]), .S(pe_1_2_0_N77) );
  FA_X1 pe_1_2_0_sub_81_U2_6 ( .A(int_data_res_2__0__6_), .B(pe_1_2_0_n75), 
        .CI(pe_1_2_0_sub_81_carry[6]), .CO(pe_1_2_0_sub_81_carry[7]), .S(
        pe_1_2_0_N76) );
  FA_X1 pe_1_2_0_sub_81_U2_5 ( .A(int_data_res_2__0__5_), .B(pe_1_2_0_n75), 
        .CI(pe_1_2_0_sub_81_carry[5]), .CO(pe_1_2_0_sub_81_carry[6]), .S(
        pe_1_2_0_N75) );
  FA_X1 pe_1_2_0_sub_81_U2_4 ( .A(int_data_res_2__0__4_), .B(pe_1_2_0_n75), 
        .CI(pe_1_2_0_sub_81_carry[4]), .CO(pe_1_2_0_sub_81_carry[5]), .S(
        pe_1_2_0_N74) );
  FA_X1 pe_1_2_0_sub_81_U2_3 ( .A(int_data_res_2__0__3_), .B(pe_1_2_0_n75), 
        .CI(pe_1_2_0_sub_81_carry[3]), .CO(pe_1_2_0_sub_81_carry[4]), .S(
        pe_1_2_0_N73) );
  FA_X1 pe_1_2_0_sub_81_U2_2 ( .A(int_data_res_2__0__2_), .B(pe_1_2_0_n74), 
        .CI(pe_1_2_0_sub_81_carry[2]), .CO(pe_1_2_0_sub_81_carry[3]), .S(
        pe_1_2_0_N72) );
  FA_X1 pe_1_2_0_sub_81_U2_1 ( .A(int_data_res_2__0__1_), .B(pe_1_2_0_n73), 
        .CI(pe_1_2_0_sub_81_carry[1]), .CO(pe_1_2_0_sub_81_carry[2]), .S(
        pe_1_2_0_N71) );
  FA_X1 pe_1_2_0_add_83_U1_7 ( .A(int_data_res_2__0__7_), .B(
        pe_1_2_0_int_data_3_), .CI(pe_1_2_0_add_83_carry[7]), .S(pe_1_2_0_N85)
         );
  FA_X1 pe_1_2_0_add_83_U1_6 ( .A(int_data_res_2__0__6_), .B(
        pe_1_2_0_int_data_3_), .CI(pe_1_2_0_add_83_carry[6]), .CO(
        pe_1_2_0_add_83_carry[7]), .S(pe_1_2_0_N84) );
  FA_X1 pe_1_2_0_add_83_U1_5 ( .A(int_data_res_2__0__5_), .B(
        pe_1_2_0_int_data_3_), .CI(pe_1_2_0_add_83_carry[5]), .CO(
        pe_1_2_0_add_83_carry[6]), .S(pe_1_2_0_N83) );
  FA_X1 pe_1_2_0_add_83_U1_4 ( .A(int_data_res_2__0__4_), .B(
        pe_1_2_0_int_data_3_), .CI(pe_1_2_0_add_83_carry[4]), .CO(
        pe_1_2_0_add_83_carry[5]), .S(pe_1_2_0_N82) );
  FA_X1 pe_1_2_0_add_83_U1_3 ( .A(int_data_res_2__0__3_), .B(
        pe_1_2_0_int_data_3_), .CI(pe_1_2_0_add_83_carry[3]), .CO(
        pe_1_2_0_add_83_carry[4]), .S(pe_1_2_0_N81) );
  FA_X1 pe_1_2_0_add_83_U1_2 ( .A(int_data_res_2__0__2_), .B(
        pe_1_2_0_int_data_2_), .CI(pe_1_2_0_add_83_carry[2]), .CO(
        pe_1_2_0_add_83_carry[3]), .S(pe_1_2_0_N80) );
  FA_X1 pe_1_2_0_add_83_U1_1 ( .A(int_data_res_2__0__1_), .B(
        pe_1_2_0_int_data_1_), .CI(pe_1_2_0_n2), .CO(pe_1_2_0_add_83_carry[2]), 
        .S(pe_1_2_0_N79) );
  NAND3_X1 pe_1_2_0_U56 ( .A1(n32), .A2(pe_1_2_0_n43), .A3(pe_1_2_0_n61), .ZN(
        pe_1_2_0_n40) );
  NAND3_X1 pe_1_2_0_U55 ( .A1(pe_1_2_0_n43), .A2(pe_1_2_0_n60), .A3(
        pe_1_2_0_n61), .ZN(pe_1_2_0_n39) );
  NAND3_X1 pe_1_2_0_U54 ( .A1(pe_1_2_0_n43), .A2(pe_1_2_0_n62), .A3(n32), .ZN(
        pe_1_2_0_n38) );
  NAND3_X1 pe_1_2_0_U53 ( .A1(pe_1_2_0_n60), .A2(pe_1_2_0_n62), .A3(
        pe_1_2_0_n43), .ZN(pe_1_2_0_n37) );
  DFFR_X1 pe_1_2_0_int_q_acc_reg_6_ ( .D(pe_1_2_0_n77), .CK(pe_1_2_0_net6304), 
        .RN(pe_1_2_0_n70), .Q(int_data_res_2__0__6_) );
  DFFR_X1 pe_1_2_0_int_q_acc_reg_5_ ( .D(pe_1_2_0_n78), .CK(pe_1_2_0_net6304), 
        .RN(pe_1_2_0_n70), .Q(int_data_res_2__0__5_) );
  DFFR_X1 pe_1_2_0_int_q_acc_reg_4_ ( .D(pe_1_2_0_n79), .CK(pe_1_2_0_net6304), 
        .RN(pe_1_2_0_n70), .Q(int_data_res_2__0__4_) );
  DFFR_X1 pe_1_2_0_int_q_acc_reg_3_ ( .D(pe_1_2_0_n80), .CK(pe_1_2_0_net6304), 
        .RN(pe_1_2_0_n70), .Q(int_data_res_2__0__3_) );
  DFFR_X1 pe_1_2_0_int_q_acc_reg_2_ ( .D(pe_1_2_0_n81), .CK(pe_1_2_0_net6304), 
        .RN(pe_1_2_0_n70), .Q(int_data_res_2__0__2_) );
  DFFR_X1 pe_1_2_0_int_q_acc_reg_1_ ( .D(pe_1_2_0_n82), .CK(pe_1_2_0_net6304), 
        .RN(pe_1_2_0_n70), .Q(int_data_res_2__0__1_) );
  DFFR_X1 pe_1_2_0_int_q_acc_reg_7_ ( .D(pe_1_2_0_n76), .CK(pe_1_2_0_net6304), 
        .RN(pe_1_2_0_n70), .Q(int_data_res_2__0__7_) );
  CLKGATETST_X1 pe_1_2_0_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_2_0_n87), .SE(1'b0), .GCK(pe_1_2_0_net6243) );
  CLKGATETST_X1 pe_1_2_0_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_2_0_n86), .SE(1'b0), .GCK(pe_1_2_0_net6249) );
  CLKGATETST_X1 pe_1_2_0_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_2_0_n85), .SE(1'b0), .GCK(pe_1_2_0_net6254) );
  CLKGATETST_X1 pe_1_2_0_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_2_0_n84), .SE(1'b0), .GCK(pe_1_2_0_net6259) );
  CLKGATETST_X1 pe_1_2_0_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_2_0_n89), .SE(1'b0), .GCK(pe_1_2_0_net6264) );
  CLKGATETST_X1 pe_1_2_0_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_2_0_n88), .SE(1'b0), .GCK(pe_1_2_0_net6269) );
  CLKGATETST_X1 pe_1_2_0_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_2_0_N64), .SE(1'b0), .GCK(pe_1_2_0_net6274) );
  CLKGATETST_X1 pe_1_2_0_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_2_0_N63), .SE(1'b0), .GCK(pe_1_2_0_net6279) );
  CLKGATETST_X1 pe_1_2_0_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_2_0_N62), .SE(1'b0), .GCK(pe_1_2_0_net6284) );
  CLKGATETST_X1 pe_1_2_0_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_2_0_N61), .SE(1'b0), .GCK(pe_1_2_0_net6289) );
  CLKGATETST_X1 pe_1_2_0_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_2_0_N60), .SE(1'b0), .GCK(pe_1_2_0_net6294) );
  CLKGATETST_X1 pe_1_2_0_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_2_0_N59), .SE(1'b0), .GCK(pe_1_2_0_net6299) );
  CLKGATETST_X1 pe_1_2_0_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_2_0_N90), .SE(1'b0), .GCK(pe_1_2_0_net6304) );
  CLKBUF_X1 pe_1_2_1_U112 ( .A(pe_1_2_1_n72), .Z(pe_1_2_1_n71) );
  INV_X1 pe_1_2_1_U111 ( .A(n74), .ZN(pe_1_2_1_n70) );
  INV_X1 pe_1_2_1_U110 ( .A(n66), .ZN(pe_1_2_1_n69) );
  INV_X1 pe_1_2_1_U109 ( .A(n66), .ZN(pe_1_2_1_n68) );
  INV_X1 pe_1_2_1_U108 ( .A(n66), .ZN(pe_1_2_1_n67) );
  INV_X1 pe_1_2_1_U107 ( .A(pe_1_2_1_n69), .ZN(pe_1_2_1_n66) );
  INV_X1 pe_1_2_1_U106 ( .A(pe_1_2_1_n63), .ZN(pe_1_2_1_n62) );
  INV_X1 pe_1_2_1_U105 ( .A(pe_1_2_1_n61), .ZN(pe_1_2_1_n60) );
  INV_X1 pe_1_2_1_U104 ( .A(n26), .ZN(pe_1_2_1_n59) );
  INV_X1 pe_1_2_1_U103 ( .A(pe_1_2_1_n59), .ZN(pe_1_2_1_n58) );
  INV_X1 pe_1_2_1_U102 ( .A(n18), .ZN(pe_1_2_1_n57) );
  MUX2_X1 pe_1_2_1_U101 ( .A(pe_1_2_1_n54), .B(pe_1_2_1_n51), .S(n46), .Z(
        int_data_x_2__1__3_) );
  MUX2_X1 pe_1_2_1_U100 ( .A(pe_1_2_1_n53), .B(pe_1_2_1_n52), .S(pe_1_2_1_n62), 
        .Z(pe_1_2_1_n54) );
  MUX2_X1 pe_1_2_1_U99 ( .A(pe_1_2_1_int_q_reg_h[23]), .B(
        pe_1_2_1_int_q_reg_h[19]), .S(pe_1_2_1_n56), .Z(pe_1_2_1_n53) );
  MUX2_X1 pe_1_2_1_U98 ( .A(pe_1_2_1_int_q_reg_h[15]), .B(
        pe_1_2_1_int_q_reg_h[11]), .S(pe_1_2_1_n56), .Z(pe_1_2_1_n52) );
  MUX2_X1 pe_1_2_1_U97 ( .A(pe_1_2_1_int_q_reg_h[7]), .B(
        pe_1_2_1_int_q_reg_h[3]), .S(pe_1_2_1_n56), .Z(pe_1_2_1_n51) );
  MUX2_X1 pe_1_2_1_U96 ( .A(pe_1_2_1_n50), .B(pe_1_2_1_n47), .S(n46), .Z(
        int_data_x_2__1__2_) );
  MUX2_X1 pe_1_2_1_U95 ( .A(pe_1_2_1_n49), .B(pe_1_2_1_n48), .S(pe_1_2_1_n62), 
        .Z(pe_1_2_1_n50) );
  MUX2_X1 pe_1_2_1_U94 ( .A(pe_1_2_1_int_q_reg_h[22]), .B(
        pe_1_2_1_int_q_reg_h[18]), .S(pe_1_2_1_n56), .Z(pe_1_2_1_n49) );
  MUX2_X1 pe_1_2_1_U93 ( .A(pe_1_2_1_int_q_reg_h[14]), .B(
        pe_1_2_1_int_q_reg_h[10]), .S(pe_1_2_1_n56), .Z(pe_1_2_1_n48) );
  MUX2_X1 pe_1_2_1_U92 ( .A(pe_1_2_1_int_q_reg_h[6]), .B(
        pe_1_2_1_int_q_reg_h[2]), .S(pe_1_2_1_n56), .Z(pe_1_2_1_n47) );
  MUX2_X1 pe_1_2_1_U91 ( .A(pe_1_2_1_n46), .B(pe_1_2_1_n24), .S(n46), .Z(
        int_data_x_2__1__1_) );
  MUX2_X1 pe_1_2_1_U90 ( .A(pe_1_2_1_n45), .B(pe_1_2_1_n25), .S(pe_1_2_1_n62), 
        .Z(pe_1_2_1_n46) );
  MUX2_X1 pe_1_2_1_U89 ( .A(pe_1_2_1_int_q_reg_h[21]), .B(
        pe_1_2_1_int_q_reg_h[17]), .S(pe_1_2_1_n56), .Z(pe_1_2_1_n45) );
  MUX2_X1 pe_1_2_1_U88 ( .A(pe_1_2_1_int_q_reg_h[13]), .B(
        pe_1_2_1_int_q_reg_h[9]), .S(pe_1_2_1_n56), .Z(pe_1_2_1_n25) );
  MUX2_X1 pe_1_2_1_U87 ( .A(pe_1_2_1_int_q_reg_h[5]), .B(
        pe_1_2_1_int_q_reg_h[1]), .S(pe_1_2_1_n56), .Z(pe_1_2_1_n24) );
  MUX2_X1 pe_1_2_1_U86 ( .A(pe_1_2_1_n23), .B(pe_1_2_1_n20), .S(n46), .Z(
        int_data_x_2__1__0_) );
  MUX2_X1 pe_1_2_1_U85 ( .A(pe_1_2_1_n22), .B(pe_1_2_1_n21), .S(pe_1_2_1_n62), 
        .Z(pe_1_2_1_n23) );
  MUX2_X1 pe_1_2_1_U84 ( .A(pe_1_2_1_int_q_reg_h[20]), .B(
        pe_1_2_1_int_q_reg_h[16]), .S(pe_1_2_1_n56), .Z(pe_1_2_1_n22) );
  MUX2_X1 pe_1_2_1_U83 ( .A(pe_1_2_1_int_q_reg_h[12]), .B(
        pe_1_2_1_int_q_reg_h[8]), .S(pe_1_2_1_n56), .Z(pe_1_2_1_n21) );
  MUX2_X1 pe_1_2_1_U82 ( .A(pe_1_2_1_int_q_reg_h[4]), .B(
        pe_1_2_1_int_q_reg_h[0]), .S(pe_1_2_1_n56), .Z(pe_1_2_1_n20) );
  MUX2_X1 pe_1_2_1_U81 ( .A(pe_1_2_1_n19), .B(pe_1_2_1_n16), .S(n46), .Z(
        int_data_y_2__1__3_) );
  MUX2_X1 pe_1_2_1_U80 ( .A(pe_1_2_1_n18), .B(pe_1_2_1_n17), .S(pe_1_2_1_n62), 
        .Z(pe_1_2_1_n19) );
  MUX2_X1 pe_1_2_1_U79 ( .A(pe_1_2_1_int_q_reg_v[23]), .B(
        pe_1_2_1_int_q_reg_v[19]), .S(pe_1_2_1_n55), .Z(pe_1_2_1_n18) );
  MUX2_X1 pe_1_2_1_U78 ( .A(pe_1_2_1_int_q_reg_v[15]), .B(
        pe_1_2_1_int_q_reg_v[11]), .S(pe_1_2_1_n55), .Z(pe_1_2_1_n17) );
  MUX2_X1 pe_1_2_1_U77 ( .A(pe_1_2_1_int_q_reg_v[7]), .B(
        pe_1_2_1_int_q_reg_v[3]), .S(pe_1_2_1_n55), .Z(pe_1_2_1_n16) );
  MUX2_X1 pe_1_2_1_U76 ( .A(pe_1_2_1_n15), .B(pe_1_2_1_n12), .S(n46), .Z(
        int_data_y_2__1__2_) );
  MUX2_X1 pe_1_2_1_U75 ( .A(pe_1_2_1_n14), .B(pe_1_2_1_n13), .S(pe_1_2_1_n62), 
        .Z(pe_1_2_1_n15) );
  MUX2_X1 pe_1_2_1_U74 ( .A(pe_1_2_1_int_q_reg_v[22]), .B(
        pe_1_2_1_int_q_reg_v[18]), .S(pe_1_2_1_n55), .Z(pe_1_2_1_n14) );
  MUX2_X1 pe_1_2_1_U73 ( .A(pe_1_2_1_int_q_reg_v[14]), .B(
        pe_1_2_1_int_q_reg_v[10]), .S(pe_1_2_1_n55), .Z(pe_1_2_1_n13) );
  MUX2_X1 pe_1_2_1_U72 ( .A(pe_1_2_1_int_q_reg_v[6]), .B(
        pe_1_2_1_int_q_reg_v[2]), .S(pe_1_2_1_n55), .Z(pe_1_2_1_n12) );
  MUX2_X1 pe_1_2_1_U71 ( .A(pe_1_2_1_n11), .B(pe_1_2_1_n8), .S(n46), .Z(
        int_data_y_2__1__1_) );
  MUX2_X1 pe_1_2_1_U70 ( .A(pe_1_2_1_n10), .B(pe_1_2_1_n9), .S(pe_1_2_1_n62), 
        .Z(pe_1_2_1_n11) );
  MUX2_X1 pe_1_2_1_U69 ( .A(pe_1_2_1_int_q_reg_v[21]), .B(
        pe_1_2_1_int_q_reg_v[17]), .S(pe_1_2_1_n55), .Z(pe_1_2_1_n10) );
  MUX2_X1 pe_1_2_1_U68 ( .A(pe_1_2_1_int_q_reg_v[13]), .B(
        pe_1_2_1_int_q_reg_v[9]), .S(pe_1_2_1_n55), .Z(pe_1_2_1_n9) );
  MUX2_X1 pe_1_2_1_U67 ( .A(pe_1_2_1_int_q_reg_v[5]), .B(
        pe_1_2_1_int_q_reg_v[1]), .S(pe_1_2_1_n55), .Z(pe_1_2_1_n8) );
  MUX2_X1 pe_1_2_1_U66 ( .A(pe_1_2_1_n7), .B(pe_1_2_1_n4), .S(n46), .Z(
        int_data_y_2__1__0_) );
  MUX2_X1 pe_1_2_1_U65 ( .A(pe_1_2_1_n6), .B(pe_1_2_1_n5), .S(pe_1_2_1_n62), 
        .Z(pe_1_2_1_n7) );
  MUX2_X1 pe_1_2_1_U64 ( .A(pe_1_2_1_int_q_reg_v[20]), .B(
        pe_1_2_1_int_q_reg_v[16]), .S(pe_1_2_1_n55), .Z(pe_1_2_1_n6) );
  MUX2_X1 pe_1_2_1_U63 ( .A(pe_1_2_1_int_q_reg_v[12]), .B(
        pe_1_2_1_int_q_reg_v[8]), .S(pe_1_2_1_n55), .Z(pe_1_2_1_n5) );
  MUX2_X1 pe_1_2_1_U62 ( .A(pe_1_2_1_int_q_reg_v[4]), .B(
        pe_1_2_1_int_q_reg_v[0]), .S(pe_1_2_1_n55), .Z(pe_1_2_1_n4) );
  AOI222_X1 pe_1_2_1_U61 ( .A1(int_data_res_3__1__2_), .A2(pe_1_2_1_n64), .B1(
        pe_1_2_1_N80), .B2(pe_1_2_1_n27), .C1(pe_1_2_1_N72), .C2(pe_1_2_1_n28), 
        .ZN(pe_1_2_1_n33) );
  INV_X1 pe_1_2_1_U60 ( .A(pe_1_2_1_n33), .ZN(pe_1_2_1_n82) );
  AOI222_X1 pe_1_2_1_U59 ( .A1(int_data_res_3__1__6_), .A2(pe_1_2_1_n64), .B1(
        pe_1_2_1_N84), .B2(pe_1_2_1_n27), .C1(pe_1_2_1_N76), .C2(pe_1_2_1_n28), 
        .ZN(pe_1_2_1_n29) );
  INV_X1 pe_1_2_1_U58 ( .A(pe_1_2_1_n29), .ZN(pe_1_2_1_n78) );
  XNOR2_X1 pe_1_2_1_U57 ( .A(pe_1_2_1_n73), .B(int_data_res_2__1__0_), .ZN(
        pe_1_2_1_N70) );
  AOI222_X1 pe_1_2_1_U52 ( .A1(int_data_res_3__1__0_), .A2(pe_1_2_1_n64), .B1(
        pe_1_2_1_n1), .B2(pe_1_2_1_n27), .C1(pe_1_2_1_N70), .C2(pe_1_2_1_n28), 
        .ZN(pe_1_2_1_n35) );
  INV_X1 pe_1_2_1_U51 ( .A(pe_1_2_1_n35), .ZN(pe_1_2_1_n84) );
  AOI222_X1 pe_1_2_1_U50 ( .A1(int_data_res_3__1__1_), .A2(pe_1_2_1_n64), .B1(
        pe_1_2_1_N79), .B2(pe_1_2_1_n27), .C1(pe_1_2_1_N71), .C2(pe_1_2_1_n28), 
        .ZN(pe_1_2_1_n34) );
  INV_X1 pe_1_2_1_U49 ( .A(pe_1_2_1_n34), .ZN(pe_1_2_1_n83) );
  AOI222_X1 pe_1_2_1_U48 ( .A1(int_data_res_3__1__3_), .A2(pe_1_2_1_n64), .B1(
        pe_1_2_1_N81), .B2(pe_1_2_1_n27), .C1(pe_1_2_1_N73), .C2(pe_1_2_1_n28), 
        .ZN(pe_1_2_1_n32) );
  INV_X1 pe_1_2_1_U47 ( .A(pe_1_2_1_n32), .ZN(pe_1_2_1_n81) );
  AOI222_X1 pe_1_2_1_U46 ( .A1(int_data_res_3__1__4_), .A2(pe_1_2_1_n64), .B1(
        pe_1_2_1_N82), .B2(pe_1_2_1_n27), .C1(pe_1_2_1_N74), .C2(pe_1_2_1_n28), 
        .ZN(pe_1_2_1_n31) );
  INV_X1 pe_1_2_1_U45 ( .A(pe_1_2_1_n31), .ZN(pe_1_2_1_n80) );
  AOI222_X1 pe_1_2_1_U44 ( .A1(int_data_res_3__1__5_), .A2(pe_1_2_1_n64), .B1(
        pe_1_2_1_N83), .B2(pe_1_2_1_n27), .C1(pe_1_2_1_N75), .C2(pe_1_2_1_n28), 
        .ZN(pe_1_2_1_n30) );
  INV_X1 pe_1_2_1_U43 ( .A(pe_1_2_1_n30), .ZN(pe_1_2_1_n79) );
  NAND2_X1 pe_1_2_1_U42 ( .A1(pe_1_2_1_int_data_0_), .A2(pe_1_2_1_n3), .ZN(
        pe_1_2_1_sub_81_carry[1]) );
  INV_X1 pe_1_2_1_U41 ( .A(pe_1_2_1_int_data_1_), .ZN(pe_1_2_1_n74) );
  INV_X1 pe_1_2_1_U40 ( .A(pe_1_2_1_int_data_2_), .ZN(pe_1_2_1_n75) );
  AND2_X1 pe_1_2_1_U39 ( .A1(pe_1_2_1_int_data_0_), .A2(int_data_res_2__1__0_), 
        .ZN(pe_1_2_1_n2) );
  AOI222_X1 pe_1_2_1_U38 ( .A1(pe_1_2_1_n64), .A2(int_data_res_3__1__7_), .B1(
        pe_1_2_1_N85), .B2(pe_1_2_1_n27), .C1(pe_1_2_1_N77), .C2(pe_1_2_1_n28), 
        .ZN(pe_1_2_1_n26) );
  INV_X1 pe_1_2_1_U37 ( .A(pe_1_2_1_n26), .ZN(pe_1_2_1_n77) );
  NOR3_X1 pe_1_2_1_U36 ( .A1(pe_1_2_1_n59), .A2(pe_1_2_1_n65), .A3(int_ckg[46]), .ZN(pe_1_2_1_n36) );
  OR2_X1 pe_1_2_1_U35 ( .A1(pe_1_2_1_n36), .A2(pe_1_2_1_n64), .ZN(pe_1_2_1_N90) );
  INV_X1 pe_1_2_1_U34 ( .A(n38), .ZN(pe_1_2_1_n63) );
  AND2_X1 pe_1_2_1_U33 ( .A1(int_data_x_2__1__2_), .A2(pe_1_2_1_n58), .ZN(
        pe_1_2_1_int_data_2_) );
  AND2_X1 pe_1_2_1_U32 ( .A1(int_data_x_2__1__1_), .A2(pe_1_2_1_n58), .ZN(
        pe_1_2_1_int_data_1_) );
  AND2_X1 pe_1_2_1_U31 ( .A1(int_data_x_2__1__3_), .A2(pe_1_2_1_n58), .ZN(
        pe_1_2_1_int_data_3_) );
  BUF_X1 pe_1_2_1_U30 ( .A(n60), .Z(pe_1_2_1_n64) );
  INV_X1 pe_1_2_1_U29 ( .A(n32), .ZN(pe_1_2_1_n61) );
  AND2_X1 pe_1_2_1_U28 ( .A1(int_data_x_2__1__0_), .A2(pe_1_2_1_n58), .ZN(
        pe_1_2_1_int_data_0_) );
  NAND2_X1 pe_1_2_1_U27 ( .A1(pe_1_2_1_n44), .A2(pe_1_2_1_n61), .ZN(
        pe_1_2_1_n41) );
  AND3_X1 pe_1_2_1_U26 ( .A1(n74), .A2(pe_1_2_1_n63), .A3(n46), .ZN(
        pe_1_2_1_n44) );
  INV_X1 pe_1_2_1_U25 ( .A(pe_1_2_1_int_data_3_), .ZN(pe_1_2_1_n76) );
  NOR2_X1 pe_1_2_1_U24 ( .A1(pe_1_2_1_n70), .A2(n46), .ZN(pe_1_2_1_n43) );
  NOR2_X1 pe_1_2_1_U23 ( .A1(pe_1_2_1_n57), .A2(pe_1_2_1_n64), .ZN(
        pe_1_2_1_n28) );
  NOR2_X1 pe_1_2_1_U22 ( .A1(n18), .A2(pe_1_2_1_n64), .ZN(pe_1_2_1_n27) );
  INV_X1 pe_1_2_1_U21 ( .A(pe_1_2_1_int_data_0_), .ZN(pe_1_2_1_n73) );
  INV_X1 pe_1_2_1_U20 ( .A(pe_1_2_1_n41), .ZN(pe_1_2_1_n90) );
  INV_X1 pe_1_2_1_U19 ( .A(pe_1_2_1_n37), .ZN(pe_1_2_1_n88) );
  INV_X1 pe_1_2_1_U18 ( .A(pe_1_2_1_n38), .ZN(pe_1_2_1_n87) );
  INV_X1 pe_1_2_1_U17 ( .A(pe_1_2_1_n39), .ZN(pe_1_2_1_n86) );
  NOR2_X1 pe_1_2_1_U16 ( .A1(pe_1_2_1_n68), .A2(pe_1_2_1_n42), .ZN(
        pe_1_2_1_N59) );
  NOR2_X1 pe_1_2_1_U15 ( .A1(pe_1_2_1_n68), .A2(pe_1_2_1_n41), .ZN(
        pe_1_2_1_N60) );
  NOR2_X1 pe_1_2_1_U14 ( .A1(pe_1_2_1_n68), .A2(pe_1_2_1_n38), .ZN(
        pe_1_2_1_N63) );
  NOR2_X1 pe_1_2_1_U13 ( .A1(pe_1_2_1_n67), .A2(pe_1_2_1_n40), .ZN(
        pe_1_2_1_N61) );
  NOR2_X1 pe_1_2_1_U12 ( .A1(pe_1_2_1_n67), .A2(pe_1_2_1_n39), .ZN(
        pe_1_2_1_N62) );
  NOR2_X1 pe_1_2_1_U11 ( .A1(pe_1_2_1_n37), .A2(pe_1_2_1_n67), .ZN(
        pe_1_2_1_N64) );
  NAND2_X1 pe_1_2_1_U10 ( .A1(pe_1_2_1_n44), .A2(pe_1_2_1_n60), .ZN(
        pe_1_2_1_n42) );
  BUF_X1 pe_1_2_1_U9 ( .A(pe_1_2_1_n60), .Z(pe_1_2_1_n55) );
  INV_X1 pe_1_2_1_U8 ( .A(pe_1_2_1_n69), .ZN(pe_1_2_1_n65) );
  BUF_X1 pe_1_2_1_U7 ( .A(pe_1_2_1_n60), .Z(pe_1_2_1_n56) );
  INV_X1 pe_1_2_1_U6 ( .A(pe_1_2_1_n42), .ZN(pe_1_2_1_n89) );
  INV_X1 pe_1_2_1_U5 ( .A(pe_1_2_1_n40), .ZN(pe_1_2_1_n85) );
  INV_X2 pe_1_2_1_U4 ( .A(n82), .ZN(pe_1_2_1_n72) );
  XOR2_X1 pe_1_2_1_U3 ( .A(pe_1_2_1_int_data_0_), .B(int_data_res_2__1__0_), 
        .Z(pe_1_2_1_n1) );
  DFFR_X1 pe_1_2_1_int_q_acc_reg_0_ ( .D(pe_1_2_1_n84), .CK(pe_1_2_1_net6226), 
        .RN(pe_1_2_1_n72), .Q(int_data_res_2__1__0_), .QN(pe_1_2_1_n3) );
  DFFR_X1 pe_1_2_1_int_q_reg_v_reg_0__0_ ( .D(int_data_y_3__1__0_), .CK(
        pe_1_2_1_net6196), .RN(pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_v[20]) );
  DFFR_X1 pe_1_2_1_int_q_reg_v_reg_0__1_ ( .D(int_data_y_3__1__1_), .CK(
        pe_1_2_1_net6196), .RN(pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_v[21]) );
  DFFR_X1 pe_1_2_1_int_q_reg_v_reg_0__2_ ( .D(int_data_y_3__1__2_), .CK(
        pe_1_2_1_net6196), .RN(pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_v[22]) );
  DFFR_X1 pe_1_2_1_int_q_reg_v_reg_0__3_ ( .D(int_data_y_3__1__3_), .CK(
        pe_1_2_1_net6196), .RN(pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_v[23]) );
  DFFR_X1 pe_1_2_1_int_q_reg_v_reg_1__0_ ( .D(int_data_y_3__1__0_), .CK(
        pe_1_2_1_net6201), .RN(pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_v[16]) );
  DFFR_X1 pe_1_2_1_int_q_reg_v_reg_1__1_ ( .D(int_data_y_3__1__1_), .CK(
        pe_1_2_1_net6201), .RN(pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_v[17]) );
  DFFR_X1 pe_1_2_1_int_q_reg_v_reg_1__2_ ( .D(int_data_y_3__1__2_), .CK(
        pe_1_2_1_net6201), .RN(pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_v[18]) );
  DFFR_X1 pe_1_2_1_int_q_reg_v_reg_1__3_ ( .D(int_data_y_3__1__3_), .CK(
        pe_1_2_1_net6201), .RN(pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_v[19]) );
  DFFR_X1 pe_1_2_1_int_q_reg_v_reg_2__0_ ( .D(int_data_y_3__1__0_), .CK(
        pe_1_2_1_net6206), .RN(pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_v[12]) );
  DFFR_X1 pe_1_2_1_int_q_reg_v_reg_2__1_ ( .D(int_data_y_3__1__1_), .CK(
        pe_1_2_1_net6206), .RN(pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_v[13]) );
  DFFR_X1 pe_1_2_1_int_q_reg_v_reg_2__2_ ( .D(int_data_y_3__1__2_), .CK(
        pe_1_2_1_net6206), .RN(pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_v[14]) );
  DFFR_X1 pe_1_2_1_int_q_reg_v_reg_2__3_ ( .D(int_data_y_3__1__3_), .CK(
        pe_1_2_1_net6206), .RN(pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_v[15]) );
  DFFR_X1 pe_1_2_1_int_q_reg_v_reg_3__0_ ( .D(int_data_y_3__1__0_), .CK(
        pe_1_2_1_net6211), .RN(pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_v[8]) );
  DFFR_X1 pe_1_2_1_int_q_reg_v_reg_3__1_ ( .D(int_data_y_3__1__1_), .CK(
        pe_1_2_1_net6211), .RN(pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_v[9]) );
  DFFR_X1 pe_1_2_1_int_q_reg_v_reg_3__2_ ( .D(int_data_y_3__1__2_), .CK(
        pe_1_2_1_net6211), .RN(pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_v[10]) );
  DFFR_X1 pe_1_2_1_int_q_reg_v_reg_3__3_ ( .D(int_data_y_3__1__3_), .CK(
        pe_1_2_1_net6211), .RN(pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_v[11]) );
  DFFR_X1 pe_1_2_1_int_q_reg_v_reg_4__0_ ( .D(int_data_y_3__1__0_), .CK(
        pe_1_2_1_net6216), .RN(pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_v[4]) );
  DFFR_X1 pe_1_2_1_int_q_reg_v_reg_4__1_ ( .D(int_data_y_3__1__1_), .CK(
        pe_1_2_1_net6216), .RN(pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_v[5]) );
  DFFR_X1 pe_1_2_1_int_q_reg_v_reg_4__2_ ( .D(int_data_y_3__1__2_), .CK(
        pe_1_2_1_net6216), .RN(pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_v[6]) );
  DFFR_X1 pe_1_2_1_int_q_reg_v_reg_4__3_ ( .D(int_data_y_3__1__3_), .CK(
        pe_1_2_1_net6216), .RN(pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_v[7]) );
  DFFR_X1 pe_1_2_1_int_q_reg_v_reg_5__0_ ( .D(int_data_y_3__1__0_), .CK(
        pe_1_2_1_net6221), .RN(pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_v[0]) );
  DFFR_X1 pe_1_2_1_int_q_reg_v_reg_5__1_ ( .D(int_data_y_3__1__1_), .CK(
        pe_1_2_1_net6221), .RN(pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_v[1]) );
  DFFR_X1 pe_1_2_1_int_q_reg_v_reg_5__2_ ( .D(int_data_y_3__1__2_), .CK(
        pe_1_2_1_net6221), .RN(pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_v[2]) );
  DFFR_X1 pe_1_2_1_int_q_reg_v_reg_5__3_ ( .D(int_data_y_3__1__3_), .CK(
        pe_1_2_1_net6221), .RN(pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_2_1_int_q_reg_h_reg_0__0_ ( .D(int_data_x_2__2__0_), .SI(
        int_data_y_3__1__0_), .SE(pe_1_2_1_n65), .CK(pe_1_2_1_net6165), .RN(
        pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_2_1_int_q_reg_h_reg_0__1_ ( .D(int_data_x_2__2__1_), .SI(
        int_data_y_3__1__1_), .SE(pe_1_2_1_n65), .CK(pe_1_2_1_net6165), .RN(
        pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_2_1_int_q_reg_h_reg_0__2_ ( .D(int_data_x_2__2__2_), .SI(
        int_data_y_3__1__2_), .SE(pe_1_2_1_n65), .CK(pe_1_2_1_net6165), .RN(
        pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_2_1_int_q_reg_h_reg_0__3_ ( .D(int_data_x_2__2__3_), .SI(
        int_data_y_3__1__3_), .SE(pe_1_2_1_n65), .CK(pe_1_2_1_net6165), .RN(
        pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_2_1_int_q_reg_h_reg_1__0_ ( .D(int_data_x_2__2__0_), .SI(
        int_data_y_3__1__0_), .SE(pe_1_2_1_n65), .CK(pe_1_2_1_net6171), .RN(
        pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_2_1_int_q_reg_h_reg_1__1_ ( .D(int_data_x_2__2__1_), .SI(
        int_data_y_3__1__1_), .SE(pe_1_2_1_n65), .CK(pe_1_2_1_net6171), .RN(
        pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_2_1_int_q_reg_h_reg_1__2_ ( .D(int_data_x_2__2__2_), .SI(
        int_data_y_3__1__2_), .SE(pe_1_2_1_n65), .CK(pe_1_2_1_net6171), .RN(
        pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_2_1_int_q_reg_h_reg_1__3_ ( .D(int_data_x_2__2__3_), .SI(
        int_data_y_3__1__3_), .SE(pe_1_2_1_n65), .CK(pe_1_2_1_net6171), .RN(
        pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_2_1_int_q_reg_h_reg_2__0_ ( .D(int_data_x_2__2__0_), .SI(
        int_data_y_3__1__0_), .SE(pe_1_2_1_n65), .CK(pe_1_2_1_net6176), .RN(
        pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_2_1_int_q_reg_h_reg_2__1_ ( .D(int_data_x_2__2__1_), .SI(
        int_data_y_3__1__1_), .SE(pe_1_2_1_n65), .CK(pe_1_2_1_net6176), .RN(
        pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_2_1_int_q_reg_h_reg_2__2_ ( .D(int_data_x_2__2__2_), .SI(
        int_data_y_3__1__2_), .SE(pe_1_2_1_n65), .CK(pe_1_2_1_net6176), .RN(
        pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_2_1_int_q_reg_h_reg_2__3_ ( .D(int_data_x_2__2__3_), .SI(
        int_data_y_3__1__3_), .SE(pe_1_2_1_n65), .CK(pe_1_2_1_net6176), .RN(
        pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_2_1_int_q_reg_h_reg_3__0_ ( .D(int_data_x_2__2__0_), .SI(
        int_data_y_3__1__0_), .SE(pe_1_2_1_n65), .CK(pe_1_2_1_net6181), .RN(
        pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_2_1_int_q_reg_h_reg_3__1_ ( .D(int_data_x_2__2__1_), .SI(
        int_data_y_3__1__1_), .SE(pe_1_2_1_n65), .CK(pe_1_2_1_net6181), .RN(
        pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_2_1_int_q_reg_h_reg_3__2_ ( .D(int_data_x_2__2__2_), .SI(
        int_data_y_3__1__2_), .SE(pe_1_2_1_n65), .CK(pe_1_2_1_net6181), .RN(
        pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_2_1_int_q_reg_h_reg_3__3_ ( .D(int_data_x_2__2__3_), .SI(
        int_data_y_3__1__3_), .SE(pe_1_2_1_n65), .CK(pe_1_2_1_net6181), .RN(
        pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_2_1_int_q_reg_h_reg_4__0_ ( .D(int_data_x_2__2__0_), .SI(
        int_data_y_3__1__0_), .SE(pe_1_2_1_n66), .CK(pe_1_2_1_net6186), .RN(
        pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_2_1_int_q_reg_h_reg_4__1_ ( .D(int_data_x_2__2__1_), .SI(
        int_data_y_3__1__1_), .SE(pe_1_2_1_n66), .CK(pe_1_2_1_net6186), .RN(
        pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_2_1_int_q_reg_h_reg_4__2_ ( .D(int_data_x_2__2__2_), .SI(
        int_data_y_3__1__2_), .SE(pe_1_2_1_n66), .CK(pe_1_2_1_net6186), .RN(
        pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_2_1_int_q_reg_h_reg_4__3_ ( .D(int_data_x_2__2__3_), .SI(
        int_data_y_3__1__3_), .SE(pe_1_2_1_n66), .CK(pe_1_2_1_net6186), .RN(
        pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_2_1_int_q_reg_h_reg_5__0_ ( .D(int_data_x_2__2__0_), .SI(
        int_data_y_3__1__0_), .SE(pe_1_2_1_n66), .CK(pe_1_2_1_net6191), .RN(
        pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_2_1_int_q_reg_h_reg_5__1_ ( .D(int_data_x_2__2__1_), .SI(
        int_data_y_3__1__1_), .SE(pe_1_2_1_n66), .CK(pe_1_2_1_net6191), .RN(
        pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_2_1_int_q_reg_h_reg_5__2_ ( .D(int_data_x_2__2__2_), .SI(
        int_data_y_3__1__2_), .SE(pe_1_2_1_n66), .CK(pe_1_2_1_net6191), .RN(
        pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_2_1_int_q_reg_h_reg_5__3_ ( .D(int_data_x_2__2__3_), .SI(
        int_data_y_3__1__3_), .SE(pe_1_2_1_n66), .CK(pe_1_2_1_net6191), .RN(
        pe_1_2_1_n72), .Q(pe_1_2_1_int_q_reg_h[3]) );
  FA_X1 pe_1_2_1_sub_81_U2_7 ( .A(int_data_res_2__1__7_), .B(pe_1_2_1_n76), 
        .CI(pe_1_2_1_sub_81_carry[7]), .S(pe_1_2_1_N77) );
  FA_X1 pe_1_2_1_sub_81_U2_6 ( .A(int_data_res_2__1__6_), .B(pe_1_2_1_n76), 
        .CI(pe_1_2_1_sub_81_carry[6]), .CO(pe_1_2_1_sub_81_carry[7]), .S(
        pe_1_2_1_N76) );
  FA_X1 pe_1_2_1_sub_81_U2_5 ( .A(int_data_res_2__1__5_), .B(pe_1_2_1_n76), 
        .CI(pe_1_2_1_sub_81_carry[5]), .CO(pe_1_2_1_sub_81_carry[6]), .S(
        pe_1_2_1_N75) );
  FA_X1 pe_1_2_1_sub_81_U2_4 ( .A(int_data_res_2__1__4_), .B(pe_1_2_1_n76), 
        .CI(pe_1_2_1_sub_81_carry[4]), .CO(pe_1_2_1_sub_81_carry[5]), .S(
        pe_1_2_1_N74) );
  FA_X1 pe_1_2_1_sub_81_U2_3 ( .A(int_data_res_2__1__3_), .B(pe_1_2_1_n76), 
        .CI(pe_1_2_1_sub_81_carry[3]), .CO(pe_1_2_1_sub_81_carry[4]), .S(
        pe_1_2_1_N73) );
  FA_X1 pe_1_2_1_sub_81_U2_2 ( .A(int_data_res_2__1__2_), .B(pe_1_2_1_n75), 
        .CI(pe_1_2_1_sub_81_carry[2]), .CO(pe_1_2_1_sub_81_carry[3]), .S(
        pe_1_2_1_N72) );
  FA_X1 pe_1_2_1_sub_81_U2_1 ( .A(int_data_res_2__1__1_), .B(pe_1_2_1_n74), 
        .CI(pe_1_2_1_sub_81_carry[1]), .CO(pe_1_2_1_sub_81_carry[2]), .S(
        pe_1_2_1_N71) );
  FA_X1 pe_1_2_1_add_83_U1_7 ( .A(int_data_res_2__1__7_), .B(
        pe_1_2_1_int_data_3_), .CI(pe_1_2_1_add_83_carry[7]), .S(pe_1_2_1_N85)
         );
  FA_X1 pe_1_2_1_add_83_U1_6 ( .A(int_data_res_2__1__6_), .B(
        pe_1_2_1_int_data_3_), .CI(pe_1_2_1_add_83_carry[6]), .CO(
        pe_1_2_1_add_83_carry[7]), .S(pe_1_2_1_N84) );
  FA_X1 pe_1_2_1_add_83_U1_5 ( .A(int_data_res_2__1__5_), .B(
        pe_1_2_1_int_data_3_), .CI(pe_1_2_1_add_83_carry[5]), .CO(
        pe_1_2_1_add_83_carry[6]), .S(pe_1_2_1_N83) );
  FA_X1 pe_1_2_1_add_83_U1_4 ( .A(int_data_res_2__1__4_), .B(
        pe_1_2_1_int_data_3_), .CI(pe_1_2_1_add_83_carry[4]), .CO(
        pe_1_2_1_add_83_carry[5]), .S(pe_1_2_1_N82) );
  FA_X1 pe_1_2_1_add_83_U1_3 ( .A(int_data_res_2__1__3_), .B(
        pe_1_2_1_int_data_3_), .CI(pe_1_2_1_add_83_carry[3]), .CO(
        pe_1_2_1_add_83_carry[4]), .S(pe_1_2_1_N81) );
  FA_X1 pe_1_2_1_add_83_U1_2 ( .A(int_data_res_2__1__2_), .B(
        pe_1_2_1_int_data_2_), .CI(pe_1_2_1_add_83_carry[2]), .CO(
        pe_1_2_1_add_83_carry[3]), .S(pe_1_2_1_N80) );
  FA_X1 pe_1_2_1_add_83_U1_1 ( .A(int_data_res_2__1__1_), .B(
        pe_1_2_1_int_data_1_), .CI(pe_1_2_1_n2), .CO(pe_1_2_1_add_83_carry[2]), 
        .S(pe_1_2_1_N79) );
  NAND3_X1 pe_1_2_1_U56 ( .A1(pe_1_2_1_n60), .A2(pe_1_2_1_n43), .A3(
        pe_1_2_1_n62), .ZN(pe_1_2_1_n40) );
  NAND3_X1 pe_1_2_1_U55 ( .A1(pe_1_2_1_n43), .A2(pe_1_2_1_n61), .A3(
        pe_1_2_1_n62), .ZN(pe_1_2_1_n39) );
  NAND3_X1 pe_1_2_1_U54 ( .A1(pe_1_2_1_n43), .A2(pe_1_2_1_n63), .A3(
        pe_1_2_1_n60), .ZN(pe_1_2_1_n38) );
  NAND3_X1 pe_1_2_1_U53 ( .A1(pe_1_2_1_n61), .A2(pe_1_2_1_n63), .A3(
        pe_1_2_1_n43), .ZN(pe_1_2_1_n37) );
  DFFR_X1 pe_1_2_1_int_q_acc_reg_6_ ( .D(pe_1_2_1_n78), .CK(pe_1_2_1_net6226), 
        .RN(pe_1_2_1_n71), .Q(int_data_res_2__1__6_) );
  DFFR_X1 pe_1_2_1_int_q_acc_reg_5_ ( .D(pe_1_2_1_n79), .CK(pe_1_2_1_net6226), 
        .RN(pe_1_2_1_n71), .Q(int_data_res_2__1__5_) );
  DFFR_X1 pe_1_2_1_int_q_acc_reg_4_ ( .D(pe_1_2_1_n80), .CK(pe_1_2_1_net6226), 
        .RN(pe_1_2_1_n71), .Q(int_data_res_2__1__4_) );
  DFFR_X1 pe_1_2_1_int_q_acc_reg_3_ ( .D(pe_1_2_1_n81), .CK(pe_1_2_1_net6226), 
        .RN(pe_1_2_1_n71), .Q(int_data_res_2__1__3_) );
  DFFR_X1 pe_1_2_1_int_q_acc_reg_2_ ( .D(pe_1_2_1_n82), .CK(pe_1_2_1_net6226), 
        .RN(pe_1_2_1_n71), .Q(int_data_res_2__1__2_) );
  DFFR_X1 pe_1_2_1_int_q_acc_reg_1_ ( .D(pe_1_2_1_n83), .CK(pe_1_2_1_net6226), 
        .RN(pe_1_2_1_n71), .Q(int_data_res_2__1__1_) );
  DFFR_X1 pe_1_2_1_int_q_acc_reg_7_ ( .D(pe_1_2_1_n77), .CK(pe_1_2_1_net6226), 
        .RN(pe_1_2_1_n71), .Q(int_data_res_2__1__7_) );
  CLKGATETST_X1 pe_1_2_1_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_2_1_n88), .SE(1'b0), .GCK(pe_1_2_1_net6165) );
  CLKGATETST_X1 pe_1_2_1_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_2_1_n87), .SE(1'b0), .GCK(pe_1_2_1_net6171) );
  CLKGATETST_X1 pe_1_2_1_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_2_1_n86), .SE(1'b0), .GCK(pe_1_2_1_net6176) );
  CLKGATETST_X1 pe_1_2_1_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_2_1_n85), .SE(1'b0), .GCK(pe_1_2_1_net6181) );
  CLKGATETST_X1 pe_1_2_1_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_2_1_n90), .SE(1'b0), .GCK(pe_1_2_1_net6186) );
  CLKGATETST_X1 pe_1_2_1_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_2_1_n89), .SE(1'b0), .GCK(pe_1_2_1_net6191) );
  CLKGATETST_X1 pe_1_2_1_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_2_1_N64), .SE(1'b0), .GCK(pe_1_2_1_net6196) );
  CLKGATETST_X1 pe_1_2_1_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_2_1_N63), .SE(1'b0), .GCK(pe_1_2_1_net6201) );
  CLKGATETST_X1 pe_1_2_1_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_2_1_N62), .SE(1'b0), .GCK(pe_1_2_1_net6206) );
  CLKGATETST_X1 pe_1_2_1_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_2_1_N61), .SE(1'b0), .GCK(pe_1_2_1_net6211) );
  CLKGATETST_X1 pe_1_2_1_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_2_1_N60), .SE(1'b0), .GCK(pe_1_2_1_net6216) );
  CLKGATETST_X1 pe_1_2_1_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_2_1_N59), .SE(1'b0), .GCK(pe_1_2_1_net6221) );
  CLKGATETST_X1 pe_1_2_1_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_2_1_N90), .SE(1'b0), .GCK(pe_1_2_1_net6226) );
  CLKBUF_X1 pe_1_2_2_U112 ( .A(pe_1_2_2_n72), .Z(pe_1_2_2_n71) );
  INV_X1 pe_1_2_2_U111 ( .A(n74), .ZN(pe_1_2_2_n70) );
  INV_X1 pe_1_2_2_U110 ( .A(n66), .ZN(pe_1_2_2_n69) );
  INV_X1 pe_1_2_2_U109 ( .A(n66), .ZN(pe_1_2_2_n68) );
  INV_X1 pe_1_2_2_U108 ( .A(n66), .ZN(pe_1_2_2_n67) );
  INV_X1 pe_1_2_2_U107 ( .A(pe_1_2_2_n69), .ZN(pe_1_2_2_n66) );
  INV_X1 pe_1_2_2_U106 ( .A(pe_1_2_2_n63), .ZN(pe_1_2_2_n62) );
  INV_X1 pe_1_2_2_U105 ( .A(pe_1_2_2_n61), .ZN(pe_1_2_2_n60) );
  INV_X1 pe_1_2_2_U104 ( .A(n26), .ZN(pe_1_2_2_n59) );
  INV_X1 pe_1_2_2_U103 ( .A(pe_1_2_2_n59), .ZN(pe_1_2_2_n58) );
  INV_X1 pe_1_2_2_U102 ( .A(n18), .ZN(pe_1_2_2_n57) );
  MUX2_X1 pe_1_2_2_U101 ( .A(pe_1_2_2_n54), .B(pe_1_2_2_n51), .S(n46), .Z(
        int_data_x_2__2__3_) );
  MUX2_X1 pe_1_2_2_U100 ( .A(pe_1_2_2_n53), .B(pe_1_2_2_n52), .S(pe_1_2_2_n62), 
        .Z(pe_1_2_2_n54) );
  MUX2_X1 pe_1_2_2_U99 ( .A(pe_1_2_2_int_q_reg_h[23]), .B(
        pe_1_2_2_int_q_reg_h[19]), .S(pe_1_2_2_n56), .Z(pe_1_2_2_n53) );
  MUX2_X1 pe_1_2_2_U98 ( .A(pe_1_2_2_int_q_reg_h[15]), .B(
        pe_1_2_2_int_q_reg_h[11]), .S(pe_1_2_2_n56), .Z(pe_1_2_2_n52) );
  MUX2_X1 pe_1_2_2_U97 ( .A(pe_1_2_2_int_q_reg_h[7]), .B(
        pe_1_2_2_int_q_reg_h[3]), .S(pe_1_2_2_n56), .Z(pe_1_2_2_n51) );
  MUX2_X1 pe_1_2_2_U96 ( .A(pe_1_2_2_n50), .B(pe_1_2_2_n47), .S(n46), .Z(
        int_data_x_2__2__2_) );
  MUX2_X1 pe_1_2_2_U95 ( .A(pe_1_2_2_n49), .B(pe_1_2_2_n48), .S(pe_1_2_2_n62), 
        .Z(pe_1_2_2_n50) );
  MUX2_X1 pe_1_2_2_U94 ( .A(pe_1_2_2_int_q_reg_h[22]), .B(
        pe_1_2_2_int_q_reg_h[18]), .S(pe_1_2_2_n56), .Z(pe_1_2_2_n49) );
  MUX2_X1 pe_1_2_2_U93 ( .A(pe_1_2_2_int_q_reg_h[14]), .B(
        pe_1_2_2_int_q_reg_h[10]), .S(pe_1_2_2_n56), .Z(pe_1_2_2_n48) );
  MUX2_X1 pe_1_2_2_U92 ( .A(pe_1_2_2_int_q_reg_h[6]), .B(
        pe_1_2_2_int_q_reg_h[2]), .S(pe_1_2_2_n56), .Z(pe_1_2_2_n47) );
  MUX2_X1 pe_1_2_2_U91 ( .A(pe_1_2_2_n46), .B(pe_1_2_2_n24), .S(n46), .Z(
        int_data_x_2__2__1_) );
  MUX2_X1 pe_1_2_2_U90 ( .A(pe_1_2_2_n45), .B(pe_1_2_2_n25), .S(pe_1_2_2_n62), 
        .Z(pe_1_2_2_n46) );
  MUX2_X1 pe_1_2_2_U89 ( .A(pe_1_2_2_int_q_reg_h[21]), .B(
        pe_1_2_2_int_q_reg_h[17]), .S(pe_1_2_2_n56), .Z(pe_1_2_2_n45) );
  MUX2_X1 pe_1_2_2_U88 ( .A(pe_1_2_2_int_q_reg_h[13]), .B(
        pe_1_2_2_int_q_reg_h[9]), .S(pe_1_2_2_n56), .Z(pe_1_2_2_n25) );
  MUX2_X1 pe_1_2_2_U87 ( .A(pe_1_2_2_int_q_reg_h[5]), .B(
        pe_1_2_2_int_q_reg_h[1]), .S(pe_1_2_2_n56), .Z(pe_1_2_2_n24) );
  MUX2_X1 pe_1_2_2_U86 ( .A(pe_1_2_2_n23), .B(pe_1_2_2_n20), .S(n46), .Z(
        int_data_x_2__2__0_) );
  MUX2_X1 pe_1_2_2_U85 ( .A(pe_1_2_2_n22), .B(pe_1_2_2_n21), .S(pe_1_2_2_n62), 
        .Z(pe_1_2_2_n23) );
  MUX2_X1 pe_1_2_2_U84 ( .A(pe_1_2_2_int_q_reg_h[20]), .B(
        pe_1_2_2_int_q_reg_h[16]), .S(pe_1_2_2_n56), .Z(pe_1_2_2_n22) );
  MUX2_X1 pe_1_2_2_U83 ( .A(pe_1_2_2_int_q_reg_h[12]), .B(
        pe_1_2_2_int_q_reg_h[8]), .S(pe_1_2_2_n56), .Z(pe_1_2_2_n21) );
  MUX2_X1 pe_1_2_2_U82 ( .A(pe_1_2_2_int_q_reg_h[4]), .B(
        pe_1_2_2_int_q_reg_h[0]), .S(pe_1_2_2_n56), .Z(pe_1_2_2_n20) );
  MUX2_X1 pe_1_2_2_U81 ( .A(pe_1_2_2_n19), .B(pe_1_2_2_n16), .S(n46), .Z(
        int_data_y_2__2__3_) );
  MUX2_X1 pe_1_2_2_U80 ( .A(pe_1_2_2_n18), .B(pe_1_2_2_n17), .S(pe_1_2_2_n62), 
        .Z(pe_1_2_2_n19) );
  MUX2_X1 pe_1_2_2_U79 ( .A(pe_1_2_2_int_q_reg_v[23]), .B(
        pe_1_2_2_int_q_reg_v[19]), .S(pe_1_2_2_n55), .Z(pe_1_2_2_n18) );
  MUX2_X1 pe_1_2_2_U78 ( .A(pe_1_2_2_int_q_reg_v[15]), .B(
        pe_1_2_2_int_q_reg_v[11]), .S(pe_1_2_2_n55), .Z(pe_1_2_2_n17) );
  MUX2_X1 pe_1_2_2_U77 ( .A(pe_1_2_2_int_q_reg_v[7]), .B(
        pe_1_2_2_int_q_reg_v[3]), .S(pe_1_2_2_n55), .Z(pe_1_2_2_n16) );
  MUX2_X1 pe_1_2_2_U76 ( .A(pe_1_2_2_n15), .B(pe_1_2_2_n12), .S(n46), .Z(
        int_data_y_2__2__2_) );
  MUX2_X1 pe_1_2_2_U75 ( .A(pe_1_2_2_n14), .B(pe_1_2_2_n13), .S(pe_1_2_2_n62), 
        .Z(pe_1_2_2_n15) );
  MUX2_X1 pe_1_2_2_U74 ( .A(pe_1_2_2_int_q_reg_v[22]), .B(
        pe_1_2_2_int_q_reg_v[18]), .S(pe_1_2_2_n55), .Z(pe_1_2_2_n14) );
  MUX2_X1 pe_1_2_2_U73 ( .A(pe_1_2_2_int_q_reg_v[14]), .B(
        pe_1_2_2_int_q_reg_v[10]), .S(pe_1_2_2_n55), .Z(pe_1_2_2_n13) );
  MUX2_X1 pe_1_2_2_U72 ( .A(pe_1_2_2_int_q_reg_v[6]), .B(
        pe_1_2_2_int_q_reg_v[2]), .S(pe_1_2_2_n55), .Z(pe_1_2_2_n12) );
  MUX2_X1 pe_1_2_2_U71 ( .A(pe_1_2_2_n11), .B(pe_1_2_2_n8), .S(n46), .Z(
        int_data_y_2__2__1_) );
  MUX2_X1 pe_1_2_2_U70 ( .A(pe_1_2_2_n10), .B(pe_1_2_2_n9), .S(pe_1_2_2_n62), 
        .Z(pe_1_2_2_n11) );
  MUX2_X1 pe_1_2_2_U69 ( .A(pe_1_2_2_int_q_reg_v[21]), .B(
        pe_1_2_2_int_q_reg_v[17]), .S(pe_1_2_2_n55), .Z(pe_1_2_2_n10) );
  MUX2_X1 pe_1_2_2_U68 ( .A(pe_1_2_2_int_q_reg_v[13]), .B(
        pe_1_2_2_int_q_reg_v[9]), .S(pe_1_2_2_n55), .Z(pe_1_2_2_n9) );
  MUX2_X1 pe_1_2_2_U67 ( .A(pe_1_2_2_int_q_reg_v[5]), .B(
        pe_1_2_2_int_q_reg_v[1]), .S(pe_1_2_2_n55), .Z(pe_1_2_2_n8) );
  MUX2_X1 pe_1_2_2_U66 ( .A(pe_1_2_2_n7), .B(pe_1_2_2_n4), .S(n46), .Z(
        int_data_y_2__2__0_) );
  MUX2_X1 pe_1_2_2_U65 ( .A(pe_1_2_2_n6), .B(pe_1_2_2_n5), .S(pe_1_2_2_n62), 
        .Z(pe_1_2_2_n7) );
  MUX2_X1 pe_1_2_2_U64 ( .A(pe_1_2_2_int_q_reg_v[20]), .B(
        pe_1_2_2_int_q_reg_v[16]), .S(pe_1_2_2_n55), .Z(pe_1_2_2_n6) );
  MUX2_X1 pe_1_2_2_U63 ( .A(pe_1_2_2_int_q_reg_v[12]), .B(
        pe_1_2_2_int_q_reg_v[8]), .S(pe_1_2_2_n55), .Z(pe_1_2_2_n5) );
  MUX2_X1 pe_1_2_2_U62 ( .A(pe_1_2_2_int_q_reg_v[4]), .B(
        pe_1_2_2_int_q_reg_v[0]), .S(pe_1_2_2_n55), .Z(pe_1_2_2_n4) );
  AOI222_X1 pe_1_2_2_U61 ( .A1(int_data_res_3__2__2_), .A2(pe_1_2_2_n64), .B1(
        pe_1_2_2_N80), .B2(pe_1_2_2_n27), .C1(pe_1_2_2_N72), .C2(pe_1_2_2_n28), 
        .ZN(pe_1_2_2_n33) );
  INV_X1 pe_1_2_2_U60 ( .A(pe_1_2_2_n33), .ZN(pe_1_2_2_n82) );
  AOI222_X1 pe_1_2_2_U59 ( .A1(int_data_res_3__2__6_), .A2(pe_1_2_2_n64), .B1(
        pe_1_2_2_N84), .B2(pe_1_2_2_n27), .C1(pe_1_2_2_N76), .C2(pe_1_2_2_n28), 
        .ZN(pe_1_2_2_n29) );
  INV_X1 pe_1_2_2_U58 ( .A(pe_1_2_2_n29), .ZN(pe_1_2_2_n78) );
  XNOR2_X1 pe_1_2_2_U57 ( .A(pe_1_2_2_n73), .B(int_data_res_2__2__0_), .ZN(
        pe_1_2_2_N70) );
  AOI222_X1 pe_1_2_2_U52 ( .A1(int_data_res_3__2__0_), .A2(pe_1_2_2_n64), .B1(
        pe_1_2_2_n1), .B2(pe_1_2_2_n27), .C1(pe_1_2_2_N70), .C2(pe_1_2_2_n28), 
        .ZN(pe_1_2_2_n35) );
  INV_X1 pe_1_2_2_U51 ( .A(pe_1_2_2_n35), .ZN(pe_1_2_2_n84) );
  AOI222_X1 pe_1_2_2_U50 ( .A1(int_data_res_3__2__1_), .A2(pe_1_2_2_n64), .B1(
        pe_1_2_2_N79), .B2(pe_1_2_2_n27), .C1(pe_1_2_2_N71), .C2(pe_1_2_2_n28), 
        .ZN(pe_1_2_2_n34) );
  INV_X1 pe_1_2_2_U49 ( .A(pe_1_2_2_n34), .ZN(pe_1_2_2_n83) );
  AOI222_X1 pe_1_2_2_U48 ( .A1(int_data_res_3__2__3_), .A2(pe_1_2_2_n64), .B1(
        pe_1_2_2_N81), .B2(pe_1_2_2_n27), .C1(pe_1_2_2_N73), .C2(pe_1_2_2_n28), 
        .ZN(pe_1_2_2_n32) );
  INV_X1 pe_1_2_2_U47 ( .A(pe_1_2_2_n32), .ZN(pe_1_2_2_n81) );
  AOI222_X1 pe_1_2_2_U46 ( .A1(int_data_res_3__2__4_), .A2(pe_1_2_2_n64), .B1(
        pe_1_2_2_N82), .B2(pe_1_2_2_n27), .C1(pe_1_2_2_N74), .C2(pe_1_2_2_n28), 
        .ZN(pe_1_2_2_n31) );
  INV_X1 pe_1_2_2_U45 ( .A(pe_1_2_2_n31), .ZN(pe_1_2_2_n80) );
  AOI222_X1 pe_1_2_2_U44 ( .A1(int_data_res_3__2__5_), .A2(pe_1_2_2_n64), .B1(
        pe_1_2_2_N83), .B2(pe_1_2_2_n27), .C1(pe_1_2_2_N75), .C2(pe_1_2_2_n28), 
        .ZN(pe_1_2_2_n30) );
  INV_X1 pe_1_2_2_U43 ( .A(pe_1_2_2_n30), .ZN(pe_1_2_2_n79) );
  NAND2_X1 pe_1_2_2_U42 ( .A1(pe_1_2_2_int_data_0_), .A2(pe_1_2_2_n3), .ZN(
        pe_1_2_2_sub_81_carry[1]) );
  INV_X1 pe_1_2_2_U41 ( .A(pe_1_2_2_int_data_1_), .ZN(pe_1_2_2_n74) );
  INV_X1 pe_1_2_2_U40 ( .A(pe_1_2_2_int_data_2_), .ZN(pe_1_2_2_n75) );
  AND2_X1 pe_1_2_2_U39 ( .A1(pe_1_2_2_int_data_0_), .A2(int_data_res_2__2__0_), 
        .ZN(pe_1_2_2_n2) );
  AOI222_X1 pe_1_2_2_U38 ( .A1(pe_1_2_2_n64), .A2(int_data_res_3__2__7_), .B1(
        pe_1_2_2_N85), .B2(pe_1_2_2_n27), .C1(pe_1_2_2_N77), .C2(pe_1_2_2_n28), 
        .ZN(pe_1_2_2_n26) );
  INV_X1 pe_1_2_2_U37 ( .A(pe_1_2_2_n26), .ZN(pe_1_2_2_n77) );
  NOR3_X1 pe_1_2_2_U36 ( .A1(pe_1_2_2_n59), .A2(pe_1_2_2_n65), .A3(int_ckg[45]), .ZN(pe_1_2_2_n36) );
  OR2_X1 pe_1_2_2_U35 ( .A1(pe_1_2_2_n36), .A2(pe_1_2_2_n64), .ZN(pe_1_2_2_N90) );
  INV_X1 pe_1_2_2_U34 ( .A(n38), .ZN(pe_1_2_2_n63) );
  AND2_X1 pe_1_2_2_U33 ( .A1(int_data_x_2__2__2_), .A2(pe_1_2_2_n58), .ZN(
        pe_1_2_2_int_data_2_) );
  AND2_X1 pe_1_2_2_U32 ( .A1(int_data_x_2__2__1_), .A2(pe_1_2_2_n58), .ZN(
        pe_1_2_2_int_data_1_) );
  AND2_X1 pe_1_2_2_U31 ( .A1(int_data_x_2__2__3_), .A2(pe_1_2_2_n58), .ZN(
        pe_1_2_2_int_data_3_) );
  BUF_X1 pe_1_2_2_U30 ( .A(n60), .Z(pe_1_2_2_n64) );
  INV_X1 pe_1_2_2_U29 ( .A(n32), .ZN(pe_1_2_2_n61) );
  AND2_X1 pe_1_2_2_U28 ( .A1(int_data_x_2__2__0_), .A2(pe_1_2_2_n58), .ZN(
        pe_1_2_2_int_data_0_) );
  NAND2_X1 pe_1_2_2_U27 ( .A1(pe_1_2_2_n44), .A2(pe_1_2_2_n61), .ZN(
        pe_1_2_2_n41) );
  AND3_X1 pe_1_2_2_U26 ( .A1(n74), .A2(pe_1_2_2_n63), .A3(n46), .ZN(
        pe_1_2_2_n44) );
  INV_X1 pe_1_2_2_U25 ( .A(pe_1_2_2_int_data_3_), .ZN(pe_1_2_2_n76) );
  NOR2_X1 pe_1_2_2_U24 ( .A1(pe_1_2_2_n70), .A2(n46), .ZN(pe_1_2_2_n43) );
  NOR2_X1 pe_1_2_2_U23 ( .A1(pe_1_2_2_n57), .A2(pe_1_2_2_n64), .ZN(
        pe_1_2_2_n28) );
  NOR2_X1 pe_1_2_2_U22 ( .A1(n18), .A2(pe_1_2_2_n64), .ZN(pe_1_2_2_n27) );
  INV_X1 pe_1_2_2_U21 ( .A(pe_1_2_2_int_data_0_), .ZN(pe_1_2_2_n73) );
  INV_X1 pe_1_2_2_U20 ( .A(pe_1_2_2_n41), .ZN(pe_1_2_2_n90) );
  INV_X1 pe_1_2_2_U19 ( .A(pe_1_2_2_n37), .ZN(pe_1_2_2_n88) );
  INV_X1 pe_1_2_2_U18 ( .A(pe_1_2_2_n38), .ZN(pe_1_2_2_n87) );
  INV_X1 pe_1_2_2_U17 ( .A(pe_1_2_2_n39), .ZN(pe_1_2_2_n86) );
  NOR2_X1 pe_1_2_2_U16 ( .A1(pe_1_2_2_n68), .A2(pe_1_2_2_n42), .ZN(
        pe_1_2_2_N59) );
  NOR2_X1 pe_1_2_2_U15 ( .A1(pe_1_2_2_n68), .A2(pe_1_2_2_n41), .ZN(
        pe_1_2_2_N60) );
  NOR2_X1 pe_1_2_2_U14 ( .A1(pe_1_2_2_n68), .A2(pe_1_2_2_n38), .ZN(
        pe_1_2_2_N63) );
  NOR2_X1 pe_1_2_2_U13 ( .A1(pe_1_2_2_n67), .A2(pe_1_2_2_n40), .ZN(
        pe_1_2_2_N61) );
  NOR2_X1 pe_1_2_2_U12 ( .A1(pe_1_2_2_n67), .A2(pe_1_2_2_n39), .ZN(
        pe_1_2_2_N62) );
  NOR2_X1 pe_1_2_2_U11 ( .A1(pe_1_2_2_n37), .A2(pe_1_2_2_n67), .ZN(
        pe_1_2_2_N64) );
  NAND2_X1 pe_1_2_2_U10 ( .A1(pe_1_2_2_n44), .A2(pe_1_2_2_n60), .ZN(
        pe_1_2_2_n42) );
  BUF_X1 pe_1_2_2_U9 ( .A(pe_1_2_2_n60), .Z(pe_1_2_2_n55) );
  INV_X1 pe_1_2_2_U8 ( .A(pe_1_2_2_n69), .ZN(pe_1_2_2_n65) );
  BUF_X1 pe_1_2_2_U7 ( .A(pe_1_2_2_n60), .Z(pe_1_2_2_n56) );
  INV_X1 pe_1_2_2_U6 ( .A(pe_1_2_2_n42), .ZN(pe_1_2_2_n89) );
  INV_X1 pe_1_2_2_U5 ( .A(pe_1_2_2_n40), .ZN(pe_1_2_2_n85) );
  INV_X2 pe_1_2_2_U4 ( .A(n82), .ZN(pe_1_2_2_n72) );
  XOR2_X1 pe_1_2_2_U3 ( .A(pe_1_2_2_int_data_0_), .B(int_data_res_2__2__0_), 
        .Z(pe_1_2_2_n1) );
  DFFR_X1 pe_1_2_2_int_q_acc_reg_0_ ( .D(pe_1_2_2_n84), .CK(pe_1_2_2_net6148), 
        .RN(pe_1_2_2_n72), .Q(int_data_res_2__2__0_), .QN(pe_1_2_2_n3) );
  DFFR_X1 pe_1_2_2_int_q_reg_v_reg_0__0_ ( .D(int_data_y_3__2__0_), .CK(
        pe_1_2_2_net6118), .RN(pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_v[20]) );
  DFFR_X1 pe_1_2_2_int_q_reg_v_reg_0__1_ ( .D(int_data_y_3__2__1_), .CK(
        pe_1_2_2_net6118), .RN(pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_v[21]) );
  DFFR_X1 pe_1_2_2_int_q_reg_v_reg_0__2_ ( .D(int_data_y_3__2__2_), .CK(
        pe_1_2_2_net6118), .RN(pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_v[22]) );
  DFFR_X1 pe_1_2_2_int_q_reg_v_reg_0__3_ ( .D(int_data_y_3__2__3_), .CK(
        pe_1_2_2_net6118), .RN(pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_v[23]) );
  DFFR_X1 pe_1_2_2_int_q_reg_v_reg_1__0_ ( .D(int_data_y_3__2__0_), .CK(
        pe_1_2_2_net6123), .RN(pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_v[16]) );
  DFFR_X1 pe_1_2_2_int_q_reg_v_reg_1__1_ ( .D(int_data_y_3__2__1_), .CK(
        pe_1_2_2_net6123), .RN(pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_v[17]) );
  DFFR_X1 pe_1_2_2_int_q_reg_v_reg_1__2_ ( .D(int_data_y_3__2__2_), .CK(
        pe_1_2_2_net6123), .RN(pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_v[18]) );
  DFFR_X1 pe_1_2_2_int_q_reg_v_reg_1__3_ ( .D(int_data_y_3__2__3_), .CK(
        pe_1_2_2_net6123), .RN(pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_v[19]) );
  DFFR_X1 pe_1_2_2_int_q_reg_v_reg_2__0_ ( .D(int_data_y_3__2__0_), .CK(
        pe_1_2_2_net6128), .RN(pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_v[12]) );
  DFFR_X1 pe_1_2_2_int_q_reg_v_reg_2__1_ ( .D(int_data_y_3__2__1_), .CK(
        pe_1_2_2_net6128), .RN(pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_v[13]) );
  DFFR_X1 pe_1_2_2_int_q_reg_v_reg_2__2_ ( .D(int_data_y_3__2__2_), .CK(
        pe_1_2_2_net6128), .RN(pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_v[14]) );
  DFFR_X1 pe_1_2_2_int_q_reg_v_reg_2__3_ ( .D(int_data_y_3__2__3_), .CK(
        pe_1_2_2_net6128), .RN(pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_v[15]) );
  DFFR_X1 pe_1_2_2_int_q_reg_v_reg_3__0_ ( .D(int_data_y_3__2__0_), .CK(
        pe_1_2_2_net6133), .RN(pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_v[8]) );
  DFFR_X1 pe_1_2_2_int_q_reg_v_reg_3__1_ ( .D(int_data_y_3__2__1_), .CK(
        pe_1_2_2_net6133), .RN(pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_v[9]) );
  DFFR_X1 pe_1_2_2_int_q_reg_v_reg_3__2_ ( .D(int_data_y_3__2__2_), .CK(
        pe_1_2_2_net6133), .RN(pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_v[10]) );
  DFFR_X1 pe_1_2_2_int_q_reg_v_reg_3__3_ ( .D(int_data_y_3__2__3_), .CK(
        pe_1_2_2_net6133), .RN(pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_v[11]) );
  DFFR_X1 pe_1_2_2_int_q_reg_v_reg_4__0_ ( .D(int_data_y_3__2__0_), .CK(
        pe_1_2_2_net6138), .RN(pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_v[4]) );
  DFFR_X1 pe_1_2_2_int_q_reg_v_reg_4__1_ ( .D(int_data_y_3__2__1_), .CK(
        pe_1_2_2_net6138), .RN(pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_v[5]) );
  DFFR_X1 pe_1_2_2_int_q_reg_v_reg_4__2_ ( .D(int_data_y_3__2__2_), .CK(
        pe_1_2_2_net6138), .RN(pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_v[6]) );
  DFFR_X1 pe_1_2_2_int_q_reg_v_reg_4__3_ ( .D(int_data_y_3__2__3_), .CK(
        pe_1_2_2_net6138), .RN(pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_v[7]) );
  DFFR_X1 pe_1_2_2_int_q_reg_v_reg_5__0_ ( .D(int_data_y_3__2__0_), .CK(
        pe_1_2_2_net6143), .RN(pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_v[0]) );
  DFFR_X1 pe_1_2_2_int_q_reg_v_reg_5__1_ ( .D(int_data_y_3__2__1_), .CK(
        pe_1_2_2_net6143), .RN(pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_v[1]) );
  DFFR_X1 pe_1_2_2_int_q_reg_v_reg_5__2_ ( .D(int_data_y_3__2__2_), .CK(
        pe_1_2_2_net6143), .RN(pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_v[2]) );
  DFFR_X1 pe_1_2_2_int_q_reg_v_reg_5__3_ ( .D(int_data_y_3__2__3_), .CK(
        pe_1_2_2_net6143), .RN(pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_2_2_int_q_reg_h_reg_0__0_ ( .D(int_data_x_2__3__0_), .SI(
        int_data_y_3__2__0_), .SE(pe_1_2_2_n65), .CK(pe_1_2_2_net6087), .RN(
        pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_2_2_int_q_reg_h_reg_0__1_ ( .D(int_data_x_2__3__1_), .SI(
        int_data_y_3__2__1_), .SE(pe_1_2_2_n65), .CK(pe_1_2_2_net6087), .RN(
        pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_2_2_int_q_reg_h_reg_0__2_ ( .D(int_data_x_2__3__2_), .SI(
        int_data_y_3__2__2_), .SE(pe_1_2_2_n65), .CK(pe_1_2_2_net6087), .RN(
        pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_2_2_int_q_reg_h_reg_0__3_ ( .D(int_data_x_2__3__3_), .SI(
        int_data_y_3__2__3_), .SE(pe_1_2_2_n65), .CK(pe_1_2_2_net6087), .RN(
        pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_2_2_int_q_reg_h_reg_1__0_ ( .D(int_data_x_2__3__0_), .SI(
        int_data_y_3__2__0_), .SE(pe_1_2_2_n65), .CK(pe_1_2_2_net6093), .RN(
        pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_2_2_int_q_reg_h_reg_1__1_ ( .D(int_data_x_2__3__1_), .SI(
        int_data_y_3__2__1_), .SE(pe_1_2_2_n65), .CK(pe_1_2_2_net6093), .RN(
        pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_2_2_int_q_reg_h_reg_1__2_ ( .D(int_data_x_2__3__2_), .SI(
        int_data_y_3__2__2_), .SE(pe_1_2_2_n65), .CK(pe_1_2_2_net6093), .RN(
        pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_2_2_int_q_reg_h_reg_1__3_ ( .D(int_data_x_2__3__3_), .SI(
        int_data_y_3__2__3_), .SE(pe_1_2_2_n65), .CK(pe_1_2_2_net6093), .RN(
        pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_2_2_int_q_reg_h_reg_2__0_ ( .D(int_data_x_2__3__0_), .SI(
        int_data_y_3__2__0_), .SE(pe_1_2_2_n65), .CK(pe_1_2_2_net6098), .RN(
        pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_2_2_int_q_reg_h_reg_2__1_ ( .D(int_data_x_2__3__1_), .SI(
        int_data_y_3__2__1_), .SE(pe_1_2_2_n65), .CK(pe_1_2_2_net6098), .RN(
        pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_2_2_int_q_reg_h_reg_2__2_ ( .D(int_data_x_2__3__2_), .SI(
        int_data_y_3__2__2_), .SE(pe_1_2_2_n65), .CK(pe_1_2_2_net6098), .RN(
        pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_2_2_int_q_reg_h_reg_2__3_ ( .D(int_data_x_2__3__3_), .SI(
        int_data_y_3__2__3_), .SE(pe_1_2_2_n65), .CK(pe_1_2_2_net6098), .RN(
        pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_2_2_int_q_reg_h_reg_3__0_ ( .D(int_data_x_2__3__0_), .SI(
        int_data_y_3__2__0_), .SE(pe_1_2_2_n65), .CK(pe_1_2_2_net6103), .RN(
        pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_2_2_int_q_reg_h_reg_3__1_ ( .D(int_data_x_2__3__1_), .SI(
        int_data_y_3__2__1_), .SE(pe_1_2_2_n65), .CK(pe_1_2_2_net6103), .RN(
        pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_2_2_int_q_reg_h_reg_3__2_ ( .D(int_data_x_2__3__2_), .SI(
        int_data_y_3__2__2_), .SE(pe_1_2_2_n65), .CK(pe_1_2_2_net6103), .RN(
        pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_2_2_int_q_reg_h_reg_3__3_ ( .D(int_data_x_2__3__3_), .SI(
        int_data_y_3__2__3_), .SE(pe_1_2_2_n65), .CK(pe_1_2_2_net6103), .RN(
        pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_2_2_int_q_reg_h_reg_4__0_ ( .D(int_data_x_2__3__0_), .SI(
        int_data_y_3__2__0_), .SE(pe_1_2_2_n66), .CK(pe_1_2_2_net6108), .RN(
        pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_2_2_int_q_reg_h_reg_4__1_ ( .D(int_data_x_2__3__1_), .SI(
        int_data_y_3__2__1_), .SE(pe_1_2_2_n66), .CK(pe_1_2_2_net6108), .RN(
        pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_2_2_int_q_reg_h_reg_4__2_ ( .D(int_data_x_2__3__2_), .SI(
        int_data_y_3__2__2_), .SE(pe_1_2_2_n66), .CK(pe_1_2_2_net6108), .RN(
        pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_2_2_int_q_reg_h_reg_4__3_ ( .D(int_data_x_2__3__3_), .SI(
        int_data_y_3__2__3_), .SE(pe_1_2_2_n66), .CK(pe_1_2_2_net6108), .RN(
        pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_2_2_int_q_reg_h_reg_5__0_ ( .D(int_data_x_2__3__0_), .SI(
        int_data_y_3__2__0_), .SE(pe_1_2_2_n66), .CK(pe_1_2_2_net6113), .RN(
        pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_2_2_int_q_reg_h_reg_5__1_ ( .D(int_data_x_2__3__1_), .SI(
        int_data_y_3__2__1_), .SE(pe_1_2_2_n66), .CK(pe_1_2_2_net6113), .RN(
        pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_2_2_int_q_reg_h_reg_5__2_ ( .D(int_data_x_2__3__2_), .SI(
        int_data_y_3__2__2_), .SE(pe_1_2_2_n66), .CK(pe_1_2_2_net6113), .RN(
        pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_2_2_int_q_reg_h_reg_5__3_ ( .D(int_data_x_2__3__3_), .SI(
        int_data_y_3__2__3_), .SE(pe_1_2_2_n66), .CK(pe_1_2_2_net6113), .RN(
        pe_1_2_2_n72), .Q(pe_1_2_2_int_q_reg_h[3]) );
  FA_X1 pe_1_2_2_sub_81_U2_7 ( .A(int_data_res_2__2__7_), .B(pe_1_2_2_n76), 
        .CI(pe_1_2_2_sub_81_carry[7]), .S(pe_1_2_2_N77) );
  FA_X1 pe_1_2_2_sub_81_U2_6 ( .A(int_data_res_2__2__6_), .B(pe_1_2_2_n76), 
        .CI(pe_1_2_2_sub_81_carry[6]), .CO(pe_1_2_2_sub_81_carry[7]), .S(
        pe_1_2_2_N76) );
  FA_X1 pe_1_2_2_sub_81_U2_5 ( .A(int_data_res_2__2__5_), .B(pe_1_2_2_n76), 
        .CI(pe_1_2_2_sub_81_carry[5]), .CO(pe_1_2_2_sub_81_carry[6]), .S(
        pe_1_2_2_N75) );
  FA_X1 pe_1_2_2_sub_81_U2_4 ( .A(int_data_res_2__2__4_), .B(pe_1_2_2_n76), 
        .CI(pe_1_2_2_sub_81_carry[4]), .CO(pe_1_2_2_sub_81_carry[5]), .S(
        pe_1_2_2_N74) );
  FA_X1 pe_1_2_2_sub_81_U2_3 ( .A(int_data_res_2__2__3_), .B(pe_1_2_2_n76), 
        .CI(pe_1_2_2_sub_81_carry[3]), .CO(pe_1_2_2_sub_81_carry[4]), .S(
        pe_1_2_2_N73) );
  FA_X1 pe_1_2_2_sub_81_U2_2 ( .A(int_data_res_2__2__2_), .B(pe_1_2_2_n75), 
        .CI(pe_1_2_2_sub_81_carry[2]), .CO(pe_1_2_2_sub_81_carry[3]), .S(
        pe_1_2_2_N72) );
  FA_X1 pe_1_2_2_sub_81_U2_1 ( .A(int_data_res_2__2__1_), .B(pe_1_2_2_n74), 
        .CI(pe_1_2_2_sub_81_carry[1]), .CO(pe_1_2_2_sub_81_carry[2]), .S(
        pe_1_2_2_N71) );
  FA_X1 pe_1_2_2_add_83_U1_7 ( .A(int_data_res_2__2__7_), .B(
        pe_1_2_2_int_data_3_), .CI(pe_1_2_2_add_83_carry[7]), .S(pe_1_2_2_N85)
         );
  FA_X1 pe_1_2_2_add_83_U1_6 ( .A(int_data_res_2__2__6_), .B(
        pe_1_2_2_int_data_3_), .CI(pe_1_2_2_add_83_carry[6]), .CO(
        pe_1_2_2_add_83_carry[7]), .S(pe_1_2_2_N84) );
  FA_X1 pe_1_2_2_add_83_U1_5 ( .A(int_data_res_2__2__5_), .B(
        pe_1_2_2_int_data_3_), .CI(pe_1_2_2_add_83_carry[5]), .CO(
        pe_1_2_2_add_83_carry[6]), .S(pe_1_2_2_N83) );
  FA_X1 pe_1_2_2_add_83_U1_4 ( .A(int_data_res_2__2__4_), .B(
        pe_1_2_2_int_data_3_), .CI(pe_1_2_2_add_83_carry[4]), .CO(
        pe_1_2_2_add_83_carry[5]), .S(pe_1_2_2_N82) );
  FA_X1 pe_1_2_2_add_83_U1_3 ( .A(int_data_res_2__2__3_), .B(
        pe_1_2_2_int_data_3_), .CI(pe_1_2_2_add_83_carry[3]), .CO(
        pe_1_2_2_add_83_carry[4]), .S(pe_1_2_2_N81) );
  FA_X1 pe_1_2_2_add_83_U1_2 ( .A(int_data_res_2__2__2_), .B(
        pe_1_2_2_int_data_2_), .CI(pe_1_2_2_add_83_carry[2]), .CO(
        pe_1_2_2_add_83_carry[3]), .S(pe_1_2_2_N80) );
  FA_X1 pe_1_2_2_add_83_U1_1 ( .A(int_data_res_2__2__1_), .B(
        pe_1_2_2_int_data_1_), .CI(pe_1_2_2_n2), .CO(pe_1_2_2_add_83_carry[2]), 
        .S(pe_1_2_2_N79) );
  NAND3_X1 pe_1_2_2_U56 ( .A1(pe_1_2_2_n60), .A2(pe_1_2_2_n43), .A3(
        pe_1_2_2_n62), .ZN(pe_1_2_2_n40) );
  NAND3_X1 pe_1_2_2_U55 ( .A1(pe_1_2_2_n43), .A2(pe_1_2_2_n61), .A3(
        pe_1_2_2_n62), .ZN(pe_1_2_2_n39) );
  NAND3_X1 pe_1_2_2_U54 ( .A1(pe_1_2_2_n43), .A2(pe_1_2_2_n63), .A3(
        pe_1_2_2_n60), .ZN(pe_1_2_2_n38) );
  NAND3_X1 pe_1_2_2_U53 ( .A1(pe_1_2_2_n61), .A2(pe_1_2_2_n63), .A3(
        pe_1_2_2_n43), .ZN(pe_1_2_2_n37) );
  DFFR_X1 pe_1_2_2_int_q_acc_reg_6_ ( .D(pe_1_2_2_n78), .CK(pe_1_2_2_net6148), 
        .RN(pe_1_2_2_n71), .Q(int_data_res_2__2__6_) );
  DFFR_X1 pe_1_2_2_int_q_acc_reg_5_ ( .D(pe_1_2_2_n79), .CK(pe_1_2_2_net6148), 
        .RN(pe_1_2_2_n71), .Q(int_data_res_2__2__5_) );
  DFFR_X1 pe_1_2_2_int_q_acc_reg_4_ ( .D(pe_1_2_2_n80), .CK(pe_1_2_2_net6148), 
        .RN(pe_1_2_2_n71), .Q(int_data_res_2__2__4_) );
  DFFR_X1 pe_1_2_2_int_q_acc_reg_3_ ( .D(pe_1_2_2_n81), .CK(pe_1_2_2_net6148), 
        .RN(pe_1_2_2_n71), .Q(int_data_res_2__2__3_) );
  DFFR_X1 pe_1_2_2_int_q_acc_reg_2_ ( .D(pe_1_2_2_n82), .CK(pe_1_2_2_net6148), 
        .RN(pe_1_2_2_n71), .Q(int_data_res_2__2__2_) );
  DFFR_X1 pe_1_2_2_int_q_acc_reg_1_ ( .D(pe_1_2_2_n83), .CK(pe_1_2_2_net6148), 
        .RN(pe_1_2_2_n71), .Q(int_data_res_2__2__1_) );
  DFFR_X1 pe_1_2_2_int_q_acc_reg_7_ ( .D(pe_1_2_2_n77), .CK(pe_1_2_2_net6148), 
        .RN(pe_1_2_2_n71), .Q(int_data_res_2__2__7_) );
  CLKGATETST_X1 pe_1_2_2_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_2_2_n88), .SE(1'b0), .GCK(pe_1_2_2_net6087) );
  CLKGATETST_X1 pe_1_2_2_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_2_2_n87), .SE(1'b0), .GCK(pe_1_2_2_net6093) );
  CLKGATETST_X1 pe_1_2_2_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_2_2_n86), .SE(1'b0), .GCK(pe_1_2_2_net6098) );
  CLKGATETST_X1 pe_1_2_2_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_2_2_n85), .SE(1'b0), .GCK(pe_1_2_2_net6103) );
  CLKGATETST_X1 pe_1_2_2_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_2_2_n90), .SE(1'b0), .GCK(pe_1_2_2_net6108) );
  CLKGATETST_X1 pe_1_2_2_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_2_2_n89), .SE(1'b0), .GCK(pe_1_2_2_net6113) );
  CLKGATETST_X1 pe_1_2_2_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_2_2_N64), .SE(1'b0), .GCK(pe_1_2_2_net6118) );
  CLKGATETST_X1 pe_1_2_2_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_2_2_N63), .SE(1'b0), .GCK(pe_1_2_2_net6123) );
  CLKGATETST_X1 pe_1_2_2_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_2_2_N62), .SE(1'b0), .GCK(pe_1_2_2_net6128) );
  CLKGATETST_X1 pe_1_2_2_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_2_2_N61), .SE(1'b0), .GCK(pe_1_2_2_net6133) );
  CLKGATETST_X1 pe_1_2_2_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_2_2_N60), .SE(1'b0), .GCK(pe_1_2_2_net6138) );
  CLKGATETST_X1 pe_1_2_2_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_2_2_N59), .SE(1'b0), .GCK(pe_1_2_2_net6143) );
  CLKGATETST_X1 pe_1_2_2_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_2_2_N90), .SE(1'b0), .GCK(pe_1_2_2_net6148) );
  CLKBUF_X1 pe_1_2_3_U112 ( .A(pe_1_2_3_n72), .Z(pe_1_2_3_n71) );
  INV_X1 pe_1_2_3_U111 ( .A(n74), .ZN(pe_1_2_3_n70) );
  INV_X1 pe_1_2_3_U110 ( .A(n66), .ZN(pe_1_2_3_n69) );
  INV_X1 pe_1_2_3_U109 ( .A(n66), .ZN(pe_1_2_3_n68) );
  INV_X1 pe_1_2_3_U108 ( .A(n66), .ZN(pe_1_2_3_n67) );
  INV_X1 pe_1_2_3_U107 ( .A(pe_1_2_3_n69), .ZN(pe_1_2_3_n66) );
  INV_X1 pe_1_2_3_U106 ( .A(pe_1_2_3_n63), .ZN(pe_1_2_3_n62) );
  INV_X1 pe_1_2_3_U105 ( .A(pe_1_2_3_n61), .ZN(pe_1_2_3_n60) );
  INV_X1 pe_1_2_3_U104 ( .A(n26), .ZN(pe_1_2_3_n59) );
  INV_X1 pe_1_2_3_U103 ( .A(pe_1_2_3_n59), .ZN(pe_1_2_3_n58) );
  INV_X1 pe_1_2_3_U102 ( .A(n18), .ZN(pe_1_2_3_n57) );
  MUX2_X1 pe_1_2_3_U101 ( .A(pe_1_2_3_n54), .B(pe_1_2_3_n51), .S(n46), .Z(
        int_data_x_2__3__3_) );
  MUX2_X1 pe_1_2_3_U100 ( .A(pe_1_2_3_n53), .B(pe_1_2_3_n52), .S(pe_1_2_3_n62), 
        .Z(pe_1_2_3_n54) );
  MUX2_X1 pe_1_2_3_U99 ( .A(pe_1_2_3_int_q_reg_h[23]), .B(
        pe_1_2_3_int_q_reg_h[19]), .S(pe_1_2_3_n56), .Z(pe_1_2_3_n53) );
  MUX2_X1 pe_1_2_3_U98 ( .A(pe_1_2_3_int_q_reg_h[15]), .B(
        pe_1_2_3_int_q_reg_h[11]), .S(pe_1_2_3_n56), .Z(pe_1_2_3_n52) );
  MUX2_X1 pe_1_2_3_U97 ( .A(pe_1_2_3_int_q_reg_h[7]), .B(
        pe_1_2_3_int_q_reg_h[3]), .S(pe_1_2_3_n56), .Z(pe_1_2_3_n51) );
  MUX2_X1 pe_1_2_3_U96 ( .A(pe_1_2_3_n50), .B(pe_1_2_3_n47), .S(n46), .Z(
        int_data_x_2__3__2_) );
  MUX2_X1 pe_1_2_3_U95 ( .A(pe_1_2_3_n49), .B(pe_1_2_3_n48), .S(pe_1_2_3_n62), 
        .Z(pe_1_2_3_n50) );
  MUX2_X1 pe_1_2_3_U94 ( .A(pe_1_2_3_int_q_reg_h[22]), .B(
        pe_1_2_3_int_q_reg_h[18]), .S(pe_1_2_3_n56), .Z(pe_1_2_3_n49) );
  MUX2_X1 pe_1_2_3_U93 ( .A(pe_1_2_3_int_q_reg_h[14]), .B(
        pe_1_2_3_int_q_reg_h[10]), .S(pe_1_2_3_n56), .Z(pe_1_2_3_n48) );
  MUX2_X1 pe_1_2_3_U92 ( .A(pe_1_2_3_int_q_reg_h[6]), .B(
        pe_1_2_3_int_q_reg_h[2]), .S(pe_1_2_3_n56), .Z(pe_1_2_3_n47) );
  MUX2_X1 pe_1_2_3_U91 ( .A(pe_1_2_3_n46), .B(pe_1_2_3_n24), .S(n46), .Z(
        int_data_x_2__3__1_) );
  MUX2_X1 pe_1_2_3_U90 ( .A(pe_1_2_3_n45), .B(pe_1_2_3_n25), .S(pe_1_2_3_n62), 
        .Z(pe_1_2_3_n46) );
  MUX2_X1 pe_1_2_3_U89 ( .A(pe_1_2_3_int_q_reg_h[21]), .B(
        pe_1_2_3_int_q_reg_h[17]), .S(pe_1_2_3_n56), .Z(pe_1_2_3_n45) );
  MUX2_X1 pe_1_2_3_U88 ( .A(pe_1_2_3_int_q_reg_h[13]), .B(
        pe_1_2_3_int_q_reg_h[9]), .S(pe_1_2_3_n56), .Z(pe_1_2_3_n25) );
  MUX2_X1 pe_1_2_3_U87 ( .A(pe_1_2_3_int_q_reg_h[5]), .B(
        pe_1_2_3_int_q_reg_h[1]), .S(pe_1_2_3_n56), .Z(pe_1_2_3_n24) );
  MUX2_X1 pe_1_2_3_U86 ( .A(pe_1_2_3_n23), .B(pe_1_2_3_n20), .S(n46), .Z(
        int_data_x_2__3__0_) );
  MUX2_X1 pe_1_2_3_U85 ( .A(pe_1_2_3_n22), .B(pe_1_2_3_n21), .S(pe_1_2_3_n62), 
        .Z(pe_1_2_3_n23) );
  MUX2_X1 pe_1_2_3_U84 ( .A(pe_1_2_3_int_q_reg_h[20]), .B(
        pe_1_2_3_int_q_reg_h[16]), .S(pe_1_2_3_n56), .Z(pe_1_2_3_n22) );
  MUX2_X1 pe_1_2_3_U83 ( .A(pe_1_2_3_int_q_reg_h[12]), .B(
        pe_1_2_3_int_q_reg_h[8]), .S(pe_1_2_3_n56), .Z(pe_1_2_3_n21) );
  MUX2_X1 pe_1_2_3_U82 ( .A(pe_1_2_3_int_q_reg_h[4]), .B(
        pe_1_2_3_int_q_reg_h[0]), .S(pe_1_2_3_n56), .Z(pe_1_2_3_n20) );
  MUX2_X1 pe_1_2_3_U81 ( .A(pe_1_2_3_n19), .B(pe_1_2_3_n16), .S(n46), .Z(
        int_data_y_2__3__3_) );
  MUX2_X1 pe_1_2_3_U80 ( .A(pe_1_2_3_n18), .B(pe_1_2_3_n17), .S(pe_1_2_3_n62), 
        .Z(pe_1_2_3_n19) );
  MUX2_X1 pe_1_2_3_U79 ( .A(pe_1_2_3_int_q_reg_v[23]), .B(
        pe_1_2_3_int_q_reg_v[19]), .S(pe_1_2_3_n55), .Z(pe_1_2_3_n18) );
  MUX2_X1 pe_1_2_3_U78 ( .A(pe_1_2_3_int_q_reg_v[15]), .B(
        pe_1_2_3_int_q_reg_v[11]), .S(pe_1_2_3_n55), .Z(pe_1_2_3_n17) );
  MUX2_X1 pe_1_2_3_U77 ( .A(pe_1_2_3_int_q_reg_v[7]), .B(
        pe_1_2_3_int_q_reg_v[3]), .S(pe_1_2_3_n55), .Z(pe_1_2_3_n16) );
  MUX2_X1 pe_1_2_3_U76 ( .A(pe_1_2_3_n15), .B(pe_1_2_3_n12), .S(n46), .Z(
        int_data_y_2__3__2_) );
  MUX2_X1 pe_1_2_3_U75 ( .A(pe_1_2_3_n14), .B(pe_1_2_3_n13), .S(pe_1_2_3_n62), 
        .Z(pe_1_2_3_n15) );
  MUX2_X1 pe_1_2_3_U74 ( .A(pe_1_2_3_int_q_reg_v[22]), .B(
        pe_1_2_3_int_q_reg_v[18]), .S(pe_1_2_3_n55), .Z(pe_1_2_3_n14) );
  MUX2_X1 pe_1_2_3_U73 ( .A(pe_1_2_3_int_q_reg_v[14]), .B(
        pe_1_2_3_int_q_reg_v[10]), .S(pe_1_2_3_n55), .Z(pe_1_2_3_n13) );
  MUX2_X1 pe_1_2_3_U72 ( .A(pe_1_2_3_int_q_reg_v[6]), .B(
        pe_1_2_3_int_q_reg_v[2]), .S(pe_1_2_3_n55), .Z(pe_1_2_3_n12) );
  MUX2_X1 pe_1_2_3_U71 ( .A(pe_1_2_3_n11), .B(pe_1_2_3_n8), .S(n46), .Z(
        int_data_y_2__3__1_) );
  MUX2_X1 pe_1_2_3_U70 ( .A(pe_1_2_3_n10), .B(pe_1_2_3_n9), .S(pe_1_2_3_n62), 
        .Z(pe_1_2_3_n11) );
  MUX2_X1 pe_1_2_3_U69 ( .A(pe_1_2_3_int_q_reg_v[21]), .B(
        pe_1_2_3_int_q_reg_v[17]), .S(pe_1_2_3_n55), .Z(pe_1_2_3_n10) );
  MUX2_X1 pe_1_2_3_U68 ( .A(pe_1_2_3_int_q_reg_v[13]), .B(
        pe_1_2_3_int_q_reg_v[9]), .S(pe_1_2_3_n55), .Z(pe_1_2_3_n9) );
  MUX2_X1 pe_1_2_3_U67 ( .A(pe_1_2_3_int_q_reg_v[5]), .B(
        pe_1_2_3_int_q_reg_v[1]), .S(pe_1_2_3_n55), .Z(pe_1_2_3_n8) );
  MUX2_X1 pe_1_2_3_U66 ( .A(pe_1_2_3_n7), .B(pe_1_2_3_n4), .S(n46), .Z(
        int_data_y_2__3__0_) );
  MUX2_X1 pe_1_2_3_U65 ( .A(pe_1_2_3_n6), .B(pe_1_2_3_n5), .S(pe_1_2_3_n62), 
        .Z(pe_1_2_3_n7) );
  MUX2_X1 pe_1_2_3_U64 ( .A(pe_1_2_3_int_q_reg_v[20]), .B(
        pe_1_2_3_int_q_reg_v[16]), .S(pe_1_2_3_n55), .Z(pe_1_2_3_n6) );
  MUX2_X1 pe_1_2_3_U63 ( .A(pe_1_2_3_int_q_reg_v[12]), .B(
        pe_1_2_3_int_q_reg_v[8]), .S(pe_1_2_3_n55), .Z(pe_1_2_3_n5) );
  MUX2_X1 pe_1_2_3_U62 ( .A(pe_1_2_3_int_q_reg_v[4]), .B(
        pe_1_2_3_int_q_reg_v[0]), .S(pe_1_2_3_n55), .Z(pe_1_2_3_n4) );
  AOI222_X1 pe_1_2_3_U61 ( .A1(int_data_res_3__3__2_), .A2(pe_1_2_3_n64), .B1(
        pe_1_2_3_N80), .B2(pe_1_2_3_n27), .C1(pe_1_2_3_N72), .C2(pe_1_2_3_n28), 
        .ZN(pe_1_2_3_n33) );
  INV_X1 pe_1_2_3_U60 ( .A(pe_1_2_3_n33), .ZN(pe_1_2_3_n82) );
  AOI222_X1 pe_1_2_3_U59 ( .A1(int_data_res_3__3__6_), .A2(pe_1_2_3_n64), .B1(
        pe_1_2_3_N84), .B2(pe_1_2_3_n27), .C1(pe_1_2_3_N76), .C2(pe_1_2_3_n28), 
        .ZN(pe_1_2_3_n29) );
  INV_X1 pe_1_2_3_U58 ( .A(pe_1_2_3_n29), .ZN(pe_1_2_3_n78) );
  XNOR2_X1 pe_1_2_3_U57 ( .A(pe_1_2_3_n73), .B(int_data_res_2__3__0_), .ZN(
        pe_1_2_3_N70) );
  AOI222_X1 pe_1_2_3_U52 ( .A1(int_data_res_3__3__0_), .A2(pe_1_2_3_n64), .B1(
        pe_1_2_3_n1), .B2(pe_1_2_3_n27), .C1(pe_1_2_3_N70), .C2(pe_1_2_3_n28), 
        .ZN(pe_1_2_3_n35) );
  INV_X1 pe_1_2_3_U51 ( .A(pe_1_2_3_n35), .ZN(pe_1_2_3_n84) );
  AOI222_X1 pe_1_2_3_U50 ( .A1(int_data_res_3__3__1_), .A2(pe_1_2_3_n64), .B1(
        pe_1_2_3_N79), .B2(pe_1_2_3_n27), .C1(pe_1_2_3_N71), .C2(pe_1_2_3_n28), 
        .ZN(pe_1_2_3_n34) );
  INV_X1 pe_1_2_3_U49 ( .A(pe_1_2_3_n34), .ZN(pe_1_2_3_n83) );
  AOI222_X1 pe_1_2_3_U48 ( .A1(int_data_res_3__3__3_), .A2(pe_1_2_3_n64), .B1(
        pe_1_2_3_N81), .B2(pe_1_2_3_n27), .C1(pe_1_2_3_N73), .C2(pe_1_2_3_n28), 
        .ZN(pe_1_2_3_n32) );
  INV_X1 pe_1_2_3_U47 ( .A(pe_1_2_3_n32), .ZN(pe_1_2_3_n81) );
  AOI222_X1 pe_1_2_3_U46 ( .A1(int_data_res_3__3__4_), .A2(pe_1_2_3_n64), .B1(
        pe_1_2_3_N82), .B2(pe_1_2_3_n27), .C1(pe_1_2_3_N74), .C2(pe_1_2_3_n28), 
        .ZN(pe_1_2_3_n31) );
  INV_X1 pe_1_2_3_U45 ( .A(pe_1_2_3_n31), .ZN(pe_1_2_3_n80) );
  AOI222_X1 pe_1_2_3_U44 ( .A1(int_data_res_3__3__5_), .A2(pe_1_2_3_n64), .B1(
        pe_1_2_3_N83), .B2(pe_1_2_3_n27), .C1(pe_1_2_3_N75), .C2(pe_1_2_3_n28), 
        .ZN(pe_1_2_3_n30) );
  INV_X1 pe_1_2_3_U43 ( .A(pe_1_2_3_n30), .ZN(pe_1_2_3_n79) );
  NAND2_X1 pe_1_2_3_U42 ( .A1(pe_1_2_3_int_data_0_), .A2(pe_1_2_3_n3), .ZN(
        pe_1_2_3_sub_81_carry[1]) );
  INV_X1 pe_1_2_3_U41 ( .A(pe_1_2_3_int_data_1_), .ZN(pe_1_2_3_n74) );
  INV_X1 pe_1_2_3_U40 ( .A(pe_1_2_3_int_data_2_), .ZN(pe_1_2_3_n75) );
  AND2_X1 pe_1_2_3_U39 ( .A1(pe_1_2_3_int_data_0_), .A2(int_data_res_2__3__0_), 
        .ZN(pe_1_2_3_n2) );
  AOI222_X1 pe_1_2_3_U38 ( .A1(pe_1_2_3_n64), .A2(int_data_res_3__3__7_), .B1(
        pe_1_2_3_N85), .B2(pe_1_2_3_n27), .C1(pe_1_2_3_N77), .C2(pe_1_2_3_n28), 
        .ZN(pe_1_2_3_n26) );
  INV_X1 pe_1_2_3_U37 ( .A(pe_1_2_3_n26), .ZN(pe_1_2_3_n77) );
  NOR3_X1 pe_1_2_3_U36 ( .A1(pe_1_2_3_n59), .A2(pe_1_2_3_n65), .A3(int_ckg[44]), .ZN(pe_1_2_3_n36) );
  OR2_X1 pe_1_2_3_U35 ( .A1(pe_1_2_3_n36), .A2(pe_1_2_3_n64), .ZN(pe_1_2_3_N90) );
  INV_X1 pe_1_2_3_U34 ( .A(n38), .ZN(pe_1_2_3_n63) );
  AND2_X1 pe_1_2_3_U33 ( .A1(int_data_x_2__3__2_), .A2(pe_1_2_3_n58), .ZN(
        pe_1_2_3_int_data_2_) );
  AND2_X1 pe_1_2_3_U32 ( .A1(int_data_x_2__3__1_), .A2(pe_1_2_3_n58), .ZN(
        pe_1_2_3_int_data_1_) );
  AND2_X1 pe_1_2_3_U31 ( .A1(int_data_x_2__3__3_), .A2(pe_1_2_3_n58), .ZN(
        pe_1_2_3_int_data_3_) );
  BUF_X1 pe_1_2_3_U30 ( .A(n60), .Z(pe_1_2_3_n64) );
  INV_X1 pe_1_2_3_U29 ( .A(n32), .ZN(pe_1_2_3_n61) );
  AND2_X1 pe_1_2_3_U28 ( .A1(int_data_x_2__3__0_), .A2(pe_1_2_3_n58), .ZN(
        pe_1_2_3_int_data_0_) );
  NAND2_X1 pe_1_2_3_U27 ( .A1(pe_1_2_3_n44), .A2(pe_1_2_3_n61), .ZN(
        pe_1_2_3_n41) );
  AND3_X1 pe_1_2_3_U26 ( .A1(n74), .A2(pe_1_2_3_n63), .A3(n46), .ZN(
        pe_1_2_3_n44) );
  INV_X1 pe_1_2_3_U25 ( .A(pe_1_2_3_int_data_3_), .ZN(pe_1_2_3_n76) );
  NOR2_X1 pe_1_2_3_U24 ( .A1(pe_1_2_3_n70), .A2(n46), .ZN(pe_1_2_3_n43) );
  NOR2_X1 pe_1_2_3_U23 ( .A1(pe_1_2_3_n57), .A2(pe_1_2_3_n64), .ZN(
        pe_1_2_3_n28) );
  NOR2_X1 pe_1_2_3_U22 ( .A1(n18), .A2(pe_1_2_3_n64), .ZN(pe_1_2_3_n27) );
  INV_X1 pe_1_2_3_U21 ( .A(pe_1_2_3_int_data_0_), .ZN(pe_1_2_3_n73) );
  INV_X1 pe_1_2_3_U20 ( .A(pe_1_2_3_n41), .ZN(pe_1_2_3_n90) );
  INV_X1 pe_1_2_3_U19 ( .A(pe_1_2_3_n37), .ZN(pe_1_2_3_n88) );
  INV_X1 pe_1_2_3_U18 ( .A(pe_1_2_3_n38), .ZN(pe_1_2_3_n87) );
  INV_X1 pe_1_2_3_U17 ( .A(pe_1_2_3_n39), .ZN(pe_1_2_3_n86) );
  NOR2_X1 pe_1_2_3_U16 ( .A1(pe_1_2_3_n68), .A2(pe_1_2_3_n42), .ZN(
        pe_1_2_3_N59) );
  NOR2_X1 pe_1_2_3_U15 ( .A1(pe_1_2_3_n68), .A2(pe_1_2_3_n41), .ZN(
        pe_1_2_3_N60) );
  NOR2_X1 pe_1_2_3_U14 ( .A1(pe_1_2_3_n68), .A2(pe_1_2_3_n38), .ZN(
        pe_1_2_3_N63) );
  NOR2_X1 pe_1_2_3_U13 ( .A1(pe_1_2_3_n67), .A2(pe_1_2_3_n40), .ZN(
        pe_1_2_3_N61) );
  NOR2_X1 pe_1_2_3_U12 ( .A1(pe_1_2_3_n67), .A2(pe_1_2_3_n39), .ZN(
        pe_1_2_3_N62) );
  NOR2_X1 pe_1_2_3_U11 ( .A1(pe_1_2_3_n37), .A2(pe_1_2_3_n67), .ZN(
        pe_1_2_3_N64) );
  NAND2_X1 pe_1_2_3_U10 ( .A1(pe_1_2_3_n44), .A2(pe_1_2_3_n60), .ZN(
        pe_1_2_3_n42) );
  BUF_X1 pe_1_2_3_U9 ( .A(pe_1_2_3_n60), .Z(pe_1_2_3_n55) );
  INV_X1 pe_1_2_3_U8 ( .A(pe_1_2_3_n69), .ZN(pe_1_2_3_n65) );
  BUF_X1 pe_1_2_3_U7 ( .A(pe_1_2_3_n60), .Z(pe_1_2_3_n56) );
  INV_X1 pe_1_2_3_U6 ( .A(pe_1_2_3_n42), .ZN(pe_1_2_3_n89) );
  INV_X1 pe_1_2_3_U5 ( .A(pe_1_2_3_n40), .ZN(pe_1_2_3_n85) );
  INV_X2 pe_1_2_3_U4 ( .A(n82), .ZN(pe_1_2_3_n72) );
  XOR2_X1 pe_1_2_3_U3 ( .A(pe_1_2_3_int_data_0_), .B(int_data_res_2__3__0_), 
        .Z(pe_1_2_3_n1) );
  DFFR_X1 pe_1_2_3_int_q_acc_reg_0_ ( .D(pe_1_2_3_n84), .CK(pe_1_2_3_net6070), 
        .RN(pe_1_2_3_n72), .Q(int_data_res_2__3__0_), .QN(pe_1_2_3_n3) );
  DFFR_X1 pe_1_2_3_int_q_reg_v_reg_0__0_ ( .D(int_data_y_3__3__0_), .CK(
        pe_1_2_3_net6040), .RN(pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_v[20]) );
  DFFR_X1 pe_1_2_3_int_q_reg_v_reg_0__1_ ( .D(int_data_y_3__3__1_), .CK(
        pe_1_2_3_net6040), .RN(pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_v[21]) );
  DFFR_X1 pe_1_2_3_int_q_reg_v_reg_0__2_ ( .D(int_data_y_3__3__2_), .CK(
        pe_1_2_3_net6040), .RN(pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_v[22]) );
  DFFR_X1 pe_1_2_3_int_q_reg_v_reg_0__3_ ( .D(int_data_y_3__3__3_), .CK(
        pe_1_2_3_net6040), .RN(pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_v[23]) );
  DFFR_X1 pe_1_2_3_int_q_reg_v_reg_1__0_ ( .D(int_data_y_3__3__0_), .CK(
        pe_1_2_3_net6045), .RN(pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_v[16]) );
  DFFR_X1 pe_1_2_3_int_q_reg_v_reg_1__1_ ( .D(int_data_y_3__3__1_), .CK(
        pe_1_2_3_net6045), .RN(pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_v[17]) );
  DFFR_X1 pe_1_2_3_int_q_reg_v_reg_1__2_ ( .D(int_data_y_3__3__2_), .CK(
        pe_1_2_3_net6045), .RN(pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_v[18]) );
  DFFR_X1 pe_1_2_3_int_q_reg_v_reg_1__3_ ( .D(int_data_y_3__3__3_), .CK(
        pe_1_2_3_net6045), .RN(pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_v[19]) );
  DFFR_X1 pe_1_2_3_int_q_reg_v_reg_2__0_ ( .D(int_data_y_3__3__0_), .CK(
        pe_1_2_3_net6050), .RN(pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_v[12]) );
  DFFR_X1 pe_1_2_3_int_q_reg_v_reg_2__1_ ( .D(int_data_y_3__3__1_), .CK(
        pe_1_2_3_net6050), .RN(pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_v[13]) );
  DFFR_X1 pe_1_2_3_int_q_reg_v_reg_2__2_ ( .D(int_data_y_3__3__2_), .CK(
        pe_1_2_3_net6050), .RN(pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_v[14]) );
  DFFR_X1 pe_1_2_3_int_q_reg_v_reg_2__3_ ( .D(int_data_y_3__3__3_), .CK(
        pe_1_2_3_net6050), .RN(pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_v[15]) );
  DFFR_X1 pe_1_2_3_int_q_reg_v_reg_3__0_ ( .D(int_data_y_3__3__0_), .CK(
        pe_1_2_3_net6055), .RN(pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_v[8]) );
  DFFR_X1 pe_1_2_3_int_q_reg_v_reg_3__1_ ( .D(int_data_y_3__3__1_), .CK(
        pe_1_2_3_net6055), .RN(pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_v[9]) );
  DFFR_X1 pe_1_2_3_int_q_reg_v_reg_3__2_ ( .D(int_data_y_3__3__2_), .CK(
        pe_1_2_3_net6055), .RN(pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_v[10]) );
  DFFR_X1 pe_1_2_3_int_q_reg_v_reg_3__3_ ( .D(int_data_y_3__3__3_), .CK(
        pe_1_2_3_net6055), .RN(pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_v[11]) );
  DFFR_X1 pe_1_2_3_int_q_reg_v_reg_4__0_ ( .D(int_data_y_3__3__0_), .CK(
        pe_1_2_3_net6060), .RN(pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_v[4]) );
  DFFR_X1 pe_1_2_3_int_q_reg_v_reg_4__1_ ( .D(int_data_y_3__3__1_), .CK(
        pe_1_2_3_net6060), .RN(pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_v[5]) );
  DFFR_X1 pe_1_2_3_int_q_reg_v_reg_4__2_ ( .D(int_data_y_3__3__2_), .CK(
        pe_1_2_3_net6060), .RN(pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_v[6]) );
  DFFR_X1 pe_1_2_3_int_q_reg_v_reg_4__3_ ( .D(int_data_y_3__3__3_), .CK(
        pe_1_2_3_net6060), .RN(pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_v[7]) );
  DFFR_X1 pe_1_2_3_int_q_reg_v_reg_5__0_ ( .D(int_data_y_3__3__0_), .CK(
        pe_1_2_3_net6065), .RN(pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_v[0]) );
  DFFR_X1 pe_1_2_3_int_q_reg_v_reg_5__1_ ( .D(int_data_y_3__3__1_), .CK(
        pe_1_2_3_net6065), .RN(pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_v[1]) );
  DFFR_X1 pe_1_2_3_int_q_reg_v_reg_5__2_ ( .D(int_data_y_3__3__2_), .CK(
        pe_1_2_3_net6065), .RN(pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_v[2]) );
  DFFR_X1 pe_1_2_3_int_q_reg_v_reg_5__3_ ( .D(int_data_y_3__3__3_), .CK(
        pe_1_2_3_net6065), .RN(pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_2_3_int_q_reg_h_reg_0__0_ ( .D(int_data_x_2__4__0_), .SI(
        int_data_y_3__3__0_), .SE(pe_1_2_3_n65), .CK(pe_1_2_3_net6009), .RN(
        pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_2_3_int_q_reg_h_reg_0__1_ ( .D(int_data_x_2__4__1_), .SI(
        int_data_y_3__3__1_), .SE(pe_1_2_3_n65), .CK(pe_1_2_3_net6009), .RN(
        pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_2_3_int_q_reg_h_reg_0__2_ ( .D(int_data_x_2__4__2_), .SI(
        int_data_y_3__3__2_), .SE(pe_1_2_3_n65), .CK(pe_1_2_3_net6009), .RN(
        pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_2_3_int_q_reg_h_reg_0__3_ ( .D(int_data_x_2__4__3_), .SI(
        int_data_y_3__3__3_), .SE(pe_1_2_3_n65), .CK(pe_1_2_3_net6009), .RN(
        pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_2_3_int_q_reg_h_reg_1__0_ ( .D(int_data_x_2__4__0_), .SI(
        int_data_y_3__3__0_), .SE(pe_1_2_3_n65), .CK(pe_1_2_3_net6015), .RN(
        pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_2_3_int_q_reg_h_reg_1__1_ ( .D(int_data_x_2__4__1_), .SI(
        int_data_y_3__3__1_), .SE(pe_1_2_3_n65), .CK(pe_1_2_3_net6015), .RN(
        pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_2_3_int_q_reg_h_reg_1__2_ ( .D(int_data_x_2__4__2_), .SI(
        int_data_y_3__3__2_), .SE(pe_1_2_3_n65), .CK(pe_1_2_3_net6015), .RN(
        pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_2_3_int_q_reg_h_reg_1__3_ ( .D(int_data_x_2__4__3_), .SI(
        int_data_y_3__3__3_), .SE(pe_1_2_3_n65), .CK(pe_1_2_3_net6015), .RN(
        pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_2_3_int_q_reg_h_reg_2__0_ ( .D(int_data_x_2__4__0_), .SI(
        int_data_y_3__3__0_), .SE(pe_1_2_3_n65), .CK(pe_1_2_3_net6020), .RN(
        pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_2_3_int_q_reg_h_reg_2__1_ ( .D(int_data_x_2__4__1_), .SI(
        int_data_y_3__3__1_), .SE(pe_1_2_3_n65), .CK(pe_1_2_3_net6020), .RN(
        pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_2_3_int_q_reg_h_reg_2__2_ ( .D(int_data_x_2__4__2_), .SI(
        int_data_y_3__3__2_), .SE(pe_1_2_3_n65), .CK(pe_1_2_3_net6020), .RN(
        pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_2_3_int_q_reg_h_reg_2__3_ ( .D(int_data_x_2__4__3_), .SI(
        int_data_y_3__3__3_), .SE(pe_1_2_3_n65), .CK(pe_1_2_3_net6020), .RN(
        pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_2_3_int_q_reg_h_reg_3__0_ ( .D(int_data_x_2__4__0_), .SI(
        int_data_y_3__3__0_), .SE(pe_1_2_3_n65), .CK(pe_1_2_3_net6025), .RN(
        pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_2_3_int_q_reg_h_reg_3__1_ ( .D(int_data_x_2__4__1_), .SI(
        int_data_y_3__3__1_), .SE(pe_1_2_3_n65), .CK(pe_1_2_3_net6025), .RN(
        pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_2_3_int_q_reg_h_reg_3__2_ ( .D(int_data_x_2__4__2_), .SI(
        int_data_y_3__3__2_), .SE(pe_1_2_3_n65), .CK(pe_1_2_3_net6025), .RN(
        pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_2_3_int_q_reg_h_reg_3__3_ ( .D(int_data_x_2__4__3_), .SI(
        int_data_y_3__3__3_), .SE(pe_1_2_3_n65), .CK(pe_1_2_3_net6025), .RN(
        pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_2_3_int_q_reg_h_reg_4__0_ ( .D(int_data_x_2__4__0_), .SI(
        int_data_y_3__3__0_), .SE(pe_1_2_3_n66), .CK(pe_1_2_3_net6030), .RN(
        pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_2_3_int_q_reg_h_reg_4__1_ ( .D(int_data_x_2__4__1_), .SI(
        int_data_y_3__3__1_), .SE(pe_1_2_3_n66), .CK(pe_1_2_3_net6030), .RN(
        pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_2_3_int_q_reg_h_reg_4__2_ ( .D(int_data_x_2__4__2_), .SI(
        int_data_y_3__3__2_), .SE(pe_1_2_3_n66), .CK(pe_1_2_3_net6030), .RN(
        pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_2_3_int_q_reg_h_reg_4__3_ ( .D(int_data_x_2__4__3_), .SI(
        int_data_y_3__3__3_), .SE(pe_1_2_3_n66), .CK(pe_1_2_3_net6030), .RN(
        pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_2_3_int_q_reg_h_reg_5__0_ ( .D(int_data_x_2__4__0_), .SI(
        int_data_y_3__3__0_), .SE(pe_1_2_3_n66), .CK(pe_1_2_3_net6035), .RN(
        pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_2_3_int_q_reg_h_reg_5__1_ ( .D(int_data_x_2__4__1_), .SI(
        int_data_y_3__3__1_), .SE(pe_1_2_3_n66), .CK(pe_1_2_3_net6035), .RN(
        pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_2_3_int_q_reg_h_reg_5__2_ ( .D(int_data_x_2__4__2_), .SI(
        int_data_y_3__3__2_), .SE(pe_1_2_3_n66), .CK(pe_1_2_3_net6035), .RN(
        pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_2_3_int_q_reg_h_reg_5__3_ ( .D(int_data_x_2__4__3_), .SI(
        int_data_y_3__3__3_), .SE(pe_1_2_3_n66), .CK(pe_1_2_3_net6035), .RN(
        pe_1_2_3_n72), .Q(pe_1_2_3_int_q_reg_h[3]) );
  FA_X1 pe_1_2_3_sub_81_U2_7 ( .A(int_data_res_2__3__7_), .B(pe_1_2_3_n76), 
        .CI(pe_1_2_3_sub_81_carry[7]), .S(pe_1_2_3_N77) );
  FA_X1 pe_1_2_3_sub_81_U2_6 ( .A(int_data_res_2__3__6_), .B(pe_1_2_3_n76), 
        .CI(pe_1_2_3_sub_81_carry[6]), .CO(pe_1_2_3_sub_81_carry[7]), .S(
        pe_1_2_3_N76) );
  FA_X1 pe_1_2_3_sub_81_U2_5 ( .A(int_data_res_2__3__5_), .B(pe_1_2_3_n76), 
        .CI(pe_1_2_3_sub_81_carry[5]), .CO(pe_1_2_3_sub_81_carry[6]), .S(
        pe_1_2_3_N75) );
  FA_X1 pe_1_2_3_sub_81_U2_4 ( .A(int_data_res_2__3__4_), .B(pe_1_2_3_n76), 
        .CI(pe_1_2_3_sub_81_carry[4]), .CO(pe_1_2_3_sub_81_carry[5]), .S(
        pe_1_2_3_N74) );
  FA_X1 pe_1_2_3_sub_81_U2_3 ( .A(int_data_res_2__3__3_), .B(pe_1_2_3_n76), 
        .CI(pe_1_2_3_sub_81_carry[3]), .CO(pe_1_2_3_sub_81_carry[4]), .S(
        pe_1_2_3_N73) );
  FA_X1 pe_1_2_3_sub_81_U2_2 ( .A(int_data_res_2__3__2_), .B(pe_1_2_3_n75), 
        .CI(pe_1_2_3_sub_81_carry[2]), .CO(pe_1_2_3_sub_81_carry[3]), .S(
        pe_1_2_3_N72) );
  FA_X1 pe_1_2_3_sub_81_U2_1 ( .A(int_data_res_2__3__1_), .B(pe_1_2_3_n74), 
        .CI(pe_1_2_3_sub_81_carry[1]), .CO(pe_1_2_3_sub_81_carry[2]), .S(
        pe_1_2_3_N71) );
  FA_X1 pe_1_2_3_add_83_U1_7 ( .A(int_data_res_2__3__7_), .B(
        pe_1_2_3_int_data_3_), .CI(pe_1_2_3_add_83_carry[7]), .S(pe_1_2_3_N85)
         );
  FA_X1 pe_1_2_3_add_83_U1_6 ( .A(int_data_res_2__3__6_), .B(
        pe_1_2_3_int_data_3_), .CI(pe_1_2_3_add_83_carry[6]), .CO(
        pe_1_2_3_add_83_carry[7]), .S(pe_1_2_3_N84) );
  FA_X1 pe_1_2_3_add_83_U1_5 ( .A(int_data_res_2__3__5_), .B(
        pe_1_2_3_int_data_3_), .CI(pe_1_2_3_add_83_carry[5]), .CO(
        pe_1_2_3_add_83_carry[6]), .S(pe_1_2_3_N83) );
  FA_X1 pe_1_2_3_add_83_U1_4 ( .A(int_data_res_2__3__4_), .B(
        pe_1_2_3_int_data_3_), .CI(pe_1_2_3_add_83_carry[4]), .CO(
        pe_1_2_3_add_83_carry[5]), .S(pe_1_2_3_N82) );
  FA_X1 pe_1_2_3_add_83_U1_3 ( .A(int_data_res_2__3__3_), .B(
        pe_1_2_3_int_data_3_), .CI(pe_1_2_3_add_83_carry[3]), .CO(
        pe_1_2_3_add_83_carry[4]), .S(pe_1_2_3_N81) );
  FA_X1 pe_1_2_3_add_83_U1_2 ( .A(int_data_res_2__3__2_), .B(
        pe_1_2_3_int_data_2_), .CI(pe_1_2_3_add_83_carry[2]), .CO(
        pe_1_2_3_add_83_carry[3]), .S(pe_1_2_3_N80) );
  FA_X1 pe_1_2_3_add_83_U1_1 ( .A(int_data_res_2__3__1_), .B(
        pe_1_2_3_int_data_1_), .CI(pe_1_2_3_n2), .CO(pe_1_2_3_add_83_carry[2]), 
        .S(pe_1_2_3_N79) );
  NAND3_X1 pe_1_2_3_U56 ( .A1(pe_1_2_3_n60), .A2(pe_1_2_3_n43), .A3(
        pe_1_2_3_n62), .ZN(pe_1_2_3_n40) );
  NAND3_X1 pe_1_2_3_U55 ( .A1(pe_1_2_3_n43), .A2(pe_1_2_3_n61), .A3(
        pe_1_2_3_n62), .ZN(pe_1_2_3_n39) );
  NAND3_X1 pe_1_2_3_U54 ( .A1(pe_1_2_3_n43), .A2(pe_1_2_3_n63), .A3(
        pe_1_2_3_n60), .ZN(pe_1_2_3_n38) );
  NAND3_X1 pe_1_2_3_U53 ( .A1(pe_1_2_3_n61), .A2(pe_1_2_3_n63), .A3(
        pe_1_2_3_n43), .ZN(pe_1_2_3_n37) );
  DFFR_X1 pe_1_2_3_int_q_acc_reg_6_ ( .D(pe_1_2_3_n78), .CK(pe_1_2_3_net6070), 
        .RN(pe_1_2_3_n71), .Q(int_data_res_2__3__6_) );
  DFFR_X1 pe_1_2_3_int_q_acc_reg_5_ ( .D(pe_1_2_3_n79), .CK(pe_1_2_3_net6070), 
        .RN(pe_1_2_3_n71), .Q(int_data_res_2__3__5_) );
  DFFR_X1 pe_1_2_3_int_q_acc_reg_4_ ( .D(pe_1_2_3_n80), .CK(pe_1_2_3_net6070), 
        .RN(pe_1_2_3_n71), .Q(int_data_res_2__3__4_) );
  DFFR_X1 pe_1_2_3_int_q_acc_reg_3_ ( .D(pe_1_2_3_n81), .CK(pe_1_2_3_net6070), 
        .RN(pe_1_2_3_n71), .Q(int_data_res_2__3__3_) );
  DFFR_X1 pe_1_2_3_int_q_acc_reg_2_ ( .D(pe_1_2_3_n82), .CK(pe_1_2_3_net6070), 
        .RN(pe_1_2_3_n71), .Q(int_data_res_2__3__2_) );
  DFFR_X1 pe_1_2_3_int_q_acc_reg_1_ ( .D(pe_1_2_3_n83), .CK(pe_1_2_3_net6070), 
        .RN(pe_1_2_3_n71), .Q(int_data_res_2__3__1_) );
  DFFR_X1 pe_1_2_3_int_q_acc_reg_7_ ( .D(pe_1_2_3_n77), .CK(pe_1_2_3_net6070), 
        .RN(pe_1_2_3_n71), .Q(int_data_res_2__3__7_) );
  CLKGATETST_X1 pe_1_2_3_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_2_3_n88), .SE(1'b0), .GCK(pe_1_2_3_net6009) );
  CLKGATETST_X1 pe_1_2_3_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_2_3_n87), .SE(1'b0), .GCK(pe_1_2_3_net6015) );
  CLKGATETST_X1 pe_1_2_3_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_2_3_n86), .SE(1'b0), .GCK(pe_1_2_3_net6020) );
  CLKGATETST_X1 pe_1_2_3_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_2_3_n85), .SE(1'b0), .GCK(pe_1_2_3_net6025) );
  CLKGATETST_X1 pe_1_2_3_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_2_3_n90), .SE(1'b0), .GCK(pe_1_2_3_net6030) );
  CLKGATETST_X1 pe_1_2_3_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_2_3_n89), .SE(1'b0), .GCK(pe_1_2_3_net6035) );
  CLKGATETST_X1 pe_1_2_3_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_2_3_N64), .SE(1'b0), .GCK(pe_1_2_3_net6040) );
  CLKGATETST_X1 pe_1_2_3_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_2_3_N63), .SE(1'b0), .GCK(pe_1_2_3_net6045) );
  CLKGATETST_X1 pe_1_2_3_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_2_3_N62), .SE(1'b0), .GCK(pe_1_2_3_net6050) );
  CLKGATETST_X1 pe_1_2_3_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_2_3_N61), .SE(1'b0), .GCK(pe_1_2_3_net6055) );
  CLKGATETST_X1 pe_1_2_3_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_2_3_N60), .SE(1'b0), .GCK(pe_1_2_3_net6060) );
  CLKGATETST_X1 pe_1_2_3_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_2_3_N59), .SE(1'b0), .GCK(pe_1_2_3_net6065) );
  CLKGATETST_X1 pe_1_2_3_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_2_3_N90), .SE(1'b0), .GCK(pe_1_2_3_net6070) );
  CLKBUF_X1 pe_1_2_4_U112 ( .A(pe_1_2_4_n72), .Z(pe_1_2_4_n71) );
  INV_X1 pe_1_2_4_U111 ( .A(n74), .ZN(pe_1_2_4_n70) );
  INV_X1 pe_1_2_4_U110 ( .A(n66), .ZN(pe_1_2_4_n69) );
  INV_X1 pe_1_2_4_U109 ( .A(n66), .ZN(pe_1_2_4_n68) );
  INV_X1 pe_1_2_4_U108 ( .A(n66), .ZN(pe_1_2_4_n67) );
  INV_X1 pe_1_2_4_U107 ( .A(pe_1_2_4_n69), .ZN(pe_1_2_4_n66) );
  INV_X1 pe_1_2_4_U106 ( .A(pe_1_2_4_n63), .ZN(pe_1_2_4_n62) );
  INV_X1 pe_1_2_4_U105 ( .A(pe_1_2_4_n61), .ZN(pe_1_2_4_n60) );
  INV_X1 pe_1_2_4_U104 ( .A(n26), .ZN(pe_1_2_4_n59) );
  INV_X1 pe_1_2_4_U103 ( .A(pe_1_2_4_n59), .ZN(pe_1_2_4_n58) );
  INV_X1 pe_1_2_4_U102 ( .A(n18), .ZN(pe_1_2_4_n57) );
  MUX2_X1 pe_1_2_4_U101 ( .A(pe_1_2_4_n54), .B(pe_1_2_4_n51), .S(n47), .Z(
        int_data_x_2__4__3_) );
  MUX2_X1 pe_1_2_4_U100 ( .A(pe_1_2_4_n53), .B(pe_1_2_4_n52), .S(pe_1_2_4_n62), 
        .Z(pe_1_2_4_n54) );
  MUX2_X1 pe_1_2_4_U99 ( .A(pe_1_2_4_int_q_reg_h[23]), .B(
        pe_1_2_4_int_q_reg_h[19]), .S(pe_1_2_4_n56), .Z(pe_1_2_4_n53) );
  MUX2_X1 pe_1_2_4_U98 ( .A(pe_1_2_4_int_q_reg_h[15]), .B(
        pe_1_2_4_int_q_reg_h[11]), .S(pe_1_2_4_n56), .Z(pe_1_2_4_n52) );
  MUX2_X1 pe_1_2_4_U97 ( .A(pe_1_2_4_int_q_reg_h[7]), .B(
        pe_1_2_4_int_q_reg_h[3]), .S(pe_1_2_4_n56), .Z(pe_1_2_4_n51) );
  MUX2_X1 pe_1_2_4_U96 ( .A(pe_1_2_4_n50), .B(pe_1_2_4_n47), .S(n47), .Z(
        int_data_x_2__4__2_) );
  MUX2_X1 pe_1_2_4_U95 ( .A(pe_1_2_4_n49), .B(pe_1_2_4_n48), .S(pe_1_2_4_n62), 
        .Z(pe_1_2_4_n50) );
  MUX2_X1 pe_1_2_4_U94 ( .A(pe_1_2_4_int_q_reg_h[22]), .B(
        pe_1_2_4_int_q_reg_h[18]), .S(pe_1_2_4_n56), .Z(pe_1_2_4_n49) );
  MUX2_X1 pe_1_2_4_U93 ( .A(pe_1_2_4_int_q_reg_h[14]), .B(
        pe_1_2_4_int_q_reg_h[10]), .S(pe_1_2_4_n56), .Z(pe_1_2_4_n48) );
  MUX2_X1 pe_1_2_4_U92 ( .A(pe_1_2_4_int_q_reg_h[6]), .B(
        pe_1_2_4_int_q_reg_h[2]), .S(pe_1_2_4_n56), .Z(pe_1_2_4_n47) );
  MUX2_X1 pe_1_2_4_U91 ( .A(pe_1_2_4_n46), .B(pe_1_2_4_n24), .S(n47), .Z(
        int_data_x_2__4__1_) );
  MUX2_X1 pe_1_2_4_U90 ( .A(pe_1_2_4_n45), .B(pe_1_2_4_n25), .S(pe_1_2_4_n62), 
        .Z(pe_1_2_4_n46) );
  MUX2_X1 pe_1_2_4_U89 ( .A(pe_1_2_4_int_q_reg_h[21]), .B(
        pe_1_2_4_int_q_reg_h[17]), .S(pe_1_2_4_n56), .Z(pe_1_2_4_n45) );
  MUX2_X1 pe_1_2_4_U88 ( .A(pe_1_2_4_int_q_reg_h[13]), .B(
        pe_1_2_4_int_q_reg_h[9]), .S(pe_1_2_4_n56), .Z(pe_1_2_4_n25) );
  MUX2_X1 pe_1_2_4_U87 ( .A(pe_1_2_4_int_q_reg_h[5]), .B(
        pe_1_2_4_int_q_reg_h[1]), .S(pe_1_2_4_n56), .Z(pe_1_2_4_n24) );
  MUX2_X1 pe_1_2_4_U86 ( .A(pe_1_2_4_n23), .B(pe_1_2_4_n20), .S(n47), .Z(
        int_data_x_2__4__0_) );
  MUX2_X1 pe_1_2_4_U85 ( .A(pe_1_2_4_n22), .B(pe_1_2_4_n21), .S(pe_1_2_4_n62), 
        .Z(pe_1_2_4_n23) );
  MUX2_X1 pe_1_2_4_U84 ( .A(pe_1_2_4_int_q_reg_h[20]), .B(
        pe_1_2_4_int_q_reg_h[16]), .S(pe_1_2_4_n56), .Z(pe_1_2_4_n22) );
  MUX2_X1 pe_1_2_4_U83 ( .A(pe_1_2_4_int_q_reg_h[12]), .B(
        pe_1_2_4_int_q_reg_h[8]), .S(pe_1_2_4_n56), .Z(pe_1_2_4_n21) );
  MUX2_X1 pe_1_2_4_U82 ( .A(pe_1_2_4_int_q_reg_h[4]), .B(
        pe_1_2_4_int_q_reg_h[0]), .S(pe_1_2_4_n56), .Z(pe_1_2_4_n20) );
  MUX2_X1 pe_1_2_4_U81 ( .A(pe_1_2_4_n19), .B(pe_1_2_4_n16), .S(n47), .Z(
        int_data_y_2__4__3_) );
  MUX2_X1 pe_1_2_4_U80 ( .A(pe_1_2_4_n18), .B(pe_1_2_4_n17), .S(pe_1_2_4_n62), 
        .Z(pe_1_2_4_n19) );
  MUX2_X1 pe_1_2_4_U79 ( .A(pe_1_2_4_int_q_reg_v[23]), .B(
        pe_1_2_4_int_q_reg_v[19]), .S(pe_1_2_4_n55), .Z(pe_1_2_4_n18) );
  MUX2_X1 pe_1_2_4_U78 ( .A(pe_1_2_4_int_q_reg_v[15]), .B(
        pe_1_2_4_int_q_reg_v[11]), .S(pe_1_2_4_n55), .Z(pe_1_2_4_n17) );
  MUX2_X1 pe_1_2_4_U77 ( .A(pe_1_2_4_int_q_reg_v[7]), .B(
        pe_1_2_4_int_q_reg_v[3]), .S(pe_1_2_4_n55), .Z(pe_1_2_4_n16) );
  MUX2_X1 pe_1_2_4_U76 ( .A(pe_1_2_4_n15), .B(pe_1_2_4_n12), .S(n47), .Z(
        int_data_y_2__4__2_) );
  MUX2_X1 pe_1_2_4_U75 ( .A(pe_1_2_4_n14), .B(pe_1_2_4_n13), .S(pe_1_2_4_n62), 
        .Z(pe_1_2_4_n15) );
  MUX2_X1 pe_1_2_4_U74 ( .A(pe_1_2_4_int_q_reg_v[22]), .B(
        pe_1_2_4_int_q_reg_v[18]), .S(pe_1_2_4_n55), .Z(pe_1_2_4_n14) );
  MUX2_X1 pe_1_2_4_U73 ( .A(pe_1_2_4_int_q_reg_v[14]), .B(
        pe_1_2_4_int_q_reg_v[10]), .S(pe_1_2_4_n55), .Z(pe_1_2_4_n13) );
  MUX2_X1 pe_1_2_4_U72 ( .A(pe_1_2_4_int_q_reg_v[6]), .B(
        pe_1_2_4_int_q_reg_v[2]), .S(pe_1_2_4_n55), .Z(pe_1_2_4_n12) );
  MUX2_X1 pe_1_2_4_U71 ( .A(pe_1_2_4_n11), .B(pe_1_2_4_n8), .S(n47), .Z(
        int_data_y_2__4__1_) );
  MUX2_X1 pe_1_2_4_U70 ( .A(pe_1_2_4_n10), .B(pe_1_2_4_n9), .S(pe_1_2_4_n62), 
        .Z(pe_1_2_4_n11) );
  MUX2_X1 pe_1_2_4_U69 ( .A(pe_1_2_4_int_q_reg_v[21]), .B(
        pe_1_2_4_int_q_reg_v[17]), .S(pe_1_2_4_n55), .Z(pe_1_2_4_n10) );
  MUX2_X1 pe_1_2_4_U68 ( .A(pe_1_2_4_int_q_reg_v[13]), .B(
        pe_1_2_4_int_q_reg_v[9]), .S(pe_1_2_4_n55), .Z(pe_1_2_4_n9) );
  MUX2_X1 pe_1_2_4_U67 ( .A(pe_1_2_4_int_q_reg_v[5]), .B(
        pe_1_2_4_int_q_reg_v[1]), .S(pe_1_2_4_n55), .Z(pe_1_2_4_n8) );
  MUX2_X1 pe_1_2_4_U66 ( .A(pe_1_2_4_n7), .B(pe_1_2_4_n4), .S(n47), .Z(
        int_data_y_2__4__0_) );
  MUX2_X1 pe_1_2_4_U65 ( .A(pe_1_2_4_n6), .B(pe_1_2_4_n5), .S(pe_1_2_4_n62), 
        .Z(pe_1_2_4_n7) );
  MUX2_X1 pe_1_2_4_U64 ( .A(pe_1_2_4_int_q_reg_v[20]), .B(
        pe_1_2_4_int_q_reg_v[16]), .S(pe_1_2_4_n55), .Z(pe_1_2_4_n6) );
  MUX2_X1 pe_1_2_4_U63 ( .A(pe_1_2_4_int_q_reg_v[12]), .B(
        pe_1_2_4_int_q_reg_v[8]), .S(pe_1_2_4_n55), .Z(pe_1_2_4_n5) );
  MUX2_X1 pe_1_2_4_U62 ( .A(pe_1_2_4_int_q_reg_v[4]), .B(
        pe_1_2_4_int_q_reg_v[0]), .S(pe_1_2_4_n55), .Z(pe_1_2_4_n4) );
  AOI222_X1 pe_1_2_4_U61 ( .A1(int_data_res_3__4__2_), .A2(pe_1_2_4_n64), .B1(
        pe_1_2_4_N80), .B2(pe_1_2_4_n27), .C1(pe_1_2_4_N72), .C2(pe_1_2_4_n28), 
        .ZN(pe_1_2_4_n33) );
  INV_X1 pe_1_2_4_U60 ( .A(pe_1_2_4_n33), .ZN(pe_1_2_4_n82) );
  AOI222_X1 pe_1_2_4_U59 ( .A1(int_data_res_3__4__6_), .A2(pe_1_2_4_n64), .B1(
        pe_1_2_4_N84), .B2(pe_1_2_4_n27), .C1(pe_1_2_4_N76), .C2(pe_1_2_4_n28), 
        .ZN(pe_1_2_4_n29) );
  INV_X1 pe_1_2_4_U58 ( .A(pe_1_2_4_n29), .ZN(pe_1_2_4_n78) );
  XNOR2_X1 pe_1_2_4_U57 ( .A(pe_1_2_4_n73), .B(int_data_res_2__4__0_), .ZN(
        pe_1_2_4_N70) );
  AOI222_X1 pe_1_2_4_U52 ( .A1(int_data_res_3__4__0_), .A2(pe_1_2_4_n64), .B1(
        pe_1_2_4_n1), .B2(pe_1_2_4_n27), .C1(pe_1_2_4_N70), .C2(pe_1_2_4_n28), 
        .ZN(pe_1_2_4_n35) );
  INV_X1 pe_1_2_4_U51 ( .A(pe_1_2_4_n35), .ZN(pe_1_2_4_n84) );
  AOI222_X1 pe_1_2_4_U50 ( .A1(int_data_res_3__4__1_), .A2(pe_1_2_4_n64), .B1(
        pe_1_2_4_N79), .B2(pe_1_2_4_n27), .C1(pe_1_2_4_N71), .C2(pe_1_2_4_n28), 
        .ZN(pe_1_2_4_n34) );
  INV_X1 pe_1_2_4_U49 ( .A(pe_1_2_4_n34), .ZN(pe_1_2_4_n83) );
  AOI222_X1 pe_1_2_4_U48 ( .A1(int_data_res_3__4__3_), .A2(pe_1_2_4_n64), .B1(
        pe_1_2_4_N81), .B2(pe_1_2_4_n27), .C1(pe_1_2_4_N73), .C2(pe_1_2_4_n28), 
        .ZN(pe_1_2_4_n32) );
  INV_X1 pe_1_2_4_U47 ( .A(pe_1_2_4_n32), .ZN(pe_1_2_4_n81) );
  AOI222_X1 pe_1_2_4_U46 ( .A1(int_data_res_3__4__4_), .A2(pe_1_2_4_n64), .B1(
        pe_1_2_4_N82), .B2(pe_1_2_4_n27), .C1(pe_1_2_4_N74), .C2(pe_1_2_4_n28), 
        .ZN(pe_1_2_4_n31) );
  INV_X1 pe_1_2_4_U45 ( .A(pe_1_2_4_n31), .ZN(pe_1_2_4_n80) );
  AOI222_X1 pe_1_2_4_U44 ( .A1(int_data_res_3__4__5_), .A2(pe_1_2_4_n64), .B1(
        pe_1_2_4_N83), .B2(pe_1_2_4_n27), .C1(pe_1_2_4_N75), .C2(pe_1_2_4_n28), 
        .ZN(pe_1_2_4_n30) );
  INV_X1 pe_1_2_4_U43 ( .A(pe_1_2_4_n30), .ZN(pe_1_2_4_n79) );
  NAND2_X1 pe_1_2_4_U42 ( .A1(pe_1_2_4_int_data_0_), .A2(pe_1_2_4_n3), .ZN(
        pe_1_2_4_sub_81_carry[1]) );
  INV_X1 pe_1_2_4_U41 ( .A(pe_1_2_4_int_data_1_), .ZN(pe_1_2_4_n74) );
  INV_X1 pe_1_2_4_U40 ( .A(pe_1_2_4_int_data_2_), .ZN(pe_1_2_4_n75) );
  AND2_X1 pe_1_2_4_U39 ( .A1(pe_1_2_4_int_data_0_), .A2(int_data_res_2__4__0_), 
        .ZN(pe_1_2_4_n2) );
  AOI222_X1 pe_1_2_4_U38 ( .A1(pe_1_2_4_n64), .A2(int_data_res_3__4__7_), .B1(
        pe_1_2_4_N85), .B2(pe_1_2_4_n27), .C1(pe_1_2_4_N77), .C2(pe_1_2_4_n28), 
        .ZN(pe_1_2_4_n26) );
  INV_X1 pe_1_2_4_U37 ( .A(pe_1_2_4_n26), .ZN(pe_1_2_4_n77) );
  NOR3_X1 pe_1_2_4_U36 ( .A1(pe_1_2_4_n59), .A2(pe_1_2_4_n65), .A3(int_ckg[43]), .ZN(pe_1_2_4_n36) );
  OR2_X1 pe_1_2_4_U35 ( .A1(pe_1_2_4_n36), .A2(pe_1_2_4_n64), .ZN(pe_1_2_4_N90) );
  INV_X1 pe_1_2_4_U34 ( .A(n38), .ZN(pe_1_2_4_n63) );
  AND2_X1 pe_1_2_4_U33 ( .A1(int_data_x_2__4__2_), .A2(pe_1_2_4_n58), .ZN(
        pe_1_2_4_int_data_2_) );
  AND2_X1 pe_1_2_4_U32 ( .A1(int_data_x_2__4__1_), .A2(pe_1_2_4_n58), .ZN(
        pe_1_2_4_int_data_1_) );
  AND2_X1 pe_1_2_4_U31 ( .A1(int_data_x_2__4__3_), .A2(pe_1_2_4_n58), .ZN(
        pe_1_2_4_int_data_3_) );
  BUF_X1 pe_1_2_4_U30 ( .A(n60), .Z(pe_1_2_4_n64) );
  INV_X1 pe_1_2_4_U29 ( .A(n32), .ZN(pe_1_2_4_n61) );
  AND2_X1 pe_1_2_4_U28 ( .A1(int_data_x_2__4__0_), .A2(pe_1_2_4_n58), .ZN(
        pe_1_2_4_int_data_0_) );
  NAND2_X1 pe_1_2_4_U27 ( .A1(pe_1_2_4_n44), .A2(pe_1_2_4_n61), .ZN(
        pe_1_2_4_n41) );
  AND3_X1 pe_1_2_4_U26 ( .A1(n74), .A2(pe_1_2_4_n63), .A3(n47), .ZN(
        pe_1_2_4_n44) );
  INV_X1 pe_1_2_4_U25 ( .A(pe_1_2_4_int_data_3_), .ZN(pe_1_2_4_n76) );
  NOR2_X1 pe_1_2_4_U24 ( .A1(pe_1_2_4_n70), .A2(n47), .ZN(pe_1_2_4_n43) );
  NOR2_X1 pe_1_2_4_U23 ( .A1(pe_1_2_4_n57), .A2(pe_1_2_4_n64), .ZN(
        pe_1_2_4_n28) );
  NOR2_X1 pe_1_2_4_U22 ( .A1(n18), .A2(pe_1_2_4_n64), .ZN(pe_1_2_4_n27) );
  INV_X1 pe_1_2_4_U21 ( .A(pe_1_2_4_int_data_0_), .ZN(pe_1_2_4_n73) );
  INV_X1 pe_1_2_4_U20 ( .A(pe_1_2_4_n41), .ZN(pe_1_2_4_n90) );
  INV_X1 pe_1_2_4_U19 ( .A(pe_1_2_4_n37), .ZN(pe_1_2_4_n88) );
  INV_X1 pe_1_2_4_U18 ( .A(pe_1_2_4_n38), .ZN(pe_1_2_4_n87) );
  INV_X1 pe_1_2_4_U17 ( .A(pe_1_2_4_n39), .ZN(pe_1_2_4_n86) );
  NOR2_X1 pe_1_2_4_U16 ( .A1(pe_1_2_4_n68), .A2(pe_1_2_4_n42), .ZN(
        pe_1_2_4_N59) );
  NOR2_X1 pe_1_2_4_U15 ( .A1(pe_1_2_4_n68), .A2(pe_1_2_4_n41), .ZN(
        pe_1_2_4_N60) );
  NOR2_X1 pe_1_2_4_U14 ( .A1(pe_1_2_4_n68), .A2(pe_1_2_4_n38), .ZN(
        pe_1_2_4_N63) );
  NOR2_X1 pe_1_2_4_U13 ( .A1(pe_1_2_4_n67), .A2(pe_1_2_4_n40), .ZN(
        pe_1_2_4_N61) );
  NOR2_X1 pe_1_2_4_U12 ( .A1(pe_1_2_4_n67), .A2(pe_1_2_4_n39), .ZN(
        pe_1_2_4_N62) );
  NOR2_X1 pe_1_2_4_U11 ( .A1(pe_1_2_4_n37), .A2(pe_1_2_4_n67), .ZN(
        pe_1_2_4_N64) );
  NAND2_X1 pe_1_2_4_U10 ( .A1(pe_1_2_4_n44), .A2(pe_1_2_4_n60), .ZN(
        pe_1_2_4_n42) );
  BUF_X1 pe_1_2_4_U9 ( .A(pe_1_2_4_n60), .Z(pe_1_2_4_n55) );
  INV_X1 pe_1_2_4_U8 ( .A(pe_1_2_4_n69), .ZN(pe_1_2_4_n65) );
  BUF_X1 pe_1_2_4_U7 ( .A(pe_1_2_4_n60), .Z(pe_1_2_4_n56) );
  INV_X1 pe_1_2_4_U6 ( .A(pe_1_2_4_n42), .ZN(pe_1_2_4_n89) );
  INV_X1 pe_1_2_4_U5 ( .A(pe_1_2_4_n40), .ZN(pe_1_2_4_n85) );
  INV_X2 pe_1_2_4_U4 ( .A(n82), .ZN(pe_1_2_4_n72) );
  XOR2_X1 pe_1_2_4_U3 ( .A(pe_1_2_4_int_data_0_), .B(int_data_res_2__4__0_), 
        .Z(pe_1_2_4_n1) );
  DFFR_X1 pe_1_2_4_int_q_acc_reg_0_ ( .D(pe_1_2_4_n84), .CK(pe_1_2_4_net5992), 
        .RN(pe_1_2_4_n72), .Q(int_data_res_2__4__0_), .QN(pe_1_2_4_n3) );
  DFFR_X1 pe_1_2_4_int_q_reg_v_reg_0__0_ ( .D(int_data_y_3__4__0_), .CK(
        pe_1_2_4_net5962), .RN(pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_v[20]) );
  DFFR_X1 pe_1_2_4_int_q_reg_v_reg_0__1_ ( .D(int_data_y_3__4__1_), .CK(
        pe_1_2_4_net5962), .RN(pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_v[21]) );
  DFFR_X1 pe_1_2_4_int_q_reg_v_reg_0__2_ ( .D(int_data_y_3__4__2_), .CK(
        pe_1_2_4_net5962), .RN(pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_v[22]) );
  DFFR_X1 pe_1_2_4_int_q_reg_v_reg_0__3_ ( .D(int_data_y_3__4__3_), .CK(
        pe_1_2_4_net5962), .RN(pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_v[23]) );
  DFFR_X1 pe_1_2_4_int_q_reg_v_reg_1__0_ ( .D(int_data_y_3__4__0_), .CK(
        pe_1_2_4_net5967), .RN(pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_v[16]) );
  DFFR_X1 pe_1_2_4_int_q_reg_v_reg_1__1_ ( .D(int_data_y_3__4__1_), .CK(
        pe_1_2_4_net5967), .RN(pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_v[17]) );
  DFFR_X1 pe_1_2_4_int_q_reg_v_reg_1__2_ ( .D(int_data_y_3__4__2_), .CK(
        pe_1_2_4_net5967), .RN(pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_v[18]) );
  DFFR_X1 pe_1_2_4_int_q_reg_v_reg_1__3_ ( .D(int_data_y_3__4__3_), .CK(
        pe_1_2_4_net5967), .RN(pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_v[19]) );
  DFFR_X1 pe_1_2_4_int_q_reg_v_reg_2__0_ ( .D(int_data_y_3__4__0_), .CK(
        pe_1_2_4_net5972), .RN(pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_v[12]) );
  DFFR_X1 pe_1_2_4_int_q_reg_v_reg_2__1_ ( .D(int_data_y_3__4__1_), .CK(
        pe_1_2_4_net5972), .RN(pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_v[13]) );
  DFFR_X1 pe_1_2_4_int_q_reg_v_reg_2__2_ ( .D(int_data_y_3__4__2_), .CK(
        pe_1_2_4_net5972), .RN(pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_v[14]) );
  DFFR_X1 pe_1_2_4_int_q_reg_v_reg_2__3_ ( .D(int_data_y_3__4__3_), .CK(
        pe_1_2_4_net5972), .RN(pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_v[15]) );
  DFFR_X1 pe_1_2_4_int_q_reg_v_reg_3__0_ ( .D(int_data_y_3__4__0_), .CK(
        pe_1_2_4_net5977), .RN(pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_v[8]) );
  DFFR_X1 pe_1_2_4_int_q_reg_v_reg_3__1_ ( .D(int_data_y_3__4__1_), .CK(
        pe_1_2_4_net5977), .RN(pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_v[9]) );
  DFFR_X1 pe_1_2_4_int_q_reg_v_reg_3__2_ ( .D(int_data_y_3__4__2_), .CK(
        pe_1_2_4_net5977), .RN(pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_v[10]) );
  DFFR_X1 pe_1_2_4_int_q_reg_v_reg_3__3_ ( .D(int_data_y_3__4__3_), .CK(
        pe_1_2_4_net5977), .RN(pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_v[11]) );
  DFFR_X1 pe_1_2_4_int_q_reg_v_reg_4__0_ ( .D(int_data_y_3__4__0_), .CK(
        pe_1_2_4_net5982), .RN(pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_v[4]) );
  DFFR_X1 pe_1_2_4_int_q_reg_v_reg_4__1_ ( .D(int_data_y_3__4__1_), .CK(
        pe_1_2_4_net5982), .RN(pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_v[5]) );
  DFFR_X1 pe_1_2_4_int_q_reg_v_reg_4__2_ ( .D(int_data_y_3__4__2_), .CK(
        pe_1_2_4_net5982), .RN(pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_v[6]) );
  DFFR_X1 pe_1_2_4_int_q_reg_v_reg_4__3_ ( .D(int_data_y_3__4__3_), .CK(
        pe_1_2_4_net5982), .RN(pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_v[7]) );
  DFFR_X1 pe_1_2_4_int_q_reg_v_reg_5__0_ ( .D(int_data_y_3__4__0_), .CK(
        pe_1_2_4_net5987), .RN(pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_v[0]) );
  DFFR_X1 pe_1_2_4_int_q_reg_v_reg_5__1_ ( .D(int_data_y_3__4__1_), .CK(
        pe_1_2_4_net5987), .RN(pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_v[1]) );
  DFFR_X1 pe_1_2_4_int_q_reg_v_reg_5__2_ ( .D(int_data_y_3__4__2_), .CK(
        pe_1_2_4_net5987), .RN(pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_v[2]) );
  DFFR_X1 pe_1_2_4_int_q_reg_v_reg_5__3_ ( .D(int_data_y_3__4__3_), .CK(
        pe_1_2_4_net5987), .RN(pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_2_4_int_q_reg_h_reg_0__0_ ( .D(int_data_x_2__5__0_), .SI(
        int_data_y_3__4__0_), .SE(pe_1_2_4_n65), .CK(pe_1_2_4_net5931), .RN(
        pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_2_4_int_q_reg_h_reg_0__1_ ( .D(int_data_x_2__5__1_), .SI(
        int_data_y_3__4__1_), .SE(pe_1_2_4_n65), .CK(pe_1_2_4_net5931), .RN(
        pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_2_4_int_q_reg_h_reg_0__2_ ( .D(int_data_x_2__5__2_), .SI(
        int_data_y_3__4__2_), .SE(pe_1_2_4_n65), .CK(pe_1_2_4_net5931), .RN(
        pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_2_4_int_q_reg_h_reg_0__3_ ( .D(int_data_x_2__5__3_), .SI(
        int_data_y_3__4__3_), .SE(pe_1_2_4_n65), .CK(pe_1_2_4_net5931), .RN(
        pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_2_4_int_q_reg_h_reg_1__0_ ( .D(int_data_x_2__5__0_), .SI(
        int_data_y_3__4__0_), .SE(pe_1_2_4_n65), .CK(pe_1_2_4_net5937), .RN(
        pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_2_4_int_q_reg_h_reg_1__1_ ( .D(int_data_x_2__5__1_), .SI(
        int_data_y_3__4__1_), .SE(pe_1_2_4_n65), .CK(pe_1_2_4_net5937), .RN(
        pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_2_4_int_q_reg_h_reg_1__2_ ( .D(int_data_x_2__5__2_), .SI(
        int_data_y_3__4__2_), .SE(pe_1_2_4_n65), .CK(pe_1_2_4_net5937), .RN(
        pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_2_4_int_q_reg_h_reg_1__3_ ( .D(int_data_x_2__5__3_), .SI(
        int_data_y_3__4__3_), .SE(pe_1_2_4_n65), .CK(pe_1_2_4_net5937), .RN(
        pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_2_4_int_q_reg_h_reg_2__0_ ( .D(int_data_x_2__5__0_), .SI(
        int_data_y_3__4__0_), .SE(pe_1_2_4_n65), .CK(pe_1_2_4_net5942), .RN(
        pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_2_4_int_q_reg_h_reg_2__1_ ( .D(int_data_x_2__5__1_), .SI(
        int_data_y_3__4__1_), .SE(pe_1_2_4_n65), .CK(pe_1_2_4_net5942), .RN(
        pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_2_4_int_q_reg_h_reg_2__2_ ( .D(int_data_x_2__5__2_), .SI(
        int_data_y_3__4__2_), .SE(pe_1_2_4_n65), .CK(pe_1_2_4_net5942), .RN(
        pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_2_4_int_q_reg_h_reg_2__3_ ( .D(int_data_x_2__5__3_), .SI(
        int_data_y_3__4__3_), .SE(pe_1_2_4_n65), .CK(pe_1_2_4_net5942), .RN(
        pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_2_4_int_q_reg_h_reg_3__0_ ( .D(int_data_x_2__5__0_), .SI(
        int_data_y_3__4__0_), .SE(pe_1_2_4_n65), .CK(pe_1_2_4_net5947), .RN(
        pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_2_4_int_q_reg_h_reg_3__1_ ( .D(int_data_x_2__5__1_), .SI(
        int_data_y_3__4__1_), .SE(pe_1_2_4_n65), .CK(pe_1_2_4_net5947), .RN(
        pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_2_4_int_q_reg_h_reg_3__2_ ( .D(int_data_x_2__5__2_), .SI(
        int_data_y_3__4__2_), .SE(pe_1_2_4_n65), .CK(pe_1_2_4_net5947), .RN(
        pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_2_4_int_q_reg_h_reg_3__3_ ( .D(int_data_x_2__5__3_), .SI(
        int_data_y_3__4__3_), .SE(pe_1_2_4_n65), .CK(pe_1_2_4_net5947), .RN(
        pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_2_4_int_q_reg_h_reg_4__0_ ( .D(int_data_x_2__5__0_), .SI(
        int_data_y_3__4__0_), .SE(pe_1_2_4_n66), .CK(pe_1_2_4_net5952), .RN(
        pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_2_4_int_q_reg_h_reg_4__1_ ( .D(int_data_x_2__5__1_), .SI(
        int_data_y_3__4__1_), .SE(pe_1_2_4_n66), .CK(pe_1_2_4_net5952), .RN(
        pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_2_4_int_q_reg_h_reg_4__2_ ( .D(int_data_x_2__5__2_), .SI(
        int_data_y_3__4__2_), .SE(pe_1_2_4_n66), .CK(pe_1_2_4_net5952), .RN(
        pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_2_4_int_q_reg_h_reg_4__3_ ( .D(int_data_x_2__5__3_), .SI(
        int_data_y_3__4__3_), .SE(pe_1_2_4_n66), .CK(pe_1_2_4_net5952), .RN(
        pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_2_4_int_q_reg_h_reg_5__0_ ( .D(int_data_x_2__5__0_), .SI(
        int_data_y_3__4__0_), .SE(pe_1_2_4_n66), .CK(pe_1_2_4_net5957), .RN(
        pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_2_4_int_q_reg_h_reg_5__1_ ( .D(int_data_x_2__5__1_), .SI(
        int_data_y_3__4__1_), .SE(pe_1_2_4_n66), .CK(pe_1_2_4_net5957), .RN(
        pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_2_4_int_q_reg_h_reg_5__2_ ( .D(int_data_x_2__5__2_), .SI(
        int_data_y_3__4__2_), .SE(pe_1_2_4_n66), .CK(pe_1_2_4_net5957), .RN(
        pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_2_4_int_q_reg_h_reg_5__3_ ( .D(int_data_x_2__5__3_), .SI(
        int_data_y_3__4__3_), .SE(pe_1_2_4_n66), .CK(pe_1_2_4_net5957), .RN(
        pe_1_2_4_n72), .Q(pe_1_2_4_int_q_reg_h[3]) );
  FA_X1 pe_1_2_4_sub_81_U2_7 ( .A(int_data_res_2__4__7_), .B(pe_1_2_4_n76), 
        .CI(pe_1_2_4_sub_81_carry[7]), .S(pe_1_2_4_N77) );
  FA_X1 pe_1_2_4_sub_81_U2_6 ( .A(int_data_res_2__4__6_), .B(pe_1_2_4_n76), 
        .CI(pe_1_2_4_sub_81_carry[6]), .CO(pe_1_2_4_sub_81_carry[7]), .S(
        pe_1_2_4_N76) );
  FA_X1 pe_1_2_4_sub_81_U2_5 ( .A(int_data_res_2__4__5_), .B(pe_1_2_4_n76), 
        .CI(pe_1_2_4_sub_81_carry[5]), .CO(pe_1_2_4_sub_81_carry[6]), .S(
        pe_1_2_4_N75) );
  FA_X1 pe_1_2_4_sub_81_U2_4 ( .A(int_data_res_2__4__4_), .B(pe_1_2_4_n76), 
        .CI(pe_1_2_4_sub_81_carry[4]), .CO(pe_1_2_4_sub_81_carry[5]), .S(
        pe_1_2_4_N74) );
  FA_X1 pe_1_2_4_sub_81_U2_3 ( .A(int_data_res_2__4__3_), .B(pe_1_2_4_n76), 
        .CI(pe_1_2_4_sub_81_carry[3]), .CO(pe_1_2_4_sub_81_carry[4]), .S(
        pe_1_2_4_N73) );
  FA_X1 pe_1_2_4_sub_81_U2_2 ( .A(int_data_res_2__4__2_), .B(pe_1_2_4_n75), 
        .CI(pe_1_2_4_sub_81_carry[2]), .CO(pe_1_2_4_sub_81_carry[3]), .S(
        pe_1_2_4_N72) );
  FA_X1 pe_1_2_4_sub_81_U2_1 ( .A(int_data_res_2__4__1_), .B(pe_1_2_4_n74), 
        .CI(pe_1_2_4_sub_81_carry[1]), .CO(pe_1_2_4_sub_81_carry[2]), .S(
        pe_1_2_4_N71) );
  FA_X1 pe_1_2_4_add_83_U1_7 ( .A(int_data_res_2__4__7_), .B(
        pe_1_2_4_int_data_3_), .CI(pe_1_2_4_add_83_carry[7]), .S(pe_1_2_4_N85)
         );
  FA_X1 pe_1_2_4_add_83_U1_6 ( .A(int_data_res_2__4__6_), .B(
        pe_1_2_4_int_data_3_), .CI(pe_1_2_4_add_83_carry[6]), .CO(
        pe_1_2_4_add_83_carry[7]), .S(pe_1_2_4_N84) );
  FA_X1 pe_1_2_4_add_83_U1_5 ( .A(int_data_res_2__4__5_), .B(
        pe_1_2_4_int_data_3_), .CI(pe_1_2_4_add_83_carry[5]), .CO(
        pe_1_2_4_add_83_carry[6]), .S(pe_1_2_4_N83) );
  FA_X1 pe_1_2_4_add_83_U1_4 ( .A(int_data_res_2__4__4_), .B(
        pe_1_2_4_int_data_3_), .CI(pe_1_2_4_add_83_carry[4]), .CO(
        pe_1_2_4_add_83_carry[5]), .S(pe_1_2_4_N82) );
  FA_X1 pe_1_2_4_add_83_U1_3 ( .A(int_data_res_2__4__3_), .B(
        pe_1_2_4_int_data_3_), .CI(pe_1_2_4_add_83_carry[3]), .CO(
        pe_1_2_4_add_83_carry[4]), .S(pe_1_2_4_N81) );
  FA_X1 pe_1_2_4_add_83_U1_2 ( .A(int_data_res_2__4__2_), .B(
        pe_1_2_4_int_data_2_), .CI(pe_1_2_4_add_83_carry[2]), .CO(
        pe_1_2_4_add_83_carry[3]), .S(pe_1_2_4_N80) );
  FA_X1 pe_1_2_4_add_83_U1_1 ( .A(int_data_res_2__4__1_), .B(
        pe_1_2_4_int_data_1_), .CI(pe_1_2_4_n2), .CO(pe_1_2_4_add_83_carry[2]), 
        .S(pe_1_2_4_N79) );
  NAND3_X1 pe_1_2_4_U56 ( .A1(pe_1_2_4_n60), .A2(pe_1_2_4_n43), .A3(
        pe_1_2_4_n62), .ZN(pe_1_2_4_n40) );
  NAND3_X1 pe_1_2_4_U55 ( .A1(pe_1_2_4_n43), .A2(pe_1_2_4_n61), .A3(
        pe_1_2_4_n62), .ZN(pe_1_2_4_n39) );
  NAND3_X1 pe_1_2_4_U54 ( .A1(pe_1_2_4_n43), .A2(pe_1_2_4_n63), .A3(
        pe_1_2_4_n60), .ZN(pe_1_2_4_n38) );
  NAND3_X1 pe_1_2_4_U53 ( .A1(pe_1_2_4_n61), .A2(pe_1_2_4_n63), .A3(
        pe_1_2_4_n43), .ZN(pe_1_2_4_n37) );
  DFFR_X1 pe_1_2_4_int_q_acc_reg_6_ ( .D(pe_1_2_4_n78), .CK(pe_1_2_4_net5992), 
        .RN(pe_1_2_4_n71), .Q(int_data_res_2__4__6_) );
  DFFR_X1 pe_1_2_4_int_q_acc_reg_5_ ( .D(pe_1_2_4_n79), .CK(pe_1_2_4_net5992), 
        .RN(pe_1_2_4_n71), .Q(int_data_res_2__4__5_) );
  DFFR_X1 pe_1_2_4_int_q_acc_reg_4_ ( .D(pe_1_2_4_n80), .CK(pe_1_2_4_net5992), 
        .RN(pe_1_2_4_n71), .Q(int_data_res_2__4__4_) );
  DFFR_X1 pe_1_2_4_int_q_acc_reg_3_ ( .D(pe_1_2_4_n81), .CK(pe_1_2_4_net5992), 
        .RN(pe_1_2_4_n71), .Q(int_data_res_2__4__3_) );
  DFFR_X1 pe_1_2_4_int_q_acc_reg_2_ ( .D(pe_1_2_4_n82), .CK(pe_1_2_4_net5992), 
        .RN(pe_1_2_4_n71), .Q(int_data_res_2__4__2_) );
  DFFR_X1 pe_1_2_4_int_q_acc_reg_1_ ( .D(pe_1_2_4_n83), .CK(pe_1_2_4_net5992), 
        .RN(pe_1_2_4_n71), .Q(int_data_res_2__4__1_) );
  DFFR_X1 pe_1_2_4_int_q_acc_reg_7_ ( .D(pe_1_2_4_n77), .CK(pe_1_2_4_net5992), 
        .RN(pe_1_2_4_n71), .Q(int_data_res_2__4__7_) );
  CLKGATETST_X1 pe_1_2_4_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_2_4_n88), .SE(1'b0), .GCK(pe_1_2_4_net5931) );
  CLKGATETST_X1 pe_1_2_4_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_2_4_n87), .SE(1'b0), .GCK(pe_1_2_4_net5937) );
  CLKGATETST_X1 pe_1_2_4_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_2_4_n86), .SE(1'b0), .GCK(pe_1_2_4_net5942) );
  CLKGATETST_X1 pe_1_2_4_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_2_4_n85), .SE(1'b0), .GCK(pe_1_2_4_net5947) );
  CLKGATETST_X1 pe_1_2_4_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_2_4_n90), .SE(1'b0), .GCK(pe_1_2_4_net5952) );
  CLKGATETST_X1 pe_1_2_4_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_2_4_n89), .SE(1'b0), .GCK(pe_1_2_4_net5957) );
  CLKGATETST_X1 pe_1_2_4_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_2_4_N64), .SE(1'b0), .GCK(pe_1_2_4_net5962) );
  CLKGATETST_X1 pe_1_2_4_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_2_4_N63), .SE(1'b0), .GCK(pe_1_2_4_net5967) );
  CLKGATETST_X1 pe_1_2_4_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_2_4_N62), .SE(1'b0), .GCK(pe_1_2_4_net5972) );
  CLKGATETST_X1 pe_1_2_4_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_2_4_N61), .SE(1'b0), .GCK(pe_1_2_4_net5977) );
  CLKGATETST_X1 pe_1_2_4_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_2_4_N60), .SE(1'b0), .GCK(pe_1_2_4_net5982) );
  CLKGATETST_X1 pe_1_2_4_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_2_4_N59), .SE(1'b0), .GCK(pe_1_2_4_net5987) );
  CLKGATETST_X1 pe_1_2_4_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_2_4_N90), .SE(1'b0), .GCK(pe_1_2_4_net5992) );
  CLKBUF_X1 pe_1_2_5_U112 ( .A(pe_1_2_5_n72), .Z(pe_1_2_5_n71) );
  INV_X1 pe_1_2_5_U111 ( .A(n74), .ZN(pe_1_2_5_n70) );
  INV_X1 pe_1_2_5_U110 ( .A(n66), .ZN(pe_1_2_5_n69) );
  INV_X1 pe_1_2_5_U109 ( .A(n66), .ZN(pe_1_2_5_n68) );
  INV_X1 pe_1_2_5_U108 ( .A(n66), .ZN(pe_1_2_5_n67) );
  INV_X1 pe_1_2_5_U107 ( .A(pe_1_2_5_n69), .ZN(pe_1_2_5_n66) );
  INV_X1 pe_1_2_5_U106 ( .A(pe_1_2_5_n63), .ZN(pe_1_2_5_n62) );
  INV_X1 pe_1_2_5_U105 ( .A(pe_1_2_5_n61), .ZN(pe_1_2_5_n60) );
  INV_X1 pe_1_2_5_U104 ( .A(n26), .ZN(pe_1_2_5_n59) );
  INV_X1 pe_1_2_5_U103 ( .A(pe_1_2_5_n59), .ZN(pe_1_2_5_n58) );
  INV_X1 pe_1_2_5_U102 ( .A(n18), .ZN(pe_1_2_5_n57) );
  MUX2_X1 pe_1_2_5_U101 ( .A(pe_1_2_5_n54), .B(pe_1_2_5_n51), .S(n47), .Z(
        int_data_x_2__5__3_) );
  MUX2_X1 pe_1_2_5_U100 ( .A(pe_1_2_5_n53), .B(pe_1_2_5_n52), .S(pe_1_2_5_n62), 
        .Z(pe_1_2_5_n54) );
  MUX2_X1 pe_1_2_5_U99 ( .A(pe_1_2_5_int_q_reg_h[23]), .B(
        pe_1_2_5_int_q_reg_h[19]), .S(pe_1_2_5_n56), .Z(pe_1_2_5_n53) );
  MUX2_X1 pe_1_2_5_U98 ( .A(pe_1_2_5_int_q_reg_h[15]), .B(
        pe_1_2_5_int_q_reg_h[11]), .S(pe_1_2_5_n56), .Z(pe_1_2_5_n52) );
  MUX2_X1 pe_1_2_5_U97 ( .A(pe_1_2_5_int_q_reg_h[7]), .B(
        pe_1_2_5_int_q_reg_h[3]), .S(pe_1_2_5_n56), .Z(pe_1_2_5_n51) );
  MUX2_X1 pe_1_2_5_U96 ( .A(pe_1_2_5_n50), .B(pe_1_2_5_n47), .S(n47), .Z(
        int_data_x_2__5__2_) );
  MUX2_X1 pe_1_2_5_U95 ( .A(pe_1_2_5_n49), .B(pe_1_2_5_n48), .S(pe_1_2_5_n62), 
        .Z(pe_1_2_5_n50) );
  MUX2_X1 pe_1_2_5_U94 ( .A(pe_1_2_5_int_q_reg_h[22]), .B(
        pe_1_2_5_int_q_reg_h[18]), .S(pe_1_2_5_n56), .Z(pe_1_2_5_n49) );
  MUX2_X1 pe_1_2_5_U93 ( .A(pe_1_2_5_int_q_reg_h[14]), .B(
        pe_1_2_5_int_q_reg_h[10]), .S(pe_1_2_5_n56), .Z(pe_1_2_5_n48) );
  MUX2_X1 pe_1_2_5_U92 ( .A(pe_1_2_5_int_q_reg_h[6]), .B(
        pe_1_2_5_int_q_reg_h[2]), .S(pe_1_2_5_n56), .Z(pe_1_2_5_n47) );
  MUX2_X1 pe_1_2_5_U91 ( .A(pe_1_2_5_n46), .B(pe_1_2_5_n24), .S(n47), .Z(
        int_data_x_2__5__1_) );
  MUX2_X1 pe_1_2_5_U90 ( .A(pe_1_2_5_n45), .B(pe_1_2_5_n25), .S(pe_1_2_5_n62), 
        .Z(pe_1_2_5_n46) );
  MUX2_X1 pe_1_2_5_U89 ( .A(pe_1_2_5_int_q_reg_h[21]), .B(
        pe_1_2_5_int_q_reg_h[17]), .S(pe_1_2_5_n56), .Z(pe_1_2_5_n45) );
  MUX2_X1 pe_1_2_5_U88 ( .A(pe_1_2_5_int_q_reg_h[13]), .B(
        pe_1_2_5_int_q_reg_h[9]), .S(pe_1_2_5_n56), .Z(pe_1_2_5_n25) );
  MUX2_X1 pe_1_2_5_U87 ( .A(pe_1_2_5_int_q_reg_h[5]), .B(
        pe_1_2_5_int_q_reg_h[1]), .S(pe_1_2_5_n56), .Z(pe_1_2_5_n24) );
  MUX2_X1 pe_1_2_5_U86 ( .A(pe_1_2_5_n23), .B(pe_1_2_5_n20), .S(n47), .Z(
        int_data_x_2__5__0_) );
  MUX2_X1 pe_1_2_5_U85 ( .A(pe_1_2_5_n22), .B(pe_1_2_5_n21), .S(pe_1_2_5_n62), 
        .Z(pe_1_2_5_n23) );
  MUX2_X1 pe_1_2_5_U84 ( .A(pe_1_2_5_int_q_reg_h[20]), .B(
        pe_1_2_5_int_q_reg_h[16]), .S(pe_1_2_5_n56), .Z(pe_1_2_5_n22) );
  MUX2_X1 pe_1_2_5_U83 ( .A(pe_1_2_5_int_q_reg_h[12]), .B(
        pe_1_2_5_int_q_reg_h[8]), .S(pe_1_2_5_n56), .Z(pe_1_2_5_n21) );
  MUX2_X1 pe_1_2_5_U82 ( .A(pe_1_2_5_int_q_reg_h[4]), .B(
        pe_1_2_5_int_q_reg_h[0]), .S(pe_1_2_5_n56), .Z(pe_1_2_5_n20) );
  MUX2_X1 pe_1_2_5_U81 ( .A(pe_1_2_5_n19), .B(pe_1_2_5_n16), .S(n47), .Z(
        int_data_y_2__5__3_) );
  MUX2_X1 pe_1_2_5_U80 ( .A(pe_1_2_5_n18), .B(pe_1_2_5_n17), .S(pe_1_2_5_n62), 
        .Z(pe_1_2_5_n19) );
  MUX2_X1 pe_1_2_5_U79 ( .A(pe_1_2_5_int_q_reg_v[23]), .B(
        pe_1_2_5_int_q_reg_v[19]), .S(pe_1_2_5_n55), .Z(pe_1_2_5_n18) );
  MUX2_X1 pe_1_2_5_U78 ( .A(pe_1_2_5_int_q_reg_v[15]), .B(
        pe_1_2_5_int_q_reg_v[11]), .S(pe_1_2_5_n55), .Z(pe_1_2_5_n17) );
  MUX2_X1 pe_1_2_5_U77 ( .A(pe_1_2_5_int_q_reg_v[7]), .B(
        pe_1_2_5_int_q_reg_v[3]), .S(pe_1_2_5_n55), .Z(pe_1_2_5_n16) );
  MUX2_X1 pe_1_2_5_U76 ( .A(pe_1_2_5_n15), .B(pe_1_2_5_n12), .S(n47), .Z(
        int_data_y_2__5__2_) );
  MUX2_X1 pe_1_2_5_U75 ( .A(pe_1_2_5_n14), .B(pe_1_2_5_n13), .S(pe_1_2_5_n62), 
        .Z(pe_1_2_5_n15) );
  MUX2_X1 pe_1_2_5_U74 ( .A(pe_1_2_5_int_q_reg_v[22]), .B(
        pe_1_2_5_int_q_reg_v[18]), .S(pe_1_2_5_n55), .Z(pe_1_2_5_n14) );
  MUX2_X1 pe_1_2_5_U73 ( .A(pe_1_2_5_int_q_reg_v[14]), .B(
        pe_1_2_5_int_q_reg_v[10]), .S(pe_1_2_5_n55), .Z(pe_1_2_5_n13) );
  MUX2_X1 pe_1_2_5_U72 ( .A(pe_1_2_5_int_q_reg_v[6]), .B(
        pe_1_2_5_int_q_reg_v[2]), .S(pe_1_2_5_n55), .Z(pe_1_2_5_n12) );
  MUX2_X1 pe_1_2_5_U71 ( .A(pe_1_2_5_n11), .B(pe_1_2_5_n8), .S(n47), .Z(
        int_data_y_2__5__1_) );
  MUX2_X1 pe_1_2_5_U70 ( .A(pe_1_2_5_n10), .B(pe_1_2_5_n9), .S(pe_1_2_5_n62), 
        .Z(pe_1_2_5_n11) );
  MUX2_X1 pe_1_2_5_U69 ( .A(pe_1_2_5_int_q_reg_v[21]), .B(
        pe_1_2_5_int_q_reg_v[17]), .S(pe_1_2_5_n55), .Z(pe_1_2_5_n10) );
  MUX2_X1 pe_1_2_5_U68 ( .A(pe_1_2_5_int_q_reg_v[13]), .B(
        pe_1_2_5_int_q_reg_v[9]), .S(pe_1_2_5_n55), .Z(pe_1_2_5_n9) );
  MUX2_X1 pe_1_2_5_U67 ( .A(pe_1_2_5_int_q_reg_v[5]), .B(
        pe_1_2_5_int_q_reg_v[1]), .S(pe_1_2_5_n55), .Z(pe_1_2_5_n8) );
  MUX2_X1 pe_1_2_5_U66 ( .A(pe_1_2_5_n7), .B(pe_1_2_5_n4), .S(n47), .Z(
        int_data_y_2__5__0_) );
  MUX2_X1 pe_1_2_5_U65 ( .A(pe_1_2_5_n6), .B(pe_1_2_5_n5), .S(pe_1_2_5_n62), 
        .Z(pe_1_2_5_n7) );
  MUX2_X1 pe_1_2_5_U64 ( .A(pe_1_2_5_int_q_reg_v[20]), .B(
        pe_1_2_5_int_q_reg_v[16]), .S(pe_1_2_5_n55), .Z(pe_1_2_5_n6) );
  MUX2_X1 pe_1_2_5_U63 ( .A(pe_1_2_5_int_q_reg_v[12]), .B(
        pe_1_2_5_int_q_reg_v[8]), .S(pe_1_2_5_n55), .Z(pe_1_2_5_n5) );
  MUX2_X1 pe_1_2_5_U62 ( .A(pe_1_2_5_int_q_reg_v[4]), .B(
        pe_1_2_5_int_q_reg_v[0]), .S(pe_1_2_5_n55), .Z(pe_1_2_5_n4) );
  AOI222_X1 pe_1_2_5_U61 ( .A1(int_data_res_3__5__2_), .A2(pe_1_2_5_n64), .B1(
        pe_1_2_5_N80), .B2(pe_1_2_5_n27), .C1(pe_1_2_5_N72), .C2(pe_1_2_5_n28), 
        .ZN(pe_1_2_5_n33) );
  INV_X1 pe_1_2_5_U60 ( .A(pe_1_2_5_n33), .ZN(pe_1_2_5_n82) );
  AOI222_X1 pe_1_2_5_U59 ( .A1(int_data_res_3__5__6_), .A2(pe_1_2_5_n64), .B1(
        pe_1_2_5_N84), .B2(pe_1_2_5_n27), .C1(pe_1_2_5_N76), .C2(pe_1_2_5_n28), 
        .ZN(pe_1_2_5_n29) );
  INV_X1 pe_1_2_5_U58 ( .A(pe_1_2_5_n29), .ZN(pe_1_2_5_n78) );
  XNOR2_X1 pe_1_2_5_U57 ( .A(pe_1_2_5_n73), .B(int_data_res_2__5__0_), .ZN(
        pe_1_2_5_N70) );
  AOI222_X1 pe_1_2_5_U52 ( .A1(int_data_res_3__5__0_), .A2(pe_1_2_5_n64), .B1(
        pe_1_2_5_n1), .B2(pe_1_2_5_n27), .C1(pe_1_2_5_N70), .C2(pe_1_2_5_n28), 
        .ZN(pe_1_2_5_n35) );
  INV_X1 pe_1_2_5_U51 ( .A(pe_1_2_5_n35), .ZN(pe_1_2_5_n84) );
  AOI222_X1 pe_1_2_5_U50 ( .A1(int_data_res_3__5__1_), .A2(pe_1_2_5_n64), .B1(
        pe_1_2_5_N79), .B2(pe_1_2_5_n27), .C1(pe_1_2_5_N71), .C2(pe_1_2_5_n28), 
        .ZN(pe_1_2_5_n34) );
  INV_X1 pe_1_2_5_U49 ( .A(pe_1_2_5_n34), .ZN(pe_1_2_5_n83) );
  AOI222_X1 pe_1_2_5_U48 ( .A1(int_data_res_3__5__3_), .A2(pe_1_2_5_n64), .B1(
        pe_1_2_5_N81), .B2(pe_1_2_5_n27), .C1(pe_1_2_5_N73), .C2(pe_1_2_5_n28), 
        .ZN(pe_1_2_5_n32) );
  INV_X1 pe_1_2_5_U47 ( .A(pe_1_2_5_n32), .ZN(pe_1_2_5_n81) );
  AOI222_X1 pe_1_2_5_U46 ( .A1(int_data_res_3__5__4_), .A2(pe_1_2_5_n64), .B1(
        pe_1_2_5_N82), .B2(pe_1_2_5_n27), .C1(pe_1_2_5_N74), .C2(pe_1_2_5_n28), 
        .ZN(pe_1_2_5_n31) );
  INV_X1 pe_1_2_5_U45 ( .A(pe_1_2_5_n31), .ZN(pe_1_2_5_n80) );
  AOI222_X1 pe_1_2_5_U44 ( .A1(int_data_res_3__5__5_), .A2(pe_1_2_5_n64), .B1(
        pe_1_2_5_N83), .B2(pe_1_2_5_n27), .C1(pe_1_2_5_N75), .C2(pe_1_2_5_n28), 
        .ZN(pe_1_2_5_n30) );
  INV_X1 pe_1_2_5_U43 ( .A(pe_1_2_5_n30), .ZN(pe_1_2_5_n79) );
  NAND2_X1 pe_1_2_5_U42 ( .A1(pe_1_2_5_int_data_0_), .A2(pe_1_2_5_n3), .ZN(
        pe_1_2_5_sub_81_carry[1]) );
  INV_X1 pe_1_2_5_U41 ( .A(pe_1_2_5_int_data_1_), .ZN(pe_1_2_5_n74) );
  INV_X1 pe_1_2_5_U40 ( .A(pe_1_2_5_int_data_2_), .ZN(pe_1_2_5_n75) );
  AND2_X1 pe_1_2_5_U39 ( .A1(pe_1_2_5_int_data_0_), .A2(int_data_res_2__5__0_), 
        .ZN(pe_1_2_5_n2) );
  AOI222_X1 pe_1_2_5_U38 ( .A1(pe_1_2_5_n64), .A2(int_data_res_3__5__7_), .B1(
        pe_1_2_5_N85), .B2(pe_1_2_5_n27), .C1(pe_1_2_5_N77), .C2(pe_1_2_5_n28), 
        .ZN(pe_1_2_5_n26) );
  INV_X1 pe_1_2_5_U37 ( .A(pe_1_2_5_n26), .ZN(pe_1_2_5_n77) );
  NOR3_X1 pe_1_2_5_U36 ( .A1(pe_1_2_5_n59), .A2(pe_1_2_5_n65), .A3(int_ckg[42]), .ZN(pe_1_2_5_n36) );
  OR2_X1 pe_1_2_5_U35 ( .A1(pe_1_2_5_n36), .A2(pe_1_2_5_n64), .ZN(pe_1_2_5_N90) );
  INV_X1 pe_1_2_5_U34 ( .A(n38), .ZN(pe_1_2_5_n63) );
  AND2_X1 pe_1_2_5_U33 ( .A1(int_data_x_2__5__2_), .A2(pe_1_2_5_n58), .ZN(
        pe_1_2_5_int_data_2_) );
  AND2_X1 pe_1_2_5_U32 ( .A1(int_data_x_2__5__1_), .A2(pe_1_2_5_n58), .ZN(
        pe_1_2_5_int_data_1_) );
  AND2_X1 pe_1_2_5_U31 ( .A1(int_data_x_2__5__3_), .A2(pe_1_2_5_n58), .ZN(
        pe_1_2_5_int_data_3_) );
  BUF_X1 pe_1_2_5_U30 ( .A(n60), .Z(pe_1_2_5_n64) );
  INV_X1 pe_1_2_5_U29 ( .A(n32), .ZN(pe_1_2_5_n61) );
  AND2_X1 pe_1_2_5_U28 ( .A1(int_data_x_2__5__0_), .A2(pe_1_2_5_n58), .ZN(
        pe_1_2_5_int_data_0_) );
  NAND2_X1 pe_1_2_5_U27 ( .A1(pe_1_2_5_n44), .A2(pe_1_2_5_n61), .ZN(
        pe_1_2_5_n41) );
  AND3_X1 pe_1_2_5_U26 ( .A1(n74), .A2(pe_1_2_5_n63), .A3(n47), .ZN(
        pe_1_2_5_n44) );
  INV_X1 pe_1_2_5_U25 ( .A(pe_1_2_5_int_data_3_), .ZN(pe_1_2_5_n76) );
  NOR2_X1 pe_1_2_5_U24 ( .A1(pe_1_2_5_n70), .A2(n47), .ZN(pe_1_2_5_n43) );
  NOR2_X1 pe_1_2_5_U23 ( .A1(pe_1_2_5_n57), .A2(pe_1_2_5_n64), .ZN(
        pe_1_2_5_n28) );
  NOR2_X1 pe_1_2_5_U22 ( .A1(n18), .A2(pe_1_2_5_n64), .ZN(pe_1_2_5_n27) );
  INV_X1 pe_1_2_5_U21 ( .A(pe_1_2_5_int_data_0_), .ZN(pe_1_2_5_n73) );
  INV_X1 pe_1_2_5_U20 ( .A(pe_1_2_5_n41), .ZN(pe_1_2_5_n90) );
  INV_X1 pe_1_2_5_U19 ( .A(pe_1_2_5_n37), .ZN(pe_1_2_5_n88) );
  INV_X1 pe_1_2_5_U18 ( .A(pe_1_2_5_n38), .ZN(pe_1_2_5_n87) );
  INV_X1 pe_1_2_5_U17 ( .A(pe_1_2_5_n39), .ZN(pe_1_2_5_n86) );
  NOR2_X1 pe_1_2_5_U16 ( .A1(pe_1_2_5_n68), .A2(pe_1_2_5_n42), .ZN(
        pe_1_2_5_N59) );
  NOR2_X1 pe_1_2_5_U15 ( .A1(pe_1_2_5_n68), .A2(pe_1_2_5_n41), .ZN(
        pe_1_2_5_N60) );
  NOR2_X1 pe_1_2_5_U14 ( .A1(pe_1_2_5_n68), .A2(pe_1_2_5_n38), .ZN(
        pe_1_2_5_N63) );
  NOR2_X1 pe_1_2_5_U13 ( .A1(pe_1_2_5_n67), .A2(pe_1_2_5_n40), .ZN(
        pe_1_2_5_N61) );
  NOR2_X1 pe_1_2_5_U12 ( .A1(pe_1_2_5_n67), .A2(pe_1_2_5_n39), .ZN(
        pe_1_2_5_N62) );
  NOR2_X1 pe_1_2_5_U11 ( .A1(pe_1_2_5_n37), .A2(pe_1_2_5_n67), .ZN(
        pe_1_2_5_N64) );
  NAND2_X1 pe_1_2_5_U10 ( .A1(pe_1_2_5_n44), .A2(pe_1_2_5_n60), .ZN(
        pe_1_2_5_n42) );
  BUF_X1 pe_1_2_5_U9 ( .A(pe_1_2_5_n60), .Z(pe_1_2_5_n55) );
  INV_X1 pe_1_2_5_U8 ( .A(pe_1_2_5_n69), .ZN(pe_1_2_5_n65) );
  BUF_X1 pe_1_2_5_U7 ( .A(pe_1_2_5_n60), .Z(pe_1_2_5_n56) );
  INV_X1 pe_1_2_5_U6 ( .A(pe_1_2_5_n42), .ZN(pe_1_2_5_n89) );
  INV_X1 pe_1_2_5_U5 ( .A(pe_1_2_5_n40), .ZN(pe_1_2_5_n85) );
  INV_X2 pe_1_2_5_U4 ( .A(n82), .ZN(pe_1_2_5_n72) );
  XOR2_X1 pe_1_2_5_U3 ( .A(pe_1_2_5_int_data_0_), .B(int_data_res_2__5__0_), 
        .Z(pe_1_2_5_n1) );
  DFFR_X1 pe_1_2_5_int_q_acc_reg_0_ ( .D(pe_1_2_5_n84), .CK(pe_1_2_5_net5914), 
        .RN(pe_1_2_5_n72), .Q(int_data_res_2__5__0_), .QN(pe_1_2_5_n3) );
  DFFR_X1 pe_1_2_5_int_q_reg_v_reg_0__0_ ( .D(int_data_y_3__5__0_), .CK(
        pe_1_2_5_net5884), .RN(pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_v[20]) );
  DFFR_X1 pe_1_2_5_int_q_reg_v_reg_0__1_ ( .D(int_data_y_3__5__1_), .CK(
        pe_1_2_5_net5884), .RN(pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_v[21]) );
  DFFR_X1 pe_1_2_5_int_q_reg_v_reg_0__2_ ( .D(int_data_y_3__5__2_), .CK(
        pe_1_2_5_net5884), .RN(pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_v[22]) );
  DFFR_X1 pe_1_2_5_int_q_reg_v_reg_0__3_ ( .D(int_data_y_3__5__3_), .CK(
        pe_1_2_5_net5884), .RN(pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_v[23]) );
  DFFR_X1 pe_1_2_5_int_q_reg_v_reg_1__0_ ( .D(int_data_y_3__5__0_), .CK(
        pe_1_2_5_net5889), .RN(pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_v[16]) );
  DFFR_X1 pe_1_2_5_int_q_reg_v_reg_1__1_ ( .D(int_data_y_3__5__1_), .CK(
        pe_1_2_5_net5889), .RN(pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_v[17]) );
  DFFR_X1 pe_1_2_5_int_q_reg_v_reg_1__2_ ( .D(int_data_y_3__5__2_), .CK(
        pe_1_2_5_net5889), .RN(pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_v[18]) );
  DFFR_X1 pe_1_2_5_int_q_reg_v_reg_1__3_ ( .D(int_data_y_3__5__3_), .CK(
        pe_1_2_5_net5889), .RN(pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_v[19]) );
  DFFR_X1 pe_1_2_5_int_q_reg_v_reg_2__0_ ( .D(int_data_y_3__5__0_), .CK(
        pe_1_2_5_net5894), .RN(pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_v[12]) );
  DFFR_X1 pe_1_2_5_int_q_reg_v_reg_2__1_ ( .D(int_data_y_3__5__1_), .CK(
        pe_1_2_5_net5894), .RN(pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_v[13]) );
  DFFR_X1 pe_1_2_5_int_q_reg_v_reg_2__2_ ( .D(int_data_y_3__5__2_), .CK(
        pe_1_2_5_net5894), .RN(pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_v[14]) );
  DFFR_X1 pe_1_2_5_int_q_reg_v_reg_2__3_ ( .D(int_data_y_3__5__3_), .CK(
        pe_1_2_5_net5894), .RN(pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_v[15]) );
  DFFR_X1 pe_1_2_5_int_q_reg_v_reg_3__0_ ( .D(int_data_y_3__5__0_), .CK(
        pe_1_2_5_net5899), .RN(pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_v[8]) );
  DFFR_X1 pe_1_2_5_int_q_reg_v_reg_3__1_ ( .D(int_data_y_3__5__1_), .CK(
        pe_1_2_5_net5899), .RN(pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_v[9]) );
  DFFR_X1 pe_1_2_5_int_q_reg_v_reg_3__2_ ( .D(int_data_y_3__5__2_), .CK(
        pe_1_2_5_net5899), .RN(pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_v[10]) );
  DFFR_X1 pe_1_2_5_int_q_reg_v_reg_3__3_ ( .D(int_data_y_3__5__3_), .CK(
        pe_1_2_5_net5899), .RN(pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_v[11]) );
  DFFR_X1 pe_1_2_5_int_q_reg_v_reg_4__0_ ( .D(int_data_y_3__5__0_), .CK(
        pe_1_2_5_net5904), .RN(pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_v[4]) );
  DFFR_X1 pe_1_2_5_int_q_reg_v_reg_4__1_ ( .D(int_data_y_3__5__1_), .CK(
        pe_1_2_5_net5904), .RN(pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_v[5]) );
  DFFR_X1 pe_1_2_5_int_q_reg_v_reg_4__2_ ( .D(int_data_y_3__5__2_), .CK(
        pe_1_2_5_net5904), .RN(pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_v[6]) );
  DFFR_X1 pe_1_2_5_int_q_reg_v_reg_4__3_ ( .D(int_data_y_3__5__3_), .CK(
        pe_1_2_5_net5904), .RN(pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_v[7]) );
  DFFR_X1 pe_1_2_5_int_q_reg_v_reg_5__0_ ( .D(int_data_y_3__5__0_), .CK(
        pe_1_2_5_net5909), .RN(pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_v[0]) );
  DFFR_X1 pe_1_2_5_int_q_reg_v_reg_5__1_ ( .D(int_data_y_3__5__1_), .CK(
        pe_1_2_5_net5909), .RN(pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_v[1]) );
  DFFR_X1 pe_1_2_5_int_q_reg_v_reg_5__2_ ( .D(int_data_y_3__5__2_), .CK(
        pe_1_2_5_net5909), .RN(pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_v[2]) );
  DFFR_X1 pe_1_2_5_int_q_reg_v_reg_5__3_ ( .D(int_data_y_3__5__3_), .CK(
        pe_1_2_5_net5909), .RN(pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_2_5_int_q_reg_h_reg_0__0_ ( .D(int_data_x_2__6__0_), .SI(
        int_data_y_3__5__0_), .SE(pe_1_2_5_n65), .CK(pe_1_2_5_net5853), .RN(
        pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_2_5_int_q_reg_h_reg_0__1_ ( .D(int_data_x_2__6__1_), .SI(
        int_data_y_3__5__1_), .SE(pe_1_2_5_n65), .CK(pe_1_2_5_net5853), .RN(
        pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_2_5_int_q_reg_h_reg_0__2_ ( .D(int_data_x_2__6__2_), .SI(
        int_data_y_3__5__2_), .SE(pe_1_2_5_n65), .CK(pe_1_2_5_net5853), .RN(
        pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_2_5_int_q_reg_h_reg_0__3_ ( .D(int_data_x_2__6__3_), .SI(
        int_data_y_3__5__3_), .SE(pe_1_2_5_n65), .CK(pe_1_2_5_net5853), .RN(
        pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_2_5_int_q_reg_h_reg_1__0_ ( .D(int_data_x_2__6__0_), .SI(
        int_data_y_3__5__0_), .SE(pe_1_2_5_n65), .CK(pe_1_2_5_net5859), .RN(
        pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_2_5_int_q_reg_h_reg_1__1_ ( .D(int_data_x_2__6__1_), .SI(
        int_data_y_3__5__1_), .SE(pe_1_2_5_n65), .CK(pe_1_2_5_net5859), .RN(
        pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_2_5_int_q_reg_h_reg_1__2_ ( .D(int_data_x_2__6__2_), .SI(
        int_data_y_3__5__2_), .SE(pe_1_2_5_n65), .CK(pe_1_2_5_net5859), .RN(
        pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_2_5_int_q_reg_h_reg_1__3_ ( .D(int_data_x_2__6__3_), .SI(
        int_data_y_3__5__3_), .SE(pe_1_2_5_n65), .CK(pe_1_2_5_net5859), .RN(
        pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_2_5_int_q_reg_h_reg_2__0_ ( .D(int_data_x_2__6__0_), .SI(
        int_data_y_3__5__0_), .SE(pe_1_2_5_n65), .CK(pe_1_2_5_net5864), .RN(
        pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_2_5_int_q_reg_h_reg_2__1_ ( .D(int_data_x_2__6__1_), .SI(
        int_data_y_3__5__1_), .SE(pe_1_2_5_n65), .CK(pe_1_2_5_net5864), .RN(
        pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_2_5_int_q_reg_h_reg_2__2_ ( .D(int_data_x_2__6__2_), .SI(
        int_data_y_3__5__2_), .SE(pe_1_2_5_n65), .CK(pe_1_2_5_net5864), .RN(
        pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_2_5_int_q_reg_h_reg_2__3_ ( .D(int_data_x_2__6__3_), .SI(
        int_data_y_3__5__3_), .SE(pe_1_2_5_n65), .CK(pe_1_2_5_net5864), .RN(
        pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_2_5_int_q_reg_h_reg_3__0_ ( .D(int_data_x_2__6__0_), .SI(
        int_data_y_3__5__0_), .SE(pe_1_2_5_n65), .CK(pe_1_2_5_net5869), .RN(
        pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_2_5_int_q_reg_h_reg_3__1_ ( .D(int_data_x_2__6__1_), .SI(
        int_data_y_3__5__1_), .SE(pe_1_2_5_n65), .CK(pe_1_2_5_net5869), .RN(
        pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_2_5_int_q_reg_h_reg_3__2_ ( .D(int_data_x_2__6__2_), .SI(
        int_data_y_3__5__2_), .SE(pe_1_2_5_n65), .CK(pe_1_2_5_net5869), .RN(
        pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_2_5_int_q_reg_h_reg_3__3_ ( .D(int_data_x_2__6__3_), .SI(
        int_data_y_3__5__3_), .SE(pe_1_2_5_n65), .CK(pe_1_2_5_net5869), .RN(
        pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_2_5_int_q_reg_h_reg_4__0_ ( .D(int_data_x_2__6__0_), .SI(
        int_data_y_3__5__0_), .SE(pe_1_2_5_n66), .CK(pe_1_2_5_net5874), .RN(
        pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_2_5_int_q_reg_h_reg_4__1_ ( .D(int_data_x_2__6__1_), .SI(
        int_data_y_3__5__1_), .SE(pe_1_2_5_n66), .CK(pe_1_2_5_net5874), .RN(
        pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_2_5_int_q_reg_h_reg_4__2_ ( .D(int_data_x_2__6__2_), .SI(
        int_data_y_3__5__2_), .SE(pe_1_2_5_n66), .CK(pe_1_2_5_net5874), .RN(
        pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_2_5_int_q_reg_h_reg_4__3_ ( .D(int_data_x_2__6__3_), .SI(
        int_data_y_3__5__3_), .SE(pe_1_2_5_n66), .CK(pe_1_2_5_net5874), .RN(
        pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_2_5_int_q_reg_h_reg_5__0_ ( .D(int_data_x_2__6__0_), .SI(
        int_data_y_3__5__0_), .SE(pe_1_2_5_n66), .CK(pe_1_2_5_net5879), .RN(
        pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_2_5_int_q_reg_h_reg_5__1_ ( .D(int_data_x_2__6__1_), .SI(
        int_data_y_3__5__1_), .SE(pe_1_2_5_n66), .CK(pe_1_2_5_net5879), .RN(
        pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_2_5_int_q_reg_h_reg_5__2_ ( .D(int_data_x_2__6__2_), .SI(
        int_data_y_3__5__2_), .SE(pe_1_2_5_n66), .CK(pe_1_2_5_net5879), .RN(
        pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_2_5_int_q_reg_h_reg_5__3_ ( .D(int_data_x_2__6__3_), .SI(
        int_data_y_3__5__3_), .SE(pe_1_2_5_n66), .CK(pe_1_2_5_net5879), .RN(
        pe_1_2_5_n72), .Q(pe_1_2_5_int_q_reg_h[3]) );
  FA_X1 pe_1_2_5_sub_81_U2_7 ( .A(int_data_res_2__5__7_), .B(pe_1_2_5_n76), 
        .CI(pe_1_2_5_sub_81_carry[7]), .S(pe_1_2_5_N77) );
  FA_X1 pe_1_2_5_sub_81_U2_6 ( .A(int_data_res_2__5__6_), .B(pe_1_2_5_n76), 
        .CI(pe_1_2_5_sub_81_carry[6]), .CO(pe_1_2_5_sub_81_carry[7]), .S(
        pe_1_2_5_N76) );
  FA_X1 pe_1_2_5_sub_81_U2_5 ( .A(int_data_res_2__5__5_), .B(pe_1_2_5_n76), 
        .CI(pe_1_2_5_sub_81_carry[5]), .CO(pe_1_2_5_sub_81_carry[6]), .S(
        pe_1_2_5_N75) );
  FA_X1 pe_1_2_5_sub_81_U2_4 ( .A(int_data_res_2__5__4_), .B(pe_1_2_5_n76), 
        .CI(pe_1_2_5_sub_81_carry[4]), .CO(pe_1_2_5_sub_81_carry[5]), .S(
        pe_1_2_5_N74) );
  FA_X1 pe_1_2_5_sub_81_U2_3 ( .A(int_data_res_2__5__3_), .B(pe_1_2_5_n76), 
        .CI(pe_1_2_5_sub_81_carry[3]), .CO(pe_1_2_5_sub_81_carry[4]), .S(
        pe_1_2_5_N73) );
  FA_X1 pe_1_2_5_sub_81_U2_2 ( .A(int_data_res_2__5__2_), .B(pe_1_2_5_n75), 
        .CI(pe_1_2_5_sub_81_carry[2]), .CO(pe_1_2_5_sub_81_carry[3]), .S(
        pe_1_2_5_N72) );
  FA_X1 pe_1_2_5_sub_81_U2_1 ( .A(int_data_res_2__5__1_), .B(pe_1_2_5_n74), 
        .CI(pe_1_2_5_sub_81_carry[1]), .CO(pe_1_2_5_sub_81_carry[2]), .S(
        pe_1_2_5_N71) );
  FA_X1 pe_1_2_5_add_83_U1_7 ( .A(int_data_res_2__5__7_), .B(
        pe_1_2_5_int_data_3_), .CI(pe_1_2_5_add_83_carry[7]), .S(pe_1_2_5_N85)
         );
  FA_X1 pe_1_2_5_add_83_U1_6 ( .A(int_data_res_2__5__6_), .B(
        pe_1_2_5_int_data_3_), .CI(pe_1_2_5_add_83_carry[6]), .CO(
        pe_1_2_5_add_83_carry[7]), .S(pe_1_2_5_N84) );
  FA_X1 pe_1_2_5_add_83_U1_5 ( .A(int_data_res_2__5__5_), .B(
        pe_1_2_5_int_data_3_), .CI(pe_1_2_5_add_83_carry[5]), .CO(
        pe_1_2_5_add_83_carry[6]), .S(pe_1_2_5_N83) );
  FA_X1 pe_1_2_5_add_83_U1_4 ( .A(int_data_res_2__5__4_), .B(
        pe_1_2_5_int_data_3_), .CI(pe_1_2_5_add_83_carry[4]), .CO(
        pe_1_2_5_add_83_carry[5]), .S(pe_1_2_5_N82) );
  FA_X1 pe_1_2_5_add_83_U1_3 ( .A(int_data_res_2__5__3_), .B(
        pe_1_2_5_int_data_3_), .CI(pe_1_2_5_add_83_carry[3]), .CO(
        pe_1_2_5_add_83_carry[4]), .S(pe_1_2_5_N81) );
  FA_X1 pe_1_2_5_add_83_U1_2 ( .A(int_data_res_2__5__2_), .B(
        pe_1_2_5_int_data_2_), .CI(pe_1_2_5_add_83_carry[2]), .CO(
        pe_1_2_5_add_83_carry[3]), .S(pe_1_2_5_N80) );
  FA_X1 pe_1_2_5_add_83_U1_1 ( .A(int_data_res_2__5__1_), .B(
        pe_1_2_5_int_data_1_), .CI(pe_1_2_5_n2), .CO(pe_1_2_5_add_83_carry[2]), 
        .S(pe_1_2_5_N79) );
  NAND3_X1 pe_1_2_5_U56 ( .A1(pe_1_2_5_n60), .A2(pe_1_2_5_n43), .A3(
        pe_1_2_5_n62), .ZN(pe_1_2_5_n40) );
  NAND3_X1 pe_1_2_5_U55 ( .A1(pe_1_2_5_n43), .A2(pe_1_2_5_n61), .A3(
        pe_1_2_5_n62), .ZN(pe_1_2_5_n39) );
  NAND3_X1 pe_1_2_5_U54 ( .A1(pe_1_2_5_n43), .A2(pe_1_2_5_n63), .A3(
        pe_1_2_5_n60), .ZN(pe_1_2_5_n38) );
  NAND3_X1 pe_1_2_5_U53 ( .A1(pe_1_2_5_n61), .A2(pe_1_2_5_n63), .A3(
        pe_1_2_5_n43), .ZN(pe_1_2_5_n37) );
  DFFR_X1 pe_1_2_5_int_q_acc_reg_6_ ( .D(pe_1_2_5_n78), .CK(pe_1_2_5_net5914), 
        .RN(pe_1_2_5_n71), .Q(int_data_res_2__5__6_) );
  DFFR_X1 pe_1_2_5_int_q_acc_reg_5_ ( .D(pe_1_2_5_n79), .CK(pe_1_2_5_net5914), 
        .RN(pe_1_2_5_n71), .Q(int_data_res_2__5__5_) );
  DFFR_X1 pe_1_2_5_int_q_acc_reg_4_ ( .D(pe_1_2_5_n80), .CK(pe_1_2_5_net5914), 
        .RN(pe_1_2_5_n71), .Q(int_data_res_2__5__4_) );
  DFFR_X1 pe_1_2_5_int_q_acc_reg_3_ ( .D(pe_1_2_5_n81), .CK(pe_1_2_5_net5914), 
        .RN(pe_1_2_5_n71), .Q(int_data_res_2__5__3_) );
  DFFR_X1 pe_1_2_5_int_q_acc_reg_2_ ( .D(pe_1_2_5_n82), .CK(pe_1_2_5_net5914), 
        .RN(pe_1_2_5_n71), .Q(int_data_res_2__5__2_) );
  DFFR_X1 pe_1_2_5_int_q_acc_reg_1_ ( .D(pe_1_2_5_n83), .CK(pe_1_2_5_net5914), 
        .RN(pe_1_2_5_n71), .Q(int_data_res_2__5__1_) );
  DFFR_X1 pe_1_2_5_int_q_acc_reg_7_ ( .D(pe_1_2_5_n77), .CK(pe_1_2_5_net5914), 
        .RN(pe_1_2_5_n71), .Q(int_data_res_2__5__7_) );
  CLKGATETST_X1 pe_1_2_5_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_2_5_n88), .SE(1'b0), .GCK(pe_1_2_5_net5853) );
  CLKGATETST_X1 pe_1_2_5_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_2_5_n87), .SE(1'b0), .GCK(pe_1_2_5_net5859) );
  CLKGATETST_X1 pe_1_2_5_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_2_5_n86), .SE(1'b0), .GCK(pe_1_2_5_net5864) );
  CLKGATETST_X1 pe_1_2_5_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_2_5_n85), .SE(1'b0), .GCK(pe_1_2_5_net5869) );
  CLKGATETST_X1 pe_1_2_5_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_2_5_n90), .SE(1'b0), .GCK(pe_1_2_5_net5874) );
  CLKGATETST_X1 pe_1_2_5_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_2_5_n89), .SE(1'b0), .GCK(pe_1_2_5_net5879) );
  CLKGATETST_X1 pe_1_2_5_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_2_5_N64), .SE(1'b0), .GCK(pe_1_2_5_net5884) );
  CLKGATETST_X1 pe_1_2_5_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_2_5_N63), .SE(1'b0), .GCK(pe_1_2_5_net5889) );
  CLKGATETST_X1 pe_1_2_5_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_2_5_N62), .SE(1'b0), .GCK(pe_1_2_5_net5894) );
  CLKGATETST_X1 pe_1_2_5_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_2_5_N61), .SE(1'b0), .GCK(pe_1_2_5_net5899) );
  CLKGATETST_X1 pe_1_2_5_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_2_5_N60), .SE(1'b0), .GCK(pe_1_2_5_net5904) );
  CLKGATETST_X1 pe_1_2_5_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_2_5_N59), .SE(1'b0), .GCK(pe_1_2_5_net5909) );
  CLKGATETST_X1 pe_1_2_5_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_2_5_N90), .SE(1'b0), .GCK(pe_1_2_5_net5914) );
  CLKBUF_X1 pe_1_2_6_U112 ( .A(pe_1_2_6_n72), .Z(pe_1_2_6_n71) );
  INV_X1 pe_1_2_6_U111 ( .A(n74), .ZN(pe_1_2_6_n70) );
  INV_X1 pe_1_2_6_U110 ( .A(n66), .ZN(pe_1_2_6_n69) );
  INV_X1 pe_1_2_6_U109 ( .A(n66), .ZN(pe_1_2_6_n68) );
  INV_X1 pe_1_2_6_U108 ( .A(n66), .ZN(pe_1_2_6_n67) );
  INV_X1 pe_1_2_6_U107 ( .A(pe_1_2_6_n69), .ZN(pe_1_2_6_n66) );
  INV_X1 pe_1_2_6_U106 ( .A(pe_1_2_6_n63), .ZN(pe_1_2_6_n62) );
  INV_X1 pe_1_2_6_U105 ( .A(pe_1_2_6_n61), .ZN(pe_1_2_6_n60) );
  INV_X1 pe_1_2_6_U104 ( .A(n26), .ZN(pe_1_2_6_n59) );
  INV_X1 pe_1_2_6_U103 ( .A(pe_1_2_6_n59), .ZN(pe_1_2_6_n58) );
  INV_X1 pe_1_2_6_U102 ( .A(n18), .ZN(pe_1_2_6_n57) );
  MUX2_X1 pe_1_2_6_U101 ( .A(pe_1_2_6_n54), .B(pe_1_2_6_n51), .S(n47), .Z(
        int_data_x_2__6__3_) );
  MUX2_X1 pe_1_2_6_U100 ( .A(pe_1_2_6_n53), .B(pe_1_2_6_n52), .S(pe_1_2_6_n62), 
        .Z(pe_1_2_6_n54) );
  MUX2_X1 pe_1_2_6_U99 ( .A(pe_1_2_6_int_q_reg_h[23]), .B(
        pe_1_2_6_int_q_reg_h[19]), .S(pe_1_2_6_n56), .Z(pe_1_2_6_n53) );
  MUX2_X1 pe_1_2_6_U98 ( .A(pe_1_2_6_int_q_reg_h[15]), .B(
        pe_1_2_6_int_q_reg_h[11]), .S(pe_1_2_6_n56), .Z(pe_1_2_6_n52) );
  MUX2_X1 pe_1_2_6_U97 ( .A(pe_1_2_6_int_q_reg_h[7]), .B(
        pe_1_2_6_int_q_reg_h[3]), .S(pe_1_2_6_n56), .Z(pe_1_2_6_n51) );
  MUX2_X1 pe_1_2_6_U96 ( .A(pe_1_2_6_n50), .B(pe_1_2_6_n47), .S(n47), .Z(
        int_data_x_2__6__2_) );
  MUX2_X1 pe_1_2_6_U95 ( .A(pe_1_2_6_n49), .B(pe_1_2_6_n48), .S(pe_1_2_6_n62), 
        .Z(pe_1_2_6_n50) );
  MUX2_X1 pe_1_2_6_U94 ( .A(pe_1_2_6_int_q_reg_h[22]), .B(
        pe_1_2_6_int_q_reg_h[18]), .S(pe_1_2_6_n56), .Z(pe_1_2_6_n49) );
  MUX2_X1 pe_1_2_6_U93 ( .A(pe_1_2_6_int_q_reg_h[14]), .B(
        pe_1_2_6_int_q_reg_h[10]), .S(pe_1_2_6_n56), .Z(pe_1_2_6_n48) );
  MUX2_X1 pe_1_2_6_U92 ( .A(pe_1_2_6_int_q_reg_h[6]), .B(
        pe_1_2_6_int_q_reg_h[2]), .S(pe_1_2_6_n56), .Z(pe_1_2_6_n47) );
  MUX2_X1 pe_1_2_6_U91 ( .A(pe_1_2_6_n46), .B(pe_1_2_6_n24), .S(n47), .Z(
        int_data_x_2__6__1_) );
  MUX2_X1 pe_1_2_6_U90 ( .A(pe_1_2_6_n45), .B(pe_1_2_6_n25), .S(pe_1_2_6_n62), 
        .Z(pe_1_2_6_n46) );
  MUX2_X1 pe_1_2_6_U89 ( .A(pe_1_2_6_int_q_reg_h[21]), .B(
        pe_1_2_6_int_q_reg_h[17]), .S(pe_1_2_6_n56), .Z(pe_1_2_6_n45) );
  MUX2_X1 pe_1_2_6_U88 ( .A(pe_1_2_6_int_q_reg_h[13]), .B(
        pe_1_2_6_int_q_reg_h[9]), .S(pe_1_2_6_n56), .Z(pe_1_2_6_n25) );
  MUX2_X1 pe_1_2_6_U87 ( .A(pe_1_2_6_int_q_reg_h[5]), .B(
        pe_1_2_6_int_q_reg_h[1]), .S(pe_1_2_6_n56), .Z(pe_1_2_6_n24) );
  MUX2_X1 pe_1_2_6_U86 ( .A(pe_1_2_6_n23), .B(pe_1_2_6_n20), .S(n47), .Z(
        int_data_x_2__6__0_) );
  MUX2_X1 pe_1_2_6_U85 ( .A(pe_1_2_6_n22), .B(pe_1_2_6_n21), .S(pe_1_2_6_n62), 
        .Z(pe_1_2_6_n23) );
  MUX2_X1 pe_1_2_6_U84 ( .A(pe_1_2_6_int_q_reg_h[20]), .B(
        pe_1_2_6_int_q_reg_h[16]), .S(pe_1_2_6_n56), .Z(pe_1_2_6_n22) );
  MUX2_X1 pe_1_2_6_U83 ( .A(pe_1_2_6_int_q_reg_h[12]), .B(
        pe_1_2_6_int_q_reg_h[8]), .S(pe_1_2_6_n56), .Z(pe_1_2_6_n21) );
  MUX2_X1 pe_1_2_6_U82 ( .A(pe_1_2_6_int_q_reg_h[4]), .B(
        pe_1_2_6_int_q_reg_h[0]), .S(pe_1_2_6_n56), .Z(pe_1_2_6_n20) );
  MUX2_X1 pe_1_2_6_U81 ( .A(pe_1_2_6_n19), .B(pe_1_2_6_n16), .S(n47), .Z(
        int_data_y_2__6__3_) );
  MUX2_X1 pe_1_2_6_U80 ( .A(pe_1_2_6_n18), .B(pe_1_2_6_n17), .S(pe_1_2_6_n62), 
        .Z(pe_1_2_6_n19) );
  MUX2_X1 pe_1_2_6_U79 ( .A(pe_1_2_6_int_q_reg_v[23]), .B(
        pe_1_2_6_int_q_reg_v[19]), .S(pe_1_2_6_n55), .Z(pe_1_2_6_n18) );
  MUX2_X1 pe_1_2_6_U78 ( .A(pe_1_2_6_int_q_reg_v[15]), .B(
        pe_1_2_6_int_q_reg_v[11]), .S(pe_1_2_6_n55), .Z(pe_1_2_6_n17) );
  MUX2_X1 pe_1_2_6_U77 ( .A(pe_1_2_6_int_q_reg_v[7]), .B(
        pe_1_2_6_int_q_reg_v[3]), .S(pe_1_2_6_n55), .Z(pe_1_2_6_n16) );
  MUX2_X1 pe_1_2_6_U76 ( .A(pe_1_2_6_n15), .B(pe_1_2_6_n12), .S(n47), .Z(
        int_data_y_2__6__2_) );
  MUX2_X1 pe_1_2_6_U75 ( .A(pe_1_2_6_n14), .B(pe_1_2_6_n13), .S(pe_1_2_6_n62), 
        .Z(pe_1_2_6_n15) );
  MUX2_X1 pe_1_2_6_U74 ( .A(pe_1_2_6_int_q_reg_v[22]), .B(
        pe_1_2_6_int_q_reg_v[18]), .S(pe_1_2_6_n55), .Z(pe_1_2_6_n14) );
  MUX2_X1 pe_1_2_6_U73 ( .A(pe_1_2_6_int_q_reg_v[14]), .B(
        pe_1_2_6_int_q_reg_v[10]), .S(pe_1_2_6_n55), .Z(pe_1_2_6_n13) );
  MUX2_X1 pe_1_2_6_U72 ( .A(pe_1_2_6_int_q_reg_v[6]), .B(
        pe_1_2_6_int_q_reg_v[2]), .S(pe_1_2_6_n55), .Z(pe_1_2_6_n12) );
  MUX2_X1 pe_1_2_6_U71 ( .A(pe_1_2_6_n11), .B(pe_1_2_6_n8), .S(n47), .Z(
        int_data_y_2__6__1_) );
  MUX2_X1 pe_1_2_6_U70 ( .A(pe_1_2_6_n10), .B(pe_1_2_6_n9), .S(pe_1_2_6_n62), 
        .Z(pe_1_2_6_n11) );
  MUX2_X1 pe_1_2_6_U69 ( .A(pe_1_2_6_int_q_reg_v[21]), .B(
        pe_1_2_6_int_q_reg_v[17]), .S(pe_1_2_6_n55), .Z(pe_1_2_6_n10) );
  MUX2_X1 pe_1_2_6_U68 ( .A(pe_1_2_6_int_q_reg_v[13]), .B(
        pe_1_2_6_int_q_reg_v[9]), .S(pe_1_2_6_n55), .Z(pe_1_2_6_n9) );
  MUX2_X1 pe_1_2_6_U67 ( .A(pe_1_2_6_int_q_reg_v[5]), .B(
        pe_1_2_6_int_q_reg_v[1]), .S(pe_1_2_6_n55), .Z(pe_1_2_6_n8) );
  MUX2_X1 pe_1_2_6_U66 ( .A(pe_1_2_6_n7), .B(pe_1_2_6_n4), .S(n47), .Z(
        int_data_y_2__6__0_) );
  MUX2_X1 pe_1_2_6_U65 ( .A(pe_1_2_6_n6), .B(pe_1_2_6_n5), .S(pe_1_2_6_n62), 
        .Z(pe_1_2_6_n7) );
  MUX2_X1 pe_1_2_6_U64 ( .A(pe_1_2_6_int_q_reg_v[20]), .B(
        pe_1_2_6_int_q_reg_v[16]), .S(pe_1_2_6_n55), .Z(pe_1_2_6_n6) );
  MUX2_X1 pe_1_2_6_U63 ( .A(pe_1_2_6_int_q_reg_v[12]), .B(
        pe_1_2_6_int_q_reg_v[8]), .S(pe_1_2_6_n55), .Z(pe_1_2_6_n5) );
  MUX2_X1 pe_1_2_6_U62 ( .A(pe_1_2_6_int_q_reg_v[4]), .B(
        pe_1_2_6_int_q_reg_v[0]), .S(pe_1_2_6_n55), .Z(pe_1_2_6_n4) );
  AOI222_X1 pe_1_2_6_U61 ( .A1(int_data_res_3__6__2_), .A2(pe_1_2_6_n64), .B1(
        pe_1_2_6_N80), .B2(pe_1_2_6_n27), .C1(pe_1_2_6_N72), .C2(pe_1_2_6_n28), 
        .ZN(pe_1_2_6_n33) );
  INV_X1 pe_1_2_6_U60 ( .A(pe_1_2_6_n33), .ZN(pe_1_2_6_n82) );
  AOI222_X1 pe_1_2_6_U59 ( .A1(int_data_res_3__6__6_), .A2(pe_1_2_6_n64), .B1(
        pe_1_2_6_N84), .B2(pe_1_2_6_n27), .C1(pe_1_2_6_N76), .C2(pe_1_2_6_n28), 
        .ZN(pe_1_2_6_n29) );
  INV_X1 pe_1_2_6_U58 ( .A(pe_1_2_6_n29), .ZN(pe_1_2_6_n78) );
  XNOR2_X1 pe_1_2_6_U57 ( .A(pe_1_2_6_n73), .B(int_data_res_2__6__0_), .ZN(
        pe_1_2_6_N70) );
  AOI222_X1 pe_1_2_6_U52 ( .A1(int_data_res_3__6__0_), .A2(pe_1_2_6_n64), .B1(
        pe_1_2_6_n1), .B2(pe_1_2_6_n27), .C1(pe_1_2_6_N70), .C2(pe_1_2_6_n28), 
        .ZN(pe_1_2_6_n35) );
  INV_X1 pe_1_2_6_U51 ( .A(pe_1_2_6_n35), .ZN(pe_1_2_6_n84) );
  AOI222_X1 pe_1_2_6_U50 ( .A1(int_data_res_3__6__1_), .A2(pe_1_2_6_n64), .B1(
        pe_1_2_6_N79), .B2(pe_1_2_6_n27), .C1(pe_1_2_6_N71), .C2(pe_1_2_6_n28), 
        .ZN(pe_1_2_6_n34) );
  INV_X1 pe_1_2_6_U49 ( .A(pe_1_2_6_n34), .ZN(pe_1_2_6_n83) );
  AOI222_X1 pe_1_2_6_U48 ( .A1(int_data_res_3__6__3_), .A2(pe_1_2_6_n64), .B1(
        pe_1_2_6_N81), .B2(pe_1_2_6_n27), .C1(pe_1_2_6_N73), .C2(pe_1_2_6_n28), 
        .ZN(pe_1_2_6_n32) );
  INV_X1 pe_1_2_6_U47 ( .A(pe_1_2_6_n32), .ZN(pe_1_2_6_n81) );
  AOI222_X1 pe_1_2_6_U46 ( .A1(int_data_res_3__6__4_), .A2(pe_1_2_6_n64), .B1(
        pe_1_2_6_N82), .B2(pe_1_2_6_n27), .C1(pe_1_2_6_N74), .C2(pe_1_2_6_n28), 
        .ZN(pe_1_2_6_n31) );
  INV_X1 pe_1_2_6_U45 ( .A(pe_1_2_6_n31), .ZN(pe_1_2_6_n80) );
  AOI222_X1 pe_1_2_6_U44 ( .A1(int_data_res_3__6__5_), .A2(pe_1_2_6_n64), .B1(
        pe_1_2_6_N83), .B2(pe_1_2_6_n27), .C1(pe_1_2_6_N75), .C2(pe_1_2_6_n28), 
        .ZN(pe_1_2_6_n30) );
  INV_X1 pe_1_2_6_U43 ( .A(pe_1_2_6_n30), .ZN(pe_1_2_6_n79) );
  NAND2_X1 pe_1_2_6_U42 ( .A1(pe_1_2_6_int_data_0_), .A2(pe_1_2_6_n3), .ZN(
        pe_1_2_6_sub_81_carry[1]) );
  INV_X1 pe_1_2_6_U41 ( .A(pe_1_2_6_int_data_1_), .ZN(pe_1_2_6_n74) );
  INV_X1 pe_1_2_6_U40 ( .A(pe_1_2_6_int_data_2_), .ZN(pe_1_2_6_n75) );
  AND2_X1 pe_1_2_6_U39 ( .A1(pe_1_2_6_int_data_0_), .A2(int_data_res_2__6__0_), 
        .ZN(pe_1_2_6_n2) );
  AOI222_X1 pe_1_2_6_U38 ( .A1(pe_1_2_6_n64), .A2(int_data_res_3__6__7_), .B1(
        pe_1_2_6_N85), .B2(pe_1_2_6_n27), .C1(pe_1_2_6_N77), .C2(pe_1_2_6_n28), 
        .ZN(pe_1_2_6_n26) );
  INV_X1 pe_1_2_6_U37 ( .A(pe_1_2_6_n26), .ZN(pe_1_2_6_n77) );
  NOR3_X1 pe_1_2_6_U36 ( .A1(pe_1_2_6_n59), .A2(pe_1_2_6_n65), .A3(int_ckg[41]), .ZN(pe_1_2_6_n36) );
  OR2_X1 pe_1_2_6_U35 ( .A1(pe_1_2_6_n36), .A2(pe_1_2_6_n64), .ZN(pe_1_2_6_N90) );
  INV_X1 pe_1_2_6_U34 ( .A(n38), .ZN(pe_1_2_6_n63) );
  AND2_X1 pe_1_2_6_U33 ( .A1(int_data_x_2__6__2_), .A2(pe_1_2_6_n58), .ZN(
        pe_1_2_6_int_data_2_) );
  AND2_X1 pe_1_2_6_U32 ( .A1(int_data_x_2__6__1_), .A2(pe_1_2_6_n58), .ZN(
        pe_1_2_6_int_data_1_) );
  AND2_X1 pe_1_2_6_U31 ( .A1(int_data_x_2__6__3_), .A2(pe_1_2_6_n58), .ZN(
        pe_1_2_6_int_data_3_) );
  BUF_X1 pe_1_2_6_U30 ( .A(n60), .Z(pe_1_2_6_n64) );
  INV_X1 pe_1_2_6_U29 ( .A(n32), .ZN(pe_1_2_6_n61) );
  AND2_X1 pe_1_2_6_U28 ( .A1(int_data_x_2__6__0_), .A2(pe_1_2_6_n58), .ZN(
        pe_1_2_6_int_data_0_) );
  NAND2_X1 pe_1_2_6_U27 ( .A1(pe_1_2_6_n44), .A2(pe_1_2_6_n61), .ZN(
        pe_1_2_6_n41) );
  AND3_X1 pe_1_2_6_U26 ( .A1(n74), .A2(pe_1_2_6_n63), .A3(n47), .ZN(
        pe_1_2_6_n44) );
  INV_X1 pe_1_2_6_U25 ( .A(pe_1_2_6_int_data_3_), .ZN(pe_1_2_6_n76) );
  NOR2_X1 pe_1_2_6_U24 ( .A1(pe_1_2_6_n70), .A2(n47), .ZN(pe_1_2_6_n43) );
  NOR2_X1 pe_1_2_6_U23 ( .A1(pe_1_2_6_n57), .A2(pe_1_2_6_n64), .ZN(
        pe_1_2_6_n28) );
  NOR2_X1 pe_1_2_6_U22 ( .A1(n18), .A2(pe_1_2_6_n64), .ZN(pe_1_2_6_n27) );
  INV_X1 pe_1_2_6_U21 ( .A(pe_1_2_6_int_data_0_), .ZN(pe_1_2_6_n73) );
  INV_X1 pe_1_2_6_U20 ( .A(pe_1_2_6_n41), .ZN(pe_1_2_6_n90) );
  INV_X1 pe_1_2_6_U19 ( .A(pe_1_2_6_n37), .ZN(pe_1_2_6_n88) );
  INV_X1 pe_1_2_6_U18 ( .A(pe_1_2_6_n38), .ZN(pe_1_2_6_n87) );
  INV_X1 pe_1_2_6_U17 ( .A(pe_1_2_6_n39), .ZN(pe_1_2_6_n86) );
  NOR2_X1 pe_1_2_6_U16 ( .A1(pe_1_2_6_n68), .A2(pe_1_2_6_n42), .ZN(
        pe_1_2_6_N59) );
  NOR2_X1 pe_1_2_6_U15 ( .A1(pe_1_2_6_n68), .A2(pe_1_2_6_n41), .ZN(
        pe_1_2_6_N60) );
  NOR2_X1 pe_1_2_6_U14 ( .A1(pe_1_2_6_n68), .A2(pe_1_2_6_n38), .ZN(
        pe_1_2_6_N63) );
  NOR2_X1 pe_1_2_6_U13 ( .A1(pe_1_2_6_n67), .A2(pe_1_2_6_n40), .ZN(
        pe_1_2_6_N61) );
  NOR2_X1 pe_1_2_6_U12 ( .A1(pe_1_2_6_n67), .A2(pe_1_2_6_n39), .ZN(
        pe_1_2_6_N62) );
  NOR2_X1 pe_1_2_6_U11 ( .A1(pe_1_2_6_n37), .A2(pe_1_2_6_n67), .ZN(
        pe_1_2_6_N64) );
  NAND2_X1 pe_1_2_6_U10 ( .A1(pe_1_2_6_n44), .A2(pe_1_2_6_n60), .ZN(
        pe_1_2_6_n42) );
  BUF_X1 pe_1_2_6_U9 ( .A(pe_1_2_6_n60), .Z(pe_1_2_6_n55) );
  INV_X1 pe_1_2_6_U8 ( .A(pe_1_2_6_n69), .ZN(pe_1_2_6_n65) );
  BUF_X1 pe_1_2_6_U7 ( .A(pe_1_2_6_n60), .Z(pe_1_2_6_n56) );
  INV_X1 pe_1_2_6_U6 ( .A(pe_1_2_6_n42), .ZN(pe_1_2_6_n89) );
  INV_X1 pe_1_2_6_U5 ( .A(pe_1_2_6_n40), .ZN(pe_1_2_6_n85) );
  INV_X2 pe_1_2_6_U4 ( .A(n82), .ZN(pe_1_2_6_n72) );
  XOR2_X1 pe_1_2_6_U3 ( .A(pe_1_2_6_int_data_0_), .B(int_data_res_2__6__0_), 
        .Z(pe_1_2_6_n1) );
  DFFR_X1 pe_1_2_6_int_q_acc_reg_0_ ( .D(pe_1_2_6_n84), .CK(pe_1_2_6_net5836), 
        .RN(pe_1_2_6_n72), .Q(int_data_res_2__6__0_), .QN(pe_1_2_6_n3) );
  DFFR_X1 pe_1_2_6_int_q_reg_v_reg_0__0_ ( .D(int_data_y_3__6__0_), .CK(
        pe_1_2_6_net5806), .RN(pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_v[20]) );
  DFFR_X1 pe_1_2_6_int_q_reg_v_reg_0__1_ ( .D(int_data_y_3__6__1_), .CK(
        pe_1_2_6_net5806), .RN(pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_v[21]) );
  DFFR_X1 pe_1_2_6_int_q_reg_v_reg_0__2_ ( .D(int_data_y_3__6__2_), .CK(
        pe_1_2_6_net5806), .RN(pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_v[22]) );
  DFFR_X1 pe_1_2_6_int_q_reg_v_reg_0__3_ ( .D(int_data_y_3__6__3_), .CK(
        pe_1_2_6_net5806), .RN(pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_v[23]) );
  DFFR_X1 pe_1_2_6_int_q_reg_v_reg_1__0_ ( .D(int_data_y_3__6__0_), .CK(
        pe_1_2_6_net5811), .RN(pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_v[16]) );
  DFFR_X1 pe_1_2_6_int_q_reg_v_reg_1__1_ ( .D(int_data_y_3__6__1_), .CK(
        pe_1_2_6_net5811), .RN(pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_v[17]) );
  DFFR_X1 pe_1_2_6_int_q_reg_v_reg_1__2_ ( .D(int_data_y_3__6__2_), .CK(
        pe_1_2_6_net5811), .RN(pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_v[18]) );
  DFFR_X1 pe_1_2_6_int_q_reg_v_reg_1__3_ ( .D(int_data_y_3__6__3_), .CK(
        pe_1_2_6_net5811), .RN(pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_v[19]) );
  DFFR_X1 pe_1_2_6_int_q_reg_v_reg_2__0_ ( .D(int_data_y_3__6__0_), .CK(
        pe_1_2_6_net5816), .RN(pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_v[12]) );
  DFFR_X1 pe_1_2_6_int_q_reg_v_reg_2__1_ ( .D(int_data_y_3__6__1_), .CK(
        pe_1_2_6_net5816), .RN(pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_v[13]) );
  DFFR_X1 pe_1_2_6_int_q_reg_v_reg_2__2_ ( .D(int_data_y_3__6__2_), .CK(
        pe_1_2_6_net5816), .RN(pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_v[14]) );
  DFFR_X1 pe_1_2_6_int_q_reg_v_reg_2__3_ ( .D(int_data_y_3__6__3_), .CK(
        pe_1_2_6_net5816), .RN(pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_v[15]) );
  DFFR_X1 pe_1_2_6_int_q_reg_v_reg_3__0_ ( .D(int_data_y_3__6__0_), .CK(
        pe_1_2_6_net5821), .RN(pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_v[8]) );
  DFFR_X1 pe_1_2_6_int_q_reg_v_reg_3__1_ ( .D(int_data_y_3__6__1_), .CK(
        pe_1_2_6_net5821), .RN(pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_v[9]) );
  DFFR_X1 pe_1_2_6_int_q_reg_v_reg_3__2_ ( .D(int_data_y_3__6__2_), .CK(
        pe_1_2_6_net5821), .RN(pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_v[10]) );
  DFFR_X1 pe_1_2_6_int_q_reg_v_reg_3__3_ ( .D(int_data_y_3__6__3_), .CK(
        pe_1_2_6_net5821), .RN(pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_v[11]) );
  DFFR_X1 pe_1_2_6_int_q_reg_v_reg_4__0_ ( .D(int_data_y_3__6__0_), .CK(
        pe_1_2_6_net5826), .RN(pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_v[4]) );
  DFFR_X1 pe_1_2_6_int_q_reg_v_reg_4__1_ ( .D(int_data_y_3__6__1_), .CK(
        pe_1_2_6_net5826), .RN(pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_v[5]) );
  DFFR_X1 pe_1_2_6_int_q_reg_v_reg_4__2_ ( .D(int_data_y_3__6__2_), .CK(
        pe_1_2_6_net5826), .RN(pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_v[6]) );
  DFFR_X1 pe_1_2_6_int_q_reg_v_reg_4__3_ ( .D(int_data_y_3__6__3_), .CK(
        pe_1_2_6_net5826), .RN(pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_v[7]) );
  DFFR_X1 pe_1_2_6_int_q_reg_v_reg_5__0_ ( .D(int_data_y_3__6__0_), .CK(
        pe_1_2_6_net5831), .RN(pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_v[0]) );
  DFFR_X1 pe_1_2_6_int_q_reg_v_reg_5__1_ ( .D(int_data_y_3__6__1_), .CK(
        pe_1_2_6_net5831), .RN(pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_v[1]) );
  DFFR_X1 pe_1_2_6_int_q_reg_v_reg_5__2_ ( .D(int_data_y_3__6__2_), .CK(
        pe_1_2_6_net5831), .RN(pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_v[2]) );
  DFFR_X1 pe_1_2_6_int_q_reg_v_reg_5__3_ ( .D(int_data_y_3__6__3_), .CK(
        pe_1_2_6_net5831), .RN(pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_2_6_int_q_reg_h_reg_0__0_ ( .D(int_data_x_2__7__0_), .SI(
        int_data_y_3__6__0_), .SE(pe_1_2_6_n65), .CK(pe_1_2_6_net5775), .RN(
        pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_2_6_int_q_reg_h_reg_0__1_ ( .D(int_data_x_2__7__1_), .SI(
        int_data_y_3__6__1_), .SE(pe_1_2_6_n65), .CK(pe_1_2_6_net5775), .RN(
        pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_2_6_int_q_reg_h_reg_0__2_ ( .D(int_data_x_2__7__2_), .SI(
        int_data_y_3__6__2_), .SE(pe_1_2_6_n65), .CK(pe_1_2_6_net5775), .RN(
        pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_2_6_int_q_reg_h_reg_0__3_ ( .D(int_data_x_2__7__3_), .SI(
        int_data_y_3__6__3_), .SE(pe_1_2_6_n65), .CK(pe_1_2_6_net5775), .RN(
        pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_2_6_int_q_reg_h_reg_1__0_ ( .D(int_data_x_2__7__0_), .SI(
        int_data_y_3__6__0_), .SE(pe_1_2_6_n65), .CK(pe_1_2_6_net5781), .RN(
        pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_2_6_int_q_reg_h_reg_1__1_ ( .D(int_data_x_2__7__1_), .SI(
        int_data_y_3__6__1_), .SE(pe_1_2_6_n65), .CK(pe_1_2_6_net5781), .RN(
        pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_2_6_int_q_reg_h_reg_1__2_ ( .D(int_data_x_2__7__2_), .SI(
        int_data_y_3__6__2_), .SE(pe_1_2_6_n65), .CK(pe_1_2_6_net5781), .RN(
        pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_2_6_int_q_reg_h_reg_1__3_ ( .D(int_data_x_2__7__3_), .SI(
        int_data_y_3__6__3_), .SE(pe_1_2_6_n65), .CK(pe_1_2_6_net5781), .RN(
        pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_2_6_int_q_reg_h_reg_2__0_ ( .D(int_data_x_2__7__0_), .SI(
        int_data_y_3__6__0_), .SE(pe_1_2_6_n65), .CK(pe_1_2_6_net5786), .RN(
        pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_2_6_int_q_reg_h_reg_2__1_ ( .D(int_data_x_2__7__1_), .SI(
        int_data_y_3__6__1_), .SE(pe_1_2_6_n65), .CK(pe_1_2_6_net5786), .RN(
        pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_2_6_int_q_reg_h_reg_2__2_ ( .D(int_data_x_2__7__2_), .SI(
        int_data_y_3__6__2_), .SE(pe_1_2_6_n65), .CK(pe_1_2_6_net5786), .RN(
        pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_2_6_int_q_reg_h_reg_2__3_ ( .D(int_data_x_2__7__3_), .SI(
        int_data_y_3__6__3_), .SE(pe_1_2_6_n65), .CK(pe_1_2_6_net5786), .RN(
        pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_2_6_int_q_reg_h_reg_3__0_ ( .D(int_data_x_2__7__0_), .SI(
        int_data_y_3__6__0_), .SE(pe_1_2_6_n65), .CK(pe_1_2_6_net5791), .RN(
        pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_2_6_int_q_reg_h_reg_3__1_ ( .D(int_data_x_2__7__1_), .SI(
        int_data_y_3__6__1_), .SE(pe_1_2_6_n65), .CK(pe_1_2_6_net5791), .RN(
        pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_2_6_int_q_reg_h_reg_3__2_ ( .D(int_data_x_2__7__2_), .SI(
        int_data_y_3__6__2_), .SE(pe_1_2_6_n65), .CK(pe_1_2_6_net5791), .RN(
        pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_2_6_int_q_reg_h_reg_3__3_ ( .D(int_data_x_2__7__3_), .SI(
        int_data_y_3__6__3_), .SE(pe_1_2_6_n65), .CK(pe_1_2_6_net5791), .RN(
        pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_2_6_int_q_reg_h_reg_4__0_ ( .D(int_data_x_2__7__0_), .SI(
        int_data_y_3__6__0_), .SE(pe_1_2_6_n66), .CK(pe_1_2_6_net5796), .RN(
        pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_2_6_int_q_reg_h_reg_4__1_ ( .D(int_data_x_2__7__1_), .SI(
        int_data_y_3__6__1_), .SE(pe_1_2_6_n66), .CK(pe_1_2_6_net5796), .RN(
        pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_2_6_int_q_reg_h_reg_4__2_ ( .D(int_data_x_2__7__2_), .SI(
        int_data_y_3__6__2_), .SE(pe_1_2_6_n66), .CK(pe_1_2_6_net5796), .RN(
        pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_2_6_int_q_reg_h_reg_4__3_ ( .D(int_data_x_2__7__3_), .SI(
        int_data_y_3__6__3_), .SE(pe_1_2_6_n66), .CK(pe_1_2_6_net5796), .RN(
        pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_2_6_int_q_reg_h_reg_5__0_ ( .D(int_data_x_2__7__0_), .SI(
        int_data_y_3__6__0_), .SE(pe_1_2_6_n66), .CK(pe_1_2_6_net5801), .RN(
        pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_2_6_int_q_reg_h_reg_5__1_ ( .D(int_data_x_2__7__1_), .SI(
        int_data_y_3__6__1_), .SE(pe_1_2_6_n66), .CK(pe_1_2_6_net5801), .RN(
        pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_2_6_int_q_reg_h_reg_5__2_ ( .D(int_data_x_2__7__2_), .SI(
        int_data_y_3__6__2_), .SE(pe_1_2_6_n66), .CK(pe_1_2_6_net5801), .RN(
        pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_2_6_int_q_reg_h_reg_5__3_ ( .D(int_data_x_2__7__3_), .SI(
        int_data_y_3__6__3_), .SE(pe_1_2_6_n66), .CK(pe_1_2_6_net5801), .RN(
        pe_1_2_6_n72), .Q(pe_1_2_6_int_q_reg_h[3]) );
  FA_X1 pe_1_2_6_sub_81_U2_7 ( .A(int_data_res_2__6__7_), .B(pe_1_2_6_n76), 
        .CI(pe_1_2_6_sub_81_carry[7]), .S(pe_1_2_6_N77) );
  FA_X1 pe_1_2_6_sub_81_U2_6 ( .A(int_data_res_2__6__6_), .B(pe_1_2_6_n76), 
        .CI(pe_1_2_6_sub_81_carry[6]), .CO(pe_1_2_6_sub_81_carry[7]), .S(
        pe_1_2_6_N76) );
  FA_X1 pe_1_2_6_sub_81_U2_5 ( .A(int_data_res_2__6__5_), .B(pe_1_2_6_n76), 
        .CI(pe_1_2_6_sub_81_carry[5]), .CO(pe_1_2_6_sub_81_carry[6]), .S(
        pe_1_2_6_N75) );
  FA_X1 pe_1_2_6_sub_81_U2_4 ( .A(int_data_res_2__6__4_), .B(pe_1_2_6_n76), 
        .CI(pe_1_2_6_sub_81_carry[4]), .CO(pe_1_2_6_sub_81_carry[5]), .S(
        pe_1_2_6_N74) );
  FA_X1 pe_1_2_6_sub_81_U2_3 ( .A(int_data_res_2__6__3_), .B(pe_1_2_6_n76), 
        .CI(pe_1_2_6_sub_81_carry[3]), .CO(pe_1_2_6_sub_81_carry[4]), .S(
        pe_1_2_6_N73) );
  FA_X1 pe_1_2_6_sub_81_U2_2 ( .A(int_data_res_2__6__2_), .B(pe_1_2_6_n75), 
        .CI(pe_1_2_6_sub_81_carry[2]), .CO(pe_1_2_6_sub_81_carry[3]), .S(
        pe_1_2_6_N72) );
  FA_X1 pe_1_2_6_sub_81_U2_1 ( .A(int_data_res_2__6__1_), .B(pe_1_2_6_n74), 
        .CI(pe_1_2_6_sub_81_carry[1]), .CO(pe_1_2_6_sub_81_carry[2]), .S(
        pe_1_2_6_N71) );
  FA_X1 pe_1_2_6_add_83_U1_7 ( .A(int_data_res_2__6__7_), .B(
        pe_1_2_6_int_data_3_), .CI(pe_1_2_6_add_83_carry[7]), .S(pe_1_2_6_N85)
         );
  FA_X1 pe_1_2_6_add_83_U1_6 ( .A(int_data_res_2__6__6_), .B(
        pe_1_2_6_int_data_3_), .CI(pe_1_2_6_add_83_carry[6]), .CO(
        pe_1_2_6_add_83_carry[7]), .S(pe_1_2_6_N84) );
  FA_X1 pe_1_2_6_add_83_U1_5 ( .A(int_data_res_2__6__5_), .B(
        pe_1_2_6_int_data_3_), .CI(pe_1_2_6_add_83_carry[5]), .CO(
        pe_1_2_6_add_83_carry[6]), .S(pe_1_2_6_N83) );
  FA_X1 pe_1_2_6_add_83_U1_4 ( .A(int_data_res_2__6__4_), .B(
        pe_1_2_6_int_data_3_), .CI(pe_1_2_6_add_83_carry[4]), .CO(
        pe_1_2_6_add_83_carry[5]), .S(pe_1_2_6_N82) );
  FA_X1 pe_1_2_6_add_83_U1_3 ( .A(int_data_res_2__6__3_), .B(
        pe_1_2_6_int_data_3_), .CI(pe_1_2_6_add_83_carry[3]), .CO(
        pe_1_2_6_add_83_carry[4]), .S(pe_1_2_6_N81) );
  FA_X1 pe_1_2_6_add_83_U1_2 ( .A(int_data_res_2__6__2_), .B(
        pe_1_2_6_int_data_2_), .CI(pe_1_2_6_add_83_carry[2]), .CO(
        pe_1_2_6_add_83_carry[3]), .S(pe_1_2_6_N80) );
  FA_X1 pe_1_2_6_add_83_U1_1 ( .A(int_data_res_2__6__1_), .B(
        pe_1_2_6_int_data_1_), .CI(pe_1_2_6_n2), .CO(pe_1_2_6_add_83_carry[2]), 
        .S(pe_1_2_6_N79) );
  NAND3_X1 pe_1_2_6_U56 ( .A1(pe_1_2_6_n60), .A2(pe_1_2_6_n43), .A3(
        pe_1_2_6_n62), .ZN(pe_1_2_6_n40) );
  NAND3_X1 pe_1_2_6_U55 ( .A1(pe_1_2_6_n43), .A2(pe_1_2_6_n61), .A3(
        pe_1_2_6_n62), .ZN(pe_1_2_6_n39) );
  NAND3_X1 pe_1_2_6_U54 ( .A1(pe_1_2_6_n43), .A2(pe_1_2_6_n63), .A3(
        pe_1_2_6_n60), .ZN(pe_1_2_6_n38) );
  NAND3_X1 pe_1_2_6_U53 ( .A1(pe_1_2_6_n61), .A2(pe_1_2_6_n63), .A3(
        pe_1_2_6_n43), .ZN(pe_1_2_6_n37) );
  DFFR_X1 pe_1_2_6_int_q_acc_reg_6_ ( .D(pe_1_2_6_n78), .CK(pe_1_2_6_net5836), 
        .RN(pe_1_2_6_n71), .Q(int_data_res_2__6__6_) );
  DFFR_X1 pe_1_2_6_int_q_acc_reg_5_ ( .D(pe_1_2_6_n79), .CK(pe_1_2_6_net5836), 
        .RN(pe_1_2_6_n71), .Q(int_data_res_2__6__5_) );
  DFFR_X1 pe_1_2_6_int_q_acc_reg_4_ ( .D(pe_1_2_6_n80), .CK(pe_1_2_6_net5836), 
        .RN(pe_1_2_6_n71), .Q(int_data_res_2__6__4_) );
  DFFR_X1 pe_1_2_6_int_q_acc_reg_3_ ( .D(pe_1_2_6_n81), .CK(pe_1_2_6_net5836), 
        .RN(pe_1_2_6_n71), .Q(int_data_res_2__6__3_) );
  DFFR_X1 pe_1_2_6_int_q_acc_reg_2_ ( .D(pe_1_2_6_n82), .CK(pe_1_2_6_net5836), 
        .RN(pe_1_2_6_n71), .Q(int_data_res_2__6__2_) );
  DFFR_X1 pe_1_2_6_int_q_acc_reg_1_ ( .D(pe_1_2_6_n83), .CK(pe_1_2_6_net5836), 
        .RN(pe_1_2_6_n71), .Q(int_data_res_2__6__1_) );
  DFFR_X1 pe_1_2_6_int_q_acc_reg_7_ ( .D(pe_1_2_6_n77), .CK(pe_1_2_6_net5836), 
        .RN(pe_1_2_6_n71), .Q(int_data_res_2__6__7_) );
  CLKGATETST_X1 pe_1_2_6_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_2_6_n88), .SE(1'b0), .GCK(pe_1_2_6_net5775) );
  CLKGATETST_X1 pe_1_2_6_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_2_6_n87), .SE(1'b0), .GCK(pe_1_2_6_net5781) );
  CLKGATETST_X1 pe_1_2_6_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_2_6_n86), .SE(1'b0), .GCK(pe_1_2_6_net5786) );
  CLKGATETST_X1 pe_1_2_6_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_2_6_n85), .SE(1'b0), .GCK(pe_1_2_6_net5791) );
  CLKGATETST_X1 pe_1_2_6_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_2_6_n90), .SE(1'b0), .GCK(pe_1_2_6_net5796) );
  CLKGATETST_X1 pe_1_2_6_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_2_6_n89), .SE(1'b0), .GCK(pe_1_2_6_net5801) );
  CLKGATETST_X1 pe_1_2_6_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_2_6_N64), .SE(1'b0), .GCK(pe_1_2_6_net5806) );
  CLKGATETST_X1 pe_1_2_6_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_2_6_N63), .SE(1'b0), .GCK(pe_1_2_6_net5811) );
  CLKGATETST_X1 pe_1_2_6_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_2_6_N62), .SE(1'b0), .GCK(pe_1_2_6_net5816) );
  CLKGATETST_X1 pe_1_2_6_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_2_6_N61), .SE(1'b0), .GCK(pe_1_2_6_net5821) );
  CLKGATETST_X1 pe_1_2_6_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_2_6_N60), .SE(1'b0), .GCK(pe_1_2_6_net5826) );
  CLKGATETST_X1 pe_1_2_6_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_2_6_N59), .SE(1'b0), .GCK(pe_1_2_6_net5831) );
  CLKGATETST_X1 pe_1_2_6_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_2_6_N90), .SE(1'b0), .GCK(pe_1_2_6_net5836) );
  CLKBUF_X1 pe_1_2_7_U112 ( .A(pe_1_2_7_n72), .Z(pe_1_2_7_n71) );
  INV_X1 pe_1_2_7_U111 ( .A(n74), .ZN(pe_1_2_7_n70) );
  INV_X1 pe_1_2_7_U110 ( .A(n66), .ZN(pe_1_2_7_n69) );
  INV_X1 pe_1_2_7_U109 ( .A(n66), .ZN(pe_1_2_7_n68) );
  INV_X1 pe_1_2_7_U108 ( .A(n66), .ZN(pe_1_2_7_n67) );
  INV_X1 pe_1_2_7_U107 ( .A(pe_1_2_7_n69), .ZN(pe_1_2_7_n66) );
  INV_X1 pe_1_2_7_U106 ( .A(pe_1_2_7_n63), .ZN(pe_1_2_7_n62) );
  INV_X1 pe_1_2_7_U105 ( .A(pe_1_2_7_n61), .ZN(pe_1_2_7_n60) );
  INV_X1 pe_1_2_7_U104 ( .A(n26), .ZN(pe_1_2_7_n59) );
  INV_X1 pe_1_2_7_U103 ( .A(pe_1_2_7_n59), .ZN(pe_1_2_7_n58) );
  INV_X1 pe_1_2_7_U102 ( .A(n18), .ZN(pe_1_2_7_n57) );
  MUX2_X1 pe_1_2_7_U101 ( .A(pe_1_2_7_n54), .B(pe_1_2_7_n51), .S(n47), .Z(
        int_data_x_2__7__3_) );
  MUX2_X1 pe_1_2_7_U100 ( .A(pe_1_2_7_n53), .B(pe_1_2_7_n52), .S(pe_1_2_7_n62), 
        .Z(pe_1_2_7_n54) );
  MUX2_X1 pe_1_2_7_U99 ( .A(pe_1_2_7_int_q_reg_h[23]), .B(
        pe_1_2_7_int_q_reg_h[19]), .S(pe_1_2_7_n56), .Z(pe_1_2_7_n53) );
  MUX2_X1 pe_1_2_7_U98 ( .A(pe_1_2_7_int_q_reg_h[15]), .B(
        pe_1_2_7_int_q_reg_h[11]), .S(pe_1_2_7_n56), .Z(pe_1_2_7_n52) );
  MUX2_X1 pe_1_2_7_U97 ( .A(pe_1_2_7_int_q_reg_h[7]), .B(
        pe_1_2_7_int_q_reg_h[3]), .S(pe_1_2_7_n56), .Z(pe_1_2_7_n51) );
  MUX2_X1 pe_1_2_7_U96 ( .A(pe_1_2_7_n50), .B(pe_1_2_7_n47), .S(n47), .Z(
        int_data_x_2__7__2_) );
  MUX2_X1 pe_1_2_7_U95 ( .A(pe_1_2_7_n49), .B(pe_1_2_7_n48), .S(pe_1_2_7_n62), 
        .Z(pe_1_2_7_n50) );
  MUX2_X1 pe_1_2_7_U94 ( .A(pe_1_2_7_int_q_reg_h[22]), .B(
        pe_1_2_7_int_q_reg_h[18]), .S(pe_1_2_7_n56), .Z(pe_1_2_7_n49) );
  MUX2_X1 pe_1_2_7_U93 ( .A(pe_1_2_7_int_q_reg_h[14]), .B(
        pe_1_2_7_int_q_reg_h[10]), .S(pe_1_2_7_n56), .Z(pe_1_2_7_n48) );
  MUX2_X1 pe_1_2_7_U92 ( .A(pe_1_2_7_int_q_reg_h[6]), .B(
        pe_1_2_7_int_q_reg_h[2]), .S(pe_1_2_7_n56), .Z(pe_1_2_7_n47) );
  MUX2_X1 pe_1_2_7_U91 ( .A(pe_1_2_7_n46), .B(pe_1_2_7_n24), .S(n47), .Z(
        int_data_x_2__7__1_) );
  MUX2_X1 pe_1_2_7_U90 ( .A(pe_1_2_7_n45), .B(pe_1_2_7_n25), .S(pe_1_2_7_n62), 
        .Z(pe_1_2_7_n46) );
  MUX2_X1 pe_1_2_7_U89 ( .A(pe_1_2_7_int_q_reg_h[21]), .B(
        pe_1_2_7_int_q_reg_h[17]), .S(pe_1_2_7_n56), .Z(pe_1_2_7_n45) );
  MUX2_X1 pe_1_2_7_U88 ( .A(pe_1_2_7_int_q_reg_h[13]), .B(
        pe_1_2_7_int_q_reg_h[9]), .S(pe_1_2_7_n56), .Z(pe_1_2_7_n25) );
  MUX2_X1 pe_1_2_7_U87 ( .A(pe_1_2_7_int_q_reg_h[5]), .B(
        pe_1_2_7_int_q_reg_h[1]), .S(pe_1_2_7_n56), .Z(pe_1_2_7_n24) );
  MUX2_X1 pe_1_2_7_U86 ( .A(pe_1_2_7_n23), .B(pe_1_2_7_n20), .S(n47), .Z(
        int_data_x_2__7__0_) );
  MUX2_X1 pe_1_2_7_U85 ( .A(pe_1_2_7_n22), .B(pe_1_2_7_n21), .S(pe_1_2_7_n62), 
        .Z(pe_1_2_7_n23) );
  MUX2_X1 pe_1_2_7_U84 ( .A(pe_1_2_7_int_q_reg_h[20]), .B(
        pe_1_2_7_int_q_reg_h[16]), .S(pe_1_2_7_n56), .Z(pe_1_2_7_n22) );
  MUX2_X1 pe_1_2_7_U83 ( .A(pe_1_2_7_int_q_reg_h[12]), .B(
        pe_1_2_7_int_q_reg_h[8]), .S(pe_1_2_7_n56), .Z(pe_1_2_7_n21) );
  MUX2_X1 pe_1_2_7_U82 ( .A(pe_1_2_7_int_q_reg_h[4]), .B(
        pe_1_2_7_int_q_reg_h[0]), .S(pe_1_2_7_n56), .Z(pe_1_2_7_n20) );
  MUX2_X1 pe_1_2_7_U81 ( .A(pe_1_2_7_n19), .B(pe_1_2_7_n16), .S(n47), .Z(
        int_data_y_2__7__3_) );
  MUX2_X1 pe_1_2_7_U80 ( .A(pe_1_2_7_n18), .B(pe_1_2_7_n17), .S(pe_1_2_7_n62), 
        .Z(pe_1_2_7_n19) );
  MUX2_X1 pe_1_2_7_U79 ( .A(pe_1_2_7_int_q_reg_v[23]), .B(
        pe_1_2_7_int_q_reg_v[19]), .S(pe_1_2_7_n55), .Z(pe_1_2_7_n18) );
  MUX2_X1 pe_1_2_7_U78 ( .A(pe_1_2_7_int_q_reg_v[15]), .B(
        pe_1_2_7_int_q_reg_v[11]), .S(pe_1_2_7_n55), .Z(pe_1_2_7_n17) );
  MUX2_X1 pe_1_2_7_U77 ( .A(pe_1_2_7_int_q_reg_v[7]), .B(
        pe_1_2_7_int_q_reg_v[3]), .S(pe_1_2_7_n55), .Z(pe_1_2_7_n16) );
  MUX2_X1 pe_1_2_7_U76 ( .A(pe_1_2_7_n15), .B(pe_1_2_7_n12), .S(n47), .Z(
        int_data_y_2__7__2_) );
  MUX2_X1 pe_1_2_7_U75 ( .A(pe_1_2_7_n14), .B(pe_1_2_7_n13), .S(pe_1_2_7_n62), 
        .Z(pe_1_2_7_n15) );
  MUX2_X1 pe_1_2_7_U74 ( .A(pe_1_2_7_int_q_reg_v[22]), .B(
        pe_1_2_7_int_q_reg_v[18]), .S(pe_1_2_7_n55), .Z(pe_1_2_7_n14) );
  MUX2_X1 pe_1_2_7_U73 ( .A(pe_1_2_7_int_q_reg_v[14]), .B(
        pe_1_2_7_int_q_reg_v[10]), .S(pe_1_2_7_n55), .Z(pe_1_2_7_n13) );
  MUX2_X1 pe_1_2_7_U72 ( .A(pe_1_2_7_int_q_reg_v[6]), .B(
        pe_1_2_7_int_q_reg_v[2]), .S(pe_1_2_7_n55), .Z(pe_1_2_7_n12) );
  MUX2_X1 pe_1_2_7_U71 ( .A(pe_1_2_7_n11), .B(pe_1_2_7_n8), .S(n47), .Z(
        int_data_y_2__7__1_) );
  MUX2_X1 pe_1_2_7_U70 ( .A(pe_1_2_7_n10), .B(pe_1_2_7_n9), .S(pe_1_2_7_n62), 
        .Z(pe_1_2_7_n11) );
  MUX2_X1 pe_1_2_7_U69 ( .A(pe_1_2_7_int_q_reg_v[21]), .B(
        pe_1_2_7_int_q_reg_v[17]), .S(pe_1_2_7_n55), .Z(pe_1_2_7_n10) );
  MUX2_X1 pe_1_2_7_U68 ( .A(pe_1_2_7_int_q_reg_v[13]), .B(
        pe_1_2_7_int_q_reg_v[9]), .S(pe_1_2_7_n55), .Z(pe_1_2_7_n9) );
  MUX2_X1 pe_1_2_7_U67 ( .A(pe_1_2_7_int_q_reg_v[5]), .B(
        pe_1_2_7_int_q_reg_v[1]), .S(pe_1_2_7_n55), .Z(pe_1_2_7_n8) );
  MUX2_X1 pe_1_2_7_U66 ( .A(pe_1_2_7_n7), .B(pe_1_2_7_n4), .S(n47), .Z(
        int_data_y_2__7__0_) );
  MUX2_X1 pe_1_2_7_U65 ( .A(pe_1_2_7_n6), .B(pe_1_2_7_n5), .S(pe_1_2_7_n62), 
        .Z(pe_1_2_7_n7) );
  MUX2_X1 pe_1_2_7_U64 ( .A(pe_1_2_7_int_q_reg_v[20]), .B(
        pe_1_2_7_int_q_reg_v[16]), .S(pe_1_2_7_n55), .Z(pe_1_2_7_n6) );
  MUX2_X1 pe_1_2_7_U63 ( .A(pe_1_2_7_int_q_reg_v[12]), .B(
        pe_1_2_7_int_q_reg_v[8]), .S(pe_1_2_7_n55), .Z(pe_1_2_7_n5) );
  MUX2_X1 pe_1_2_7_U62 ( .A(pe_1_2_7_int_q_reg_v[4]), .B(
        pe_1_2_7_int_q_reg_v[0]), .S(pe_1_2_7_n55), .Z(pe_1_2_7_n4) );
  AOI222_X1 pe_1_2_7_U61 ( .A1(int_data_res_3__7__2_), .A2(pe_1_2_7_n64), .B1(
        pe_1_2_7_N80), .B2(pe_1_2_7_n27), .C1(pe_1_2_7_N72), .C2(pe_1_2_7_n28), 
        .ZN(pe_1_2_7_n33) );
  INV_X1 pe_1_2_7_U60 ( .A(pe_1_2_7_n33), .ZN(pe_1_2_7_n82) );
  AOI222_X1 pe_1_2_7_U59 ( .A1(int_data_res_3__7__6_), .A2(pe_1_2_7_n64), .B1(
        pe_1_2_7_N84), .B2(pe_1_2_7_n27), .C1(pe_1_2_7_N76), .C2(pe_1_2_7_n28), 
        .ZN(pe_1_2_7_n29) );
  INV_X1 pe_1_2_7_U58 ( .A(pe_1_2_7_n29), .ZN(pe_1_2_7_n78) );
  XNOR2_X1 pe_1_2_7_U57 ( .A(pe_1_2_7_n73), .B(int_data_res_2__7__0_), .ZN(
        pe_1_2_7_N70) );
  AOI222_X1 pe_1_2_7_U52 ( .A1(int_data_res_3__7__0_), .A2(pe_1_2_7_n64), .B1(
        pe_1_2_7_n1), .B2(pe_1_2_7_n27), .C1(pe_1_2_7_N70), .C2(pe_1_2_7_n28), 
        .ZN(pe_1_2_7_n35) );
  INV_X1 pe_1_2_7_U51 ( .A(pe_1_2_7_n35), .ZN(pe_1_2_7_n84) );
  AOI222_X1 pe_1_2_7_U50 ( .A1(int_data_res_3__7__1_), .A2(pe_1_2_7_n64), .B1(
        pe_1_2_7_N79), .B2(pe_1_2_7_n27), .C1(pe_1_2_7_N71), .C2(pe_1_2_7_n28), 
        .ZN(pe_1_2_7_n34) );
  INV_X1 pe_1_2_7_U49 ( .A(pe_1_2_7_n34), .ZN(pe_1_2_7_n83) );
  AOI222_X1 pe_1_2_7_U48 ( .A1(int_data_res_3__7__3_), .A2(pe_1_2_7_n64), .B1(
        pe_1_2_7_N81), .B2(pe_1_2_7_n27), .C1(pe_1_2_7_N73), .C2(pe_1_2_7_n28), 
        .ZN(pe_1_2_7_n32) );
  INV_X1 pe_1_2_7_U47 ( .A(pe_1_2_7_n32), .ZN(pe_1_2_7_n81) );
  AOI222_X1 pe_1_2_7_U46 ( .A1(int_data_res_3__7__4_), .A2(pe_1_2_7_n64), .B1(
        pe_1_2_7_N82), .B2(pe_1_2_7_n27), .C1(pe_1_2_7_N74), .C2(pe_1_2_7_n28), 
        .ZN(pe_1_2_7_n31) );
  INV_X1 pe_1_2_7_U45 ( .A(pe_1_2_7_n31), .ZN(pe_1_2_7_n80) );
  AOI222_X1 pe_1_2_7_U44 ( .A1(int_data_res_3__7__5_), .A2(pe_1_2_7_n64), .B1(
        pe_1_2_7_N83), .B2(pe_1_2_7_n27), .C1(pe_1_2_7_N75), .C2(pe_1_2_7_n28), 
        .ZN(pe_1_2_7_n30) );
  INV_X1 pe_1_2_7_U43 ( .A(pe_1_2_7_n30), .ZN(pe_1_2_7_n79) );
  NAND2_X1 pe_1_2_7_U42 ( .A1(pe_1_2_7_int_data_0_), .A2(pe_1_2_7_n3), .ZN(
        pe_1_2_7_sub_81_carry[1]) );
  INV_X1 pe_1_2_7_U41 ( .A(pe_1_2_7_int_data_1_), .ZN(pe_1_2_7_n74) );
  INV_X1 pe_1_2_7_U40 ( .A(pe_1_2_7_int_data_2_), .ZN(pe_1_2_7_n75) );
  AND2_X1 pe_1_2_7_U39 ( .A1(pe_1_2_7_int_data_0_), .A2(int_data_res_2__7__0_), 
        .ZN(pe_1_2_7_n2) );
  AOI222_X1 pe_1_2_7_U38 ( .A1(pe_1_2_7_n64), .A2(int_data_res_3__7__7_), .B1(
        pe_1_2_7_N85), .B2(pe_1_2_7_n27), .C1(pe_1_2_7_N77), .C2(pe_1_2_7_n28), 
        .ZN(pe_1_2_7_n26) );
  INV_X1 pe_1_2_7_U37 ( .A(pe_1_2_7_n26), .ZN(pe_1_2_7_n77) );
  NOR3_X1 pe_1_2_7_U36 ( .A1(pe_1_2_7_n59), .A2(pe_1_2_7_n65), .A3(int_ckg[40]), .ZN(pe_1_2_7_n36) );
  OR2_X1 pe_1_2_7_U35 ( .A1(pe_1_2_7_n36), .A2(pe_1_2_7_n64), .ZN(pe_1_2_7_N90) );
  INV_X1 pe_1_2_7_U34 ( .A(n38), .ZN(pe_1_2_7_n63) );
  AND2_X1 pe_1_2_7_U33 ( .A1(int_data_x_2__7__2_), .A2(pe_1_2_7_n58), .ZN(
        pe_1_2_7_int_data_2_) );
  AND2_X1 pe_1_2_7_U32 ( .A1(int_data_x_2__7__1_), .A2(pe_1_2_7_n58), .ZN(
        pe_1_2_7_int_data_1_) );
  AND2_X1 pe_1_2_7_U31 ( .A1(int_data_x_2__7__3_), .A2(pe_1_2_7_n58), .ZN(
        pe_1_2_7_int_data_3_) );
  BUF_X1 pe_1_2_7_U30 ( .A(n60), .Z(pe_1_2_7_n64) );
  INV_X1 pe_1_2_7_U29 ( .A(n32), .ZN(pe_1_2_7_n61) );
  AND2_X1 pe_1_2_7_U28 ( .A1(int_data_x_2__7__0_), .A2(pe_1_2_7_n58), .ZN(
        pe_1_2_7_int_data_0_) );
  NAND2_X1 pe_1_2_7_U27 ( .A1(pe_1_2_7_n44), .A2(pe_1_2_7_n61), .ZN(
        pe_1_2_7_n41) );
  AND3_X1 pe_1_2_7_U26 ( .A1(n74), .A2(pe_1_2_7_n63), .A3(n47), .ZN(
        pe_1_2_7_n44) );
  INV_X1 pe_1_2_7_U25 ( .A(pe_1_2_7_int_data_3_), .ZN(pe_1_2_7_n76) );
  NOR2_X1 pe_1_2_7_U24 ( .A1(pe_1_2_7_n70), .A2(n47), .ZN(pe_1_2_7_n43) );
  NOR2_X1 pe_1_2_7_U23 ( .A1(pe_1_2_7_n57), .A2(pe_1_2_7_n64), .ZN(
        pe_1_2_7_n28) );
  NOR2_X1 pe_1_2_7_U22 ( .A1(n18), .A2(pe_1_2_7_n64), .ZN(pe_1_2_7_n27) );
  INV_X1 pe_1_2_7_U21 ( .A(pe_1_2_7_int_data_0_), .ZN(pe_1_2_7_n73) );
  INV_X1 pe_1_2_7_U20 ( .A(pe_1_2_7_n41), .ZN(pe_1_2_7_n90) );
  INV_X1 pe_1_2_7_U19 ( .A(pe_1_2_7_n37), .ZN(pe_1_2_7_n88) );
  INV_X1 pe_1_2_7_U18 ( .A(pe_1_2_7_n38), .ZN(pe_1_2_7_n87) );
  INV_X1 pe_1_2_7_U17 ( .A(pe_1_2_7_n39), .ZN(pe_1_2_7_n86) );
  NOR2_X1 pe_1_2_7_U16 ( .A1(pe_1_2_7_n68), .A2(pe_1_2_7_n42), .ZN(
        pe_1_2_7_N59) );
  NOR2_X1 pe_1_2_7_U15 ( .A1(pe_1_2_7_n68), .A2(pe_1_2_7_n41), .ZN(
        pe_1_2_7_N60) );
  NOR2_X1 pe_1_2_7_U14 ( .A1(pe_1_2_7_n68), .A2(pe_1_2_7_n38), .ZN(
        pe_1_2_7_N63) );
  NOR2_X1 pe_1_2_7_U13 ( .A1(pe_1_2_7_n67), .A2(pe_1_2_7_n40), .ZN(
        pe_1_2_7_N61) );
  NOR2_X1 pe_1_2_7_U12 ( .A1(pe_1_2_7_n67), .A2(pe_1_2_7_n39), .ZN(
        pe_1_2_7_N62) );
  NOR2_X1 pe_1_2_7_U11 ( .A1(pe_1_2_7_n37), .A2(pe_1_2_7_n67), .ZN(
        pe_1_2_7_N64) );
  NAND2_X1 pe_1_2_7_U10 ( .A1(pe_1_2_7_n44), .A2(pe_1_2_7_n60), .ZN(
        pe_1_2_7_n42) );
  BUF_X1 pe_1_2_7_U9 ( .A(pe_1_2_7_n60), .Z(pe_1_2_7_n55) );
  INV_X1 pe_1_2_7_U8 ( .A(pe_1_2_7_n69), .ZN(pe_1_2_7_n65) );
  BUF_X1 pe_1_2_7_U7 ( .A(pe_1_2_7_n60), .Z(pe_1_2_7_n56) );
  INV_X1 pe_1_2_7_U6 ( .A(pe_1_2_7_n42), .ZN(pe_1_2_7_n89) );
  INV_X1 pe_1_2_7_U5 ( .A(pe_1_2_7_n40), .ZN(pe_1_2_7_n85) );
  INV_X2 pe_1_2_7_U4 ( .A(n82), .ZN(pe_1_2_7_n72) );
  XOR2_X1 pe_1_2_7_U3 ( .A(pe_1_2_7_int_data_0_), .B(int_data_res_2__7__0_), 
        .Z(pe_1_2_7_n1) );
  DFFR_X1 pe_1_2_7_int_q_acc_reg_0_ ( .D(pe_1_2_7_n84), .CK(pe_1_2_7_net5758), 
        .RN(pe_1_2_7_n72), .Q(int_data_res_2__7__0_), .QN(pe_1_2_7_n3) );
  DFFR_X1 pe_1_2_7_int_q_reg_v_reg_0__0_ ( .D(int_data_y_3__7__0_), .CK(
        pe_1_2_7_net5728), .RN(pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_v[20]) );
  DFFR_X1 pe_1_2_7_int_q_reg_v_reg_0__1_ ( .D(int_data_y_3__7__1_), .CK(
        pe_1_2_7_net5728), .RN(pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_v[21]) );
  DFFR_X1 pe_1_2_7_int_q_reg_v_reg_0__2_ ( .D(int_data_y_3__7__2_), .CK(
        pe_1_2_7_net5728), .RN(pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_v[22]) );
  DFFR_X1 pe_1_2_7_int_q_reg_v_reg_0__3_ ( .D(int_data_y_3__7__3_), .CK(
        pe_1_2_7_net5728), .RN(pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_v[23]) );
  DFFR_X1 pe_1_2_7_int_q_reg_v_reg_1__0_ ( .D(int_data_y_3__7__0_), .CK(
        pe_1_2_7_net5733), .RN(pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_v[16]) );
  DFFR_X1 pe_1_2_7_int_q_reg_v_reg_1__1_ ( .D(int_data_y_3__7__1_), .CK(
        pe_1_2_7_net5733), .RN(pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_v[17]) );
  DFFR_X1 pe_1_2_7_int_q_reg_v_reg_1__2_ ( .D(int_data_y_3__7__2_), .CK(
        pe_1_2_7_net5733), .RN(pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_v[18]) );
  DFFR_X1 pe_1_2_7_int_q_reg_v_reg_1__3_ ( .D(int_data_y_3__7__3_), .CK(
        pe_1_2_7_net5733), .RN(pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_v[19]) );
  DFFR_X1 pe_1_2_7_int_q_reg_v_reg_2__0_ ( .D(int_data_y_3__7__0_), .CK(
        pe_1_2_7_net5738), .RN(pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_v[12]) );
  DFFR_X1 pe_1_2_7_int_q_reg_v_reg_2__1_ ( .D(int_data_y_3__7__1_), .CK(
        pe_1_2_7_net5738), .RN(pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_v[13]) );
  DFFR_X1 pe_1_2_7_int_q_reg_v_reg_2__2_ ( .D(int_data_y_3__7__2_), .CK(
        pe_1_2_7_net5738), .RN(pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_v[14]) );
  DFFR_X1 pe_1_2_7_int_q_reg_v_reg_2__3_ ( .D(int_data_y_3__7__3_), .CK(
        pe_1_2_7_net5738), .RN(pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_v[15]) );
  DFFR_X1 pe_1_2_7_int_q_reg_v_reg_3__0_ ( .D(int_data_y_3__7__0_), .CK(
        pe_1_2_7_net5743), .RN(pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_v[8]) );
  DFFR_X1 pe_1_2_7_int_q_reg_v_reg_3__1_ ( .D(int_data_y_3__7__1_), .CK(
        pe_1_2_7_net5743), .RN(pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_v[9]) );
  DFFR_X1 pe_1_2_7_int_q_reg_v_reg_3__2_ ( .D(int_data_y_3__7__2_), .CK(
        pe_1_2_7_net5743), .RN(pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_v[10]) );
  DFFR_X1 pe_1_2_7_int_q_reg_v_reg_3__3_ ( .D(int_data_y_3__7__3_), .CK(
        pe_1_2_7_net5743), .RN(pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_v[11]) );
  DFFR_X1 pe_1_2_7_int_q_reg_v_reg_4__0_ ( .D(int_data_y_3__7__0_), .CK(
        pe_1_2_7_net5748), .RN(pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_v[4]) );
  DFFR_X1 pe_1_2_7_int_q_reg_v_reg_4__1_ ( .D(int_data_y_3__7__1_), .CK(
        pe_1_2_7_net5748), .RN(pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_v[5]) );
  DFFR_X1 pe_1_2_7_int_q_reg_v_reg_4__2_ ( .D(int_data_y_3__7__2_), .CK(
        pe_1_2_7_net5748), .RN(pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_v[6]) );
  DFFR_X1 pe_1_2_7_int_q_reg_v_reg_4__3_ ( .D(int_data_y_3__7__3_), .CK(
        pe_1_2_7_net5748), .RN(pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_v[7]) );
  DFFR_X1 pe_1_2_7_int_q_reg_v_reg_5__0_ ( .D(int_data_y_3__7__0_), .CK(
        pe_1_2_7_net5753), .RN(pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_v[0]) );
  DFFR_X1 pe_1_2_7_int_q_reg_v_reg_5__1_ ( .D(int_data_y_3__7__1_), .CK(
        pe_1_2_7_net5753), .RN(pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_v[1]) );
  DFFR_X1 pe_1_2_7_int_q_reg_v_reg_5__2_ ( .D(int_data_y_3__7__2_), .CK(
        pe_1_2_7_net5753), .RN(pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_v[2]) );
  DFFR_X1 pe_1_2_7_int_q_reg_v_reg_5__3_ ( .D(int_data_y_3__7__3_), .CK(
        pe_1_2_7_net5753), .RN(pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_2_7_int_q_reg_h_reg_0__0_ ( .D(i_data_conv_h[20]), .SI(
        int_data_y_3__7__0_), .SE(pe_1_2_7_n65), .CK(pe_1_2_7_net5697), .RN(
        pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_2_7_int_q_reg_h_reg_0__1_ ( .D(i_data_conv_h[21]), .SI(
        int_data_y_3__7__1_), .SE(pe_1_2_7_n65), .CK(pe_1_2_7_net5697), .RN(
        pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_2_7_int_q_reg_h_reg_0__2_ ( .D(i_data_conv_h[22]), .SI(
        int_data_y_3__7__2_), .SE(pe_1_2_7_n65), .CK(pe_1_2_7_net5697), .RN(
        pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_2_7_int_q_reg_h_reg_0__3_ ( .D(i_data_conv_h[23]), .SI(
        int_data_y_3__7__3_), .SE(pe_1_2_7_n65), .CK(pe_1_2_7_net5697), .RN(
        pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_2_7_int_q_reg_h_reg_1__0_ ( .D(i_data_conv_h[20]), .SI(
        int_data_y_3__7__0_), .SE(pe_1_2_7_n65), .CK(pe_1_2_7_net5703), .RN(
        pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_2_7_int_q_reg_h_reg_1__1_ ( .D(i_data_conv_h[21]), .SI(
        int_data_y_3__7__1_), .SE(pe_1_2_7_n65), .CK(pe_1_2_7_net5703), .RN(
        pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_2_7_int_q_reg_h_reg_1__2_ ( .D(i_data_conv_h[22]), .SI(
        int_data_y_3__7__2_), .SE(pe_1_2_7_n65), .CK(pe_1_2_7_net5703), .RN(
        pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_2_7_int_q_reg_h_reg_1__3_ ( .D(i_data_conv_h[23]), .SI(
        int_data_y_3__7__3_), .SE(pe_1_2_7_n65), .CK(pe_1_2_7_net5703), .RN(
        pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_2_7_int_q_reg_h_reg_2__0_ ( .D(i_data_conv_h[20]), .SI(
        int_data_y_3__7__0_), .SE(pe_1_2_7_n65), .CK(pe_1_2_7_net5708), .RN(
        pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_2_7_int_q_reg_h_reg_2__1_ ( .D(i_data_conv_h[21]), .SI(
        int_data_y_3__7__1_), .SE(pe_1_2_7_n65), .CK(pe_1_2_7_net5708), .RN(
        pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_2_7_int_q_reg_h_reg_2__2_ ( .D(i_data_conv_h[22]), .SI(
        int_data_y_3__7__2_), .SE(pe_1_2_7_n65), .CK(pe_1_2_7_net5708), .RN(
        pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_2_7_int_q_reg_h_reg_2__3_ ( .D(i_data_conv_h[23]), .SI(
        int_data_y_3__7__3_), .SE(pe_1_2_7_n65), .CK(pe_1_2_7_net5708), .RN(
        pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_2_7_int_q_reg_h_reg_3__0_ ( .D(i_data_conv_h[20]), .SI(
        int_data_y_3__7__0_), .SE(pe_1_2_7_n65), .CK(pe_1_2_7_net5713), .RN(
        pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_2_7_int_q_reg_h_reg_3__1_ ( .D(i_data_conv_h[21]), .SI(
        int_data_y_3__7__1_), .SE(pe_1_2_7_n65), .CK(pe_1_2_7_net5713), .RN(
        pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_2_7_int_q_reg_h_reg_3__2_ ( .D(i_data_conv_h[22]), .SI(
        int_data_y_3__7__2_), .SE(pe_1_2_7_n65), .CK(pe_1_2_7_net5713), .RN(
        pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_2_7_int_q_reg_h_reg_3__3_ ( .D(i_data_conv_h[23]), .SI(
        int_data_y_3__7__3_), .SE(pe_1_2_7_n65), .CK(pe_1_2_7_net5713), .RN(
        pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_2_7_int_q_reg_h_reg_4__0_ ( .D(i_data_conv_h[20]), .SI(
        int_data_y_3__7__0_), .SE(pe_1_2_7_n66), .CK(pe_1_2_7_net5718), .RN(
        pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_2_7_int_q_reg_h_reg_4__1_ ( .D(i_data_conv_h[21]), .SI(
        int_data_y_3__7__1_), .SE(pe_1_2_7_n66), .CK(pe_1_2_7_net5718), .RN(
        pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_2_7_int_q_reg_h_reg_4__2_ ( .D(i_data_conv_h[22]), .SI(
        int_data_y_3__7__2_), .SE(pe_1_2_7_n66), .CK(pe_1_2_7_net5718), .RN(
        pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_2_7_int_q_reg_h_reg_4__3_ ( .D(i_data_conv_h[23]), .SI(
        int_data_y_3__7__3_), .SE(pe_1_2_7_n66), .CK(pe_1_2_7_net5718), .RN(
        pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_2_7_int_q_reg_h_reg_5__0_ ( .D(i_data_conv_h[20]), .SI(
        int_data_y_3__7__0_), .SE(pe_1_2_7_n66), .CK(pe_1_2_7_net5723), .RN(
        pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_2_7_int_q_reg_h_reg_5__1_ ( .D(i_data_conv_h[21]), .SI(
        int_data_y_3__7__1_), .SE(pe_1_2_7_n66), .CK(pe_1_2_7_net5723), .RN(
        pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_2_7_int_q_reg_h_reg_5__2_ ( .D(i_data_conv_h[22]), .SI(
        int_data_y_3__7__2_), .SE(pe_1_2_7_n66), .CK(pe_1_2_7_net5723), .RN(
        pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_2_7_int_q_reg_h_reg_5__3_ ( .D(i_data_conv_h[23]), .SI(
        int_data_y_3__7__3_), .SE(pe_1_2_7_n66), .CK(pe_1_2_7_net5723), .RN(
        pe_1_2_7_n72), .Q(pe_1_2_7_int_q_reg_h[3]) );
  FA_X1 pe_1_2_7_sub_81_U2_7 ( .A(int_data_res_2__7__7_), .B(pe_1_2_7_n76), 
        .CI(pe_1_2_7_sub_81_carry[7]), .S(pe_1_2_7_N77) );
  FA_X1 pe_1_2_7_sub_81_U2_6 ( .A(int_data_res_2__7__6_), .B(pe_1_2_7_n76), 
        .CI(pe_1_2_7_sub_81_carry[6]), .CO(pe_1_2_7_sub_81_carry[7]), .S(
        pe_1_2_7_N76) );
  FA_X1 pe_1_2_7_sub_81_U2_5 ( .A(int_data_res_2__7__5_), .B(pe_1_2_7_n76), 
        .CI(pe_1_2_7_sub_81_carry[5]), .CO(pe_1_2_7_sub_81_carry[6]), .S(
        pe_1_2_7_N75) );
  FA_X1 pe_1_2_7_sub_81_U2_4 ( .A(int_data_res_2__7__4_), .B(pe_1_2_7_n76), 
        .CI(pe_1_2_7_sub_81_carry[4]), .CO(pe_1_2_7_sub_81_carry[5]), .S(
        pe_1_2_7_N74) );
  FA_X1 pe_1_2_7_sub_81_U2_3 ( .A(int_data_res_2__7__3_), .B(pe_1_2_7_n76), 
        .CI(pe_1_2_7_sub_81_carry[3]), .CO(pe_1_2_7_sub_81_carry[4]), .S(
        pe_1_2_7_N73) );
  FA_X1 pe_1_2_7_sub_81_U2_2 ( .A(int_data_res_2__7__2_), .B(pe_1_2_7_n75), 
        .CI(pe_1_2_7_sub_81_carry[2]), .CO(pe_1_2_7_sub_81_carry[3]), .S(
        pe_1_2_7_N72) );
  FA_X1 pe_1_2_7_sub_81_U2_1 ( .A(int_data_res_2__7__1_), .B(pe_1_2_7_n74), 
        .CI(pe_1_2_7_sub_81_carry[1]), .CO(pe_1_2_7_sub_81_carry[2]), .S(
        pe_1_2_7_N71) );
  FA_X1 pe_1_2_7_add_83_U1_7 ( .A(int_data_res_2__7__7_), .B(
        pe_1_2_7_int_data_3_), .CI(pe_1_2_7_add_83_carry[7]), .S(pe_1_2_7_N85)
         );
  FA_X1 pe_1_2_7_add_83_U1_6 ( .A(int_data_res_2__7__6_), .B(
        pe_1_2_7_int_data_3_), .CI(pe_1_2_7_add_83_carry[6]), .CO(
        pe_1_2_7_add_83_carry[7]), .S(pe_1_2_7_N84) );
  FA_X1 pe_1_2_7_add_83_U1_5 ( .A(int_data_res_2__7__5_), .B(
        pe_1_2_7_int_data_3_), .CI(pe_1_2_7_add_83_carry[5]), .CO(
        pe_1_2_7_add_83_carry[6]), .S(pe_1_2_7_N83) );
  FA_X1 pe_1_2_7_add_83_U1_4 ( .A(int_data_res_2__7__4_), .B(
        pe_1_2_7_int_data_3_), .CI(pe_1_2_7_add_83_carry[4]), .CO(
        pe_1_2_7_add_83_carry[5]), .S(pe_1_2_7_N82) );
  FA_X1 pe_1_2_7_add_83_U1_3 ( .A(int_data_res_2__7__3_), .B(
        pe_1_2_7_int_data_3_), .CI(pe_1_2_7_add_83_carry[3]), .CO(
        pe_1_2_7_add_83_carry[4]), .S(pe_1_2_7_N81) );
  FA_X1 pe_1_2_7_add_83_U1_2 ( .A(int_data_res_2__7__2_), .B(
        pe_1_2_7_int_data_2_), .CI(pe_1_2_7_add_83_carry[2]), .CO(
        pe_1_2_7_add_83_carry[3]), .S(pe_1_2_7_N80) );
  FA_X1 pe_1_2_7_add_83_U1_1 ( .A(int_data_res_2__7__1_), .B(
        pe_1_2_7_int_data_1_), .CI(pe_1_2_7_n2), .CO(pe_1_2_7_add_83_carry[2]), 
        .S(pe_1_2_7_N79) );
  NAND3_X1 pe_1_2_7_U56 ( .A1(pe_1_2_7_n60), .A2(pe_1_2_7_n43), .A3(
        pe_1_2_7_n62), .ZN(pe_1_2_7_n40) );
  NAND3_X1 pe_1_2_7_U55 ( .A1(pe_1_2_7_n43), .A2(pe_1_2_7_n61), .A3(
        pe_1_2_7_n62), .ZN(pe_1_2_7_n39) );
  NAND3_X1 pe_1_2_7_U54 ( .A1(pe_1_2_7_n43), .A2(pe_1_2_7_n63), .A3(
        pe_1_2_7_n60), .ZN(pe_1_2_7_n38) );
  NAND3_X1 pe_1_2_7_U53 ( .A1(pe_1_2_7_n61), .A2(pe_1_2_7_n63), .A3(
        pe_1_2_7_n43), .ZN(pe_1_2_7_n37) );
  DFFR_X1 pe_1_2_7_int_q_acc_reg_6_ ( .D(pe_1_2_7_n78), .CK(pe_1_2_7_net5758), 
        .RN(pe_1_2_7_n71), .Q(int_data_res_2__7__6_) );
  DFFR_X1 pe_1_2_7_int_q_acc_reg_5_ ( .D(pe_1_2_7_n79), .CK(pe_1_2_7_net5758), 
        .RN(pe_1_2_7_n71), .Q(int_data_res_2__7__5_) );
  DFFR_X1 pe_1_2_7_int_q_acc_reg_4_ ( .D(pe_1_2_7_n80), .CK(pe_1_2_7_net5758), 
        .RN(pe_1_2_7_n71), .Q(int_data_res_2__7__4_) );
  DFFR_X1 pe_1_2_7_int_q_acc_reg_3_ ( .D(pe_1_2_7_n81), .CK(pe_1_2_7_net5758), 
        .RN(pe_1_2_7_n71), .Q(int_data_res_2__7__3_) );
  DFFR_X1 pe_1_2_7_int_q_acc_reg_2_ ( .D(pe_1_2_7_n82), .CK(pe_1_2_7_net5758), 
        .RN(pe_1_2_7_n71), .Q(int_data_res_2__7__2_) );
  DFFR_X1 pe_1_2_7_int_q_acc_reg_1_ ( .D(pe_1_2_7_n83), .CK(pe_1_2_7_net5758), 
        .RN(pe_1_2_7_n71), .Q(int_data_res_2__7__1_) );
  DFFR_X1 pe_1_2_7_int_q_acc_reg_7_ ( .D(pe_1_2_7_n77), .CK(pe_1_2_7_net5758), 
        .RN(pe_1_2_7_n71), .Q(int_data_res_2__7__7_) );
  CLKGATETST_X1 pe_1_2_7_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_2_7_n88), .SE(1'b0), .GCK(pe_1_2_7_net5697) );
  CLKGATETST_X1 pe_1_2_7_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_2_7_n87), .SE(1'b0), .GCK(pe_1_2_7_net5703) );
  CLKGATETST_X1 pe_1_2_7_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_2_7_n86), .SE(1'b0), .GCK(pe_1_2_7_net5708) );
  CLKGATETST_X1 pe_1_2_7_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_2_7_n85), .SE(1'b0), .GCK(pe_1_2_7_net5713) );
  CLKGATETST_X1 pe_1_2_7_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_2_7_n90), .SE(1'b0), .GCK(pe_1_2_7_net5718) );
  CLKGATETST_X1 pe_1_2_7_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_2_7_n89), .SE(1'b0), .GCK(pe_1_2_7_net5723) );
  CLKGATETST_X1 pe_1_2_7_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_2_7_N64), .SE(1'b0), .GCK(pe_1_2_7_net5728) );
  CLKGATETST_X1 pe_1_2_7_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_2_7_N63), .SE(1'b0), .GCK(pe_1_2_7_net5733) );
  CLKGATETST_X1 pe_1_2_7_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_2_7_N62), .SE(1'b0), .GCK(pe_1_2_7_net5738) );
  CLKGATETST_X1 pe_1_2_7_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_2_7_N61), .SE(1'b0), .GCK(pe_1_2_7_net5743) );
  CLKGATETST_X1 pe_1_2_7_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_2_7_N60), .SE(1'b0), .GCK(pe_1_2_7_net5748) );
  CLKGATETST_X1 pe_1_2_7_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_2_7_N59), .SE(1'b0), .GCK(pe_1_2_7_net5753) );
  CLKGATETST_X1 pe_1_2_7_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_2_7_N90), .SE(1'b0), .GCK(pe_1_2_7_net5758) );
  CLKBUF_X1 pe_1_3_0_U109 ( .A(pe_1_3_0_n69), .Z(pe_1_3_0_n68) );
  INV_X1 pe_1_3_0_U108 ( .A(n75), .ZN(pe_1_3_0_n67) );
  INV_X1 pe_1_3_0_U107 ( .A(n67), .ZN(pe_1_3_0_n66) );
  INV_X1 pe_1_3_0_U106 ( .A(n67), .ZN(pe_1_3_0_n65) );
  INV_X1 pe_1_3_0_U105 ( .A(pe_1_3_0_n66), .ZN(pe_1_3_0_n64) );
  INV_X1 pe_1_3_0_U104 ( .A(pe_1_3_0_n61), .ZN(pe_1_3_0_n60) );
  INV_X1 pe_1_3_0_U103 ( .A(n27), .ZN(pe_1_3_0_n58) );
  INV_X1 pe_1_3_0_U102 ( .A(n19), .ZN(pe_1_3_0_n57) );
  MUX2_X1 pe_1_3_0_U101 ( .A(pe_1_3_0_n54), .B(pe_1_3_0_n51), .S(n47), .Z(
        pe_1_3_0_o_data_h_3_) );
  MUX2_X1 pe_1_3_0_U100 ( .A(pe_1_3_0_n53), .B(pe_1_3_0_n52), .S(pe_1_3_0_n60), 
        .Z(pe_1_3_0_n54) );
  MUX2_X1 pe_1_3_0_U99 ( .A(pe_1_3_0_int_q_reg_h[23]), .B(
        pe_1_3_0_int_q_reg_h[19]), .S(pe_1_3_0_n56), .Z(pe_1_3_0_n53) );
  MUX2_X1 pe_1_3_0_U98 ( .A(pe_1_3_0_int_q_reg_h[15]), .B(
        pe_1_3_0_int_q_reg_h[11]), .S(pe_1_3_0_n56), .Z(pe_1_3_0_n52) );
  MUX2_X1 pe_1_3_0_U97 ( .A(pe_1_3_0_int_q_reg_h[7]), .B(
        pe_1_3_0_int_q_reg_h[3]), .S(pe_1_3_0_n56), .Z(pe_1_3_0_n51) );
  MUX2_X1 pe_1_3_0_U96 ( .A(pe_1_3_0_n50), .B(pe_1_3_0_n47), .S(n47), .Z(
        pe_1_3_0_o_data_h_2_) );
  MUX2_X1 pe_1_3_0_U95 ( .A(pe_1_3_0_n49), .B(pe_1_3_0_n48), .S(pe_1_3_0_n60), 
        .Z(pe_1_3_0_n50) );
  MUX2_X1 pe_1_3_0_U94 ( .A(pe_1_3_0_int_q_reg_h[22]), .B(
        pe_1_3_0_int_q_reg_h[18]), .S(pe_1_3_0_n56), .Z(pe_1_3_0_n49) );
  MUX2_X1 pe_1_3_0_U93 ( .A(pe_1_3_0_int_q_reg_h[14]), .B(
        pe_1_3_0_int_q_reg_h[10]), .S(pe_1_3_0_n56), .Z(pe_1_3_0_n48) );
  MUX2_X1 pe_1_3_0_U92 ( .A(pe_1_3_0_int_q_reg_h[6]), .B(
        pe_1_3_0_int_q_reg_h[2]), .S(pe_1_3_0_n56), .Z(pe_1_3_0_n47) );
  MUX2_X1 pe_1_3_0_U91 ( .A(pe_1_3_0_n46), .B(pe_1_3_0_n24), .S(n47), .Z(
        pe_1_3_0_o_data_h_1_) );
  MUX2_X1 pe_1_3_0_U90 ( .A(pe_1_3_0_n45), .B(pe_1_3_0_n25), .S(pe_1_3_0_n60), 
        .Z(pe_1_3_0_n46) );
  MUX2_X1 pe_1_3_0_U89 ( .A(pe_1_3_0_int_q_reg_h[21]), .B(
        pe_1_3_0_int_q_reg_h[17]), .S(pe_1_3_0_n56), .Z(pe_1_3_0_n45) );
  MUX2_X1 pe_1_3_0_U88 ( .A(pe_1_3_0_int_q_reg_h[13]), .B(
        pe_1_3_0_int_q_reg_h[9]), .S(pe_1_3_0_n56), .Z(pe_1_3_0_n25) );
  MUX2_X1 pe_1_3_0_U87 ( .A(pe_1_3_0_int_q_reg_h[5]), .B(
        pe_1_3_0_int_q_reg_h[1]), .S(pe_1_3_0_n56), .Z(pe_1_3_0_n24) );
  MUX2_X1 pe_1_3_0_U86 ( .A(pe_1_3_0_n23), .B(pe_1_3_0_n20), .S(n47), .Z(
        pe_1_3_0_o_data_h_0_) );
  MUX2_X1 pe_1_3_0_U85 ( .A(pe_1_3_0_n22), .B(pe_1_3_0_n21), .S(pe_1_3_0_n60), 
        .Z(pe_1_3_0_n23) );
  MUX2_X1 pe_1_3_0_U84 ( .A(pe_1_3_0_int_q_reg_h[20]), .B(
        pe_1_3_0_int_q_reg_h[16]), .S(pe_1_3_0_n56), .Z(pe_1_3_0_n22) );
  MUX2_X1 pe_1_3_0_U83 ( .A(pe_1_3_0_int_q_reg_h[12]), .B(
        pe_1_3_0_int_q_reg_h[8]), .S(pe_1_3_0_n56), .Z(pe_1_3_0_n21) );
  MUX2_X1 pe_1_3_0_U82 ( .A(pe_1_3_0_int_q_reg_h[4]), .B(
        pe_1_3_0_int_q_reg_h[0]), .S(pe_1_3_0_n56), .Z(pe_1_3_0_n20) );
  MUX2_X1 pe_1_3_0_U81 ( .A(pe_1_3_0_n19), .B(pe_1_3_0_n16), .S(n47), .Z(
        int_data_y_3__0__3_) );
  MUX2_X1 pe_1_3_0_U80 ( .A(pe_1_3_0_n18), .B(pe_1_3_0_n17), .S(pe_1_3_0_n60), 
        .Z(pe_1_3_0_n19) );
  MUX2_X1 pe_1_3_0_U79 ( .A(pe_1_3_0_int_q_reg_v[23]), .B(
        pe_1_3_0_int_q_reg_v[19]), .S(pe_1_3_0_n55), .Z(pe_1_3_0_n18) );
  MUX2_X1 pe_1_3_0_U78 ( .A(pe_1_3_0_int_q_reg_v[15]), .B(
        pe_1_3_0_int_q_reg_v[11]), .S(pe_1_3_0_n55), .Z(pe_1_3_0_n17) );
  MUX2_X1 pe_1_3_0_U77 ( .A(pe_1_3_0_int_q_reg_v[7]), .B(
        pe_1_3_0_int_q_reg_v[3]), .S(pe_1_3_0_n55), .Z(pe_1_3_0_n16) );
  MUX2_X1 pe_1_3_0_U76 ( .A(pe_1_3_0_n15), .B(pe_1_3_0_n12), .S(n47), .Z(
        int_data_y_3__0__2_) );
  MUX2_X1 pe_1_3_0_U75 ( .A(pe_1_3_0_n14), .B(pe_1_3_0_n13), .S(pe_1_3_0_n60), 
        .Z(pe_1_3_0_n15) );
  MUX2_X1 pe_1_3_0_U74 ( .A(pe_1_3_0_int_q_reg_v[22]), .B(
        pe_1_3_0_int_q_reg_v[18]), .S(pe_1_3_0_n55), .Z(pe_1_3_0_n14) );
  MUX2_X1 pe_1_3_0_U73 ( .A(pe_1_3_0_int_q_reg_v[14]), .B(
        pe_1_3_0_int_q_reg_v[10]), .S(pe_1_3_0_n55), .Z(pe_1_3_0_n13) );
  MUX2_X1 pe_1_3_0_U72 ( .A(pe_1_3_0_int_q_reg_v[6]), .B(
        pe_1_3_0_int_q_reg_v[2]), .S(pe_1_3_0_n55), .Z(pe_1_3_0_n12) );
  MUX2_X1 pe_1_3_0_U71 ( .A(pe_1_3_0_n11), .B(pe_1_3_0_n8), .S(n47), .Z(
        int_data_y_3__0__1_) );
  MUX2_X1 pe_1_3_0_U70 ( .A(pe_1_3_0_n10), .B(pe_1_3_0_n9), .S(pe_1_3_0_n60), 
        .Z(pe_1_3_0_n11) );
  MUX2_X1 pe_1_3_0_U69 ( .A(pe_1_3_0_int_q_reg_v[21]), .B(
        pe_1_3_0_int_q_reg_v[17]), .S(pe_1_3_0_n55), .Z(pe_1_3_0_n10) );
  MUX2_X1 pe_1_3_0_U68 ( .A(pe_1_3_0_int_q_reg_v[13]), .B(
        pe_1_3_0_int_q_reg_v[9]), .S(pe_1_3_0_n55), .Z(pe_1_3_0_n9) );
  MUX2_X1 pe_1_3_0_U67 ( .A(pe_1_3_0_int_q_reg_v[5]), .B(
        pe_1_3_0_int_q_reg_v[1]), .S(pe_1_3_0_n55), .Z(pe_1_3_0_n8) );
  MUX2_X1 pe_1_3_0_U66 ( .A(pe_1_3_0_n7), .B(pe_1_3_0_n4), .S(n47), .Z(
        int_data_y_3__0__0_) );
  MUX2_X1 pe_1_3_0_U65 ( .A(pe_1_3_0_n6), .B(pe_1_3_0_n5), .S(pe_1_3_0_n60), 
        .Z(pe_1_3_0_n7) );
  MUX2_X1 pe_1_3_0_U64 ( .A(pe_1_3_0_int_q_reg_v[20]), .B(
        pe_1_3_0_int_q_reg_v[16]), .S(pe_1_3_0_n55), .Z(pe_1_3_0_n6) );
  MUX2_X1 pe_1_3_0_U63 ( .A(pe_1_3_0_int_q_reg_v[12]), .B(
        pe_1_3_0_int_q_reg_v[8]), .S(pe_1_3_0_n55), .Z(pe_1_3_0_n5) );
  MUX2_X1 pe_1_3_0_U62 ( .A(pe_1_3_0_int_q_reg_v[4]), .B(
        pe_1_3_0_int_q_reg_v[0]), .S(pe_1_3_0_n55), .Z(pe_1_3_0_n4) );
  AND2_X1 pe_1_3_0_U61 ( .A1(pe_1_3_0_o_data_h_3_), .A2(n27), .ZN(
        pe_1_3_0_int_data_3_) );
  NAND2_X1 pe_1_3_0_U60 ( .A1(pe_1_3_0_int_data_0_), .A2(pe_1_3_0_n3), .ZN(
        pe_1_3_0_sub_81_carry[1]) );
  INV_X1 pe_1_3_0_U59 ( .A(pe_1_3_0_int_data_1_), .ZN(pe_1_3_0_n71) );
  AOI222_X1 pe_1_3_0_U58 ( .A1(pe_1_3_0_n62), .A2(int_data_res_4__0__7_), .B1(
        pe_1_3_0_N85), .B2(pe_1_3_0_n27), .C1(pe_1_3_0_N77), .C2(pe_1_3_0_n28), 
        .ZN(pe_1_3_0_n26) );
  INV_X1 pe_1_3_0_U57 ( .A(pe_1_3_0_n26), .ZN(pe_1_3_0_n74) );
  AOI222_X1 pe_1_3_0_U52 ( .A1(int_data_res_4__0__1_), .A2(pe_1_3_0_n62), .B1(
        pe_1_3_0_N79), .B2(pe_1_3_0_n27), .C1(pe_1_3_0_N71), .C2(pe_1_3_0_n28), 
        .ZN(pe_1_3_0_n34) );
  INV_X1 pe_1_3_0_U51 ( .A(pe_1_3_0_n34), .ZN(pe_1_3_0_n80) );
  AOI222_X1 pe_1_3_0_U50 ( .A1(int_data_res_4__0__2_), .A2(pe_1_3_0_n62), .B1(
        pe_1_3_0_N80), .B2(pe_1_3_0_n27), .C1(pe_1_3_0_N72), .C2(pe_1_3_0_n28), 
        .ZN(pe_1_3_0_n33) );
  INV_X1 pe_1_3_0_U49 ( .A(pe_1_3_0_n33), .ZN(pe_1_3_0_n79) );
  AOI222_X1 pe_1_3_0_U48 ( .A1(int_data_res_4__0__6_), .A2(pe_1_3_0_n62), .B1(
        pe_1_3_0_N84), .B2(pe_1_3_0_n27), .C1(pe_1_3_0_N76), .C2(pe_1_3_0_n28), 
        .ZN(pe_1_3_0_n29) );
  INV_X1 pe_1_3_0_U47 ( .A(pe_1_3_0_n29), .ZN(pe_1_3_0_n75) );
  AND2_X1 pe_1_3_0_U46 ( .A1(pe_1_3_0_o_data_h_2_), .A2(n27), .ZN(
        pe_1_3_0_int_data_2_) );
  AND2_X1 pe_1_3_0_U45 ( .A1(pe_1_3_0_o_data_h_1_), .A2(n27), .ZN(
        pe_1_3_0_int_data_1_) );
  INV_X1 pe_1_3_0_U44 ( .A(pe_1_3_0_int_data_2_), .ZN(pe_1_3_0_n72) );
  AND2_X1 pe_1_3_0_U43 ( .A1(pe_1_3_0_int_data_0_), .A2(int_data_res_3__0__0_), 
        .ZN(pe_1_3_0_n2) );
  AND2_X1 pe_1_3_0_U42 ( .A1(pe_1_3_0_o_data_h_0_), .A2(n27), .ZN(
        pe_1_3_0_int_data_0_) );
  XNOR2_X1 pe_1_3_0_U41 ( .A(pe_1_3_0_n70), .B(int_data_res_3__0__0_), .ZN(
        pe_1_3_0_N70) );
  AOI222_X1 pe_1_3_0_U40 ( .A1(int_data_res_4__0__0_), .A2(pe_1_3_0_n62), .B1(
        pe_1_3_0_n1), .B2(pe_1_3_0_n27), .C1(pe_1_3_0_N70), .C2(pe_1_3_0_n28), 
        .ZN(pe_1_3_0_n35) );
  INV_X1 pe_1_3_0_U39 ( .A(pe_1_3_0_n35), .ZN(pe_1_3_0_n81) );
  AOI222_X1 pe_1_3_0_U38 ( .A1(int_data_res_4__0__3_), .A2(pe_1_3_0_n62), .B1(
        pe_1_3_0_N81), .B2(pe_1_3_0_n27), .C1(pe_1_3_0_N73), .C2(pe_1_3_0_n28), 
        .ZN(pe_1_3_0_n32) );
  INV_X1 pe_1_3_0_U37 ( .A(pe_1_3_0_n32), .ZN(pe_1_3_0_n78) );
  AOI222_X1 pe_1_3_0_U36 ( .A1(int_data_res_4__0__4_), .A2(pe_1_3_0_n62), .B1(
        pe_1_3_0_N82), .B2(pe_1_3_0_n27), .C1(pe_1_3_0_N74), .C2(pe_1_3_0_n28), 
        .ZN(pe_1_3_0_n31) );
  INV_X1 pe_1_3_0_U35 ( .A(pe_1_3_0_n31), .ZN(pe_1_3_0_n77) );
  AOI222_X1 pe_1_3_0_U34 ( .A1(int_data_res_4__0__5_), .A2(pe_1_3_0_n62), .B1(
        pe_1_3_0_N83), .B2(pe_1_3_0_n27), .C1(pe_1_3_0_N75), .C2(pe_1_3_0_n28), 
        .ZN(pe_1_3_0_n30) );
  INV_X1 pe_1_3_0_U33 ( .A(pe_1_3_0_n30), .ZN(pe_1_3_0_n76) );
  NOR3_X1 pe_1_3_0_U32 ( .A1(pe_1_3_0_n58), .A2(pe_1_3_0_n63), .A3(int_ckg[39]), .ZN(pe_1_3_0_n36) );
  OR2_X1 pe_1_3_0_U31 ( .A1(pe_1_3_0_n36), .A2(pe_1_3_0_n62), .ZN(pe_1_3_0_N90) );
  INV_X1 pe_1_3_0_U30 ( .A(pe_1_3_0_int_data_0_), .ZN(pe_1_3_0_n70) );
  INV_X1 pe_1_3_0_U29 ( .A(n39), .ZN(pe_1_3_0_n61) );
  INV_X1 pe_1_3_0_U28 ( .A(n33), .ZN(pe_1_3_0_n59) );
  INV_X1 pe_1_3_0_U27 ( .A(pe_1_3_0_int_data_3_), .ZN(pe_1_3_0_n73) );
  BUF_X1 pe_1_3_0_U26 ( .A(n61), .Z(pe_1_3_0_n62) );
  NAND2_X1 pe_1_3_0_U25 ( .A1(pe_1_3_0_n44), .A2(pe_1_3_0_n59), .ZN(
        pe_1_3_0_n41) );
  AND3_X1 pe_1_3_0_U24 ( .A1(n75), .A2(pe_1_3_0_n61), .A3(n47), .ZN(
        pe_1_3_0_n44) );
  NOR2_X1 pe_1_3_0_U23 ( .A1(pe_1_3_0_n67), .A2(n47), .ZN(pe_1_3_0_n43) );
  NOR2_X1 pe_1_3_0_U22 ( .A1(pe_1_3_0_n57), .A2(pe_1_3_0_n62), .ZN(
        pe_1_3_0_n28) );
  NOR2_X1 pe_1_3_0_U21 ( .A1(n19), .A2(pe_1_3_0_n62), .ZN(pe_1_3_0_n27) );
  INV_X1 pe_1_3_0_U20 ( .A(pe_1_3_0_n41), .ZN(pe_1_3_0_n87) );
  INV_X1 pe_1_3_0_U19 ( .A(pe_1_3_0_n37), .ZN(pe_1_3_0_n85) );
  INV_X1 pe_1_3_0_U18 ( .A(pe_1_3_0_n38), .ZN(pe_1_3_0_n84) );
  INV_X1 pe_1_3_0_U17 ( .A(pe_1_3_0_n39), .ZN(pe_1_3_0_n83) );
  NOR2_X1 pe_1_3_0_U16 ( .A1(pe_1_3_0_n65), .A2(pe_1_3_0_n42), .ZN(
        pe_1_3_0_N59) );
  NOR2_X1 pe_1_3_0_U15 ( .A1(pe_1_3_0_n65), .A2(pe_1_3_0_n41), .ZN(
        pe_1_3_0_N60) );
  NOR2_X1 pe_1_3_0_U14 ( .A1(pe_1_3_0_n65), .A2(pe_1_3_0_n38), .ZN(
        pe_1_3_0_N63) );
  NOR2_X1 pe_1_3_0_U13 ( .A1(pe_1_3_0_n65), .A2(pe_1_3_0_n40), .ZN(
        pe_1_3_0_N61) );
  NOR2_X1 pe_1_3_0_U12 ( .A1(pe_1_3_0_n65), .A2(pe_1_3_0_n39), .ZN(
        pe_1_3_0_N62) );
  NOR2_X1 pe_1_3_0_U11 ( .A1(pe_1_3_0_n37), .A2(pe_1_3_0_n65), .ZN(
        pe_1_3_0_N64) );
  NAND2_X1 pe_1_3_0_U10 ( .A1(pe_1_3_0_n44), .A2(n33), .ZN(pe_1_3_0_n42) );
  BUF_X1 pe_1_3_0_U9 ( .A(n33), .Z(pe_1_3_0_n55) );
  BUF_X1 pe_1_3_0_U8 ( .A(n33), .Z(pe_1_3_0_n56) );
  INV_X1 pe_1_3_0_U7 ( .A(pe_1_3_0_n66), .ZN(pe_1_3_0_n63) );
  INV_X1 pe_1_3_0_U6 ( .A(pe_1_3_0_n42), .ZN(pe_1_3_0_n86) );
  INV_X1 pe_1_3_0_U5 ( .A(pe_1_3_0_n40), .ZN(pe_1_3_0_n82) );
  INV_X2 pe_1_3_0_U4 ( .A(n83), .ZN(pe_1_3_0_n69) );
  XOR2_X1 pe_1_3_0_U3 ( .A(pe_1_3_0_int_data_0_), .B(int_data_res_3__0__0_), 
        .Z(pe_1_3_0_n1) );
  DFFR_X1 pe_1_3_0_int_q_acc_reg_0_ ( .D(pe_1_3_0_n81), .CK(pe_1_3_0_net5680), 
        .RN(pe_1_3_0_n69), .Q(int_data_res_3__0__0_), .QN(pe_1_3_0_n3) );
  DFFR_X1 pe_1_3_0_int_q_reg_v_reg_0__0_ ( .D(int_data_y_4__0__0_), .CK(
        pe_1_3_0_net5650), .RN(pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_v[20]) );
  DFFR_X1 pe_1_3_0_int_q_reg_v_reg_0__1_ ( .D(int_data_y_4__0__1_), .CK(
        pe_1_3_0_net5650), .RN(pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_v[21]) );
  DFFR_X1 pe_1_3_0_int_q_reg_v_reg_0__2_ ( .D(int_data_y_4__0__2_), .CK(
        pe_1_3_0_net5650), .RN(pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_v[22]) );
  DFFR_X1 pe_1_3_0_int_q_reg_v_reg_0__3_ ( .D(int_data_y_4__0__3_), .CK(
        pe_1_3_0_net5650), .RN(pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_v[23]) );
  DFFR_X1 pe_1_3_0_int_q_reg_v_reg_1__0_ ( .D(int_data_y_4__0__0_), .CK(
        pe_1_3_0_net5655), .RN(pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_v[16]) );
  DFFR_X1 pe_1_3_0_int_q_reg_v_reg_1__1_ ( .D(int_data_y_4__0__1_), .CK(
        pe_1_3_0_net5655), .RN(pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_v[17]) );
  DFFR_X1 pe_1_3_0_int_q_reg_v_reg_1__2_ ( .D(int_data_y_4__0__2_), .CK(
        pe_1_3_0_net5655), .RN(pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_v[18]) );
  DFFR_X1 pe_1_3_0_int_q_reg_v_reg_1__3_ ( .D(int_data_y_4__0__3_), .CK(
        pe_1_3_0_net5655), .RN(pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_v[19]) );
  DFFR_X1 pe_1_3_0_int_q_reg_v_reg_2__0_ ( .D(int_data_y_4__0__0_), .CK(
        pe_1_3_0_net5660), .RN(pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_v[12]) );
  DFFR_X1 pe_1_3_0_int_q_reg_v_reg_2__1_ ( .D(int_data_y_4__0__1_), .CK(
        pe_1_3_0_net5660), .RN(pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_v[13]) );
  DFFR_X1 pe_1_3_0_int_q_reg_v_reg_2__2_ ( .D(int_data_y_4__0__2_), .CK(
        pe_1_3_0_net5660), .RN(pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_v[14]) );
  DFFR_X1 pe_1_3_0_int_q_reg_v_reg_2__3_ ( .D(int_data_y_4__0__3_), .CK(
        pe_1_3_0_net5660), .RN(pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_v[15]) );
  DFFR_X1 pe_1_3_0_int_q_reg_v_reg_3__0_ ( .D(int_data_y_4__0__0_), .CK(
        pe_1_3_0_net5665), .RN(pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_v[8]) );
  DFFR_X1 pe_1_3_0_int_q_reg_v_reg_3__1_ ( .D(int_data_y_4__0__1_), .CK(
        pe_1_3_0_net5665), .RN(pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_v[9]) );
  DFFR_X1 pe_1_3_0_int_q_reg_v_reg_3__2_ ( .D(int_data_y_4__0__2_), .CK(
        pe_1_3_0_net5665), .RN(pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_v[10]) );
  DFFR_X1 pe_1_3_0_int_q_reg_v_reg_3__3_ ( .D(int_data_y_4__0__3_), .CK(
        pe_1_3_0_net5665), .RN(pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_v[11]) );
  DFFR_X1 pe_1_3_0_int_q_reg_v_reg_4__0_ ( .D(int_data_y_4__0__0_), .CK(
        pe_1_3_0_net5670), .RN(pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_v[4]) );
  DFFR_X1 pe_1_3_0_int_q_reg_v_reg_4__1_ ( .D(int_data_y_4__0__1_), .CK(
        pe_1_3_0_net5670), .RN(pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_v[5]) );
  DFFR_X1 pe_1_3_0_int_q_reg_v_reg_4__2_ ( .D(int_data_y_4__0__2_), .CK(
        pe_1_3_0_net5670), .RN(pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_v[6]) );
  DFFR_X1 pe_1_3_0_int_q_reg_v_reg_4__3_ ( .D(int_data_y_4__0__3_), .CK(
        pe_1_3_0_net5670), .RN(pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_v[7]) );
  DFFR_X1 pe_1_3_0_int_q_reg_v_reg_5__0_ ( .D(int_data_y_4__0__0_), .CK(
        pe_1_3_0_net5675), .RN(pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_v[0]) );
  DFFR_X1 pe_1_3_0_int_q_reg_v_reg_5__1_ ( .D(int_data_y_4__0__1_), .CK(
        pe_1_3_0_net5675), .RN(pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_v[1]) );
  DFFR_X1 pe_1_3_0_int_q_reg_v_reg_5__2_ ( .D(int_data_y_4__0__2_), .CK(
        pe_1_3_0_net5675), .RN(pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_v[2]) );
  DFFR_X1 pe_1_3_0_int_q_reg_v_reg_5__3_ ( .D(int_data_y_4__0__3_), .CK(
        pe_1_3_0_net5675), .RN(pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_3_0_int_q_reg_h_reg_0__0_ ( .D(int_data_x_3__1__0_), .SI(
        int_data_y_4__0__0_), .SE(pe_1_3_0_n63), .CK(pe_1_3_0_net5619), .RN(
        pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_3_0_int_q_reg_h_reg_0__1_ ( .D(int_data_x_3__1__1_), .SI(
        int_data_y_4__0__1_), .SE(pe_1_3_0_n63), .CK(pe_1_3_0_net5619), .RN(
        pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_3_0_int_q_reg_h_reg_0__2_ ( .D(int_data_x_3__1__2_), .SI(
        int_data_y_4__0__2_), .SE(pe_1_3_0_n63), .CK(pe_1_3_0_net5619), .RN(
        pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_3_0_int_q_reg_h_reg_0__3_ ( .D(int_data_x_3__1__3_), .SI(
        int_data_y_4__0__3_), .SE(pe_1_3_0_n63), .CK(pe_1_3_0_net5619), .RN(
        pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_3_0_int_q_reg_h_reg_1__0_ ( .D(int_data_x_3__1__0_), .SI(
        int_data_y_4__0__0_), .SE(pe_1_3_0_n63), .CK(pe_1_3_0_net5625), .RN(
        pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_3_0_int_q_reg_h_reg_1__1_ ( .D(int_data_x_3__1__1_), .SI(
        int_data_y_4__0__1_), .SE(pe_1_3_0_n63), .CK(pe_1_3_0_net5625), .RN(
        pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_3_0_int_q_reg_h_reg_1__2_ ( .D(int_data_x_3__1__2_), .SI(
        int_data_y_4__0__2_), .SE(pe_1_3_0_n63), .CK(pe_1_3_0_net5625), .RN(
        pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_3_0_int_q_reg_h_reg_1__3_ ( .D(int_data_x_3__1__3_), .SI(
        int_data_y_4__0__3_), .SE(pe_1_3_0_n63), .CK(pe_1_3_0_net5625), .RN(
        pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_3_0_int_q_reg_h_reg_2__0_ ( .D(int_data_x_3__1__0_), .SI(
        int_data_y_4__0__0_), .SE(pe_1_3_0_n63), .CK(pe_1_3_0_net5630), .RN(
        pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_3_0_int_q_reg_h_reg_2__1_ ( .D(int_data_x_3__1__1_), .SI(
        int_data_y_4__0__1_), .SE(pe_1_3_0_n63), .CK(pe_1_3_0_net5630), .RN(
        pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_3_0_int_q_reg_h_reg_2__2_ ( .D(int_data_x_3__1__2_), .SI(
        int_data_y_4__0__2_), .SE(pe_1_3_0_n63), .CK(pe_1_3_0_net5630), .RN(
        pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_3_0_int_q_reg_h_reg_2__3_ ( .D(int_data_x_3__1__3_), .SI(
        int_data_y_4__0__3_), .SE(pe_1_3_0_n63), .CK(pe_1_3_0_net5630), .RN(
        pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_3_0_int_q_reg_h_reg_3__0_ ( .D(int_data_x_3__1__0_), .SI(
        int_data_y_4__0__0_), .SE(pe_1_3_0_n63), .CK(pe_1_3_0_net5635), .RN(
        pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_3_0_int_q_reg_h_reg_3__1_ ( .D(int_data_x_3__1__1_), .SI(
        int_data_y_4__0__1_), .SE(pe_1_3_0_n63), .CK(pe_1_3_0_net5635), .RN(
        pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_3_0_int_q_reg_h_reg_3__2_ ( .D(int_data_x_3__1__2_), .SI(
        int_data_y_4__0__2_), .SE(pe_1_3_0_n63), .CK(pe_1_3_0_net5635), .RN(
        pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_3_0_int_q_reg_h_reg_3__3_ ( .D(int_data_x_3__1__3_), .SI(
        int_data_y_4__0__3_), .SE(pe_1_3_0_n63), .CK(pe_1_3_0_net5635), .RN(
        pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_3_0_int_q_reg_h_reg_4__0_ ( .D(int_data_x_3__1__0_), .SI(
        int_data_y_4__0__0_), .SE(pe_1_3_0_n64), .CK(pe_1_3_0_net5640), .RN(
        pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_3_0_int_q_reg_h_reg_4__1_ ( .D(int_data_x_3__1__1_), .SI(
        int_data_y_4__0__1_), .SE(pe_1_3_0_n64), .CK(pe_1_3_0_net5640), .RN(
        pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_3_0_int_q_reg_h_reg_4__2_ ( .D(int_data_x_3__1__2_), .SI(
        int_data_y_4__0__2_), .SE(pe_1_3_0_n64), .CK(pe_1_3_0_net5640), .RN(
        pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_3_0_int_q_reg_h_reg_4__3_ ( .D(int_data_x_3__1__3_), .SI(
        int_data_y_4__0__3_), .SE(pe_1_3_0_n64), .CK(pe_1_3_0_net5640), .RN(
        pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_3_0_int_q_reg_h_reg_5__0_ ( .D(int_data_x_3__1__0_), .SI(
        int_data_y_4__0__0_), .SE(pe_1_3_0_n64), .CK(pe_1_3_0_net5645), .RN(
        pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_3_0_int_q_reg_h_reg_5__1_ ( .D(int_data_x_3__1__1_), .SI(
        int_data_y_4__0__1_), .SE(pe_1_3_0_n64), .CK(pe_1_3_0_net5645), .RN(
        pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_3_0_int_q_reg_h_reg_5__2_ ( .D(int_data_x_3__1__2_), .SI(
        int_data_y_4__0__2_), .SE(pe_1_3_0_n64), .CK(pe_1_3_0_net5645), .RN(
        pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_3_0_int_q_reg_h_reg_5__3_ ( .D(int_data_x_3__1__3_), .SI(
        int_data_y_4__0__3_), .SE(pe_1_3_0_n64), .CK(pe_1_3_0_net5645), .RN(
        pe_1_3_0_n69), .Q(pe_1_3_0_int_q_reg_h[3]) );
  FA_X1 pe_1_3_0_sub_81_U2_7 ( .A(int_data_res_3__0__7_), .B(pe_1_3_0_n73), 
        .CI(pe_1_3_0_sub_81_carry[7]), .S(pe_1_3_0_N77) );
  FA_X1 pe_1_3_0_sub_81_U2_6 ( .A(int_data_res_3__0__6_), .B(pe_1_3_0_n73), 
        .CI(pe_1_3_0_sub_81_carry[6]), .CO(pe_1_3_0_sub_81_carry[7]), .S(
        pe_1_3_0_N76) );
  FA_X1 pe_1_3_0_sub_81_U2_5 ( .A(int_data_res_3__0__5_), .B(pe_1_3_0_n73), 
        .CI(pe_1_3_0_sub_81_carry[5]), .CO(pe_1_3_0_sub_81_carry[6]), .S(
        pe_1_3_0_N75) );
  FA_X1 pe_1_3_0_sub_81_U2_4 ( .A(int_data_res_3__0__4_), .B(pe_1_3_0_n73), 
        .CI(pe_1_3_0_sub_81_carry[4]), .CO(pe_1_3_0_sub_81_carry[5]), .S(
        pe_1_3_0_N74) );
  FA_X1 pe_1_3_0_sub_81_U2_3 ( .A(int_data_res_3__0__3_), .B(pe_1_3_0_n73), 
        .CI(pe_1_3_0_sub_81_carry[3]), .CO(pe_1_3_0_sub_81_carry[4]), .S(
        pe_1_3_0_N73) );
  FA_X1 pe_1_3_0_sub_81_U2_2 ( .A(int_data_res_3__0__2_), .B(pe_1_3_0_n72), 
        .CI(pe_1_3_0_sub_81_carry[2]), .CO(pe_1_3_0_sub_81_carry[3]), .S(
        pe_1_3_0_N72) );
  FA_X1 pe_1_3_0_sub_81_U2_1 ( .A(int_data_res_3__0__1_), .B(pe_1_3_0_n71), 
        .CI(pe_1_3_0_sub_81_carry[1]), .CO(pe_1_3_0_sub_81_carry[2]), .S(
        pe_1_3_0_N71) );
  FA_X1 pe_1_3_0_add_83_U1_7 ( .A(int_data_res_3__0__7_), .B(
        pe_1_3_0_int_data_3_), .CI(pe_1_3_0_add_83_carry[7]), .S(pe_1_3_0_N85)
         );
  FA_X1 pe_1_3_0_add_83_U1_6 ( .A(int_data_res_3__0__6_), .B(
        pe_1_3_0_int_data_3_), .CI(pe_1_3_0_add_83_carry[6]), .CO(
        pe_1_3_0_add_83_carry[7]), .S(pe_1_3_0_N84) );
  FA_X1 pe_1_3_0_add_83_U1_5 ( .A(int_data_res_3__0__5_), .B(
        pe_1_3_0_int_data_3_), .CI(pe_1_3_0_add_83_carry[5]), .CO(
        pe_1_3_0_add_83_carry[6]), .S(pe_1_3_0_N83) );
  FA_X1 pe_1_3_0_add_83_U1_4 ( .A(int_data_res_3__0__4_), .B(
        pe_1_3_0_int_data_3_), .CI(pe_1_3_0_add_83_carry[4]), .CO(
        pe_1_3_0_add_83_carry[5]), .S(pe_1_3_0_N82) );
  FA_X1 pe_1_3_0_add_83_U1_3 ( .A(int_data_res_3__0__3_), .B(
        pe_1_3_0_int_data_3_), .CI(pe_1_3_0_add_83_carry[3]), .CO(
        pe_1_3_0_add_83_carry[4]), .S(pe_1_3_0_N81) );
  FA_X1 pe_1_3_0_add_83_U1_2 ( .A(int_data_res_3__0__2_), .B(
        pe_1_3_0_int_data_2_), .CI(pe_1_3_0_add_83_carry[2]), .CO(
        pe_1_3_0_add_83_carry[3]), .S(pe_1_3_0_N80) );
  FA_X1 pe_1_3_0_add_83_U1_1 ( .A(int_data_res_3__0__1_), .B(
        pe_1_3_0_int_data_1_), .CI(pe_1_3_0_n2), .CO(pe_1_3_0_add_83_carry[2]), 
        .S(pe_1_3_0_N79) );
  NAND3_X1 pe_1_3_0_U56 ( .A1(n33), .A2(pe_1_3_0_n43), .A3(pe_1_3_0_n60), .ZN(
        pe_1_3_0_n40) );
  NAND3_X1 pe_1_3_0_U55 ( .A1(pe_1_3_0_n43), .A2(pe_1_3_0_n59), .A3(
        pe_1_3_0_n60), .ZN(pe_1_3_0_n39) );
  NAND3_X1 pe_1_3_0_U54 ( .A1(pe_1_3_0_n43), .A2(pe_1_3_0_n61), .A3(n33), .ZN(
        pe_1_3_0_n38) );
  NAND3_X1 pe_1_3_0_U53 ( .A1(pe_1_3_0_n59), .A2(pe_1_3_0_n61), .A3(
        pe_1_3_0_n43), .ZN(pe_1_3_0_n37) );
  DFFR_X1 pe_1_3_0_int_q_acc_reg_6_ ( .D(pe_1_3_0_n75), .CK(pe_1_3_0_net5680), 
        .RN(pe_1_3_0_n68), .Q(int_data_res_3__0__6_) );
  DFFR_X1 pe_1_3_0_int_q_acc_reg_5_ ( .D(pe_1_3_0_n76), .CK(pe_1_3_0_net5680), 
        .RN(pe_1_3_0_n68), .Q(int_data_res_3__0__5_) );
  DFFR_X1 pe_1_3_0_int_q_acc_reg_4_ ( .D(pe_1_3_0_n77), .CK(pe_1_3_0_net5680), 
        .RN(pe_1_3_0_n68), .Q(int_data_res_3__0__4_) );
  DFFR_X1 pe_1_3_0_int_q_acc_reg_3_ ( .D(pe_1_3_0_n78), .CK(pe_1_3_0_net5680), 
        .RN(pe_1_3_0_n68), .Q(int_data_res_3__0__3_) );
  DFFR_X1 pe_1_3_0_int_q_acc_reg_2_ ( .D(pe_1_3_0_n79), .CK(pe_1_3_0_net5680), 
        .RN(pe_1_3_0_n68), .Q(int_data_res_3__0__2_) );
  DFFR_X1 pe_1_3_0_int_q_acc_reg_1_ ( .D(pe_1_3_0_n80), .CK(pe_1_3_0_net5680), 
        .RN(pe_1_3_0_n68), .Q(int_data_res_3__0__1_) );
  DFFR_X1 pe_1_3_0_int_q_acc_reg_7_ ( .D(pe_1_3_0_n74), .CK(pe_1_3_0_net5680), 
        .RN(pe_1_3_0_n68), .Q(int_data_res_3__0__7_) );
  CLKGATETST_X1 pe_1_3_0_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_3_0_n85), .SE(1'b0), .GCK(pe_1_3_0_net5619) );
  CLKGATETST_X1 pe_1_3_0_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_3_0_n84), .SE(1'b0), .GCK(pe_1_3_0_net5625) );
  CLKGATETST_X1 pe_1_3_0_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_3_0_n83), .SE(1'b0), .GCK(pe_1_3_0_net5630) );
  CLKGATETST_X1 pe_1_3_0_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_3_0_n82), .SE(1'b0), .GCK(pe_1_3_0_net5635) );
  CLKGATETST_X1 pe_1_3_0_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_3_0_n87), .SE(1'b0), .GCK(pe_1_3_0_net5640) );
  CLKGATETST_X1 pe_1_3_0_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_3_0_n86), .SE(1'b0), .GCK(pe_1_3_0_net5645) );
  CLKGATETST_X1 pe_1_3_0_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_3_0_N64), .SE(1'b0), .GCK(pe_1_3_0_net5650) );
  CLKGATETST_X1 pe_1_3_0_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_3_0_N63), .SE(1'b0), .GCK(pe_1_3_0_net5655) );
  CLKGATETST_X1 pe_1_3_0_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_3_0_N62), .SE(1'b0), .GCK(pe_1_3_0_net5660) );
  CLKGATETST_X1 pe_1_3_0_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_3_0_N61), .SE(1'b0), .GCK(pe_1_3_0_net5665) );
  CLKGATETST_X1 pe_1_3_0_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_3_0_N60), .SE(1'b0), .GCK(pe_1_3_0_net5670) );
  CLKGATETST_X1 pe_1_3_0_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_3_0_N59), .SE(1'b0), .GCK(pe_1_3_0_net5675) );
  CLKGATETST_X1 pe_1_3_0_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_3_0_N90), .SE(1'b0), .GCK(pe_1_3_0_net5680) );
  CLKBUF_X1 pe_1_3_1_U108 ( .A(pe_1_3_1_n68), .Z(pe_1_3_1_n67) );
  INV_X1 pe_1_3_1_U107 ( .A(n75), .ZN(pe_1_3_1_n66) );
  INV_X1 pe_1_3_1_U106 ( .A(n67), .ZN(pe_1_3_1_n65) );
  INV_X1 pe_1_3_1_U105 ( .A(n67), .ZN(pe_1_3_1_n64) );
  INV_X1 pe_1_3_1_U104 ( .A(pe_1_3_1_n65), .ZN(pe_1_3_1_n63) );
  INV_X1 pe_1_3_1_U103 ( .A(n27), .ZN(pe_1_3_1_n58) );
  INV_X1 pe_1_3_1_U102 ( .A(n19), .ZN(pe_1_3_1_n57) );
  MUX2_X1 pe_1_3_1_U101 ( .A(pe_1_3_1_n54), .B(pe_1_3_1_n51), .S(n48), .Z(
        int_data_x_3__1__3_) );
  MUX2_X1 pe_1_3_1_U100 ( .A(pe_1_3_1_n53), .B(pe_1_3_1_n52), .S(n39), .Z(
        pe_1_3_1_n54) );
  MUX2_X1 pe_1_3_1_U99 ( .A(pe_1_3_1_int_q_reg_h[23]), .B(
        pe_1_3_1_int_q_reg_h[19]), .S(pe_1_3_1_n56), .Z(pe_1_3_1_n53) );
  MUX2_X1 pe_1_3_1_U98 ( .A(pe_1_3_1_int_q_reg_h[15]), .B(
        pe_1_3_1_int_q_reg_h[11]), .S(pe_1_3_1_n56), .Z(pe_1_3_1_n52) );
  MUX2_X1 pe_1_3_1_U97 ( .A(pe_1_3_1_int_q_reg_h[7]), .B(
        pe_1_3_1_int_q_reg_h[3]), .S(pe_1_3_1_n56), .Z(pe_1_3_1_n51) );
  MUX2_X1 pe_1_3_1_U96 ( .A(pe_1_3_1_n50), .B(pe_1_3_1_n47), .S(n48), .Z(
        int_data_x_3__1__2_) );
  MUX2_X1 pe_1_3_1_U95 ( .A(pe_1_3_1_n49), .B(pe_1_3_1_n48), .S(n39), .Z(
        pe_1_3_1_n50) );
  MUX2_X1 pe_1_3_1_U94 ( .A(pe_1_3_1_int_q_reg_h[22]), .B(
        pe_1_3_1_int_q_reg_h[18]), .S(pe_1_3_1_n56), .Z(pe_1_3_1_n49) );
  MUX2_X1 pe_1_3_1_U93 ( .A(pe_1_3_1_int_q_reg_h[14]), .B(
        pe_1_3_1_int_q_reg_h[10]), .S(pe_1_3_1_n56), .Z(pe_1_3_1_n48) );
  MUX2_X1 pe_1_3_1_U92 ( .A(pe_1_3_1_int_q_reg_h[6]), .B(
        pe_1_3_1_int_q_reg_h[2]), .S(pe_1_3_1_n56), .Z(pe_1_3_1_n47) );
  MUX2_X1 pe_1_3_1_U91 ( .A(pe_1_3_1_n46), .B(pe_1_3_1_n24), .S(n48), .Z(
        int_data_x_3__1__1_) );
  MUX2_X1 pe_1_3_1_U90 ( .A(pe_1_3_1_n45), .B(pe_1_3_1_n25), .S(n39), .Z(
        pe_1_3_1_n46) );
  MUX2_X1 pe_1_3_1_U89 ( .A(pe_1_3_1_int_q_reg_h[21]), .B(
        pe_1_3_1_int_q_reg_h[17]), .S(pe_1_3_1_n56), .Z(pe_1_3_1_n45) );
  MUX2_X1 pe_1_3_1_U88 ( .A(pe_1_3_1_int_q_reg_h[13]), .B(
        pe_1_3_1_int_q_reg_h[9]), .S(pe_1_3_1_n56), .Z(pe_1_3_1_n25) );
  MUX2_X1 pe_1_3_1_U87 ( .A(pe_1_3_1_int_q_reg_h[5]), .B(
        pe_1_3_1_int_q_reg_h[1]), .S(pe_1_3_1_n56), .Z(pe_1_3_1_n24) );
  MUX2_X1 pe_1_3_1_U86 ( .A(pe_1_3_1_n23), .B(pe_1_3_1_n20), .S(n48), .Z(
        int_data_x_3__1__0_) );
  MUX2_X1 pe_1_3_1_U85 ( .A(pe_1_3_1_n22), .B(pe_1_3_1_n21), .S(n39), .Z(
        pe_1_3_1_n23) );
  MUX2_X1 pe_1_3_1_U84 ( .A(pe_1_3_1_int_q_reg_h[20]), .B(
        pe_1_3_1_int_q_reg_h[16]), .S(pe_1_3_1_n56), .Z(pe_1_3_1_n22) );
  MUX2_X1 pe_1_3_1_U83 ( .A(pe_1_3_1_int_q_reg_h[12]), .B(
        pe_1_3_1_int_q_reg_h[8]), .S(pe_1_3_1_n56), .Z(pe_1_3_1_n21) );
  MUX2_X1 pe_1_3_1_U82 ( .A(pe_1_3_1_int_q_reg_h[4]), .B(
        pe_1_3_1_int_q_reg_h[0]), .S(pe_1_3_1_n56), .Z(pe_1_3_1_n20) );
  MUX2_X1 pe_1_3_1_U81 ( .A(pe_1_3_1_n19), .B(pe_1_3_1_n16), .S(n48), .Z(
        int_data_y_3__1__3_) );
  MUX2_X1 pe_1_3_1_U80 ( .A(pe_1_3_1_n18), .B(pe_1_3_1_n17), .S(n39), .Z(
        pe_1_3_1_n19) );
  MUX2_X1 pe_1_3_1_U79 ( .A(pe_1_3_1_int_q_reg_v[23]), .B(
        pe_1_3_1_int_q_reg_v[19]), .S(pe_1_3_1_n55), .Z(pe_1_3_1_n18) );
  MUX2_X1 pe_1_3_1_U78 ( .A(pe_1_3_1_int_q_reg_v[15]), .B(
        pe_1_3_1_int_q_reg_v[11]), .S(pe_1_3_1_n55), .Z(pe_1_3_1_n17) );
  MUX2_X1 pe_1_3_1_U77 ( .A(pe_1_3_1_int_q_reg_v[7]), .B(
        pe_1_3_1_int_q_reg_v[3]), .S(pe_1_3_1_n55), .Z(pe_1_3_1_n16) );
  MUX2_X1 pe_1_3_1_U76 ( .A(pe_1_3_1_n15), .B(pe_1_3_1_n12), .S(n48), .Z(
        int_data_y_3__1__2_) );
  MUX2_X1 pe_1_3_1_U75 ( .A(pe_1_3_1_n14), .B(pe_1_3_1_n13), .S(n39), .Z(
        pe_1_3_1_n15) );
  MUX2_X1 pe_1_3_1_U74 ( .A(pe_1_3_1_int_q_reg_v[22]), .B(
        pe_1_3_1_int_q_reg_v[18]), .S(pe_1_3_1_n55), .Z(pe_1_3_1_n14) );
  MUX2_X1 pe_1_3_1_U73 ( .A(pe_1_3_1_int_q_reg_v[14]), .B(
        pe_1_3_1_int_q_reg_v[10]), .S(pe_1_3_1_n55), .Z(pe_1_3_1_n13) );
  MUX2_X1 pe_1_3_1_U72 ( .A(pe_1_3_1_int_q_reg_v[6]), .B(
        pe_1_3_1_int_q_reg_v[2]), .S(pe_1_3_1_n55), .Z(pe_1_3_1_n12) );
  MUX2_X1 pe_1_3_1_U71 ( .A(pe_1_3_1_n11), .B(pe_1_3_1_n8), .S(n48), .Z(
        int_data_y_3__1__1_) );
  MUX2_X1 pe_1_3_1_U70 ( .A(pe_1_3_1_n10), .B(pe_1_3_1_n9), .S(n39), .Z(
        pe_1_3_1_n11) );
  MUX2_X1 pe_1_3_1_U69 ( .A(pe_1_3_1_int_q_reg_v[21]), .B(
        pe_1_3_1_int_q_reg_v[17]), .S(pe_1_3_1_n55), .Z(pe_1_3_1_n10) );
  MUX2_X1 pe_1_3_1_U68 ( .A(pe_1_3_1_int_q_reg_v[13]), .B(
        pe_1_3_1_int_q_reg_v[9]), .S(pe_1_3_1_n55), .Z(pe_1_3_1_n9) );
  MUX2_X1 pe_1_3_1_U67 ( .A(pe_1_3_1_int_q_reg_v[5]), .B(
        pe_1_3_1_int_q_reg_v[1]), .S(pe_1_3_1_n55), .Z(pe_1_3_1_n8) );
  MUX2_X1 pe_1_3_1_U66 ( .A(pe_1_3_1_n7), .B(pe_1_3_1_n4), .S(n48), .Z(
        int_data_y_3__1__0_) );
  MUX2_X1 pe_1_3_1_U65 ( .A(pe_1_3_1_n6), .B(pe_1_3_1_n5), .S(n39), .Z(
        pe_1_3_1_n7) );
  MUX2_X1 pe_1_3_1_U64 ( .A(pe_1_3_1_int_q_reg_v[20]), .B(
        pe_1_3_1_int_q_reg_v[16]), .S(pe_1_3_1_n55), .Z(pe_1_3_1_n6) );
  MUX2_X1 pe_1_3_1_U63 ( .A(pe_1_3_1_int_q_reg_v[12]), .B(
        pe_1_3_1_int_q_reg_v[8]), .S(pe_1_3_1_n55), .Z(pe_1_3_1_n5) );
  MUX2_X1 pe_1_3_1_U62 ( .A(pe_1_3_1_int_q_reg_v[4]), .B(
        pe_1_3_1_int_q_reg_v[0]), .S(pe_1_3_1_n55), .Z(pe_1_3_1_n4) );
  AOI222_X1 pe_1_3_1_U61 ( .A1(int_data_res_4__1__2_), .A2(pe_1_3_1_n61), .B1(
        pe_1_3_1_N80), .B2(pe_1_3_1_n27), .C1(pe_1_3_1_N72), .C2(pe_1_3_1_n28), 
        .ZN(pe_1_3_1_n33) );
  INV_X1 pe_1_3_1_U60 ( .A(pe_1_3_1_n33), .ZN(pe_1_3_1_n78) );
  AOI222_X1 pe_1_3_1_U59 ( .A1(int_data_res_4__1__6_), .A2(pe_1_3_1_n61), .B1(
        pe_1_3_1_N84), .B2(pe_1_3_1_n27), .C1(pe_1_3_1_N76), .C2(pe_1_3_1_n28), 
        .ZN(pe_1_3_1_n29) );
  INV_X1 pe_1_3_1_U58 ( .A(pe_1_3_1_n29), .ZN(pe_1_3_1_n74) );
  XNOR2_X1 pe_1_3_1_U57 ( .A(pe_1_3_1_n69), .B(int_data_res_3__1__0_), .ZN(
        pe_1_3_1_N70) );
  AOI222_X1 pe_1_3_1_U52 ( .A1(int_data_res_4__1__0_), .A2(pe_1_3_1_n61), .B1(
        pe_1_3_1_n1), .B2(pe_1_3_1_n27), .C1(pe_1_3_1_N70), .C2(pe_1_3_1_n28), 
        .ZN(pe_1_3_1_n35) );
  INV_X1 pe_1_3_1_U51 ( .A(pe_1_3_1_n35), .ZN(pe_1_3_1_n80) );
  AOI222_X1 pe_1_3_1_U50 ( .A1(int_data_res_4__1__1_), .A2(pe_1_3_1_n61), .B1(
        pe_1_3_1_N79), .B2(pe_1_3_1_n27), .C1(pe_1_3_1_N71), .C2(pe_1_3_1_n28), 
        .ZN(pe_1_3_1_n34) );
  INV_X1 pe_1_3_1_U49 ( .A(pe_1_3_1_n34), .ZN(pe_1_3_1_n79) );
  AOI222_X1 pe_1_3_1_U48 ( .A1(int_data_res_4__1__3_), .A2(pe_1_3_1_n61), .B1(
        pe_1_3_1_N81), .B2(pe_1_3_1_n27), .C1(pe_1_3_1_N73), .C2(pe_1_3_1_n28), 
        .ZN(pe_1_3_1_n32) );
  INV_X1 pe_1_3_1_U47 ( .A(pe_1_3_1_n32), .ZN(pe_1_3_1_n77) );
  AOI222_X1 pe_1_3_1_U46 ( .A1(int_data_res_4__1__4_), .A2(pe_1_3_1_n61), .B1(
        pe_1_3_1_N82), .B2(pe_1_3_1_n27), .C1(pe_1_3_1_N74), .C2(pe_1_3_1_n28), 
        .ZN(pe_1_3_1_n31) );
  INV_X1 pe_1_3_1_U45 ( .A(pe_1_3_1_n31), .ZN(pe_1_3_1_n76) );
  AOI222_X1 pe_1_3_1_U44 ( .A1(int_data_res_4__1__5_), .A2(pe_1_3_1_n61), .B1(
        pe_1_3_1_N83), .B2(pe_1_3_1_n27), .C1(pe_1_3_1_N75), .C2(pe_1_3_1_n28), 
        .ZN(pe_1_3_1_n30) );
  INV_X1 pe_1_3_1_U43 ( .A(pe_1_3_1_n30), .ZN(pe_1_3_1_n75) );
  NAND2_X1 pe_1_3_1_U42 ( .A1(pe_1_3_1_int_data_0_), .A2(pe_1_3_1_n3), .ZN(
        pe_1_3_1_sub_81_carry[1]) );
  INV_X1 pe_1_3_1_U41 ( .A(pe_1_3_1_int_data_1_), .ZN(pe_1_3_1_n70) );
  INV_X1 pe_1_3_1_U40 ( .A(pe_1_3_1_int_data_2_), .ZN(pe_1_3_1_n71) );
  AND2_X1 pe_1_3_1_U39 ( .A1(pe_1_3_1_int_data_0_), .A2(int_data_res_3__1__0_), 
        .ZN(pe_1_3_1_n2) );
  AOI222_X1 pe_1_3_1_U38 ( .A1(pe_1_3_1_n61), .A2(int_data_res_4__1__7_), .B1(
        pe_1_3_1_N85), .B2(pe_1_3_1_n27), .C1(pe_1_3_1_N77), .C2(pe_1_3_1_n28), 
        .ZN(pe_1_3_1_n26) );
  INV_X1 pe_1_3_1_U37 ( .A(pe_1_3_1_n26), .ZN(pe_1_3_1_n73) );
  NOR3_X1 pe_1_3_1_U36 ( .A1(pe_1_3_1_n58), .A2(pe_1_3_1_n62), .A3(int_ckg[38]), .ZN(pe_1_3_1_n36) );
  OR2_X1 pe_1_3_1_U35 ( .A1(pe_1_3_1_n36), .A2(pe_1_3_1_n61), .ZN(pe_1_3_1_N90) );
  INV_X1 pe_1_3_1_U34 ( .A(n39), .ZN(pe_1_3_1_n60) );
  AND2_X1 pe_1_3_1_U33 ( .A1(int_data_x_3__1__2_), .A2(n27), .ZN(
        pe_1_3_1_int_data_2_) );
  AND2_X1 pe_1_3_1_U32 ( .A1(int_data_x_3__1__1_), .A2(n27), .ZN(
        pe_1_3_1_int_data_1_) );
  AND2_X1 pe_1_3_1_U31 ( .A1(int_data_x_3__1__3_), .A2(n27), .ZN(
        pe_1_3_1_int_data_3_) );
  BUF_X1 pe_1_3_1_U30 ( .A(n61), .Z(pe_1_3_1_n61) );
  INV_X1 pe_1_3_1_U29 ( .A(n33), .ZN(pe_1_3_1_n59) );
  AND2_X1 pe_1_3_1_U28 ( .A1(int_data_x_3__1__0_), .A2(n27), .ZN(
        pe_1_3_1_int_data_0_) );
  NAND2_X1 pe_1_3_1_U27 ( .A1(pe_1_3_1_n44), .A2(pe_1_3_1_n59), .ZN(
        pe_1_3_1_n41) );
  AND3_X1 pe_1_3_1_U26 ( .A1(n75), .A2(pe_1_3_1_n60), .A3(n48), .ZN(
        pe_1_3_1_n44) );
  INV_X1 pe_1_3_1_U25 ( .A(pe_1_3_1_int_data_3_), .ZN(pe_1_3_1_n72) );
  NOR2_X1 pe_1_3_1_U24 ( .A1(pe_1_3_1_n66), .A2(n48), .ZN(pe_1_3_1_n43) );
  NOR2_X1 pe_1_3_1_U23 ( .A1(pe_1_3_1_n57), .A2(pe_1_3_1_n61), .ZN(
        pe_1_3_1_n28) );
  NOR2_X1 pe_1_3_1_U22 ( .A1(n19), .A2(pe_1_3_1_n61), .ZN(pe_1_3_1_n27) );
  INV_X1 pe_1_3_1_U21 ( .A(pe_1_3_1_int_data_0_), .ZN(pe_1_3_1_n69) );
  INV_X1 pe_1_3_1_U20 ( .A(pe_1_3_1_n41), .ZN(pe_1_3_1_n86) );
  INV_X1 pe_1_3_1_U19 ( .A(pe_1_3_1_n37), .ZN(pe_1_3_1_n84) );
  INV_X1 pe_1_3_1_U18 ( .A(pe_1_3_1_n38), .ZN(pe_1_3_1_n83) );
  INV_X1 pe_1_3_1_U17 ( .A(pe_1_3_1_n39), .ZN(pe_1_3_1_n82) );
  NOR2_X1 pe_1_3_1_U16 ( .A1(pe_1_3_1_n64), .A2(pe_1_3_1_n42), .ZN(
        pe_1_3_1_N59) );
  NOR2_X1 pe_1_3_1_U15 ( .A1(pe_1_3_1_n64), .A2(pe_1_3_1_n41), .ZN(
        pe_1_3_1_N60) );
  NOR2_X1 pe_1_3_1_U14 ( .A1(pe_1_3_1_n64), .A2(pe_1_3_1_n38), .ZN(
        pe_1_3_1_N63) );
  NOR2_X1 pe_1_3_1_U13 ( .A1(pe_1_3_1_n64), .A2(pe_1_3_1_n40), .ZN(
        pe_1_3_1_N61) );
  NOR2_X1 pe_1_3_1_U12 ( .A1(pe_1_3_1_n64), .A2(pe_1_3_1_n39), .ZN(
        pe_1_3_1_N62) );
  NOR2_X1 pe_1_3_1_U11 ( .A1(pe_1_3_1_n37), .A2(pe_1_3_1_n64), .ZN(
        pe_1_3_1_N64) );
  NAND2_X1 pe_1_3_1_U10 ( .A1(pe_1_3_1_n44), .A2(n33), .ZN(pe_1_3_1_n42) );
  BUF_X1 pe_1_3_1_U9 ( .A(n33), .Z(pe_1_3_1_n55) );
  INV_X1 pe_1_3_1_U8 ( .A(pe_1_3_1_n65), .ZN(pe_1_3_1_n62) );
  BUF_X1 pe_1_3_1_U7 ( .A(n33), .Z(pe_1_3_1_n56) );
  INV_X1 pe_1_3_1_U6 ( .A(pe_1_3_1_n42), .ZN(pe_1_3_1_n85) );
  INV_X1 pe_1_3_1_U5 ( .A(pe_1_3_1_n40), .ZN(pe_1_3_1_n81) );
  INV_X2 pe_1_3_1_U4 ( .A(n83), .ZN(pe_1_3_1_n68) );
  XOR2_X1 pe_1_3_1_U3 ( .A(pe_1_3_1_int_data_0_), .B(int_data_res_3__1__0_), 
        .Z(pe_1_3_1_n1) );
  DFFR_X1 pe_1_3_1_int_q_acc_reg_0_ ( .D(pe_1_3_1_n80), .CK(pe_1_3_1_net5602), 
        .RN(pe_1_3_1_n68), .Q(int_data_res_3__1__0_), .QN(pe_1_3_1_n3) );
  DFFR_X1 pe_1_3_1_int_q_reg_v_reg_0__0_ ( .D(int_data_y_4__1__0_), .CK(
        pe_1_3_1_net5572), .RN(pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_v[20]) );
  DFFR_X1 pe_1_3_1_int_q_reg_v_reg_0__1_ ( .D(int_data_y_4__1__1_), .CK(
        pe_1_3_1_net5572), .RN(pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_v[21]) );
  DFFR_X1 pe_1_3_1_int_q_reg_v_reg_0__2_ ( .D(int_data_y_4__1__2_), .CK(
        pe_1_3_1_net5572), .RN(pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_v[22]) );
  DFFR_X1 pe_1_3_1_int_q_reg_v_reg_0__3_ ( .D(int_data_y_4__1__3_), .CK(
        pe_1_3_1_net5572), .RN(pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_v[23]) );
  DFFR_X1 pe_1_3_1_int_q_reg_v_reg_1__0_ ( .D(int_data_y_4__1__0_), .CK(
        pe_1_3_1_net5577), .RN(pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_v[16]) );
  DFFR_X1 pe_1_3_1_int_q_reg_v_reg_1__1_ ( .D(int_data_y_4__1__1_), .CK(
        pe_1_3_1_net5577), .RN(pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_v[17]) );
  DFFR_X1 pe_1_3_1_int_q_reg_v_reg_1__2_ ( .D(int_data_y_4__1__2_), .CK(
        pe_1_3_1_net5577), .RN(pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_v[18]) );
  DFFR_X1 pe_1_3_1_int_q_reg_v_reg_1__3_ ( .D(int_data_y_4__1__3_), .CK(
        pe_1_3_1_net5577), .RN(pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_v[19]) );
  DFFR_X1 pe_1_3_1_int_q_reg_v_reg_2__0_ ( .D(int_data_y_4__1__0_), .CK(
        pe_1_3_1_net5582), .RN(pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_v[12]) );
  DFFR_X1 pe_1_3_1_int_q_reg_v_reg_2__1_ ( .D(int_data_y_4__1__1_), .CK(
        pe_1_3_1_net5582), .RN(pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_v[13]) );
  DFFR_X1 pe_1_3_1_int_q_reg_v_reg_2__2_ ( .D(int_data_y_4__1__2_), .CK(
        pe_1_3_1_net5582), .RN(pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_v[14]) );
  DFFR_X1 pe_1_3_1_int_q_reg_v_reg_2__3_ ( .D(int_data_y_4__1__3_), .CK(
        pe_1_3_1_net5582), .RN(pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_v[15]) );
  DFFR_X1 pe_1_3_1_int_q_reg_v_reg_3__0_ ( .D(int_data_y_4__1__0_), .CK(
        pe_1_3_1_net5587), .RN(pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_v[8]) );
  DFFR_X1 pe_1_3_1_int_q_reg_v_reg_3__1_ ( .D(int_data_y_4__1__1_), .CK(
        pe_1_3_1_net5587), .RN(pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_v[9]) );
  DFFR_X1 pe_1_3_1_int_q_reg_v_reg_3__2_ ( .D(int_data_y_4__1__2_), .CK(
        pe_1_3_1_net5587), .RN(pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_v[10]) );
  DFFR_X1 pe_1_3_1_int_q_reg_v_reg_3__3_ ( .D(int_data_y_4__1__3_), .CK(
        pe_1_3_1_net5587), .RN(pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_v[11]) );
  DFFR_X1 pe_1_3_1_int_q_reg_v_reg_4__0_ ( .D(int_data_y_4__1__0_), .CK(
        pe_1_3_1_net5592), .RN(pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_v[4]) );
  DFFR_X1 pe_1_3_1_int_q_reg_v_reg_4__1_ ( .D(int_data_y_4__1__1_), .CK(
        pe_1_3_1_net5592), .RN(pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_v[5]) );
  DFFR_X1 pe_1_3_1_int_q_reg_v_reg_4__2_ ( .D(int_data_y_4__1__2_), .CK(
        pe_1_3_1_net5592), .RN(pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_v[6]) );
  DFFR_X1 pe_1_3_1_int_q_reg_v_reg_4__3_ ( .D(int_data_y_4__1__3_), .CK(
        pe_1_3_1_net5592), .RN(pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_v[7]) );
  DFFR_X1 pe_1_3_1_int_q_reg_v_reg_5__0_ ( .D(int_data_y_4__1__0_), .CK(
        pe_1_3_1_net5597), .RN(pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_v[0]) );
  DFFR_X1 pe_1_3_1_int_q_reg_v_reg_5__1_ ( .D(int_data_y_4__1__1_), .CK(
        pe_1_3_1_net5597), .RN(pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_v[1]) );
  DFFR_X1 pe_1_3_1_int_q_reg_v_reg_5__2_ ( .D(int_data_y_4__1__2_), .CK(
        pe_1_3_1_net5597), .RN(pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_v[2]) );
  DFFR_X1 pe_1_3_1_int_q_reg_v_reg_5__3_ ( .D(int_data_y_4__1__3_), .CK(
        pe_1_3_1_net5597), .RN(pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_3_1_int_q_reg_h_reg_0__0_ ( .D(int_data_x_3__2__0_), .SI(
        int_data_y_4__1__0_), .SE(pe_1_3_1_n62), .CK(pe_1_3_1_net5541), .RN(
        pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_3_1_int_q_reg_h_reg_0__1_ ( .D(int_data_x_3__2__1_), .SI(
        int_data_y_4__1__1_), .SE(pe_1_3_1_n62), .CK(pe_1_3_1_net5541), .RN(
        pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_3_1_int_q_reg_h_reg_0__2_ ( .D(int_data_x_3__2__2_), .SI(
        int_data_y_4__1__2_), .SE(pe_1_3_1_n62), .CK(pe_1_3_1_net5541), .RN(
        pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_3_1_int_q_reg_h_reg_0__3_ ( .D(int_data_x_3__2__3_), .SI(
        int_data_y_4__1__3_), .SE(pe_1_3_1_n62), .CK(pe_1_3_1_net5541), .RN(
        pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_3_1_int_q_reg_h_reg_1__0_ ( .D(int_data_x_3__2__0_), .SI(
        int_data_y_4__1__0_), .SE(pe_1_3_1_n62), .CK(pe_1_3_1_net5547), .RN(
        pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_3_1_int_q_reg_h_reg_1__1_ ( .D(int_data_x_3__2__1_), .SI(
        int_data_y_4__1__1_), .SE(pe_1_3_1_n62), .CK(pe_1_3_1_net5547), .RN(
        pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_3_1_int_q_reg_h_reg_1__2_ ( .D(int_data_x_3__2__2_), .SI(
        int_data_y_4__1__2_), .SE(pe_1_3_1_n62), .CK(pe_1_3_1_net5547), .RN(
        pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_3_1_int_q_reg_h_reg_1__3_ ( .D(int_data_x_3__2__3_), .SI(
        int_data_y_4__1__3_), .SE(pe_1_3_1_n62), .CK(pe_1_3_1_net5547), .RN(
        pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_3_1_int_q_reg_h_reg_2__0_ ( .D(int_data_x_3__2__0_), .SI(
        int_data_y_4__1__0_), .SE(pe_1_3_1_n62), .CK(pe_1_3_1_net5552), .RN(
        pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_3_1_int_q_reg_h_reg_2__1_ ( .D(int_data_x_3__2__1_), .SI(
        int_data_y_4__1__1_), .SE(pe_1_3_1_n62), .CK(pe_1_3_1_net5552), .RN(
        pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_3_1_int_q_reg_h_reg_2__2_ ( .D(int_data_x_3__2__2_), .SI(
        int_data_y_4__1__2_), .SE(pe_1_3_1_n62), .CK(pe_1_3_1_net5552), .RN(
        pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_3_1_int_q_reg_h_reg_2__3_ ( .D(int_data_x_3__2__3_), .SI(
        int_data_y_4__1__3_), .SE(pe_1_3_1_n62), .CK(pe_1_3_1_net5552), .RN(
        pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_3_1_int_q_reg_h_reg_3__0_ ( .D(int_data_x_3__2__0_), .SI(
        int_data_y_4__1__0_), .SE(pe_1_3_1_n62), .CK(pe_1_3_1_net5557), .RN(
        pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_3_1_int_q_reg_h_reg_3__1_ ( .D(int_data_x_3__2__1_), .SI(
        int_data_y_4__1__1_), .SE(pe_1_3_1_n62), .CK(pe_1_3_1_net5557), .RN(
        pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_3_1_int_q_reg_h_reg_3__2_ ( .D(int_data_x_3__2__2_), .SI(
        int_data_y_4__1__2_), .SE(pe_1_3_1_n62), .CK(pe_1_3_1_net5557), .RN(
        pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_3_1_int_q_reg_h_reg_3__3_ ( .D(int_data_x_3__2__3_), .SI(
        int_data_y_4__1__3_), .SE(pe_1_3_1_n62), .CK(pe_1_3_1_net5557), .RN(
        pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_3_1_int_q_reg_h_reg_4__0_ ( .D(int_data_x_3__2__0_), .SI(
        int_data_y_4__1__0_), .SE(pe_1_3_1_n63), .CK(pe_1_3_1_net5562), .RN(
        pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_3_1_int_q_reg_h_reg_4__1_ ( .D(int_data_x_3__2__1_), .SI(
        int_data_y_4__1__1_), .SE(pe_1_3_1_n63), .CK(pe_1_3_1_net5562), .RN(
        pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_3_1_int_q_reg_h_reg_4__2_ ( .D(int_data_x_3__2__2_), .SI(
        int_data_y_4__1__2_), .SE(pe_1_3_1_n63), .CK(pe_1_3_1_net5562), .RN(
        pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_3_1_int_q_reg_h_reg_4__3_ ( .D(int_data_x_3__2__3_), .SI(
        int_data_y_4__1__3_), .SE(pe_1_3_1_n63), .CK(pe_1_3_1_net5562), .RN(
        pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_3_1_int_q_reg_h_reg_5__0_ ( .D(int_data_x_3__2__0_), .SI(
        int_data_y_4__1__0_), .SE(pe_1_3_1_n63), .CK(pe_1_3_1_net5567), .RN(
        pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_3_1_int_q_reg_h_reg_5__1_ ( .D(int_data_x_3__2__1_), .SI(
        int_data_y_4__1__1_), .SE(pe_1_3_1_n63), .CK(pe_1_3_1_net5567), .RN(
        pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_3_1_int_q_reg_h_reg_5__2_ ( .D(int_data_x_3__2__2_), .SI(
        int_data_y_4__1__2_), .SE(pe_1_3_1_n63), .CK(pe_1_3_1_net5567), .RN(
        pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_3_1_int_q_reg_h_reg_5__3_ ( .D(int_data_x_3__2__3_), .SI(
        int_data_y_4__1__3_), .SE(pe_1_3_1_n63), .CK(pe_1_3_1_net5567), .RN(
        pe_1_3_1_n68), .Q(pe_1_3_1_int_q_reg_h[3]) );
  FA_X1 pe_1_3_1_sub_81_U2_7 ( .A(int_data_res_3__1__7_), .B(pe_1_3_1_n72), 
        .CI(pe_1_3_1_sub_81_carry[7]), .S(pe_1_3_1_N77) );
  FA_X1 pe_1_3_1_sub_81_U2_6 ( .A(int_data_res_3__1__6_), .B(pe_1_3_1_n72), 
        .CI(pe_1_3_1_sub_81_carry[6]), .CO(pe_1_3_1_sub_81_carry[7]), .S(
        pe_1_3_1_N76) );
  FA_X1 pe_1_3_1_sub_81_U2_5 ( .A(int_data_res_3__1__5_), .B(pe_1_3_1_n72), 
        .CI(pe_1_3_1_sub_81_carry[5]), .CO(pe_1_3_1_sub_81_carry[6]), .S(
        pe_1_3_1_N75) );
  FA_X1 pe_1_3_1_sub_81_U2_4 ( .A(int_data_res_3__1__4_), .B(pe_1_3_1_n72), 
        .CI(pe_1_3_1_sub_81_carry[4]), .CO(pe_1_3_1_sub_81_carry[5]), .S(
        pe_1_3_1_N74) );
  FA_X1 pe_1_3_1_sub_81_U2_3 ( .A(int_data_res_3__1__3_), .B(pe_1_3_1_n72), 
        .CI(pe_1_3_1_sub_81_carry[3]), .CO(pe_1_3_1_sub_81_carry[4]), .S(
        pe_1_3_1_N73) );
  FA_X1 pe_1_3_1_sub_81_U2_2 ( .A(int_data_res_3__1__2_), .B(pe_1_3_1_n71), 
        .CI(pe_1_3_1_sub_81_carry[2]), .CO(pe_1_3_1_sub_81_carry[3]), .S(
        pe_1_3_1_N72) );
  FA_X1 pe_1_3_1_sub_81_U2_1 ( .A(int_data_res_3__1__1_), .B(pe_1_3_1_n70), 
        .CI(pe_1_3_1_sub_81_carry[1]), .CO(pe_1_3_1_sub_81_carry[2]), .S(
        pe_1_3_1_N71) );
  FA_X1 pe_1_3_1_add_83_U1_7 ( .A(int_data_res_3__1__7_), .B(
        pe_1_3_1_int_data_3_), .CI(pe_1_3_1_add_83_carry[7]), .S(pe_1_3_1_N85)
         );
  FA_X1 pe_1_3_1_add_83_U1_6 ( .A(int_data_res_3__1__6_), .B(
        pe_1_3_1_int_data_3_), .CI(pe_1_3_1_add_83_carry[6]), .CO(
        pe_1_3_1_add_83_carry[7]), .S(pe_1_3_1_N84) );
  FA_X1 pe_1_3_1_add_83_U1_5 ( .A(int_data_res_3__1__5_), .B(
        pe_1_3_1_int_data_3_), .CI(pe_1_3_1_add_83_carry[5]), .CO(
        pe_1_3_1_add_83_carry[6]), .S(pe_1_3_1_N83) );
  FA_X1 pe_1_3_1_add_83_U1_4 ( .A(int_data_res_3__1__4_), .B(
        pe_1_3_1_int_data_3_), .CI(pe_1_3_1_add_83_carry[4]), .CO(
        pe_1_3_1_add_83_carry[5]), .S(pe_1_3_1_N82) );
  FA_X1 pe_1_3_1_add_83_U1_3 ( .A(int_data_res_3__1__3_), .B(
        pe_1_3_1_int_data_3_), .CI(pe_1_3_1_add_83_carry[3]), .CO(
        pe_1_3_1_add_83_carry[4]), .S(pe_1_3_1_N81) );
  FA_X1 pe_1_3_1_add_83_U1_2 ( .A(int_data_res_3__1__2_), .B(
        pe_1_3_1_int_data_2_), .CI(pe_1_3_1_add_83_carry[2]), .CO(
        pe_1_3_1_add_83_carry[3]), .S(pe_1_3_1_N80) );
  FA_X1 pe_1_3_1_add_83_U1_1 ( .A(int_data_res_3__1__1_), .B(
        pe_1_3_1_int_data_1_), .CI(pe_1_3_1_n2), .CO(pe_1_3_1_add_83_carry[2]), 
        .S(pe_1_3_1_N79) );
  NAND3_X1 pe_1_3_1_U56 ( .A1(n33), .A2(pe_1_3_1_n43), .A3(n39), .ZN(
        pe_1_3_1_n40) );
  NAND3_X1 pe_1_3_1_U55 ( .A1(pe_1_3_1_n43), .A2(pe_1_3_1_n59), .A3(n39), .ZN(
        pe_1_3_1_n39) );
  NAND3_X1 pe_1_3_1_U54 ( .A1(pe_1_3_1_n43), .A2(pe_1_3_1_n60), .A3(n33), .ZN(
        pe_1_3_1_n38) );
  NAND3_X1 pe_1_3_1_U53 ( .A1(pe_1_3_1_n59), .A2(pe_1_3_1_n60), .A3(
        pe_1_3_1_n43), .ZN(pe_1_3_1_n37) );
  DFFR_X1 pe_1_3_1_int_q_acc_reg_6_ ( .D(pe_1_3_1_n74), .CK(pe_1_3_1_net5602), 
        .RN(pe_1_3_1_n67), .Q(int_data_res_3__1__6_) );
  DFFR_X1 pe_1_3_1_int_q_acc_reg_5_ ( .D(pe_1_3_1_n75), .CK(pe_1_3_1_net5602), 
        .RN(pe_1_3_1_n67), .Q(int_data_res_3__1__5_) );
  DFFR_X1 pe_1_3_1_int_q_acc_reg_4_ ( .D(pe_1_3_1_n76), .CK(pe_1_3_1_net5602), 
        .RN(pe_1_3_1_n67), .Q(int_data_res_3__1__4_) );
  DFFR_X1 pe_1_3_1_int_q_acc_reg_3_ ( .D(pe_1_3_1_n77), .CK(pe_1_3_1_net5602), 
        .RN(pe_1_3_1_n67), .Q(int_data_res_3__1__3_) );
  DFFR_X1 pe_1_3_1_int_q_acc_reg_2_ ( .D(pe_1_3_1_n78), .CK(pe_1_3_1_net5602), 
        .RN(pe_1_3_1_n67), .Q(int_data_res_3__1__2_) );
  DFFR_X1 pe_1_3_1_int_q_acc_reg_1_ ( .D(pe_1_3_1_n79), .CK(pe_1_3_1_net5602), 
        .RN(pe_1_3_1_n67), .Q(int_data_res_3__1__1_) );
  DFFR_X1 pe_1_3_1_int_q_acc_reg_7_ ( .D(pe_1_3_1_n73), .CK(pe_1_3_1_net5602), 
        .RN(pe_1_3_1_n67), .Q(int_data_res_3__1__7_) );
  CLKGATETST_X1 pe_1_3_1_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_3_1_n84), .SE(1'b0), .GCK(pe_1_3_1_net5541) );
  CLKGATETST_X1 pe_1_3_1_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_3_1_n83), .SE(1'b0), .GCK(pe_1_3_1_net5547) );
  CLKGATETST_X1 pe_1_3_1_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_3_1_n82), .SE(1'b0), .GCK(pe_1_3_1_net5552) );
  CLKGATETST_X1 pe_1_3_1_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_3_1_n81), .SE(1'b0), .GCK(pe_1_3_1_net5557) );
  CLKGATETST_X1 pe_1_3_1_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_3_1_n86), .SE(1'b0), .GCK(pe_1_3_1_net5562) );
  CLKGATETST_X1 pe_1_3_1_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_3_1_n85), .SE(1'b0), .GCK(pe_1_3_1_net5567) );
  CLKGATETST_X1 pe_1_3_1_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_3_1_N64), .SE(1'b0), .GCK(pe_1_3_1_net5572) );
  CLKGATETST_X1 pe_1_3_1_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_3_1_N63), .SE(1'b0), .GCK(pe_1_3_1_net5577) );
  CLKGATETST_X1 pe_1_3_1_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_3_1_N62), .SE(1'b0), .GCK(pe_1_3_1_net5582) );
  CLKGATETST_X1 pe_1_3_1_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_3_1_N61), .SE(1'b0), .GCK(pe_1_3_1_net5587) );
  CLKGATETST_X1 pe_1_3_1_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_3_1_N60), .SE(1'b0), .GCK(pe_1_3_1_net5592) );
  CLKGATETST_X1 pe_1_3_1_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_3_1_N59), .SE(1'b0), .GCK(pe_1_3_1_net5597) );
  CLKGATETST_X1 pe_1_3_1_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_3_1_N90), .SE(1'b0), .GCK(pe_1_3_1_net5602) );
  CLKBUF_X1 pe_1_3_2_U109 ( .A(pe_1_3_2_n69), .Z(pe_1_3_2_n68) );
  INV_X1 pe_1_3_2_U108 ( .A(n75), .ZN(pe_1_3_2_n67) );
  INV_X1 pe_1_3_2_U107 ( .A(n67), .ZN(pe_1_3_2_n66) );
  INV_X1 pe_1_3_2_U106 ( .A(n67), .ZN(pe_1_3_2_n65) );
  INV_X1 pe_1_3_2_U105 ( .A(pe_1_3_2_n66), .ZN(pe_1_3_2_n64) );
  INV_X1 pe_1_3_2_U104 ( .A(pe_1_3_2_n61), .ZN(pe_1_3_2_n60) );
  INV_X1 pe_1_3_2_U103 ( .A(n27), .ZN(pe_1_3_2_n58) );
  INV_X1 pe_1_3_2_U102 ( .A(n19), .ZN(pe_1_3_2_n57) );
  MUX2_X1 pe_1_3_2_U101 ( .A(pe_1_3_2_n54), .B(pe_1_3_2_n51), .S(n48), .Z(
        int_data_x_3__2__3_) );
  MUX2_X1 pe_1_3_2_U100 ( .A(pe_1_3_2_n53), .B(pe_1_3_2_n52), .S(pe_1_3_2_n60), 
        .Z(pe_1_3_2_n54) );
  MUX2_X1 pe_1_3_2_U99 ( .A(pe_1_3_2_int_q_reg_h[23]), .B(
        pe_1_3_2_int_q_reg_h[19]), .S(pe_1_3_2_n56), .Z(pe_1_3_2_n53) );
  MUX2_X1 pe_1_3_2_U98 ( .A(pe_1_3_2_int_q_reg_h[15]), .B(
        pe_1_3_2_int_q_reg_h[11]), .S(pe_1_3_2_n56), .Z(pe_1_3_2_n52) );
  MUX2_X1 pe_1_3_2_U97 ( .A(pe_1_3_2_int_q_reg_h[7]), .B(
        pe_1_3_2_int_q_reg_h[3]), .S(pe_1_3_2_n56), .Z(pe_1_3_2_n51) );
  MUX2_X1 pe_1_3_2_U96 ( .A(pe_1_3_2_n50), .B(pe_1_3_2_n47), .S(n48), .Z(
        int_data_x_3__2__2_) );
  MUX2_X1 pe_1_3_2_U95 ( .A(pe_1_3_2_n49), .B(pe_1_3_2_n48), .S(pe_1_3_2_n60), 
        .Z(pe_1_3_2_n50) );
  MUX2_X1 pe_1_3_2_U94 ( .A(pe_1_3_2_int_q_reg_h[22]), .B(
        pe_1_3_2_int_q_reg_h[18]), .S(pe_1_3_2_n56), .Z(pe_1_3_2_n49) );
  MUX2_X1 pe_1_3_2_U93 ( .A(pe_1_3_2_int_q_reg_h[14]), .B(
        pe_1_3_2_int_q_reg_h[10]), .S(pe_1_3_2_n56), .Z(pe_1_3_2_n48) );
  MUX2_X1 pe_1_3_2_U92 ( .A(pe_1_3_2_int_q_reg_h[6]), .B(
        pe_1_3_2_int_q_reg_h[2]), .S(pe_1_3_2_n56), .Z(pe_1_3_2_n47) );
  MUX2_X1 pe_1_3_2_U91 ( .A(pe_1_3_2_n46), .B(pe_1_3_2_n24), .S(n48), .Z(
        int_data_x_3__2__1_) );
  MUX2_X1 pe_1_3_2_U90 ( .A(pe_1_3_2_n45), .B(pe_1_3_2_n25), .S(pe_1_3_2_n60), 
        .Z(pe_1_3_2_n46) );
  MUX2_X1 pe_1_3_2_U89 ( .A(pe_1_3_2_int_q_reg_h[21]), .B(
        pe_1_3_2_int_q_reg_h[17]), .S(pe_1_3_2_n56), .Z(pe_1_3_2_n45) );
  MUX2_X1 pe_1_3_2_U88 ( .A(pe_1_3_2_int_q_reg_h[13]), .B(
        pe_1_3_2_int_q_reg_h[9]), .S(pe_1_3_2_n56), .Z(pe_1_3_2_n25) );
  MUX2_X1 pe_1_3_2_U87 ( .A(pe_1_3_2_int_q_reg_h[5]), .B(
        pe_1_3_2_int_q_reg_h[1]), .S(pe_1_3_2_n56), .Z(pe_1_3_2_n24) );
  MUX2_X1 pe_1_3_2_U86 ( .A(pe_1_3_2_n23), .B(pe_1_3_2_n20), .S(n48), .Z(
        int_data_x_3__2__0_) );
  MUX2_X1 pe_1_3_2_U85 ( .A(pe_1_3_2_n22), .B(pe_1_3_2_n21), .S(pe_1_3_2_n60), 
        .Z(pe_1_3_2_n23) );
  MUX2_X1 pe_1_3_2_U84 ( .A(pe_1_3_2_int_q_reg_h[20]), .B(
        pe_1_3_2_int_q_reg_h[16]), .S(pe_1_3_2_n56), .Z(pe_1_3_2_n22) );
  MUX2_X1 pe_1_3_2_U83 ( .A(pe_1_3_2_int_q_reg_h[12]), .B(
        pe_1_3_2_int_q_reg_h[8]), .S(pe_1_3_2_n56), .Z(pe_1_3_2_n21) );
  MUX2_X1 pe_1_3_2_U82 ( .A(pe_1_3_2_int_q_reg_h[4]), .B(
        pe_1_3_2_int_q_reg_h[0]), .S(pe_1_3_2_n56), .Z(pe_1_3_2_n20) );
  MUX2_X1 pe_1_3_2_U81 ( .A(pe_1_3_2_n19), .B(pe_1_3_2_n16), .S(n48), .Z(
        int_data_y_3__2__3_) );
  MUX2_X1 pe_1_3_2_U80 ( .A(pe_1_3_2_n18), .B(pe_1_3_2_n17), .S(pe_1_3_2_n60), 
        .Z(pe_1_3_2_n19) );
  MUX2_X1 pe_1_3_2_U79 ( .A(pe_1_3_2_int_q_reg_v[23]), .B(
        pe_1_3_2_int_q_reg_v[19]), .S(pe_1_3_2_n55), .Z(pe_1_3_2_n18) );
  MUX2_X1 pe_1_3_2_U78 ( .A(pe_1_3_2_int_q_reg_v[15]), .B(
        pe_1_3_2_int_q_reg_v[11]), .S(pe_1_3_2_n55), .Z(pe_1_3_2_n17) );
  MUX2_X1 pe_1_3_2_U77 ( .A(pe_1_3_2_int_q_reg_v[7]), .B(
        pe_1_3_2_int_q_reg_v[3]), .S(pe_1_3_2_n55), .Z(pe_1_3_2_n16) );
  MUX2_X1 pe_1_3_2_U76 ( .A(pe_1_3_2_n15), .B(pe_1_3_2_n12), .S(n48), .Z(
        int_data_y_3__2__2_) );
  MUX2_X1 pe_1_3_2_U75 ( .A(pe_1_3_2_n14), .B(pe_1_3_2_n13), .S(pe_1_3_2_n60), 
        .Z(pe_1_3_2_n15) );
  MUX2_X1 pe_1_3_2_U74 ( .A(pe_1_3_2_int_q_reg_v[22]), .B(
        pe_1_3_2_int_q_reg_v[18]), .S(pe_1_3_2_n55), .Z(pe_1_3_2_n14) );
  MUX2_X1 pe_1_3_2_U73 ( .A(pe_1_3_2_int_q_reg_v[14]), .B(
        pe_1_3_2_int_q_reg_v[10]), .S(pe_1_3_2_n55), .Z(pe_1_3_2_n13) );
  MUX2_X1 pe_1_3_2_U72 ( .A(pe_1_3_2_int_q_reg_v[6]), .B(
        pe_1_3_2_int_q_reg_v[2]), .S(pe_1_3_2_n55), .Z(pe_1_3_2_n12) );
  MUX2_X1 pe_1_3_2_U71 ( .A(pe_1_3_2_n11), .B(pe_1_3_2_n8), .S(n48), .Z(
        int_data_y_3__2__1_) );
  MUX2_X1 pe_1_3_2_U70 ( .A(pe_1_3_2_n10), .B(pe_1_3_2_n9), .S(pe_1_3_2_n60), 
        .Z(pe_1_3_2_n11) );
  MUX2_X1 pe_1_3_2_U69 ( .A(pe_1_3_2_int_q_reg_v[21]), .B(
        pe_1_3_2_int_q_reg_v[17]), .S(pe_1_3_2_n55), .Z(pe_1_3_2_n10) );
  MUX2_X1 pe_1_3_2_U68 ( .A(pe_1_3_2_int_q_reg_v[13]), .B(
        pe_1_3_2_int_q_reg_v[9]), .S(pe_1_3_2_n55), .Z(pe_1_3_2_n9) );
  MUX2_X1 pe_1_3_2_U67 ( .A(pe_1_3_2_int_q_reg_v[5]), .B(
        pe_1_3_2_int_q_reg_v[1]), .S(pe_1_3_2_n55), .Z(pe_1_3_2_n8) );
  MUX2_X1 pe_1_3_2_U66 ( .A(pe_1_3_2_n7), .B(pe_1_3_2_n4), .S(n48), .Z(
        int_data_y_3__2__0_) );
  MUX2_X1 pe_1_3_2_U65 ( .A(pe_1_3_2_n6), .B(pe_1_3_2_n5), .S(pe_1_3_2_n60), 
        .Z(pe_1_3_2_n7) );
  MUX2_X1 pe_1_3_2_U64 ( .A(pe_1_3_2_int_q_reg_v[20]), .B(
        pe_1_3_2_int_q_reg_v[16]), .S(pe_1_3_2_n55), .Z(pe_1_3_2_n6) );
  MUX2_X1 pe_1_3_2_U63 ( .A(pe_1_3_2_int_q_reg_v[12]), .B(
        pe_1_3_2_int_q_reg_v[8]), .S(pe_1_3_2_n55), .Z(pe_1_3_2_n5) );
  MUX2_X1 pe_1_3_2_U62 ( .A(pe_1_3_2_int_q_reg_v[4]), .B(
        pe_1_3_2_int_q_reg_v[0]), .S(pe_1_3_2_n55), .Z(pe_1_3_2_n4) );
  AOI222_X1 pe_1_3_2_U61 ( .A1(int_data_res_4__2__2_), .A2(pe_1_3_2_n62), .B1(
        pe_1_3_2_N80), .B2(pe_1_3_2_n27), .C1(pe_1_3_2_N72), .C2(pe_1_3_2_n28), 
        .ZN(pe_1_3_2_n33) );
  INV_X1 pe_1_3_2_U60 ( .A(pe_1_3_2_n33), .ZN(pe_1_3_2_n79) );
  AOI222_X1 pe_1_3_2_U59 ( .A1(int_data_res_4__2__6_), .A2(pe_1_3_2_n62), .B1(
        pe_1_3_2_N84), .B2(pe_1_3_2_n27), .C1(pe_1_3_2_N76), .C2(pe_1_3_2_n28), 
        .ZN(pe_1_3_2_n29) );
  INV_X1 pe_1_3_2_U58 ( .A(pe_1_3_2_n29), .ZN(pe_1_3_2_n75) );
  XNOR2_X1 pe_1_3_2_U57 ( .A(pe_1_3_2_n70), .B(int_data_res_3__2__0_), .ZN(
        pe_1_3_2_N70) );
  AOI222_X1 pe_1_3_2_U52 ( .A1(int_data_res_4__2__0_), .A2(pe_1_3_2_n62), .B1(
        pe_1_3_2_n1), .B2(pe_1_3_2_n27), .C1(pe_1_3_2_N70), .C2(pe_1_3_2_n28), 
        .ZN(pe_1_3_2_n35) );
  INV_X1 pe_1_3_2_U51 ( .A(pe_1_3_2_n35), .ZN(pe_1_3_2_n81) );
  AOI222_X1 pe_1_3_2_U50 ( .A1(int_data_res_4__2__1_), .A2(pe_1_3_2_n62), .B1(
        pe_1_3_2_N79), .B2(pe_1_3_2_n27), .C1(pe_1_3_2_N71), .C2(pe_1_3_2_n28), 
        .ZN(pe_1_3_2_n34) );
  INV_X1 pe_1_3_2_U49 ( .A(pe_1_3_2_n34), .ZN(pe_1_3_2_n80) );
  AOI222_X1 pe_1_3_2_U48 ( .A1(int_data_res_4__2__3_), .A2(pe_1_3_2_n62), .B1(
        pe_1_3_2_N81), .B2(pe_1_3_2_n27), .C1(pe_1_3_2_N73), .C2(pe_1_3_2_n28), 
        .ZN(pe_1_3_2_n32) );
  INV_X1 pe_1_3_2_U47 ( .A(pe_1_3_2_n32), .ZN(pe_1_3_2_n78) );
  AOI222_X1 pe_1_3_2_U46 ( .A1(int_data_res_4__2__4_), .A2(pe_1_3_2_n62), .B1(
        pe_1_3_2_N82), .B2(pe_1_3_2_n27), .C1(pe_1_3_2_N74), .C2(pe_1_3_2_n28), 
        .ZN(pe_1_3_2_n31) );
  INV_X1 pe_1_3_2_U45 ( .A(pe_1_3_2_n31), .ZN(pe_1_3_2_n77) );
  AOI222_X1 pe_1_3_2_U44 ( .A1(int_data_res_4__2__5_), .A2(pe_1_3_2_n62), .B1(
        pe_1_3_2_N83), .B2(pe_1_3_2_n27), .C1(pe_1_3_2_N75), .C2(pe_1_3_2_n28), 
        .ZN(pe_1_3_2_n30) );
  INV_X1 pe_1_3_2_U43 ( .A(pe_1_3_2_n30), .ZN(pe_1_3_2_n76) );
  NAND2_X1 pe_1_3_2_U42 ( .A1(pe_1_3_2_int_data_0_), .A2(pe_1_3_2_n3), .ZN(
        pe_1_3_2_sub_81_carry[1]) );
  INV_X1 pe_1_3_2_U41 ( .A(pe_1_3_2_int_data_1_), .ZN(pe_1_3_2_n71) );
  INV_X1 pe_1_3_2_U40 ( .A(pe_1_3_2_int_data_2_), .ZN(pe_1_3_2_n72) );
  AND2_X1 pe_1_3_2_U39 ( .A1(pe_1_3_2_int_data_0_), .A2(int_data_res_3__2__0_), 
        .ZN(pe_1_3_2_n2) );
  AOI222_X1 pe_1_3_2_U38 ( .A1(pe_1_3_2_n62), .A2(int_data_res_4__2__7_), .B1(
        pe_1_3_2_N85), .B2(pe_1_3_2_n27), .C1(pe_1_3_2_N77), .C2(pe_1_3_2_n28), 
        .ZN(pe_1_3_2_n26) );
  INV_X1 pe_1_3_2_U37 ( .A(pe_1_3_2_n26), .ZN(pe_1_3_2_n74) );
  NOR3_X1 pe_1_3_2_U36 ( .A1(pe_1_3_2_n58), .A2(pe_1_3_2_n63), .A3(int_ckg[37]), .ZN(pe_1_3_2_n36) );
  OR2_X1 pe_1_3_2_U35 ( .A1(pe_1_3_2_n36), .A2(pe_1_3_2_n62), .ZN(pe_1_3_2_N90) );
  INV_X1 pe_1_3_2_U34 ( .A(n39), .ZN(pe_1_3_2_n61) );
  AND2_X1 pe_1_3_2_U33 ( .A1(int_data_x_3__2__2_), .A2(n27), .ZN(
        pe_1_3_2_int_data_2_) );
  AND2_X1 pe_1_3_2_U32 ( .A1(int_data_x_3__2__1_), .A2(n27), .ZN(
        pe_1_3_2_int_data_1_) );
  AND2_X1 pe_1_3_2_U31 ( .A1(int_data_x_3__2__3_), .A2(n27), .ZN(
        pe_1_3_2_int_data_3_) );
  BUF_X1 pe_1_3_2_U30 ( .A(n61), .Z(pe_1_3_2_n62) );
  INV_X1 pe_1_3_2_U29 ( .A(n33), .ZN(pe_1_3_2_n59) );
  AND2_X1 pe_1_3_2_U28 ( .A1(int_data_x_3__2__0_), .A2(n27), .ZN(
        pe_1_3_2_int_data_0_) );
  NAND2_X1 pe_1_3_2_U27 ( .A1(pe_1_3_2_n44), .A2(pe_1_3_2_n59), .ZN(
        pe_1_3_2_n41) );
  AND3_X1 pe_1_3_2_U26 ( .A1(n75), .A2(pe_1_3_2_n61), .A3(n48), .ZN(
        pe_1_3_2_n44) );
  INV_X1 pe_1_3_2_U25 ( .A(pe_1_3_2_int_data_3_), .ZN(pe_1_3_2_n73) );
  NOR2_X1 pe_1_3_2_U24 ( .A1(pe_1_3_2_n67), .A2(n48), .ZN(pe_1_3_2_n43) );
  NOR2_X1 pe_1_3_2_U23 ( .A1(pe_1_3_2_n57), .A2(pe_1_3_2_n62), .ZN(
        pe_1_3_2_n28) );
  NOR2_X1 pe_1_3_2_U22 ( .A1(n19), .A2(pe_1_3_2_n62), .ZN(pe_1_3_2_n27) );
  INV_X1 pe_1_3_2_U21 ( .A(pe_1_3_2_int_data_0_), .ZN(pe_1_3_2_n70) );
  INV_X1 pe_1_3_2_U20 ( .A(pe_1_3_2_n41), .ZN(pe_1_3_2_n87) );
  INV_X1 pe_1_3_2_U19 ( .A(pe_1_3_2_n37), .ZN(pe_1_3_2_n85) );
  INV_X1 pe_1_3_2_U18 ( .A(pe_1_3_2_n38), .ZN(pe_1_3_2_n84) );
  INV_X1 pe_1_3_2_U17 ( .A(pe_1_3_2_n39), .ZN(pe_1_3_2_n83) );
  NOR2_X1 pe_1_3_2_U16 ( .A1(pe_1_3_2_n65), .A2(pe_1_3_2_n42), .ZN(
        pe_1_3_2_N59) );
  NOR2_X1 pe_1_3_2_U15 ( .A1(pe_1_3_2_n65), .A2(pe_1_3_2_n41), .ZN(
        pe_1_3_2_N60) );
  NOR2_X1 pe_1_3_2_U14 ( .A1(pe_1_3_2_n65), .A2(pe_1_3_2_n38), .ZN(
        pe_1_3_2_N63) );
  NOR2_X1 pe_1_3_2_U13 ( .A1(pe_1_3_2_n65), .A2(pe_1_3_2_n40), .ZN(
        pe_1_3_2_N61) );
  NOR2_X1 pe_1_3_2_U12 ( .A1(pe_1_3_2_n65), .A2(pe_1_3_2_n39), .ZN(
        pe_1_3_2_N62) );
  NOR2_X1 pe_1_3_2_U11 ( .A1(pe_1_3_2_n37), .A2(pe_1_3_2_n65), .ZN(
        pe_1_3_2_N64) );
  NAND2_X1 pe_1_3_2_U10 ( .A1(pe_1_3_2_n44), .A2(n33), .ZN(pe_1_3_2_n42) );
  BUF_X1 pe_1_3_2_U9 ( .A(n33), .Z(pe_1_3_2_n55) );
  INV_X1 pe_1_3_2_U8 ( .A(pe_1_3_2_n66), .ZN(pe_1_3_2_n63) );
  BUF_X1 pe_1_3_2_U7 ( .A(n33), .Z(pe_1_3_2_n56) );
  INV_X1 pe_1_3_2_U6 ( .A(pe_1_3_2_n42), .ZN(pe_1_3_2_n86) );
  INV_X1 pe_1_3_2_U5 ( .A(pe_1_3_2_n40), .ZN(pe_1_3_2_n82) );
  INV_X2 pe_1_3_2_U4 ( .A(n83), .ZN(pe_1_3_2_n69) );
  XOR2_X1 pe_1_3_2_U3 ( .A(pe_1_3_2_int_data_0_), .B(int_data_res_3__2__0_), 
        .Z(pe_1_3_2_n1) );
  DFFR_X1 pe_1_3_2_int_q_acc_reg_0_ ( .D(pe_1_3_2_n81), .CK(pe_1_3_2_net5524), 
        .RN(pe_1_3_2_n69), .Q(int_data_res_3__2__0_), .QN(pe_1_3_2_n3) );
  DFFR_X1 pe_1_3_2_int_q_reg_v_reg_0__0_ ( .D(int_data_y_4__2__0_), .CK(
        pe_1_3_2_net5494), .RN(pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_v[20]) );
  DFFR_X1 pe_1_3_2_int_q_reg_v_reg_0__1_ ( .D(int_data_y_4__2__1_), .CK(
        pe_1_3_2_net5494), .RN(pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_v[21]) );
  DFFR_X1 pe_1_3_2_int_q_reg_v_reg_0__2_ ( .D(int_data_y_4__2__2_), .CK(
        pe_1_3_2_net5494), .RN(pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_v[22]) );
  DFFR_X1 pe_1_3_2_int_q_reg_v_reg_0__3_ ( .D(int_data_y_4__2__3_), .CK(
        pe_1_3_2_net5494), .RN(pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_v[23]) );
  DFFR_X1 pe_1_3_2_int_q_reg_v_reg_1__0_ ( .D(int_data_y_4__2__0_), .CK(
        pe_1_3_2_net5499), .RN(pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_v[16]) );
  DFFR_X1 pe_1_3_2_int_q_reg_v_reg_1__1_ ( .D(int_data_y_4__2__1_), .CK(
        pe_1_3_2_net5499), .RN(pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_v[17]) );
  DFFR_X1 pe_1_3_2_int_q_reg_v_reg_1__2_ ( .D(int_data_y_4__2__2_), .CK(
        pe_1_3_2_net5499), .RN(pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_v[18]) );
  DFFR_X1 pe_1_3_2_int_q_reg_v_reg_1__3_ ( .D(int_data_y_4__2__3_), .CK(
        pe_1_3_2_net5499), .RN(pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_v[19]) );
  DFFR_X1 pe_1_3_2_int_q_reg_v_reg_2__0_ ( .D(int_data_y_4__2__0_), .CK(
        pe_1_3_2_net5504), .RN(pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_v[12]) );
  DFFR_X1 pe_1_3_2_int_q_reg_v_reg_2__1_ ( .D(int_data_y_4__2__1_), .CK(
        pe_1_3_2_net5504), .RN(pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_v[13]) );
  DFFR_X1 pe_1_3_2_int_q_reg_v_reg_2__2_ ( .D(int_data_y_4__2__2_), .CK(
        pe_1_3_2_net5504), .RN(pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_v[14]) );
  DFFR_X1 pe_1_3_2_int_q_reg_v_reg_2__3_ ( .D(int_data_y_4__2__3_), .CK(
        pe_1_3_2_net5504), .RN(pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_v[15]) );
  DFFR_X1 pe_1_3_2_int_q_reg_v_reg_3__0_ ( .D(int_data_y_4__2__0_), .CK(
        pe_1_3_2_net5509), .RN(pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_v[8]) );
  DFFR_X1 pe_1_3_2_int_q_reg_v_reg_3__1_ ( .D(int_data_y_4__2__1_), .CK(
        pe_1_3_2_net5509), .RN(pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_v[9]) );
  DFFR_X1 pe_1_3_2_int_q_reg_v_reg_3__2_ ( .D(int_data_y_4__2__2_), .CK(
        pe_1_3_2_net5509), .RN(pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_v[10]) );
  DFFR_X1 pe_1_3_2_int_q_reg_v_reg_3__3_ ( .D(int_data_y_4__2__3_), .CK(
        pe_1_3_2_net5509), .RN(pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_v[11]) );
  DFFR_X1 pe_1_3_2_int_q_reg_v_reg_4__0_ ( .D(int_data_y_4__2__0_), .CK(
        pe_1_3_2_net5514), .RN(pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_v[4]) );
  DFFR_X1 pe_1_3_2_int_q_reg_v_reg_4__1_ ( .D(int_data_y_4__2__1_), .CK(
        pe_1_3_2_net5514), .RN(pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_v[5]) );
  DFFR_X1 pe_1_3_2_int_q_reg_v_reg_4__2_ ( .D(int_data_y_4__2__2_), .CK(
        pe_1_3_2_net5514), .RN(pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_v[6]) );
  DFFR_X1 pe_1_3_2_int_q_reg_v_reg_4__3_ ( .D(int_data_y_4__2__3_), .CK(
        pe_1_3_2_net5514), .RN(pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_v[7]) );
  DFFR_X1 pe_1_3_2_int_q_reg_v_reg_5__0_ ( .D(int_data_y_4__2__0_), .CK(
        pe_1_3_2_net5519), .RN(pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_v[0]) );
  DFFR_X1 pe_1_3_2_int_q_reg_v_reg_5__1_ ( .D(int_data_y_4__2__1_), .CK(
        pe_1_3_2_net5519), .RN(pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_v[1]) );
  DFFR_X1 pe_1_3_2_int_q_reg_v_reg_5__2_ ( .D(int_data_y_4__2__2_), .CK(
        pe_1_3_2_net5519), .RN(pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_v[2]) );
  DFFR_X1 pe_1_3_2_int_q_reg_v_reg_5__3_ ( .D(int_data_y_4__2__3_), .CK(
        pe_1_3_2_net5519), .RN(pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_3_2_int_q_reg_h_reg_0__0_ ( .D(int_data_x_3__3__0_), .SI(
        int_data_y_4__2__0_), .SE(pe_1_3_2_n63), .CK(pe_1_3_2_net5463), .RN(
        pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_3_2_int_q_reg_h_reg_0__1_ ( .D(int_data_x_3__3__1_), .SI(
        int_data_y_4__2__1_), .SE(pe_1_3_2_n63), .CK(pe_1_3_2_net5463), .RN(
        pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_3_2_int_q_reg_h_reg_0__2_ ( .D(int_data_x_3__3__2_), .SI(
        int_data_y_4__2__2_), .SE(pe_1_3_2_n63), .CK(pe_1_3_2_net5463), .RN(
        pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_3_2_int_q_reg_h_reg_0__3_ ( .D(int_data_x_3__3__3_), .SI(
        int_data_y_4__2__3_), .SE(pe_1_3_2_n63), .CK(pe_1_3_2_net5463), .RN(
        pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_3_2_int_q_reg_h_reg_1__0_ ( .D(int_data_x_3__3__0_), .SI(
        int_data_y_4__2__0_), .SE(pe_1_3_2_n63), .CK(pe_1_3_2_net5469), .RN(
        pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_3_2_int_q_reg_h_reg_1__1_ ( .D(int_data_x_3__3__1_), .SI(
        int_data_y_4__2__1_), .SE(pe_1_3_2_n63), .CK(pe_1_3_2_net5469), .RN(
        pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_3_2_int_q_reg_h_reg_1__2_ ( .D(int_data_x_3__3__2_), .SI(
        int_data_y_4__2__2_), .SE(pe_1_3_2_n63), .CK(pe_1_3_2_net5469), .RN(
        pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_3_2_int_q_reg_h_reg_1__3_ ( .D(int_data_x_3__3__3_), .SI(
        int_data_y_4__2__3_), .SE(pe_1_3_2_n63), .CK(pe_1_3_2_net5469), .RN(
        pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_3_2_int_q_reg_h_reg_2__0_ ( .D(int_data_x_3__3__0_), .SI(
        int_data_y_4__2__0_), .SE(pe_1_3_2_n63), .CK(pe_1_3_2_net5474), .RN(
        pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_3_2_int_q_reg_h_reg_2__1_ ( .D(int_data_x_3__3__1_), .SI(
        int_data_y_4__2__1_), .SE(pe_1_3_2_n63), .CK(pe_1_3_2_net5474), .RN(
        pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_3_2_int_q_reg_h_reg_2__2_ ( .D(int_data_x_3__3__2_), .SI(
        int_data_y_4__2__2_), .SE(pe_1_3_2_n63), .CK(pe_1_3_2_net5474), .RN(
        pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_3_2_int_q_reg_h_reg_2__3_ ( .D(int_data_x_3__3__3_), .SI(
        int_data_y_4__2__3_), .SE(pe_1_3_2_n63), .CK(pe_1_3_2_net5474), .RN(
        pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_3_2_int_q_reg_h_reg_3__0_ ( .D(int_data_x_3__3__0_), .SI(
        int_data_y_4__2__0_), .SE(pe_1_3_2_n63), .CK(pe_1_3_2_net5479), .RN(
        pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_3_2_int_q_reg_h_reg_3__1_ ( .D(int_data_x_3__3__1_), .SI(
        int_data_y_4__2__1_), .SE(pe_1_3_2_n63), .CK(pe_1_3_2_net5479), .RN(
        pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_3_2_int_q_reg_h_reg_3__2_ ( .D(int_data_x_3__3__2_), .SI(
        int_data_y_4__2__2_), .SE(pe_1_3_2_n63), .CK(pe_1_3_2_net5479), .RN(
        pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_3_2_int_q_reg_h_reg_3__3_ ( .D(int_data_x_3__3__3_), .SI(
        int_data_y_4__2__3_), .SE(pe_1_3_2_n63), .CK(pe_1_3_2_net5479), .RN(
        pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_3_2_int_q_reg_h_reg_4__0_ ( .D(int_data_x_3__3__0_), .SI(
        int_data_y_4__2__0_), .SE(pe_1_3_2_n64), .CK(pe_1_3_2_net5484), .RN(
        pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_3_2_int_q_reg_h_reg_4__1_ ( .D(int_data_x_3__3__1_), .SI(
        int_data_y_4__2__1_), .SE(pe_1_3_2_n64), .CK(pe_1_3_2_net5484), .RN(
        pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_3_2_int_q_reg_h_reg_4__2_ ( .D(int_data_x_3__3__2_), .SI(
        int_data_y_4__2__2_), .SE(pe_1_3_2_n64), .CK(pe_1_3_2_net5484), .RN(
        pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_3_2_int_q_reg_h_reg_4__3_ ( .D(int_data_x_3__3__3_), .SI(
        int_data_y_4__2__3_), .SE(pe_1_3_2_n64), .CK(pe_1_3_2_net5484), .RN(
        pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_3_2_int_q_reg_h_reg_5__0_ ( .D(int_data_x_3__3__0_), .SI(
        int_data_y_4__2__0_), .SE(pe_1_3_2_n64), .CK(pe_1_3_2_net5489), .RN(
        pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_3_2_int_q_reg_h_reg_5__1_ ( .D(int_data_x_3__3__1_), .SI(
        int_data_y_4__2__1_), .SE(pe_1_3_2_n64), .CK(pe_1_3_2_net5489), .RN(
        pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_3_2_int_q_reg_h_reg_5__2_ ( .D(int_data_x_3__3__2_), .SI(
        int_data_y_4__2__2_), .SE(pe_1_3_2_n64), .CK(pe_1_3_2_net5489), .RN(
        pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_3_2_int_q_reg_h_reg_5__3_ ( .D(int_data_x_3__3__3_), .SI(
        int_data_y_4__2__3_), .SE(pe_1_3_2_n64), .CK(pe_1_3_2_net5489), .RN(
        pe_1_3_2_n69), .Q(pe_1_3_2_int_q_reg_h[3]) );
  FA_X1 pe_1_3_2_sub_81_U2_7 ( .A(int_data_res_3__2__7_), .B(pe_1_3_2_n73), 
        .CI(pe_1_3_2_sub_81_carry[7]), .S(pe_1_3_2_N77) );
  FA_X1 pe_1_3_2_sub_81_U2_6 ( .A(int_data_res_3__2__6_), .B(pe_1_3_2_n73), 
        .CI(pe_1_3_2_sub_81_carry[6]), .CO(pe_1_3_2_sub_81_carry[7]), .S(
        pe_1_3_2_N76) );
  FA_X1 pe_1_3_2_sub_81_U2_5 ( .A(int_data_res_3__2__5_), .B(pe_1_3_2_n73), 
        .CI(pe_1_3_2_sub_81_carry[5]), .CO(pe_1_3_2_sub_81_carry[6]), .S(
        pe_1_3_2_N75) );
  FA_X1 pe_1_3_2_sub_81_U2_4 ( .A(int_data_res_3__2__4_), .B(pe_1_3_2_n73), 
        .CI(pe_1_3_2_sub_81_carry[4]), .CO(pe_1_3_2_sub_81_carry[5]), .S(
        pe_1_3_2_N74) );
  FA_X1 pe_1_3_2_sub_81_U2_3 ( .A(int_data_res_3__2__3_), .B(pe_1_3_2_n73), 
        .CI(pe_1_3_2_sub_81_carry[3]), .CO(pe_1_3_2_sub_81_carry[4]), .S(
        pe_1_3_2_N73) );
  FA_X1 pe_1_3_2_sub_81_U2_2 ( .A(int_data_res_3__2__2_), .B(pe_1_3_2_n72), 
        .CI(pe_1_3_2_sub_81_carry[2]), .CO(pe_1_3_2_sub_81_carry[3]), .S(
        pe_1_3_2_N72) );
  FA_X1 pe_1_3_2_sub_81_U2_1 ( .A(int_data_res_3__2__1_), .B(pe_1_3_2_n71), 
        .CI(pe_1_3_2_sub_81_carry[1]), .CO(pe_1_3_2_sub_81_carry[2]), .S(
        pe_1_3_2_N71) );
  FA_X1 pe_1_3_2_add_83_U1_7 ( .A(int_data_res_3__2__7_), .B(
        pe_1_3_2_int_data_3_), .CI(pe_1_3_2_add_83_carry[7]), .S(pe_1_3_2_N85)
         );
  FA_X1 pe_1_3_2_add_83_U1_6 ( .A(int_data_res_3__2__6_), .B(
        pe_1_3_2_int_data_3_), .CI(pe_1_3_2_add_83_carry[6]), .CO(
        pe_1_3_2_add_83_carry[7]), .S(pe_1_3_2_N84) );
  FA_X1 pe_1_3_2_add_83_U1_5 ( .A(int_data_res_3__2__5_), .B(
        pe_1_3_2_int_data_3_), .CI(pe_1_3_2_add_83_carry[5]), .CO(
        pe_1_3_2_add_83_carry[6]), .S(pe_1_3_2_N83) );
  FA_X1 pe_1_3_2_add_83_U1_4 ( .A(int_data_res_3__2__4_), .B(
        pe_1_3_2_int_data_3_), .CI(pe_1_3_2_add_83_carry[4]), .CO(
        pe_1_3_2_add_83_carry[5]), .S(pe_1_3_2_N82) );
  FA_X1 pe_1_3_2_add_83_U1_3 ( .A(int_data_res_3__2__3_), .B(
        pe_1_3_2_int_data_3_), .CI(pe_1_3_2_add_83_carry[3]), .CO(
        pe_1_3_2_add_83_carry[4]), .S(pe_1_3_2_N81) );
  FA_X1 pe_1_3_2_add_83_U1_2 ( .A(int_data_res_3__2__2_), .B(
        pe_1_3_2_int_data_2_), .CI(pe_1_3_2_add_83_carry[2]), .CO(
        pe_1_3_2_add_83_carry[3]), .S(pe_1_3_2_N80) );
  FA_X1 pe_1_3_2_add_83_U1_1 ( .A(int_data_res_3__2__1_), .B(
        pe_1_3_2_int_data_1_), .CI(pe_1_3_2_n2), .CO(pe_1_3_2_add_83_carry[2]), 
        .S(pe_1_3_2_N79) );
  NAND3_X1 pe_1_3_2_U56 ( .A1(n33), .A2(pe_1_3_2_n43), .A3(pe_1_3_2_n60), .ZN(
        pe_1_3_2_n40) );
  NAND3_X1 pe_1_3_2_U55 ( .A1(pe_1_3_2_n43), .A2(pe_1_3_2_n59), .A3(
        pe_1_3_2_n60), .ZN(pe_1_3_2_n39) );
  NAND3_X1 pe_1_3_2_U54 ( .A1(pe_1_3_2_n43), .A2(pe_1_3_2_n61), .A3(n33), .ZN(
        pe_1_3_2_n38) );
  NAND3_X1 pe_1_3_2_U53 ( .A1(pe_1_3_2_n59), .A2(pe_1_3_2_n61), .A3(
        pe_1_3_2_n43), .ZN(pe_1_3_2_n37) );
  DFFR_X1 pe_1_3_2_int_q_acc_reg_6_ ( .D(pe_1_3_2_n75), .CK(pe_1_3_2_net5524), 
        .RN(pe_1_3_2_n68), .Q(int_data_res_3__2__6_) );
  DFFR_X1 pe_1_3_2_int_q_acc_reg_5_ ( .D(pe_1_3_2_n76), .CK(pe_1_3_2_net5524), 
        .RN(pe_1_3_2_n68), .Q(int_data_res_3__2__5_) );
  DFFR_X1 pe_1_3_2_int_q_acc_reg_4_ ( .D(pe_1_3_2_n77), .CK(pe_1_3_2_net5524), 
        .RN(pe_1_3_2_n68), .Q(int_data_res_3__2__4_) );
  DFFR_X1 pe_1_3_2_int_q_acc_reg_3_ ( .D(pe_1_3_2_n78), .CK(pe_1_3_2_net5524), 
        .RN(pe_1_3_2_n68), .Q(int_data_res_3__2__3_) );
  DFFR_X1 pe_1_3_2_int_q_acc_reg_2_ ( .D(pe_1_3_2_n79), .CK(pe_1_3_2_net5524), 
        .RN(pe_1_3_2_n68), .Q(int_data_res_3__2__2_) );
  DFFR_X1 pe_1_3_2_int_q_acc_reg_1_ ( .D(pe_1_3_2_n80), .CK(pe_1_3_2_net5524), 
        .RN(pe_1_3_2_n68), .Q(int_data_res_3__2__1_) );
  DFFR_X1 pe_1_3_2_int_q_acc_reg_7_ ( .D(pe_1_3_2_n74), .CK(pe_1_3_2_net5524), 
        .RN(pe_1_3_2_n68), .Q(int_data_res_3__2__7_) );
  CLKGATETST_X1 pe_1_3_2_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_3_2_n85), .SE(1'b0), .GCK(pe_1_3_2_net5463) );
  CLKGATETST_X1 pe_1_3_2_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_3_2_n84), .SE(1'b0), .GCK(pe_1_3_2_net5469) );
  CLKGATETST_X1 pe_1_3_2_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_3_2_n83), .SE(1'b0), .GCK(pe_1_3_2_net5474) );
  CLKGATETST_X1 pe_1_3_2_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_3_2_n82), .SE(1'b0), .GCK(pe_1_3_2_net5479) );
  CLKGATETST_X1 pe_1_3_2_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_3_2_n87), .SE(1'b0), .GCK(pe_1_3_2_net5484) );
  CLKGATETST_X1 pe_1_3_2_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_3_2_n86), .SE(1'b0), .GCK(pe_1_3_2_net5489) );
  CLKGATETST_X1 pe_1_3_2_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_3_2_N64), .SE(1'b0), .GCK(pe_1_3_2_net5494) );
  CLKGATETST_X1 pe_1_3_2_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_3_2_N63), .SE(1'b0), .GCK(pe_1_3_2_net5499) );
  CLKGATETST_X1 pe_1_3_2_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_3_2_N62), .SE(1'b0), .GCK(pe_1_3_2_net5504) );
  CLKGATETST_X1 pe_1_3_2_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_3_2_N61), .SE(1'b0), .GCK(pe_1_3_2_net5509) );
  CLKGATETST_X1 pe_1_3_2_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_3_2_N60), .SE(1'b0), .GCK(pe_1_3_2_net5514) );
  CLKGATETST_X1 pe_1_3_2_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_3_2_N59), .SE(1'b0), .GCK(pe_1_3_2_net5519) );
  CLKGATETST_X1 pe_1_3_2_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_3_2_N90), .SE(1'b0), .GCK(pe_1_3_2_net5524) );
  CLKBUF_X1 pe_1_3_3_U110 ( .A(pe_1_3_3_n70), .Z(pe_1_3_3_n69) );
  INV_X1 pe_1_3_3_U109 ( .A(n75), .ZN(pe_1_3_3_n68) );
  INV_X1 pe_1_3_3_U108 ( .A(n67), .ZN(pe_1_3_3_n67) );
  INV_X1 pe_1_3_3_U107 ( .A(n67), .ZN(pe_1_3_3_n66) );
  INV_X1 pe_1_3_3_U106 ( .A(pe_1_3_3_n67), .ZN(pe_1_3_3_n65) );
  INV_X1 pe_1_3_3_U105 ( .A(pe_1_3_3_n62), .ZN(pe_1_3_3_n61) );
  INV_X1 pe_1_3_3_U104 ( .A(pe_1_3_3_n60), .ZN(pe_1_3_3_n59) );
  INV_X1 pe_1_3_3_U103 ( .A(n27), .ZN(pe_1_3_3_n58) );
  INV_X1 pe_1_3_3_U102 ( .A(n19), .ZN(pe_1_3_3_n57) );
  MUX2_X1 pe_1_3_3_U101 ( .A(pe_1_3_3_n54), .B(pe_1_3_3_n51), .S(n48), .Z(
        int_data_x_3__3__3_) );
  MUX2_X1 pe_1_3_3_U100 ( .A(pe_1_3_3_n53), .B(pe_1_3_3_n52), .S(pe_1_3_3_n61), 
        .Z(pe_1_3_3_n54) );
  MUX2_X1 pe_1_3_3_U99 ( .A(pe_1_3_3_int_q_reg_h[23]), .B(
        pe_1_3_3_int_q_reg_h[19]), .S(pe_1_3_3_n56), .Z(pe_1_3_3_n53) );
  MUX2_X1 pe_1_3_3_U98 ( .A(pe_1_3_3_int_q_reg_h[15]), .B(
        pe_1_3_3_int_q_reg_h[11]), .S(pe_1_3_3_n56), .Z(pe_1_3_3_n52) );
  MUX2_X1 pe_1_3_3_U97 ( .A(pe_1_3_3_int_q_reg_h[7]), .B(
        pe_1_3_3_int_q_reg_h[3]), .S(pe_1_3_3_n56), .Z(pe_1_3_3_n51) );
  MUX2_X1 pe_1_3_3_U96 ( .A(pe_1_3_3_n50), .B(pe_1_3_3_n47), .S(n48), .Z(
        int_data_x_3__3__2_) );
  MUX2_X1 pe_1_3_3_U95 ( .A(pe_1_3_3_n49), .B(pe_1_3_3_n48), .S(pe_1_3_3_n61), 
        .Z(pe_1_3_3_n50) );
  MUX2_X1 pe_1_3_3_U94 ( .A(pe_1_3_3_int_q_reg_h[22]), .B(
        pe_1_3_3_int_q_reg_h[18]), .S(pe_1_3_3_n56), .Z(pe_1_3_3_n49) );
  MUX2_X1 pe_1_3_3_U93 ( .A(pe_1_3_3_int_q_reg_h[14]), .B(
        pe_1_3_3_int_q_reg_h[10]), .S(pe_1_3_3_n56), .Z(pe_1_3_3_n48) );
  MUX2_X1 pe_1_3_3_U92 ( .A(pe_1_3_3_int_q_reg_h[6]), .B(
        pe_1_3_3_int_q_reg_h[2]), .S(pe_1_3_3_n56), .Z(pe_1_3_3_n47) );
  MUX2_X1 pe_1_3_3_U91 ( .A(pe_1_3_3_n46), .B(pe_1_3_3_n24), .S(n48), .Z(
        int_data_x_3__3__1_) );
  MUX2_X1 pe_1_3_3_U90 ( .A(pe_1_3_3_n45), .B(pe_1_3_3_n25), .S(pe_1_3_3_n61), 
        .Z(pe_1_3_3_n46) );
  MUX2_X1 pe_1_3_3_U89 ( .A(pe_1_3_3_int_q_reg_h[21]), .B(
        pe_1_3_3_int_q_reg_h[17]), .S(pe_1_3_3_n56), .Z(pe_1_3_3_n45) );
  MUX2_X1 pe_1_3_3_U88 ( .A(pe_1_3_3_int_q_reg_h[13]), .B(
        pe_1_3_3_int_q_reg_h[9]), .S(pe_1_3_3_n56), .Z(pe_1_3_3_n25) );
  MUX2_X1 pe_1_3_3_U87 ( .A(pe_1_3_3_int_q_reg_h[5]), .B(
        pe_1_3_3_int_q_reg_h[1]), .S(pe_1_3_3_n56), .Z(pe_1_3_3_n24) );
  MUX2_X1 pe_1_3_3_U86 ( .A(pe_1_3_3_n23), .B(pe_1_3_3_n20), .S(n48), .Z(
        int_data_x_3__3__0_) );
  MUX2_X1 pe_1_3_3_U85 ( .A(pe_1_3_3_n22), .B(pe_1_3_3_n21), .S(pe_1_3_3_n61), 
        .Z(pe_1_3_3_n23) );
  MUX2_X1 pe_1_3_3_U84 ( .A(pe_1_3_3_int_q_reg_h[20]), .B(
        pe_1_3_3_int_q_reg_h[16]), .S(pe_1_3_3_n56), .Z(pe_1_3_3_n22) );
  MUX2_X1 pe_1_3_3_U83 ( .A(pe_1_3_3_int_q_reg_h[12]), .B(
        pe_1_3_3_int_q_reg_h[8]), .S(pe_1_3_3_n56), .Z(pe_1_3_3_n21) );
  MUX2_X1 pe_1_3_3_U82 ( .A(pe_1_3_3_int_q_reg_h[4]), .B(
        pe_1_3_3_int_q_reg_h[0]), .S(pe_1_3_3_n56), .Z(pe_1_3_3_n20) );
  MUX2_X1 pe_1_3_3_U81 ( .A(pe_1_3_3_n19), .B(pe_1_3_3_n16), .S(n48), .Z(
        int_data_y_3__3__3_) );
  MUX2_X1 pe_1_3_3_U80 ( .A(pe_1_3_3_n18), .B(pe_1_3_3_n17), .S(pe_1_3_3_n61), 
        .Z(pe_1_3_3_n19) );
  MUX2_X1 pe_1_3_3_U79 ( .A(pe_1_3_3_int_q_reg_v[23]), .B(
        pe_1_3_3_int_q_reg_v[19]), .S(pe_1_3_3_n55), .Z(pe_1_3_3_n18) );
  MUX2_X1 pe_1_3_3_U78 ( .A(pe_1_3_3_int_q_reg_v[15]), .B(
        pe_1_3_3_int_q_reg_v[11]), .S(pe_1_3_3_n55), .Z(pe_1_3_3_n17) );
  MUX2_X1 pe_1_3_3_U77 ( .A(pe_1_3_3_int_q_reg_v[7]), .B(
        pe_1_3_3_int_q_reg_v[3]), .S(pe_1_3_3_n55), .Z(pe_1_3_3_n16) );
  MUX2_X1 pe_1_3_3_U76 ( .A(pe_1_3_3_n15), .B(pe_1_3_3_n12), .S(n48), .Z(
        int_data_y_3__3__2_) );
  MUX2_X1 pe_1_3_3_U75 ( .A(pe_1_3_3_n14), .B(pe_1_3_3_n13), .S(pe_1_3_3_n61), 
        .Z(pe_1_3_3_n15) );
  MUX2_X1 pe_1_3_3_U74 ( .A(pe_1_3_3_int_q_reg_v[22]), .B(
        pe_1_3_3_int_q_reg_v[18]), .S(pe_1_3_3_n55), .Z(pe_1_3_3_n14) );
  MUX2_X1 pe_1_3_3_U73 ( .A(pe_1_3_3_int_q_reg_v[14]), .B(
        pe_1_3_3_int_q_reg_v[10]), .S(pe_1_3_3_n55), .Z(pe_1_3_3_n13) );
  MUX2_X1 pe_1_3_3_U72 ( .A(pe_1_3_3_int_q_reg_v[6]), .B(
        pe_1_3_3_int_q_reg_v[2]), .S(pe_1_3_3_n55), .Z(pe_1_3_3_n12) );
  MUX2_X1 pe_1_3_3_U71 ( .A(pe_1_3_3_n11), .B(pe_1_3_3_n8), .S(n48), .Z(
        int_data_y_3__3__1_) );
  MUX2_X1 pe_1_3_3_U70 ( .A(pe_1_3_3_n10), .B(pe_1_3_3_n9), .S(pe_1_3_3_n61), 
        .Z(pe_1_3_3_n11) );
  MUX2_X1 pe_1_3_3_U69 ( .A(pe_1_3_3_int_q_reg_v[21]), .B(
        pe_1_3_3_int_q_reg_v[17]), .S(pe_1_3_3_n55), .Z(pe_1_3_3_n10) );
  MUX2_X1 pe_1_3_3_U68 ( .A(pe_1_3_3_int_q_reg_v[13]), .B(
        pe_1_3_3_int_q_reg_v[9]), .S(pe_1_3_3_n55), .Z(pe_1_3_3_n9) );
  MUX2_X1 pe_1_3_3_U67 ( .A(pe_1_3_3_int_q_reg_v[5]), .B(
        pe_1_3_3_int_q_reg_v[1]), .S(pe_1_3_3_n55), .Z(pe_1_3_3_n8) );
  MUX2_X1 pe_1_3_3_U66 ( .A(pe_1_3_3_n7), .B(pe_1_3_3_n4), .S(n48), .Z(
        int_data_y_3__3__0_) );
  MUX2_X1 pe_1_3_3_U65 ( .A(pe_1_3_3_n6), .B(pe_1_3_3_n5), .S(pe_1_3_3_n61), 
        .Z(pe_1_3_3_n7) );
  MUX2_X1 pe_1_3_3_U64 ( .A(pe_1_3_3_int_q_reg_v[20]), .B(
        pe_1_3_3_int_q_reg_v[16]), .S(pe_1_3_3_n55), .Z(pe_1_3_3_n6) );
  MUX2_X1 pe_1_3_3_U63 ( .A(pe_1_3_3_int_q_reg_v[12]), .B(
        pe_1_3_3_int_q_reg_v[8]), .S(pe_1_3_3_n55), .Z(pe_1_3_3_n5) );
  MUX2_X1 pe_1_3_3_U62 ( .A(pe_1_3_3_int_q_reg_v[4]), .B(
        pe_1_3_3_int_q_reg_v[0]), .S(pe_1_3_3_n55), .Z(pe_1_3_3_n4) );
  AOI222_X1 pe_1_3_3_U61 ( .A1(int_data_res_4__3__2_), .A2(pe_1_3_3_n63), .B1(
        pe_1_3_3_N80), .B2(pe_1_3_3_n27), .C1(pe_1_3_3_N72), .C2(pe_1_3_3_n28), 
        .ZN(pe_1_3_3_n33) );
  INV_X1 pe_1_3_3_U60 ( .A(pe_1_3_3_n33), .ZN(pe_1_3_3_n80) );
  AOI222_X1 pe_1_3_3_U59 ( .A1(int_data_res_4__3__6_), .A2(pe_1_3_3_n63), .B1(
        pe_1_3_3_N84), .B2(pe_1_3_3_n27), .C1(pe_1_3_3_N76), .C2(pe_1_3_3_n28), 
        .ZN(pe_1_3_3_n29) );
  INV_X1 pe_1_3_3_U58 ( .A(pe_1_3_3_n29), .ZN(pe_1_3_3_n76) );
  XNOR2_X1 pe_1_3_3_U57 ( .A(pe_1_3_3_n71), .B(int_data_res_3__3__0_), .ZN(
        pe_1_3_3_N70) );
  AOI222_X1 pe_1_3_3_U52 ( .A1(int_data_res_4__3__0_), .A2(pe_1_3_3_n63), .B1(
        pe_1_3_3_n1), .B2(pe_1_3_3_n27), .C1(pe_1_3_3_N70), .C2(pe_1_3_3_n28), 
        .ZN(pe_1_3_3_n35) );
  INV_X1 pe_1_3_3_U51 ( .A(pe_1_3_3_n35), .ZN(pe_1_3_3_n82) );
  AOI222_X1 pe_1_3_3_U50 ( .A1(int_data_res_4__3__1_), .A2(pe_1_3_3_n63), .B1(
        pe_1_3_3_N79), .B2(pe_1_3_3_n27), .C1(pe_1_3_3_N71), .C2(pe_1_3_3_n28), 
        .ZN(pe_1_3_3_n34) );
  INV_X1 pe_1_3_3_U49 ( .A(pe_1_3_3_n34), .ZN(pe_1_3_3_n81) );
  AOI222_X1 pe_1_3_3_U48 ( .A1(int_data_res_4__3__3_), .A2(pe_1_3_3_n63), .B1(
        pe_1_3_3_N81), .B2(pe_1_3_3_n27), .C1(pe_1_3_3_N73), .C2(pe_1_3_3_n28), 
        .ZN(pe_1_3_3_n32) );
  INV_X1 pe_1_3_3_U47 ( .A(pe_1_3_3_n32), .ZN(pe_1_3_3_n79) );
  AOI222_X1 pe_1_3_3_U46 ( .A1(int_data_res_4__3__4_), .A2(pe_1_3_3_n63), .B1(
        pe_1_3_3_N82), .B2(pe_1_3_3_n27), .C1(pe_1_3_3_N74), .C2(pe_1_3_3_n28), 
        .ZN(pe_1_3_3_n31) );
  INV_X1 pe_1_3_3_U45 ( .A(pe_1_3_3_n31), .ZN(pe_1_3_3_n78) );
  AOI222_X1 pe_1_3_3_U44 ( .A1(int_data_res_4__3__5_), .A2(pe_1_3_3_n63), .B1(
        pe_1_3_3_N83), .B2(pe_1_3_3_n27), .C1(pe_1_3_3_N75), .C2(pe_1_3_3_n28), 
        .ZN(pe_1_3_3_n30) );
  INV_X1 pe_1_3_3_U43 ( .A(pe_1_3_3_n30), .ZN(pe_1_3_3_n77) );
  NAND2_X1 pe_1_3_3_U42 ( .A1(pe_1_3_3_int_data_0_), .A2(pe_1_3_3_n3), .ZN(
        pe_1_3_3_sub_81_carry[1]) );
  INV_X1 pe_1_3_3_U41 ( .A(pe_1_3_3_int_data_1_), .ZN(pe_1_3_3_n72) );
  INV_X1 pe_1_3_3_U40 ( .A(pe_1_3_3_int_data_2_), .ZN(pe_1_3_3_n73) );
  AND2_X1 pe_1_3_3_U39 ( .A1(pe_1_3_3_int_data_0_), .A2(int_data_res_3__3__0_), 
        .ZN(pe_1_3_3_n2) );
  AOI222_X1 pe_1_3_3_U38 ( .A1(pe_1_3_3_n63), .A2(int_data_res_4__3__7_), .B1(
        pe_1_3_3_N85), .B2(pe_1_3_3_n27), .C1(pe_1_3_3_N77), .C2(pe_1_3_3_n28), 
        .ZN(pe_1_3_3_n26) );
  INV_X1 pe_1_3_3_U37 ( .A(pe_1_3_3_n26), .ZN(pe_1_3_3_n75) );
  NOR3_X1 pe_1_3_3_U36 ( .A1(pe_1_3_3_n58), .A2(pe_1_3_3_n64), .A3(int_ckg[36]), .ZN(pe_1_3_3_n36) );
  OR2_X1 pe_1_3_3_U35 ( .A1(pe_1_3_3_n36), .A2(pe_1_3_3_n63), .ZN(pe_1_3_3_N90) );
  INV_X1 pe_1_3_3_U34 ( .A(n39), .ZN(pe_1_3_3_n62) );
  AND2_X1 pe_1_3_3_U33 ( .A1(int_data_x_3__3__2_), .A2(n27), .ZN(
        pe_1_3_3_int_data_2_) );
  AND2_X1 pe_1_3_3_U32 ( .A1(int_data_x_3__3__1_), .A2(n27), .ZN(
        pe_1_3_3_int_data_1_) );
  AND2_X1 pe_1_3_3_U31 ( .A1(int_data_x_3__3__3_), .A2(n27), .ZN(
        pe_1_3_3_int_data_3_) );
  BUF_X1 pe_1_3_3_U30 ( .A(n61), .Z(pe_1_3_3_n63) );
  INV_X1 pe_1_3_3_U29 ( .A(n33), .ZN(pe_1_3_3_n60) );
  AND2_X1 pe_1_3_3_U28 ( .A1(int_data_x_3__3__0_), .A2(n27), .ZN(
        pe_1_3_3_int_data_0_) );
  NAND2_X1 pe_1_3_3_U27 ( .A1(pe_1_3_3_n44), .A2(pe_1_3_3_n60), .ZN(
        pe_1_3_3_n41) );
  AND3_X1 pe_1_3_3_U26 ( .A1(n75), .A2(pe_1_3_3_n62), .A3(n48), .ZN(
        pe_1_3_3_n44) );
  INV_X1 pe_1_3_3_U25 ( .A(pe_1_3_3_int_data_3_), .ZN(pe_1_3_3_n74) );
  NOR2_X1 pe_1_3_3_U24 ( .A1(pe_1_3_3_n68), .A2(n48), .ZN(pe_1_3_3_n43) );
  NOR2_X1 pe_1_3_3_U23 ( .A1(pe_1_3_3_n57), .A2(pe_1_3_3_n63), .ZN(
        pe_1_3_3_n28) );
  NOR2_X1 pe_1_3_3_U22 ( .A1(n19), .A2(pe_1_3_3_n63), .ZN(pe_1_3_3_n27) );
  INV_X1 pe_1_3_3_U21 ( .A(pe_1_3_3_int_data_0_), .ZN(pe_1_3_3_n71) );
  INV_X1 pe_1_3_3_U20 ( .A(pe_1_3_3_n41), .ZN(pe_1_3_3_n88) );
  INV_X1 pe_1_3_3_U19 ( .A(pe_1_3_3_n37), .ZN(pe_1_3_3_n86) );
  INV_X1 pe_1_3_3_U18 ( .A(pe_1_3_3_n38), .ZN(pe_1_3_3_n85) );
  INV_X1 pe_1_3_3_U17 ( .A(pe_1_3_3_n39), .ZN(pe_1_3_3_n84) );
  NOR2_X1 pe_1_3_3_U16 ( .A1(pe_1_3_3_n66), .A2(pe_1_3_3_n42), .ZN(
        pe_1_3_3_N59) );
  NOR2_X1 pe_1_3_3_U15 ( .A1(pe_1_3_3_n66), .A2(pe_1_3_3_n41), .ZN(
        pe_1_3_3_N60) );
  NOR2_X1 pe_1_3_3_U14 ( .A1(pe_1_3_3_n66), .A2(pe_1_3_3_n38), .ZN(
        pe_1_3_3_N63) );
  NOR2_X1 pe_1_3_3_U13 ( .A1(pe_1_3_3_n66), .A2(pe_1_3_3_n40), .ZN(
        pe_1_3_3_N61) );
  NOR2_X1 pe_1_3_3_U12 ( .A1(pe_1_3_3_n66), .A2(pe_1_3_3_n39), .ZN(
        pe_1_3_3_N62) );
  NOR2_X1 pe_1_3_3_U11 ( .A1(pe_1_3_3_n37), .A2(pe_1_3_3_n66), .ZN(
        pe_1_3_3_N64) );
  NAND2_X1 pe_1_3_3_U10 ( .A1(pe_1_3_3_n44), .A2(pe_1_3_3_n59), .ZN(
        pe_1_3_3_n42) );
  BUF_X1 pe_1_3_3_U9 ( .A(pe_1_3_3_n59), .Z(pe_1_3_3_n55) );
  INV_X1 pe_1_3_3_U8 ( .A(pe_1_3_3_n67), .ZN(pe_1_3_3_n64) );
  BUF_X1 pe_1_3_3_U7 ( .A(pe_1_3_3_n59), .Z(pe_1_3_3_n56) );
  INV_X1 pe_1_3_3_U6 ( .A(pe_1_3_3_n42), .ZN(pe_1_3_3_n87) );
  INV_X1 pe_1_3_3_U5 ( .A(pe_1_3_3_n40), .ZN(pe_1_3_3_n83) );
  INV_X2 pe_1_3_3_U4 ( .A(n83), .ZN(pe_1_3_3_n70) );
  XOR2_X1 pe_1_3_3_U3 ( .A(pe_1_3_3_int_data_0_), .B(int_data_res_3__3__0_), 
        .Z(pe_1_3_3_n1) );
  DFFR_X1 pe_1_3_3_int_q_acc_reg_0_ ( .D(pe_1_3_3_n82), .CK(pe_1_3_3_net5446), 
        .RN(pe_1_3_3_n70), .Q(int_data_res_3__3__0_), .QN(pe_1_3_3_n3) );
  DFFR_X1 pe_1_3_3_int_q_reg_v_reg_0__0_ ( .D(int_data_y_4__3__0_), .CK(
        pe_1_3_3_net5416), .RN(pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_v[20]) );
  DFFR_X1 pe_1_3_3_int_q_reg_v_reg_0__1_ ( .D(int_data_y_4__3__1_), .CK(
        pe_1_3_3_net5416), .RN(pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_v[21]) );
  DFFR_X1 pe_1_3_3_int_q_reg_v_reg_0__2_ ( .D(int_data_y_4__3__2_), .CK(
        pe_1_3_3_net5416), .RN(pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_v[22]) );
  DFFR_X1 pe_1_3_3_int_q_reg_v_reg_0__3_ ( .D(int_data_y_4__3__3_), .CK(
        pe_1_3_3_net5416), .RN(pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_v[23]) );
  DFFR_X1 pe_1_3_3_int_q_reg_v_reg_1__0_ ( .D(int_data_y_4__3__0_), .CK(
        pe_1_3_3_net5421), .RN(pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_v[16]) );
  DFFR_X1 pe_1_3_3_int_q_reg_v_reg_1__1_ ( .D(int_data_y_4__3__1_), .CK(
        pe_1_3_3_net5421), .RN(pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_v[17]) );
  DFFR_X1 pe_1_3_3_int_q_reg_v_reg_1__2_ ( .D(int_data_y_4__3__2_), .CK(
        pe_1_3_3_net5421), .RN(pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_v[18]) );
  DFFR_X1 pe_1_3_3_int_q_reg_v_reg_1__3_ ( .D(int_data_y_4__3__3_), .CK(
        pe_1_3_3_net5421), .RN(pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_v[19]) );
  DFFR_X1 pe_1_3_3_int_q_reg_v_reg_2__0_ ( .D(int_data_y_4__3__0_), .CK(
        pe_1_3_3_net5426), .RN(pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_v[12]) );
  DFFR_X1 pe_1_3_3_int_q_reg_v_reg_2__1_ ( .D(int_data_y_4__3__1_), .CK(
        pe_1_3_3_net5426), .RN(pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_v[13]) );
  DFFR_X1 pe_1_3_3_int_q_reg_v_reg_2__2_ ( .D(int_data_y_4__3__2_), .CK(
        pe_1_3_3_net5426), .RN(pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_v[14]) );
  DFFR_X1 pe_1_3_3_int_q_reg_v_reg_2__3_ ( .D(int_data_y_4__3__3_), .CK(
        pe_1_3_3_net5426), .RN(pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_v[15]) );
  DFFR_X1 pe_1_3_3_int_q_reg_v_reg_3__0_ ( .D(int_data_y_4__3__0_), .CK(
        pe_1_3_3_net5431), .RN(pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_v[8]) );
  DFFR_X1 pe_1_3_3_int_q_reg_v_reg_3__1_ ( .D(int_data_y_4__3__1_), .CK(
        pe_1_3_3_net5431), .RN(pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_v[9]) );
  DFFR_X1 pe_1_3_3_int_q_reg_v_reg_3__2_ ( .D(int_data_y_4__3__2_), .CK(
        pe_1_3_3_net5431), .RN(pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_v[10]) );
  DFFR_X1 pe_1_3_3_int_q_reg_v_reg_3__3_ ( .D(int_data_y_4__3__3_), .CK(
        pe_1_3_3_net5431), .RN(pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_v[11]) );
  DFFR_X1 pe_1_3_3_int_q_reg_v_reg_4__0_ ( .D(int_data_y_4__3__0_), .CK(
        pe_1_3_3_net5436), .RN(pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_v[4]) );
  DFFR_X1 pe_1_3_3_int_q_reg_v_reg_4__1_ ( .D(int_data_y_4__3__1_), .CK(
        pe_1_3_3_net5436), .RN(pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_v[5]) );
  DFFR_X1 pe_1_3_3_int_q_reg_v_reg_4__2_ ( .D(int_data_y_4__3__2_), .CK(
        pe_1_3_3_net5436), .RN(pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_v[6]) );
  DFFR_X1 pe_1_3_3_int_q_reg_v_reg_4__3_ ( .D(int_data_y_4__3__3_), .CK(
        pe_1_3_3_net5436), .RN(pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_v[7]) );
  DFFR_X1 pe_1_3_3_int_q_reg_v_reg_5__0_ ( .D(int_data_y_4__3__0_), .CK(
        pe_1_3_3_net5441), .RN(pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_v[0]) );
  DFFR_X1 pe_1_3_3_int_q_reg_v_reg_5__1_ ( .D(int_data_y_4__3__1_), .CK(
        pe_1_3_3_net5441), .RN(pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_v[1]) );
  DFFR_X1 pe_1_3_3_int_q_reg_v_reg_5__2_ ( .D(int_data_y_4__3__2_), .CK(
        pe_1_3_3_net5441), .RN(pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_v[2]) );
  DFFR_X1 pe_1_3_3_int_q_reg_v_reg_5__3_ ( .D(int_data_y_4__3__3_), .CK(
        pe_1_3_3_net5441), .RN(pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_3_3_int_q_reg_h_reg_0__0_ ( .D(int_data_x_3__4__0_), .SI(
        int_data_y_4__3__0_), .SE(pe_1_3_3_n64), .CK(pe_1_3_3_net5385), .RN(
        pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_3_3_int_q_reg_h_reg_0__1_ ( .D(int_data_x_3__4__1_), .SI(
        int_data_y_4__3__1_), .SE(pe_1_3_3_n64), .CK(pe_1_3_3_net5385), .RN(
        pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_3_3_int_q_reg_h_reg_0__2_ ( .D(int_data_x_3__4__2_), .SI(
        int_data_y_4__3__2_), .SE(pe_1_3_3_n64), .CK(pe_1_3_3_net5385), .RN(
        pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_3_3_int_q_reg_h_reg_0__3_ ( .D(int_data_x_3__4__3_), .SI(
        int_data_y_4__3__3_), .SE(pe_1_3_3_n64), .CK(pe_1_3_3_net5385), .RN(
        pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_3_3_int_q_reg_h_reg_1__0_ ( .D(int_data_x_3__4__0_), .SI(
        int_data_y_4__3__0_), .SE(pe_1_3_3_n64), .CK(pe_1_3_3_net5391), .RN(
        pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_3_3_int_q_reg_h_reg_1__1_ ( .D(int_data_x_3__4__1_), .SI(
        int_data_y_4__3__1_), .SE(pe_1_3_3_n64), .CK(pe_1_3_3_net5391), .RN(
        pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_3_3_int_q_reg_h_reg_1__2_ ( .D(int_data_x_3__4__2_), .SI(
        int_data_y_4__3__2_), .SE(pe_1_3_3_n64), .CK(pe_1_3_3_net5391), .RN(
        pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_3_3_int_q_reg_h_reg_1__3_ ( .D(int_data_x_3__4__3_), .SI(
        int_data_y_4__3__3_), .SE(pe_1_3_3_n64), .CK(pe_1_3_3_net5391), .RN(
        pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_3_3_int_q_reg_h_reg_2__0_ ( .D(int_data_x_3__4__0_), .SI(
        int_data_y_4__3__0_), .SE(pe_1_3_3_n64), .CK(pe_1_3_3_net5396), .RN(
        pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_3_3_int_q_reg_h_reg_2__1_ ( .D(int_data_x_3__4__1_), .SI(
        int_data_y_4__3__1_), .SE(pe_1_3_3_n64), .CK(pe_1_3_3_net5396), .RN(
        pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_3_3_int_q_reg_h_reg_2__2_ ( .D(int_data_x_3__4__2_), .SI(
        int_data_y_4__3__2_), .SE(pe_1_3_3_n64), .CK(pe_1_3_3_net5396), .RN(
        pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_3_3_int_q_reg_h_reg_2__3_ ( .D(int_data_x_3__4__3_), .SI(
        int_data_y_4__3__3_), .SE(pe_1_3_3_n64), .CK(pe_1_3_3_net5396), .RN(
        pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_3_3_int_q_reg_h_reg_3__0_ ( .D(int_data_x_3__4__0_), .SI(
        int_data_y_4__3__0_), .SE(pe_1_3_3_n64), .CK(pe_1_3_3_net5401), .RN(
        pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_3_3_int_q_reg_h_reg_3__1_ ( .D(int_data_x_3__4__1_), .SI(
        int_data_y_4__3__1_), .SE(pe_1_3_3_n64), .CK(pe_1_3_3_net5401), .RN(
        pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_3_3_int_q_reg_h_reg_3__2_ ( .D(int_data_x_3__4__2_), .SI(
        int_data_y_4__3__2_), .SE(pe_1_3_3_n64), .CK(pe_1_3_3_net5401), .RN(
        pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_3_3_int_q_reg_h_reg_3__3_ ( .D(int_data_x_3__4__3_), .SI(
        int_data_y_4__3__3_), .SE(pe_1_3_3_n64), .CK(pe_1_3_3_net5401), .RN(
        pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_3_3_int_q_reg_h_reg_4__0_ ( .D(int_data_x_3__4__0_), .SI(
        int_data_y_4__3__0_), .SE(pe_1_3_3_n65), .CK(pe_1_3_3_net5406), .RN(
        pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_3_3_int_q_reg_h_reg_4__1_ ( .D(int_data_x_3__4__1_), .SI(
        int_data_y_4__3__1_), .SE(pe_1_3_3_n65), .CK(pe_1_3_3_net5406), .RN(
        pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_3_3_int_q_reg_h_reg_4__2_ ( .D(int_data_x_3__4__2_), .SI(
        int_data_y_4__3__2_), .SE(pe_1_3_3_n65), .CK(pe_1_3_3_net5406), .RN(
        pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_3_3_int_q_reg_h_reg_4__3_ ( .D(int_data_x_3__4__3_), .SI(
        int_data_y_4__3__3_), .SE(pe_1_3_3_n65), .CK(pe_1_3_3_net5406), .RN(
        pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_3_3_int_q_reg_h_reg_5__0_ ( .D(int_data_x_3__4__0_), .SI(
        int_data_y_4__3__0_), .SE(pe_1_3_3_n65), .CK(pe_1_3_3_net5411), .RN(
        pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_3_3_int_q_reg_h_reg_5__1_ ( .D(int_data_x_3__4__1_), .SI(
        int_data_y_4__3__1_), .SE(pe_1_3_3_n65), .CK(pe_1_3_3_net5411), .RN(
        pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_3_3_int_q_reg_h_reg_5__2_ ( .D(int_data_x_3__4__2_), .SI(
        int_data_y_4__3__2_), .SE(pe_1_3_3_n65), .CK(pe_1_3_3_net5411), .RN(
        pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_3_3_int_q_reg_h_reg_5__3_ ( .D(int_data_x_3__4__3_), .SI(
        int_data_y_4__3__3_), .SE(pe_1_3_3_n65), .CK(pe_1_3_3_net5411), .RN(
        pe_1_3_3_n70), .Q(pe_1_3_3_int_q_reg_h[3]) );
  FA_X1 pe_1_3_3_sub_81_U2_7 ( .A(int_data_res_3__3__7_), .B(pe_1_3_3_n74), 
        .CI(pe_1_3_3_sub_81_carry[7]), .S(pe_1_3_3_N77) );
  FA_X1 pe_1_3_3_sub_81_U2_6 ( .A(int_data_res_3__3__6_), .B(pe_1_3_3_n74), 
        .CI(pe_1_3_3_sub_81_carry[6]), .CO(pe_1_3_3_sub_81_carry[7]), .S(
        pe_1_3_3_N76) );
  FA_X1 pe_1_3_3_sub_81_U2_5 ( .A(int_data_res_3__3__5_), .B(pe_1_3_3_n74), 
        .CI(pe_1_3_3_sub_81_carry[5]), .CO(pe_1_3_3_sub_81_carry[6]), .S(
        pe_1_3_3_N75) );
  FA_X1 pe_1_3_3_sub_81_U2_4 ( .A(int_data_res_3__3__4_), .B(pe_1_3_3_n74), 
        .CI(pe_1_3_3_sub_81_carry[4]), .CO(pe_1_3_3_sub_81_carry[5]), .S(
        pe_1_3_3_N74) );
  FA_X1 pe_1_3_3_sub_81_U2_3 ( .A(int_data_res_3__3__3_), .B(pe_1_3_3_n74), 
        .CI(pe_1_3_3_sub_81_carry[3]), .CO(pe_1_3_3_sub_81_carry[4]), .S(
        pe_1_3_3_N73) );
  FA_X1 pe_1_3_3_sub_81_U2_2 ( .A(int_data_res_3__3__2_), .B(pe_1_3_3_n73), 
        .CI(pe_1_3_3_sub_81_carry[2]), .CO(pe_1_3_3_sub_81_carry[3]), .S(
        pe_1_3_3_N72) );
  FA_X1 pe_1_3_3_sub_81_U2_1 ( .A(int_data_res_3__3__1_), .B(pe_1_3_3_n72), 
        .CI(pe_1_3_3_sub_81_carry[1]), .CO(pe_1_3_3_sub_81_carry[2]), .S(
        pe_1_3_3_N71) );
  FA_X1 pe_1_3_3_add_83_U1_7 ( .A(int_data_res_3__3__7_), .B(
        pe_1_3_3_int_data_3_), .CI(pe_1_3_3_add_83_carry[7]), .S(pe_1_3_3_N85)
         );
  FA_X1 pe_1_3_3_add_83_U1_6 ( .A(int_data_res_3__3__6_), .B(
        pe_1_3_3_int_data_3_), .CI(pe_1_3_3_add_83_carry[6]), .CO(
        pe_1_3_3_add_83_carry[7]), .S(pe_1_3_3_N84) );
  FA_X1 pe_1_3_3_add_83_U1_5 ( .A(int_data_res_3__3__5_), .B(
        pe_1_3_3_int_data_3_), .CI(pe_1_3_3_add_83_carry[5]), .CO(
        pe_1_3_3_add_83_carry[6]), .S(pe_1_3_3_N83) );
  FA_X1 pe_1_3_3_add_83_U1_4 ( .A(int_data_res_3__3__4_), .B(
        pe_1_3_3_int_data_3_), .CI(pe_1_3_3_add_83_carry[4]), .CO(
        pe_1_3_3_add_83_carry[5]), .S(pe_1_3_3_N82) );
  FA_X1 pe_1_3_3_add_83_U1_3 ( .A(int_data_res_3__3__3_), .B(
        pe_1_3_3_int_data_3_), .CI(pe_1_3_3_add_83_carry[3]), .CO(
        pe_1_3_3_add_83_carry[4]), .S(pe_1_3_3_N81) );
  FA_X1 pe_1_3_3_add_83_U1_2 ( .A(int_data_res_3__3__2_), .B(
        pe_1_3_3_int_data_2_), .CI(pe_1_3_3_add_83_carry[2]), .CO(
        pe_1_3_3_add_83_carry[3]), .S(pe_1_3_3_N80) );
  FA_X1 pe_1_3_3_add_83_U1_1 ( .A(int_data_res_3__3__1_), .B(
        pe_1_3_3_int_data_1_), .CI(pe_1_3_3_n2), .CO(pe_1_3_3_add_83_carry[2]), 
        .S(pe_1_3_3_N79) );
  NAND3_X1 pe_1_3_3_U56 ( .A1(pe_1_3_3_n59), .A2(pe_1_3_3_n43), .A3(
        pe_1_3_3_n61), .ZN(pe_1_3_3_n40) );
  NAND3_X1 pe_1_3_3_U55 ( .A1(pe_1_3_3_n43), .A2(pe_1_3_3_n60), .A3(
        pe_1_3_3_n61), .ZN(pe_1_3_3_n39) );
  NAND3_X1 pe_1_3_3_U54 ( .A1(pe_1_3_3_n43), .A2(pe_1_3_3_n62), .A3(
        pe_1_3_3_n59), .ZN(pe_1_3_3_n38) );
  NAND3_X1 pe_1_3_3_U53 ( .A1(pe_1_3_3_n60), .A2(pe_1_3_3_n62), .A3(
        pe_1_3_3_n43), .ZN(pe_1_3_3_n37) );
  DFFR_X1 pe_1_3_3_int_q_acc_reg_6_ ( .D(pe_1_3_3_n76), .CK(pe_1_3_3_net5446), 
        .RN(pe_1_3_3_n69), .Q(int_data_res_3__3__6_) );
  DFFR_X1 pe_1_3_3_int_q_acc_reg_5_ ( .D(pe_1_3_3_n77), .CK(pe_1_3_3_net5446), 
        .RN(pe_1_3_3_n69), .Q(int_data_res_3__3__5_) );
  DFFR_X1 pe_1_3_3_int_q_acc_reg_4_ ( .D(pe_1_3_3_n78), .CK(pe_1_3_3_net5446), 
        .RN(pe_1_3_3_n69), .Q(int_data_res_3__3__4_) );
  DFFR_X1 pe_1_3_3_int_q_acc_reg_3_ ( .D(pe_1_3_3_n79), .CK(pe_1_3_3_net5446), 
        .RN(pe_1_3_3_n69), .Q(int_data_res_3__3__3_) );
  DFFR_X1 pe_1_3_3_int_q_acc_reg_2_ ( .D(pe_1_3_3_n80), .CK(pe_1_3_3_net5446), 
        .RN(pe_1_3_3_n69), .Q(int_data_res_3__3__2_) );
  DFFR_X1 pe_1_3_3_int_q_acc_reg_1_ ( .D(pe_1_3_3_n81), .CK(pe_1_3_3_net5446), 
        .RN(pe_1_3_3_n69), .Q(int_data_res_3__3__1_) );
  DFFR_X1 pe_1_3_3_int_q_acc_reg_7_ ( .D(pe_1_3_3_n75), .CK(pe_1_3_3_net5446), 
        .RN(pe_1_3_3_n69), .Q(int_data_res_3__3__7_) );
  CLKGATETST_X1 pe_1_3_3_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_3_3_n86), .SE(1'b0), .GCK(pe_1_3_3_net5385) );
  CLKGATETST_X1 pe_1_3_3_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_3_3_n85), .SE(1'b0), .GCK(pe_1_3_3_net5391) );
  CLKGATETST_X1 pe_1_3_3_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_3_3_n84), .SE(1'b0), .GCK(pe_1_3_3_net5396) );
  CLKGATETST_X1 pe_1_3_3_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_3_3_n83), .SE(1'b0), .GCK(pe_1_3_3_net5401) );
  CLKGATETST_X1 pe_1_3_3_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_3_3_n88), .SE(1'b0), .GCK(pe_1_3_3_net5406) );
  CLKGATETST_X1 pe_1_3_3_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_3_3_n87), .SE(1'b0), .GCK(pe_1_3_3_net5411) );
  CLKGATETST_X1 pe_1_3_3_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_3_3_N64), .SE(1'b0), .GCK(pe_1_3_3_net5416) );
  CLKGATETST_X1 pe_1_3_3_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_3_3_N63), .SE(1'b0), .GCK(pe_1_3_3_net5421) );
  CLKGATETST_X1 pe_1_3_3_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_3_3_N62), .SE(1'b0), .GCK(pe_1_3_3_net5426) );
  CLKGATETST_X1 pe_1_3_3_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_3_3_N61), .SE(1'b0), .GCK(pe_1_3_3_net5431) );
  CLKGATETST_X1 pe_1_3_3_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_3_3_N60), .SE(1'b0), .GCK(pe_1_3_3_net5436) );
  CLKGATETST_X1 pe_1_3_3_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_3_3_N59), .SE(1'b0), .GCK(pe_1_3_3_net5441) );
  CLKGATETST_X1 pe_1_3_3_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_3_3_N90), .SE(1'b0), .GCK(pe_1_3_3_net5446) );
  CLKBUF_X1 pe_1_3_4_U112 ( .A(pe_1_3_4_n72), .Z(pe_1_3_4_n71) );
  INV_X1 pe_1_3_4_U111 ( .A(n75), .ZN(pe_1_3_4_n70) );
  INV_X1 pe_1_3_4_U110 ( .A(n67), .ZN(pe_1_3_4_n69) );
  INV_X1 pe_1_3_4_U109 ( .A(n67), .ZN(pe_1_3_4_n68) );
  INV_X1 pe_1_3_4_U108 ( .A(n67), .ZN(pe_1_3_4_n67) );
  INV_X1 pe_1_3_4_U107 ( .A(pe_1_3_4_n69), .ZN(pe_1_3_4_n66) );
  INV_X1 pe_1_3_4_U106 ( .A(pe_1_3_4_n63), .ZN(pe_1_3_4_n62) );
  INV_X1 pe_1_3_4_U105 ( .A(pe_1_3_4_n61), .ZN(pe_1_3_4_n60) );
  INV_X1 pe_1_3_4_U104 ( .A(n27), .ZN(pe_1_3_4_n59) );
  INV_X1 pe_1_3_4_U103 ( .A(pe_1_3_4_n59), .ZN(pe_1_3_4_n58) );
  INV_X1 pe_1_3_4_U102 ( .A(n19), .ZN(pe_1_3_4_n57) );
  MUX2_X1 pe_1_3_4_U101 ( .A(pe_1_3_4_n54), .B(pe_1_3_4_n51), .S(n48), .Z(
        int_data_x_3__4__3_) );
  MUX2_X1 pe_1_3_4_U100 ( .A(pe_1_3_4_n53), .B(pe_1_3_4_n52), .S(pe_1_3_4_n62), 
        .Z(pe_1_3_4_n54) );
  MUX2_X1 pe_1_3_4_U99 ( .A(pe_1_3_4_int_q_reg_h[23]), .B(
        pe_1_3_4_int_q_reg_h[19]), .S(pe_1_3_4_n56), .Z(pe_1_3_4_n53) );
  MUX2_X1 pe_1_3_4_U98 ( .A(pe_1_3_4_int_q_reg_h[15]), .B(
        pe_1_3_4_int_q_reg_h[11]), .S(pe_1_3_4_n56), .Z(pe_1_3_4_n52) );
  MUX2_X1 pe_1_3_4_U97 ( .A(pe_1_3_4_int_q_reg_h[7]), .B(
        pe_1_3_4_int_q_reg_h[3]), .S(pe_1_3_4_n56), .Z(pe_1_3_4_n51) );
  MUX2_X1 pe_1_3_4_U96 ( .A(pe_1_3_4_n50), .B(pe_1_3_4_n47), .S(n48), .Z(
        int_data_x_3__4__2_) );
  MUX2_X1 pe_1_3_4_U95 ( .A(pe_1_3_4_n49), .B(pe_1_3_4_n48), .S(pe_1_3_4_n62), 
        .Z(pe_1_3_4_n50) );
  MUX2_X1 pe_1_3_4_U94 ( .A(pe_1_3_4_int_q_reg_h[22]), .B(
        pe_1_3_4_int_q_reg_h[18]), .S(pe_1_3_4_n56), .Z(pe_1_3_4_n49) );
  MUX2_X1 pe_1_3_4_U93 ( .A(pe_1_3_4_int_q_reg_h[14]), .B(
        pe_1_3_4_int_q_reg_h[10]), .S(pe_1_3_4_n56), .Z(pe_1_3_4_n48) );
  MUX2_X1 pe_1_3_4_U92 ( .A(pe_1_3_4_int_q_reg_h[6]), .B(
        pe_1_3_4_int_q_reg_h[2]), .S(pe_1_3_4_n56), .Z(pe_1_3_4_n47) );
  MUX2_X1 pe_1_3_4_U91 ( .A(pe_1_3_4_n46), .B(pe_1_3_4_n24), .S(n48), .Z(
        int_data_x_3__4__1_) );
  MUX2_X1 pe_1_3_4_U90 ( .A(pe_1_3_4_n45), .B(pe_1_3_4_n25), .S(pe_1_3_4_n62), 
        .Z(pe_1_3_4_n46) );
  MUX2_X1 pe_1_3_4_U89 ( .A(pe_1_3_4_int_q_reg_h[21]), .B(
        pe_1_3_4_int_q_reg_h[17]), .S(pe_1_3_4_n56), .Z(pe_1_3_4_n45) );
  MUX2_X1 pe_1_3_4_U88 ( .A(pe_1_3_4_int_q_reg_h[13]), .B(
        pe_1_3_4_int_q_reg_h[9]), .S(pe_1_3_4_n56), .Z(pe_1_3_4_n25) );
  MUX2_X1 pe_1_3_4_U87 ( .A(pe_1_3_4_int_q_reg_h[5]), .B(
        pe_1_3_4_int_q_reg_h[1]), .S(pe_1_3_4_n56), .Z(pe_1_3_4_n24) );
  MUX2_X1 pe_1_3_4_U86 ( .A(pe_1_3_4_n23), .B(pe_1_3_4_n20), .S(n48), .Z(
        int_data_x_3__4__0_) );
  MUX2_X1 pe_1_3_4_U85 ( .A(pe_1_3_4_n22), .B(pe_1_3_4_n21), .S(pe_1_3_4_n62), 
        .Z(pe_1_3_4_n23) );
  MUX2_X1 pe_1_3_4_U84 ( .A(pe_1_3_4_int_q_reg_h[20]), .B(
        pe_1_3_4_int_q_reg_h[16]), .S(pe_1_3_4_n56), .Z(pe_1_3_4_n22) );
  MUX2_X1 pe_1_3_4_U83 ( .A(pe_1_3_4_int_q_reg_h[12]), .B(
        pe_1_3_4_int_q_reg_h[8]), .S(pe_1_3_4_n56), .Z(pe_1_3_4_n21) );
  MUX2_X1 pe_1_3_4_U82 ( .A(pe_1_3_4_int_q_reg_h[4]), .B(
        pe_1_3_4_int_q_reg_h[0]), .S(pe_1_3_4_n56), .Z(pe_1_3_4_n20) );
  MUX2_X1 pe_1_3_4_U81 ( .A(pe_1_3_4_n19), .B(pe_1_3_4_n16), .S(n48), .Z(
        int_data_y_3__4__3_) );
  MUX2_X1 pe_1_3_4_U80 ( .A(pe_1_3_4_n18), .B(pe_1_3_4_n17), .S(pe_1_3_4_n62), 
        .Z(pe_1_3_4_n19) );
  MUX2_X1 pe_1_3_4_U79 ( .A(pe_1_3_4_int_q_reg_v[23]), .B(
        pe_1_3_4_int_q_reg_v[19]), .S(pe_1_3_4_n55), .Z(pe_1_3_4_n18) );
  MUX2_X1 pe_1_3_4_U78 ( .A(pe_1_3_4_int_q_reg_v[15]), .B(
        pe_1_3_4_int_q_reg_v[11]), .S(pe_1_3_4_n55), .Z(pe_1_3_4_n17) );
  MUX2_X1 pe_1_3_4_U77 ( .A(pe_1_3_4_int_q_reg_v[7]), .B(
        pe_1_3_4_int_q_reg_v[3]), .S(pe_1_3_4_n55), .Z(pe_1_3_4_n16) );
  MUX2_X1 pe_1_3_4_U76 ( .A(pe_1_3_4_n15), .B(pe_1_3_4_n12), .S(n48), .Z(
        int_data_y_3__4__2_) );
  MUX2_X1 pe_1_3_4_U75 ( .A(pe_1_3_4_n14), .B(pe_1_3_4_n13), .S(pe_1_3_4_n62), 
        .Z(pe_1_3_4_n15) );
  MUX2_X1 pe_1_3_4_U74 ( .A(pe_1_3_4_int_q_reg_v[22]), .B(
        pe_1_3_4_int_q_reg_v[18]), .S(pe_1_3_4_n55), .Z(pe_1_3_4_n14) );
  MUX2_X1 pe_1_3_4_U73 ( .A(pe_1_3_4_int_q_reg_v[14]), .B(
        pe_1_3_4_int_q_reg_v[10]), .S(pe_1_3_4_n55), .Z(pe_1_3_4_n13) );
  MUX2_X1 pe_1_3_4_U72 ( .A(pe_1_3_4_int_q_reg_v[6]), .B(
        pe_1_3_4_int_q_reg_v[2]), .S(pe_1_3_4_n55), .Z(pe_1_3_4_n12) );
  MUX2_X1 pe_1_3_4_U71 ( .A(pe_1_3_4_n11), .B(pe_1_3_4_n8), .S(n48), .Z(
        int_data_y_3__4__1_) );
  MUX2_X1 pe_1_3_4_U70 ( .A(pe_1_3_4_n10), .B(pe_1_3_4_n9), .S(pe_1_3_4_n62), 
        .Z(pe_1_3_4_n11) );
  MUX2_X1 pe_1_3_4_U69 ( .A(pe_1_3_4_int_q_reg_v[21]), .B(
        pe_1_3_4_int_q_reg_v[17]), .S(pe_1_3_4_n55), .Z(pe_1_3_4_n10) );
  MUX2_X1 pe_1_3_4_U68 ( .A(pe_1_3_4_int_q_reg_v[13]), .B(
        pe_1_3_4_int_q_reg_v[9]), .S(pe_1_3_4_n55), .Z(pe_1_3_4_n9) );
  MUX2_X1 pe_1_3_4_U67 ( .A(pe_1_3_4_int_q_reg_v[5]), .B(
        pe_1_3_4_int_q_reg_v[1]), .S(pe_1_3_4_n55), .Z(pe_1_3_4_n8) );
  MUX2_X1 pe_1_3_4_U66 ( .A(pe_1_3_4_n7), .B(pe_1_3_4_n4), .S(n48), .Z(
        int_data_y_3__4__0_) );
  MUX2_X1 pe_1_3_4_U65 ( .A(pe_1_3_4_n6), .B(pe_1_3_4_n5), .S(pe_1_3_4_n62), 
        .Z(pe_1_3_4_n7) );
  MUX2_X1 pe_1_3_4_U64 ( .A(pe_1_3_4_int_q_reg_v[20]), .B(
        pe_1_3_4_int_q_reg_v[16]), .S(pe_1_3_4_n55), .Z(pe_1_3_4_n6) );
  MUX2_X1 pe_1_3_4_U63 ( .A(pe_1_3_4_int_q_reg_v[12]), .B(
        pe_1_3_4_int_q_reg_v[8]), .S(pe_1_3_4_n55), .Z(pe_1_3_4_n5) );
  MUX2_X1 pe_1_3_4_U62 ( .A(pe_1_3_4_int_q_reg_v[4]), .B(
        pe_1_3_4_int_q_reg_v[0]), .S(pe_1_3_4_n55), .Z(pe_1_3_4_n4) );
  AOI222_X1 pe_1_3_4_U61 ( .A1(int_data_res_4__4__2_), .A2(pe_1_3_4_n64), .B1(
        pe_1_3_4_N80), .B2(pe_1_3_4_n27), .C1(pe_1_3_4_N72), .C2(pe_1_3_4_n28), 
        .ZN(pe_1_3_4_n33) );
  INV_X1 pe_1_3_4_U60 ( .A(pe_1_3_4_n33), .ZN(pe_1_3_4_n82) );
  AOI222_X1 pe_1_3_4_U59 ( .A1(int_data_res_4__4__6_), .A2(pe_1_3_4_n64), .B1(
        pe_1_3_4_N84), .B2(pe_1_3_4_n27), .C1(pe_1_3_4_N76), .C2(pe_1_3_4_n28), 
        .ZN(pe_1_3_4_n29) );
  INV_X1 pe_1_3_4_U58 ( .A(pe_1_3_4_n29), .ZN(pe_1_3_4_n78) );
  XNOR2_X1 pe_1_3_4_U57 ( .A(pe_1_3_4_n73), .B(int_data_res_3__4__0_), .ZN(
        pe_1_3_4_N70) );
  AOI222_X1 pe_1_3_4_U52 ( .A1(int_data_res_4__4__0_), .A2(pe_1_3_4_n64), .B1(
        pe_1_3_4_n1), .B2(pe_1_3_4_n27), .C1(pe_1_3_4_N70), .C2(pe_1_3_4_n28), 
        .ZN(pe_1_3_4_n35) );
  INV_X1 pe_1_3_4_U51 ( .A(pe_1_3_4_n35), .ZN(pe_1_3_4_n84) );
  AOI222_X1 pe_1_3_4_U50 ( .A1(int_data_res_4__4__1_), .A2(pe_1_3_4_n64), .B1(
        pe_1_3_4_N79), .B2(pe_1_3_4_n27), .C1(pe_1_3_4_N71), .C2(pe_1_3_4_n28), 
        .ZN(pe_1_3_4_n34) );
  INV_X1 pe_1_3_4_U49 ( .A(pe_1_3_4_n34), .ZN(pe_1_3_4_n83) );
  AOI222_X1 pe_1_3_4_U48 ( .A1(int_data_res_4__4__3_), .A2(pe_1_3_4_n64), .B1(
        pe_1_3_4_N81), .B2(pe_1_3_4_n27), .C1(pe_1_3_4_N73), .C2(pe_1_3_4_n28), 
        .ZN(pe_1_3_4_n32) );
  INV_X1 pe_1_3_4_U47 ( .A(pe_1_3_4_n32), .ZN(pe_1_3_4_n81) );
  AOI222_X1 pe_1_3_4_U46 ( .A1(int_data_res_4__4__4_), .A2(pe_1_3_4_n64), .B1(
        pe_1_3_4_N82), .B2(pe_1_3_4_n27), .C1(pe_1_3_4_N74), .C2(pe_1_3_4_n28), 
        .ZN(pe_1_3_4_n31) );
  INV_X1 pe_1_3_4_U45 ( .A(pe_1_3_4_n31), .ZN(pe_1_3_4_n80) );
  AOI222_X1 pe_1_3_4_U44 ( .A1(int_data_res_4__4__5_), .A2(pe_1_3_4_n64), .B1(
        pe_1_3_4_N83), .B2(pe_1_3_4_n27), .C1(pe_1_3_4_N75), .C2(pe_1_3_4_n28), 
        .ZN(pe_1_3_4_n30) );
  INV_X1 pe_1_3_4_U43 ( .A(pe_1_3_4_n30), .ZN(pe_1_3_4_n79) );
  NAND2_X1 pe_1_3_4_U42 ( .A1(pe_1_3_4_int_data_0_), .A2(pe_1_3_4_n3), .ZN(
        pe_1_3_4_sub_81_carry[1]) );
  INV_X1 pe_1_3_4_U41 ( .A(pe_1_3_4_int_data_1_), .ZN(pe_1_3_4_n74) );
  INV_X1 pe_1_3_4_U40 ( .A(pe_1_3_4_int_data_2_), .ZN(pe_1_3_4_n75) );
  AND2_X1 pe_1_3_4_U39 ( .A1(pe_1_3_4_int_data_0_), .A2(int_data_res_3__4__0_), 
        .ZN(pe_1_3_4_n2) );
  AOI222_X1 pe_1_3_4_U38 ( .A1(pe_1_3_4_n64), .A2(int_data_res_4__4__7_), .B1(
        pe_1_3_4_N85), .B2(pe_1_3_4_n27), .C1(pe_1_3_4_N77), .C2(pe_1_3_4_n28), 
        .ZN(pe_1_3_4_n26) );
  INV_X1 pe_1_3_4_U37 ( .A(pe_1_3_4_n26), .ZN(pe_1_3_4_n77) );
  NOR3_X1 pe_1_3_4_U36 ( .A1(pe_1_3_4_n59), .A2(pe_1_3_4_n65), .A3(int_ckg[35]), .ZN(pe_1_3_4_n36) );
  OR2_X1 pe_1_3_4_U35 ( .A1(pe_1_3_4_n36), .A2(pe_1_3_4_n64), .ZN(pe_1_3_4_N90) );
  INV_X1 pe_1_3_4_U34 ( .A(n39), .ZN(pe_1_3_4_n63) );
  AND2_X1 pe_1_3_4_U33 ( .A1(int_data_x_3__4__2_), .A2(pe_1_3_4_n58), .ZN(
        pe_1_3_4_int_data_2_) );
  AND2_X1 pe_1_3_4_U32 ( .A1(int_data_x_3__4__1_), .A2(pe_1_3_4_n58), .ZN(
        pe_1_3_4_int_data_1_) );
  AND2_X1 pe_1_3_4_U31 ( .A1(int_data_x_3__4__3_), .A2(pe_1_3_4_n58), .ZN(
        pe_1_3_4_int_data_3_) );
  BUF_X1 pe_1_3_4_U30 ( .A(n61), .Z(pe_1_3_4_n64) );
  INV_X1 pe_1_3_4_U29 ( .A(n33), .ZN(pe_1_3_4_n61) );
  AND2_X1 pe_1_3_4_U28 ( .A1(int_data_x_3__4__0_), .A2(pe_1_3_4_n58), .ZN(
        pe_1_3_4_int_data_0_) );
  NAND2_X1 pe_1_3_4_U27 ( .A1(pe_1_3_4_n44), .A2(pe_1_3_4_n61), .ZN(
        pe_1_3_4_n41) );
  AND3_X1 pe_1_3_4_U26 ( .A1(n75), .A2(pe_1_3_4_n63), .A3(n48), .ZN(
        pe_1_3_4_n44) );
  INV_X1 pe_1_3_4_U25 ( .A(pe_1_3_4_int_data_3_), .ZN(pe_1_3_4_n76) );
  NOR2_X1 pe_1_3_4_U24 ( .A1(pe_1_3_4_n70), .A2(n48), .ZN(pe_1_3_4_n43) );
  NOR2_X1 pe_1_3_4_U23 ( .A1(pe_1_3_4_n57), .A2(pe_1_3_4_n64), .ZN(
        pe_1_3_4_n28) );
  NOR2_X1 pe_1_3_4_U22 ( .A1(n19), .A2(pe_1_3_4_n64), .ZN(pe_1_3_4_n27) );
  INV_X1 pe_1_3_4_U21 ( .A(pe_1_3_4_int_data_0_), .ZN(pe_1_3_4_n73) );
  INV_X1 pe_1_3_4_U20 ( .A(pe_1_3_4_n41), .ZN(pe_1_3_4_n90) );
  INV_X1 pe_1_3_4_U19 ( .A(pe_1_3_4_n37), .ZN(pe_1_3_4_n88) );
  INV_X1 pe_1_3_4_U18 ( .A(pe_1_3_4_n38), .ZN(pe_1_3_4_n87) );
  INV_X1 pe_1_3_4_U17 ( .A(pe_1_3_4_n39), .ZN(pe_1_3_4_n86) );
  NOR2_X1 pe_1_3_4_U16 ( .A1(pe_1_3_4_n68), .A2(pe_1_3_4_n42), .ZN(
        pe_1_3_4_N59) );
  NOR2_X1 pe_1_3_4_U15 ( .A1(pe_1_3_4_n68), .A2(pe_1_3_4_n41), .ZN(
        pe_1_3_4_N60) );
  NOR2_X1 pe_1_3_4_U14 ( .A1(pe_1_3_4_n68), .A2(pe_1_3_4_n38), .ZN(
        pe_1_3_4_N63) );
  NOR2_X1 pe_1_3_4_U13 ( .A1(pe_1_3_4_n67), .A2(pe_1_3_4_n40), .ZN(
        pe_1_3_4_N61) );
  NOR2_X1 pe_1_3_4_U12 ( .A1(pe_1_3_4_n67), .A2(pe_1_3_4_n39), .ZN(
        pe_1_3_4_N62) );
  NOR2_X1 pe_1_3_4_U11 ( .A1(pe_1_3_4_n37), .A2(pe_1_3_4_n67), .ZN(
        pe_1_3_4_N64) );
  NAND2_X1 pe_1_3_4_U10 ( .A1(pe_1_3_4_n44), .A2(pe_1_3_4_n60), .ZN(
        pe_1_3_4_n42) );
  BUF_X1 pe_1_3_4_U9 ( .A(pe_1_3_4_n60), .Z(pe_1_3_4_n55) );
  INV_X1 pe_1_3_4_U8 ( .A(pe_1_3_4_n69), .ZN(pe_1_3_4_n65) );
  BUF_X1 pe_1_3_4_U7 ( .A(pe_1_3_4_n60), .Z(pe_1_3_4_n56) );
  INV_X1 pe_1_3_4_U6 ( .A(pe_1_3_4_n42), .ZN(pe_1_3_4_n89) );
  INV_X1 pe_1_3_4_U5 ( .A(pe_1_3_4_n40), .ZN(pe_1_3_4_n85) );
  INV_X2 pe_1_3_4_U4 ( .A(n83), .ZN(pe_1_3_4_n72) );
  XOR2_X1 pe_1_3_4_U3 ( .A(pe_1_3_4_int_data_0_), .B(int_data_res_3__4__0_), 
        .Z(pe_1_3_4_n1) );
  DFFR_X1 pe_1_3_4_int_q_acc_reg_0_ ( .D(pe_1_3_4_n84), .CK(pe_1_3_4_net5368), 
        .RN(pe_1_3_4_n72), .Q(int_data_res_3__4__0_), .QN(pe_1_3_4_n3) );
  DFFR_X1 pe_1_3_4_int_q_reg_v_reg_0__0_ ( .D(int_data_y_4__4__0_), .CK(
        pe_1_3_4_net5338), .RN(pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_v[20]) );
  DFFR_X1 pe_1_3_4_int_q_reg_v_reg_0__1_ ( .D(int_data_y_4__4__1_), .CK(
        pe_1_3_4_net5338), .RN(pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_v[21]) );
  DFFR_X1 pe_1_3_4_int_q_reg_v_reg_0__2_ ( .D(int_data_y_4__4__2_), .CK(
        pe_1_3_4_net5338), .RN(pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_v[22]) );
  DFFR_X1 pe_1_3_4_int_q_reg_v_reg_0__3_ ( .D(int_data_y_4__4__3_), .CK(
        pe_1_3_4_net5338), .RN(pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_v[23]) );
  DFFR_X1 pe_1_3_4_int_q_reg_v_reg_1__0_ ( .D(int_data_y_4__4__0_), .CK(
        pe_1_3_4_net5343), .RN(pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_v[16]) );
  DFFR_X1 pe_1_3_4_int_q_reg_v_reg_1__1_ ( .D(int_data_y_4__4__1_), .CK(
        pe_1_3_4_net5343), .RN(pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_v[17]) );
  DFFR_X1 pe_1_3_4_int_q_reg_v_reg_1__2_ ( .D(int_data_y_4__4__2_), .CK(
        pe_1_3_4_net5343), .RN(pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_v[18]) );
  DFFR_X1 pe_1_3_4_int_q_reg_v_reg_1__3_ ( .D(int_data_y_4__4__3_), .CK(
        pe_1_3_4_net5343), .RN(pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_v[19]) );
  DFFR_X1 pe_1_3_4_int_q_reg_v_reg_2__0_ ( .D(int_data_y_4__4__0_), .CK(
        pe_1_3_4_net5348), .RN(pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_v[12]) );
  DFFR_X1 pe_1_3_4_int_q_reg_v_reg_2__1_ ( .D(int_data_y_4__4__1_), .CK(
        pe_1_3_4_net5348), .RN(pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_v[13]) );
  DFFR_X1 pe_1_3_4_int_q_reg_v_reg_2__2_ ( .D(int_data_y_4__4__2_), .CK(
        pe_1_3_4_net5348), .RN(pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_v[14]) );
  DFFR_X1 pe_1_3_4_int_q_reg_v_reg_2__3_ ( .D(int_data_y_4__4__3_), .CK(
        pe_1_3_4_net5348), .RN(pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_v[15]) );
  DFFR_X1 pe_1_3_4_int_q_reg_v_reg_3__0_ ( .D(int_data_y_4__4__0_), .CK(
        pe_1_3_4_net5353), .RN(pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_v[8]) );
  DFFR_X1 pe_1_3_4_int_q_reg_v_reg_3__1_ ( .D(int_data_y_4__4__1_), .CK(
        pe_1_3_4_net5353), .RN(pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_v[9]) );
  DFFR_X1 pe_1_3_4_int_q_reg_v_reg_3__2_ ( .D(int_data_y_4__4__2_), .CK(
        pe_1_3_4_net5353), .RN(pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_v[10]) );
  DFFR_X1 pe_1_3_4_int_q_reg_v_reg_3__3_ ( .D(int_data_y_4__4__3_), .CK(
        pe_1_3_4_net5353), .RN(pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_v[11]) );
  DFFR_X1 pe_1_3_4_int_q_reg_v_reg_4__0_ ( .D(int_data_y_4__4__0_), .CK(
        pe_1_3_4_net5358), .RN(pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_v[4]) );
  DFFR_X1 pe_1_3_4_int_q_reg_v_reg_4__1_ ( .D(int_data_y_4__4__1_), .CK(
        pe_1_3_4_net5358), .RN(pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_v[5]) );
  DFFR_X1 pe_1_3_4_int_q_reg_v_reg_4__2_ ( .D(int_data_y_4__4__2_), .CK(
        pe_1_3_4_net5358), .RN(pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_v[6]) );
  DFFR_X1 pe_1_3_4_int_q_reg_v_reg_4__3_ ( .D(int_data_y_4__4__3_), .CK(
        pe_1_3_4_net5358), .RN(pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_v[7]) );
  DFFR_X1 pe_1_3_4_int_q_reg_v_reg_5__0_ ( .D(int_data_y_4__4__0_), .CK(
        pe_1_3_4_net5363), .RN(pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_v[0]) );
  DFFR_X1 pe_1_3_4_int_q_reg_v_reg_5__1_ ( .D(int_data_y_4__4__1_), .CK(
        pe_1_3_4_net5363), .RN(pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_v[1]) );
  DFFR_X1 pe_1_3_4_int_q_reg_v_reg_5__2_ ( .D(int_data_y_4__4__2_), .CK(
        pe_1_3_4_net5363), .RN(pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_v[2]) );
  DFFR_X1 pe_1_3_4_int_q_reg_v_reg_5__3_ ( .D(int_data_y_4__4__3_), .CK(
        pe_1_3_4_net5363), .RN(pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_3_4_int_q_reg_h_reg_0__0_ ( .D(int_data_x_3__5__0_), .SI(
        int_data_y_4__4__0_), .SE(pe_1_3_4_n65), .CK(pe_1_3_4_net5307), .RN(
        pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_3_4_int_q_reg_h_reg_0__1_ ( .D(int_data_x_3__5__1_), .SI(
        int_data_y_4__4__1_), .SE(pe_1_3_4_n65), .CK(pe_1_3_4_net5307), .RN(
        pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_3_4_int_q_reg_h_reg_0__2_ ( .D(int_data_x_3__5__2_), .SI(
        int_data_y_4__4__2_), .SE(pe_1_3_4_n65), .CK(pe_1_3_4_net5307), .RN(
        pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_3_4_int_q_reg_h_reg_0__3_ ( .D(int_data_x_3__5__3_), .SI(
        int_data_y_4__4__3_), .SE(pe_1_3_4_n65), .CK(pe_1_3_4_net5307), .RN(
        pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_3_4_int_q_reg_h_reg_1__0_ ( .D(int_data_x_3__5__0_), .SI(
        int_data_y_4__4__0_), .SE(pe_1_3_4_n65), .CK(pe_1_3_4_net5313), .RN(
        pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_3_4_int_q_reg_h_reg_1__1_ ( .D(int_data_x_3__5__1_), .SI(
        int_data_y_4__4__1_), .SE(pe_1_3_4_n65), .CK(pe_1_3_4_net5313), .RN(
        pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_3_4_int_q_reg_h_reg_1__2_ ( .D(int_data_x_3__5__2_), .SI(
        int_data_y_4__4__2_), .SE(pe_1_3_4_n65), .CK(pe_1_3_4_net5313), .RN(
        pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_3_4_int_q_reg_h_reg_1__3_ ( .D(int_data_x_3__5__3_), .SI(
        int_data_y_4__4__3_), .SE(pe_1_3_4_n65), .CK(pe_1_3_4_net5313), .RN(
        pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_3_4_int_q_reg_h_reg_2__0_ ( .D(int_data_x_3__5__0_), .SI(
        int_data_y_4__4__0_), .SE(pe_1_3_4_n65), .CK(pe_1_3_4_net5318), .RN(
        pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_3_4_int_q_reg_h_reg_2__1_ ( .D(int_data_x_3__5__1_), .SI(
        int_data_y_4__4__1_), .SE(pe_1_3_4_n65), .CK(pe_1_3_4_net5318), .RN(
        pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_3_4_int_q_reg_h_reg_2__2_ ( .D(int_data_x_3__5__2_), .SI(
        int_data_y_4__4__2_), .SE(pe_1_3_4_n65), .CK(pe_1_3_4_net5318), .RN(
        pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_3_4_int_q_reg_h_reg_2__3_ ( .D(int_data_x_3__5__3_), .SI(
        int_data_y_4__4__3_), .SE(pe_1_3_4_n65), .CK(pe_1_3_4_net5318), .RN(
        pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_3_4_int_q_reg_h_reg_3__0_ ( .D(int_data_x_3__5__0_), .SI(
        int_data_y_4__4__0_), .SE(pe_1_3_4_n65), .CK(pe_1_3_4_net5323), .RN(
        pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_3_4_int_q_reg_h_reg_3__1_ ( .D(int_data_x_3__5__1_), .SI(
        int_data_y_4__4__1_), .SE(pe_1_3_4_n65), .CK(pe_1_3_4_net5323), .RN(
        pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_3_4_int_q_reg_h_reg_3__2_ ( .D(int_data_x_3__5__2_), .SI(
        int_data_y_4__4__2_), .SE(pe_1_3_4_n65), .CK(pe_1_3_4_net5323), .RN(
        pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_3_4_int_q_reg_h_reg_3__3_ ( .D(int_data_x_3__5__3_), .SI(
        int_data_y_4__4__3_), .SE(pe_1_3_4_n65), .CK(pe_1_3_4_net5323), .RN(
        pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_3_4_int_q_reg_h_reg_4__0_ ( .D(int_data_x_3__5__0_), .SI(
        int_data_y_4__4__0_), .SE(pe_1_3_4_n66), .CK(pe_1_3_4_net5328), .RN(
        pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_3_4_int_q_reg_h_reg_4__1_ ( .D(int_data_x_3__5__1_), .SI(
        int_data_y_4__4__1_), .SE(pe_1_3_4_n66), .CK(pe_1_3_4_net5328), .RN(
        pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_3_4_int_q_reg_h_reg_4__2_ ( .D(int_data_x_3__5__2_), .SI(
        int_data_y_4__4__2_), .SE(pe_1_3_4_n66), .CK(pe_1_3_4_net5328), .RN(
        pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_3_4_int_q_reg_h_reg_4__3_ ( .D(int_data_x_3__5__3_), .SI(
        int_data_y_4__4__3_), .SE(pe_1_3_4_n66), .CK(pe_1_3_4_net5328), .RN(
        pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_3_4_int_q_reg_h_reg_5__0_ ( .D(int_data_x_3__5__0_), .SI(
        int_data_y_4__4__0_), .SE(pe_1_3_4_n66), .CK(pe_1_3_4_net5333), .RN(
        pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_3_4_int_q_reg_h_reg_5__1_ ( .D(int_data_x_3__5__1_), .SI(
        int_data_y_4__4__1_), .SE(pe_1_3_4_n66), .CK(pe_1_3_4_net5333), .RN(
        pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_3_4_int_q_reg_h_reg_5__2_ ( .D(int_data_x_3__5__2_), .SI(
        int_data_y_4__4__2_), .SE(pe_1_3_4_n66), .CK(pe_1_3_4_net5333), .RN(
        pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_3_4_int_q_reg_h_reg_5__3_ ( .D(int_data_x_3__5__3_), .SI(
        int_data_y_4__4__3_), .SE(pe_1_3_4_n66), .CK(pe_1_3_4_net5333), .RN(
        pe_1_3_4_n72), .Q(pe_1_3_4_int_q_reg_h[3]) );
  FA_X1 pe_1_3_4_sub_81_U2_7 ( .A(int_data_res_3__4__7_), .B(pe_1_3_4_n76), 
        .CI(pe_1_3_4_sub_81_carry[7]), .S(pe_1_3_4_N77) );
  FA_X1 pe_1_3_4_sub_81_U2_6 ( .A(int_data_res_3__4__6_), .B(pe_1_3_4_n76), 
        .CI(pe_1_3_4_sub_81_carry[6]), .CO(pe_1_3_4_sub_81_carry[7]), .S(
        pe_1_3_4_N76) );
  FA_X1 pe_1_3_4_sub_81_U2_5 ( .A(int_data_res_3__4__5_), .B(pe_1_3_4_n76), 
        .CI(pe_1_3_4_sub_81_carry[5]), .CO(pe_1_3_4_sub_81_carry[6]), .S(
        pe_1_3_4_N75) );
  FA_X1 pe_1_3_4_sub_81_U2_4 ( .A(int_data_res_3__4__4_), .B(pe_1_3_4_n76), 
        .CI(pe_1_3_4_sub_81_carry[4]), .CO(pe_1_3_4_sub_81_carry[5]), .S(
        pe_1_3_4_N74) );
  FA_X1 pe_1_3_4_sub_81_U2_3 ( .A(int_data_res_3__4__3_), .B(pe_1_3_4_n76), 
        .CI(pe_1_3_4_sub_81_carry[3]), .CO(pe_1_3_4_sub_81_carry[4]), .S(
        pe_1_3_4_N73) );
  FA_X1 pe_1_3_4_sub_81_U2_2 ( .A(int_data_res_3__4__2_), .B(pe_1_3_4_n75), 
        .CI(pe_1_3_4_sub_81_carry[2]), .CO(pe_1_3_4_sub_81_carry[3]), .S(
        pe_1_3_4_N72) );
  FA_X1 pe_1_3_4_sub_81_U2_1 ( .A(int_data_res_3__4__1_), .B(pe_1_3_4_n74), 
        .CI(pe_1_3_4_sub_81_carry[1]), .CO(pe_1_3_4_sub_81_carry[2]), .S(
        pe_1_3_4_N71) );
  FA_X1 pe_1_3_4_add_83_U1_7 ( .A(int_data_res_3__4__7_), .B(
        pe_1_3_4_int_data_3_), .CI(pe_1_3_4_add_83_carry[7]), .S(pe_1_3_4_N85)
         );
  FA_X1 pe_1_3_4_add_83_U1_6 ( .A(int_data_res_3__4__6_), .B(
        pe_1_3_4_int_data_3_), .CI(pe_1_3_4_add_83_carry[6]), .CO(
        pe_1_3_4_add_83_carry[7]), .S(pe_1_3_4_N84) );
  FA_X1 pe_1_3_4_add_83_U1_5 ( .A(int_data_res_3__4__5_), .B(
        pe_1_3_4_int_data_3_), .CI(pe_1_3_4_add_83_carry[5]), .CO(
        pe_1_3_4_add_83_carry[6]), .S(pe_1_3_4_N83) );
  FA_X1 pe_1_3_4_add_83_U1_4 ( .A(int_data_res_3__4__4_), .B(
        pe_1_3_4_int_data_3_), .CI(pe_1_3_4_add_83_carry[4]), .CO(
        pe_1_3_4_add_83_carry[5]), .S(pe_1_3_4_N82) );
  FA_X1 pe_1_3_4_add_83_U1_3 ( .A(int_data_res_3__4__3_), .B(
        pe_1_3_4_int_data_3_), .CI(pe_1_3_4_add_83_carry[3]), .CO(
        pe_1_3_4_add_83_carry[4]), .S(pe_1_3_4_N81) );
  FA_X1 pe_1_3_4_add_83_U1_2 ( .A(int_data_res_3__4__2_), .B(
        pe_1_3_4_int_data_2_), .CI(pe_1_3_4_add_83_carry[2]), .CO(
        pe_1_3_4_add_83_carry[3]), .S(pe_1_3_4_N80) );
  FA_X1 pe_1_3_4_add_83_U1_1 ( .A(int_data_res_3__4__1_), .B(
        pe_1_3_4_int_data_1_), .CI(pe_1_3_4_n2), .CO(pe_1_3_4_add_83_carry[2]), 
        .S(pe_1_3_4_N79) );
  NAND3_X1 pe_1_3_4_U56 ( .A1(pe_1_3_4_n60), .A2(pe_1_3_4_n43), .A3(
        pe_1_3_4_n62), .ZN(pe_1_3_4_n40) );
  NAND3_X1 pe_1_3_4_U55 ( .A1(pe_1_3_4_n43), .A2(pe_1_3_4_n61), .A3(
        pe_1_3_4_n62), .ZN(pe_1_3_4_n39) );
  NAND3_X1 pe_1_3_4_U54 ( .A1(pe_1_3_4_n43), .A2(pe_1_3_4_n63), .A3(
        pe_1_3_4_n60), .ZN(pe_1_3_4_n38) );
  NAND3_X1 pe_1_3_4_U53 ( .A1(pe_1_3_4_n61), .A2(pe_1_3_4_n63), .A3(
        pe_1_3_4_n43), .ZN(pe_1_3_4_n37) );
  DFFR_X1 pe_1_3_4_int_q_acc_reg_6_ ( .D(pe_1_3_4_n78), .CK(pe_1_3_4_net5368), 
        .RN(pe_1_3_4_n71), .Q(int_data_res_3__4__6_) );
  DFFR_X1 pe_1_3_4_int_q_acc_reg_5_ ( .D(pe_1_3_4_n79), .CK(pe_1_3_4_net5368), 
        .RN(pe_1_3_4_n71), .Q(int_data_res_3__4__5_) );
  DFFR_X1 pe_1_3_4_int_q_acc_reg_4_ ( .D(pe_1_3_4_n80), .CK(pe_1_3_4_net5368), 
        .RN(pe_1_3_4_n71), .Q(int_data_res_3__4__4_) );
  DFFR_X1 pe_1_3_4_int_q_acc_reg_3_ ( .D(pe_1_3_4_n81), .CK(pe_1_3_4_net5368), 
        .RN(pe_1_3_4_n71), .Q(int_data_res_3__4__3_) );
  DFFR_X1 pe_1_3_4_int_q_acc_reg_2_ ( .D(pe_1_3_4_n82), .CK(pe_1_3_4_net5368), 
        .RN(pe_1_3_4_n71), .Q(int_data_res_3__4__2_) );
  DFFR_X1 pe_1_3_4_int_q_acc_reg_1_ ( .D(pe_1_3_4_n83), .CK(pe_1_3_4_net5368), 
        .RN(pe_1_3_4_n71), .Q(int_data_res_3__4__1_) );
  DFFR_X1 pe_1_3_4_int_q_acc_reg_7_ ( .D(pe_1_3_4_n77), .CK(pe_1_3_4_net5368), 
        .RN(pe_1_3_4_n71), .Q(int_data_res_3__4__7_) );
  CLKGATETST_X1 pe_1_3_4_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_3_4_n88), .SE(1'b0), .GCK(pe_1_3_4_net5307) );
  CLKGATETST_X1 pe_1_3_4_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_3_4_n87), .SE(1'b0), .GCK(pe_1_3_4_net5313) );
  CLKGATETST_X1 pe_1_3_4_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_3_4_n86), .SE(1'b0), .GCK(pe_1_3_4_net5318) );
  CLKGATETST_X1 pe_1_3_4_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_3_4_n85), .SE(1'b0), .GCK(pe_1_3_4_net5323) );
  CLKGATETST_X1 pe_1_3_4_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_3_4_n90), .SE(1'b0), .GCK(pe_1_3_4_net5328) );
  CLKGATETST_X1 pe_1_3_4_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_3_4_n89), .SE(1'b0), .GCK(pe_1_3_4_net5333) );
  CLKGATETST_X1 pe_1_3_4_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_3_4_N64), .SE(1'b0), .GCK(pe_1_3_4_net5338) );
  CLKGATETST_X1 pe_1_3_4_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_3_4_N63), .SE(1'b0), .GCK(pe_1_3_4_net5343) );
  CLKGATETST_X1 pe_1_3_4_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_3_4_N62), .SE(1'b0), .GCK(pe_1_3_4_net5348) );
  CLKGATETST_X1 pe_1_3_4_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_3_4_N61), .SE(1'b0), .GCK(pe_1_3_4_net5353) );
  CLKGATETST_X1 pe_1_3_4_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_3_4_N60), .SE(1'b0), .GCK(pe_1_3_4_net5358) );
  CLKGATETST_X1 pe_1_3_4_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_3_4_N59), .SE(1'b0), .GCK(pe_1_3_4_net5363) );
  CLKGATETST_X1 pe_1_3_4_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_3_4_N90), .SE(1'b0), .GCK(pe_1_3_4_net5368) );
  CLKBUF_X1 pe_1_3_5_U112 ( .A(pe_1_3_5_n72), .Z(pe_1_3_5_n71) );
  INV_X1 pe_1_3_5_U111 ( .A(n75), .ZN(pe_1_3_5_n70) );
  INV_X1 pe_1_3_5_U110 ( .A(n67), .ZN(pe_1_3_5_n69) );
  INV_X1 pe_1_3_5_U109 ( .A(n67), .ZN(pe_1_3_5_n68) );
  INV_X1 pe_1_3_5_U108 ( .A(n67), .ZN(pe_1_3_5_n67) );
  INV_X1 pe_1_3_5_U107 ( .A(pe_1_3_5_n69), .ZN(pe_1_3_5_n66) );
  INV_X1 pe_1_3_5_U106 ( .A(pe_1_3_5_n63), .ZN(pe_1_3_5_n62) );
  INV_X1 pe_1_3_5_U105 ( .A(pe_1_3_5_n61), .ZN(pe_1_3_5_n60) );
  INV_X1 pe_1_3_5_U104 ( .A(n27), .ZN(pe_1_3_5_n59) );
  INV_X1 pe_1_3_5_U103 ( .A(pe_1_3_5_n59), .ZN(pe_1_3_5_n58) );
  INV_X1 pe_1_3_5_U102 ( .A(n19), .ZN(pe_1_3_5_n57) );
  MUX2_X1 pe_1_3_5_U101 ( .A(pe_1_3_5_n54), .B(pe_1_3_5_n51), .S(n48), .Z(
        int_data_x_3__5__3_) );
  MUX2_X1 pe_1_3_5_U100 ( .A(pe_1_3_5_n53), .B(pe_1_3_5_n52), .S(pe_1_3_5_n62), 
        .Z(pe_1_3_5_n54) );
  MUX2_X1 pe_1_3_5_U99 ( .A(pe_1_3_5_int_q_reg_h[23]), .B(
        pe_1_3_5_int_q_reg_h[19]), .S(pe_1_3_5_n56), .Z(pe_1_3_5_n53) );
  MUX2_X1 pe_1_3_5_U98 ( .A(pe_1_3_5_int_q_reg_h[15]), .B(
        pe_1_3_5_int_q_reg_h[11]), .S(pe_1_3_5_n56), .Z(pe_1_3_5_n52) );
  MUX2_X1 pe_1_3_5_U97 ( .A(pe_1_3_5_int_q_reg_h[7]), .B(
        pe_1_3_5_int_q_reg_h[3]), .S(pe_1_3_5_n56), .Z(pe_1_3_5_n51) );
  MUX2_X1 pe_1_3_5_U96 ( .A(pe_1_3_5_n50), .B(pe_1_3_5_n47), .S(n48), .Z(
        int_data_x_3__5__2_) );
  MUX2_X1 pe_1_3_5_U95 ( .A(pe_1_3_5_n49), .B(pe_1_3_5_n48), .S(pe_1_3_5_n62), 
        .Z(pe_1_3_5_n50) );
  MUX2_X1 pe_1_3_5_U94 ( .A(pe_1_3_5_int_q_reg_h[22]), .B(
        pe_1_3_5_int_q_reg_h[18]), .S(pe_1_3_5_n56), .Z(pe_1_3_5_n49) );
  MUX2_X1 pe_1_3_5_U93 ( .A(pe_1_3_5_int_q_reg_h[14]), .B(
        pe_1_3_5_int_q_reg_h[10]), .S(pe_1_3_5_n56), .Z(pe_1_3_5_n48) );
  MUX2_X1 pe_1_3_5_U92 ( .A(pe_1_3_5_int_q_reg_h[6]), .B(
        pe_1_3_5_int_q_reg_h[2]), .S(pe_1_3_5_n56), .Z(pe_1_3_5_n47) );
  MUX2_X1 pe_1_3_5_U91 ( .A(pe_1_3_5_n46), .B(pe_1_3_5_n24), .S(n48), .Z(
        int_data_x_3__5__1_) );
  MUX2_X1 pe_1_3_5_U90 ( .A(pe_1_3_5_n45), .B(pe_1_3_5_n25), .S(pe_1_3_5_n62), 
        .Z(pe_1_3_5_n46) );
  MUX2_X1 pe_1_3_5_U89 ( .A(pe_1_3_5_int_q_reg_h[21]), .B(
        pe_1_3_5_int_q_reg_h[17]), .S(pe_1_3_5_n56), .Z(pe_1_3_5_n45) );
  MUX2_X1 pe_1_3_5_U88 ( .A(pe_1_3_5_int_q_reg_h[13]), .B(
        pe_1_3_5_int_q_reg_h[9]), .S(pe_1_3_5_n56), .Z(pe_1_3_5_n25) );
  MUX2_X1 pe_1_3_5_U87 ( .A(pe_1_3_5_int_q_reg_h[5]), .B(
        pe_1_3_5_int_q_reg_h[1]), .S(pe_1_3_5_n56), .Z(pe_1_3_5_n24) );
  MUX2_X1 pe_1_3_5_U86 ( .A(pe_1_3_5_n23), .B(pe_1_3_5_n20), .S(n48), .Z(
        int_data_x_3__5__0_) );
  MUX2_X1 pe_1_3_5_U85 ( .A(pe_1_3_5_n22), .B(pe_1_3_5_n21), .S(pe_1_3_5_n62), 
        .Z(pe_1_3_5_n23) );
  MUX2_X1 pe_1_3_5_U84 ( .A(pe_1_3_5_int_q_reg_h[20]), .B(
        pe_1_3_5_int_q_reg_h[16]), .S(pe_1_3_5_n56), .Z(pe_1_3_5_n22) );
  MUX2_X1 pe_1_3_5_U83 ( .A(pe_1_3_5_int_q_reg_h[12]), .B(
        pe_1_3_5_int_q_reg_h[8]), .S(pe_1_3_5_n56), .Z(pe_1_3_5_n21) );
  MUX2_X1 pe_1_3_5_U82 ( .A(pe_1_3_5_int_q_reg_h[4]), .B(
        pe_1_3_5_int_q_reg_h[0]), .S(pe_1_3_5_n56), .Z(pe_1_3_5_n20) );
  MUX2_X1 pe_1_3_5_U81 ( .A(pe_1_3_5_n19), .B(pe_1_3_5_n16), .S(n48), .Z(
        int_data_y_3__5__3_) );
  MUX2_X1 pe_1_3_5_U80 ( .A(pe_1_3_5_n18), .B(pe_1_3_5_n17), .S(pe_1_3_5_n62), 
        .Z(pe_1_3_5_n19) );
  MUX2_X1 pe_1_3_5_U79 ( .A(pe_1_3_5_int_q_reg_v[23]), .B(
        pe_1_3_5_int_q_reg_v[19]), .S(pe_1_3_5_n55), .Z(pe_1_3_5_n18) );
  MUX2_X1 pe_1_3_5_U78 ( .A(pe_1_3_5_int_q_reg_v[15]), .B(
        pe_1_3_5_int_q_reg_v[11]), .S(pe_1_3_5_n55), .Z(pe_1_3_5_n17) );
  MUX2_X1 pe_1_3_5_U77 ( .A(pe_1_3_5_int_q_reg_v[7]), .B(
        pe_1_3_5_int_q_reg_v[3]), .S(pe_1_3_5_n55), .Z(pe_1_3_5_n16) );
  MUX2_X1 pe_1_3_5_U76 ( .A(pe_1_3_5_n15), .B(pe_1_3_5_n12), .S(n48), .Z(
        int_data_y_3__5__2_) );
  MUX2_X1 pe_1_3_5_U75 ( .A(pe_1_3_5_n14), .B(pe_1_3_5_n13), .S(pe_1_3_5_n62), 
        .Z(pe_1_3_5_n15) );
  MUX2_X1 pe_1_3_5_U74 ( .A(pe_1_3_5_int_q_reg_v[22]), .B(
        pe_1_3_5_int_q_reg_v[18]), .S(pe_1_3_5_n55), .Z(pe_1_3_5_n14) );
  MUX2_X1 pe_1_3_5_U73 ( .A(pe_1_3_5_int_q_reg_v[14]), .B(
        pe_1_3_5_int_q_reg_v[10]), .S(pe_1_3_5_n55), .Z(pe_1_3_5_n13) );
  MUX2_X1 pe_1_3_5_U72 ( .A(pe_1_3_5_int_q_reg_v[6]), .B(
        pe_1_3_5_int_q_reg_v[2]), .S(pe_1_3_5_n55), .Z(pe_1_3_5_n12) );
  MUX2_X1 pe_1_3_5_U71 ( .A(pe_1_3_5_n11), .B(pe_1_3_5_n8), .S(n48), .Z(
        int_data_y_3__5__1_) );
  MUX2_X1 pe_1_3_5_U70 ( .A(pe_1_3_5_n10), .B(pe_1_3_5_n9), .S(pe_1_3_5_n62), 
        .Z(pe_1_3_5_n11) );
  MUX2_X1 pe_1_3_5_U69 ( .A(pe_1_3_5_int_q_reg_v[21]), .B(
        pe_1_3_5_int_q_reg_v[17]), .S(pe_1_3_5_n55), .Z(pe_1_3_5_n10) );
  MUX2_X1 pe_1_3_5_U68 ( .A(pe_1_3_5_int_q_reg_v[13]), .B(
        pe_1_3_5_int_q_reg_v[9]), .S(pe_1_3_5_n55), .Z(pe_1_3_5_n9) );
  MUX2_X1 pe_1_3_5_U67 ( .A(pe_1_3_5_int_q_reg_v[5]), .B(
        pe_1_3_5_int_q_reg_v[1]), .S(pe_1_3_5_n55), .Z(pe_1_3_5_n8) );
  MUX2_X1 pe_1_3_5_U66 ( .A(pe_1_3_5_n7), .B(pe_1_3_5_n4), .S(n48), .Z(
        int_data_y_3__5__0_) );
  MUX2_X1 pe_1_3_5_U65 ( .A(pe_1_3_5_n6), .B(pe_1_3_5_n5), .S(pe_1_3_5_n62), 
        .Z(pe_1_3_5_n7) );
  MUX2_X1 pe_1_3_5_U64 ( .A(pe_1_3_5_int_q_reg_v[20]), .B(
        pe_1_3_5_int_q_reg_v[16]), .S(pe_1_3_5_n55), .Z(pe_1_3_5_n6) );
  MUX2_X1 pe_1_3_5_U63 ( .A(pe_1_3_5_int_q_reg_v[12]), .B(
        pe_1_3_5_int_q_reg_v[8]), .S(pe_1_3_5_n55), .Z(pe_1_3_5_n5) );
  MUX2_X1 pe_1_3_5_U62 ( .A(pe_1_3_5_int_q_reg_v[4]), .B(
        pe_1_3_5_int_q_reg_v[0]), .S(pe_1_3_5_n55), .Z(pe_1_3_5_n4) );
  AOI222_X1 pe_1_3_5_U61 ( .A1(int_data_res_4__5__2_), .A2(pe_1_3_5_n64), .B1(
        pe_1_3_5_N80), .B2(pe_1_3_5_n27), .C1(pe_1_3_5_N72), .C2(pe_1_3_5_n28), 
        .ZN(pe_1_3_5_n33) );
  INV_X1 pe_1_3_5_U60 ( .A(pe_1_3_5_n33), .ZN(pe_1_3_5_n82) );
  AOI222_X1 pe_1_3_5_U59 ( .A1(int_data_res_4__5__6_), .A2(pe_1_3_5_n64), .B1(
        pe_1_3_5_N84), .B2(pe_1_3_5_n27), .C1(pe_1_3_5_N76), .C2(pe_1_3_5_n28), 
        .ZN(pe_1_3_5_n29) );
  INV_X1 pe_1_3_5_U58 ( .A(pe_1_3_5_n29), .ZN(pe_1_3_5_n78) );
  XNOR2_X1 pe_1_3_5_U57 ( .A(pe_1_3_5_n73), .B(int_data_res_3__5__0_), .ZN(
        pe_1_3_5_N70) );
  AOI222_X1 pe_1_3_5_U52 ( .A1(int_data_res_4__5__0_), .A2(pe_1_3_5_n64), .B1(
        pe_1_3_5_n1), .B2(pe_1_3_5_n27), .C1(pe_1_3_5_N70), .C2(pe_1_3_5_n28), 
        .ZN(pe_1_3_5_n35) );
  INV_X1 pe_1_3_5_U51 ( .A(pe_1_3_5_n35), .ZN(pe_1_3_5_n84) );
  AOI222_X1 pe_1_3_5_U50 ( .A1(int_data_res_4__5__1_), .A2(pe_1_3_5_n64), .B1(
        pe_1_3_5_N79), .B2(pe_1_3_5_n27), .C1(pe_1_3_5_N71), .C2(pe_1_3_5_n28), 
        .ZN(pe_1_3_5_n34) );
  INV_X1 pe_1_3_5_U49 ( .A(pe_1_3_5_n34), .ZN(pe_1_3_5_n83) );
  AOI222_X1 pe_1_3_5_U48 ( .A1(int_data_res_4__5__3_), .A2(pe_1_3_5_n64), .B1(
        pe_1_3_5_N81), .B2(pe_1_3_5_n27), .C1(pe_1_3_5_N73), .C2(pe_1_3_5_n28), 
        .ZN(pe_1_3_5_n32) );
  INV_X1 pe_1_3_5_U47 ( .A(pe_1_3_5_n32), .ZN(pe_1_3_5_n81) );
  AOI222_X1 pe_1_3_5_U46 ( .A1(int_data_res_4__5__4_), .A2(pe_1_3_5_n64), .B1(
        pe_1_3_5_N82), .B2(pe_1_3_5_n27), .C1(pe_1_3_5_N74), .C2(pe_1_3_5_n28), 
        .ZN(pe_1_3_5_n31) );
  INV_X1 pe_1_3_5_U45 ( .A(pe_1_3_5_n31), .ZN(pe_1_3_5_n80) );
  AOI222_X1 pe_1_3_5_U44 ( .A1(int_data_res_4__5__5_), .A2(pe_1_3_5_n64), .B1(
        pe_1_3_5_N83), .B2(pe_1_3_5_n27), .C1(pe_1_3_5_N75), .C2(pe_1_3_5_n28), 
        .ZN(pe_1_3_5_n30) );
  INV_X1 pe_1_3_5_U43 ( .A(pe_1_3_5_n30), .ZN(pe_1_3_5_n79) );
  NAND2_X1 pe_1_3_5_U42 ( .A1(pe_1_3_5_int_data_0_), .A2(pe_1_3_5_n3), .ZN(
        pe_1_3_5_sub_81_carry[1]) );
  INV_X1 pe_1_3_5_U41 ( .A(pe_1_3_5_int_data_1_), .ZN(pe_1_3_5_n74) );
  INV_X1 pe_1_3_5_U40 ( .A(pe_1_3_5_int_data_2_), .ZN(pe_1_3_5_n75) );
  AND2_X1 pe_1_3_5_U39 ( .A1(pe_1_3_5_int_data_0_), .A2(int_data_res_3__5__0_), 
        .ZN(pe_1_3_5_n2) );
  AOI222_X1 pe_1_3_5_U38 ( .A1(pe_1_3_5_n64), .A2(int_data_res_4__5__7_), .B1(
        pe_1_3_5_N85), .B2(pe_1_3_5_n27), .C1(pe_1_3_5_N77), .C2(pe_1_3_5_n28), 
        .ZN(pe_1_3_5_n26) );
  INV_X1 pe_1_3_5_U37 ( .A(pe_1_3_5_n26), .ZN(pe_1_3_5_n77) );
  NOR3_X1 pe_1_3_5_U36 ( .A1(pe_1_3_5_n59), .A2(pe_1_3_5_n65), .A3(int_ckg[34]), .ZN(pe_1_3_5_n36) );
  OR2_X1 pe_1_3_5_U35 ( .A1(pe_1_3_5_n36), .A2(pe_1_3_5_n64), .ZN(pe_1_3_5_N90) );
  INV_X1 pe_1_3_5_U34 ( .A(n39), .ZN(pe_1_3_5_n63) );
  AND2_X1 pe_1_3_5_U33 ( .A1(int_data_x_3__5__2_), .A2(pe_1_3_5_n58), .ZN(
        pe_1_3_5_int_data_2_) );
  AND2_X1 pe_1_3_5_U32 ( .A1(int_data_x_3__5__1_), .A2(pe_1_3_5_n58), .ZN(
        pe_1_3_5_int_data_1_) );
  AND2_X1 pe_1_3_5_U31 ( .A1(int_data_x_3__5__3_), .A2(pe_1_3_5_n58), .ZN(
        pe_1_3_5_int_data_3_) );
  BUF_X1 pe_1_3_5_U30 ( .A(n61), .Z(pe_1_3_5_n64) );
  INV_X1 pe_1_3_5_U29 ( .A(n33), .ZN(pe_1_3_5_n61) );
  AND2_X1 pe_1_3_5_U28 ( .A1(int_data_x_3__5__0_), .A2(pe_1_3_5_n58), .ZN(
        pe_1_3_5_int_data_0_) );
  NAND2_X1 pe_1_3_5_U27 ( .A1(pe_1_3_5_n44), .A2(pe_1_3_5_n61), .ZN(
        pe_1_3_5_n41) );
  AND3_X1 pe_1_3_5_U26 ( .A1(n75), .A2(pe_1_3_5_n63), .A3(n48), .ZN(
        pe_1_3_5_n44) );
  INV_X1 pe_1_3_5_U25 ( .A(pe_1_3_5_int_data_3_), .ZN(pe_1_3_5_n76) );
  NOR2_X1 pe_1_3_5_U24 ( .A1(pe_1_3_5_n70), .A2(n48), .ZN(pe_1_3_5_n43) );
  NOR2_X1 pe_1_3_5_U23 ( .A1(pe_1_3_5_n57), .A2(pe_1_3_5_n64), .ZN(
        pe_1_3_5_n28) );
  NOR2_X1 pe_1_3_5_U22 ( .A1(n19), .A2(pe_1_3_5_n64), .ZN(pe_1_3_5_n27) );
  INV_X1 pe_1_3_5_U21 ( .A(pe_1_3_5_int_data_0_), .ZN(pe_1_3_5_n73) );
  INV_X1 pe_1_3_5_U20 ( .A(pe_1_3_5_n41), .ZN(pe_1_3_5_n90) );
  INV_X1 pe_1_3_5_U19 ( .A(pe_1_3_5_n37), .ZN(pe_1_3_5_n88) );
  INV_X1 pe_1_3_5_U18 ( .A(pe_1_3_5_n38), .ZN(pe_1_3_5_n87) );
  INV_X1 pe_1_3_5_U17 ( .A(pe_1_3_5_n39), .ZN(pe_1_3_5_n86) );
  NOR2_X1 pe_1_3_5_U16 ( .A1(pe_1_3_5_n68), .A2(pe_1_3_5_n42), .ZN(
        pe_1_3_5_N59) );
  NOR2_X1 pe_1_3_5_U15 ( .A1(pe_1_3_5_n68), .A2(pe_1_3_5_n41), .ZN(
        pe_1_3_5_N60) );
  NOR2_X1 pe_1_3_5_U14 ( .A1(pe_1_3_5_n68), .A2(pe_1_3_5_n38), .ZN(
        pe_1_3_5_N63) );
  NOR2_X1 pe_1_3_5_U13 ( .A1(pe_1_3_5_n67), .A2(pe_1_3_5_n40), .ZN(
        pe_1_3_5_N61) );
  NOR2_X1 pe_1_3_5_U12 ( .A1(pe_1_3_5_n67), .A2(pe_1_3_5_n39), .ZN(
        pe_1_3_5_N62) );
  NOR2_X1 pe_1_3_5_U11 ( .A1(pe_1_3_5_n37), .A2(pe_1_3_5_n67), .ZN(
        pe_1_3_5_N64) );
  NAND2_X1 pe_1_3_5_U10 ( .A1(pe_1_3_5_n44), .A2(pe_1_3_5_n60), .ZN(
        pe_1_3_5_n42) );
  BUF_X1 pe_1_3_5_U9 ( .A(pe_1_3_5_n60), .Z(pe_1_3_5_n55) );
  INV_X1 pe_1_3_5_U8 ( .A(pe_1_3_5_n69), .ZN(pe_1_3_5_n65) );
  BUF_X1 pe_1_3_5_U7 ( .A(pe_1_3_5_n60), .Z(pe_1_3_5_n56) );
  INV_X1 pe_1_3_5_U6 ( .A(pe_1_3_5_n42), .ZN(pe_1_3_5_n89) );
  INV_X1 pe_1_3_5_U5 ( .A(pe_1_3_5_n40), .ZN(pe_1_3_5_n85) );
  INV_X2 pe_1_3_5_U4 ( .A(n83), .ZN(pe_1_3_5_n72) );
  XOR2_X1 pe_1_3_5_U3 ( .A(pe_1_3_5_int_data_0_), .B(int_data_res_3__5__0_), 
        .Z(pe_1_3_5_n1) );
  DFFR_X1 pe_1_3_5_int_q_acc_reg_0_ ( .D(pe_1_3_5_n84), .CK(pe_1_3_5_net5290), 
        .RN(pe_1_3_5_n72), .Q(int_data_res_3__5__0_), .QN(pe_1_3_5_n3) );
  DFFR_X1 pe_1_3_5_int_q_reg_v_reg_0__0_ ( .D(int_data_y_4__5__0_), .CK(
        pe_1_3_5_net5260), .RN(pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_v[20]) );
  DFFR_X1 pe_1_3_5_int_q_reg_v_reg_0__1_ ( .D(int_data_y_4__5__1_), .CK(
        pe_1_3_5_net5260), .RN(pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_v[21]) );
  DFFR_X1 pe_1_3_5_int_q_reg_v_reg_0__2_ ( .D(int_data_y_4__5__2_), .CK(
        pe_1_3_5_net5260), .RN(pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_v[22]) );
  DFFR_X1 pe_1_3_5_int_q_reg_v_reg_0__3_ ( .D(int_data_y_4__5__3_), .CK(
        pe_1_3_5_net5260), .RN(pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_v[23]) );
  DFFR_X1 pe_1_3_5_int_q_reg_v_reg_1__0_ ( .D(int_data_y_4__5__0_), .CK(
        pe_1_3_5_net5265), .RN(pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_v[16]) );
  DFFR_X1 pe_1_3_5_int_q_reg_v_reg_1__1_ ( .D(int_data_y_4__5__1_), .CK(
        pe_1_3_5_net5265), .RN(pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_v[17]) );
  DFFR_X1 pe_1_3_5_int_q_reg_v_reg_1__2_ ( .D(int_data_y_4__5__2_), .CK(
        pe_1_3_5_net5265), .RN(pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_v[18]) );
  DFFR_X1 pe_1_3_5_int_q_reg_v_reg_1__3_ ( .D(int_data_y_4__5__3_), .CK(
        pe_1_3_5_net5265), .RN(pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_v[19]) );
  DFFR_X1 pe_1_3_5_int_q_reg_v_reg_2__0_ ( .D(int_data_y_4__5__0_), .CK(
        pe_1_3_5_net5270), .RN(pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_v[12]) );
  DFFR_X1 pe_1_3_5_int_q_reg_v_reg_2__1_ ( .D(int_data_y_4__5__1_), .CK(
        pe_1_3_5_net5270), .RN(pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_v[13]) );
  DFFR_X1 pe_1_3_5_int_q_reg_v_reg_2__2_ ( .D(int_data_y_4__5__2_), .CK(
        pe_1_3_5_net5270), .RN(pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_v[14]) );
  DFFR_X1 pe_1_3_5_int_q_reg_v_reg_2__3_ ( .D(int_data_y_4__5__3_), .CK(
        pe_1_3_5_net5270), .RN(pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_v[15]) );
  DFFR_X1 pe_1_3_5_int_q_reg_v_reg_3__0_ ( .D(int_data_y_4__5__0_), .CK(
        pe_1_3_5_net5275), .RN(pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_v[8]) );
  DFFR_X1 pe_1_3_5_int_q_reg_v_reg_3__1_ ( .D(int_data_y_4__5__1_), .CK(
        pe_1_3_5_net5275), .RN(pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_v[9]) );
  DFFR_X1 pe_1_3_5_int_q_reg_v_reg_3__2_ ( .D(int_data_y_4__5__2_), .CK(
        pe_1_3_5_net5275), .RN(pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_v[10]) );
  DFFR_X1 pe_1_3_5_int_q_reg_v_reg_3__3_ ( .D(int_data_y_4__5__3_), .CK(
        pe_1_3_5_net5275), .RN(pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_v[11]) );
  DFFR_X1 pe_1_3_5_int_q_reg_v_reg_4__0_ ( .D(int_data_y_4__5__0_), .CK(
        pe_1_3_5_net5280), .RN(pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_v[4]) );
  DFFR_X1 pe_1_3_5_int_q_reg_v_reg_4__1_ ( .D(int_data_y_4__5__1_), .CK(
        pe_1_3_5_net5280), .RN(pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_v[5]) );
  DFFR_X1 pe_1_3_5_int_q_reg_v_reg_4__2_ ( .D(int_data_y_4__5__2_), .CK(
        pe_1_3_5_net5280), .RN(pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_v[6]) );
  DFFR_X1 pe_1_3_5_int_q_reg_v_reg_4__3_ ( .D(int_data_y_4__5__3_), .CK(
        pe_1_3_5_net5280), .RN(pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_v[7]) );
  DFFR_X1 pe_1_3_5_int_q_reg_v_reg_5__0_ ( .D(int_data_y_4__5__0_), .CK(
        pe_1_3_5_net5285), .RN(pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_v[0]) );
  DFFR_X1 pe_1_3_5_int_q_reg_v_reg_5__1_ ( .D(int_data_y_4__5__1_), .CK(
        pe_1_3_5_net5285), .RN(pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_v[1]) );
  DFFR_X1 pe_1_3_5_int_q_reg_v_reg_5__2_ ( .D(int_data_y_4__5__2_), .CK(
        pe_1_3_5_net5285), .RN(pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_v[2]) );
  DFFR_X1 pe_1_3_5_int_q_reg_v_reg_5__3_ ( .D(int_data_y_4__5__3_), .CK(
        pe_1_3_5_net5285), .RN(pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_3_5_int_q_reg_h_reg_0__0_ ( .D(int_data_x_3__6__0_), .SI(
        int_data_y_4__5__0_), .SE(pe_1_3_5_n65), .CK(pe_1_3_5_net5229), .RN(
        pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_3_5_int_q_reg_h_reg_0__1_ ( .D(int_data_x_3__6__1_), .SI(
        int_data_y_4__5__1_), .SE(pe_1_3_5_n65), .CK(pe_1_3_5_net5229), .RN(
        pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_3_5_int_q_reg_h_reg_0__2_ ( .D(int_data_x_3__6__2_), .SI(
        int_data_y_4__5__2_), .SE(pe_1_3_5_n65), .CK(pe_1_3_5_net5229), .RN(
        pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_3_5_int_q_reg_h_reg_0__3_ ( .D(int_data_x_3__6__3_), .SI(
        int_data_y_4__5__3_), .SE(pe_1_3_5_n65), .CK(pe_1_3_5_net5229), .RN(
        pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_3_5_int_q_reg_h_reg_1__0_ ( .D(int_data_x_3__6__0_), .SI(
        int_data_y_4__5__0_), .SE(pe_1_3_5_n65), .CK(pe_1_3_5_net5235), .RN(
        pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_3_5_int_q_reg_h_reg_1__1_ ( .D(int_data_x_3__6__1_), .SI(
        int_data_y_4__5__1_), .SE(pe_1_3_5_n65), .CK(pe_1_3_5_net5235), .RN(
        pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_3_5_int_q_reg_h_reg_1__2_ ( .D(int_data_x_3__6__2_), .SI(
        int_data_y_4__5__2_), .SE(pe_1_3_5_n65), .CK(pe_1_3_5_net5235), .RN(
        pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_3_5_int_q_reg_h_reg_1__3_ ( .D(int_data_x_3__6__3_), .SI(
        int_data_y_4__5__3_), .SE(pe_1_3_5_n65), .CK(pe_1_3_5_net5235), .RN(
        pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_3_5_int_q_reg_h_reg_2__0_ ( .D(int_data_x_3__6__0_), .SI(
        int_data_y_4__5__0_), .SE(pe_1_3_5_n65), .CK(pe_1_3_5_net5240), .RN(
        pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_3_5_int_q_reg_h_reg_2__1_ ( .D(int_data_x_3__6__1_), .SI(
        int_data_y_4__5__1_), .SE(pe_1_3_5_n65), .CK(pe_1_3_5_net5240), .RN(
        pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_3_5_int_q_reg_h_reg_2__2_ ( .D(int_data_x_3__6__2_), .SI(
        int_data_y_4__5__2_), .SE(pe_1_3_5_n65), .CK(pe_1_3_5_net5240), .RN(
        pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_3_5_int_q_reg_h_reg_2__3_ ( .D(int_data_x_3__6__3_), .SI(
        int_data_y_4__5__3_), .SE(pe_1_3_5_n65), .CK(pe_1_3_5_net5240), .RN(
        pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_3_5_int_q_reg_h_reg_3__0_ ( .D(int_data_x_3__6__0_), .SI(
        int_data_y_4__5__0_), .SE(pe_1_3_5_n65), .CK(pe_1_3_5_net5245), .RN(
        pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_3_5_int_q_reg_h_reg_3__1_ ( .D(int_data_x_3__6__1_), .SI(
        int_data_y_4__5__1_), .SE(pe_1_3_5_n65), .CK(pe_1_3_5_net5245), .RN(
        pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_3_5_int_q_reg_h_reg_3__2_ ( .D(int_data_x_3__6__2_), .SI(
        int_data_y_4__5__2_), .SE(pe_1_3_5_n65), .CK(pe_1_3_5_net5245), .RN(
        pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_3_5_int_q_reg_h_reg_3__3_ ( .D(int_data_x_3__6__3_), .SI(
        int_data_y_4__5__3_), .SE(pe_1_3_5_n65), .CK(pe_1_3_5_net5245), .RN(
        pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_3_5_int_q_reg_h_reg_4__0_ ( .D(int_data_x_3__6__0_), .SI(
        int_data_y_4__5__0_), .SE(pe_1_3_5_n66), .CK(pe_1_3_5_net5250), .RN(
        pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_3_5_int_q_reg_h_reg_4__1_ ( .D(int_data_x_3__6__1_), .SI(
        int_data_y_4__5__1_), .SE(pe_1_3_5_n66), .CK(pe_1_3_5_net5250), .RN(
        pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_3_5_int_q_reg_h_reg_4__2_ ( .D(int_data_x_3__6__2_), .SI(
        int_data_y_4__5__2_), .SE(pe_1_3_5_n66), .CK(pe_1_3_5_net5250), .RN(
        pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_3_5_int_q_reg_h_reg_4__3_ ( .D(int_data_x_3__6__3_), .SI(
        int_data_y_4__5__3_), .SE(pe_1_3_5_n66), .CK(pe_1_3_5_net5250), .RN(
        pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_3_5_int_q_reg_h_reg_5__0_ ( .D(int_data_x_3__6__0_), .SI(
        int_data_y_4__5__0_), .SE(pe_1_3_5_n66), .CK(pe_1_3_5_net5255), .RN(
        pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_3_5_int_q_reg_h_reg_5__1_ ( .D(int_data_x_3__6__1_), .SI(
        int_data_y_4__5__1_), .SE(pe_1_3_5_n66), .CK(pe_1_3_5_net5255), .RN(
        pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_3_5_int_q_reg_h_reg_5__2_ ( .D(int_data_x_3__6__2_), .SI(
        int_data_y_4__5__2_), .SE(pe_1_3_5_n66), .CK(pe_1_3_5_net5255), .RN(
        pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_3_5_int_q_reg_h_reg_5__3_ ( .D(int_data_x_3__6__3_), .SI(
        int_data_y_4__5__3_), .SE(pe_1_3_5_n66), .CK(pe_1_3_5_net5255), .RN(
        pe_1_3_5_n72), .Q(pe_1_3_5_int_q_reg_h[3]) );
  FA_X1 pe_1_3_5_sub_81_U2_7 ( .A(int_data_res_3__5__7_), .B(pe_1_3_5_n76), 
        .CI(pe_1_3_5_sub_81_carry[7]), .S(pe_1_3_5_N77) );
  FA_X1 pe_1_3_5_sub_81_U2_6 ( .A(int_data_res_3__5__6_), .B(pe_1_3_5_n76), 
        .CI(pe_1_3_5_sub_81_carry[6]), .CO(pe_1_3_5_sub_81_carry[7]), .S(
        pe_1_3_5_N76) );
  FA_X1 pe_1_3_5_sub_81_U2_5 ( .A(int_data_res_3__5__5_), .B(pe_1_3_5_n76), 
        .CI(pe_1_3_5_sub_81_carry[5]), .CO(pe_1_3_5_sub_81_carry[6]), .S(
        pe_1_3_5_N75) );
  FA_X1 pe_1_3_5_sub_81_U2_4 ( .A(int_data_res_3__5__4_), .B(pe_1_3_5_n76), 
        .CI(pe_1_3_5_sub_81_carry[4]), .CO(pe_1_3_5_sub_81_carry[5]), .S(
        pe_1_3_5_N74) );
  FA_X1 pe_1_3_5_sub_81_U2_3 ( .A(int_data_res_3__5__3_), .B(pe_1_3_5_n76), 
        .CI(pe_1_3_5_sub_81_carry[3]), .CO(pe_1_3_5_sub_81_carry[4]), .S(
        pe_1_3_5_N73) );
  FA_X1 pe_1_3_5_sub_81_U2_2 ( .A(int_data_res_3__5__2_), .B(pe_1_3_5_n75), 
        .CI(pe_1_3_5_sub_81_carry[2]), .CO(pe_1_3_5_sub_81_carry[3]), .S(
        pe_1_3_5_N72) );
  FA_X1 pe_1_3_5_sub_81_U2_1 ( .A(int_data_res_3__5__1_), .B(pe_1_3_5_n74), 
        .CI(pe_1_3_5_sub_81_carry[1]), .CO(pe_1_3_5_sub_81_carry[2]), .S(
        pe_1_3_5_N71) );
  FA_X1 pe_1_3_5_add_83_U1_7 ( .A(int_data_res_3__5__7_), .B(
        pe_1_3_5_int_data_3_), .CI(pe_1_3_5_add_83_carry[7]), .S(pe_1_3_5_N85)
         );
  FA_X1 pe_1_3_5_add_83_U1_6 ( .A(int_data_res_3__5__6_), .B(
        pe_1_3_5_int_data_3_), .CI(pe_1_3_5_add_83_carry[6]), .CO(
        pe_1_3_5_add_83_carry[7]), .S(pe_1_3_5_N84) );
  FA_X1 pe_1_3_5_add_83_U1_5 ( .A(int_data_res_3__5__5_), .B(
        pe_1_3_5_int_data_3_), .CI(pe_1_3_5_add_83_carry[5]), .CO(
        pe_1_3_5_add_83_carry[6]), .S(pe_1_3_5_N83) );
  FA_X1 pe_1_3_5_add_83_U1_4 ( .A(int_data_res_3__5__4_), .B(
        pe_1_3_5_int_data_3_), .CI(pe_1_3_5_add_83_carry[4]), .CO(
        pe_1_3_5_add_83_carry[5]), .S(pe_1_3_5_N82) );
  FA_X1 pe_1_3_5_add_83_U1_3 ( .A(int_data_res_3__5__3_), .B(
        pe_1_3_5_int_data_3_), .CI(pe_1_3_5_add_83_carry[3]), .CO(
        pe_1_3_5_add_83_carry[4]), .S(pe_1_3_5_N81) );
  FA_X1 pe_1_3_5_add_83_U1_2 ( .A(int_data_res_3__5__2_), .B(
        pe_1_3_5_int_data_2_), .CI(pe_1_3_5_add_83_carry[2]), .CO(
        pe_1_3_5_add_83_carry[3]), .S(pe_1_3_5_N80) );
  FA_X1 pe_1_3_5_add_83_U1_1 ( .A(int_data_res_3__5__1_), .B(
        pe_1_3_5_int_data_1_), .CI(pe_1_3_5_n2), .CO(pe_1_3_5_add_83_carry[2]), 
        .S(pe_1_3_5_N79) );
  NAND3_X1 pe_1_3_5_U56 ( .A1(pe_1_3_5_n60), .A2(pe_1_3_5_n43), .A3(
        pe_1_3_5_n62), .ZN(pe_1_3_5_n40) );
  NAND3_X1 pe_1_3_5_U55 ( .A1(pe_1_3_5_n43), .A2(pe_1_3_5_n61), .A3(
        pe_1_3_5_n62), .ZN(pe_1_3_5_n39) );
  NAND3_X1 pe_1_3_5_U54 ( .A1(pe_1_3_5_n43), .A2(pe_1_3_5_n63), .A3(
        pe_1_3_5_n60), .ZN(pe_1_3_5_n38) );
  NAND3_X1 pe_1_3_5_U53 ( .A1(pe_1_3_5_n61), .A2(pe_1_3_5_n63), .A3(
        pe_1_3_5_n43), .ZN(pe_1_3_5_n37) );
  DFFR_X1 pe_1_3_5_int_q_acc_reg_6_ ( .D(pe_1_3_5_n78), .CK(pe_1_3_5_net5290), 
        .RN(pe_1_3_5_n71), .Q(int_data_res_3__5__6_) );
  DFFR_X1 pe_1_3_5_int_q_acc_reg_5_ ( .D(pe_1_3_5_n79), .CK(pe_1_3_5_net5290), 
        .RN(pe_1_3_5_n71), .Q(int_data_res_3__5__5_) );
  DFFR_X1 pe_1_3_5_int_q_acc_reg_4_ ( .D(pe_1_3_5_n80), .CK(pe_1_3_5_net5290), 
        .RN(pe_1_3_5_n71), .Q(int_data_res_3__5__4_) );
  DFFR_X1 pe_1_3_5_int_q_acc_reg_3_ ( .D(pe_1_3_5_n81), .CK(pe_1_3_5_net5290), 
        .RN(pe_1_3_5_n71), .Q(int_data_res_3__5__3_) );
  DFFR_X1 pe_1_3_5_int_q_acc_reg_2_ ( .D(pe_1_3_5_n82), .CK(pe_1_3_5_net5290), 
        .RN(pe_1_3_5_n71), .Q(int_data_res_3__5__2_) );
  DFFR_X1 pe_1_3_5_int_q_acc_reg_1_ ( .D(pe_1_3_5_n83), .CK(pe_1_3_5_net5290), 
        .RN(pe_1_3_5_n71), .Q(int_data_res_3__5__1_) );
  DFFR_X1 pe_1_3_5_int_q_acc_reg_7_ ( .D(pe_1_3_5_n77), .CK(pe_1_3_5_net5290), 
        .RN(pe_1_3_5_n71), .Q(int_data_res_3__5__7_) );
  CLKGATETST_X1 pe_1_3_5_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_3_5_n88), .SE(1'b0), .GCK(pe_1_3_5_net5229) );
  CLKGATETST_X1 pe_1_3_5_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_3_5_n87), .SE(1'b0), .GCK(pe_1_3_5_net5235) );
  CLKGATETST_X1 pe_1_3_5_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_3_5_n86), .SE(1'b0), .GCK(pe_1_3_5_net5240) );
  CLKGATETST_X1 pe_1_3_5_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_3_5_n85), .SE(1'b0), .GCK(pe_1_3_5_net5245) );
  CLKGATETST_X1 pe_1_3_5_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_3_5_n90), .SE(1'b0), .GCK(pe_1_3_5_net5250) );
  CLKGATETST_X1 pe_1_3_5_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_3_5_n89), .SE(1'b0), .GCK(pe_1_3_5_net5255) );
  CLKGATETST_X1 pe_1_3_5_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_3_5_N64), .SE(1'b0), .GCK(pe_1_3_5_net5260) );
  CLKGATETST_X1 pe_1_3_5_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_3_5_N63), .SE(1'b0), .GCK(pe_1_3_5_net5265) );
  CLKGATETST_X1 pe_1_3_5_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_3_5_N62), .SE(1'b0), .GCK(pe_1_3_5_net5270) );
  CLKGATETST_X1 pe_1_3_5_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_3_5_N61), .SE(1'b0), .GCK(pe_1_3_5_net5275) );
  CLKGATETST_X1 pe_1_3_5_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_3_5_N60), .SE(1'b0), .GCK(pe_1_3_5_net5280) );
  CLKGATETST_X1 pe_1_3_5_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_3_5_N59), .SE(1'b0), .GCK(pe_1_3_5_net5285) );
  CLKGATETST_X1 pe_1_3_5_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_3_5_N90), .SE(1'b0), .GCK(pe_1_3_5_net5290) );
  CLKBUF_X1 pe_1_3_6_U112 ( .A(pe_1_3_6_n72), .Z(pe_1_3_6_n71) );
  INV_X1 pe_1_3_6_U111 ( .A(n75), .ZN(pe_1_3_6_n70) );
  INV_X1 pe_1_3_6_U110 ( .A(n67), .ZN(pe_1_3_6_n69) );
  INV_X1 pe_1_3_6_U109 ( .A(n67), .ZN(pe_1_3_6_n68) );
  INV_X1 pe_1_3_6_U108 ( .A(n67), .ZN(pe_1_3_6_n67) );
  INV_X1 pe_1_3_6_U107 ( .A(pe_1_3_6_n69), .ZN(pe_1_3_6_n66) );
  INV_X1 pe_1_3_6_U106 ( .A(pe_1_3_6_n63), .ZN(pe_1_3_6_n62) );
  INV_X1 pe_1_3_6_U105 ( .A(pe_1_3_6_n61), .ZN(pe_1_3_6_n60) );
  INV_X1 pe_1_3_6_U104 ( .A(n27), .ZN(pe_1_3_6_n59) );
  INV_X1 pe_1_3_6_U103 ( .A(pe_1_3_6_n59), .ZN(pe_1_3_6_n58) );
  INV_X1 pe_1_3_6_U102 ( .A(n19), .ZN(pe_1_3_6_n57) );
  MUX2_X1 pe_1_3_6_U101 ( .A(pe_1_3_6_n54), .B(pe_1_3_6_n51), .S(n49), .Z(
        int_data_x_3__6__3_) );
  MUX2_X1 pe_1_3_6_U100 ( .A(pe_1_3_6_n53), .B(pe_1_3_6_n52), .S(pe_1_3_6_n62), 
        .Z(pe_1_3_6_n54) );
  MUX2_X1 pe_1_3_6_U99 ( .A(pe_1_3_6_int_q_reg_h[23]), .B(
        pe_1_3_6_int_q_reg_h[19]), .S(pe_1_3_6_n56), .Z(pe_1_3_6_n53) );
  MUX2_X1 pe_1_3_6_U98 ( .A(pe_1_3_6_int_q_reg_h[15]), .B(
        pe_1_3_6_int_q_reg_h[11]), .S(pe_1_3_6_n56), .Z(pe_1_3_6_n52) );
  MUX2_X1 pe_1_3_6_U97 ( .A(pe_1_3_6_int_q_reg_h[7]), .B(
        pe_1_3_6_int_q_reg_h[3]), .S(pe_1_3_6_n56), .Z(pe_1_3_6_n51) );
  MUX2_X1 pe_1_3_6_U96 ( .A(pe_1_3_6_n50), .B(pe_1_3_6_n47), .S(n49), .Z(
        int_data_x_3__6__2_) );
  MUX2_X1 pe_1_3_6_U95 ( .A(pe_1_3_6_n49), .B(pe_1_3_6_n48), .S(pe_1_3_6_n62), 
        .Z(pe_1_3_6_n50) );
  MUX2_X1 pe_1_3_6_U94 ( .A(pe_1_3_6_int_q_reg_h[22]), .B(
        pe_1_3_6_int_q_reg_h[18]), .S(pe_1_3_6_n56), .Z(pe_1_3_6_n49) );
  MUX2_X1 pe_1_3_6_U93 ( .A(pe_1_3_6_int_q_reg_h[14]), .B(
        pe_1_3_6_int_q_reg_h[10]), .S(pe_1_3_6_n56), .Z(pe_1_3_6_n48) );
  MUX2_X1 pe_1_3_6_U92 ( .A(pe_1_3_6_int_q_reg_h[6]), .B(
        pe_1_3_6_int_q_reg_h[2]), .S(pe_1_3_6_n56), .Z(pe_1_3_6_n47) );
  MUX2_X1 pe_1_3_6_U91 ( .A(pe_1_3_6_n46), .B(pe_1_3_6_n24), .S(n49), .Z(
        int_data_x_3__6__1_) );
  MUX2_X1 pe_1_3_6_U90 ( .A(pe_1_3_6_n45), .B(pe_1_3_6_n25), .S(pe_1_3_6_n62), 
        .Z(pe_1_3_6_n46) );
  MUX2_X1 pe_1_3_6_U89 ( .A(pe_1_3_6_int_q_reg_h[21]), .B(
        pe_1_3_6_int_q_reg_h[17]), .S(pe_1_3_6_n56), .Z(pe_1_3_6_n45) );
  MUX2_X1 pe_1_3_6_U88 ( .A(pe_1_3_6_int_q_reg_h[13]), .B(
        pe_1_3_6_int_q_reg_h[9]), .S(pe_1_3_6_n56), .Z(pe_1_3_6_n25) );
  MUX2_X1 pe_1_3_6_U87 ( .A(pe_1_3_6_int_q_reg_h[5]), .B(
        pe_1_3_6_int_q_reg_h[1]), .S(pe_1_3_6_n56), .Z(pe_1_3_6_n24) );
  MUX2_X1 pe_1_3_6_U86 ( .A(pe_1_3_6_n23), .B(pe_1_3_6_n20), .S(n49), .Z(
        int_data_x_3__6__0_) );
  MUX2_X1 pe_1_3_6_U85 ( .A(pe_1_3_6_n22), .B(pe_1_3_6_n21), .S(pe_1_3_6_n62), 
        .Z(pe_1_3_6_n23) );
  MUX2_X1 pe_1_3_6_U84 ( .A(pe_1_3_6_int_q_reg_h[20]), .B(
        pe_1_3_6_int_q_reg_h[16]), .S(pe_1_3_6_n56), .Z(pe_1_3_6_n22) );
  MUX2_X1 pe_1_3_6_U83 ( .A(pe_1_3_6_int_q_reg_h[12]), .B(
        pe_1_3_6_int_q_reg_h[8]), .S(pe_1_3_6_n56), .Z(pe_1_3_6_n21) );
  MUX2_X1 pe_1_3_6_U82 ( .A(pe_1_3_6_int_q_reg_h[4]), .B(
        pe_1_3_6_int_q_reg_h[0]), .S(pe_1_3_6_n56), .Z(pe_1_3_6_n20) );
  MUX2_X1 pe_1_3_6_U81 ( .A(pe_1_3_6_n19), .B(pe_1_3_6_n16), .S(n49), .Z(
        int_data_y_3__6__3_) );
  MUX2_X1 pe_1_3_6_U80 ( .A(pe_1_3_6_n18), .B(pe_1_3_6_n17), .S(pe_1_3_6_n62), 
        .Z(pe_1_3_6_n19) );
  MUX2_X1 pe_1_3_6_U79 ( .A(pe_1_3_6_int_q_reg_v[23]), .B(
        pe_1_3_6_int_q_reg_v[19]), .S(pe_1_3_6_n55), .Z(pe_1_3_6_n18) );
  MUX2_X1 pe_1_3_6_U78 ( .A(pe_1_3_6_int_q_reg_v[15]), .B(
        pe_1_3_6_int_q_reg_v[11]), .S(pe_1_3_6_n55), .Z(pe_1_3_6_n17) );
  MUX2_X1 pe_1_3_6_U77 ( .A(pe_1_3_6_int_q_reg_v[7]), .B(
        pe_1_3_6_int_q_reg_v[3]), .S(pe_1_3_6_n55), .Z(pe_1_3_6_n16) );
  MUX2_X1 pe_1_3_6_U76 ( .A(pe_1_3_6_n15), .B(pe_1_3_6_n12), .S(n49), .Z(
        int_data_y_3__6__2_) );
  MUX2_X1 pe_1_3_6_U75 ( .A(pe_1_3_6_n14), .B(pe_1_3_6_n13), .S(pe_1_3_6_n62), 
        .Z(pe_1_3_6_n15) );
  MUX2_X1 pe_1_3_6_U74 ( .A(pe_1_3_6_int_q_reg_v[22]), .B(
        pe_1_3_6_int_q_reg_v[18]), .S(pe_1_3_6_n55), .Z(pe_1_3_6_n14) );
  MUX2_X1 pe_1_3_6_U73 ( .A(pe_1_3_6_int_q_reg_v[14]), .B(
        pe_1_3_6_int_q_reg_v[10]), .S(pe_1_3_6_n55), .Z(pe_1_3_6_n13) );
  MUX2_X1 pe_1_3_6_U72 ( .A(pe_1_3_6_int_q_reg_v[6]), .B(
        pe_1_3_6_int_q_reg_v[2]), .S(pe_1_3_6_n55), .Z(pe_1_3_6_n12) );
  MUX2_X1 pe_1_3_6_U71 ( .A(pe_1_3_6_n11), .B(pe_1_3_6_n8), .S(n49), .Z(
        int_data_y_3__6__1_) );
  MUX2_X1 pe_1_3_6_U70 ( .A(pe_1_3_6_n10), .B(pe_1_3_6_n9), .S(pe_1_3_6_n62), 
        .Z(pe_1_3_6_n11) );
  MUX2_X1 pe_1_3_6_U69 ( .A(pe_1_3_6_int_q_reg_v[21]), .B(
        pe_1_3_6_int_q_reg_v[17]), .S(pe_1_3_6_n55), .Z(pe_1_3_6_n10) );
  MUX2_X1 pe_1_3_6_U68 ( .A(pe_1_3_6_int_q_reg_v[13]), .B(
        pe_1_3_6_int_q_reg_v[9]), .S(pe_1_3_6_n55), .Z(pe_1_3_6_n9) );
  MUX2_X1 pe_1_3_6_U67 ( .A(pe_1_3_6_int_q_reg_v[5]), .B(
        pe_1_3_6_int_q_reg_v[1]), .S(pe_1_3_6_n55), .Z(pe_1_3_6_n8) );
  MUX2_X1 pe_1_3_6_U66 ( .A(pe_1_3_6_n7), .B(pe_1_3_6_n4), .S(n49), .Z(
        int_data_y_3__6__0_) );
  MUX2_X1 pe_1_3_6_U65 ( .A(pe_1_3_6_n6), .B(pe_1_3_6_n5), .S(pe_1_3_6_n62), 
        .Z(pe_1_3_6_n7) );
  MUX2_X1 pe_1_3_6_U64 ( .A(pe_1_3_6_int_q_reg_v[20]), .B(
        pe_1_3_6_int_q_reg_v[16]), .S(pe_1_3_6_n55), .Z(pe_1_3_6_n6) );
  MUX2_X1 pe_1_3_6_U63 ( .A(pe_1_3_6_int_q_reg_v[12]), .B(
        pe_1_3_6_int_q_reg_v[8]), .S(pe_1_3_6_n55), .Z(pe_1_3_6_n5) );
  MUX2_X1 pe_1_3_6_U62 ( .A(pe_1_3_6_int_q_reg_v[4]), .B(
        pe_1_3_6_int_q_reg_v[0]), .S(pe_1_3_6_n55), .Z(pe_1_3_6_n4) );
  AOI222_X1 pe_1_3_6_U61 ( .A1(int_data_res_4__6__2_), .A2(pe_1_3_6_n64), .B1(
        pe_1_3_6_N80), .B2(pe_1_3_6_n27), .C1(pe_1_3_6_N72), .C2(pe_1_3_6_n28), 
        .ZN(pe_1_3_6_n33) );
  INV_X1 pe_1_3_6_U60 ( .A(pe_1_3_6_n33), .ZN(pe_1_3_6_n82) );
  AOI222_X1 pe_1_3_6_U59 ( .A1(int_data_res_4__6__6_), .A2(pe_1_3_6_n64), .B1(
        pe_1_3_6_N84), .B2(pe_1_3_6_n27), .C1(pe_1_3_6_N76), .C2(pe_1_3_6_n28), 
        .ZN(pe_1_3_6_n29) );
  INV_X1 pe_1_3_6_U58 ( .A(pe_1_3_6_n29), .ZN(pe_1_3_6_n78) );
  XNOR2_X1 pe_1_3_6_U57 ( .A(pe_1_3_6_n73), .B(int_data_res_3__6__0_), .ZN(
        pe_1_3_6_N70) );
  AOI222_X1 pe_1_3_6_U52 ( .A1(int_data_res_4__6__0_), .A2(pe_1_3_6_n64), .B1(
        pe_1_3_6_n1), .B2(pe_1_3_6_n27), .C1(pe_1_3_6_N70), .C2(pe_1_3_6_n28), 
        .ZN(pe_1_3_6_n35) );
  INV_X1 pe_1_3_6_U51 ( .A(pe_1_3_6_n35), .ZN(pe_1_3_6_n84) );
  AOI222_X1 pe_1_3_6_U50 ( .A1(int_data_res_4__6__1_), .A2(pe_1_3_6_n64), .B1(
        pe_1_3_6_N79), .B2(pe_1_3_6_n27), .C1(pe_1_3_6_N71), .C2(pe_1_3_6_n28), 
        .ZN(pe_1_3_6_n34) );
  INV_X1 pe_1_3_6_U49 ( .A(pe_1_3_6_n34), .ZN(pe_1_3_6_n83) );
  AOI222_X1 pe_1_3_6_U48 ( .A1(int_data_res_4__6__3_), .A2(pe_1_3_6_n64), .B1(
        pe_1_3_6_N81), .B2(pe_1_3_6_n27), .C1(pe_1_3_6_N73), .C2(pe_1_3_6_n28), 
        .ZN(pe_1_3_6_n32) );
  INV_X1 pe_1_3_6_U47 ( .A(pe_1_3_6_n32), .ZN(pe_1_3_6_n81) );
  AOI222_X1 pe_1_3_6_U46 ( .A1(int_data_res_4__6__4_), .A2(pe_1_3_6_n64), .B1(
        pe_1_3_6_N82), .B2(pe_1_3_6_n27), .C1(pe_1_3_6_N74), .C2(pe_1_3_6_n28), 
        .ZN(pe_1_3_6_n31) );
  INV_X1 pe_1_3_6_U45 ( .A(pe_1_3_6_n31), .ZN(pe_1_3_6_n80) );
  AOI222_X1 pe_1_3_6_U44 ( .A1(int_data_res_4__6__5_), .A2(pe_1_3_6_n64), .B1(
        pe_1_3_6_N83), .B2(pe_1_3_6_n27), .C1(pe_1_3_6_N75), .C2(pe_1_3_6_n28), 
        .ZN(pe_1_3_6_n30) );
  INV_X1 pe_1_3_6_U43 ( .A(pe_1_3_6_n30), .ZN(pe_1_3_6_n79) );
  NAND2_X1 pe_1_3_6_U42 ( .A1(pe_1_3_6_int_data_0_), .A2(pe_1_3_6_n3), .ZN(
        pe_1_3_6_sub_81_carry[1]) );
  INV_X1 pe_1_3_6_U41 ( .A(pe_1_3_6_int_data_1_), .ZN(pe_1_3_6_n74) );
  INV_X1 pe_1_3_6_U40 ( .A(pe_1_3_6_int_data_2_), .ZN(pe_1_3_6_n75) );
  AND2_X1 pe_1_3_6_U39 ( .A1(pe_1_3_6_int_data_0_), .A2(int_data_res_3__6__0_), 
        .ZN(pe_1_3_6_n2) );
  AOI222_X1 pe_1_3_6_U38 ( .A1(pe_1_3_6_n64), .A2(int_data_res_4__6__7_), .B1(
        pe_1_3_6_N85), .B2(pe_1_3_6_n27), .C1(pe_1_3_6_N77), .C2(pe_1_3_6_n28), 
        .ZN(pe_1_3_6_n26) );
  INV_X1 pe_1_3_6_U37 ( .A(pe_1_3_6_n26), .ZN(pe_1_3_6_n77) );
  NOR3_X1 pe_1_3_6_U36 ( .A1(pe_1_3_6_n59), .A2(pe_1_3_6_n65), .A3(int_ckg[33]), .ZN(pe_1_3_6_n36) );
  OR2_X1 pe_1_3_6_U35 ( .A1(pe_1_3_6_n36), .A2(pe_1_3_6_n64), .ZN(pe_1_3_6_N90) );
  INV_X1 pe_1_3_6_U34 ( .A(n39), .ZN(pe_1_3_6_n63) );
  AND2_X1 pe_1_3_6_U33 ( .A1(int_data_x_3__6__2_), .A2(pe_1_3_6_n58), .ZN(
        pe_1_3_6_int_data_2_) );
  AND2_X1 pe_1_3_6_U32 ( .A1(int_data_x_3__6__1_), .A2(pe_1_3_6_n58), .ZN(
        pe_1_3_6_int_data_1_) );
  AND2_X1 pe_1_3_6_U31 ( .A1(int_data_x_3__6__3_), .A2(pe_1_3_6_n58), .ZN(
        pe_1_3_6_int_data_3_) );
  BUF_X1 pe_1_3_6_U30 ( .A(n61), .Z(pe_1_3_6_n64) );
  INV_X1 pe_1_3_6_U29 ( .A(n33), .ZN(pe_1_3_6_n61) );
  AND2_X1 pe_1_3_6_U28 ( .A1(int_data_x_3__6__0_), .A2(pe_1_3_6_n58), .ZN(
        pe_1_3_6_int_data_0_) );
  NAND2_X1 pe_1_3_6_U27 ( .A1(pe_1_3_6_n44), .A2(pe_1_3_6_n61), .ZN(
        pe_1_3_6_n41) );
  AND3_X1 pe_1_3_6_U26 ( .A1(n75), .A2(pe_1_3_6_n63), .A3(n49), .ZN(
        pe_1_3_6_n44) );
  INV_X1 pe_1_3_6_U25 ( .A(pe_1_3_6_int_data_3_), .ZN(pe_1_3_6_n76) );
  NOR2_X1 pe_1_3_6_U24 ( .A1(pe_1_3_6_n70), .A2(n49), .ZN(pe_1_3_6_n43) );
  NOR2_X1 pe_1_3_6_U23 ( .A1(pe_1_3_6_n57), .A2(pe_1_3_6_n64), .ZN(
        pe_1_3_6_n28) );
  NOR2_X1 pe_1_3_6_U22 ( .A1(n19), .A2(pe_1_3_6_n64), .ZN(pe_1_3_6_n27) );
  INV_X1 pe_1_3_6_U21 ( .A(pe_1_3_6_int_data_0_), .ZN(pe_1_3_6_n73) );
  INV_X1 pe_1_3_6_U20 ( .A(pe_1_3_6_n41), .ZN(pe_1_3_6_n90) );
  INV_X1 pe_1_3_6_U19 ( .A(pe_1_3_6_n37), .ZN(pe_1_3_6_n88) );
  INV_X1 pe_1_3_6_U18 ( .A(pe_1_3_6_n38), .ZN(pe_1_3_6_n87) );
  INV_X1 pe_1_3_6_U17 ( .A(pe_1_3_6_n39), .ZN(pe_1_3_6_n86) );
  NOR2_X1 pe_1_3_6_U16 ( .A1(pe_1_3_6_n68), .A2(pe_1_3_6_n42), .ZN(
        pe_1_3_6_N59) );
  NOR2_X1 pe_1_3_6_U15 ( .A1(pe_1_3_6_n68), .A2(pe_1_3_6_n41), .ZN(
        pe_1_3_6_N60) );
  NOR2_X1 pe_1_3_6_U14 ( .A1(pe_1_3_6_n68), .A2(pe_1_3_6_n38), .ZN(
        pe_1_3_6_N63) );
  NOR2_X1 pe_1_3_6_U13 ( .A1(pe_1_3_6_n67), .A2(pe_1_3_6_n40), .ZN(
        pe_1_3_6_N61) );
  NOR2_X1 pe_1_3_6_U12 ( .A1(pe_1_3_6_n67), .A2(pe_1_3_6_n39), .ZN(
        pe_1_3_6_N62) );
  NOR2_X1 pe_1_3_6_U11 ( .A1(pe_1_3_6_n37), .A2(pe_1_3_6_n67), .ZN(
        pe_1_3_6_N64) );
  NAND2_X1 pe_1_3_6_U10 ( .A1(pe_1_3_6_n44), .A2(pe_1_3_6_n60), .ZN(
        pe_1_3_6_n42) );
  BUF_X1 pe_1_3_6_U9 ( .A(pe_1_3_6_n60), .Z(pe_1_3_6_n55) );
  INV_X1 pe_1_3_6_U8 ( .A(pe_1_3_6_n69), .ZN(pe_1_3_6_n65) );
  BUF_X1 pe_1_3_6_U7 ( .A(pe_1_3_6_n60), .Z(pe_1_3_6_n56) );
  INV_X1 pe_1_3_6_U6 ( .A(pe_1_3_6_n42), .ZN(pe_1_3_6_n89) );
  INV_X1 pe_1_3_6_U5 ( .A(pe_1_3_6_n40), .ZN(pe_1_3_6_n85) );
  INV_X2 pe_1_3_6_U4 ( .A(n83), .ZN(pe_1_3_6_n72) );
  XOR2_X1 pe_1_3_6_U3 ( .A(pe_1_3_6_int_data_0_), .B(int_data_res_3__6__0_), 
        .Z(pe_1_3_6_n1) );
  DFFR_X1 pe_1_3_6_int_q_acc_reg_0_ ( .D(pe_1_3_6_n84), .CK(pe_1_3_6_net5212), 
        .RN(pe_1_3_6_n72), .Q(int_data_res_3__6__0_), .QN(pe_1_3_6_n3) );
  DFFR_X1 pe_1_3_6_int_q_reg_v_reg_0__0_ ( .D(int_data_y_4__6__0_), .CK(
        pe_1_3_6_net5182), .RN(pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_v[20]) );
  DFFR_X1 pe_1_3_6_int_q_reg_v_reg_0__1_ ( .D(int_data_y_4__6__1_), .CK(
        pe_1_3_6_net5182), .RN(pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_v[21]) );
  DFFR_X1 pe_1_3_6_int_q_reg_v_reg_0__2_ ( .D(int_data_y_4__6__2_), .CK(
        pe_1_3_6_net5182), .RN(pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_v[22]) );
  DFFR_X1 pe_1_3_6_int_q_reg_v_reg_0__3_ ( .D(int_data_y_4__6__3_), .CK(
        pe_1_3_6_net5182), .RN(pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_v[23]) );
  DFFR_X1 pe_1_3_6_int_q_reg_v_reg_1__0_ ( .D(int_data_y_4__6__0_), .CK(
        pe_1_3_6_net5187), .RN(pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_v[16]) );
  DFFR_X1 pe_1_3_6_int_q_reg_v_reg_1__1_ ( .D(int_data_y_4__6__1_), .CK(
        pe_1_3_6_net5187), .RN(pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_v[17]) );
  DFFR_X1 pe_1_3_6_int_q_reg_v_reg_1__2_ ( .D(int_data_y_4__6__2_), .CK(
        pe_1_3_6_net5187), .RN(pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_v[18]) );
  DFFR_X1 pe_1_3_6_int_q_reg_v_reg_1__3_ ( .D(int_data_y_4__6__3_), .CK(
        pe_1_3_6_net5187), .RN(pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_v[19]) );
  DFFR_X1 pe_1_3_6_int_q_reg_v_reg_2__0_ ( .D(int_data_y_4__6__0_), .CK(
        pe_1_3_6_net5192), .RN(pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_v[12]) );
  DFFR_X1 pe_1_3_6_int_q_reg_v_reg_2__1_ ( .D(int_data_y_4__6__1_), .CK(
        pe_1_3_6_net5192), .RN(pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_v[13]) );
  DFFR_X1 pe_1_3_6_int_q_reg_v_reg_2__2_ ( .D(int_data_y_4__6__2_), .CK(
        pe_1_3_6_net5192), .RN(pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_v[14]) );
  DFFR_X1 pe_1_3_6_int_q_reg_v_reg_2__3_ ( .D(int_data_y_4__6__3_), .CK(
        pe_1_3_6_net5192), .RN(pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_v[15]) );
  DFFR_X1 pe_1_3_6_int_q_reg_v_reg_3__0_ ( .D(int_data_y_4__6__0_), .CK(
        pe_1_3_6_net5197), .RN(pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_v[8]) );
  DFFR_X1 pe_1_3_6_int_q_reg_v_reg_3__1_ ( .D(int_data_y_4__6__1_), .CK(
        pe_1_3_6_net5197), .RN(pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_v[9]) );
  DFFR_X1 pe_1_3_6_int_q_reg_v_reg_3__2_ ( .D(int_data_y_4__6__2_), .CK(
        pe_1_3_6_net5197), .RN(pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_v[10]) );
  DFFR_X1 pe_1_3_6_int_q_reg_v_reg_3__3_ ( .D(int_data_y_4__6__3_), .CK(
        pe_1_3_6_net5197), .RN(pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_v[11]) );
  DFFR_X1 pe_1_3_6_int_q_reg_v_reg_4__0_ ( .D(int_data_y_4__6__0_), .CK(
        pe_1_3_6_net5202), .RN(pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_v[4]) );
  DFFR_X1 pe_1_3_6_int_q_reg_v_reg_4__1_ ( .D(int_data_y_4__6__1_), .CK(
        pe_1_3_6_net5202), .RN(pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_v[5]) );
  DFFR_X1 pe_1_3_6_int_q_reg_v_reg_4__2_ ( .D(int_data_y_4__6__2_), .CK(
        pe_1_3_6_net5202), .RN(pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_v[6]) );
  DFFR_X1 pe_1_3_6_int_q_reg_v_reg_4__3_ ( .D(int_data_y_4__6__3_), .CK(
        pe_1_3_6_net5202), .RN(pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_v[7]) );
  DFFR_X1 pe_1_3_6_int_q_reg_v_reg_5__0_ ( .D(int_data_y_4__6__0_), .CK(
        pe_1_3_6_net5207), .RN(pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_v[0]) );
  DFFR_X1 pe_1_3_6_int_q_reg_v_reg_5__1_ ( .D(int_data_y_4__6__1_), .CK(
        pe_1_3_6_net5207), .RN(pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_v[1]) );
  DFFR_X1 pe_1_3_6_int_q_reg_v_reg_5__2_ ( .D(int_data_y_4__6__2_), .CK(
        pe_1_3_6_net5207), .RN(pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_v[2]) );
  DFFR_X1 pe_1_3_6_int_q_reg_v_reg_5__3_ ( .D(int_data_y_4__6__3_), .CK(
        pe_1_3_6_net5207), .RN(pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_3_6_int_q_reg_h_reg_0__0_ ( .D(int_data_x_3__7__0_), .SI(
        int_data_y_4__6__0_), .SE(pe_1_3_6_n65), .CK(pe_1_3_6_net5151), .RN(
        pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_3_6_int_q_reg_h_reg_0__1_ ( .D(int_data_x_3__7__1_), .SI(
        int_data_y_4__6__1_), .SE(pe_1_3_6_n65), .CK(pe_1_3_6_net5151), .RN(
        pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_3_6_int_q_reg_h_reg_0__2_ ( .D(int_data_x_3__7__2_), .SI(
        int_data_y_4__6__2_), .SE(pe_1_3_6_n65), .CK(pe_1_3_6_net5151), .RN(
        pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_3_6_int_q_reg_h_reg_0__3_ ( .D(int_data_x_3__7__3_), .SI(
        int_data_y_4__6__3_), .SE(pe_1_3_6_n65), .CK(pe_1_3_6_net5151), .RN(
        pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_3_6_int_q_reg_h_reg_1__0_ ( .D(int_data_x_3__7__0_), .SI(
        int_data_y_4__6__0_), .SE(pe_1_3_6_n65), .CK(pe_1_3_6_net5157), .RN(
        pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_3_6_int_q_reg_h_reg_1__1_ ( .D(int_data_x_3__7__1_), .SI(
        int_data_y_4__6__1_), .SE(pe_1_3_6_n65), .CK(pe_1_3_6_net5157), .RN(
        pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_3_6_int_q_reg_h_reg_1__2_ ( .D(int_data_x_3__7__2_), .SI(
        int_data_y_4__6__2_), .SE(pe_1_3_6_n65), .CK(pe_1_3_6_net5157), .RN(
        pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_3_6_int_q_reg_h_reg_1__3_ ( .D(int_data_x_3__7__3_), .SI(
        int_data_y_4__6__3_), .SE(pe_1_3_6_n65), .CK(pe_1_3_6_net5157), .RN(
        pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_3_6_int_q_reg_h_reg_2__0_ ( .D(int_data_x_3__7__0_), .SI(
        int_data_y_4__6__0_), .SE(pe_1_3_6_n65), .CK(pe_1_3_6_net5162), .RN(
        pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_3_6_int_q_reg_h_reg_2__1_ ( .D(int_data_x_3__7__1_), .SI(
        int_data_y_4__6__1_), .SE(pe_1_3_6_n65), .CK(pe_1_3_6_net5162), .RN(
        pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_3_6_int_q_reg_h_reg_2__2_ ( .D(int_data_x_3__7__2_), .SI(
        int_data_y_4__6__2_), .SE(pe_1_3_6_n65), .CK(pe_1_3_6_net5162), .RN(
        pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_3_6_int_q_reg_h_reg_2__3_ ( .D(int_data_x_3__7__3_), .SI(
        int_data_y_4__6__3_), .SE(pe_1_3_6_n65), .CK(pe_1_3_6_net5162), .RN(
        pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_3_6_int_q_reg_h_reg_3__0_ ( .D(int_data_x_3__7__0_), .SI(
        int_data_y_4__6__0_), .SE(pe_1_3_6_n65), .CK(pe_1_3_6_net5167), .RN(
        pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_3_6_int_q_reg_h_reg_3__1_ ( .D(int_data_x_3__7__1_), .SI(
        int_data_y_4__6__1_), .SE(pe_1_3_6_n65), .CK(pe_1_3_6_net5167), .RN(
        pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_3_6_int_q_reg_h_reg_3__2_ ( .D(int_data_x_3__7__2_), .SI(
        int_data_y_4__6__2_), .SE(pe_1_3_6_n65), .CK(pe_1_3_6_net5167), .RN(
        pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_3_6_int_q_reg_h_reg_3__3_ ( .D(int_data_x_3__7__3_), .SI(
        int_data_y_4__6__3_), .SE(pe_1_3_6_n65), .CK(pe_1_3_6_net5167), .RN(
        pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_3_6_int_q_reg_h_reg_4__0_ ( .D(int_data_x_3__7__0_), .SI(
        int_data_y_4__6__0_), .SE(pe_1_3_6_n66), .CK(pe_1_3_6_net5172), .RN(
        pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_3_6_int_q_reg_h_reg_4__1_ ( .D(int_data_x_3__7__1_), .SI(
        int_data_y_4__6__1_), .SE(pe_1_3_6_n66), .CK(pe_1_3_6_net5172), .RN(
        pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_3_6_int_q_reg_h_reg_4__2_ ( .D(int_data_x_3__7__2_), .SI(
        int_data_y_4__6__2_), .SE(pe_1_3_6_n66), .CK(pe_1_3_6_net5172), .RN(
        pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_3_6_int_q_reg_h_reg_4__3_ ( .D(int_data_x_3__7__3_), .SI(
        int_data_y_4__6__3_), .SE(pe_1_3_6_n66), .CK(pe_1_3_6_net5172), .RN(
        pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_3_6_int_q_reg_h_reg_5__0_ ( .D(int_data_x_3__7__0_), .SI(
        int_data_y_4__6__0_), .SE(pe_1_3_6_n66), .CK(pe_1_3_6_net5177), .RN(
        pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_3_6_int_q_reg_h_reg_5__1_ ( .D(int_data_x_3__7__1_), .SI(
        int_data_y_4__6__1_), .SE(pe_1_3_6_n66), .CK(pe_1_3_6_net5177), .RN(
        pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_3_6_int_q_reg_h_reg_5__2_ ( .D(int_data_x_3__7__2_), .SI(
        int_data_y_4__6__2_), .SE(pe_1_3_6_n66), .CK(pe_1_3_6_net5177), .RN(
        pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_3_6_int_q_reg_h_reg_5__3_ ( .D(int_data_x_3__7__3_), .SI(
        int_data_y_4__6__3_), .SE(pe_1_3_6_n66), .CK(pe_1_3_6_net5177), .RN(
        pe_1_3_6_n72), .Q(pe_1_3_6_int_q_reg_h[3]) );
  FA_X1 pe_1_3_6_sub_81_U2_7 ( .A(int_data_res_3__6__7_), .B(pe_1_3_6_n76), 
        .CI(pe_1_3_6_sub_81_carry[7]), .S(pe_1_3_6_N77) );
  FA_X1 pe_1_3_6_sub_81_U2_6 ( .A(int_data_res_3__6__6_), .B(pe_1_3_6_n76), 
        .CI(pe_1_3_6_sub_81_carry[6]), .CO(pe_1_3_6_sub_81_carry[7]), .S(
        pe_1_3_6_N76) );
  FA_X1 pe_1_3_6_sub_81_U2_5 ( .A(int_data_res_3__6__5_), .B(pe_1_3_6_n76), 
        .CI(pe_1_3_6_sub_81_carry[5]), .CO(pe_1_3_6_sub_81_carry[6]), .S(
        pe_1_3_6_N75) );
  FA_X1 pe_1_3_6_sub_81_U2_4 ( .A(int_data_res_3__6__4_), .B(pe_1_3_6_n76), 
        .CI(pe_1_3_6_sub_81_carry[4]), .CO(pe_1_3_6_sub_81_carry[5]), .S(
        pe_1_3_6_N74) );
  FA_X1 pe_1_3_6_sub_81_U2_3 ( .A(int_data_res_3__6__3_), .B(pe_1_3_6_n76), 
        .CI(pe_1_3_6_sub_81_carry[3]), .CO(pe_1_3_6_sub_81_carry[4]), .S(
        pe_1_3_6_N73) );
  FA_X1 pe_1_3_6_sub_81_U2_2 ( .A(int_data_res_3__6__2_), .B(pe_1_3_6_n75), 
        .CI(pe_1_3_6_sub_81_carry[2]), .CO(pe_1_3_6_sub_81_carry[3]), .S(
        pe_1_3_6_N72) );
  FA_X1 pe_1_3_6_sub_81_U2_1 ( .A(int_data_res_3__6__1_), .B(pe_1_3_6_n74), 
        .CI(pe_1_3_6_sub_81_carry[1]), .CO(pe_1_3_6_sub_81_carry[2]), .S(
        pe_1_3_6_N71) );
  FA_X1 pe_1_3_6_add_83_U1_7 ( .A(int_data_res_3__6__7_), .B(
        pe_1_3_6_int_data_3_), .CI(pe_1_3_6_add_83_carry[7]), .S(pe_1_3_6_N85)
         );
  FA_X1 pe_1_3_6_add_83_U1_6 ( .A(int_data_res_3__6__6_), .B(
        pe_1_3_6_int_data_3_), .CI(pe_1_3_6_add_83_carry[6]), .CO(
        pe_1_3_6_add_83_carry[7]), .S(pe_1_3_6_N84) );
  FA_X1 pe_1_3_6_add_83_U1_5 ( .A(int_data_res_3__6__5_), .B(
        pe_1_3_6_int_data_3_), .CI(pe_1_3_6_add_83_carry[5]), .CO(
        pe_1_3_6_add_83_carry[6]), .S(pe_1_3_6_N83) );
  FA_X1 pe_1_3_6_add_83_U1_4 ( .A(int_data_res_3__6__4_), .B(
        pe_1_3_6_int_data_3_), .CI(pe_1_3_6_add_83_carry[4]), .CO(
        pe_1_3_6_add_83_carry[5]), .S(pe_1_3_6_N82) );
  FA_X1 pe_1_3_6_add_83_U1_3 ( .A(int_data_res_3__6__3_), .B(
        pe_1_3_6_int_data_3_), .CI(pe_1_3_6_add_83_carry[3]), .CO(
        pe_1_3_6_add_83_carry[4]), .S(pe_1_3_6_N81) );
  FA_X1 pe_1_3_6_add_83_U1_2 ( .A(int_data_res_3__6__2_), .B(
        pe_1_3_6_int_data_2_), .CI(pe_1_3_6_add_83_carry[2]), .CO(
        pe_1_3_6_add_83_carry[3]), .S(pe_1_3_6_N80) );
  FA_X1 pe_1_3_6_add_83_U1_1 ( .A(int_data_res_3__6__1_), .B(
        pe_1_3_6_int_data_1_), .CI(pe_1_3_6_n2), .CO(pe_1_3_6_add_83_carry[2]), 
        .S(pe_1_3_6_N79) );
  NAND3_X1 pe_1_3_6_U56 ( .A1(pe_1_3_6_n60), .A2(pe_1_3_6_n43), .A3(
        pe_1_3_6_n62), .ZN(pe_1_3_6_n40) );
  NAND3_X1 pe_1_3_6_U55 ( .A1(pe_1_3_6_n43), .A2(pe_1_3_6_n61), .A3(
        pe_1_3_6_n62), .ZN(pe_1_3_6_n39) );
  NAND3_X1 pe_1_3_6_U54 ( .A1(pe_1_3_6_n43), .A2(pe_1_3_6_n63), .A3(
        pe_1_3_6_n60), .ZN(pe_1_3_6_n38) );
  NAND3_X1 pe_1_3_6_U53 ( .A1(pe_1_3_6_n61), .A2(pe_1_3_6_n63), .A3(
        pe_1_3_6_n43), .ZN(pe_1_3_6_n37) );
  DFFR_X1 pe_1_3_6_int_q_acc_reg_6_ ( .D(pe_1_3_6_n78), .CK(pe_1_3_6_net5212), 
        .RN(pe_1_3_6_n71), .Q(int_data_res_3__6__6_) );
  DFFR_X1 pe_1_3_6_int_q_acc_reg_5_ ( .D(pe_1_3_6_n79), .CK(pe_1_3_6_net5212), 
        .RN(pe_1_3_6_n71), .Q(int_data_res_3__6__5_) );
  DFFR_X1 pe_1_3_6_int_q_acc_reg_4_ ( .D(pe_1_3_6_n80), .CK(pe_1_3_6_net5212), 
        .RN(pe_1_3_6_n71), .Q(int_data_res_3__6__4_) );
  DFFR_X1 pe_1_3_6_int_q_acc_reg_3_ ( .D(pe_1_3_6_n81), .CK(pe_1_3_6_net5212), 
        .RN(pe_1_3_6_n71), .Q(int_data_res_3__6__3_) );
  DFFR_X1 pe_1_3_6_int_q_acc_reg_2_ ( .D(pe_1_3_6_n82), .CK(pe_1_3_6_net5212), 
        .RN(pe_1_3_6_n71), .Q(int_data_res_3__6__2_) );
  DFFR_X1 pe_1_3_6_int_q_acc_reg_1_ ( .D(pe_1_3_6_n83), .CK(pe_1_3_6_net5212), 
        .RN(pe_1_3_6_n71), .Q(int_data_res_3__6__1_) );
  DFFR_X1 pe_1_3_6_int_q_acc_reg_7_ ( .D(pe_1_3_6_n77), .CK(pe_1_3_6_net5212), 
        .RN(pe_1_3_6_n71), .Q(int_data_res_3__6__7_) );
  CLKGATETST_X1 pe_1_3_6_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_3_6_n88), .SE(1'b0), .GCK(pe_1_3_6_net5151) );
  CLKGATETST_X1 pe_1_3_6_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_3_6_n87), .SE(1'b0), .GCK(pe_1_3_6_net5157) );
  CLKGATETST_X1 pe_1_3_6_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_3_6_n86), .SE(1'b0), .GCK(pe_1_3_6_net5162) );
  CLKGATETST_X1 pe_1_3_6_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_3_6_n85), .SE(1'b0), .GCK(pe_1_3_6_net5167) );
  CLKGATETST_X1 pe_1_3_6_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_3_6_n90), .SE(1'b0), .GCK(pe_1_3_6_net5172) );
  CLKGATETST_X1 pe_1_3_6_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_3_6_n89), .SE(1'b0), .GCK(pe_1_3_6_net5177) );
  CLKGATETST_X1 pe_1_3_6_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_3_6_N64), .SE(1'b0), .GCK(pe_1_3_6_net5182) );
  CLKGATETST_X1 pe_1_3_6_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_3_6_N63), .SE(1'b0), .GCK(pe_1_3_6_net5187) );
  CLKGATETST_X1 pe_1_3_6_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_3_6_N62), .SE(1'b0), .GCK(pe_1_3_6_net5192) );
  CLKGATETST_X1 pe_1_3_6_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_3_6_N61), .SE(1'b0), .GCK(pe_1_3_6_net5197) );
  CLKGATETST_X1 pe_1_3_6_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_3_6_N60), .SE(1'b0), .GCK(pe_1_3_6_net5202) );
  CLKGATETST_X1 pe_1_3_6_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_3_6_N59), .SE(1'b0), .GCK(pe_1_3_6_net5207) );
  CLKGATETST_X1 pe_1_3_6_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_3_6_N90), .SE(1'b0), .GCK(pe_1_3_6_net5212) );
  CLKBUF_X1 pe_1_3_7_U112 ( .A(pe_1_3_7_n72), .Z(pe_1_3_7_n71) );
  INV_X1 pe_1_3_7_U111 ( .A(n75), .ZN(pe_1_3_7_n70) );
  INV_X1 pe_1_3_7_U110 ( .A(n67), .ZN(pe_1_3_7_n69) );
  INV_X1 pe_1_3_7_U109 ( .A(n67), .ZN(pe_1_3_7_n68) );
  INV_X1 pe_1_3_7_U108 ( .A(n67), .ZN(pe_1_3_7_n67) );
  INV_X1 pe_1_3_7_U107 ( .A(pe_1_3_7_n69), .ZN(pe_1_3_7_n66) );
  INV_X1 pe_1_3_7_U106 ( .A(pe_1_3_7_n63), .ZN(pe_1_3_7_n62) );
  INV_X1 pe_1_3_7_U105 ( .A(pe_1_3_7_n61), .ZN(pe_1_3_7_n60) );
  INV_X1 pe_1_3_7_U104 ( .A(n27), .ZN(pe_1_3_7_n59) );
  INV_X1 pe_1_3_7_U103 ( .A(pe_1_3_7_n59), .ZN(pe_1_3_7_n58) );
  INV_X1 pe_1_3_7_U102 ( .A(n19), .ZN(pe_1_3_7_n57) );
  MUX2_X1 pe_1_3_7_U101 ( .A(pe_1_3_7_n54), .B(pe_1_3_7_n51), .S(n49), .Z(
        int_data_x_3__7__3_) );
  MUX2_X1 pe_1_3_7_U100 ( .A(pe_1_3_7_n53), .B(pe_1_3_7_n52), .S(pe_1_3_7_n62), 
        .Z(pe_1_3_7_n54) );
  MUX2_X1 pe_1_3_7_U99 ( .A(pe_1_3_7_int_q_reg_h[23]), .B(
        pe_1_3_7_int_q_reg_h[19]), .S(pe_1_3_7_n56), .Z(pe_1_3_7_n53) );
  MUX2_X1 pe_1_3_7_U98 ( .A(pe_1_3_7_int_q_reg_h[15]), .B(
        pe_1_3_7_int_q_reg_h[11]), .S(pe_1_3_7_n56), .Z(pe_1_3_7_n52) );
  MUX2_X1 pe_1_3_7_U97 ( .A(pe_1_3_7_int_q_reg_h[7]), .B(
        pe_1_3_7_int_q_reg_h[3]), .S(pe_1_3_7_n56), .Z(pe_1_3_7_n51) );
  MUX2_X1 pe_1_3_7_U96 ( .A(pe_1_3_7_n50), .B(pe_1_3_7_n47), .S(n49), .Z(
        int_data_x_3__7__2_) );
  MUX2_X1 pe_1_3_7_U95 ( .A(pe_1_3_7_n49), .B(pe_1_3_7_n48), .S(pe_1_3_7_n62), 
        .Z(pe_1_3_7_n50) );
  MUX2_X1 pe_1_3_7_U94 ( .A(pe_1_3_7_int_q_reg_h[22]), .B(
        pe_1_3_7_int_q_reg_h[18]), .S(pe_1_3_7_n56), .Z(pe_1_3_7_n49) );
  MUX2_X1 pe_1_3_7_U93 ( .A(pe_1_3_7_int_q_reg_h[14]), .B(
        pe_1_3_7_int_q_reg_h[10]), .S(pe_1_3_7_n56), .Z(pe_1_3_7_n48) );
  MUX2_X1 pe_1_3_7_U92 ( .A(pe_1_3_7_int_q_reg_h[6]), .B(
        pe_1_3_7_int_q_reg_h[2]), .S(pe_1_3_7_n56), .Z(pe_1_3_7_n47) );
  MUX2_X1 pe_1_3_7_U91 ( .A(pe_1_3_7_n46), .B(pe_1_3_7_n24), .S(n49), .Z(
        int_data_x_3__7__1_) );
  MUX2_X1 pe_1_3_7_U90 ( .A(pe_1_3_7_n45), .B(pe_1_3_7_n25), .S(pe_1_3_7_n62), 
        .Z(pe_1_3_7_n46) );
  MUX2_X1 pe_1_3_7_U89 ( .A(pe_1_3_7_int_q_reg_h[21]), .B(
        pe_1_3_7_int_q_reg_h[17]), .S(pe_1_3_7_n56), .Z(pe_1_3_7_n45) );
  MUX2_X1 pe_1_3_7_U88 ( .A(pe_1_3_7_int_q_reg_h[13]), .B(
        pe_1_3_7_int_q_reg_h[9]), .S(pe_1_3_7_n56), .Z(pe_1_3_7_n25) );
  MUX2_X1 pe_1_3_7_U87 ( .A(pe_1_3_7_int_q_reg_h[5]), .B(
        pe_1_3_7_int_q_reg_h[1]), .S(pe_1_3_7_n56), .Z(pe_1_3_7_n24) );
  MUX2_X1 pe_1_3_7_U86 ( .A(pe_1_3_7_n23), .B(pe_1_3_7_n20), .S(n49), .Z(
        int_data_x_3__7__0_) );
  MUX2_X1 pe_1_3_7_U85 ( .A(pe_1_3_7_n22), .B(pe_1_3_7_n21), .S(pe_1_3_7_n62), 
        .Z(pe_1_3_7_n23) );
  MUX2_X1 pe_1_3_7_U84 ( .A(pe_1_3_7_int_q_reg_h[20]), .B(
        pe_1_3_7_int_q_reg_h[16]), .S(pe_1_3_7_n56), .Z(pe_1_3_7_n22) );
  MUX2_X1 pe_1_3_7_U83 ( .A(pe_1_3_7_int_q_reg_h[12]), .B(
        pe_1_3_7_int_q_reg_h[8]), .S(pe_1_3_7_n56), .Z(pe_1_3_7_n21) );
  MUX2_X1 pe_1_3_7_U82 ( .A(pe_1_3_7_int_q_reg_h[4]), .B(
        pe_1_3_7_int_q_reg_h[0]), .S(pe_1_3_7_n56), .Z(pe_1_3_7_n20) );
  MUX2_X1 pe_1_3_7_U81 ( .A(pe_1_3_7_n19), .B(pe_1_3_7_n16), .S(n49), .Z(
        int_data_y_3__7__3_) );
  MUX2_X1 pe_1_3_7_U80 ( .A(pe_1_3_7_n18), .B(pe_1_3_7_n17), .S(pe_1_3_7_n62), 
        .Z(pe_1_3_7_n19) );
  MUX2_X1 pe_1_3_7_U79 ( .A(pe_1_3_7_int_q_reg_v[23]), .B(
        pe_1_3_7_int_q_reg_v[19]), .S(pe_1_3_7_n55), .Z(pe_1_3_7_n18) );
  MUX2_X1 pe_1_3_7_U78 ( .A(pe_1_3_7_int_q_reg_v[15]), .B(
        pe_1_3_7_int_q_reg_v[11]), .S(pe_1_3_7_n55), .Z(pe_1_3_7_n17) );
  MUX2_X1 pe_1_3_7_U77 ( .A(pe_1_3_7_int_q_reg_v[7]), .B(
        pe_1_3_7_int_q_reg_v[3]), .S(pe_1_3_7_n55), .Z(pe_1_3_7_n16) );
  MUX2_X1 pe_1_3_7_U76 ( .A(pe_1_3_7_n15), .B(pe_1_3_7_n12), .S(n49), .Z(
        int_data_y_3__7__2_) );
  MUX2_X1 pe_1_3_7_U75 ( .A(pe_1_3_7_n14), .B(pe_1_3_7_n13), .S(pe_1_3_7_n62), 
        .Z(pe_1_3_7_n15) );
  MUX2_X1 pe_1_3_7_U74 ( .A(pe_1_3_7_int_q_reg_v[22]), .B(
        pe_1_3_7_int_q_reg_v[18]), .S(pe_1_3_7_n55), .Z(pe_1_3_7_n14) );
  MUX2_X1 pe_1_3_7_U73 ( .A(pe_1_3_7_int_q_reg_v[14]), .B(
        pe_1_3_7_int_q_reg_v[10]), .S(pe_1_3_7_n55), .Z(pe_1_3_7_n13) );
  MUX2_X1 pe_1_3_7_U72 ( .A(pe_1_3_7_int_q_reg_v[6]), .B(
        pe_1_3_7_int_q_reg_v[2]), .S(pe_1_3_7_n55), .Z(pe_1_3_7_n12) );
  MUX2_X1 pe_1_3_7_U71 ( .A(pe_1_3_7_n11), .B(pe_1_3_7_n8), .S(n49), .Z(
        int_data_y_3__7__1_) );
  MUX2_X1 pe_1_3_7_U70 ( .A(pe_1_3_7_n10), .B(pe_1_3_7_n9), .S(pe_1_3_7_n62), 
        .Z(pe_1_3_7_n11) );
  MUX2_X1 pe_1_3_7_U69 ( .A(pe_1_3_7_int_q_reg_v[21]), .B(
        pe_1_3_7_int_q_reg_v[17]), .S(pe_1_3_7_n55), .Z(pe_1_3_7_n10) );
  MUX2_X1 pe_1_3_7_U68 ( .A(pe_1_3_7_int_q_reg_v[13]), .B(
        pe_1_3_7_int_q_reg_v[9]), .S(pe_1_3_7_n55), .Z(pe_1_3_7_n9) );
  MUX2_X1 pe_1_3_7_U67 ( .A(pe_1_3_7_int_q_reg_v[5]), .B(
        pe_1_3_7_int_q_reg_v[1]), .S(pe_1_3_7_n55), .Z(pe_1_3_7_n8) );
  MUX2_X1 pe_1_3_7_U66 ( .A(pe_1_3_7_n7), .B(pe_1_3_7_n4), .S(n49), .Z(
        int_data_y_3__7__0_) );
  MUX2_X1 pe_1_3_7_U65 ( .A(pe_1_3_7_n6), .B(pe_1_3_7_n5), .S(pe_1_3_7_n62), 
        .Z(pe_1_3_7_n7) );
  MUX2_X1 pe_1_3_7_U64 ( .A(pe_1_3_7_int_q_reg_v[20]), .B(
        pe_1_3_7_int_q_reg_v[16]), .S(pe_1_3_7_n55), .Z(pe_1_3_7_n6) );
  MUX2_X1 pe_1_3_7_U63 ( .A(pe_1_3_7_int_q_reg_v[12]), .B(
        pe_1_3_7_int_q_reg_v[8]), .S(pe_1_3_7_n55), .Z(pe_1_3_7_n5) );
  MUX2_X1 pe_1_3_7_U62 ( .A(pe_1_3_7_int_q_reg_v[4]), .B(
        pe_1_3_7_int_q_reg_v[0]), .S(pe_1_3_7_n55), .Z(pe_1_3_7_n4) );
  AOI222_X1 pe_1_3_7_U61 ( .A1(int_data_res_4__7__2_), .A2(pe_1_3_7_n64), .B1(
        pe_1_3_7_N80), .B2(pe_1_3_7_n27), .C1(pe_1_3_7_N72), .C2(pe_1_3_7_n28), 
        .ZN(pe_1_3_7_n33) );
  INV_X1 pe_1_3_7_U60 ( .A(pe_1_3_7_n33), .ZN(pe_1_3_7_n82) );
  AOI222_X1 pe_1_3_7_U59 ( .A1(int_data_res_4__7__6_), .A2(pe_1_3_7_n64), .B1(
        pe_1_3_7_N84), .B2(pe_1_3_7_n27), .C1(pe_1_3_7_N76), .C2(pe_1_3_7_n28), 
        .ZN(pe_1_3_7_n29) );
  INV_X1 pe_1_3_7_U58 ( .A(pe_1_3_7_n29), .ZN(pe_1_3_7_n78) );
  XNOR2_X1 pe_1_3_7_U57 ( .A(pe_1_3_7_n73), .B(int_data_res_3__7__0_), .ZN(
        pe_1_3_7_N70) );
  AOI222_X1 pe_1_3_7_U52 ( .A1(int_data_res_4__7__0_), .A2(pe_1_3_7_n64), .B1(
        pe_1_3_7_n1), .B2(pe_1_3_7_n27), .C1(pe_1_3_7_N70), .C2(pe_1_3_7_n28), 
        .ZN(pe_1_3_7_n35) );
  INV_X1 pe_1_3_7_U51 ( .A(pe_1_3_7_n35), .ZN(pe_1_3_7_n84) );
  AOI222_X1 pe_1_3_7_U50 ( .A1(int_data_res_4__7__1_), .A2(pe_1_3_7_n64), .B1(
        pe_1_3_7_N79), .B2(pe_1_3_7_n27), .C1(pe_1_3_7_N71), .C2(pe_1_3_7_n28), 
        .ZN(pe_1_3_7_n34) );
  INV_X1 pe_1_3_7_U49 ( .A(pe_1_3_7_n34), .ZN(pe_1_3_7_n83) );
  AOI222_X1 pe_1_3_7_U48 ( .A1(int_data_res_4__7__3_), .A2(pe_1_3_7_n64), .B1(
        pe_1_3_7_N81), .B2(pe_1_3_7_n27), .C1(pe_1_3_7_N73), .C2(pe_1_3_7_n28), 
        .ZN(pe_1_3_7_n32) );
  INV_X1 pe_1_3_7_U47 ( .A(pe_1_3_7_n32), .ZN(pe_1_3_7_n81) );
  AOI222_X1 pe_1_3_7_U46 ( .A1(int_data_res_4__7__4_), .A2(pe_1_3_7_n64), .B1(
        pe_1_3_7_N82), .B2(pe_1_3_7_n27), .C1(pe_1_3_7_N74), .C2(pe_1_3_7_n28), 
        .ZN(pe_1_3_7_n31) );
  INV_X1 pe_1_3_7_U45 ( .A(pe_1_3_7_n31), .ZN(pe_1_3_7_n80) );
  AOI222_X1 pe_1_3_7_U44 ( .A1(int_data_res_4__7__5_), .A2(pe_1_3_7_n64), .B1(
        pe_1_3_7_N83), .B2(pe_1_3_7_n27), .C1(pe_1_3_7_N75), .C2(pe_1_3_7_n28), 
        .ZN(pe_1_3_7_n30) );
  INV_X1 pe_1_3_7_U43 ( .A(pe_1_3_7_n30), .ZN(pe_1_3_7_n79) );
  NAND2_X1 pe_1_3_7_U42 ( .A1(pe_1_3_7_int_data_0_), .A2(pe_1_3_7_n3), .ZN(
        pe_1_3_7_sub_81_carry[1]) );
  INV_X1 pe_1_3_7_U41 ( .A(pe_1_3_7_int_data_1_), .ZN(pe_1_3_7_n74) );
  INV_X1 pe_1_3_7_U40 ( .A(pe_1_3_7_int_data_2_), .ZN(pe_1_3_7_n75) );
  AND2_X1 pe_1_3_7_U39 ( .A1(pe_1_3_7_int_data_0_), .A2(int_data_res_3__7__0_), 
        .ZN(pe_1_3_7_n2) );
  AOI222_X1 pe_1_3_7_U38 ( .A1(pe_1_3_7_n64), .A2(int_data_res_4__7__7_), .B1(
        pe_1_3_7_N85), .B2(pe_1_3_7_n27), .C1(pe_1_3_7_N77), .C2(pe_1_3_7_n28), 
        .ZN(pe_1_3_7_n26) );
  INV_X1 pe_1_3_7_U37 ( .A(pe_1_3_7_n26), .ZN(pe_1_3_7_n77) );
  NOR3_X1 pe_1_3_7_U36 ( .A1(pe_1_3_7_n59), .A2(pe_1_3_7_n65), .A3(int_ckg[32]), .ZN(pe_1_3_7_n36) );
  OR2_X1 pe_1_3_7_U35 ( .A1(pe_1_3_7_n36), .A2(pe_1_3_7_n64), .ZN(pe_1_3_7_N90) );
  INV_X1 pe_1_3_7_U34 ( .A(n39), .ZN(pe_1_3_7_n63) );
  AND2_X1 pe_1_3_7_U33 ( .A1(int_data_x_3__7__2_), .A2(pe_1_3_7_n58), .ZN(
        pe_1_3_7_int_data_2_) );
  AND2_X1 pe_1_3_7_U32 ( .A1(int_data_x_3__7__1_), .A2(pe_1_3_7_n58), .ZN(
        pe_1_3_7_int_data_1_) );
  AND2_X1 pe_1_3_7_U31 ( .A1(int_data_x_3__7__3_), .A2(pe_1_3_7_n58), .ZN(
        pe_1_3_7_int_data_3_) );
  BUF_X1 pe_1_3_7_U30 ( .A(n61), .Z(pe_1_3_7_n64) );
  INV_X1 pe_1_3_7_U29 ( .A(n33), .ZN(pe_1_3_7_n61) );
  AND2_X1 pe_1_3_7_U28 ( .A1(int_data_x_3__7__0_), .A2(pe_1_3_7_n58), .ZN(
        pe_1_3_7_int_data_0_) );
  NAND2_X1 pe_1_3_7_U27 ( .A1(pe_1_3_7_n44), .A2(pe_1_3_7_n61), .ZN(
        pe_1_3_7_n41) );
  AND3_X1 pe_1_3_7_U26 ( .A1(n75), .A2(pe_1_3_7_n63), .A3(n49), .ZN(
        pe_1_3_7_n44) );
  INV_X1 pe_1_3_7_U25 ( .A(pe_1_3_7_int_data_3_), .ZN(pe_1_3_7_n76) );
  NOR2_X1 pe_1_3_7_U24 ( .A1(pe_1_3_7_n70), .A2(n49), .ZN(pe_1_3_7_n43) );
  NOR2_X1 pe_1_3_7_U23 ( .A1(pe_1_3_7_n57), .A2(pe_1_3_7_n64), .ZN(
        pe_1_3_7_n28) );
  NOR2_X1 pe_1_3_7_U22 ( .A1(n19), .A2(pe_1_3_7_n64), .ZN(pe_1_3_7_n27) );
  INV_X1 pe_1_3_7_U21 ( .A(pe_1_3_7_int_data_0_), .ZN(pe_1_3_7_n73) );
  INV_X1 pe_1_3_7_U20 ( .A(pe_1_3_7_n41), .ZN(pe_1_3_7_n90) );
  INV_X1 pe_1_3_7_U19 ( .A(pe_1_3_7_n37), .ZN(pe_1_3_7_n88) );
  INV_X1 pe_1_3_7_U18 ( .A(pe_1_3_7_n38), .ZN(pe_1_3_7_n87) );
  INV_X1 pe_1_3_7_U17 ( .A(pe_1_3_7_n39), .ZN(pe_1_3_7_n86) );
  NOR2_X1 pe_1_3_7_U16 ( .A1(pe_1_3_7_n68), .A2(pe_1_3_7_n42), .ZN(
        pe_1_3_7_N59) );
  NOR2_X1 pe_1_3_7_U15 ( .A1(pe_1_3_7_n68), .A2(pe_1_3_7_n41), .ZN(
        pe_1_3_7_N60) );
  NOR2_X1 pe_1_3_7_U14 ( .A1(pe_1_3_7_n68), .A2(pe_1_3_7_n38), .ZN(
        pe_1_3_7_N63) );
  NOR2_X1 pe_1_3_7_U13 ( .A1(pe_1_3_7_n67), .A2(pe_1_3_7_n40), .ZN(
        pe_1_3_7_N61) );
  NOR2_X1 pe_1_3_7_U12 ( .A1(pe_1_3_7_n67), .A2(pe_1_3_7_n39), .ZN(
        pe_1_3_7_N62) );
  NOR2_X1 pe_1_3_7_U11 ( .A1(pe_1_3_7_n37), .A2(pe_1_3_7_n67), .ZN(
        pe_1_3_7_N64) );
  NAND2_X1 pe_1_3_7_U10 ( .A1(pe_1_3_7_n44), .A2(pe_1_3_7_n60), .ZN(
        pe_1_3_7_n42) );
  BUF_X1 pe_1_3_7_U9 ( .A(pe_1_3_7_n60), .Z(pe_1_3_7_n55) );
  INV_X1 pe_1_3_7_U8 ( .A(pe_1_3_7_n69), .ZN(pe_1_3_7_n65) );
  BUF_X1 pe_1_3_7_U7 ( .A(pe_1_3_7_n60), .Z(pe_1_3_7_n56) );
  INV_X1 pe_1_3_7_U6 ( .A(pe_1_3_7_n42), .ZN(pe_1_3_7_n89) );
  INV_X1 pe_1_3_7_U5 ( .A(pe_1_3_7_n40), .ZN(pe_1_3_7_n85) );
  INV_X2 pe_1_3_7_U4 ( .A(n83), .ZN(pe_1_3_7_n72) );
  XOR2_X1 pe_1_3_7_U3 ( .A(pe_1_3_7_int_data_0_), .B(int_data_res_3__7__0_), 
        .Z(pe_1_3_7_n1) );
  DFFR_X1 pe_1_3_7_int_q_acc_reg_0_ ( .D(pe_1_3_7_n84), .CK(pe_1_3_7_net5134), 
        .RN(pe_1_3_7_n72), .Q(int_data_res_3__7__0_), .QN(pe_1_3_7_n3) );
  DFFR_X1 pe_1_3_7_int_q_reg_v_reg_0__0_ ( .D(int_data_y_4__7__0_), .CK(
        pe_1_3_7_net5104), .RN(pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_v[20]) );
  DFFR_X1 pe_1_3_7_int_q_reg_v_reg_0__1_ ( .D(int_data_y_4__7__1_), .CK(
        pe_1_3_7_net5104), .RN(pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_v[21]) );
  DFFR_X1 pe_1_3_7_int_q_reg_v_reg_0__2_ ( .D(int_data_y_4__7__2_), .CK(
        pe_1_3_7_net5104), .RN(pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_v[22]) );
  DFFR_X1 pe_1_3_7_int_q_reg_v_reg_0__3_ ( .D(int_data_y_4__7__3_), .CK(
        pe_1_3_7_net5104), .RN(pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_v[23]) );
  DFFR_X1 pe_1_3_7_int_q_reg_v_reg_1__0_ ( .D(int_data_y_4__7__0_), .CK(
        pe_1_3_7_net5109), .RN(pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_v[16]) );
  DFFR_X1 pe_1_3_7_int_q_reg_v_reg_1__1_ ( .D(int_data_y_4__7__1_), .CK(
        pe_1_3_7_net5109), .RN(pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_v[17]) );
  DFFR_X1 pe_1_3_7_int_q_reg_v_reg_1__2_ ( .D(int_data_y_4__7__2_), .CK(
        pe_1_3_7_net5109), .RN(pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_v[18]) );
  DFFR_X1 pe_1_3_7_int_q_reg_v_reg_1__3_ ( .D(int_data_y_4__7__3_), .CK(
        pe_1_3_7_net5109), .RN(pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_v[19]) );
  DFFR_X1 pe_1_3_7_int_q_reg_v_reg_2__0_ ( .D(int_data_y_4__7__0_), .CK(
        pe_1_3_7_net5114), .RN(pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_v[12]) );
  DFFR_X1 pe_1_3_7_int_q_reg_v_reg_2__1_ ( .D(int_data_y_4__7__1_), .CK(
        pe_1_3_7_net5114), .RN(pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_v[13]) );
  DFFR_X1 pe_1_3_7_int_q_reg_v_reg_2__2_ ( .D(int_data_y_4__7__2_), .CK(
        pe_1_3_7_net5114), .RN(pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_v[14]) );
  DFFR_X1 pe_1_3_7_int_q_reg_v_reg_2__3_ ( .D(int_data_y_4__7__3_), .CK(
        pe_1_3_7_net5114), .RN(pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_v[15]) );
  DFFR_X1 pe_1_3_7_int_q_reg_v_reg_3__0_ ( .D(int_data_y_4__7__0_), .CK(
        pe_1_3_7_net5119), .RN(pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_v[8]) );
  DFFR_X1 pe_1_3_7_int_q_reg_v_reg_3__1_ ( .D(int_data_y_4__7__1_), .CK(
        pe_1_3_7_net5119), .RN(pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_v[9]) );
  DFFR_X1 pe_1_3_7_int_q_reg_v_reg_3__2_ ( .D(int_data_y_4__7__2_), .CK(
        pe_1_3_7_net5119), .RN(pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_v[10]) );
  DFFR_X1 pe_1_3_7_int_q_reg_v_reg_3__3_ ( .D(int_data_y_4__7__3_), .CK(
        pe_1_3_7_net5119), .RN(pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_v[11]) );
  DFFR_X1 pe_1_3_7_int_q_reg_v_reg_4__0_ ( .D(int_data_y_4__7__0_), .CK(
        pe_1_3_7_net5124), .RN(pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_v[4]) );
  DFFR_X1 pe_1_3_7_int_q_reg_v_reg_4__1_ ( .D(int_data_y_4__7__1_), .CK(
        pe_1_3_7_net5124), .RN(pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_v[5]) );
  DFFR_X1 pe_1_3_7_int_q_reg_v_reg_4__2_ ( .D(int_data_y_4__7__2_), .CK(
        pe_1_3_7_net5124), .RN(pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_v[6]) );
  DFFR_X1 pe_1_3_7_int_q_reg_v_reg_4__3_ ( .D(int_data_y_4__7__3_), .CK(
        pe_1_3_7_net5124), .RN(pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_v[7]) );
  DFFR_X1 pe_1_3_7_int_q_reg_v_reg_5__0_ ( .D(int_data_y_4__7__0_), .CK(
        pe_1_3_7_net5129), .RN(pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_v[0]) );
  DFFR_X1 pe_1_3_7_int_q_reg_v_reg_5__1_ ( .D(int_data_y_4__7__1_), .CK(
        pe_1_3_7_net5129), .RN(pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_v[1]) );
  DFFR_X1 pe_1_3_7_int_q_reg_v_reg_5__2_ ( .D(int_data_y_4__7__2_), .CK(
        pe_1_3_7_net5129), .RN(pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_v[2]) );
  DFFR_X1 pe_1_3_7_int_q_reg_v_reg_5__3_ ( .D(int_data_y_4__7__3_), .CK(
        pe_1_3_7_net5129), .RN(pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_3_7_int_q_reg_h_reg_0__0_ ( .D(i_data_conv_h[16]), .SI(
        int_data_y_4__7__0_), .SE(pe_1_3_7_n65), .CK(pe_1_3_7_net5073), .RN(
        pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_3_7_int_q_reg_h_reg_0__1_ ( .D(i_data_conv_h[17]), .SI(
        int_data_y_4__7__1_), .SE(pe_1_3_7_n65), .CK(pe_1_3_7_net5073), .RN(
        pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_3_7_int_q_reg_h_reg_0__2_ ( .D(i_data_conv_h[18]), .SI(
        int_data_y_4__7__2_), .SE(pe_1_3_7_n65), .CK(pe_1_3_7_net5073), .RN(
        pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_3_7_int_q_reg_h_reg_0__3_ ( .D(i_data_conv_h[19]), .SI(
        int_data_y_4__7__3_), .SE(pe_1_3_7_n65), .CK(pe_1_3_7_net5073), .RN(
        pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_3_7_int_q_reg_h_reg_1__0_ ( .D(i_data_conv_h[16]), .SI(
        int_data_y_4__7__0_), .SE(pe_1_3_7_n65), .CK(pe_1_3_7_net5079), .RN(
        pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_3_7_int_q_reg_h_reg_1__1_ ( .D(i_data_conv_h[17]), .SI(
        int_data_y_4__7__1_), .SE(pe_1_3_7_n65), .CK(pe_1_3_7_net5079), .RN(
        pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_3_7_int_q_reg_h_reg_1__2_ ( .D(i_data_conv_h[18]), .SI(
        int_data_y_4__7__2_), .SE(pe_1_3_7_n65), .CK(pe_1_3_7_net5079), .RN(
        pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_3_7_int_q_reg_h_reg_1__3_ ( .D(i_data_conv_h[19]), .SI(
        int_data_y_4__7__3_), .SE(pe_1_3_7_n65), .CK(pe_1_3_7_net5079), .RN(
        pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_3_7_int_q_reg_h_reg_2__0_ ( .D(i_data_conv_h[16]), .SI(
        int_data_y_4__7__0_), .SE(pe_1_3_7_n65), .CK(pe_1_3_7_net5084), .RN(
        pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_3_7_int_q_reg_h_reg_2__1_ ( .D(i_data_conv_h[17]), .SI(
        int_data_y_4__7__1_), .SE(pe_1_3_7_n65), .CK(pe_1_3_7_net5084), .RN(
        pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_3_7_int_q_reg_h_reg_2__2_ ( .D(i_data_conv_h[18]), .SI(
        int_data_y_4__7__2_), .SE(pe_1_3_7_n65), .CK(pe_1_3_7_net5084), .RN(
        pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_3_7_int_q_reg_h_reg_2__3_ ( .D(i_data_conv_h[19]), .SI(
        int_data_y_4__7__3_), .SE(pe_1_3_7_n65), .CK(pe_1_3_7_net5084), .RN(
        pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_3_7_int_q_reg_h_reg_3__0_ ( .D(i_data_conv_h[16]), .SI(
        int_data_y_4__7__0_), .SE(pe_1_3_7_n65), .CK(pe_1_3_7_net5089), .RN(
        pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_3_7_int_q_reg_h_reg_3__1_ ( .D(i_data_conv_h[17]), .SI(
        int_data_y_4__7__1_), .SE(pe_1_3_7_n65), .CK(pe_1_3_7_net5089), .RN(
        pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_3_7_int_q_reg_h_reg_3__2_ ( .D(i_data_conv_h[18]), .SI(
        int_data_y_4__7__2_), .SE(pe_1_3_7_n65), .CK(pe_1_3_7_net5089), .RN(
        pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_3_7_int_q_reg_h_reg_3__3_ ( .D(i_data_conv_h[19]), .SI(
        int_data_y_4__7__3_), .SE(pe_1_3_7_n65), .CK(pe_1_3_7_net5089), .RN(
        pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_3_7_int_q_reg_h_reg_4__0_ ( .D(i_data_conv_h[16]), .SI(
        int_data_y_4__7__0_), .SE(pe_1_3_7_n66), .CK(pe_1_3_7_net5094), .RN(
        pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_3_7_int_q_reg_h_reg_4__1_ ( .D(i_data_conv_h[17]), .SI(
        int_data_y_4__7__1_), .SE(pe_1_3_7_n66), .CK(pe_1_3_7_net5094), .RN(
        pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_3_7_int_q_reg_h_reg_4__2_ ( .D(i_data_conv_h[18]), .SI(
        int_data_y_4__7__2_), .SE(pe_1_3_7_n66), .CK(pe_1_3_7_net5094), .RN(
        pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_3_7_int_q_reg_h_reg_4__3_ ( .D(i_data_conv_h[19]), .SI(
        int_data_y_4__7__3_), .SE(pe_1_3_7_n66), .CK(pe_1_3_7_net5094), .RN(
        pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_3_7_int_q_reg_h_reg_5__0_ ( .D(i_data_conv_h[16]), .SI(
        int_data_y_4__7__0_), .SE(pe_1_3_7_n66), .CK(pe_1_3_7_net5099), .RN(
        pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_3_7_int_q_reg_h_reg_5__1_ ( .D(i_data_conv_h[17]), .SI(
        int_data_y_4__7__1_), .SE(pe_1_3_7_n66), .CK(pe_1_3_7_net5099), .RN(
        pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_3_7_int_q_reg_h_reg_5__2_ ( .D(i_data_conv_h[18]), .SI(
        int_data_y_4__7__2_), .SE(pe_1_3_7_n66), .CK(pe_1_3_7_net5099), .RN(
        pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_3_7_int_q_reg_h_reg_5__3_ ( .D(i_data_conv_h[19]), .SI(
        int_data_y_4__7__3_), .SE(pe_1_3_7_n66), .CK(pe_1_3_7_net5099), .RN(
        pe_1_3_7_n72), .Q(pe_1_3_7_int_q_reg_h[3]) );
  FA_X1 pe_1_3_7_sub_81_U2_7 ( .A(int_data_res_3__7__7_), .B(pe_1_3_7_n76), 
        .CI(pe_1_3_7_sub_81_carry[7]), .S(pe_1_3_7_N77) );
  FA_X1 pe_1_3_7_sub_81_U2_6 ( .A(int_data_res_3__7__6_), .B(pe_1_3_7_n76), 
        .CI(pe_1_3_7_sub_81_carry[6]), .CO(pe_1_3_7_sub_81_carry[7]), .S(
        pe_1_3_7_N76) );
  FA_X1 pe_1_3_7_sub_81_U2_5 ( .A(int_data_res_3__7__5_), .B(pe_1_3_7_n76), 
        .CI(pe_1_3_7_sub_81_carry[5]), .CO(pe_1_3_7_sub_81_carry[6]), .S(
        pe_1_3_7_N75) );
  FA_X1 pe_1_3_7_sub_81_U2_4 ( .A(int_data_res_3__7__4_), .B(pe_1_3_7_n76), 
        .CI(pe_1_3_7_sub_81_carry[4]), .CO(pe_1_3_7_sub_81_carry[5]), .S(
        pe_1_3_7_N74) );
  FA_X1 pe_1_3_7_sub_81_U2_3 ( .A(int_data_res_3__7__3_), .B(pe_1_3_7_n76), 
        .CI(pe_1_3_7_sub_81_carry[3]), .CO(pe_1_3_7_sub_81_carry[4]), .S(
        pe_1_3_7_N73) );
  FA_X1 pe_1_3_7_sub_81_U2_2 ( .A(int_data_res_3__7__2_), .B(pe_1_3_7_n75), 
        .CI(pe_1_3_7_sub_81_carry[2]), .CO(pe_1_3_7_sub_81_carry[3]), .S(
        pe_1_3_7_N72) );
  FA_X1 pe_1_3_7_sub_81_U2_1 ( .A(int_data_res_3__7__1_), .B(pe_1_3_7_n74), 
        .CI(pe_1_3_7_sub_81_carry[1]), .CO(pe_1_3_7_sub_81_carry[2]), .S(
        pe_1_3_7_N71) );
  FA_X1 pe_1_3_7_add_83_U1_7 ( .A(int_data_res_3__7__7_), .B(
        pe_1_3_7_int_data_3_), .CI(pe_1_3_7_add_83_carry[7]), .S(pe_1_3_7_N85)
         );
  FA_X1 pe_1_3_7_add_83_U1_6 ( .A(int_data_res_3__7__6_), .B(
        pe_1_3_7_int_data_3_), .CI(pe_1_3_7_add_83_carry[6]), .CO(
        pe_1_3_7_add_83_carry[7]), .S(pe_1_3_7_N84) );
  FA_X1 pe_1_3_7_add_83_U1_5 ( .A(int_data_res_3__7__5_), .B(
        pe_1_3_7_int_data_3_), .CI(pe_1_3_7_add_83_carry[5]), .CO(
        pe_1_3_7_add_83_carry[6]), .S(pe_1_3_7_N83) );
  FA_X1 pe_1_3_7_add_83_U1_4 ( .A(int_data_res_3__7__4_), .B(
        pe_1_3_7_int_data_3_), .CI(pe_1_3_7_add_83_carry[4]), .CO(
        pe_1_3_7_add_83_carry[5]), .S(pe_1_3_7_N82) );
  FA_X1 pe_1_3_7_add_83_U1_3 ( .A(int_data_res_3__7__3_), .B(
        pe_1_3_7_int_data_3_), .CI(pe_1_3_7_add_83_carry[3]), .CO(
        pe_1_3_7_add_83_carry[4]), .S(pe_1_3_7_N81) );
  FA_X1 pe_1_3_7_add_83_U1_2 ( .A(int_data_res_3__7__2_), .B(
        pe_1_3_7_int_data_2_), .CI(pe_1_3_7_add_83_carry[2]), .CO(
        pe_1_3_7_add_83_carry[3]), .S(pe_1_3_7_N80) );
  FA_X1 pe_1_3_7_add_83_U1_1 ( .A(int_data_res_3__7__1_), .B(
        pe_1_3_7_int_data_1_), .CI(pe_1_3_7_n2), .CO(pe_1_3_7_add_83_carry[2]), 
        .S(pe_1_3_7_N79) );
  NAND3_X1 pe_1_3_7_U56 ( .A1(pe_1_3_7_n60), .A2(pe_1_3_7_n43), .A3(
        pe_1_3_7_n62), .ZN(pe_1_3_7_n40) );
  NAND3_X1 pe_1_3_7_U55 ( .A1(pe_1_3_7_n43), .A2(pe_1_3_7_n61), .A3(
        pe_1_3_7_n62), .ZN(pe_1_3_7_n39) );
  NAND3_X1 pe_1_3_7_U54 ( .A1(pe_1_3_7_n43), .A2(pe_1_3_7_n63), .A3(
        pe_1_3_7_n60), .ZN(pe_1_3_7_n38) );
  NAND3_X1 pe_1_3_7_U53 ( .A1(pe_1_3_7_n61), .A2(pe_1_3_7_n63), .A3(
        pe_1_3_7_n43), .ZN(pe_1_3_7_n37) );
  DFFR_X1 pe_1_3_7_int_q_acc_reg_6_ ( .D(pe_1_3_7_n78), .CK(pe_1_3_7_net5134), 
        .RN(pe_1_3_7_n71), .Q(int_data_res_3__7__6_) );
  DFFR_X1 pe_1_3_7_int_q_acc_reg_5_ ( .D(pe_1_3_7_n79), .CK(pe_1_3_7_net5134), 
        .RN(pe_1_3_7_n71), .Q(int_data_res_3__7__5_) );
  DFFR_X1 pe_1_3_7_int_q_acc_reg_4_ ( .D(pe_1_3_7_n80), .CK(pe_1_3_7_net5134), 
        .RN(pe_1_3_7_n71), .Q(int_data_res_3__7__4_) );
  DFFR_X1 pe_1_3_7_int_q_acc_reg_3_ ( .D(pe_1_3_7_n81), .CK(pe_1_3_7_net5134), 
        .RN(pe_1_3_7_n71), .Q(int_data_res_3__7__3_) );
  DFFR_X1 pe_1_3_7_int_q_acc_reg_2_ ( .D(pe_1_3_7_n82), .CK(pe_1_3_7_net5134), 
        .RN(pe_1_3_7_n71), .Q(int_data_res_3__7__2_) );
  DFFR_X1 pe_1_3_7_int_q_acc_reg_1_ ( .D(pe_1_3_7_n83), .CK(pe_1_3_7_net5134), 
        .RN(pe_1_3_7_n71), .Q(int_data_res_3__7__1_) );
  DFFR_X1 pe_1_3_7_int_q_acc_reg_7_ ( .D(pe_1_3_7_n77), .CK(pe_1_3_7_net5134), 
        .RN(pe_1_3_7_n71), .Q(int_data_res_3__7__7_) );
  CLKGATETST_X1 pe_1_3_7_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_3_7_n88), .SE(1'b0), .GCK(pe_1_3_7_net5073) );
  CLKGATETST_X1 pe_1_3_7_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_3_7_n87), .SE(1'b0), .GCK(pe_1_3_7_net5079) );
  CLKGATETST_X1 pe_1_3_7_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_3_7_n86), .SE(1'b0), .GCK(pe_1_3_7_net5084) );
  CLKGATETST_X1 pe_1_3_7_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_3_7_n85), .SE(1'b0), .GCK(pe_1_3_7_net5089) );
  CLKGATETST_X1 pe_1_3_7_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_3_7_n90), .SE(1'b0), .GCK(pe_1_3_7_net5094) );
  CLKGATETST_X1 pe_1_3_7_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_3_7_n89), .SE(1'b0), .GCK(pe_1_3_7_net5099) );
  CLKGATETST_X1 pe_1_3_7_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_3_7_N64), .SE(1'b0), .GCK(pe_1_3_7_net5104) );
  CLKGATETST_X1 pe_1_3_7_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_3_7_N63), .SE(1'b0), .GCK(pe_1_3_7_net5109) );
  CLKGATETST_X1 pe_1_3_7_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_3_7_N62), .SE(1'b0), .GCK(pe_1_3_7_net5114) );
  CLKGATETST_X1 pe_1_3_7_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_3_7_N61), .SE(1'b0), .GCK(pe_1_3_7_net5119) );
  CLKGATETST_X1 pe_1_3_7_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_3_7_N60), .SE(1'b0), .GCK(pe_1_3_7_net5124) );
  CLKGATETST_X1 pe_1_3_7_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_3_7_N59), .SE(1'b0), .GCK(pe_1_3_7_net5129) );
  CLKGATETST_X1 pe_1_3_7_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_3_7_N90), .SE(1'b0), .GCK(pe_1_3_7_net5134) );
  CLKBUF_X1 pe_1_4_0_U112 ( .A(pe_1_4_0_n72), .Z(pe_1_4_0_n71) );
  INV_X1 pe_1_4_0_U111 ( .A(n75), .ZN(pe_1_4_0_n70) );
  INV_X1 pe_1_4_0_U110 ( .A(n67), .ZN(pe_1_4_0_n69) );
  INV_X1 pe_1_4_0_U109 ( .A(n67), .ZN(pe_1_4_0_n68) );
  INV_X1 pe_1_4_0_U108 ( .A(n67), .ZN(pe_1_4_0_n67) );
  INV_X1 pe_1_4_0_U107 ( .A(pe_1_4_0_n69), .ZN(pe_1_4_0_n66) );
  INV_X1 pe_1_4_0_U106 ( .A(pe_1_4_0_n63), .ZN(pe_1_4_0_n62) );
  INV_X1 pe_1_4_0_U105 ( .A(pe_1_4_0_n61), .ZN(pe_1_4_0_n60) );
  INV_X1 pe_1_4_0_U104 ( .A(n27), .ZN(pe_1_4_0_n59) );
  INV_X1 pe_1_4_0_U103 ( .A(pe_1_4_0_n59), .ZN(pe_1_4_0_n58) );
  INV_X1 pe_1_4_0_U102 ( .A(n19), .ZN(pe_1_4_0_n57) );
  MUX2_X1 pe_1_4_0_U101 ( .A(pe_1_4_0_n54), .B(pe_1_4_0_n51), .S(n49), .Z(
        pe_1_4_0_o_data_h_3_) );
  MUX2_X1 pe_1_4_0_U100 ( .A(pe_1_4_0_n53), .B(pe_1_4_0_n52), .S(pe_1_4_0_n62), 
        .Z(pe_1_4_0_n54) );
  MUX2_X1 pe_1_4_0_U99 ( .A(pe_1_4_0_int_q_reg_h[23]), .B(
        pe_1_4_0_int_q_reg_h[19]), .S(pe_1_4_0_n56), .Z(pe_1_4_0_n53) );
  MUX2_X1 pe_1_4_0_U98 ( .A(pe_1_4_0_int_q_reg_h[15]), .B(
        pe_1_4_0_int_q_reg_h[11]), .S(pe_1_4_0_n56), .Z(pe_1_4_0_n52) );
  MUX2_X1 pe_1_4_0_U97 ( .A(pe_1_4_0_int_q_reg_h[7]), .B(
        pe_1_4_0_int_q_reg_h[3]), .S(pe_1_4_0_n56), .Z(pe_1_4_0_n51) );
  MUX2_X1 pe_1_4_0_U96 ( .A(pe_1_4_0_n50), .B(pe_1_4_0_n47), .S(n49), .Z(
        pe_1_4_0_o_data_h_2_) );
  MUX2_X1 pe_1_4_0_U95 ( .A(pe_1_4_0_n49), .B(pe_1_4_0_n48), .S(pe_1_4_0_n62), 
        .Z(pe_1_4_0_n50) );
  MUX2_X1 pe_1_4_0_U94 ( .A(pe_1_4_0_int_q_reg_h[22]), .B(
        pe_1_4_0_int_q_reg_h[18]), .S(pe_1_4_0_n56), .Z(pe_1_4_0_n49) );
  MUX2_X1 pe_1_4_0_U93 ( .A(pe_1_4_0_int_q_reg_h[14]), .B(
        pe_1_4_0_int_q_reg_h[10]), .S(pe_1_4_0_n56), .Z(pe_1_4_0_n48) );
  MUX2_X1 pe_1_4_0_U92 ( .A(pe_1_4_0_int_q_reg_h[6]), .B(
        pe_1_4_0_int_q_reg_h[2]), .S(pe_1_4_0_n56), .Z(pe_1_4_0_n47) );
  MUX2_X1 pe_1_4_0_U91 ( .A(pe_1_4_0_n46), .B(pe_1_4_0_n24), .S(n49), .Z(
        pe_1_4_0_o_data_h_1_) );
  MUX2_X1 pe_1_4_0_U90 ( .A(pe_1_4_0_n45), .B(pe_1_4_0_n25), .S(pe_1_4_0_n62), 
        .Z(pe_1_4_0_n46) );
  MUX2_X1 pe_1_4_0_U89 ( .A(pe_1_4_0_int_q_reg_h[21]), .B(
        pe_1_4_0_int_q_reg_h[17]), .S(pe_1_4_0_n56), .Z(pe_1_4_0_n45) );
  MUX2_X1 pe_1_4_0_U88 ( .A(pe_1_4_0_int_q_reg_h[13]), .B(
        pe_1_4_0_int_q_reg_h[9]), .S(pe_1_4_0_n56), .Z(pe_1_4_0_n25) );
  MUX2_X1 pe_1_4_0_U87 ( .A(pe_1_4_0_int_q_reg_h[5]), .B(
        pe_1_4_0_int_q_reg_h[1]), .S(pe_1_4_0_n56), .Z(pe_1_4_0_n24) );
  MUX2_X1 pe_1_4_0_U86 ( .A(pe_1_4_0_n23), .B(pe_1_4_0_n20), .S(n49), .Z(
        pe_1_4_0_o_data_h_0_) );
  MUX2_X1 pe_1_4_0_U85 ( .A(pe_1_4_0_n22), .B(pe_1_4_0_n21), .S(pe_1_4_0_n62), 
        .Z(pe_1_4_0_n23) );
  MUX2_X1 pe_1_4_0_U84 ( .A(pe_1_4_0_int_q_reg_h[20]), .B(
        pe_1_4_0_int_q_reg_h[16]), .S(pe_1_4_0_n56), .Z(pe_1_4_0_n22) );
  MUX2_X1 pe_1_4_0_U83 ( .A(pe_1_4_0_int_q_reg_h[12]), .B(
        pe_1_4_0_int_q_reg_h[8]), .S(pe_1_4_0_n56), .Z(pe_1_4_0_n21) );
  MUX2_X1 pe_1_4_0_U82 ( .A(pe_1_4_0_int_q_reg_h[4]), .B(
        pe_1_4_0_int_q_reg_h[0]), .S(pe_1_4_0_n56), .Z(pe_1_4_0_n20) );
  MUX2_X1 pe_1_4_0_U81 ( .A(pe_1_4_0_n19), .B(pe_1_4_0_n16), .S(n49), .Z(
        int_data_y_4__0__3_) );
  MUX2_X1 pe_1_4_0_U80 ( .A(pe_1_4_0_n18), .B(pe_1_4_0_n17), .S(pe_1_4_0_n62), 
        .Z(pe_1_4_0_n19) );
  MUX2_X1 pe_1_4_0_U79 ( .A(pe_1_4_0_int_q_reg_v[23]), .B(
        pe_1_4_0_int_q_reg_v[19]), .S(pe_1_4_0_n55), .Z(pe_1_4_0_n18) );
  MUX2_X1 pe_1_4_0_U78 ( .A(pe_1_4_0_int_q_reg_v[15]), .B(
        pe_1_4_0_int_q_reg_v[11]), .S(pe_1_4_0_n55), .Z(pe_1_4_0_n17) );
  MUX2_X1 pe_1_4_0_U77 ( .A(pe_1_4_0_int_q_reg_v[7]), .B(
        pe_1_4_0_int_q_reg_v[3]), .S(pe_1_4_0_n55), .Z(pe_1_4_0_n16) );
  MUX2_X1 pe_1_4_0_U76 ( .A(pe_1_4_0_n15), .B(pe_1_4_0_n12), .S(n49), .Z(
        int_data_y_4__0__2_) );
  MUX2_X1 pe_1_4_0_U75 ( .A(pe_1_4_0_n14), .B(pe_1_4_0_n13), .S(pe_1_4_0_n62), 
        .Z(pe_1_4_0_n15) );
  MUX2_X1 pe_1_4_0_U74 ( .A(pe_1_4_0_int_q_reg_v[22]), .B(
        pe_1_4_0_int_q_reg_v[18]), .S(pe_1_4_0_n55), .Z(pe_1_4_0_n14) );
  MUX2_X1 pe_1_4_0_U73 ( .A(pe_1_4_0_int_q_reg_v[14]), .B(
        pe_1_4_0_int_q_reg_v[10]), .S(pe_1_4_0_n55), .Z(pe_1_4_0_n13) );
  MUX2_X1 pe_1_4_0_U72 ( .A(pe_1_4_0_int_q_reg_v[6]), .B(
        pe_1_4_0_int_q_reg_v[2]), .S(pe_1_4_0_n55), .Z(pe_1_4_0_n12) );
  MUX2_X1 pe_1_4_0_U71 ( .A(pe_1_4_0_n11), .B(pe_1_4_0_n8), .S(n49), .Z(
        int_data_y_4__0__1_) );
  MUX2_X1 pe_1_4_0_U70 ( .A(pe_1_4_0_n10), .B(pe_1_4_0_n9), .S(pe_1_4_0_n62), 
        .Z(pe_1_4_0_n11) );
  MUX2_X1 pe_1_4_0_U69 ( .A(pe_1_4_0_int_q_reg_v[21]), .B(
        pe_1_4_0_int_q_reg_v[17]), .S(pe_1_4_0_n55), .Z(pe_1_4_0_n10) );
  MUX2_X1 pe_1_4_0_U68 ( .A(pe_1_4_0_int_q_reg_v[13]), .B(
        pe_1_4_0_int_q_reg_v[9]), .S(pe_1_4_0_n55), .Z(pe_1_4_0_n9) );
  MUX2_X1 pe_1_4_0_U67 ( .A(pe_1_4_0_int_q_reg_v[5]), .B(
        pe_1_4_0_int_q_reg_v[1]), .S(pe_1_4_0_n55), .Z(pe_1_4_0_n8) );
  MUX2_X1 pe_1_4_0_U66 ( .A(pe_1_4_0_n7), .B(pe_1_4_0_n4), .S(n49), .Z(
        int_data_y_4__0__0_) );
  MUX2_X1 pe_1_4_0_U65 ( .A(pe_1_4_0_n6), .B(pe_1_4_0_n5), .S(pe_1_4_0_n62), 
        .Z(pe_1_4_0_n7) );
  MUX2_X1 pe_1_4_0_U64 ( .A(pe_1_4_0_int_q_reg_v[20]), .B(
        pe_1_4_0_int_q_reg_v[16]), .S(pe_1_4_0_n55), .Z(pe_1_4_0_n6) );
  MUX2_X1 pe_1_4_0_U63 ( .A(pe_1_4_0_int_q_reg_v[12]), .B(
        pe_1_4_0_int_q_reg_v[8]), .S(pe_1_4_0_n55), .Z(pe_1_4_0_n5) );
  MUX2_X1 pe_1_4_0_U62 ( .A(pe_1_4_0_int_q_reg_v[4]), .B(
        pe_1_4_0_int_q_reg_v[0]), .S(pe_1_4_0_n55), .Z(pe_1_4_0_n4) );
  AND2_X1 pe_1_4_0_U61 ( .A1(pe_1_4_0_o_data_h_3_), .A2(pe_1_4_0_n58), .ZN(
        pe_1_4_0_int_data_3_) );
  NAND2_X1 pe_1_4_0_U60 ( .A1(pe_1_4_0_int_data_0_), .A2(pe_1_4_0_n3), .ZN(
        pe_1_4_0_sub_81_carry[1]) );
  INV_X1 pe_1_4_0_U59 ( .A(pe_1_4_0_int_data_1_), .ZN(pe_1_4_0_n74) );
  AOI222_X1 pe_1_4_0_U58 ( .A1(pe_1_4_0_n64), .A2(int_data_res_5__0__7_), .B1(
        pe_1_4_0_N85), .B2(pe_1_4_0_n27), .C1(pe_1_4_0_N77), .C2(pe_1_4_0_n28), 
        .ZN(pe_1_4_0_n26) );
  INV_X1 pe_1_4_0_U57 ( .A(pe_1_4_0_n26), .ZN(pe_1_4_0_n77) );
  AOI222_X1 pe_1_4_0_U52 ( .A1(int_data_res_5__0__1_), .A2(pe_1_4_0_n64), .B1(
        pe_1_4_0_N79), .B2(pe_1_4_0_n27), .C1(pe_1_4_0_N71), .C2(pe_1_4_0_n28), 
        .ZN(pe_1_4_0_n34) );
  INV_X1 pe_1_4_0_U51 ( .A(pe_1_4_0_n34), .ZN(pe_1_4_0_n83) );
  AOI222_X1 pe_1_4_0_U50 ( .A1(int_data_res_5__0__2_), .A2(pe_1_4_0_n64), .B1(
        pe_1_4_0_N80), .B2(pe_1_4_0_n27), .C1(pe_1_4_0_N72), .C2(pe_1_4_0_n28), 
        .ZN(pe_1_4_0_n33) );
  INV_X1 pe_1_4_0_U49 ( .A(pe_1_4_0_n33), .ZN(pe_1_4_0_n82) );
  AOI222_X1 pe_1_4_0_U48 ( .A1(int_data_res_5__0__6_), .A2(pe_1_4_0_n64), .B1(
        pe_1_4_0_N84), .B2(pe_1_4_0_n27), .C1(pe_1_4_0_N76), .C2(pe_1_4_0_n28), 
        .ZN(pe_1_4_0_n29) );
  INV_X1 pe_1_4_0_U47 ( .A(pe_1_4_0_n29), .ZN(pe_1_4_0_n78) );
  AND2_X1 pe_1_4_0_U46 ( .A1(pe_1_4_0_o_data_h_2_), .A2(pe_1_4_0_n58), .ZN(
        pe_1_4_0_int_data_2_) );
  AND2_X1 pe_1_4_0_U45 ( .A1(pe_1_4_0_o_data_h_1_), .A2(pe_1_4_0_n58), .ZN(
        pe_1_4_0_int_data_1_) );
  INV_X1 pe_1_4_0_U44 ( .A(pe_1_4_0_int_data_2_), .ZN(pe_1_4_0_n75) );
  AND2_X1 pe_1_4_0_U43 ( .A1(pe_1_4_0_int_data_0_), .A2(int_data_res_4__0__0_), 
        .ZN(pe_1_4_0_n2) );
  AND2_X1 pe_1_4_0_U42 ( .A1(pe_1_4_0_o_data_h_0_), .A2(pe_1_4_0_n58), .ZN(
        pe_1_4_0_int_data_0_) );
  XNOR2_X1 pe_1_4_0_U41 ( .A(pe_1_4_0_n73), .B(int_data_res_4__0__0_), .ZN(
        pe_1_4_0_N70) );
  AOI222_X1 pe_1_4_0_U40 ( .A1(int_data_res_5__0__0_), .A2(pe_1_4_0_n64), .B1(
        pe_1_4_0_n1), .B2(pe_1_4_0_n27), .C1(pe_1_4_0_N70), .C2(pe_1_4_0_n28), 
        .ZN(pe_1_4_0_n35) );
  INV_X1 pe_1_4_0_U39 ( .A(pe_1_4_0_n35), .ZN(pe_1_4_0_n84) );
  AOI222_X1 pe_1_4_0_U38 ( .A1(int_data_res_5__0__3_), .A2(pe_1_4_0_n64), .B1(
        pe_1_4_0_N81), .B2(pe_1_4_0_n27), .C1(pe_1_4_0_N73), .C2(pe_1_4_0_n28), 
        .ZN(pe_1_4_0_n32) );
  INV_X1 pe_1_4_0_U37 ( .A(pe_1_4_0_n32), .ZN(pe_1_4_0_n81) );
  AOI222_X1 pe_1_4_0_U36 ( .A1(int_data_res_5__0__4_), .A2(pe_1_4_0_n64), .B1(
        pe_1_4_0_N82), .B2(pe_1_4_0_n27), .C1(pe_1_4_0_N74), .C2(pe_1_4_0_n28), 
        .ZN(pe_1_4_0_n31) );
  INV_X1 pe_1_4_0_U35 ( .A(pe_1_4_0_n31), .ZN(pe_1_4_0_n80) );
  AOI222_X1 pe_1_4_0_U34 ( .A1(int_data_res_5__0__5_), .A2(pe_1_4_0_n64), .B1(
        pe_1_4_0_N83), .B2(pe_1_4_0_n27), .C1(pe_1_4_0_N75), .C2(pe_1_4_0_n28), 
        .ZN(pe_1_4_0_n30) );
  INV_X1 pe_1_4_0_U33 ( .A(pe_1_4_0_n30), .ZN(pe_1_4_0_n79) );
  NOR3_X1 pe_1_4_0_U32 ( .A1(pe_1_4_0_n59), .A2(pe_1_4_0_n65), .A3(int_ckg[31]), .ZN(pe_1_4_0_n36) );
  OR2_X1 pe_1_4_0_U31 ( .A1(pe_1_4_0_n36), .A2(pe_1_4_0_n64), .ZN(pe_1_4_0_N90) );
  INV_X1 pe_1_4_0_U30 ( .A(pe_1_4_0_int_data_0_), .ZN(pe_1_4_0_n73) );
  INV_X1 pe_1_4_0_U29 ( .A(n39), .ZN(pe_1_4_0_n63) );
  INV_X1 pe_1_4_0_U28 ( .A(n33), .ZN(pe_1_4_0_n61) );
  INV_X1 pe_1_4_0_U27 ( .A(pe_1_4_0_int_data_3_), .ZN(pe_1_4_0_n76) );
  BUF_X1 pe_1_4_0_U26 ( .A(n61), .Z(pe_1_4_0_n64) );
  NAND2_X1 pe_1_4_0_U25 ( .A1(pe_1_4_0_n44), .A2(pe_1_4_0_n61), .ZN(
        pe_1_4_0_n41) );
  AND3_X1 pe_1_4_0_U24 ( .A1(n75), .A2(pe_1_4_0_n63), .A3(n49), .ZN(
        pe_1_4_0_n44) );
  NOR2_X1 pe_1_4_0_U23 ( .A1(pe_1_4_0_n70), .A2(n49), .ZN(pe_1_4_0_n43) );
  NOR2_X1 pe_1_4_0_U22 ( .A1(pe_1_4_0_n57), .A2(pe_1_4_0_n64), .ZN(
        pe_1_4_0_n28) );
  NOR2_X1 pe_1_4_0_U21 ( .A1(n19), .A2(pe_1_4_0_n64), .ZN(pe_1_4_0_n27) );
  INV_X1 pe_1_4_0_U20 ( .A(pe_1_4_0_n41), .ZN(pe_1_4_0_n90) );
  INV_X1 pe_1_4_0_U19 ( .A(pe_1_4_0_n37), .ZN(pe_1_4_0_n88) );
  INV_X1 pe_1_4_0_U18 ( .A(pe_1_4_0_n38), .ZN(pe_1_4_0_n87) );
  INV_X1 pe_1_4_0_U17 ( .A(pe_1_4_0_n39), .ZN(pe_1_4_0_n86) );
  NOR2_X1 pe_1_4_0_U16 ( .A1(pe_1_4_0_n68), .A2(pe_1_4_0_n42), .ZN(
        pe_1_4_0_N59) );
  NOR2_X1 pe_1_4_0_U15 ( .A1(pe_1_4_0_n68), .A2(pe_1_4_0_n41), .ZN(
        pe_1_4_0_N60) );
  NOR2_X1 pe_1_4_0_U14 ( .A1(pe_1_4_0_n68), .A2(pe_1_4_0_n38), .ZN(
        pe_1_4_0_N63) );
  NOR2_X1 pe_1_4_0_U13 ( .A1(pe_1_4_0_n67), .A2(pe_1_4_0_n40), .ZN(
        pe_1_4_0_N61) );
  NOR2_X1 pe_1_4_0_U12 ( .A1(pe_1_4_0_n67), .A2(pe_1_4_0_n39), .ZN(
        pe_1_4_0_N62) );
  NOR2_X1 pe_1_4_0_U11 ( .A1(pe_1_4_0_n37), .A2(pe_1_4_0_n67), .ZN(
        pe_1_4_0_N64) );
  NAND2_X1 pe_1_4_0_U10 ( .A1(pe_1_4_0_n44), .A2(pe_1_4_0_n60), .ZN(
        pe_1_4_0_n42) );
  BUF_X1 pe_1_4_0_U9 ( .A(pe_1_4_0_n60), .Z(pe_1_4_0_n55) );
  BUF_X1 pe_1_4_0_U8 ( .A(pe_1_4_0_n60), .Z(pe_1_4_0_n56) );
  INV_X1 pe_1_4_0_U7 ( .A(pe_1_4_0_n69), .ZN(pe_1_4_0_n65) );
  INV_X1 pe_1_4_0_U6 ( .A(pe_1_4_0_n42), .ZN(pe_1_4_0_n89) );
  INV_X1 pe_1_4_0_U5 ( .A(pe_1_4_0_n40), .ZN(pe_1_4_0_n85) );
  INV_X2 pe_1_4_0_U4 ( .A(n83), .ZN(pe_1_4_0_n72) );
  XOR2_X1 pe_1_4_0_U3 ( .A(pe_1_4_0_int_data_0_), .B(int_data_res_4__0__0_), 
        .Z(pe_1_4_0_n1) );
  DFFR_X1 pe_1_4_0_int_q_acc_reg_0_ ( .D(pe_1_4_0_n84), .CK(pe_1_4_0_net5056), 
        .RN(pe_1_4_0_n72), .Q(int_data_res_4__0__0_), .QN(pe_1_4_0_n3) );
  DFFR_X1 pe_1_4_0_int_q_reg_v_reg_0__0_ ( .D(int_data_y_5__0__0_), .CK(
        pe_1_4_0_net5026), .RN(pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_v[20]) );
  DFFR_X1 pe_1_4_0_int_q_reg_v_reg_0__1_ ( .D(int_data_y_5__0__1_), .CK(
        pe_1_4_0_net5026), .RN(pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_v[21]) );
  DFFR_X1 pe_1_4_0_int_q_reg_v_reg_0__2_ ( .D(int_data_y_5__0__2_), .CK(
        pe_1_4_0_net5026), .RN(pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_v[22]) );
  DFFR_X1 pe_1_4_0_int_q_reg_v_reg_0__3_ ( .D(int_data_y_5__0__3_), .CK(
        pe_1_4_0_net5026), .RN(pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_v[23]) );
  DFFR_X1 pe_1_4_0_int_q_reg_v_reg_1__0_ ( .D(int_data_y_5__0__0_), .CK(
        pe_1_4_0_net5031), .RN(pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_v[16]) );
  DFFR_X1 pe_1_4_0_int_q_reg_v_reg_1__1_ ( .D(int_data_y_5__0__1_), .CK(
        pe_1_4_0_net5031), .RN(pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_v[17]) );
  DFFR_X1 pe_1_4_0_int_q_reg_v_reg_1__2_ ( .D(int_data_y_5__0__2_), .CK(
        pe_1_4_0_net5031), .RN(pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_v[18]) );
  DFFR_X1 pe_1_4_0_int_q_reg_v_reg_1__3_ ( .D(int_data_y_5__0__3_), .CK(
        pe_1_4_0_net5031), .RN(pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_v[19]) );
  DFFR_X1 pe_1_4_0_int_q_reg_v_reg_2__0_ ( .D(int_data_y_5__0__0_), .CK(
        pe_1_4_0_net5036), .RN(pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_v[12]) );
  DFFR_X1 pe_1_4_0_int_q_reg_v_reg_2__1_ ( .D(int_data_y_5__0__1_), .CK(
        pe_1_4_0_net5036), .RN(pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_v[13]) );
  DFFR_X1 pe_1_4_0_int_q_reg_v_reg_2__2_ ( .D(int_data_y_5__0__2_), .CK(
        pe_1_4_0_net5036), .RN(pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_v[14]) );
  DFFR_X1 pe_1_4_0_int_q_reg_v_reg_2__3_ ( .D(int_data_y_5__0__3_), .CK(
        pe_1_4_0_net5036), .RN(pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_v[15]) );
  DFFR_X1 pe_1_4_0_int_q_reg_v_reg_3__0_ ( .D(int_data_y_5__0__0_), .CK(
        pe_1_4_0_net5041), .RN(pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_v[8]) );
  DFFR_X1 pe_1_4_0_int_q_reg_v_reg_3__1_ ( .D(int_data_y_5__0__1_), .CK(
        pe_1_4_0_net5041), .RN(pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_v[9]) );
  DFFR_X1 pe_1_4_0_int_q_reg_v_reg_3__2_ ( .D(int_data_y_5__0__2_), .CK(
        pe_1_4_0_net5041), .RN(pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_v[10]) );
  DFFR_X1 pe_1_4_0_int_q_reg_v_reg_3__3_ ( .D(int_data_y_5__0__3_), .CK(
        pe_1_4_0_net5041), .RN(pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_v[11]) );
  DFFR_X1 pe_1_4_0_int_q_reg_v_reg_4__0_ ( .D(int_data_y_5__0__0_), .CK(
        pe_1_4_0_net5046), .RN(pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_v[4]) );
  DFFR_X1 pe_1_4_0_int_q_reg_v_reg_4__1_ ( .D(int_data_y_5__0__1_), .CK(
        pe_1_4_0_net5046), .RN(pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_v[5]) );
  DFFR_X1 pe_1_4_0_int_q_reg_v_reg_4__2_ ( .D(int_data_y_5__0__2_), .CK(
        pe_1_4_0_net5046), .RN(pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_v[6]) );
  DFFR_X1 pe_1_4_0_int_q_reg_v_reg_4__3_ ( .D(int_data_y_5__0__3_), .CK(
        pe_1_4_0_net5046), .RN(pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_v[7]) );
  DFFR_X1 pe_1_4_0_int_q_reg_v_reg_5__0_ ( .D(int_data_y_5__0__0_), .CK(
        pe_1_4_0_net5051), .RN(pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_v[0]) );
  DFFR_X1 pe_1_4_0_int_q_reg_v_reg_5__1_ ( .D(int_data_y_5__0__1_), .CK(
        pe_1_4_0_net5051), .RN(pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_v[1]) );
  DFFR_X1 pe_1_4_0_int_q_reg_v_reg_5__2_ ( .D(int_data_y_5__0__2_), .CK(
        pe_1_4_0_net5051), .RN(pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_v[2]) );
  DFFR_X1 pe_1_4_0_int_q_reg_v_reg_5__3_ ( .D(int_data_y_5__0__3_), .CK(
        pe_1_4_0_net5051), .RN(pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_4_0_int_q_reg_h_reg_0__0_ ( .D(int_data_x_4__1__0_), .SI(
        int_data_y_5__0__0_), .SE(pe_1_4_0_n65), .CK(pe_1_4_0_net4995), .RN(
        pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_4_0_int_q_reg_h_reg_0__1_ ( .D(int_data_x_4__1__1_), .SI(
        int_data_y_5__0__1_), .SE(pe_1_4_0_n65), .CK(pe_1_4_0_net4995), .RN(
        pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_4_0_int_q_reg_h_reg_0__2_ ( .D(int_data_x_4__1__2_), .SI(
        int_data_y_5__0__2_), .SE(pe_1_4_0_n65), .CK(pe_1_4_0_net4995), .RN(
        pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_4_0_int_q_reg_h_reg_0__3_ ( .D(int_data_x_4__1__3_), .SI(
        int_data_y_5__0__3_), .SE(pe_1_4_0_n65), .CK(pe_1_4_0_net4995), .RN(
        pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_4_0_int_q_reg_h_reg_1__0_ ( .D(int_data_x_4__1__0_), .SI(
        int_data_y_5__0__0_), .SE(pe_1_4_0_n65), .CK(pe_1_4_0_net5001), .RN(
        pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_4_0_int_q_reg_h_reg_1__1_ ( .D(int_data_x_4__1__1_), .SI(
        int_data_y_5__0__1_), .SE(pe_1_4_0_n65), .CK(pe_1_4_0_net5001), .RN(
        pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_4_0_int_q_reg_h_reg_1__2_ ( .D(int_data_x_4__1__2_), .SI(
        int_data_y_5__0__2_), .SE(pe_1_4_0_n65), .CK(pe_1_4_0_net5001), .RN(
        pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_4_0_int_q_reg_h_reg_1__3_ ( .D(int_data_x_4__1__3_), .SI(
        int_data_y_5__0__3_), .SE(pe_1_4_0_n65), .CK(pe_1_4_0_net5001), .RN(
        pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_4_0_int_q_reg_h_reg_2__0_ ( .D(int_data_x_4__1__0_), .SI(
        int_data_y_5__0__0_), .SE(pe_1_4_0_n65), .CK(pe_1_4_0_net5006), .RN(
        pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_4_0_int_q_reg_h_reg_2__1_ ( .D(int_data_x_4__1__1_), .SI(
        int_data_y_5__0__1_), .SE(pe_1_4_0_n65), .CK(pe_1_4_0_net5006), .RN(
        pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_4_0_int_q_reg_h_reg_2__2_ ( .D(int_data_x_4__1__2_), .SI(
        int_data_y_5__0__2_), .SE(pe_1_4_0_n65), .CK(pe_1_4_0_net5006), .RN(
        pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_4_0_int_q_reg_h_reg_2__3_ ( .D(int_data_x_4__1__3_), .SI(
        int_data_y_5__0__3_), .SE(pe_1_4_0_n65), .CK(pe_1_4_0_net5006), .RN(
        pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_4_0_int_q_reg_h_reg_3__0_ ( .D(int_data_x_4__1__0_), .SI(
        int_data_y_5__0__0_), .SE(pe_1_4_0_n65), .CK(pe_1_4_0_net5011), .RN(
        pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_4_0_int_q_reg_h_reg_3__1_ ( .D(int_data_x_4__1__1_), .SI(
        int_data_y_5__0__1_), .SE(pe_1_4_0_n65), .CK(pe_1_4_0_net5011), .RN(
        pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_4_0_int_q_reg_h_reg_3__2_ ( .D(int_data_x_4__1__2_), .SI(
        int_data_y_5__0__2_), .SE(pe_1_4_0_n65), .CK(pe_1_4_0_net5011), .RN(
        pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_4_0_int_q_reg_h_reg_3__3_ ( .D(int_data_x_4__1__3_), .SI(
        int_data_y_5__0__3_), .SE(pe_1_4_0_n65), .CK(pe_1_4_0_net5011), .RN(
        pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_4_0_int_q_reg_h_reg_4__0_ ( .D(int_data_x_4__1__0_), .SI(
        int_data_y_5__0__0_), .SE(pe_1_4_0_n66), .CK(pe_1_4_0_net5016), .RN(
        pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_4_0_int_q_reg_h_reg_4__1_ ( .D(int_data_x_4__1__1_), .SI(
        int_data_y_5__0__1_), .SE(pe_1_4_0_n66), .CK(pe_1_4_0_net5016), .RN(
        pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_4_0_int_q_reg_h_reg_4__2_ ( .D(int_data_x_4__1__2_), .SI(
        int_data_y_5__0__2_), .SE(pe_1_4_0_n66), .CK(pe_1_4_0_net5016), .RN(
        pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_4_0_int_q_reg_h_reg_4__3_ ( .D(int_data_x_4__1__3_), .SI(
        int_data_y_5__0__3_), .SE(pe_1_4_0_n66), .CK(pe_1_4_0_net5016), .RN(
        pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_4_0_int_q_reg_h_reg_5__0_ ( .D(int_data_x_4__1__0_), .SI(
        int_data_y_5__0__0_), .SE(pe_1_4_0_n66), .CK(pe_1_4_0_net5021), .RN(
        pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_4_0_int_q_reg_h_reg_5__1_ ( .D(int_data_x_4__1__1_), .SI(
        int_data_y_5__0__1_), .SE(pe_1_4_0_n66), .CK(pe_1_4_0_net5021), .RN(
        pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_4_0_int_q_reg_h_reg_5__2_ ( .D(int_data_x_4__1__2_), .SI(
        int_data_y_5__0__2_), .SE(pe_1_4_0_n66), .CK(pe_1_4_0_net5021), .RN(
        pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_4_0_int_q_reg_h_reg_5__3_ ( .D(int_data_x_4__1__3_), .SI(
        int_data_y_5__0__3_), .SE(pe_1_4_0_n66), .CK(pe_1_4_0_net5021), .RN(
        pe_1_4_0_n72), .Q(pe_1_4_0_int_q_reg_h[3]) );
  FA_X1 pe_1_4_0_sub_81_U2_7 ( .A(int_data_res_4__0__7_), .B(pe_1_4_0_n76), 
        .CI(pe_1_4_0_sub_81_carry[7]), .S(pe_1_4_0_N77) );
  FA_X1 pe_1_4_0_sub_81_U2_6 ( .A(int_data_res_4__0__6_), .B(pe_1_4_0_n76), 
        .CI(pe_1_4_0_sub_81_carry[6]), .CO(pe_1_4_0_sub_81_carry[7]), .S(
        pe_1_4_0_N76) );
  FA_X1 pe_1_4_0_sub_81_U2_5 ( .A(int_data_res_4__0__5_), .B(pe_1_4_0_n76), 
        .CI(pe_1_4_0_sub_81_carry[5]), .CO(pe_1_4_0_sub_81_carry[6]), .S(
        pe_1_4_0_N75) );
  FA_X1 pe_1_4_0_sub_81_U2_4 ( .A(int_data_res_4__0__4_), .B(pe_1_4_0_n76), 
        .CI(pe_1_4_0_sub_81_carry[4]), .CO(pe_1_4_0_sub_81_carry[5]), .S(
        pe_1_4_0_N74) );
  FA_X1 pe_1_4_0_sub_81_U2_3 ( .A(int_data_res_4__0__3_), .B(pe_1_4_0_n76), 
        .CI(pe_1_4_0_sub_81_carry[3]), .CO(pe_1_4_0_sub_81_carry[4]), .S(
        pe_1_4_0_N73) );
  FA_X1 pe_1_4_0_sub_81_U2_2 ( .A(int_data_res_4__0__2_), .B(pe_1_4_0_n75), 
        .CI(pe_1_4_0_sub_81_carry[2]), .CO(pe_1_4_0_sub_81_carry[3]), .S(
        pe_1_4_0_N72) );
  FA_X1 pe_1_4_0_sub_81_U2_1 ( .A(int_data_res_4__0__1_), .B(pe_1_4_0_n74), 
        .CI(pe_1_4_0_sub_81_carry[1]), .CO(pe_1_4_0_sub_81_carry[2]), .S(
        pe_1_4_0_N71) );
  FA_X1 pe_1_4_0_add_83_U1_7 ( .A(int_data_res_4__0__7_), .B(
        pe_1_4_0_int_data_3_), .CI(pe_1_4_0_add_83_carry[7]), .S(pe_1_4_0_N85)
         );
  FA_X1 pe_1_4_0_add_83_U1_6 ( .A(int_data_res_4__0__6_), .B(
        pe_1_4_0_int_data_3_), .CI(pe_1_4_0_add_83_carry[6]), .CO(
        pe_1_4_0_add_83_carry[7]), .S(pe_1_4_0_N84) );
  FA_X1 pe_1_4_0_add_83_U1_5 ( .A(int_data_res_4__0__5_), .B(
        pe_1_4_0_int_data_3_), .CI(pe_1_4_0_add_83_carry[5]), .CO(
        pe_1_4_0_add_83_carry[6]), .S(pe_1_4_0_N83) );
  FA_X1 pe_1_4_0_add_83_U1_4 ( .A(int_data_res_4__0__4_), .B(
        pe_1_4_0_int_data_3_), .CI(pe_1_4_0_add_83_carry[4]), .CO(
        pe_1_4_0_add_83_carry[5]), .S(pe_1_4_0_N82) );
  FA_X1 pe_1_4_0_add_83_U1_3 ( .A(int_data_res_4__0__3_), .B(
        pe_1_4_0_int_data_3_), .CI(pe_1_4_0_add_83_carry[3]), .CO(
        pe_1_4_0_add_83_carry[4]), .S(pe_1_4_0_N81) );
  FA_X1 pe_1_4_0_add_83_U1_2 ( .A(int_data_res_4__0__2_), .B(
        pe_1_4_0_int_data_2_), .CI(pe_1_4_0_add_83_carry[2]), .CO(
        pe_1_4_0_add_83_carry[3]), .S(pe_1_4_0_N80) );
  FA_X1 pe_1_4_0_add_83_U1_1 ( .A(int_data_res_4__0__1_), .B(
        pe_1_4_0_int_data_1_), .CI(pe_1_4_0_n2), .CO(pe_1_4_0_add_83_carry[2]), 
        .S(pe_1_4_0_N79) );
  NAND3_X1 pe_1_4_0_U56 ( .A1(pe_1_4_0_n60), .A2(pe_1_4_0_n43), .A3(
        pe_1_4_0_n62), .ZN(pe_1_4_0_n40) );
  NAND3_X1 pe_1_4_0_U55 ( .A1(pe_1_4_0_n43), .A2(pe_1_4_0_n61), .A3(
        pe_1_4_0_n62), .ZN(pe_1_4_0_n39) );
  NAND3_X1 pe_1_4_0_U54 ( .A1(pe_1_4_0_n43), .A2(pe_1_4_0_n63), .A3(
        pe_1_4_0_n60), .ZN(pe_1_4_0_n38) );
  NAND3_X1 pe_1_4_0_U53 ( .A1(pe_1_4_0_n61), .A2(pe_1_4_0_n63), .A3(
        pe_1_4_0_n43), .ZN(pe_1_4_0_n37) );
  DFFR_X1 pe_1_4_0_int_q_acc_reg_6_ ( .D(pe_1_4_0_n78), .CK(pe_1_4_0_net5056), 
        .RN(pe_1_4_0_n71), .Q(int_data_res_4__0__6_) );
  DFFR_X1 pe_1_4_0_int_q_acc_reg_5_ ( .D(pe_1_4_0_n79), .CK(pe_1_4_0_net5056), 
        .RN(pe_1_4_0_n71), .Q(int_data_res_4__0__5_) );
  DFFR_X1 pe_1_4_0_int_q_acc_reg_4_ ( .D(pe_1_4_0_n80), .CK(pe_1_4_0_net5056), 
        .RN(pe_1_4_0_n71), .Q(int_data_res_4__0__4_) );
  DFFR_X1 pe_1_4_0_int_q_acc_reg_3_ ( .D(pe_1_4_0_n81), .CK(pe_1_4_0_net5056), 
        .RN(pe_1_4_0_n71), .Q(int_data_res_4__0__3_) );
  DFFR_X1 pe_1_4_0_int_q_acc_reg_2_ ( .D(pe_1_4_0_n82), .CK(pe_1_4_0_net5056), 
        .RN(pe_1_4_0_n71), .Q(int_data_res_4__0__2_) );
  DFFR_X1 pe_1_4_0_int_q_acc_reg_1_ ( .D(pe_1_4_0_n83), .CK(pe_1_4_0_net5056), 
        .RN(pe_1_4_0_n71), .Q(int_data_res_4__0__1_) );
  DFFR_X1 pe_1_4_0_int_q_acc_reg_7_ ( .D(pe_1_4_0_n77), .CK(pe_1_4_0_net5056), 
        .RN(pe_1_4_0_n71), .Q(int_data_res_4__0__7_) );
  CLKGATETST_X1 pe_1_4_0_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_4_0_n88), .SE(1'b0), .GCK(pe_1_4_0_net4995) );
  CLKGATETST_X1 pe_1_4_0_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_4_0_n87), .SE(1'b0), .GCK(pe_1_4_0_net5001) );
  CLKGATETST_X1 pe_1_4_0_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_4_0_n86), .SE(1'b0), .GCK(pe_1_4_0_net5006) );
  CLKGATETST_X1 pe_1_4_0_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_4_0_n85), .SE(1'b0), .GCK(pe_1_4_0_net5011) );
  CLKGATETST_X1 pe_1_4_0_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_4_0_n90), .SE(1'b0), .GCK(pe_1_4_0_net5016) );
  CLKGATETST_X1 pe_1_4_0_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_4_0_n89), .SE(1'b0), .GCK(pe_1_4_0_net5021) );
  CLKGATETST_X1 pe_1_4_0_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_4_0_N64), .SE(1'b0), .GCK(pe_1_4_0_net5026) );
  CLKGATETST_X1 pe_1_4_0_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_4_0_N63), .SE(1'b0), .GCK(pe_1_4_0_net5031) );
  CLKGATETST_X1 pe_1_4_0_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_4_0_N62), .SE(1'b0), .GCK(pe_1_4_0_net5036) );
  CLKGATETST_X1 pe_1_4_0_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_4_0_N61), .SE(1'b0), .GCK(pe_1_4_0_net5041) );
  CLKGATETST_X1 pe_1_4_0_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_4_0_N60), .SE(1'b0), .GCK(pe_1_4_0_net5046) );
  CLKGATETST_X1 pe_1_4_0_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_4_0_N59), .SE(1'b0), .GCK(pe_1_4_0_net5051) );
  CLKGATETST_X1 pe_1_4_0_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_4_0_N90), .SE(1'b0), .GCK(pe_1_4_0_net5056) );
  CLKBUF_X1 pe_1_4_1_U112 ( .A(pe_1_4_1_n72), .Z(pe_1_4_1_n71) );
  INV_X1 pe_1_4_1_U111 ( .A(n75), .ZN(pe_1_4_1_n70) );
  INV_X1 pe_1_4_1_U110 ( .A(n67), .ZN(pe_1_4_1_n69) );
  INV_X1 pe_1_4_1_U109 ( .A(n67), .ZN(pe_1_4_1_n68) );
  INV_X1 pe_1_4_1_U108 ( .A(n67), .ZN(pe_1_4_1_n67) );
  INV_X1 pe_1_4_1_U107 ( .A(pe_1_4_1_n69), .ZN(pe_1_4_1_n66) );
  INV_X1 pe_1_4_1_U106 ( .A(pe_1_4_1_n63), .ZN(pe_1_4_1_n62) );
  INV_X1 pe_1_4_1_U105 ( .A(pe_1_4_1_n61), .ZN(pe_1_4_1_n60) );
  INV_X1 pe_1_4_1_U104 ( .A(n27), .ZN(pe_1_4_1_n59) );
  INV_X1 pe_1_4_1_U103 ( .A(pe_1_4_1_n59), .ZN(pe_1_4_1_n58) );
  INV_X1 pe_1_4_1_U102 ( .A(n19), .ZN(pe_1_4_1_n57) );
  MUX2_X1 pe_1_4_1_U101 ( .A(pe_1_4_1_n54), .B(pe_1_4_1_n51), .S(n49), .Z(
        int_data_x_4__1__3_) );
  MUX2_X1 pe_1_4_1_U100 ( .A(pe_1_4_1_n53), .B(pe_1_4_1_n52), .S(pe_1_4_1_n62), 
        .Z(pe_1_4_1_n54) );
  MUX2_X1 pe_1_4_1_U99 ( .A(pe_1_4_1_int_q_reg_h[23]), .B(
        pe_1_4_1_int_q_reg_h[19]), .S(pe_1_4_1_n56), .Z(pe_1_4_1_n53) );
  MUX2_X1 pe_1_4_1_U98 ( .A(pe_1_4_1_int_q_reg_h[15]), .B(
        pe_1_4_1_int_q_reg_h[11]), .S(pe_1_4_1_n56), .Z(pe_1_4_1_n52) );
  MUX2_X1 pe_1_4_1_U97 ( .A(pe_1_4_1_int_q_reg_h[7]), .B(
        pe_1_4_1_int_q_reg_h[3]), .S(pe_1_4_1_n56), .Z(pe_1_4_1_n51) );
  MUX2_X1 pe_1_4_1_U96 ( .A(pe_1_4_1_n50), .B(pe_1_4_1_n47), .S(n49), .Z(
        int_data_x_4__1__2_) );
  MUX2_X1 pe_1_4_1_U95 ( .A(pe_1_4_1_n49), .B(pe_1_4_1_n48), .S(pe_1_4_1_n62), 
        .Z(pe_1_4_1_n50) );
  MUX2_X1 pe_1_4_1_U94 ( .A(pe_1_4_1_int_q_reg_h[22]), .B(
        pe_1_4_1_int_q_reg_h[18]), .S(pe_1_4_1_n56), .Z(pe_1_4_1_n49) );
  MUX2_X1 pe_1_4_1_U93 ( .A(pe_1_4_1_int_q_reg_h[14]), .B(
        pe_1_4_1_int_q_reg_h[10]), .S(pe_1_4_1_n56), .Z(pe_1_4_1_n48) );
  MUX2_X1 pe_1_4_1_U92 ( .A(pe_1_4_1_int_q_reg_h[6]), .B(
        pe_1_4_1_int_q_reg_h[2]), .S(pe_1_4_1_n56), .Z(pe_1_4_1_n47) );
  MUX2_X1 pe_1_4_1_U91 ( .A(pe_1_4_1_n46), .B(pe_1_4_1_n24), .S(n49), .Z(
        int_data_x_4__1__1_) );
  MUX2_X1 pe_1_4_1_U90 ( .A(pe_1_4_1_n45), .B(pe_1_4_1_n25), .S(pe_1_4_1_n62), 
        .Z(pe_1_4_1_n46) );
  MUX2_X1 pe_1_4_1_U89 ( .A(pe_1_4_1_int_q_reg_h[21]), .B(
        pe_1_4_1_int_q_reg_h[17]), .S(pe_1_4_1_n56), .Z(pe_1_4_1_n45) );
  MUX2_X1 pe_1_4_1_U88 ( .A(pe_1_4_1_int_q_reg_h[13]), .B(
        pe_1_4_1_int_q_reg_h[9]), .S(pe_1_4_1_n56), .Z(pe_1_4_1_n25) );
  MUX2_X1 pe_1_4_1_U87 ( .A(pe_1_4_1_int_q_reg_h[5]), .B(
        pe_1_4_1_int_q_reg_h[1]), .S(pe_1_4_1_n56), .Z(pe_1_4_1_n24) );
  MUX2_X1 pe_1_4_1_U86 ( .A(pe_1_4_1_n23), .B(pe_1_4_1_n20), .S(n49), .Z(
        int_data_x_4__1__0_) );
  MUX2_X1 pe_1_4_1_U85 ( .A(pe_1_4_1_n22), .B(pe_1_4_1_n21), .S(pe_1_4_1_n62), 
        .Z(pe_1_4_1_n23) );
  MUX2_X1 pe_1_4_1_U84 ( .A(pe_1_4_1_int_q_reg_h[20]), .B(
        pe_1_4_1_int_q_reg_h[16]), .S(pe_1_4_1_n56), .Z(pe_1_4_1_n22) );
  MUX2_X1 pe_1_4_1_U83 ( .A(pe_1_4_1_int_q_reg_h[12]), .B(
        pe_1_4_1_int_q_reg_h[8]), .S(pe_1_4_1_n56), .Z(pe_1_4_1_n21) );
  MUX2_X1 pe_1_4_1_U82 ( .A(pe_1_4_1_int_q_reg_h[4]), .B(
        pe_1_4_1_int_q_reg_h[0]), .S(pe_1_4_1_n56), .Z(pe_1_4_1_n20) );
  MUX2_X1 pe_1_4_1_U81 ( .A(pe_1_4_1_n19), .B(pe_1_4_1_n16), .S(n49), .Z(
        int_data_y_4__1__3_) );
  MUX2_X1 pe_1_4_1_U80 ( .A(pe_1_4_1_n18), .B(pe_1_4_1_n17), .S(pe_1_4_1_n62), 
        .Z(pe_1_4_1_n19) );
  MUX2_X1 pe_1_4_1_U79 ( .A(pe_1_4_1_int_q_reg_v[23]), .B(
        pe_1_4_1_int_q_reg_v[19]), .S(pe_1_4_1_n55), .Z(pe_1_4_1_n18) );
  MUX2_X1 pe_1_4_1_U78 ( .A(pe_1_4_1_int_q_reg_v[15]), .B(
        pe_1_4_1_int_q_reg_v[11]), .S(pe_1_4_1_n55), .Z(pe_1_4_1_n17) );
  MUX2_X1 pe_1_4_1_U77 ( .A(pe_1_4_1_int_q_reg_v[7]), .B(
        pe_1_4_1_int_q_reg_v[3]), .S(pe_1_4_1_n55), .Z(pe_1_4_1_n16) );
  MUX2_X1 pe_1_4_1_U76 ( .A(pe_1_4_1_n15), .B(pe_1_4_1_n12), .S(n49), .Z(
        int_data_y_4__1__2_) );
  MUX2_X1 pe_1_4_1_U75 ( .A(pe_1_4_1_n14), .B(pe_1_4_1_n13), .S(pe_1_4_1_n62), 
        .Z(pe_1_4_1_n15) );
  MUX2_X1 pe_1_4_1_U74 ( .A(pe_1_4_1_int_q_reg_v[22]), .B(
        pe_1_4_1_int_q_reg_v[18]), .S(pe_1_4_1_n55), .Z(pe_1_4_1_n14) );
  MUX2_X1 pe_1_4_1_U73 ( .A(pe_1_4_1_int_q_reg_v[14]), .B(
        pe_1_4_1_int_q_reg_v[10]), .S(pe_1_4_1_n55), .Z(pe_1_4_1_n13) );
  MUX2_X1 pe_1_4_1_U72 ( .A(pe_1_4_1_int_q_reg_v[6]), .B(
        pe_1_4_1_int_q_reg_v[2]), .S(pe_1_4_1_n55), .Z(pe_1_4_1_n12) );
  MUX2_X1 pe_1_4_1_U71 ( .A(pe_1_4_1_n11), .B(pe_1_4_1_n8), .S(n49), .Z(
        int_data_y_4__1__1_) );
  MUX2_X1 pe_1_4_1_U70 ( .A(pe_1_4_1_n10), .B(pe_1_4_1_n9), .S(pe_1_4_1_n62), 
        .Z(pe_1_4_1_n11) );
  MUX2_X1 pe_1_4_1_U69 ( .A(pe_1_4_1_int_q_reg_v[21]), .B(
        pe_1_4_1_int_q_reg_v[17]), .S(pe_1_4_1_n55), .Z(pe_1_4_1_n10) );
  MUX2_X1 pe_1_4_1_U68 ( .A(pe_1_4_1_int_q_reg_v[13]), .B(
        pe_1_4_1_int_q_reg_v[9]), .S(pe_1_4_1_n55), .Z(pe_1_4_1_n9) );
  MUX2_X1 pe_1_4_1_U67 ( .A(pe_1_4_1_int_q_reg_v[5]), .B(
        pe_1_4_1_int_q_reg_v[1]), .S(pe_1_4_1_n55), .Z(pe_1_4_1_n8) );
  MUX2_X1 pe_1_4_1_U66 ( .A(pe_1_4_1_n7), .B(pe_1_4_1_n4), .S(n49), .Z(
        int_data_y_4__1__0_) );
  MUX2_X1 pe_1_4_1_U65 ( .A(pe_1_4_1_n6), .B(pe_1_4_1_n5), .S(pe_1_4_1_n62), 
        .Z(pe_1_4_1_n7) );
  MUX2_X1 pe_1_4_1_U64 ( .A(pe_1_4_1_int_q_reg_v[20]), .B(
        pe_1_4_1_int_q_reg_v[16]), .S(pe_1_4_1_n55), .Z(pe_1_4_1_n6) );
  MUX2_X1 pe_1_4_1_U63 ( .A(pe_1_4_1_int_q_reg_v[12]), .B(
        pe_1_4_1_int_q_reg_v[8]), .S(pe_1_4_1_n55), .Z(pe_1_4_1_n5) );
  MUX2_X1 pe_1_4_1_U62 ( .A(pe_1_4_1_int_q_reg_v[4]), .B(
        pe_1_4_1_int_q_reg_v[0]), .S(pe_1_4_1_n55), .Z(pe_1_4_1_n4) );
  AOI222_X1 pe_1_4_1_U61 ( .A1(int_data_res_5__1__2_), .A2(pe_1_4_1_n64), .B1(
        pe_1_4_1_N80), .B2(pe_1_4_1_n27), .C1(pe_1_4_1_N72), .C2(pe_1_4_1_n28), 
        .ZN(pe_1_4_1_n33) );
  INV_X1 pe_1_4_1_U60 ( .A(pe_1_4_1_n33), .ZN(pe_1_4_1_n82) );
  AOI222_X1 pe_1_4_1_U59 ( .A1(int_data_res_5__1__6_), .A2(pe_1_4_1_n64), .B1(
        pe_1_4_1_N84), .B2(pe_1_4_1_n27), .C1(pe_1_4_1_N76), .C2(pe_1_4_1_n28), 
        .ZN(pe_1_4_1_n29) );
  INV_X1 pe_1_4_1_U58 ( .A(pe_1_4_1_n29), .ZN(pe_1_4_1_n78) );
  XNOR2_X1 pe_1_4_1_U57 ( .A(pe_1_4_1_n73), .B(int_data_res_4__1__0_), .ZN(
        pe_1_4_1_N70) );
  AOI222_X1 pe_1_4_1_U52 ( .A1(int_data_res_5__1__0_), .A2(pe_1_4_1_n64), .B1(
        pe_1_4_1_n1), .B2(pe_1_4_1_n27), .C1(pe_1_4_1_N70), .C2(pe_1_4_1_n28), 
        .ZN(pe_1_4_1_n35) );
  INV_X1 pe_1_4_1_U51 ( .A(pe_1_4_1_n35), .ZN(pe_1_4_1_n84) );
  AOI222_X1 pe_1_4_1_U50 ( .A1(int_data_res_5__1__1_), .A2(pe_1_4_1_n64), .B1(
        pe_1_4_1_N79), .B2(pe_1_4_1_n27), .C1(pe_1_4_1_N71), .C2(pe_1_4_1_n28), 
        .ZN(pe_1_4_1_n34) );
  INV_X1 pe_1_4_1_U49 ( .A(pe_1_4_1_n34), .ZN(pe_1_4_1_n83) );
  AOI222_X1 pe_1_4_1_U48 ( .A1(int_data_res_5__1__3_), .A2(pe_1_4_1_n64), .B1(
        pe_1_4_1_N81), .B2(pe_1_4_1_n27), .C1(pe_1_4_1_N73), .C2(pe_1_4_1_n28), 
        .ZN(pe_1_4_1_n32) );
  INV_X1 pe_1_4_1_U47 ( .A(pe_1_4_1_n32), .ZN(pe_1_4_1_n81) );
  AOI222_X1 pe_1_4_1_U46 ( .A1(int_data_res_5__1__4_), .A2(pe_1_4_1_n64), .B1(
        pe_1_4_1_N82), .B2(pe_1_4_1_n27), .C1(pe_1_4_1_N74), .C2(pe_1_4_1_n28), 
        .ZN(pe_1_4_1_n31) );
  INV_X1 pe_1_4_1_U45 ( .A(pe_1_4_1_n31), .ZN(pe_1_4_1_n80) );
  AOI222_X1 pe_1_4_1_U44 ( .A1(int_data_res_5__1__5_), .A2(pe_1_4_1_n64), .B1(
        pe_1_4_1_N83), .B2(pe_1_4_1_n27), .C1(pe_1_4_1_N75), .C2(pe_1_4_1_n28), 
        .ZN(pe_1_4_1_n30) );
  INV_X1 pe_1_4_1_U43 ( .A(pe_1_4_1_n30), .ZN(pe_1_4_1_n79) );
  NAND2_X1 pe_1_4_1_U42 ( .A1(pe_1_4_1_int_data_0_), .A2(pe_1_4_1_n3), .ZN(
        pe_1_4_1_sub_81_carry[1]) );
  INV_X1 pe_1_4_1_U41 ( .A(pe_1_4_1_int_data_1_), .ZN(pe_1_4_1_n74) );
  INV_X1 pe_1_4_1_U40 ( .A(pe_1_4_1_int_data_2_), .ZN(pe_1_4_1_n75) );
  AND2_X1 pe_1_4_1_U39 ( .A1(pe_1_4_1_int_data_0_), .A2(int_data_res_4__1__0_), 
        .ZN(pe_1_4_1_n2) );
  AOI222_X1 pe_1_4_1_U38 ( .A1(pe_1_4_1_n64), .A2(int_data_res_5__1__7_), .B1(
        pe_1_4_1_N85), .B2(pe_1_4_1_n27), .C1(pe_1_4_1_N77), .C2(pe_1_4_1_n28), 
        .ZN(pe_1_4_1_n26) );
  INV_X1 pe_1_4_1_U37 ( .A(pe_1_4_1_n26), .ZN(pe_1_4_1_n77) );
  NOR3_X1 pe_1_4_1_U36 ( .A1(pe_1_4_1_n59), .A2(pe_1_4_1_n65), .A3(int_ckg[30]), .ZN(pe_1_4_1_n36) );
  OR2_X1 pe_1_4_1_U35 ( .A1(pe_1_4_1_n36), .A2(pe_1_4_1_n64), .ZN(pe_1_4_1_N90) );
  INV_X1 pe_1_4_1_U34 ( .A(n39), .ZN(pe_1_4_1_n63) );
  AND2_X1 pe_1_4_1_U33 ( .A1(int_data_x_4__1__2_), .A2(pe_1_4_1_n58), .ZN(
        pe_1_4_1_int_data_2_) );
  AND2_X1 pe_1_4_1_U32 ( .A1(int_data_x_4__1__1_), .A2(pe_1_4_1_n58), .ZN(
        pe_1_4_1_int_data_1_) );
  AND2_X1 pe_1_4_1_U31 ( .A1(int_data_x_4__1__3_), .A2(pe_1_4_1_n58), .ZN(
        pe_1_4_1_int_data_3_) );
  BUF_X1 pe_1_4_1_U30 ( .A(n61), .Z(pe_1_4_1_n64) );
  INV_X1 pe_1_4_1_U29 ( .A(n33), .ZN(pe_1_4_1_n61) );
  AND2_X1 pe_1_4_1_U28 ( .A1(int_data_x_4__1__0_), .A2(pe_1_4_1_n58), .ZN(
        pe_1_4_1_int_data_0_) );
  NAND2_X1 pe_1_4_1_U27 ( .A1(pe_1_4_1_n44), .A2(pe_1_4_1_n61), .ZN(
        pe_1_4_1_n41) );
  AND3_X1 pe_1_4_1_U26 ( .A1(n75), .A2(pe_1_4_1_n63), .A3(n49), .ZN(
        pe_1_4_1_n44) );
  INV_X1 pe_1_4_1_U25 ( .A(pe_1_4_1_int_data_3_), .ZN(pe_1_4_1_n76) );
  NOR2_X1 pe_1_4_1_U24 ( .A1(pe_1_4_1_n70), .A2(n49), .ZN(pe_1_4_1_n43) );
  NOR2_X1 pe_1_4_1_U23 ( .A1(pe_1_4_1_n57), .A2(pe_1_4_1_n64), .ZN(
        pe_1_4_1_n28) );
  NOR2_X1 pe_1_4_1_U22 ( .A1(n19), .A2(pe_1_4_1_n64), .ZN(pe_1_4_1_n27) );
  INV_X1 pe_1_4_1_U21 ( .A(pe_1_4_1_int_data_0_), .ZN(pe_1_4_1_n73) );
  INV_X1 pe_1_4_1_U20 ( .A(pe_1_4_1_n41), .ZN(pe_1_4_1_n90) );
  INV_X1 pe_1_4_1_U19 ( .A(pe_1_4_1_n37), .ZN(pe_1_4_1_n88) );
  INV_X1 pe_1_4_1_U18 ( .A(pe_1_4_1_n38), .ZN(pe_1_4_1_n87) );
  INV_X1 pe_1_4_1_U17 ( .A(pe_1_4_1_n39), .ZN(pe_1_4_1_n86) );
  NOR2_X1 pe_1_4_1_U16 ( .A1(pe_1_4_1_n68), .A2(pe_1_4_1_n42), .ZN(
        pe_1_4_1_N59) );
  NOR2_X1 pe_1_4_1_U15 ( .A1(pe_1_4_1_n68), .A2(pe_1_4_1_n41), .ZN(
        pe_1_4_1_N60) );
  NOR2_X1 pe_1_4_1_U14 ( .A1(pe_1_4_1_n68), .A2(pe_1_4_1_n38), .ZN(
        pe_1_4_1_N63) );
  NOR2_X1 pe_1_4_1_U13 ( .A1(pe_1_4_1_n67), .A2(pe_1_4_1_n40), .ZN(
        pe_1_4_1_N61) );
  NOR2_X1 pe_1_4_1_U12 ( .A1(pe_1_4_1_n67), .A2(pe_1_4_1_n39), .ZN(
        pe_1_4_1_N62) );
  NOR2_X1 pe_1_4_1_U11 ( .A1(pe_1_4_1_n37), .A2(pe_1_4_1_n67), .ZN(
        pe_1_4_1_N64) );
  NAND2_X1 pe_1_4_1_U10 ( .A1(pe_1_4_1_n44), .A2(pe_1_4_1_n60), .ZN(
        pe_1_4_1_n42) );
  BUF_X1 pe_1_4_1_U9 ( .A(pe_1_4_1_n60), .Z(pe_1_4_1_n55) );
  INV_X1 pe_1_4_1_U8 ( .A(pe_1_4_1_n69), .ZN(pe_1_4_1_n65) );
  BUF_X1 pe_1_4_1_U7 ( .A(pe_1_4_1_n60), .Z(pe_1_4_1_n56) );
  INV_X1 pe_1_4_1_U6 ( .A(pe_1_4_1_n42), .ZN(pe_1_4_1_n89) );
  INV_X1 pe_1_4_1_U5 ( .A(pe_1_4_1_n40), .ZN(pe_1_4_1_n85) );
  INV_X2 pe_1_4_1_U4 ( .A(n83), .ZN(pe_1_4_1_n72) );
  XOR2_X1 pe_1_4_1_U3 ( .A(pe_1_4_1_int_data_0_), .B(int_data_res_4__1__0_), 
        .Z(pe_1_4_1_n1) );
  DFFR_X1 pe_1_4_1_int_q_acc_reg_0_ ( .D(pe_1_4_1_n84), .CK(pe_1_4_1_net4978), 
        .RN(pe_1_4_1_n72), .Q(int_data_res_4__1__0_), .QN(pe_1_4_1_n3) );
  DFFR_X1 pe_1_4_1_int_q_reg_v_reg_0__0_ ( .D(int_data_y_5__1__0_), .CK(
        pe_1_4_1_net4948), .RN(pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_v[20]) );
  DFFR_X1 pe_1_4_1_int_q_reg_v_reg_0__1_ ( .D(int_data_y_5__1__1_), .CK(
        pe_1_4_1_net4948), .RN(pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_v[21]) );
  DFFR_X1 pe_1_4_1_int_q_reg_v_reg_0__2_ ( .D(int_data_y_5__1__2_), .CK(
        pe_1_4_1_net4948), .RN(pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_v[22]) );
  DFFR_X1 pe_1_4_1_int_q_reg_v_reg_0__3_ ( .D(int_data_y_5__1__3_), .CK(
        pe_1_4_1_net4948), .RN(pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_v[23]) );
  DFFR_X1 pe_1_4_1_int_q_reg_v_reg_1__0_ ( .D(int_data_y_5__1__0_), .CK(
        pe_1_4_1_net4953), .RN(pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_v[16]) );
  DFFR_X1 pe_1_4_1_int_q_reg_v_reg_1__1_ ( .D(int_data_y_5__1__1_), .CK(
        pe_1_4_1_net4953), .RN(pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_v[17]) );
  DFFR_X1 pe_1_4_1_int_q_reg_v_reg_1__2_ ( .D(int_data_y_5__1__2_), .CK(
        pe_1_4_1_net4953), .RN(pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_v[18]) );
  DFFR_X1 pe_1_4_1_int_q_reg_v_reg_1__3_ ( .D(int_data_y_5__1__3_), .CK(
        pe_1_4_1_net4953), .RN(pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_v[19]) );
  DFFR_X1 pe_1_4_1_int_q_reg_v_reg_2__0_ ( .D(int_data_y_5__1__0_), .CK(
        pe_1_4_1_net4958), .RN(pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_v[12]) );
  DFFR_X1 pe_1_4_1_int_q_reg_v_reg_2__1_ ( .D(int_data_y_5__1__1_), .CK(
        pe_1_4_1_net4958), .RN(pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_v[13]) );
  DFFR_X1 pe_1_4_1_int_q_reg_v_reg_2__2_ ( .D(int_data_y_5__1__2_), .CK(
        pe_1_4_1_net4958), .RN(pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_v[14]) );
  DFFR_X1 pe_1_4_1_int_q_reg_v_reg_2__3_ ( .D(int_data_y_5__1__3_), .CK(
        pe_1_4_1_net4958), .RN(pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_v[15]) );
  DFFR_X1 pe_1_4_1_int_q_reg_v_reg_3__0_ ( .D(int_data_y_5__1__0_), .CK(
        pe_1_4_1_net4963), .RN(pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_v[8]) );
  DFFR_X1 pe_1_4_1_int_q_reg_v_reg_3__1_ ( .D(int_data_y_5__1__1_), .CK(
        pe_1_4_1_net4963), .RN(pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_v[9]) );
  DFFR_X1 pe_1_4_1_int_q_reg_v_reg_3__2_ ( .D(int_data_y_5__1__2_), .CK(
        pe_1_4_1_net4963), .RN(pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_v[10]) );
  DFFR_X1 pe_1_4_1_int_q_reg_v_reg_3__3_ ( .D(int_data_y_5__1__3_), .CK(
        pe_1_4_1_net4963), .RN(pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_v[11]) );
  DFFR_X1 pe_1_4_1_int_q_reg_v_reg_4__0_ ( .D(int_data_y_5__1__0_), .CK(
        pe_1_4_1_net4968), .RN(pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_v[4]) );
  DFFR_X1 pe_1_4_1_int_q_reg_v_reg_4__1_ ( .D(int_data_y_5__1__1_), .CK(
        pe_1_4_1_net4968), .RN(pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_v[5]) );
  DFFR_X1 pe_1_4_1_int_q_reg_v_reg_4__2_ ( .D(int_data_y_5__1__2_), .CK(
        pe_1_4_1_net4968), .RN(pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_v[6]) );
  DFFR_X1 pe_1_4_1_int_q_reg_v_reg_4__3_ ( .D(int_data_y_5__1__3_), .CK(
        pe_1_4_1_net4968), .RN(pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_v[7]) );
  DFFR_X1 pe_1_4_1_int_q_reg_v_reg_5__0_ ( .D(int_data_y_5__1__0_), .CK(
        pe_1_4_1_net4973), .RN(pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_v[0]) );
  DFFR_X1 pe_1_4_1_int_q_reg_v_reg_5__1_ ( .D(int_data_y_5__1__1_), .CK(
        pe_1_4_1_net4973), .RN(pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_v[1]) );
  DFFR_X1 pe_1_4_1_int_q_reg_v_reg_5__2_ ( .D(int_data_y_5__1__2_), .CK(
        pe_1_4_1_net4973), .RN(pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_v[2]) );
  DFFR_X1 pe_1_4_1_int_q_reg_v_reg_5__3_ ( .D(int_data_y_5__1__3_), .CK(
        pe_1_4_1_net4973), .RN(pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_4_1_int_q_reg_h_reg_0__0_ ( .D(int_data_x_4__2__0_), .SI(
        int_data_y_5__1__0_), .SE(pe_1_4_1_n65), .CK(pe_1_4_1_net4917), .RN(
        pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_4_1_int_q_reg_h_reg_0__1_ ( .D(int_data_x_4__2__1_), .SI(
        int_data_y_5__1__1_), .SE(pe_1_4_1_n65), .CK(pe_1_4_1_net4917), .RN(
        pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_4_1_int_q_reg_h_reg_0__2_ ( .D(int_data_x_4__2__2_), .SI(
        int_data_y_5__1__2_), .SE(pe_1_4_1_n65), .CK(pe_1_4_1_net4917), .RN(
        pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_4_1_int_q_reg_h_reg_0__3_ ( .D(int_data_x_4__2__3_), .SI(
        int_data_y_5__1__3_), .SE(pe_1_4_1_n65), .CK(pe_1_4_1_net4917), .RN(
        pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_4_1_int_q_reg_h_reg_1__0_ ( .D(int_data_x_4__2__0_), .SI(
        int_data_y_5__1__0_), .SE(pe_1_4_1_n65), .CK(pe_1_4_1_net4923), .RN(
        pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_4_1_int_q_reg_h_reg_1__1_ ( .D(int_data_x_4__2__1_), .SI(
        int_data_y_5__1__1_), .SE(pe_1_4_1_n65), .CK(pe_1_4_1_net4923), .RN(
        pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_4_1_int_q_reg_h_reg_1__2_ ( .D(int_data_x_4__2__2_), .SI(
        int_data_y_5__1__2_), .SE(pe_1_4_1_n65), .CK(pe_1_4_1_net4923), .RN(
        pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_4_1_int_q_reg_h_reg_1__3_ ( .D(int_data_x_4__2__3_), .SI(
        int_data_y_5__1__3_), .SE(pe_1_4_1_n65), .CK(pe_1_4_1_net4923), .RN(
        pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_4_1_int_q_reg_h_reg_2__0_ ( .D(int_data_x_4__2__0_), .SI(
        int_data_y_5__1__0_), .SE(pe_1_4_1_n65), .CK(pe_1_4_1_net4928), .RN(
        pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_4_1_int_q_reg_h_reg_2__1_ ( .D(int_data_x_4__2__1_), .SI(
        int_data_y_5__1__1_), .SE(pe_1_4_1_n65), .CK(pe_1_4_1_net4928), .RN(
        pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_4_1_int_q_reg_h_reg_2__2_ ( .D(int_data_x_4__2__2_), .SI(
        int_data_y_5__1__2_), .SE(pe_1_4_1_n65), .CK(pe_1_4_1_net4928), .RN(
        pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_4_1_int_q_reg_h_reg_2__3_ ( .D(int_data_x_4__2__3_), .SI(
        int_data_y_5__1__3_), .SE(pe_1_4_1_n65), .CK(pe_1_4_1_net4928), .RN(
        pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_4_1_int_q_reg_h_reg_3__0_ ( .D(int_data_x_4__2__0_), .SI(
        int_data_y_5__1__0_), .SE(pe_1_4_1_n65), .CK(pe_1_4_1_net4933), .RN(
        pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_4_1_int_q_reg_h_reg_3__1_ ( .D(int_data_x_4__2__1_), .SI(
        int_data_y_5__1__1_), .SE(pe_1_4_1_n65), .CK(pe_1_4_1_net4933), .RN(
        pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_4_1_int_q_reg_h_reg_3__2_ ( .D(int_data_x_4__2__2_), .SI(
        int_data_y_5__1__2_), .SE(pe_1_4_1_n65), .CK(pe_1_4_1_net4933), .RN(
        pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_4_1_int_q_reg_h_reg_3__3_ ( .D(int_data_x_4__2__3_), .SI(
        int_data_y_5__1__3_), .SE(pe_1_4_1_n65), .CK(pe_1_4_1_net4933), .RN(
        pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_4_1_int_q_reg_h_reg_4__0_ ( .D(int_data_x_4__2__0_), .SI(
        int_data_y_5__1__0_), .SE(pe_1_4_1_n66), .CK(pe_1_4_1_net4938), .RN(
        pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_4_1_int_q_reg_h_reg_4__1_ ( .D(int_data_x_4__2__1_), .SI(
        int_data_y_5__1__1_), .SE(pe_1_4_1_n66), .CK(pe_1_4_1_net4938), .RN(
        pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_4_1_int_q_reg_h_reg_4__2_ ( .D(int_data_x_4__2__2_), .SI(
        int_data_y_5__1__2_), .SE(pe_1_4_1_n66), .CK(pe_1_4_1_net4938), .RN(
        pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_4_1_int_q_reg_h_reg_4__3_ ( .D(int_data_x_4__2__3_), .SI(
        int_data_y_5__1__3_), .SE(pe_1_4_1_n66), .CK(pe_1_4_1_net4938), .RN(
        pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_4_1_int_q_reg_h_reg_5__0_ ( .D(int_data_x_4__2__0_), .SI(
        int_data_y_5__1__0_), .SE(pe_1_4_1_n66), .CK(pe_1_4_1_net4943), .RN(
        pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_4_1_int_q_reg_h_reg_5__1_ ( .D(int_data_x_4__2__1_), .SI(
        int_data_y_5__1__1_), .SE(pe_1_4_1_n66), .CK(pe_1_4_1_net4943), .RN(
        pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_4_1_int_q_reg_h_reg_5__2_ ( .D(int_data_x_4__2__2_), .SI(
        int_data_y_5__1__2_), .SE(pe_1_4_1_n66), .CK(pe_1_4_1_net4943), .RN(
        pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_4_1_int_q_reg_h_reg_5__3_ ( .D(int_data_x_4__2__3_), .SI(
        int_data_y_5__1__3_), .SE(pe_1_4_1_n66), .CK(pe_1_4_1_net4943), .RN(
        pe_1_4_1_n72), .Q(pe_1_4_1_int_q_reg_h[3]) );
  FA_X1 pe_1_4_1_sub_81_U2_7 ( .A(int_data_res_4__1__7_), .B(pe_1_4_1_n76), 
        .CI(pe_1_4_1_sub_81_carry[7]), .S(pe_1_4_1_N77) );
  FA_X1 pe_1_4_1_sub_81_U2_6 ( .A(int_data_res_4__1__6_), .B(pe_1_4_1_n76), 
        .CI(pe_1_4_1_sub_81_carry[6]), .CO(pe_1_4_1_sub_81_carry[7]), .S(
        pe_1_4_1_N76) );
  FA_X1 pe_1_4_1_sub_81_U2_5 ( .A(int_data_res_4__1__5_), .B(pe_1_4_1_n76), 
        .CI(pe_1_4_1_sub_81_carry[5]), .CO(pe_1_4_1_sub_81_carry[6]), .S(
        pe_1_4_1_N75) );
  FA_X1 pe_1_4_1_sub_81_U2_4 ( .A(int_data_res_4__1__4_), .B(pe_1_4_1_n76), 
        .CI(pe_1_4_1_sub_81_carry[4]), .CO(pe_1_4_1_sub_81_carry[5]), .S(
        pe_1_4_1_N74) );
  FA_X1 pe_1_4_1_sub_81_U2_3 ( .A(int_data_res_4__1__3_), .B(pe_1_4_1_n76), 
        .CI(pe_1_4_1_sub_81_carry[3]), .CO(pe_1_4_1_sub_81_carry[4]), .S(
        pe_1_4_1_N73) );
  FA_X1 pe_1_4_1_sub_81_U2_2 ( .A(int_data_res_4__1__2_), .B(pe_1_4_1_n75), 
        .CI(pe_1_4_1_sub_81_carry[2]), .CO(pe_1_4_1_sub_81_carry[3]), .S(
        pe_1_4_1_N72) );
  FA_X1 pe_1_4_1_sub_81_U2_1 ( .A(int_data_res_4__1__1_), .B(pe_1_4_1_n74), 
        .CI(pe_1_4_1_sub_81_carry[1]), .CO(pe_1_4_1_sub_81_carry[2]), .S(
        pe_1_4_1_N71) );
  FA_X1 pe_1_4_1_add_83_U1_7 ( .A(int_data_res_4__1__7_), .B(
        pe_1_4_1_int_data_3_), .CI(pe_1_4_1_add_83_carry[7]), .S(pe_1_4_1_N85)
         );
  FA_X1 pe_1_4_1_add_83_U1_6 ( .A(int_data_res_4__1__6_), .B(
        pe_1_4_1_int_data_3_), .CI(pe_1_4_1_add_83_carry[6]), .CO(
        pe_1_4_1_add_83_carry[7]), .S(pe_1_4_1_N84) );
  FA_X1 pe_1_4_1_add_83_U1_5 ( .A(int_data_res_4__1__5_), .B(
        pe_1_4_1_int_data_3_), .CI(pe_1_4_1_add_83_carry[5]), .CO(
        pe_1_4_1_add_83_carry[6]), .S(pe_1_4_1_N83) );
  FA_X1 pe_1_4_1_add_83_U1_4 ( .A(int_data_res_4__1__4_), .B(
        pe_1_4_1_int_data_3_), .CI(pe_1_4_1_add_83_carry[4]), .CO(
        pe_1_4_1_add_83_carry[5]), .S(pe_1_4_1_N82) );
  FA_X1 pe_1_4_1_add_83_U1_3 ( .A(int_data_res_4__1__3_), .B(
        pe_1_4_1_int_data_3_), .CI(pe_1_4_1_add_83_carry[3]), .CO(
        pe_1_4_1_add_83_carry[4]), .S(pe_1_4_1_N81) );
  FA_X1 pe_1_4_1_add_83_U1_2 ( .A(int_data_res_4__1__2_), .B(
        pe_1_4_1_int_data_2_), .CI(pe_1_4_1_add_83_carry[2]), .CO(
        pe_1_4_1_add_83_carry[3]), .S(pe_1_4_1_N80) );
  FA_X1 pe_1_4_1_add_83_U1_1 ( .A(int_data_res_4__1__1_), .B(
        pe_1_4_1_int_data_1_), .CI(pe_1_4_1_n2), .CO(pe_1_4_1_add_83_carry[2]), 
        .S(pe_1_4_1_N79) );
  NAND3_X1 pe_1_4_1_U56 ( .A1(pe_1_4_1_n60), .A2(pe_1_4_1_n43), .A3(
        pe_1_4_1_n62), .ZN(pe_1_4_1_n40) );
  NAND3_X1 pe_1_4_1_U55 ( .A1(pe_1_4_1_n43), .A2(pe_1_4_1_n61), .A3(
        pe_1_4_1_n62), .ZN(pe_1_4_1_n39) );
  NAND3_X1 pe_1_4_1_U54 ( .A1(pe_1_4_1_n43), .A2(pe_1_4_1_n63), .A3(
        pe_1_4_1_n60), .ZN(pe_1_4_1_n38) );
  NAND3_X1 pe_1_4_1_U53 ( .A1(pe_1_4_1_n61), .A2(pe_1_4_1_n63), .A3(
        pe_1_4_1_n43), .ZN(pe_1_4_1_n37) );
  DFFR_X1 pe_1_4_1_int_q_acc_reg_6_ ( .D(pe_1_4_1_n78), .CK(pe_1_4_1_net4978), 
        .RN(pe_1_4_1_n71), .Q(int_data_res_4__1__6_) );
  DFFR_X1 pe_1_4_1_int_q_acc_reg_5_ ( .D(pe_1_4_1_n79), .CK(pe_1_4_1_net4978), 
        .RN(pe_1_4_1_n71), .Q(int_data_res_4__1__5_) );
  DFFR_X1 pe_1_4_1_int_q_acc_reg_4_ ( .D(pe_1_4_1_n80), .CK(pe_1_4_1_net4978), 
        .RN(pe_1_4_1_n71), .Q(int_data_res_4__1__4_) );
  DFFR_X1 pe_1_4_1_int_q_acc_reg_3_ ( .D(pe_1_4_1_n81), .CK(pe_1_4_1_net4978), 
        .RN(pe_1_4_1_n71), .Q(int_data_res_4__1__3_) );
  DFFR_X1 pe_1_4_1_int_q_acc_reg_2_ ( .D(pe_1_4_1_n82), .CK(pe_1_4_1_net4978), 
        .RN(pe_1_4_1_n71), .Q(int_data_res_4__1__2_) );
  DFFR_X1 pe_1_4_1_int_q_acc_reg_1_ ( .D(pe_1_4_1_n83), .CK(pe_1_4_1_net4978), 
        .RN(pe_1_4_1_n71), .Q(int_data_res_4__1__1_) );
  DFFR_X1 pe_1_4_1_int_q_acc_reg_7_ ( .D(pe_1_4_1_n77), .CK(pe_1_4_1_net4978), 
        .RN(pe_1_4_1_n71), .Q(int_data_res_4__1__7_) );
  CLKGATETST_X1 pe_1_4_1_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_4_1_n88), .SE(1'b0), .GCK(pe_1_4_1_net4917) );
  CLKGATETST_X1 pe_1_4_1_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_4_1_n87), .SE(1'b0), .GCK(pe_1_4_1_net4923) );
  CLKGATETST_X1 pe_1_4_1_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_4_1_n86), .SE(1'b0), .GCK(pe_1_4_1_net4928) );
  CLKGATETST_X1 pe_1_4_1_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_4_1_n85), .SE(1'b0), .GCK(pe_1_4_1_net4933) );
  CLKGATETST_X1 pe_1_4_1_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_4_1_n90), .SE(1'b0), .GCK(pe_1_4_1_net4938) );
  CLKGATETST_X1 pe_1_4_1_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_4_1_n89), .SE(1'b0), .GCK(pe_1_4_1_net4943) );
  CLKGATETST_X1 pe_1_4_1_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_4_1_N64), .SE(1'b0), .GCK(pe_1_4_1_net4948) );
  CLKGATETST_X1 pe_1_4_1_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_4_1_N63), .SE(1'b0), .GCK(pe_1_4_1_net4953) );
  CLKGATETST_X1 pe_1_4_1_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_4_1_N62), .SE(1'b0), .GCK(pe_1_4_1_net4958) );
  CLKGATETST_X1 pe_1_4_1_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_4_1_N61), .SE(1'b0), .GCK(pe_1_4_1_net4963) );
  CLKGATETST_X1 pe_1_4_1_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_4_1_N60), .SE(1'b0), .GCK(pe_1_4_1_net4968) );
  CLKGATETST_X1 pe_1_4_1_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_4_1_N59), .SE(1'b0), .GCK(pe_1_4_1_net4973) );
  CLKGATETST_X1 pe_1_4_1_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_4_1_N90), .SE(1'b0), .GCK(pe_1_4_1_net4978) );
  CLKBUF_X1 pe_1_4_2_U112 ( .A(pe_1_4_2_n72), .Z(pe_1_4_2_n71) );
  INV_X1 pe_1_4_2_U111 ( .A(n75), .ZN(pe_1_4_2_n70) );
  INV_X1 pe_1_4_2_U110 ( .A(n67), .ZN(pe_1_4_2_n69) );
  INV_X1 pe_1_4_2_U109 ( .A(n67), .ZN(pe_1_4_2_n68) );
  INV_X1 pe_1_4_2_U108 ( .A(n67), .ZN(pe_1_4_2_n67) );
  INV_X1 pe_1_4_2_U107 ( .A(pe_1_4_2_n69), .ZN(pe_1_4_2_n66) );
  INV_X1 pe_1_4_2_U106 ( .A(pe_1_4_2_n63), .ZN(pe_1_4_2_n62) );
  INV_X1 pe_1_4_2_U105 ( .A(pe_1_4_2_n61), .ZN(pe_1_4_2_n60) );
  INV_X1 pe_1_4_2_U104 ( .A(n27), .ZN(pe_1_4_2_n59) );
  INV_X1 pe_1_4_2_U103 ( .A(pe_1_4_2_n59), .ZN(pe_1_4_2_n58) );
  INV_X1 pe_1_4_2_U102 ( .A(n19), .ZN(pe_1_4_2_n57) );
  MUX2_X1 pe_1_4_2_U101 ( .A(pe_1_4_2_n54), .B(pe_1_4_2_n51), .S(n49), .Z(
        int_data_x_4__2__3_) );
  MUX2_X1 pe_1_4_2_U100 ( .A(pe_1_4_2_n53), .B(pe_1_4_2_n52), .S(pe_1_4_2_n62), 
        .Z(pe_1_4_2_n54) );
  MUX2_X1 pe_1_4_2_U99 ( .A(pe_1_4_2_int_q_reg_h[23]), .B(
        pe_1_4_2_int_q_reg_h[19]), .S(pe_1_4_2_n56), .Z(pe_1_4_2_n53) );
  MUX2_X1 pe_1_4_2_U98 ( .A(pe_1_4_2_int_q_reg_h[15]), .B(
        pe_1_4_2_int_q_reg_h[11]), .S(pe_1_4_2_n56), .Z(pe_1_4_2_n52) );
  MUX2_X1 pe_1_4_2_U97 ( .A(pe_1_4_2_int_q_reg_h[7]), .B(
        pe_1_4_2_int_q_reg_h[3]), .S(pe_1_4_2_n56), .Z(pe_1_4_2_n51) );
  MUX2_X1 pe_1_4_2_U96 ( .A(pe_1_4_2_n50), .B(pe_1_4_2_n47), .S(n49), .Z(
        int_data_x_4__2__2_) );
  MUX2_X1 pe_1_4_2_U95 ( .A(pe_1_4_2_n49), .B(pe_1_4_2_n48), .S(pe_1_4_2_n62), 
        .Z(pe_1_4_2_n50) );
  MUX2_X1 pe_1_4_2_U94 ( .A(pe_1_4_2_int_q_reg_h[22]), .B(
        pe_1_4_2_int_q_reg_h[18]), .S(pe_1_4_2_n56), .Z(pe_1_4_2_n49) );
  MUX2_X1 pe_1_4_2_U93 ( .A(pe_1_4_2_int_q_reg_h[14]), .B(
        pe_1_4_2_int_q_reg_h[10]), .S(pe_1_4_2_n56), .Z(pe_1_4_2_n48) );
  MUX2_X1 pe_1_4_2_U92 ( .A(pe_1_4_2_int_q_reg_h[6]), .B(
        pe_1_4_2_int_q_reg_h[2]), .S(pe_1_4_2_n56), .Z(pe_1_4_2_n47) );
  MUX2_X1 pe_1_4_2_U91 ( .A(pe_1_4_2_n46), .B(pe_1_4_2_n24), .S(n49), .Z(
        int_data_x_4__2__1_) );
  MUX2_X1 pe_1_4_2_U90 ( .A(pe_1_4_2_n45), .B(pe_1_4_2_n25), .S(pe_1_4_2_n62), 
        .Z(pe_1_4_2_n46) );
  MUX2_X1 pe_1_4_2_U89 ( .A(pe_1_4_2_int_q_reg_h[21]), .B(
        pe_1_4_2_int_q_reg_h[17]), .S(pe_1_4_2_n56), .Z(pe_1_4_2_n45) );
  MUX2_X1 pe_1_4_2_U88 ( .A(pe_1_4_2_int_q_reg_h[13]), .B(
        pe_1_4_2_int_q_reg_h[9]), .S(pe_1_4_2_n56), .Z(pe_1_4_2_n25) );
  MUX2_X1 pe_1_4_2_U87 ( .A(pe_1_4_2_int_q_reg_h[5]), .B(
        pe_1_4_2_int_q_reg_h[1]), .S(pe_1_4_2_n56), .Z(pe_1_4_2_n24) );
  MUX2_X1 pe_1_4_2_U86 ( .A(pe_1_4_2_n23), .B(pe_1_4_2_n20), .S(n49), .Z(
        int_data_x_4__2__0_) );
  MUX2_X1 pe_1_4_2_U85 ( .A(pe_1_4_2_n22), .B(pe_1_4_2_n21), .S(pe_1_4_2_n62), 
        .Z(pe_1_4_2_n23) );
  MUX2_X1 pe_1_4_2_U84 ( .A(pe_1_4_2_int_q_reg_h[20]), .B(
        pe_1_4_2_int_q_reg_h[16]), .S(pe_1_4_2_n56), .Z(pe_1_4_2_n22) );
  MUX2_X1 pe_1_4_2_U83 ( .A(pe_1_4_2_int_q_reg_h[12]), .B(
        pe_1_4_2_int_q_reg_h[8]), .S(pe_1_4_2_n56), .Z(pe_1_4_2_n21) );
  MUX2_X1 pe_1_4_2_U82 ( .A(pe_1_4_2_int_q_reg_h[4]), .B(
        pe_1_4_2_int_q_reg_h[0]), .S(pe_1_4_2_n56), .Z(pe_1_4_2_n20) );
  MUX2_X1 pe_1_4_2_U81 ( .A(pe_1_4_2_n19), .B(pe_1_4_2_n16), .S(n49), .Z(
        int_data_y_4__2__3_) );
  MUX2_X1 pe_1_4_2_U80 ( .A(pe_1_4_2_n18), .B(pe_1_4_2_n17), .S(pe_1_4_2_n62), 
        .Z(pe_1_4_2_n19) );
  MUX2_X1 pe_1_4_2_U79 ( .A(pe_1_4_2_int_q_reg_v[23]), .B(
        pe_1_4_2_int_q_reg_v[19]), .S(pe_1_4_2_n55), .Z(pe_1_4_2_n18) );
  MUX2_X1 pe_1_4_2_U78 ( .A(pe_1_4_2_int_q_reg_v[15]), .B(
        pe_1_4_2_int_q_reg_v[11]), .S(pe_1_4_2_n55), .Z(pe_1_4_2_n17) );
  MUX2_X1 pe_1_4_2_U77 ( .A(pe_1_4_2_int_q_reg_v[7]), .B(
        pe_1_4_2_int_q_reg_v[3]), .S(pe_1_4_2_n55), .Z(pe_1_4_2_n16) );
  MUX2_X1 pe_1_4_2_U76 ( .A(pe_1_4_2_n15), .B(pe_1_4_2_n12), .S(n49), .Z(
        int_data_y_4__2__2_) );
  MUX2_X1 pe_1_4_2_U75 ( .A(pe_1_4_2_n14), .B(pe_1_4_2_n13), .S(pe_1_4_2_n62), 
        .Z(pe_1_4_2_n15) );
  MUX2_X1 pe_1_4_2_U74 ( .A(pe_1_4_2_int_q_reg_v[22]), .B(
        pe_1_4_2_int_q_reg_v[18]), .S(pe_1_4_2_n55), .Z(pe_1_4_2_n14) );
  MUX2_X1 pe_1_4_2_U73 ( .A(pe_1_4_2_int_q_reg_v[14]), .B(
        pe_1_4_2_int_q_reg_v[10]), .S(pe_1_4_2_n55), .Z(pe_1_4_2_n13) );
  MUX2_X1 pe_1_4_2_U72 ( .A(pe_1_4_2_int_q_reg_v[6]), .B(
        pe_1_4_2_int_q_reg_v[2]), .S(pe_1_4_2_n55), .Z(pe_1_4_2_n12) );
  MUX2_X1 pe_1_4_2_U71 ( .A(pe_1_4_2_n11), .B(pe_1_4_2_n8), .S(n49), .Z(
        int_data_y_4__2__1_) );
  MUX2_X1 pe_1_4_2_U70 ( .A(pe_1_4_2_n10), .B(pe_1_4_2_n9), .S(pe_1_4_2_n62), 
        .Z(pe_1_4_2_n11) );
  MUX2_X1 pe_1_4_2_U69 ( .A(pe_1_4_2_int_q_reg_v[21]), .B(
        pe_1_4_2_int_q_reg_v[17]), .S(pe_1_4_2_n55), .Z(pe_1_4_2_n10) );
  MUX2_X1 pe_1_4_2_U68 ( .A(pe_1_4_2_int_q_reg_v[13]), .B(
        pe_1_4_2_int_q_reg_v[9]), .S(pe_1_4_2_n55), .Z(pe_1_4_2_n9) );
  MUX2_X1 pe_1_4_2_U67 ( .A(pe_1_4_2_int_q_reg_v[5]), .B(
        pe_1_4_2_int_q_reg_v[1]), .S(pe_1_4_2_n55), .Z(pe_1_4_2_n8) );
  MUX2_X1 pe_1_4_2_U66 ( .A(pe_1_4_2_n7), .B(pe_1_4_2_n4), .S(n49), .Z(
        int_data_y_4__2__0_) );
  MUX2_X1 pe_1_4_2_U65 ( .A(pe_1_4_2_n6), .B(pe_1_4_2_n5), .S(pe_1_4_2_n62), 
        .Z(pe_1_4_2_n7) );
  MUX2_X1 pe_1_4_2_U64 ( .A(pe_1_4_2_int_q_reg_v[20]), .B(
        pe_1_4_2_int_q_reg_v[16]), .S(pe_1_4_2_n55), .Z(pe_1_4_2_n6) );
  MUX2_X1 pe_1_4_2_U63 ( .A(pe_1_4_2_int_q_reg_v[12]), .B(
        pe_1_4_2_int_q_reg_v[8]), .S(pe_1_4_2_n55), .Z(pe_1_4_2_n5) );
  MUX2_X1 pe_1_4_2_U62 ( .A(pe_1_4_2_int_q_reg_v[4]), .B(
        pe_1_4_2_int_q_reg_v[0]), .S(pe_1_4_2_n55), .Z(pe_1_4_2_n4) );
  AOI222_X1 pe_1_4_2_U61 ( .A1(int_data_res_5__2__2_), .A2(pe_1_4_2_n64), .B1(
        pe_1_4_2_N80), .B2(pe_1_4_2_n27), .C1(pe_1_4_2_N72), .C2(pe_1_4_2_n28), 
        .ZN(pe_1_4_2_n33) );
  INV_X1 pe_1_4_2_U60 ( .A(pe_1_4_2_n33), .ZN(pe_1_4_2_n82) );
  AOI222_X1 pe_1_4_2_U59 ( .A1(int_data_res_5__2__6_), .A2(pe_1_4_2_n64), .B1(
        pe_1_4_2_N84), .B2(pe_1_4_2_n27), .C1(pe_1_4_2_N76), .C2(pe_1_4_2_n28), 
        .ZN(pe_1_4_2_n29) );
  INV_X1 pe_1_4_2_U58 ( .A(pe_1_4_2_n29), .ZN(pe_1_4_2_n78) );
  XNOR2_X1 pe_1_4_2_U57 ( .A(pe_1_4_2_n73), .B(int_data_res_4__2__0_), .ZN(
        pe_1_4_2_N70) );
  AOI222_X1 pe_1_4_2_U52 ( .A1(int_data_res_5__2__0_), .A2(pe_1_4_2_n64), .B1(
        pe_1_4_2_n1), .B2(pe_1_4_2_n27), .C1(pe_1_4_2_N70), .C2(pe_1_4_2_n28), 
        .ZN(pe_1_4_2_n35) );
  INV_X1 pe_1_4_2_U51 ( .A(pe_1_4_2_n35), .ZN(pe_1_4_2_n84) );
  AOI222_X1 pe_1_4_2_U50 ( .A1(int_data_res_5__2__1_), .A2(pe_1_4_2_n64), .B1(
        pe_1_4_2_N79), .B2(pe_1_4_2_n27), .C1(pe_1_4_2_N71), .C2(pe_1_4_2_n28), 
        .ZN(pe_1_4_2_n34) );
  INV_X1 pe_1_4_2_U49 ( .A(pe_1_4_2_n34), .ZN(pe_1_4_2_n83) );
  AOI222_X1 pe_1_4_2_U48 ( .A1(int_data_res_5__2__3_), .A2(pe_1_4_2_n64), .B1(
        pe_1_4_2_N81), .B2(pe_1_4_2_n27), .C1(pe_1_4_2_N73), .C2(pe_1_4_2_n28), 
        .ZN(pe_1_4_2_n32) );
  INV_X1 pe_1_4_2_U47 ( .A(pe_1_4_2_n32), .ZN(pe_1_4_2_n81) );
  AOI222_X1 pe_1_4_2_U46 ( .A1(int_data_res_5__2__4_), .A2(pe_1_4_2_n64), .B1(
        pe_1_4_2_N82), .B2(pe_1_4_2_n27), .C1(pe_1_4_2_N74), .C2(pe_1_4_2_n28), 
        .ZN(pe_1_4_2_n31) );
  INV_X1 pe_1_4_2_U45 ( .A(pe_1_4_2_n31), .ZN(pe_1_4_2_n80) );
  AOI222_X1 pe_1_4_2_U44 ( .A1(int_data_res_5__2__5_), .A2(pe_1_4_2_n64), .B1(
        pe_1_4_2_N83), .B2(pe_1_4_2_n27), .C1(pe_1_4_2_N75), .C2(pe_1_4_2_n28), 
        .ZN(pe_1_4_2_n30) );
  INV_X1 pe_1_4_2_U43 ( .A(pe_1_4_2_n30), .ZN(pe_1_4_2_n79) );
  NAND2_X1 pe_1_4_2_U42 ( .A1(pe_1_4_2_int_data_0_), .A2(pe_1_4_2_n3), .ZN(
        pe_1_4_2_sub_81_carry[1]) );
  INV_X1 pe_1_4_2_U41 ( .A(pe_1_4_2_int_data_1_), .ZN(pe_1_4_2_n74) );
  INV_X1 pe_1_4_2_U40 ( .A(pe_1_4_2_int_data_2_), .ZN(pe_1_4_2_n75) );
  AND2_X1 pe_1_4_2_U39 ( .A1(pe_1_4_2_int_data_0_), .A2(int_data_res_4__2__0_), 
        .ZN(pe_1_4_2_n2) );
  AOI222_X1 pe_1_4_2_U38 ( .A1(pe_1_4_2_n64), .A2(int_data_res_5__2__7_), .B1(
        pe_1_4_2_N85), .B2(pe_1_4_2_n27), .C1(pe_1_4_2_N77), .C2(pe_1_4_2_n28), 
        .ZN(pe_1_4_2_n26) );
  INV_X1 pe_1_4_2_U37 ( .A(pe_1_4_2_n26), .ZN(pe_1_4_2_n77) );
  NOR3_X1 pe_1_4_2_U36 ( .A1(pe_1_4_2_n59), .A2(pe_1_4_2_n65), .A3(int_ckg[29]), .ZN(pe_1_4_2_n36) );
  OR2_X1 pe_1_4_2_U35 ( .A1(pe_1_4_2_n36), .A2(pe_1_4_2_n64), .ZN(pe_1_4_2_N90) );
  INV_X1 pe_1_4_2_U34 ( .A(n39), .ZN(pe_1_4_2_n63) );
  AND2_X1 pe_1_4_2_U33 ( .A1(int_data_x_4__2__2_), .A2(pe_1_4_2_n58), .ZN(
        pe_1_4_2_int_data_2_) );
  AND2_X1 pe_1_4_2_U32 ( .A1(int_data_x_4__2__1_), .A2(pe_1_4_2_n58), .ZN(
        pe_1_4_2_int_data_1_) );
  AND2_X1 pe_1_4_2_U31 ( .A1(int_data_x_4__2__3_), .A2(pe_1_4_2_n58), .ZN(
        pe_1_4_2_int_data_3_) );
  BUF_X1 pe_1_4_2_U30 ( .A(n61), .Z(pe_1_4_2_n64) );
  INV_X1 pe_1_4_2_U29 ( .A(n33), .ZN(pe_1_4_2_n61) );
  AND2_X1 pe_1_4_2_U28 ( .A1(int_data_x_4__2__0_), .A2(pe_1_4_2_n58), .ZN(
        pe_1_4_2_int_data_0_) );
  NAND2_X1 pe_1_4_2_U27 ( .A1(pe_1_4_2_n44), .A2(pe_1_4_2_n61), .ZN(
        pe_1_4_2_n41) );
  AND3_X1 pe_1_4_2_U26 ( .A1(n75), .A2(pe_1_4_2_n63), .A3(n49), .ZN(
        pe_1_4_2_n44) );
  INV_X1 pe_1_4_2_U25 ( .A(pe_1_4_2_int_data_3_), .ZN(pe_1_4_2_n76) );
  NOR2_X1 pe_1_4_2_U24 ( .A1(pe_1_4_2_n70), .A2(n49), .ZN(pe_1_4_2_n43) );
  NOR2_X1 pe_1_4_2_U23 ( .A1(pe_1_4_2_n57), .A2(pe_1_4_2_n64), .ZN(
        pe_1_4_2_n28) );
  NOR2_X1 pe_1_4_2_U22 ( .A1(n19), .A2(pe_1_4_2_n64), .ZN(pe_1_4_2_n27) );
  INV_X1 pe_1_4_2_U21 ( .A(pe_1_4_2_int_data_0_), .ZN(pe_1_4_2_n73) );
  INV_X1 pe_1_4_2_U20 ( .A(pe_1_4_2_n41), .ZN(pe_1_4_2_n90) );
  INV_X1 pe_1_4_2_U19 ( .A(pe_1_4_2_n37), .ZN(pe_1_4_2_n88) );
  INV_X1 pe_1_4_2_U18 ( .A(pe_1_4_2_n38), .ZN(pe_1_4_2_n87) );
  INV_X1 pe_1_4_2_U17 ( .A(pe_1_4_2_n39), .ZN(pe_1_4_2_n86) );
  NOR2_X1 pe_1_4_2_U16 ( .A1(pe_1_4_2_n68), .A2(pe_1_4_2_n42), .ZN(
        pe_1_4_2_N59) );
  NOR2_X1 pe_1_4_2_U15 ( .A1(pe_1_4_2_n68), .A2(pe_1_4_2_n41), .ZN(
        pe_1_4_2_N60) );
  NOR2_X1 pe_1_4_2_U14 ( .A1(pe_1_4_2_n68), .A2(pe_1_4_2_n38), .ZN(
        pe_1_4_2_N63) );
  NOR2_X1 pe_1_4_2_U13 ( .A1(pe_1_4_2_n67), .A2(pe_1_4_2_n40), .ZN(
        pe_1_4_2_N61) );
  NOR2_X1 pe_1_4_2_U12 ( .A1(pe_1_4_2_n67), .A2(pe_1_4_2_n39), .ZN(
        pe_1_4_2_N62) );
  NOR2_X1 pe_1_4_2_U11 ( .A1(pe_1_4_2_n37), .A2(pe_1_4_2_n67), .ZN(
        pe_1_4_2_N64) );
  NAND2_X1 pe_1_4_2_U10 ( .A1(pe_1_4_2_n44), .A2(pe_1_4_2_n60), .ZN(
        pe_1_4_2_n42) );
  BUF_X1 pe_1_4_2_U9 ( .A(pe_1_4_2_n60), .Z(pe_1_4_2_n55) );
  INV_X1 pe_1_4_2_U8 ( .A(pe_1_4_2_n69), .ZN(pe_1_4_2_n65) );
  BUF_X1 pe_1_4_2_U7 ( .A(pe_1_4_2_n60), .Z(pe_1_4_2_n56) );
  INV_X1 pe_1_4_2_U6 ( .A(pe_1_4_2_n42), .ZN(pe_1_4_2_n89) );
  INV_X1 pe_1_4_2_U5 ( .A(pe_1_4_2_n40), .ZN(pe_1_4_2_n85) );
  INV_X2 pe_1_4_2_U4 ( .A(n83), .ZN(pe_1_4_2_n72) );
  XOR2_X1 pe_1_4_2_U3 ( .A(pe_1_4_2_int_data_0_), .B(int_data_res_4__2__0_), 
        .Z(pe_1_4_2_n1) );
  DFFR_X1 pe_1_4_2_int_q_acc_reg_0_ ( .D(pe_1_4_2_n84), .CK(pe_1_4_2_net4900), 
        .RN(pe_1_4_2_n72), .Q(int_data_res_4__2__0_), .QN(pe_1_4_2_n3) );
  DFFR_X1 pe_1_4_2_int_q_reg_v_reg_0__0_ ( .D(int_data_y_5__2__0_), .CK(
        pe_1_4_2_net4870), .RN(pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_v[20]) );
  DFFR_X1 pe_1_4_2_int_q_reg_v_reg_0__1_ ( .D(int_data_y_5__2__1_), .CK(
        pe_1_4_2_net4870), .RN(pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_v[21]) );
  DFFR_X1 pe_1_4_2_int_q_reg_v_reg_0__2_ ( .D(int_data_y_5__2__2_), .CK(
        pe_1_4_2_net4870), .RN(pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_v[22]) );
  DFFR_X1 pe_1_4_2_int_q_reg_v_reg_0__3_ ( .D(int_data_y_5__2__3_), .CK(
        pe_1_4_2_net4870), .RN(pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_v[23]) );
  DFFR_X1 pe_1_4_2_int_q_reg_v_reg_1__0_ ( .D(int_data_y_5__2__0_), .CK(
        pe_1_4_2_net4875), .RN(pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_v[16]) );
  DFFR_X1 pe_1_4_2_int_q_reg_v_reg_1__1_ ( .D(int_data_y_5__2__1_), .CK(
        pe_1_4_2_net4875), .RN(pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_v[17]) );
  DFFR_X1 pe_1_4_2_int_q_reg_v_reg_1__2_ ( .D(int_data_y_5__2__2_), .CK(
        pe_1_4_2_net4875), .RN(pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_v[18]) );
  DFFR_X1 pe_1_4_2_int_q_reg_v_reg_1__3_ ( .D(int_data_y_5__2__3_), .CK(
        pe_1_4_2_net4875), .RN(pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_v[19]) );
  DFFR_X1 pe_1_4_2_int_q_reg_v_reg_2__0_ ( .D(int_data_y_5__2__0_), .CK(
        pe_1_4_2_net4880), .RN(pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_v[12]) );
  DFFR_X1 pe_1_4_2_int_q_reg_v_reg_2__1_ ( .D(int_data_y_5__2__1_), .CK(
        pe_1_4_2_net4880), .RN(pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_v[13]) );
  DFFR_X1 pe_1_4_2_int_q_reg_v_reg_2__2_ ( .D(int_data_y_5__2__2_), .CK(
        pe_1_4_2_net4880), .RN(pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_v[14]) );
  DFFR_X1 pe_1_4_2_int_q_reg_v_reg_2__3_ ( .D(int_data_y_5__2__3_), .CK(
        pe_1_4_2_net4880), .RN(pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_v[15]) );
  DFFR_X1 pe_1_4_2_int_q_reg_v_reg_3__0_ ( .D(int_data_y_5__2__0_), .CK(
        pe_1_4_2_net4885), .RN(pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_v[8]) );
  DFFR_X1 pe_1_4_2_int_q_reg_v_reg_3__1_ ( .D(int_data_y_5__2__1_), .CK(
        pe_1_4_2_net4885), .RN(pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_v[9]) );
  DFFR_X1 pe_1_4_2_int_q_reg_v_reg_3__2_ ( .D(int_data_y_5__2__2_), .CK(
        pe_1_4_2_net4885), .RN(pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_v[10]) );
  DFFR_X1 pe_1_4_2_int_q_reg_v_reg_3__3_ ( .D(int_data_y_5__2__3_), .CK(
        pe_1_4_2_net4885), .RN(pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_v[11]) );
  DFFR_X1 pe_1_4_2_int_q_reg_v_reg_4__0_ ( .D(int_data_y_5__2__0_), .CK(
        pe_1_4_2_net4890), .RN(pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_v[4]) );
  DFFR_X1 pe_1_4_2_int_q_reg_v_reg_4__1_ ( .D(int_data_y_5__2__1_), .CK(
        pe_1_4_2_net4890), .RN(pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_v[5]) );
  DFFR_X1 pe_1_4_2_int_q_reg_v_reg_4__2_ ( .D(int_data_y_5__2__2_), .CK(
        pe_1_4_2_net4890), .RN(pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_v[6]) );
  DFFR_X1 pe_1_4_2_int_q_reg_v_reg_4__3_ ( .D(int_data_y_5__2__3_), .CK(
        pe_1_4_2_net4890), .RN(pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_v[7]) );
  DFFR_X1 pe_1_4_2_int_q_reg_v_reg_5__0_ ( .D(int_data_y_5__2__0_), .CK(
        pe_1_4_2_net4895), .RN(pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_v[0]) );
  DFFR_X1 pe_1_4_2_int_q_reg_v_reg_5__1_ ( .D(int_data_y_5__2__1_), .CK(
        pe_1_4_2_net4895), .RN(pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_v[1]) );
  DFFR_X1 pe_1_4_2_int_q_reg_v_reg_5__2_ ( .D(int_data_y_5__2__2_), .CK(
        pe_1_4_2_net4895), .RN(pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_v[2]) );
  DFFR_X1 pe_1_4_2_int_q_reg_v_reg_5__3_ ( .D(int_data_y_5__2__3_), .CK(
        pe_1_4_2_net4895), .RN(pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_4_2_int_q_reg_h_reg_0__0_ ( .D(int_data_x_4__3__0_), .SI(
        int_data_y_5__2__0_), .SE(pe_1_4_2_n65), .CK(pe_1_4_2_net4839), .RN(
        pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_4_2_int_q_reg_h_reg_0__1_ ( .D(int_data_x_4__3__1_), .SI(
        int_data_y_5__2__1_), .SE(pe_1_4_2_n65), .CK(pe_1_4_2_net4839), .RN(
        pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_4_2_int_q_reg_h_reg_0__2_ ( .D(int_data_x_4__3__2_), .SI(
        int_data_y_5__2__2_), .SE(pe_1_4_2_n65), .CK(pe_1_4_2_net4839), .RN(
        pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_4_2_int_q_reg_h_reg_0__3_ ( .D(int_data_x_4__3__3_), .SI(
        int_data_y_5__2__3_), .SE(pe_1_4_2_n65), .CK(pe_1_4_2_net4839), .RN(
        pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_4_2_int_q_reg_h_reg_1__0_ ( .D(int_data_x_4__3__0_), .SI(
        int_data_y_5__2__0_), .SE(pe_1_4_2_n65), .CK(pe_1_4_2_net4845), .RN(
        pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_4_2_int_q_reg_h_reg_1__1_ ( .D(int_data_x_4__3__1_), .SI(
        int_data_y_5__2__1_), .SE(pe_1_4_2_n65), .CK(pe_1_4_2_net4845), .RN(
        pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_4_2_int_q_reg_h_reg_1__2_ ( .D(int_data_x_4__3__2_), .SI(
        int_data_y_5__2__2_), .SE(pe_1_4_2_n65), .CK(pe_1_4_2_net4845), .RN(
        pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_4_2_int_q_reg_h_reg_1__3_ ( .D(int_data_x_4__3__3_), .SI(
        int_data_y_5__2__3_), .SE(pe_1_4_2_n65), .CK(pe_1_4_2_net4845), .RN(
        pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_4_2_int_q_reg_h_reg_2__0_ ( .D(int_data_x_4__3__0_), .SI(
        int_data_y_5__2__0_), .SE(pe_1_4_2_n65), .CK(pe_1_4_2_net4850), .RN(
        pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_4_2_int_q_reg_h_reg_2__1_ ( .D(int_data_x_4__3__1_), .SI(
        int_data_y_5__2__1_), .SE(pe_1_4_2_n65), .CK(pe_1_4_2_net4850), .RN(
        pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_4_2_int_q_reg_h_reg_2__2_ ( .D(int_data_x_4__3__2_), .SI(
        int_data_y_5__2__2_), .SE(pe_1_4_2_n65), .CK(pe_1_4_2_net4850), .RN(
        pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_4_2_int_q_reg_h_reg_2__3_ ( .D(int_data_x_4__3__3_), .SI(
        int_data_y_5__2__3_), .SE(pe_1_4_2_n65), .CK(pe_1_4_2_net4850), .RN(
        pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_4_2_int_q_reg_h_reg_3__0_ ( .D(int_data_x_4__3__0_), .SI(
        int_data_y_5__2__0_), .SE(pe_1_4_2_n65), .CK(pe_1_4_2_net4855), .RN(
        pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_4_2_int_q_reg_h_reg_3__1_ ( .D(int_data_x_4__3__1_), .SI(
        int_data_y_5__2__1_), .SE(pe_1_4_2_n65), .CK(pe_1_4_2_net4855), .RN(
        pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_4_2_int_q_reg_h_reg_3__2_ ( .D(int_data_x_4__3__2_), .SI(
        int_data_y_5__2__2_), .SE(pe_1_4_2_n65), .CK(pe_1_4_2_net4855), .RN(
        pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_4_2_int_q_reg_h_reg_3__3_ ( .D(int_data_x_4__3__3_), .SI(
        int_data_y_5__2__3_), .SE(pe_1_4_2_n65), .CK(pe_1_4_2_net4855), .RN(
        pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_4_2_int_q_reg_h_reg_4__0_ ( .D(int_data_x_4__3__0_), .SI(
        int_data_y_5__2__0_), .SE(pe_1_4_2_n66), .CK(pe_1_4_2_net4860), .RN(
        pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_4_2_int_q_reg_h_reg_4__1_ ( .D(int_data_x_4__3__1_), .SI(
        int_data_y_5__2__1_), .SE(pe_1_4_2_n66), .CK(pe_1_4_2_net4860), .RN(
        pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_4_2_int_q_reg_h_reg_4__2_ ( .D(int_data_x_4__3__2_), .SI(
        int_data_y_5__2__2_), .SE(pe_1_4_2_n66), .CK(pe_1_4_2_net4860), .RN(
        pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_4_2_int_q_reg_h_reg_4__3_ ( .D(int_data_x_4__3__3_), .SI(
        int_data_y_5__2__3_), .SE(pe_1_4_2_n66), .CK(pe_1_4_2_net4860), .RN(
        pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_4_2_int_q_reg_h_reg_5__0_ ( .D(int_data_x_4__3__0_), .SI(
        int_data_y_5__2__0_), .SE(pe_1_4_2_n66), .CK(pe_1_4_2_net4865), .RN(
        pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_4_2_int_q_reg_h_reg_5__1_ ( .D(int_data_x_4__3__1_), .SI(
        int_data_y_5__2__1_), .SE(pe_1_4_2_n66), .CK(pe_1_4_2_net4865), .RN(
        pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_4_2_int_q_reg_h_reg_5__2_ ( .D(int_data_x_4__3__2_), .SI(
        int_data_y_5__2__2_), .SE(pe_1_4_2_n66), .CK(pe_1_4_2_net4865), .RN(
        pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_4_2_int_q_reg_h_reg_5__3_ ( .D(int_data_x_4__3__3_), .SI(
        int_data_y_5__2__3_), .SE(pe_1_4_2_n66), .CK(pe_1_4_2_net4865), .RN(
        pe_1_4_2_n72), .Q(pe_1_4_2_int_q_reg_h[3]) );
  FA_X1 pe_1_4_2_sub_81_U2_7 ( .A(int_data_res_4__2__7_), .B(pe_1_4_2_n76), 
        .CI(pe_1_4_2_sub_81_carry[7]), .S(pe_1_4_2_N77) );
  FA_X1 pe_1_4_2_sub_81_U2_6 ( .A(int_data_res_4__2__6_), .B(pe_1_4_2_n76), 
        .CI(pe_1_4_2_sub_81_carry[6]), .CO(pe_1_4_2_sub_81_carry[7]), .S(
        pe_1_4_2_N76) );
  FA_X1 pe_1_4_2_sub_81_U2_5 ( .A(int_data_res_4__2__5_), .B(pe_1_4_2_n76), 
        .CI(pe_1_4_2_sub_81_carry[5]), .CO(pe_1_4_2_sub_81_carry[6]), .S(
        pe_1_4_2_N75) );
  FA_X1 pe_1_4_2_sub_81_U2_4 ( .A(int_data_res_4__2__4_), .B(pe_1_4_2_n76), 
        .CI(pe_1_4_2_sub_81_carry[4]), .CO(pe_1_4_2_sub_81_carry[5]), .S(
        pe_1_4_2_N74) );
  FA_X1 pe_1_4_2_sub_81_U2_3 ( .A(int_data_res_4__2__3_), .B(pe_1_4_2_n76), 
        .CI(pe_1_4_2_sub_81_carry[3]), .CO(pe_1_4_2_sub_81_carry[4]), .S(
        pe_1_4_2_N73) );
  FA_X1 pe_1_4_2_sub_81_U2_2 ( .A(int_data_res_4__2__2_), .B(pe_1_4_2_n75), 
        .CI(pe_1_4_2_sub_81_carry[2]), .CO(pe_1_4_2_sub_81_carry[3]), .S(
        pe_1_4_2_N72) );
  FA_X1 pe_1_4_2_sub_81_U2_1 ( .A(int_data_res_4__2__1_), .B(pe_1_4_2_n74), 
        .CI(pe_1_4_2_sub_81_carry[1]), .CO(pe_1_4_2_sub_81_carry[2]), .S(
        pe_1_4_2_N71) );
  FA_X1 pe_1_4_2_add_83_U1_7 ( .A(int_data_res_4__2__7_), .B(
        pe_1_4_2_int_data_3_), .CI(pe_1_4_2_add_83_carry[7]), .S(pe_1_4_2_N85)
         );
  FA_X1 pe_1_4_2_add_83_U1_6 ( .A(int_data_res_4__2__6_), .B(
        pe_1_4_2_int_data_3_), .CI(pe_1_4_2_add_83_carry[6]), .CO(
        pe_1_4_2_add_83_carry[7]), .S(pe_1_4_2_N84) );
  FA_X1 pe_1_4_2_add_83_U1_5 ( .A(int_data_res_4__2__5_), .B(
        pe_1_4_2_int_data_3_), .CI(pe_1_4_2_add_83_carry[5]), .CO(
        pe_1_4_2_add_83_carry[6]), .S(pe_1_4_2_N83) );
  FA_X1 pe_1_4_2_add_83_U1_4 ( .A(int_data_res_4__2__4_), .B(
        pe_1_4_2_int_data_3_), .CI(pe_1_4_2_add_83_carry[4]), .CO(
        pe_1_4_2_add_83_carry[5]), .S(pe_1_4_2_N82) );
  FA_X1 pe_1_4_2_add_83_U1_3 ( .A(int_data_res_4__2__3_), .B(
        pe_1_4_2_int_data_3_), .CI(pe_1_4_2_add_83_carry[3]), .CO(
        pe_1_4_2_add_83_carry[4]), .S(pe_1_4_2_N81) );
  FA_X1 pe_1_4_2_add_83_U1_2 ( .A(int_data_res_4__2__2_), .B(
        pe_1_4_2_int_data_2_), .CI(pe_1_4_2_add_83_carry[2]), .CO(
        pe_1_4_2_add_83_carry[3]), .S(pe_1_4_2_N80) );
  FA_X1 pe_1_4_2_add_83_U1_1 ( .A(int_data_res_4__2__1_), .B(
        pe_1_4_2_int_data_1_), .CI(pe_1_4_2_n2), .CO(pe_1_4_2_add_83_carry[2]), 
        .S(pe_1_4_2_N79) );
  NAND3_X1 pe_1_4_2_U56 ( .A1(pe_1_4_2_n60), .A2(pe_1_4_2_n43), .A3(
        pe_1_4_2_n62), .ZN(pe_1_4_2_n40) );
  NAND3_X1 pe_1_4_2_U55 ( .A1(pe_1_4_2_n43), .A2(pe_1_4_2_n61), .A3(
        pe_1_4_2_n62), .ZN(pe_1_4_2_n39) );
  NAND3_X1 pe_1_4_2_U54 ( .A1(pe_1_4_2_n43), .A2(pe_1_4_2_n63), .A3(
        pe_1_4_2_n60), .ZN(pe_1_4_2_n38) );
  NAND3_X1 pe_1_4_2_U53 ( .A1(pe_1_4_2_n61), .A2(pe_1_4_2_n63), .A3(
        pe_1_4_2_n43), .ZN(pe_1_4_2_n37) );
  DFFR_X1 pe_1_4_2_int_q_acc_reg_6_ ( .D(pe_1_4_2_n78), .CK(pe_1_4_2_net4900), 
        .RN(pe_1_4_2_n71), .Q(int_data_res_4__2__6_) );
  DFFR_X1 pe_1_4_2_int_q_acc_reg_5_ ( .D(pe_1_4_2_n79), .CK(pe_1_4_2_net4900), 
        .RN(pe_1_4_2_n71), .Q(int_data_res_4__2__5_) );
  DFFR_X1 pe_1_4_2_int_q_acc_reg_4_ ( .D(pe_1_4_2_n80), .CK(pe_1_4_2_net4900), 
        .RN(pe_1_4_2_n71), .Q(int_data_res_4__2__4_) );
  DFFR_X1 pe_1_4_2_int_q_acc_reg_3_ ( .D(pe_1_4_2_n81), .CK(pe_1_4_2_net4900), 
        .RN(pe_1_4_2_n71), .Q(int_data_res_4__2__3_) );
  DFFR_X1 pe_1_4_2_int_q_acc_reg_2_ ( .D(pe_1_4_2_n82), .CK(pe_1_4_2_net4900), 
        .RN(pe_1_4_2_n71), .Q(int_data_res_4__2__2_) );
  DFFR_X1 pe_1_4_2_int_q_acc_reg_1_ ( .D(pe_1_4_2_n83), .CK(pe_1_4_2_net4900), 
        .RN(pe_1_4_2_n71), .Q(int_data_res_4__2__1_) );
  DFFR_X1 pe_1_4_2_int_q_acc_reg_7_ ( .D(pe_1_4_2_n77), .CK(pe_1_4_2_net4900), 
        .RN(pe_1_4_2_n71), .Q(int_data_res_4__2__7_) );
  CLKGATETST_X1 pe_1_4_2_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_4_2_n88), .SE(1'b0), .GCK(pe_1_4_2_net4839) );
  CLKGATETST_X1 pe_1_4_2_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_4_2_n87), .SE(1'b0), .GCK(pe_1_4_2_net4845) );
  CLKGATETST_X1 pe_1_4_2_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_4_2_n86), .SE(1'b0), .GCK(pe_1_4_2_net4850) );
  CLKGATETST_X1 pe_1_4_2_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_4_2_n85), .SE(1'b0), .GCK(pe_1_4_2_net4855) );
  CLKGATETST_X1 pe_1_4_2_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_4_2_n90), .SE(1'b0), .GCK(pe_1_4_2_net4860) );
  CLKGATETST_X1 pe_1_4_2_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_4_2_n89), .SE(1'b0), .GCK(pe_1_4_2_net4865) );
  CLKGATETST_X1 pe_1_4_2_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_4_2_N64), .SE(1'b0), .GCK(pe_1_4_2_net4870) );
  CLKGATETST_X1 pe_1_4_2_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_4_2_N63), .SE(1'b0), .GCK(pe_1_4_2_net4875) );
  CLKGATETST_X1 pe_1_4_2_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_4_2_N62), .SE(1'b0), .GCK(pe_1_4_2_net4880) );
  CLKGATETST_X1 pe_1_4_2_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_4_2_N61), .SE(1'b0), .GCK(pe_1_4_2_net4885) );
  CLKGATETST_X1 pe_1_4_2_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_4_2_N60), .SE(1'b0), .GCK(pe_1_4_2_net4890) );
  CLKGATETST_X1 pe_1_4_2_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_4_2_N59), .SE(1'b0), .GCK(pe_1_4_2_net4895) );
  CLKGATETST_X1 pe_1_4_2_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_4_2_N90), .SE(1'b0), .GCK(pe_1_4_2_net4900) );
  CLKBUF_X1 pe_1_4_3_U112 ( .A(pe_1_4_3_n72), .Z(pe_1_4_3_n71) );
  INV_X1 pe_1_4_3_U111 ( .A(n75), .ZN(pe_1_4_3_n70) );
  INV_X1 pe_1_4_3_U110 ( .A(n67), .ZN(pe_1_4_3_n69) );
  INV_X1 pe_1_4_3_U109 ( .A(n67), .ZN(pe_1_4_3_n68) );
  INV_X1 pe_1_4_3_U108 ( .A(n67), .ZN(pe_1_4_3_n67) );
  INV_X1 pe_1_4_3_U107 ( .A(pe_1_4_3_n69), .ZN(pe_1_4_3_n66) );
  INV_X1 pe_1_4_3_U106 ( .A(pe_1_4_3_n63), .ZN(pe_1_4_3_n62) );
  INV_X1 pe_1_4_3_U105 ( .A(pe_1_4_3_n61), .ZN(pe_1_4_3_n60) );
  INV_X1 pe_1_4_3_U104 ( .A(n27), .ZN(pe_1_4_3_n59) );
  INV_X1 pe_1_4_3_U103 ( .A(pe_1_4_3_n59), .ZN(pe_1_4_3_n58) );
  INV_X1 pe_1_4_3_U102 ( .A(n19), .ZN(pe_1_4_3_n57) );
  MUX2_X1 pe_1_4_3_U101 ( .A(pe_1_4_3_n54), .B(pe_1_4_3_n51), .S(n50), .Z(
        int_data_x_4__3__3_) );
  MUX2_X1 pe_1_4_3_U100 ( .A(pe_1_4_3_n53), .B(pe_1_4_3_n52), .S(pe_1_4_3_n62), 
        .Z(pe_1_4_3_n54) );
  MUX2_X1 pe_1_4_3_U99 ( .A(pe_1_4_3_int_q_reg_h[23]), .B(
        pe_1_4_3_int_q_reg_h[19]), .S(pe_1_4_3_n56), .Z(pe_1_4_3_n53) );
  MUX2_X1 pe_1_4_3_U98 ( .A(pe_1_4_3_int_q_reg_h[15]), .B(
        pe_1_4_3_int_q_reg_h[11]), .S(pe_1_4_3_n56), .Z(pe_1_4_3_n52) );
  MUX2_X1 pe_1_4_3_U97 ( .A(pe_1_4_3_int_q_reg_h[7]), .B(
        pe_1_4_3_int_q_reg_h[3]), .S(pe_1_4_3_n56), .Z(pe_1_4_3_n51) );
  MUX2_X1 pe_1_4_3_U96 ( .A(pe_1_4_3_n50), .B(pe_1_4_3_n47), .S(n50), .Z(
        int_data_x_4__3__2_) );
  MUX2_X1 pe_1_4_3_U95 ( .A(pe_1_4_3_n49), .B(pe_1_4_3_n48), .S(pe_1_4_3_n62), 
        .Z(pe_1_4_3_n50) );
  MUX2_X1 pe_1_4_3_U94 ( .A(pe_1_4_3_int_q_reg_h[22]), .B(
        pe_1_4_3_int_q_reg_h[18]), .S(pe_1_4_3_n56), .Z(pe_1_4_3_n49) );
  MUX2_X1 pe_1_4_3_U93 ( .A(pe_1_4_3_int_q_reg_h[14]), .B(
        pe_1_4_3_int_q_reg_h[10]), .S(pe_1_4_3_n56), .Z(pe_1_4_3_n48) );
  MUX2_X1 pe_1_4_3_U92 ( .A(pe_1_4_3_int_q_reg_h[6]), .B(
        pe_1_4_3_int_q_reg_h[2]), .S(pe_1_4_3_n56), .Z(pe_1_4_3_n47) );
  MUX2_X1 pe_1_4_3_U91 ( .A(pe_1_4_3_n46), .B(pe_1_4_3_n24), .S(n50), .Z(
        int_data_x_4__3__1_) );
  MUX2_X1 pe_1_4_3_U90 ( .A(pe_1_4_3_n45), .B(pe_1_4_3_n25), .S(pe_1_4_3_n62), 
        .Z(pe_1_4_3_n46) );
  MUX2_X1 pe_1_4_3_U89 ( .A(pe_1_4_3_int_q_reg_h[21]), .B(
        pe_1_4_3_int_q_reg_h[17]), .S(pe_1_4_3_n56), .Z(pe_1_4_3_n45) );
  MUX2_X1 pe_1_4_3_U88 ( .A(pe_1_4_3_int_q_reg_h[13]), .B(
        pe_1_4_3_int_q_reg_h[9]), .S(pe_1_4_3_n56), .Z(pe_1_4_3_n25) );
  MUX2_X1 pe_1_4_3_U87 ( .A(pe_1_4_3_int_q_reg_h[5]), .B(
        pe_1_4_3_int_q_reg_h[1]), .S(pe_1_4_3_n56), .Z(pe_1_4_3_n24) );
  MUX2_X1 pe_1_4_3_U86 ( .A(pe_1_4_3_n23), .B(pe_1_4_3_n20), .S(n50), .Z(
        int_data_x_4__3__0_) );
  MUX2_X1 pe_1_4_3_U85 ( .A(pe_1_4_3_n22), .B(pe_1_4_3_n21), .S(pe_1_4_3_n62), 
        .Z(pe_1_4_3_n23) );
  MUX2_X1 pe_1_4_3_U84 ( .A(pe_1_4_3_int_q_reg_h[20]), .B(
        pe_1_4_3_int_q_reg_h[16]), .S(pe_1_4_3_n56), .Z(pe_1_4_3_n22) );
  MUX2_X1 pe_1_4_3_U83 ( .A(pe_1_4_3_int_q_reg_h[12]), .B(
        pe_1_4_3_int_q_reg_h[8]), .S(pe_1_4_3_n56), .Z(pe_1_4_3_n21) );
  MUX2_X1 pe_1_4_3_U82 ( .A(pe_1_4_3_int_q_reg_h[4]), .B(
        pe_1_4_3_int_q_reg_h[0]), .S(pe_1_4_3_n56), .Z(pe_1_4_3_n20) );
  MUX2_X1 pe_1_4_3_U81 ( .A(pe_1_4_3_n19), .B(pe_1_4_3_n16), .S(n50), .Z(
        int_data_y_4__3__3_) );
  MUX2_X1 pe_1_4_3_U80 ( .A(pe_1_4_3_n18), .B(pe_1_4_3_n17), .S(pe_1_4_3_n62), 
        .Z(pe_1_4_3_n19) );
  MUX2_X1 pe_1_4_3_U79 ( .A(pe_1_4_3_int_q_reg_v[23]), .B(
        pe_1_4_3_int_q_reg_v[19]), .S(pe_1_4_3_n55), .Z(pe_1_4_3_n18) );
  MUX2_X1 pe_1_4_3_U78 ( .A(pe_1_4_3_int_q_reg_v[15]), .B(
        pe_1_4_3_int_q_reg_v[11]), .S(pe_1_4_3_n55), .Z(pe_1_4_3_n17) );
  MUX2_X1 pe_1_4_3_U77 ( .A(pe_1_4_3_int_q_reg_v[7]), .B(
        pe_1_4_3_int_q_reg_v[3]), .S(pe_1_4_3_n55), .Z(pe_1_4_3_n16) );
  MUX2_X1 pe_1_4_3_U76 ( .A(pe_1_4_3_n15), .B(pe_1_4_3_n12), .S(n50), .Z(
        int_data_y_4__3__2_) );
  MUX2_X1 pe_1_4_3_U75 ( .A(pe_1_4_3_n14), .B(pe_1_4_3_n13), .S(pe_1_4_3_n62), 
        .Z(pe_1_4_3_n15) );
  MUX2_X1 pe_1_4_3_U74 ( .A(pe_1_4_3_int_q_reg_v[22]), .B(
        pe_1_4_3_int_q_reg_v[18]), .S(pe_1_4_3_n55), .Z(pe_1_4_3_n14) );
  MUX2_X1 pe_1_4_3_U73 ( .A(pe_1_4_3_int_q_reg_v[14]), .B(
        pe_1_4_3_int_q_reg_v[10]), .S(pe_1_4_3_n55), .Z(pe_1_4_3_n13) );
  MUX2_X1 pe_1_4_3_U72 ( .A(pe_1_4_3_int_q_reg_v[6]), .B(
        pe_1_4_3_int_q_reg_v[2]), .S(pe_1_4_3_n55), .Z(pe_1_4_3_n12) );
  MUX2_X1 pe_1_4_3_U71 ( .A(pe_1_4_3_n11), .B(pe_1_4_3_n8), .S(n50), .Z(
        int_data_y_4__3__1_) );
  MUX2_X1 pe_1_4_3_U70 ( .A(pe_1_4_3_n10), .B(pe_1_4_3_n9), .S(pe_1_4_3_n62), 
        .Z(pe_1_4_3_n11) );
  MUX2_X1 pe_1_4_3_U69 ( .A(pe_1_4_3_int_q_reg_v[21]), .B(
        pe_1_4_3_int_q_reg_v[17]), .S(pe_1_4_3_n55), .Z(pe_1_4_3_n10) );
  MUX2_X1 pe_1_4_3_U68 ( .A(pe_1_4_3_int_q_reg_v[13]), .B(
        pe_1_4_3_int_q_reg_v[9]), .S(pe_1_4_3_n55), .Z(pe_1_4_3_n9) );
  MUX2_X1 pe_1_4_3_U67 ( .A(pe_1_4_3_int_q_reg_v[5]), .B(
        pe_1_4_3_int_q_reg_v[1]), .S(pe_1_4_3_n55), .Z(pe_1_4_3_n8) );
  MUX2_X1 pe_1_4_3_U66 ( .A(pe_1_4_3_n7), .B(pe_1_4_3_n4), .S(n50), .Z(
        int_data_y_4__3__0_) );
  MUX2_X1 pe_1_4_3_U65 ( .A(pe_1_4_3_n6), .B(pe_1_4_3_n5), .S(pe_1_4_3_n62), 
        .Z(pe_1_4_3_n7) );
  MUX2_X1 pe_1_4_3_U64 ( .A(pe_1_4_3_int_q_reg_v[20]), .B(
        pe_1_4_3_int_q_reg_v[16]), .S(pe_1_4_3_n55), .Z(pe_1_4_3_n6) );
  MUX2_X1 pe_1_4_3_U63 ( .A(pe_1_4_3_int_q_reg_v[12]), .B(
        pe_1_4_3_int_q_reg_v[8]), .S(pe_1_4_3_n55), .Z(pe_1_4_3_n5) );
  MUX2_X1 pe_1_4_3_U62 ( .A(pe_1_4_3_int_q_reg_v[4]), .B(
        pe_1_4_3_int_q_reg_v[0]), .S(pe_1_4_3_n55), .Z(pe_1_4_3_n4) );
  AOI222_X1 pe_1_4_3_U61 ( .A1(int_data_res_5__3__2_), .A2(pe_1_4_3_n64), .B1(
        pe_1_4_3_N80), .B2(pe_1_4_3_n27), .C1(pe_1_4_3_N72), .C2(pe_1_4_3_n28), 
        .ZN(pe_1_4_3_n33) );
  INV_X1 pe_1_4_3_U60 ( .A(pe_1_4_3_n33), .ZN(pe_1_4_3_n82) );
  AOI222_X1 pe_1_4_3_U59 ( .A1(int_data_res_5__3__6_), .A2(pe_1_4_3_n64), .B1(
        pe_1_4_3_N84), .B2(pe_1_4_3_n27), .C1(pe_1_4_3_N76), .C2(pe_1_4_3_n28), 
        .ZN(pe_1_4_3_n29) );
  INV_X1 pe_1_4_3_U58 ( .A(pe_1_4_3_n29), .ZN(pe_1_4_3_n78) );
  XNOR2_X1 pe_1_4_3_U57 ( .A(pe_1_4_3_n73), .B(int_data_res_4__3__0_), .ZN(
        pe_1_4_3_N70) );
  AOI222_X1 pe_1_4_3_U52 ( .A1(int_data_res_5__3__0_), .A2(pe_1_4_3_n64), .B1(
        pe_1_4_3_n1), .B2(pe_1_4_3_n27), .C1(pe_1_4_3_N70), .C2(pe_1_4_3_n28), 
        .ZN(pe_1_4_3_n35) );
  INV_X1 pe_1_4_3_U51 ( .A(pe_1_4_3_n35), .ZN(pe_1_4_3_n84) );
  AOI222_X1 pe_1_4_3_U50 ( .A1(int_data_res_5__3__1_), .A2(pe_1_4_3_n64), .B1(
        pe_1_4_3_N79), .B2(pe_1_4_3_n27), .C1(pe_1_4_3_N71), .C2(pe_1_4_3_n28), 
        .ZN(pe_1_4_3_n34) );
  INV_X1 pe_1_4_3_U49 ( .A(pe_1_4_3_n34), .ZN(pe_1_4_3_n83) );
  AOI222_X1 pe_1_4_3_U48 ( .A1(int_data_res_5__3__3_), .A2(pe_1_4_3_n64), .B1(
        pe_1_4_3_N81), .B2(pe_1_4_3_n27), .C1(pe_1_4_3_N73), .C2(pe_1_4_3_n28), 
        .ZN(pe_1_4_3_n32) );
  INV_X1 pe_1_4_3_U47 ( .A(pe_1_4_3_n32), .ZN(pe_1_4_3_n81) );
  AOI222_X1 pe_1_4_3_U46 ( .A1(int_data_res_5__3__4_), .A2(pe_1_4_3_n64), .B1(
        pe_1_4_3_N82), .B2(pe_1_4_3_n27), .C1(pe_1_4_3_N74), .C2(pe_1_4_3_n28), 
        .ZN(pe_1_4_3_n31) );
  INV_X1 pe_1_4_3_U45 ( .A(pe_1_4_3_n31), .ZN(pe_1_4_3_n80) );
  AOI222_X1 pe_1_4_3_U44 ( .A1(int_data_res_5__3__5_), .A2(pe_1_4_3_n64), .B1(
        pe_1_4_3_N83), .B2(pe_1_4_3_n27), .C1(pe_1_4_3_N75), .C2(pe_1_4_3_n28), 
        .ZN(pe_1_4_3_n30) );
  INV_X1 pe_1_4_3_U43 ( .A(pe_1_4_3_n30), .ZN(pe_1_4_3_n79) );
  NAND2_X1 pe_1_4_3_U42 ( .A1(pe_1_4_3_int_data_0_), .A2(pe_1_4_3_n3), .ZN(
        pe_1_4_3_sub_81_carry[1]) );
  INV_X1 pe_1_4_3_U41 ( .A(pe_1_4_3_int_data_1_), .ZN(pe_1_4_3_n74) );
  INV_X1 pe_1_4_3_U40 ( .A(pe_1_4_3_int_data_2_), .ZN(pe_1_4_3_n75) );
  AND2_X1 pe_1_4_3_U39 ( .A1(pe_1_4_3_int_data_0_), .A2(int_data_res_4__3__0_), 
        .ZN(pe_1_4_3_n2) );
  AOI222_X1 pe_1_4_3_U38 ( .A1(pe_1_4_3_n64), .A2(int_data_res_5__3__7_), .B1(
        pe_1_4_3_N85), .B2(pe_1_4_3_n27), .C1(pe_1_4_3_N77), .C2(pe_1_4_3_n28), 
        .ZN(pe_1_4_3_n26) );
  INV_X1 pe_1_4_3_U37 ( .A(pe_1_4_3_n26), .ZN(pe_1_4_3_n77) );
  NOR3_X1 pe_1_4_3_U36 ( .A1(pe_1_4_3_n59), .A2(pe_1_4_3_n65), .A3(int_ckg[28]), .ZN(pe_1_4_3_n36) );
  OR2_X1 pe_1_4_3_U35 ( .A1(pe_1_4_3_n36), .A2(pe_1_4_3_n64), .ZN(pe_1_4_3_N90) );
  INV_X1 pe_1_4_3_U34 ( .A(n39), .ZN(pe_1_4_3_n63) );
  AND2_X1 pe_1_4_3_U33 ( .A1(int_data_x_4__3__2_), .A2(pe_1_4_3_n58), .ZN(
        pe_1_4_3_int_data_2_) );
  AND2_X1 pe_1_4_3_U32 ( .A1(int_data_x_4__3__1_), .A2(pe_1_4_3_n58), .ZN(
        pe_1_4_3_int_data_1_) );
  AND2_X1 pe_1_4_3_U31 ( .A1(int_data_x_4__3__3_), .A2(pe_1_4_3_n58), .ZN(
        pe_1_4_3_int_data_3_) );
  BUF_X1 pe_1_4_3_U30 ( .A(n61), .Z(pe_1_4_3_n64) );
  INV_X1 pe_1_4_3_U29 ( .A(n33), .ZN(pe_1_4_3_n61) );
  AND2_X1 pe_1_4_3_U28 ( .A1(int_data_x_4__3__0_), .A2(pe_1_4_3_n58), .ZN(
        pe_1_4_3_int_data_0_) );
  NAND2_X1 pe_1_4_3_U27 ( .A1(pe_1_4_3_n44), .A2(pe_1_4_3_n61), .ZN(
        pe_1_4_3_n41) );
  AND3_X1 pe_1_4_3_U26 ( .A1(n75), .A2(pe_1_4_3_n63), .A3(n50), .ZN(
        pe_1_4_3_n44) );
  INV_X1 pe_1_4_3_U25 ( .A(pe_1_4_3_int_data_3_), .ZN(pe_1_4_3_n76) );
  NOR2_X1 pe_1_4_3_U24 ( .A1(pe_1_4_3_n70), .A2(n50), .ZN(pe_1_4_3_n43) );
  NOR2_X1 pe_1_4_3_U23 ( .A1(pe_1_4_3_n57), .A2(pe_1_4_3_n64), .ZN(
        pe_1_4_3_n28) );
  NOR2_X1 pe_1_4_3_U22 ( .A1(n19), .A2(pe_1_4_3_n64), .ZN(pe_1_4_3_n27) );
  INV_X1 pe_1_4_3_U21 ( .A(pe_1_4_3_int_data_0_), .ZN(pe_1_4_3_n73) );
  INV_X1 pe_1_4_3_U20 ( .A(pe_1_4_3_n41), .ZN(pe_1_4_3_n90) );
  INV_X1 pe_1_4_3_U19 ( .A(pe_1_4_3_n37), .ZN(pe_1_4_3_n88) );
  INV_X1 pe_1_4_3_U18 ( .A(pe_1_4_3_n38), .ZN(pe_1_4_3_n87) );
  INV_X1 pe_1_4_3_U17 ( .A(pe_1_4_3_n39), .ZN(pe_1_4_3_n86) );
  NOR2_X1 pe_1_4_3_U16 ( .A1(pe_1_4_3_n68), .A2(pe_1_4_3_n42), .ZN(
        pe_1_4_3_N59) );
  NOR2_X1 pe_1_4_3_U15 ( .A1(pe_1_4_3_n68), .A2(pe_1_4_3_n41), .ZN(
        pe_1_4_3_N60) );
  NOR2_X1 pe_1_4_3_U14 ( .A1(pe_1_4_3_n68), .A2(pe_1_4_3_n38), .ZN(
        pe_1_4_3_N63) );
  NOR2_X1 pe_1_4_3_U13 ( .A1(pe_1_4_3_n67), .A2(pe_1_4_3_n40), .ZN(
        pe_1_4_3_N61) );
  NOR2_X1 pe_1_4_3_U12 ( .A1(pe_1_4_3_n67), .A2(pe_1_4_3_n39), .ZN(
        pe_1_4_3_N62) );
  NOR2_X1 pe_1_4_3_U11 ( .A1(pe_1_4_3_n37), .A2(pe_1_4_3_n67), .ZN(
        pe_1_4_3_N64) );
  NAND2_X1 pe_1_4_3_U10 ( .A1(pe_1_4_3_n44), .A2(pe_1_4_3_n60), .ZN(
        pe_1_4_3_n42) );
  BUF_X1 pe_1_4_3_U9 ( .A(pe_1_4_3_n60), .Z(pe_1_4_3_n55) );
  INV_X1 pe_1_4_3_U8 ( .A(pe_1_4_3_n69), .ZN(pe_1_4_3_n65) );
  BUF_X1 pe_1_4_3_U7 ( .A(pe_1_4_3_n60), .Z(pe_1_4_3_n56) );
  INV_X1 pe_1_4_3_U6 ( .A(pe_1_4_3_n42), .ZN(pe_1_4_3_n89) );
  INV_X1 pe_1_4_3_U5 ( .A(pe_1_4_3_n40), .ZN(pe_1_4_3_n85) );
  INV_X2 pe_1_4_3_U4 ( .A(n83), .ZN(pe_1_4_3_n72) );
  XOR2_X1 pe_1_4_3_U3 ( .A(pe_1_4_3_int_data_0_), .B(int_data_res_4__3__0_), 
        .Z(pe_1_4_3_n1) );
  DFFR_X1 pe_1_4_3_int_q_acc_reg_0_ ( .D(pe_1_4_3_n84), .CK(pe_1_4_3_net4822), 
        .RN(pe_1_4_3_n72), .Q(int_data_res_4__3__0_), .QN(pe_1_4_3_n3) );
  DFFR_X1 pe_1_4_3_int_q_reg_v_reg_0__0_ ( .D(int_data_y_5__3__0_), .CK(
        pe_1_4_3_net4792), .RN(pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_v[20]) );
  DFFR_X1 pe_1_4_3_int_q_reg_v_reg_0__1_ ( .D(int_data_y_5__3__1_), .CK(
        pe_1_4_3_net4792), .RN(pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_v[21]) );
  DFFR_X1 pe_1_4_3_int_q_reg_v_reg_0__2_ ( .D(int_data_y_5__3__2_), .CK(
        pe_1_4_3_net4792), .RN(pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_v[22]) );
  DFFR_X1 pe_1_4_3_int_q_reg_v_reg_0__3_ ( .D(int_data_y_5__3__3_), .CK(
        pe_1_4_3_net4792), .RN(pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_v[23]) );
  DFFR_X1 pe_1_4_3_int_q_reg_v_reg_1__0_ ( .D(int_data_y_5__3__0_), .CK(
        pe_1_4_3_net4797), .RN(pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_v[16]) );
  DFFR_X1 pe_1_4_3_int_q_reg_v_reg_1__1_ ( .D(int_data_y_5__3__1_), .CK(
        pe_1_4_3_net4797), .RN(pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_v[17]) );
  DFFR_X1 pe_1_4_3_int_q_reg_v_reg_1__2_ ( .D(int_data_y_5__3__2_), .CK(
        pe_1_4_3_net4797), .RN(pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_v[18]) );
  DFFR_X1 pe_1_4_3_int_q_reg_v_reg_1__3_ ( .D(int_data_y_5__3__3_), .CK(
        pe_1_4_3_net4797), .RN(pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_v[19]) );
  DFFR_X1 pe_1_4_3_int_q_reg_v_reg_2__0_ ( .D(int_data_y_5__3__0_), .CK(
        pe_1_4_3_net4802), .RN(pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_v[12]) );
  DFFR_X1 pe_1_4_3_int_q_reg_v_reg_2__1_ ( .D(int_data_y_5__3__1_), .CK(
        pe_1_4_3_net4802), .RN(pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_v[13]) );
  DFFR_X1 pe_1_4_3_int_q_reg_v_reg_2__2_ ( .D(int_data_y_5__3__2_), .CK(
        pe_1_4_3_net4802), .RN(pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_v[14]) );
  DFFR_X1 pe_1_4_3_int_q_reg_v_reg_2__3_ ( .D(int_data_y_5__3__3_), .CK(
        pe_1_4_3_net4802), .RN(pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_v[15]) );
  DFFR_X1 pe_1_4_3_int_q_reg_v_reg_3__0_ ( .D(int_data_y_5__3__0_), .CK(
        pe_1_4_3_net4807), .RN(pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_v[8]) );
  DFFR_X1 pe_1_4_3_int_q_reg_v_reg_3__1_ ( .D(int_data_y_5__3__1_), .CK(
        pe_1_4_3_net4807), .RN(pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_v[9]) );
  DFFR_X1 pe_1_4_3_int_q_reg_v_reg_3__2_ ( .D(int_data_y_5__3__2_), .CK(
        pe_1_4_3_net4807), .RN(pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_v[10]) );
  DFFR_X1 pe_1_4_3_int_q_reg_v_reg_3__3_ ( .D(int_data_y_5__3__3_), .CK(
        pe_1_4_3_net4807), .RN(pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_v[11]) );
  DFFR_X1 pe_1_4_3_int_q_reg_v_reg_4__0_ ( .D(int_data_y_5__3__0_), .CK(
        pe_1_4_3_net4812), .RN(pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_v[4]) );
  DFFR_X1 pe_1_4_3_int_q_reg_v_reg_4__1_ ( .D(int_data_y_5__3__1_), .CK(
        pe_1_4_3_net4812), .RN(pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_v[5]) );
  DFFR_X1 pe_1_4_3_int_q_reg_v_reg_4__2_ ( .D(int_data_y_5__3__2_), .CK(
        pe_1_4_3_net4812), .RN(pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_v[6]) );
  DFFR_X1 pe_1_4_3_int_q_reg_v_reg_4__3_ ( .D(int_data_y_5__3__3_), .CK(
        pe_1_4_3_net4812), .RN(pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_v[7]) );
  DFFR_X1 pe_1_4_3_int_q_reg_v_reg_5__0_ ( .D(int_data_y_5__3__0_), .CK(
        pe_1_4_3_net4817), .RN(pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_v[0]) );
  DFFR_X1 pe_1_4_3_int_q_reg_v_reg_5__1_ ( .D(int_data_y_5__3__1_), .CK(
        pe_1_4_3_net4817), .RN(pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_v[1]) );
  DFFR_X1 pe_1_4_3_int_q_reg_v_reg_5__2_ ( .D(int_data_y_5__3__2_), .CK(
        pe_1_4_3_net4817), .RN(pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_v[2]) );
  DFFR_X1 pe_1_4_3_int_q_reg_v_reg_5__3_ ( .D(int_data_y_5__3__3_), .CK(
        pe_1_4_3_net4817), .RN(pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_4_3_int_q_reg_h_reg_0__0_ ( .D(int_data_x_4__4__0_), .SI(
        int_data_y_5__3__0_), .SE(pe_1_4_3_n65), .CK(pe_1_4_3_net4761), .RN(
        pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_4_3_int_q_reg_h_reg_0__1_ ( .D(int_data_x_4__4__1_), .SI(
        int_data_y_5__3__1_), .SE(pe_1_4_3_n65), .CK(pe_1_4_3_net4761), .RN(
        pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_4_3_int_q_reg_h_reg_0__2_ ( .D(int_data_x_4__4__2_), .SI(
        int_data_y_5__3__2_), .SE(pe_1_4_3_n65), .CK(pe_1_4_3_net4761), .RN(
        pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_4_3_int_q_reg_h_reg_0__3_ ( .D(int_data_x_4__4__3_), .SI(
        int_data_y_5__3__3_), .SE(pe_1_4_3_n65), .CK(pe_1_4_3_net4761), .RN(
        pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_4_3_int_q_reg_h_reg_1__0_ ( .D(int_data_x_4__4__0_), .SI(
        int_data_y_5__3__0_), .SE(pe_1_4_3_n65), .CK(pe_1_4_3_net4767), .RN(
        pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_4_3_int_q_reg_h_reg_1__1_ ( .D(int_data_x_4__4__1_), .SI(
        int_data_y_5__3__1_), .SE(pe_1_4_3_n65), .CK(pe_1_4_3_net4767), .RN(
        pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_4_3_int_q_reg_h_reg_1__2_ ( .D(int_data_x_4__4__2_), .SI(
        int_data_y_5__3__2_), .SE(pe_1_4_3_n65), .CK(pe_1_4_3_net4767), .RN(
        pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_4_3_int_q_reg_h_reg_1__3_ ( .D(int_data_x_4__4__3_), .SI(
        int_data_y_5__3__3_), .SE(pe_1_4_3_n65), .CK(pe_1_4_3_net4767), .RN(
        pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_4_3_int_q_reg_h_reg_2__0_ ( .D(int_data_x_4__4__0_), .SI(
        int_data_y_5__3__0_), .SE(pe_1_4_3_n65), .CK(pe_1_4_3_net4772), .RN(
        pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_4_3_int_q_reg_h_reg_2__1_ ( .D(int_data_x_4__4__1_), .SI(
        int_data_y_5__3__1_), .SE(pe_1_4_3_n65), .CK(pe_1_4_3_net4772), .RN(
        pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_4_3_int_q_reg_h_reg_2__2_ ( .D(int_data_x_4__4__2_), .SI(
        int_data_y_5__3__2_), .SE(pe_1_4_3_n65), .CK(pe_1_4_3_net4772), .RN(
        pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_4_3_int_q_reg_h_reg_2__3_ ( .D(int_data_x_4__4__3_), .SI(
        int_data_y_5__3__3_), .SE(pe_1_4_3_n65), .CK(pe_1_4_3_net4772), .RN(
        pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_4_3_int_q_reg_h_reg_3__0_ ( .D(int_data_x_4__4__0_), .SI(
        int_data_y_5__3__0_), .SE(pe_1_4_3_n65), .CK(pe_1_4_3_net4777), .RN(
        pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_4_3_int_q_reg_h_reg_3__1_ ( .D(int_data_x_4__4__1_), .SI(
        int_data_y_5__3__1_), .SE(pe_1_4_3_n65), .CK(pe_1_4_3_net4777), .RN(
        pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_4_3_int_q_reg_h_reg_3__2_ ( .D(int_data_x_4__4__2_), .SI(
        int_data_y_5__3__2_), .SE(pe_1_4_3_n65), .CK(pe_1_4_3_net4777), .RN(
        pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_4_3_int_q_reg_h_reg_3__3_ ( .D(int_data_x_4__4__3_), .SI(
        int_data_y_5__3__3_), .SE(pe_1_4_3_n65), .CK(pe_1_4_3_net4777), .RN(
        pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_4_3_int_q_reg_h_reg_4__0_ ( .D(int_data_x_4__4__0_), .SI(
        int_data_y_5__3__0_), .SE(pe_1_4_3_n66), .CK(pe_1_4_3_net4782), .RN(
        pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_4_3_int_q_reg_h_reg_4__1_ ( .D(int_data_x_4__4__1_), .SI(
        int_data_y_5__3__1_), .SE(pe_1_4_3_n66), .CK(pe_1_4_3_net4782), .RN(
        pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_4_3_int_q_reg_h_reg_4__2_ ( .D(int_data_x_4__4__2_), .SI(
        int_data_y_5__3__2_), .SE(pe_1_4_3_n66), .CK(pe_1_4_3_net4782), .RN(
        pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_4_3_int_q_reg_h_reg_4__3_ ( .D(int_data_x_4__4__3_), .SI(
        int_data_y_5__3__3_), .SE(pe_1_4_3_n66), .CK(pe_1_4_3_net4782), .RN(
        pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_4_3_int_q_reg_h_reg_5__0_ ( .D(int_data_x_4__4__0_), .SI(
        int_data_y_5__3__0_), .SE(pe_1_4_3_n66), .CK(pe_1_4_3_net4787), .RN(
        pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_4_3_int_q_reg_h_reg_5__1_ ( .D(int_data_x_4__4__1_), .SI(
        int_data_y_5__3__1_), .SE(pe_1_4_3_n66), .CK(pe_1_4_3_net4787), .RN(
        pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_4_3_int_q_reg_h_reg_5__2_ ( .D(int_data_x_4__4__2_), .SI(
        int_data_y_5__3__2_), .SE(pe_1_4_3_n66), .CK(pe_1_4_3_net4787), .RN(
        pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_4_3_int_q_reg_h_reg_5__3_ ( .D(int_data_x_4__4__3_), .SI(
        int_data_y_5__3__3_), .SE(pe_1_4_3_n66), .CK(pe_1_4_3_net4787), .RN(
        pe_1_4_3_n72), .Q(pe_1_4_3_int_q_reg_h[3]) );
  FA_X1 pe_1_4_3_sub_81_U2_7 ( .A(int_data_res_4__3__7_), .B(pe_1_4_3_n76), 
        .CI(pe_1_4_3_sub_81_carry[7]), .S(pe_1_4_3_N77) );
  FA_X1 pe_1_4_3_sub_81_U2_6 ( .A(int_data_res_4__3__6_), .B(pe_1_4_3_n76), 
        .CI(pe_1_4_3_sub_81_carry[6]), .CO(pe_1_4_3_sub_81_carry[7]), .S(
        pe_1_4_3_N76) );
  FA_X1 pe_1_4_3_sub_81_U2_5 ( .A(int_data_res_4__3__5_), .B(pe_1_4_3_n76), 
        .CI(pe_1_4_3_sub_81_carry[5]), .CO(pe_1_4_3_sub_81_carry[6]), .S(
        pe_1_4_3_N75) );
  FA_X1 pe_1_4_3_sub_81_U2_4 ( .A(int_data_res_4__3__4_), .B(pe_1_4_3_n76), 
        .CI(pe_1_4_3_sub_81_carry[4]), .CO(pe_1_4_3_sub_81_carry[5]), .S(
        pe_1_4_3_N74) );
  FA_X1 pe_1_4_3_sub_81_U2_3 ( .A(int_data_res_4__3__3_), .B(pe_1_4_3_n76), 
        .CI(pe_1_4_3_sub_81_carry[3]), .CO(pe_1_4_3_sub_81_carry[4]), .S(
        pe_1_4_3_N73) );
  FA_X1 pe_1_4_3_sub_81_U2_2 ( .A(int_data_res_4__3__2_), .B(pe_1_4_3_n75), 
        .CI(pe_1_4_3_sub_81_carry[2]), .CO(pe_1_4_3_sub_81_carry[3]), .S(
        pe_1_4_3_N72) );
  FA_X1 pe_1_4_3_sub_81_U2_1 ( .A(int_data_res_4__3__1_), .B(pe_1_4_3_n74), 
        .CI(pe_1_4_3_sub_81_carry[1]), .CO(pe_1_4_3_sub_81_carry[2]), .S(
        pe_1_4_3_N71) );
  FA_X1 pe_1_4_3_add_83_U1_7 ( .A(int_data_res_4__3__7_), .B(
        pe_1_4_3_int_data_3_), .CI(pe_1_4_3_add_83_carry[7]), .S(pe_1_4_3_N85)
         );
  FA_X1 pe_1_4_3_add_83_U1_6 ( .A(int_data_res_4__3__6_), .B(
        pe_1_4_3_int_data_3_), .CI(pe_1_4_3_add_83_carry[6]), .CO(
        pe_1_4_3_add_83_carry[7]), .S(pe_1_4_3_N84) );
  FA_X1 pe_1_4_3_add_83_U1_5 ( .A(int_data_res_4__3__5_), .B(
        pe_1_4_3_int_data_3_), .CI(pe_1_4_3_add_83_carry[5]), .CO(
        pe_1_4_3_add_83_carry[6]), .S(pe_1_4_3_N83) );
  FA_X1 pe_1_4_3_add_83_U1_4 ( .A(int_data_res_4__3__4_), .B(
        pe_1_4_3_int_data_3_), .CI(pe_1_4_3_add_83_carry[4]), .CO(
        pe_1_4_3_add_83_carry[5]), .S(pe_1_4_3_N82) );
  FA_X1 pe_1_4_3_add_83_U1_3 ( .A(int_data_res_4__3__3_), .B(
        pe_1_4_3_int_data_3_), .CI(pe_1_4_3_add_83_carry[3]), .CO(
        pe_1_4_3_add_83_carry[4]), .S(pe_1_4_3_N81) );
  FA_X1 pe_1_4_3_add_83_U1_2 ( .A(int_data_res_4__3__2_), .B(
        pe_1_4_3_int_data_2_), .CI(pe_1_4_3_add_83_carry[2]), .CO(
        pe_1_4_3_add_83_carry[3]), .S(pe_1_4_3_N80) );
  FA_X1 pe_1_4_3_add_83_U1_1 ( .A(int_data_res_4__3__1_), .B(
        pe_1_4_3_int_data_1_), .CI(pe_1_4_3_n2), .CO(pe_1_4_3_add_83_carry[2]), 
        .S(pe_1_4_3_N79) );
  NAND3_X1 pe_1_4_3_U56 ( .A1(pe_1_4_3_n60), .A2(pe_1_4_3_n43), .A3(
        pe_1_4_3_n62), .ZN(pe_1_4_3_n40) );
  NAND3_X1 pe_1_4_3_U55 ( .A1(pe_1_4_3_n43), .A2(pe_1_4_3_n61), .A3(
        pe_1_4_3_n62), .ZN(pe_1_4_3_n39) );
  NAND3_X1 pe_1_4_3_U54 ( .A1(pe_1_4_3_n43), .A2(pe_1_4_3_n63), .A3(
        pe_1_4_3_n60), .ZN(pe_1_4_3_n38) );
  NAND3_X1 pe_1_4_3_U53 ( .A1(pe_1_4_3_n61), .A2(pe_1_4_3_n63), .A3(
        pe_1_4_3_n43), .ZN(pe_1_4_3_n37) );
  DFFR_X1 pe_1_4_3_int_q_acc_reg_6_ ( .D(pe_1_4_3_n78), .CK(pe_1_4_3_net4822), 
        .RN(pe_1_4_3_n71), .Q(int_data_res_4__3__6_) );
  DFFR_X1 pe_1_4_3_int_q_acc_reg_5_ ( .D(pe_1_4_3_n79), .CK(pe_1_4_3_net4822), 
        .RN(pe_1_4_3_n71), .Q(int_data_res_4__3__5_) );
  DFFR_X1 pe_1_4_3_int_q_acc_reg_4_ ( .D(pe_1_4_3_n80), .CK(pe_1_4_3_net4822), 
        .RN(pe_1_4_3_n71), .Q(int_data_res_4__3__4_) );
  DFFR_X1 pe_1_4_3_int_q_acc_reg_3_ ( .D(pe_1_4_3_n81), .CK(pe_1_4_3_net4822), 
        .RN(pe_1_4_3_n71), .Q(int_data_res_4__3__3_) );
  DFFR_X1 pe_1_4_3_int_q_acc_reg_2_ ( .D(pe_1_4_3_n82), .CK(pe_1_4_3_net4822), 
        .RN(pe_1_4_3_n71), .Q(int_data_res_4__3__2_) );
  DFFR_X1 pe_1_4_3_int_q_acc_reg_1_ ( .D(pe_1_4_3_n83), .CK(pe_1_4_3_net4822), 
        .RN(pe_1_4_3_n71), .Q(int_data_res_4__3__1_) );
  DFFR_X1 pe_1_4_3_int_q_acc_reg_7_ ( .D(pe_1_4_3_n77), .CK(pe_1_4_3_net4822), 
        .RN(pe_1_4_3_n71), .Q(int_data_res_4__3__7_) );
  CLKGATETST_X1 pe_1_4_3_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_4_3_n88), .SE(1'b0), .GCK(pe_1_4_3_net4761) );
  CLKGATETST_X1 pe_1_4_3_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_4_3_n87), .SE(1'b0), .GCK(pe_1_4_3_net4767) );
  CLKGATETST_X1 pe_1_4_3_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_4_3_n86), .SE(1'b0), .GCK(pe_1_4_3_net4772) );
  CLKGATETST_X1 pe_1_4_3_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_4_3_n85), .SE(1'b0), .GCK(pe_1_4_3_net4777) );
  CLKGATETST_X1 pe_1_4_3_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_4_3_n90), .SE(1'b0), .GCK(pe_1_4_3_net4782) );
  CLKGATETST_X1 pe_1_4_3_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_4_3_n89), .SE(1'b0), .GCK(pe_1_4_3_net4787) );
  CLKGATETST_X1 pe_1_4_3_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_4_3_N64), .SE(1'b0), .GCK(pe_1_4_3_net4792) );
  CLKGATETST_X1 pe_1_4_3_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_4_3_N63), .SE(1'b0), .GCK(pe_1_4_3_net4797) );
  CLKGATETST_X1 pe_1_4_3_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_4_3_N62), .SE(1'b0), .GCK(pe_1_4_3_net4802) );
  CLKGATETST_X1 pe_1_4_3_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_4_3_N61), .SE(1'b0), .GCK(pe_1_4_3_net4807) );
  CLKGATETST_X1 pe_1_4_3_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_4_3_N60), .SE(1'b0), .GCK(pe_1_4_3_net4812) );
  CLKGATETST_X1 pe_1_4_3_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_4_3_N59), .SE(1'b0), .GCK(pe_1_4_3_net4817) );
  CLKGATETST_X1 pe_1_4_3_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_4_3_N90), .SE(1'b0), .GCK(pe_1_4_3_net4822) );
  CLKBUF_X1 pe_1_4_4_U108 ( .A(pe_1_4_4_n68), .Z(pe_1_4_4_n67) );
  INV_X1 pe_1_4_4_U107 ( .A(n76), .ZN(pe_1_4_4_n66) );
  INV_X1 pe_1_4_4_U106 ( .A(n68), .ZN(pe_1_4_4_n65) );
  INV_X1 pe_1_4_4_U105 ( .A(n68), .ZN(pe_1_4_4_n64) );
  INV_X1 pe_1_4_4_U104 ( .A(pe_1_4_4_n65), .ZN(pe_1_4_4_n63) );
  INV_X1 pe_1_4_4_U103 ( .A(n28), .ZN(pe_1_4_4_n58) );
  INV_X1 pe_1_4_4_U102 ( .A(n20), .ZN(pe_1_4_4_n57) );
  MUX2_X1 pe_1_4_4_U101 ( .A(pe_1_4_4_n54), .B(pe_1_4_4_n51), .S(n50), .Z(
        int_data_x_4__4__3_) );
  MUX2_X1 pe_1_4_4_U100 ( .A(pe_1_4_4_n53), .B(pe_1_4_4_n52), .S(n40), .Z(
        pe_1_4_4_n54) );
  MUX2_X1 pe_1_4_4_U99 ( .A(pe_1_4_4_int_q_reg_h[23]), .B(
        pe_1_4_4_int_q_reg_h[19]), .S(pe_1_4_4_n56), .Z(pe_1_4_4_n53) );
  MUX2_X1 pe_1_4_4_U98 ( .A(pe_1_4_4_int_q_reg_h[15]), .B(
        pe_1_4_4_int_q_reg_h[11]), .S(pe_1_4_4_n56), .Z(pe_1_4_4_n52) );
  MUX2_X1 pe_1_4_4_U97 ( .A(pe_1_4_4_int_q_reg_h[7]), .B(
        pe_1_4_4_int_q_reg_h[3]), .S(pe_1_4_4_n56), .Z(pe_1_4_4_n51) );
  MUX2_X1 pe_1_4_4_U96 ( .A(pe_1_4_4_n50), .B(pe_1_4_4_n47), .S(n50), .Z(
        int_data_x_4__4__2_) );
  MUX2_X1 pe_1_4_4_U95 ( .A(pe_1_4_4_n49), .B(pe_1_4_4_n48), .S(n40), .Z(
        pe_1_4_4_n50) );
  MUX2_X1 pe_1_4_4_U94 ( .A(pe_1_4_4_int_q_reg_h[22]), .B(
        pe_1_4_4_int_q_reg_h[18]), .S(pe_1_4_4_n56), .Z(pe_1_4_4_n49) );
  MUX2_X1 pe_1_4_4_U93 ( .A(pe_1_4_4_int_q_reg_h[14]), .B(
        pe_1_4_4_int_q_reg_h[10]), .S(pe_1_4_4_n56), .Z(pe_1_4_4_n48) );
  MUX2_X1 pe_1_4_4_U92 ( .A(pe_1_4_4_int_q_reg_h[6]), .B(
        pe_1_4_4_int_q_reg_h[2]), .S(pe_1_4_4_n56), .Z(pe_1_4_4_n47) );
  MUX2_X1 pe_1_4_4_U91 ( .A(pe_1_4_4_n46), .B(pe_1_4_4_n24), .S(n50), .Z(
        int_data_x_4__4__1_) );
  MUX2_X1 pe_1_4_4_U90 ( .A(pe_1_4_4_n45), .B(pe_1_4_4_n25), .S(n40), .Z(
        pe_1_4_4_n46) );
  MUX2_X1 pe_1_4_4_U89 ( .A(pe_1_4_4_int_q_reg_h[21]), .B(
        pe_1_4_4_int_q_reg_h[17]), .S(pe_1_4_4_n56), .Z(pe_1_4_4_n45) );
  MUX2_X1 pe_1_4_4_U88 ( .A(pe_1_4_4_int_q_reg_h[13]), .B(
        pe_1_4_4_int_q_reg_h[9]), .S(pe_1_4_4_n56), .Z(pe_1_4_4_n25) );
  MUX2_X1 pe_1_4_4_U87 ( .A(pe_1_4_4_int_q_reg_h[5]), .B(
        pe_1_4_4_int_q_reg_h[1]), .S(pe_1_4_4_n56), .Z(pe_1_4_4_n24) );
  MUX2_X1 pe_1_4_4_U86 ( .A(pe_1_4_4_n23), .B(pe_1_4_4_n20), .S(n50), .Z(
        int_data_x_4__4__0_) );
  MUX2_X1 pe_1_4_4_U85 ( .A(pe_1_4_4_n22), .B(pe_1_4_4_n21), .S(n40), .Z(
        pe_1_4_4_n23) );
  MUX2_X1 pe_1_4_4_U84 ( .A(pe_1_4_4_int_q_reg_h[20]), .B(
        pe_1_4_4_int_q_reg_h[16]), .S(pe_1_4_4_n56), .Z(pe_1_4_4_n22) );
  MUX2_X1 pe_1_4_4_U83 ( .A(pe_1_4_4_int_q_reg_h[12]), .B(
        pe_1_4_4_int_q_reg_h[8]), .S(pe_1_4_4_n56), .Z(pe_1_4_4_n21) );
  MUX2_X1 pe_1_4_4_U82 ( .A(pe_1_4_4_int_q_reg_h[4]), .B(
        pe_1_4_4_int_q_reg_h[0]), .S(pe_1_4_4_n56), .Z(pe_1_4_4_n20) );
  MUX2_X1 pe_1_4_4_U81 ( .A(pe_1_4_4_n19), .B(pe_1_4_4_n16), .S(n50), .Z(
        int_data_y_4__4__3_) );
  MUX2_X1 pe_1_4_4_U80 ( .A(pe_1_4_4_n18), .B(pe_1_4_4_n17), .S(n40), .Z(
        pe_1_4_4_n19) );
  MUX2_X1 pe_1_4_4_U79 ( .A(pe_1_4_4_int_q_reg_v[23]), .B(
        pe_1_4_4_int_q_reg_v[19]), .S(pe_1_4_4_n55), .Z(pe_1_4_4_n18) );
  MUX2_X1 pe_1_4_4_U78 ( .A(pe_1_4_4_int_q_reg_v[15]), .B(
        pe_1_4_4_int_q_reg_v[11]), .S(pe_1_4_4_n55), .Z(pe_1_4_4_n17) );
  MUX2_X1 pe_1_4_4_U77 ( .A(pe_1_4_4_int_q_reg_v[7]), .B(
        pe_1_4_4_int_q_reg_v[3]), .S(pe_1_4_4_n55), .Z(pe_1_4_4_n16) );
  MUX2_X1 pe_1_4_4_U76 ( .A(pe_1_4_4_n15), .B(pe_1_4_4_n12), .S(n50), .Z(
        int_data_y_4__4__2_) );
  MUX2_X1 pe_1_4_4_U75 ( .A(pe_1_4_4_n14), .B(pe_1_4_4_n13), .S(n40), .Z(
        pe_1_4_4_n15) );
  MUX2_X1 pe_1_4_4_U74 ( .A(pe_1_4_4_int_q_reg_v[22]), .B(
        pe_1_4_4_int_q_reg_v[18]), .S(pe_1_4_4_n55), .Z(pe_1_4_4_n14) );
  MUX2_X1 pe_1_4_4_U73 ( .A(pe_1_4_4_int_q_reg_v[14]), .B(
        pe_1_4_4_int_q_reg_v[10]), .S(pe_1_4_4_n55), .Z(pe_1_4_4_n13) );
  MUX2_X1 pe_1_4_4_U72 ( .A(pe_1_4_4_int_q_reg_v[6]), .B(
        pe_1_4_4_int_q_reg_v[2]), .S(pe_1_4_4_n55), .Z(pe_1_4_4_n12) );
  MUX2_X1 pe_1_4_4_U71 ( .A(pe_1_4_4_n11), .B(pe_1_4_4_n8), .S(n50), .Z(
        int_data_y_4__4__1_) );
  MUX2_X1 pe_1_4_4_U70 ( .A(pe_1_4_4_n10), .B(pe_1_4_4_n9), .S(n40), .Z(
        pe_1_4_4_n11) );
  MUX2_X1 pe_1_4_4_U69 ( .A(pe_1_4_4_int_q_reg_v[21]), .B(
        pe_1_4_4_int_q_reg_v[17]), .S(pe_1_4_4_n55), .Z(pe_1_4_4_n10) );
  MUX2_X1 pe_1_4_4_U68 ( .A(pe_1_4_4_int_q_reg_v[13]), .B(
        pe_1_4_4_int_q_reg_v[9]), .S(pe_1_4_4_n55), .Z(pe_1_4_4_n9) );
  MUX2_X1 pe_1_4_4_U67 ( .A(pe_1_4_4_int_q_reg_v[5]), .B(
        pe_1_4_4_int_q_reg_v[1]), .S(pe_1_4_4_n55), .Z(pe_1_4_4_n8) );
  MUX2_X1 pe_1_4_4_U66 ( .A(pe_1_4_4_n7), .B(pe_1_4_4_n4), .S(n50), .Z(
        int_data_y_4__4__0_) );
  MUX2_X1 pe_1_4_4_U65 ( .A(pe_1_4_4_n6), .B(pe_1_4_4_n5), .S(n40), .Z(
        pe_1_4_4_n7) );
  MUX2_X1 pe_1_4_4_U64 ( .A(pe_1_4_4_int_q_reg_v[20]), .B(
        pe_1_4_4_int_q_reg_v[16]), .S(pe_1_4_4_n55), .Z(pe_1_4_4_n6) );
  MUX2_X1 pe_1_4_4_U63 ( .A(pe_1_4_4_int_q_reg_v[12]), .B(
        pe_1_4_4_int_q_reg_v[8]), .S(pe_1_4_4_n55), .Z(pe_1_4_4_n5) );
  MUX2_X1 pe_1_4_4_U62 ( .A(pe_1_4_4_int_q_reg_v[4]), .B(
        pe_1_4_4_int_q_reg_v[0]), .S(pe_1_4_4_n55), .Z(pe_1_4_4_n4) );
  AOI222_X1 pe_1_4_4_U61 ( .A1(int_data_res_5__4__2_), .A2(pe_1_4_4_n61), .B1(
        pe_1_4_4_N80), .B2(pe_1_4_4_n27), .C1(pe_1_4_4_N72), .C2(pe_1_4_4_n28), 
        .ZN(pe_1_4_4_n33) );
  INV_X1 pe_1_4_4_U60 ( .A(pe_1_4_4_n33), .ZN(pe_1_4_4_n78) );
  AOI222_X1 pe_1_4_4_U59 ( .A1(int_data_res_5__4__6_), .A2(pe_1_4_4_n61), .B1(
        pe_1_4_4_N84), .B2(pe_1_4_4_n27), .C1(pe_1_4_4_N76), .C2(pe_1_4_4_n28), 
        .ZN(pe_1_4_4_n29) );
  INV_X1 pe_1_4_4_U58 ( .A(pe_1_4_4_n29), .ZN(pe_1_4_4_n74) );
  XNOR2_X1 pe_1_4_4_U57 ( .A(pe_1_4_4_n69), .B(int_data_res_4__4__0_), .ZN(
        pe_1_4_4_N70) );
  AOI222_X1 pe_1_4_4_U52 ( .A1(int_data_res_5__4__0_), .A2(pe_1_4_4_n61), .B1(
        pe_1_4_4_n1), .B2(pe_1_4_4_n27), .C1(pe_1_4_4_N70), .C2(pe_1_4_4_n28), 
        .ZN(pe_1_4_4_n35) );
  INV_X1 pe_1_4_4_U51 ( .A(pe_1_4_4_n35), .ZN(pe_1_4_4_n80) );
  AOI222_X1 pe_1_4_4_U50 ( .A1(int_data_res_5__4__1_), .A2(pe_1_4_4_n61), .B1(
        pe_1_4_4_N79), .B2(pe_1_4_4_n27), .C1(pe_1_4_4_N71), .C2(pe_1_4_4_n28), 
        .ZN(pe_1_4_4_n34) );
  INV_X1 pe_1_4_4_U49 ( .A(pe_1_4_4_n34), .ZN(pe_1_4_4_n79) );
  AOI222_X1 pe_1_4_4_U48 ( .A1(int_data_res_5__4__3_), .A2(pe_1_4_4_n61), .B1(
        pe_1_4_4_N81), .B2(pe_1_4_4_n27), .C1(pe_1_4_4_N73), .C2(pe_1_4_4_n28), 
        .ZN(pe_1_4_4_n32) );
  INV_X1 pe_1_4_4_U47 ( .A(pe_1_4_4_n32), .ZN(pe_1_4_4_n77) );
  AOI222_X1 pe_1_4_4_U46 ( .A1(int_data_res_5__4__4_), .A2(pe_1_4_4_n61), .B1(
        pe_1_4_4_N82), .B2(pe_1_4_4_n27), .C1(pe_1_4_4_N74), .C2(pe_1_4_4_n28), 
        .ZN(pe_1_4_4_n31) );
  INV_X1 pe_1_4_4_U45 ( .A(pe_1_4_4_n31), .ZN(pe_1_4_4_n76) );
  AOI222_X1 pe_1_4_4_U44 ( .A1(int_data_res_5__4__5_), .A2(pe_1_4_4_n61), .B1(
        pe_1_4_4_N83), .B2(pe_1_4_4_n27), .C1(pe_1_4_4_N75), .C2(pe_1_4_4_n28), 
        .ZN(pe_1_4_4_n30) );
  INV_X1 pe_1_4_4_U43 ( .A(pe_1_4_4_n30), .ZN(pe_1_4_4_n75) );
  NAND2_X1 pe_1_4_4_U42 ( .A1(pe_1_4_4_int_data_0_), .A2(pe_1_4_4_n3), .ZN(
        pe_1_4_4_sub_81_carry[1]) );
  INV_X1 pe_1_4_4_U41 ( .A(pe_1_4_4_int_data_1_), .ZN(pe_1_4_4_n70) );
  INV_X1 pe_1_4_4_U40 ( .A(pe_1_4_4_int_data_2_), .ZN(pe_1_4_4_n71) );
  AND2_X1 pe_1_4_4_U39 ( .A1(pe_1_4_4_int_data_0_), .A2(int_data_res_4__4__0_), 
        .ZN(pe_1_4_4_n2) );
  AOI222_X1 pe_1_4_4_U38 ( .A1(pe_1_4_4_n61), .A2(int_data_res_5__4__7_), .B1(
        pe_1_4_4_N85), .B2(pe_1_4_4_n27), .C1(pe_1_4_4_N77), .C2(pe_1_4_4_n28), 
        .ZN(pe_1_4_4_n26) );
  INV_X1 pe_1_4_4_U37 ( .A(pe_1_4_4_n26), .ZN(pe_1_4_4_n73) );
  NOR3_X1 pe_1_4_4_U36 ( .A1(pe_1_4_4_n58), .A2(pe_1_4_4_n62), .A3(int_ckg[27]), .ZN(pe_1_4_4_n36) );
  OR2_X1 pe_1_4_4_U35 ( .A1(pe_1_4_4_n36), .A2(pe_1_4_4_n61), .ZN(pe_1_4_4_N90) );
  INV_X1 pe_1_4_4_U34 ( .A(n40), .ZN(pe_1_4_4_n60) );
  AND2_X1 pe_1_4_4_U33 ( .A1(int_data_x_4__4__2_), .A2(n28), .ZN(
        pe_1_4_4_int_data_2_) );
  AND2_X1 pe_1_4_4_U32 ( .A1(int_data_x_4__4__1_), .A2(n28), .ZN(
        pe_1_4_4_int_data_1_) );
  AND2_X1 pe_1_4_4_U31 ( .A1(int_data_x_4__4__3_), .A2(n28), .ZN(
        pe_1_4_4_int_data_3_) );
  BUF_X1 pe_1_4_4_U30 ( .A(n62), .Z(pe_1_4_4_n61) );
  INV_X1 pe_1_4_4_U29 ( .A(n34), .ZN(pe_1_4_4_n59) );
  AND2_X1 pe_1_4_4_U28 ( .A1(int_data_x_4__4__0_), .A2(n28), .ZN(
        pe_1_4_4_int_data_0_) );
  NAND2_X1 pe_1_4_4_U27 ( .A1(pe_1_4_4_n44), .A2(pe_1_4_4_n59), .ZN(
        pe_1_4_4_n41) );
  AND3_X1 pe_1_4_4_U26 ( .A1(n76), .A2(pe_1_4_4_n60), .A3(n50), .ZN(
        pe_1_4_4_n44) );
  INV_X1 pe_1_4_4_U25 ( .A(pe_1_4_4_int_data_3_), .ZN(pe_1_4_4_n72) );
  NOR2_X1 pe_1_4_4_U24 ( .A1(pe_1_4_4_n66), .A2(n50), .ZN(pe_1_4_4_n43) );
  NOR2_X1 pe_1_4_4_U23 ( .A1(pe_1_4_4_n57), .A2(pe_1_4_4_n61), .ZN(
        pe_1_4_4_n28) );
  NOR2_X1 pe_1_4_4_U22 ( .A1(n20), .A2(pe_1_4_4_n61), .ZN(pe_1_4_4_n27) );
  INV_X1 pe_1_4_4_U21 ( .A(pe_1_4_4_int_data_0_), .ZN(pe_1_4_4_n69) );
  INV_X1 pe_1_4_4_U20 ( .A(pe_1_4_4_n41), .ZN(pe_1_4_4_n86) );
  INV_X1 pe_1_4_4_U19 ( .A(pe_1_4_4_n37), .ZN(pe_1_4_4_n84) );
  INV_X1 pe_1_4_4_U18 ( .A(pe_1_4_4_n38), .ZN(pe_1_4_4_n83) );
  INV_X1 pe_1_4_4_U17 ( .A(pe_1_4_4_n39), .ZN(pe_1_4_4_n82) );
  NOR2_X1 pe_1_4_4_U16 ( .A1(pe_1_4_4_n64), .A2(pe_1_4_4_n42), .ZN(
        pe_1_4_4_N59) );
  NOR2_X1 pe_1_4_4_U15 ( .A1(pe_1_4_4_n64), .A2(pe_1_4_4_n41), .ZN(
        pe_1_4_4_N60) );
  NOR2_X1 pe_1_4_4_U14 ( .A1(pe_1_4_4_n64), .A2(pe_1_4_4_n38), .ZN(
        pe_1_4_4_N63) );
  NOR2_X1 pe_1_4_4_U13 ( .A1(pe_1_4_4_n64), .A2(pe_1_4_4_n40), .ZN(
        pe_1_4_4_N61) );
  NOR2_X1 pe_1_4_4_U12 ( .A1(pe_1_4_4_n64), .A2(pe_1_4_4_n39), .ZN(
        pe_1_4_4_N62) );
  NOR2_X1 pe_1_4_4_U11 ( .A1(pe_1_4_4_n37), .A2(pe_1_4_4_n64), .ZN(
        pe_1_4_4_N64) );
  NAND2_X1 pe_1_4_4_U10 ( .A1(pe_1_4_4_n44), .A2(n34), .ZN(pe_1_4_4_n42) );
  BUF_X1 pe_1_4_4_U9 ( .A(n34), .Z(pe_1_4_4_n55) );
  INV_X1 pe_1_4_4_U8 ( .A(pe_1_4_4_n65), .ZN(pe_1_4_4_n62) );
  BUF_X1 pe_1_4_4_U7 ( .A(n34), .Z(pe_1_4_4_n56) );
  INV_X1 pe_1_4_4_U6 ( .A(pe_1_4_4_n42), .ZN(pe_1_4_4_n85) );
  INV_X1 pe_1_4_4_U5 ( .A(pe_1_4_4_n40), .ZN(pe_1_4_4_n81) );
  INV_X2 pe_1_4_4_U4 ( .A(n84), .ZN(pe_1_4_4_n68) );
  XOR2_X1 pe_1_4_4_U3 ( .A(pe_1_4_4_int_data_0_), .B(int_data_res_4__4__0_), 
        .Z(pe_1_4_4_n1) );
  DFFR_X1 pe_1_4_4_int_q_acc_reg_0_ ( .D(pe_1_4_4_n80), .CK(pe_1_4_4_net4744), 
        .RN(pe_1_4_4_n68), .Q(int_data_res_4__4__0_), .QN(pe_1_4_4_n3) );
  DFFR_X1 pe_1_4_4_int_q_reg_v_reg_0__0_ ( .D(int_data_y_5__4__0_), .CK(
        pe_1_4_4_net4714), .RN(pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_v[20]) );
  DFFR_X1 pe_1_4_4_int_q_reg_v_reg_0__1_ ( .D(int_data_y_5__4__1_), .CK(
        pe_1_4_4_net4714), .RN(pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_v[21]) );
  DFFR_X1 pe_1_4_4_int_q_reg_v_reg_0__2_ ( .D(int_data_y_5__4__2_), .CK(
        pe_1_4_4_net4714), .RN(pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_v[22]) );
  DFFR_X1 pe_1_4_4_int_q_reg_v_reg_0__3_ ( .D(int_data_y_5__4__3_), .CK(
        pe_1_4_4_net4714), .RN(pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_v[23]) );
  DFFR_X1 pe_1_4_4_int_q_reg_v_reg_1__0_ ( .D(int_data_y_5__4__0_), .CK(
        pe_1_4_4_net4719), .RN(pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_v[16]) );
  DFFR_X1 pe_1_4_4_int_q_reg_v_reg_1__1_ ( .D(int_data_y_5__4__1_), .CK(
        pe_1_4_4_net4719), .RN(pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_v[17]) );
  DFFR_X1 pe_1_4_4_int_q_reg_v_reg_1__2_ ( .D(int_data_y_5__4__2_), .CK(
        pe_1_4_4_net4719), .RN(pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_v[18]) );
  DFFR_X1 pe_1_4_4_int_q_reg_v_reg_1__3_ ( .D(int_data_y_5__4__3_), .CK(
        pe_1_4_4_net4719), .RN(pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_v[19]) );
  DFFR_X1 pe_1_4_4_int_q_reg_v_reg_2__0_ ( .D(int_data_y_5__4__0_), .CK(
        pe_1_4_4_net4724), .RN(pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_v[12]) );
  DFFR_X1 pe_1_4_4_int_q_reg_v_reg_2__1_ ( .D(int_data_y_5__4__1_), .CK(
        pe_1_4_4_net4724), .RN(pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_v[13]) );
  DFFR_X1 pe_1_4_4_int_q_reg_v_reg_2__2_ ( .D(int_data_y_5__4__2_), .CK(
        pe_1_4_4_net4724), .RN(pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_v[14]) );
  DFFR_X1 pe_1_4_4_int_q_reg_v_reg_2__3_ ( .D(int_data_y_5__4__3_), .CK(
        pe_1_4_4_net4724), .RN(pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_v[15]) );
  DFFR_X1 pe_1_4_4_int_q_reg_v_reg_3__0_ ( .D(int_data_y_5__4__0_), .CK(
        pe_1_4_4_net4729), .RN(pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_v[8]) );
  DFFR_X1 pe_1_4_4_int_q_reg_v_reg_3__1_ ( .D(int_data_y_5__4__1_), .CK(
        pe_1_4_4_net4729), .RN(pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_v[9]) );
  DFFR_X1 pe_1_4_4_int_q_reg_v_reg_3__2_ ( .D(int_data_y_5__4__2_), .CK(
        pe_1_4_4_net4729), .RN(pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_v[10]) );
  DFFR_X1 pe_1_4_4_int_q_reg_v_reg_3__3_ ( .D(int_data_y_5__4__3_), .CK(
        pe_1_4_4_net4729), .RN(pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_v[11]) );
  DFFR_X1 pe_1_4_4_int_q_reg_v_reg_4__0_ ( .D(int_data_y_5__4__0_), .CK(
        pe_1_4_4_net4734), .RN(pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_v[4]) );
  DFFR_X1 pe_1_4_4_int_q_reg_v_reg_4__1_ ( .D(int_data_y_5__4__1_), .CK(
        pe_1_4_4_net4734), .RN(pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_v[5]) );
  DFFR_X1 pe_1_4_4_int_q_reg_v_reg_4__2_ ( .D(int_data_y_5__4__2_), .CK(
        pe_1_4_4_net4734), .RN(pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_v[6]) );
  DFFR_X1 pe_1_4_4_int_q_reg_v_reg_4__3_ ( .D(int_data_y_5__4__3_), .CK(
        pe_1_4_4_net4734), .RN(pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_v[7]) );
  DFFR_X1 pe_1_4_4_int_q_reg_v_reg_5__0_ ( .D(int_data_y_5__4__0_), .CK(
        pe_1_4_4_net4739), .RN(pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_v[0]) );
  DFFR_X1 pe_1_4_4_int_q_reg_v_reg_5__1_ ( .D(int_data_y_5__4__1_), .CK(
        pe_1_4_4_net4739), .RN(pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_v[1]) );
  DFFR_X1 pe_1_4_4_int_q_reg_v_reg_5__2_ ( .D(int_data_y_5__4__2_), .CK(
        pe_1_4_4_net4739), .RN(pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_v[2]) );
  DFFR_X1 pe_1_4_4_int_q_reg_v_reg_5__3_ ( .D(int_data_y_5__4__3_), .CK(
        pe_1_4_4_net4739), .RN(pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_4_4_int_q_reg_h_reg_0__0_ ( .D(int_data_x_4__5__0_), .SI(
        int_data_y_5__4__0_), .SE(pe_1_4_4_n62), .CK(pe_1_4_4_net4683), .RN(
        pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_4_4_int_q_reg_h_reg_0__1_ ( .D(int_data_x_4__5__1_), .SI(
        int_data_y_5__4__1_), .SE(pe_1_4_4_n62), .CK(pe_1_4_4_net4683), .RN(
        pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_4_4_int_q_reg_h_reg_0__2_ ( .D(int_data_x_4__5__2_), .SI(
        int_data_y_5__4__2_), .SE(pe_1_4_4_n62), .CK(pe_1_4_4_net4683), .RN(
        pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_4_4_int_q_reg_h_reg_0__3_ ( .D(int_data_x_4__5__3_), .SI(
        int_data_y_5__4__3_), .SE(pe_1_4_4_n62), .CK(pe_1_4_4_net4683), .RN(
        pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_4_4_int_q_reg_h_reg_1__0_ ( .D(int_data_x_4__5__0_), .SI(
        int_data_y_5__4__0_), .SE(pe_1_4_4_n62), .CK(pe_1_4_4_net4689), .RN(
        pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_4_4_int_q_reg_h_reg_1__1_ ( .D(int_data_x_4__5__1_), .SI(
        int_data_y_5__4__1_), .SE(pe_1_4_4_n62), .CK(pe_1_4_4_net4689), .RN(
        pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_4_4_int_q_reg_h_reg_1__2_ ( .D(int_data_x_4__5__2_), .SI(
        int_data_y_5__4__2_), .SE(pe_1_4_4_n62), .CK(pe_1_4_4_net4689), .RN(
        pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_4_4_int_q_reg_h_reg_1__3_ ( .D(int_data_x_4__5__3_), .SI(
        int_data_y_5__4__3_), .SE(pe_1_4_4_n62), .CK(pe_1_4_4_net4689), .RN(
        pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_4_4_int_q_reg_h_reg_2__0_ ( .D(int_data_x_4__5__0_), .SI(
        int_data_y_5__4__0_), .SE(pe_1_4_4_n62), .CK(pe_1_4_4_net4694), .RN(
        pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_4_4_int_q_reg_h_reg_2__1_ ( .D(int_data_x_4__5__1_), .SI(
        int_data_y_5__4__1_), .SE(pe_1_4_4_n62), .CK(pe_1_4_4_net4694), .RN(
        pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_4_4_int_q_reg_h_reg_2__2_ ( .D(int_data_x_4__5__2_), .SI(
        int_data_y_5__4__2_), .SE(pe_1_4_4_n62), .CK(pe_1_4_4_net4694), .RN(
        pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_4_4_int_q_reg_h_reg_2__3_ ( .D(int_data_x_4__5__3_), .SI(
        int_data_y_5__4__3_), .SE(pe_1_4_4_n62), .CK(pe_1_4_4_net4694), .RN(
        pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_4_4_int_q_reg_h_reg_3__0_ ( .D(int_data_x_4__5__0_), .SI(
        int_data_y_5__4__0_), .SE(pe_1_4_4_n62), .CK(pe_1_4_4_net4699), .RN(
        pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_4_4_int_q_reg_h_reg_3__1_ ( .D(int_data_x_4__5__1_), .SI(
        int_data_y_5__4__1_), .SE(pe_1_4_4_n62), .CK(pe_1_4_4_net4699), .RN(
        pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_4_4_int_q_reg_h_reg_3__2_ ( .D(int_data_x_4__5__2_), .SI(
        int_data_y_5__4__2_), .SE(pe_1_4_4_n62), .CK(pe_1_4_4_net4699), .RN(
        pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_4_4_int_q_reg_h_reg_3__3_ ( .D(int_data_x_4__5__3_), .SI(
        int_data_y_5__4__3_), .SE(pe_1_4_4_n62), .CK(pe_1_4_4_net4699), .RN(
        pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_4_4_int_q_reg_h_reg_4__0_ ( .D(int_data_x_4__5__0_), .SI(
        int_data_y_5__4__0_), .SE(pe_1_4_4_n63), .CK(pe_1_4_4_net4704), .RN(
        pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_4_4_int_q_reg_h_reg_4__1_ ( .D(int_data_x_4__5__1_), .SI(
        int_data_y_5__4__1_), .SE(pe_1_4_4_n63), .CK(pe_1_4_4_net4704), .RN(
        pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_4_4_int_q_reg_h_reg_4__2_ ( .D(int_data_x_4__5__2_), .SI(
        int_data_y_5__4__2_), .SE(pe_1_4_4_n63), .CK(pe_1_4_4_net4704), .RN(
        pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_4_4_int_q_reg_h_reg_4__3_ ( .D(int_data_x_4__5__3_), .SI(
        int_data_y_5__4__3_), .SE(pe_1_4_4_n63), .CK(pe_1_4_4_net4704), .RN(
        pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_4_4_int_q_reg_h_reg_5__0_ ( .D(int_data_x_4__5__0_), .SI(
        int_data_y_5__4__0_), .SE(pe_1_4_4_n63), .CK(pe_1_4_4_net4709), .RN(
        pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_4_4_int_q_reg_h_reg_5__1_ ( .D(int_data_x_4__5__1_), .SI(
        int_data_y_5__4__1_), .SE(pe_1_4_4_n63), .CK(pe_1_4_4_net4709), .RN(
        pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_4_4_int_q_reg_h_reg_5__2_ ( .D(int_data_x_4__5__2_), .SI(
        int_data_y_5__4__2_), .SE(pe_1_4_4_n63), .CK(pe_1_4_4_net4709), .RN(
        pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_4_4_int_q_reg_h_reg_5__3_ ( .D(int_data_x_4__5__3_), .SI(
        int_data_y_5__4__3_), .SE(pe_1_4_4_n63), .CK(pe_1_4_4_net4709), .RN(
        pe_1_4_4_n68), .Q(pe_1_4_4_int_q_reg_h[3]) );
  FA_X1 pe_1_4_4_sub_81_U2_7 ( .A(int_data_res_4__4__7_), .B(pe_1_4_4_n72), 
        .CI(pe_1_4_4_sub_81_carry[7]), .S(pe_1_4_4_N77) );
  FA_X1 pe_1_4_4_sub_81_U2_6 ( .A(int_data_res_4__4__6_), .B(pe_1_4_4_n72), 
        .CI(pe_1_4_4_sub_81_carry[6]), .CO(pe_1_4_4_sub_81_carry[7]), .S(
        pe_1_4_4_N76) );
  FA_X1 pe_1_4_4_sub_81_U2_5 ( .A(int_data_res_4__4__5_), .B(pe_1_4_4_n72), 
        .CI(pe_1_4_4_sub_81_carry[5]), .CO(pe_1_4_4_sub_81_carry[6]), .S(
        pe_1_4_4_N75) );
  FA_X1 pe_1_4_4_sub_81_U2_4 ( .A(int_data_res_4__4__4_), .B(pe_1_4_4_n72), 
        .CI(pe_1_4_4_sub_81_carry[4]), .CO(pe_1_4_4_sub_81_carry[5]), .S(
        pe_1_4_4_N74) );
  FA_X1 pe_1_4_4_sub_81_U2_3 ( .A(int_data_res_4__4__3_), .B(pe_1_4_4_n72), 
        .CI(pe_1_4_4_sub_81_carry[3]), .CO(pe_1_4_4_sub_81_carry[4]), .S(
        pe_1_4_4_N73) );
  FA_X1 pe_1_4_4_sub_81_U2_2 ( .A(int_data_res_4__4__2_), .B(pe_1_4_4_n71), 
        .CI(pe_1_4_4_sub_81_carry[2]), .CO(pe_1_4_4_sub_81_carry[3]), .S(
        pe_1_4_4_N72) );
  FA_X1 pe_1_4_4_sub_81_U2_1 ( .A(int_data_res_4__4__1_), .B(pe_1_4_4_n70), 
        .CI(pe_1_4_4_sub_81_carry[1]), .CO(pe_1_4_4_sub_81_carry[2]), .S(
        pe_1_4_4_N71) );
  FA_X1 pe_1_4_4_add_83_U1_7 ( .A(int_data_res_4__4__7_), .B(
        pe_1_4_4_int_data_3_), .CI(pe_1_4_4_add_83_carry[7]), .S(pe_1_4_4_N85)
         );
  FA_X1 pe_1_4_4_add_83_U1_6 ( .A(int_data_res_4__4__6_), .B(
        pe_1_4_4_int_data_3_), .CI(pe_1_4_4_add_83_carry[6]), .CO(
        pe_1_4_4_add_83_carry[7]), .S(pe_1_4_4_N84) );
  FA_X1 pe_1_4_4_add_83_U1_5 ( .A(int_data_res_4__4__5_), .B(
        pe_1_4_4_int_data_3_), .CI(pe_1_4_4_add_83_carry[5]), .CO(
        pe_1_4_4_add_83_carry[6]), .S(pe_1_4_4_N83) );
  FA_X1 pe_1_4_4_add_83_U1_4 ( .A(int_data_res_4__4__4_), .B(
        pe_1_4_4_int_data_3_), .CI(pe_1_4_4_add_83_carry[4]), .CO(
        pe_1_4_4_add_83_carry[5]), .S(pe_1_4_4_N82) );
  FA_X1 pe_1_4_4_add_83_U1_3 ( .A(int_data_res_4__4__3_), .B(
        pe_1_4_4_int_data_3_), .CI(pe_1_4_4_add_83_carry[3]), .CO(
        pe_1_4_4_add_83_carry[4]), .S(pe_1_4_4_N81) );
  FA_X1 pe_1_4_4_add_83_U1_2 ( .A(int_data_res_4__4__2_), .B(
        pe_1_4_4_int_data_2_), .CI(pe_1_4_4_add_83_carry[2]), .CO(
        pe_1_4_4_add_83_carry[3]), .S(pe_1_4_4_N80) );
  FA_X1 pe_1_4_4_add_83_U1_1 ( .A(int_data_res_4__4__1_), .B(
        pe_1_4_4_int_data_1_), .CI(pe_1_4_4_n2), .CO(pe_1_4_4_add_83_carry[2]), 
        .S(pe_1_4_4_N79) );
  NAND3_X1 pe_1_4_4_U56 ( .A1(n34), .A2(pe_1_4_4_n43), .A3(n40), .ZN(
        pe_1_4_4_n40) );
  NAND3_X1 pe_1_4_4_U55 ( .A1(pe_1_4_4_n43), .A2(pe_1_4_4_n59), .A3(n40), .ZN(
        pe_1_4_4_n39) );
  NAND3_X1 pe_1_4_4_U54 ( .A1(pe_1_4_4_n43), .A2(pe_1_4_4_n60), .A3(n34), .ZN(
        pe_1_4_4_n38) );
  NAND3_X1 pe_1_4_4_U53 ( .A1(pe_1_4_4_n59), .A2(pe_1_4_4_n60), .A3(
        pe_1_4_4_n43), .ZN(pe_1_4_4_n37) );
  DFFR_X1 pe_1_4_4_int_q_acc_reg_6_ ( .D(pe_1_4_4_n74), .CK(pe_1_4_4_net4744), 
        .RN(pe_1_4_4_n67), .Q(int_data_res_4__4__6_) );
  DFFR_X1 pe_1_4_4_int_q_acc_reg_5_ ( .D(pe_1_4_4_n75), .CK(pe_1_4_4_net4744), 
        .RN(pe_1_4_4_n67), .Q(int_data_res_4__4__5_) );
  DFFR_X1 pe_1_4_4_int_q_acc_reg_4_ ( .D(pe_1_4_4_n76), .CK(pe_1_4_4_net4744), 
        .RN(pe_1_4_4_n67), .Q(int_data_res_4__4__4_) );
  DFFR_X1 pe_1_4_4_int_q_acc_reg_3_ ( .D(pe_1_4_4_n77), .CK(pe_1_4_4_net4744), 
        .RN(pe_1_4_4_n67), .Q(int_data_res_4__4__3_) );
  DFFR_X1 pe_1_4_4_int_q_acc_reg_2_ ( .D(pe_1_4_4_n78), .CK(pe_1_4_4_net4744), 
        .RN(pe_1_4_4_n67), .Q(int_data_res_4__4__2_) );
  DFFR_X1 pe_1_4_4_int_q_acc_reg_1_ ( .D(pe_1_4_4_n79), .CK(pe_1_4_4_net4744), 
        .RN(pe_1_4_4_n67), .Q(int_data_res_4__4__1_) );
  DFFR_X1 pe_1_4_4_int_q_acc_reg_7_ ( .D(pe_1_4_4_n73), .CK(pe_1_4_4_net4744), 
        .RN(pe_1_4_4_n67), .Q(int_data_res_4__4__7_) );
  CLKGATETST_X1 pe_1_4_4_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_4_4_n84), .SE(1'b0), .GCK(pe_1_4_4_net4683) );
  CLKGATETST_X1 pe_1_4_4_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_4_4_n83), .SE(1'b0), .GCK(pe_1_4_4_net4689) );
  CLKGATETST_X1 pe_1_4_4_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_4_4_n82), .SE(1'b0), .GCK(pe_1_4_4_net4694) );
  CLKGATETST_X1 pe_1_4_4_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_4_4_n81), .SE(1'b0), .GCK(pe_1_4_4_net4699) );
  CLKGATETST_X1 pe_1_4_4_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_4_4_n86), .SE(1'b0), .GCK(pe_1_4_4_net4704) );
  CLKGATETST_X1 pe_1_4_4_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_4_4_n85), .SE(1'b0), .GCK(pe_1_4_4_net4709) );
  CLKGATETST_X1 pe_1_4_4_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_4_4_N64), .SE(1'b0), .GCK(pe_1_4_4_net4714) );
  CLKGATETST_X1 pe_1_4_4_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_4_4_N63), .SE(1'b0), .GCK(pe_1_4_4_net4719) );
  CLKGATETST_X1 pe_1_4_4_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_4_4_N62), .SE(1'b0), .GCK(pe_1_4_4_net4724) );
  CLKGATETST_X1 pe_1_4_4_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_4_4_N61), .SE(1'b0), .GCK(pe_1_4_4_net4729) );
  CLKGATETST_X1 pe_1_4_4_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_4_4_N60), .SE(1'b0), .GCK(pe_1_4_4_net4734) );
  CLKGATETST_X1 pe_1_4_4_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_4_4_N59), .SE(1'b0), .GCK(pe_1_4_4_net4739) );
  CLKGATETST_X1 pe_1_4_4_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_4_4_N90), .SE(1'b0), .GCK(pe_1_4_4_net4744) );
  CLKBUF_X1 pe_1_4_5_U109 ( .A(pe_1_4_5_n69), .Z(pe_1_4_5_n68) );
  INV_X1 pe_1_4_5_U108 ( .A(n76), .ZN(pe_1_4_5_n67) );
  INV_X1 pe_1_4_5_U107 ( .A(n68), .ZN(pe_1_4_5_n66) );
  INV_X1 pe_1_4_5_U106 ( .A(n68), .ZN(pe_1_4_5_n65) );
  INV_X1 pe_1_4_5_U105 ( .A(pe_1_4_5_n66), .ZN(pe_1_4_5_n64) );
  INV_X1 pe_1_4_5_U104 ( .A(pe_1_4_5_n61), .ZN(pe_1_4_5_n60) );
  INV_X1 pe_1_4_5_U103 ( .A(n28), .ZN(pe_1_4_5_n58) );
  INV_X1 pe_1_4_5_U102 ( .A(n20), .ZN(pe_1_4_5_n57) );
  MUX2_X1 pe_1_4_5_U101 ( .A(pe_1_4_5_n54), .B(pe_1_4_5_n51), .S(n50), .Z(
        int_data_x_4__5__3_) );
  MUX2_X1 pe_1_4_5_U100 ( .A(pe_1_4_5_n53), .B(pe_1_4_5_n52), .S(pe_1_4_5_n60), 
        .Z(pe_1_4_5_n54) );
  MUX2_X1 pe_1_4_5_U99 ( .A(pe_1_4_5_int_q_reg_h[23]), .B(
        pe_1_4_5_int_q_reg_h[19]), .S(pe_1_4_5_n56), .Z(pe_1_4_5_n53) );
  MUX2_X1 pe_1_4_5_U98 ( .A(pe_1_4_5_int_q_reg_h[15]), .B(
        pe_1_4_5_int_q_reg_h[11]), .S(pe_1_4_5_n56), .Z(pe_1_4_5_n52) );
  MUX2_X1 pe_1_4_5_U97 ( .A(pe_1_4_5_int_q_reg_h[7]), .B(
        pe_1_4_5_int_q_reg_h[3]), .S(pe_1_4_5_n56), .Z(pe_1_4_5_n51) );
  MUX2_X1 pe_1_4_5_U96 ( .A(pe_1_4_5_n50), .B(pe_1_4_5_n47), .S(n50), .Z(
        int_data_x_4__5__2_) );
  MUX2_X1 pe_1_4_5_U95 ( .A(pe_1_4_5_n49), .B(pe_1_4_5_n48), .S(pe_1_4_5_n60), 
        .Z(pe_1_4_5_n50) );
  MUX2_X1 pe_1_4_5_U94 ( .A(pe_1_4_5_int_q_reg_h[22]), .B(
        pe_1_4_5_int_q_reg_h[18]), .S(pe_1_4_5_n56), .Z(pe_1_4_5_n49) );
  MUX2_X1 pe_1_4_5_U93 ( .A(pe_1_4_5_int_q_reg_h[14]), .B(
        pe_1_4_5_int_q_reg_h[10]), .S(pe_1_4_5_n56), .Z(pe_1_4_5_n48) );
  MUX2_X1 pe_1_4_5_U92 ( .A(pe_1_4_5_int_q_reg_h[6]), .B(
        pe_1_4_5_int_q_reg_h[2]), .S(pe_1_4_5_n56), .Z(pe_1_4_5_n47) );
  MUX2_X1 pe_1_4_5_U91 ( .A(pe_1_4_5_n46), .B(pe_1_4_5_n24), .S(n50), .Z(
        int_data_x_4__5__1_) );
  MUX2_X1 pe_1_4_5_U90 ( .A(pe_1_4_5_n45), .B(pe_1_4_5_n25), .S(pe_1_4_5_n60), 
        .Z(pe_1_4_5_n46) );
  MUX2_X1 pe_1_4_5_U89 ( .A(pe_1_4_5_int_q_reg_h[21]), .B(
        pe_1_4_5_int_q_reg_h[17]), .S(pe_1_4_5_n56), .Z(pe_1_4_5_n45) );
  MUX2_X1 pe_1_4_5_U88 ( .A(pe_1_4_5_int_q_reg_h[13]), .B(
        pe_1_4_5_int_q_reg_h[9]), .S(pe_1_4_5_n56), .Z(pe_1_4_5_n25) );
  MUX2_X1 pe_1_4_5_U87 ( .A(pe_1_4_5_int_q_reg_h[5]), .B(
        pe_1_4_5_int_q_reg_h[1]), .S(pe_1_4_5_n56), .Z(pe_1_4_5_n24) );
  MUX2_X1 pe_1_4_5_U86 ( .A(pe_1_4_5_n23), .B(pe_1_4_5_n20), .S(n50), .Z(
        int_data_x_4__5__0_) );
  MUX2_X1 pe_1_4_5_U85 ( .A(pe_1_4_5_n22), .B(pe_1_4_5_n21), .S(pe_1_4_5_n60), 
        .Z(pe_1_4_5_n23) );
  MUX2_X1 pe_1_4_5_U84 ( .A(pe_1_4_5_int_q_reg_h[20]), .B(
        pe_1_4_5_int_q_reg_h[16]), .S(pe_1_4_5_n56), .Z(pe_1_4_5_n22) );
  MUX2_X1 pe_1_4_5_U83 ( .A(pe_1_4_5_int_q_reg_h[12]), .B(
        pe_1_4_5_int_q_reg_h[8]), .S(pe_1_4_5_n56), .Z(pe_1_4_5_n21) );
  MUX2_X1 pe_1_4_5_U82 ( .A(pe_1_4_5_int_q_reg_h[4]), .B(
        pe_1_4_5_int_q_reg_h[0]), .S(pe_1_4_5_n56), .Z(pe_1_4_5_n20) );
  MUX2_X1 pe_1_4_5_U81 ( .A(pe_1_4_5_n19), .B(pe_1_4_5_n16), .S(n50), .Z(
        int_data_y_4__5__3_) );
  MUX2_X1 pe_1_4_5_U80 ( .A(pe_1_4_5_n18), .B(pe_1_4_5_n17), .S(pe_1_4_5_n60), 
        .Z(pe_1_4_5_n19) );
  MUX2_X1 pe_1_4_5_U79 ( .A(pe_1_4_5_int_q_reg_v[23]), .B(
        pe_1_4_5_int_q_reg_v[19]), .S(pe_1_4_5_n55), .Z(pe_1_4_5_n18) );
  MUX2_X1 pe_1_4_5_U78 ( .A(pe_1_4_5_int_q_reg_v[15]), .B(
        pe_1_4_5_int_q_reg_v[11]), .S(pe_1_4_5_n55), .Z(pe_1_4_5_n17) );
  MUX2_X1 pe_1_4_5_U77 ( .A(pe_1_4_5_int_q_reg_v[7]), .B(
        pe_1_4_5_int_q_reg_v[3]), .S(pe_1_4_5_n55), .Z(pe_1_4_5_n16) );
  MUX2_X1 pe_1_4_5_U76 ( .A(pe_1_4_5_n15), .B(pe_1_4_5_n12), .S(n50), .Z(
        int_data_y_4__5__2_) );
  MUX2_X1 pe_1_4_5_U75 ( .A(pe_1_4_5_n14), .B(pe_1_4_5_n13), .S(pe_1_4_5_n60), 
        .Z(pe_1_4_5_n15) );
  MUX2_X1 pe_1_4_5_U74 ( .A(pe_1_4_5_int_q_reg_v[22]), .B(
        pe_1_4_5_int_q_reg_v[18]), .S(pe_1_4_5_n55), .Z(pe_1_4_5_n14) );
  MUX2_X1 pe_1_4_5_U73 ( .A(pe_1_4_5_int_q_reg_v[14]), .B(
        pe_1_4_5_int_q_reg_v[10]), .S(pe_1_4_5_n55), .Z(pe_1_4_5_n13) );
  MUX2_X1 pe_1_4_5_U72 ( .A(pe_1_4_5_int_q_reg_v[6]), .B(
        pe_1_4_5_int_q_reg_v[2]), .S(pe_1_4_5_n55), .Z(pe_1_4_5_n12) );
  MUX2_X1 pe_1_4_5_U71 ( .A(pe_1_4_5_n11), .B(pe_1_4_5_n8), .S(n50), .Z(
        int_data_y_4__5__1_) );
  MUX2_X1 pe_1_4_5_U70 ( .A(pe_1_4_5_n10), .B(pe_1_4_5_n9), .S(pe_1_4_5_n60), 
        .Z(pe_1_4_5_n11) );
  MUX2_X1 pe_1_4_5_U69 ( .A(pe_1_4_5_int_q_reg_v[21]), .B(
        pe_1_4_5_int_q_reg_v[17]), .S(pe_1_4_5_n55), .Z(pe_1_4_5_n10) );
  MUX2_X1 pe_1_4_5_U68 ( .A(pe_1_4_5_int_q_reg_v[13]), .B(
        pe_1_4_5_int_q_reg_v[9]), .S(pe_1_4_5_n55), .Z(pe_1_4_5_n9) );
  MUX2_X1 pe_1_4_5_U67 ( .A(pe_1_4_5_int_q_reg_v[5]), .B(
        pe_1_4_5_int_q_reg_v[1]), .S(pe_1_4_5_n55), .Z(pe_1_4_5_n8) );
  MUX2_X1 pe_1_4_5_U66 ( .A(pe_1_4_5_n7), .B(pe_1_4_5_n4), .S(n50), .Z(
        int_data_y_4__5__0_) );
  MUX2_X1 pe_1_4_5_U65 ( .A(pe_1_4_5_n6), .B(pe_1_4_5_n5), .S(pe_1_4_5_n60), 
        .Z(pe_1_4_5_n7) );
  MUX2_X1 pe_1_4_5_U64 ( .A(pe_1_4_5_int_q_reg_v[20]), .B(
        pe_1_4_5_int_q_reg_v[16]), .S(pe_1_4_5_n55), .Z(pe_1_4_5_n6) );
  MUX2_X1 pe_1_4_5_U63 ( .A(pe_1_4_5_int_q_reg_v[12]), .B(
        pe_1_4_5_int_q_reg_v[8]), .S(pe_1_4_5_n55), .Z(pe_1_4_5_n5) );
  MUX2_X1 pe_1_4_5_U62 ( .A(pe_1_4_5_int_q_reg_v[4]), .B(
        pe_1_4_5_int_q_reg_v[0]), .S(pe_1_4_5_n55), .Z(pe_1_4_5_n4) );
  AOI222_X1 pe_1_4_5_U61 ( .A1(int_data_res_5__5__2_), .A2(pe_1_4_5_n62), .B1(
        pe_1_4_5_N80), .B2(pe_1_4_5_n27), .C1(pe_1_4_5_N72), .C2(pe_1_4_5_n28), 
        .ZN(pe_1_4_5_n33) );
  INV_X1 pe_1_4_5_U60 ( .A(pe_1_4_5_n33), .ZN(pe_1_4_5_n79) );
  AOI222_X1 pe_1_4_5_U59 ( .A1(int_data_res_5__5__6_), .A2(pe_1_4_5_n62), .B1(
        pe_1_4_5_N84), .B2(pe_1_4_5_n27), .C1(pe_1_4_5_N76), .C2(pe_1_4_5_n28), 
        .ZN(pe_1_4_5_n29) );
  INV_X1 pe_1_4_5_U58 ( .A(pe_1_4_5_n29), .ZN(pe_1_4_5_n75) );
  XNOR2_X1 pe_1_4_5_U57 ( .A(pe_1_4_5_n70), .B(int_data_res_4__5__0_), .ZN(
        pe_1_4_5_N70) );
  AOI222_X1 pe_1_4_5_U52 ( .A1(int_data_res_5__5__0_), .A2(pe_1_4_5_n62), .B1(
        pe_1_4_5_n1), .B2(pe_1_4_5_n27), .C1(pe_1_4_5_N70), .C2(pe_1_4_5_n28), 
        .ZN(pe_1_4_5_n35) );
  INV_X1 pe_1_4_5_U51 ( .A(pe_1_4_5_n35), .ZN(pe_1_4_5_n81) );
  AOI222_X1 pe_1_4_5_U50 ( .A1(int_data_res_5__5__1_), .A2(pe_1_4_5_n62), .B1(
        pe_1_4_5_N79), .B2(pe_1_4_5_n27), .C1(pe_1_4_5_N71), .C2(pe_1_4_5_n28), 
        .ZN(pe_1_4_5_n34) );
  INV_X1 pe_1_4_5_U49 ( .A(pe_1_4_5_n34), .ZN(pe_1_4_5_n80) );
  AOI222_X1 pe_1_4_5_U48 ( .A1(int_data_res_5__5__3_), .A2(pe_1_4_5_n62), .B1(
        pe_1_4_5_N81), .B2(pe_1_4_5_n27), .C1(pe_1_4_5_N73), .C2(pe_1_4_5_n28), 
        .ZN(pe_1_4_5_n32) );
  INV_X1 pe_1_4_5_U47 ( .A(pe_1_4_5_n32), .ZN(pe_1_4_5_n78) );
  AOI222_X1 pe_1_4_5_U46 ( .A1(int_data_res_5__5__4_), .A2(pe_1_4_5_n62), .B1(
        pe_1_4_5_N82), .B2(pe_1_4_5_n27), .C1(pe_1_4_5_N74), .C2(pe_1_4_5_n28), 
        .ZN(pe_1_4_5_n31) );
  INV_X1 pe_1_4_5_U45 ( .A(pe_1_4_5_n31), .ZN(pe_1_4_5_n77) );
  AOI222_X1 pe_1_4_5_U44 ( .A1(int_data_res_5__5__5_), .A2(pe_1_4_5_n62), .B1(
        pe_1_4_5_N83), .B2(pe_1_4_5_n27), .C1(pe_1_4_5_N75), .C2(pe_1_4_5_n28), 
        .ZN(pe_1_4_5_n30) );
  INV_X1 pe_1_4_5_U43 ( .A(pe_1_4_5_n30), .ZN(pe_1_4_5_n76) );
  NAND2_X1 pe_1_4_5_U42 ( .A1(pe_1_4_5_int_data_0_), .A2(pe_1_4_5_n3), .ZN(
        pe_1_4_5_sub_81_carry[1]) );
  INV_X1 pe_1_4_5_U41 ( .A(pe_1_4_5_int_data_1_), .ZN(pe_1_4_5_n71) );
  INV_X1 pe_1_4_5_U40 ( .A(pe_1_4_5_int_data_2_), .ZN(pe_1_4_5_n72) );
  AND2_X1 pe_1_4_5_U39 ( .A1(pe_1_4_5_int_data_0_), .A2(int_data_res_4__5__0_), 
        .ZN(pe_1_4_5_n2) );
  AOI222_X1 pe_1_4_5_U38 ( .A1(pe_1_4_5_n62), .A2(int_data_res_5__5__7_), .B1(
        pe_1_4_5_N85), .B2(pe_1_4_5_n27), .C1(pe_1_4_5_N77), .C2(pe_1_4_5_n28), 
        .ZN(pe_1_4_5_n26) );
  INV_X1 pe_1_4_5_U37 ( .A(pe_1_4_5_n26), .ZN(pe_1_4_5_n74) );
  NOR3_X1 pe_1_4_5_U36 ( .A1(pe_1_4_5_n58), .A2(pe_1_4_5_n63), .A3(int_ckg[26]), .ZN(pe_1_4_5_n36) );
  OR2_X1 pe_1_4_5_U35 ( .A1(pe_1_4_5_n36), .A2(pe_1_4_5_n62), .ZN(pe_1_4_5_N90) );
  INV_X1 pe_1_4_5_U34 ( .A(n40), .ZN(pe_1_4_5_n61) );
  AND2_X1 pe_1_4_5_U33 ( .A1(int_data_x_4__5__2_), .A2(n28), .ZN(
        pe_1_4_5_int_data_2_) );
  AND2_X1 pe_1_4_5_U32 ( .A1(int_data_x_4__5__1_), .A2(n28), .ZN(
        pe_1_4_5_int_data_1_) );
  AND2_X1 pe_1_4_5_U31 ( .A1(int_data_x_4__5__3_), .A2(n28), .ZN(
        pe_1_4_5_int_data_3_) );
  BUF_X1 pe_1_4_5_U30 ( .A(n62), .Z(pe_1_4_5_n62) );
  INV_X1 pe_1_4_5_U29 ( .A(n34), .ZN(pe_1_4_5_n59) );
  AND2_X1 pe_1_4_5_U28 ( .A1(int_data_x_4__5__0_), .A2(n28), .ZN(
        pe_1_4_5_int_data_0_) );
  NAND2_X1 pe_1_4_5_U27 ( .A1(pe_1_4_5_n44), .A2(pe_1_4_5_n59), .ZN(
        pe_1_4_5_n41) );
  AND3_X1 pe_1_4_5_U26 ( .A1(n76), .A2(pe_1_4_5_n61), .A3(n50), .ZN(
        pe_1_4_5_n44) );
  INV_X1 pe_1_4_5_U25 ( .A(pe_1_4_5_int_data_3_), .ZN(pe_1_4_5_n73) );
  NOR2_X1 pe_1_4_5_U24 ( .A1(pe_1_4_5_n67), .A2(n50), .ZN(pe_1_4_5_n43) );
  NOR2_X1 pe_1_4_5_U23 ( .A1(pe_1_4_5_n57), .A2(pe_1_4_5_n62), .ZN(
        pe_1_4_5_n28) );
  NOR2_X1 pe_1_4_5_U22 ( .A1(n20), .A2(pe_1_4_5_n62), .ZN(pe_1_4_5_n27) );
  INV_X1 pe_1_4_5_U21 ( .A(pe_1_4_5_int_data_0_), .ZN(pe_1_4_5_n70) );
  INV_X1 pe_1_4_5_U20 ( .A(pe_1_4_5_n41), .ZN(pe_1_4_5_n87) );
  INV_X1 pe_1_4_5_U19 ( .A(pe_1_4_5_n37), .ZN(pe_1_4_5_n85) );
  INV_X1 pe_1_4_5_U18 ( .A(pe_1_4_5_n38), .ZN(pe_1_4_5_n84) );
  INV_X1 pe_1_4_5_U17 ( .A(pe_1_4_5_n39), .ZN(pe_1_4_5_n83) );
  NOR2_X1 pe_1_4_5_U16 ( .A1(pe_1_4_5_n65), .A2(pe_1_4_5_n42), .ZN(
        pe_1_4_5_N59) );
  NOR2_X1 pe_1_4_5_U15 ( .A1(pe_1_4_5_n65), .A2(pe_1_4_5_n41), .ZN(
        pe_1_4_5_N60) );
  NOR2_X1 pe_1_4_5_U14 ( .A1(pe_1_4_5_n65), .A2(pe_1_4_5_n38), .ZN(
        pe_1_4_5_N63) );
  NOR2_X1 pe_1_4_5_U13 ( .A1(pe_1_4_5_n65), .A2(pe_1_4_5_n40), .ZN(
        pe_1_4_5_N61) );
  NOR2_X1 pe_1_4_5_U12 ( .A1(pe_1_4_5_n65), .A2(pe_1_4_5_n39), .ZN(
        pe_1_4_5_N62) );
  NOR2_X1 pe_1_4_5_U11 ( .A1(pe_1_4_5_n37), .A2(pe_1_4_5_n65), .ZN(
        pe_1_4_5_N64) );
  NAND2_X1 pe_1_4_5_U10 ( .A1(pe_1_4_5_n44), .A2(n34), .ZN(pe_1_4_5_n42) );
  BUF_X1 pe_1_4_5_U9 ( .A(n34), .Z(pe_1_4_5_n55) );
  INV_X1 pe_1_4_5_U8 ( .A(pe_1_4_5_n66), .ZN(pe_1_4_5_n63) );
  BUF_X1 pe_1_4_5_U7 ( .A(n34), .Z(pe_1_4_5_n56) );
  INV_X1 pe_1_4_5_U6 ( .A(pe_1_4_5_n42), .ZN(pe_1_4_5_n86) );
  INV_X1 pe_1_4_5_U5 ( .A(pe_1_4_5_n40), .ZN(pe_1_4_5_n82) );
  INV_X2 pe_1_4_5_U4 ( .A(n84), .ZN(pe_1_4_5_n69) );
  XOR2_X1 pe_1_4_5_U3 ( .A(pe_1_4_5_int_data_0_), .B(int_data_res_4__5__0_), 
        .Z(pe_1_4_5_n1) );
  DFFR_X1 pe_1_4_5_int_q_acc_reg_0_ ( .D(pe_1_4_5_n81), .CK(pe_1_4_5_net4666), 
        .RN(pe_1_4_5_n69), .Q(int_data_res_4__5__0_), .QN(pe_1_4_5_n3) );
  DFFR_X1 pe_1_4_5_int_q_reg_v_reg_0__0_ ( .D(int_data_y_5__5__0_), .CK(
        pe_1_4_5_net4636), .RN(pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_v[20]) );
  DFFR_X1 pe_1_4_5_int_q_reg_v_reg_0__1_ ( .D(int_data_y_5__5__1_), .CK(
        pe_1_4_5_net4636), .RN(pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_v[21]) );
  DFFR_X1 pe_1_4_5_int_q_reg_v_reg_0__2_ ( .D(int_data_y_5__5__2_), .CK(
        pe_1_4_5_net4636), .RN(pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_v[22]) );
  DFFR_X1 pe_1_4_5_int_q_reg_v_reg_0__3_ ( .D(int_data_y_5__5__3_), .CK(
        pe_1_4_5_net4636), .RN(pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_v[23]) );
  DFFR_X1 pe_1_4_5_int_q_reg_v_reg_1__0_ ( .D(int_data_y_5__5__0_), .CK(
        pe_1_4_5_net4641), .RN(pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_v[16]) );
  DFFR_X1 pe_1_4_5_int_q_reg_v_reg_1__1_ ( .D(int_data_y_5__5__1_), .CK(
        pe_1_4_5_net4641), .RN(pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_v[17]) );
  DFFR_X1 pe_1_4_5_int_q_reg_v_reg_1__2_ ( .D(int_data_y_5__5__2_), .CK(
        pe_1_4_5_net4641), .RN(pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_v[18]) );
  DFFR_X1 pe_1_4_5_int_q_reg_v_reg_1__3_ ( .D(int_data_y_5__5__3_), .CK(
        pe_1_4_5_net4641), .RN(pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_v[19]) );
  DFFR_X1 pe_1_4_5_int_q_reg_v_reg_2__0_ ( .D(int_data_y_5__5__0_), .CK(
        pe_1_4_5_net4646), .RN(pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_v[12]) );
  DFFR_X1 pe_1_4_5_int_q_reg_v_reg_2__1_ ( .D(int_data_y_5__5__1_), .CK(
        pe_1_4_5_net4646), .RN(pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_v[13]) );
  DFFR_X1 pe_1_4_5_int_q_reg_v_reg_2__2_ ( .D(int_data_y_5__5__2_), .CK(
        pe_1_4_5_net4646), .RN(pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_v[14]) );
  DFFR_X1 pe_1_4_5_int_q_reg_v_reg_2__3_ ( .D(int_data_y_5__5__3_), .CK(
        pe_1_4_5_net4646), .RN(pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_v[15]) );
  DFFR_X1 pe_1_4_5_int_q_reg_v_reg_3__0_ ( .D(int_data_y_5__5__0_), .CK(
        pe_1_4_5_net4651), .RN(pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_v[8]) );
  DFFR_X1 pe_1_4_5_int_q_reg_v_reg_3__1_ ( .D(int_data_y_5__5__1_), .CK(
        pe_1_4_5_net4651), .RN(pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_v[9]) );
  DFFR_X1 pe_1_4_5_int_q_reg_v_reg_3__2_ ( .D(int_data_y_5__5__2_), .CK(
        pe_1_4_5_net4651), .RN(pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_v[10]) );
  DFFR_X1 pe_1_4_5_int_q_reg_v_reg_3__3_ ( .D(int_data_y_5__5__3_), .CK(
        pe_1_4_5_net4651), .RN(pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_v[11]) );
  DFFR_X1 pe_1_4_5_int_q_reg_v_reg_4__0_ ( .D(int_data_y_5__5__0_), .CK(
        pe_1_4_5_net4656), .RN(pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_v[4]) );
  DFFR_X1 pe_1_4_5_int_q_reg_v_reg_4__1_ ( .D(int_data_y_5__5__1_), .CK(
        pe_1_4_5_net4656), .RN(pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_v[5]) );
  DFFR_X1 pe_1_4_5_int_q_reg_v_reg_4__2_ ( .D(int_data_y_5__5__2_), .CK(
        pe_1_4_5_net4656), .RN(pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_v[6]) );
  DFFR_X1 pe_1_4_5_int_q_reg_v_reg_4__3_ ( .D(int_data_y_5__5__3_), .CK(
        pe_1_4_5_net4656), .RN(pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_v[7]) );
  DFFR_X1 pe_1_4_5_int_q_reg_v_reg_5__0_ ( .D(int_data_y_5__5__0_), .CK(
        pe_1_4_5_net4661), .RN(pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_v[0]) );
  DFFR_X1 pe_1_4_5_int_q_reg_v_reg_5__1_ ( .D(int_data_y_5__5__1_), .CK(
        pe_1_4_5_net4661), .RN(pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_v[1]) );
  DFFR_X1 pe_1_4_5_int_q_reg_v_reg_5__2_ ( .D(int_data_y_5__5__2_), .CK(
        pe_1_4_5_net4661), .RN(pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_v[2]) );
  DFFR_X1 pe_1_4_5_int_q_reg_v_reg_5__3_ ( .D(int_data_y_5__5__3_), .CK(
        pe_1_4_5_net4661), .RN(pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_4_5_int_q_reg_h_reg_0__0_ ( .D(int_data_x_4__6__0_), .SI(
        int_data_y_5__5__0_), .SE(pe_1_4_5_n63), .CK(pe_1_4_5_net4605), .RN(
        pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_4_5_int_q_reg_h_reg_0__1_ ( .D(int_data_x_4__6__1_), .SI(
        int_data_y_5__5__1_), .SE(pe_1_4_5_n63), .CK(pe_1_4_5_net4605), .RN(
        pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_4_5_int_q_reg_h_reg_0__2_ ( .D(int_data_x_4__6__2_), .SI(
        int_data_y_5__5__2_), .SE(pe_1_4_5_n63), .CK(pe_1_4_5_net4605), .RN(
        pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_4_5_int_q_reg_h_reg_0__3_ ( .D(int_data_x_4__6__3_), .SI(
        int_data_y_5__5__3_), .SE(pe_1_4_5_n63), .CK(pe_1_4_5_net4605), .RN(
        pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_4_5_int_q_reg_h_reg_1__0_ ( .D(int_data_x_4__6__0_), .SI(
        int_data_y_5__5__0_), .SE(pe_1_4_5_n63), .CK(pe_1_4_5_net4611), .RN(
        pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_4_5_int_q_reg_h_reg_1__1_ ( .D(int_data_x_4__6__1_), .SI(
        int_data_y_5__5__1_), .SE(pe_1_4_5_n63), .CK(pe_1_4_5_net4611), .RN(
        pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_4_5_int_q_reg_h_reg_1__2_ ( .D(int_data_x_4__6__2_), .SI(
        int_data_y_5__5__2_), .SE(pe_1_4_5_n63), .CK(pe_1_4_5_net4611), .RN(
        pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_4_5_int_q_reg_h_reg_1__3_ ( .D(int_data_x_4__6__3_), .SI(
        int_data_y_5__5__3_), .SE(pe_1_4_5_n63), .CK(pe_1_4_5_net4611), .RN(
        pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_4_5_int_q_reg_h_reg_2__0_ ( .D(int_data_x_4__6__0_), .SI(
        int_data_y_5__5__0_), .SE(pe_1_4_5_n63), .CK(pe_1_4_5_net4616), .RN(
        pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_4_5_int_q_reg_h_reg_2__1_ ( .D(int_data_x_4__6__1_), .SI(
        int_data_y_5__5__1_), .SE(pe_1_4_5_n63), .CK(pe_1_4_5_net4616), .RN(
        pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_4_5_int_q_reg_h_reg_2__2_ ( .D(int_data_x_4__6__2_), .SI(
        int_data_y_5__5__2_), .SE(pe_1_4_5_n63), .CK(pe_1_4_5_net4616), .RN(
        pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_4_5_int_q_reg_h_reg_2__3_ ( .D(int_data_x_4__6__3_), .SI(
        int_data_y_5__5__3_), .SE(pe_1_4_5_n63), .CK(pe_1_4_5_net4616), .RN(
        pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_4_5_int_q_reg_h_reg_3__0_ ( .D(int_data_x_4__6__0_), .SI(
        int_data_y_5__5__0_), .SE(pe_1_4_5_n63), .CK(pe_1_4_5_net4621), .RN(
        pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_4_5_int_q_reg_h_reg_3__1_ ( .D(int_data_x_4__6__1_), .SI(
        int_data_y_5__5__1_), .SE(pe_1_4_5_n63), .CK(pe_1_4_5_net4621), .RN(
        pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_4_5_int_q_reg_h_reg_3__2_ ( .D(int_data_x_4__6__2_), .SI(
        int_data_y_5__5__2_), .SE(pe_1_4_5_n63), .CK(pe_1_4_5_net4621), .RN(
        pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_4_5_int_q_reg_h_reg_3__3_ ( .D(int_data_x_4__6__3_), .SI(
        int_data_y_5__5__3_), .SE(pe_1_4_5_n63), .CK(pe_1_4_5_net4621), .RN(
        pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_4_5_int_q_reg_h_reg_4__0_ ( .D(int_data_x_4__6__0_), .SI(
        int_data_y_5__5__0_), .SE(pe_1_4_5_n64), .CK(pe_1_4_5_net4626), .RN(
        pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_4_5_int_q_reg_h_reg_4__1_ ( .D(int_data_x_4__6__1_), .SI(
        int_data_y_5__5__1_), .SE(pe_1_4_5_n64), .CK(pe_1_4_5_net4626), .RN(
        pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_4_5_int_q_reg_h_reg_4__2_ ( .D(int_data_x_4__6__2_), .SI(
        int_data_y_5__5__2_), .SE(pe_1_4_5_n64), .CK(pe_1_4_5_net4626), .RN(
        pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_4_5_int_q_reg_h_reg_4__3_ ( .D(int_data_x_4__6__3_), .SI(
        int_data_y_5__5__3_), .SE(pe_1_4_5_n64), .CK(pe_1_4_5_net4626), .RN(
        pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_4_5_int_q_reg_h_reg_5__0_ ( .D(int_data_x_4__6__0_), .SI(
        int_data_y_5__5__0_), .SE(pe_1_4_5_n64), .CK(pe_1_4_5_net4631), .RN(
        pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_4_5_int_q_reg_h_reg_5__1_ ( .D(int_data_x_4__6__1_), .SI(
        int_data_y_5__5__1_), .SE(pe_1_4_5_n64), .CK(pe_1_4_5_net4631), .RN(
        pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_4_5_int_q_reg_h_reg_5__2_ ( .D(int_data_x_4__6__2_), .SI(
        int_data_y_5__5__2_), .SE(pe_1_4_5_n64), .CK(pe_1_4_5_net4631), .RN(
        pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_4_5_int_q_reg_h_reg_5__3_ ( .D(int_data_x_4__6__3_), .SI(
        int_data_y_5__5__3_), .SE(pe_1_4_5_n64), .CK(pe_1_4_5_net4631), .RN(
        pe_1_4_5_n69), .Q(pe_1_4_5_int_q_reg_h[3]) );
  FA_X1 pe_1_4_5_sub_81_U2_7 ( .A(int_data_res_4__5__7_), .B(pe_1_4_5_n73), 
        .CI(pe_1_4_5_sub_81_carry[7]), .S(pe_1_4_5_N77) );
  FA_X1 pe_1_4_5_sub_81_U2_6 ( .A(int_data_res_4__5__6_), .B(pe_1_4_5_n73), 
        .CI(pe_1_4_5_sub_81_carry[6]), .CO(pe_1_4_5_sub_81_carry[7]), .S(
        pe_1_4_5_N76) );
  FA_X1 pe_1_4_5_sub_81_U2_5 ( .A(int_data_res_4__5__5_), .B(pe_1_4_5_n73), 
        .CI(pe_1_4_5_sub_81_carry[5]), .CO(pe_1_4_5_sub_81_carry[6]), .S(
        pe_1_4_5_N75) );
  FA_X1 pe_1_4_5_sub_81_U2_4 ( .A(int_data_res_4__5__4_), .B(pe_1_4_5_n73), 
        .CI(pe_1_4_5_sub_81_carry[4]), .CO(pe_1_4_5_sub_81_carry[5]), .S(
        pe_1_4_5_N74) );
  FA_X1 pe_1_4_5_sub_81_U2_3 ( .A(int_data_res_4__5__3_), .B(pe_1_4_5_n73), 
        .CI(pe_1_4_5_sub_81_carry[3]), .CO(pe_1_4_5_sub_81_carry[4]), .S(
        pe_1_4_5_N73) );
  FA_X1 pe_1_4_5_sub_81_U2_2 ( .A(int_data_res_4__5__2_), .B(pe_1_4_5_n72), 
        .CI(pe_1_4_5_sub_81_carry[2]), .CO(pe_1_4_5_sub_81_carry[3]), .S(
        pe_1_4_5_N72) );
  FA_X1 pe_1_4_5_sub_81_U2_1 ( .A(int_data_res_4__5__1_), .B(pe_1_4_5_n71), 
        .CI(pe_1_4_5_sub_81_carry[1]), .CO(pe_1_4_5_sub_81_carry[2]), .S(
        pe_1_4_5_N71) );
  FA_X1 pe_1_4_5_add_83_U1_7 ( .A(int_data_res_4__5__7_), .B(
        pe_1_4_5_int_data_3_), .CI(pe_1_4_5_add_83_carry[7]), .S(pe_1_4_5_N85)
         );
  FA_X1 pe_1_4_5_add_83_U1_6 ( .A(int_data_res_4__5__6_), .B(
        pe_1_4_5_int_data_3_), .CI(pe_1_4_5_add_83_carry[6]), .CO(
        pe_1_4_5_add_83_carry[7]), .S(pe_1_4_5_N84) );
  FA_X1 pe_1_4_5_add_83_U1_5 ( .A(int_data_res_4__5__5_), .B(
        pe_1_4_5_int_data_3_), .CI(pe_1_4_5_add_83_carry[5]), .CO(
        pe_1_4_5_add_83_carry[6]), .S(pe_1_4_5_N83) );
  FA_X1 pe_1_4_5_add_83_U1_4 ( .A(int_data_res_4__5__4_), .B(
        pe_1_4_5_int_data_3_), .CI(pe_1_4_5_add_83_carry[4]), .CO(
        pe_1_4_5_add_83_carry[5]), .S(pe_1_4_5_N82) );
  FA_X1 pe_1_4_5_add_83_U1_3 ( .A(int_data_res_4__5__3_), .B(
        pe_1_4_5_int_data_3_), .CI(pe_1_4_5_add_83_carry[3]), .CO(
        pe_1_4_5_add_83_carry[4]), .S(pe_1_4_5_N81) );
  FA_X1 pe_1_4_5_add_83_U1_2 ( .A(int_data_res_4__5__2_), .B(
        pe_1_4_5_int_data_2_), .CI(pe_1_4_5_add_83_carry[2]), .CO(
        pe_1_4_5_add_83_carry[3]), .S(pe_1_4_5_N80) );
  FA_X1 pe_1_4_5_add_83_U1_1 ( .A(int_data_res_4__5__1_), .B(
        pe_1_4_5_int_data_1_), .CI(pe_1_4_5_n2), .CO(pe_1_4_5_add_83_carry[2]), 
        .S(pe_1_4_5_N79) );
  NAND3_X1 pe_1_4_5_U56 ( .A1(n34), .A2(pe_1_4_5_n43), .A3(pe_1_4_5_n60), .ZN(
        pe_1_4_5_n40) );
  NAND3_X1 pe_1_4_5_U55 ( .A1(pe_1_4_5_n43), .A2(pe_1_4_5_n59), .A3(
        pe_1_4_5_n60), .ZN(pe_1_4_5_n39) );
  NAND3_X1 pe_1_4_5_U54 ( .A1(pe_1_4_5_n43), .A2(pe_1_4_5_n61), .A3(n34), .ZN(
        pe_1_4_5_n38) );
  NAND3_X1 pe_1_4_5_U53 ( .A1(pe_1_4_5_n59), .A2(pe_1_4_5_n61), .A3(
        pe_1_4_5_n43), .ZN(pe_1_4_5_n37) );
  DFFR_X1 pe_1_4_5_int_q_acc_reg_6_ ( .D(pe_1_4_5_n75), .CK(pe_1_4_5_net4666), 
        .RN(pe_1_4_5_n68), .Q(int_data_res_4__5__6_) );
  DFFR_X1 pe_1_4_5_int_q_acc_reg_5_ ( .D(pe_1_4_5_n76), .CK(pe_1_4_5_net4666), 
        .RN(pe_1_4_5_n68), .Q(int_data_res_4__5__5_) );
  DFFR_X1 pe_1_4_5_int_q_acc_reg_4_ ( .D(pe_1_4_5_n77), .CK(pe_1_4_5_net4666), 
        .RN(pe_1_4_5_n68), .Q(int_data_res_4__5__4_) );
  DFFR_X1 pe_1_4_5_int_q_acc_reg_3_ ( .D(pe_1_4_5_n78), .CK(pe_1_4_5_net4666), 
        .RN(pe_1_4_5_n68), .Q(int_data_res_4__5__3_) );
  DFFR_X1 pe_1_4_5_int_q_acc_reg_2_ ( .D(pe_1_4_5_n79), .CK(pe_1_4_5_net4666), 
        .RN(pe_1_4_5_n68), .Q(int_data_res_4__5__2_) );
  DFFR_X1 pe_1_4_5_int_q_acc_reg_1_ ( .D(pe_1_4_5_n80), .CK(pe_1_4_5_net4666), 
        .RN(pe_1_4_5_n68), .Q(int_data_res_4__5__1_) );
  DFFR_X1 pe_1_4_5_int_q_acc_reg_7_ ( .D(pe_1_4_5_n74), .CK(pe_1_4_5_net4666), 
        .RN(pe_1_4_5_n68), .Q(int_data_res_4__5__7_) );
  CLKGATETST_X1 pe_1_4_5_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_4_5_n85), .SE(1'b0), .GCK(pe_1_4_5_net4605) );
  CLKGATETST_X1 pe_1_4_5_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_4_5_n84), .SE(1'b0), .GCK(pe_1_4_5_net4611) );
  CLKGATETST_X1 pe_1_4_5_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_4_5_n83), .SE(1'b0), .GCK(pe_1_4_5_net4616) );
  CLKGATETST_X1 pe_1_4_5_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_4_5_n82), .SE(1'b0), .GCK(pe_1_4_5_net4621) );
  CLKGATETST_X1 pe_1_4_5_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_4_5_n87), .SE(1'b0), .GCK(pe_1_4_5_net4626) );
  CLKGATETST_X1 pe_1_4_5_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_4_5_n86), .SE(1'b0), .GCK(pe_1_4_5_net4631) );
  CLKGATETST_X1 pe_1_4_5_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_4_5_N64), .SE(1'b0), .GCK(pe_1_4_5_net4636) );
  CLKGATETST_X1 pe_1_4_5_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_4_5_N63), .SE(1'b0), .GCK(pe_1_4_5_net4641) );
  CLKGATETST_X1 pe_1_4_5_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_4_5_N62), .SE(1'b0), .GCK(pe_1_4_5_net4646) );
  CLKGATETST_X1 pe_1_4_5_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_4_5_N61), .SE(1'b0), .GCK(pe_1_4_5_net4651) );
  CLKGATETST_X1 pe_1_4_5_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_4_5_N60), .SE(1'b0), .GCK(pe_1_4_5_net4656) );
  CLKGATETST_X1 pe_1_4_5_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_4_5_N59), .SE(1'b0), .GCK(pe_1_4_5_net4661) );
  CLKGATETST_X1 pe_1_4_5_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_4_5_N90), .SE(1'b0), .GCK(pe_1_4_5_net4666) );
  CLKBUF_X1 pe_1_4_6_U110 ( .A(pe_1_4_6_n70), .Z(pe_1_4_6_n69) );
  INV_X1 pe_1_4_6_U109 ( .A(n76), .ZN(pe_1_4_6_n68) );
  INV_X1 pe_1_4_6_U108 ( .A(n68), .ZN(pe_1_4_6_n67) );
  INV_X1 pe_1_4_6_U107 ( .A(n68), .ZN(pe_1_4_6_n66) );
  INV_X1 pe_1_4_6_U106 ( .A(pe_1_4_6_n67), .ZN(pe_1_4_6_n65) );
  INV_X1 pe_1_4_6_U105 ( .A(pe_1_4_6_n62), .ZN(pe_1_4_6_n61) );
  INV_X1 pe_1_4_6_U104 ( .A(pe_1_4_6_n60), .ZN(pe_1_4_6_n59) );
  INV_X1 pe_1_4_6_U103 ( .A(n28), .ZN(pe_1_4_6_n58) );
  INV_X1 pe_1_4_6_U102 ( .A(n20), .ZN(pe_1_4_6_n57) );
  MUX2_X1 pe_1_4_6_U101 ( .A(pe_1_4_6_n54), .B(pe_1_4_6_n51), .S(n50), .Z(
        int_data_x_4__6__3_) );
  MUX2_X1 pe_1_4_6_U100 ( .A(pe_1_4_6_n53), .B(pe_1_4_6_n52), .S(pe_1_4_6_n61), 
        .Z(pe_1_4_6_n54) );
  MUX2_X1 pe_1_4_6_U99 ( .A(pe_1_4_6_int_q_reg_h[23]), .B(
        pe_1_4_6_int_q_reg_h[19]), .S(pe_1_4_6_n56), .Z(pe_1_4_6_n53) );
  MUX2_X1 pe_1_4_6_U98 ( .A(pe_1_4_6_int_q_reg_h[15]), .B(
        pe_1_4_6_int_q_reg_h[11]), .S(pe_1_4_6_n56), .Z(pe_1_4_6_n52) );
  MUX2_X1 pe_1_4_6_U97 ( .A(pe_1_4_6_int_q_reg_h[7]), .B(
        pe_1_4_6_int_q_reg_h[3]), .S(pe_1_4_6_n56), .Z(pe_1_4_6_n51) );
  MUX2_X1 pe_1_4_6_U96 ( .A(pe_1_4_6_n50), .B(pe_1_4_6_n47), .S(n50), .Z(
        int_data_x_4__6__2_) );
  MUX2_X1 pe_1_4_6_U95 ( .A(pe_1_4_6_n49), .B(pe_1_4_6_n48), .S(pe_1_4_6_n61), 
        .Z(pe_1_4_6_n50) );
  MUX2_X1 pe_1_4_6_U94 ( .A(pe_1_4_6_int_q_reg_h[22]), .B(
        pe_1_4_6_int_q_reg_h[18]), .S(pe_1_4_6_n56), .Z(pe_1_4_6_n49) );
  MUX2_X1 pe_1_4_6_U93 ( .A(pe_1_4_6_int_q_reg_h[14]), .B(
        pe_1_4_6_int_q_reg_h[10]), .S(pe_1_4_6_n56), .Z(pe_1_4_6_n48) );
  MUX2_X1 pe_1_4_6_U92 ( .A(pe_1_4_6_int_q_reg_h[6]), .B(
        pe_1_4_6_int_q_reg_h[2]), .S(pe_1_4_6_n56), .Z(pe_1_4_6_n47) );
  MUX2_X1 pe_1_4_6_U91 ( .A(pe_1_4_6_n46), .B(pe_1_4_6_n24), .S(n50), .Z(
        int_data_x_4__6__1_) );
  MUX2_X1 pe_1_4_6_U90 ( .A(pe_1_4_6_n45), .B(pe_1_4_6_n25), .S(pe_1_4_6_n61), 
        .Z(pe_1_4_6_n46) );
  MUX2_X1 pe_1_4_6_U89 ( .A(pe_1_4_6_int_q_reg_h[21]), .B(
        pe_1_4_6_int_q_reg_h[17]), .S(pe_1_4_6_n56), .Z(pe_1_4_6_n45) );
  MUX2_X1 pe_1_4_6_U88 ( .A(pe_1_4_6_int_q_reg_h[13]), .B(
        pe_1_4_6_int_q_reg_h[9]), .S(pe_1_4_6_n56), .Z(pe_1_4_6_n25) );
  MUX2_X1 pe_1_4_6_U87 ( .A(pe_1_4_6_int_q_reg_h[5]), .B(
        pe_1_4_6_int_q_reg_h[1]), .S(pe_1_4_6_n56), .Z(pe_1_4_6_n24) );
  MUX2_X1 pe_1_4_6_U86 ( .A(pe_1_4_6_n23), .B(pe_1_4_6_n20), .S(n50), .Z(
        int_data_x_4__6__0_) );
  MUX2_X1 pe_1_4_6_U85 ( .A(pe_1_4_6_n22), .B(pe_1_4_6_n21), .S(pe_1_4_6_n61), 
        .Z(pe_1_4_6_n23) );
  MUX2_X1 pe_1_4_6_U84 ( .A(pe_1_4_6_int_q_reg_h[20]), .B(
        pe_1_4_6_int_q_reg_h[16]), .S(pe_1_4_6_n56), .Z(pe_1_4_6_n22) );
  MUX2_X1 pe_1_4_6_U83 ( .A(pe_1_4_6_int_q_reg_h[12]), .B(
        pe_1_4_6_int_q_reg_h[8]), .S(pe_1_4_6_n56), .Z(pe_1_4_6_n21) );
  MUX2_X1 pe_1_4_6_U82 ( .A(pe_1_4_6_int_q_reg_h[4]), .B(
        pe_1_4_6_int_q_reg_h[0]), .S(pe_1_4_6_n56), .Z(pe_1_4_6_n20) );
  MUX2_X1 pe_1_4_6_U81 ( .A(pe_1_4_6_n19), .B(pe_1_4_6_n16), .S(n50), .Z(
        int_data_y_4__6__3_) );
  MUX2_X1 pe_1_4_6_U80 ( .A(pe_1_4_6_n18), .B(pe_1_4_6_n17), .S(pe_1_4_6_n61), 
        .Z(pe_1_4_6_n19) );
  MUX2_X1 pe_1_4_6_U79 ( .A(pe_1_4_6_int_q_reg_v[23]), .B(
        pe_1_4_6_int_q_reg_v[19]), .S(pe_1_4_6_n55), .Z(pe_1_4_6_n18) );
  MUX2_X1 pe_1_4_6_U78 ( .A(pe_1_4_6_int_q_reg_v[15]), .B(
        pe_1_4_6_int_q_reg_v[11]), .S(pe_1_4_6_n55), .Z(pe_1_4_6_n17) );
  MUX2_X1 pe_1_4_6_U77 ( .A(pe_1_4_6_int_q_reg_v[7]), .B(
        pe_1_4_6_int_q_reg_v[3]), .S(pe_1_4_6_n55), .Z(pe_1_4_6_n16) );
  MUX2_X1 pe_1_4_6_U76 ( .A(pe_1_4_6_n15), .B(pe_1_4_6_n12), .S(n50), .Z(
        int_data_y_4__6__2_) );
  MUX2_X1 pe_1_4_6_U75 ( .A(pe_1_4_6_n14), .B(pe_1_4_6_n13), .S(pe_1_4_6_n61), 
        .Z(pe_1_4_6_n15) );
  MUX2_X1 pe_1_4_6_U74 ( .A(pe_1_4_6_int_q_reg_v[22]), .B(
        pe_1_4_6_int_q_reg_v[18]), .S(pe_1_4_6_n55), .Z(pe_1_4_6_n14) );
  MUX2_X1 pe_1_4_6_U73 ( .A(pe_1_4_6_int_q_reg_v[14]), .B(
        pe_1_4_6_int_q_reg_v[10]), .S(pe_1_4_6_n55), .Z(pe_1_4_6_n13) );
  MUX2_X1 pe_1_4_6_U72 ( .A(pe_1_4_6_int_q_reg_v[6]), .B(
        pe_1_4_6_int_q_reg_v[2]), .S(pe_1_4_6_n55), .Z(pe_1_4_6_n12) );
  MUX2_X1 pe_1_4_6_U71 ( .A(pe_1_4_6_n11), .B(pe_1_4_6_n8), .S(n50), .Z(
        int_data_y_4__6__1_) );
  MUX2_X1 pe_1_4_6_U70 ( .A(pe_1_4_6_n10), .B(pe_1_4_6_n9), .S(pe_1_4_6_n61), 
        .Z(pe_1_4_6_n11) );
  MUX2_X1 pe_1_4_6_U69 ( .A(pe_1_4_6_int_q_reg_v[21]), .B(
        pe_1_4_6_int_q_reg_v[17]), .S(pe_1_4_6_n55), .Z(pe_1_4_6_n10) );
  MUX2_X1 pe_1_4_6_U68 ( .A(pe_1_4_6_int_q_reg_v[13]), .B(
        pe_1_4_6_int_q_reg_v[9]), .S(pe_1_4_6_n55), .Z(pe_1_4_6_n9) );
  MUX2_X1 pe_1_4_6_U67 ( .A(pe_1_4_6_int_q_reg_v[5]), .B(
        pe_1_4_6_int_q_reg_v[1]), .S(pe_1_4_6_n55), .Z(pe_1_4_6_n8) );
  MUX2_X1 pe_1_4_6_U66 ( .A(pe_1_4_6_n7), .B(pe_1_4_6_n4), .S(n50), .Z(
        int_data_y_4__6__0_) );
  MUX2_X1 pe_1_4_6_U65 ( .A(pe_1_4_6_n6), .B(pe_1_4_6_n5), .S(pe_1_4_6_n61), 
        .Z(pe_1_4_6_n7) );
  MUX2_X1 pe_1_4_6_U64 ( .A(pe_1_4_6_int_q_reg_v[20]), .B(
        pe_1_4_6_int_q_reg_v[16]), .S(pe_1_4_6_n55), .Z(pe_1_4_6_n6) );
  MUX2_X1 pe_1_4_6_U63 ( .A(pe_1_4_6_int_q_reg_v[12]), .B(
        pe_1_4_6_int_q_reg_v[8]), .S(pe_1_4_6_n55), .Z(pe_1_4_6_n5) );
  MUX2_X1 pe_1_4_6_U62 ( .A(pe_1_4_6_int_q_reg_v[4]), .B(
        pe_1_4_6_int_q_reg_v[0]), .S(pe_1_4_6_n55), .Z(pe_1_4_6_n4) );
  AOI222_X1 pe_1_4_6_U61 ( .A1(int_data_res_5__6__2_), .A2(pe_1_4_6_n63), .B1(
        pe_1_4_6_N80), .B2(pe_1_4_6_n27), .C1(pe_1_4_6_N72), .C2(pe_1_4_6_n28), 
        .ZN(pe_1_4_6_n33) );
  INV_X1 pe_1_4_6_U60 ( .A(pe_1_4_6_n33), .ZN(pe_1_4_6_n80) );
  AOI222_X1 pe_1_4_6_U59 ( .A1(int_data_res_5__6__6_), .A2(pe_1_4_6_n63), .B1(
        pe_1_4_6_N84), .B2(pe_1_4_6_n27), .C1(pe_1_4_6_N76), .C2(pe_1_4_6_n28), 
        .ZN(pe_1_4_6_n29) );
  INV_X1 pe_1_4_6_U58 ( .A(pe_1_4_6_n29), .ZN(pe_1_4_6_n76) );
  XNOR2_X1 pe_1_4_6_U57 ( .A(pe_1_4_6_n71), .B(int_data_res_4__6__0_), .ZN(
        pe_1_4_6_N70) );
  AOI222_X1 pe_1_4_6_U52 ( .A1(int_data_res_5__6__0_), .A2(pe_1_4_6_n63), .B1(
        pe_1_4_6_n1), .B2(pe_1_4_6_n27), .C1(pe_1_4_6_N70), .C2(pe_1_4_6_n28), 
        .ZN(pe_1_4_6_n35) );
  INV_X1 pe_1_4_6_U51 ( .A(pe_1_4_6_n35), .ZN(pe_1_4_6_n82) );
  AOI222_X1 pe_1_4_6_U50 ( .A1(int_data_res_5__6__1_), .A2(pe_1_4_6_n63), .B1(
        pe_1_4_6_N79), .B2(pe_1_4_6_n27), .C1(pe_1_4_6_N71), .C2(pe_1_4_6_n28), 
        .ZN(pe_1_4_6_n34) );
  INV_X1 pe_1_4_6_U49 ( .A(pe_1_4_6_n34), .ZN(pe_1_4_6_n81) );
  AOI222_X1 pe_1_4_6_U48 ( .A1(int_data_res_5__6__3_), .A2(pe_1_4_6_n63), .B1(
        pe_1_4_6_N81), .B2(pe_1_4_6_n27), .C1(pe_1_4_6_N73), .C2(pe_1_4_6_n28), 
        .ZN(pe_1_4_6_n32) );
  INV_X1 pe_1_4_6_U47 ( .A(pe_1_4_6_n32), .ZN(pe_1_4_6_n79) );
  AOI222_X1 pe_1_4_6_U46 ( .A1(int_data_res_5__6__4_), .A2(pe_1_4_6_n63), .B1(
        pe_1_4_6_N82), .B2(pe_1_4_6_n27), .C1(pe_1_4_6_N74), .C2(pe_1_4_6_n28), 
        .ZN(pe_1_4_6_n31) );
  INV_X1 pe_1_4_6_U45 ( .A(pe_1_4_6_n31), .ZN(pe_1_4_6_n78) );
  AOI222_X1 pe_1_4_6_U44 ( .A1(int_data_res_5__6__5_), .A2(pe_1_4_6_n63), .B1(
        pe_1_4_6_N83), .B2(pe_1_4_6_n27), .C1(pe_1_4_6_N75), .C2(pe_1_4_6_n28), 
        .ZN(pe_1_4_6_n30) );
  INV_X1 pe_1_4_6_U43 ( .A(pe_1_4_6_n30), .ZN(pe_1_4_6_n77) );
  NAND2_X1 pe_1_4_6_U42 ( .A1(pe_1_4_6_int_data_0_), .A2(pe_1_4_6_n3), .ZN(
        pe_1_4_6_sub_81_carry[1]) );
  INV_X1 pe_1_4_6_U41 ( .A(pe_1_4_6_int_data_1_), .ZN(pe_1_4_6_n72) );
  INV_X1 pe_1_4_6_U40 ( .A(pe_1_4_6_int_data_2_), .ZN(pe_1_4_6_n73) );
  AND2_X1 pe_1_4_6_U39 ( .A1(pe_1_4_6_int_data_0_), .A2(int_data_res_4__6__0_), 
        .ZN(pe_1_4_6_n2) );
  AOI222_X1 pe_1_4_6_U38 ( .A1(pe_1_4_6_n63), .A2(int_data_res_5__6__7_), .B1(
        pe_1_4_6_N85), .B2(pe_1_4_6_n27), .C1(pe_1_4_6_N77), .C2(pe_1_4_6_n28), 
        .ZN(pe_1_4_6_n26) );
  INV_X1 pe_1_4_6_U37 ( .A(pe_1_4_6_n26), .ZN(pe_1_4_6_n75) );
  NOR3_X1 pe_1_4_6_U36 ( .A1(pe_1_4_6_n58), .A2(pe_1_4_6_n64), .A3(int_ckg[25]), .ZN(pe_1_4_6_n36) );
  OR2_X1 pe_1_4_6_U35 ( .A1(pe_1_4_6_n36), .A2(pe_1_4_6_n63), .ZN(pe_1_4_6_N90) );
  INV_X1 pe_1_4_6_U34 ( .A(n40), .ZN(pe_1_4_6_n62) );
  AND2_X1 pe_1_4_6_U33 ( .A1(int_data_x_4__6__2_), .A2(n28), .ZN(
        pe_1_4_6_int_data_2_) );
  AND2_X1 pe_1_4_6_U32 ( .A1(int_data_x_4__6__1_), .A2(n28), .ZN(
        pe_1_4_6_int_data_1_) );
  AND2_X1 pe_1_4_6_U31 ( .A1(int_data_x_4__6__3_), .A2(n28), .ZN(
        pe_1_4_6_int_data_3_) );
  BUF_X1 pe_1_4_6_U30 ( .A(n62), .Z(pe_1_4_6_n63) );
  INV_X1 pe_1_4_6_U29 ( .A(n34), .ZN(pe_1_4_6_n60) );
  AND2_X1 pe_1_4_6_U28 ( .A1(int_data_x_4__6__0_), .A2(n28), .ZN(
        pe_1_4_6_int_data_0_) );
  NAND2_X1 pe_1_4_6_U27 ( .A1(pe_1_4_6_n44), .A2(pe_1_4_6_n60), .ZN(
        pe_1_4_6_n41) );
  AND3_X1 pe_1_4_6_U26 ( .A1(n76), .A2(pe_1_4_6_n62), .A3(n50), .ZN(
        pe_1_4_6_n44) );
  INV_X1 pe_1_4_6_U25 ( .A(pe_1_4_6_int_data_3_), .ZN(pe_1_4_6_n74) );
  NOR2_X1 pe_1_4_6_U24 ( .A1(pe_1_4_6_n68), .A2(n50), .ZN(pe_1_4_6_n43) );
  NOR2_X1 pe_1_4_6_U23 ( .A1(pe_1_4_6_n57), .A2(pe_1_4_6_n63), .ZN(
        pe_1_4_6_n28) );
  NOR2_X1 pe_1_4_6_U22 ( .A1(n20), .A2(pe_1_4_6_n63), .ZN(pe_1_4_6_n27) );
  INV_X1 pe_1_4_6_U21 ( .A(pe_1_4_6_int_data_0_), .ZN(pe_1_4_6_n71) );
  INV_X1 pe_1_4_6_U20 ( .A(pe_1_4_6_n41), .ZN(pe_1_4_6_n88) );
  INV_X1 pe_1_4_6_U19 ( .A(pe_1_4_6_n37), .ZN(pe_1_4_6_n86) );
  INV_X1 pe_1_4_6_U18 ( .A(pe_1_4_6_n38), .ZN(pe_1_4_6_n85) );
  INV_X1 pe_1_4_6_U17 ( .A(pe_1_4_6_n39), .ZN(pe_1_4_6_n84) );
  NOR2_X1 pe_1_4_6_U16 ( .A1(pe_1_4_6_n66), .A2(pe_1_4_6_n42), .ZN(
        pe_1_4_6_N59) );
  NOR2_X1 pe_1_4_6_U15 ( .A1(pe_1_4_6_n66), .A2(pe_1_4_6_n41), .ZN(
        pe_1_4_6_N60) );
  NOR2_X1 pe_1_4_6_U14 ( .A1(pe_1_4_6_n66), .A2(pe_1_4_6_n38), .ZN(
        pe_1_4_6_N63) );
  NOR2_X1 pe_1_4_6_U13 ( .A1(pe_1_4_6_n66), .A2(pe_1_4_6_n40), .ZN(
        pe_1_4_6_N61) );
  NOR2_X1 pe_1_4_6_U12 ( .A1(pe_1_4_6_n66), .A2(pe_1_4_6_n39), .ZN(
        pe_1_4_6_N62) );
  NOR2_X1 pe_1_4_6_U11 ( .A1(pe_1_4_6_n37), .A2(pe_1_4_6_n66), .ZN(
        pe_1_4_6_N64) );
  NAND2_X1 pe_1_4_6_U10 ( .A1(pe_1_4_6_n44), .A2(pe_1_4_6_n59), .ZN(
        pe_1_4_6_n42) );
  BUF_X1 pe_1_4_6_U9 ( .A(pe_1_4_6_n59), .Z(pe_1_4_6_n55) );
  INV_X1 pe_1_4_6_U8 ( .A(pe_1_4_6_n67), .ZN(pe_1_4_6_n64) );
  BUF_X1 pe_1_4_6_U7 ( .A(pe_1_4_6_n59), .Z(pe_1_4_6_n56) );
  INV_X1 pe_1_4_6_U6 ( .A(pe_1_4_6_n42), .ZN(pe_1_4_6_n87) );
  INV_X1 pe_1_4_6_U5 ( .A(pe_1_4_6_n40), .ZN(pe_1_4_6_n83) );
  INV_X2 pe_1_4_6_U4 ( .A(n84), .ZN(pe_1_4_6_n70) );
  XOR2_X1 pe_1_4_6_U3 ( .A(pe_1_4_6_int_data_0_), .B(int_data_res_4__6__0_), 
        .Z(pe_1_4_6_n1) );
  DFFR_X1 pe_1_4_6_int_q_acc_reg_0_ ( .D(pe_1_4_6_n82), .CK(pe_1_4_6_net4588), 
        .RN(pe_1_4_6_n70), .Q(int_data_res_4__6__0_), .QN(pe_1_4_6_n3) );
  DFFR_X1 pe_1_4_6_int_q_reg_v_reg_0__0_ ( .D(int_data_y_5__6__0_), .CK(
        pe_1_4_6_net4558), .RN(pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_v[20]) );
  DFFR_X1 pe_1_4_6_int_q_reg_v_reg_0__1_ ( .D(int_data_y_5__6__1_), .CK(
        pe_1_4_6_net4558), .RN(pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_v[21]) );
  DFFR_X1 pe_1_4_6_int_q_reg_v_reg_0__2_ ( .D(int_data_y_5__6__2_), .CK(
        pe_1_4_6_net4558), .RN(pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_v[22]) );
  DFFR_X1 pe_1_4_6_int_q_reg_v_reg_0__3_ ( .D(int_data_y_5__6__3_), .CK(
        pe_1_4_6_net4558), .RN(pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_v[23]) );
  DFFR_X1 pe_1_4_6_int_q_reg_v_reg_1__0_ ( .D(int_data_y_5__6__0_), .CK(
        pe_1_4_6_net4563), .RN(pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_v[16]) );
  DFFR_X1 pe_1_4_6_int_q_reg_v_reg_1__1_ ( .D(int_data_y_5__6__1_), .CK(
        pe_1_4_6_net4563), .RN(pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_v[17]) );
  DFFR_X1 pe_1_4_6_int_q_reg_v_reg_1__2_ ( .D(int_data_y_5__6__2_), .CK(
        pe_1_4_6_net4563), .RN(pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_v[18]) );
  DFFR_X1 pe_1_4_6_int_q_reg_v_reg_1__3_ ( .D(int_data_y_5__6__3_), .CK(
        pe_1_4_6_net4563), .RN(pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_v[19]) );
  DFFR_X1 pe_1_4_6_int_q_reg_v_reg_2__0_ ( .D(int_data_y_5__6__0_), .CK(
        pe_1_4_6_net4568), .RN(pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_v[12]) );
  DFFR_X1 pe_1_4_6_int_q_reg_v_reg_2__1_ ( .D(int_data_y_5__6__1_), .CK(
        pe_1_4_6_net4568), .RN(pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_v[13]) );
  DFFR_X1 pe_1_4_6_int_q_reg_v_reg_2__2_ ( .D(int_data_y_5__6__2_), .CK(
        pe_1_4_6_net4568), .RN(pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_v[14]) );
  DFFR_X1 pe_1_4_6_int_q_reg_v_reg_2__3_ ( .D(int_data_y_5__6__3_), .CK(
        pe_1_4_6_net4568), .RN(pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_v[15]) );
  DFFR_X1 pe_1_4_6_int_q_reg_v_reg_3__0_ ( .D(int_data_y_5__6__0_), .CK(
        pe_1_4_6_net4573), .RN(pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_v[8]) );
  DFFR_X1 pe_1_4_6_int_q_reg_v_reg_3__1_ ( .D(int_data_y_5__6__1_), .CK(
        pe_1_4_6_net4573), .RN(pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_v[9]) );
  DFFR_X1 pe_1_4_6_int_q_reg_v_reg_3__2_ ( .D(int_data_y_5__6__2_), .CK(
        pe_1_4_6_net4573), .RN(pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_v[10]) );
  DFFR_X1 pe_1_4_6_int_q_reg_v_reg_3__3_ ( .D(int_data_y_5__6__3_), .CK(
        pe_1_4_6_net4573), .RN(pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_v[11]) );
  DFFR_X1 pe_1_4_6_int_q_reg_v_reg_4__0_ ( .D(int_data_y_5__6__0_), .CK(
        pe_1_4_6_net4578), .RN(pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_v[4]) );
  DFFR_X1 pe_1_4_6_int_q_reg_v_reg_4__1_ ( .D(int_data_y_5__6__1_), .CK(
        pe_1_4_6_net4578), .RN(pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_v[5]) );
  DFFR_X1 pe_1_4_6_int_q_reg_v_reg_4__2_ ( .D(int_data_y_5__6__2_), .CK(
        pe_1_4_6_net4578), .RN(pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_v[6]) );
  DFFR_X1 pe_1_4_6_int_q_reg_v_reg_4__3_ ( .D(int_data_y_5__6__3_), .CK(
        pe_1_4_6_net4578), .RN(pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_v[7]) );
  DFFR_X1 pe_1_4_6_int_q_reg_v_reg_5__0_ ( .D(int_data_y_5__6__0_), .CK(
        pe_1_4_6_net4583), .RN(pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_v[0]) );
  DFFR_X1 pe_1_4_6_int_q_reg_v_reg_5__1_ ( .D(int_data_y_5__6__1_), .CK(
        pe_1_4_6_net4583), .RN(pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_v[1]) );
  DFFR_X1 pe_1_4_6_int_q_reg_v_reg_5__2_ ( .D(int_data_y_5__6__2_), .CK(
        pe_1_4_6_net4583), .RN(pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_v[2]) );
  DFFR_X1 pe_1_4_6_int_q_reg_v_reg_5__3_ ( .D(int_data_y_5__6__3_), .CK(
        pe_1_4_6_net4583), .RN(pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_4_6_int_q_reg_h_reg_0__0_ ( .D(int_data_x_4__7__0_), .SI(
        int_data_y_5__6__0_), .SE(pe_1_4_6_n64), .CK(pe_1_4_6_net4527), .RN(
        pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_4_6_int_q_reg_h_reg_0__1_ ( .D(int_data_x_4__7__1_), .SI(
        int_data_y_5__6__1_), .SE(pe_1_4_6_n64), .CK(pe_1_4_6_net4527), .RN(
        pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_4_6_int_q_reg_h_reg_0__2_ ( .D(int_data_x_4__7__2_), .SI(
        int_data_y_5__6__2_), .SE(pe_1_4_6_n64), .CK(pe_1_4_6_net4527), .RN(
        pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_4_6_int_q_reg_h_reg_0__3_ ( .D(int_data_x_4__7__3_), .SI(
        int_data_y_5__6__3_), .SE(pe_1_4_6_n64), .CK(pe_1_4_6_net4527), .RN(
        pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_4_6_int_q_reg_h_reg_1__0_ ( .D(int_data_x_4__7__0_), .SI(
        int_data_y_5__6__0_), .SE(pe_1_4_6_n64), .CK(pe_1_4_6_net4533), .RN(
        pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_4_6_int_q_reg_h_reg_1__1_ ( .D(int_data_x_4__7__1_), .SI(
        int_data_y_5__6__1_), .SE(pe_1_4_6_n64), .CK(pe_1_4_6_net4533), .RN(
        pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_4_6_int_q_reg_h_reg_1__2_ ( .D(int_data_x_4__7__2_), .SI(
        int_data_y_5__6__2_), .SE(pe_1_4_6_n64), .CK(pe_1_4_6_net4533), .RN(
        pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_4_6_int_q_reg_h_reg_1__3_ ( .D(int_data_x_4__7__3_), .SI(
        int_data_y_5__6__3_), .SE(pe_1_4_6_n64), .CK(pe_1_4_6_net4533), .RN(
        pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_4_6_int_q_reg_h_reg_2__0_ ( .D(int_data_x_4__7__0_), .SI(
        int_data_y_5__6__0_), .SE(pe_1_4_6_n64), .CK(pe_1_4_6_net4538), .RN(
        pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_4_6_int_q_reg_h_reg_2__1_ ( .D(int_data_x_4__7__1_), .SI(
        int_data_y_5__6__1_), .SE(pe_1_4_6_n64), .CK(pe_1_4_6_net4538), .RN(
        pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_4_6_int_q_reg_h_reg_2__2_ ( .D(int_data_x_4__7__2_), .SI(
        int_data_y_5__6__2_), .SE(pe_1_4_6_n64), .CK(pe_1_4_6_net4538), .RN(
        pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_4_6_int_q_reg_h_reg_2__3_ ( .D(int_data_x_4__7__3_), .SI(
        int_data_y_5__6__3_), .SE(pe_1_4_6_n64), .CK(pe_1_4_6_net4538), .RN(
        pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_4_6_int_q_reg_h_reg_3__0_ ( .D(int_data_x_4__7__0_), .SI(
        int_data_y_5__6__0_), .SE(pe_1_4_6_n64), .CK(pe_1_4_6_net4543), .RN(
        pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_4_6_int_q_reg_h_reg_3__1_ ( .D(int_data_x_4__7__1_), .SI(
        int_data_y_5__6__1_), .SE(pe_1_4_6_n64), .CK(pe_1_4_6_net4543), .RN(
        pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_4_6_int_q_reg_h_reg_3__2_ ( .D(int_data_x_4__7__2_), .SI(
        int_data_y_5__6__2_), .SE(pe_1_4_6_n64), .CK(pe_1_4_6_net4543), .RN(
        pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_4_6_int_q_reg_h_reg_3__3_ ( .D(int_data_x_4__7__3_), .SI(
        int_data_y_5__6__3_), .SE(pe_1_4_6_n64), .CK(pe_1_4_6_net4543), .RN(
        pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_4_6_int_q_reg_h_reg_4__0_ ( .D(int_data_x_4__7__0_), .SI(
        int_data_y_5__6__0_), .SE(pe_1_4_6_n65), .CK(pe_1_4_6_net4548), .RN(
        pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_4_6_int_q_reg_h_reg_4__1_ ( .D(int_data_x_4__7__1_), .SI(
        int_data_y_5__6__1_), .SE(pe_1_4_6_n65), .CK(pe_1_4_6_net4548), .RN(
        pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_4_6_int_q_reg_h_reg_4__2_ ( .D(int_data_x_4__7__2_), .SI(
        int_data_y_5__6__2_), .SE(pe_1_4_6_n65), .CK(pe_1_4_6_net4548), .RN(
        pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_4_6_int_q_reg_h_reg_4__3_ ( .D(int_data_x_4__7__3_), .SI(
        int_data_y_5__6__3_), .SE(pe_1_4_6_n65), .CK(pe_1_4_6_net4548), .RN(
        pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_4_6_int_q_reg_h_reg_5__0_ ( .D(int_data_x_4__7__0_), .SI(
        int_data_y_5__6__0_), .SE(pe_1_4_6_n65), .CK(pe_1_4_6_net4553), .RN(
        pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_4_6_int_q_reg_h_reg_5__1_ ( .D(int_data_x_4__7__1_), .SI(
        int_data_y_5__6__1_), .SE(pe_1_4_6_n65), .CK(pe_1_4_6_net4553), .RN(
        pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_4_6_int_q_reg_h_reg_5__2_ ( .D(int_data_x_4__7__2_), .SI(
        int_data_y_5__6__2_), .SE(pe_1_4_6_n65), .CK(pe_1_4_6_net4553), .RN(
        pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_4_6_int_q_reg_h_reg_5__3_ ( .D(int_data_x_4__7__3_), .SI(
        int_data_y_5__6__3_), .SE(pe_1_4_6_n65), .CK(pe_1_4_6_net4553), .RN(
        pe_1_4_6_n70), .Q(pe_1_4_6_int_q_reg_h[3]) );
  FA_X1 pe_1_4_6_sub_81_U2_7 ( .A(int_data_res_4__6__7_), .B(pe_1_4_6_n74), 
        .CI(pe_1_4_6_sub_81_carry[7]), .S(pe_1_4_6_N77) );
  FA_X1 pe_1_4_6_sub_81_U2_6 ( .A(int_data_res_4__6__6_), .B(pe_1_4_6_n74), 
        .CI(pe_1_4_6_sub_81_carry[6]), .CO(pe_1_4_6_sub_81_carry[7]), .S(
        pe_1_4_6_N76) );
  FA_X1 pe_1_4_6_sub_81_U2_5 ( .A(int_data_res_4__6__5_), .B(pe_1_4_6_n74), 
        .CI(pe_1_4_6_sub_81_carry[5]), .CO(pe_1_4_6_sub_81_carry[6]), .S(
        pe_1_4_6_N75) );
  FA_X1 pe_1_4_6_sub_81_U2_4 ( .A(int_data_res_4__6__4_), .B(pe_1_4_6_n74), 
        .CI(pe_1_4_6_sub_81_carry[4]), .CO(pe_1_4_6_sub_81_carry[5]), .S(
        pe_1_4_6_N74) );
  FA_X1 pe_1_4_6_sub_81_U2_3 ( .A(int_data_res_4__6__3_), .B(pe_1_4_6_n74), 
        .CI(pe_1_4_6_sub_81_carry[3]), .CO(pe_1_4_6_sub_81_carry[4]), .S(
        pe_1_4_6_N73) );
  FA_X1 pe_1_4_6_sub_81_U2_2 ( .A(int_data_res_4__6__2_), .B(pe_1_4_6_n73), 
        .CI(pe_1_4_6_sub_81_carry[2]), .CO(pe_1_4_6_sub_81_carry[3]), .S(
        pe_1_4_6_N72) );
  FA_X1 pe_1_4_6_sub_81_U2_1 ( .A(int_data_res_4__6__1_), .B(pe_1_4_6_n72), 
        .CI(pe_1_4_6_sub_81_carry[1]), .CO(pe_1_4_6_sub_81_carry[2]), .S(
        pe_1_4_6_N71) );
  FA_X1 pe_1_4_6_add_83_U1_7 ( .A(int_data_res_4__6__7_), .B(
        pe_1_4_6_int_data_3_), .CI(pe_1_4_6_add_83_carry[7]), .S(pe_1_4_6_N85)
         );
  FA_X1 pe_1_4_6_add_83_U1_6 ( .A(int_data_res_4__6__6_), .B(
        pe_1_4_6_int_data_3_), .CI(pe_1_4_6_add_83_carry[6]), .CO(
        pe_1_4_6_add_83_carry[7]), .S(pe_1_4_6_N84) );
  FA_X1 pe_1_4_6_add_83_U1_5 ( .A(int_data_res_4__6__5_), .B(
        pe_1_4_6_int_data_3_), .CI(pe_1_4_6_add_83_carry[5]), .CO(
        pe_1_4_6_add_83_carry[6]), .S(pe_1_4_6_N83) );
  FA_X1 pe_1_4_6_add_83_U1_4 ( .A(int_data_res_4__6__4_), .B(
        pe_1_4_6_int_data_3_), .CI(pe_1_4_6_add_83_carry[4]), .CO(
        pe_1_4_6_add_83_carry[5]), .S(pe_1_4_6_N82) );
  FA_X1 pe_1_4_6_add_83_U1_3 ( .A(int_data_res_4__6__3_), .B(
        pe_1_4_6_int_data_3_), .CI(pe_1_4_6_add_83_carry[3]), .CO(
        pe_1_4_6_add_83_carry[4]), .S(pe_1_4_6_N81) );
  FA_X1 pe_1_4_6_add_83_U1_2 ( .A(int_data_res_4__6__2_), .B(
        pe_1_4_6_int_data_2_), .CI(pe_1_4_6_add_83_carry[2]), .CO(
        pe_1_4_6_add_83_carry[3]), .S(pe_1_4_6_N80) );
  FA_X1 pe_1_4_6_add_83_U1_1 ( .A(int_data_res_4__6__1_), .B(
        pe_1_4_6_int_data_1_), .CI(pe_1_4_6_n2), .CO(pe_1_4_6_add_83_carry[2]), 
        .S(pe_1_4_6_N79) );
  NAND3_X1 pe_1_4_6_U56 ( .A1(pe_1_4_6_n59), .A2(pe_1_4_6_n43), .A3(
        pe_1_4_6_n61), .ZN(pe_1_4_6_n40) );
  NAND3_X1 pe_1_4_6_U55 ( .A1(pe_1_4_6_n43), .A2(pe_1_4_6_n60), .A3(
        pe_1_4_6_n61), .ZN(pe_1_4_6_n39) );
  NAND3_X1 pe_1_4_6_U54 ( .A1(pe_1_4_6_n43), .A2(pe_1_4_6_n62), .A3(
        pe_1_4_6_n59), .ZN(pe_1_4_6_n38) );
  NAND3_X1 pe_1_4_6_U53 ( .A1(pe_1_4_6_n60), .A2(pe_1_4_6_n62), .A3(
        pe_1_4_6_n43), .ZN(pe_1_4_6_n37) );
  DFFR_X1 pe_1_4_6_int_q_acc_reg_6_ ( .D(pe_1_4_6_n76), .CK(pe_1_4_6_net4588), 
        .RN(pe_1_4_6_n69), .Q(int_data_res_4__6__6_) );
  DFFR_X1 pe_1_4_6_int_q_acc_reg_5_ ( .D(pe_1_4_6_n77), .CK(pe_1_4_6_net4588), 
        .RN(pe_1_4_6_n69), .Q(int_data_res_4__6__5_) );
  DFFR_X1 pe_1_4_6_int_q_acc_reg_4_ ( .D(pe_1_4_6_n78), .CK(pe_1_4_6_net4588), 
        .RN(pe_1_4_6_n69), .Q(int_data_res_4__6__4_) );
  DFFR_X1 pe_1_4_6_int_q_acc_reg_3_ ( .D(pe_1_4_6_n79), .CK(pe_1_4_6_net4588), 
        .RN(pe_1_4_6_n69), .Q(int_data_res_4__6__3_) );
  DFFR_X1 pe_1_4_6_int_q_acc_reg_2_ ( .D(pe_1_4_6_n80), .CK(pe_1_4_6_net4588), 
        .RN(pe_1_4_6_n69), .Q(int_data_res_4__6__2_) );
  DFFR_X1 pe_1_4_6_int_q_acc_reg_1_ ( .D(pe_1_4_6_n81), .CK(pe_1_4_6_net4588), 
        .RN(pe_1_4_6_n69), .Q(int_data_res_4__6__1_) );
  DFFR_X1 pe_1_4_6_int_q_acc_reg_7_ ( .D(pe_1_4_6_n75), .CK(pe_1_4_6_net4588), 
        .RN(pe_1_4_6_n69), .Q(int_data_res_4__6__7_) );
  CLKGATETST_X1 pe_1_4_6_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_4_6_n86), .SE(1'b0), .GCK(pe_1_4_6_net4527) );
  CLKGATETST_X1 pe_1_4_6_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_4_6_n85), .SE(1'b0), .GCK(pe_1_4_6_net4533) );
  CLKGATETST_X1 pe_1_4_6_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_4_6_n84), .SE(1'b0), .GCK(pe_1_4_6_net4538) );
  CLKGATETST_X1 pe_1_4_6_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_4_6_n83), .SE(1'b0), .GCK(pe_1_4_6_net4543) );
  CLKGATETST_X1 pe_1_4_6_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_4_6_n88), .SE(1'b0), .GCK(pe_1_4_6_net4548) );
  CLKGATETST_X1 pe_1_4_6_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_4_6_n87), .SE(1'b0), .GCK(pe_1_4_6_net4553) );
  CLKGATETST_X1 pe_1_4_6_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_4_6_N64), .SE(1'b0), .GCK(pe_1_4_6_net4558) );
  CLKGATETST_X1 pe_1_4_6_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_4_6_N63), .SE(1'b0), .GCK(pe_1_4_6_net4563) );
  CLKGATETST_X1 pe_1_4_6_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_4_6_N62), .SE(1'b0), .GCK(pe_1_4_6_net4568) );
  CLKGATETST_X1 pe_1_4_6_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_4_6_N61), .SE(1'b0), .GCK(pe_1_4_6_net4573) );
  CLKGATETST_X1 pe_1_4_6_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_4_6_N60), .SE(1'b0), .GCK(pe_1_4_6_net4578) );
  CLKGATETST_X1 pe_1_4_6_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_4_6_N59), .SE(1'b0), .GCK(pe_1_4_6_net4583) );
  CLKGATETST_X1 pe_1_4_6_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_4_6_N90), .SE(1'b0), .GCK(pe_1_4_6_net4588) );
  CLKBUF_X1 pe_1_4_7_U110 ( .A(pe_1_4_7_n70), .Z(pe_1_4_7_n69) );
  INV_X1 pe_1_4_7_U109 ( .A(n76), .ZN(pe_1_4_7_n68) );
  INV_X1 pe_1_4_7_U108 ( .A(n68), .ZN(pe_1_4_7_n67) );
  INV_X1 pe_1_4_7_U107 ( .A(n68), .ZN(pe_1_4_7_n66) );
  INV_X1 pe_1_4_7_U106 ( .A(pe_1_4_7_n67), .ZN(pe_1_4_7_n65) );
  INV_X1 pe_1_4_7_U105 ( .A(pe_1_4_7_n62), .ZN(pe_1_4_7_n61) );
  INV_X1 pe_1_4_7_U104 ( .A(pe_1_4_7_n60), .ZN(pe_1_4_7_n59) );
  INV_X1 pe_1_4_7_U103 ( .A(n28), .ZN(pe_1_4_7_n58) );
  INV_X1 pe_1_4_7_U102 ( .A(n20), .ZN(pe_1_4_7_n57) );
  MUX2_X1 pe_1_4_7_U101 ( .A(pe_1_4_7_n54), .B(pe_1_4_7_n51), .S(n50), .Z(
        int_data_x_4__7__3_) );
  MUX2_X1 pe_1_4_7_U100 ( .A(pe_1_4_7_n53), .B(pe_1_4_7_n52), .S(pe_1_4_7_n61), 
        .Z(pe_1_4_7_n54) );
  MUX2_X1 pe_1_4_7_U99 ( .A(pe_1_4_7_int_q_reg_h[23]), .B(
        pe_1_4_7_int_q_reg_h[19]), .S(pe_1_4_7_n56), .Z(pe_1_4_7_n53) );
  MUX2_X1 pe_1_4_7_U98 ( .A(pe_1_4_7_int_q_reg_h[15]), .B(
        pe_1_4_7_int_q_reg_h[11]), .S(pe_1_4_7_n56), .Z(pe_1_4_7_n52) );
  MUX2_X1 pe_1_4_7_U97 ( .A(pe_1_4_7_int_q_reg_h[7]), .B(
        pe_1_4_7_int_q_reg_h[3]), .S(pe_1_4_7_n56), .Z(pe_1_4_7_n51) );
  MUX2_X1 pe_1_4_7_U96 ( .A(pe_1_4_7_n50), .B(pe_1_4_7_n47), .S(n50), .Z(
        int_data_x_4__7__2_) );
  MUX2_X1 pe_1_4_7_U95 ( .A(pe_1_4_7_n49), .B(pe_1_4_7_n48), .S(pe_1_4_7_n61), 
        .Z(pe_1_4_7_n50) );
  MUX2_X1 pe_1_4_7_U94 ( .A(pe_1_4_7_int_q_reg_h[22]), .B(
        pe_1_4_7_int_q_reg_h[18]), .S(pe_1_4_7_n56), .Z(pe_1_4_7_n49) );
  MUX2_X1 pe_1_4_7_U93 ( .A(pe_1_4_7_int_q_reg_h[14]), .B(
        pe_1_4_7_int_q_reg_h[10]), .S(pe_1_4_7_n56), .Z(pe_1_4_7_n48) );
  MUX2_X1 pe_1_4_7_U92 ( .A(pe_1_4_7_int_q_reg_h[6]), .B(
        pe_1_4_7_int_q_reg_h[2]), .S(pe_1_4_7_n56), .Z(pe_1_4_7_n47) );
  MUX2_X1 pe_1_4_7_U91 ( .A(pe_1_4_7_n46), .B(pe_1_4_7_n24), .S(n50), .Z(
        int_data_x_4__7__1_) );
  MUX2_X1 pe_1_4_7_U90 ( .A(pe_1_4_7_n45), .B(pe_1_4_7_n25), .S(pe_1_4_7_n61), 
        .Z(pe_1_4_7_n46) );
  MUX2_X1 pe_1_4_7_U89 ( .A(pe_1_4_7_int_q_reg_h[21]), .B(
        pe_1_4_7_int_q_reg_h[17]), .S(pe_1_4_7_n56), .Z(pe_1_4_7_n45) );
  MUX2_X1 pe_1_4_7_U88 ( .A(pe_1_4_7_int_q_reg_h[13]), .B(
        pe_1_4_7_int_q_reg_h[9]), .S(pe_1_4_7_n56), .Z(pe_1_4_7_n25) );
  MUX2_X1 pe_1_4_7_U87 ( .A(pe_1_4_7_int_q_reg_h[5]), .B(
        pe_1_4_7_int_q_reg_h[1]), .S(pe_1_4_7_n56), .Z(pe_1_4_7_n24) );
  MUX2_X1 pe_1_4_7_U86 ( .A(pe_1_4_7_n23), .B(pe_1_4_7_n20), .S(n50), .Z(
        int_data_x_4__7__0_) );
  MUX2_X1 pe_1_4_7_U85 ( .A(pe_1_4_7_n22), .B(pe_1_4_7_n21), .S(pe_1_4_7_n61), 
        .Z(pe_1_4_7_n23) );
  MUX2_X1 pe_1_4_7_U84 ( .A(pe_1_4_7_int_q_reg_h[20]), .B(
        pe_1_4_7_int_q_reg_h[16]), .S(pe_1_4_7_n56), .Z(pe_1_4_7_n22) );
  MUX2_X1 pe_1_4_7_U83 ( .A(pe_1_4_7_int_q_reg_h[12]), .B(
        pe_1_4_7_int_q_reg_h[8]), .S(pe_1_4_7_n56), .Z(pe_1_4_7_n21) );
  MUX2_X1 pe_1_4_7_U82 ( .A(pe_1_4_7_int_q_reg_h[4]), .B(
        pe_1_4_7_int_q_reg_h[0]), .S(pe_1_4_7_n56), .Z(pe_1_4_7_n20) );
  MUX2_X1 pe_1_4_7_U81 ( .A(pe_1_4_7_n19), .B(pe_1_4_7_n16), .S(n50), .Z(
        int_data_y_4__7__3_) );
  MUX2_X1 pe_1_4_7_U80 ( .A(pe_1_4_7_n18), .B(pe_1_4_7_n17), .S(pe_1_4_7_n61), 
        .Z(pe_1_4_7_n19) );
  MUX2_X1 pe_1_4_7_U79 ( .A(pe_1_4_7_int_q_reg_v[23]), .B(
        pe_1_4_7_int_q_reg_v[19]), .S(pe_1_4_7_n55), .Z(pe_1_4_7_n18) );
  MUX2_X1 pe_1_4_7_U78 ( .A(pe_1_4_7_int_q_reg_v[15]), .B(
        pe_1_4_7_int_q_reg_v[11]), .S(pe_1_4_7_n55), .Z(pe_1_4_7_n17) );
  MUX2_X1 pe_1_4_7_U77 ( .A(pe_1_4_7_int_q_reg_v[7]), .B(
        pe_1_4_7_int_q_reg_v[3]), .S(pe_1_4_7_n55), .Z(pe_1_4_7_n16) );
  MUX2_X1 pe_1_4_7_U76 ( .A(pe_1_4_7_n15), .B(pe_1_4_7_n12), .S(n50), .Z(
        int_data_y_4__7__2_) );
  MUX2_X1 pe_1_4_7_U75 ( .A(pe_1_4_7_n14), .B(pe_1_4_7_n13), .S(pe_1_4_7_n61), 
        .Z(pe_1_4_7_n15) );
  MUX2_X1 pe_1_4_7_U74 ( .A(pe_1_4_7_int_q_reg_v[22]), .B(
        pe_1_4_7_int_q_reg_v[18]), .S(pe_1_4_7_n55), .Z(pe_1_4_7_n14) );
  MUX2_X1 pe_1_4_7_U73 ( .A(pe_1_4_7_int_q_reg_v[14]), .B(
        pe_1_4_7_int_q_reg_v[10]), .S(pe_1_4_7_n55), .Z(pe_1_4_7_n13) );
  MUX2_X1 pe_1_4_7_U72 ( .A(pe_1_4_7_int_q_reg_v[6]), .B(
        pe_1_4_7_int_q_reg_v[2]), .S(pe_1_4_7_n55), .Z(pe_1_4_7_n12) );
  MUX2_X1 pe_1_4_7_U71 ( .A(pe_1_4_7_n11), .B(pe_1_4_7_n8), .S(n50), .Z(
        int_data_y_4__7__1_) );
  MUX2_X1 pe_1_4_7_U70 ( .A(pe_1_4_7_n10), .B(pe_1_4_7_n9), .S(pe_1_4_7_n61), 
        .Z(pe_1_4_7_n11) );
  MUX2_X1 pe_1_4_7_U69 ( .A(pe_1_4_7_int_q_reg_v[21]), .B(
        pe_1_4_7_int_q_reg_v[17]), .S(pe_1_4_7_n55), .Z(pe_1_4_7_n10) );
  MUX2_X1 pe_1_4_7_U68 ( .A(pe_1_4_7_int_q_reg_v[13]), .B(
        pe_1_4_7_int_q_reg_v[9]), .S(pe_1_4_7_n55), .Z(pe_1_4_7_n9) );
  MUX2_X1 pe_1_4_7_U67 ( .A(pe_1_4_7_int_q_reg_v[5]), .B(
        pe_1_4_7_int_q_reg_v[1]), .S(pe_1_4_7_n55), .Z(pe_1_4_7_n8) );
  MUX2_X1 pe_1_4_7_U66 ( .A(pe_1_4_7_n7), .B(pe_1_4_7_n4), .S(n50), .Z(
        int_data_y_4__7__0_) );
  MUX2_X1 pe_1_4_7_U65 ( .A(pe_1_4_7_n6), .B(pe_1_4_7_n5), .S(pe_1_4_7_n61), 
        .Z(pe_1_4_7_n7) );
  MUX2_X1 pe_1_4_7_U64 ( .A(pe_1_4_7_int_q_reg_v[20]), .B(
        pe_1_4_7_int_q_reg_v[16]), .S(pe_1_4_7_n55), .Z(pe_1_4_7_n6) );
  MUX2_X1 pe_1_4_7_U63 ( .A(pe_1_4_7_int_q_reg_v[12]), .B(
        pe_1_4_7_int_q_reg_v[8]), .S(pe_1_4_7_n55), .Z(pe_1_4_7_n5) );
  MUX2_X1 pe_1_4_7_U62 ( .A(pe_1_4_7_int_q_reg_v[4]), .B(
        pe_1_4_7_int_q_reg_v[0]), .S(pe_1_4_7_n55), .Z(pe_1_4_7_n4) );
  AOI222_X1 pe_1_4_7_U61 ( .A1(int_data_res_5__7__2_), .A2(pe_1_4_7_n63), .B1(
        pe_1_4_7_N80), .B2(pe_1_4_7_n27), .C1(pe_1_4_7_N72), .C2(pe_1_4_7_n28), 
        .ZN(pe_1_4_7_n33) );
  INV_X1 pe_1_4_7_U60 ( .A(pe_1_4_7_n33), .ZN(pe_1_4_7_n80) );
  AOI222_X1 pe_1_4_7_U59 ( .A1(int_data_res_5__7__6_), .A2(pe_1_4_7_n63), .B1(
        pe_1_4_7_N84), .B2(pe_1_4_7_n27), .C1(pe_1_4_7_N76), .C2(pe_1_4_7_n28), 
        .ZN(pe_1_4_7_n29) );
  INV_X1 pe_1_4_7_U58 ( .A(pe_1_4_7_n29), .ZN(pe_1_4_7_n76) );
  XNOR2_X1 pe_1_4_7_U57 ( .A(pe_1_4_7_n71), .B(int_data_res_4__7__0_), .ZN(
        pe_1_4_7_N70) );
  AOI222_X1 pe_1_4_7_U52 ( .A1(int_data_res_5__7__0_), .A2(pe_1_4_7_n63), .B1(
        pe_1_4_7_n1), .B2(pe_1_4_7_n27), .C1(pe_1_4_7_N70), .C2(pe_1_4_7_n28), 
        .ZN(pe_1_4_7_n35) );
  INV_X1 pe_1_4_7_U51 ( .A(pe_1_4_7_n35), .ZN(pe_1_4_7_n82) );
  AOI222_X1 pe_1_4_7_U50 ( .A1(int_data_res_5__7__1_), .A2(pe_1_4_7_n63), .B1(
        pe_1_4_7_N79), .B2(pe_1_4_7_n27), .C1(pe_1_4_7_N71), .C2(pe_1_4_7_n28), 
        .ZN(pe_1_4_7_n34) );
  INV_X1 pe_1_4_7_U49 ( .A(pe_1_4_7_n34), .ZN(pe_1_4_7_n81) );
  AOI222_X1 pe_1_4_7_U48 ( .A1(int_data_res_5__7__3_), .A2(pe_1_4_7_n63), .B1(
        pe_1_4_7_N81), .B2(pe_1_4_7_n27), .C1(pe_1_4_7_N73), .C2(pe_1_4_7_n28), 
        .ZN(pe_1_4_7_n32) );
  INV_X1 pe_1_4_7_U47 ( .A(pe_1_4_7_n32), .ZN(pe_1_4_7_n79) );
  AOI222_X1 pe_1_4_7_U46 ( .A1(int_data_res_5__7__4_), .A2(pe_1_4_7_n63), .B1(
        pe_1_4_7_N82), .B2(pe_1_4_7_n27), .C1(pe_1_4_7_N74), .C2(pe_1_4_7_n28), 
        .ZN(pe_1_4_7_n31) );
  INV_X1 pe_1_4_7_U45 ( .A(pe_1_4_7_n31), .ZN(pe_1_4_7_n78) );
  AOI222_X1 pe_1_4_7_U44 ( .A1(int_data_res_5__7__5_), .A2(pe_1_4_7_n63), .B1(
        pe_1_4_7_N83), .B2(pe_1_4_7_n27), .C1(pe_1_4_7_N75), .C2(pe_1_4_7_n28), 
        .ZN(pe_1_4_7_n30) );
  INV_X1 pe_1_4_7_U43 ( .A(pe_1_4_7_n30), .ZN(pe_1_4_7_n77) );
  NAND2_X1 pe_1_4_7_U42 ( .A1(pe_1_4_7_int_data_0_), .A2(pe_1_4_7_n3), .ZN(
        pe_1_4_7_sub_81_carry[1]) );
  INV_X1 pe_1_4_7_U41 ( .A(pe_1_4_7_int_data_1_), .ZN(pe_1_4_7_n72) );
  INV_X1 pe_1_4_7_U40 ( .A(pe_1_4_7_int_data_2_), .ZN(pe_1_4_7_n73) );
  AND2_X1 pe_1_4_7_U39 ( .A1(pe_1_4_7_int_data_0_), .A2(int_data_res_4__7__0_), 
        .ZN(pe_1_4_7_n2) );
  AOI222_X1 pe_1_4_7_U38 ( .A1(pe_1_4_7_n63), .A2(int_data_res_5__7__7_), .B1(
        pe_1_4_7_N85), .B2(pe_1_4_7_n27), .C1(pe_1_4_7_N77), .C2(pe_1_4_7_n28), 
        .ZN(pe_1_4_7_n26) );
  INV_X1 pe_1_4_7_U37 ( .A(pe_1_4_7_n26), .ZN(pe_1_4_7_n75) );
  NOR3_X1 pe_1_4_7_U36 ( .A1(pe_1_4_7_n58), .A2(pe_1_4_7_n64), .A3(int_ckg[24]), .ZN(pe_1_4_7_n36) );
  OR2_X1 pe_1_4_7_U35 ( .A1(pe_1_4_7_n36), .A2(pe_1_4_7_n63), .ZN(pe_1_4_7_N90) );
  INV_X1 pe_1_4_7_U34 ( .A(n40), .ZN(pe_1_4_7_n62) );
  AND2_X1 pe_1_4_7_U33 ( .A1(int_data_x_4__7__2_), .A2(n28), .ZN(
        pe_1_4_7_int_data_2_) );
  AND2_X1 pe_1_4_7_U32 ( .A1(int_data_x_4__7__1_), .A2(n28), .ZN(
        pe_1_4_7_int_data_1_) );
  AND2_X1 pe_1_4_7_U31 ( .A1(int_data_x_4__7__3_), .A2(n28), .ZN(
        pe_1_4_7_int_data_3_) );
  BUF_X1 pe_1_4_7_U30 ( .A(n62), .Z(pe_1_4_7_n63) );
  INV_X1 pe_1_4_7_U29 ( .A(n34), .ZN(pe_1_4_7_n60) );
  AND2_X1 pe_1_4_7_U28 ( .A1(int_data_x_4__7__0_), .A2(n28), .ZN(
        pe_1_4_7_int_data_0_) );
  NAND2_X1 pe_1_4_7_U27 ( .A1(pe_1_4_7_n44), .A2(pe_1_4_7_n60), .ZN(
        pe_1_4_7_n41) );
  AND3_X1 pe_1_4_7_U26 ( .A1(n76), .A2(pe_1_4_7_n62), .A3(n50), .ZN(
        pe_1_4_7_n44) );
  INV_X1 pe_1_4_7_U25 ( .A(pe_1_4_7_int_data_3_), .ZN(pe_1_4_7_n74) );
  NOR2_X1 pe_1_4_7_U24 ( .A1(pe_1_4_7_n68), .A2(n50), .ZN(pe_1_4_7_n43) );
  NOR2_X1 pe_1_4_7_U23 ( .A1(pe_1_4_7_n57), .A2(pe_1_4_7_n63), .ZN(
        pe_1_4_7_n28) );
  NOR2_X1 pe_1_4_7_U22 ( .A1(n20), .A2(pe_1_4_7_n63), .ZN(pe_1_4_7_n27) );
  INV_X1 pe_1_4_7_U21 ( .A(pe_1_4_7_int_data_0_), .ZN(pe_1_4_7_n71) );
  INV_X1 pe_1_4_7_U20 ( .A(pe_1_4_7_n41), .ZN(pe_1_4_7_n88) );
  INV_X1 pe_1_4_7_U19 ( .A(pe_1_4_7_n37), .ZN(pe_1_4_7_n86) );
  INV_X1 pe_1_4_7_U18 ( .A(pe_1_4_7_n38), .ZN(pe_1_4_7_n85) );
  INV_X1 pe_1_4_7_U17 ( .A(pe_1_4_7_n39), .ZN(pe_1_4_7_n84) );
  NOR2_X1 pe_1_4_7_U16 ( .A1(pe_1_4_7_n66), .A2(pe_1_4_7_n42), .ZN(
        pe_1_4_7_N59) );
  NOR2_X1 pe_1_4_7_U15 ( .A1(pe_1_4_7_n66), .A2(pe_1_4_7_n41), .ZN(
        pe_1_4_7_N60) );
  NOR2_X1 pe_1_4_7_U14 ( .A1(pe_1_4_7_n66), .A2(pe_1_4_7_n38), .ZN(
        pe_1_4_7_N63) );
  NOR2_X1 pe_1_4_7_U13 ( .A1(pe_1_4_7_n66), .A2(pe_1_4_7_n40), .ZN(
        pe_1_4_7_N61) );
  NOR2_X1 pe_1_4_7_U12 ( .A1(pe_1_4_7_n66), .A2(pe_1_4_7_n39), .ZN(
        pe_1_4_7_N62) );
  NOR2_X1 pe_1_4_7_U11 ( .A1(pe_1_4_7_n37), .A2(pe_1_4_7_n66), .ZN(
        pe_1_4_7_N64) );
  NAND2_X1 pe_1_4_7_U10 ( .A1(pe_1_4_7_n44), .A2(pe_1_4_7_n59), .ZN(
        pe_1_4_7_n42) );
  BUF_X1 pe_1_4_7_U9 ( .A(pe_1_4_7_n59), .Z(pe_1_4_7_n55) );
  INV_X1 pe_1_4_7_U8 ( .A(pe_1_4_7_n67), .ZN(pe_1_4_7_n64) );
  BUF_X1 pe_1_4_7_U7 ( .A(pe_1_4_7_n59), .Z(pe_1_4_7_n56) );
  INV_X1 pe_1_4_7_U6 ( .A(pe_1_4_7_n42), .ZN(pe_1_4_7_n87) );
  INV_X1 pe_1_4_7_U5 ( .A(pe_1_4_7_n40), .ZN(pe_1_4_7_n83) );
  INV_X2 pe_1_4_7_U4 ( .A(n84), .ZN(pe_1_4_7_n70) );
  XOR2_X1 pe_1_4_7_U3 ( .A(pe_1_4_7_int_data_0_), .B(int_data_res_4__7__0_), 
        .Z(pe_1_4_7_n1) );
  DFFR_X1 pe_1_4_7_int_q_acc_reg_0_ ( .D(pe_1_4_7_n82), .CK(pe_1_4_7_net4510), 
        .RN(pe_1_4_7_n70), .Q(int_data_res_4__7__0_), .QN(pe_1_4_7_n3) );
  DFFR_X1 pe_1_4_7_int_q_reg_v_reg_0__0_ ( .D(int_data_y_5__7__0_), .CK(
        pe_1_4_7_net4480), .RN(pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_v[20]) );
  DFFR_X1 pe_1_4_7_int_q_reg_v_reg_0__1_ ( .D(int_data_y_5__7__1_), .CK(
        pe_1_4_7_net4480), .RN(pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_v[21]) );
  DFFR_X1 pe_1_4_7_int_q_reg_v_reg_0__2_ ( .D(int_data_y_5__7__2_), .CK(
        pe_1_4_7_net4480), .RN(pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_v[22]) );
  DFFR_X1 pe_1_4_7_int_q_reg_v_reg_0__3_ ( .D(int_data_y_5__7__3_), .CK(
        pe_1_4_7_net4480), .RN(pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_v[23]) );
  DFFR_X1 pe_1_4_7_int_q_reg_v_reg_1__0_ ( .D(int_data_y_5__7__0_), .CK(
        pe_1_4_7_net4485), .RN(pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_v[16]) );
  DFFR_X1 pe_1_4_7_int_q_reg_v_reg_1__1_ ( .D(int_data_y_5__7__1_), .CK(
        pe_1_4_7_net4485), .RN(pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_v[17]) );
  DFFR_X1 pe_1_4_7_int_q_reg_v_reg_1__2_ ( .D(int_data_y_5__7__2_), .CK(
        pe_1_4_7_net4485), .RN(pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_v[18]) );
  DFFR_X1 pe_1_4_7_int_q_reg_v_reg_1__3_ ( .D(int_data_y_5__7__3_), .CK(
        pe_1_4_7_net4485), .RN(pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_v[19]) );
  DFFR_X1 pe_1_4_7_int_q_reg_v_reg_2__0_ ( .D(int_data_y_5__7__0_), .CK(
        pe_1_4_7_net4490), .RN(pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_v[12]) );
  DFFR_X1 pe_1_4_7_int_q_reg_v_reg_2__1_ ( .D(int_data_y_5__7__1_), .CK(
        pe_1_4_7_net4490), .RN(pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_v[13]) );
  DFFR_X1 pe_1_4_7_int_q_reg_v_reg_2__2_ ( .D(int_data_y_5__7__2_), .CK(
        pe_1_4_7_net4490), .RN(pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_v[14]) );
  DFFR_X1 pe_1_4_7_int_q_reg_v_reg_2__3_ ( .D(int_data_y_5__7__3_), .CK(
        pe_1_4_7_net4490), .RN(pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_v[15]) );
  DFFR_X1 pe_1_4_7_int_q_reg_v_reg_3__0_ ( .D(int_data_y_5__7__0_), .CK(
        pe_1_4_7_net4495), .RN(pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_v[8]) );
  DFFR_X1 pe_1_4_7_int_q_reg_v_reg_3__1_ ( .D(int_data_y_5__7__1_), .CK(
        pe_1_4_7_net4495), .RN(pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_v[9]) );
  DFFR_X1 pe_1_4_7_int_q_reg_v_reg_3__2_ ( .D(int_data_y_5__7__2_), .CK(
        pe_1_4_7_net4495), .RN(pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_v[10]) );
  DFFR_X1 pe_1_4_7_int_q_reg_v_reg_3__3_ ( .D(int_data_y_5__7__3_), .CK(
        pe_1_4_7_net4495), .RN(pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_v[11]) );
  DFFR_X1 pe_1_4_7_int_q_reg_v_reg_4__0_ ( .D(int_data_y_5__7__0_), .CK(
        pe_1_4_7_net4500), .RN(pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_v[4]) );
  DFFR_X1 pe_1_4_7_int_q_reg_v_reg_4__1_ ( .D(int_data_y_5__7__1_), .CK(
        pe_1_4_7_net4500), .RN(pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_v[5]) );
  DFFR_X1 pe_1_4_7_int_q_reg_v_reg_4__2_ ( .D(int_data_y_5__7__2_), .CK(
        pe_1_4_7_net4500), .RN(pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_v[6]) );
  DFFR_X1 pe_1_4_7_int_q_reg_v_reg_4__3_ ( .D(int_data_y_5__7__3_), .CK(
        pe_1_4_7_net4500), .RN(pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_v[7]) );
  DFFR_X1 pe_1_4_7_int_q_reg_v_reg_5__0_ ( .D(int_data_y_5__7__0_), .CK(
        pe_1_4_7_net4505), .RN(pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_v[0]) );
  DFFR_X1 pe_1_4_7_int_q_reg_v_reg_5__1_ ( .D(int_data_y_5__7__1_), .CK(
        pe_1_4_7_net4505), .RN(pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_v[1]) );
  DFFR_X1 pe_1_4_7_int_q_reg_v_reg_5__2_ ( .D(int_data_y_5__7__2_), .CK(
        pe_1_4_7_net4505), .RN(pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_v[2]) );
  DFFR_X1 pe_1_4_7_int_q_reg_v_reg_5__3_ ( .D(int_data_y_5__7__3_), .CK(
        pe_1_4_7_net4505), .RN(pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_4_7_int_q_reg_h_reg_0__0_ ( .D(i_data_conv_h[12]), .SI(
        int_data_y_5__7__0_), .SE(pe_1_4_7_n64), .CK(pe_1_4_7_net4449), .RN(
        pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_4_7_int_q_reg_h_reg_0__1_ ( .D(i_data_conv_h[13]), .SI(
        int_data_y_5__7__1_), .SE(pe_1_4_7_n64), .CK(pe_1_4_7_net4449), .RN(
        pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_4_7_int_q_reg_h_reg_0__2_ ( .D(i_data_conv_h[14]), .SI(
        int_data_y_5__7__2_), .SE(pe_1_4_7_n64), .CK(pe_1_4_7_net4449), .RN(
        pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_4_7_int_q_reg_h_reg_0__3_ ( .D(i_data_conv_h[15]), .SI(
        int_data_y_5__7__3_), .SE(pe_1_4_7_n64), .CK(pe_1_4_7_net4449), .RN(
        pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_4_7_int_q_reg_h_reg_1__0_ ( .D(i_data_conv_h[12]), .SI(
        int_data_y_5__7__0_), .SE(pe_1_4_7_n64), .CK(pe_1_4_7_net4455), .RN(
        pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_4_7_int_q_reg_h_reg_1__1_ ( .D(i_data_conv_h[13]), .SI(
        int_data_y_5__7__1_), .SE(pe_1_4_7_n64), .CK(pe_1_4_7_net4455), .RN(
        pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_4_7_int_q_reg_h_reg_1__2_ ( .D(i_data_conv_h[14]), .SI(
        int_data_y_5__7__2_), .SE(pe_1_4_7_n64), .CK(pe_1_4_7_net4455), .RN(
        pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_4_7_int_q_reg_h_reg_1__3_ ( .D(i_data_conv_h[15]), .SI(
        int_data_y_5__7__3_), .SE(pe_1_4_7_n64), .CK(pe_1_4_7_net4455), .RN(
        pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_4_7_int_q_reg_h_reg_2__0_ ( .D(i_data_conv_h[12]), .SI(
        int_data_y_5__7__0_), .SE(pe_1_4_7_n64), .CK(pe_1_4_7_net4460), .RN(
        pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_4_7_int_q_reg_h_reg_2__1_ ( .D(i_data_conv_h[13]), .SI(
        int_data_y_5__7__1_), .SE(pe_1_4_7_n64), .CK(pe_1_4_7_net4460), .RN(
        pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_4_7_int_q_reg_h_reg_2__2_ ( .D(i_data_conv_h[14]), .SI(
        int_data_y_5__7__2_), .SE(pe_1_4_7_n64), .CK(pe_1_4_7_net4460), .RN(
        pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_4_7_int_q_reg_h_reg_2__3_ ( .D(i_data_conv_h[15]), .SI(
        int_data_y_5__7__3_), .SE(pe_1_4_7_n64), .CK(pe_1_4_7_net4460), .RN(
        pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_4_7_int_q_reg_h_reg_3__0_ ( .D(i_data_conv_h[12]), .SI(
        int_data_y_5__7__0_), .SE(pe_1_4_7_n64), .CK(pe_1_4_7_net4465), .RN(
        pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_4_7_int_q_reg_h_reg_3__1_ ( .D(i_data_conv_h[13]), .SI(
        int_data_y_5__7__1_), .SE(pe_1_4_7_n64), .CK(pe_1_4_7_net4465), .RN(
        pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_4_7_int_q_reg_h_reg_3__2_ ( .D(i_data_conv_h[14]), .SI(
        int_data_y_5__7__2_), .SE(pe_1_4_7_n64), .CK(pe_1_4_7_net4465), .RN(
        pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_4_7_int_q_reg_h_reg_3__3_ ( .D(i_data_conv_h[15]), .SI(
        int_data_y_5__7__3_), .SE(pe_1_4_7_n64), .CK(pe_1_4_7_net4465), .RN(
        pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_4_7_int_q_reg_h_reg_4__0_ ( .D(i_data_conv_h[12]), .SI(
        int_data_y_5__7__0_), .SE(pe_1_4_7_n65), .CK(pe_1_4_7_net4470), .RN(
        pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_4_7_int_q_reg_h_reg_4__1_ ( .D(i_data_conv_h[13]), .SI(
        int_data_y_5__7__1_), .SE(pe_1_4_7_n65), .CK(pe_1_4_7_net4470), .RN(
        pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_4_7_int_q_reg_h_reg_4__2_ ( .D(i_data_conv_h[14]), .SI(
        int_data_y_5__7__2_), .SE(pe_1_4_7_n65), .CK(pe_1_4_7_net4470), .RN(
        pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_4_7_int_q_reg_h_reg_4__3_ ( .D(i_data_conv_h[15]), .SI(
        int_data_y_5__7__3_), .SE(pe_1_4_7_n65), .CK(pe_1_4_7_net4470), .RN(
        pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_4_7_int_q_reg_h_reg_5__0_ ( .D(i_data_conv_h[12]), .SI(
        int_data_y_5__7__0_), .SE(pe_1_4_7_n65), .CK(pe_1_4_7_net4475), .RN(
        pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_4_7_int_q_reg_h_reg_5__1_ ( .D(i_data_conv_h[13]), .SI(
        int_data_y_5__7__1_), .SE(pe_1_4_7_n65), .CK(pe_1_4_7_net4475), .RN(
        pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_4_7_int_q_reg_h_reg_5__2_ ( .D(i_data_conv_h[14]), .SI(
        int_data_y_5__7__2_), .SE(pe_1_4_7_n65), .CK(pe_1_4_7_net4475), .RN(
        pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_4_7_int_q_reg_h_reg_5__3_ ( .D(i_data_conv_h[15]), .SI(
        int_data_y_5__7__3_), .SE(pe_1_4_7_n65), .CK(pe_1_4_7_net4475), .RN(
        pe_1_4_7_n70), .Q(pe_1_4_7_int_q_reg_h[3]) );
  FA_X1 pe_1_4_7_sub_81_U2_7 ( .A(int_data_res_4__7__7_), .B(pe_1_4_7_n74), 
        .CI(pe_1_4_7_sub_81_carry[7]), .S(pe_1_4_7_N77) );
  FA_X1 pe_1_4_7_sub_81_U2_6 ( .A(int_data_res_4__7__6_), .B(pe_1_4_7_n74), 
        .CI(pe_1_4_7_sub_81_carry[6]), .CO(pe_1_4_7_sub_81_carry[7]), .S(
        pe_1_4_7_N76) );
  FA_X1 pe_1_4_7_sub_81_U2_5 ( .A(int_data_res_4__7__5_), .B(pe_1_4_7_n74), 
        .CI(pe_1_4_7_sub_81_carry[5]), .CO(pe_1_4_7_sub_81_carry[6]), .S(
        pe_1_4_7_N75) );
  FA_X1 pe_1_4_7_sub_81_U2_4 ( .A(int_data_res_4__7__4_), .B(pe_1_4_7_n74), 
        .CI(pe_1_4_7_sub_81_carry[4]), .CO(pe_1_4_7_sub_81_carry[5]), .S(
        pe_1_4_7_N74) );
  FA_X1 pe_1_4_7_sub_81_U2_3 ( .A(int_data_res_4__7__3_), .B(pe_1_4_7_n74), 
        .CI(pe_1_4_7_sub_81_carry[3]), .CO(pe_1_4_7_sub_81_carry[4]), .S(
        pe_1_4_7_N73) );
  FA_X1 pe_1_4_7_sub_81_U2_2 ( .A(int_data_res_4__7__2_), .B(pe_1_4_7_n73), 
        .CI(pe_1_4_7_sub_81_carry[2]), .CO(pe_1_4_7_sub_81_carry[3]), .S(
        pe_1_4_7_N72) );
  FA_X1 pe_1_4_7_sub_81_U2_1 ( .A(int_data_res_4__7__1_), .B(pe_1_4_7_n72), 
        .CI(pe_1_4_7_sub_81_carry[1]), .CO(pe_1_4_7_sub_81_carry[2]), .S(
        pe_1_4_7_N71) );
  FA_X1 pe_1_4_7_add_83_U1_7 ( .A(int_data_res_4__7__7_), .B(
        pe_1_4_7_int_data_3_), .CI(pe_1_4_7_add_83_carry[7]), .S(pe_1_4_7_N85)
         );
  FA_X1 pe_1_4_7_add_83_U1_6 ( .A(int_data_res_4__7__6_), .B(
        pe_1_4_7_int_data_3_), .CI(pe_1_4_7_add_83_carry[6]), .CO(
        pe_1_4_7_add_83_carry[7]), .S(pe_1_4_7_N84) );
  FA_X1 pe_1_4_7_add_83_U1_5 ( .A(int_data_res_4__7__5_), .B(
        pe_1_4_7_int_data_3_), .CI(pe_1_4_7_add_83_carry[5]), .CO(
        pe_1_4_7_add_83_carry[6]), .S(pe_1_4_7_N83) );
  FA_X1 pe_1_4_7_add_83_U1_4 ( .A(int_data_res_4__7__4_), .B(
        pe_1_4_7_int_data_3_), .CI(pe_1_4_7_add_83_carry[4]), .CO(
        pe_1_4_7_add_83_carry[5]), .S(pe_1_4_7_N82) );
  FA_X1 pe_1_4_7_add_83_U1_3 ( .A(int_data_res_4__7__3_), .B(
        pe_1_4_7_int_data_3_), .CI(pe_1_4_7_add_83_carry[3]), .CO(
        pe_1_4_7_add_83_carry[4]), .S(pe_1_4_7_N81) );
  FA_X1 pe_1_4_7_add_83_U1_2 ( .A(int_data_res_4__7__2_), .B(
        pe_1_4_7_int_data_2_), .CI(pe_1_4_7_add_83_carry[2]), .CO(
        pe_1_4_7_add_83_carry[3]), .S(pe_1_4_7_N80) );
  FA_X1 pe_1_4_7_add_83_U1_1 ( .A(int_data_res_4__7__1_), .B(
        pe_1_4_7_int_data_1_), .CI(pe_1_4_7_n2), .CO(pe_1_4_7_add_83_carry[2]), 
        .S(pe_1_4_7_N79) );
  NAND3_X1 pe_1_4_7_U56 ( .A1(pe_1_4_7_n59), .A2(pe_1_4_7_n43), .A3(
        pe_1_4_7_n61), .ZN(pe_1_4_7_n40) );
  NAND3_X1 pe_1_4_7_U55 ( .A1(pe_1_4_7_n43), .A2(pe_1_4_7_n60), .A3(
        pe_1_4_7_n61), .ZN(pe_1_4_7_n39) );
  NAND3_X1 pe_1_4_7_U54 ( .A1(pe_1_4_7_n43), .A2(pe_1_4_7_n62), .A3(
        pe_1_4_7_n59), .ZN(pe_1_4_7_n38) );
  NAND3_X1 pe_1_4_7_U53 ( .A1(pe_1_4_7_n60), .A2(pe_1_4_7_n62), .A3(
        pe_1_4_7_n43), .ZN(pe_1_4_7_n37) );
  DFFR_X1 pe_1_4_7_int_q_acc_reg_6_ ( .D(pe_1_4_7_n76), .CK(pe_1_4_7_net4510), 
        .RN(pe_1_4_7_n69), .Q(int_data_res_4__7__6_) );
  DFFR_X1 pe_1_4_7_int_q_acc_reg_5_ ( .D(pe_1_4_7_n77), .CK(pe_1_4_7_net4510), 
        .RN(pe_1_4_7_n69), .Q(int_data_res_4__7__5_) );
  DFFR_X1 pe_1_4_7_int_q_acc_reg_4_ ( .D(pe_1_4_7_n78), .CK(pe_1_4_7_net4510), 
        .RN(pe_1_4_7_n69), .Q(int_data_res_4__7__4_) );
  DFFR_X1 pe_1_4_7_int_q_acc_reg_3_ ( .D(pe_1_4_7_n79), .CK(pe_1_4_7_net4510), 
        .RN(pe_1_4_7_n69), .Q(int_data_res_4__7__3_) );
  DFFR_X1 pe_1_4_7_int_q_acc_reg_2_ ( .D(pe_1_4_7_n80), .CK(pe_1_4_7_net4510), 
        .RN(pe_1_4_7_n69), .Q(int_data_res_4__7__2_) );
  DFFR_X1 pe_1_4_7_int_q_acc_reg_1_ ( .D(pe_1_4_7_n81), .CK(pe_1_4_7_net4510), 
        .RN(pe_1_4_7_n69), .Q(int_data_res_4__7__1_) );
  DFFR_X1 pe_1_4_7_int_q_acc_reg_7_ ( .D(pe_1_4_7_n75), .CK(pe_1_4_7_net4510), 
        .RN(pe_1_4_7_n69), .Q(int_data_res_4__7__7_) );
  CLKGATETST_X1 pe_1_4_7_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_4_7_n86), .SE(1'b0), .GCK(pe_1_4_7_net4449) );
  CLKGATETST_X1 pe_1_4_7_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_4_7_n85), .SE(1'b0), .GCK(pe_1_4_7_net4455) );
  CLKGATETST_X1 pe_1_4_7_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_4_7_n84), .SE(1'b0), .GCK(pe_1_4_7_net4460) );
  CLKGATETST_X1 pe_1_4_7_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_4_7_n83), .SE(1'b0), .GCK(pe_1_4_7_net4465) );
  CLKGATETST_X1 pe_1_4_7_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_4_7_n88), .SE(1'b0), .GCK(pe_1_4_7_net4470) );
  CLKGATETST_X1 pe_1_4_7_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_4_7_n87), .SE(1'b0), .GCK(pe_1_4_7_net4475) );
  CLKGATETST_X1 pe_1_4_7_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_4_7_N64), .SE(1'b0), .GCK(pe_1_4_7_net4480) );
  CLKGATETST_X1 pe_1_4_7_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_4_7_N63), .SE(1'b0), .GCK(pe_1_4_7_net4485) );
  CLKGATETST_X1 pe_1_4_7_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_4_7_N62), .SE(1'b0), .GCK(pe_1_4_7_net4490) );
  CLKGATETST_X1 pe_1_4_7_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_4_7_N61), .SE(1'b0), .GCK(pe_1_4_7_net4495) );
  CLKGATETST_X1 pe_1_4_7_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_4_7_N60), .SE(1'b0), .GCK(pe_1_4_7_net4500) );
  CLKGATETST_X1 pe_1_4_7_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_4_7_N59), .SE(1'b0), .GCK(pe_1_4_7_net4505) );
  CLKGATETST_X1 pe_1_4_7_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_4_7_N90), .SE(1'b0), .GCK(pe_1_4_7_net4510) );
  CLKBUF_X1 pe_1_5_0_U111 ( .A(pe_1_5_0_n71), .Z(pe_1_5_0_n70) );
  INV_X1 pe_1_5_0_U110 ( .A(n76), .ZN(pe_1_5_0_n69) );
  INV_X1 pe_1_5_0_U109 ( .A(n68), .ZN(pe_1_5_0_n68) );
  INV_X1 pe_1_5_0_U108 ( .A(n68), .ZN(pe_1_5_0_n67) );
  INV_X1 pe_1_5_0_U107 ( .A(n68), .ZN(pe_1_5_0_n66) );
  INV_X1 pe_1_5_0_U106 ( .A(pe_1_5_0_n68), .ZN(pe_1_5_0_n65) );
  INV_X1 pe_1_5_0_U105 ( .A(pe_1_5_0_n62), .ZN(pe_1_5_0_n61) );
  INV_X1 pe_1_5_0_U104 ( .A(n28), .ZN(pe_1_5_0_n59) );
  INV_X1 pe_1_5_0_U103 ( .A(pe_1_5_0_n59), .ZN(pe_1_5_0_n58) );
  INV_X1 pe_1_5_0_U102 ( .A(n20), .ZN(pe_1_5_0_n57) );
  MUX2_X1 pe_1_5_0_U101 ( .A(pe_1_5_0_n54), .B(pe_1_5_0_n51), .S(n51), .Z(
        pe_1_5_0_o_data_h_3_) );
  MUX2_X1 pe_1_5_0_U100 ( .A(pe_1_5_0_n53), .B(pe_1_5_0_n52), .S(pe_1_5_0_n61), 
        .Z(pe_1_5_0_n54) );
  MUX2_X1 pe_1_5_0_U99 ( .A(pe_1_5_0_int_q_reg_h[23]), .B(
        pe_1_5_0_int_q_reg_h[19]), .S(pe_1_5_0_n56), .Z(pe_1_5_0_n53) );
  MUX2_X1 pe_1_5_0_U98 ( .A(pe_1_5_0_int_q_reg_h[15]), .B(
        pe_1_5_0_int_q_reg_h[11]), .S(pe_1_5_0_n56), .Z(pe_1_5_0_n52) );
  MUX2_X1 pe_1_5_0_U97 ( .A(pe_1_5_0_int_q_reg_h[7]), .B(
        pe_1_5_0_int_q_reg_h[3]), .S(pe_1_5_0_n56), .Z(pe_1_5_0_n51) );
  MUX2_X1 pe_1_5_0_U96 ( .A(pe_1_5_0_n50), .B(pe_1_5_0_n47), .S(n51), .Z(
        pe_1_5_0_o_data_h_2_) );
  MUX2_X1 pe_1_5_0_U95 ( .A(pe_1_5_0_n49), .B(pe_1_5_0_n48), .S(pe_1_5_0_n61), 
        .Z(pe_1_5_0_n50) );
  MUX2_X1 pe_1_5_0_U94 ( .A(pe_1_5_0_int_q_reg_h[22]), .B(
        pe_1_5_0_int_q_reg_h[18]), .S(pe_1_5_0_n56), .Z(pe_1_5_0_n49) );
  MUX2_X1 pe_1_5_0_U93 ( .A(pe_1_5_0_int_q_reg_h[14]), .B(
        pe_1_5_0_int_q_reg_h[10]), .S(pe_1_5_0_n56), .Z(pe_1_5_0_n48) );
  MUX2_X1 pe_1_5_0_U92 ( .A(pe_1_5_0_int_q_reg_h[6]), .B(
        pe_1_5_0_int_q_reg_h[2]), .S(pe_1_5_0_n56), .Z(pe_1_5_0_n47) );
  MUX2_X1 pe_1_5_0_U91 ( .A(pe_1_5_0_n46), .B(pe_1_5_0_n24), .S(n51), .Z(
        pe_1_5_0_o_data_h_1_) );
  MUX2_X1 pe_1_5_0_U90 ( .A(pe_1_5_0_n45), .B(pe_1_5_0_n25), .S(pe_1_5_0_n61), 
        .Z(pe_1_5_0_n46) );
  MUX2_X1 pe_1_5_0_U89 ( .A(pe_1_5_0_int_q_reg_h[21]), .B(
        pe_1_5_0_int_q_reg_h[17]), .S(pe_1_5_0_n56), .Z(pe_1_5_0_n45) );
  MUX2_X1 pe_1_5_0_U88 ( .A(pe_1_5_0_int_q_reg_h[13]), .B(
        pe_1_5_0_int_q_reg_h[9]), .S(pe_1_5_0_n56), .Z(pe_1_5_0_n25) );
  MUX2_X1 pe_1_5_0_U87 ( .A(pe_1_5_0_int_q_reg_h[5]), .B(
        pe_1_5_0_int_q_reg_h[1]), .S(pe_1_5_0_n56), .Z(pe_1_5_0_n24) );
  MUX2_X1 pe_1_5_0_U86 ( .A(pe_1_5_0_n23), .B(pe_1_5_0_n20), .S(n51), .Z(
        pe_1_5_0_o_data_h_0_) );
  MUX2_X1 pe_1_5_0_U85 ( .A(pe_1_5_0_n22), .B(pe_1_5_0_n21), .S(pe_1_5_0_n61), 
        .Z(pe_1_5_0_n23) );
  MUX2_X1 pe_1_5_0_U84 ( .A(pe_1_5_0_int_q_reg_h[20]), .B(
        pe_1_5_0_int_q_reg_h[16]), .S(pe_1_5_0_n56), .Z(pe_1_5_0_n22) );
  MUX2_X1 pe_1_5_0_U83 ( .A(pe_1_5_0_int_q_reg_h[12]), .B(
        pe_1_5_0_int_q_reg_h[8]), .S(pe_1_5_0_n56), .Z(pe_1_5_0_n21) );
  MUX2_X1 pe_1_5_0_U82 ( .A(pe_1_5_0_int_q_reg_h[4]), .B(
        pe_1_5_0_int_q_reg_h[0]), .S(pe_1_5_0_n56), .Z(pe_1_5_0_n20) );
  MUX2_X1 pe_1_5_0_U81 ( .A(pe_1_5_0_n19), .B(pe_1_5_0_n16), .S(n51), .Z(
        int_data_y_5__0__3_) );
  MUX2_X1 pe_1_5_0_U80 ( .A(pe_1_5_0_n18), .B(pe_1_5_0_n17), .S(pe_1_5_0_n61), 
        .Z(pe_1_5_0_n19) );
  MUX2_X1 pe_1_5_0_U79 ( .A(pe_1_5_0_int_q_reg_v[23]), .B(
        pe_1_5_0_int_q_reg_v[19]), .S(pe_1_5_0_n55), .Z(pe_1_5_0_n18) );
  MUX2_X1 pe_1_5_0_U78 ( .A(pe_1_5_0_int_q_reg_v[15]), .B(
        pe_1_5_0_int_q_reg_v[11]), .S(pe_1_5_0_n55), .Z(pe_1_5_0_n17) );
  MUX2_X1 pe_1_5_0_U77 ( .A(pe_1_5_0_int_q_reg_v[7]), .B(
        pe_1_5_0_int_q_reg_v[3]), .S(pe_1_5_0_n55), .Z(pe_1_5_0_n16) );
  MUX2_X1 pe_1_5_0_U76 ( .A(pe_1_5_0_n15), .B(pe_1_5_0_n12), .S(n51), .Z(
        int_data_y_5__0__2_) );
  MUX2_X1 pe_1_5_0_U75 ( .A(pe_1_5_0_n14), .B(pe_1_5_0_n13), .S(pe_1_5_0_n61), 
        .Z(pe_1_5_0_n15) );
  MUX2_X1 pe_1_5_0_U74 ( .A(pe_1_5_0_int_q_reg_v[22]), .B(
        pe_1_5_0_int_q_reg_v[18]), .S(pe_1_5_0_n55), .Z(pe_1_5_0_n14) );
  MUX2_X1 pe_1_5_0_U73 ( .A(pe_1_5_0_int_q_reg_v[14]), .B(
        pe_1_5_0_int_q_reg_v[10]), .S(pe_1_5_0_n55), .Z(pe_1_5_0_n13) );
  MUX2_X1 pe_1_5_0_U72 ( .A(pe_1_5_0_int_q_reg_v[6]), .B(
        pe_1_5_0_int_q_reg_v[2]), .S(pe_1_5_0_n55), .Z(pe_1_5_0_n12) );
  MUX2_X1 pe_1_5_0_U71 ( .A(pe_1_5_0_n11), .B(pe_1_5_0_n8), .S(n51), .Z(
        int_data_y_5__0__1_) );
  MUX2_X1 pe_1_5_0_U70 ( .A(pe_1_5_0_n10), .B(pe_1_5_0_n9), .S(pe_1_5_0_n61), 
        .Z(pe_1_5_0_n11) );
  MUX2_X1 pe_1_5_0_U69 ( .A(pe_1_5_0_int_q_reg_v[21]), .B(
        pe_1_5_0_int_q_reg_v[17]), .S(pe_1_5_0_n55), .Z(pe_1_5_0_n10) );
  MUX2_X1 pe_1_5_0_U68 ( .A(pe_1_5_0_int_q_reg_v[13]), .B(
        pe_1_5_0_int_q_reg_v[9]), .S(pe_1_5_0_n55), .Z(pe_1_5_0_n9) );
  MUX2_X1 pe_1_5_0_U67 ( .A(pe_1_5_0_int_q_reg_v[5]), .B(
        pe_1_5_0_int_q_reg_v[1]), .S(pe_1_5_0_n55), .Z(pe_1_5_0_n8) );
  MUX2_X1 pe_1_5_0_U66 ( .A(pe_1_5_0_n7), .B(pe_1_5_0_n4), .S(n51), .Z(
        int_data_y_5__0__0_) );
  MUX2_X1 pe_1_5_0_U65 ( .A(pe_1_5_0_n6), .B(pe_1_5_0_n5), .S(pe_1_5_0_n61), 
        .Z(pe_1_5_0_n7) );
  MUX2_X1 pe_1_5_0_U64 ( .A(pe_1_5_0_int_q_reg_v[20]), .B(
        pe_1_5_0_int_q_reg_v[16]), .S(pe_1_5_0_n55), .Z(pe_1_5_0_n6) );
  MUX2_X1 pe_1_5_0_U63 ( .A(pe_1_5_0_int_q_reg_v[12]), .B(
        pe_1_5_0_int_q_reg_v[8]), .S(pe_1_5_0_n55), .Z(pe_1_5_0_n5) );
  MUX2_X1 pe_1_5_0_U62 ( .A(pe_1_5_0_int_q_reg_v[4]), .B(
        pe_1_5_0_int_q_reg_v[0]), .S(pe_1_5_0_n55), .Z(pe_1_5_0_n4) );
  AND2_X1 pe_1_5_0_U61 ( .A1(pe_1_5_0_o_data_h_3_), .A2(pe_1_5_0_n58), .ZN(
        pe_1_5_0_int_data_3_) );
  NAND2_X1 pe_1_5_0_U60 ( .A1(pe_1_5_0_int_data_0_), .A2(pe_1_5_0_n3), .ZN(
        pe_1_5_0_sub_81_carry[1]) );
  INV_X1 pe_1_5_0_U59 ( .A(pe_1_5_0_int_data_1_), .ZN(pe_1_5_0_n73) );
  AOI222_X1 pe_1_5_0_U58 ( .A1(pe_1_5_0_n63), .A2(int_data_res_6__0__7_), .B1(
        pe_1_5_0_N85), .B2(pe_1_5_0_n27), .C1(pe_1_5_0_N77), .C2(pe_1_5_0_n28), 
        .ZN(pe_1_5_0_n26) );
  INV_X1 pe_1_5_0_U57 ( .A(pe_1_5_0_n26), .ZN(pe_1_5_0_n76) );
  AOI222_X1 pe_1_5_0_U52 ( .A1(int_data_res_6__0__1_), .A2(pe_1_5_0_n63), .B1(
        pe_1_5_0_N79), .B2(pe_1_5_0_n27), .C1(pe_1_5_0_N71), .C2(pe_1_5_0_n28), 
        .ZN(pe_1_5_0_n34) );
  INV_X1 pe_1_5_0_U51 ( .A(pe_1_5_0_n34), .ZN(pe_1_5_0_n82) );
  AOI222_X1 pe_1_5_0_U50 ( .A1(int_data_res_6__0__2_), .A2(pe_1_5_0_n63), .B1(
        pe_1_5_0_N80), .B2(pe_1_5_0_n27), .C1(pe_1_5_0_N72), .C2(pe_1_5_0_n28), 
        .ZN(pe_1_5_0_n33) );
  INV_X1 pe_1_5_0_U49 ( .A(pe_1_5_0_n33), .ZN(pe_1_5_0_n81) );
  AOI222_X1 pe_1_5_0_U48 ( .A1(int_data_res_6__0__6_), .A2(pe_1_5_0_n63), .B1(
        pe_1_5_0_N84), .B2(pe_1_5_0_n27), .C1(pe_1_5_0_N76), .C2(pe_1_5_0_n28), 
        .ZN(pe_1_5_0_n29) );
  INV_X1 pe_1_5_0_U47 ( .A(pe_1_5_0_n29), .ZN(pe_1_5_0_n77) );
  AND2_X1 pe_1_5_0_U46 ( .A1(pe_1_5_0_o_data_h_2_), .A2(pe_1_5_0_n58), .ZN(
        pe_1_5_0_int_data_2_) );
  AND2_X1 pe_1_5_0_U45 ( .A1(pe_1_5_0_o_data_h_1_), .A2(pe_1_5_0_n58), .ZN(
        pe_1_5_0_int_data_1_) );
  INV_X1 pe_1_5_0_U44 ( .A(pe_1_5_0_int_data_2_), .ZN(pe_1_5_0_n74) );
  AND2_X1 pe_1_5_0_U43 ( .A1(pe_1_5_0_int_data_0_), .A2(int_data_res_5__0__0_), 
        .ZN(pe_1_5_0_n2) );
  AND2_X1 pe_1_5_0_U42 ( .A1(pe_1_5_0_o_data_h_0_), .A2(pe_1_5_0_n58), .ZN(
        pe_1_5_0_int_data_0_) );
  XNOR2_X1 pe_1_5_0_U41 ( .A(pe_1_5_0_n72), .B(int_data_res_5__0__0_), .ZN(
        pe_1_5_0_N70) );
  AOI222_X1 pe_1_5_0_U40 ( .A1(int_data_res_6__0__0_), .A2(pe_1_5_0_n63), .B1(
        pe_1_5_0_n1), .B2(pe_1_5_0_n27), .C1(pe_1_5_0_N70), .C2(pe_1_5_0_n28), 
        .ZN(pe_1_5_0_n35) );
  INV_X1 pe_1_5_0_U39 ( .A(pe_1_5_0_n35), .ZN(pe_1_5_0_n83) );
  AOI222_X1 pe_1_5_0_U38 ( .A1(int_data_res_6__0__3_), .A2(pe_1_5_0_n63), .B1(
        pe_1_5_0_N81), .B2(pe_1_5_0_n27), .C1(pe_1_5_0_N73), .C2(pe_1_5_0_n28), 
        .ZN(pe_1_5_0_n32) );
  INV_X1 pe_1_5_0_U37 ( .A(pe_1_5_0_n32), .ZN(pe_1_5_0_n80) );
  AOI222_X1 pe_1_5_0_U36 ( .A1(int_data_res_6__0__4_), .A2(pe_1_5_0_n63), .B1(
        pe_1_5_0_N82), .B2(pe_1_5_0_n27), .C1(pe_1_5_0_N74), .C2(pe_1_5_0_n28), 
        .ZN(pe_1_5_0_n31) );
  INV_X1 pe_1_5_0_U35 ( .A(pe_1_5_0_n31), .ZN(pe_1_5_0_n79) );
  AOI222_X1 pe_1_5_0_U34 ( .A1(int_data_res_6__0__5_), .A2(pe_1_5_0_n63), .B1(
        pe_1_5_0_N83), .B2(pe_1_5_0_n27), .C1(pe_1_5_0_N75), .C2(pe_1_5_0_n28), 
        .ZN(pe_1_5_0_n30) );
  INV_X1 pe_1_5_0_U33 ( .A(pe_1_5_0_n30), .ZN(pe_1_5_0_n78) );
  NOR3_X1 pe_1_5_0_U32 ( .A1(pe_1_5_0_n59), .A2(pe_1_5_0_n64), .A3(int_ckg[23]), .ZN(pe_1_5_0_n36) );
  OR2_X1 pe_1_5_0_U31 ( .A1(pe_1_5_0_n36), .A2(pe_1_5_0_n63), .ZN(pe_1_5_0_N90) );
  INV_X1 pe_1_5_0_U30 ( .A(pe_1_5_0_int_data_0_), .ZN(pe_1_5_0_n72) );
  INV_X1 pe_1_5_0_U29 ( .A(n40), .ZN(pe_1_5_0_n62) );
  INV_X1 pe_1_5_0_U28 ( .A(n34), .ZN(pe_1_5_0_n60) );
  INV_X1 pe_1_5_0_U27 ( .A(pe_1_5_0_int_data_3_), .ZN(pe_1_5_0_n75) );
  BUF_X1 pe_1_5_0_U26 ( .A(n62), .Z(pe_1_5_0_n63) );
  NAND2_X1 pe_1_5_0_U25 ( .A1(pe_1_5_0_n44), .A2(pe_1_5_0_n60), .ZN(
        pe_1_5_0_n41) );
  AND3_X1 pe_1_5_0_U24 ( .A1(n76), .A2(pe_1_5_0_n62), .A3(n51), .ZN(
        pe_1_5_0_n44) );
  NOR2_X1 pe_1_5_0_U23 ( .A1(pe_1_5_0_n69), .A2(n51), .ZN(pe_1_5_0_n43) );
  NOR2_X1 pe_1_5_0_U22 ( .A1(pe_1_5_0_n57), .A2(pe_1_5_0_n63), .ZN(
        pe_1_5_0_n28) );
  NOR2_X1 pe_1_5_0_U21 ( .A1(n20), .A2(pe_1_5_0_n63), .ZN(pe_1_5_0_n27) );
  INV_X1 pe_1_5_0_U20 ( .A(pe_1_5_0_n41), .ZN(pe_1_5_0_n89) );
  INV_X1 pe_1_5_0_U19 ( .A(pe_1_5_0_n37), .ZN(pe_1_5_0_n87) );
  INV_X1 pe_1_5_0_U18 ( .A(pe_1_5_0_n38), .ZN(pe_1_5_0_n86) );
  INV_X1 pe_1_5_0_U17 ( .A(pe_1_5_0_n39), .ZN(pe_1_5_0_n85) );
  NOR2_X1 pe_1_5_0_U16 ( .A1(pe_1_5_0_n67), .A2(pe_1_5_0_n42), .ZN(
        pe_1_5_0_N59) );
  NOR2_X1 pe_1_5_0_U15 ( .A1(pe_1_5_0_n67), .A2(pe_1_5_0_n41), .ZN(
        pe_1_5_0_N60) );
  NOR2_X1 pe_1_5_0_U14 ( .A1(pe_1_5_0_n67), .A2(pe_1_5_0_n38), .ZN(
        pe_1_5_0_N63) );
  NOR2_X1 pe_1_5_0_U13 ( .A1(pe_1_5_0_n66), .A2(pe_1_5_0_n40), .ZN(
        pe_1_5_0_N61) );
  NOR2_X1 pe_1_5_0_U12 ( .A1(pe_1_5_0_n66), .A2(pe_1_5_0_n39), .ZN(
        pe_1_5_0_N62) );
  NOR2_X1 pe_1_5_0_U11 ( .A1(pe_1_5_0_n37), .A2(pe_1_5_0_n66), .ZN(
        pe_1_5_0_N64) );
  NAND2_X1 pe_1_5_0_U10 ( .A1(pe_1_5_0_n44), .A2(n34), .ZN(pe_1_5_0_n42) );
  BUF_X1 pe_1_5_0_U9 ( .A(n34), .Z(pe_1_5_0_n55) );
  BUF_X1 pe_1_5_0_U8 ( .A(n34), .Z(pe_1_5_0_n56) );
  INV_X1 pe_1_5_0_U7 ( .A(pe_1_5_0_n68), .ZN(pe_1_5_0_n64) );
  INV_X1 pe_1_5_0_U6 ( .A(pe_1_5_0_n42), .ZN(pe_1_5_0_n88) );
  INV_X1 pe_1_5_0_U5 ( .A(pe_1_5_0_n40), .ZN(pe_1_5_0_n84) );
  INV_X2 pe_1_5_0_U4 ( .A(n84), .ZN(pe_1_5_0_n71) );
  XOR2_X1 pe_1_5_0_U3 ( .A(pe_1_5_0_int_data_0_), .B(int_data_res_5__0__0_), 
        .Z(pe_1_5_0_n1) );
  DFFR_X1 pe_1_5_0_int_q_acc_reg_0_ ( .D(pe_1_5_0_n83), .CK(pe_1_5_0_net4432), 
        .RN(pe_1_5_0_n71), .Q(int_data_res_5__0__0_), .QN(pe_1_5_0_n3) );
  DFFR_X1 pe_1_5_0_int_q_reg_v_reg_0__0_ ( .D(int_data_y_6__0__0_), .CK(
        pe_1_5_0_net4402), .RN(pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_v[20]) );
  DFFR_X1 pe_1_5_0_int_q_reg_v_reg_0__1_ ( .D(int_data_y_6__0__1_), .CK(
        pe_1_5_0_net4402), .RN(pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_v[21]) );
  DFFR_X1 pe_1_5_0_int_q_reg_v_reg_0__2_ ( .D(int_data_y_6__0__2_), .CK(
        pe_1_5_0_net4402), .RN(pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_v[22]) );
  DFFR_X1 pe_1_5_0_int_q_reg_v_reg_0__3_ ( .D(int_data_y_6__0__3_), .CK(
        pe_1_5_0_net4402), .RN(pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_v[23]) );
  DFFR_X1 pe_1_5_0_int_q_reg_v_reg_1__0_ ( .D(int_data_y_6__0__0_), .CK(
        pe_1_5_0_net4407), .RN(pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_v[16]) );
  DFFR_X1 pe_1_5_0_int_q_reg_v_reg_1__1_ ( .D(int_data_y_6__0__1_), .CK(
        pe_1_5_0_net4407), .RN(pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_v[17]) );
  DFFR_X1 pe_1_5_0_int_q_reg_v_reg_1__2_ ( .D(int_data_y_6__0__2_), .CK(
        pe_1_5_0_net4407), .RN(pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_v[18]) );
  DFFR_X1 pe_1_5_0_int_q_reg_v_reg_1__3_ ( .D(int_data_y_6__0__3_), .CK(
        pe_1_5_0_net4407), .RN(pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_v[19]) );
  DFFR_X1 pe_1_5_0_int_q_reg_v_reg_2__0_ ( .D(int_data_y_6__0__0_), .CK(
        pe_1_5_0_net4412), .RN(pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_v[12]) );
  DFFR_X1 pe_1_5_0_int_q_reg_v_reg_2__1_ ( .D(int_data_y_6__0__1_), .CK(
        pe_1_5_0_net4412), .RN(pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_v[13]) );
  DFFR_X1 pe_1_5_0_int_q_reg_v_reg_2__2_ ( .D(int_data_y_6__0__2_), .CK(
        pe_1_5_0_net4412), .RN(pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_v[14]) );
  DFFR_X1 pe_1_5_0_int_q_reg_v_reg_2__3_ ( .D(int_data_y_6__0__3_), .CK(
        pe_1_5_0_net4412), .RN(pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_v[15]) );
  DFFR_X1 pe_1_5_0_int_q_reg_v_reg_3__0_ ( .D(int_data_y_6__0__0_), .CK(
        pe_1_5_0_net4417), .RN(pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_v[8]) );
  DFFR_X1 pe_1_5_0_int_q_reg_v_reg_3__1_ ( .D(int_data_y_6__0__1_), .CK(
        pe_1_5_0_net4417), .RN(pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_v[9]) );
  DFFR_X1 pe_1_5_0_int_q_reg_v_reg_3__2_ ( .D(int_data_y_6__0__2_), .CK(
        pe_1_5_0_net4417), .RN(pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_v[10]) );
  DFFR_X1 pe_1_5_0_int_q_reg_v_reg_3__3_ ( .D(int_data_y_6__0__3_), .CK(
        pe_1_5_0_net4417), .RN(pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_v[11]) );
  DFFR_X1 pe_1_5_0_int_q_reg_v_reg_4__0_ ( .D(int_data_y_6__0__0_), .CK(
        pe_1_5_0_net4422), .RN(pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_v[4]) );
  DFFR_X1 pe_1_5_0_int_q_reg_v_reg_4__1_ ( .D(int_data_y_6__0__1_), .CK(
        pe_1_5_0_net4422), .RN(pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_v[5]) );
  DFFR_X1 pe_1_5_0_int_q_reg_v_reg_4__2_ ( .D(int_data_y_6__0__2_), .CK(
        pe_1_5_0_net4422), .RN(pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_v[6]) );
  DFFR_X1 pe_1_5_0_int_q_reg_v_reg_4__3_ ( .D(int_data_y_6__0__3_), .CK(
        pe_1_5_0_net4422), .RN(pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_v[7]) );
  DFFR_X1 pe_1_5_0_int_q_reg_v_reg_5__0_ ( .D(int_data_y_6__0__0_), .CK(
        pe_1_5_0_net4427), .RN(pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_v[0]) );
  DFFR_X1 pe_1_5_0_int_q_reg_v_reg_5__1_ ( .D(int_data_y_6__0__1_), .CK(
        pe_1_5_0_net4427), .RN(pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_v[1]) );
  DFFR_X1 pe_1_5_0_int_q_reg_v_reg_5__2_ ( .D(int_data_y_6__0__2_), .CK(
        pe_1_5_0_net4427), .RN(pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_v[2]) );
  DFFR_X1 pe_1_5_0_int_q_reg_v_reg_5__3_ ( .D(int_data_y_6__0__3_), .CK(
        pe_1_5_0_net4427), .RN(pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_5_0_int_q_reg_h_reg_0__0_ ( .D(int_data_x_5__1__0_), .SI(
        int_data_y_6__0__0_), .SE(pe_1_5_0_n64), .CK(pe_1_5_0_net4371), .RN(
        pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_5_0_int_q_reg_h_reg_0__1_ ( .D(int_data_x_5__1__1_), .SI(
        int_data_y_6__0__1_), .SE(pe_1_5_0_n64), .CK(pe_1_5_0_net4371), .RN(
        pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_5_0_int_q_reg_h_reg_0__2_ ( .D(int_data_x_5__1__2_), .SI(
        int_data_y_6__0__2_), .SE(pe_1_5_0_n64), .CK(pe_1_5_0_net4371), .RN(
        pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_5_0_int_q_reg_h_reg_0__3_ ( .D(int_data_x_5__1__3_), .SI(
        int_data_y_6__0__3_), .SE(pe_1_5_0_n64), .CK(pe_1_5_0_net4371), .RN(
        pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_5_0_int_q_reg_h_reg_1__0_ ( .D(int_data_x_5__1__0_), .SI(
        int_data_y_6__0__0_), .SE(pe_1_5_0_n64), .CK(pe_1_5_0_net4377), .RN(
        pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_5_0_int_q_reg_h_reg_1__1_ ( .D(int_data_x_5__1__1_), .SI(
        int_data_y_6__0__1_), .SE(pe_1_5_0_n64), .CK(pe_1_5_0_net4377), .RN(
        pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_5_0_int_q_reg_h_reg_1__2_ ( .D(int_data_x_5__1__2_), .SI(
        int_data_y_6__0__2_), .SE(pe_1_5_0_n64), .CK(pe_1_5_0_net4377), .RN(
        pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_5_0_int_q_reg_h_reg_1__3_ ( .D(int_data_x_5__1__3_), .SI(
        int_data_y_6__0__3_), .SE(pe_1_5_0_n64), .CK(pe_1_5_0_net4377), .RN(
        pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_5_0_int_q_reg_h_reg_2__0_ ( .D(int_data_x_5__1__0_), .SI(
        int_data_y_6__0__0_), .SE(pe_1_5_0_n64), .CK(pe_1_5_0_net4382), .RN(
        pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_5_0_int_q_reg_h_reg_2__1_ ( .D(int_data_x_5__1__1_), .SI(
        int_data_y_6__0__1_), .SE(pe_1_5_0_n64), .CK(pe_1_5_0_net4382), .RN(
        pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_5_0_int_q_reg_h_reg_2__2_ ( .D(int_data_x_5__1__2_), .SI(
        int_data_y_6__0__2_), .SE(pe_1_5_0_n64), .CK(pe_1_5_0_net4382), .RN(
        pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_5_0_int_q_reg_h_reg_2__3_ ( .D(int_data_x_5__1__3_), .SI(
        int_data_y_6__0__3_), .SE(pe_1_5_0_n64), .CK(pe_1_5_0_net4382), .RN(
        pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_5_0_int_q_reg_h_reg_3__0_ ( .D(int_data_x_5__1__0_), .SI(
        int_data_y_6__0__0_), .SE(pe_1_5_0_n64), .CK(pe_1_5_0_net4387), .RN(
        pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_5_0_int_q_reg_h_reg_3__1_ ( .D(int_data_x_5__1__1_), .SI(
        int_data_y_6__0__1_), .SE(pe_1_5_0_n64), .CK(pe_1_5_0_net4387), .RN(
        pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_5_0_int_q_reg_h_reg_3__2_ ( .D(int_data_x_5__1__2_), .SI(
        int_data_y_6__0__2_), .SE(pe_1_5_0_n64), .CK(pe_1_5_0_net4387), .RN(
        pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_5_0_int_q_reg_h_reg_3__3_ ( .D(int_data_x_5__1__3_), .SI(
        int_data_y_6__0__3_), .SE(pe_1_5_0_n64), .CK(pe_1_5_0_net4387), .RN(
        pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_5_0_int_q_reg_h_reg_4__0_ ( .D(int_data_x_5__1__0_), .SI(
        int_data_y_6__0__0_), .SE(pe_1_5_0_n65), .CK(pe_1_5_0_net4392), .RN(
        pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_5_0_int_q_reg_h_reg_4__1_ ( .D(int_data_x_5__1__1_), .SI(
        int_data_y_6__0__1_), .SE(pe_1_5_0_n65), .CK(pe_1_5_0_net4392), .RN(
        pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_5_0_int_q_reg_h_reg_4__2_ ( .D(int_data_x_5__1__2_), .SI(
        int_data_y_6__0__2_), .SE(pe_1_5_0_n65), .CK(pe_1_5_0_net4392), .RN(
        pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_5_0_int_q_reg_h_reg_4__3_ ( .D(int_data_x_5__1__3_), .SI(
        int_data_y_6__0__3_), .SE(pe_1_5_0_n65), .CK(pe_1_5_0_net4392), .RN(
        pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_5_0_int_q_reg_h_reg_5__0_ ( .D(int_data_x_5__1__0_), .SI(
        int_data_y_6__0__0_), .SE(pe_1_5_0_n65), .CK(pe_1_5_0_net4397), .RN(
        pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_5_0_int_q_reg_h_reg_5__1_ ( .D(int_data_x_5__1__1_), .SI(
        int_data_y_6__0__1_), .SE(pe_1_5_0_n65), .CK(pe_1_5_0_net4397), .RN(
        pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_5_0_int_q_reg_h_reg_5__2_ ( .D(int_data_x_5__1__2_), .SI(
        int_data_y_6__0__2_), .SE(pe_1_5_0_n65), .CK(pe_1_5_0_net4397), .RN(
        pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_5_0_int_q_reg_h_reg_5__3_ ( .D(int_data_x_5__1__3_), .SI(
        int_data_y_6__0__3_), .SE(pe_1_5_0_n65), .CK(pe_1_5_0_net4397), .RN(
        pe_1_5_0_n71), .Q(pe_1_5_0_int_q_reg_h[3]) );
  FA_X1 pe_1_5_0_sub_81_U2_7 ( .A(int_data_res_5__0__7_), .B(pe_1_5_0_n75), 
        .CI(pe_1_5_0_sub_81_carry[7]), .S(pe_1_5_0_N77) );
  FA_X1 pe_1_5_0_sub_81_U2_6 ( .A(int_data_res_5__0__6_), .B(pe_1_5_0_n75), 
        .CI(pe_1_5_0_sub_81_carry[6]), .CO(pe_1_5_0_sub_81_carry[7]), .S(
        pe_1_5_0_N76) );
  FA_X1 pe_1_5_0_sub_81_U2_5 ( .A(int_data_res_5__0__5_), .B(pe_1_5_0_n75), 
        .CI(pe_1_5_0_sub_81_carry[5]), .CO(pe_1_5_0_sub_81_carry[6]), .S(
        pe_1_5_0_N75) );
  FA_X1 pe_1_5_0_sub_81_U2_4 ( .A(int_data_res_5__0__4_), .B(pe_1_5_0_n75), 
        .CI(pe_1_5_0_sub_81_carry[4]), .CO(pe_1_5_0_sub_81_carry[5]), .S(
        pe_1_5_0_N74) );
  FA_X1 pe_1_5_0_sub_81_U2_3 ( .A(int_data_res_5__0__3_), .B(pe_1_5_0_n75), 
        .CI(pe_1_5_0_sub_81_carry[3]), .CO(pe_1_5_0_sub_81_carry[4]), .S(
        pe_1_5_0_N73) );
  FA_X1 pe_1_5_0_sub_81_U2_2 ( .A(int_data_res_5__0__2_), .B(pe_1_5_0_n74), 
        .CI(pe_1_5_0_sub_81_carry[2]), .CO(pe_1_5_0_sub_81_carry[3]), .S(
        pe_1_5_0_N72) );
  FA_X1 pe_1_5_0_sub_81_U2_1 ( .A(int_data_res_5__0__1_), .B(pe_1_5_0_n73), 
        .CI(pe_1_5_0_sub_81_carry[1]), .CO(pe_1_5_0_sub_81_carry[2]), .S(
        pe_1_5_0_N71) );
  FA_X1 pe_1_5_0_add_83_U1_7 ( .A(int_data_res_5__0__7_), .B(
        pe_1_5_0_int_data_3_), .CI(pe_1_5_0_add_83_carry[7]), .S(pe_1_5_0_N85)
         );
  FA_X1 pe_1_5_0_add_83_U1_6 ( .A(int_data_res_5__0__6_), .B(
        pe_1_5_0_int_data_3_), .CI(pe_1_5_0_add_83_carry[6]), .CO(
        pe_1_5_0_add_83_carry[7]), .S(pe_1_5_0_N84) );
  FA_X1 pe_1_5_0_add_83_U1_5 ( .A(int_data_res_5__0__5_), .B(
        pe_1_5_0_int_data_3_), .CI(pe_1_5_0_add_83_carry[5]), .CO(
        pe_1_5_0_add_83_carry[6]), .S(pe_1_5_0_N83) );
  FA_X1 pe_1_5_0_add_83_U1_4 ( .A(int_data_res_5__0__4_), .B(
        pe_1_5_0_int_data_3_), .CI(pe_1_5_0_add_83_carry[4]), .CO(
        pe_1_5_0_add_83_carry[5]), .S(pe_1_5_0_N82) );
  FA_X1 pe_1_5_0_add_83_U1_3 ( .A(int_data_res_5__0__3_), .B(
        pe_1_5_0_int_data_3_), .CI(pe_1_5_0_add_83_carry[3]), .CO(
        pe_1_5_0_add_83_carry[4]), .S(pe_1_5_0_N81) );
  FA_X1 pe_1_5_0_add_83_U1_2 ( .A(int_data_res_5__0__2_), .B(
        pe_1_5_0_int_data_2_), .CI(pe_1_5_0_add_83_carry[2]), .CO(
        pe_1_5_0_add_83_carry[3]), .S(pe_1_5_0_N80) );
  FA_X1 pe_1_5_0_add_83_U1_1 ( .A(int_data_res_5__0__1_), .B(
        pe_1_5_0_int_data_1_), .CI(pe_1_5_0_n2), .CO(pe_1_5_0_add_83_carry[2]), 
        .S(pe_1_5_0_N79) );
  NAND3_X1 pe_1_5_0_U56 ( .A1(n34), .A2(pe_1_5_0_n43), .A3(pe_1_5_0_n61), .ZN(
        pe_1_5_0_n40) );
  NAND3_X1 pe_1_5_0_U55 ( .A1(pe_1_5_0_n43), .A2(pe_1_5_0_n60), .A3(
        pe_1_5_0_n61), .ZN(pe_1_5_0_n39) );
  NAND3_X1 pe_1_5_0_U54 ( .A1(pe_1_5_0_n43), .A2(pe_1_5_0_n62), .A3(n34), .ZN(
        pe_1_5_0_n38) );
  NAND3_X1 pe_1_5_0_U53 ( .A1(pe_1_5_0_n60), .A2(pe_1_5_0_n62), .A3(
        pe_1_5_0_n43), .ZN(pe_1_5_0_n37) );
  DFFR_X1 pe_1_5_0_int_q_acc_reg_6_ ( .D(pe_1_5_0_n77), .CK(pe_1_5_0_net4432), 
        .RN(pe_1_5_0_n70), .Q(int_data_res_5__0__6_) );
  DFFR_X1 pe_1_5_0_int_q_acc_reg_5_ ( .D(pe_1_5_0_n78), .CK(pe_1_5_0_net4432), 
        .RN(pe_1_5_0_n70), .Q(int_data_res_5__0__5_) );
  DFFR_X1 pe_1_5_0_int_q_acc_reg_4_ ( .D(pe_1_5_0_n79), .CK(pe_1_5_0_net4432), 
        .RN(pe_1_5_0_n70), .Q(int_data_res_5__0__4_) );
  DFFR_X1 pe_1_5_0_int_q_acc_reg_3_ ( .D(pe_1_5_0_n80), .CK(pe_1_5_0_net4432), 
        .RN(pe_1_5_0_n70), .Q(int_data_res_5__0__3_) );
  DFFR_X1 pe_1_5_0_int_q_acc_reg_2_ ( .D(pe_1_5_0_n81), .CK(pe_1_5_0_net4432), 
        .RN(pe_1_5_0_n70), .Q(int_data_res_5__0__2_) );
  DFFR_X1 pe_1_5_0_int_q_acc_reg_1_ ( .D(pe_1_5_0_n82), .CK(pe_1_5_0_net4432), 
        .RN(pe_1_5_0_n70), .Q(int_data_res_5__0__1_) );
  DFFR_X1 pe_1_5_0_int_q_acc_reg_7_ ( .D(pe_1_5_0_n76), .CK(pe_1_5_0_net4432), 
        .RN(pe_1_5_0_n70), .Q(int_data_res_5__0__7_) );
  CLKGATETST_X1 pe_1_5_0_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_5_0_n87), .SE(1'b0), .GCK(pe_1_5_0_net4371) );
  CLKGATETST_X1 pe_1_5_0_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_5_0_n86), .SE(1'b0), .GCK(pe_1_5_0_net4377) );
  CLKGATETST_X1 pe_1_5_0_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_5_0_n85), .SE(1'b0), .GCK(pe_1_5_0_net4382) );
  CLKGATETST_X1 pe_1_5_0_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_5_0_n84), .SE(1'b0), .GCK(pe_1_5_0_net4387) );
  CLKGATETST_X1 pe_1_5_0_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_5_0_n89), .SE(1'b0), .GCK(pe_1_5_0_net4392) );
  CLKGATETST_X1 pe_1_5_0_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_5_0_n88), .SE(1'b0), .GCK(pe_1_5_0_net4397) );
  CLKGATETST_X1 pe_1_5_0_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_5_0_N64), .SE(1'b0), .GCK(pe_1_5_0_net4402) );
  CLKGATETST_X1 pe_1_5_0_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_5_0_N63), .SE(1'b0), .GCK(pe_1_5_0_net4407) );
  CLKGATETST_X1 pe_1_5_0_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_5_0_N62), .SE(1'b0), .GCK(pe_1_5_0_net4412) );
  CLKGATETST_X1 pe_1_5_0_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_5_0_N61), .SE(1'b0), .GCK(pe_1_5_0_net4417) );
  CLKGATETST_X1 pe_1_5_0_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_5_0_N60), .SE(1'b0), .GCK(pe_1_5_0_net4422) );
  CLKGATETST_X1 pe_1_5_0_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_5_0_N59), .SE(1'b0), .GCK(pe_1_5_0_net4427) );
  CLKGATETST_X1 pe_1_5_0_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_5_0_N90), .SE(1'b0), .GCK(pe_1_5_0_net4432) );
  CLKBUF_X1 pe_1_5_1_U112 ( .A(pe_1_5_1_n72), .Z(pe_1_5_1_n71) );
  INV_X1 pe_1_5_1_U111 ( .A(n76), .ZN(pe_1_5_1_n70) );
  INV_X1 pe_1_5_1_U110 ( .A(n68), .ZN(pe_1_5_1_n69) );
  INV_X1 pe_1_5_1_U109 ( .A(n68), .ZN(pe_1_5_1_n68) );
  INV_X1 pe_1_5_1_U108 ( .A(n68), .ZN(pe_1_5_1_n67) );
  INV_X1 pe_1_5_1_U107 ( .A(pe_1_5_1_n69), .ZN(pe_1_5_1_n66) );
  INV_X1 pe_1_5_1_U106 ( .A(pe_1_5_1_n63), .ZN(pe_1_5_1_n62) );
  INV_X1 pe_1_5_1_U105 ( .A(pe_1_5_1_n61), .ZN(pe_1_5_1_n60) );
  INV_X1 pe_1_5_1_U104 ( .A(n28), .ZN(pe_1_5_1_n59) );
  INV_X1 pe_1_5_1_U103 ( .A(pe_1_5_1_n59), .ZN(pe_1_5_1_n58) );
  INV_X1 pe_1_5_1_U102 ( .A(n20), .ZN(pe_1_5_1_n57) );
  MUX2_X1 pe_1_5_1_U101 ( .A(pe_1_5_1_n54), .B(pe_1_5_1_n51), .S(n51), .Z(
        int_data_x_5__1__3_) );
  MUX2_X1 pe_1_5_1_U100 ( .A(pe_1_5_1_n53), .B(pe_1_5_1_n52), .S(pe_1_5_1_n62), 
        .Z(pe_1_5_1_n54) );
  MUX2_X1 pe_1_5_1_U99 ( .A(pe_1_5_1_int_q_reg_h[23]), .B(
        pe_1_5_1_int_q_reg_h[19]), .S(pe_1_5_1_n56), .Z(pe_1_5_1_n53) );
  MUX2_X1 pe_1_5_1_U98 ( .A(pe_1_5_1_int_q_reg_h[15]), .B(
        pe_1_5_1_int_q_reg_h[11]), .S(pe_1_5_1_n56), .Z(pe_1_5_1_n52) );
  MUX2_X1 pe_1_5_1_U97 ( .A(pe_1_5_1_int_q_reg_h[7]), .B(
        pe_1_5_1_int_q_reg_h[3]), .S(pe_1_5_1_n56), .Z(pe_1_5_1_n51) );
  MUX2_X1 pe_1_5_1_U96 ( .A(pe_1_5_1_n50), .B(pe_1_5_1_n47), .S(n51), .Z(
        int_data_x_5__1__2_) );
  MUX2_X1 pe_1_5_1_U95 ( .A(pe_1_5_1_n49), .B(pe_1_5_1_n48), .S(pe_1_5_1_n62), 
        .Z(pe_1_5_1_n50) );
  MUX2_X1 pe_1_5_1_U94 ( .A(pe_1_5_1_int_q_reg_h[22]), .B(
        pe_1_5_1_int_q_reg_h[18]), .S(pe_1_5_1_n56), .Z(pe_1_5_1_n49) );
  MUX2_X1 pe_1_5_1_U93 ( .A(pe_1_5_1_int_q_reg_h[14]), .B(
        pe_1_5_1_int_q_reg_h[10]), .S(pe_1_5_1_n56), .Z(pe_1_5_1_n48) );
  MUX2_X1 pe_1_5_1_U92 ( .A(pe_1_5_1_int_q_reg_h[6]), .B(
        pe_1_5_1_int_q_reg_h[2]), .S(pe_1_5_1_n56), .Z(pe_1_5_1_n47) );
  MUX2_X1 pe_1_5_1_U91 ( .A(pe_1_5_1_n46), .B(pe_1_5_1_n24), .S(n51), .Z(
        int_data_x_5__1__1_) );
  MUX2_X1 pe_1_5_1_U90 ( .A(pe_1_5_1_n45), .B(pe_1_5_1_n25), .S(pe_1_5_1_n62), 
        .Z(pe_1_5_1_n46) );
  MUX2_X1 pe_1_5_1_U89 ( .A(pe_1_5_1_int_q_reg_h[21]), .B(
        pe_1_5_1_int_q_reg_h[17]), .S(pe_1_5_1_n56), .Z(pe_1_5_1_n45) );
  MUX2_X1 pe_1_5_1_U88 ( .A(pe_1_5_1_int_q_reg_h[13]), .B(
        pe_1_5_1_int_q_reg_h[9]), .S(pe_1_5_1_n56), .Z(pe_1_5_1_n25) );
  MUX2_X1 pe_1_5_1_U87 ( .A(pe_1_5_1_int_q_reg_h[5]), .B(
        pe_1_5_1_int_q_reg_h[1]), .S(pe_1_5_1_n56), .Z(pe_1_5_1_n24) );
  MUX2_X1 pe_1_5_1_U86 ( .A(pe_1_5_1_n23), .B(pe_1_5_1_n20), .S(n51), .Z(
        int_data_x_5__1__0_) );
  MUX2_X1 pe_1_5_1_U85 ( .A(pe_1_5_1_n22), .B(pe_1_5_1_n21), .S(pe_1_5_1_n62), 
        .Z(pe_1_5_1_n23) );
  MUX2_X1 pe_1_5_1_U84 ( .A(pe_1_5_1_int_q_reg_h[20]), .B(
        pe_1_5_1_int_q_reg_h[16]), .S(pe_1_5_1_n56), .Z(pe_1_5_1_n22) );
  MUX2_X1 pe_1_5_1_U83 ( .A(pe_1_5_1_int_q_reg_h[12]), .B(
        pe_1_5_1_int_q_reg_h[8]), .S(pe_1_5_1_n56), .Z(pe_1_5_1_n21) );
  MUX2_X1 pe_1_5_1_U82 ( .A(pe_1_5_1_int_q_reg_h[4]), .B(
        pe_1_5_1_int_q_reg_h[0]), .S(pe_1_5_1_n56), .Z(pe_1_5_1_n20) );
  MUX2_X1 pe_1_5_1_U81 ( .A(pe_1_5_1_n19), .B(pe_1_5_1_n16), .S(n51), .Z(
        int_data_y_5__1__3_) );
  MUX2_X1 pe_1_5_1_U80 ( .A(pe_1_5_1_n18), .B(pe_1_5_1_n17), .S(pe_1_5_1_n62), 
        .Z(pe_1_5_1_n19) );
  MUX2_X1 pe_1_5_1_U79 ( .A(pe_1_5_1_int_q_reg_v[23]), .B(
        pe_1_5_1_int_q_reg_v[19]), .S(pe_1_5_1_n55), .Z(pe_1_5_1_n18) );
  MUX2_X1 pe_1_5_1_U78 ( .A(pe_1_5_1_int_q_reg_v[15]), .B(
        pe_1_5_1_int_q_reg_v[11]), .S(pe_1_5_1_n55), .Z(pe_1_5_1_n17) );
  MUX2_X1 pe_1_5_1_U77 ( .A(pe_1_5_1_int_q_reg_v[7]), .B(
        pe_1_5_1_int_q_reg_v[3]), .S(pe_1_5_1_n55), .Z(pe_1_5_1_n16) );
  MUX2_X1 pe_1_5_1_U76 ( .A(pe_1_5_1_n15), .B(pe_1_5_1_n12), .S(n51), .Z(
        int_data_y_5__1__2_) );
  MUX2_X1 pe_1_5_1_U75 ( .A(pe_1_5_1_n14), .B(pe_1_5_1_n13), .S(pe_1_5_1_n62), 
        .Z(pe_1_5_1_n15) );
  MUX2_X1 pe_1_5_1_U74 ( .A(pe_1_5_1_int_q_reg_v[22]), .B(
        pe_1_5_1_int_q_reg_v[18]), .S(pe_1_5_1_n55), .Z(pe_1_5_1_n14) );
  MUX2_X1 pe_1_5_1_U73 ( .A(pe_1_5_1_int_q_reg_v[14]), .B(
        pe_1_5_1_int_q_reg_v[10]), .S(pe_1_5_1_n55), .Z(pe_1_5_1_n13) );
  MUX2_X1 pe_1_5_1_U72 ( .A(pe_1_5_1_int_q_reg_v[6]), .B(
        pe_1_5_1_int_q_reg_v[2]), .S(pe_1_5_1_n55), .Z(pe_1_5_1_n12) );
  MUX2_X1 pe_1_5_1_U71 ( .A(pe_1_5_1_n11), .B(pe_1_5_1_n8), .S(n51), .Z(
        int_data_y_5__1__1_) );
  MUX2_X1 pe_1_5_1_U70 ( .A(pe_1_5_1_n10), .B(pe_1_5_1_n9), .S(pe_1_5_1_n62), 
        .Z(pe_1_5_1_n11) );
  MUX2_X1 pe_1_5_1_U69 ( .A(pe_1_5_1_int_q_reg_v[21]), .B(
        pe_1_5_1_int_q_reg_v[17]), .S(pe_1_5_1_n55), .Z(pe_1_5_1_n10) );
  MUX2_X1 pe_1_5_1_U68 ( .A(pe_1_5_1_int_q_reg_v[13]), .B(
        pe_1_5_1_int_q_reg_v[9]), .S(pe_1_5_1_n55), .Z(pe_1_5_1_n9) );
  MUX2_X1 pe_1_5_1_U67 ( .A(pe_1_5_1_int_q_reg_v[5]), .B(
        pe_1_5_1_int_q_reg_v[1]), .S(pe_1_5_1_n55), .Z(pe_1_5_1_n8) );
  MUX2_X1 pe_1_5_1_U66 ( .A(pe_1_5_1_n7), .B(pe_1_5_1_n4), .S(n51), .Z(
        int_data_y_5__1__0_) );
  MUX2_X1 pe_1_5_1_U65 ( .A(pe_1_5_1_n6), .B(pe_1_5_1_n5), .S(pe_1_5_1_n62), 
        .Z(pe_1_5_1_n7) );
  MUX2_X1 pe_1_5_1_U64 ( .A(pe_1_5_1_int_q_reg_v[20]), .B(
        pe_1_5_1_int_q_reg_v[16]), .S(pe_1_5_1_n55), .Z(pe_1_5_1_n6) );
  MUX2_X1 pe_1_5_1_U63 ( .A(pe_1_5_1_int_q_reg_v[12]), .B(
        pe_1_5_1_int_q_reg_v[8]), .S(pe_1_5_1_n55), .Z(pe_1_5_1_n5) );
  MUX2_X1 pe_1_5_1_U62 ( .A(pe_1_5_1_int_q_reg_v[4]), .B(
        pe_1_5_1_int_q_reg_v[0]), .S(pe_1_5_1_n55), .Z(pe_1_5_1_n4) );
  AOI222_X1 pe_1_5_1_U61 ( .A1(int_data_res_6__1__2_), .A2(pe_1_5_1_n64), .B1(
        pe_1_5_1_N80), .B2(pe_1_5_1_n27), .C1(pe_1_5_1_N72), .C2(pe_1_5_1_n28), 
        .ZN(pe_1_5_1_n33) );
  INV_X1 pe_1_5_1_U60 ( .A(pe_1_5_1_n33), .ZN(pe_1_5_1_n82) );
  AOI222_X1 pe_1_5_1_U59 ( .A1(int_data_res_6__1__6_), .A2(pe_1_5_1_n64), .B1(
        pe_1_5_1_N84), .B2(pe_1_5_1_n27), .C1(pe_1_5_1_N76), .C2(pe_1_5_1_n28), 
        .ZN(pe_1_5_1_n29) );
  INV_X1 pe_1_5_1_U58 ( .A(pe_1_5_1_n29), .ZN(pe_1_5_1_n78) );
  XNOR2_X1 pe_1_5_1_U57 ( .A(pe_1_5_1_n73), .B(int_data_res_5__1__0_), .ZN(
        pe_1_5_1_N70) );
  AOI222_X1 pe_1_5_1_U52 ( .A1(int_data_res_6__1__0_), .A2(pe_1_5_1_n64), .B1(
        pe_1_5_1_n1), .B2(pe_1_5_1_n27), .C1(pe_1_5_1_N70), .C2(pe_1_5_1_n28), 
        .ZN(pe_1_5_1_n35) );
  INV_X1 pe_1_5_1_U51 ( .A(pe_1_5_1_n35), .ZN(pe_1_5_1_n84) );
  AOI222_X1 pe_1_5_1_U50 ( .A1(int_data_res_6__1__1_), .A2(pe_1_5_1_n64), .B1(
        pe_1_5_1_N79), .B2(pe_1_5_1_n27), .C1(pe_1_5_1_N71), .C2(pe_1_5_1_n28), 
        .ZN(pe_1_5_1_n34) );
  INV_X1 pe_1_5_1_U49 ( .A(pe_1_5_1_n34), .ZN(pe_1_5_1_n83) );
  AOI222_X1 pe_1_5_1_U48 ( .A1(int_data_res_6__1__3_), .A2(pe_1_5_1_n64), .B1(
        pe_1_5_1_N81), .B2(pe_1_5_1_n27), .C1(pe_1_5_1_N73), .C2(pe_1_5_1_n28), 
        .ZN(pe_1_5_1_n32) );
  INV_X1 pe_1_5_1_U47 ( .A(pe_1_5_1_n32), .ZN(pe_1_5_1_n81) );
  AOI222_X1 pe_1_5_1_U46 ( .A1(int_data_res_6__1__4_), .A2(pe_1_5_1_n64), .B1(
        pe_1_5_1_N82), .B2(pe_1_5_1_n27), .C1(pe_1_5_1_N74), .C2(pe_1_5_1_n28), 
        .ZN(pe_1_5_1_n31) );
  INV_X1 pe_1_5_1_U45 ( .A(pe_1_5_1_n31), .ZN(pe_1_5_1_n80) );
  AOI222_X1 pe_1_5_1_U44 ( .A1(int_data_res_6__1__5_), .A2(pe_1_5_1_n64), .B1(
        pe_1_5_1_N83), .B2(pe_1_5_1_n27), .C1(pe_1_5_1_N75), .C2(pe_1_5_1_n28), 
        .ZN(pe_1_5_1_n30) );
  INV_X1 pe_1_5_1_U43 ( .A(pe_1_5_1_n30), .ZN(pe_1_5_1_n79) );
  NAND2_X1 pe_1_5_1_U42 ( .A1(pe_1_5_1_int_data_0_), .A2(pe_1_5_1_n3), .ZN(
        pe_1_5_1_sub_81_carry[1]) );
  INV_X1 pe_1_5_1_U41 ( .A(pe_1_5_1_int_data_1_), .ZN(pe_1_5_1_n74) );
  INV_X1 pe_1_5_1_U40 ( .A(pe_1_5_1_int_data_2_), .ZN(pe_1_5_1_n75) );
  AND2_X1 pe_1_5_1_U39 ( .A1(pe_1_5_1_int_data_0_), .A2(int_data_res_5__1__0_), 
        .ZN(pe_1_5_1_n2) );
  AOI222_X1 pe_1_5_1_U38 ( .A1(pe_1_5_1_n64), .A2(int_data_res_6__1__7_), .B1(
        pe_1_5_1_N85), .B2(pe_1_5_1_n27), .C1(pe_1_5_1_N77), .C2(pe_1_5_1_n28), 
        .ZN(pe_1_5_1_n26) );
  INV_X1 pe_1_5_1_U37 ( .A(pe_1_5_1_n26), .ZN(pe_1_5_1_n77) );
  NOR3_X1 pe_1_5_1_U36 ( .A1(pe_1_5_1_n59), .A2(pe_1_5_1_n65), .A3(int_ckg[22]), .ZN(pe_1_5_1_n36) );
  OR2_X1 pe_1_5_1_U35 ( .A1(pe_1_5_1_n36), .A2(pe_1_5_1_n64), .ZN(pe_1_5_1_N90) );
  INV_X1 pe_1_5_1_U34 ( .A(n40), .ZN(pe_1_5_1_n63) );
  AND2_X1 pe_1_5_1_U33 ( .A1(int_data_x_5__1__2_), .A2(pe_1_5_1_n58), .ZN(
        pe_1_5_1_int_data_2_) );
  AND2_X1 pe_1_5_1_U32 ( .A1(int_data_x_5__1__1_), .A2(pe_1_5_1_n58), .ZN(
        pe_1_5_1_int_data_1_) );
  AND2_X1 pe_1_5_1_U31 ( .A1(int_data_x_5__1__3_), .A2(pe_1_5_1_n58), .ZN(
        pe_1_5_1_int_data_3_) );
  BUF_X1 pe_1_5_1_U30 ( .A(n62), .Z(pe_1_5_1_n64) );
  INV_X1 pe_1_5_1_U29 ( .A(n34), .ZN(pe_1_5_1_n61) );
  AND2_X1 pe_1_5_1_U28 ( .A1(int_data_x_5__1__0_), .A2(pe_1_5_1_n58), .ZN(
        pe_1_5_1_int_data_0_) );
  NAND2_X1 pe_1_5_1_U27 ( .A1(pe_1_5_1_n44), .A2(pe_1_5_1_n61), .ZN(
        pe_1_5_1_n41) );
  AND3_X1 pe_1_5_1_U26 ( .A1(n76), .A2(pe_1_5_1_n63), .A3(n51), .ZN(
        pe_1_5_1_n44) );
  INV_X1 pe_1_5_1_U25 ( .A(pe_1_5_1_int_data_3_), .ZN(pe_1_5_1_n76) );
  NOR2_X1 pe_1_5_1_U24 ( .A1(pe_1_5_1_n70), .A2(n51), .ZN(pe_1_5_1_n43) );
  NOR2_X1 pe_1_5_1_U23 ( .A1(pe_1_5_1_n57), .A2(pe_1_5_1_n64), .ZN(
        pe_1_5_1_n28) );
  NOR2_X1 pe_1_5_1_U22 ( .A1(n20), .A2(pe_1_5_1_n64), .ZN(pe_1_5_1_n27) );
  INV_X1 pe_1_5_1_U21 ( .A(pe_1_5_1_int_data_0_), .ZN(pe_1_5_1_n73) );
  INV_X1 pe_1_5_1_U20 ( .A(pe_1_5_1_n41), .ZN(pe_1_5_1_n90) );
  INV_X1 pe_1_5_1_U19 ( .A(pe_1_5_1_n37), .ZN(pe_1_5_1_n88) );
  INV_X1 pe_1_5_1_U18 ( .A(pe_1_5_1_n38), .ZN(pe_1_5_1_n87) );
  INV_X1 pe_1_5_1_U17 ( .A(pe_1_5_1_n39), .ZN(pe_1_5_1_n86) );
  NOR2_X1 pe_1_5_1_U16 ( .A1(pe_1_5_1_n68), .A2(pe_1_5_1_n42), .ZN(
        pe_1_5_1_N59) );
  NOR2_X1 pe_1_5_1_U15 ( .A1(pe_1_5_1_n68), .A2(pe_1_5_1_n41), .ZN(
        pe_1_5_1_N60) );
  NOR2_X1 pe_1_5_1_U14 ( .A1(pe_1_5_1_n68), .A2(pe_1_5_1_n38), .ZN(
        pe_1_5_1_N63) );
  NOR2_X1 pe_1_5_1_U13 ( .A1(pe_1_5_1_n67), .A2(pe_1_5_1_n40), .ZN(
        pe_1_5_1_N61) );
  NOR2_X1 pe_1_5_1_U12 ( .A1(pe_1_5_1_n67), .A2(pe_1_5_1_n39), .ZN(
        pe_1_5_1_N62) );
  NOR2_X1 pe_1_5_1_U11 ( .A1(pe_1_5_1_n37), .A2(pe_1_5_1_n67), .ZN(
        pe_1_5_1_N64) );
  NAND2_X1 pe_1_5_1_U10 ( .A1(pe_1_5_1_n44), .A2(pe_1_5_1_n60), .ZN(
        pe_1_5_1_n42) );
  BUF_X1 pe_1_5_1_U9 ( .A(pe_1_5_1_n60), .Z(pe_1_5_1_n55) );
  INV_X1 pe_1_5_1_U8 ( .A(pe_1_5_1_n69), .ZN(pe_1_5_1_n65) );
  BUF_X1 pe_1_5_1_U7 ( .A(pe_1_5_1_n60), .Z(pe_1_5_1_n56) );
  INV_X1 pe_1_5_1_U6 ( .A(pe_1_5_1_n42), .ZN(pe_1_5_1_n89) );
  INV_X1 pe_1_5_1_U5 ( .A(pe_1_5_1_n40), .ZN(pe_1_5_1_n85) );
  INV_X2 pe_1_5_1_U4 ( .A(n84), .ZN(pe_1_5_1_n72) );
  XOR2_X1 pe_1_5_1_U3 ( .A(pe_1_5_1_int_data_0_), .B(int_data_res_5__1__0_), 
        .Z(pe_1_5_1_n1) );
  DFFR_X1 pe_1_5_1_int_q_acc_reg_0_ ( .D(pe_1_5_1_n84), .CK(pe_1_5_1_net4354), 
        .RN(pe_1_5_1_n72), .Q(int_data_res_5__1__0_), .QN(pe_1_5_1_n3) );
  DFFR_X1 pe_1_5_1_int_q_reg_v_reg_0__0_ ( .D(int_data_y_6__1__0_), .CK(
        pe_1_5_1_net4324), .RN(pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_v[20]) );
  DFFR_X1 pe_1_5_1_int_q_reg_v_reg_0__1_ ( .D(int_data_y_6__1__1_), .CK(
        pe_1_5_1_net4324), .RN(pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_v[21]) );
  DFFR_X1 pe_1_5_1_int_q_reg_v_reg_0__2_ ( .D(int_data_y_6__1__2_), .CK(
        pe_1_5_1_net4324), .RN(pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_v[22]) );
  DFFR_X1 pe_1_5_1_int_q_reg_v_reg_0__3_ ( .D(int_data_y_6__1__3_), .CK(
        pe_1_5_1_net4324), .RN(pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_v[23]) );
  DFFR_X1 pe_1_5_1_int_q_reg_v_reg_1__0_ ( .D(int_data_y_6__1__0_), .CK(
        pe_1_5_1_net4329), .RN(pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_v[16]) );
  DFFR_X1 pe_1_5_1_int_q_reg_v_reg_1__1_ ( .D(int_data_y_6__1__1_), .CK(
        pe_1_5_1_net4329), .RN(pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_v[17]) );
  DFFR_X1 pe_1_5_1_int_q_reg_v_reg_1__2_ ( .D(int_data_y_6__1__2_), .CK(
        pe_1_5_1_net4329), .RN(pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_v[18]) );
  DFFR_X1 pe_1_5_1_int_q_reg_v_reg_1__3_ ( .D(int_data_y_6__1__3_), .CK(
        pe_1_5_1_net4329), .RN(pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_v[19]) );
  DFFR_X1 pe_1_5_1_int_q_reg_v_reg_2__0_ ( .D(int_data_y_6__1__0_), .CK(
        pe_1_5_1_net4334), .RN(pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_v[12]) );
  DFFR_X1 pe_1_5_1_int_q_reg_v_reg_2__1_ ( .D(int_data_y_6__1__1_), .CK(
        pe_1_5_1_net4334), .RN(pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_v[13]) );
  DFFR_X1 pe_1_5_1_int_q_reg_v_reg_2__2_ ( .D(int_data_y_6__1__2_), .CK(
        pe_1_5_1_net4334), .RN(pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_v[14]) );
  DFFR_X1 pe_1_5_1_int_q_reg_v_reg_2__3_ ( .D(int_data_y_6__1__3_), .CK(
        pe_1_5_1_net4334), .RN(pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_v[15]) );
  DFFR_X1 pe_1_5_1_int_q_reg_v_reg_3__0_ ( .D(int_data_y_6__1__0_), .CK(
        pe_1_5_1_net4339), .RN(pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_v[8]) );
  DFFR_X1 pe_1_5_1_int_q_reg_v_reg_3__1_ ( .D(int_data_y_6__1__1_), .CK(
        pe_1_5_1_net4339), .RN(pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_v[9]) );
  DFFR_X1 pe_1_5_1_int_q_reg_v_reg_3__2_ ( .D(int_data_y_6__1__2_), .CK(
        pe_1_5_1_net4339), .RN(pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_v[10]) );
  DFFR_X1 pe_1_5_1_int_q_reg_v_reg_3__3_ ( .D(int_data_y_6__1__3_), .CK(
        pe_1_5_1_net4339), .RN(pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_v[11]) );
  DFFR_X1 pe_1_5_1_int_q_reg_v_reg_4__0_ ( .D(int_data_y_6__1__0_), .CK(
        pe_1_5_1_net4344), .RN(pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_v[4]) );
  DFFR_X1 pe_1_5_1_int_q_reg_v_reg_4__1_ ( .D(int_data_y_6__1__1_), .CK(
        pe_1_5_1_net4344), .RN(pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_v[5]) );
  DFFR_X1 pe_1_5_1_int_q_reg_v_reg_4__2_ ( .D(int_data_y_6__1__2_), .CK(
        pe_1_5_1_net4344), .RN(pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_v[6]) );
  DFFR_X1 pe_1_5_1_int_q_reg_v_reg_4__3_ ( .D(int_data_y_6__1__3_), .CK(
        pe_1_5_1_net4344), .RN(pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_v[7]) );
  DFFR_X1 pe_1_5_1_int_q_reg_v_reg_5__0_ ( .D(int_data_y_6__1__0_), .CK(
        pe_1_5_1_net4349), .RN(pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_v[0]) );
  DFFR_X1 pe_1_5_1_int_q_reg_v_reg_5__1_ ( .D(int_data_y_6__1__1_), .CK(
        pe_1_5_1_net4349), .RN(pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_v[1]) );
  DFFR_X1 pe_1_5_1_int_q_reg_v_reg_5__2_ ( .D(int_data_y_6__1__2_), .CK(
        pe_1_5_1_net4349), .RN(pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_v[2]) );
  DFFR_X1 pe_1_5_1_int_q_reg_v_reg_5__3_ ( .D(int_data_y_6__1__3_), .CK(
        pe_1_5_1_net4349), .RN(pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_5_1_int_q_reg_h_reg_0__0_ ( .D(int_data_x_5__2__0_), .SI(
        int_data_y_6__1__0_), .SE(pe_1_5_1_n65), .CK(pe_1_5_1_net4293), .RN(
        pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_5_1_int_q_reg_h_reg_0__1_ ( .D(int_data_x_5__2__1_), .SI(
        int_data_y_6__1__1_), .SE(pe_1_5_1_n65), .CK(pe_1_5_1_net4293), .RN(
        pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_5_1_int_q_reg_h_reg_0__2_ ( .D(int_data_x_5__2__2_), .SI(
        int_data_y_6__1__2_), .SE(pe_1_5_1_n65), .CK(pe_1_5_1_net4293), .RN(
        pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_5_1_int_q_reg_h_reg_0__3_ ( .D(int_data_x_5__2__3_), .SI(
        int_data_y_6__1__3_), .SE(pe_1_5_1_n65), .CK(pe_1_5_1_net4293), .RN(
        pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_5_1_int_q_reg_h_reg_1__0_ ( .D(int_data_x_5__2__0_), .SI(
        int_data_y_6__1__0_), .SE(pe_1_5_1_n65), .CK(pe_1_5_1_net4299), .RN(
        pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_5_1_int_q_reg_h_reg_1__1_ ( .D(int_data_x_5__2__1_), .SI(
        int_data_y_6__1__1_), .SE(pe_1_5_1_n65), .CK(pe_1_5_1_net4299), .RN(
        pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_5_1_int_q_reg_h_reg_1__2_ ( .D(int_data_x_5__2__2_), .SI(
        int_data_y_6__1__2_), .SE(pe_1_5_1_n65), .CK(pe_1_5_1_net4299), .RN(
        pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_5_1_int_q_reg_h_reg_1__3_ ( .D(int_data_x_5__2__3_), .SI(
        int_data_y_6__1__3_), .SE(pe_1_5_1_n65), .CK(pe_1_5_1_net4299), .RN(
        pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_5_1_int_q_reg_h_reg_2__0_ ( .D(int_data_x_5__2__0_), .SI(
        int_data_y_6__1__0_), .SE(pe_1_5_1_n65), .CK(pe_1_5_1_net4304), .RN(
        pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_5_1_int_q_reg_h_reg_2__1_ ( .D(int_data_x_5__2__1_), .SI(
        int_data_y_6__1__1_), .SE(pe_1_5_1_n65), .CK(pe_1_5_1_net4304), .RN(
        pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_5_1_int_q_reg_h_reg_2__2_ ( .D(int_data_x_5__2__2_), .SI(
        int_data_y_6__1__2_), .SE(pe_1_5_1_n65), .CK(pe_1_5_1_net4304), .RN(
        pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_5_1_int_q_reg_h_reg_2__3_ ( .D(int_data_x_5__2__3_), .SI(
        int_data_y_6__1__3_), .SE(pe_1_5_1_n65), .CK(pe_1_5_1_net4304), .RN(
        pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_5_1_int_q_reg_h_reg_3__0_ ( .D(int_data_x_5__2__0_), .SI(
        int_data_y_6__1__0_), .SE(pe_1_5_1_n65), .CK(pe_1_5_1_net4309), .RN(
        pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_5_1_int_q_reg_h_reg_3__1_ ( .D(int_data_x_5__2__1_), .SI(
        int_data_y_6__1__1_), .SE(pe_1_5_1_n65), .CK(pe_1_5_1_net4309), .RN(
        pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_5_1_int_q_reg_h_reg_3__2_ ( .D(int_data_x_5__2__2_), .SI(
        int_data_y_6__1__2_), .SE(pe_1_5_1_n65), .CK(pe_1_5_1_net4309), .RN(
        pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_5_1_int_q_reg_h_reg_3__3_ ( .D(int_data_x_5__2__3_), .SI(
        int_data_y_6__1__3_), .SE(pe_1_5_1_n65), .CK(pe_1_5_1_net4309), .RN(
        pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_5_1_int_q_reg_h_reg_4__0_ ( .D(int_data_x_5__2__0_), .SI(
        int_data_y_6__1__0_), .SE(pe_1_5_1_n66), .CK(pe_1_5_1_net4314), .RN(
        pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_5_1_int_q_reg_h_reg_4__1_ ( .D(int_data_x_5__2__1_), .SI(
        int_data_y_6__1__1_), .SE(pe_1_5_1_n66), .CK(pe_1_5_1_net4314), .RN(
        pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_5_1_int_q_reg_h_reg_4__2_ ( .D(int_data_x_5__2__2_), .SI(
        int_data_y_6__1__2_), .SE(pe_1_5_1_n66), .CK(pe_1_5_1_net4314), .RN(
        pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_5_1_int_q_reg_h_reg_4__3_ ( .D(int_data_x_5__2__3_), .SI(
        int_data_y_6__1__3_), .SE(pe_1_5_1_n66), .CK(pe_1_5_1_net4314), .RN(
        pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_5_1_int_q_reg_h_reg_5__0_ ( .D(int_data_x_5__2__0_), .SI(
        int_data_y_6__1__0_), .SE(pe_1_5_1_n66), .CK(pe_1_5_1_net4319), .RN(
        pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_5_1_int_q_reg_h_reg_5__1_ ( .D(int_data_x_5__2__1_), .SI(
        int_data_y_6__1__1_), .SE(pe_1_5_1_n66), .CK(pe_1_5_1_net4319), .RN(
        pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_5_1_int_q_reg_h_reg_5__2_ ( .D(int_data_x_5__2__2_), .SI(
        int_data_y_6__1__2_), .SE(pe_1_5_1_n66), .CK(pe_1_5_1_net4319), .RN(
        pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_5_1_int_q_reg_h_reg_5__3_ ( .D(int_data_x_5__2__3_), .SI(
        int_data_y_6__1__3_), .SE(pe_1_5_1_n66), .CK(pe_1_5_1_net4319), .RN(
        pe_1_5_1_n72), .Q(pe_1_5_1_int_q_reg_h[3]) );
  FA_X1 pe_1_5_1_sub_81_U2_7 ( .A(int_data_res_5__1__7_), .B(pe_1_5_1_n76), 
        .CI(pe_1_5_1_sub_81_carry[7]), .S(pe_1_5_1_N77) );
  FA_X1 pe_1_5_1_sub_81_U2_6 ( .A(int_data_res_5__1__6_), .B(pe_1_5_1_n76), 
        .CI(pe_1_5_1_sub_81_carry[6]), .CO(pe_1_5_1_sub_81_carry[7]), .S(
        pe_1_5_1_N76) );
  FA_X1 pe_1_5_1_sub_81_U2_5 ( .A(int_data_res_5__1__5_), .B(pe_1_5_1_n76), 
        .CI(pe_1_5_1_sub_81_carry[5]), .CO(pe_1_5_1_sub_81_carry[6]), .S(
        pe_1_5_1_N75) );
  FA_X1 pe_1_5_1_sub_81_U2_4 ( .A(int_data_res_5__1__4_), .B(pe_1_5_1_n76), 
        .CI(pe_1_5_1_sub_81_carry[4]), .CO(pe_1_5_1_sub_81_carry[5]), .S(
        pe_1_5_1_N74) );
  FA_X1 pe_1_5_1_sub_81_U2_3 ( .A(int_data_res_5__1__3_), .B(pe_1_5_1_n76), 
        .CI(pe_1_5_1_sub_81_carry[3]), .CO(pe_1_5_1_sub_81_carry[4]), .S(
        pe_1_5_1_N73) );
  FA_X1 pe_1_5_1_sub_81_U2_2 ( .A(int_data_res_5__1__2_), .B(pe_1_5_1_n75), 
        .CI(pe_1_5_1_sub_81_carry[2]), .CO(pe_1_5_1_sub_81_carry[3]), .S(
        pe_1_5_1_N72) );
  FA_X1 pe_1_5_1_sub_81_U2_1 ( .A(int_data_res_5__1__1_), .B(pe_1_5_1_n74), 
        .CI(pe_1_5_1_sub_81_carry[1]), .CO(pe_1_5_1_sub_81_carry[2]), .S(
        pe_1_5_1_N71) );
  FA_X1 pe_1_5_1_add_83_U1_7 ( .A(int_data_res_5__1__7_), .B(
        pe_1_5_1_int_data_3_), .CI(pe_1_5_1_add_83_carry[7]), .S(pe_1_5_1_N85)
         );
  FA_X1 pe_1_5_1_add_83_U1_6 ( .A(int_data_res_5__1__6_), .B(
        pe_1_5_1_int_data_3_), .CI(pe_1_5_1_add_83_carry[6]), .CO(
        pe_1_5_1_add_83_carry[7]), .S(pe_1_5_1_N84) );
  FA_X1 pe_1_5_1_add_83_U1_5 ( .A(int_data_res_5__1__5_), .B(
        pe_1_5_1_int_data_3_), .CI(pe_1_5_1_add_83_carry[5]), .CO(
        pe_1_5_1_add_83_carry[6]), .S(pe_1_5_1_N83) );
  FA_X1 pe_1_5_1_add_83_U1_4 ( .A(int_data_res_5__1__4_), .B(
        pe_1_5_1_int_data_3_), .CI(pe_1_5_1_add_83_carry[4]), .CO(
        pe_1_5_1_add_83_carry[5]), .S(pe_1_5_1_N82) );
  FA_X1 pe_1_5_1_add_83_U1_3 ( .A(int_data_res_5__1__3_), .B(
        pe_1_5_1_int_data_3_), .CI(pe_1_5_1_add_83_carry[3]), .CO(
        pe_1_5_1_add_83_carry[4]), .S(pe_1_5_1_N81) );
  FA_X1 pe_1_5_1_add_83_U1_2 ( .A(int_data_res_5__1__2_), .B(
        pe_1_5_1_int_data_2_), .CI(pe_1_5_1_add_83_carry[2]), .CO(
        pe_1_5_1_add_83_carry[3]), .S(pe_1_5_1_N80) );
  FA_X1 pe_1_5_1_add_83_U1_1 ( .A(int_data_res_5__1__1_), .B(
        pe_1_5_1_int_data_1_), .CI(pe_1_5_1_n2), .CO(pe_1_5_1_add_83_carry[2]), 
        .S(pe_1_5_1_N79) );
  NAND3_X1 pe_1_5_1_U56 ( .A1(pe_1_5_1_n60), .A2(pe_1_5_1_n43), .A3(
        pe_1_5_1_n62), .ZN(pe_1_5_1_n40) );
  NAND3_X1 pe_1_5_1_U55 ( .A1(pe_1_5_1_n43), .A2(pe_1_5_1_n61), .A3(
        pe_1_5_1_n62), .ZN(pe_1_5_1_n39) );
  NAND3_X1 pe_1_5_1_U54 ( .A1(pe_1_5_1_n43), .A2(pe_1_5_1_n63), .A3(
        pe_1_5_1_n60), .ZN(pe_1_5_1_n38) );
  NAND3_X1 pe_1_5_1_U53 ( .A1(pe_1_5_1_n61), .A2(pe_1_5_1_n63), .A3(
        pe_1_5_1_n43), .ZN(pe_1_5_1_n37) );
  DFFR_X1 pe_1_5_1_int_q_acc_reg_6_ ( .D(pe_1_5_1_n78), .CK(pe_1_5_1_net4354), 
        .RN(pe_1_5_1_n71), .Q(int_data_res_5__1__6_) );
  DFFR_X1 pe_1_5_1_int_q_acc_reg_5_ ( .D(pe_1_5_1_n79), .CK(pe_1_5_1_net4354), 
        .RN(pe_1_5_1_n71), .Q(int_data_res_5__1__5_) );
  DFFR_X1 pe_1_5_1_int_q_acc_reg_4_ ( .D(pe_1_5_1_n80), .CK(pe_1_5_1_net4354), 
        .RN(pe_1_5_1_n71), .Q(int_data_res_5__1__4_) );
  DFFR_X1 pe_1_5_1_int_q_acc_reg_3_ ( .D(pe_1_5_1_n81), .CK(pe_1_5_1_net4354), 
        .RN(pe_1_5_1_n71), .Q(int_data_res_5__1__3_) );
  DFFR_X1 pe_1_5_1_int_q_acc_reg_2_ ( .D(pe_1_5_1_n82), .CK(pe_1_5_1_net4354), 
        .RN(pe_1_5_1_n71), .Q(int_data_res_5__1__2_) );
  DFFR_X1 pe_1_5_1_int_q_acc_reg_1_ ( .D(pe_1_5_1_n83), .CK(pe_1_5_1_net4354), 
        .RN(pe_1_5_1_n71), .Q(int_data_res_5__1__1_) );
  DFFR_X1 pe_1_5_1_int_q_acc_reg_7_ ( .D(pe_1_5_1_n77), .CK(pe_1_5_1_net4354), 
        .RN(pe_1_5_1_n71), .Q(int_data_res_5__1__7_) );
  CLKGATETST_X1 pe_1_5_1_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_5_1_n88), .SE(1'b0), .GCK(pe_1_5_1_net4293) );
  CLKGATETST_X1 pe_1_5_1_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_5_1_n87), .SE(1'b0), .GCK(pe_1_5_1_net4299) );
  CLKGATETST_X1 pe_1_5_1_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_5_1_n86), .SE(1'b0), .GCK(pe_1_5_1_net4304) );
  CLKGATETST_X1 pe_1_5_1_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_5_1_n85), .SE(1'b0), .GCK(pe_1_5_1_net4309) );
  CLKGATETST_X1 pe_1_5_1_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_5_1_n90), .SE(1'b0), .GCK(pe_1_5_1_net4314) );
  CLKGATETST_X1 pe_1_5_1_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_5_1_n89), .SE(1'b0), .GCK(pe_1_5_1_net4319) );
  CLKGATETST_X1 pe_1_5_1_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_5_1_N64), .SE(1'b0), .GCK(pe_1_5_1_net4324) );
  CLKGATETST_X1 pe_1_5_1_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_5_1_N63), .SE(1'b0), .GCK(pe_1_5_1_net4329) );
  CLKGATETST_X1 pe_1_5_1_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_5_1_N62), .SE(1'b0), .GCK(pe_1_5_1_net4334) );
  CLKGATETST_X1 pe_1_5_1_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_5_1_N61), .SE(1'b0), .GCK(pe_1_5_1_net4339) );
  CLKGATETST_X1 pe_1_5_1_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_5_1_N60), .SE(1'b0), .GCK(pe_1_5_1_net4344) );
  CLKGATETST_X1 pe_1_5_1_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_5_1_N59), .SE(1'b0), .GCK(pe_1_5_1_net4349) );
  CLKGATETST_X1 pe_1_5_1_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_5_1_N90), .SE(1'b0), .GCK(pe_1_5_1_net4354) );
  CLKBUF_X1 pe_1_5_2_U112 ( .A(pe_1_5_2_n72), .Z(pe_1_5_2_n71) );
  INV_X1 pe_1_5_2_U111 ( .A(n76), .ZN(pe_1_5_2_n70) );
  INV_X1 pe_1_5_2_U110 ( .A(n68), .ZN(pe_1_5_2_n69) );
  INV_X1 pe_1_5_2_U109 ( .A(n68), .ZN(pe_1_5_2_n68) );
  INV_X1 pe_1_5_2_U108 ( .A(n68), .ZN(pe_1_5_2_n67) );
  INV_X1 pe_1_5_2_U107 ( .A(pe_1_5_2_n69), .ZN(pe_1_5_2_n66) );
  INV_X1 pe_1_5_2_U106 ( .A(pe_1_5_2_n63), .ZN(pe_1_5_2_n62) );
  INV_X1 pe_1_5_2_U105 ( .A(pe_1_5_2_n61), .ZN(pe_1_5_2_n60) );
  INV_X1 pe_1_5_2_U104 ( .A(n28), .ZN(pe_1_5_2_n59) );
  INV_X1 pe_1_5_2_U103 ( .A(pe_1_5_2_n59), .ZN(pe_1_5_2_n58) );
  INV_X1 pe_1_5_2_U102 ( .A(n20), .ZN(pe_1_5_2_n57) );
  MUX2_X1 pe_1_5_2_U101 ( .A(pe_1_5_2_n54), .B(pe_1_5_2_n51), .S(n51), .Z(
        int_data_x_5__2__3_) );
  MUX2_X1 pe_1_5_2_U100 ( .A(pe_1_5_2_n53), .B(pe_1_5_2_n52), .S(pe_1_5_2_n62), 
        .Z(pe_1_5_2_n54) );
  MUX2_X1 pe_1_5_2_U99 ( .A(pe_1_5_2_int_q_reg_h[23]), .B(
        pe_1_5_2_int_q_reg_h[19]), .S(pe_1_5_2_n56), .Z(pe_1_5_2_n53) );
  MUX2_X1 pe_1_5_2_U98 ( .A(pe_1_5_2_int_q_reg_h[15]), .B(
        pe_1_5_2_int_q_reg_h[11]), .S(pe_1_5_2_n56), .Z(pe_1_5_2_n52) );
  MUX2_X1 pe_1_5_2_U97 ( .A(pe_1_5_2_int_q_reg_h[7]), .B(
        pe_1_5_2_int_q_reg_h[3]), .S(pe_1_5_2_n56), .Z(pe_1_5_2_n51) );
  MUX2_X1 pe_1_5_2_U96 ( .A(pe_1_5_2_n50), .B(pe_1_5_2_n47), .S(n51), .Z(
        int_data_x_5__2__2_) );
  MUX2_X1 pe_1_5_2_U95 ( .A(pe_1_5_2_n49), .B(pe_1_5_2_n48), .S(pe_1_5_2_n62), 
        .Z(pe_1_5_2_n50) );
  MUX2_X1 pe_1_5_2_U94 ( .A(pe_1_5_2_int_q_reg_h[22]), .B(
        pe_1_5_2_int_q_reg_h[18]), .S(pe_1_5_2_n56), .Z(pe_1_5_2_n49) );
  MUX2_X1 pe_1_5_2_U93 ( .A(pe_1_5_2_int_q_reg_h[14]), .B(
        pe_1_5_2_int_q_reg_h[10]), .S(pe_1_5_2_n56), .Z(pe_1_5_2_n48) );
  MUX2_X1 pe_1_5_2_U92 ( .A(pe_1_5_2_int_q_reg_h[6]), .B(
        pe_1_5_2_int_q_reg_h[2]), .S(pe_1_5_2_n56), .Z(pe_1_5_2_n47) );
  MUX2_X1 pe_1_5_2_U91 ( .A(pe_1_5_2_n46), .B(pe_1_5_2_n24), .S(n51), .Z(
        int_data_x_5__2__1_) );
  MUX2_X1 pe_1_5_2_U90 ( .A(pe_1_5_2_n45), .B(pe_1_5_2_n25), .S(pe_1_5_2_n62), 
        .Z(pe_1_5_2_n46) );
  MUX2_X1 pe_1_5_2_U89 ( .A(pe_1_5_2_int_q_reg_h[21]), .B(
        pe_1_5_2_int_q_reg_h[17]), .S(pe_1_5_2_n56), .Z(pe_1_5_2_n45) );
  MUX2_X1 pe_1_5_2_U88 ( .A(pe_1_5_2_int_q_reg_h[13]), .B(
        pe_1_5_2_int_q_reg_h[9]), .S(pe_1_5_2_n56), .Z(pe_1_5_2_n25) );
  MUX2_X1 pe_1_5_2_U87 ( .A(pe_1_5_2_int_q_reg_h[5]), .B(
        pe_1_5_2_int_q_reg_h[1]), .S(pe_1_5_2_n56), .Z(pe_1_5_2_n24) );
  MUX2_X1 pe_1_5_2_U86 ( .A(pe_1_5_2_n23), .B(pe_1_5_2_n20), .S(n51), .Z(
        int_data_x_5__2__0_) );
  MUX2_X1 pe_1_5_2_U85 ( .A(pe_1_5_2_n22), .B(pe_1_5_2_n21), .S(pe_1_5_2_n62), 
        .Z(pe_1_5_2_n23) );
  MUX2_X1 pe_1_5_2_U84 ( .A(pe_1_5_2_int_q_reg_h[20]), .B(
        pe_1_5_2_int_q_reg_h[16]), .S(pe_1_5_2_n56), .Z(pe_1_5_2_n22) );
  MUX2_X1 pe_1_5_2_U83 ( .A(pe_1_5_2_int_q_reg_h[12]), .B(
        pe_1_5_2_int_q_reg_h[8]), .S(pe_1_5_2_n56), .Z(pe_1_5_2_n21) );
  MUX2_X1 pe_1_5_2_U82 ( .A(pe_1_5_2_int_q_reg_h[4]), .B(
        pe_1_5_2_int_q_reg_h[0]), .S(pe_1_5_2_n56), .Z(pe_1_5_2_n20) );
  MUX2_X1 pe_1_5_2_U81 ( .A(pe_1_5_2_n19), .B(pe_1_5_2_n16), .S(n51), .Z(
        int_data_y_5__2__3_) );
  MUX2_X1 pe_1_5_2_U80 ( .A(pe_1_5_2_n18), .B(pe_1_5_2_n17), .S(pe_1_5_2_n62), 
        .Z(pe_1_5_2_n19) );
  MUX2_X1 pe_1_5_2_U79 ( .A(pe_1_5_2_int_q_reg_v[23]), .B(
        pe_1_5_2_int_q_reg_v[19]), .S(pe_1_5_2_n55), .Z(pe_1_5_2_n18) );
  MUX2_X1 pe_1_5_2_U78 ( .A(pe_1_5_2_int_q_reg_v[15]), .B(
        pe_1_5_2_int_q_reg_v[11]), .S(pe_1_5_2_n55), .Z(pe_1_5_2_n17) );
  MUX2_X1 pe_1_5_2_U77 ( .A(pe_1_5_2_int_q_reg_v[7]), .B(
        pe_1_5_2_int_q_reg_v[3]), .S(pe_1_5_2_n55), .Z(pe_1_5_2_n16) );
  MUX2_X1 pe_1_5_2_U76 ( .A(pe_1_5_2_n15), .B(pe_1_5_2_n12), .S(n51), .Z(
        int_data_y_5__2__2_) );
  MUX2_X1 pe_1_5_2_U75 ( .A(pe_1_5_2_n14), .B(pe_1_5_2_n13), .S(pe_1_5_2_n62), 
        .Z(pe_1_5_2_n15) );
  MUX2_X1 pe_1_5_2_U74 ( .A(pe_1_5_2_int_q_reg_v[22]), .B(
        pe_1_5_2_int_q_reg_v[18]), .S(pe_1_5_2_n55), .Z(pe_1_5_2_n14) );
  MUX2_X1 pe_1_5_2_U73 ( .A(pe_1_5_2_int_q_reg_v[14]), .B(
        pe_1_5_2_int_q_reg_v[10]), .S(pe_1_5_2_n55), .Z(pe_1_5_2_n13) );
  MUX2_X1 pe_1_5_2_U72 ( .A(pe_1_5_2_int_q_reg_v[6]), .B(
        pe_1_5_2_int_q_reg_v[2]), .S(pe_1_5_2_n55), .Z(pe_1_5_2_n12) );
  MUX2_X1 pe_1_5_2_U71 ( .A(pe_1_5_2_n11), .B(pe_1_5_2_n8), .S(n51), .Z(
        int_data_y_5__2__1_) );
  MUX2_X1 pe_1_5_2_U70 ( .A(pe_1_5_2_n10), .B(pe_1_5_2_n9), .S(pe_1_5_2_n62), 
        .Z(pe_1_5_2_n11) );
  MUX2_X1 pe_1_5_2_U69 ( .A(pe_1_5_2_int_q_reg_v[21]), .B(
        pe_1_5_2_int_q_reg_v[17]), .S(pe_1_5_2_n55), .Z(pe_1_5_2_n10) );
  MUX2_X1 pe_1_5_2_U68 ( .A(pe_1_5_2_int_q_reg_v[13]), .B(
        pe_1_5_2_int_q_reg_v[9]), .S(pe_1_5_2_n55), .Z(pe_1_5_2_n9) );
  MUX2_X1 pe_1_5_2_U67 ( .A(pe_1_5_2_int_q_reg_v[5]), .B(
        pe_1_5_2_int_q_reg_v[1]), .S(pe_1_5_2_n55), .Z(pe_1_5_2_n8) );
  MUX2_X1 pe_1_5_2_U66 ( .A(pe_1_5_2_n7), .B(pe_1_5_2_n4), .S(n51), .Z(
        int_data_y_5__2__0_) );
  MUX2_X1 pe_1_5_2_U65 ( .A(pe_1_5_2_n6), .B(pe_1_5_2_n5), .S(pe_1_5_2_n62), 
        .Z(pe_1_5_2_n7) );
  MUX2_X1 pe_1_5_2_U64 ( .A(pe_1_5_2_int_q_reg_v[20]), .B(
        pe_1_5_2_int_q_reg_v[16]), .S(pe_1_5_2_n55), .Z(pe_1_5_2_n6) );
  MUX2_X1 pe_1_5_2_U63 ( .A(pe_1_5_2_int_q_reg_v[12]), .B(
        pe_1_5_2_int_q_reg_v[8]), .S(pe_1_5_2_n55), .Z(pe_1_5_2_n5) );
  MUX2_X1 pe_1_5_2_U62 ( .A(pe_1_5_2_int_q_reg_v[4]), .B(
        pe_1_5_2_int_q_reg_v[0]), .S(pe_1_5_2_n55), .Z(pe_1_5_2_n4) );
  AOI222_X1 pe_1_5_2_U61 ( .A1(int_data_res_6__2__2_), .A2(pe_1_5_2_n64), .B1(
        pe_1_5_2_N80), .B2(pe_1_5_2_n27), .C1(pe_1_5_2_N72), .C2(pe_1_5_2_n28), 
        .ZN(pe_1_5_2_n33) );
  INV_X1 pe_1_5_2_U60 ( .A(pe_1_5_2_n33), .ZN(pe_1_5_2_n82) );
  AOI222_X1 pe_1_5_2_U59 ( .A1(int_data_res_6__2__6_), .A2(pe_1_5_2_n64), .B1(
        pe_1_5_2_N84), .B2(pe_1_5_2_n27), .C1(pe_1_5_2_N76), .C2(pe_1_5_2_n28), 
        .ZN(pe_1_5_2_n29) );
  INV_X1 pe_1_5_2_U58 ( .A(pe_1_5_2_n29), .ZN(pe_1_5_2_n78) );
  XNOR2_X1 pe_1_5_2_U57 ( .A(pe_1_5_2_n73), .B(int_data_res_5__2__0_), .ZN(
        pe_1_5_2_N70) );
  AOI222_X1 pe_1_5_2_U52 ( .A1(int_data_res_6__2__0_), .A2(pe_1_5_2_n64), .B1(
        pe_1_5_2_n1), .B2(pe_1_5_2_n27), .C1(pe_1_5_2_N70), .C2(pe_1_5_2_n28), 
        .ZN(pe_1_5_2_n35) );
  INV_X1 pe_1_5_2_U51 ( .A(pe_1_5_2_n35), .ZN(pe_1_5_2_n84) );
  AOI222_X1 pe_1_5_2_U50 ( .A1(int_data_res_6__2__1_), .A2(pe_1_5_2_n64), .B1(
        pe_1_5_2_N79), .B2(pe_1_5_2_n27), .C1(pe_1_5_2_N71), .C2(pe_1_5_2_n28), 
        .ZN(pe_1_5_2_n34) );
  INV_X1 pe_1_5_2_U49 ( .A(pe_1_5_2_n34), .ZN(pe_1_5_2_n83) );
  AOI222_X1 pe_1_5_2_U48 ( .A1(int_data_res_6__2__3_), .A2(pe_1_5_2_n64), .B1(
        pe_1_5_2_N81), .B2(pe_1_5_2_n27), .C1(pe_1_5_2_N73), .C2(pe_1_5_2_n28), 
        .ZN(pe_1_5_2_n32) );
  INV_X1 pe_1_5_2_U47 ( .A(pe_1_5_2_n32), .ZN(pe_1_5_2_n81) );
  AOI222_X1 pe_1_5_2_U46 ( .A1(int_data_res_6__2__4_), .A2(pe_1_5_2_n64), .B1(
        pe_1_5_2_N82), .B2(pe_1_5_2_n27), .C1(pe_1_5_2_N74), .C2(pe_1_5_2_n28), 
        .ZN(pe_1_5_2_n31) );
  INV_X1 pe_1_5_2_U45 ( .A(pe_1_5_2_n31), .ZN(pe_1_5_2_n80) );
  AOI222_X1 pe_1_5_2_U44 ( .A1(int_data_res_6__2__5_), .A2(pe_1_5_2_n64), .B1(
        pe_1_5_2_N83), .B2(pe_1_5_2_n27), .C1(pe_1_5_2_N75), .C2(pe_1_5_2_n28), 
        .ZN(pe_1_5_2_n30) );
  INV_X1 pe_1_5_2_U43 ( .A(pe_1_5_2_n30), .ZN(pe_1_5_2_n79) );
  NAND2_X1 pe_1_5_2_U42 ( .A1(pe_1_5_2_int_data_0_), .A2(pe_1_5_2_n3), .ZN(
        pe_1_5_2_sub_81_carry[1]) );
  INV_X1 pe_1_5_2_U41 ( .A(pe_1_5_2_int_data_1_), .ZN(pe_1_5_2_n74) );
  INV_X1 pe_1_5_2_U40 ( .A(pe_1_5_2_int_data_2_), .ZN(pe_1_5_2_n75) );
  AND2_X1 pe_1_5_2_U39 ( .A1(pe_1_5_2_int_data_0_), .A2(int_data_res_5__2__0_), 
        .ZN(pe_1_5_2_n2) );
  AOI222_X1 pe_1_5_2_U38 ( .A1(pe_1_5_2_n64), .A2(int_data_res_6__2__7_), .B1(
        pe_1_5_2_N85), .B2(pe_1_5_2_n27), .C1(pe_1_5_2_N77), .C2(pe_1_5_2_n28), 
        .ZN(pe_1_5_2_n26) );
  INV_X1 pe_1_5_2_U37 ( .A(pe_1_5_2_n26), .ZN(pe_1_5_2_n77) );
  NOR3_X1 pe_1_5_2_U36 ( .A1(pe_1_5_2_n59), .A2(pe_1_5_2_n65), .A3(int_ckg[21]), .ZN(pe_1_5_2_n36) );
  OR2_X1 pe_1_5_2_U35 ( .A1(pe_1_5_2_n36), .A2(pe_1_5_2_n64), .ZN(pe_1_5_2_N90) );
  INV_X1 pe_1_5_2_U34 ( .A(n40), .ZN(pe_1_5_2_n63) );
  AND2_X1 pe_1_5_2_U33 ( .A1(int_data_x_5__2__2_), .A2(pe_1_5_2_n58), .ZN(
        pe_1_5_2_int_data_2_) );
  AND2_X1 pe_1_5_2_U32 ( .A1(int_data_x_5__2__1_), .A2(pe_1_5_2_n58), .ZN(
        pe_1_5_2_int_data_1_) );
  AND2_X1 pe_1_5_2_U31 ( .A1(int_data_x_5__2__3_), .A2(pe_1_5_2_n58), .ZN(
        pe_1_5_2_int_data_3_) );
  BUF_X1 pe_1_5_2_U30 ( .A(n62), .Z(pe_1_5_2_n64) );
  INV_X1 pe_1_5_2_U29 ( .A(n34), .ZN(pe_1_5_2_n61) );
  AND2_X1 pe_1_5_2_U28 ( .A1(int_data_x_5__2__0_), .A2(pe_1_5_2_n58), .ZN(
        pe_1_5_2_int_data_0_) );
  NAND2_X1 pe_1_5_2_U27 ( .A1(pe_1_5_2_n44), .A2(pe_1_5_2_n61), .ZN(
        pe_1_5_2_n41) );
  AND3_X1 pe_1_5_2_U26 ( .A1(n76), .A2(pe_1_5_2_n63), .A3(n51), .ZN(
        pe_1_5_2_n44) );
  INV_X1 pe_1_5_2_U25 ( .A(pe_1_5_2_int_data_3_), .ZN(pe_1_5_2_n76) );
  NOR2_X1 pe_1_5_2_U24 ( .A1(pe_1_5_2_n70), .A2(n51), .ZN(pe_1_5_2_n43) );
  NOR2_X1 pe_1_5_2_U23 ( .A1(pe_1_5_2_n57), .A2(pe_1_5_2_n64), .ZN(
        pe_1_5_2_n28) );
  NOR2_X1 pe_1_5_2_U22 ( .A1(n20), .A2(pe_1_5_2_n64), .ZN(pe_1_5_2_n27) );
  INV_X1 pe_1_5_2_U21 ( .A(pe_1_5_2_int_data_0_), .ZN(pe_1_5_2_n73) );
  INV_X1 pe_1_5_2_U20 ( .A(pe_1_5_2_n41), .ZN(pe_1_5_2_n90) );
  INV_X1 pe_1_5_2_U19 ( .A(pe_1_5_2_n37), .ZN(pe_1_5_2_n88) );
  INV_X1 pe_1_5_2_U18 ( .A(pe_1_5_2_n38), .ZN(pe_1_5_2_n87) );
  INV_X1 pe_1_5_2_U17 ( .A(pe_1_5_2_n39), .ZN(pe_1_5_2_n86) );
  NOR2_X1 pe_1_5_2_U16 ( .A1(pe_1_5_2_n68), .A2(pe_1_5_2_n42), .ZN(
        pe_1_5_2_N59) );
  NOR2_X1 pe_1_5_2_U15 ( .A1(pe_1_5_2_n68), .A2(pe_1_5_2_n41), .ZN(
        pe_1_5_2_N60) );
  NOR2_X1 pe_1_5_2_U14 ( .A1(pe_1_5_2_n68), .A2(pe_1_5_2_n38), .ZN(
        pe_1_5_2_N63) );
  NOR2_X1 pe_1_5_2_U13 ( .A1(pe_1_5_2_n67), .A2(pe_1_5_2_n40), .ZN(
        pe_1_5_2_N61) );
  NOR2_X1 pe_1_5_2_U12 ( .A1(pe_1_5_2_n67), .A2(pe_1_5_2_n39), .ZN(
        pe_1_5_2_N62) );
  NOR2_X1 pe_1_5_2_U11 ( .A1(pe_1_5_2_n37), .A2(pe_1_5_2_n67), .ZN(
        pe_1_5_2_N64) );
  NAND2_X1 pe_1_5_2_U10 ( .A1(pe_1_5_2_n44), .A2(pe_1_5_2_n60), .ZN(
        pe_1_5_2_n42) );
  BUF_X1 pe_1_5_2_U9 ( .A(pe_1_5_2_n60), .Z(pe_1_5_2_n55) );
  INV_X1 pe_1_5_2_U8 ( .A(pe_1_5_2_n69), .ZN(pe_1_5_2_n65) );
  BUF_X1 pe_1_5_2_U7 ( .A(pe_1_5_2_n60), .Z(pe_1_5_2_n56) );
  INV_X1 pe_1_5_2_U6 ( .A(pe_1_5_2_n42), .ZN(pe_1_5_2_n89) );
  INV_X1 pe_1_5_2_U5 ( .A(pe_1_5_2_n40), .ZN(pe_1_5_2_n85) );
  INV_X2 pe_1_5_2_U4 ( .A(n84), .ZN(pe_1_5_2_n72) );
  XOR2_X1 pe_1_5_2_U3 ( .A(pe_1_5_2_int_data_0_), .B(int_data_res_5__2__0_), 
        .Z(pe_1_5_2_n1) );
  DFFR_X1 pe_1_5_2_int_q_acc_reg_0_ ( .D(pe_1_5_2_n84), .CK(pe_1_5_2_net4276), 
        .RN(pe_1_5_2_n72), .Q(int_data_res_5__2__0_), .QN(pe_1_5_2_n3) );
  DFFR_X1 pe_1_5_2_int_q_reg_v_reg_0__0_ ( .D(int_data_y_6__2__0_), .CK(
        pe_1_5_2_net4246), .RN(pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_v[20]) );
  DFFR_X1 pe_1_5_2_int_q_reg_v_reg_0__1_ ( .D(int_data_y_6__2__1_), .CK(
        pe_1_5_2_net4246), .RN(pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_v[21]) );
  DFFR_X1 pe_1_5_2_int_q_reg_v_reg_0__2_ ( .D(int_data_y_6__2__2_), .CK(
        pe_1_5_2_net4246), .RN(pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_v[22]) );
  DFFR_X1 pe_1_5_2_int_q_reg_v_reg_0__3_ ( .D(int_data_y_6__2__3_), .CK(
        pe_1_5_2_net4246), .RN(pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_v[23]) );
  DFFR_X1 pe_1_5_2_int_q_reg_v_reg_1__0_ ( .D(int_data_y_6__2__0_), .CK(
        pe_1_5_2_net4251), .RN(pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_v[16]) );
  DFFR_X1 pe_1_5_2_int_q_reg_v_reg_1__1_ ( .D(int_data_y_6__2__1_), .CK(
        pe_1_5_2_net4251), .RN(pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_v[17]) );
  DFFR_X1 pe_1_5_2_int_q_reg_v_reg_1__2_ ( .D(int_data_y_6__2__2_), .CK(
        pe_1_5_2_net4251), .RN(pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_v[18]) );
  DFFR_X1 pe_1_5_2_int_q_reg_v_reg_1__3_ ( .D(int_data_y_6__2__3_), .CK(
        pe_1_5_2_net4251), .RN(pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_v[19]) );
  DFFR_X1 pe_1_5_2_int_q_reg_v_reg_2__0_ ( .D(int_data_y_6__2__0_), .CK(
        pe_1_5_2_net4256), .RN(pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_v[12]) );
  DFFR_X1 pe_1_5_2_int_q_reg_v_reg_2__1_ ( .D(int_data_y_6__2__1_), .CK(
        pe_1_5_2_net4256), .RN(pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_v[13]) );
  DFFR_X1 pe_1_5_2_int_q_reg_v_reg_2__2_ ( .D(int_data_y_6__2__2_), .CK(
        pe_1_5_2_net4256), .RN(pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_v[14]) );
  DFFR_X1 pe_1_5_2_int_q_reg_v_reg_2__3_ ( .D(int_data_y_6__2__3_), .CK(
        pe_1_5_2_net4256), .RN(pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_v[15]) );
  DFFR_X1 pe_1_5_2_int_q_reg_v_reg_3__0_ ( .D(int_data_y_6__2__0_), .CK(
        pe_1_5_2_net4261), .RN(pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_v[8]) );
  DFFR_X1 pe_1_5_2_int_q_reg_v_reg_3__1_ ( .D(int_data_y_6__2__1_), .CK(
        pe_1_5_2_net4261), .RN(pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_v[9]) );
  DFFR_X1 pe_1_5_2_int_q_reg_v_reg_3__2_ ( .D(int_data_y_6__2__2_), .CK(
        pe_1_5_2_net4261), .RN(pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_v[10]) );
  DFFR_X1 pe_1_5_2_int_q_reg_v_reg_3__3_ ( .D(int_data_y_6__2__3_), .CK(
        pe_1_5_2_net4261), .RN(pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_v[11]) );
  DFFR_X1 pe_1_5_2_int_q_reg_v_reg_4__0_ ( .D(int_data_y_6__2__0_), .CK(
        pe_1_5_2_net4266), .RN(pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_v[4]) );
  DFFR_X1 pe_1_5_2_int_q_reg_v_reg_4__1_ ( .D(int_data_y_6__2__1_), .CK(
        pe_1_5_2_net4266), .RN(pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_v[5]) );
  DFFR_X1 pe_1_5_2_int_q_reg_v_reg_4__2_ ( .D(int_data_y_6__2__2_), .CK(
        pe_1_5_2_net4266), .RN(pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_v[6]) );
  DFFR_X1 pe_1_5_2_int_q_reg_v_reg_4__3_ ( .D(int_data_y_6__2__3_), .CK(
        pe_1_5_2_net4266), .RN(pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_v[7]) );
  DFFR_X1 pe_1_5_2_int_q_reg_v_reg_5__0_ ( .D(int_data_y_6__2__0_), .CK(
        pe_1_5_2_net4271), .RN(pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_v[0]) );
  DFFR_X1 pe_1_5_2_int_q_reg_v_reg_5__1_ ( .D(int_data_y_6__2__1_), .CK(
        pe_1_5_2_net4271), .RN(pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_v[1]) );
  DFFR_X1 pe_1_5_2_int_q_reg_v_reg_5__2_ ( .D(int_data_y_6__2__2_), .CK(
        pe_1_5_2_net4271), .RN(pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_v[2]) );
  DFFR_X1 pe_1_5_2_int_q_reg_v_reg_5__3_ ( .D(int_data_y_6__2__3_), .CK(
        pe_1_5_2_net4271), .RN(pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_5_2_int_q_reg_h_reg_0__0_ ( .D(int_data_x_5__3__0_), .SI(
        int_data_y_6__2__0_), .SE(pe_1_5_2_n65), .CK(pe_1_5_2_net4215), .RN(
        pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_5_2_int_q_reg_h_reg_0__1_ ( .D(int_data_x_5__3__1_), .SI(
        int_data_y_6__2__1_), .SE(pe_1_5_2_n65), .CK(pe_1_5_2_net4215), .RN(
        pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_5_2_int_q_reg_h_reg_0__2_ ( .D(int_data_x_5__3__2_), .SI(
        int_data_y_6__2__2_), .SE(pe_1_5_2_n65), .CK(pe_1_5_2_net4215), .RN(
        pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_5_2_int_q_reg_h_reg_0__3_ ( .D(int_data_x_5__3__3_), .SI(
        int_data_y_6__2__3_), .SE(pe_1_5_2_n65), .CK(pe_1_5_2_net4215), .RN(
        pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_5_2_int_q_reg_h_reg_1__0_ ( .D(int_data_x_5__3__0_), .SI(
        int_data_y_6__2__0_), .SE(pe_1_5_2_n65), .CK(pe_1_5_2_net4221), .RN(
        pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_5_2_int_q_reg_h_reg_1__1_ ( .D(int_data_x_5__3__1_), .SI(
        int_data_y_6__2__1_), .SE(pe_1_5_2_n65), .CK(pe_1_5_2_net4221), .RN(
        pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_5_2_int_q_reg_h_reg_1__2_ ( .D(int_data_x_5__3__2_), .SI(
        int_data_y_6__2__2_), .SE(pe_1_5_2_n65), .CK(pe_1_5_2_net4221), .RN(
        pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_5_2_int_q_reg_h_reg_1__3_ ( .D(int_data_x_5__3__3_), .SI(
        int_data_y_6__2__3_), .SE(pe_1_5_2_n65), .CK(pe_1_5_2_net4221), .RN(
        pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_5_2_int_q_reg_h_reg_2__0_ ( .D(int_data_x_5__3__0_), .SI(
        int_data_y_6__2__0_), .SE(pe_1_5_2_n65), .CK(pe_1_5_2_net4226), .RN(
        pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_5_2_int_q_reg_h_reg_2__1_ ( .D(int_data_x_5__3__1_), .SI(
        int_data_y_6__2__1_), .SE(pe_1_5_2_n65), .CK(pe_1_5_2_net4226), .RN(
        pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_5_2_int_q_reg_h_reg_2__2_ ( .D(int_data_x_5__3__2_), .SI(
        int_data_y_6__2__2_), .SE(pe_1_5_2_n65), .CK(pe_1_5_2_net4226), .RN(
        pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_5_2_int_q_reg_h_reg_2__3_ ( .D(int_data_x_5__3__3_), .SI(
        int_data_y_6__2__3_), .SE(pe_1_5_2_n65), .CK(pe_1_5_2_net4226), .RN(
        pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_5_2_int_q_reg_h_reg_3__0_ ( .D(int_data_x_5__3__0_), .SI(
        int_data_y_6__2__0_), .SE(pe_1_5_2_n65), .CK(pe_1_5_2_net4231), .RN(
        pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_5_2_int_q_reg_h_reg_3__1_ ( .D(int_data_x_5__3__1_), .SI(
        int_data_y_6__2__1_), .SE(pe_1_5_2_n65), .CK(pe_1_5_2_net4231), .RN(
        pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_5_2_int_q_reg_h_reg_3__2_ ( .D(int_data_x_5__3__2_), .SI(
        int_data_y_6__2__2_), .SE(pe_1_5_2_n65), .CK(pe_1_5_2_net4231), .RN(
        pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_5_2_int_q_reg_h_reg_3__3_ ( .D(int_data_x_5__3__3_), .SI(
        int_data_y_6__2__3_), .SE(pe_1_5_2_n65), .CK(pe_1_5_2_net4231), .RN(
        pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_5_2_int_q_reg_h_reg_4__0_ ( .D(int_data_x_5__3__0_), .SI(
        int_data_y_6__2__0_), .SE(pe_1_5_2_n66), .CK(pe_1_5_2_net4236), .RN(
        pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_5_2_int_q_reg_h_reg_4__1_ ( .D(int_data_x_5__3__1_), .SI(
        int_data_y_6__2__1_), .SE(pe_1_5_2_n66), .CK(pe_1_5_2_net4236), .RN(
        pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_5_2_int_q_reg_h_reg_4__2_ ( .D(int_data_x_5__3__2_), .SI(
        int_data_y_6__2__2_), .SE(pe_1_5_2_n66), .CK(pe_1_5_2_net4236), .RN(
        pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_5_2_int_q_reg_h_reg_4__3_ ( .D(int_data_x_5__3__3_), .SI(
        int_data_y_6__2__3_), .SE(pe_1_5_2_n66), .CK(pe_1_5_2_net4236), .RN(
        pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_5_2_int_q_reg_h_reg_5__0_ ( .D(int_data_x_5__3__0_), .SI(
        int_data_y_6__2__0_), .SE(pe_1_5_2_n66), .CK(pe_1_5_2_net4241), .RN(
        pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_5_2_int_q_reg_h_reg_5__1_ ( .D(int_data_x_5__3__1_), .SI(
        int_data_y_6__2__1_), .SE(pe_1_5_2_n66), .CK(pe_1_5_2_net4241), .RN(
        pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_5_2_int_q_reg_h_reg_5__2_ ( .D(int_data_x_5__3__2_), .SI(
        int_data_y_6__2__2_), .SE(pe_1_5_2_n66), .CK(pe_1_5_2_net4241), .RN(
        pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_5_2_int_q_reg_h_reg_5__3_ ( .D(int_data_x_5__3__3_), .SI(
        int_data_y_6__2__3_), .SE(pe_1_5_2_n66), .CK(pe_1_5_2_net4241), .RN(
        pe_1_5_2_n72), .Q(pe_1_5_2_int_q_reg_h[3]) );
  FA_X1 pe_1_5_2_sub_81_U2_7 ( .A(int_data_res_5__2__7_), .B(pe_1_5_2_n76), 
        .CI(pe_1_5_2_sub_81_carry[7]), .S(pe_1_5_2_N77) );
  FA_X1 pe_1_5_2_sub_81_U2_6 ( .A(int_data_res_5__2__6_), .B(pe_1_5_2_n76), 
        .CI(pe_1_5_2_sub_81_carry[6]), .CO(pe_1_5_2_sub_81_carry[7]), .S(
        pe_1_5_2_N76) );
  FA_X1 pe_1_5_2_sub_81_U2_5 ( .A(int_data_res_5__2__5_), .B(pe_1_5_2_n76), 
        .CI(pe_1_5_2_sub_81_carry[5]), .CO(pe_1_5_2_sub_81_carry[6]), .S(
        pe_1_5_2_N75) );
  FA_X1 pe_1_5_2_sub_81_U2_4 ( .A(int_data_res_5__2__4_), .B(pe_1_5_2_n76), 
        .CI(pe_1_5_2_sub_81_carry[4]), .CO(pe_1_5_2_sub_81_carry[5]), .S(
        pe_1_5_2_N74) );
  FA_X1 pe_1_5_2_sub_81_U2_3 ( .A(int_data_res_5__2__3_), .B(pe_1_5_2_n76), 
        .CI(pe_1_5_2_sub_81_carry[3]), .CO(pe_1_5_2_sub_81_carry[4]), .S(
        pe_1_5_2_N73) );
  FA_X1 pe_1_5_2_sub_81_U2_2 ( .A(int_data_res_5__2__2_), .B(pe_1_5_2_n75), 
        .CI(pe_1_5_2_sub_81_carry[2]), .CO(pe_1_5_2_sub_81_carry[3]), .S(
        pe_1_5_2_N72) );
  FA_X1 pe_1_5_2_sub_81_U2_1 ( .A(int_data_res_5__2__1_), .B(pe_1_5_2_n74), 
        .CI(pe_1_5_2_sub_81_carry[1]), .CO(pe_1_5_2_sub_81_carry[2]), .S(
        pe_1_5_2_N71) );
  FA_X1 pe_1_5_2_add_83_U1_7 ( .A(int_data_res_5__2__7_), .B(
        pe_1_5_2_int_data_3_), .CI(pe_1_5_2_add_83_carry[7]), .S(pe_1_5_2_N85)
         );
  FA_X1 pe_1_5_2_add_83_U1_6 ( .A(int_data_res_5__2__6_), .B(
        pe_1_5_2_int_data_3_), .CI(pe_1_5_2_add_83_carry[6]), .CO(
        pe_1_5_2_add_83_carry[7]), .S(pe_1_5_2_N84) );
  FA_X1 pe_1_5_2_add_83_U1_5 ( .A(int_data_res_5__2__5_), .B(
        pe_1_5_2_int_data_3_), .CI(pe_1_5_2_add_83_carry[5]), .CO(
        pe_1_5_2_add_83_carry[6]), .S(pe_1_5_2_N83) );
  FA_X1 pe_1_5_2_add_83_U1_4 ( .A(int_data_res_5__2__4_), .B(
        pe_1_5_2_int_data_3_), .CI(pe_1_5_2_add_83_carry[4]), .CO(
        pe_1_5_2_add_83_carry[5]), .S(pe_1_5_2_N82) );
  FA_X1 pe_1_5_2_add_83_U1_3 ( .A(int_data_res_5__2__3_), .B(
        pe_1_5_2_int_data_3_), .CI(pe_1_5_2_add_83_carry[3]), .CO(
        pe_1_5_2_add_83_carry[4]), .S(pe_1_5_2_N81) );
  FA_X1 pe_1_5_2_add_83_U1_2 ( .A(int_data_res_5__2__2_), .B(
        pe_1_5_2_int_data_2_), .CI(pe_1_5_2_add_83_carry[2]), .CO(
        pe_1_5_2_add_83_carry[3]), .S(pe_1_5_2_N80) );
  FA_X1 pe_1_5_2_add_83_U1_1 ( .A(int_data_res_5__2__1_), .B(
        pe_1_5_2_int_data_1_), .CI(pe_1_5_2_n2), .CO(pe_1_5_2_add_83_carry[2]), 
        .S(pe_1_5_2_N79) );
  NAND3_X1 pe_1_5_2_U56 ( .A1(pe_1_5_2_n60), .A2(pe_1_5_2_n43), .A3(
        pe_1_5_2_n62), .ZN(pe_1_5_2_n40) );
  NAND3_X1 pe_1_5_2_U55 ( .A1(pe_1_5_2_n43), .A2(pe_1_5_2_n61), .A3(
        pe_1_5_2_n62), .ZN(pe_1_5_2_n39) );
  NAND3_X1 pe_1_5_2_U54 ( .A1(pe_1_5_2_n43), .A2(pe_1_5_2_n63), .A3(
        pe_1_5_2_n60), .ZN(pe_1_5_2_n38) );
  NAND3_X1 pe_1_5_2_U53 ( .A1(pe_1_5_2_n61), .A2(pe_1_5_2_n63), .A3(
        pe_1_5_2_n43), .ZN(pe_1_5_2_n37) );
  DFFR_X1 pe_1_5_2_int_q_acc_reg_6_ ( .D(pe_1_5_2_n78), .CK(pe_1_5_2_net4276), 
        .RN(pe_1_5_2_n71), .Q(int_data_res_5__2__6_) );
  DFFR_X1 pe_1_5_2_int_q_acc_reg_5_ ( .D(pe_1_5_2_n79), .CK(pe_1_5_2_net4276), 
        .RN(pe_1_5_2_n71), .Q(int_data_res_5__2__5_) );
  DFFR_X1 pe_1_5_2_int_q_acc_reg_4_ ( .D(pe_1_5_2_n80), .CK(pe_1_5_2_net4276), 
        .RN(pe_1_5_2_n71), .Q(int_data_res_5__2__4_) );
  DFFR_X1 pe_1_5_2_int_q_acc_reg_3_ ( .D(pe_1_5_2_n81), .CK(pe_1_5_2_net4276), 
        .RN(pe_1_5_2_n71), .Q(int_data_res_5__2__3_) );
  DFFR_X1 pe_1_5_2_int_q_acc_reg_2_ ( .D(pe_1_5_2_n82), .CK(pe_1_5_2_net4276), 
        .RN(pe_1_5_2_n71), .Q(int_data_res_5__2__2_) );
  DFFR_X1 pe_1_5_2_int_q_acc_reg_1_ ( .D(pe_1_5_2_n83), .CK(pe_1_5_2_net4276), 
        .RN(pe_1_5_2_n71), .Q(int_data_res_5__2__1_) );
  DFFR_X1 pe_1_5_2_int_q_acc_reg_7_ ( .D(pe_1_5_2_n77), .CK(pe_1_5_2_net4276), 
        .RN(pe_1_5_2_n71), .Q(int_data_res_5__2__7_) );
  CLKGATETST_X1 pe_1_5_2_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_5_2_n88), .SE(1'b0), .GCK(pe_1_5_2_net4215) );
  CLKGATETST_X1 pe_1_5_2_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_5_2_n87), .SE(1'b0), .GCK(pe_1_5_2_net4221) );
  CLKGATETST_X1 pe_1_5_2_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_5_2_n86), .SE(1'b0), .GCK(pe_1_5_2_net4226) );
  CLKGATETST_X1 pe_1_5_2_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_5_2_n85), .SE(1'b0), .GCK(pe_1_5_2_net4231) );
  CLKGATETST_X1 pe_1_5_2_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_5_2_n90), .SE(1'b0), .GCK(pe_1_5_2_net4236) );
  CLKGATETST_X1 pe_1_5_2_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_5_2_n89), .SE(1'b0), .GCK(pe_1_5_2_net4241) );
  CLKGATETST_X1 pe_1_5_2_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_5_2_N64), .SE(1'b0), .GCK(pe_1_5_2_net4246) );
  CLKGATETST_X1 pe_1_5_2_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_5_2_N63), .SE(1'b0), .GCK(pe_1_5_2_net4251) );
  CLKGATETST_X1 pe_1_5_2_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_5_2_N62), .SE(1'b0), .GCK(pe_1_5_2_net4256) );
  CLKGATETST_X1 pe_1_5_2_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_5_2_N61), .SE(1'b0), .GCK(pe_1_5_2_net4261) );
  CLKGATETST_X1 pe_1_5_2_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_5_2_N60), .SE(1'b0), .GCK(pe_1_5_2_net4266) );
  CLKGATETST_X1 pe_1_5_2_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_5_2_N59), .SE(1'b0), .GCK(pe_1_5_2_net4271) );
  CLKGATETST_X1 pe_1_5_2_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_5_2_N90), .SE(1'b0), .GCK(pe_1_5_2_net4276) );
  CLKBUF_X1 pe_1_5_3_U112 ( .A(pe_1_5_3_n72), .Z(pe_1_5_3_n71) );
  INV_X1 pe_1_5_3_U111 ( .A(n76), .ZN(pe_1_5_3_n70) );
  INV_X1 pe_1_5_3_U110 ( .A(n68), .ZN(pe_1_5_3_n69) );
  INV_X1 pe_1_5_3_U109 ( .A(n68), .ZN(pe_1_5_3_n68) );
  INV_X1 pe_1_5_3_U108 ( .A(n68), .ZN(pe_1_5_3_n67) );
  INV_X1 pe_1_5_3_U107 ( .A(pe_1_5_3_n69), .ZN(pe_1_5_3_n66) );
  INV_X1 pe_1_5_3_U106 ( .A(pe_1_5_3_n63), .ZN(pe_1_5_3_n62) );
  INV_X1 pe_1_5_3_U105 ( .A(pe_1_5_3_n61), .ZN(pe_1_5_3_n60) );
  INV_X1 pe_1_5_3_U104 ( .A(n28), .ZN(pe_1_5_3_n59) );
  INV_X1 pe_1_5_3_U103 ( .A(pe_1_5_3_n59), .ZN(pe_1_5_3_n58) );
  INV_X1 pe_1_5_3_U102 ( .A(n20), .ZN(pe_1_5_3_n57) );
  MUX2_X1 pe_1_5_3_U101 ( .A(pe_1_5_3_n54), .B(pe_1_5_3_n51), .S(n51), .Z(
        int_data_x_5__3__3_) );
  MUX2_X1 pe_1_5_3_U100 ( .A(pe_1_5_3_n53), .B(pe_1_5_3_n52), .S(pe_1_5_3_n62), 
        .Z(pe_1_5_3_n54) );
  MUX2_X1 pe_1_5_3_U99 ( .A(pe_1_5_3_int_q_reg_h[23]), .B(
        pe_1_5_3_int_q_reg_h[19]), .S(pe_1_5_3_n56), .Z(pe_1_5_3_n53) );
  MUX2_X1 pe_1_5_3_U98 ( .A(pe_1_5_3_int_q_reg_h[15]), .B(
        pe_1_5_3_int_q_reg_h[11]), .S(pe_1_5_3_n56), .Z(pe_1_5_3_n52) );
  MUX2_X1 pe_1_5_3_U97 ( .A(pe_1_5_3_int_q_reg_h[7]), .B(
        pe_1_5_3_int_q_reg_h[3]), .S(pe_1_5_3_n56), .Z(pe_1_5_3_n51) );
  MUX2_X1 pe_1_5_3_U96 ( .A(pe_1_5_3_n50), .B(pe_1_5_3_n47), .S(n51), .Z(
        int_data_x_5__3__2_) );
  MUX2_X1 pe_1_5_3_U95 ( .A(pe_1_5_3_n49), .B(pe_1_5_3_n48), .S(pe_1_5_3_n62), 
        .Z(pe_1_5_3_n50) );
  MUX2_X1 pe_1_5_3_U94 ( .A(pe_1_5_3_int_q_reg_h[22]), .B(
        pe_1_5_3_int_q_reg_h[18]), .S(pe_1_5_3_n56), .Z(pe_1_5_3_n49) );
  MUX2_X1 pe_1_5_3_U93 ( .A(pe_1_5_3_int_q_reg_h[14]), .B(
        pe_1_5_3_int_q_reg_h[10]), .S(pe_1_5_3_n56), .Z(pe_1_5_3_n48) );
  MUX2_X1 pe_1_5_3_U92 ( .A(pe_1_5_3_int_q_reg_h[6]), .B(
        pe_1_5_3_int_q_reg_h[2]), .S(pe_1_5_3_n56), .Z(pe_1_5_3_n47) );
  MUX2_X1 pe_1_5_3_U91 ( .A(pe_1_5_3_n46), .B(pe_1_5_3_n24), .S(n51), .Z(
        int_data_x_5__3__1_) );
  MUX2_X1 pe_1_5_3_U90 ( .A(pe_1_5_3_n45), .B(pe_1_5_3_n25), .S(pe_1_5_3_n62), 
        .Z(pe_1_5_3_n46) );
  MUX2_X1 pe_1_5_3_U89 ( .A(pe_1_5_3_int_q_reg_h[21]), .B(
        pe_1_5_3_int_q_reg_h[17]), .S(pe_1_5_3_n56), .Z(pe_1_5_3_n45) );
  MUX2_X1 pe_1_5_3_U88 ( .A(pe_1_5_3_int_q_reg_h[13]), .B(
        pe_1_5_3_int_q_reg_h[9]), .S(pe_1_5_3_n56), .Z(pe_1_5_3_n25) );
  MUX2_X1 pe_1_5_3_U87 ( .A(pe_1_5_3_int_q_reg_h[5]), .B(
        pe_1_5_3_int_q_reg_h[1]), .S(pe_1_5_3_n56), .Z(pe_1_5_3_n24) );
  MUX2_X1 pe_1_5_3_U86 ( .A(pe_1_5_3_n23), .B(pe_1_5_3_n20), .S(n51), .Z(
        int_data_x_5__3__0_) );
  MUX2_X1 pe_1_5_3_U85 ( .A(pe_1_5_3_n22), .B(pe_1_5_3_n21), .S(pe_1_5_3_n62), 
        .Z(pe_1_5_3_n23) );
  MUX2_X1 pe_1_5_3_U84 ( .A(pe_1_5_3_int_q_reg_h[20]), .B(
        pe_1_5_3_int_q_reg_h[16]), .S(pe_1_5_3_n56), .Z(pe_1_5_3_n22) );
  MUX2_X1 pe_1_5_3_U83 ( .A(pe_1_5_3_int_q_reg_h[12]), .B(
        pe_1_5_3_int_q_reg_h[8]), .S(pe_1_5_3_n56), .Z(pe_1_5_3_n21) );
  MUX2_X1 pe_1_5_3_U82 ( .A(pe_1_5_3_int_q_reg_h[4]), .B(
        pe_1_5_3_int_q_reg_h[0]), .S(pe_1_5_3_n56), .Z(pe_1_5_3_n20) );
  MUX2_X1 pe_1_5_3_U81 ( .A(pe_1_5_3_n19), .B(pe_1_5_3_n16), .S(n51), .Z(
        int_data_y_5__3__3_) );
  MUX2_X1 pe_1_5_3_U80 ( .A(pe_1_5_3_n18), .B(pe_1_5_3_n17), .S(pe_1_5_3_n62), 
        .Z(pe_1_5_3_n19) );
  MUX2_X1 pe_1_5_3_U79 ( .A(pe_1_5_3_int_q_reg_v[23]), .B(
        pe_1_5_3_int_q_reg_v[19]), .S(pe_1_5_3_n55), .Z(pe_1_5_3_n18) );
  MUX2_X1 pe_1_5_3_U78 ( .A(pe_1_5_3_int_q_reg_v[15]), .B(
        pe_1_5_3_int_q_reg_v[11]), .S(pe_1_5_3_n55), .Z(pe_1_5_3_n17) );
  MUX2_X1 pe_1_5_3_U77 ( .A(pe_1_5_3_int_q_reg_v[7]), .B(
        pe_1_5_3_int_q_reg_v[3]), .S(pe_1_5_3_n55), .Z(pe_1_5_3_n16) );
  MUX2_X1 pe_1_5_3_U76 ( .A(pe_1_5_3_n15), .B(pe_1_5_3_n12), .S(n51), .Z(
        int_data_y_5__3__2_) );
  MUX2_X1 pe_1_5_3_U75 ( .A(pe_1_5_3_n14), .B(pe_1_5_3_n13), .S(pe_1_5_3_n62), 
        .Z(pe_1_5_3_n15) );
  MUX2_X1 pe_1_5_3_U74 ( .A(pe_1_5_3_int_q_reg_v[22]), .B(
        pe_1_5_3_int_q_reg_v[18]), .S(pe_1_5_3_n55), .Z(pe_1_5_3_n14) );
  MUX2_X1 pe_1_5_3_U73 ( .A(pe_1_5_3_int_q_reg_v[14]), .B(
        pe_1_5_3_int_q_reg_v[10]), .S(pe_1_5_3_n55), .Z(pe_1_5_3_n13) );
  MUX2_X1 pe_1_5_3_U72 ( .A(pe_1_5_3_int_q_reg_v[6]), .B(
        pe_1_5_3_int_q_reg_v[2]), .S(pe_1_5_3_n55), .Z(pe_1_5_3_n12) );
  MUX2_X1 pe_1_5_3_U71 ( .A(pe_1_5_3_n11), .B(pe_1_5_3_n8), .S(n51), .Z(
        int_data_y_5__3__1_) );
  MUX2_X1 pe_1_5_3_U70 ( .A(pe_1_5_3_n10), .B(pe_1_5_3_n9), .S(pe_1_5_3_n62), 
        .Z(pe_1_5_3_n11) );
  MUX2_X1 pe_1_5_3_U69 ( .A(pe_1_5_3_int_q_reg_v[21]), .B(
        pe_1_5_3_int_q_reg_v[17]), .S(pe_1_5_3_n55), .Z(pe_1_5_3_n10) );
  MUX2_X1 pe_1_5_3_U68 ( .A(pe_1_5_3_int_q_reg_v[13]), .B(
        pe_1_5_3_int_q_reg_v[9]), .S(pe_1_5_3_n55), .Z(pe_1_5_3_n9) );
  MUX2_X1 pe_1_5_3_U67 ( .A(pe_1_5_3_int_q_reg_v[5]), .B(
        pe_1_5_3_int_q_reg_v[1]), .S(pe_1_5_3_n55), .Z(pe_1_5_3_n8) );
  MUX2_X1 pe_1_5_3_U66 ( .A(pe_1_5_3_n7), .B(pe_1_5_3_n4), .S(n51), .Z(
        int_data_y_5__3__0_) );
  MUX2_X1 pe_1_5_3_U65 ( .A(pe_1_5_3_n6), .B(pe_1_5_3_n5), .S(pe_1_5_3_n62), 
        .Z(pe_1_5_3_n7) );
  MUX2_X1 pe_1_5_3_U64 ( .A(pe_1_5_3_int_q_reg_v[20]), .B(
        pe_1_5_3_int_q_reg_v[16]), .S(pe_1_5_3_n55), .Z(pe_1_5_3_n6) );
  MUX2_X1 pe_1_5_3_U63 ( .A(pe_1_5_3_int_q_reg_v[12]), .B(
        pe_1_5_3_int_q_reg_v[8]), .S(pe_1_5_3_n55), .Z(pe_1_5_3_n5) );
  MUX2_X1 pe_1_5_3_U62 ( .A(pe_1_5_3_int_q_reg_v[4]), .B(
        pe_1_5_3_int_q_reg_v[0]), .S(pe_1_5_3_n55), .Z(pe_1_5_3_n4) );
  AOI222_X1 pe_1_5_3_U61 ( .A1(int_data_res_6__3__2_), .A2(pe_1_5_3_n64), .B1(
        pe_1_5_3_N80), .B2(pe_1_5_3_n27), .C1(pe_1_5_3_N72), .C2(pe_1_5_3_n28), 
        .ZN(pe_1_5_3_n33) );
  INV_X1 pe_1_5_3_U60 ( .A(pe_1_5_3_n33), .ZN(pe_1_5_3_n82) );
  AOI222_X1 pe_1_5_3_U59 ( .A1(int_data_res_6__3__6_), .A2(pe_1_5_3_n64), .B1(
        pe_1_5_3_N84), .B2(pe_1_5_3_n27), .C1(pe_1_5_3_N76), .C2(pe_1_5_3_n28), 
        .ZN(pe_1_5_3_n29) );
  INV_X1 pe_1_5_3_U58 ( .A(pe_1_5_3_n29), .ZN(pe_1_5_3_n78) );
  XNOR2_X1 pe_1_5_3_U57 ( .A(pe_1_5_3_n73), .B(int_data_res_5__3__0_), .ZN(
        pe_1_5_3_N70) );
  AOI222_X1 pe_1_5_3_U52 ( .A1(int_data_res_6__3__0_), .A2(pe_1_5_3_n64), .B1(
        pe_1_5_3_n1), .B2(pe_1_5_3_n27), .C1(pe_1_5_3_N70), .C2(pe_1_5_3_n28), 
        .ZN(pe_1_5_3_n35) );
  INV_X1 pe_1_5_3_U51 ( .A(pe_1_5_3_n35), .ZN(pe_1_5_3_n84) );
  AOI222_X1 pe_1_5_3_U50 ( .A1(int_data_res_6__3__1_), .A2(pe_1_5_3_n64), .B1(
        pe_1_5_3_N79), .B2(pe_1_5_3_n27), .C1(pe_1_5_3_N71), .C2(pe_1_5_3_n28), 
        .ZN(pe_1_5_3_n34) );
  INV_X1 pe_1_5_3_U49 ( .A(pe_1_5_3_n34), .ZN(pe_1_5_3_n83) );
  AOI222_X1 pe_1_5_3_U48 ( .A1(int_data_res_6__3__3_), .A2(pe_1_5_3_n64), .B1(
        pe_1_5_3_N81), .B2(pe_1_5_3_n27), .C1(pe_1_5_3_N73), .C2(pe_1_5_3_n28), 
        .ZN(pe_1_5_3_n32) );
  INV_X1 pe_1_5_3_U47 ( .A(pe_1_5_3_n32), .ZN(pe_1_5_3_n81) );
  AOI222_X1 pe_1_5_3_U46 ( .A1(int_data_res_6__3__4_), .A2(pe_1_5_3_n64), .B1(
        pe_1_5_3_N82), .B2(pe_1_5_3_n27), .C1(pe_1_5_3_N74), .C2(pe_1_5_3_n28), 
        .ZN(pe_1_5_3_n31) );
  INV_X1 pe_1_5_3_U45 ( .A(pe_1_5_3_n31), .ZN(pe_1_5_3_n80) );
  AOI222_X1 pe_1_5_3_U44 ( .A1(int_data_res_6__3__5_), .A2(pe_1_5_3_n64), .B1(
        pe_1_5_3_N83), .B2(pe_1_5_3_n27), .C1(pe_1_5_3_N75), .C2(pe_1_5_3_n28), 
        .ZN(pe_1_5_3_n30) );
  INV_X1 pe_1_5_3_U43 ( .A(pe_1_5_3_n30), .ZN(pe_1_5_3_n79) );
  NAND2_X1 pe_1_5_3_U42 ( .A1(pe_1_5_3_int_data_0_), .A2(pe_1_5_3_n3), .ZN(
        pe_1_5_3_sub_81_carry[1]) );
  INV_X1 pe_1_5_3_U41 ( .A(pe_1_5_3_int_data_1_), .ZN(pe_1_5_3_n74) );
  INV_X1 pe_1_5_3_U40 ( .A(pe_1_5_3_int_data_2_), .ZN(pe_1_5_3_n75) );
  AND2_X1 pe_1_5_3_U39 ( .A1(pe_1_5_3_int_data_0_), .A2(int_data_res_5__3__0_), 
        .ZN(pe_1_5_3_n2) );
  AOI222_X1 pe_1_5_3_U38 ( .A1(pe_1_5_3_n64), .A2(int_data_res_6__3__7_), .B1(
        pe_1_5_3_N85), .B2(pe_1_5_3_n27), .C1(pe_1_5_3_N77), .C2(pe_1_5_3_n28), 
        .ZN(pe_1_5_3_n26) );
  INV_X1 pe_1_5_3_U37 ( .A(pe_1_5_3_n26), .ZN(pe_1_5_3_n77) );
  NOR3_X1 pe_1_5_3_U36 ( .A1(pe_1_5_3_n59), .A2(pe_1_5_3_n65), .A3(int_ckg[20]), .ZN(pe_1_5_3_n36) );
  OR2_X1 pe_1_5_3_U35 ( .A1(pe_1_5_3_n36), .A2(pe_1_5_3_n64), .ZN(pe_1_5_3_N90) );
  INV_X1 pe_1_5_3_U34 ( .A(n40), .ZN(pe_1_5_3_n63) );
  AND2_X1 pe_1_5_3_U33 ( .A1(int_data_x_5__3__2_), .A2(pe_1_5_3_n58), .ZN(
        pe_1_5_3_int_data_2_) );
  AND2_X1 pe_1_5_3_U32 ( .A1(int_data_x_5__3__1_), .A2(pe_1_5_3_n58), .ZN(
        pe_1_5_3_int_data_1_) );
  AND2_X1 pe_1_5_3_U31 ( .A1(int_data_x_5__3__3_), .A2(pe_1_5_3_n58), .ZN(
        pe_1_5_3_int_data_3_) );
  BUF_X1 pe_1_5_3_U30 ( .A(n62), .Z(pe_1_5_3_n64) );
  INV_X1 pe_1_5_3_U29 ( .A(n34), .ZN(pe_1_5_3_n61) );
  AND2_X1 pe_1_5_3_U28 ( .A1(int_data_x_5__3__0_), .A2(pe_1_5_3_n58), .ZN(
        pe_1_5_3_int_data_0_) );
  NAND2_X1 pe_1_5_3_U27 ( .A1(pe_1_5_3_n44), .A2(pe_1_5_3_n61), .ZN(
        pe_1_5_3_n41) );
  AND3_X1 pe_1_5_3_U26 ( .A1(n76), .A2(pe_1_5_3_n63), .A3(n51), .ZN(
        pe_1_5_3_n44) );
  INV_X1 pe_1_5_3_U25 ( .A(pe_1_5_3_int_data_3_), .ZN(pe_1_5_3_n76) );
  NOR2_X1 pe_1_5_3_U24 ( .A1(pe_1_5_3_n70), .A2(n51), .ZN(pe_1_5_3_n43) );
  NOR2_X1 pe_1_5_3_U23 ( .A1(pe_1_5_3_n57), .A2(pe_1_5_3_n64), .ZN(
        pe_1_5_3_n28) );
  NOR2_X1 pe_1_5_3_U22 ( .A1(n20), .A2(pe_1_5_3_n64), .ZN(pe_1_5_3_n27) );
  INV_X1 pe_1_5_3_U21 ( .A(pe_1_5_3_int_data_0_), .ZN(pe_1_5_3_n73) );
  INV_X1 pe_1_5_3_U20 ( .A(pe_1_5_3_n41), .ZN(pe_1_5_3_n90) );
  INV_X1 pe_1_5_3_U19 ( .A(pe_1_5_3_n37), .ZN(pe_1_5_3_n88) );
  INV_X1 pe_1_5_3_U18 ( .A(pe_1_5_3_n38), .ZN(pe_1_5_3_n87) );
  INV_X1 pe_1_5_3_U17 ( .A(pe_1_5_3_n39), .ZN(pe_1_5_3_n86) );
  NOR2_X1 pe_1_5_3_U16 ( .A1(pe_1_5_3_n68), .A2(pe_1_5_3_n42), .ZN(
        pe_1_5_3_N59) );
  NOR2_X1 pe_1_5_3_U15 ( .A1(pe_1_5_3_n68), .A2(pe_1_5_3_n41), .ZN(
        pe_1_5_3_N60) );
  NOR2_X1 pe_1_5_3_U14 ( .A1(pe_1_5_3_n68), .A2(pe_1_5_3_n38), .ZN(
        pe_1_5_3_N63) );
  NOR2_X1 pe_1_5_3_U13 ( .A1(pe_1_5_3_n67), .A2(pe_1_5_3_n40), .ZN(
        pe_1_5_3_N61) );
  NOR2_X1 pe_1_5_3_U12 ( .A1(pe_1_5_3_n67), .A2(pe_1_5_3_n39), .ZN(
        pe_1_5_3_N62) );
  NOR2_X1 pe_1_5_3_U11 ( .A1(pe_1_5_3_n37), .A2(pe_1_5_3_n67), .ZN(
        pe_1_5_3_N64) );
  NAND2_X1 pe_1_5_3_U10 ( .A1(pe_1_5_3_n44), .A2(pe_1_5_3_n60), .ZN(
        pe_1_5_3_n42) );
  BUF_X1 pe_1_5_3_U9 ( .A(pe_1_5_3_n60), .Z(pe_1_5_3_n55) );
  INV_X1 pe_1_5_3_U8 ( .A(pe_1_5_3_n69), .ZN(pe_1_5_3_n65) );
  BUF_X1 pe_1_5_3_U7 ( .A(pe_1_5_3_n60), .Z(pe_1_5_3_n56) );
  INV_X1 pe_1_5_3_U6 ( .A(pe_1_5_3_n42), .ZN(pe_1_5_3_n89) );
  INV_X1 pe_1_5_3_U5 ( .A(pe_1_5_3_n40), .ZN(pe_1_5_3_n85) );
  INV_X2 pe_1_5_3_U4 ( .A(n84), .ZN(pe_1_5_3_n72) );
  XOR2_X1 pe_1_5_3_U3 ( .A(pe_1_5_3_int_data_0_), .B(int_data_res_5__3__0_), 
        .Z(pe_1_5_3_n1) );
  DFFR_X1 pe_1_5_3_int_q_acc_reg_0_ ( .D(pe_1_5_3_n84), .CK(pe_1_5_3_net4198), 
        .RN(pe_1_5_3_n72), .Q(int_data_res_5__3__0_), .QN(pe_1_5_3_n3) );
  DFFR_X1 pe_1_5_3_int_q_reg_v_reg_0__0_ ( .D(int_data_y_6__3__0_), .CK(
        pe_1_5_3_net4168), .RN(pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_v[20]) );
  DFFR_X1 pe_1_5_3_int_q_reg_v_reg_0__1_ ( .D(int_data_y_6__3__1_), .CK(
        pe_1_5_3_net4168), .RN(pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_v[21]) );
  DFFR_X1 pe_1_5_3_int_q_reg_v_reg_0__2_ ( .D(int_data_y_6__3__2_), .CK(
        pe_1_5_3_net4168), .RN(pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_v[22]) );
  DFFR_X1 pe_1_5_3_int_q_reg_v_reg_0__3_ ( .D(int_data_y_6__3__3_), .CK(
        pe_1_5_3_net4168), .RN(pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_v[23]) );
  DFFR_X1 pe_1_5_3_int_q_reg_v_reg_1__0_ ( .D(int_data_y_6__3__0_), .CK(
        pe_1_5_3_net4173), .RN(pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_v[16]) );
  DFFR_X1 pe_1_5_3_int_q_reg_v_reg_1__1_ ( .D(int_data_y_6__3__1_), .CK(
        pe_1_5_3_net4173), .RN(pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_v[17]) );
  DFFR_X1 pe_1_5_3_int_q_reg_v_reg_1__2_ ( .D(int_data_y_6__3__2_), .CK(
        pe_1_5_3_net4173), .RN(pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_v[18]) );
  DFFR_X1 pe_1_5_3_int_q_reg_v_reg_1__3_ ( .D(int_data_y_6__3__3_), .CK(
        pe_1_5_3_net4173), .RN(pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_v[19]) );
  DFFR_X1 pe_1_5_3_int_q_reg_v_reg_2__0_ ( .D(int_data_y_6__3__0_), .CK(
        pe_1_5_3_net4178), .RN(pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_v[12]) );
  DFFR_X1 pe_1_5_3_int_q_reg_v_reg_2__1_ ( .D(int_data_y_6__3__1_), .CK(
        pe_1_5_3_net4178), .RN(pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_v[13]) );
  DFFR_X1 pe_1_5_3_int_q_reg_v_reg_2__2_ ( .D(int_data_y_6__3__2_), .CK(
        pe_1_5_3_net4178), .RN(pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_v[14]) );
  DFFR_X1 pe_1_5_3_int_q_reg_v_reg_2__3_ ( .D(int_data_y_6__3__3_), .CK(
        pe_1_5_3_net4178), .RN(pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_v[15]) );
  DFFR_X1 pe_1_5_3_int_q_reg_v_reg_3__0_ ( .D(int_data_y_6__3__0_), .CK(
        pe_1_5_3_net4183), .RN(pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_v[8]) );
  DFFR_X1 pe_1_5_3_int_q_reg_v_reg_3__1_ ( .D(int_data_y_6__3__1_), .CK(
        pe_1_5_3_net4183), .RN(pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_v[9]) );
  DFFR_X1 pe_1_5_3_int_q_reg_v_reg_3__2_ ( .D(int_data_y_6__3__2_), .CK(
        pe_1_5_3_net4183), .RN(pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_v[10]) );
  DFFR_X1 pe_1_5_3_int_q_reg_v_reg_3__3_ ( .D(int_data_y_6__3__3_), .CK(
        pe_1_5_3_net4183), .RN(pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_v[11]) );
  DFFR_X1 pe_1_5_3_int_q_reg_v_reg_4__0_ ( .D(int_data_y_6__3__0_), .CK(
        pe_1_5_3_net4188), .RN(pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_v[4]) );
  DFFR_X1 pe_1_5_3_int_q_reg_v_reg_4__1_ ( .D(int_data_y_6__3__1_), .CK(
        pe_1_5_3_net4188), .RN(pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_v[5]) );
  DFFR_X1 pe_1_5_3_int_q_reg_v_reg_4__2_ ( .D(int_data_y_6__3__2_), .CK(
        pe_1_5_3_net4188), .RN(pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_v[6]) );
  DFFR_X1 pe_1_5_3_int_q_reg_v_reg_4__3_ ( .D(int_data_y_6__3__3_), .CK(
        pe_1_5_3_net4188), .RN(pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_v[7]) );
  DFFR_X1 pe_1_5_3_int_q_reg_v_reg_5__0_ ( .D(int_data_y_6__3__0_), .CK(
        pe_1_5_3_net4193), .RN(pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_v[0]) );
  DFFR_X1 pe_1_5_3_int_q_reg_v_reg_5__1_ ( .D(int_data_y_6__3__1_), .CK(
        pe_1_5_3_net4193), .RN(pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_v[1]) );
  DFFR_X1 pe_1_5_3_int_q_reg_v_reg_5__2_ ( .D(int_data_y_6__3__2_), .CK(
        pe_1_5_3_net4193), .RN(pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_v[2]) );
  DFFR_X1 pe_1_5_3_int_q_reg_v_reg_5__3_ ( .D(int_data_y_6__3__3_), .CK(
        pe_1_5_3_net4193), .RN(pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_5_3_int_q_reg_h_reg_0__0_ ( .D(int_data_x_5__4__0_), .SI(
        int_data_y_6__3__0_), .SE(pe_1_5_3_n65), .CK(pe_1_5_3_net4137), .RN(
        pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_5_3_int_q_reg_h_reg_0__1_ ( .D(int_data_x_5__4__1_), .SI(
        int_data_y_6__3__1_), .SE(pe_1_5_3_n65), .CK(pe_1_5_3_net4137), .RN(
        pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_5_3_int_q_reg_h_reg_0__2_ ( .D(int_data_x_5__4__2_), .SI(
        int_data_y_6__3__2_), .SE(pe_1_5_3_n65), .CK(pe_1_5_3_net4137), .RN(
        pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_5_3_int_q_reg_h_reg_0__3_ ( .D(int_data_x_5__4__3_), .SI(
        int_data_y_6__3__3_), .SE(pe_1_5_3_n65), .CK(pe_1_5_3_net4137), .RN(
        pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_5_3_int_q_reg_h_reg_1__0_ ( .D(int_data_x_5__4__0_), .SI(
        int_data_y_6__3__0_), .SE(pe_1_5_3_n65), .CK(pe_1_5_3_net4143), .RN(
        pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_5_3_int_q_reg_h_reg_1__1_ ( .D(int_data_x_5__4__1_), .SI(
        int_data_y_6__3__1_), .SE(pe_1_5_3_n65), .CK(pe_1_5_3_net4143), .RN(
        pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_5_3_int_q_reg_h_reg_1__2_ ( .D(int_data_x_5__4__2_), .SI(
        int_data_y_6__3__2_), .SE(pe_1_5_3_n65), .CK(pe_1_5_3_net4143), .RN(
        pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_5_3_int_q_reg_h_reg_1__3_ ( .D(int_data_x_5__4__3_), .SI(
        int_data_y_6__3__3_), .SE(pe_1_5_3_n65), .CK(pe_1_5_3_net4143), .RN(
        pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_5_3_int_q_reg_h_reg_2__0_ ( .D(int_data_x_5__4__0_), .SI(
        int_data_y_6__3__0_), .SE(pe_1_5_3_n65), .CK(pe_1_5_3_net4148), .RN(
        pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_5_3_int_q_reg_h_reg_2__1_ ( .D(int_data_x_5__4__1_), .SI(
        int_data_y_6__3__1_), .SE(pe_1_5_3_n65), .CK(pe_1_5_3_net4148), .RN(
        pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_5_3_int_q_reg_h_reg_2__2_ ( .D(int_data_x_5__4__2_), .SI(
        int_data_y_6__3__2_), .SE(pe_1_5_3_n65), .CK(pe_1_5_3_net4148), .RN(
        pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_5_3_int_q_reg_h_reg_2__3_ ( .D(int_data_x_5__4__3_), .SI(
        int_data_y_6__3__3_), .SE(pe_1_5_3_n65), .CK(pe_1_5_3_net4148), .RN(
        pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_5_3_int_q_reg_h_reg_3__0_ ( .D(int_data_x_5__4__0_), .SI(
        int_data_y_6__3__0_), .SE(pe_1_5_3_n65), .CK(pe_1_5_3_net4153), .RN(
        pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_5_3_int_q_reg_h_reg_3__1_ ( .D(int_data_x_5__4__1_), .SI(
        int_data_y_6__3__1_), .SE(pe_1_5_3_n65), .CK(pe_1_5_3_net4153), .RN(
        pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_5_3_int_q_reg_h_reg_3__2_ ( .D(int_data_x_5__4__2_), .SI(
        int_data_y_6__3__2_), .SE(pe_1_5_3_n65), .CK(pe_1_5_3_net4153), .RN(
        pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_5_3_int_q_reg_h_reg_3__3_ ( .D(int_data_x_5__4__3_), .SI(
        int_data_y_6__3__3_), .SE(pe_1_5_3_n65), .CK(pe_1_5_3_net4153), .RN(
        pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_5_3_int_q_reg_h_reg_4__0_ ( .D(int_data_x_5__4__0_), .SI(
        int_data_y_6__3__0_), .SE(pe_1_5_3_n66), .CK(pe_1_5_3_net4158), .RN(
        pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_5_3_int_q_reg_h_reg_4__1_ ( .D(int_data_x_5__4__1_), .SI(
        int_data_y_6__3__1_), .SE(pe_1_5_3_n66), .CK(pe_1_5_3_net4158), .RN(
        pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_5_3_int_q_reg_h_reg_4__2_ ( .D(int_data_x_5__4__2_), .SI(
        int_data_y_6__3__2_), .SE(pe_1_5_3_n66), .CK(pe_1_5_3_net4158), .RN(
        pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_5_3_int_q_reg_h_reg_4__3_ ( .D(int_data_x_5__4__3_), .SI(
        int_data_y_6__3__3_), .SE(pe_1_5_3_n66), .CK(pe_1_5_3_net4158), .RN(
        pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_5_3_int_q_reg_h_reg_5__0_ ( .D(int_data_x_5__4__0_), .SI(
        int_data_y_6__3__0_), .SE(pe_1_5_3_n66), .CK(pe_1_5_3_net4163), .RN(
        pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_5_3_int_q_reg_h_reg_5__1_ ( .D(int_data_x_5__4__1_), .SI(
        int_data_y_6__3__1_), .SE(pe_1_5_3_n66), .CK(pe_1_5_3_net4163), .RN(
        pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_5_3_int_q_reg_h_reg_5__2_ ( .D(int_data_x_5__4__2_), .SI(
        int_data_y_6__3__2_), .SE(pe_1_5_3_n66), .CK(pe_1_5_3_net4163), .RN(
        pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_5_3_int_q_reg_h_reg_5__3_ ( .D(int_data_x_5__4__3_), .SI(
        int_data_y_6__3__3_), .SE(pe_1_5_3_n66), .CK(pe_1_5_3_net4163), .RN(
        pe_1_5_3_n72), .Q(pe_1_5_3_int_q_reg_h[3]) );
  FA_X1 pe_1_5_3_sub_81_U2_7 ( .A(int_data_res_5__3__7_), .B(pe_1_5_3_n76), 
        .CI(pe_1_5_3_sub_81_carry[7]), .S(pe_1_5_3_N77) );
  FA_X1 pe_1_5_3_sub_81_U2_6 ( .A(int_data_res_5__3__6_), .B(pe_1_5_3_n76), 
        .CI(pe_1_5_3_sub_81_carry[6]), .CO(pe_1_5_3_sub_81_carry[7]), .S(
        pe_1_5_3_N76) );
  FA_X1 pe_1_5_3_sub_81_U2_5 ( .A(int_data_res_5__3__5_), .B(pe_1_5_3_n76), 
        .CI(pe_1_5_3_sub_81_carry[5]), .CO(pe_1_5_3_sub_81_carry[6]), .S(
        pe_1_5_3_N75) );
  FA_X1 pe_1_5_3_sub_81_U2_4 ( .A(int_data_res_5__3__4_), .B(pe_1_5_3_n76), 
        .CI(pe_1_5_3_sub_81_carry[4]), .CO(pe_1_5_3_sub_81_carry[5]), .S(
        pe_1_5_3_N74) );
  FA_X1 pe_1_5_3_sub_81_U2_3 ( .A(int_data_res_5__3__3_), .B(pe_1_5_3_n76), 
        .CI(pe_1_5_3_sub_81_carry[3]), .CO(pe_1_5_3_sub_81_carry[4]), .S(
        pe_1_5_3_N73) );
  FA_X1 pe_1_5_3_sub_81_U2_2 ( .A(int_data_res_5__3__2_), .B(pe_1_5_3_n75), 
        .CI(pe_1_5_3_sub_81_carry[2]), .CO(pe_1_5_3_sub_81_carry[3]), .S(
        pe_1_5_3_N72) );
  FA_X1 pe_1_5_3_sub_81_U2_1 ( .A(int_data_res_5__3__1_), .B(pe_1_5_3_n74), 
        .CI(pe_1_5_3_sub_81_carry[1]), .CO(pe_1_5_3_sub_81_carry[2]), .S(
        pe_1_5_3_N71) );
  FA_X1 pe_1_5_3_add_83_U1_7 ( .A(int_data_res_5__3__7_), .B(
        pe_1_5_3_int_data_3_), .CI(pe_1_5_3_add_83_carry[7]), .S(pe_1_5_3_N85)
         );
  FA_X1 pe_1_5_3_add_83_U1_6 ( .A(int_data_res_5__3__6_), .B(
        pe_1_5_3_int_data_3_), .CI(pe_1_5_3_add_83_carry[6]), .CO(
        pe_1_5_3_add_83_carry[7]), .S(pe_1_5_3_N84) );
  FA_X1 pe_1_5_3_add_83_U1_5 ( .A(int_data_res_5__3__5_), .B(
        pe_1_5_3_int_data_3_), .CI(pe_1_5_3_add_83_carry[5]), .CO(
        pe_1_5_3_add_83_carry[6]), .S(pe_1_5_3_N83) );
  FA_X1 pe_1_5_3_add_83_U1_4 ( .A(int_data_res_5__3__4_), .B(
        pe_1_5_3_int_data_3_), .CI(pe_1_5_3_add_83_carry[4]), .CO(
        pe_1_5_3_add_83_carry[5]), .S(pe_1_5_3_N82) );
  FA_X1 pe_1_5_3_add_83_U1_3 ( .A(int_data_res_5__3__3_), .B(
        pe_1_5_3_int_data_3_), .CI(pe_1_5_3_add_83_carry[3]), .CO(
        pe_1_5_3_add_83_carry[4]), .S(pe_1_5_3_N81) );
  FA_X1 pe_1_5_3_add_83_U1_2 ( .A(int_data_res_5__3__2_), .B(
        pe_1_5_3_int_data_2_), .CI(pe_1_5_3_add_83_carry[2]), .CO(
        pe_1_5_3_add_83_carry[3]), .S(pe_1_5_3_N80) );
  FA_X1 pe_1_5_3_add_83_U1_1 ( .A(int_data_res_5__3__1_), .B(
        pe_1_5_3_int_data_1_), .CI(pe_1_5_3_n2), .CO(pe_1_5_3_add_83_carry[2]), 
        .S(pe_1_5_3_N79) );
  NAND3_X1 pe_1_5_3_U56 ( .A1(pe_1_5_3_n60), .A2(pe_1_5_3_n43), .A3(
        pe_1_5_3_n62), .ZN(pe_1_5_3_n40) );
  NAND3_X1 pe_1_5_3_U55 ( .A1(pe_1_5_3_n43), .A2(pe_1_5_3_n61), .A3(
        pe_1_5_3_n62), .ZN(pe_1_5_3_n39) );
  NAND3_X1 pe_1_5_3_U54 ( .A1(pe_1_5_3_n43), .A2(pe_1_5_3_n63), .A3(
        pe_1_5_3_n60), .ZN(pe_1_5_3_n38) );
  NAND3_X1 pe_1_5_3_U53 ( .A1(pe_1_5_3_n61), .A2(pe_1_5_3_n63), .A3(
        pe_1_5_3_n43), .ZN(pe_1_5_3_n37) );
  DFFR_X1 pe_1_5_3_int_q_acc_reg_6_ ( .D(pe_1_5_3_n78), .CK(pe_1_5_3_net4198), 
        .RN(pe_1_5_3_n71), .Q(int_data_res_5__3__6_) );
  DFFR_X1 pe_1_5_3_int_q_acc_reg_5_ ( .D(pe_1_5_3_n79), .CK(pe_1_5_3_net4198), 
        .RN(pe_1_5_3_n71), .Q(int_data_res_5__3__5_) );
  DFFR_X1 pe_1_5_3_int_q_acc_reg_4_ ( .D(pe_1_5_3_n80), .CK(pe_1_5_3_net4198), 
        .RN(pe_1_5_3_n71), .Q(int_data_res_5__3__4_) );
  DFFR_X1 pe_1_5_3_int_q_acc_reg_3_ ( .D(pe_1_5_3_n81), .CK(pe_1_5_3_net4198), 
        .RN(pe_1_5_3_n71), .Q(int_data_res_5__3__3_) );
  DFFR_X1 pe_1_5_3_int_q_acc_reg_2_ ( .D(pe_1_5_3_n82), .CK(pe_1_5_3_net4198), 
        .RN(pe_1_5_3_n71), .Q(int_data_res_5__3__2_) );
  DFFR_X1 pe_1_5_3_int_q_acc_reg_1_ ( .D(pe_1_5_3_n83), .CK(pe_1_5_3_net4198), 
        .RN(pe_1_5_3_n71), .Q(int_data_res_5__3__1_) );
  DFFR_X1 pe_1_5_3_int_q_acc_reg_7_ ( .D(pe_1_5_3_n77), .CK(pe_1_5_3_net4198), 
        .RN(pe_1_5_3_n71), .Q(int_data_res_5__3__7_) );
  CLKGATETST_X1 pe_1_5_3_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_5_3_n88), .SE(1'b0), .GCK(pe_1_5_3_net4137) );
  CLKGATETST_X1 pe_1_5_3_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_5_3_n87), .SE(1'b0), .GCK(pe_1_5_3_net4143) );
  CLKGATETST_X1 pe_1_5_3_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_5_3_n86), .SE(1'b0), .GCK(pe_1_5_3_net4148) );
  CLKGATETST_X1 pe_1_5_3_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_5_3_n85), .SE(1'b0), .GCK(pe_1_5_3_net4153) );
  CLKGATETST_X1 pe_1_5_3_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_5_3_n90), .SE(1'b0), .GCK(pe_1_5_3_net4158) );
  CLKGATETST_X1 pe_1_5_3_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_5_3_n89), .SE(1'b0), .GCK(pe_1_5_3_net4163) );
  CLKGATETST_X1 pe_1_5_3_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_5_3_N64), .SE(1'b0), .GCK(pe_1_5_3_net4168) );
  CLKGATETST_X1 pe_1_5_3_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_5_3_N63), .SE(1'b0), .GCK(pe_1_5_3_net4173) );
  CLKGATETST_X1 pe_1_5_3_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_5_3_N62), .SE(1'b0), .GCK(pe_1_5_3_net4178) );
  CLKGATETST_X1 pe_1_5_3_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_5_3_N61), .SE(1'b0), .GCK(pe_1_5_3_net4183) );
  CLKGATETST_X1 pe_1_5_3_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_5_3_N60), .SE(1'b0), .GCK(pe_1_5_3_net4188) );
  CLKGATETST_X1 pe_1_5_3_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_5_3_N59), .SE(1'b0), .GCK(pe_1_5_3_net4193) );
  CLKGATETST_X1 pe_1_5_3_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_5_3_N90), .SE(1'b0), .GCK(pe_1_5_3_net4198) );
  CLKBUF_X1 pe_1_5_4_U112 ( .A(pe_1_5_4_n72), .Z(pe_1_5_4_n71) );
  INV_X1 pe_1_5_4_U111 ( .A(n76), .ZN(pe_1_5_4_n70) );
  INV_X1 pe_1_5_4_U110 ( .A(n68), .ZN(pe_1_5_4_n69) );
  INV_X1 pe_1_5_4_U109 ( .A(n68), .ZN(pe_1_5_4_n68) );
  INV_X1 pe_1_5_4_U108 ( .A(n68), .ZN(pe_1_5_4_n67) );
  INV_X1 pe_1_5_4_U107 ( .A(pe_1_5_4_n69), .ZN(pe_1_5_4_n66) );
  INV_X1 pe_1_5_4_U106 ( .A(pe_1_5_4_n63), .ZN(pe_1_5_4_n62) );
  INV_X1 pe_1_5_4_U105 ( .A(pe_1_5_4_n61), .ZN(pe_1_5_4_n60) );
  INV_X1 pe_1_5_4_U104 ( .A(n28), .ZN(pe_1_5_4_n59) );
  INV_X1 pe_1_5_4_U103 ( .A(pe_1_5_4_n59), .ZN(pe_1_5_4_n58) );
  INV_X1 pe_1_5_4_U102 ( .A(n20), .ZN(pe_1_5_4_n57) );
  MUX2_X1 pe_1_5_4_U101 ( .A(pe_1_5_4_n54), .B(pe_1_5_4_n51), .S(n51), .Z(
        int_data_x_5__4__3_) );
  MUX2_X1 pe_1_5_4_U100 ( .A(pe_1_5_4_n53), .B(pe_1_5_4_n52), .S(pe_1_5_4_n62), 
        .Z(pe_1_5_4_n54) );
  MUX2_X1 pe_1_5_4_U99 ( .A(pe_1_5_4_int_q_reg_h[23]), .B(
        pe_1_5_4_int_q_reg_h[19]), .S(pe_1_5_4_n56), .Z(pe_1_5_4_n53) );
  MUX2_X1 pe_1_5_4_U98 ( .A(pe_1_5_4_int_q_reg_h[15]), .B(
        pe_1_5_4_int_q_reg_h[11]), .S(pe_1_5_4_n56), .Z(pe_1_5_4_n52) );
  MUX2_X1 pe_1_5_4_U97 ( .A(pe_1_5_4_int_q_reg_h[7]), .B(
        pe_1_5_4_int_q_reg_h[3]), .S(pe_1_5_4_n56), .Z(pe_1_5_4_n51) );
  MUX2_X1 pe_1_5_4_U96 ( .A(pe_1_5_4_n50), .B(pe_1_5_4_n47), .S(n51), .Z(
        int_data_x_5__4__2_) );
  MUX2_X1 pe_1_5_4_U95 ( .A(pe_1_5_4_n49), .B(pe_1_5_4_n48), .S(pe_1_5_4_n62), 
        .Z(pe_1_5_4_n50) );
  MUX2_X1 pe_1_5_4_U94 ( .A(pe_1_5_4_int_q_reg_h[22]), .B(
        pe_1_5_4_int_q_reg_h[18]), .S(pe_1_5_4_n56), .Z(pe_1_5_4_n49) );
  MUX2_X1 pe_1_5_4_U93 ( .A(pe_1_5_4_int_q_reg_h[14]), .B(
        pe_1_5_4_int_q_reg_h[10]), .S(pe_1_5_4_n56), .Z(pe_1_5_4_n48) );
  MUX2_X1 pe_1_5_4_U92 ( .A(pe_1_5_4_int_q_reg_h[6]), .B(
        pe_1_5_4_int_q_reg_h[2]), .S(pe_1_5_4_n56), .Z(pe_1_5_4_n47) );
  MUX2_X1 pe_1_5_4_U91 ( .A(pe_1_5_4_n46), .B(pe_1_5_4_n24), .S(n51), .Z(
        int_data_x_5__4__1_) );
  MUX2_X1 pe_1_5_4_U90 ( .A(pe_1_5_4_n45), .B(pe_1_5_4_n25), .S(pe_1_5_4_n62), 
        .Z(pe_1_5_4_n46) );
  MUX2_X1 pe_1_5_4_U89 ( .A(pe_1_5_4_int_q_reg_h[21]), .B(
        pe_1_5_4_int_q_reg_h[17]), .S(pe_1_5_4_n56), .Z(pe_1_5_4_n45) );
  MUX2_X1 pe_1_5_4_U88 ( .A(pe_1_5_4_int_q_reg_h[13]), .B(
        pe_1_5_4_int_q_reg_h[9]), .S(pe_1_5_4_n56), .Z(pe_1_5_4_n25) );
  MUX2_X1 pe_1_5_4_U87 ( .A(pe_1_5_4_int_q_reg_h[5]), .B(
        pe_1_5_4_int_q_reg_h[1]), .S(pe_1_5_4_n56), .Z(pe_1_5_4_n24) );
  MUX2_X1 pe_1_5_4_U86 ( .A(pe_1_5_4_n23), .B(pe_1_5_4_n20), .S(n51), .Z(
        int_data_x_5__4__0_) );
  MUX2_X1 pe_1_5_4_U85 ( .A(pe_1_5_4_n22), .B(pe_1_5_4_n21), .S(pe_1_5_4_n62), 
        .Z(pe_1_5_4_n23) );
  MUX2_X1 pe_1_5_4_U84 ( .A(pe_1_5_4_int_q_reg_h[20]), .B(
        pe_1_5_4_int_q_reg_h[16]), .S(pe_1_5_4_n56), .Z(pe_1_5_4_n22) );
  MUX2_X1 pe_1_5_4_U83 ( .A(pe_1_5_4_int_q_reg_h[12]), .B(
        pe_1_5_4_int_q_reg_h[8]), .S(pe_1_5_4_n56), .Z(pe_1_5_4_n21) );
  MUX2_X1 pe_1_5_4_U82 ( .A(pe_1_5_4_int_q_reg_h[4]), .B(
        pe_1_5_4_int_q_reg_h[0]), .S(pe_1_5_4_n56), .Z(pe_1_5_4_n20) );
  MUX2_X1 pe_1_5_4_U81 ( .A(pe_1_5_4_n19), .B(pe_1_5_4_n16), .S(n51), .Z(
        int_data_y_5__4__3_) );
  MUX2_X1 pe_1_5_4_U80 ( .A(pe_1_5_4_n18), .B(pe_1_5_4_n17), .S(pe_1_5_4_n62), 
        .Z(pe_1_5_4_n19) );
  MUX2_X1 pe_1_5_4_U79 ( .A(pe_1_5_4_int_q_reg_v[23]), .B(
        pe_1_5_4_int_q_reg_v[19]), .S(pe_1_5_4_n55), .Z(pe_1_5_4_n18) );
  MUX2_X1 pe_1_5_4_U78 ( .A(pe_1_5_4_int_q_reg_v[15]), .B(
        pe_1_5_4_int_q_reg_v[11]), .S(pe_1_5_4_n55), .Z(pe_1_5_4_n17) );
  MUX2_X1 pe_1_5_4_U77 ( .A(pe_1_5_4_int_q_reg_v[7]), .B(
        pe_1_5_4_int_q_reg_v[3]), .S(pe_1_5_4_n55), .Z(pe_1_5_4_n16) );
  MUX2_X1 pe_1_5_4_U76 ( .A(pe_1_5_4_n15), .B(pe_1_5_4_n12), .S(n51), .Z(
        int_data_y_5__4__2_) );
  MUX2_X1 pe_1_5_4_U75 ( .A(pe_1_5_4_n14), .B(pe_1_5_4_n13), .S(pe_1_5_4_n62), 
        .Z(pe_1_5_4_n15) );
  MUX2_X1 pe_1_5_4_U74 ( .A(pe_1_5_4_int_q_reg_v[22]), .B(
        pe_1_5_4_int_q_reg_v[18]), .S(pe_1_5_4_n55), .Z(pe_1_5_4_n14) );
  MUX2_X1 pe_1_5_4_U73 ( .A(pe_1_5_4_int_q_reg_v[14]), .B(
        pe_1_5_4_int_q_reg_v[10]), .S(pe_1_5_4_n55), .Z(pe_1_5_4_n13) );
  MUX2_X1 pe_1_5_4_U72 ( .A(pe_1_5_4_int_q_reg_v[6]), .B(
        pe_1_5_4_int_q_reg_v[2]), .S(pe_1_5_4_n55), .Z(pe_1_5_4_n12) );
  MUX2_X1 pe_1_5_4_U71 ( .A(pe_1_5_4_n11), .B(pe_1_5_4_n8), .S(n51), .Z(
        int_data_y_5__4__1_) );
  MUX2_X1 pe_1_5_4_U70 ( .A(pe_1_5_4_n10), .B(pe_1_5_4_n9), .S(pe_1_5_4_n62), 
        .Z(pe_1_5_4_n11) );
  MUX2_X1 pe_1_5_4_U69 ( .A(pe_1_5_4_int_q_reg_v[21]), .B(
        pe_1_5_4_int_q_reg_v[17]), .S(pe_1_5_4_n55), .Z(pe_1_5_4_n10) );
  MUX2_X1 pe_1_5_4_U68 ( .A(pe_1_5_4_int_q_reg_v[13]), .B(
        pe_1_5_4_int_q_reg_v[9]), .S(pe_1_5_4_n55), .Z(pe_1_5_4_n9) );
  MUX2_X1 pe_1_5_4_U67 ( .A(pe_1_5_4_int_q_reg_v[5]), .B(
        pe_1_5_4_int_q_reg_v[1]), .S(pe_1_5_4_n55), .Z(pe_1_5_4_n8) );
  MUX2_X1 pe_1_5_4_U66 ( .A(pe_1_5_4_n7), .B(pe_1_5_4_n4), .S(n51), .Z(
        int_data_y_5__4__0_) );
  MUX2_X1 pe_1_5_4_U65 ( .A(pe_1_5_4_n6), .B(pe_1_5_4_n5), .S(pe_1_5_4_n62), 
        .Z(pe_1_5_4_n7) );
  MUX2_X1 pe_1_5_4_U64 ( .A(pe_1_5_4_int_q_reg_v[20]), .B(
        pe_1_5_4_int_q_reg_v[16]), .S(pe_1_5_4_n55), .Z(pe_1_5_4_n6) );
  MUX2_X1 pe_1_5_4_U63 ( .A(pe_1_5_4_int_q_reg_v[12]), .B(
        pe_1_5_4_int_q_reg_v[8]), .S(pe_1_5_4_n55), .Z(pe_1_5_4_n5) );
  MUX2_X1 pe_1_5_4_U62 ( .A(pe_1_5_4_int_q_reg_v[4]), .B(
        pe_1_5_4_int_q_reg_v[0]), .S(pe_1_5_4_n55), .Z(pe_1_5_4_n4) );
  AOI222_X1 pe_1_5_4_U61 ( .A1(int_data_res_6__4__2_), .A2(pe_1_5_4_n64), .B1(
        pe_1_5_4_N80), .B2(pe_1_5_4_n27), .C1(pe_1_5_4_N72), .C2(pe_1_5_4_n28), 
        .ZN(pe_1_5_4_n33) );
  INV_X1 pe_1_5_4_U60 ( .A(pe_1_5_4_n33), .ZN(pe_1_5_4_n82) );
  AOI222_X1 pe_1_5_4_U59 ( .A1(int_data_res_6__4__6_), .A2(pe_1_5_4_n64), .B1(
        pe_1_5_4_N84), .B2(pe_1_5_4_n27), .C1(pe_1_5_4_N76), .C2(pe_1_5_4_n28), 
        .ZN(pe_1_5_4_n29) );
  INV_X1 pe_1_5_4_U58 ( .A(pe_1_5_4_n29), .ZN(pe_1_5_4_n78) );
  XNOR2_X1 pe_1_5_4_U57 ( .A(pe_1_5_4_n73), .B(int_data_res_5__4__0_), .ZN(
        pe_1_5_4_N70) );
  AOI222_X1 pe_1_5_4_U52 ( .A1(int_data_res_6__4__0_), .A2(pe_1_5_4_n64), .B1(
        pe_1_5_4_n1), .B2(pe_1_5_4_n27), .C1(pe_1_5_4_N70), .C2(pe_1_5_4_n28), 
        .ZN(pe_1_5_4_n35) );
  INV_X1 pe_1_5_4_U51 ( .A(pe_1_5_4_n35), .ZN(pe_1_5_4_n84) );
  AOI222_X1 pe_1_5_4_U50 ( .A1(int_data_res_6__4__1_), .A2(pe_1_5_4_n64), .B1(
        pe_1_5_4_N79), .B2(pe_1_5_4_n27), .C1(pe_1_5_4_N71), .C2(pe_1_5_4_n28), 
        .ZN(pe_1_5_4_n34) );
  INV_X1 pe_1_5_4_U49 ( .A(pe_1_5_4_n34), .ZN(pe_1_5_4_n83) );
  AOI222_X1 pe_1_5_4_U48 ( .A1(int_data_res_6__4__3_), .A2(pe_1_5_4_n64), .B1(
        pe_1_5_4_N81), .B2(pe_1_5_4_n27), .C1(pe_1_5_4_N73), .C2(pe_1_5_4_n28), 
        .ZN(pe_1_5_4_n32) );
  INV_X1 pe_1_5_4_U47 ( .A(pe_1_5_4_n32), .ZN(pe_1_5_4_n81) );
  AOI222_X1 pe_1_5_4_U46 ( .A1(int_data_res_6__4__4_), .A2(pe_1_5_4_n64), .B1(
        pe_1_5_4_N82), .B2(pe_1_5_4_n27), .C1(pe_1_5_4_N74), .C2(pe_1_5_4_n28), 
        .ZN(pe_1_5_4_n31) );
  INV_X1 pe_1_5_4_U45 ( .A(pe_1_5_4_n31), .ZN(pe_1_5_4_n80) );
  AOI222_X1 pe_1_5_4_U44 ( .A1(int_data_res_6__4__5_), .A2(pe_1_5_4_n64), .B1(
        pe_1_5_4_N83), .B2(pe_1_5_4_n27), .C1(pe_1_5_4_N75), .C2(pe_1_5_4_n28), 
        .ZN(pe_1_5_4_n30) );
  INV_X1 pe_1_5_4_U43 ( .A(pe_1_5_4_n30), .ZN(pe_1_5_4_n79) );
  NAND2_X1 pe_1_5_4_U42 ( .A1(pe_1_5_4_int_data_0_), .A2(pe_1_5_4_n3), .ZN(
        pe_1_5_4_sub_81_carry[1]) );
  INV_X1 pe_1_5_4_U41 ( .A(pe_1_5_4_int_data_1_), .ZN(pe_1_5_4_n74) );
  INV_X1 pe_1_5_4_U40 ( .A(pe_1_5_4_int_data_2_), .ZN(pe_1_5_4_n75) );
  AND2_X1 pe_1_5_4_U39 ( .A1(pe_1_5_4_int_data_0_), .A2(int_data_res_5__4__0_), 
        .ZN(pe_1_5_4_n2) );
  AOI222_X1 pe_1_5_4_U38 ( .A1(pe_1_5_4_n64), .A2(int_data_res_6__4__7_), .B1(
        pe_1_5_4_N85), .B2(pe_1_5_4_n27), .C1(pe_1_5_4_N77), .C2(pe_1_5_4_n28), 
        .ZN(pe_1_5_4_n26) );
  INV_X1 pe_1_5_4_U37 ( .A(pe_1_5_4_n26), .ZN(pe_1_5_4_n77) );
  NOR3_X1 pe_1_5_4_U36 ( .A1(pe_1_5_4_n59), .A2(pe_1_5_4_n65), .A3(int_ckg[19]), .ZN(pe_1_5_4_n36) );
  OR2_X1 pe_1_5_4_U35 ( .A1(pe_1_5_4_n36), .A2(pe_1_5_4_n64), .ZN(pe_1_5_4_N90) );
  INV_X1 pe_1_5_4_U34 ( .A(n40), .ZN(pe_1_5_4_n63) );
  AND2_X1 pe_1_5_4_U33 ( .A1(int_data_x_5__4__2_), .A2(pe_1_5_4_n58), .ZN(
        pe_1_5_4_int_data_2_) );
  AND2_X1 pe_1_5_4_U32 ( .A1(int_data_x_5__4__1_), .A2(pe_1_5_4_n58), .ZN(
        pe_1_5_4_int_data_1_) );
  AND2_X1 pe_1_5_4_U31 ( .A1(int_data_x_5__4__3_), .A2(pe_1_5_4_n58), .ZN(
        pe_1_5_4_int_data_3_) );
  BUF_X1 pe_1_5_4_U30 ( .A(n62), .Z(pe_1_5_4_n64) );
  INV_X1 pe_1_5_4_U29 ( .A(n34), .ZN(pe_1_5_4_n61) );
  AND2_X1 pe_1_5_4_U28 ( .A1(int_data_x_5__4__0_), .A2(pe_1_5_4_n58), .ZN(
        pe_1_5_4_int_data_0_) );
  NAND2_X1 pe_1_5_4_U27 ( .A1(pe_1_5_4_n44), .A2(pe_1_5_4_n61), .ZN(
        pe_1_5_4_n41) );
  AND3_X1 pe_1_5_4_U26 ( .A1(n76), .A2(pe_1_5_4_n63), .A3(n51), .ZN(
        pe_1_5_4_n44) );
  INV_X1 pe_1_5_4_U25 ( .A(pe_1_5_4_int_data_3_), .ZN(pe_1_5_4_n76) );
  NOR2_X1 pe_1_5_4_U24 ( .A1(pe_1_5_4_n70), .A2(n51), .ZN(pe_1_5_4_n43) );
  NOR2_X1 pe_1_5_4_U23 ( .A1(pe_1_5_4_n57), .A2(pe_1_5_4_n64), .ZN(
        pe_1_5_4_n28) );
  NOR2_X1 pe_1_5_4_U22 ( .A1(n20), .A2(pe_1_5_4_n64), .ZN(pe_1_5_4_n27) );
  INV_X1 pe_1_5_4_U21 ( .A(pe_1_5_4_int_data_0_), .ZN(pe_1_5_4_n73) );
  INV_X1 pe_1_5_4_U20 ( .A(pe_1_5_4_n41), .ZN(pe_1_5_4_n90) );
  INV_X1 pe_1_5_4_U19 ( .A(pe_1_5_4_n37), .ZN(pe_1_5_4_n88) );
  INV_X1 pe_1_5_4_U18 ( .A(pe_1_5_4_n38), .ZN(pe_1_5_4_n87) );
  INV_X1 pe_1_5_4_U17 ( .A(pe_1_5_4_n39), .ZN(pe_1_5_4_n86) );
  NOR2_X1 pe_1_5_4_U16 ( .A1(pe_1_5_4_n68), .A2(pe_1_5_4_n42), .ZN(
        pe_1_5_4_N59) );
  NOR2_X1 pe_1_5_4_U15 ( .A1(pe_1_5_4_n68), .A2(pe_1_5_4_n41), .ZN(
        pe_1_5_4_N60) );
  NOR2_X1 pe_1_5_4_U14 ( .A1(pe_1_5_4_n68), .A2(pe_1_5_4_n38), .ZN(
        pe_1_5_4_N63) );
  NOR2_X1 pe_1_5_4_U13 ( .A1(pe_1_5_4_n67), .A2(pe_1_5_4_n40), .ZN(
        pe_1_5_4_N61) );
  NOR2_X1 pe_1_5_4_U12 ( .A1(pe_1_5_4_n67), .A2(pe_1_5_4_n39), .ZN(
        pe_1_5_4_N62) );
  NOR2_X1 pe_1_5_4_U11 ( .A1(pe_1_5_4_n37), .A2(pe_1_5_4_n67), .ZN(
        pe_1_5_4_N64) );
  NAND2_X1 pe_1_5_4_U10 ( .A1(pe_1_5_4_n44), .A2(pe_1_5_4_n60), .ZN(
        pe_1_5_4_n42) );
  BUF_X1 pe_1_5_4_U9 ( .A(pe_1_5_4_n60), .Z(pe_1_5_4_n55) );
  INV_X1 pe_1_5_4_U8 ( .A(pe_1_5_4_n69), .ZN(pe_1_5_4_n65) );
  BUF_X1 pe_1_5_4_U7 ( .A(pe_1_5_4_n60), .Z(pe_1_5_4_n56) );
  INV_X1 pe_1_5_4_U6 ( .A(pe_1_5_4_n42), .ZN(pe_1_5_4_n89) );
  INV_X1 pe_1_5_4_U5 ( .A(pe_1_5_4_n40), .ZN(pe_1_5_4_n85) );
  INV_X2 pe_1_5_4_U4 ( .A(n84), .ZN(pe_1_5_4_n72) );
  XOR2_X1 pe_1_5_4_U3 ( .A(pe_1_5_4_int_data_0_), .B(int_data_res_5__4__0_), 
        .Z(pe_1_5_4_n1) );
  DFFR_X1 pe_1_5_4_int_q_acc_reg_0_ ( .D(pe_1_5_4_n84), .CK(pe_1_5_4_net4120), 
        .RN(pe_1_5_4_n72), .Q(int_data_res_5__4__0_), .QN(pe_1_5_4_n3) );
  DFFR_X1 pe_1_5_4_int_q_reg_v_reg_0__0_ ( .D(int_data_y_6__4__0_), .CK(
        pe_1_5_4_net4090), .RN(pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_v[20]) );
  DFFR_X1 pe_1_5_4_int_q_reg_v_reg_0__1_ ( .D(int_data_y_6__4__1_), .CK(
        pe_1_5_4_net4090), .RN(pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_v[21]) );
  DFFR_X1 pe_1_5_4_int_q_reg_v_reg_0__2_ ( .D(int_data_y_6__4__2_), .CK(
        pe_1_5_4_net4090), .RN(pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_v[22]) );
  DFFR_X1 pe_1_5_4_int_q_reg_v_reg_0__3_ ( .D(int_data_y_6__4__3_), .CK(
        pe_1_5_4_net4090), .RN(pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_v[23]) );
  DFFR_X1 pe_1_5_4_int_q_reg_v_reg_1__0_ ( .D(int_data_y_6__4__0_), .CK(
        pe_1_5_4_net4095), .RN(pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_v[16]) );
  DFFR_X1 pe_1_5_4_int_q_reg_v_reg_1__1_ ( .D(int_data_y_6__4__1_), .CK(
        pe_1_5_4_net4095), .RN(pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_v[17]) );
  DFFR_X1 pe_1_5_4_int_q_reg_v_reg_1__2_ ( .D(int_data_y_6__4__2_), .CK(
        pe_1_5_4_net4095), .RN(pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_v[18]) );
  DFFR_X1 pe_1_5_4_int_q_reg_v_reg_1__3_ ( .D(int_data_y_6__4__3_), .CK(
        pe_1_5_4_net4095), .RN(pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_v[19]) );
  DFFR_X1 pe_1_5_4_int_q_reg_v_reg_2__0_ ( .D(int_data_y_6__4__0_), .CK(
        pe_1_5_4_net4100), .RN(pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_v[12]) );
  DFFR_X1 pe_1_5_4_int_q_reg_v_reg_2__1_ ( .D(int_data_y_6__4__1_), .CK(
        pe_1_5_4_net4100), .RN(pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_v[13]) );
  DFFR_X1 pe_1_5_4_int_q_reg_v_reg_2__2_ ( .D(int_data_y_6__4__2_), .CK(
        pe_1_5_4_net4100), .RN(pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_v[14]) );
  DFFR_X1 pe_1_5_4_int_q_reg_v_reg_2__3_ ( .D(int_data_y_6__4__3_), .CK(
        pe_1_5_4_net4100), .RN(pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_v[15]) );
  DFFR_X1 pe_1_5_4_int_q_reg_v_reg_3__0_ ( .D(int_data_y_6__4__0_), .CK(
        pe_1_5_4_net4105), .RN(pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_v[8]) );
  DFFR_X1 pe_1_5_4_int_q_reg_v_reg_3__1_ ( .D(int_data_y_6__4__1_), .CK(
        pe_1_5_4_net4105), .RN(pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_v[9]) );
  DFFR_X1 pe_1_5_4_int_q_reg_v_reg_3__2_ ( .D(int_data_y_6__4__2_), .CK(
        pe_1_5_4_net4105), .RN(pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_v[10]) );
  DFFR_X1 pe_1_5_4_int_q_reg_v_reg_3__3_ ( .D(int_data_y_6__4__3_), .CK(
        pe_1_5_4_net4105), .RN(pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_v[11]) );
  DFFR_X1 pe_1_5_4_int_q_reg_v_reg_4__0_ ( .D(int_data_y_6__4__0_), .CK(
        pe_1_5_4_net4110), .RN(pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_v[4]) );
  DFFR_X1 pe_1_5_4_int_q_reg_v_reg_4__1_ ( .D(int_data_y_6__4__1_), .CK(
        pe_1_5_4_net4110), .RN(pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_v[5]) );
  DFFR_X1 pe_1_5_4_int_q_reg_v_reg_4__2_ ( .D(int_data_y_6__4__2_), .CK(
        pe_1_5_4_net4110), .RN(pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_v[6]) );
  DFFR_X1 pe_1_5_4_int_q_reg_v_reg_4__3_ ( .D(int_data_y_6__4__3_), .CK(
        pe_1_5_4_net4110), .RN(pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_v[7]) );
  DFFR_X1 pe_1_5_4_int_q_reg_v_reg_5__0_ ( .D(int_data_y_6__4__0_), .CK(
        pe_1_5_4_net4115), .RN(pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_v[0]) );
  DFFR_X1 pe_1_5_4_int_q_reg_v_reg_5__1_ ( .D(int_data_y_6__4__1_), .CK(
        pe_1_5_4_net4115), .RN(pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_v[1]) );
  DFFR_X1 pe_1_5_4_int_q_reg_v_reg_5__2_ ( .D(int_data_y_6__4__2_), .CK(
        pe_1_5_4_net4115), .RN(pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_v[2]) );
  DFFR_X1 pe_1_5_4_int_q_reg_v_reg_5__3_ ( .D(int_data_y_6__4__3_), .CK(
        pe_1_5_4_net4115), .RN(pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_5_4_int_q_reg_h_reg_0__0_ ( .D(int_data_x_5__5__0_), .SI(
        int_data_y_6__4__0_), .SE(pe_1_5_4_n65), .CK(pe_1_5_4_net4059), .RN(
        pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_5_4_int_q_reg_h_reg_0__1_ ( .D(int_data_x_5__5__1_), .SI(
        int_data_y_6__4__1_), .SE(pe_1_5_4_n65), .CK(pe_1_5_4_net4059), .RN(
        pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_5_4_int_q_reg_h_reg_0__2_ ( .D(int_data_x_5__5__2_), .SI(
        int_data_y_6__4__2_), .SE(pe_1_5_4_n65), .CK(pe_1_5_4_net4059), .RN(
        pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_5_4_int_q_reg_h_reg_0__3_ ( .D(int_data_x_5__5__3_), .SI(
        int_data_y_6__4__3_), .SE(pe_1_5_4_n65), .CK(pe_1_5_4_net4059), .RN(
        pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_5_4_int_q_reg_h_reg_1__0_ ( .D(int_data_x_5__5__0_), .SI(
        int_data_y_6__4__0_), .SE(pe_1_5_4_n65), .CK(pe_1_5_4_net4065), .RN(
        pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_5_4_int_q_reg_h_reg_1__1_ ( .D(int_data_x_5__5__1_), .SI(
        int_data_y_6__4__1_), .SE(pe_1_5_4_n65), .CK(pe_1_5_4_net4065), .RN(
        pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_5_4_int_q_reg_h_reg_1__2_ ( .D(int_data_x_5__5__2_), .SI(
        int_data_y_6__4__2_), .SE(pe_1_5_4_n65), .CK(pe_1_5_4_net4065), .RN(
        pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_5_4_int_q_reg_h_reg_1__3_ ( .D(int_data_x_5__5__3_), .SI(
        int_data_y_6__4__3_), .SE(pe_1_5_4_n65), .CK(pe_1_5_4_net4065), .RN(
        pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_5_4_int_q_reg_h_reg_2__0_ ( .D(int_data_x_5__5__0_), .SI(
        int_data_y_6__4__0_), .SE(pe_1_5_4_n65), .CK(pe_1_5_4_net4070), .RN(
        pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_5_4_int_q_reg_h_reg_2__1_ ( .D(int_data_x_5__5__1_), .SI(
        int_data_y_6__4__1_), .SE(pe_1_5_4_n65), .CK(pe_1_5_4_net4070), .RN(
        pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_5_4_int_q_reg_h_reg_2__2_ ( .D(int_data_x_5__5__2_), .SI(
        int_data_y_6__4__2_), .SE(pe_1_5_4_n65), .CK(pe_1_5_4_net4070), .RN(
        pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_5_4_int_q_reg_h_reg_2__3_ ( .D(int_data_x_5__5__3_), .SI(
        int_data_y_6__4__3_), .SE(pe_1_5_4_n65), .CK(pe_1_5_4_net4070), .RN(
        pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_5_4_int_q_reg_h_reg_3__0_ ( .D(int_data_x_5__5__0_), .SI(
        int_data_y_6__4__0_), .SE(pe_1_5_4_n65), .CK(pe_1_5_4_net4075), .RN(
        pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_5_4_int_q_reg_h_reg_3__1_ ( .D(int_data_x_5__5__1_), .SI(
        int_data_y_6__4__1_), .SE(pe_1_5_4_n65), .CK(pe_1_5_4_net4075), .RN(
        pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_5_4_int_q_reg_h_reg_3__2_ ( .D(int_data_x_5__5__2_), .SI(
        int_data_y_6__4__2_), .SE(pe_1_5_4_n65), .CK(pe_1_5_4_net4075), .RN(
        pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_5_4_int_q_reg_h_reg_3__3_ ( .D(int_data_x_5__5__3_), .SI(
        int_data_y_6__4__3_), .SE(pe_1_5_4_n65), .CK(pe_1_5_4_net4075), .RN(
        pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_5_4_int_q_reg_h_reg_4__0_ ( .D(int_data_x_5__5__0_), .SI(
        int_data_y_6__4__0_), .SE(pe_1_5_4_n66), .CK(pe_1_5_4_net4080), .RN(
        pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_5_4_int_q_reg_h_reg_4__1_ ( .D(int_data_x_5__5__1_), .SI(
        int_data_y_6__4__1_), .SE(pe_1_5_4_n66), .CK(pe_1_5_4_net4080), .RN(
        pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_5_4_int_q_reg_h_reg_4__2_ ( .D(int_data_x_5__5__2_), .SI(
        int_data_y_6__4__2_), .SE(pe_1_5_4_n66), .CK(pe_1_5_4_net4080), .RN(
        pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_5_4_int_q_reg_h_reg_4__3_ ( .D(int_data_x_5__5__3_), .SI(
        int_data_y_6__4__3_), .SE(pe_1_5_4_n66), .CK(pe_1_5_4_net4080), .RN(
        pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_5_4_int_q_reg_h_reg_5__0_ ( .D(int_data_x_5__5__0_), .SI(
        int_data_y_6__4__0_), .SE(pe_1_5_4_n66), .CK(pe_1_5_4_net4085), .RN(
        pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_5_4_int_q_reg_h_reg_5__1_ ( .D(int_data_x_5__5__1_), .SI(
        int_data_y_6__4__1_), .SE(pe_1_5_4_n66), .CK(pe_1_5_4_net4085), .RN(
        pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_5_4_int_q_reg_h_reg_5__2_ ( .D(int_data_x_5__5__2_), .SI(
        int_data_y_6__4__2_), .SE(pe_1_5_4_n66), .CK(pe_1_5_4_net4085), .RN(
        pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_5_4_int_q_reg_h_reg_5__3_ ( .D(int_data_x_5__5__3_), .SI(
        int_data_y_6__4__3_), .SE(pe_1_5_4_n66), .CK(pe_1_5_4_net4085), .RN(
        pe_1_5_4_n72), .Q(pe_1_5_4_int_q_reg_h[3]) );
  FA_X1 pe_1_5_4_sub_81_U2_7 ( .A(int_data_res_5__4__7_), .B(pe_1_5_4_n76), 
        .CI(pe_1_5_4_sub_81_carry[7]), .S(pe_1_5_4_N77) );
  FA_X1 pe_1_5_4_sub_81_U2_6 ( .A(int_data_res_5__4__6_), .B(pe_1_5_4_n76), 
        .CI(pe_1_5_4_sub_81_carry[6]), .CO(pe_1_5_4_sub_81_carry[7]), .S(
        pe_1_5_4_N76) );
  FA_X1 pe_1_5_4_sub_81_U2_5 ( .A(int_data_res_5__4__5_), .B(pe_1_5_4_n76), 
        .CI(pe_1_5_4_sub_81_carry[5]), .CO(pe_1_5_4_sub_81_carry[6]), .S(
        pe_1_5_4_N75) );
  FA_X1 pe_1_5_4_sub_81_U2_4 ( .A(int_data_res_5__4__4_), .B(pe_1_5_4_n76), 
        .CI(pe_1_5_4_sub_81_carry[4]), .CO(pe_1_5_4_sub_81_carry[5]), .S(
        pe_1_5_4_N74) );
  FA_X1 pe_1_5_4_sub_81_U2_3 ( .A(int_data_res_5__4__3_), .B(pe_1_5_4_n76), 
        .CI(pe_1_5_4_sub_81_carry[3]), .CO(pe_1_5_4_sub_81_carry[4]), .S(
        pe_1_5_4_N73) );
  FA_X1 pe_1_5_4_sub_81_U2_2 ( .A(int_data_res_5__4__2_), .B(pe_1_5_4_n75), 
        .CI(pe_1_5_4_sub_81_carry[2]), .CO(pe_1_5_4_sub_81_carry[3]), .S(
        pe_1_5_4_N72) );
  FA_X1 pe_1_5_4_sub_81_U2_1 ( .A(int_data_res_5__4__1_), .B(pe_1_5_4_n74), 
        .CI(pe_1_5_4_sub_81_carry[1]), .CO(pe_1_5_4_sub_81_carry[2]), .S(
        pe_1_5_4_N71) );
  FA_X1 pe_1_5_4_add_83_U1_7 ( .A(int_data_res_5__4__7_), .B(
        pe_1_5_4_int_data_3_), .CI(pe_1_5_4_add_83_carry[7]), .S(pe_1_5_4_N85)
         );
  FA_X1 pe_1_5_4_add_83_U1_6 ( .A(int_data_res_5__4__6_), .B(
        pe_1_5_4_int_data_3_), .CI(pe_1_5_4_add_83_carry[6]), .CO(
        pe_1_5_4_add_83_carry[7]), .S(pe_1_5_4_N84) );
  FA_X1 pe_1_5_4_add_83_U1_5 ( .A(int_data_res_5__4__5_), .B(
        pe_1_5_4_int_data_3_), .CI(pe_1_5_4_add_83_carry[5]), .CO(
        pe_1_5_4_add_83_carry[6]), .S(pe_1_5_4_N83) );
  FA_X1 pe_1_5_4_add_83_U1_4 ( .A(int_data_res_5__4__4_), .B(
        pe_1_5_4_int_data_3_), .CI(pe_1_5_4_add_83_carry[4]), .CO(
        pe_1_5_4_add_83_carry[5]), .S(pe_1_5_4_N82) );
  FA_X1 pe_1_5_4_add_83_U1_3 ( .A(int_data_res_5__4__3_), .B(
        pe_1_5_4_int_data_3_), .CI(pe_1_5_4_add_83_carry[3]), .CO(
        pe_1_5_4_add_83_carry[4]), .S(pe_1_5_4_N81) );
  FA_X1 pe_1_5_4_add_83_U1_2 ( .A(int_data_res_5__4__2_), .B(
        pe_1_5_4_int_data_2_), .CI(pe_1_5_4_add_83_carry[2]), .CO(
        pe_1_5_4_add_83_carry[3]), .S(pe_1_5_4_N80) );
  FA_X1 pe_1_5_4_add_83_U1_1 ( .A(int_data_res_5__4__1_), .B(
        pe_1_5_4_int_data_1_), .CI(pe_1_5_4_n2), .CO(pe_1_5_4_add_83_carry[2]), 
        .S(pe_1_5_4_N79) );
  NAND3_X1 pe_1_5_4_U56 ( .A1(pe_1_5_4_n60), .A2(pe_1_5_4_n43), .A3(
        pe_1_5_4_n62), .ZN(pe_1_5_4_n40) );
  NAND3_X1 pe_1_5_4_U55 ( .A1(pe_1_5_4_n43), .A2(pe_1_5_4_n61), .A3(
        pe_1_5_4_n62), .ZN(pe_1_5_4_n39) );
  NAND3_X1 pe_1_5_4_U54 ( .A1(pe_1_5_4_n43), .A2(pe_1_5_4_n63), .A3(
        pe_1_5_4_n60), .ZN(pe_1_5_4_n38) );
  NAND3_X1 pe_1_5_4_U53 ( .A1(pe_1_5_4_n61), .A2(pe_1_5_4_n63), .A3(
        pe_1_5_4_n43), .ZN(pe_1_5_4_n37) );
  DFFR_X1 pe_1_5_4_int_q_acc_reg_6_ ( .D(pe_1_5_4_n78), .CK(pe_1_5_4_net4120), 
        .RN(pe_1_5_4_n71), .Q(int_data_res_5__4__6_) );
  DFFR_X1 pe_1_5_4_int_q_acc_reg_5_ ( .D(pe_1_5_4_n79), .CK(pe_1_5_4_net4120), 
        .RN(pe_1_5_4_n71), .Q(int_data_res_5__4__5_) );
  DFFR_X1 pe_1_5_4_int_q_acc_reg_4_ ( .D(pe_1_5_4_n80), .CK(pe_1_5_4_net4120), 
        .RN(pe_1_5_4_n71), .Q(int_data_res_5__4__4_) );
  DFFR_X1 pe_1_5_4_int_q_acc_reg_3_ ( .D(pe_1_5_4_n81), .CK(pe_1_5_4_net4120), 
        .RN(pe_1_5_4_n71), .Q(int_data_res_5__4__3_) );
  DFFR_X1 pe_1_5_4_int_q_acc_reg_2_ ( .D(pe_1_5_4_n82), .CK(pe_1_5_4_net4120), 
        .RN(pe_1_5_4_n71), .Q(int_data_res_5__4__2_) );
  DFFR_X1 pe_1_5_4_int_q_acc_reg_1_ ( .D(pe_1_5_4_n83), .CK(pe_1_5_4_net4120), 
        .RN(pe_1_5_4_n71), .Q(int_data_res_5__4__1_) );
  DFFR_X1 pe_1_5_4_int_q_acc_reg_7_ ( .D(pe_1_5_4_n77), .CK(pe_1_5_4_net4120), 
        .RN(pe_1_5_4_n71), .Q(int_data_res_5__4__7_) );
  CLKGATETST_X1 pe_1_5_4_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_5_4_n88), .SE(1'b0), .GCK(pe_1_5_4_net4059) );
  CLKGATETST_X1 pe_1_5_4_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_5_4_n87), .SE(1'b0), .GCK(pe_1_5_4_net4065) );
  CLKGATETST_X1 pe_1_5_4_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_5_4_n86), .SE(1'b0), .GCK(pe_1_5_4_net4070) );
  CLKGATETST_X1 pe_1_5_4_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_5_4_n85), .SE(1'b0), .GCK(pe_1_5_4_net4075) );
  CLKGATETST_X1 pe_1_5_4_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_5_4_n90), .SE(1'b0), .GCK(pe_1_5_4_net4080) );
  CLKGATETST_X1 pe_1_5_4_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_5_4_n89), .SE(1'b0), .GCK(pe_1_5_4_net4085) );
  CLKGATETST_X1 pe_1_5_4_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_5_4_N64), .SE(1'b0), .GCK(pe_1_5_4_net4090) );
  CLKGATETST_X1 pe_1_5_4_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_5_4_N63), .SE(1'b0), .GCK(pe_1_5_4_net4095) );
  CLKGATETST_X1 pe_1_5_4_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_5_4_N62), .SE(1'b0), .GCK(pe_1_5_4_net4100) );
  CLKGATETST_X1 pe_1_5_4_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_5_4_N61), .SE(1'b0), .GCK(pe_1_5_4_net4105) );
  CLKGATETST_X1 pe_1_5_4_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_5_4_N60), .SE(1'b0), .GCK(pe_1_5_4_net4110) );
  CLKGATETST_X1 pe_1_5_4_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_5_4_N59), .SE(1'b0), .GCK(pe_1_5_4_net4115) );
  CLKGATETST_X1 pe_1_5_4_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_5_4_N90), .SE(1'b0), .GCK(pe_1_5_4_net4120) );
  CLKBUF_X1 pe_1_5_5_U112 ( .A(pe_1_5_5_n72), .Z(pe_1_5_5_n71) );
  INV_X1 pe_1_5_5_U111 ( .A(n76), .ZN(pe_1_5_5_n70) );
  INV_X1 pe_1_5_5_U110 ( .A(n68), .ZN(pe_1_5_5_n69) );
  INV_X1 pe_1_5_5_U109 ( .A(n68), .ZN(pe_1_5_5_n68) );
  INV_X1 pe_1_5_5_U108 ( .A(n68), .ZN(pe_1_5_5_n67) );
  INV_X1 pe_1_5_5_U107 ( .A(pe_1_5_5_n69), .ZN(pe_1_5_5_n66) );
  INV_X1 pe_1_5_5_U106 ( .A(pe_1_5_5_n63), .ZN(pe_1_5_5_n62) );
  INV_X1 pe_1_5_5_U105 ( .A(pe_1_5_5_n61), .ZN(pe_1_5_5_n60) );
  INV_X1 pe_1_5_5_U104 ( .A(n28), .ZN(pe_1_5_5_n59) );
  INV_X1 pe_1_5_5_U103 ( .A(pe_1_5_5_n59), .ZN(pe_1_5_5_n58) );
  INV_X1 pe_1_5_5_U102 ( .A(n20), .ZN(pe_1_5_5_n57) );
  MUX2_X1 pe_1_5_5_U101 ( .A(pe_1_5_5_n54), .B(pe_1_5_5_n51), .S(n52), .Z(
        int_data_x_5__5__3_) );
  MUX2_X1 pe_1_5_5_U100 ( .A(pe_1_5_5_n53), .B(pe_1_5_5_n52), .S(pe_1_5_5_n62), 
        .Z(pe_1_5_5_n54) );
  MUX2_X1 pe_1_5_5_U99 ( .A(pe_1_5_5_int_q_reg_h[23]), .B(
        pe_1_5_5_int_q_reg_h[19]), .S(pe_1_5_5_n56), .Z(pe_1_5_5_n53) );
  MUX2_X1 pe_1_5_5_U98 ( .A(pe_1_5_5_int_q_reg_h[15]), .B(
        pe_1_5_5_int_q_reg_h[11]), .S(pe_1_5_5_n56), .Z(pe_1_5_5_n52) );
  MUX2_X1 pe_1_5_5_U97 ( .A(pe_1_5_5_int_q_reg_h[7]), .B(
        pe_1_5_5_int_q_reg_h[3]), .S(pe_1_5_5_n56), .Z(pe_1_5_5_n51) );
  MUX2_X1 pe_1_5_5_U96 ( .A(pe_1_5_5_n50), .B(pe_1_5_5_n47), .S(n52), .Z(
        int_data_x_5__5__2_) );
  MUX2_X1 pe_1_5_5_U95 ( .A(pe_1_5_5_n49), .B(pe_1_5_5_n48), .S(pe_1_5_5_n62), 
        .Z(pe_1_5_5_n50) );
  MUX2_X1 pe_1_5_5_U94 ( .A(pe_1_5_5_int_q_reg_h[22]), .B(
        pe_1_5_5_int_q_reg_h[18]), .S(pe_1_5_5_n56), .Z(pe_1_5_5_n49) );
  MUX2_X1 pe_1_5_5_U93 ( .A(pe_1_5_5_int_q_reg_h[14]), .B(
        pe_1_5_5_int_q_reg_h[10]), .S(pe_1_5_5_n56), .Z(pe_1_5_5_n48) );
  MUX2_X1 pe_1_5_5_U92 ( .A(pe_1_5_5_int_q_reg_h[6]), .B(
        pe_1_5_5_int_q_reg_h[2]), .S(pe_1_5_5_n56), .Z(pe_1_5_5_n47) );
  MUX2_X1 pe_1_5_5_U91 ( .A(pe_1_5_5_n46), .B(pe_1_5_5_n24), .S(n52), .Z(
        int_data_x_5__5__1_) );
  MUX2_X1 pe_1_5_5_U90 ( .A(pe_1_5_5_n45), .B(pe_1_5_5_n25), .S(pe_1_5_5_n62), 
        .Z(pe_1_5_5_n46) );
  MUX2_X1 pe_1_5_5_U89 ( .A(pe_1_5_5_int_q_reg_h[21]), .B(
        pe_1_5_5_int_q_reg_h[17]), .S(pe_1_5_5_n56), .Z(pe_1_5_5_n45) );
  MUX2_X1 pe_1_5_5_U88 ( .A(pe_1_5_5_int_q_reg_h[13]), .B(
        pe_1_5_5_int_q_reg_h[9]), .S(pe_1_5_5_n56), .Z(pe_1_5_5_n25) );
  MUX2_X1 pe_1_5_5_U87 ( .A(pe_1_5_5_int_q_reg_h[5]), .B(
        pe_1_5_5_int_q_reg_h[1]), .S(pe_1_5_5_n56), .Z(pe_1_5_5_n24) );
  MUX2_X1 pe_1_5_5_U86 ( .A(pe_1_5_5_n23), .B(pe_1_5_5_n20), .S(n52), .Z(
        int_data_x_5__5__0_) );
  MUX2_X1 pe_1_5_5_U85 ( .A(pe_1_5_5_n22), .B(pe_1_5_5_n21), .S(pe_1_5_5_n62), 
        .Z(pe_1_5_5_n23) );
  MUX2_X1 pe_1_5_5_U84 ( .A(pe_1_5_5_int_q_reg_h[20]), .B(
        pe_1_5_5_int_q_reg_h[16]), .S(pe_1_5_5_n56), .Z(pe_1_5_5_n22) );
  MUX2_X1 pe_1_5_5_U83 ( .A(pe_1_5_5_int_q_reg_h[12]), .B(
        pe_1_5_5_int_q_reg_h[8]), .S(pe_1_5_5_n56), .Z(pe_1_5_5_n21) );
  MUX2_X1 pe_1_5_5_U82 ( .A(pe_1_5_5_int_q_reg_h[4]), .B(
        pe_1_5_5_int_q_reg_h[0]), .S(pe_1_5_5_n56), .Z(pe_1_5_5_n20) );
  MUX2_X1 pe_1_5_5_U81 ( .A(pe_1_5_5_n19), .B(pe_1_5_5_n16), .S(n52), .Z(
        int_data_y_5__5__3_) );
  MUX2_X1 pe_1_5_5_U80 ( .A(pe_1_5_5_n18), .B(pe_1_5_5_n17), .S(pe_1_5_5_n62), 
        .Z(pe_1_5_5_n19) );
  MUX2_X1 pe_1_5_5_U79 ( .A(pe_1_5_5_int_q_reg_v[23]), .B(
        pe_1_5_5_int_q_reg_v[19]), .S(pe_1_5_5_n55), .Z(pe_1_5_5_n18) );
  MUX2_X1 pe_1_5_5_U78 ( .A(pe_1_5_5_int_q_reg_v[15]), .B(
        pe_1_5_5_int_q_reg_v[11]), .S(pe_1_5_5_n55), .Z(pe_1_5_5_n17) );
  MUX2_X1 pe_1_5_5_U77 ( .A(pe_1_5_5_int_q_reg_v[7]), .B(
        pe_1_5_5_int_q_reg_v[3]), .S(pe_1_5_5_n55), .Z(pe_1_5_5_n16) );
  MUX2_X1 pe_1_5_5_U76 ( .A(pe_1_5_5_n15), .B(pe_1_5_5_n12), .S(n52), .Z(
        int_data_y_5__5__2_) );
  MUX2_X1 pe_1_5_5_U75 ( .A(pe_1_5_5_n14), .B(pe_1_5_5_n13), .S(pe_1_5_5_n62), 
        .Z(pe_1_5_5_n15) );
  MUX2_X1 pe_1_5_5_U74 ( .A(pe_1_5_5_int_q_reg_v[22]), .B(
        pe_1_5_5_int_q_reg_v[18]), .S(pe_1_5_5_n55), .Z(pe_1_5_5_n14) );
  MUX2_X1 pe_1_5_5_U73 ( .A(pe_1_5_5_int_q_reg_v[14]), .B(
        pe_1_5_5_int_q_reg_v[10]), .S(pe_1_5_5_n55), .Z(pe_1_5_5_n13) );
  MUX2_X1 pe_1_5_5_U72 ( .A(pe_1_5_5_int_q_reg_v[6]), .B(
        pe_1_5_5_int_q_reg_v[2]), .S(pe_1_5_5_n55), .Z(pe_1_5_5_n12) );
  MUX2_X1 pe_1_5_5_U71 ( .A(pe_1_5_5_n11), .B(pe_1_5_5_n8), .S(n52), .Z(
        int_data_y_5__5__1_) );
  MUX2_X1 pe_1_5_5_U70 ( .A(pe_1_5_5_n10), .B(pe_1_5_5_n9), .S(pe_1_5_5_n62), 
        .Z(pe_1_5_5_n11) );
  MUX2_X1 pe_1_5_5_U69 ( .A(pe_1_5_5_int_q_reg_v[21]), .B(
        pe_1_5_5_int_q_reg_v[17]), .S(pe_1_5_5_n55), .Z(pe_1_5_5_n10) );
  MUX2_X1 pe_1_5_5_U68 ( .A(pe_1_5_5_int_q_reg_v[13]), .B(
        pe_1_5_5_int_q_reg_v[9]), .S(pe_1_5_5_n55), .Z(pe_1_5_5_n9) );
  MUX2_X1 pe_1_5_5_U67 ( .A(pe_1_5_5_int_q_reg_v[5]), .B(
        pe_1_5_5_int_q_reg_v[1]), .S(pe_1_5_5_n55), .Z(pe_1_5_5_n8) );
  MUX2_X1 pe_1_5_5_U66 ( .A(pe_1_5_5_n7), .B(pe_1_5_5_n4), .S(n52), .Z(
        int_data_y_5__5__0_) );
  MUX2_X1 pe_1_5_5_U65 ( .A(pe_1_5_5_n6), .B(pe_1_5_5_n5), .S(pe_1_5_5_n62), 
        .Z(pe_1_5_5_n7) );
  MUX2_X1 pe_1_5_5_U64 ( .A(pe_1_5_5_int_q_reg_v[20]), .B(
        pe_1_5_5_int_q_reg_v[16]), .S(pe_1_5_5_n55), .Z(pe_1_5_5_n6) );
  MUX2_X1 pe_1_5_5_U63 ( .A(pe_1_5_5_int_q_reg_v[12]), .B(
        pe_1_5_5_int_q_reg_v[8]), .S(pe_1_5_5_n55), .Z(pe_1_5_5_n5) );
  MUX2_X1 pe_1_5_5_U62 ( .A(pe_1_5_5_int_q_reg_v[4]), .B(
        pe_1_5_5_int_q_reg_v[0]), .S(pe_1_5_5_n55), .Z(pe_1_5_5_n4) );
  AOI222_X1 pe_1_5_5_U61 ( .A1(int_data_res_6__5__2_), .A2(pe_1_5_5_n64), .B1(
        pe_1_5_5_N80), .B2(pe_1_5_5_n27), .C1(pe_1_5_5_N72), .C2(pe_1_5_5_n28), 
        .ZN(pe_1_5_5_n33) );
  INV_X1 pe_1_5_5_U60 ( .A(pe_1_5_5_n33), .ZN(pe_1_5_5_n82) );
  AOI222_X1 pe_1_5_5_U59 ( .A1(int_data_res_6__5__6_), .A2(pe_1_5_5_n64), .B1(
        pe_1_5_5_N84), .B2(pe_1_5_5_n27), .C1(pe_1_5_5_N76), .C2(pe_1_5_5_n28), 
        .ZN(pe_1_5_5_n29) );
  INV_X1 pe_1_5_5_U58 ( .A(pe_1_5_5_n29), .ZN(pe_1_5_5_n78) );
  XNOR2_X1 pe_1_5_5_U57 ( .A(pe_1_5_5_n73), .B(int_data_res_5__5__0_), .ZN(
        pe_1_5_5_N70) );
  AOI222_X1 pe_1_5_5_U52 ( .A1(int_data_res_6__5__0_), .A2(pe_1_5_5_n64), .B1(
        pe_1_5_5_n1), .B2(pe_1_5_5_n27), .C1(pe_1_5_5_N70), .C2(pe_1_5_5_n28), 
        .ZN(pe_1_5_5_n35) );
  INV_X1 pe_1_5_5_U51 ( .A(pe_1_5_5_n35), .ZN(pe_1_5_5_n84) );
  AOI222_X1 pe_1_5_5_U50 ( .A1(int_data_res_6__5__1_), .A2(pe_1_5_5_n64), .B1(
        pe_1_5_5_N79), .B2(pe_1_5_5_n27), .C1(pe_1_5_5_N71), .C2(pe_1_5_5_n28), 
        .ZN(pe_1_5_5_n34) );
  INV_X1 pe_1_5_5_U49 ( .A(pe_1_5_5_n34), .ZN(pe_1_5_5_n83) );
  AOI222_X1 pe_1_5_5_U48 ( .A1(int_data_res_6__5__3_), .A2(pe_1_5_5_n64), .B1(
        pe_1_5_5_N81), .B2(pe_1_5_5_n27), .C1(pe_1_5_5_N73), .C2(pe_1_5_5_n28), 
        .ZN(pe_1_5_5_n32) );
  INV_X1 pe_1_5_5_U47 ( .A(pe_1_5_5_n32), .ZN(pe_1_5_5_n81) );
  AOI222_X1 pe_1_5_5_U46 ( .A1(int_data_res_6__5__4_), .A2(pe_1_5_5_n64), .B1(
        pe_1_5_5_N82), .B2(pe_1_5_5_n27), .C1(pe_1_5_5_N74), .C2(pe_1_5_5_n28), 
        .ZN(pe_1_5_5_n31) );
  INV_X1 pe_1_5_5_U45 ( .A(pe_1_5_5_n31), .ZN(pe_1_5_5_n80) );
  AOI222_X1 pe_1_5_5_U44 ( .A1(int_data_res_6__5__5_), .A2(pe_1_5_5_n64), .B1(
        pe_1_5_5_N83), .B2(pe_1_5_5_n27), .C1(pe_1_5_5_N75), .C2(pe_1_5_5_n28), 
        .ZN(pe_1_5_5_n30) );
  INV_X1 pe_1_5_5_U43 ( .A(pe_1_5_5_n30), .ZN(pe_1_5_5_n79) );
  NAND2_X1 pe_1_5_5_U42 ( .A1(pe_1_5_5_int_data_0_), .A2(pe_1_5_5_n3), .ZN(
        pe_1_5_5_sub_81_carry[1]) );
  INV_X1 pe_1_5_5_U41 ( .A(pe_1_5_5_int_data_1_), .ZN(pe_1_5_5_n74) );
  INV_X1 pe_1_5_5_U40 ( .A(pe_1_5_5_int_data_2_), .ZN(pe_1_5_5_n75) );
  AND2_X1 pe_1_5_5_U39 ( .A1(pe_1_5_5_int_data_0_), .A2(int_data_res_5__5__0_), 
        .ZN(pe_1_5_5_n2) );
  AOI222_X1 pe_1_5_5_U38 ( .A1(pe_1_5_5_n64), .A2(int_data_res_6__5__7_), .B1(
        pe_1_5_5_N85), .B2(pe_1_5_5_n27), .C1(pe_1_5_5_N77), .C2(pe_1_5_5_n28), 
        .ZN(pe_1_5_5_n26) );
  INV_X1 pe_1_5_5_U37 ( .A(pe_1_5_5_n26), .ZN(pe_1_5_5_n77) );
  NOR3_X1 pe_1_5_5_U36 ( .A1(pe_1_5_5_n59), .A2(pe_1_5_5_n65), .A3(int_ckg[18]), .ZN(pe_1_5_5_n36) );
  OR2_X1 pe_1_5_5_U35 ( .A1(pe_1_5_5_n36), .A2(pe_1_5_5_n64), .ZN(pe_1_5_5_N90) );
  INV_X1 pe_1_5_5_U34 ( .A(n40), .ZN(pe_1_5_5_n63) );
  AND2_X1 pe_1_5_5_U33 ( .A1(int_data_x_5__5__2_), .A2(pe_1_5_5_n58), .ZN(
        pe_1_5_5_int_data_2_) );
  AND2_X1 pe_1_5_5_U32 ( .A1(int_data_x_5__5__1_), .A2(pe_1_5_5_n58), .ZN(
        pe_1_5_5_int_data_1_) );
  AND2_X1 pe_1_5_5_U31 ( .A1(int_data_x_5__5__3_), .A2(pe_1_5_5_n58), .ZN(
        pe_1_5_5_int_data_3_) );
  BUF_X1 pe_1_5_5_U30 ( .A(n62), .Z(pe_1_5_5_n64) );
  INV_X1 pe_1_5_5_U29 ( .A(n34), .ZN(pe_1_5_5_n61) );
  AND2_X1 pe_1_5_5_U28 ( .A1(int_data_x_5__5__0_), .A2(pe_1_5_5_n58), .ZN(
        pe_1_5_5_int_data_0_) );
  NAND2_X1 pe_1_5_5_U27 ( .A1(pe_1_5_5_n44), .A2(pe_1_5_5_n61), .ZN(
        pe_1_5_5_n41) );
  AND3_X1 pe_1_5_5_U26 ( .A1(n76), .A2(pe_1_5_5_n63), .A3(n52), .ZN(
        pe_1_5_5_n44) );
  INV_X1 pe_1_5_5_U25 ( .A(pe_1_5_5_int_data_3_), .ZN(pe_1_5_5_n76) );
  NOR2_X1 pe_1_5_5_U24 ( .A1(pe_1_5_5_n70), .A2(n52), .ZN(pe_1_5_5_n43) );
  NOR2_X1 pe_1_5_5_U23 ( .A1(pe_1_5_5_n57), .A2(pe_1_5_5_n64), .ZN(
        pe_1_5_5_n28) );
  NOR2_X1 pe_1_5_5_U22 ( .A1(n20), .A2(pe_1_5_5_n64), .ZN(pe_1_5_5_n27) );
  INV_X1 pe_1_5_5_U21 ( .A(pe_1_5_5_int_data_0_), .ZN(pe_1_5_5_n73) );
  INV_X1 pe_1_5_5_U20 ( .A(pe_1_5_5_n41), .ZN(pe_1_5_5_n90) );
  INV_X1 pe_1_5_5_U19 ( .A(pe_1_5_5_n37), .ZN(pe_1_5_5_n88) );
  INV_X1 pe_1_5_5_U18 ( .A(pe_1_5_5_n38), .ZN(pe_1_5_5_n87) );
  INV_X1 pe_1_5_5_U17 ( .A(pe_1_5_5_n39), .ZN(pe_1_5_5_n86) );
  NOR2_X1 pe_1_5_5_U16 ( .A1(pe_1_5_5_n68), .A2(pe_1_5_5_n42), .ZN(
        pe_1_5_5_N59) );
  NOR2_X1 pe_1_5_5_U15 ( .A1(pe_1_5_5_n68), .A2(pe_1_5_5_n41), .ZN(
        pe_1_5_5_N60) );
  NOR2_X1 pe_1_5_5_U14 ( .A1(pe_1_5_5_n68), .A2(pe_1_5_5_n38), .ZN(
        pe_1_5_5_N63) );
  NOR2_X1 pe_1_5_5_U13 ( .A1(pe_1_5_5_n67), .A2(pe_1_5_5_n40), .ZN(
        pe_1_5_5_N61) );
  NOR2_X1 pe_1_5_5_U12 ( .A1(pe_1_5_5_n67), .A2(pe_1_5_5_n39), .ZN(
        pe_1_5_5_N62) );
  NOR2_X1 pe_1_5_5_U11 ( .A1(pe_1_5_5_n37), .A2(pe_1_5_5_n67), .ZN(
        pe_1_5_5_N64) );
  NAND2_X1 pe_1_5_5_U10 ( .A1(pe_1_5_5_n44), .A2(pe_1_5_5_n60), .ZN(
        pe_1_5_5_n42) );
  BUF_X1 pe_1_5_5_U9 ( .A(pe_1_5_5_n60), .Z(pe_1_5_5_n55) );
  INV_X1 pe_1_5_5_U8 ( .A(pe_1_5_5_n69), .ZN(pe_1_5_5_n65) );
  BUF_X1 pe_1_5_5_U7 ( .A(pe_1_5_5_n60), .Z(pe_1_5_5_n56) );
  INV_X1 pe_1_5_5_U6 ( .A(pe_1_5_5_n42), .ZN(pe_1_5_5_n89) );
  INV_X1 pe_1_5_5_U5 ( .A(pe_1_5_5_n40), .ZN(pe_1_5_5_n85) );
  INV_X2 pe_1_5_5_U4 ( .A(n84), .ZN(pe_1_5_5_n72) );
  XOR2_X1 pe_1_5_5_U3 ( .A(pe_1_5_5_int_data_0_), .B(int_data_res_5__5__0_), 
        .Z(pe_1_5_5_n1) );
  DFFR_X1 pe_1_5_5_int_q_acc_reg_0_ ( .D(pe_1_5_5_n84), .CK(pe_1_5_5_net4042), 
        .RN(pe_1_5_5_n72), .Q(int_data_res_5__5__0_), .QN(pe_1_5_5_n3) );
  DFFR_X1 pe_1_5_5_int_q_reg_v_reg_0__0_ ( .D(int_data_y_6__5__0_), .CK(
        pe_1_5_5_net4012), .RN(pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_v[20]) );
  DFFR_X1 pe_1_5_5_int_q_reg_v_reg_0__1_ ( .D(int_data_y_6__5__1_), .CK(
        pe_1_5_5_net4012), .RN(pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_v[21]) );
  DFFR_X1 pe_1_5_5_int_q_reg_v_reg_0__2_ ( .D(int_data_y_6__5__2_), .CK(
        pe_1_5_5_net4012), .RN(pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_v[22]) );
  DFFR_X1 pe_1_5_5_int_q_reg_v_reg_0__3_ ( .D(int_data_y_6__5__3_), .CK(
        pe_1_5_5_net4012), .RN(pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_v[23]) );
  DFFR_X1 pe_1_5_5_int_q_reg_v_reg_1__0_ ( .D(int_data_y_6__5__0_), .CK(
        pe_1_5_5_net4017), .RN(pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_v[16]) );
  DFFR_X1 pe_1_5_5_int_q_reg_v_reg_1__1_ ( .D(int_data_y_6__5__1_), .CK(
        pe_1_5_5_net4017), .RN(pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_v[17]) );
  DFFR_X1 pe_1_5_5_int_q_reg_v_reg_1__2_ ( .D(int_data_y_6__5__2_), .CK(
        pe_1_5_5_net4017), .RN(pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_v[18]) );
  DFFR_X1 pe_1_5_5_int_q_reg_v_reg_1__3_ ( .D(int_data_y_6__5__3_), .CK(
        pe_1_5_5_net4017), .RN(pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_v[19]) );
  DFFR_X1 pe_1_5_5_int_q_reg_v_reg_2__0_ ( .D(int_data_y_6__5__0_), .CK(
        pe_1_5_5_net4022), .RN(pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_v[12]) );
  DFFR_X1 pe_1_5_5_int_q_reg_v_reg_2__1_ ( .D(int_data_y_6__5__1_), .CK(
        pe_1_5_5_net4022), .RN(pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_v[13]) );
  DFFR_X1 pe_1_5_5_int_q_reg_v_reg_2__2_ ( .D(int_data_y_6__5__2_), .CK(
        pe_1_5_5_net4022), .RN(pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_v[14]) );
  DFFR_X1 pe_1_5_5_int_q_reg_v_reg_2__3_ ( .D(int_data_y_6__5__3_), .CK(
        pe_1_5_5_net4022), .RN(pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_v[15]) );
  DFFR_X1 pe_1_5_5_int_q_reg_v_reg_3__0_ ( .D(int_data_y_6__5__0_), .CK(
        pe_1_5_5_net4027), .RN(pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_v[8]) );
  DFFR_X1 pe_1_5_5_int_q_reg_v_reg_3__1_ ( .D(int_data_y_6__5__1_), .CK(
        pe_1_5_5_net4027), .RN(pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_v[9]) );
  DFFR_X1 pe_1_5_5_int_q_reg_v_reg_3__2_ ( .D(int_data_y_6__5__2_), .CK(
        pe_1_5_5_net4027), .RN(pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_v[10]) );
  DFFR_X1 pe_1_5_5_int_q_reg_v_reg_3__3_ ( .D(int_data_y_6__5__3_), .CK(
        pe_1_5_5_net4027), .RN(pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_v[11]) );
  DFFR_X1 pe_1_5_5_int_q_reg_v_reg_4__0_ ( .D(int_data_y_6__5__0_), .CK(
        pe_1_5_5_net4032), .RN(pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_v[4]) );
  DFFR_X1 pe_1_5_5_int_q_reg_v_reg_4__1_ ( .D(int_data_y_6__5__1_), .CK(
        pe_1_5_5_net4032), .RN(pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_v[5]) );
  DFFR_X1 pe_1_5_5_int_q_reg_v_reg_4__2_ ( .D(int_data_y_6__5__2_), .CK(
        pe_1_5_5_net4032), .RN(pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_v[6]) );
  DFFR_X1 pe_1_5_5_int_q_reg_v_reg_4__3_ ( .D(int_data_y_6__5__3_), .CK(
        pe_1_5_5_net4032), .RN(pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_v[7]) );
  DFFR_X1 pe_1_5_5_int_q_reg_v_reg_5__0_ ( .D(int_data_y_6__5__0_), .CK(
        pe_1_5_5_net4037), .RN(pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_v[0]) );
  DFFR_X1 pe_1_5_5_int_q_reg_v_reg_5__1_ ( .D(int_data_y_6__5__1_), .CK(
        pe_1_5_5_net4037), .RN(pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_v[1]) );
  DFFR_X1 pe_1_5_5_int_q_reg_v_reg_5__2_ ( .D(int_data_y_6__5__2_), .CK(
        pe_1_5_5_net4037), .RN(pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_v[2]) );
  DFFR_X1 pe_1_5_5_int_q_reg_v_reg_5__3_ ( .D(int_data_y_6__5__3_), .CK(
        pe_1_5_5_net4037), .RN(pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_5_5_int_q_reg_h_reg_0__0_ ( .D(int_data_x_5__6__0_), .SI(
        int_data_y_6__5__0_), .SE(pe_1_5_5_n65), .CK(pe_1_5_5_net3981), .RN(
        pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_5_5_int_q_reg_h_reg_0__1_ ( .D(int_data_x_5__6__1_), .SI(
        int_data_y_6__5__1_), .SE(pe_1_5_5_n65), .CK(pe_1_5_5_net3981), .RN(
        pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_5_5_int_q_reg_h_reg_0__2_ ( .D(int_data_x_5__6__2_), .SI(
        int_data_y_6__5__2_), .SE(pe_1_5_5_n65), .CK(pe_1_5_5_net3981), .RN(
        pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_5_5_int_q_reg_h_reg_0__3_ ( .D(int_data_x_5__6__3_), .SI(
        int_data_y_6__5__3_), .SE(pe_1_5_5_n65), .CK(pe_1_5_5_net3981), .RN(
        pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_5_5_int_q_reg_h_reg_1__0_ ( .D(int_data_x_5__6__0_), .SI(
        int_data_y_6__5__0_), .SE(pe_1_5_5_n65), .CK(pe_1_5_5_net3987), .RN(
        pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_5_5_int_q_reg_h_reg_1__1_ ( .D(int_data_x_5__6__1_), .SI(
        int_data_y_6__5__1_), .SE(pe_1_5_5_n65), .CK(pe_1_5_5_net3987), .RN(
        pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_5_5_int_q_reg_h_reg_1__2_ ( .D(int_data_x_5__6__2_), .SI(
        int_data_y_6__5__2_), .SE(pe_1_5_5_n65), .CK(pe_1_5_5_net3987), .RN(
        pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_5_5_int_q_reg_h_reg_1__3_ ( .D(int_data_x_5__6__3_), .SI(
        int_data_y_6__5__3_), .SE(pe_1_5_5_n65), .CK(pe_1_5_5_net3987), .RN(
        pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_5_5_int_q_reg_h_reg_2__0_ ( .D(int_data_x_5__6__0_), .SI(
        int_data_y_6__5__0_), .SE(pe_1_5_5_n65), .CK(pe_1_5_5_net3992), .RN(
        pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_5_5_int_q_reg_h_reg_2__1_ ( .D(int_data_x_5__6__1_), .SI(
        int_data_y_6__5__1_), .SE(pe_1_5_5_n65), .CK(pe_1_5_5_net3992), .RN(
        pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_5_5_int_q_reg_h_reg_2__2_ ( .D(int_data_x_5__6__2_), .SI(
        int_data_y_6__5__2_), .SE(pe_1_5_5_n65), .CK(pe_1_5_5_net3992), .RN(
        pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_5_5_int_q_reg_h_reg_2__3_ ( .D(int_data_x_5__6__3_), .SI(
        int_data_y_6__5__3_), .SE(pe_1_5_5_n65), .CK(pe_1_5_5_net3992), .RN(
        pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_5_5_int_q_reg_h_reg_3__0_ ( .D(int_data_x_5__6__0_), .SI(
        int_data_y_6__5__0_), .SE(pe_1_5_5_n65), .CK(pe_1_5_5_net3997), .RN(
        pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_5_5_int_q_reg_h_reg_3__1_ ( .D(int_data_x_5__6__1_), .SI(
        int_data_y_6__5__1_), .SE(pe_1_5_5_n65), .CK(pe_1_5_5_net3997), .RN(
        pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_5_5_int_q_reg_h_reg_3__2_ ( .D(int_data_x_5__6__2_), .SI(
        int_data_y_6__5__2_), .SE(pe_1_5_5_n65), .CK(pe_1_5_5_net3997), .RN(
        pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_5_5_int_q_reg_h_reg_3__3_ ( .D(int_data_x_5__6__3_), .SI(
        int_data_y_6__5__3_), .SE(pe_1_5_5_n65), .CK(pe_1_5_5_net3997), .RN(
        pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_5_5_int_q_reg_h_reg_4__0_ ( .D(int_data_x_5__6__0_), .SI(
        int_data_y_6__5__0_), .SE(pe_1_5_5_n66), .CK(pe_1_5_5_net4002), .RN(
        pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_5_5_int_q_reg_h_reg_4__1_ ( .D(int_data_x_5__6__1_), .SI(
        int_data_y_6__5__1_), .SE(pe_1_5_5_n66), .CK(pe_1_5_5_net4002), .RN(
        pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_5_5_int_q_reg_h_reg_4__2_ ( .D(int_data_x_5__6__2_), .SI(
        int_data_y_6__5__2_), .SE(pe_1_5_5_n66), .CK(pe_1_5_5_net4002), .RN(
        pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_5_5_int_q_reg_h_reg_4__3_ ( .D(int_data_x_5__6__3_), .SI(
        int_data_y_6__5__3_), .SE(pe_1_5_5_n66), .CK(pe_1_5_5_net4002), .RN(
        pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_5_5_int_q_reg_h_reg_5__0_ ( .D(int_data_x_5__6__0_), .SI(
        int_data_y_6__5__0_), .SE(pe_1_5_5_n66), .CK(pe_1_5_5_net4007), .RN(
        pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_5_5_int_q_reg_h_reg_5__1_ ( .D(int_data_x_5__6__1_), .SI(
        int_data_y_6__5__1_), .SE(pe_1_5_5_n66), .CK(pe_1_5_5_net4007), .RN(
        pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_5_5_int_q_reg_h_reg_5__2_ ( .D(int_data_x_5__6__2_), .SI(
        int_data_y_6__5__2_), .SE(pe_1_5_5_n66), .CK(pe_1_5_5_net4007), .RN(
        pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_5_5_int_q_reg_h_reg_5__3_ ( .D(int_data_x_5__6__3_), .SI(
        int_data_y_6__5__3_), .SE(pe_1_5_5_n66), .CK(pe_1_5_5_net4007), .RN(
        pe_1_5_5_n72), .Q(pe_1_5_5_int_q_reg_h[3]) );
  FA_X1 pe_1_5_5_sub_81_U2_7 ( .A(int_data_res_5__5__7_), .B(pe_1_5_5_n76), 
        .CI(pe_1_5_5_sub_81_carry[7]), .S(pe_1_5_5_N77) );
  FA_X1 pe_1_5_5_sub_81_U2_6 ( .A(int_data_res_5__5__6_), .B(pe_1_5_5_n76), 
        .CI(pe_1_5_5_sub_81_carry[6]), .CO(pe_1_5_5_sub_81_carry[7]), .S(
        pe_1_5_5_N76) );
  FA_X1 pe_1_5_5_sub_81_U2_5 ( .A(int_data_res_5__5__5_), .B(pe_1_5_5_n76), 
        .CI(pe_1_5_5_sub_81_carry[5]), .CO(pe_1_5_5_sub_81_carry[6]), .S(
        pe_1_5_5_N75) );
  FA_X1 pe_1_5_5_sub_81_U2_4 ( .A(int_data_res_5__5__4_), .B(pe_1_5_5_n76), 
        .CI(pe_1_5_5_sub_81_carry[4]), .CO(pe_1_5_5_sub_81_carry[5]), .S(
        pe_1_5_5_N74) );
  FA_X1 pe_1_5_5_sub_81_U2_3 ( .A(int_data_res_5__5__3_), .B(pe_1_5_5_n76), 
        .CI(pe_1_5_5_sub_81_carry[3]), .CO(pe_1_5_5_sub_81_carry[4]), .S(
        pe_1_5_5_N73) );
  FA_X1 pe_1_5_5_sub_81_U2_2 ( .A(int_data_res_5__5__2_), .B(pe_1_5_5_n75), 
        .CI(pe_1_5_5_sub_81_carry[2]), .CO(pe_1_5_5_sub_81_carry[3]), .S(
        pe_1_5_5_N72) );
  FA_X1 pe_1_5_5_sub_81_U2_1 ( .A(int_data_res_5__5__1_), .B(pe_1_5_5_n74), 
        .CI(pe_1_5_5_sub_81_carry[1]), .CO(pe_1_5_5_sub_81_carry[2]), .S(
        pe_1_5_5_N71) );
  FA_X1 pe_1_5_5_add_83_U1_7 ( .A(int_data_res_5__5__7_), .B(
        pe_1_5_5_int_data_3_), .CI(pe_1_5_5_add_83_carry[7]), .S(pe_1_5_5_N85)
         );
  FA_X1 pe_1_5_5_add_83_U1_6 ( .A(int_data_res_5__5__6_), .B(
        pe_1_5_5_int_data_3_), .CI(pe_1_5_5_add_83_carry[6]), .CO(
        pe_1_5_5_add_83_carry[7]), .S(pe_1_5_5_N84) );
  FA_X1 pe_1_5_5_add_83_U1_5 ( .A(int_data_res_5__5__5_), .B(
        pe_1_5_5_int_data_3_), .CI(pe_1_5_5_add_83_carry[5]), .CO(
        pe_1_5_5_add_83_carry[6]), .S(pe_1_5_5_N83) );
  FA_X1 pe_1_5_5_add_83_U1_4 ( .A(int_data_res_5__5__4_), .B(
        pe_1_5_5_int_data_3_), .CI(pe_1_5_5_add_83_carry[4]), .CO(
        pe_1_5_5_add_83_carry[5]), .S(pe_1_5_5_N82) );
  FA_X1 pe_1_5_5_add_83_U1_3 ( .A(int_data_res_5__5__3_), .B(
        pe_1_5_5_int_data_3_), .CI(pe_1_5_5_add_83_carry[3]), .CO(
        pe_1_5_5_add_83_carry[4]), .S(pe_1_5_5_N81) );
  FA_X1 pe_1_5_5_add_83_U1_2 ( .A(int_data_res_5__5__2_), .B(
        pe_1_5_5_int_data_2_), .CI(pe_1_5_5_add_83_carry[2]), .CO(
        pe_1_5_5_add_83_carry[3]), .S(pe_1_5_5_N80) );
  FA_X1 pe_1_5_5_add_83_U1_1 ( .A(int_data_res_5__5__1_), .B(
        pe_1_5_5_int_data_1_), .CI(pe_1_5_5_n2), .CO(pe_1_5_5_add_83_carry[2]), 
        .S(pe_1_5_5_N79) );
  NAND3_X1 pe_1_5_5_U56 ( .A1(pe_1_5_5_n60), .A2(pe_1_5_5_n43), .A3(
        pe_1_5_5_n62), .ZN(pe_1_5_5_n40) );
  NAND3_X1 pe_1_5_5_U55 ( .A1(pe_1_5_5_n43), .A2(pe_1_5_5_n61), .A3(
        pe_1_5_5_n62), .ZN(pe_1_5_5_n39) );
  NAND3_X1 pe_1_5_5_U54 ( .A1(pe_1_5_5_n43), .A2(pe_1_5_5_n63), .A3(
        pe_1_5_5_n60), .ZN(pe_1_5_5_n38) );
  NAND3_X1 pe_1_5_5_U53 ( .A1(pe_1_5_5_n61), .A2(pe_1_5_5_n63), .A3(
        pe_1_5_5_n43), .ZN(pe_1_5_5_n37) );
  DFFR_X1 pe_1_5_5_int_q_acc_reg_6_ ( .D(pe_1_5_5_n78), .CK(pe_1_5_5_net4042), 
        .RN(pe_1_5_5_n71), .Q(int_data_res_5__5__6_) );
  DFFR_X1 pe_1_5_5_int_q_acc_reg_5_ ( .D(pe_1_5_5_n79), .CK(pe_1_5_5_net4042), 
        .RN(pe_1_5_5_n71), .Q(int_data_res_5__5__5_) );
  DFFR_X1 pe_1_5_5_int_q_acc_reg_4_ ( .D(pe_1_5_5_n80), .CK(pe_1_5_5_net4042), 
        .RN(pe_1_5_5_n71), .Q(int_data_res_5__5__4_) );
  DFFR_X1 pe_1_5_5_int_q_acc_reg_3_ ( .D(pe_1_5_5_n81), .CK(pe_1_5_5_net4042), 
        .RN(pe_1_5_5_n71), .Q(int_data_res_5__5__3_) );
  DFFR_X1 pe_1_5_5_int_q_acc_reg_2_ ( .D(pe_1_5_5_n82), .CK(pe_1_5_5_net4042), 
        .RN(pe_1_5_5_n71), .Q(int_data_res_5__5__2_) );
  DFFR_X1 pe_1_5_5_int_q_acc_reg_1_ ( .D(pe_1_5_5_n83), .CK(pe_1_5_5_net4042), 
        .RN(pe_1_5_5_n71), .Q(int_data_res_5__5__1_) );
  DFFR_X1 pe_1_5_5_int_q_acc_reg_7_ ( .D(pe_1_5_5_n77), .CK(pe_1_5_5_net4042), 
        .RN(pe_1_5_5_n71), .Q(int_data_res_5__5__7_) );
  CLKGATETST_X1 pe_1_5_5_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_5_5_n88), .SE(1'b0), .GCK(pe_1_5_5_net3981) );
  CLKGATETST_X1 pe_1_5_5_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_5_5_n87), .SE(1'b0), .GCK(pe_1_5_5_net3987) );
  CLKGATETST_X1 pe_1_5_5_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_5_5_n86), .SE(1'b0), .GCK(pe_1_5_5_net3992) );
  CLKGATETST_X1 pe_1_5_5_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_5_5_n85), .SE(1'b0), .GCK(pe_1_5_5_net3997) );
  CLKGATETST_X1 pe_1_5_5_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_5_5_n90), .SE(1'b0), .GCK(pe_1_5_5_net4002) );
  CLKGATETST_X1 pe_1_5_5_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_5_5_n89), .SE(1'b0), .GCK(pe_1_5_5_net4007) );
  CLKGATETST_X1 pe_1_5_5_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_5_5_N64), .SE(1'b0), .GCK(pe_1_5_5_net4012) );
  CLKGATETST_X1 pe_1_5_5_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_5_5_N63), .SE(1'b0), .GCK(pe_1_5_5_net4017) );
  CLKGATETST_X1 pe_1_5_5_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_5_5_N62), .SE(1'b0), .GCK(pe_1_5_5_net4022) );
  CLKGATETST_X1 pe_1_5_5_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_5_5_N61), .SE(1'b0), .GCK(pe_1_5_5_net4027) );
  CLKGATETST_X1 pe_1_5_5_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_5_5_N60), .SE(1'b0), .GCK(pe_1_5_5_net4032) );
  CLKGATETST_X1 pe_1_5_5_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_5_5_N59), .SE(1'b0), .GCK(pe_1_5_5_net4037) );
  CLKGATETST_X1 pe_1_5_5_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_5_5_N90), .SE(1'b0), .GCK(pe_1_5_5_net4042) );
  CLKBUF_X1 pe_1_5_6_U112 ( .A(pe_1_5_6_n72), .Z(pe_1_5_6_n71) );
  INV_X1 pe_1_5_6_U111 ( .A(n76), .ZN(pe_1_5_6_n70) );
  INV_X1 pe_1_5_6_U110 ( .A(n68), .ZN(pe_1_5_6_n69) );
  INV_X1 pe_1_5_6_U109 ( .A(n68), .ZN(pe_1_5_6_n68) );
  INV_X1 pe_1_5_6_U108 ( .A(n68), .ZN(pe_1_5_6_n67) );
  INV_X1 pe_1_5_6_U107 ( .A(pe_1_5_6_n69), .ZN(pe_1_5_6_n66) );
  INV_X1 pe_1_5_6_U106 ( .A(pe_1_5_6_n63), .ZN(pe_1_5_6_n62) );
  INV_X1 pe_1_5_6_U105 ( .A(pe_1_5_6_n61), .ZN(pe_1_5_6_n60) );
  INV_X1 pe_1_5_6_U104 ( .A(n28), .ZN(pe_1_5_6_n59) );
  INV_X1 pe_1_5_6_U103 ( .A(pe_1_5_6_n59), .ZN(pe_1_5_6_n58) );
  INV_X1 pe_1_5_6_U102 ( .A(n20), .ZN(pe_1_5_6_n57) );
  MUX2_X1 pe_1_5_6_U101 ( .A(pe_1_5_6_n54), .B(pe_1_5_6_n51), .S(n52), .Z(
        int_data_x_5__6__3_) );
  MUX2_X1 pe_1_5_6_U100 ( .A(pe_1_5_6_n53), .B(pe_1_5_6_n52), .S(pe_1_5_6_n62), 
        .Z(pe_1_5_6_n54) );
  MUX2_X1 pe_1_5_6_U99 ( .A(pe_1_5_6_int_q_reg_h[23]), .B(
        pe_1_5_6_int_q_reg_h[19]), .S(pe_1_5_6_n56), .Z(pe_1_5_6_n53) );
  MUX2_X1 pe_1_5_6_U98 ( .A(pe_1_5_6_int_q_reg_h[15]), .B(
        pe_1_5_6_int_q_reg_h[11]), .S(pe_1_5_6_n56), .Z(pe_1_5_6_n52) );
  MUX2_X1 pe_1_5_6_U97 ( .A(pe_1_5_6_int_q_reg_h[7]), .B(
        pe_1_5_6_int_q_reg_h[3]), .S(pe_1_5_6_n56), .Z(pe_1_5_6_n51) );
  MUX2_X1 pe_1_5_6_U96 ( .A(pe_1_5_6_n50), .B(pe_1_5_6_n47), .S(n52), .Z(
        int_data_x_5__6__2_) );
  MUX2_X1 pe_1_5_6_U95 ( .A(pe_1_5_6_n49), .B(pe_1_5_6_n48), .S(pe_1_5_6_n62), 
        .Z(pe_1_5_6_n50) );
  MUX2_X1 pe_1_5_6_U94 ( .A(pe_1_5_6_int_q_reg_h[22]), .B(
        pe_1_5_6_int_q_reg_h[18]), .S(pe_1_5_6_n56), .Z(pe_1_5_6_n49) );
  MUX2_X1 pe_1_5_6_U93 ( .A(pe_1_5_6_int_q_reg_h[14]), .B(
        pe_1_5_6_int_q_reg_h[10]), .S(pe_1_5_6_n56), .Z(pe_1_5_6_n48) );
  MUX2_X1 pe_1_5_6_U92 ( .A(pe_1_5_6_int_q_reg_h[6]), .B(
        pe_1_5_6_int_q_reg_h[2]), .S(pe_1_5_6_n56), .Z(pe_1_5_6_n47) );
  MUX2_X1 pe_1_5_6_U91 ( .A(pe_1_5_6_n46), .B(pe_1_5_6_n24), .S(n52), .Z(
        int_data_x_5__6__1_) );
  MUX2_X1 pe_1_5_6_U90 ( .A(pe_1_5_6_n45), .B(pe_1_5_6_n25), .S(pe_1_5_6_n62), 
        .Z(pe_1_5_6_n46) );
  MUX2_X1 pe_1_5_6_U89 ( .A(pe_1_5_6_int_q_reg_h[21]), .B(
        pe_1_5_6_int_q_reg_h[17]), .S(pe_1_5_6_n56), .Z(pe_1_5_6_n45) );
  MUX2_X1 pe_1_5_6_U88 ( .A(pe_1_5_6_int_q_reg_h[13]), .B(
        pe_1_5_6_int_q_reg_h[9]), .S(pe_1_5_6_n56), .Z(pe_1_5_6_n25) );
  MUX2_X1 pe_1_5_6_U87 ( .A(pe_1_5_6_int_q_reg_h[5]), .B(
        pe_1_5_6_int_q_reg_h[1]), .S(pe_1_5_6_n56), .Z(pe_1_5_6_n24) );
  MUX2_X1 pe_1_5_6_U86 ( .A(pe_1_5_6_n23), .B(pe_1_5_6_n20), .S(n52), .Z(
        int_data_x_5__6__0_) );
  MUX2_X1 pe_1_5_6_U85 ( .A(pe_1_5_6_n22), .B(pe_1_5_6_n21), .S(pe_1_5_6_n62), 
        .Z(pe_1_5_6_n23) );
  MUX2_X1 pe_1_5_6_U84 ( .A(pe_1_5_6_int_q_reg_h[20]), .B(
        pe_1_5_6_int_q_reg_h[16]), .S(pe_1_5_6_n56), .Z(pe_1_5_6_n22) );
  MUX2_X1 pe_1_5_6_U83 ( .A(pe_1_5_6_int_q_reg_h[12]), .B(
        pe_1_5_6_int_q_reg_h[8]), .S(pe_1_5_6_n56), .Z(pe_1_5_6_n21) );
  MUX2_X1 pe_1_5_6_U82 ( .A(pe_1_5_6_int_q_reg_h[4]), .B(
        pe_1_5_6_int_q_reg_h[0]), .S(pe_1_5_6_n56), .Z(pe_1_5_6_n20) );
  MUX2_X1 pe_1_5_6_U81 ( .A(pe_1_5_6_n19), .B(pe_1_5_6_n16), .S(n52), .Z(
        int_data_y_5__6__3_) );
  MUX2_X1 pe_1_5_6_U80 ( .A(pe_1_5_6_n18), .B(pe_1_5_6_n17), .S(pe_1_5_6_n62), 
        .Z(pe_1_5_6_n19) );
  MUX2_X1 pe_1_5_6_U79 ( .A(pe_1_5_6_int_q_reg_v[23]), .B(
        pe_1_5_6_int_q_reg_v[19]), .S(pe_1_5_6_n55), .Z(pe_1_5_6_n18) );
  MUX2_X1 pe_1_5_6_U78 ( .A(pe_1_5_6_int_q_reg_v[15]), .B(
        pe_1_5_6_int_q_reg_v[11]), .S(pe_1_5_6_n55), .Z(pe_1_5_6_n17) );
  MUX2_X1 pe_1_5_6_U77 ( .A(pe_1_5_6_int_q_reg_v[7]), .B(
        pe_1_5_6_int_q_reg_v[3]), .S(pe_1_5_6_n55), .Z(pe_1_5_6_n16) );
  MUX2_X1 pe_1_5_6_U76 ( .A(pe_1_5_6_n15), .B(pe_1_5_6_n12), .S(n52), .Z(
        int_data_y_5__6__2_) );
  MUX2_X1 pe_1_5_6_U75 ( .A(pe_1_5_6_n14), .B(pe_1_5_6_n13), .S(pe_1_5_6_n62), 
        .Z(pe_1_5_6_n15) );
  MUX2_X1 pe_1_5_6_U74 ( .A(pe_1_5_6_int_q_reg_v[22]), .B(
        pe_1_5_6_int_q_reg_v[18]), .S(pe_1_5_6_n55), .Z(pe_1_5_6_n14) );
  MUX2_X1 pe_1_5_6_U73 ( .A(pe_1_5_6_int_q_reg_v[14]), .B(
        pe_1_5_6_int_q_reg_v[10]), .S(pe_1_5_6_n55), .Z(pe_1_5_6_n13) );
  MUX2_X1 pe_1_5_6_U72 ( .A(pe_1_5_6_int_q_reg_v[6]), .B(
        pe_1_5_6_int_q_reg_v[2]), .S(pe_1_5_6_n55), .Z(pe_1_5_6_n12) );
  MUX2_X1 pe_1_5_6_U71 ( .A(pe_1_5_6_n11), .B(pe_1_5_6_n8), .S(n52), .Z(
        int_data_y_5__6__1_) );
  MUX2_X1 pe_1_5_6_U70 ( .A(pe_1_5_6_n10), .B(pe_1_5_6_n9), .S(pe_1_5_6_n62), 
        .Z(pe_1_5_6_n11) );
  MUX2_X1 pe_1_5_6_U69 ( .A(pe_1_5_6_int_q_reg_v[21]), .B(
        pe_1_5_6_int_q_reg_v[17]), .S(pe_1_5_6_n55), .Z(pe_1_5_6_n10) );
  MUX2_X1 pe_1_5_6_U68 ( .A(pe_1_5_6_int_q_reg_v[13]), .B(
        pe_1_5_6_int_q_reg_v[9]), .S(pe_1_5_6_n55), .Z(pe_1_5_6_n9) );
  MUX2_X1 pe_1_5_6_U67 ( .A(pe_1_5_6_int_q_reg_v[5]), .B(
        pe_1_5_6_int_q_reg_v[1]), .S(pe_1_5_6_n55), .Z(pe_1_5_6_n8) );
  MUX2_X1 pe_1_5_6_U66 ( .A(pe_1_5_6_n7), .B(pe_1_5_6_n4), .S(n52), .Z(
        int_data_y_5__6__0_) );
  MUX2_X1 pe_1_5_6_U65 ( .A(pe_1_5_6_n6), .B(pe_1_5_6_n5), .S(pe_1_5_6_n62), 
        .Z(pe_1_5_6_n7) );
  MUX2_X1 pe_1_5_6_U64 ( .A(pe_1_5_6_int_q_reg_v[20]), .B(
        pe_1_5_6_int_q_reg_v[16]), .S(pe_1_5_6_n55), .Z(pe_1_5_6_n6) );
  MUX2_X1 pe_1_5_6_U63 ( .A(pe_1_5_6_int_q_reg_v[12]), .B(
        pe_1_5_6_int_q_reg_v[8]), .S(pe_1_5_6_n55), .Z(pe_1_5_6_n5) );
  MUX2_X1 pe_1_5_6_U62 ( .A(pe_1_5_6_int_q_reg_v[4]), .B(
        pe_1_5_6_int_q_reg_v[0]), .S(pe_1_5_6_n55), .Z(pe_1_5_6_n4) );
  AOI222_X1 pe_1_5_6_U61 ( .A1(int_data_res_6__6__2_), .A2(pe_1_5_6_n64), .B1(
        pe_1_5_6_N80), .B2(pe_1_5_6_n27), .C1(pe_1_5_6_N72), .C2(pe_1_5_6_n28), 
        .ZN(pe_1_5_6_n33) );
  INV_X1 pe_1_5_6_U60 ( .A(pe_1_5_6_n33), .ZN(pe_1_5_6_n82) );
  AOI222_X1 pe_1_5_6_U59 ( .A1(int_data_res_6__6__6_), .A2(pe_1_5_6_n64), .B1(
        pe_1_5_6_N84), .B2(pe_1_5_6_n27), .C1(pe_1_5_6_N76), .C2(pe_1_5_6_n28), 
        .ZN(pe_1_5_6_n29) );
  INV_X1 pe_1_5_6_U58 ( .A(pe_1_5_6_n29), .ZN(pe_1_5_6_n78) );
  XNOR2_X1 pe_1_5_6_U57 ( .A(pe_1_5_6_n73), .B(int_data_res_5__6__0_), .ZN(
        pe_1_5_6_N70) );
  AOI222_X1 pe_1_5_6_U52 ( .A1(int_data_res_6__6__0_), .A2(pe_1_5_6_n64), .B1(
        pe_1_5_6_n1), .B2(pe_1_5_6_n27), .C1(pe_1_5_6_N70), .C2(pe_1_5_6_n28), 
        .ZN(pe_1_5_6_n35) );
  INV_X1 pe_1_5_6_U51 ( .A(pe_1_5_6_n35), .ZN(pe_1_5_6_n84) );
  AOI222_X1 pe_1_5_6_U50 ( .A1(int_data_res_6__6__1_), .A2(pe_1_5_6_n64), .B1(
        pe_1_5_6_N79), .B2(pe_1_5_6_n27), .C1(pe_1_5_6_N71), .C2(pe_1_5_6_n28), 
        .ZN(pe_1_5_6_n34) );
  INV_X1 pe_1_5_6_U49 ( .A(pe_1_5_6_n34), .ZN(pe_1_5_6_n83) );
  AOI222_X1 pe_1_5_6_U48 ( .A1(int_data_res_6__6__3_), .A2(pe_1_5_6_n64), .B1(
        pe_1_5_6_N81), .B2(pe_1_5_6_n27), .C1(pe_1_5_6_N73), .C2(pe_1_5_6_n28), 
        .ZN(pe_1_5_6_n32) );
  INV_X1 pe_1_5_6_U47 ( .A(pe_1_5_6_n32), .ZN(pe_1_5_6_n81) );
  AOI222_X1 pe_1_5_6_U46 ( .A1(int_data_res_6__6__4_), .A2(pe_1_5_6_n64), .B1(
        pe_1_5_6_N82), .B2(pe_1_5_6_n27), .C1(pe_1_5_6_N74), .C2(pe_1_5_6_n28), 
        .ZN(pe_1_5_6_n31) );
  INV_X1 pe_1_5_6_U45 ( .A(pe_1_5_6_n31), .ZN(pe_1_5_6_n80) );
  AOI222_X1 pe_1_5_6_U44 ( .A1(int_data_res_6__6__5_), .A2(pe_1_5_6_n64), .B1(
        pe_1_5_6_N83), .B2(pe_1_5_6_n27), .C1(pe_1_5_6_N75), .C2(pe_1_5_6_n28), 
        .ZN(pe_1_5_6_n30) );
  INV_X1 pe_1_5_6_U43 ( .A(pe_1_5_6_n30), .ZN(pe_1_5_6_n79) );
  NAND2_X1 pe_1_5_6_U42 ( .A1(pe_1_5_6_int_data_0_), .A2(pe_1_5_6_n3), .ZN(
        pe_1_5_6_sub_81_carry[1]) );
  INV_X1 pe_1_5_6_U41 ( .A(pe_1_5_6_int_data_1_), .ZN(pe_1_5_6_n74) );
  INV_X1 pe_1_5_6_U40 ( .A(pe_1_5_6_int_data_2_), .ZN(pe_1_5_6_n75) );
  AND2_X1 pe_1_5_6_U39 ( .A1(pe_1_5_6_int_data_0_), .A2(int_data_res_5__6__0_), 
        .ZN(pe_1_5_6_n2) );
  AOI222_X1 pe_1_5_6_U38 ( .A1(pe_1_5_6_n64), .A2(int_data_res_6__6__7_), .B1(
        pe_1_5_6_N85), .B2(pe_1_5_6_n27), .C1(pe_1_5_6_N77), .C2(pe_1_5_6_n28), 
        .ZN(pe_1_5_6_n26) );
  INV_X1 pe_1_5_6_U37 ( .A(pe_1_5_6_n26), .ZN(pe_1_5_6_n77) );
  NOR3_X1 pe_1_5_6_U36 ( .A1(pe_1_5_6_n59), .A2(pe_1_5_6_n65), .A3(int_ckg[17]), .ZN(pe_1_5_6_n36) );
  OR2_X1 pe_1_5_6_U35 ( .A1(pe_1_5_6_n36), .A2(pe_1_5_6_n64), .ZN(pe_1_5_6_N90) );
  INV_X1 pe_1_5_6_U34 ( .A(n40), .ZN(pe_1_5_6_n63) );
  AND2_X1 pe_1_5_6_U33 ( .A1(int_data_x_5__6__2_), .A2(pe_1_5_6_n58), .ZN(
        pe_1_5_6_int_data_2_) );
  AND2_X1 pe_1_5_6_U32 ( .A1(int_data_x_5__6__1_), .A2(pe_1_5_6_n58), .ZN(
        pe_1_5_6_int_data_1_) );
  AND2_X1 pe_1_5_6_U31 ( .A1(int_data_x_5__6__3_), .A2(pe_1_5_6_n58), .ZN(
        pe_1_5_6_int_data_3_) );
  BUF_X1 pe_1_5_6_U30 ( .A(n62), .Z(pe_1_5_6_n64) );
  INV_X1 pe_1_5_6_U29 ( .A(n34), .ZN(pe_1_5_6_n61) );
  AND2_X1 pe_1_5_6_U28 ( .A1(int_data_x_5__6__0_), .A2(pe_1_5_6_n58), .ZN(
        pe_1_5_6_int_data_0_) );
  NAND2_X1 pe_1_5_6_U27 ( .A1(pe_1_5_6_n44), .A2(pe_1_5_6_n61), .ZN(
        pe_1_5_6_n41) );
  AND3_X1 pe_1_5_6_U26 ( .A1(n76), .A2(pe_1_5_6_n63), .A3(n52), .ZN(
        pe_1_5_6_n44) );
  INV_X1 pe_1_5_6_U25 ( .A(pe_1_5_6_int_data_3_), .ZN(pe_1_5_6_n76) );
  NOR2_X1 pe_1_5_6_U24 ( .A1(pe_1_5_6_n70), .A2(n52), .ZN(pe_1_5_6_n43) );
  NOR2_X1 pe_1_5_6_U23 ( .A1(pe_1_5_6_n57), .A2(pe_1_5_6_n64), .ZN(
        pe_1_5_6_n28) );
  NOR2_X1 pe_1_5_6_U22 ( .A1(n20), .A2(pe_1_5_6_n64), .ZN(pe_1_5_6_n27) );
  INV_X1 pe_1_5_6_U21 ( .A(pe_1_5_6_int_data_0_), .ZN(pe_1_5_6_n73) );
  INV_X1 pe_1_5_6_U20 ( .A(pe_1_5_6_n41), .ZN(pe_1_5_6_n90) );
  INV_X1 pe_1_5_6_U19 ( .A(pe_1_5_6_n37), .ZN(pe_1_5_6_n88) );
  INV_X1 pe_1_5_6_U18 ( .A(pe_1_5_6_n38), .ZN(pe_1_5_6_n87) );
  INV_X1 pe_1_5_6_U17 ( .A(pe_1_5_6_n39), .ZN(pe_1_5_6_n86) );
  NOR2_X1 pe_1_5_6_U16 ( .A1(pe_1_5_6_n68), .A2(pe_1_5_6_n42), .ZN(
        pe_1_5_6_N59) );
  NOR2_X1 pe_1_5_6_U15 ( .A1(pe_1_5_6_n68), .A2(pe_1_5_6_n41), .ZN(
        pe_1_5_6_N60) );
  NOR2_X1 pe_1_5_6_U14 ( .A1(pe_1_5_6_n68), .A2(pe_1_5_6_n38), .ZN(
        pe_1_5_6_N63) );
  NOR2_X1 pe_1_5_6_U13 ( .A1(pe_1_5_6_n67), .A2(pe_1_5_6_n40), .ZN(
        pe_1_5_6_N61) );
  NOR2_X1 pe_1_5_6_U12 ( .A1(pe_1_5_6_n67), .A2(pe_1_5_6_n39), .ZN(
        pe_1_5_6_N62) );
  NOR2_X1 pe_1_5_6_U11 ( .A1(pe_1_5_6_n37), .A2(pe_1_5_6_n67), .ZN(
        pe_1_5_6_N64) );
  NAND2_X1 pe_1_5_6_U10 ( .A1(pe_1_5_6_n44), .A2(pe_1_5_6_n60), .ZN(
        pe_1_5_6_n42) );
  BUF_X1 pe_1_5_6_U9 ( .A(pe_1_5_6_n60), .Z(pe_1_5_6_n55) );
  INV_X1 pe_1_5_6_U8 ( .A(pe_1_5_6_n69), .ZN(pe_1_5_6_n65) );
  BUF_X1 pe_1_5_6_U7 ( .A(pe_1_5_6_n60), .Z(pe_1_5_6_n56) );
  INV_X1 pe_1_5_6_U6 ( .A(pe_1_5_6_n42), .ZN(pe_1_5_6_n89) );
  INV_X1 pe_1_5_6_U5 ( .A(pe_1_5_6_n40), .ZN(pe_1_5_6_n85) );
  INV_X2 pe_1_5_6_U4 ( .A(n84), .ZN(pe_1_5_6_n72) );
  XOR2_X1 pe_1_5_6_U3 ( .A(pe_1_5_6_int_data_0_), .B(int_data_res_5__6__0_), 
        .Z(pe_1_5_6_n1) );
  DFFR_X1 pe_1_5_6_int_q_acc_reg_0_ ( .D(pe_1_5_6_n84), .CK(pe_1_5_6_net3964), 
        .RN(pe_1_5_6_n72), .Q(int_data_res_5__6__0_), .QN(pe_1_5_6_n3) );
  DFFR_X1 pe_1_5_6_int_q_reg_v_reg_0__0_ ( .D(int_data_y_6__6__0_), .CK(
        pe_1_5_6_net3934), .RN(pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_v[20]) );
  DFFR_X1 pe_1_5_6_int_q_reg_v_reg_0__1_ ( .D(int_data_y_6__6__1_), .CK(
        pe_1_5_6_net3934), .RN(pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_v[21]) );
  DFFR_X1 pe_1_5_6_int_q_reg_v_reg_0__2_ ( .D(int_data_y_6__6__2_), .CK(
        pe_1_5_6_net3934), .RN(pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_v[22]) );
  DFFR_X1 pe_1_5_6_int_q_reg_v_reg_0__3_ ( .D(int_data_y_6__6__3_), .CK(
        pe_1_5_6_net3934), .RN(pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_v[23]) );
  DFFR_X1 pe_1_5_6_int_q_reg_v_reg_1__0_ ( .D(int_data_y_6__6__0_), .CK(
        pe_1_5_6_net3939), .RN(pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_v[16]) );
  DFFR_X1 pe_1_5_6_int_q_reg_v_reg_1__1_ ( .D(int_data_y_6__6__1_), .CK(
        pe_1_5_6_net3939), .RN(pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_v[17]) );
  DFFR_X1 pe_1_5_6_int_q_reg_v_reg_1__2_ ( .D(int_data_y_6__6__2_), .CK(
        pe_1_5_6_net3939), .RN(pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_v[18]) );
  DFFR_X1 pe_1_5_6_int_q_reg_v_reg_1__3_ ( .D(int_data_y_6__6__3_), .CK(
        pe_1_5_6_net3939), .RN(pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_v[19]) );
  DFFR_X1 pe_1_5_6_int_q_reg_v_reg_2__0_ ( .D(int_data_y_6__6__0_), .CK(
        pe_1_5_6_net3944), .RN(pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_v[12]) );
  DFFR_X1 pe_1_5_6_int_q_reg_v_reg_2__1_ ( .D(int_data_y_6__6__1_), .CK(
        pe_1_5_6_net3944), .RN(pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_v[13]) );
  DFFR_X1 pe_1_5_6_int_q_reg_v_reg_2__2_ ( .D(int_data_y_6__6__2_), .CK(
        pe_1_5_6_net3944), .RN(pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_v[14]) );
  DFFR_X1 pe_1_5_6_int_q_reg_v_reg_2__3_ ( .D(int_data_y_6__6__3_), .CK(
        pe_1_5_6_net3944), .RN(pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_v[15]) );
  DFFR_X1 pe_1_5_6_int_q_reg_v_reg_3__0_ ( .D(int_data_y_6__6__0_), .CK(
        pe_1_5_6_net3949), .RN(pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_v[8]) );
  DFFR_X1 pe_1_5_6_int_q_reg_v_reg_3__1_ ( .D(int_data_y_6__6__1_), .CK(
        pe_1_5_6_net3949), .RN(pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_v[9]) );
  DFFR_X1 pe_1_5_6_int_q_reg_v_reg_3__2_ ( .D(int_data_y_6__6__2_), .CK(
        pe_1_5_6_net3949), .RN(pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_v[10]) );
  DFFR_X1 pe_1_5_6_int_q_reg_v_reg_3__3_ ( .D(int_data_y_6__6__3_), .CK(
        pe_1_5_6_net3949), .RN(pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_v[11]) );
  DFFR_X1 pe_1_5_6_int_q_reg_v_reg_4__0_ ( .D(int_data_y_6__6__0_), .CK(
        pe_1_5_6_net3954), .RN(pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_v[4]) );
  DFFR_X1 pe_1_5_6_int_q_reg_v_reg_4__1_ ( .D(int_data_y_6__6__1_), .CK(
        pe_1_5_6_net3954), .RN(pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_v[5]) );
  DFFR_X1 pe_1_5_6_int_q_reg_v_reg_4__2_ ( .D(int_data_y_6__6__2_), .CK(
        pe_1_5_6_net3954), .RN(pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_v[6]) );
  DFFR_X1 pe_1_5_6_int_q_reg_v_reg_4__3_ ( .D(int_data_y_6__6__3_), .CK(
        pe_1_5_6_net3954), .RN(pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_v[7]) );
  DFFR_X1 pe_1_5_6_int_q_reg_v_reg_5__0_ ( .D(int_data_y_6__6__0_), .CK(
        pe_1_5_6_net3959), .RN(pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_v[0]) );
  DFFR_X1 pe_1_5_6_int_q_reg_v_reg_5__1_ ( .D(int_data_y_6__6__1_), .CK(
        pe_1_5_6_net3959), .RN(pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_v[1]) );
  DFFR_X1 pe_1_5_6_int_q_reg_v_reg_5__2_ ( .D(int_data_y_6__6__2_), .CK(
        pe_1_5_6_net3959), .RN(pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_v[2]) );
  DFFR_X1 pe_1_5_6_int_q_reg_v_reg_5__3_ ( .D(int_data_y_6__6__3_), .CK(
        pe_1_5_6_net3959), .RN(pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_5_6_int_q_reg_h_reg_0__0_ ( .D(int_data_x_5__7__0_), .SI(
        int_data_y_6__6__0_), .SE(pe_1_5_6_n65), .CK(pe_1_5_6_net3903), .RN(
        pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_5_6_int_q_reg_h_reg_0__1_ ( .D(int_data_x_5__7__1_), .SI(
        int_data_y_6__6__1_), .SE(pe_1_5_6_n65), .CK(pe_1_5_6_net3903), .RN(
        pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_5_6_int_q_reg_h_reg_0__2_ ( .D(int_data_x_5__7__2_), .SI(
        int_data_y_6__6__2_), .SE(pe_1_5_6_n65), .CK(pe_1_5_6_net3903), .RN(
        pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_5_6_int_q_reg_h_reg_0__3_ ( .D(int_data_x_5__7__3_), .SI(
        int_data_y_6__6__3_), .SE(pe_1_5_6_n65), .CK(pe_1_5_6_net3903), .RN(
        pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_5_6_int_q_reg_h_reg_1__0_ ( .D(int_data_x_5__7__0_), .SI(
        int_data_y_6__6__0_), .SE(pe_1_5_6_n65), .CK(pe_1_5_6_net3909), .RN(
        pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_5_6_int_q_reg_h_reg_1__1_ ( .D(int_data_x_5__7__1_), .SI(
        int_data_y_6__6__1_), .SE(pe_1_5_6_n65), .CK(pe_1_5_6_net3909), .RN(
        pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_5_6_int_q_reg_h_reg_1__2_ ( .D(int_data_x_5__7__2_), .SI(
        int_data_y_6__6__2_), .SE(pe_1_5_6_n65), .CK(pe_1_5_6_net3909), .RN(
        pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_5_6_int_q_reg_h_reg_1__3_ ( .D(int_data_x_5__7__3_), .SI(
        int_data_y_6__6__3_), .SE(pe_1_5_6_n65), .CK(pe_1_5_6_net3909), .RN(
        pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_5_6_int_q_reg_h_reg_2__0_ ( .D(int_data_x_5__7__0_), .SI(
        int_data_y_6__6__0_), .SE(pe_1_5_6_n65), .CK(pe_1_5_6_net3914), .RN(
        pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_5_6_int_q_reg_h_reg_2__1_ ( .D(int_data_x_5__7__1_), .SI(
        int_data_y_6__6__1_), .SE(pe_1_5_6_n65), .CK(pe_1_5_6_net3914), .RN(
        pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_5_6_int_q_reg_h_reg_2__2_ ( .D(int_data_x_5__7__2_), .SI(
        int_data_y_6__6__2_), .SE(pe_1_5_6_n65), .CK(pe_1_5_6_net3914), .RN(
        pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_5_6_int_q_reg_h_reg_2__3_ ( .D(int_data_x_5__7__3_), .SI(
        int_data_y_6__6__3_), .SE(pe_1_5_6_n65), .CK(pe_1_5_6_net3914), .RN(
        pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_5_6_int_q_reg_h_reg_3__0_ ( .D(int_data_x_5__7__0_), .SI(
        int_data_y_6__6__0_), .SE(pe_1_5_6_n65), .CK(pe_1_5_6_net3919), .RN(
        pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_5_6_int_q_reg_h_reg_3__1_ ( .D(int_data_x_5__7__1_), .SI(
        int_data_y_6__6__1_), .SE(pe_1_5_6_n65), .CK(pe_1_5_6_net3919), .RN(
        pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_5_6_int_q_reg_h_reg_3__2_ ( .D(int_data_x_5__7__2_), .SI(
        int_data_y_6__6__2_), .SE(pe_1_5_6_n65), .CK(pe_1_5_6_net3919), .RN(
        pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_5_6_int_q_reg_h_reg_3__3_ ( .D(int_data_x_5__7__3_), .SI(
        int_data_y_6__6__3_), .SE(pe_1_5_6_n65), .CK(pe_1_5_6_net3919), .RN(
        pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_5_6_int_q_reg_h_reg_4__0_ ( .D(int_data_x_5__7__0_), .SI(
        int_data_y_6__6__0_), .SE(pe_1_5_6_n66), .CK(pe_1_5_6_net3924), .RN(
        pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_5_6_int_q_reg_h_reg_4__1_ ( .D(int_data_x_5__7__1_), .SI(
        int_data_y_6__6__1_), .SE(pe_1_5_6_n66), .CK(pe_1_5_6_net3924), .RN(
        pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_5_6_int_q_reg_h_reg_4__2_ ( .D(int_data_x_5__7__2_), .SI(
        int_data_y_6__6__2_), .SE(pe_1_5_6_n66), .CK(pe_1_5_6_net3924), .RN(
        pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_5_6_int_q_reg_h_reg_4__3_ ( .D(int_data_x_5__7__3_), .SI(
        int_data_y_6__6__3_), .SE(pe_1_5_6_n66), .CK(pe_1_5_6_net3924), .RN(
        pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_5_6_int_q_reg_h_reg_5__0_ ( .D(int_data_x_5__7__0_), .SI(
        int_data_y_6__6__0_), .SE(pe_1_5_6_n66), .CK(pe_1_5_6_net3929), .RN(
        pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_5_6_int_q_reg_h_reg_5__1_ ( .D(int_data_x_5__7__1_), .SI(
        int_data_y_6__6__1_), .SE(pe_1_5_6_n66), .CK(pe_1_5_6_net3929), .RN(
        pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_5_6_int_q_reg_h_reg_5__2_ ( .D(int_data_x_5__7__2_), .SI(
        int_data_y_6__6__2_), .SE(pe_1_5_6_n66), .CK(pe_1_5_6_net3929), .RN(
        pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_5_6_int_q_reg_h_reg_5__3_ ( .D(int_data_x_5__7__3_), .SI(
        int_data_y_6__6__3_), .SE(pe_1_5_6_n66), .CK(pe_1_5_6_net3929), .RN(
        pe_1_5_6_n72), .Q(pe_1_5_6_int_q_reg_h[3]) );
  FA_X1 pe_1_5_6_sub_81_U2_7 ( .A(int_data_res_5__6__7_), .B(pe_1_5_6_n76), 
        .CI(pe_1_5_6_sub_81_carry[7]), .S(pe_1_5_6_N77) );
  FA_X1 pe_1_5_6_sub_81_U2_6 ( .A(int_data_res_5__6__6_), .B(pe_1_5_6_n76), 
        .CI(pe_1_5_6_sub_81_carry[6]), .CO(pe_1_5_6_sub_81_carry[7]), .S(
        pe_1_5_6_N76) );
  FA_X1 pe_1_5_6_sub_81_U2_5 ( .A(int_data_res_5__6__5_), .B(pe_1_5_6_n76), 
        .CI(pe_1_5_6_sub_81_carry[5]), .CO(pe_1_5_6_sub_81_carry[6]), .S(
        pe_1_5_6_N75) );
  FA_X1 pe_1_5_6_sub_81_U2_4 ( .A(int_data_res_5__6__4_), .B(pe_1_5_6_n76), 
        .CI(pe_1_5_6_sub_81_carry[4]), .CO(pe_1_5_6_sub_81_carry[5]), .S(
        pe_1_5_6_N74) );
  FA_X1 pe_1_5_6_sub_81_U2_3 ( .A(int_data_res_5__6__3_), .B(pe_1_5_6_n76), 
        .CI(pe_1_5_6_sub_81_carry[3]), .CO(pe_1_5_6_sub_81_carry[4]), .S(
        pe_1_5_6_N73) );
  FA_X1 pe_1_5_6_sub_81_U2_2 ( .A(int_data_res_5__6__2_), .B(pe_1_5_6_n75), 
        .CI(pe_1_5_6_sub_81_carry[2]), .CO(pe_1_5_6_sub_81_carry[3]), .S(
        pe_1_5_6_N72) );
  FA_X1 pe_1_5_6_sub_81_U2_1 ( .A(int_data_res_5__6__1_), .B(pe_1_5_6_n74), 
        .CI(pe_1_5_6_sub_81_carry[1]), .CO(pe_1_5_6_sub_81_carry[2]), .S(
        pe_1_5_6_N71) );
  FA_X1 pe_1_5_6_add_83_U1_7 ( .A(int_data_res_5__6__7_), .B(
        pe_1_5_6_int_data_3_), .CI(pe_1_5_6_add_83_carry[7]), .S(pe_1_5_6_N85)
         );
  FA_X1 pe_1_5_6_add_83_U1_6 ( .A(int_data_res_5__6__6_), .B(
        pe_1_5_6_int_data_3_), .CI(pe_1_5_6_add_83_carry[6]), .CO(
        pe_1_5_6_add_83_carry[7]), .S(pe_1_5_6_N84) );
  FA_X1 pe_1_5_6_add_83_U1_5 ( .A(int_data_res_5__6__5_), .B(
        pe_1_5_6_int_data_3_), .CI(pe_1_5_6_add_83_carry[5]), .CO(
        pe_1_5_6_add_83_carry[6]), .S(pe_1_5_6_N83) );
  FA_X1 pe_1_5_6_add_83_U1_4 ( .A(int_data_res_5__6__4_), .B(
        pe_1_5_6_int_data_3_), .CI(pe_1_5_6_add_83_carry[4]), .CO(
        pe_1_5_6_add_83_carry[5]), .S(pe_1_5_6_N82) );
  FA_X1 pe_1_5_6_add_83_U1_3 ( .A(int_data_res_5__6__3_), .B(
        pe_1_5_6_int_data_3_), .CI(pe_1_5_6_add_83_carry[3]), .CO(
        pe_1_5_6_add_83_carry[4]), .S(pe_1_5_6_N81) );
  FA_X1 pe_1_5_6_add_83_U1_2 ( .A(int_data_res_5__6__2_), .B(
        pe_1_5_6_int_data_2_), .CI(pe_1_5_6_add_83_carry[2]), .CO(
        pe_1_5_6_add_83_carry[3]), .S(pe_1_5_6_N80) );
  FA_X1 pe_1_5_6_add_83_U1_1 ( .A(int_data_res_5__6__1_), .B(
        pe_1_5_6_int_data_1_), .CI(pe_1_5_6_n2), .CO(pe_1_5_6_add_83_carry[2]), 
        .S(pe_1_5_6_N79) );
  NAND3_X1 pe_1_5_6_U56 ( .A1(pe_1_5_6_n60), .A2(pe_1_5_6_n43), .A3(
        pe_1_5_6_n62), .ZN(pe_1_5_6_n40) );
  NAND3_X1 pe_1_5_6_U55 ( .A1(pe_1_5_6_n43), .A2(pe_1_5_6_n61), .A3(
        pe_1_5_6_n62), .ZN(pe_1_5_6_n39) );
  NAND3_X1 pe_1_5_6_U54 ( .A1(pe_1_5_6_n43), .A2(pe_1_5_6_n63), .A3(
        pe_1_5_6_n60), .ZN(pe_1_5_6_n38) );
  NAND3_X1 pe_1_5_6_U53 ( .A1(pe_1_5_6_n61), .A2(pe_1_5_6_n63), .A3(
        pe_1_5_6_n43), .ZN(pe_1_5_6_n37) );
  DFFR_X1 pe_1_5_6_int_q_acc_reg_6_ ( .D(pe_1_5_6_n78), .CK(pe_1_5_6_net3964), 
        .RN(pe_1_5_6_n71), .Q(int_data_res_5__6__6_) );
  DFFR_X1 pe_1_5_6_int_q_acc_reg_5_ ( .D(pe_1_5_6_n79), .CK(pe_1_5_6_net3964), 
        .RN(pe_1_5_6_n71), .Q(int_data_res_5__6__5_) );
  DFFR_X1 pe_1_5_6_int_q_acc_reg_4_ ( .D(pe_1_5_6_n80), .CK(pe_1_5_6_net3964), 
        .RN(pe_1_5_6_n71), .Q(int_data_res_5__6__4_) );
  DFFR_X1 pe_1_5_6_int_q_acc_reg_3_ ( .D(pe_1_5_6_n81), .CK(pe_1_5_6_net3964), 
        .RN(pe_1_5_6_n71), .Q(int_data_res_5__6__3_) );
  DFFR_X1 pe_1_5_6_int_q_acc_reg_2_ ( .D(pe_1_5_6_n82), .CK(pe_1_5_6_net3964), 
        .RN(pe_1_5_6_n71), .Q(int_data_res_5__6__2_) );
  DFFR_X1 pe_1_5_6_int_q_acc_reg_1_ ( .D(pe_1_5_6_n83), .CK(pe_1_5_6_net3964), 
        .RN(pe_1_5_6_n71), .Q(int_data_res_5__6__1_) );
  DFFR_X1 pe_1_5_6_int_q_acc_reg_7_ ( .D(pe_1_5_6_n77), .CK(pe_1_5_6_net3964), 
        .RN(pe_1_5_6_n71), .Q(int_data_res_5__6__7_) );
  CLKGATETST_X1 pe_1_5_6_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_5_6_n88), .SE(1'b0), .GCK(pe_1_5_6_net3903) );
  CLKGATETST_X1 pe_1_5_6_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_5_6_n87), .SE(1'b0), .GCK(pe_1_5_6_net3909) );
  CLKGATETST_X1 pe_1_5_6_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_5_6_n86), .SE(1'b0), .GCK(pe_1_5_6_net3914) );
  CLKGATETST_X1 pe_1_5_6_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_5_6_n85), .SE(1'b0), .GCK(pe_1_5_6_net3919) );
  CLKGATETST_X1 pe_1_5_6_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_5_6_n90), .SE(1'b0), .GCK(pe_1_5_6_net3924) );
  CLKGATETST_X1 pe_1_5_6_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_5_6_n89), .SE(1'b0), .GCK(pe_1_5_6_net3929) );
  CLKGATETST_X1 pe_1_5_6_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_5_6_N64), .SE(1'b0), .GCK(pe_1_5_6_net3934) );
  CLKGATETST_X1 pe_1_5_6_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_5_6_N63), .SE(1'b0), .GCK(pe_1_5_6_net3939) );
  CLKGATETST_X1 pe_1_5_6_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_5_6_N62), .SE(1'b0), .GCK(pe_1_5_6_net3944) );
  CLKGATETST_X1 pe_1_5_6_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_5_6_N61), .SE(1'b0), .GCK(pe_1_5_6_net3949) );
  CLKGATETST_X1 pe_1_5_6_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_5_6_N60), .SE(1'b0), .GCK(pe_1_5_6_net3954) );
  CLKGATETST_X1 pe_1_5_6_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_5_6_N59), .SE(1'b0), .GCK(pe_1_5_6_net3959) );
  CLKGATETST_X1 pe_1_5_6_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_5_6_N90), .SE(1'b0), .GCK(pe_1_5_6_net3964) );
  CLKBUF_X1 pe_1_5_7_U112 ( .A(pe_1_5_7_n72), .Z(pe_1_5_7_n71) );
  INV_X1 pe_1_5_7_U111 ( .A(n76), .ZN(pe_1_5_7_n70) );
  INV_X1 pe_1_5_7_U110 ( .A(n68), .ZN(pe_1_5_7_n69) );
  INV_X1 pe_1_5_7_U109 ( .A(n68), .ZN(pe_1_5_7_n68) );
  INV_X1 pe_1_5_7_U108 ( .A(n68), .ZN(pe_1_5_7_n67) );
  INV_X1 pe_1_5_7_U107 ( .A(pe_1_5_7_n69), .ZN(pe_1_5_7_n66) );
  INV_X1 pe_1_5_7_U106 ( .A(pe_1_5_7_n63), .ZN(pe_1_5_7_n62) );
  INV_X1 pe_1_5_7_U105 ( .A(pe_1_5_7_n61), .ZN(pe_1_5_7_n60) );
  INV_X1 pe_1_5_7_U104 ( .A(n28), .ZN(pe_1_5_7_n59) );
  INV_X1 pe_1_5_7_U103 ( .A(pe_1_5_7_n59), .ZN(pe_1_5_7_n58) );
  INV_X1 pe_1_5_7_U102 ( .A(n20), .ZN(pe_1_5_7_n57) );
  MUX2_X1 pe_1_5_7_U101 ( .A(pe_1_5_7_n54), .B(pe_1_5_7_n51), .S(n52), .Z(
        int_data_x_5__7__3_) );
  MUX2_X1 pe_1_5_7_U100 ( .A(pe_1_5_7_n53), .B(pe_1_5_7_n52), .S(pe_1_5_7_n62), 
        .Z(pe_1_5_7_n54) );
  MUX2_X1 pe_1_5_7_U99 ( .A(pe_1_5_7_int_q_reg_h[23]), .B(
        pe_1_5_7_int_q_reg_h[19]), .S(pe_1_5_7_n56), .Z(pe_1_5_7_n53) );
  MUX2_X1 pe_1_5_7_U98 ( .A(pe_1_5_7_int_q_reg_h[15]), .B(
        pe_1_5_7_int_q_reg_h[11]), .S(pe_1_5_7_n56), .Z(pe_1_5_7_n52) );
  MUX2_X1 pe_1_5_7_U97 ( .A(pe_1_5_7_int_q_reg_h[7]), .B(
        pe_1_5_7_int_q_reg_h[3]), .S(pe_1_5_7_n56), .Z(pe_1_5_7_n51) );
  MUX2_X1 pe_1_5_7_U96 ( .A(pe_1_5_7_n50), .B(pe_1_5_7_n47), .S(n52), .Z(
        int_data_x_5__7__2_) );
  MUX2_X1 pe_1_5_7_U95 ( .A(pe_1_5_7_n49), .B(pe_1_5_7_n48), .S(pe_1_5_7_n62), 
        .Z(pe_1_5_7_n50) );
  MUX2_X1 pe_1_5_7_U94 ( .A(pe_1_5_7_int_q_reg_h[22]), .B(
        pe_1_5_7_int_q_reg_h[18]), .S(pe_1_5_7_n56), .Z(pe_1_5_7_n49) );
  MUX2_X1 pe_1_5_7_U93 ( .A(pe_1_5_7_int_q_reg_h[14]), .B(
        pe_1_5_7_int_q_reg_h[10]), .S(pe_1_5_7_n56), .Z(pe_1_5_7_n48) );
  MUX2_X1 pe_1_5_7_U92 ( .A(pe_1_5_7_int_q_reg_h[6]), .B(
        pe_1_5_7_int_q_reg_h[2]), .S(pe_1_5_7_n56), .Z(pe_1_5_7_n47) );
  MUX2_X1 pe_1_5_7_U91 ( .A(pe_1_5_7_n46), .B(pe_1_5_7_n24), .S(n52), .Z(
        int_data_x_5__7__1_) );
  MUX2_X1 pe_1_5_7_U90 ( .A(pe_1_5_7_n45), .B(pe_1_5_7_n25), .S(pe_1_5_7_n62), 
        .Z(pe_1_5_7_n46) );
  MUX2_X1 pe_1_5_7_U89 ( .A(pe_1_5_7_int_q_reg_h[21]), .B(
        pe_1_5_7_int_q_reg_h[17]), .S(pe_1_5_7_n56), .Z(pe_1_5_7_n45) );
  MUX2_X1 pe_1_5_7_U88 ( .A(pe_1_5_7_int_q_reg_h[13]), .B(
        pe_1_5_7_int_q_reg_h[9]), .S(pe_1_5_7_n56), .Z(pe_1_5_7_n25) );
  MUX2_X1 pe_1_5_7_U87 ( .A(pe_1_5_7_int_q_reg_h[5]), .B(
        pe_1_5_7_int_q_reg_h[1]), .S(pe_1_5_7_n56), .Z(pe_1_5_7_n24) );
  MUX2_X1 pe_1_5_7_U86 ( .A(pe_1_5_7_n23), .B(pe_1_5_7_n20), .S(n52), .Z(
        int_data_x_5__7__0_) );
  MUX2_X1 pe_1_5_7_U85 ( .A(pe_1_5_7_n22), .B(pe_1_5_7_n21), .S(pe_1_5_7_n62), 
        .Z(pe_1_5_7_n23) );
  MUX2_X1 pe_1_5_7_U84 ( .A(pe_1_5_7_int_q_reg_h[20]), .B(
        pe_1_5_7_int_q_reg_h[16]), .S(pe_1_5_7_n56), .Z(pe_1_5_7_n22) );
  MUX2_X1 pe_1_5_7_U83 ( .A(pe_1_5_7_int_q_reg_h[12]), .B(
        pe_1_5_7_int_q_reg_h[8]), .S(pe_1_5_7_n56), .Z(pe_1_5_7_n21) );
  MUX2_X1 pe_1_5_7_U82 ( .A(pe_1_5_7_int_q_reg_h[4]), .B(
        pe_1_5_7_int_q_reg_h[0]), .S(pe_1_5_7_n56), .Z(pe_1_5_7_n20) );
  MUX2_X1 pe_1_5_7_U81 ( .A(pe_1_5_7_n19), .B(pe_1_5_7_n16), .S(n52), .Z(
        int_data_y_5__7__3_) );
  MUX2_X1 pe_1_5_7_U80 ( .A(pe_1_5_7_n18), .B(pe_1_5_7_n17), .S(pe_1_5_7_n62), 
        .Z(pe_1_5_7_n19) );
  MUX2_X1 pe_1_5_7_U79 ( .A(pe_1_5_7_int_q_reg_v[23]), .B(
        pe_1_5_7_int_q_reg_v[19]), .S(pe_1_5_7_n55), .Z(pe_1_5_7_n18) );
  MUX2_X1 pe_1_5_7_U78 ( .A(pe_1_5_7_int_q_reg_v[15]), .B(
        pe_1_5_7_int_q_reg_v[11]), .S(pe_1_5_7_n55), .Z(pe_1_5_7_n17) );
  MUX2_X1 pe_1_5_7_U77 ( .A(pe_1_5_7_int_q_reg_v[7]), .B(
        pe_1_5_7_int_q_reg_v[3]), .S(pe_1_5_7_n55), .Z(pe_1_5_7_n16) );
  MUX2_X1 pe_1_5_7_U76 ( .A(pe_1_5_7_n15), .B(pe_1_5_7_n12), .S(n52), .Z(
        int_data_y_5__7__2_) );
  MUX2_X1 pe_1_5_7_U75 ( .A(pe_1_5_7_n14), .B(pe_1_5_7_n13), .S(pe_1_5_7_n62), 
        .Z(pe_1_5_7_n15) );
  MUX2_X1 pe_1_5_7_U74 ( .A(pe_1_5_7_int_q_reg_v[22]), .B(
        pe_1_5_7_int_q_reg_v[18]), .S(pe_1_5_7_n55), .Z(pe_1_5_7_n14) );
  MUX2_X1 pe_1_5_7_U73 ( .A(pe_1_5_7_int_q_reg_v[14]), .B(
        pe_1_5_7_int_q_reg_v[10]), .S(pe_1_5_7_n55), .Z(pe_1_5_7_n13) );
  MUX2_X1 pe_1_5_7_U72 ( .A(pe_1_5_7_int_q_reg_v[6]), .B(
        pe_1_5_7_int_q_reg_v[2]), .S(pe_1_5_7_n55), .Z(pe_1_5_7_n12) );
  MUX2_X1 pe_1_5_7_U71 ( .A(pe_1_5_7_n11), .B(pe_1_5_7_n8), .S(n52), .Z(
        int_data_y_5__7__1_) );
  MUX2_X1 pe_1_5_7_U70 ( .A(pe_1_5_7_n10), .B(pe_1_5_7_n9), .S(pe_1_5_7_n62), 
        .Z(pe_1_5_7_n11) );
  MUX2_X1 pe_1_5_7_U69 ( .A(pe_1_5_7_int_q_reg_v[21]), .B(
        pe_1_5_7_int_q_reg_v[17]), .S(pe_1_5_7_n55), .Z(pe_1_5_7_n10) );
  MUX2_X1 pe_1_5_7_U68 ( .A(pe_1_5_7_int_q_reg_v[13]), .B(
        pe_1_5_7_int_q_reg_v[9]), .S(pe_1_5_7_n55), .Z(pe_1_5_7_n9) );
  MUX2_X1 pe_1_5_7_U67 ( .A(pe_1_5_7_int_q_reg_v[5]), .B(
        pe_1_5_7_int_q_reg_v[1]), .S(pe_1_5_7_n55), .Z(pe_1_5_7_n8) );
  MUX2_X1 pe_1_5_7_U66 ( .A(pe_1_5_7_n7), .B(pe_1_5_7_n4), .S(n52), .Z(
        int_data_y_5__7__0_) );
  MUX2_X1 pe_1_5_7_U65 ( .A(pe_1_5_7_n6), .B(pe_1_5_7_n5), .S(pe_1_5_7_n62), 
        .Z(pe_1_5_7_n7) );
  MUX2_X1 pe_1_5_7_U64 ( .A(pe_1_5_7_int_q_reg_v[20]), .B(
        pe_1_5_7_int_q_reg_v[16]), .S(pe_1_5_7_n55), .Z(pe_1_5_7_n6) );
  MUX2_X1 pe_1_5_7_U63 ( .A(pe_1_5_7_int_q_reg_v[12]), .B(
        pe_1_5_7_int_q_reg_v[8]), .S(pe_1_5_7_n55), .Z(pe_1_5_7_n5) );
  MUX2_X1 pe_1_5_7_U62 ( .A(pe_1_5_7_int_q_reg_v[4]), .B(
        pe_1_5_7_int_q_reg_v[0]), .S(pe_1_5_7_n55), .Z(pe_1_5_7_n4) );
  AOI222_X1 pe_1_5_7_U61 ( .A1(int_data_res_6__7__2_), .A2(pe_1_5_7_n64), .B1(
        pe_1_5_7_N80), .B2(pe_1_5_7_n27), .C1(pe_1_5_7_N72), .C2(pe_1_5_7_n28), 
        .ZN(pe_1_5_7_n33) );
  INV_X1 pe_1_5_7_U60 ( .A(pe_1_5_7_n33), .ZN(pe_1_5_7_n82) );
  AOI222_X1 pe_1_5_7_U59 ( .A1(int_data_res_6__7__6_), .A2(pe_1_5_7_n64), .B1(
        pe_1_5_7_N84), .B2(pe_1_5_7_n27), .C1(pe_1_5_7_N76), .C2(pe_1_5_7_n28), 
        .ZN(pe_1_5_7_n29) );
  INV_X1 pe_1_5_7_U58 ( .A(pe_1_5_7_n29), .ZN(pe_1_5_7_n78) );
  XNOR2_X1 pe_1_5_7_U57 ( .A(pe_1_5_7_n73), .B(int_data_res_5__7__0_), .ZN(
        pe_1_5_7_N70) );
  AOI222_X1 pe_1_5_7_U52 ( .A1(int_data_res_6__7__0_), .A2(pe_1_5_7_n64), .B1(
        pe_1_5_7_n1), .B2(pe_1_5_7_n27), .C1(pe_1_5_7_N70), .C2(pe_1_5_7_n28), 
        .ZN(pe_1_5_7_n35) );
  INV_X1 pe_1_5_7_U51 ( .A(pe_1_5_7_n35), .ZN(pe_1_5_7_n84) );
  AOI222_X1 pe_1_5_7_U50 ( .A1(int_data_res_6__7__1_), .A2(pe_1_5_7_n64), .B1(
        pe_1_5_7_N79), .B2(pe_1_5_7_n27), .C1(pe_1_5_7_N71), .C2(pe_1_5_7_n28), 
        .ZN(pe_1_5_7_n34) );
  INV_X1 pe_1_5_7_U49 ( .A(pe_1_5_7_n34), .ZN(pe_1_5_7_n83) );
  AOI222_X1 pe_1_5_7_U48 ( .A1(int_data_res_6__7__3_), .A2(pe_1_5_7_n64), .B1(
        pe_1_5_7_N81), .B2(pe_1_5_7_n27), .C1(pe_1_5_7_N73), .C2(pe_1_5_7_n28), 
        .ZN(pe_1_5_7_n32) );
  INV_X1 pe_1_5_7_U47 ( .A(pe_1_5_7_n32), .ZN(pe_1_5_7_n81) );
  AOI222_X1 pe_1_5_7_U46 ( .A1(int_data_res_6__7__4_), .A2(pe_1_5_7_n64), .B1(
        pe_1_5_7_N82), .B2(pe_1_5_7_n27), .C1(pe_1_5_7_N74), .C2(pe_1_5_7_n28), 
        .ZN(pe_1_5_7_n31) );
  INV_X1 pe_1_5_7_U45 ( .A(pe_1_5_7_n31), .ZN(pe_1_5_7_n80) );
  AOI222_X1 pe_1_5_7_U44 ( .A1(int_data_res_6__7__5_), .A2(pe_1_5_7_n64), .B1(
        pe_1_5_7_N83), .B2(pe_1_5_7_n27), .C1(pe_1_5_7_N75), .C2(pe_1_5_7_n28), 
        .ZN(pe_1_5_7_n30) );
  INV_X1 pe_1_5_7_U43 ( .A(pe_1_5_7_n30), .ZN(pe_1_5_7_n79) );
  NAND2_X1 pe_1_5_7_U42 ( .A1(pe_1_5_7_int_data_0_), .A2(pe_1_5_7_n3), .ZN(
        pe_1_5_7_sub_81_carry[1]) );
  INV_X1 pe_1_5_7_U41 ( .A(pe_1_5_7_int_data_1_), .ZN(pe_1_5_7_n74) );
  INV_X1 pe_1_5_7_U40 ( .A(pe_1_5_7_int_data_2_), .ZN(pe_1_5_7_n75) );
  AND2_X1 pe_1_5_7_U39 ( .A1(pe_1_5_7_int_data_0_), .A2(int_data_res_5__7__0_), 
        .ZN(pe_1_5_7_n2) );
  AOI222_X1 pe_1_5_7_U38 ( .A1(pe_1_5_7_n64), .A2(int_data_res_6__7__7_), .B1(
        pe_1_5_7_N85), .B2(pe_1_5_7_n27), .C1(pe_1_5_7_N77), .C2(pe_1_5_7_n28), 
        .ZN(pe_1_5_7_n26) );
  INV_X1 pe_1_5_7_U37 ( .A(pe_1_5_7_n26), .ZN(pe_1_5_7_n77) );
  NOR3_X1 pe_1_5_7_U36 ( .A1(pe_1_5_7_n59), .A2(pe_1_5_7_n65), .A3(int_ckg[16]), .ZN(pe_1_5_7_n36) );
  OR2_X1 pe_1_5_7_U35 ( .A1(pe_1_5_7_n36), .A2(pe_1_5_7_n64), .ZN(pe_1_5_7_N90) );
  INV_X1 pe_1_5_7_U34 ( .A(n40), .ZN(pe_1_5_7_n63) );
  AND2_X1 pe_1_5_7_U33 ( .A1(int_data_x_5__7__2_), .A2(pe_1_5_7_n58), .ZN(
        pe_1_5_7_int_data_2_) );
  AND2_X1 pe_1_5_7_U32 ( .A1(int_data_x_5__7__1_), .A2(pe_1_5_7_n58), .ZN(
        pe_1_5_7_int_data_1_) );
  AND2_X1 pe_1_5_7_U31 ( .A1(int_data_x_5__7__3_), .A2(pe_1_5_7_n58), .ZN(
        pe_1_5_7_int_data_3_) );
  BUF_X1 pe_1_5_7_U30 ( .A(n62), .Z(pe_1_5_7_n64) );
  INV_X1 pe_1_5_7_U29 ( .A(n34), .ZN(pe_1_5_7_n61) );
  AND2_X1 pe_1_5_7_U28 ( .A1(int_data_x_5__7__0_), .A2(pe_1_5_7_n58), .ZN(
        pe_1_5_7_int_data_0_) );
  NAND2_X1 pe_1_5_7_U27 ( .A1(pe_1_5_7_n44), .A2(pe_1_5_7_n61), .ZN(
        pe_1_5_7_n41) );
  AND3_X1 pe_1_5_7_U26 ( .A1(n76), .A2(pe_1_5_7_n63), .A3(n52), .ZN(
        pe_1_5_7_n44) );
  INV_X1 pe_1_5_7_U25 ( .A(pe_1_5_7_int_data_3_), .ZN(pe_1_5_7_n76) );
  NOR2_X1 pe_1_5_7_U24 ( .A1(pe_1_5_7_n70), .A2(n52), .ZN(pe_1_5_7_n43) );
  NOR2_X1 pe_1_5_7_U23 ( .A1(pe_1_5_7_n57), .A2(pe_1_5_7_n64), .ZN(
        pe_1_5_7_n28) );
  NOR2_X1 pe_1_5_7_U22 ( .A1(n20), .A2(pe_1_5_7_n64), .ZN(pe_1_5_7_n27) );
  INV_X1 pe_1_5_7_U21 ( .A(pe_1_5_7_int_data_0_), .ZN(pe_1_5_7_n73) );
  INV_X1 pe_1_5_7_U20 ( .A(pe_1_5_7_n41), .ZN(pe_1_5_7_n90) );
  INV_X1 pe_1_5_7_U19 ( .A(pe_1_5_7_n37), .ZN(pe_1_5_7_n88) );
  INV_X1 pe_1_5_7_U18 ( .A(pe_1_5_7_n38), .ZN(pe_1_5_7_n87) );
  INV_X1 pe_1_5_7_U17 ( .A(pe_1_5_7_n39), .ZN(pe_1_5_7_n86) );
  NOR2_X1 pe_1_5_7_U16 ( .A1(pe_1_5_7_n68), .A2(pe_1_5_7_n42), .ZN(
        pe_1_5_7_N59) );
  NOR2_X1 pe_1_5_7_U15 ( .A1(pe_1_5_7_n68), .A2(pe_1_5_7_n41), .ZN(
        pe_1_5_7_N60) );
  NOR2_X1 pe_1_5_7_U14 ( .A1(pe_1_5_7_n68), .A2(pe_1_5_7_n38), .ZN(
        pe_1_5_7_N63) );
  NOR2_X1 pe_1_5_7_U13 ( .A1(pe_1_5_7_n67), .A2(pe_1_5_7_n40), .ZN(
        pe_1_5_7_N61) );
  NOR2_X1 pe_1_5_7_U12 ( .A1(pe_1_5_7_n67), .A2(pe_1_5_7_n39), .ZN(
        pe_1_5_7_N62) );
  NOR2_X1 pe_1_5_7_U11 ( .A1(pe_1_5_7_n37), .A2(pe_1_5_7_n67), .ZN(
        pe_1_5_7_N64) );
  NAND2_X1 pe_1_5_7_U10 ( .A1(pe_1_5_7_n44), .A2(pe_1_5_7_n60), .ZN(
        pe_1_5_7_n42) );
  BUF_X1 pe_1_5_7_U9 ( .A(pe_1_5_7_n60), .Z(pe_1_5_7_n55) );
  INV_X1 pe_1_5_7_U8 ( .A(pe_1_5_7_n69), .ZN(pe_1_5_7_n65) );
  BUF_X1 pe_1_5_7_U7 ( .A(pe_1_5_7_n60), .Z(pe_1_5_7_n56) );
  INV_X1 pe_1_5_7_U6 ( .A(pe_1_5_7_n42), .ZN(pe_1_5_7_n89) );
  INV_X1 pe_1_5_7_U5 ( .A(pe_1_5_7_n40), .ZN(pe_1_5_7_n85) );
  INV_X2 pe_1_5_7_U4 ( .A(n84), .ZN(pe_1_5_7_n72) );
  XOR2_X1 pe_1_5_7_U3 ( .A(pe_1_5_7_int_data_0_), .B(int_data_res_5__7__0_), 
        .Z(pe_1_5_7_n1) );
  DFFR_X1 pe_1_5_7_int_q_acc_reg_0_ ( .D(pe_1_5_7_n84), .CK(pe_1_5_7_net3886), 
        .RN(pe_1_5_7_n72), .Q(int_data_res_5__7__0_), .QN(pe_1_5_7_n3) );
  DFFR_X1 pe_1_5_7_int_q_reg_v_reg_0__0_ ( .D(int_data_y_6__7__0_), .CK(
        pe_1_5_7_net3856), .RN(pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_v[20]) );
  DFFR_X1 pe_1_5_7_int_q_reg_v_reg_0__1_ ( .D(int_data_y_6__7__1_), .CK(
        pe_1_5_7_net3856), .RN(pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_v[21]) );
  DFFR_X1 pe_1_5_7_int_q_reg_v_reg_0__2_ ( .D(int_data_y_6__7__2_), .CK(
        pe_1_5_7_net3856), .RN(pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_v[22]) );
  DFFR_X1 pe_1_5_7_int_q_reg_v_reg_0__3_ ( .D(int_data_y_6__7__3_), .CK(
        pe_1_5_7_net3856), .RN(pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_v[23]) );
  DFFR_X1 pe_1_5_7_int_q_reg_v_reg_1__0_ ( .D(int_data_y_6__7__0_), .CK(
        pe_1_5_7_net3861), .RN(pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_v[16]) );
  DFFR_X1 pe_1_5_7_int_q_reg_v_reg_1__1_ ( .D(int_data_y_6__7__1_), .CK(
        pe_1_5_7_net3861), .RN(pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_v[17]) );
  DFFR_X1 pe_1_5_7_int_q_reg_v_reg_1__2_ ( .D(int_data_y_6__7__2_), .CK(
        pe_1_5_7_net3861), .RN(pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_v[18]) );
  DFFR_X1 pe_1_5_7_int_q_reg_v_reg_1__3_ ( .D(int_data_y_6__7__3_), .CK(
        pe_1_5_7_net3861), .RN(pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_v[19]) );
  DFFR_X1 pe_1_5_7_int_q_reg_v_reg_2__0_ ( .D(int_data_y_6__7__0_), .CK(
        pe_1_5_7_net3866), .RN(pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_v[12]) );
  DFFR_X1 pe_1_5_7_int_q_reg_v_reg_2__1_ ( .D(int_data_y_6__7__1_), .CK(
        pe_1_5_7_net3866), .RN(pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_v[13]) );
  DFFR_X1 pe_1_5_7_int_q_reg_v_reg_2__2_ ( .D(int_data_y_6__7__2_), .CK(
        pe_1_5_7_net3866), .RN(pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_v[14]) );
  DFFR_X1 pe_1_5_7_int_q_reg_v_reg_2__3_ ( .D(int_data_y_6__7__3_), .CK(
        pe_1_5_7_net3866), .RN(pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_v[15]) );
  DFFR_X1 pe_1_5_7_int_q_reg_v_reg_3__0_ ( .D(int_data_y_6__7__0_), .CK(
        pe_1_5_7_net3871), .RN(pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_v[8]) );
  DFFR_X1 pe_1_5_7_int_q_reg_v_reg_3__1_ ( .D(int_data_y_6__7__1_), .CK(
        pe_1_5_7_net3871), .RN(pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_v[9]) );
  DFFR_X1 pe_1_5_7_int_q_reg_v_reg_3__2_ ( .D(int_data_y_6__7__2_), .CK(
        pe_1_5_7_net3871), .RN(pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_v[10]) );
  DFFR_X1 pe_1_5_7_int_q_reg_v_reg_3__3_ ( .D(int_data_y_6__7__3_), .CK(
        pe_1_5_7_net3871), .RN(pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_v[11]) );
  DFFR_X1 pe_1_5_7_int_q_reg_v_reg_4__0_ ( .D(int_data_y_6__7__0_), .CK(
        pe_1_5_7_net3876), .RN(pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_v[4]) );
  DFFR_X1 pe_1_5_7_int_q_reg_v_reg_4__1_ ( .D(int_data_y_6__7__1_), .CK(
        pe_1_5_7_net3876), .RN(pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_v[5]) );
  DFFR_X1 pe_1_5_7_int_q_reg_v_reg_4__2_ ( .D(int_data_y_6__7__2_), .CK(
        pe_1_5_7_net3876), .RN(pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_v[6]) );
  DFFR_X1 pe_1_5_7_int_q_reg_v_reg_4__3_ ( .D(int_data_y_6__7__3_), .CK(
        pe_1_5_7_net3876), .RN(pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_v[7]) );
  DFFR_X1 pe_1_5_7_int_q_reg_v_reg_5__0_ ( .D(int_data_y_6__7__0_), .CK(
        pe_1_5_7_net3881), .RN(pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_v[0]) );
  DFFR_X1 pe_1_5_7_int_q_reg_v_reg_5__1_ ( .D(int_data_y_6__7__1_), .CK(
        pe_1_5_7_net3881), .RN(pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_v[1]) );
  DFFR_X1 pe_1_5_7_int_q_reg_v_reg_5__2_ ( .D(int_data_y_6__7__2_), .CK(
        pe_1_5_7_net3881), .RN(pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_v[2]) );
  DFFR_X1 pe_1_5_7_int_q_reg_v_reg_5__3_ ( .D(int_data_y_6__7__3_), .CK(
        pe_1_5_7_net3881), .RN(pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_5_7_int_q_reg_h_reg_0__0_ ( .D(i_data_conv_h[8]), .SI(
        int_data_y_6__7__0_), .SE(pe_1_5_7_n65), .CK(pe_1_5_7_net3825), .RN(
        pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_5_7_int_q_reg_h_reg_0__1_ ( .D(i_data_conv_h[9]), .SI(
        int_data_y_6__7__1_), .SE(pe_1_5_7_n65), .CK(pe_1_5_7_net3825), .RN(
        pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_5_7_int_q_reg_h_reg_0__2_ ( .D(i_data_conv_h[10]), .SI(
        int_data_y_6__7__2_), .SE(pe_1_5_7_n65), .CK(pe_1_5_7_net3825), .RN(
        pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_5_7_int_q_reg_h_reg_0__3_ ( .D(i_data_conv_h[11]), .SI(
        int_data_y_6__7__3_), .SE(pe_1_5_7_n65), .CK(pe_1_5_7_net3825), .RN(
        pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_5_7_int_q_reg_h_reg_1__0_ ( .D(i_data_conv_h[8]), .SI(
        int_data_y_6__7__0_), .SE(pe_1_5_7_n65), .CK(pe_1_5_7_net3831), .RN(
        pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_5_7_int_q_reg_h_reg_1__1_ ( .D(i_data_conv_h[9]), .SI(
        int_data_y_6__7__1_), .SE(pe_1_5_7_n65), .CK(pe_1_5_7_net3831), .RN(
        pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_5_7_int_q_reg_h_reg_1__2_ ( .D(i_data_conv_h[10]), .SI(
        int_data_y_6__7__2_), .SE(pe_1_5_7_n65), .CK(pe_1_5_7_net3831), .RN(
        pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_5_7_int_q_reg_h_reg_1__3_ ( .D(i_data_conv_h[11]), .SI(
        int_data_y_6__7__3_), .SE(pe_1_5_7_n65), .CK(pe_1_5_7_net3831), .RN(
        pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_5_7_int_q_reg_h_reg_2__0_ ( .D(i_data_conv_h[8]), .SI(
        int_data_y_6__7__0_), .SE(pe_1_5_7_n65), .CK(pe_1_5_7_net3836), .RN(
        pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_5_7_int_q_reg_h_reg_2__1_ ( .D(i_data_conv_h[9]), .SI(
        int_data_y_6__7__1_), .SE(pe_1_5_7_n65), .CK(pe_1_5_7_net3836), .RN(
        pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_5_7_int_q_reg_h_reg_2__2_ ( .D(i_data_conv_h[10]), .SI(
        int_data_y_6__7__2_), .SE(pe_1_5_7_n65), .CK(pe_1_5_7_net3836), .RN(
        pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_5_7_int_q_reg_h_reg_2__3_ ( .D(i_data_conv_h[11]), .SI(
        int_data_y_6__7__3_), .SE(pe_1_5_7_n65), .CK(pe_1_5_7_net3836), .RN(
        pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_5_7_int_q_reg_h_reg_3__0_ ( .D(i_data_conv_h[8]), .SI(
        int_data_y_6__7__0_), .SE(pe_1_5_7_n65), .CK(pe_1_5_7_net3841), .RN(
        pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_5_7_int_q_reg_h_reg_3__1_ ( .D(i_data_conv_h[9]), .SI(
        int_data_y_6__7__1_), .SE(pe_1_5_7_n65), .CK(pe_1_5_7_net3841), .RN(
        pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_5_7_int_q_reg_h_reg_3__2_ ( .D(i_data_conv_h[10]), .SI(
        int_data_y_6__7__2_), .SE(pe_1_5_7_n65), .CK(pe_1_5_7_net3841), .RN(
        pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_5_7_int_q_reg_h_reg_3__3_ ( .D(i_data_conv_h[11]), .SI(
        int_data_y_6__7__3_), .SE(pe_1_5_7_n65), .CK(pe_1_5_7_net3841), .RN(
        pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_5_7_int_q_reg_h_reg_4__0_ ( .D(i_data_conv_h[8]), .SI(
        int_data_y_6__7__0_), .SE(pe_1_5_7_n66), .CK(pe_1_5_7_net3846), .RN(
        pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_5_7_int_q_reg_h_reg_4__1_ ( .D(i_data_conv_h[9]), .SI(
        int_data_y_6__7__1_), .SE(pe_1_5_7_n66), .CK(pe_1_5_7_net3846), .RN(
        pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_5_7_int_q_reg_h_reg_4__2_ ( .D(i_data_conv_h[10]), .SI(
        int_data_y_6__7__2_), .SE(pe_1_5_7_n66), .CK(pe_1_5_7_net3846), .RN(
        pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_5_7_int_q_reg_h_reg_4__3_ ( .D(i_data_conv_h[11]), .SI(
        int_data_y_6__7__3_), .SE(pe_1_5_7_n66), .CK(pe_1_5_7_net3846), .RN(
        pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_5_7_int_q_reg_h_reg_5__0_ ( .D(i_data_conv_h[8]), .SI(
        int_data_y_6__7__0_), .SE(pe_1_5_7_n66), .CK(pe_1_5_7_net3851), .RN(
        pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_5_7_int_q_reg_h_reg_5__1_ ( .D(i_data_conv_h[9]), .SI(
        int_data_y_6__7__1_), .SE(pe_1_5_7_n66), .CK(pe_1_5_7_net3851), .RN(
        pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_5_7_int_q_reg_h_reg_5__2_ ( .D(i_data_conv_h[10]), .SI(
        int_data_y_6__7__2_), .SE(pe_1_5_7_n66), .CK(pe_1_5_7_net3851), .RN(
        pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_5_7_int_q_reg_h_reg_5__3_ ( .D(i_data_conv_h[11]), .SI(
        int_data_y_6__7__3_), .SE(pe_1_5_7_n66), .CK(pe_1_5_7_net3851), .RN(
        pe_1_5_7_n72), .Q(pe_1_5_7_int_q_reg_h[3]) );
  FA_X1 pe_1_5_7_sub_81_U2_7 ( .A(int_data_res_5__7__7_), .B(pe_1_5_7_n76), 
        .CI(pe_1_5_7_sub_81_carry[7]), .S(pe_1_5_7_N77) );
  FA_X1 pe_1_5_7_sub_81_U2_6 ( .A(int_data_res_5__7__6_), .B(pe_1_5_7_n76), 
        .CI(pe_1_5_7_sub_81_carry[6]), .CO(pe_1_5_7_sub_81_carry[7]), .S(
        pe_1_5_7_N76) );
  FA_X1 pe_1_5_7_sub_81_U2_5 ( .A(int_data_res_5__7__5_), .B(pe_1_5_7_n76), 
        .CI(pe_1_5_7_sub_81_carry[5]), .CO(pe_1_5_7_sub_81_carry[6]), .S(
        pe_1_5_7_N75) );
  FA_X1 pe_1_5_7_sub_81_U2_4 ( .A(int_data_res_5__7__4_), .B(pe_1_5_7_n76), 
        .CI(pe_1_5_7_sub_81_carry[4]), .CO(pe_1_5_7_sub_81_carry[5]), .S(
        pe_1_5_7_N74) );
  FA_X1 pe_1_5_7_sub_81_U2_3 ( .A(int_data_res_5__7__3_), .B(pe_1_5_7_n76), 
        .CI(pe_1_5_7_sub_81_carry[3]), .CO(pe_1_5_7_sub_81_carry[4]), .S(
        pe_1_5_7_N73) );
  FA_X1 pe_1_5_7_sub_81_U2_2 ( .A(int_data_res_5__7__2_), .B(pe_1_5_7_n75), 
        .CI(pe_1_5_7_sub_81_carry[2]), .CO(pe_1_5_7_sub_81_carry[3]), .S(
        pe_1_5_7_N72) );
  FA_X1 pe_1_5_7_sub_81_U2_1 ( .A(int_data_res_5__7__1_), .B(pe_1_5_7_n74), 
        .CI(pe_1_5_7_sub_81_carry[1]), .CO(pe_1_5_7_sub_81_carry[2]), .S(
        pe_1_5_7_N71) );
  FA_X1 pe_1_5_7_add_83_U1_7 ( .A(int_data_res_5__7__7_), .B(
        pe_1_5_7_int_data_3_), .CI(pe_1_5_7_add_83_carry[7]), .S(pe_1_5_7_N85)
         );
  FA_X1 pe_1_5_7_add_83_U1_6 ( .A(int_data_res_5__7__6_), .B(
        pe_1_5_7_int_data_3_), .CI(pe_1_5_7_add_83_carry[6]), .CO(
        pe_1_5_7_add_83_carry[7]), .S(pe_1_5_7_N84) );
  FA_X1 pe_1_5_7_add_83_U1_5 ( .A(int_data_res_5__7__5_), .B(
        pe_1_5_7_int_data_3_), .CI(pe_1_5_7_add_83_carry[5]), .CO(
        pe_1_5_7_add_83_carry[6]), .S(pe_1_5_7_N83) );
  FA_X1 pe_1_5_7_add_83_U1_4 ( .A(int_data_res_5__7__4_), .B(
        pe_1_5_7_int_data_3_), .CI(pe_1_5_7_add_83_carry[4]), .CO(
        pe_1_5_7_add_83_carry[5]), .S(pe_1_5_7_N82) );
  FA_X1 pe_1_5_7_add_83_U1_3 ( .A(int_data_res_5__7__3_), .B(
        pe_1_5_7_int_data_3_), .CI(pe_1_5_7_add_83_carry[3]), .CO(
        pe_1_5_7_add_83_carry[4]), .S(pe_1_5_7_N81) );
  FA_X1 pe_1_5_7_add_83_U1_2 ( .A(int_data_res_5__7__2_), .B(
        pe_1_5_7_int_data_2_), .CI(pe_1_5_7_add_83_carry[2]), .CO(
        pe_1_5_7_add_83_carry[3]), .S(pe_1_5_7_N80) );
  FA_X1 pe_1_5_7_add_83_U1_1 ( .A(int_data_res_5__7__1_), .B(
        pe_1_5_7_int_data_1_), .CI(pe_1_5_7_n2), .CO(pe_1_5_7_add_83_carry[2]), 
        .S(pe_1_5_7_N79) );
  NAND3_X1 pe_1_5_7_U56 ( .A1(pe_1_5_7_n60), .A2(pe_1_5_7_n43), .A3(
        pe_1_5_7_n62), .ZN(pe_1_5_7_n40) );
  NAND3_X1 pe_1_5_7_U55 ( .A1(pe_1_5_7_n43), .A2(pe_1_5_7_n61), .A3(
        pe_1_5_7_n62), .ZN(pe_1_5_7_n39) );
  NAND3_X1 pe_1_5_7_U54 ( .A1(pe_1_5_7_n43), .A2(pe_1_5_7_n63), .A3(
        pe_1_5_7_n60), .ZN(pe_1_5_7_n38) );
  NAND3_X1 pe_1_5_7_U53 ( .A1(pe_1_5_7_n61), .A2(pe_1_5_7_n63), .A3(
        pe_1_5_7_n43), .ZN(pe_1_5_7_n37) );
  DFFR_X1 pe_1_5_7_int_q_acc_reg_6_ ( .D(pe_1_5_7_n78), .CK(pe_1_5_7_net3886), 
        .RN(pe_1_5_7_n71), .Q(int_data_res_5__7__6_) );
  DFFR_X1 pe_1_5_7_int_q_acc_reg_5_ ( .D(pe_1_5_7_n79), .CK(pe_1_5_7_net3886), 
        .RN(pe_1_5_7_n71), .Q(int_data_res_5__7__5_) );
  DFFR_X1 pe_1_5_7_int_q_acc_reg_4_ ( .D(pe_1_5_7_n80), .CK(pe_1_5_7_net3886), 
        .RN(pe_1_5_7_n71), .Q(int_data_res_5__7__4_) );
  DFFR_X1 pe_1_5_7_int_q_acc_reg_3_ ( .D(pe_1_5_7_n81), .CK(pe_1_5_7_net3886), 
        .RN(pe_1_5_7_n71), .Q(int_data_res_5__7__3_) );
  DFFR_X1 pe_1_5_7_int_q_acc_reg_2_ ( .D(pe_1_5_7_n82), .CK(pe_1_5_7_net3886), 
        .RN(pe_1_5_7_n71), .Q(int_data_res_5__7__2_) );
  DFFR_X1 pe_1_5_7_int_q_acc_reg_1_ ( .D(pe_1_5_7_n83), .CK(pe_1_5_7_net3886), 
        .RN(pe_1_5_7_n71), .Q(int_data_res_5__7__1_) );
  DFFR_X1 pe_1_5_7_int_q_acc_reg_7_ ( .D(pe_1_5_7_n77), .CK(pe_1_5_7_net3886), 
        .RN(pe_1_5_7_n71), .Q(int_data_res_5__7__7_) );
  CLKGATETST_X1 pe_1_5_7_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_5_7_n88), .SE(1'b0), .GCK(pe_1_5_7_net3825) );
  CLKGATETST_X1 pe_1_5_7_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_5_7_n87), .SE(1'b0), .GCK(pe_1_5_7_net3831) );
  CLKGATETST_X1 pe_1_5_7_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_5_7_n86), .SE(1'b0), .GCK(pe_1_5_7_net3836) );
  CLKGATETST_X1 pe_1_5_7_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_5_7_n85), .SE(1'b0), .GCK(pe_1_5_7_net3841) );
  CLKGATETST_X1 pe_1_5_7_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_5_7_n90), .SE(1'b0), .GCK(pe_1_5_7_net3846) );
  CLKGATETST_X1 pe_1_5_7_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_5_7_n89), .SE(1'b0), .GCK(pe_1_5_7_net3851) );
  CLKGATETST_X1 pe_1_5_7_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_5_7_N64), .SE(1'b0), .GCK(pe_1_5_7_net3856) );
  CLKGATETST_X1 pe_1_5_7_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_5_7_N63), .SE(1'b0), .GCK(pe_1_5_7_net3861) );
  CLKGATETST_X1 pe_1_5_7_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_5_7_N62), .SE(1'b0), .GCK(pe_1_5_7_net3866) );
  CLKGATETST_X1 pe_1_5_7_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_5_7_N61), .SE(1'b0), .GCK(pe_1_5_7_net3871) );
  CLKGATETST_X1 pe_1_5_7_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_5_7_N60), .SE(1'b0), .GCK(pe_1_5_7_net3876) );
  CLKGATETST_X1 pe_1_5_7_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_5_7_N59), .SE(1'b0), .GCK(pe_1_5_7_net3881) );
  CLKGATETST_X1 pe_1_5_7_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_5_7_N90), .SE(1'b0), .GCK(pe_1_5_7_net3886) );
  CLKBUF_X1 pe_1_6_0_U109 ( .A(pe_1_6_0_n69), .Z(pe_1_6_0_n68) );
  INV_X1 pe_1_6_0_U108 ( .A(n77), .ZN(pe_1_6_0_n67) );
  INV_X1 pe_1_6_0_U107 ( .A(n69), .ZN(pe_1_6_0_n66) );
  INV_X1 pe_1_6_0_U106 ( .A(n69), .ZN(pe_1_6_0_n65) );
  INV_X1 pe_1_6_0_U105 ( .A(pe_1_6_0_n66), .ZN(pe_1_6_0_n64) );
  INV_X1 pe_1_6_0_U104 ( .A(pe_1_6_0_n61), .ZN(pe_1_6_0_n60) );
  INV_X1 pe_1_6_0_U103 ( .A(n29), .ZN(pe_1_6_0_n58) );
  INV_X1 pe_1_6_0_U102 ( .A(n21), .ZN(pe_1_6_0_n57) );
  MUX2_X1 pe_1_6_0_U101 ( .A(pe_1_6_0_n54), .B(pe_1_6_0_n51), .S(n52), .Z(
        pe_1_6_0_o_data_h_3_) );
  MUX2_X1 pe_1_6_0_U100 ( .A(pe_1_6_0_n53), .B(pe_1_6_0_n52), .S(pe_1_6_0_n60), 
        .Z(pe_1_6_0_n54) );
  MUX2_X1 pe_1_6_0_U99 ( .A(pe_1_6_0_int_q_reg_h[23]), .B(
        pe_1_6_0_int_q_reg_h[19]), .S(pe_1_6_0_n56), .Z(pe_1_6_0_n53) );
  MUX2_X1 pe_1_6_0_U98 ( .A(pe_1_6_0_int_q_reg_h[15]), .B(
        pe_1_6_0_int_q_reg_h[11]), .S(pe_1_6_0_n56), .Z(pe_1_6_0_n52) );
  MUX2_X1 pe_1_6_0_U97 ( .A(pe_1_6_0_int_q_reg_h[7]), .B(
        pe_1_6_0_int_q_reg_h[3]), .S(pe_1_6_0_n56), .Z(pe_1_6_0_n51) );
  MUX2_X1 pe_1_6_0_U96 ( .A(pe_1_6_0_n50), .B(pe_1_6_0_n47), .S(n52), .Z(
        pe_1_6_0_o_data_h_2_) );
  MUX2_X1 pe_1_6_0_U95 ( .A(pe_1_6_0_n49), .B(pe_1_6_0_n48), .S(pe_1_6_0_n60), 
        .Z(pe_1_6_0_n50) );
  MUX2_X1 pe_1_6_0_U94 ( .A(pe_1_6_0_int_q_reg_h[22]), .B(
        pe_1_6_0_int_q_reg_h[18]), .S(pe_1_6_0_n56), .Z(pe_1_6_0_n49) );
  MUX2_X1 pe_1_6_0_U93 ( .A(pe_1_6_0_int_q_reg_h[14]), .B(
        pe_1_6_0_int_q_reg_h[10]), .S(pe_1_6_0_n56), .Z(pe_1_6_0_n48) );
  MUX2_X1 pe_1_6_0_U92 ( .A(pe_1_6_0_int_q_reg_h[6]), .B(
        pe_1_6_0_int_q_reg_h[2]), .S(pe_1_6_0_n56), .Z(pe_1_6_0_n47) );
  MUX2_X1 pe_1_6_0_U91 ( .A(pe_1_6_0_n46), .B(pe_1_6_0_n24), .S(n52), .Z(
        pe_1_6_0_o_data_h_1_) );
  MUX2_X1 pe_1_6_0_U90 ( .A(pe_1_6_0_n45), .B(pe_1_6_0_n25), .S(pe_1_6_0_n60), 
        .Z(pe_1_6_0_n46) );
  MUX2_X1 pe_1_6_0_U89 ( .A(pe_1_6_0_int_q_reg_h[21]), .B(
        pe_1_6_0_int_q_reg_h[17]), .S(pe_1_6_0_n56), .Z(pe_1_6_0_n45) );
  MUX2_X1 pe_1_6_0_U88 ( .A(pe_1_6_0_int_q_reg_h[13]), .B(
        pe_1_6_0_int_q_reg_h[9]), .S(pe_1_6_0_n56), .Z(pe_1_6_0_n25) );
  MUX2_X1 pe_1_6_0_U87 ( .A(pe_1_6_0_int_q_reg_h[5]), .B(
        pe_1_6_0_int_q_reg_h[1]), .S(pe_1_6_0_n56), .Z(pe_1_6_0_n24) );
  MUX2_X1 pe_1_6_0_U86 ( .A(pe_1_6_0_n23), .B(pe_1_6_0_n20), .S(n52), .Z(
        pe_1_6_0_o_data_h_0_) );
  MUX2_X1 pe_1_6_0_U85 ( .A(pe_1_6_0_n22), .B(pe_1_6_0_n21), .S(pe_1_6_0_n60), 
        .Z(pe_1_6_0_n23) );
  MUX2_X1 pe_1_6_0_U84 ( .A(pe_1_6_0_int_q_reg_h[20]), .B(
        pe_1_6_0_int_q_reg_h[16]), .S(pe_1_6_0_n56), .Z(pe_1_6_0_n22) );
  MUX2_X1 pe_1_6_0_U83 ( .A(pe_1_6_0_int_q_reg_h[12]), .B(
        pe_1_6_0_int_q_reg_h[8]), .S(pe_1_6_0_n56), .Z(pe_1_6_0_n21) );
  MUX2_X1 pe_1_6_0_U82 ( .A(pe_1_6_0_int_q_reg_h[4]), .B(
        pe_1_6_0_int_q_reg_h[0]), .S(pe_1_6_0_n56), .Z(pe_1_6_0_n20) );
  MUX2_X1 pe_1_6_0_U81 ( .A(pe_1_6_0_n19), .B(pe_1_6_0_n16), .S(n52), .Z(
        int_data_y_6__0__3_) );
  MUX2_X1 pe_1_6_0_U80 ( .A(pe_1_6_0_n18), .B(pe_1_6_0_n17), .S(pe_1_6_0_n60), 
        .Z(pe_1_6_0_n19) );
  MUX2_X1 pe_1_6_0_U79 ( .A(pe_1_6_0_int_q_reg_v[23]), .B(
        pe_1_6_0_int_q_reg_v[19]), .S(pe_1_6_0_n55), .Z(pe_1_6_0_n18) );
  MUX2_X1 pe_1_6_0_U78 ( .A(pe_1_6_0_int_q_reg_v[15]), .B(
        pe_1_6_0_int_q_reg_v[11]), .S(pe_1_6_0_n55), .Z(pe_1_6_0_n17) );
  MUX2_X1 pe_1_6_0_U77 ( .A(pe_1_6_0_int_q_reg_v[7]), .B(
        pe_1_6_0_int_q_reg_v[3]), .S(pe_1_6_0_n55), .Z(pe_1_6_0_n16) );
  MUX2_X1 pe_1_6_0_U76 ( .A(pe_1_6_0_n15), .B(pe_1_6_0_n12), .S(n52), .Z(
        int_data_y_6__0__2_) );
  MUX2_X1 pe_1_6_0_U75 ( .A(pe_1_6_0_n14), .B(pe_1_6_0_n13), .S(pe_1_6_0_n60), 
        .Z(pe_1_6_0_n15) );
  MUX2_X1 pe_1_6_0_U74 ( .A(pe_1_6_0_int_q_reg_v[22]), .B(
        pe_1_6_0_int_q_reg_v[18]), .S(pe_1_6_0_n55), .Z(pe_1_6_0_n14) );
  MUX2_X1 pe_1_6_0_U73 ( .A(pe_1_6_0_int_q_reg_v[14]), .B(
        pe_1_6_0_int_q_reg_v[10]), .S(pe_1_6_0_n55), .Z(pe_1_6_0_n13) );
  MUX2_X1 pe_1_6_0_U72 ( .A(pe_1_6_0_int_q_reg_v[6]), .B(
        pe_1_6_0_int_q_reg_v[2]), .S(pe_1_6_0_n55), .Z(pe_1_6_0_n12) );
  MUX2_X1 pe_1_6_0_U71 ( .A(pe_1_6_0_n11), .B(pe_1_6_0_n8), .S(n52), .Z(
        int_data_y_6__0__1_) );
  MUX2_X1 pe_1_6_0_U70 ( .A(pe_1_6_0_n10), .B(pe_1_6_0_n9), .S(pe_1_6_0_n60), 
        .Z(pe_1_6_0_n11) );
  MUX2_X1 pe_1_6_0_U69 ( .A(pe_1_6_0_int_q_reg_v[21]), .B(
        pe_1_6_0_int_q_reg_v[17]), .S(pe_1_6_0_n55), .Z(pe_1_6_0_n10) );
  MUX2_X1 pe_1_6_0_U68 ( .A(pe_1_6_0_int_q_reg_v[13]), .B(
        pe_1_6_0_int_q_reg_v[9]), .S(pe_1_6_0_n55), .Z(pe_1_6_0_n9) );
  MUX2_X1 pe_1_6_0_U67 ( .A(pe_1_6_0_int_q_reg_v[5]), .B(
        pe_1_6_0_int_q_reg_v[1]), .S(pe_1_6_0_n55), .Z(pe_1_6_0_n8) );
  MUX2_X1 pe_1_6_0_U66 ( .A(pe_1_6_0_n7), .B(pe_1_6_0_n4), .S(n52), .Z(
        int_data_y_6__0__0_) );
  MUX2_X1 pe_1_6_0_U65 ( .A(pe_1_6_0_n6), .B(pe_1_6_0_n5), .S(pe_1_6_0_n60), 
        .Z(pe_1_6_0_n7) );
  MUX2_X1 pe_1_6_0_U64 ( .A(pe_1_6_0_int_q_reg_v[20]), .B(
        pe_1_6_0_int_q_reg_v[16]), .S(pe_1_6_0_n55), .Z(pe_1_6_0_n6) );
  MUX2_X1 pe_1_6_0_U63 ( .A(pe_1_6_0_int_q_reg_v[12]), .B(
        pe_1_6_0_int_q_reg_v[8]), .S(pe_1_6_0_n55), .Z(pe_1_6_0_n5) );
  MUX2_X1 pe_1_6_0_U62 ( .A(pe_1_6_0_int_q_reg_v[4]), .B(
        pe_1_6_0_int_q_reg_v[0]), .S(pe_1_6_0_n55), .Z(pe_1_6_0_n4) );
  AND2_X1 pe_1_6_0_U61 ( .A1(pe_1_6_0_o_data_h_3_), .A2(n29), .ZN(
        pe_1_6_0_int_data_3_) );
  NAND2_X1 pe_1_6_0_U60 ( .A1(pe_1_6_0_int_data_0_), .A2(pe_1_6_0_n3), .ZN(
        pe_1_6_0_sub_81_carry[1]) );
  INV_X1 pe_1_6_0_U59 ( .A(pe_1_6_0_int_data_1_), .ZN(pe_1_6_0_n71) );
  AOI222_X1 pe_1_6_0_U58 ( .A1(pe_1_6_0_n62), .A2(int_data_res_7__0__7_), .B1(
        pe_1_6_0_N85), .B2(pe_1_6_0_n27), .C1(pe_1_6_0_N77), .C2(pe_1_6_0_n28), 
        .ZN(pe_1_6_0_n26) );
  INV_X1 pe_1_6_0_U57 ( .A(pe_1_6_0_n26), .ZN(pe_1_6_0_n74) );
  AOI222_X1 pe_1_6_0_U52 ( .A1(int_data_res_7__0__1_), .A2(pe_1_6_0_n62), .B1(
        pe_1_6_0_N79), .B2(pe_1_6_0_n27), .C1(pe_1_6_0_N71), .C2(pe_1_6_0_n28), 
        .ZN(pe_1_6_0_n34) );
  INV_X1 pe_1_6_0_U51 ( .A(pe_1_6_0_n34), .ZN(pe_1_6_0_n80) );
  AOI222_X1 pe_1_6_0_U50 ( .A1(int_data_res_7__0__2_), .A2(pe_1_6_0_n62), .B1(
        pe_1_6_0_N80), .B2(pe_1_6_0_n27), .C1(pe_1_6_0_N72), .C2(pe_1_6_0_n28), 
        .ZN(pe_1_6_0_n33) );
  INV_X1 pe_1_6_0_U49 ( .A(pe_1_6_0_n33), .ZN(pe_1_6_0_n79) );
  AOI222_X1 pe_1_6_0_U48 ( .A1(int_data_res_7__0__6_), .A2(pe_1_6_0_n62), .B1(
        pe_1_6_0_N84), .B2(pe_1_6_0_n27), .C1(pe_1_6_0_N76), .C2(pe_1_6_0_n28), 
        .ZN(pe_1_6_0_n29) );
  INV_X1 pe_1_6_0_U47 ( .A(pe_1_6_0_n29), .ZN(pe_1_6_0_n75) );
  AND2_X1 pe_1_6_0_U46 ( .A1(pe_1_6_0_o_data_h_2_), .A2(n29), .ZN(
        pe_1_6_0_int_data_2_) );
  AND2_X1 pe_1_6_0_U45 ( .A1(pe_1_6_0_o_data_h_1_), .A2(n29), .ZN(
        pe_1_6_0_int_data_1_) );
  INV_X1 pe_1_6_0_U44 ( .A(pe_1_6_0_int_data_2_), .ZN(pe_1_6_0_n72) );
  AND2_X1 pe_1_6_0_U43 ( .A1(pe_1_6_0_int_data_0_), .A2(int_data_res_6__0__0_), 
        .ZN(pe_1_6_0_n2) );
  AND2_X1 pe_1_6_0_U42 ( .A1(pe_1_6_0_o_data_h_0_), .A2(n29), .ZN(
        pe_1_6_0_int_data_0_) );
  XNOR2_X1 pe_1_6_0_U41 ( .A(pe_1_6_0_n70), .B(int_data_res_6__0__0_), .ZN(
        pe_1_6_0_N70) );
  AOI222_X1 pe_1_6_0_U40 ( .A1(int_data_res_7__0__0_), .A2(pe_1_6_0_n62), .B1(
        pe_1_6_0_n1), .B2(pe_1_6_0_n27), .C1(pe_1_6_0_N70), .C2(pe_1_6_0_n28), 
        .ZN(pe_1_6_0_n35) );
  INV_X1 pe_1_6_0_U39 ( .A(pe_1_6_0_n35), .ZN(pe_1_6_0_n81) );
  AOI222_X1 pe_1_6_0_U38 ( .A1(int_data_res_7__0__3_), .A2(pe_1_6_0_n62), .B1(
        pe_1_6_0_N81), .B2(pe_1_6_0_n27), .C1(pe_1_6_0_N73), .C2(pe_1_6_0_n28), 
        .ZN(pe_1_6_0_n32) );
  INV_X1 pe_1_6_0_U37 ( .A(pe_1_6_0_n32), .ZN(pe_1_6_0_n78) );
  AOI222_X1 pe_1_6_0_U36 ( .A1(int_data_res_7__0__4_), .A2(pe_1_6_0_n62), .B1(
        pe_1_6_0_N82), .B2(pe_1_6_0_n27), .C1(pe_1_6_0_N74), .C2(pe_1_6_0_n28), 
        .ZN(pe_1_6_0_n31) );
  INV_X1 pe_1_6_0_U35 ( .A(pe_1_6_0_n31), .ZN(pe_1_6_0_n77) );
  AOI222_X1 pe_1_6_0_U34 ( .A1(int_data_res_7__0__5_), .A2(pe_1_6_0_n62), .B1(
        pe_1_6_0_N83), .B2(pe_1_6_0_n27), .C1(pe_1_6_0_N75), .C2(pe_1_6_0_n28), 
        .ZN(pe_1_6_0_n30) );
  INV_X1 pe_1_6_0_U33 ( .A(pe_1_6_0_n30), .ZN(pe_1_6_0_n76) );
  NOR3_X1 pe_1_6_0_U32 ( .A1(pe_1_6_0_n58), .A2(pe_1_6_0_n63), .A3(int_ckg[15]), .ZN(pe_1_6_0_n36) );
  OR2_X1 pe_1_6_0_U31 ( .A1(pe_1_6_0_n36), .A2(pe_1_6_0_n62), .ZN(pe_1_6_0_N90) );
  INV_X1 pe_1_6_0_U30 ( .A(pe_1_6_0_int_data_0_), .ZN(pe_1_6_0_n70) );
  INV_X1 pe_1_6_0_U29 ( .A(n41), .ZN(pe_1_6_0_n61) );
  INV_X1 pe_1_6_0_U28 ( .A(n35), .ZN(pe_1_6_0_n59) );
  INV_X1 pe_1_6_0_U27 ( .A(pe_1_6_0_int_data_3_), .ZN(pe_1_6_0_n73) );
  BUF_X1 pe_1_6_0_U26 ( .A(n63), .Z(pe_1_6_0_n62) );
  NAND2_X1 pe_1_6_0_U25 ( .A1(pe_1_6_0_n44), .A2(pe_1_6_0_n59), .ZN(
        pe_1_6_0_n41) );
  AND3_X1 pe_1_6_0_U24 ( .A1(n77), .A2(pe_1_6_0_n61), .A3(n52), .ZN(
        pe_1_6_0_n44) );
  NOR2_X1 pe_1_6_0_U23 ( .A1(pe_1_6_0_n67), .A2(n52), .ZN(pe_1_6_0_n43) );
  NOR2_X1 pe_1_6_0_U22 ( .A1(pe_1_6_0_n57), .A2(pe_1_6_0_n62), .ZN(
        pe_1_6_0_n28) );
  NOR2_X1 pe_1_6_0_U21 ( .A1(n21), .A2(pe_1_6_0_n62), .ZN(pe_1_6_0_n27) );
  INV_X1 pe_1_6_0_U20 ( .A(pe_1_6_0_n41), .ZN(pe_1_6_0_n87) );
  INV_X1 pe_1_6_0_U19 ( .A(pe_1_6_0_n37), .ZN(pe_1_6_0_n85) );
  INV_X1 pe_1_6_0_U18 ( .A(pe_1_6_0_n38), .ZN(pe_1_6_0_n84) );
  INV_X1 pe_1_6_0_U17 ( .A(pe_1_6_0_n39), .ZN(pe_1_6_0_n83) );
  NOR2_X1 pe_1_6_0_U16 ( .A1(pe_1_6_0_n65), .A2(pe_1_6_0_n42), .ZN(
        pe_1_6_0_N59) );
  NOR2_X1 pe_1_6_0_U15 ( .A1(pe_1_6_0_n65), .A2(pe_1_6_0_n41), .ZN(
        pe_1_6_0_N60) );
  NOR2_X1 pe_1_6_0_U14 ( .A1(pe_1_6_0_n65), .A2(pe_1_6_0_n38), .ZN(
        pe_1_6_0_N63) );
  NOR2_X1 pe_1_6_0_U13 ( .A1(pe_1_6_0_n65), .A2(pe_1_6_0_n40), .ZN(
        pe_1_6_0_N61) );
  NOR2_X1 pe_1_6_0_U12 ( .A1(pe_1_6_0_n65), .A2(pe_1_6_0_n39), .ZN(
        pe_1_6_0_N62) );
  NOR2_X1 pe_1_6_0_U11 ( .A1(pe_1_6_0_n37), .A2(pe_1_6_0_n65), .ZN(
        pe_1_6_0_N64) );
  NAND2_X1 pe_1_6_0_U10 ( .A1(pe_1_6_0_n44), .A2(n35), .ZN(pe_1_6_0_n42) );
  BUF_X1 pe_1_6_0_U9 ( .A(n35), .Z(pe_1_6_0_n55) );
  BUF_X1 pe_1_6_0_U8 ( .A(n35), .Z(pe_1_6_0_n56) );
  INV_X1 pe_1_6_0_U7 ( .A(pe_1_6_0_n66), .ZN(pe_1_6_0_n63) );
  INV_X1 pe_1_6_0_U6 ( .A(pe_1_6_0_n42), .ZN(pe_1_6_0_n86) );
  INV_X1 pe_1_6_0_U5 ( .A(pe_1_6_0_n40), .ZN(pe_1_6_0_n82) );
  INV_X2 pe_1_6_0_U4 ( .A(n85), .ZN(pe_1_6_0_n69) );
  XOR2_X1 pe_1_6_0_U3 ( .A(pe_1_6_0_int_data_0_), .B(int_data_res_6__0__0_), 
        .Z(pe_1_6_0_n1) );
  DFFR_X1 pe_1_6_0_int_q_acc_reg_0_ ( .D(pe_1_6_0_n81), .CK(pe_1_6_0_net3808), 
        .RN(pe_1_6_0_n69), .Q(int_data_res_6__0__0_), .QN(pe_1_6_0_n3) );
  DFFR_X1 pe_1_6_0_int_q_reg_v_reg_0__0_ ( .D(int_data_y_7__0__0_), .CK(
        pe_1_6_0_net3778), .RN(pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_v[20]) );
  DFFR_X1 pe_1_6_0_int_q_reg_v_reg_0__1_ ( .D(int_data_y_7__0__1_), .CK(
        pe_1_6_0_net3778), .RN(pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_v[21]) );
  DFFR_X1 pe_1_6_0_int_q_reg_v_reg_0__2_ ( .D(int_data_y_7__0__2_), .CK(
        pe_1_6_0_net3778), .RN(pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_v[22]) );
  DFFR_X1 pe_1_6_0_int_q_reg_v_reg_0__3_ ( .D(int_data_y_7__0__3_), .CK(
        pe_1_6_0_net3778), .RN(pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_v[23]) );
  DFFR_X1 pe_1_6_0_int_q_reg_v_reg_1__0_ ( .D(int_data_y_7__0__0_), .CK(
        pe_1_6_0_net3783), .RN(pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_v[16]) );
  DFFR_X1 pe_1_6_0_int_q_reg_v_reg_1__1_ ( .D(int_data_y_7__0__1_), .CK(
        pe_1_6_0_net3783), .RN(pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_v[17]) );
  DFFR_X1 pe_1_6_0_int_q_reg_v_reg_1__2_ ( .D(int_data_y_7__0__2_), .CK(
        pe_1_6_0_net3783), .RN(pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_v[18]) );
  DFFR_X1 pe_1_6_0_int_q_reg_v_reg_1__3_ ( .D(int_data_y_7__0__3_), .CK(
        pe_1_6_0_net3783), .RN(pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_v[19]) );
  DFFR_X1 pe_1_6_0_int_q_reg_v_reg_2__0_ ( .D(int_data_y_7__0__0_), .CK(
        pe_1_6_0_net3788), .RN(pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_v[12]) );
  DFFR_X1 pe_1_6_0_int_q_reg_v_reg_2__1_ ( .D(int_data_y_7__0__1_), .CK(
        pe_1_6_0_net3788), .RN(pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_v[13]) );
  DFFR_X1 pe_1_6_0_int_q_reg_v_reg_2__2_ ( .D(int_data_y_7__0__2_), .CK(
        pe_1_6_0_net3788), .RN(pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_v[14]) );
  DFFR_X1 pe_1_6_0_int_q_reg_v_reg_2__3_ ( .D(int_data_y_7__0__3_), .CK(
        pe_1_6_0_net3788), .RN(pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_v[15]) );
  DFFR_X1 pe_1_6_0_int_q_reg_v_reg_3__0_ ( .D(int_data_y_7__0__0_), .CK(
        pe_1_6_0_net3793), .RN(pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_v[8]) );
  DFFR_X1 pe_1_6_0_int_q_reg_v_reg_3__1_ ( .D(int_data_y_7__0__1_), .CK(
        pe_1_6_0_net3793), .RN(pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_v[9]) );
  DFFR_X1 pe_1_6_0_int_q_reg_v_reg_3__2_ ( .D(int_data_y_7__0__2_), .CK(
        pe_1_6_0_net3793), .RN(pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_v[10]) );
  DFFR_X1 pe_1_6_0_int_q_reg_v_reg_3__3_ ( .D(int_data_y_7__0__3_), .CK(
        pe_1_6_0_net3793), .RN(pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_v[11]) );
  DFFR_X1 pe_1_6_0_int_q_reg_v_reg_4__0_ ( .D(int_data_y_7__0__0_), .CK(
        pe_1_6_0_net3798), .RN(pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_v[4]) );
  DFFR_X1 pe_1_6_0_int_q_reg_v_reg_4__1_ ( .D(int_data_y_7__0__1_), .CK(
        pe_1_6_0_net3798), .RN(pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_v[5]) );
  DFFR_X1 pe_1_6_0_int_q_reg_v_reg_4__2_ ( .D(int_data_y_7__0__2_), .CK(
        pe_1_6_0_net3798), .RN(pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_v[6]) );
  DFFR_X1 pe_1_6_0_int_q_reg_v_reg_4__3_ ( .D(int_data_y_7__0__3_), .CK(
        pe_1_6_0_net3798), .RN(pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_v[7]) );
  DFFR_X1 pe_1_6_0_int_q_reg_v_reg_5__0_ ( .D(int_data_y_7__0__0_), .CK(
        pe_1_6_0_net3803), .RN(pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_v[0]) );
  DFFR_X1 pe_1_6_0_int_q_reg_v_reg_5__1_ ( .D(int_data_y_7__0__1_), .CK(
        pe_1_6_0_net3803), .RN(pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_v[1]) );
  DFFR_X1 pe_1_6_0_int_q_reg_v_reg_5__2_ ( .D(int_data_y_7__0__2_), .CK(
        pe_1_6_0_net3803), .RN(pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_v[2]) );
  DFFR_X1 pe_1_6_0_int_q_reg_v_reg_5__3_ ( .D(int_data_y_7__0__3_), .CK(
        pe_1_6_0_net3803), .RN(pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_6_0_int_q_reg_h_reg_0__0_ ( .D(int_data_x_6__1__0_), .SI(
        int_data_y_7__0__0_), .SE(pe_1_6_0_n63), .CK(pe_1_6_0_net3747), .RN(
        pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_6_0_int_q_reg_h_reg_0__1_ ( .D(int_data_x_6__1__1_), .SI(
        int_data_y_7__0__1_), .SE(pe_1_6_0_n63), .CK(pe_1_6_0_net3747), .RN(
        pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_6_0_int_q_reg_h_reg_0__2_ ( .D(int_data_x_6__1__2_), .SI(
        int_data_y_7__0__2_), .SE(pe_1_6_0_n63), .CK(pe_1_6_0_net3747), .RN(
        pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_6_0_int_q_reg_h_reg_0__3_ ( .D(int_data_x_6__1__3_), .SI(
        int_data_y_7__0__3_), .SE(pe_1_6_0_n63), .CK(pe_1_6_0_net3747), .RN(
        pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_6_0_int_q_reg_h_reg_1__0_ ( .D(int_data_x_6__1__0_), .SI(
        int_data_y_7__0__0_), .SE(pe_1_6_0_n63), .CK(pe_1_6_0_net3753), .RN(
        pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_6_0_int_q_reg_h_reg_1__1_ ( .D(int_data_x_6__1__1_), .SI(
        int_data_y_7__0__1_), .SE(pe_1_6_0_n63), .CK(pe_1_6_0_net3753), .RN(
        pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_6_0_int_q_reg_h_reg_1__2_ ( .D(int_data_x_6__1__2_), .SI(
        int_data_y_7__0__2_), .SE(pe_1_6_0_n63), .CK(pe_1_6_0_net3753), .RN(
        pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_6_0_int_q_reg_h_reg_1__3_ ( .D(int_data_x_6__1__3_), .SI(
        int_data_y_7__0__3_), .SE(pe_1_6_0_n63), .CK(pe_1_6_0_net3753), .RN(
        pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_6_0_int_q_reg_h_reg_2__0_ ( .D(int_data_x_6__1__0_), .SI(
        int_data_y_7__0__0_), .SE(pe_1_6_0_n63), .CK(pe_1_6_0_net3758), .RN(
        pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_6_0_int_q_reg_h_reg_2__1_ ( .D(int_data_x_6__1__1_), .SI(
        int_data_y_7__0__1_), .SE(pe_1_6_0_n63), .CK(pe_1_6_0_net3758), .RN(
        pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_6_0_int_q_reg_h_reg_2__2_ ( .D(int_data_x_6__1__2_), .SI(
        int_data_y_7__0__2_), .SE(pe_1_6_0_n63), .CK(pe_1_6_0_net3758), .RN(
        pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_6_0_int_q_reg_h_reg_2__3_ ( .D(int_data_x_6__1__3_), .SI(
        int_data_y_7__0__3_), .SE(pe_1_6_0_n63), .CK(pe_1_6_0_net3758), .RN(
        pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_6_0_int_q_reg_h_reg_3__0_ ( .D(int_data_x_6__1__0_), .SI(
        int_data_y_7__0__0_), .SE(pe_1_6_0_n63), .CK(pe_1_6_0_net3763), .RN(
        pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_6_0_int_q_reg_h_reg_3__1_ ( .D(int_data_x_6__1__1_), .SI(
        int_data_y_7__0__1_), .SE(pe_1_6_0_n63), .CK(pe_1_6_0_net3763), .RN(
        pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_6_0_int_q_reg_h_reg_3__2_ ( .D(int_data_x_6__1__2_), .SI(
        int_data_y_7__0__2_), .SE(pe_1_6_0_n63), .CK(pe_1_6_0_net3763), .RN(
        pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_6_0_int_q_reg_h_reg_3__3_ ( .D(int_data_x_6__1__3_), .SI(
        int_data_y_7__0__3_), .SE(pe_1_6_0_n63), .CK(pe_1_6_0_net3763), .RN(
        pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_6_0_int_q_reg_h_reg_4__0_ ( .D(int_data_x_6__1__0_), .SI(
        int_data_y_7__0__0_), .SE(pe_1_6_0_n64), .CK(pe_1_6_0_net3768), .RN(
        pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_6_0_int_q_reg_h_reg_4__1_ ( .D(int_data_x_6__1__1_), .SI(
        int_data_y_7__0__1_), .SE(pe_1_6_0_n64), .CK(pe_1_6_0_net3768), .RN(
        pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_6_0_int_q_reg_h_reg_4__2_ ( .D(int_data_x_6__1__2_), .SI(
        int_data_y_7__0__2_), .SE(pe_1_6_0_n64), .CK(pe_1_6_0_net3768), .RN(
        pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_6_0_int_q_reg_h_reg_4__3_ ( .D(int_data_x_6__1__3_), .SI(
        int_data_y_7__0__3_), .SE(pe_1_6_0_n64), .CK(pe_1_6_0_net3768), .RN(
        pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_6_0_int_q_reg_h_reg_5__0_ ( .D(int_data_x_6__1__0_), .SI(
        int_data_y_7__0__0_), .SE(pe_1_6_0_n64), .CK(pe_1_6_0_net3773), .RN(
        pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_6_0_int_q_reg_h_reg_5__1_ ( .D(int_data_x_6__1__1_), .SI(
        int_data_y_7__0__1_), .SE(pe_1_6_0_n64), .CK(pe_1_6_0_net3773), .RN(
        pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_6_0_int_q_reg_h_reg_5__2_ ( .D(int_data_x_6__1__2_), .SI(
        int_data_y_7__0__2_), .SE(pe_1_6_0_n64), .CK(pe_1_6_0_net3773), .RN(
        pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_6_0_int_q_reg_h_reg_5__3_ ( .D(int_data_x_6__1__3_), .SI(
        int_data_y_7__0__3_), .SE(pe_1_6_0_n64), .CK(pe_1_6_0_net3773), .RN(
        pe_1_6_0_n69), .Q(pe_1_6_0_int_q_reg_h[3]) );
  FA_X1 pe_1_6_0_sub_81_U2_7 ( .A(int_data_res_6__0__7_), .B(pe_1_6_0_n73), 
        .CI(pe_1_6_0_sub_81_carry[7]), .S(pe_1_6_0_N77) );
  FA_X1 pe_1_6_0_sub_81_U2_6 ( .A(int_data_res_6__0__6_), .B(pe_1_6_0_n73), 
        .CI(pe_1_6_0_sub_81_carry[6]), .CO(pe_1_6_0_sub_81_carry[7]), .S(
        pe_1_6_0_N76) );
  FA_X1 pe_1_6_0_sub_81_U2_5 ( .A(int_data_res_6__0__5_), .B(pe_1_6_0_n73), 
        .CI(pe_1_6_0_sub_81_carry[5]), .CO(pe_1_6_0_sub_81_carry[6]), .S(
        pe_1_6_0_N75) );
  FA_X1 pe_1_6_0_sub_81_U2_4 ( .A(int_data_res_6__0__4_), .B(pe_1_6_0_n73), 
        .CI(pe_1_6_0_sub_81_carry[4]), .CO(pe_1_6_0_sub_81_carry[5]), .S(
        pe_1_6_0_N74) );
  FA_X1 pe_1_6_0_sub_81_U2_3 ( .A(int_data_res_6__0__3_), .B(pe_1_6_0_n73), 
        .CI(pe_1_6_0_sub_81_carry[3]), .CO(pe_1_6_0_sub_81_carry[4]), .S(
        pe_1_6_0_N73) );
  FA_X1 pe_1_6_0_sub_81_U2_2 ( .A(int_data_res_6__0__2_), .B(pe_1_6_0_n72), 
        .CI(pe_1_6_0_sub_81_carry[2]), .CO(pe_1_6_0_sub_81_carry[3]), .S(
        pe_1_6_0_N72) );
  FA_X1 pe_1_6_0_sub_81_U2_1 ( .A(int_data_res_6__0__1_), .B(pe_1_6_0_n71), 
        .CI(pe_1_6_0_sub_81_carry[1]), .CO(pe_1_6_0_sub_81_carry[2]), .S(
        pe_1_6_0_N71) );
  FA_X1 pe_1_6_0_add_83_U1_7 ( .A(int_data_res_6__0__7_), .B(
        pe_1_6_0_int_data_3_), .CI(pe_1_6_0_add_83_carry[7]), .S(pe_1_6_0_N85)
         );
  FA_X1 pe_1_6_0_add_83_U1_6 ( .A(int_data_res_6__0__6_), .B(
        pe_1_6_0_int_data_3_), .CI(pe_1_6_0_add_83_carry[6]), .CO(
        pe_1_6_0_add_83_carry[7]), .S(pe_1_6_0_N84) );
  FA_X1 pe_1_6_0_add_83_U1_5 ( .A(int_data_res_6__0__5_), .B(
        pe_1_6_0_int_data_3_), .CI(pe_1_6_0_add_83_carry[5]), .CO(
        pe_1_6_0_add_83_carry[6]), .S(pe_1_6_0_N83) );
  FA_X1 pe_1_6_0_add_83_U1_4 ( .A(int_data_res_6__0__4_), .B(
        pe_1_6_0_int_data_3_), .CI(pe_1_6_0_add_83_carry[4]), .CO(
        pe_1_6_0_add_83_carry[5]), .S(pe_1_6_0_N82) );
  FA_X1 pe_1_6_0_add_83_U1_3 ( .A(int_data_res_6__0__3_), .B(
        pe_1_6_0_int_data_3_), .CI(pe_1_6_0_add_83_carry[3]), .CO(
        pe_1_6_0_add_83_carry[4]), .S(pe_1_6_0_N81) );
  FA_X1 pe_1_6_0_add_83_U1_2 ( .A(int_data_res_6__0__2_), .B(
        pe_1_6_0_int_data_2_), .CI(pe_1_6_0_add_83_carry[2]), .CO(
        pe_1_6_0_add_83_carry[3]), .S(pe_1_6_0_N80) );
  FA_X1 pe_1_6_0_add_83_U1_1 ( .A(int_data_res_6__0__1_), .B(
        pe_1_6_0_int_data_1_), .CI(pe_1_6_0_n2), .CO(pe_1_6_0_add_83_carry[2]), 
        .S(pe_1_6_0_N79) );
  NAND3_X1 pe_1_6_0_U56 ( .A1(n35), .A2(pe_1_6_0_n43), .A3(pe_1_6_0_n60), .ZN(
        pe_1_6_0_n40) );
  NAND3_X1 pe_1_6_0_U55 ( .A1(pe_1_6_0_n43), .A2(pe_1_6_0_n59), .A3(
        pe_1_6_0_n60), .ZN(pe_1_6_0_n39) );
  NAND3_X1 pe_1_6_0_U54 ( .A1(pe_1_6_0_n43), .A2(pe_1_6_0_n61), .A3(n35), .ZN(
        pe_1_6_0_n38) );
  NAND3_X1 pe_1_6_0_U53 ( .A1(pe_1_6_0_n59), .A2(pe_1_6_0_n61), .A3(
        pe_1_6_0_n43), .ZN(pe_1_6_0_n37) );
  DFFR_X1 pe_1_6_0_int_q_acc_reg_6_ ( .D(pe_1_6_0_n75), .CK(pe_1_6_0_net3808), 
        .RN(pe_1_6_0_n68), .Q(int_data_res_6__0__6_) );
  DFFR_X1 pe_1_6_0_int_q_acc_reg_5_ ( .D(pe_1_6_0_n76), .CK(pe_1_6_0_net3808), 
        .RN(pe_1_6_0_n68), .Q(int_data_res_6__0__5_) );
  DFFR_X1 pe_1_6_0_int_q_acc_reg_4_ ( .D(pe_1_6_0_n77), .CK(pe_1_6_0_net3808), 
        .RN(pe_1_6_0_n68), .Q(int_data_res_6__0__4_) );
  DFFR_X1 pe_1_6_0_int_q_acc_reg_3_ ( .D(pe_1_6_0_n78), .CK(pe_1_6_0_net3808), 
        .RN(pe_1_6_0_n68), .Q(int_data_res_6__0__3_) );
  DFFR_X1 pe_1_6_0_int_q_acc_reg_2_ ( .D(pe_1_6_0_n79), .CK(pe_1_6_0_net3808), 
        .RN(pe_1_6_0_n68), .Q(int_data_res_6__0__2_) );
  DFFR_X1 pe_1_6_0_int_q_acc_reg_1_ ( .D(pe_1_6_0_n80), .CK(pe_1_6_0_net3808), 
        .RN(pe_1_6_0_n68), .Q(int_data_res_6__0__1_) );
  DFFR_X1 pe_1_6_0_int_q_acc_reg_7_ ( .D(pe_1_6_0_n74), .CK(pe_1_6_0_net3808), 
        .RN(pe_1_6_0_n68), .Q(int_data_res_6__0__7_) );
  CLKGATETST_X1 pe_1_6_0_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_6_0_n85), .SE(1'b0), .GCK(pe_1_6_0_net3747) );
  CLKGATETST_X1 pe_1_6_0_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_6_0_n84), .SE(1'b0), .GCK(pe_1_6_0_net3753) );
  CLKGATETST_X1 pe_1_6_0_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_6_0_n83), .SE(1'b0), .GCK(pe_1_6_0_net3758) );
  CLKGATETST_X1 pe_1_6_0_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_6_0_n82), .SE(1'b0), .GCK(pe_1_6_0_net3763) );
  CLKGATETST_X1 pe_1_6_0_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_6_0_n87), .SE(1'b0), .GCK(pe_1_6_0_net3768) );
  CLKGATETST_X1 pe_1_6_0_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_6_0_n86), .SE(1'b0), .GCK(pe_1_6_0_net3773) );
  CLKGATETST_X1 pe_1_6_0_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_6_0_N64), .SE(1'b0), .GCK(pe_1_6_0_net3778) );
  CLKGATETST_X1 pe_1_6_0_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_6_0_N63), .SE(1'b0), .GCK(pe_1_6_0_net3783) );
  CLKGATETST_X1 pe_1_6_0_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_6_0_N62), .SE(1'b0), .GCK(pe_1_6_0_net3788) );
  CLKGATETST_X1 pe_1_6_0_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_6_0_N61), .SE(1'b0), .GCK(pe_1_6_0_net3793) );
  CLKGATETST_X1 pe_1_6_0_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_6_0_N60), .SE(1'b0), .GCK(pe_1_6_0_net3798) );
  CLKGATETST_X1 pe_1_6_0_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_6_0_N59), .SE(1'b0), .GCK(pe_1_6_0_net3803) );
  CLKGATETST_X1 pe_1_6_0_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_6_0_N90), .SE(1'b0), .GCK(pe_1_6_0_net3808) );
  CLKBUF_X1 pe_1_6_1_U108 ( .A(pe_1_6_1_n68), .Z(pe_1_6_1_n67) );
  INV_X1 pe_1_6_1_U107 ( .A(n77), .ZN(pe_1_6_1_n66) );
  INV_X1 pe_1_6_1_U106 ( .A(n69), .ZN(pe_1_6_1_n65) );
  INV_X1 pe_1_6_1_U105 ( .A(n69), .ZN(pe_1_6_1_n64) );
  INV_X1 pe_1_6_1_U104 ( .A(pe_1_6_1_n65), .ZN(pe_1_6_1_n63) );
  INV_X1 pe_1_6_1_U103 ( .A(n29), .ZN(pe_1_6_1_n58) );
  INV_X1 pe_1_6_1_U102 ( .A(n21), .ZN(pe_1_6_1_n57) );
  MUX2_X1 pe_1_6_1_U101 ( .A(pe_1_6_1_n54), .B(pe_1_6_1_n51), .S(n52), .Z(
        int_data_x_6__1__3_) );
  MUX2_X1 pe_1_6_1_U100 ( .A(pe_1_6_1_n53), .B(pe_1_6_1_n52), .S(n41), .Z(
        pe_1_6_1_n54) );
  MUX2_X1 pe_1_6_1_U99 ( .A(pe_1_6_1_int_q_reg_h[23]), .B(
        pe_1_6_1_int_q_reg_h[19]), .S(pe_1_6_1_n56), .Z(pe_1_6_1_n53) );
  MUX2_X1 pe_1_6_1_U98 ( .A(pe_1_6_1_int_q_reg_h[15]), .B(
        pe_1_6_1_int_q_reg_h[11]), .S(pe_1_6_1_n56), .Z(pe_1_6_1_n52) );
  MUX2_X1 pe_1_6_1_U97 ( .A(pe_1_6_1_int_q_reg_h[7]), .B(
        pe_1_6_1_int_q_reg_h[3]), .S(pe_1_6_1_n56), .Z(pe_1_6_1_n51) );
  MUX2_X1 pe_1_6_1_U96 ( .A(pe_1_6_1_n50), .B(pe_1_6_1_n47), .S(n52), .Z(
        int_data_x_6__1__2_) );
  MUX2_X1 pe_1_6_1_U95 ( .A(pe_1_6_1_n49), .B(pe_1_6_1_n48), .S(n41), .Z(
        pe_1_6_1_n50) );
  MUX2_X1 pe_1_6_1_U94 ( .A(pe_1_6_1_int_q_reg_h[22]), .B(
        pe_1_6_1_int_q_reg_h[18]), .S(pe_1_6_1_n56), .Z(pe_1_6_1_n49) );
  MUX2_X1 pe_1_6_1_U93 ( .A(pe_1_6_1_int_q_reg_h[14]), .B(
        pe_1_6_1_int_q_reg_h[10]), .S(pe_1_6_1_n56), .Z(pe_1_6_1_n48) );
  MUX2_X1 pe_1_6_1_U92 ( .A(pe_1_6_1_int_q_reg_h[6]), .B(
        pe_1_6_1_int_q_reg_h[2]), .S(pe_1_6_1_n56), .Z(pe_1_6_1_n47) );
  MUX2_X1 pe_1_6_1_U91 ( .A(pe_1_6_1_n46), .B(pe_1_6_1_n24), .S(n52), .Z(
        int_data_x_6__1__1_) );
  MUX2_X1 pe_1_6_1_U90 ( .A(pe_1_6_1_n45), .B(pe_1_6_1_n25), .S(n41), .Z(
        pe_1_6_1_n46) );
  MUX2_X1 pe_1_6_1_U89 ( .A(pe_1_6_1_int_q_reg_h[21]), .B(
        pe_1_6_1_int_q_reg_h[17]), .S(pe_1_6_1_n56), .Z(pe_1_6_1_n45) );
  MUX2_X1 pe_1_6_1_U88 ( .A(pe_1_6_1_int_q_reg_h[13]), .B(
        pe_1_6_1_int_q_reg_h[9]), .S(pe_1_6_1_n56), .Z(pe_1_6_1_n25) );
  MUX2_X1 pe_1_6_1_U87 ( .A(pe_1_6_1_int_q_reg_h[5]), .B(
        pe_1_6_1_int_q_reg_h[1]), .S(pe_1_6_1_n56), .Z(pe_1_6_1_n24) );
  MUX2_X1 pe_1_6_1_U86 ( .A(pe_1_6_1_n23), .B(pe_1_6_1_n20), .S(n52), .Z(
        int_data_x_6__1__0_) );
  MUX2_X1 pe_1_6_1_U85 ( .A(pe_1_6_1_n22), .B(pe_1_6_1_n21), .S(n41), .Z(
        pe_1_6_1_n23) );
  MUX2_X1 pe_1_6_1_U84 ( .A(pe_1_6_1_int_q_reg_h[20]), .B(
        pe_1_6_1_int_q_reg_h[16]), .S(pe_1_6_1_n56), .Z(pe_1_6_1_n22) );
  MUX2_X1 pe_1_6_1_U83 ( .A(pe_1_6_1_int_q_reg_h[12]), .B(
        pe_1_6_1_int_q_reg_h[8]), .S(pe_1_6_1_n56), .Z(pe_1_6_1_n21) );
  MUX2_X1 pe_1_6_1_U82 ( .A(pe_1_6_1_int_q_reg_h[4]), .B(
        pe_1_6_1_int_q_reg_h[0]), .S(pe_1_6_1_n56), .Z(pe_1_6_1_n20) );
  MUX2_X1 pe_1_6_1_U81 ( .A(pe_1_6_1_n19), .B(pe_1_6_1_n16), .S(n52), .Z(
        int_data_y_6__1__3_) );
  MUX2_X1 pe_1_6_1_U80 ( .A(pe_1_6_1_n18), .B(pe_1_6_1_n17), .S(n41), .Z(
        pe_1_6_1_n19) );
  MUX2_X1 pe_1_6_1_U79 ( .A(pe_1_6_1_int_q_reg_v[23]), .B(
        pe_1_6_1_int_q_reg_v[19]), .S(pe_1_6_1_n55), .Z(pe_1_6_1_n18) );
  MUX2_X1 pe_1_6_1_U78 ( .A(pe_1_6_1_int_q_reg_v[15]), .B(
        pe_1_6_1_int_q_reg_v[11]), .S(pe_1_6_1_n55), .Z(pe_1_6_1_n17) );
  MUX2_X1 pe_1_6_1_U77 ( .A(pe_1_6_1_int_q_reg_v[7]), .B(
        pe_1_6_1_int_q_reg_v[3]), .S(pe_1_6_1_n55), .Z(pe_1_6_1_n16) );
  MUX2_X1 pe_1_6_1_U76 ( .A(pe_1_6_1_n15), .B(pe_1_6_1_n12), .S(n52), .Z(
        int_data_y_6__1__2_) );
  MUX2_X1 pe_1_6_1_U75 ( .A(pe_1_6_1_n14), .B(pe_1_6_1_n13), .S(n41), .Z(
        pe_1_6_1_n15) );
  MUX2_X1 pe_1_6_1_U74 ( .A(pe_1_6_1_int_q_reg_v[22]), .B(
        pe_1_6_1_int_q_reg_v[18]), .S(pe_1_6_1_n55), .Z(pe_1_6_1_n14) );
  MUX2_X1 pe_1_6_1_U73 ( .A(pe_1_6_1_int_q_reg_v[14]), .B(
        pe_1_6_1_int_q_reg_v[10]), .S(pe_1_6_1_n55), .Z(pe_1_6_1_n13) );
  MUX2_X1 pe_1_6_1_U72 ( .A(pe_1_6_1_int_q_reg_v[6]), .B(
        pe_1_6_1_int_q_reg_v[2]), .S(pe_1_6_1_n55), .Z(pe_1_6_1_n12) );
  MUX2_X1 pe_1_6_1_U71 ( .A(pe_1_6_1_n11), .B(pe_1_6_1_n8), .S(n52), .Z(
        int_data_y_6__1__1_) );
  MUX2_X1 pe_1_6_1_U70 ( .A(pe_1_6_1_n10), .B(pe_1_6_1_n9), .S(n41), .Z(
        pe_1_6_1_n11) );
  MUX2_X1 pe_1_6_1_U69 ( .A(pe_1_6_1_int_q_reg_v[21]), .B(
        pe_1_6_1_int_q_reg_v[17]), .S(pe_1_6_1_n55), .Z(pe_1_6_1_n10) );
  MUX2_X1 pe_1_6_1_U68 ( .A(pe_1_6_1_int_q_reg_v[13]), .B(
        pe_1_6_1_int_q_reg_v[9]), .S(pe_1_6_1_n55), .Z(pe_1_6_1_n9) );
  MUX2_X1 pe_1_6_1_U67 ( .A(pe_1_6_1_int_q_reg_v[5]), .B(
        pe_1_6_1_int_q_reg_v[1]), .S(pe_1_6_1_n55), .Z(pe_1_6_1_n8) );
  MUX2_X1 pe_1_6_1_U66 ( .A(pe_1_6_1_n7), .B(pe_1_6_1_n4), .S(n52), .Z(
        int_data_y_6__1__0_) );
  MUX2_X1 pe_1_6_1_U65 ( .A(pe_1_6_1_n6), .B(pe_1_6_1_n5), .S(n41), .Z(
        pe_1_6_1_n7) );
  MUX2_X1 pe_1_6_1_U64 ( .A(pe_1_6_1_int_q_reg_v[20]), .B(
        pe_1_6_1_int_q_reg_v[16]), .S(pe_1_6_1_n55), .Z(pe_1_6_1_n6) );
  MUX2_X1 pe_1_6_1_U63 ( .A(pe_1_6_1_int_q_reg_v[12]), .B(
        pe_1_6_1_int_q_reg_v[8]), .S(pe_1_6_1_n55), .Z(pe_1_6_1_n5) );
  MUX2_X1 pe_1_6_1_U62 ( .A(pe_1_6_1_int_q_reg_v[4]), .B(
        pe_1_6_1_int_q_reg_v[0]), .S(pe_1_6_1_n55), .Z(pe_1_6_1_n4) );
  AOI222_X1 pe_1_6_1_U61 ( .A1(int_data_res_7__1__2_), .A2(pe_1_6_1_n61), .B1(
        pe_1_6_1_N80), .B2(pe_1_6_1_n27), .C1(pe_1_6_1_N72), .C2(pe_1_6_1_n28), 
        .ZN(pe_1_6_1_n33) );
  INV_X1 pe_1_6_1_U60 ( .A(pe_1_6_1_n33), .ZN(pe_1_6_1_n78) );
  AOI222_X1 pe_1_6_1_U59 ( .A1(int_data_res_7__1__6_), .A2(pe_1_6_1_n61), .B1(
        pe_1_6_1_N84), .B2(pe_1_6_1_n27), .C1(pe_1_6_1_N76), .C2(pe_1_6_1_n28), 
        .ZN(pe_1_6_1_n29) );
  INV_X1 pe_1_6_1_U58 ( .A(pe_1_6_1_n29), .ZN(pe_1_6_1_n74) );
  XNOR2_X1 pe_1_6_1_U57 ( .A(pe_1_6_1_n69), .B(int_data_res_6__1__0_), .ZN(
        pe_1_6_1_N70) );
  AOI222_X1 pe_1_6_1_U52 ( .A1(int_data_res_7__1__0_), .A2(pe_1_6_1_n61), .B1(
        pe_1_6_1_n1), .B2(pe_1_6_1_n27), .C1(pe_1_6_1_N70), .C2(pe_1_6_1_n28), 
        .ZN(pe_1_6_1_n35) );
  INV_X1 pe_1_6_1_U51 ( .A(pe_1_6_1_n35), .ZN(pe_1_6_1_n80) );
  AOI222_X1 pe_1_6_1_U50 ( .A1(int_data_res_7__1__1_), .A2(pe_1_6_1_n61), .B1(
        pe_1_6_1_N79), .B2(pe_1_6_1_n27), .C1(pe_1_6_1_N71), .C2(pe_1_6_1_n28), 
        .ZN(pe_1_6_1_n34) );
  INV_X1 pe_1_6_1_U49 ( .A(pe_1_6_1_n34), .ZN(pe_1_6_1_n79) );
  AOI222_X1 pe_1_6_1_U48 ( .A1(int_data_res_7__1__3_), .A2(pe_1_6_1_n61), .B1(
        pe_1_6_1_N81), .B2(pe_1_6_1_n27), .C1(pe_1_6_1_N73), .C2(pe_1_6_1_n28), 
        .ZN(pe_1_6_1_n32) );
  INV_X1 pe_1_6_1_U47 ( .A(pe_1_6_1_n32), .ZN(pe_1_6_1_n77) );
  AOI222_X1 pe_1_6_1_U46 ( .A1(int_data_res_7__1__4_), .A2(pe_1_6_1_n61), .B1(
        pe_1_6_1_N82), .B2(pe_1_6_1_n27), .C1(pe_1_6_1_N74), .C2(pe_1_6_1_n28), 
        .ZN(pe_1_6_1_n31) );
  INV_X1 pe_1_6_1_U45 ( .A(pe_1_6_1_n31), .ZN(pe_1_6_1_n76) );
  AOI222_X1 pe_1_6_1_U44 ( .A1(int_data_res_7__1__5_), .A2(pe_1_6_1_n61), .B1(
        pe_1_6_1_N83), .B2(pe_1_6_1_n27), .C1(pe_1_6_1_N75), .C2(pe_1_6_1_n28), 
        .ZN(pe_1_6_1_n30) );
  INV_X1 pe_1_6_1_U43 ( .A(pe_1_6_1_n30), .ZN(pe_1_6_1_n75) );
  NAND2_X1 pe_1_6_1_U42 ( .A1(pe_1_6_1_int_data_0_), .A2(pe_1_6_1_n3), .ZN(
        pe_1_6_1_sub_81_carry[1]) );
  INV_X1 pe_1_6_1_U41 ( .A(pe_1_6_1_int_data_1_), .ZN(pe_1_6_1_n70) );
  INV_X1 pe_1_6_1_U40 ( .A(pe_1_6_1_int_data_2_), .ZN(pe_1_6_1_n71) );
  AND2_X1 pe_1_6_1_U39 ( .A1(pe_1_6_1_int_data_0_), .A2(int_data_res_6__1__0_), 
        .ZN(pe_1_6_1_n2) );
  AOI222_X1 pe_1_6_1_U38 ( .A1(pe_1_6_1_n61), .A2(int_data_res_7__1__7_), .B1(
        pe_1_6_1_N85), .B2(pe_1_6_1_n27), .C1(pe_1_6_1_N77), .C2(pe_1_6_1_n28), 
        .ZN(pe_1_6_1_n26) );
  INV_X1 pe_1_6_1_U37 ( .A(pe_1_6_1_n26), .ZN(pe_1_6_1_n73) );
  NOR3_X1 pe_1_6_1_U36 ( .A1(pe_1_6_1_n58), .A2(pe_1_6_1_n62), .A3(int_ckg[14]), .ZN(pe_1_6_1_n36) );
  OR2_X1 pe_1_6_1_U35 ( .A1(pe_1_6_1_n36), .A2(pe_1_6_1_n61), .ZN(pe_1_6_1_N90) );
  INV_X1 pe_1_6_1_U34 ( .A(n41), .ZN(pe_1_6_1_n60) );
  AND2_X1 pe_1_6_1_U33 ( .A1(int_data_x_6__1__2_), .A2(n29), .ZN(
        pe_1_6_1_int_data_2_) );
  AND2_X1 pe_1_6_1_U32 ( .A1(int_data_x_6__1__1_), .A2(n29), .ZN(
        pe_1_6_1_int_data_1_) );
  AND2_X1 pe_1_6_1_U31 ( .A1(int_data_x_6__1__3_), .A2(n29), .ZN(
        pe_1_6_1_int_data_3_) );
  BUF_X1 pe_1_6_1_U30 ( .A(n63), .Z(pe_1_6_1_n61) );
  INV_X1 pe_1_6_1_U29 ( .A(n35), .ZN(pe_1_6_1_n59) );
  AND2_X1 pe_1_6_1_U28 ( .A1(int_data_x_6__1__0_), .A2(n29), .ZN(
        pe_1_6_1_int_data_0_) );
  NAND2_X1 pe_1_6_1_U27 ( .A1(pe_1_6_1_n44), .A2(pe_1_6_1_n59), .ZN(
        pe_1_6_1_n41) );
  AND3_X1 pe_1_6_1_U26 ( .A1(n77), .A2(pe_1_6_1_n60), .A3(n52), .ZN(
        pe_1_6_1_n44) );
  INV_X1 pe_1_6_1_U25 ( .A(pe_1_6_1_int_data_3_), .ZN(pe_1_6_1_n72) );
  NOR2_X1 pe_1_6_1_U24 ( .A1(pe_1_6_1_n66), .A2(n52), .ZN(pe_1_6_1_n43) );
  NOR2_X1 pe_1_6_1_U23 ( .A1(pe_1_6_1_n57), .A2(pe_1_6_1_n61), .ZN(
        pe_1_6_1_n28) );
  NOR2_X1 pe_1_6_1_U22 ( .A1(n21), .A2(pe_1_6_1_n61), .ZN(pe_1_6_1_n27) );
  INV_X1 pe_1_6_1_U21 ( .A(pe_1_6_1_int_data_0_), .ZN(pe_1_6_1_n69) );
  INV_X1 pe_1_6_1_U20 ( .A(pe_1_6_1_n41), .ZN(pe_1_6_1_n86) );
  INV_X1 pe_1_6_1_U19 ( .A(pe_1_6_1_n37), .ZN(pe_1_6_1_n84) );
  INV_X1 pe_1_6_1_U18 ( .A(pe_1_6_1_n38), .ZN(pe_1_6_1_n83) );
  INV_X1 pe_1_6_1_U17 ( .A(pe_1_6_1_n39), .ZN(pe_1_6_1_n82) );
  NOR2_X1 pe_1_6_1_U16 ( .A1(pe_1_6_1_n64), .A2(pe_1_6_1_n42), .ZN(
        pe_1_6_1_N59) );
  NOR2_X1 pe_1_6_1_U15 ( .A1(pe_1_6_1_n64), .A2(pe_1_6_1_n41), .ZN(
        pe_1_6_1_N60) );
  NOR2_X1 pe_1_6_1_U14 ( .A1(pe_1_6_1_n64), .A2(pe_1_6_1_n38), .ZN(
        pe_1_6_1_N63) );
  NOR2_X1 pe_1_6_1_U13 ( .A1(pe_1_6_1_n64), .A2(pe_1_6_1_n40), .ZN(
        pe_1_6_1_N61) );
  NOR2_X1 pe_1_6_1_U12 ( .A1(pe_1_6_1_n64), .A2(pe_1_6_1_n39), .ZN(
        pe_1_6_1_N62) );
  NOR2_X1 pe_1_6_1_U11 ( .A1(pe_1_6_1_n37), .A2(pe_1_6_1_n64), .ZN(
        pe_1_6_1_N64) );
  NAND2_X1 pe_1_6_1_U10 ( .A1(pe_1_6_1_n44), .A2(n35), .ZN(pe_1_6_1_n42) );
  BUF_X1 pe_1_6_1_U9 ( .A(n35), .Z(pe_1_6_1_n55) );
  INV_X1 pe_1_6_1_U8 ( .A(pe_1_6_1_n65), .ZN(pe_1_6_1_n62) );
  BUF_X1 pe_1_6_1_U7 ( .A(n35), .Z(pe_1_6_1_n56) );
  INV_X1 pe_1_6_1_U6 ( .A(pe_1_6_1_n42), .ZN(pe_1_6_1_n85) );
  INV_X1 pe_1_6_1_U5 ( .A(pe_1_6_1_n40), .ZN(pe_1_6_1_n81) );
  INV_X2 pe_1_6_1_U4 ( .A(n85), .ZN(pe_1_6_1_n68) );
  XOR2_X1 pe_1_6_1_U3 ( .A(pe_1_6_1_int_data_0_), .B(int_data_res_6__1__0_), 
        .Z(pe_1_6_1_n1) );
  DFFR_X1 pe_1_6_1_int_q_acc_reg_0_ ( .D(pe_1_6_1_n80), .CK(pe_1_6_1_net3730), 
        .RN(pe_1_6_1_n68), .Q(int_data_res_6__1__0_), .QN(pe_1_6_1_n3) );
  DFFR_X1 pe_1_6_1_int_q_reg_v_reg_0__0_ ( .D(int_data_y_7__1__0_), .CK(
        pe_1_6_1_net3700), .RN(pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_v[20]) );
  DFFR_X1 pe_1_6_1_int_q_reg_v_reg_0__1_ ( .D(int_data_y_7__1__1_), .CK(
        pe_1_6_1_net3700), .RN(pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_v[21]) );
  DFFR_X1 pe_1_6_1_int_q_reg_v_reg_0__2_ ( .D(int_data_y_7__1__2_), .CK(
        pe_1_6_1_net3700), .RN(pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_v[22]) );
  DFFR_X1 pe_1_6_1_int_q_reg_v_reg_0__3_ ( .D(int_data_y_7__1__3_), .CK(
        pe_1_6_1_net3700), .RN(pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_v[23]) );
  DFFR_X1 pe_1_6_1_int_q_reg_v_reg_1__0_ ( .D(int_data_y_7__1__0_), .CK(
        pe_1_6_1_net3705), .RN(pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_v[16]) );
  DFFR_X1 pe_1_6_1_int_q_reg_v_reg_1__1_ ( .D(int_data_y_7__1__1_), .CK(
        pe_1_6_1_net3705), .RN(pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_v[17]) );
  DFFR_X1 pe_1_6_1_int_q_reg_v_reg_1__2_ ( .D(int_data_y_7__1__2_), .CK(
        pe_1_6_1_net3705), .RN(pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_v[18]) );
  DFFR_X1 pe_1_6_1_int_q_reg_v_reg_1__3_ ( .D(int_data_y_7__1__3_), .CK(
        pe_1_6_1_net3705), .RN(pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_v[19]) );
  DFFR_X1 pe_1_6_1_int_q_reg_v_reg_2__0_ ( .D(int_data_y_7__1__0_), .CK(
        pe_1_6_1_net3710), .RN(pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_v[12]) );
  DFFR_X1 pe_1_6_1_int_q_reg_v_reg_2__1_ ( .D(int_data_y_7__1__1_), .CK(
        pe_1_6_1_net3710), .RN(pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_v[13]) );
  DFFR_X1 pe_1_6_1_int_q_reg_v_reg_2__2_ ( .D(int_data_y_7__1__2_), .CK(
        pe_1_6_1_net3710), .RN(pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_v[14]) );
  DFFR_X1 pe_1_6_1_int_q_reg_v_reg_2__3_ ( .D(int_data_y_7__1__3_), .CK(
        pe_1_6_1_net3710), .RN(pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_v[15]) );
  DFFR_X1 pe_1_6_1_int_q_reg_v_reg_3__0_ ( .D(int_data_y_7__1__0_), .CK(
        pe_1_6_1_net3715), .RN(pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_v[8]) );
  DFFR_X1 pe_1_6_1_int_q_reg_v_reg_3__1_ ( .D(int_data_y_7__1__1_), .CK(
        pe_1_6_1_net3715), .RN(pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_v[9]) );
  DFFR_X1 pe_1_6_1_int_q_reg_v_reg_3__2_ ( .D(int_data_y_7__1__2_), .CK(
        pe_1_6_1_net3715), .RN(pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_v[10]) );
  DFFR_X1 pe_1_6_1_int_q_reg_v_reg_3__3_ ( .D(int_data_y_7__1__3_), .CK(
        pe_1_6_1_net3715), .RN(pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_v[11]) );
  DFFR_X1 pe_1_6_1_int_q_reg_v_reg_4__0_ ( .D(int_data_y_7__1__0_), .CK(
        pe_1_6_1_net3720), .RN(pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_v[4]) );
  DFFR_X1 pe_1_6_1_int_q_reg_v_reg_4__1_ ( .D(int_data_y_7__1__1_), .CK(
        pe_1_6_1_net3720), .RN(pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_v[5]) );
  DFFR_X1 pe_1_6_1_int_q_reg_v_reg_4__2_ ( .D(int_data_y_7__1__2_), .CK(
        pe_1_6_1_net3720), .RN(pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_v[6]) );
  DFFR_X1 pe_1_6_1_int_q_reg_v_reg_4__3_ ( .D(int_data_y_7__1__3_), .CK(
        pe_1_6_1_net3720), .RN(pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_v[7]) );
  DFFR_X1 pe_1_6_1_int_q_reg_v_reg_5__0_ ( .D(int_data_y_7__1__0_), .CK(
        pe_1_6_1_net3725), .RN(pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_v[0]) );
  DFFR_X1 pe_1_6_1_int_q_reg_v_reg_5__1_ ( .D(int_data_y_7__1__1_), .CK(
        pe_1_6_1_net3725), .RN(pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_v[1]) );
  DFFR_X1 pe_1_6_1_int_q_reg_v_reg_5__2_ ( .D(int_data_y_7__1__2_), .CK(
        pe_1_6_1_net3725), .RN(pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_v[2]) );
  DFFR_X1 pe_1_6_1_int_q_reg_v_reg_5__3_ ( .D(int_data_y_7__1__3_), .CK(
        pe_1_6_1_net3725), .RN(pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_6_1_int_q_reg_h_reg_0__0_ ( .D(int_data_x_6__2__0_), .SI(
        int_data_y_7__1__0_), .SE(pe_1_6_1_n62), .CK(pe_1_6_1_net3669), .RN(
        pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_6_1_int_q_reg_h_reg_0__1_ ( .D(int_data_x_6__2__1_), .SI(
        int_data_y_7__1__1_), .SE(pe_1_6_1_n62), .CK(pe_1_6_1_net3669), .RN(
        pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_6_1_int_q_reg_h_reg_0__2_ ( .D(int_data_x_6__2__2_), .SI(
        int_data_y_7__1__2_), .SE(pe_1_6_1_n62), .CK(pe_1_6_1_net3669), .RN(
        pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_6_1_int_q_reg_h_reg_0__3_ ( .D(int_data_x_6__2__3_), .SI(
        int_data_y_7__1__3_), .SE(pe_1_6_1_n62), .CK(pe_1_6_1_net3669), .RN(
        pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_6_1_int_q_reg_h_reg_1__0_ ( .D(int_data_x_6__2__0_), .SI(
        int_data_y_7__1__0_), .SE(pe_1_6_1_n62), .CK(pe_1_6_1_net3675), .RN(
        pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_6_1_int_q_reg_h_reg_1__1_ ( .D(int_data_x_6__2__1_), .SI(
        int_data_y_7__1__1_), .SE(pe_1_6_1_n62), .CK(pe_1_6_1_net3675), .RN(
        pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_6_1_int_q_reg_h_reg_1__2_ ( .D(int_data_x_6__2__2_), .SI(
        int_data_y_7__1__2_), .SE(pe_1_6_1_n62), .CK(pe_1_6_1_net3675), .RN(
        pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_6_1_int_q_reg_h_reg_1__3_ ( .D(int_data_x_6__2__3_), .SI(
        int_data_y_7__1__3_), .SE(pe_1_6_1_n62), .CK(pe_1_6_1_net3675), .RN(
        pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_6_1_int_q_reg_h_reg_2__0_ ( .D(int_data_x_6__2__0_), .SI(
        int_data_y_7__1__0_), .SE(pe_1_6_1_n62), .CK(pe_1_6_1_net3680), .RN(
        pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_6_1_int_q_reg_h_reg_2__1_ ( .D(int_data_x_6__2__1_), .SI(
        int_data_y_7__1__1_), .SE(pe_1_6_1_n62), .CK(pe_1_6_1_net3680), .RN(
        pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_6_1_int_q_reg_h_reg_2__2_ ( .D(int_data_x_6__2__2_), .SI(
        int_data_y_7__1__2_), .SE(pe_1_6_1_n62), .CK(pe_1_6_1_net3680), .RN(
        pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_6_1_int_q_reg_h_reg_2__3_ ( .D(int_data_x_6__2__3_), .SI(
        int_data_y_7__1__3_), .SE(pe_1_6_1_n62), .CK(pe_1_6_1_net3680), .RN(
        pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_6_1_int_q_reg_h_reg_3__0_ ( .D(int_data_x_6__2__0_), .SI(
        int_data_y_7__1__0_), .SE(pe_1_6_1_n62), .CK(pe_1_6_1_net3685), .RN(
        pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_6_1_int_q_reg_h_reg_3__1_ ( .D(int_data_x_6__2__1_), .SI(
        int_data_y_7__1__1_), .SE(pe_1_6_1_n62), .CK(pe_1_6_1_net3685), .RN(
        pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_6_1_int_q_reg_h_reg_3__2_ ( .D(int_data_x_6__2__2_), .SI(
        int_data_y_7__1__2_), .SE(pe_1_6_1_n62), .CK(pe_1_6_1_net3685), .RN(
        pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_6_1_int_q_reg_h_reg_3__3_ ( .D(int_data_x_6__2__3_), .SI(
        int_data_y_7__1__3_), .SE(pe_1_6_1_n62), .CK(pe_1_6_1_net3685), .RN(
        pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_6_1_int_q_reg_h_reg_4__0_ ( .D(int_data_x_6__2__0_), .SI(
        int_data_y_7__1__0_), .SE(pe_1_6_1_n63), .CK(pe_1_6_1_net3690), .RN(
        pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_6_1_int_q_reg_h_reg_4__1_ ( .D(int_data_x_6__2__1_), .SI(
        int_data_y_7__1__1_), .SE(pe_1_6_1_n63), .CK(pe_1_6_1_net3690), .RN(
        pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_6_1_int_q_reg_h_reg_4__2_ ( .D(int_data_x_6__2__2_), .SI(
        int_data_y_7__1__2_), .SE(pe_1_6_1_n63), .CK(pe_1_6_1_net3690), .RN(
        pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_6_1_int_q_reg_h_reg_4__3_ ( .D(int_data_x_6__2__3_), .SI(
        int_data_y_7__1__3_), .SE(pe_1_6_1_n63), .CK(pe_1_6_1_net3690), .RN(
        pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_6_1_int_q_reg_h_reg_5__0_ ( .D(int_data_x_6__2__0_), .SI(
        int_data_y_7__1__0_), .SE(pe_1_6_1_n63), .CK(pe_1_6_1_net3695), .RN(
        pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_6_1_int_q_reg_h_reg_5__1_ ( .D(int_data_x_6__2__1_), .SI(
        int_data_y_7__1__1_), .SE(pe_1_6_1_n63), .CK(pe_1_6_1_net3695), .RN(
        pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_6_1_int_q_reg_h_reg_5__2_ ( .D(int_data_x_6__2__2_), .SI(
        int_data_y_7__1__2_), .SE(pe_1_6_1_n63), .CK(pe_1_6_1_net3695), .RN(
        pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_6_1_int_q_reg_h_reg_5__3_ ( .D(int_data_x_6__2__3_), .SI(
        int_data_y_7__1__3_), .SE(pe_1_6_1_n63), .CK(pe_1_6_1_net3695), .RN(
        pe_1_6_1_n68), .Q(pe_1_6_1_int_q_reg_h[3]) );
  FA_X1 pe_1_6_1_sub_81_U2_7 ( .A(int_data_res_6__1__7_), .B(pe_1_6_1_n72), 
        .CI(pe_1_6_1_sub_81_carry[7]), .S(pe_1_6_1_N77) );
  FA_X1 pe_1_6_1_sub_81_U2_6 ( .A(int_data_res_6__1__6_), .B(pe_1_6_1_n72), 
        .CI(pe_1_6_1_sub_81_carry[6]), .CO(pe_1_6_1_sub_81_carry[7]), .S(
        pe_1_6_1_N76) );
  FA_X1 pe_1_6_1_sub_81_U2_5 ( .A(int_data_res_6__1__5_), .B(pe_1_6_1_n72), 
        .CI(pe_1_6_1_sub_81_carry[5]), .CO(pe_1_6_1_sub_81_carry[6]), .S(
        pe_1_6_1_N75) );
  FA_X1 pe_1_6_1_sub_81_U2_4 ( .A(int_data_res_6__1__4_), .B(pe_1_6_1_n72), 
        .CI(pe_1_6_1_sub_81_carry[4]), .CO(pe_1_6_1_sub_81_carry[5]), .S(
        pe_1_6_1_N74) );
  FA_X1 pe_1_6_1_sub_81_U2_3 ( .A(int_data_res_6__1__3_), .B(pe_1_6_1_n72), 
        .CI(pe_1_6_1_sub_81_carry[3]), .CO(pe_1_6_1_sub_81_carry[4]), .S(
        pe_1_6_1_N73) );
  FA_X1 pe_1_6_1_sub_81_U2_2 ( .A(int_data_res_6__1__2_), .B(pe_1_6_1_n71), 
        .CI(pe_1_6_1_sub_81_carry[2]), .CO(pe_1_6_1_sub_81_carry[3]), .S(
        pe_1_6_1_N72) );
  FA_X1 pe_1_6_1_sub_81_U2_1 ( .A(int_data_res_6__1__1_), .B(pe_1_6_1_n70), 
        .CI(pe_1_6_1_sub_81_carry[1]), .CO(pe_1_6_1_sub_81_carry[2]), .S(
        pe_1_6_1_N71) );
  FA_X1 pe_1_6_1_add_83_U1_7 ( .A(int_data_res_6__1__7_), .B(
        pe_1_6_1_int_data_3_), .CI(pe_1_6_1_add_83_carry[7]), .S(pe_1_6_1_N85)
         );
  FA_X1 pe_1_6_1_add_83_U1_6 ( .A(int_data_res_6__1__6_), .B(
        pe_1_6_1_int_data_3_), .CI(pe_1_6_1_add_83_carry[6]), .CO(
        pe_1_6_1_add_83_carry[7]), .S(pe_1_6_1_N84) );
  FA_X1 pe_1_6_1_add_83_U1_5 ( .A(int_data_res_6__1__5_), .B(
        pe_1_6_1_int_data_3_), .CI(pe_1_6_1_add_83_carry[5]), .CO(
        pe_1_6_1_add_83_carry[6]), .S(pe_1_6_1_N83) );
  FA_X1 pe_1_6_1_add_83_U1_4 ( .A(int_data_res_6__1__4_), .B(
        pe_1_6_1_int_data_3_), .CI(pe_1_6_1_add_83_carry[4]), .CO(
        pe_1_6_1_add_83_carry[5]), .S(pe_1_6_1_N82) );
  FA_X1 pe_1_6_1_add_83_U1_3 ( .A(int_data_res_6__1__3_), .B(
        pe_1_6_1_int_data_3_), .CI(pe_1_6_1_add_83_carry[3]), .CO(
        pe_1_6_1_add_83_carry[4]), .S(pe_1_6_1_N81) );
  FA_X1 pe_1_6_1_add_83_U1_2 ( .A(int_data_res_6__1__2_), .B(
        pe_1_6_1_int_data_2_), .CI(pe_1_6_1_add_83_carry[2]), .CO(
        pe_1_6_1_add_83_carry[3]), .S(pe_1_6_1_N80) );
  FA_X1 pe_1_6_1_add_83_U1_1 ( .A(int_data_res_6__1__1_), .B(
        pe_1_6_1_int_data_1_), .CI(pe_1_6_1_n2), .CO(pe_1_6_1_add_83_carry[2]), 
        .S(pe_1_6_1_N79) );
  NAND3_X1 pe_1_6_1_U56 ( .A1(n35), .A2(pe_1_6_1_n43), .A3(n41), .ZN(
        pe_1_6_1_n40) );
  NAND3_X1 pe_1_6_1_U55 ( .A1(pe_1_6_1_n43), .A2(pe_1_6_1_n59), .A3(n41), .ZN(
        pe_1_6_1_n39) );
  NAND3_X1 pe_1_6_1_U54 ( .A1(pe_1_6_1_n43), .A2(pe_1_6_1_n60), .A3(n35), .ZN(
        pe_1_6_1_n38) );
  NAND3_X1 pe_1_6_1_U53 ( .A1(pe_1_6_1_n59), .A2(pe_1_6_1_n60), .A3(
        pe_1_6_1_n43), .ZN(pe_1_6_1_n37) );
  DFFR_X1 pe_1_6_1_int_q_acc_reg_6_ ( .D(pe_1_6_1_n74), .CK(pe_1_6_1_net3730), 
        .RN(pe_1_6_1_n67), .Q(int_data_res_6__1__6_) );
  DFFR_X1 pe_1_6_1_int_q_acc_reg_5_ ( .D(pe_1_6_1_n75), .CK(pe_1_6_1_net3730), 
        .RN(pe_1_6_1_n67), .Q(int_data_res_6__1__5_) );
  DFFR_X1 pe_1_6_1_int_q_acc_reg_4_ ( .D(pe_1_6_1_n76), .CK(pe_1_6_1_net3730), 
        .RN(pe_1_6_1_n67), .Q(int_data_res_6__1__4_) );
  DFFR_X1 pe_1_6_1_int_q_acc_reg_3_ ( .D(pe_1_6_1_n77), .CK(pe_1_6_1_net3730), 
        .RN(pe_1_6_1_n67), .Q(int_data_res_6__1__3_) );
  DFFR_X1 pe_1_6_1_int_q_acc_reg_2_ ( .D(pe_1_6_1_n78), .CK(pe_1_6_1_net3730), 
        .RN(pe_1_6_1_n67), .Q(int_data_res_6__1__2_) );
  DFFR_X1 pe_1_6_1_int_q_acc_reg_1_ ( .D(pe_1_6_1_n79), .CK(pe_1_6_1_net3730), 
        .RN(pe_1_6_1_n67), .Q(int_data_res_6__1__1_) );
  DFFR_X1 pe_1_6_1_int_q_acc_reg_7_ ( .D(pe_1_6_1_n73), .CK(pe_1_6_1_net3730), 
        .RN(pe_1_6_1_n67), .Q(int_data_res_6__1__7_) );
  CLKGATETST_X1 pe_1_6_1_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_6_1_n84), .SE(1'b0), .GCK(pe_1_6_1_net3669) );
  CLKGATETST_X1 pe_1_6_1_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_6_1_n83), .SE(1'b0), .GCK(pe_1_6_1_net3675) );
  CLKGATETST_X1 pe_1_6_1_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_6_1_n82), .SE(1'b0), .GCK(pe_1_6_1_net3680) );
  CLKGATETST_X1 pe_1_6_1_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_6_1_n81), .SE(1'b0), .GCK(pe_1_6_1_net3685) );
  CLKGATETST_X1 pe_1_6_1_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_6_1_n86), .SE(1'b0), .GCK(pe_1_6_1_net3690) );
  CLKGATETST_X1 pe_1_6_1_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_6_1_n85), .SE(1'b0), .GCK(pe_1_6_1_net3695) );
  CLKGATETST_X1 pe_1_6_1_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_6_1_N64), .SE(1'b0), .GCK(pe_1_6_1_net3700) );
  CLKGATETST_X1 pe_1_6_1_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_6_1_N63), .SE(1'b0), .GCK(pe_1_6_1_net3705) );
  CLKGATETST_X1 pe_1_6_1_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_6_1_N62), .SE(1'b0), .GCK(pe_1_6_1_net3710) );
  CLKGATETST_X1 pe_1_6_1_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_6_1_N61), .SE(1'b0), .GCK(pe_1_6_1_net3715) );
  CLKGATETST_X1 pe_1_6_1_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_6_1_N60), .SE(1'b0), .GCK(pe_1_6_1_net3720) );
  CLKGATETST_X1 pe_1_6_1_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_6_1_N59), .SE(1'b0), .GCK(pe_1_6_1_net3725) );
  CLKGATETST_X1 pe_1_6_1_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_6_1_N90), .SE(1'b0), .GCK(pe_1_6_1_net3730) );
  CLKBUF_X1 pe_1_6_2_U109 ( .A(pe_1_6_2_n69), .Z(pe_1_6_2_n68) );
  INV_X1 pe_1_6_2_U108 ( .A(n77), .ZN(pe_1_6_2_n67) );
  INV_X1 pe_1_6_2_U107 ( .A(n69), .ZN(pe_1_6_2_n66) );
  INV_X1 pe_1_6_2_U106 ( .A(n69), .ZN(pe_1_6_2_n65) );
  INV_X1 pe_1_6_2_U105 ( .A(pe_1_6_2_n66), .ZN(pe_1_6_2_n64) );
  INV_X1 pe_1_6_2_U104 ( .A(pe_1_6_2_n61), .ZN(pe_1_6_2_n60) );
  INV_X1 pe_1_6_2_U103 ( .A(n29), .ZN(pe_1_6_2_n58) );
  INV_X1 pe_1_6_2_U102 ( .A(n21), .ZN(pe_1_6_2_n57) );
  MUX2_X1 pe_1_6_2_U101 ( .A(pe_1_6_2_n54), .B(pe_1_6_2_n51), .S(n53), .Z(
        int_data_x_6__2__3_) );
  MUX2_X1 pe_1_6_2_U100 ( .A(pe_1_6_2_n53), .B(pe_1_6_2_n52), .S(pe_1_6_2_n60), 
        .Z(pe_1_6_2_n54) );
  MUX2_X1 pe_1_6_2_U99 ( .A(pe_1_6_2_int_q_reg_h[23]), .B(
        pe_1_6_2_int_q_reg_h[19]), .S(pe_1_6_2_n56), .Z(pe_1_6_2_n53) );
  MUX2_X1 pe_1_6_2_U98 ( .A(pe_1_6_2_int_q_reg_h[15]), .B(
        pe_1_6_2_int_q_reg_h[11]), .S(pe_1_6_2_n56), .Z(pe_1_6_2_n52) );
  MUX2_X1 pe_1_6_2_U97 ( .A(pe_1_6_2_int_q_reg_h[7]), .B(
        pe_1_6_2_int_q_reg_h[3]), .S(pe_1_6_2_n56), .Z(pe_1_6_2_n51) );
  MUX2_X1 pe_1_6_2_U96 ( .A(pe_1_6_2_n50), .B(pe_1_6_2_n47), .S(n53), .Z(
        int_data_x_6__2__2_) );
  MUX2_X1 pe_1_6_2_U95 ( .A(pe_1_6_2_n49), .B(pe_1_6_2_n48), .S(pe_1_6_2_n60), 
        .Z(pe_1_6_2_n50) );
  MUX2_X1 pe_1_6_2_U94 ( .A(pe_1_6_2_int_q_reg_h[22]), .B(
        pe_1_6_2_int_q_reg_h[18]), .S(pe_1_6_2_n56), .Z(pe_1_6_2_n49) );
  MUX2_X1 pe_1_6_2_U93 ( .A(pe_1_6_2_int_q_reg_h[14]), .B(
        pe_1_6_2_int_q_reg_h[10]), .S(pe_1_6_2_n56), .Z(pe_1_6_2_n48) );
  MUX2_X1 pe_1_6_2_U92 ( .A(pe_1_6_2_int_q_reg_h[6]), .B(
        pe_1_6_2_int_q_reg_h[2]), .S(pe_1_6_2_n56), .Z(pe_1_6_2_n47) );
  MUX2_X1 pe_1_6_2_U91 ( .A(pe_1_6_2_n46), .B(pe_1_6_2_n24), .S(n53), .Z(
        int_data_x_6__2__1_) );
  MUX2_X1 pe_1_6_2_U90 ( .A(pe_1_6_2_n45), .B(pe_1_6_2_n25), .S(pe_1_6_2_n60), 
        .Z(pe_1_6_2_n46) );
  MUX2_X1 pe_1_6_2_U89 ( .A(pe_1_6_2_int_q_reg_h[21]), .B(
        pe_1_6_2_int_q_reg_h[17]), .S(pe_1_6_2_n56), .Z(pe_1_6_2_n45) );
  MUX2_X1 pe_1_6_2_U88 ( .A(pe_1_6_2_int_q_reg_h[13]), .B(
        pe_1_6_2_int_q_reg_h[9]), .S(pe_1_6_2_n56), .Z(pe_1_6_2_n25) );
  MUX2_X1 pe_1_6_2_U87 ( .A(pe_1_6_2_int_q_reg_h[5]), .B(
        pe_1_6_2_int_q_reg_h[1]), .S(pe_1_6_2_n56), .Z(pe_1_6_2_n24) );
  MUX2_X1 pe_1_6_2_U86 ( .A(pe_1_6_2_n23), .B(pe_1_6_2_n20), .S(n53), .Z(
        int_data_x_6__2__0_) );
  MUX2_X1 pe_1_6_2_U85 ( .A(pe_1_6_2_n22), .B(pe_1_6_2_n21), .S(pe_1_6_2_n60), 
        .Z(pe_1_6_2_n23) );
  MUX2_X1 pe_1_6_2_U84 ( .A(pe_1_6_2_int_q_reg_h[20]), .B(
        pe_1_6_2_int_q_reg_h[16]), .S(pe_1_6_2_n56), .Z(pe_1_6_2_n22) );
  MUX2_X1 pe_1_6_2_U83 ( .A(pe_1_6_2_int_q_reg_h[12]), .B(
        pe_1_6_2_int_q_reg_h[8]), .S(pe_1_6_2_n56), .Z(pe_1_6_2_n21) );
  MUX2_X1 pe_1_6_2_U82 ( .A(pe_1_6_2_int_q_reg_h[4]), .B(
        pe_1_6_2_int_q_reg_h[0]), .S(pe_1_6_2_n56), .Z(pe_1_6_2_n20) );
  MUX2_X1 pe_1_6_2_U81 ( .A(pe_1_6_2_n19), .B(pe_1_6_2_n16), .S(n53), .Z(
        int_data_y_6__2__3_) );
  MUX2_X1 pe_1_6_2_U80 ( .A(pe_1_6_2_n18), .B(pe_1_6_2_n17), .S(pe_1_6_2_n60), 
        .Z(pe_1_6_2_n19) );
  MUX2_X1 pe_1_6_2_U79 ( .A(pe_1_6_2_int_q_reg_v[23]), .B(
        pe_1_6_2_int_q_reg_v[19]), .S(pe_1_6_2_n55), .Z(pe_1_6_2_n18) );
  MUX2_X1 pe_1_6_2_U78 ( .A(pe_1_6_2_int_q_reg_v[15]), .B(
        pe_1_6_2_int_q_reg_v[11]), .S(pe_1_6_2_n55), .Z(pe_1_6_2_n17) );
  MUX2_X1 pe_1_6_2_U77 ( .A(pe_1_6_2_int_q_reg_v[7]), .B(
        pe_1_6_2_int_q_reg_v[3]), .S(pe_1_6_2_n55), .Z(pe_1_6_2_n16) );
  MUX2_X1 pe_1_6_2_U76 ( .A(pe_1_6_2_n15), .B(pe_1_6_2_n12), .S(n53), .Z(
        int_data_y_6__2__2_) );
  MUX2_X1 pe_1_6_2_U75 ( .A(pe_1_6_2_n14), .B(pe_1_6_2_n13), .S(pe_1_6_2_n60), 
        .Z(pe_1_6_2_n15) );
  MUX2_X1 pe_1_6_2_U74 ( .A(pe_1_6_2_int_q_reg_v[22]), .B(
        pe_1_6_2_int_q_reg_v[18]), .S(pe_1_6_2_n55), .Z(pe_1_6_2_n14) );
  MUX2_X1 pe_1_6_2_U73 ( .A(pe_1_6_2_int_q_reg_v[14]), .B(
        pe_1_6_2_int_q_reg_v[10]), .S(pe_1_6_2_n55), .Z(pe_1_6_2_n13) );
  MUX2_X1 pe_1_6_2_U72 ( .A(pe_1_6_2_int_q_reg_v[6]), .B(
        pe_1_6_2_int_q_reg_v[2]), .S(pe_1_6_2_n55), .Z(pe_1_6_2_n12) );
  MUX2_X1 pe_1_6_2_U71 ( .A(pe_1_6_2_n11), .B(pe_1_6_2_n8), .S(n53), .Z(
        int_data_y_6__2__1_) );
  MUX2_X1 pe_1_6_2_U70 ( .A(pe_1_6_2_n10), .B(pe_1_6_2_n9), .S(pe_1_6_2_n60), 
        .Z(pe_1_6_2_n11) );
  MUX2_X1 pe_1_6_2_U69 ( .A(pe_1_6_2_int_q_reg_v[21]), .B(
        pe_1_6_2_int_q_reg_v[17]), .S(pe_1_6_2_n55), .Z(pe_1_6_2_n10) );
  MUX2_X1 pe_1_6_2_U68 ( .A(pe_1_6_2_int_q_reg_v[13]), .B(
        pe_1_6_2_int_q_reg_v[9]), .S(pe_1_6_2_n55), .Z(pe_1_6_2_n9) );
  MUX2_X1 pe_1_6_2_U67 ( .A(pe_1_6_2_int_q_reg_v[5]), .B(
        pe_1_6_2_int_q_reg_v[1]), .S(pe_1_6_2_n55), .Z(pe_1_6_2_n8) );
  MUX2_X1 pe_1_6_2_U66 ( .A(pe_1_6_2_n7), .B(pe_1_6_2_n4), .S(n53), .Z(
        int_data_y_6__2__0_) );
  MUX2_X1 pe_1_6_2_U65 ( .A(pe_1_6_2_n6), .B(pe_1_6_2_n5), .S(pe_1_6_2_n60), 
        .Z(pe_1_6_2_n7) );
  MUX2_X1 pe_1_6_2_U64 ( .A(pe_1_6_2_int_q_reg_v[20]), .B(
        pe_1_6_2_int_q_reg_v[16]), .S(pe_1_6_2_n55), .Z(pe_1_6_2_n6) );
  MUX2_X1 pe_1_6_2_U63 ( .A(pe_1_6_2_int_q_reg_v[12]), .B(
        pe_1_6_2_int_q_reg_v[8]), .S(pe_1_6_2_n55), .Z(pe_1_6_2_n5) );
  MUX2_X1 pe_1_6_2_U62 ( .A(pe_1_6_2_int_q_reg_v[4]), .B(
        pe_1_6_2_int_q_reg_v[0]), .S(pe_1_6_2_n55), .Z(pe_1_6_2_n4) );
  AOI222_X1 pe_1_6_2_U61 ( .A1(int_data_res_7__2__2_), .A2(pe_1_6_2_n62), .B1(
        pe_1_6_2_N80), .B2(pe_1_6_2_n27), .C1(pe_1_6_2_N72), .C2(pe_1_6_2_n28), 
        .ZN(pe_1_6_2_n33) );
  INV_X1 pe_1_6_2_U60 ( .A(pe_1_6_2_n33), .ZN(pe_1_6_2_n79) );
  AOI222_X1 pe_1_6_2_U59 ( .A1(int_data_res_7__2__6_), .A2(pe_1_6_2_n62), .B1(
        pe_1_6_2_N84), .B2(pe_1_6_2_n27), .C1(pe_1_6_2_N76), .C2(pe_1_6_2_n28), 
        .ZN(pe_1_6_2_n29) );
  INV_X1 pe_1_6_2_U58 ( .A(pe_1_6_2_n29), .ZN(pe_1_6_2_n75) );
  XNOR2_X1 pe_1_6_2_U57 ( .A(pe_1_6_2_n70), .B(int_data_res_6__2__0_), .ZN(
        pe_1_6_2_N70) );
  AOI222_X1 pe_1_6_2_U52 ( .A1(int_data_res_7__2__0_), .A2(pe_1_6_2_n62), .B1(
        pe_1_6_2_n1), .B2(pe_1_6_2_n27), .C1(pe_1_6_2_N70), .C2(pe_1_6_2_n28), 
        .ZN(pe_1_6_2_n35) );
  INV_X1 pe_1_6_2_U51 ( .A(pe_1_6_2_n35), .ZN(pe_1_6_2_n81) );
  AOI222_X1 pe_1_6_2_U50 ( .A1(int_data_res_7__2__1_), .A2(pe_1_6_2_n62), .B1(
        pe_1_6_2_N79), .B2(pe_1_6_2_n27), .C1(pe_1_6_2_N71), .C2(pe_1_6_2_n28), 
        .ZN(pe_1_6_2_n34) );
  INV_X1 pe_1_6_2_U49 ( .A(pe_1_6_2_n34), .ZN(pe_1_6_2_n80) );
  AOI222_X1 pe_1_6_2_U48 ( .A1(int_data_res_7__2__3_), .A2(pe_1_6_2_n62), .B1(
        pe_1_6_2_N81), .B2(pe_1_6_2_n27), .C1(pe_1_6_2_N73), .C2(pe_1_6_2_n28), 
        .ZN(pe_1_6_2_n32) );
  INV_X1 pe_1_6_2_U47 ( .A(pe_1_6_2_n32), .ZN(pe_1_6_2_n78) );
  AOI222_X1 pe_1_6_2_U46 ( .A1(int_data_res_7__2__4_), .A2(pe_1_6_2_n62), .B1(
        pe_1_6_2_N82), .B2(pe_1_6_2_n27), .C1(pe_1_6_2_N74), .C2(pe_1_6_2_n28), 
        .ZN(pe_1_6_2_n31) );
  INV_X1 pe_1_6_2_U45 ( .A(pe_1_6_2_n31), .ZN(pe_1_6_2_n77) );
  AOI222_X1 pe_1_6_2_U44 ( .A1(int_data_res_7__2__5_), .A2(pe_1_6_2_n62), .B1(
        pe_1_6_2_N83), .B2(pe_1_6_2_n27), .C1(pe_1_6_2_N75), .C2(pe_1_6_2_n28), 
        .ZN(pe_1_6_2_n30) );
  INV_X1 pe_1_6_2_U43 ( .A(pe_1_6_2_n30), .ZN(pe_1_6_2_n76) );
  NAND2_X1 pe_1_6_2_U42 ( .A1(pe_1_6_2_int_data_0_), .A2(pe_1_6_2_n3), .ZN(
        pe_1_6_2_sub_81_carry[1]) );
  INV_X1 pe_1_6_2_U41 ( .A(pe_1_6_2_int_data_1_), .ZN(pe_1_6_2_n71) );
  INV_X1 pe_1_6_2_U40 ( .A(pe_1_6_2_int_data_2_), .ZN(pe_1_6_2_n72) );
  AND2_X1 pe_1_6_2_U39 ( .A1(pe_1_6_2_int_data_0_), .A2(int_data_res_6__2__0_), 
        .ZN(pe_1_6_2_n2) );
  AOI222_X1 pe_1_6_2_U38 ( .A1(pe_1_6_2_n62), .A2(int_data_res_7__2__7_), .B1(
        pe_1_6_2_N85), .B2(pe_1_6_2_n27), .C1(pe_1_6_2_N77), .C2(pe_1_6_2_n28), 
        .ZN(pe_1_6_2_n26) );
  INV_X1 pe_1_6_2_U37 ( .A(pe_1_6_2_n26), .ZN(pe_1_6_2_n74) );
  NOR3_X1 pe_1_6_2_U36 ( .A1(pe_1_6_2_n58), .A2(pe_1_6_2_n63), .A3(int_ckg[13]), .ZN(pe_1_6_2_n36) );
  OR2_X1 pe_1_6_2_U35 ( .A1(pe_1_6_2_n36), .A2(pe_1_6_2_n62), .ZN(pe_1_6_2_N90) );
  INV_X1 pe_1_6_2_U34 ( .A(n41), .ZN(pe_1_6_2_n61) );
  AND2_X1 pe_1_6_2_U33 ( .A1(int_data_x_6__2__2_), .A2(n29), .ZN(
        pe_1_6_2_int_data_2_) );
  AND2_X1 pe_1_6_2_U32 ( .A1(int_data_x_6__2__1_), .A2(n29), .ZN(
        pe_1_6_2_int_data_1_) );
  AND2_X1 pe_1_6_2_U31 ( .A1(int_data_x_6__2__3_), .A2(n29), .ZN(
        pe_1_6_2_int_data_3_) );
  BUF_X1 pe_1_6_2_U30 ( .A(n63), .Z(pe_1_6_2_n62) );
  INV_X1 pe_1_6_2_U29 ( .A(n35), .ZN(pe_1_6_2_n59) );
  AND2_X1 pe_1_6_2_U28 ( .A1(int_data_x_6__2__0_), .A2(n29), .ZN(
        pe_1_6_2_int_data_0_) );
  NAND2_X1 pe_1_6_2_U27 ( .A1(pe_1_6_2_n44), .A2(pe_1_6_2_n59), .ZN(
        pe_1_6_2_n41) );
  AND3_X1 pe_1_6_2_U26 ( .A1(n77), .A2(pe_1_6_2_n61), .A3(n53), .ZN(
        pe_1_6_2_n44) );
  INV_X1 pe_1_6_2_U25 ( .A(pe_1_6_2_int_data_3_), .ZN(pe_1_6_2_n73) );
  NOR2_X1 pe_1_6_2_U24 ( .A1(pe_1_6_2_n67), .A2(n53), .ZN(pe_1_6_2_n43) );
  NOR2_X1 pe_1_6_2_U23 ( .A1(pe_1_6_2_n57), .A2(pe_1_6_2_n62), .ZN(
        pe_1_6_2_n28) );
  NOR2_X1 pe_1_6_2_U22 ( .A1(n21), .A2(pe_1_6_2_n62), .ZN(pe_1_6_2_n27) );
  INV_X1 pe_1_6_2_U21 ( .A(pe_1_6_2_int_data_0_), .ZN(pe_1_6_2_n70) );
  INV_X1 pe_1_6_2_U20 ( .A(pe_1_6_2_n41), .ZN(pe_1_6_2_n87) );
  INV_X1 pe_1_6_2_U19 ( .A(pe_1_6_2_n37), .ZN(pe_1_6_2_n85) );
  INV_X1 pe_1_6_2_U18 ( .A(pe_1_6_2_n38), .ZN(pe_1_6_2_n84) );
  INV_X1 pe_1_6_2_U17 ( .A(pe_1_6_2_n39), .ZN(pe_1_6_2_n83) );
  NOR2_X1 pe_1_6_2_U16 ( .A1(pe_1_6_2_n65), .A2(pe_1_6_2_n42), .ZN(
        pe_1_6_2_N59) );
  NOR2_X1 pe_1_6_2_U15 ( .A1(pe_1_6_2_n65), .A2(pe_1_6_2_n41), .ZN(
        pe_1_6_2_N60) );
  NOR2_X1 pe_1_6_2_U14 ( .A1(pe_1_6_2_n65), .A2(pe_1_6_2_n38), .ZN(
        pe_1_6_2_N63) );
  NOR2_X1 pe_1_6_2_U13 ( .A1(pe_1_6_2_n65), .A2(pe_1_6_2_n40), .ZN(
        pe_1_6_2_N61) );
  NOR2_X1 pe_1_6_2_U12 ( .A1(pe_1_6_2_n65), .A2(pe_1_6_2_n39), .ZN(
        pe_1_6_2_N62) );
  NOR2_X1 pe_1_6_2_U11 ( .A1(pe_1_6_2_n37), .A2(pe_1_6_2_n65), .ZN(
        pe_1_6_2_N64) );
  NAND2_X1 pe_1_6_2_U10 ( .A1(pe_1_6_2_n44), .A2(n35), .ZN(pe_1_6_2_n42) );
  BUF_X1 pe_1_6_2_U9 ( .A(n35), .Z(pe_1_6_2_n55) );
  INV_X1 pe_1_6_2_U8 ( .A(pe_1_6_2_n66), .ZN(pe_1_6_2_n63) );
  BUF_X1 pe_1_6_2_U7 ( .A(n35), .Z(pe_1_6_2_n56) );
  INV_X1 pe_1_6_2_U6 ( .A(pe_1_6_2_n42), .ZN(pe_1_6_2_n86) );
  INV_X1 pe_1_6_2_U5 ( .A(pe_1_6_2_n40), .ZN(pe_1_6_2_n82) );
  INV_X2 pe_1_6_2_U4 ( .A(n85), .ZN(pe_1_6_2_n69) );
  XOR2_X1 pe_1_6_2_U3 ( .A(pe_1_6_2_int_data_0_), .B(int_data_res_6__2__0_), 
        .Z(pe_1_6_2_n1) );
  DFFR_X1 pe_1_6_2_int_q_acc_reg_0_ ( .D(pe_1_6_2_n81), .CK(pe_1_6_2_net3652), 
        .RN(pe_1_6_2_n69), .Q(int_data_res_6__2__0_), .QN(pe_1_6_2_n3) );
  DFFR_X1 pe_1_6_2_int_q_reg_v_reg_0__0_ ( .D(int_data_y_7__2__0_), .CK(
        pe_1_6_2_net3622), .RN(pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_v[20]) );
  DFFR_X1 pe_1_6_2_int_q_reg_v_reg_0__1_ ( .D(int_data_y_7__2__1_), .CK(
        pe_1_6_2_net3622), .RN(pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_v[21]) );
  DFFR_X1 pe_1_6_2_int_q_reg_v_reg_0__2_ ( .D(int_data_y_7__2__2_), .CK(
        pe_1_6_2_net3622), .RN(pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_v[22]) );
  DFFR_X1 pe_1_6_2_int_q_reg_v_reg_0__3_ ( .D(int_data_y_7__2__3_), .CK(
        pe_1_6_2_net3622), .RN(pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_v[23]) );
  DFFR_X1 pe_1_6_2_int_q_reg_v_reg_1__0_ ( .D(int_data_y_7__2__0_), .CK(
        pe_1_6_2_net3627), .RN(pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_v[16]) );
  DFFR_X1 pe_1_6_2_int_q_reg_v_reg_1__1_ ( .D(int_data_y_7__2__1_), .CK(
        pe_1_6_2_net3627), .RN(pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_v[17]) );
  DFFR_X1 pe_1_6_2_int_q_reg_v_reg_1__2_ ( .D(int_data_y_7__2__2_), .CK(
        pe_1_6_2_net3627), .RN(pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_v[18]) );
  DFFR_X1 pe_1_6_2_int_q_reg_v_reg_1__3_ ( .D(int_data_y_7__2__3_), .CK(
        pe_1_6_2_net3627), .RN(pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_v[19]) );
  DFFR_X1 pe_1_6_2_int_q_reg_v_reg_2__0_ ( .D(int_data_y_7__2__0_), .CK(
        pe_1_6_2_net3632), .RN(pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_v[12]) );
  DFFR_X1 pe_1_6_2_int_q_reg_v_reg_2__1_ ( .D(int_data_y_7__2__1_), .CK(
        pe_1_6_2_net3632), .RN(pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_v[13]) );
  DFFR_X1 pe_1_6_2_int_q_reg_v_reg_2__2_ ( .D(int_data_y_7__2__2_), .CK(
        pe_1_6_2_net3632), .RN(pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_v[14]) );
  DFFR_X1 pe_1_6_2_int_q_reg_v_reg_2__3_ ( .D(int_data_y_7__2__3_), .CK(
        pe_1_6_2_net3632), .RN(pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_v[15]) );
  DFFR_X1 pe_1_6_2_int_q_reg_v_reg_3__0_ ( .D(int_data_y_7__2__0_), .CK(
        pe_1_6_2_net3637), .RN(pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_v[8]) );
  DFFR_X1 pe_1_6_2_int_q_reg_v_reg_3__1_ ( .D(int_data_y_7__2__1_), .CK(
        pe_1_6_2_net3637), .RN(pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_v[9]) );
  DFFR_X1 pe_1_6_2_int_q_reg_v_reg_3__2_ ( .D(int_data_y_7__2__2_), .CK(
        pe_1_6_2_net3637), .RN(pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_v[10]) );
  DFFR_X1 pe_1_6_2_int_q_reg_v_reg_3__3_ ( .D(int_data_y_7__2__3_), .CK(
        pe_1_6_2_net3637), .RN(pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_v[11]) );
  DFFR_X1 pe_1_6_2_int_q_reg_v_reg_4__0_ ( .D(int_data_y_7__2__0_), .CK(
        pe_1_6_2_net3642), .RN(pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_v[4]) );
  DFFR_X1 pe_1_6_2_int_q_reg_v_reg_4__1_ ( .D(int_data_y_7__2__1_), .CK(
        pe_1_6_2_net3642), .RN(pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_v[5]) );
  DFFR_X1 pe_1_6_2_int_q_reg_v_reg_4__2_ ( .D(int_data_y_7__2__2_), .CK(
        pe_1_6_2_net3642), .RN(pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_v[6]) );
  DFFR_X1 pe_1_6_2_int_q_reg_v_reg_4__3_ ( .D(int_data_y_7__2__3_), .CK(
        pe_1_6_2_net3642), .RN(pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_v[7]) );
  DFFR_X1 pe_1_6_2_int_q_reg_v_reg_5__0_ ( .D(int_data_y_7__2__0_), .CK(
        pe_1_6_2_net3647), .RN(pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_v[0]) );
  DFFR_X1 pe_1_6_2_int_q_reg_v_reg_5__1_ ( .D(int_data_y_7__2__1_), .CK(
        pe_1_6_2_net3647), .RN(pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_v[1]) );
  DFFR_X1 pe_1_6_2_int_q_reg_v_reg_5__2_ ( .D(int_data_y_7__2__2_), .CK(
        pe_1_6_2_net3647), .RN(pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_v[2]) );
  DFFR_X1 pe_1_6_2_int_q_reg_v_reg_5__3_ ( .D(int_data_y_7__2__3_), .CK(
        pe_1_6_2_net3647), .RN(pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_6_2_int_q_reg_h_reg_0__0_ ( .D(int_data_x_6__3__0_), .SI(
        int_data_y_7__2__0_), .SE(pe_1_6_2_n63), .CK(pe_1_6_2_net3591), .RN(
        pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_6_2_int_q_reg_h_reg_0__1_ ( .D(int_data_x_6__3__1_), .SI(
        int_data_y_7__2__1_), .SE(pe_1_6_2_n63), .CK(pe_1_6_2_net3591), .RN(
        pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_6_2_int_q_reg_h_reg_0__2_ ( .D(int_data_x_6__3__2_), .SI(
        int_data_y_7__2__2_), .SE(pe_1_6_2_n63), .CK(pe_1_6_2_net3591), .RN(
        pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_6_2_int_q_reg_h_reg_0__3_ ( .D(int_data_x_6__3__3_), .SI(
        int_data_y_7__2__3_), .SE(pe_1_6_2_n63), .CK(pe_1_6_2_net3591), .RN(
        pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_6_2_int_q_reg_h_reg_1__0_ ( .D(int_data_x_6__3__0_), .SI(
        int_data_y_7__2__0_), .SE(pe_1_6_2_n63), .CK(pe_1_6_2_net3597), .RN(
        pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_6_2_int_q_reg_h_reg_1__1_ ( .D(int_data_x_6__3__1_), .SI(
        int_data_y_7__2__1_), .SE(pe_1_6_2_n63), .CK(pe_1_6_2_net3597), .RN(
        pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_6_2_int_q_reg_h_reg_1__2_ ( .D(int_data_x_6__3__2_), .SI(
        int_data_y_7__2__2_), .SE(pe_1_6_2_n63), .CK(pe_1_6_2_net3597), .RN(
        pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_6_2_int_q_reg_h_reg_1__3_ ( .D(int_data_x_6__3__3_), .SI(
        int_data_y_7__2__3_), .SE(pe_1_6_2_n63), .CK(pe_1_6_2_net3597), .RN(
        pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_6_2_int_q_reg_h_reg_2__0_ ( .D(int_data_x_6__3__0_), .SI(
        int_data_y_7__2__0_), .SE(pe_1_6_2_n63), .CK(pe_1_6_2_net3602), .RN(
        pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_6_2_int_q_reg_h_reg_2__1_ ( .D(int_data_x_6__3__1_), .SI(
        int_data_y_7__2__1_), .SE(pe_1_6_2_n63), .CK(pe_1_6_2_net3602), .RN(
        pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_6_2_int_q_reg_h_reg_2__2_ ( .D(int_data_x_6__3__2_), .SI(
        int_data_y_7__2__2_), .SE(pe_1_6_2_n63), .CK(pe_1_6_2_net3602), .RN(
        pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_6_2_int_q_reg_h_reg_2__3_ ( .D(int_data_x_6__3__3_), .SI(
        int_data_y_7__2__3_), .SE(pe_1_6_2_n63), .CK(pe_1_6_2_net3602), .RN(
        pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_6_2_int_q_reg_h_reg_3__0_ ( .D(int_data_x_6__3__0_), .SI(
        int_data_y_7__2__0_), .SE(pe_1_6_2_n63), .CK(pe_1_6_2_net3607), .RN(
        pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_6_2_int_q_reg_h_reg_3__1_ ( .D(int_data_x_6__3__1_), .SI(
        int_data_y_7__2__1_), .SE(pe_1_6_2_n63), .CK(pe_1_6_2_net3607), .RN(
        pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_6_2_int_q_reg_h_reg_3__2_ ( .D(int_data_x_6__3__2_), .SI(
        int_data_y_7__2__2_), .SE(pe_1_6_2_n63), .CK(pe_1_6_2_net3607), .RN(
        pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_6_2_int_q_reg_h_reg_3__3_ ( .D(int_data_x_6__3__3_), .SI(
        int_data_y_7__2__3_), .SE(pe_1_6_2_n63), .CK(pe_1_6_2_net3607), .RN(
        pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_6_2_int_q_reg_h_reg_4__0_ ( .D(int_data_x_6__3__0_), .SI(
        int_data_y_7__2__0_), .SE(pe_1_6_2_n64), .CK(pe_1_6_2_net3612), .RN(
        pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_6_2_int_q_reg_h_reg_4__1_ ( .D(int_data_x_6__3__1_), .SI(
        int_data_y_7__2__1_), .SE(pe_1_6_2_n64), .CK(pe_1_6_2_net3612), .RN(
        pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_6_2_int_q_reg_h_reg_4__2_ ( .D(int_data_x_6__3__2_), .SI(
        int_data_y_7__2__2_), .SE(pe_1_6_2_n64), .CK(pe_1_6_2_net3612), .RN(
        pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_6_2_int_q_reg_h_reg_4__3_ ( .D(int_data_x_6__3__3_), .SI(
        int_data_y_7__2__3_), .SE(pe_1_6_2_n64), .CK(pe_1_6_2_net3612), .RN(
        pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_6_2_int_q_reg_h_reg_5__0_ ( .D(int_data_x_6__3__0_), .SI(
        int_data_y_7__2__0_), .SE(pe_1_6_2_n64), .CK(pe_1_6_2_net3617), .RN(
        pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_6_2_int_q_reg_h_reg_5__1_ ( .D(int_data_x_6__3__1_), .SI(
        int_data_y_7__2__1_), .SE(pe_1_6_2_n64), .CK(pe_1_6_2_net3617), .RN(
        pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_6_2_int_q_reg_h_reg_5__2_ ( .D(int_data_x_6__3__2_), .SI(
        int_data_y_7__2__2_), .SE(pe_1_6_2_n64), .CK(pe_1_6_2_net3617), .RN(
        pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_6_2_int_q_reg_h_reg_5__3_ ( .D(int_data_x_6__3__3_), .SI(
        int_data_y_7__2__3_), .SE(pe_1_6_2_n64), .CK(pe_1_6_2_net3617), .RN(
        pe_1_6_2_n69), .Q(pe_1_6_2_int_q_reg_h[3]) );
  FA_X1 pe_1_6_2_sub_81_U2_7 ( .A(int_data_res_6__2__7_), .B(pe_1_6_2_n73), 
        .CI(pe_1_6_2_sub_81_carry[7]), .S(pe_1_6_2_N77) );
  FA_X1 pe_1_6_2_sub_81_U2_6 ( .A(int_data_res_6__2__6_), .B(pe_1_6_2_n73), 
        .CI(pe_1_6_2_sub_81_carry[6]), .CO(pe_1_6_2_sub_81_carry[7]), .S(
        pe_1_6_2_N76) );
  FA_X1 pe_1_6_2_sub_81_U2_5 ( .A(int_data_res_6__2__5_), .B(pe_1_6_2_n73), 
        .CI(pe_1_6_2_sub_81_carry[5]), .CO(pe_1_6_2_sub_81_carry[6]), .S(
        pe_1_6_2_N75) );
  FA_X1 pe_1_6_2_sub_81_U2_4 ( .A(int_data_res_6__2__4_), .B(pe_1_6_2_n73), 
        .CI(pe_1_6_2_sub_81_carry[4]), .CO(pe_1_6_2_sub_81_carry[5]), .S(
        pe_1_6_2_N74) );
  FA_X1 pe_1_6_2_sub_81_U2_3 ( .A(int_data_res_6__2__3_), .B(pe_1_6_2_n73), 
        .CI(pe_1_6_2_sub_81_carry[3]), .CO(pe_1_6_2_sub_81_carry[4]), .S(
        pe_1_6_2_N73) );
  FA_X1 pe_1_6_2_sub_81_U2_2 ( .A(int_data_res_6__2__2_), .B(pe_1_6_2_n72), 
        .CI(pe_1_6_2_sub_81_carry[2]), .CO(pe_1_6_2_sub_81_carry[3]), .S(
        pe_1_6_2_N72) );
  FA_X1 pe_1_6_2_sub_81_U2_1 ( .A(int_data_res_6__2__1_), .B(pe_1_6_2_n71), 
        .CI(pe_1_6_2_sub_81_carry[1]), .CO(pe_1_6_2_sub_81_carry[2]), .S(
        pe_1_6_2_N71) );
  FA_X1 pe_1_6_2_add_83_U1_7 ( .A(int_data_res_6__2__7_), .B(
        pe_1_6_2_int_data_3_), .CI(pe_1_6_2_add_83_carry[7]), .S(pe_1_6_2_N85)
         );
  FA_X1 pe_1_6_2_add_83_U1_6 ( .A(int_data_res_6__2__6_), .B(
        pe_1_6_2_int_data_3_), .CI(pe_1_6_2_add_83_carry[6]), .CO(
        pe_1_6_2_add_83_carry[7]), .S(pe_1_6_2_N84) );
  FA_X1 pe_1_6_2_add_83_U1_5 ( .A(int_data_res_6__2__5_), .B(
        pe_1_6_2_int_data_3_), .CI(pe_1_6_2_add_83_carry[5]), .CO(
        pe_1_6_2_add_83_carry[6]), .S(pe_1_6_2_N83) );
  FA_X1 pe_1_6_2_add_83_U1_4 ( .A(int_data_res_6__2__4_), .B(
        pe_1_6_2_int_data_3_), .CI(pe_1_6_2_add_83_carry[4]), .CO(
        pe_1_6_2_add_83_carry[5]), .S(pe_1_6_2_N82) );
  FA_X1 pe_1_6_2_add_83_U1_3 ( .A(int_data_res_6__2__3_), .B(
        pe_1_6_2_int_data_3_), .CI(pe_1_6_2_add_83_carry[3]), .CO(
        pe_1_6_2_add_83_carry[4]), .S(pe_1_6_2_N81) );
  FA_X1 pe_1_6_2_add_83_U1_2 ( .A(int_data_res_6__2__2_), .B(
        pe_1_6_2_int_data_2_), .CI(pe_1_6_2_add_83_carry[2]), .CO(
        pe_1_6_2_add_83_carry[3]), .S(pe_1_6_2_N80) );
  FA_X1 pe_1_6_2_add_83_U1_1 ( .A(int_data_res_6__2__1_), .B(
        pe_1_6_2_int_data_1_), .CI(pe_1_6_2_n2), .CO(pe_1_6_2_add_83_carry[2]), 
        .S(pe_1_6_2_N79) );
  NAND3_X1 pe_1_6_2_U56 ( .A1(n35), .A2(pe_1_6_2_n43), .A3(pe_1_6_2_n60), .ZN(
        pe_1_6_2_n40) );
  NAND3_X1 pe_1_6_2_U55 ( .A1(pe_1_6_2_n43), .A2(pe_1_6_2_n59), .A3(
        pe_1_6_2_n60), .ZN(pe_1_6_2_n39) );
  NAND3_X1 pe_1_6_2_U54 ( .A1(pe_1_6_2_n43), .A2(pe_1_6_2_n61), .A3(n35), .ZN(
        pe_1_6_2_n38) );
  NAND3_X1 pe_1_6_2_U53 ( .A1(pe_1_6_2_n59), .A2(pe_1_6_2_n61), .A3(
        pe_1_6_2_n43), .ZN(pe_1_6_2_n37) );
  DFFR_X1 pe_1_6_2_int_q_acc_reg_6_ ( .D(pe_1_6_2_n75), .CK(pe_1_6_2_net3652), 
        .RN(pe_1_6_2_n68), .Q(int_data_res_6__2__6_) );
  DFFR_X1 pe_1_6_2_int_q_acc_reg_5_ ( .D(pe_1_6_2_n76), .CK(pe_1_6_2_net3652), 
        .RN(pe_1_6_2_n68), .Q(int_data_res_6__2__5_) );
  DFFR_X1 pe_1_6_2_int_q_acc_reg_4_ ( .D(pe_1_6_2_n77), .CK(pe_1_6_2_net3652), 
        .RN(pe_1_6_2_n68), .Q(int_data_res_6__2__4_) );
  DFFR_X1 pe_1_6_2_int_q_acc_reg_3_ ( .D(pe_1_6_2_n78), .CK(pe_1_6_2_net3652), 
        .RN(pe_1_6_2_n68), .Q(int_data_res_6__2__3_) );
  DFFR_X1 pe_1_6_2_int_q_acc_reg_2_ ( .D(pe_1_6_2_n79), .CK(pe_1_6_2_net3652), 
        .RN(pe_1_6_2_n68), .Q(int_data_res_6__2__2_) );
  DFFR_X1 pe_1_6_2_int_q_acc_reg_1_ ( .D(pe_1_6_2_n80), .CK(pe_1_6_2_net3652), 
        .RN(pe_1_6_2_n68), .Q(int_data_res_6__2__1_) );
  DFFR_X1 pe_1_6_2_int_q_acc_reg_7_ ( .D(pe_1_6_2_n74), .CK(pe_1_6_2_net3652), 
        .RN(pe_1_6_2_n68), .Q(int_data_res_6__2__7_) );
  CLKGATETST_X1 pe_1_6_2_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_6_2_n85), .SE(1'b0), .GCK(pe_1_6_2_net3591) );
  CLKGATETST_X1 pe_1_6_2_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_6_2_n84), .SE(1'b0), .GCK(pe_1_6_2_net3597) );
  CLKGATETST_X1 pe_1_6_2_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_6_2_n83), .SE(1'b0), .GCK(pe_1_6_2_net3602) );
  CLKGATETST_X1 pe_1_6_2_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_6_2_n82), .SE(1'b0), .GCK(pe_1_6_2_net3607) );
  CLKGATETST_X1 pe_1_6_2_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_6_2_n87), .SE(1'b0), .GCK(pe_1_6_2_net3612) );
  CLKGATETST_X1 pe_1_6_2_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_6_2_n86), .SE(1'b0), .GCK(pe_1_6_2_net3617) );
  CLKGATETST_X1 pe_1_6_2_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_6_2_N64), .SE(1'b0), .GCK(pe_1_6_2_net3622) );
  CLKGATETST_X1 pe_1_6_2_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_6_2_N63), .SE(1'b0), .GCK(pe_1_6_2_net3627) );
  CLKGATETST_X1 pe_1_6_2_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_6_2_N62), .SE(1'b0), .GCK(pe_1_6_2_net3632) );
  CLKGATETST_X1 pe_1_6_2_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_6_2_N61), .SE(1'b0), .GCK(pe_1_6_2_net3637) );
  CLKGATETST_X1 pe_1_6_2_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_6_2_N60), .SE(1'b0), .GCK(pe_1_6_2_net3642) );
  CLKGATETST_X1 pe_1_6_2_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_6_2_N59), .SE(1'b0), .GCK(pe_1_6_2_net3647) );
  CLKGATETST_X1 pe_1_6_2_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_6_2_N90), .SE(1'b0), .GCK(pe_1_6_2_net3652) );
  CLKBUF_X1 pe_1_6_3_U110 ( .A(pe_1_6_3_n70), .Z(pe_1_6_3_n69) );
  INV_X1 pe_1_6_3_U109 ( .A(n77), .ZN(pe_1_6_3_n68) );
  INV_X1 pe_1_6_3_U108 ( .A(n69), .ZN(pe_1_6_3_n67) );
  INV_X1 pe_1_6_3_U107 ( .A(n69), .ZN(pe_1_6_3_n66) );
  INV_X1 pe_1_6_3_U106 ( .A(pe_1_6_3_n67), .ZN(pe_1_6_3_n65) );
  INV_X1 pe_1_6_3_U105 ( .A(pe_1_6_3_n62), .ZN(pe_1_6_3_n61) );
  INV_X1 pe_1_6_3_U104 ( .A(pe_1_6_3_n60), .ZN(pe_1_6_3_n59) );
  INV_X1 pe_1_6_3_U103 ( .A(n29), .ZN(pe_1_6_3_n58) );
  INV_X1 pe_1_6_3_U102 ( .A(n21), .ZN(pe_1_6_3_n57) );
  MUX2_X1 pe_1_6_3_U101 ( .A(pe_1_6_3_n54), .B(pe_1_6_3_n51), .S(n53), .Z(
        int_data_x_6__3__3_) );
  MUX2_X1 pe_1_6_3_U100 ( .A(pe_1_6_3_n53), .B(pe_1_6_3_n52), .S(pe_1_6_3_n61), 
        .Z(pe_1_6_3_n54) );
  MUX2_X1 pe_1_6_3_U99 ( .A(pe_1_6_3_int_q_reg_h[23]), .B(
        pe_1_6_3_int_q_reg_h[19]), .S(pe_1_6_3_n56), .Z(pe_1_6_3_n53) );
  MUX2_X1 pe_1_6_3_U98 ( .A(pe_1_6_3_int_q_reg_h[15]), .B(
        pe_1_6_3_int_q_reg_h[11]), .S(pe_1_6_3_n56), .Z(pe_1_6_3_n52) );
  MUX2_X1 pe_1_6_3_U97 ( .A(pe_1_6_3_int_q_reg_h[7]), .B(
        pe_1_6_3_int_q_reg_h[3]), .S(pe_1_6_3_n56), .Z(pe_1_6_3_n51) );
  MUX2_X1 pe_1_6_3_U96 ( .A(pe_1_6_3_n50), .B(pe_1_6_3_n47), .S(n53), .Z(
        int_data_x_6__3__2_) );
  MUX2_X1 pe_1_6_3_U95 ( .A(pe_1_6_3_n49), .B(pe_1_6_3_n48), .S(pe_1_6_3_n61), 
        .Z(pe_1_6_3_n50) );
  MUX2_X1 pe_1_6_3_U94 ( .A(pe_1_6_3_int_q_reg_h[22]), .B(
        pe_1_6_3_int_q_reg_h[18]), .S(pe_1_6_3_n56), .Z(pe_1_6_3_n49) );
  MUX2_X1 pe_1_6_3_U93 ( .A(pe_1_6_3_int_q_reg_h[14]), .B(
        pe_1_6_3_int_q_reg_h[10]), .S(pe_1_6_3_n56), .Z(pe_1_6_3_n48) );
  MUX2_X1 pe_1_6_3_U92 ( .A(pe_1_6_3_int_q_reg_h[6]), .B(
        pe_1_6_3_int_q_reg_h[2]), .S(pe_1_6_3_n56), .Z(pe_1_6_3_n47) );
  MUX2_X1 pe_1_6_3_U91 ( .A(pe_1_6_3_n46), .B(pe_1_6_3_n24), .S(n53), .Z(
        int_data_x_6__3__1_) );
  MUX2_X1 pe_1_6_3_U90 ( .A(pe_1_6_3_n45), .B(pe_1_6_3_n25), .S(pe_1_6_3_n61), 
        .Z(pe_1_6_3_n46) );
  MUX2_X1 pe_1_6_3_U89 ( .A(pe_1_6_3_int_q_reg_h[21]), .B(
        pe_1_6_3_int_q_reg_h[17]), .S(pe_1_6_3_n56), .Z(pe_1_6_3_n45) );
  MUX2_X1 pe_1_6_3_U88 ( .A(pe_1_6_3_int_q_reg_h[13]), .B(
        pe_1_6_3_int_q_reg_h[9]), .S(pe_1_6_3_n56), .Z(pe_1_6_3_n25) );
  MUX2_X1 pe_1_6_3_U87 ( .A(pe_1_6_3_int_q_reg_h[5]), .B(
        pe_1_6_3_int_q_reg_h[1]), .S(pe_1_6_3_n56), .Z(pe_1_6_3_n24) );
  MUX2_X1 pe_1_6_3_U86 ( .A(pe_1_6_3_n23), .B(pe_1_6_3_n20), .S(n53), .Z(
        int_data_x_6__3__0_) );
  MUX2_X1 pe_1_6_3_U85 ( .A(pe_1_6_3_n22), .B(pe_1_6_3_n21), .S(pe_1_6_3_n61), 
        .Z(pe_1_6_3_n23) );
  MUX2_X1 pe_1_6_3_U84 ( .A(pe_1_6_3_int_q_reg_h[20]), .B(
        pe_1_6_3_int_q_reg_h[16]), .S(pe_1_6_3_n56), .Z(pe_1_6_3_n22) );
  MUX2_X1 pe_1_6_3_U83 ( .A(pe_1_6_3_int_q_reg_h[12]), .B(
        pe_1_6_3_int_q_reg_h[8]), .S(pe_1_6_3_n56), .Z(pe_1_6_3_n21) );
  MUX2_X1 pe_1_6_3_U82 ( .A(pe_1_6_3_int_q_reg_h[4]), .B(
        pe_1_6_3_int_q_reg_h[0]), .S(pe_1_6_3_n56), .Z(pe_1_6_3_n20) );
  MUX2_X1 pe_1_6_3_U81 ( .A(pe_1_6_3_n19), .B(pe_1_6_3_n16), .S(n53), .Z(
        int_data_y_6__3__3_) );
  MUX2_X1 pe_1_6_3_U80 ( .A(pe_1_6_3_n18), .B(pe_1_6_3_n17), .S(pe_1_6_3_n61), 
        .Z(pe_1_6_3_n19) );
  MUX2_X1 pe_1_6_3_U79 ( .A(pe_1_6_3_int_q_reg_v[23]), .B(
        pe_1_6_3_int_q_reg_v[19]), .S(pe_1_6_3_n55), .Z(pe_1_6_3_n18) );
  MUX2_X1 pe_1_6_3_U78 ( .A(pe_1_6_3_int_q_reg_v[15]), .B(
        pe_1_6_3_int_q_reg_v[11]), .S(pe_1_6_3_n55), .Z(pe_1_6_3_n17) );
  MUX2_X1 pe_1_6_3_U77 ( .A(pe_1_6_3_int_q_reg_v[7]), .B(
        pe_1_6_3_int_q_reg_v[3]), .S(pe_1_6_3_n55), .Z(pe_1_6_3_n16) );
  MUX2_X1 pe_1_6_3_U76 ( .A(pe_1_6_3_n15), .B(pe_1_6_3_n12), .S(n53), .Z(
        int_data_y_6__3__2_) );
  MUX2_X1 pe_1_6_3_U75 ( .A(pe_1_6_3_n14), .B(pe_1_6_3_n13), .S(pe_1_6_3_n61), 
        .Z(pe_1_6_3_n15) );
  MUX2_X1 pe_1_6_3_U74 ( .A(pe_1_6_3_int_q_reg_v[22]), .B(
        pe_1_6_3_int_q_reg_v[18]), .S(pe_1_6_3_n55), .Z(pe_1_6_3_n14) );
  MUX2_X1 pe_1_6_3_U73 ( .A(pe_1_6_3_int_q_reg_v[14]), .B(
        pe_1_6_3_int_q_reg_v[10]), .S(pe_1_6_3_n55), .Z(pe_1_6_3_n13) );
  MUX2_X1 pe_1_6_3_U72 ( .A(pe_1_6_3_int_q_reg_v[6]), .B(
        pe_1_6_3_int_q_reg_v[2]), .S(pe_1_6_3_n55), .Z(pe_1_6_3_n12) );
  MUX2_X1 pe_1_6_3_U71 ( .A(pe_1_6_3_n11), .B(pe_1_6_3_n8), .S(n53), .Z(
        int_data_y_6__3__1_) );
  MUX2_X1 pe_1_6_3_U70 ( .A(pe_1_6_3_n10), .B(pe_1_6_3_n9), .S(pe_1_6_3_n61), 
        .Z(pe_1_6_3_n11) );
  MUX2_X1 pe_1_6_3_U69 ( .A(pe_1_6_3_int_q_reg_v[21]), .B(
        pe_1_6_3_int_q_reg_v[17]), .S(pe_1_6_3_n55), .Z(pe_1_6_3_n10) );
  MUX2_X1 pe_1_6_3_U68 ( .A(pe_1_6_3_int_q_reg_v[13]), .B(
        pe_1_6_3_int_q_reg_v[9]), .S(pe_1_6_3_n55), .Z(pe_1_6_3_n9) );
  MUX2_X1 pe_1_6_3_U67 ( .A(pe_1_6_3_int_q_reg_v[5]), .B(
        pe_1_6_3_int_q_reg_v[1]), .S(pe_1_6_3_n55), .Z(pe_1_6_3_n8) );
  MUX2_X1 pe_1_6_3_U66 ( .A(pe_1_6_3_n7), .B(pe_1_6_3_n4), .S(n53), .Z(
        int_data_y_6__3__0_) );
  MUX2_X1 pe_1_6_3_U65 ( .A(pe_1_6_3_n6), .B(pe_1_6_3_n5), .S(pe_1_6_3_n61), 
        .Z(pe_1_6_3_n7) );
  MUX2_X1 pe_1_6_3_U64 ( .A(pe_1_6_3_int_q_reg_v[20]), .B(
        pe_1_6_3_int_q_reg_v[16]), .S(pe_1_6_3_n55), .Z(pe_1_6_3_n6) );
  MUX2_X1 pe_1_6_3_U63 ( .A(pe_1_6_3_int_q_reg_v[12]), .B(
        pe_1_6_3_int_q_reg_v[8]), .S(pe_1_6_3_n55), .Z(pe_1_6_3_n5) );
  MUX2_X1 pe_1_6_3_U62 ( .A(pe_1_6_3_int_q_reg_v[4]), .B(
        pe_1_6_3_int_q_reg_v[0]), .S(pe_1_6_3_n55), .Z(pe_1_6_3_n4) );
  AOI222_X1 pe_1_6_3_U61 ( .A1(int_data_res_7__3__2_), .A2(pe_1_6_3_n63), .B1(
        pe_1_6_3_N80), .B2(pe_1_6_3_n27), .C1(pe_1_6_3_N72), .C2(pe_1_6_3_n28), 
        .ZN(pe_1_6_3_n33) );
  INV_X1 pe_1_6_3_U60 ( .A(pe_1_6_3_n33), .ZN(pe_1_6_3_n80) );
  AOI222_X1 pe_1_6_3_U59 ( .A1(int_data_res_7__3__6_), .A2(pe_1_6_3_n63), .B1(
        pe_1_6_3_N84), .B2(pe_1_6_3_n27), .C1(pe_1_6_3_N76), .C2(pe_1_6_3_n28), 
        .ZN(pe_1_6_3_n29) );
  INV_X1 pe_1_6_3_U58 ( .A(pe_1_6_3_n29), .ZN(pe_1_6_3_n76) );
  XNOR2_X1 pe_1_6_3_U57 ( .A(pe_1_6_3_n71), .B(int_data_res_6__3__0_), .ZN(
        pe_1_6_3_N70) );
  AOI222_X1 pe_1_6_3_U52 ( .A1(int_data_res_7__3__0_), .A2(pe_1_6_3_n63), .B1(
        pe_1_6_3_n1), .B2(pe_1_6_3_n27), .C1(pe_1_6_3_N70), .C2(pe_1_6_3_n28), 
        .ZN(pe_1_6_3_n35) );
  INV_X1 pe_1_6_3_U51 ( .A(pe_1_6_3_n35), .ZN(pe_1_6_3_n82) );
  AOI222_X1 pe_1_6_3_U50 ( .A1(int_data_res_7__3__1_), .A2(pe_1_6_3_n63), .B1(
        pe_1_6_3_N79), .B2(pe_1_6_3_n27), .C1(pe_1_6_3_N71), .C2(pe_1_6_3_n28), 
        .ZN(pe_1_6_3_n34) );
  INV_X1 pe_1_6_3_U49 ( .A(pe_1_6_3_n34), .ZN(pe_1_6_3_n81) );
  AOI222_X1 pe_1_6_3_U48 ( .A1(int_data_res_7__3__3_), .A2(pe_1_6_3_n63), .B1(
        pe_1_6_3_N81), .B2(pe_1_6_3_n27), .C1(pe_1_6_3_N73), .C2(pe_1_6_3_n28), 
        .ZN(pe_1_6_3_n32) );
  INV_X1 pe_1_6_3_U47 ( .A(pe_1_6_3_n32), .ZN(pe_1_6_3_n79) );
  AOI222_X1 pe_1_6_3_U46 ( .A1(int_data_res_7__3__4_), .A2(pe_1_6_3_n63), .B1(
        pe_1_6_3_N82), .B2(pe_1_6_3_n27), .C1(pe_1_6_3_N74), .C2(pe_1_6_3_n28), 
        .ZN(pe_1_6_3_n31) );
  INV_X1 pe_1_6_3_U45 ( .A(pe_1_6_3_n31), .ZN(pe_1_6_3_n78) );
  AOI222_X1 pe_1_6_3_U44 ( .A1(int_data_res_7__3__5_), .A2(pe_1_6_3_n63), .B1(
        pe_1_6_3_N83), .B2(pe_1_6_3_n27), .C1(pe_1_6_3_N75), .C2(pe_1_6_3_n28), 
        .ZN(pe_1_6_3_n30) );
  INV_X1 pe_1_6_3_U43 ( .A(pe_1_6_3_n30), .ZN(pe_1_6_3_n77) );
  NAND2_X1 pe_1_6_3_U42 ( .A1(pe_1_6_3_int_data_0_), .A2(pe_1_6_3_n3), .ZN(
        pe_1_6_3_sub_81_carry[1]) );
  INV_X1 pe_1_6_3_U41 ( .A(pe_1_6_3_int_data_1_), .ZN(pe_1_6_3_n72) );
  INV_X1 pe_1_6_3_U40 ( .A(pe_1_6_3_int_data_2_), .ZN(pe_1_6_3_n73) );
  AND2_X1 pe_1_6_3_U39 ( .A1(pe_1_6_3_int_data_0_), .A2(int_data_res_6__3__0_), 
        .ZN(pe_1_6_3_n2) );
  AOI222_X1 pe_1_6_3_U38 ( .A1(pe_1_6_3_n63), .A2(int_data_res_7__3__7_), .B1(
        pe_1_6_3_N85), .B2(pe_1_6_3_n27), .C1(pe_1_6_3_N77), .C2(pe_1_6_3_n28), 
        .ZN(pe_1_6_3_n26) );
  INV_X1 pe_1_6_3_U37 ( .A(pe_1_6_3_n26), .ZN(pe_1_6_3_n75) );
  NOR3_X1 pe_1_6_3_U36 ( .A1(pe_1_6_3_n58), .A2(pe_1_6_3_n64), .A3(int_ckg[12]), .ZN(pe_1_6_3_n36) );
  OR2_X1 pe_1_6_3_U35 ( .A1(pe_1_6_3_n36), .A2(pe_1_6_3_n63), .ZN(pe_1_6_3_N90) );
  INV_X1 pe_1_6_3_U34 ( .A(n41), .ZN(pe_1_6_3_n62) );
  AND2_X1 pe_1_6_3_U33 ( .A1(int_data_x_6__3__2_), .A2(n29), .ZN(
        pe_1_6_3_int_data_2_) );
  AND2_X1 pe_1_6_3_U32 ( .A1(int_data_x_6__3__1_), .A2(n29), .ZN(
        pe_1_6_3_int_data_1_) );
  AND2_X1 pe_1_6_3_U31 ( .A1(int_data_x_6__3__3_), .A2(n29), .ZN(
        pe_1_6_3_int_data_3_) );
  BUF_X1 pe_1_6_3_U30 ( .A(n63), .Z(pe_1_6_3_n63) );
  INV_X1 pe_1_6_3_U29 ( .A(n35), .ZN(pe_1_6_3_n60) );
  AND2_X1 pe_1_6_3_U28 ( .A1(int_data_x_6__3__0_), .A2(n29), .ZN(
        pe_1_6_3_int_data_0_) );
  NAND2_X1 pe_1_6_3_U27 ( .A1(pe_1_6_3_n44), .A2(pe_1_6_3_n60), .ZN(
        pe_1_6_3_n41) );
  AND3_X1 pe_1_6_3_U26 ( .A1(n77), .A2(pe_1_6_3_n62), .A3(n53), .ZN(
        pe_1_6_3_n44) );
  INV_X1 pe_1_6_3_U25 ( .A(pe_1_6_3_int_data_3_), .ZN(pe_1_6_3_n74) );
  NOR2_X1 pe_1_6_3_U24 ( .A1(pe_1_6_3_n68), .A2(n53), .ZN(pe_1_6_3_n43) );
  NOR2_X1 pe_1_6_3_U23 ( .A1(pe_1_6_3_n57), .A2(pe_1_6_3_n63), .ZN(
        pe_1_6_3_n28) );
  NOR2_X1 pe_1_6_3_U22 ( .A1(n21), .A2(pe_1_6_3_n63), .ZN(pe_1_6_3_n27) );
  INV_X1 pe_1_6_3_U21 ( .A(pe_1_6_3_int_data_0_), .ZN(pe_1_6_3_n71) );
  INV_X1 pe_1_6_3_U20 ( .A(pe_1_6_3_n41), .ZN(pe_1_6_3_n88) );
  INV_X1 pe_1_6_3_U19 ( .A(pe_1_6_3_n37), .ZN(pe_1_6_3_n86) );
  INV_X1 pe_1_6_3_U18 ( .A(pe_1_6_3_n38), .ZN(pe_1_6_3_n85) );
  INV_X1 pe_1_6_3_U17 ( .A(pe_1_6_3_n39), .ZN(pe_1_6_3_n84) );
  NOR2_X1 pe_1_6_3_U16 ( .A1(pe_1_6_3_n66), .A2(pe_1_6_3_n42), .ZN(
        pe_1_6_3_N59) );
  NOR2_X1 pe_1_6_3_U15 ( .A1(pe_1_6_3_n66), .A2(pe_1_6_3_n41), .ZN(
        pe_1_6_3_N60) );
  NOR2_X1 pe_1_6_3_U14 ( .A1(pe_1_6_3_n66), .A2(pe_1_6_3_n38), .ZN(
        pe_1_6_3_N63) );
  NOR2_X1 pe_1_6_3_U13 ( .A1(pe_1_6_3_n66), .A2(pe_1_6_3_n40), .ZN(
        pe_1_6_3_N61) );
  NOR2_X1 pe_1_6_3_U12 ( .A1(pe_1_6_3_n66), .A2(pe_1_6_3_n39), .ZN(
        pe_1_6_3_N62) );
  NOR2_X1 pe_1_6_3_U11 ( .A1(pe_1_6_3_n37), .A2(pe_1_6_3_n66), .ZN(
        pe_1_6_3_N64) );
  NAND2_X1 pe_1_6_3_U10 ( .A1(pe_1_6_3_n44), .A2(pe_1_6_3_n59), .ZN(
        pe_1_6_3_n42) );
  BUF_X1 pe_1_6_3_U9 ( .A(pe_1_6_3_n59), .Z(pe_1_6_3_n55) );
  INV_X1 pe_1_6_3_U8 ( .A(pe_1_6_3_n67), .ZN(pe_1_6_3_n64) );
  BUF_X1 pe_1_6_3_U7 ( .A(pe_1_6_3_n59), .Z(pe_1_6_3_n56) );
  INV_X1 pe_1_6_3_U6 ( .A(pe_1_6_3_n42), .ZN(pe_1_6_3_n87) );
  INV_X1 pe_1_6_3_U5 ( .A(pe_1_6_3_n40), .ZN(pe_1_6_3_n83) );
  INV_X2 pe_1_6_3_U4 ( .A(n85), .ZN(pe_1_6_3_n70) );
  XOR2_X1 pe_1_6_3_U3 ( .A(pe_1_6_3_int_data_0_), .B(int_data_res_6__3__0_), 
        .Z(pe_1_6_3_n1) );
  DFFR_X1 pe_1_6_3_int_q_acc_reg_0_ ( .D(pe_1_6_3_n82), .CK(pe_1_6_3_net3574), 
        .RN(pe_1_6_3_n70), .Q(int_data_res_6__3__0_), .QN(pe_1_6_3_n3) );
  DFFR_X1 pe_1_6_3_int_q_reg_v_reg_0__0_ ( .D(int_data_y_7__3__0_), .CK(
        pe_1_6_3_net3544), .RN(pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_v[20]) );
  DFFR_X1 pe_1_6_3_int_q_reg_v_reg_0__1_ ( .D(int_data_y_7__3__1_), .CK(
        pe_1_6_3_net3544), .RN(pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_v[21]) );
  DFFR_X1 pe_1_6_3_int_q_reg_v_reg_0__2_ ( .D(int_data_y_7__3__2_), .CK(
        pe_1_6_3_net3544), .RN(pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_v[22]) );
  DFFR_X1 pe_1_6_3_int_q_reg_v_reg_0__3_ ( .D(int_data_y_7__3__3_), .CK(
        pe_1_6_3_net3544), .RN(pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_v[23]) );
  DFFR_X1 pe_1_6_3_int_q_reg_v_reg_1__0_ ( .D(int_data_y_7__3__0_), .CK(
        pe_1_6_3_net3549), .RN(pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_v[16]) );
  DFFR_X1 pe_1_6_3_int_q_reg_v_reg_1__1_ ( .D(int_data_y_7__3__1_), .CK(
        pe_1_6_3_net3549), .RN(pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_v[17]) );
  DFFR_X1 pe_1_6_3_int_q_reg_v_reg_1__2_ ( .D(int_data_y_7__3__2_), .CK(
        pe_1_6_3_net3549), .RN(pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_v[18]) );
  DFFR_X1 pe_1_6_3_int_q_reg_v_reg_1__3_ ( .D(int_data_y_7__3__3_), .CK(
        pe_1_6_3_net3549), .RN(pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_v[19]) );
  DFFR_X1 pe_1_6_3_int_q_reg_v_reg_2__0_ ( .D(int_data_y_7__3__0_), .CK(
        pe_1_6_3_net3554), .RN(pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_v[12]) );
  DFFR_X1 pe_1_6_3_int_q_reg_v_reg_2__1_ ( .D(int_data_y_7__3__1_), .CK(
        pe_1_6_3_net3554), .RN(pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_v[13]) );
  DFFR_X1 pe_1_6_3_int_q_reg_v_reg_2__2_ ( .D(int_data_y_7__3__2_), .CK(
        pe_1_6_3_net3554), .RN(pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_v[14]) );
  DFFR_X1 pe_1_6_3_int_q_reg_v_reg_2__3_ ( .D(int_data_y_7__3__3_), .CK(
        pe_1_6_3_net3554), .RN(pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_v[15]) );
  DFFR_X1 pe_1_6_3_int_q_reg_v_reg_3__0_ ( .D(int_data_y_7__3__0_), .CK(
        pe_1_6_3_net3559), .RN(pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_v[8]) );
  DFFR_X1 pe_1_6_3_int_q_reg_v_reg_3__1_ ( .D(int_data_y_7__3__1_), .CK(
        pe_1_6_3_net3559), .RN(pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_v[9]) );
  DFFR_X1 pe_1_6_3_int_q_reg_v_reg_3__2_ ( .D(int_data_y_7__3__2_), .CK(
        pe_1_6_3_net3559), .RN(pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_v[10]) );
  DFFR_X1 pe_1_6_3_int_q_reg_v_reg_3__3_ ( .D(int_data_y_7__3__3_), .CK(
        pe_1_6_3_net3559), .RN(pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_v[11]) );
  DFFR_X1 pe_1_6_3_int_q_reg_v_reg_4__0_ ( .D(int_data_y_7__3__0_), .CK(
        pe_1_6_3_net3564), .RN(pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_v[4]) );
  DFFR_X1 pe_1_6_3_int_q_reg_v_reg_4__1_ ( .D(int_data_y_7__3__1_), .CK(
        pe_1_6_3_net3564), .RN(pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_v[5]) );
  DFFR_X1 pe_1_6_3_int_q_reg_v_reg_4__2_ ( .D(int_data_y_7__3__2_), .CK(
        pe_1_6_3_net3564), .RN(pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_v[6]) );
  DFFR_X1 pe_1_6_3_int_q_reg_v_reg_4__3_ ( .D(int_data_y_7__3__3_), .CK(
        pe_1_6_3_net3564), .RN(pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_v[7]) );
  DFFR_X1 pe_1_6_3_int_q_reg_v_reg_5__0_ ( .D(int_data_y_7__3__0_), .CK(
        pe_1_6_3_net3569), .RN(pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_v[0]) );
  DFFR_X1 pe_1_6_3_int_q_reg_v_reg_5__1_ ( .D(int_data_y_7__3__1_), .CK(
        pe_1_6_3_net3569), .RN(pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_v[1]) );
  DFFR_X1 pe_1_6_3_int_q_reg_v_reg_5__2_ ( .D(int_data_y_7__3__2_), .CK(
        pe_1_6_3_net3569), .RN(pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_v[2]) );
  DFFR_X1 pe_1_6_3_int_q_reg_v_reg_5__3_ ( .D(int_data_y_7__3__3_), .CK(
        pe_1_6_3_net3569), .RN(pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_6_3_int_q_reg_h_reg_0__0_ ( .D(int_data_x_6__4__0_), .SI(
        int_data_y_7__3__0_), .SE(pe_1_6_3_n64), .CK(pe_1_6_3_net3513), .RN(
        pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_6_3_int_q_reg_h_reg_0__1_ ( .D(int_data_x_6__4__1_), .SI(
        int_data_y_7__3__1_), .SE(pe_1_6_3_n64), .CK(pe_1_6_3_net3513), .RN(
        pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_6_3_int_q_reg_h_reg_0__2_ ( .D(int_data_x_6__4__2_), .SI(
        int_data_y_7__3__2_), .SE(pe_1_6_3_n64), .CK(pe_1_6_3_net3513), .RN(
        pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_6_3_int_q_reg_h_reg_0__3_ ( .D(int_data_x_6__4__3_), .SI(
        int_data_y_7__3__3_), .SE(pe_1_6_3_n64), .CK(pe_1_6_3_net3513), .RN(
        pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_6_3_int_q_reg_h_reg_1__0_ ( .D(int_data_x_6__4__0_), .SI(
        int_data_y_7__3__0_), .SE(pe_1_6_3_n64), .CK(pe_1_6_3_net3519), .RN(
        pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_6_3_int_q_reg_h_reg_1__1_ ( .D(int_data_x_6__4__1_), .SI(
        int_data_y_7__3__1_), .SE(pe_1_6_3_n64), .CK(pe_1_6_3_net3519), .RN(
        pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_6_3_int_q_reg_h_reg_1__2_ ( .D(int_data_x_6__4__2_), .SI(
        int_data_y_7__3__2_), .SE(pe_1_6_3_n64), .CK(pe_1_6_3_net3519), .RN(
        pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_6_3_int_q_reg_h_reg_1__3_ ( .D(int_data_x_6__4__3_), .SI(
        int_data_y_7__3__3_), .SE(pe_1_6_3_n64), .CK(pe_1_6_3_net3519), .RN(
        pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_6_3_int_q_reg_h_reg_2__0_ ( .D(int_data_x_6__4__0_), .SI(
        int_data_y_7__3__0_), .SE(pe_1_6_3_n64), .CK(pe_1_6_3_net3524), .RN(
        pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_6_3_int_q_reg_h_reg_2__1_ ( .D(int_data_x_6__4__1_), .SI(
        int_data_y_7__3__1_), .SE(pe_1_6_3_n64), .CK(pe_1_6_3_net3524), .RN(
        pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_6_3_int_q_reg_h_reg_2__2_ ( .D(int_data_x_6__4__2_), .SI(
        int_data_y_7__3__2_), .SE(pe_1_6_3_n64), .CK(pe_1_6_3_net3524), .RN(
        pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_6_3_int_q_reg_h_reg_2__3_ ( .D(int_data_x_6__4__3_), .SI(
        int_data_y_7__3__3_), .SE(pe_1_6_3_n64), .CK(pe_1_6_3_net3524), .RN(
        pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_6_3_int_q_reg_h_reg_3__0_ ( .D(int_data_x_6__4__0_), .SI(
        int_data_y_7__3__0_), .SE(pe_1_6_3_n64), .CK(pe_1_6_3_net3529), .RN(
        pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_6_3_int_q_reg_h_reg_3__1_ ( .D(int_data_x_6__4__1_), .SI(
        int_data_y_7__3__1_), .SE(pe_1_6_3_n64), .CK(pe_1_6_3_net3529), .RN(
        pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_6_3_int_q_reg_h_reg_3__2_ ( .D(int_data_x_6__4__2_), .SI(
        int_data_y_7__3__2_), .SE(pe_1_6_3_n64), .CK(pe_1_6_3_net3529), .RN(
        pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_6_3_int_q_reg_h_reg_3__3_ ( .D(int_data_x_6__4__3_), .SI(
        int_data_y_7__3__3_), .SE(pe_1_6_3_n64), .CK(pe_1_6_3_net3529), .RN(
        pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_6_3_int_q_reg_h_reg_4__0_ ( .D(int_data_x_6__4__0_), .SI(
        int_data_y_7__3__0_), .SE(pe_1_6_3_n65), .CK(pe_1_6_3_net3534), .RN(
        pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_6_3_int_q_reg_h_reg_4__1_ ( .D(int_data_x_6__4__1_), .SI(
        int_data_y_7__3__1_), .SE(pe_1_6_3_n65), .CK(pe_1_6_3_net3534), .RN(
        pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_6_3_int_q_reg_h_reg_4__2_ ( .D(int_data_x_6__4__2_), .SI(
        int_data_y_7__3__2_), .SE(pe_1_6_3_n65), .CK(pe_1_6_3_net3534), .RN(
        pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_6_3_int_q_reg_h_reg_4__3_ ( .D(int_data_x_6__4__3_), .SI(
        int_data_y_7__3__3_), .SE(pe_1_6_3_n65), .CK(pe_1_6_3_net3534), .RN(
        pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_6_3_int_q_reg_h_reg_5__0_ ( .D(int_data_x_6__4__0_), .SI(
        int_data_y_7__3__0_), .SE(pe_1_6_3_n65), .CK(pe_1_6_3_net3539), .RN(
        pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_6_3_int_q_reg_h_reg_5__1_ ( .D(int_data_x_6__4__1_), .SI(
        int_data_y_7__3__1_), .SE(pe_1_6_3_n65), .CK(pe_1_6_3_net3539), .RN(
        pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_6_3_int_q_reg_h_reg_5__2_ ( .D(int_data_x_6__4__2_), .SI(
        int_data_y_7__3__2_), .SE(pe_1_6_3_n65), .CK(pe_1_6_3_net3539), .RN(
        pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_6_3_int_q_reg_h_reg_5__3_ ( .D(int_data_x_6__4__3_), .SI(
        int_data_y_7__3__3_), .SE(pe_1_6_3_n65), .CK(pe_1_6_3_net3539), .RN(
        pe_1_6_3_n70), .Q(pe_1_6_3_int_q_reg_h[3]) );
  FA_X1 pe_1_6_3_sub_81_U2_7 ( .A(int_data_res_6__3__7_), .B(pe_1_6_3_n74), 
        .CI(pe_1_6_3_sub_81_carry[7]), .S(pe_1_6_3_N77) );
  FA_X1 pe_1_6_3_sub_81_U2_6 ( .A(int_data_res_6__3__6_), .B(pe_1_6_3_n74), 
        .CI(pe_1_6_3_sub_81_carry[6]), .CO(pe_1_6_3_sub_81_carry[7]), .S(
        pe_1_6_3_N76) );
  FA_X1 pe_1_6_3_sub_81_U2_5 ( .A(int_data_res_6__3__5_), .B(pe_1_6_3_n74), 
        .CI(pe_1_6_3_sub_81_carry[5]), .CO(pe_1_6_3_sub_81_carry[6]), .S(
        pe_1_6_3_N75) );
  FA_X1 pe_1_6_3_sub_81_U2_4 ( .A(int_data_res_6__3__4_), .B(pe_1_6_3_n74), 
        .CI(pe_1_6_3_sub_81_carry[4]), .CO(pe_1_6_3_sub_81_carry[5]), .S(
        pe_1_6_3_N74) );
  FA_X1 pe_1_6_3_sub_81_U2_3 ( .A(int_data_res_6__3__3_), .B(pe_1_6_3_n74), 
        .CI(pe_1_6_3_sub_81_carry[3]), .CO(pe_1_6_3_sub_81_carry[4]), .S(
        pe_1_6_3_N73) );
  FA_X1 pe_1_6_3_sub_81_U2_2 ( .A(int_data_res_6__3__2_), .B(pe_1_6_3_n73), 
        .CI(pe_1_6_3_sub_81_carry[2]), .CO(pe_1_6_3_sub_81_carry[3]), .S(
        pe_1_6_3_N72) );
  FA_X1 pe_1_6_3_sub_81_U2_1 ( .A(int_data_res_6__3__1_), .B(pe_1_6_3_n72), 
        .CI(pe_1_6_3_sub_81_carry[1]), .CO(pe_1_6_3_sub_81_carry[2]), .S(
        pe_1_6_3_N71) );
  FA_X1 pe_1_6_3_add_83_U1_7 ( .A(int_data_res_6__3__7_), .B(
        pe_1_6_3_int_data_3_), .CI(pe_1_6_3_add_83_carry[7]), .S(pe_1_6_3_N85)
         );
  FA_X1 pe_1_6_3_add_83_U1_6 ( .A(int_data_res_6__3__6_), .B(
        pe_1_6_3_int_data_3_), .CI(pe_1_6_3_add_83_carry[6]), .CO(
        pe_1_6_3_add_83_carry[7]), .S(pe_1_6_3_N84) );
  FA_X1 pe_1_6_3_add_83_U1_5 ( .A(int_data_res_6__3__5_), .B(
        pe_1_6_3_int_data_3_), .CI(pe_1_6_3_add_83_carry[5]), .CO(
        pe_1_6_3_add_83_carry[6]), .S(pe_1_6_3_N83) );
  FA_X1 pe_1_6_3_add_83_U1_4 ( .A(int_data_res_6__3__4_), .B(
        pe_1_6_3_int_data_3_), .CI(pe_1_6_3_add_83_carry[4]), .CO(
        pe_1_6_3_add_83_carry[5]), .S(pe_1_6_3_N82) );
  FA_X1 pe_1_6_3_add_83_U1_3 ( .A(int_data_res_6__3__3_), .B(
        pe_1_6_3_int_data_3_), .CI(pe_1_6_3_add_83_carry[3]), .CO(
        pe_1_6_3_add_83_carry[4]), .S(pe_1_6_3_N81) );
  FA_X1 pe_1_6_3_add_83_U1_2 ( .A(int_data_res_6__3__2_), .B(
        pe_1_6_3_int_data_2_), .CI(pe_1_6_3_add_83_carry[2]), .CO(
        pe_1_6_3_add_83_carry[3]), .S(pe_1_6_3_N80) );
  FA_X1 pe_1_6_3_add_83_U1_1 ( .A(int_data_res_6__3__1_), .B(
        pe_1_6_3_int_data_1_), .CI(pe_1_6_3_n2), .CO(pe_1_6_3_add_83_carry[2]), 
        .S(pe_1_6_3_N79) );
  NAND3_X1 pe_1_6_3_U56 ( .A1(pe_1_6_3_n59), .A2(pe_1_6_3_n43), .A3(
        pe_1_6_3_n61), .ZN(pe_1_6_3_n40) );
  NAND3_X1 pe_1_6_3_U55 ( .A1(pe_1_6_3_n43), .A2(pe_1_6_3_n60), .A3(
        pe_1_6_3_n61), .ZN(pe_1_6_3_n39) );
  NAND3_X1 pe_1_6_3_U54 ( .A1(pe_1_6_3_n43), .A2(pe_1_6_3_n62), .A3(
        pe_1_6_3_n59), .ZN(pe_1_6_3_n38) );
  NAND3_X1 pe_1_6_3_U53 ( .A1(pe_1_6_3_n60), .A2(pe_1_6_3_n62), .A3(
        pe_1_6_3_n43), .ZN(pe_1_6_3_n37) );
  DFFR_X1 pe_1_6_3_int_q_acc_reg_6_ ( .D(pe_1_6_3_n76), .CK(pe_1_6_3_net3574), 
        .RN(pe_1_6_3_n69), .Q(int_data_res_6__3__6_) );
  DFFR_X1 pe_1_6_3_int_q_acc_reg_5_ ( .D(pe_1_6_3_n77), .CK(pe_1_6_3_net3574), 
        .RN(pe_1_6_3_n69), .Q(int_data_res_6__3__5_) );
  DFFR_X1 pe_1_6_3_int_q_acc_reg_4_ ( .D(pe_1_6_3_n78), .CK(pe_1_6_3_net3574), 
        .RN(pe_1_6_3_n69), .Q(int_data_res_6__3__4_) );
  DFFR_X1 pe_1_6_3_int_q_acc_reg_3_ ( .D(pe_1_6_3_n79), .CK(pe_1_6_3_net3574), 
        .RN(pe_1_6_3_n69), .Q(int_data_res_6__3__3_) );
  DFFR_X1 pe_1_6_3_int_q_acc_reg_2_ ( .D(pe_1_6_3_n80), .CK(pe_1_6_3_net3574), 
        .RN(pe_1_6_3_n69), .Q(int_data_res_6__3__2_) );
  DFFR_X1 pe_1_6_3_int_q_acc_reg_1_ ( .D(pe_1_6_3_n81), .CK(pe_1_6_3_net3574), 
        .RN(pe_1_6_3_n69), .Q(int_data_res_6__3__1_) );
  DFFR_X1 pe_1_6_3_int_q_acc_reg_7_ ( .D(pe_1_6_3_n75), .CK(pe_1_6_3_net3574), 
        .RN(pe_1_6_3_n69), .Q(int_data_res_6__3__7_) );
  CLKGATETST_X1 pe_1_6_3_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_6_3_n86), .SE(1'b0), .GCK(pe_1_6_3_net3513) );
  CLKGATETST_X1 pe_1_6_3_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_6_3_n85), .SE(1'b0), .GCK(pe_1_6_3_net3519) );
  CLKGATETST_X1 pe_1_6_3_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_6_3_n84), .SE(1'b0), .GCK(pe_1_6_3_net3524) );
  CLKGATETST_X1 pe_1_6_3_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_6_3_n83), .SE(1'b0), .GCK(pe_1_6_3_net3529) );
  CLKGATETST_X1 pe_1_6_3_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_6_3_n88), .SE(1'b0), .GCK(pe_1_6_3_net3534) );
  CLKGATETST_X1 pe_1_6_3_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_6_3_n87), .SE(1'b0), .GCK(pe_1_6_3_net3539) );
  CLKGATETST_X1 pe_1_6_3_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_6_3_N64), .SE(1'b0), .GCK(pe_1_6_3_net3544) );
  CLKGATETST_X1 pe_1_6_3_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_6_3_N63), .SE(1'b0), .GCK(pe_1_6_3_net3549) );
  CLKGATETST_X1 pe_1_6_3_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_6_3_N62), .SE(1'b0), .GCK(pe_1_6_3_net3554) );
  CLKGATETST_X1 pe_1_6_3_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_6_3_N61), .SE(1'b0), .GCK(pe_1_6_3_net3559) );
  CLKGATETST_X1 pe_1_6_3_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_6_3_N60), .SE(1'b0), .GCK(pe_1_6_3_net3564) );
  CLKGATETST_X1 pe_1_6_3_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_6_3_N59), .SE(1'b0), .GCK(pe_1_6_3_net3569) );
  CLKGATETST_X1 pe_1_6_3_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_6_3_N90), .SE(1'b0), .GCK(pe_1_6_3_net3574) );
  CLKBUF_X1 pe_1_6_4_U112 ( .A(pe_1_6_4_n72), .Z(pe_1_6_4_n71) );
  INV_X1 pe_1_6_4_U111 ( .A(n77), .ZN(pe_1_6_4_n70) );
  INV_X1 pe_1_6_4_U110 ( .A(n69), .ZN(pe_1_6_4_n69) );
  INV_X1 pe_1_6_4_U109 ( .A(n69), .ZN(pe_1_6_4_n68) );
  INV_X1 pe_1_6_4_U108 ( .A(n69), .ZN(pe_1_6_4_n67) );
  INV_X1 pe_1_6_4_U107 ( .A(pe_1_6_4_n69), .ZN(pe_1_6_4_n66) );
  INV_X1 pe_1_6_4_U106 ( .A(pe_1_6_4_n63), .ZN(pe_1_6_4_n62) );
  INV_X1 pe_1_6_4_U105 ( .A(pe_1_6_4_n61), .ZN(pe_1_6_4_n60) );
  INV_X1 pe_1_6_4_U104 ( .A(n29), .ZN(pe_1_6_4_n59) );
  INV_X1 pe_1_6_4_U103 ( .A(pe_1_6_4_n59), .ZN(pe_1_6_4_n58) );
  INV_X1 pe_1_6_4_U102 ( .A(n21), .ZN(pe_1_6_4_n57) );
  MUX2_X1 pe_1_6_4_U101 ( .A(pe_1_6_4_n54), .B(pe_1_6_4_n51), .S(n53), .Z(
        int_data_x_6__4__3_) );
  MUX2_X1 pe_1_6_4_U100 ( .A(pe_1_6_4_n53), .B(pe_1_6_4_n52), .S(pe_1_6_4_n62), 
        .Z(pe_1_6_4_n54) );
  MUX2_X1 pe_1_6_4_U99 ( .A(pe_1_6_4_int_q_reg_h[23]), .B(
        pe_1_6_4_int_q_reg_h[19]), .S(pe_1_6_4_n56), .Z(pe_1_6_4_n53) );
  MUX2_X1 pe_1_6_4_U98 ( .A(pe_1_6_4_int_q_reg_h[15]), .B(
        pe_1_6_4_int_q_reg_h[11]), .S(pe_1_6_4_n56), .Z(pe_1_6_4_n52) );
  MUX2_X1 pe_1_6_4_U97 ( .A(pe_1_6_4_int_q_reg_h[7]), .B(
        pe_1_6_4_int_q_reg_h[3]), .S(pe_1_6_4_n56), .Z(pe_1_6_4_n51) );
  MUX2_X1 pe_1_6_4_U96 ( .A(pe_1_6_4_n50), .B(pe_1_6_4_n47), .S(n53), .Z(
        int_data_x_6__4__2_) );
  MUX2_X1 pe_1_6_4_U95 ( .A(pe_1_6_4_n49), .B(pe_1_6_4_n48), .S(pe_1_6_4_n62), 
        .Z(pe_1_6_4_n50) );
  MUX2_X1 pe_1_6_4_U94 ( .A(pe_1_6_4_int_q_reg_h[22]), .B(
        pe_1_6_4_int_q_reg_h[18]), .S(pe_1_6_4_n56), .Z(pe_1_6_4_n49) );
  MUX2_X1 pe_1_6_4_U93 ( .A(pe_1_6_4_int_q_reg_h[14]), .B(
        pe_1_6_4_int_q_reg_h[10]), .S(pe_1_6_4_n56), .Z(pe_1_6_4_n48) );
  MUX2_X1 pe_1_6_4_U92 ( .A(pe_1_6_4_int_q_reg_h[6]), .B(
        pe_1_6_4_int_q_reg_h[2]), .S(pe_1_6_4_n56), .Z(pe_1_6_4_n47) );
  MUX2_X1 pe_1_6_4_U91 ( .A(pe_1_6_4_n46), .B(pe_1_6_4_n24), .S(n53), .Z(
        int_data_x_6__4__1_) );
  MUX2_X1 pe_1_6_4_U90 ( .A(pe_1_6_4_n45), .B(pe_1_6_4_n25), .S(pe_1_6_4_n62), 
        .Z(pe_1_6_4_n46) );
  MUX2_X1 pe_1_6_4_U89 ( .A(pe_1_6_4_int_q_reg_h[21]), .B(
        pe_1_6_4_int_q_reg_h[17]), .S(pe_1_6_4_n56), .Z(pe_1_6_4_n45) );
  MUX2_X1 pe_1_6_4_U88 ( .A(pe_1_6_4_int_q_reg_h[13]), .B(
        pe_1_6_4_int_q_reg_h[9]), .S(pe_1_6_4_n56), .Z(pe_1_6_4_n25) );
  MUX2_X1 pe_1_6_4_U87 ( .A(pe_1_6_4_int_q_reg_h[5]), .B(
        pe_1_6_4_int_q_reg_h[1]), .S(pe_1_6_4_n56), .Z(pe_1_6_4_n24) );
  MUX2_X1 pe_1_6_4_U86 ( .A(pe_1_6_4_n23), .B(pe_1_6_4_n20), .S(n53), .Z(
        int_data_x_6__4__0_) );
  MUX2_X1 pe_1_6_4_U85 ( .A(pe_1_6_4_n22), .B(pe_1_6_4_n21), .S(pe_1_6_4_n62), 
        .Z(pe_1_6_4_n23) );
  MUX2_X1 pe_1_6_4_U84 ( .A(pe_1_6_4_int_q_reg_h[20]), .B(
        pe_1_6_4_int_q_reg_h[16]), .S(pe_1_6_4_n56), .Z(pe_1_6_4_n22) );
  MUX2_X1 pe_1_6_4_U83 ( .A(pe_1_6_4_int_q_reg_h[12]), .B(
        pe_1_6_4_int_q_reg_h[8]), .S(pe_1_6_4_n56), .Z(pe_1_6_4_n21) );
  MUX2_X1 pe_1_6_4_U82 ( .A(pe_1_6_4_int_q_reg_h[4]), .B(
        pe_1_6_4_int_q_reg_h[0]), .S(pe_1_6_4_n56), .Z(pe_1_6_4_n20) );
  MUX2_X1 pe_1_6_4_U81 ( .A(pe_1_6_4_n19), .B(pe_1_6_4_n16), .S(n53), .Z(
        int_data_y_6__4__3_) );
  MUX2_X1 pe_1_6_4_U80 ( .A(pe_1_6_4_n18), .B(pe_1_6_4_n17), .S(pe_1_6_4_n62), 
        .Z(pe_1_6_4_n19) );
  MUX2_X1 pe_1_6_4_U79 ( .A(pe_1_6_4_int_q_reg_v[23]), .B(
        pe_1_6_4_int_q_reg_v[19]), .S(pe_1_6_4_n55), .Z(pe_1_6_4_n18) );
  MUX2_X1 pe_1_6_4_U78 ( .A(pe_1_6_4_int_q_reg_v[15]), .B(
        pe_1_6_4_int_q_reg_v[11]), .S(pe_1_6_4_n55), .Z(pe_1_6_4_n17) );
  MUX2_X1 pe_1_6_4_U77 ( .A(pe_1_6_4_int_q_reg_v[7]), .B(
        pe_1_6_4_int_q_reg_v[3]), .S(pe_1_6_4_n55), .Z(pe_1_6_4_n16) );
  MUX2_X1 pe_1_6_4_U76 ( .A(pe_1_6_4_n15), .B(pe_1_6_4_n12), .S(n53), .Z(
        int_data_y_6__4__2_) );
  MUX2_X1 pe_1_6_4_U75 ( .A(pe_1_6_4_n14), .B(pe_1_6_4_n13), .S(pe_1_6_4_n62), 
        .Z(pe_1_6_4_n15) );
  MUX2_X1 pe_1_6_4_U74 ( .A(pe_1_6_4_int_q_reg_v[22]), .B(
        pe_1_6_4_int_q_reg_v[18]), .S(pe_1_6_4_n55), .Z(pe_1_6_4_n14) );
  MUX2_X1 pe_1_6_4_U73 ( .A(pe_1_6_4_int_q_reg_v[14]), .B(
        pe_1_6_4_int_q_reg_v[10]), .S(pe_1_6_4_n55), .Z(pe_1_6_4_n13) );
  MUX2_X1 pe_1_6_4_U72 ( .A(pe_1_6_4_int_q_reg_v[6]), .B(
        pe_1_6_4_int_q_reg_v[2]), .S(pe_1_6_4_n55), .Z(pe_1_6_4_n12) );
  MUX2_X1 pe_1_6_4_U71 ( .A(pe_1_6_4_n11), .B(pe_1_6_4_n8), .S(n53), .Z(
        int_data_y_6__4__1_) );
  MUX2_X1 pe_1_6_4_U70 ( .A(pe_1_6_4_n10), .B(pe_1_6_4_n9), .S(pe_1_6_4_n62), 
        .Z(pe_1_6_4_n11) );
  MUX2_X1 pe_1_6_4_U69 ( .A(pe_1_6_4_int_q_reg_v[21]), .B(
        pe_1_6_4_int_q_reg_v[17]), .S(pe_1_6_4_n55), .Z(pe_1_6_4_n10) );
  MUX2_X1 pe_1_6_4_U68 ( .A(pe_1_6_4_int_q_reg_v[13]), .B(
        pe_1_6_4_int_q_reg_v[9]), .S(pe_1_6_4_n55), .Z(pe_1_6_4_n9) );
  MUX2_X1 pe_1_6_4_U67 ( .A(pe_1_6_4_int_q_reg_v[5]), .B(
        pe_1_6_4_int_q_reg_v[1]), .S(pe_1_6_4_n55), .Z(pe_1_6_4_n8) );
  MUX2_X1 pe_1_6_4_U66 ( .A(pe_1_6_4_n7), .B(pe_1_6_4_n4), .S(n53), .Z(
        int_data_y_6__4__0_) );
  MUX2_X1 pe_1_6_4_U65 ( .A(pe_1_6_4_n6), .B(pe_1_6_4_n5), .S(pe_1_6_4_n62), 
        .Z(pe_1_6_4_n7) );
  MUX2_X1 pe_1_6_4_U64 ( .A(pe_1_6_4_int_q_reg_v[20]), .B(
        pe_1_6_4_int_q_reg_v[16]), .S(pe_1_6_4_n55), .Z(pe_1_6_4_n6) );
  MUX2_X1 pe_1_6_4_U63 ( .A(pe_1_6_4_int_q_reg_v[12]), .B(
        pe_1_6_4_int_q_reg_v[8]), .S(pe_1_6_4_n55), .Z(pe_1_6_4_n5) );
  MUX2_X1 pe_1_6_4_U62 ( .A(pe_1_6_4_int_q_reg_v[4]), .B(
        pe_1_6_4_int_q_reg_v[0]), .S(pe_1_6_4_n55), .Z(pe_1_6_4_n4) );
  AOI222_X1 pe_1_6_4_U61 ( .A1(int_data_res_7__4__2_), .A2(pe_1_6_4_n64), .B1(
        pe_1_6_4_N80), .B2(pe_1_6_4_n27), .C1(pe_1_6_4_N72), .C2(pe_1_6_4_n28), 
        .ZN(pe_1_6_4_n33) );
  INV_X1 pe_1_6_4_U60 ( .A(pe_1_6_4_n33), .ZN(pe_1_6_4_n82) );
  AOI222_X1 pe_1_6_4_U59 ( .A1(int_data_res_7__4__6_), .A2(pe_1_6_4_n64), .B1(
        pe_1_6_4_N84), .B2(pe_1_6_4_n27), .C1(pe_1_6_4_N76), .C2(pe_1_6_4_n28), 
        .ZN(pe_1_6_4_n29) );
  INV_X1 pe_1_6_4_U58 ( .A(pe_1_6_4_n29), .ZN(pe_1_6_4_n78) );
  XNOR2_X1 pe_1_6_4_U57 ( .A(pe_1_6_4_n73), .B(int_data_res_6__4__0_), .ZN(
        pe_1_6_4_N70) );
  AOI222_X1 pe_1_6_4_U52 ( .A1(int_data_res_7__4__0_), .A2(pe_1_6_4_n64), .B1(
        pe_1_6_4_n1), .B2(pe_1_6_4_n27), .C1(pe_1_6_4_N70), .C2(pe_1_6_4_n28), 
        .ZN(pe_1_6_4_n35) );
  INV_X1 pe_1_6_4_U51 ( .A(pe_1_6_4_n35), .ZN(pe_1_6_4_n84) );
  AOI222_X1 pe_1_6_4_U50 ( .A1(int_data_res_7__4__1_), .A2(pe_1_6_4_n64), .B1(
        pe_1_6_4_N79), .B2(pe_1_6_4_n27), .C1(pe_1_6_4_N71), .C2(pe_1_6_4_n28), 
        .ZN(pe_1_6_4_n34) );
  INV_X1 pe_1_6_4_U49 ( .A(pe_1_6_4_n34), .ZN(pe_1_6_4_n83) );
  AOI222_X1 pe_1_6_4_U48 ( .A1(int_data_res_7__4__3_), .A2(pe_1_6_4_n64), .B1(
        pe_1_6_4_N81), .B2(pe_1_6_4_n27), .C1(pe_1_6_4_N73), .C2(pe_1_6_4_n28), 
        .ZN(pe_1_6_4_n32) );
  INV_X1 pe_1_6_4_U47 ( .A(pe_1_6_4_n32), .ZN(pe_1_6_4_n81) );
  AOI222_X1 pe_1_6_4_U46 ( .A1(int_data_res_7__4__4_), .A2(pe_1_6_4_n64), .B1(
        pe_1_6_4_N82), .B2(pe_1_6_4_n27), .C1(pe_1_6_4_N74), .C2(pe_1_6_4_n28), 
        .ZN(pe_1_6_4_n31) );
  INV_X1 pe_1_6_4_U45 ( .A(pe_1_6_4_n31), .ZN(pe_1_6_4_n80) );
  AOI222_X1 pe_1_6_4_U44 ( .A1(int_data_res_7__4__5_), .A2(pe_1_6_4_n64), .B1(
        pe_1_6_4_N83), .B2(pe_1_6_4_n27), .C1(pe_1_6_4_N75), .C2(pe_1_6_4_n28), 
        .ZN(pe_1_6_4_n30) );
  INV_X1 pe_1_6_4_U43 ( .A(pe_1_6_4_n30), .ZN(pe_1_6_4_n79) );
  NAND2_X1 pe_1_6_4_U42 ( .A1(pe_1_6_4_int_data_0_), .A2(pe_1_6_4_n3), .ZN(
        pe_1_6_4_sub_81_carry[1]) );
  INV_X1 pe_1_6_4_U41 ( .A(pe_1_6_4_int_data_1_), .ZN(pe_1_6_4_n74) );
  INV_X1 pe_1_6_4_U40 ( .A(pe_1_6_4_int_data_2_), .ZN(pe_1_6_4_n75) );
  AND2_X1 pe_1_6_4_U39 ( .A1(pe_1_6_4_int_data_0_), .A2(int_data_res_6__4__0_), 
        .ZN(pe_1_6_4_n2) );
  AOI222_X1 pe_1_6_4_U38 ( .A1(pe_1_6_4_n64), .A2(int_data_res_7__4__7_), .B1(
        pe_1_6_4_N85), .B2(pe_1_6_4_n27), .C1(pe_1_6_4_N77), .C2(pe_1_6_4_n28), 
        .ZN(pe_1_6_4_n26) );
  INV_X1 pe_1_6_4_U37 ( .A(pe_1_6_4_n26), .ZN(pe_1_6_4_n77) );
  NOR3_X1 pe_1_6_4_U36 ( .A1(pe_1_6_4_n59), .A2(pe_1_6_4_n65), .A3(int_ckg[11]), .ZN(pe_1_6_4_n36) );
  OR2_X1 pe_1_6_4_U35 ( .A1(pe_1_6_4_n36), .A2(pe_1_6_4_n64), .ZN(pe_1_6_4_N90) );
  INV_X1 pe_1_6_4_U34 ( .A(n41), .ZN(pe_1_6_4_n63) );
  AND2_X1 pe_1_6_4_U33 ( .A1(int_data_x_6__4__2_), .A2(pe_1_6_4_n58), .ZN(
        pe_1_6_4_int_data_2_) );
  AND2_X1 pe_1_6_4_U32 ( .A1(int_data_x_6__4__1_), .A2(pe_1_6_4_n58), .ZN(
        pe_1_6_4_int_data_1_) );
  AND2_X1 pe_1_6_4_U31 ( .A1(int_data_x_6__4__3_), .A2(pe_1_6_4_n58), .ZN(
        pe_1_6_4_int_data_3_) );
  BUF_X1 pe_1_6_4_U30 ( .A(n63), .Z(pe_1_6_4_n64) );
  INV_X1 pe_1_6_4_U29 ( .A(n35), .ZN(pe_1_6_4_n61) );
  AND2_X1 pe_1_6_4_U28 ( .A1(int_data_x_6__4__0_), .A2(pe_1_6_4_n58), .ZN(
        pe_1_6_4_int_data_0_) );
  NAND2_X1 pe_1_6_4_U27 ( .A1(pe_1_6_4_n44), .A2(pe_1_6_4_n61), .ZN(
        pe_1_6_4_n41) );
  AND3_X1 pe_1_6_4_U26 ( .A1(n77), .A2(pe_1_6_4_n63), .A3(n53), .ZN(
        pe_1_6_4_n44) );
  INV_X1 pe_1_6_4_U25 ( .A(pe_1_6_4_int_data_3_), .ZN(pe_1_6_4_n76) );
  NOR2_X1 pe_1_6_4_U24 ( .A1(pe_1_6_4_n70), .A2(n53), .ZN(pe_1_6_4_n43) );
  NOR2_X1 pe_1_6_4_U23 ( .A1(pe_1_6_4_n57), .A2(pe_1_6_4_n64), .ZN(
        pe_1_6_4_n28) );
  NOR2_X1 pe_1_6_4_U22 ( .A1(n21), .A2(pe_1_6_4_n64), .ZN(pe_1_6_4_n27) );
  INV_X1 pe_1_6_4_U21 ( .A(pe_1_6_4_int_data_0_), .ZN(pe_1_6_4_n73) );
  INV_X1 pe_1_6_4_U20 ( .A(pe_1_6_4_n41), .ZN(pe_1_6_4_n90) );
  INV_X1 pe_1_6_4_U19 ( .A(pe_1_6_4_n37), .ZN(pe_1_6_4_n88) );
  INV_X1 pe_1_6_4_U18 ( .A(pe_1_6_4_n38), .ZN(pe_1_6_4_n87) );
  INV_X1 pe_1_6_4_U17 ( .A(pe_1_6_4_n39), .ZN(pe_1_6_4_n86) );
  NOR2_X1 pe_1_6_4_U16 ( .A1(pe_1_6_4_n68), .A2(pe_1_6_4_n42), .ZN(
        pe_1_6_4_N59) );
  NOR2_X1 pe_1_6_4_U15 ( .A1(pe_1_6_4_n68), .A2(pe_1_6_4_n41), .ZN(
        pe_1_6_4_N60) );
  NOR2_X1 pe_1_6_4_U14 ( .A1(pe_1_6_4_n68), .A2(pe_1_6_4_n38), .ZN(
        pe_1_6_4_N63) );
  NOR2_X1 pe_1_6_4_U13 ( .A1(pe_1_6_4_n67), .A2(pe_1_6_4_n40), .ZN(
        pe_1_6_4_N61) );
  NOR2_X1 pe_1_6_4_U12 ( .A1(pe_1_6_4_n67), .A2(pe_1_6_4_n39), .ZN(
        pe_1_6_4_N62) );
  NOR2_X1 pe_1_6_4_U11 ( .A1(pe_1_6_4_n37), .A2(pe_1_6_4_n67), .ZN(
        pe_1_6_4_N64) );
  NAND2_X1 pe_1_6_4_U10 ( .A1(pe_1_6_4_n44), .A2(pe_1_6_4_n60), .ZN(
        pe_1_6_4_n42) );
  BUF_X1 pe_1_6_4_U9 ( .A(pe_1_6_4_n60), .Z(pe_1_6_4_n55) );
  INV_X1 pe_1_6_4_U8 ( .A(pe_1_6_4_n69), .ZN(pe_1_6_4_n65) );
  BUF_X1 pe_1_6_4_U7 ( .A(pe_1_6_4_n60), .Z(pe_1_6_4_n56) );
  INV_X1 pe_1_6_4_U6 ( .A(pe_1_6_4_n42), .ZN(pe_1_6_4_n89) );
  INV_X1 pe_1_6_4_U5 ( .A(pe_1_6_4_n40), .ZN(pe_1_6_4_n85) );
  INV_X2 pe_1_6_4_U4 ( .A(n85), .ZN(pe_1_6_4_n72) );
  XOR2_X1 pe_1_6_4_U3 ( .A(pe_1_6_4_int_data_0_), .B(int_data_res_6__4__0_), 
        .Z(pe_1_6_4_n1) );
  DFFR_X1 pe_1_6_4_int_q_acc_reg_0_ ( .D(pe_1_6_4_n84), .CK(pe_1_6_4_net3496), 
        .RN(pe_1_6_4_n72), .Q(int_data_res_6__4__0_), .QN(pe_1_6_4_n3) );
  DFFR_X1 pe_1_6_4_int_q_reg_v_reg_0__0_ ( .D(int_data_y_7__4__0_), .CK(
        pe_1_6_4_net3466), .RN(pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_v[20]) );
  DFFR_X1 pe_1_6_4_int_q_reg_v_reg_0__1_ ( .D(int_data_y_7__4__1_), .CK(
        pe_1_6_4_net3466), .RN(pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_v[21]) );
  DFFR_X1 pe_1_6_4_int_q_reg_v_reg_0__2_ ( .D(int_data_y_7__4__2_), .CK(
        pe_1_6_4_net3466), .RN(pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_v[22]) );
  DFFR_X1 pe_1_6_4_int_q_reg_v_reg_0__3_ ( .D(int_data_y_7__4__3_), .CK(
        pe_1_6_4_net3466), .RN(pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_v[23]) );
  DFFR_X1 pe_1_6_4_int_q_reg_v_reg_1__0_ ( .D(int_data_y_7__4__0_), .CK(
        pe_1_6_4_net3471), .RN(pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_v[16]) );
  DFFR_X1 pe_1_6_4_int_q_reg_v_reg_1__1_ ( .D(int_data_y_7__4__1_), .CK(
        pe_1_6_4_net3471), .RN(pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_v[17]) );
  DFFR_X1 pe_1_6_4_int_q_reg_v_reg_1__2_ ( .D(int_data_y_7__4__2_), .CK(
        pe_1_6_4_net3471), .RN(pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_v[18]) );
  DFFR_X1 pe_1_6_4_int_q_reg_v_reg_1__3_ ( .D(int_data_y_7__4__3_), .CK(
        pe_1_6_4_net3471), .RN(pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_v[19]) );
  DFFR_X1 pe_1_6_4_int_q_reg_v_reg_2__0_ ( .D(int_data_y_7__4__0_), .CK(
        pe_1_6_4_net3476), .RN(pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_v[12]) );
  DFFR_X1 pe_1_6_4_int_q_reg_v_reg_2__1_ ( .D(int_data_y_7__4__1_), .CK(
        pe_1_6_4_net3476), .RN(pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_v[13]) );
  DFFR_X1 pe_1_6_4_int_q_reg_v_reg_2__2_ ( .D(int_data_y_7__4__2_), .CK(
        pe_1_6_4_net3476), .RN(pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_v[14]) );
  DFFR_X1 pe_1_6_4_int_q_reg_v_reg_2__3_ ( .D(int_data_y_7__4__3_), .CK(
        pe_1_6_4_net3476), .RN(pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_v[15]) );
  DFFR_X1 pe_1_6_4_int_q_reg_v_reg_3__0_ ( .D(int_data_y_7__4__0_), .CK(
        pe_1_6_4_net3481), .RN(pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_v[8]) );
  DFFR_X1 pe_1_6_4_int_q_reg_v_reg_3__1_ ( .D(int_data_y_7__4__1_), .CK(
        pe_1_6_4_net3481), .RN(pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_v[9]) );
  DFFR_X1 pe_1_6_4_int_q_reg_v_reg_3__2_ ( .D(int_data_y_7__4__2_), .CK(
        pe_1_6_4_net3481), .RN(pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_v[10]) );
  DFFR_X1 pe_1_6_4_int_q_reg_v_reg_3__3_ ( .D(int_data_y_7__4__3_), .CK(
        pe_1_6_4_net3481), .RN(pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_v[11]) );
  DFFR_X1 pe_1_6_4_int_q_reg_v_reg_4__0_ ( .D(int_data_y_7__4__0_), .CK(
        pe_1_6_4_net3486), .RN(pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_v[4]) );
  DFFR_X1 pe_1_6_4_int_q_reg_v_reg_4__1_ ( .D(int_data_y_7__4__1_), .CK(
        pe_1_6_4_net3486), .RN(pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_v[5]) );
  DFFR_X1 pe_1_6_4_int_q_reg_v_reg_4__2_ ( .D(int_data_y_7__4__2_), .CK(
        pe_1_6_4_net3486), .RN(pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_v[6]) );
  DFFR_X1 pe_1_6_4_int_q_reg_v_reg_4__3_ ( .D(int_data_y_7__4__3_), .CK(
        pe_1_6_4_net3486), .RN(pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_v[7]) );
  DFFR_X1 pe_1_6_4_int_q_reg_v_reg_5__0_ ( .D(int_data_y_7__4__0_), .CK(
        pe_1_6_4_net3491), .RN(pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_v[0]) );
  DFFR_X1 pe_1_6_4_int_q_reg_v_reg_5__1_ ( .D(int_data_y_7__4__1_), .CK(
        pe_1_6_4_net3491), .RN(pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_v[1]) );
  DFFR_X1 pe_1_6_4_int_q_reg_v_reg_5__2_ ( .D(int_data_y_7__4__2_), .CK(
        pe_1_6_4_net3491), .RN(pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_v[2]) );
  DFFR_X1 pe_1_6_4_int_q_reg_v_reg_5__3_ ( .D(int_data_y_7__4__3_), .CK(
        pe_1_6_4_net3491), .RN(pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_6_4_int_q_reg_h_reg_0__0_ ( .D(int_data_x_6__5__0_), .SI(
        int_data_y_7__4__0_), .SE(pe_1_6_4_n65), .CK(pe_1_6_4_net3435), .RN(
        pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_6_4_int_q_reg_h_reg_0__1_ ( .D(int_data_x_6__5__1_), .SI(
        int_data_y_7__4__1_), .SE(pe_1_6_4_n65), .CK(pe_1_6_4_net3435), .RN(
        pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_6_4_int_q_reg_h_reg_0__2_ ( .D(int_data_x_6__5__2_), .SI(
        int_data_y_7__4__2_), .SE(pe_1_6_4_n65), .CK(pe_1_6_4_net3435), .RN(
        pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_6_4_int_q_reg_h_reg_0__3_ ( .D(int_data_x_6__5__3_), .SI(
        int_data_y_7__4__3_), .SE(pe_1_6_4_n65), .CK(pe_1_6_4_net3435), .RN(
        pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_6_4_int_q_reg_h_reg_1__0_ ( .D(int_data_x_6__5__0_), .SI(
        int_data_y_7__4__0_), .SE(pe_1_6_4_n65), .CK(pe_1_6_4_net3441), .RN(
        pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_6_4_int_q_reg_h_reg_1__1_ ( .D(int_data_x_6__5__1_), .SI(
        int_data_y_7__4__1_), .SE(pe_1_6_4_n65), .CK(pe_1_6_4_net3441), .RN(
        pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_6_4_int_q_reg_h_reg_1__2_ ( .D(int_data_x_6__5__2_), .SI(
        int_data_y_7__4__2_), .SE(pe_1_6_4_n65), .CK(pe_1_6_4_net3441), .RN(
        pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_6_4_int_q_reg_h_reg_1__3_ ( .D(int_data_x_6__5__3_), .SI(
        int_data_y_7__4__3_), .SE(pe_1_6_4_n65), .CK(pe_1_6_4_net3441), .RN(
        pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_6_4_int_q_reg_h_reg_2__0_ ( .D(int_data_x_6__5__0_), .SI(
        int_data_y_7__4__0_), .SE(pe_1_6_4_n65), .CK(pe_1_6_4_net3446), .RN(
        pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_6_4_int_q_reg_h_reg_2__1_ ( .D(int_data_x_6__5__1_), .SI(
        int_data_y_7__4__1_), .SE(pe_1_6_4_n65), .CK(pe_1_6_4_net3446), .RN(
        pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_6_4_int_q_reg_h_reg_2__2_ ( .D(int_data_x_6__5__2_), .SI(
        int_data_y_7__4__2_), .SE(pe_1_6_4_n65), .CK(pe_1_6_4_net3446), .RN(
        pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_6_4_int_q_reg_h_reg_2__3_ ( .D(int_data_x_6__5__3_), .SI(
        int_data_y_7__4__3_), .SE(pe_1_6_4_n65), .CK(pe_1_6_4_net3446), .RN(
        pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_6_4_int_q_reg_h_reg_3__0_ ( .D(int_data_x_6__5__0_), .SI(
        int_data_y_7__4__0_), .SE(pe_1_6_4_n65), .CK(pe_1_6_4_net3451), .RN(
        pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_6_4_int_q_reg_h_reg_3__1_ ( .D(int_data_x_6__5__1_), .SI(
        int_data_y_7__4__1_), .SE(pe_1_6_4_n65), .CK(pe_1_6_4_net3451), .RN(
        pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_6_4_int_q_reg_h_reg_3__2_ ( .D(int_data_x_6__5__2_), .SI(
        int_data_y_7__4__2_), .SE(pe_1_6_4_n65), .CK(pe_1_6_4_net3451), .RN(
        pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_6_4_int_q_reg_h_reg_3__3_ ( .D(int_data_x_6__5__3_), .SI(
        int_data_y_7__4__3_), .SE(pe_1_6_4_n65), .CK(pe_1_6_4_net3451), .RN(
        pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_6_4_int_q_reg_h_reg_4__0_ ( .D(int_data_x_6__5__0_), .SI(
        int_data_y_7__4__0_), .SE(pe_1_6_4_n66), .CK(pe_1_6_4_net3456), .RN(
        pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_6_4_int_q_reg_h_reg_4__1_ ( .D(int_data_x_6__5__1_), .SI(
        int_data_y_7__4__1_), .SE(pe_1_6_4_n66), .CK(pe_1_6_4_net3456), .RN(
        pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_6_4_int_q_reg_h_reg_4__2_ ( .D(int_data_x_6__5__2_), .SI(
        int_data_y_7__4__2_), .SE(pe_1_6_4_n66), .CK(pe_1_6_4_net3456), .RN(
        pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_6_4_int_q_reg_h_reg_4__3_ ( .D(int_data_x_6__5__3_), .SI(
        int_data_y_7__4__3_), .SE(pe_1_6_4_n66), .CK(pe_1_6_4_net3456), .RN(
        pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_6_4_int_q_reg_h_reg_5__0_ ( .D(int_data_x_6__5__0_), .SI(
        int_data_y_7__4__0_), .SE(pe_1_6_4_n66), .CK(pe_1_6_4_net3461), .RN(
        pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_6_4_int_q_reg_h_reg_5__1_ ( .D(int_data_x_6__5__1_), .SI(
        int_data_y_7__4__1_), .SE(pe_1_6_4_n66), .CK(pe_1_6_4_net3461), .RN(
        pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_6_4_int_q_reg_h_reg_5__2_ ( .D(int_data_x_6__5__2_), .SI(
        int_data_y_7__4__2_), .SE(pe_1_6_4_n66), .CK(pe_1_6_4_net3461), .RN(
        pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_6_4_int_q_reg_h_reg_5__3_ ( .D(int_data_x_6__5__3_), .SI(
        int_data_y_7__4__3_), .SE(pe_1_6_4_n66), .CK(pe_1_6_4_net3461), .RN(
        pe_1_6_4_n72), .Q(pe_1_6_4_int_q_reg_h[3]) );
  FA_X1 pe_1_6_4_sub_81_U2_7 ( .A(int_data_res_6__4__7_), .B(pe_1_6_4_n76), 
        .CI(pe_1_6_4_sub_81_carry[7]), .S(pe_1_6_4_N77) );
  FA_X1 pe_1_6_4_sub_81_U2_6 ( .A(int_data_res_6__4__6_), .B(pe_1_6_4_n76), 
        .CI(pe_1_6_4_sub_81_carry[6]), .CO(pe_1_6_4_sub_81_carry[7]), .S(
        pe_1_6_4_N76) );
  FA_X1 pe_1_6_4_sub_81_U2_5 ( .A(int_data_res_6__4__5_), .B(pe_1_6_4_n76), 
        .CI(pe_1_6_4_sub_81_carry[5]), .CO(pe_1_6_4_sub_81_carry[6]), .S(
        pe_1_6_4_N75) );
  FA_X1 pe_1_6_4_sub_81_U2_4 ( .A(int_data_res_6__4__4_), .B(pe_1_6_4_n76), 
        .CI(pe_1_6_4_sub_81_carry[4]), .CO(pe_1_6_4_sub_81_carry[5]), .S(
        pe_1_6_4_N74) );
  FA_X1 pe_1_6_4_sub_81_U2_3 ( .A(int_data_res_6__4__3_), .B(pe_1_6_4_n76), 
        .CI(pe_1_6_4_sub_81_carry[3]), .CO(pe_1_6_4_sub_81_carry[4]), .S(
        pe_1_6_4_N73) );
  FA_X1 pe_1_6_4_sub_81_U2_2 ( .A(int_data_res_6__4__2_), .B(pe_1_6_4_n75), 
        .CI(pe_1_6_4_sub_81_carry[2]), .CO(pe_1_6_4_sub_81_carry[3]), .S(
        pe_1_6_4_N72) );
  FA_X1 pe_1_6_4_sub_81_U2_1 ( .A(int_data_res_6__4__1_), .B(pe_1_6_4_n74), 
        .CI(pe_1_6_4_sub_81_carry[1]), .CO(pe_1_6_4_sub_81_carry[2]), .S(
        pe_1_6_4_N71) );
  FA_X1 pe_1_6_4_add_83_U1_7 ( .A(int_data_res_6__4__7_), .B(
        pe_1_6_4_int_data_3_), .CI(pe_1_6_4_add_83_carry[7]), .S(pe_1_6_4_N85)
         );
  FA_X1 pe_1_6_4_add_83_U1_6 ( .A(int_data_res_6__4__6_), .B(
        pe_1_6_4_int_data_3_), .CI(pe_1_6_4_add_83_carry[6]), .CO(
        pe_1_6_4_add_83_carry[7]), .S(pe_1_6_4_N84) );
  FA_X1 pe_1_6_4_add_83_U1_5 ( .A(int_data_res_6__4__5_), .B(
        pe_1_6_4_int_data_3_), .CI(pe_1_6_4_add_83_carry[5]), .CO(
        pe_1_6_4_add_83_carry[6]), .S(pe_1_6_4_N83) );
  FA_X1 pe_1_6_4_add_83_U1_4 ( .A(int_data_res_6__4__4_), .B(
        pe_1_6_4_int_data_3_), .CI(pe_1_6_4_add_83_carry[4]), .CO(
        pe_1_6_4_add_83_carry[5]), .S(pe_1_6_4_N82) );
  FA_X1 pe_1_6_4_add_83_U1_3 ( .A(int_data_res_6__4__3_), .B(
        pe_1_6_4_int_data_3_), .CI(pe_1_6_4_add_83_carry[3]), .CO(
        pe_1_6_4_add_83_carry[4]), .S(pe_1_6_4_N81) );
  FA_X1 pe_1_6_4_add_83_U1_2 ( .A(int_data_res_6__4__2_), .B(
        pe_1_6_4_int_data_2_), .CI(pe_1_6_4_add_83_carry[2]), .CO(
        pe_1_6_4_add_83_carry[3]), .S(pe_1_6_4_N80) );
  FA_X1 pe_1_6_4_add_83_U1_1 ( .A(int_data_res_6__4__1_), .B(
        pe_1_6_4_int_data_1_), .CI(pe_1_6_4_n2), .CO(pe_1_6_4_add_83_carry[2]), 
        .S(pe_1_6_4_N79) );
  NAND3_X1 pe_1_6_4_U56 ( .A1(pe_1_6_4_n60), .A2(pe_1_6_4_n43), .A3(
        pe_1_6_4_n62), .ZN(pe_1_6_4_n40) );
  NAND3_X1 pe_1_6_4_U55 ( .A1(pe_1_6_4_n43), .A2(pe_1_6_4_n61), .A3(
        pe_1_6_4_n62), .ZN(pe_1_6_4_n39) );
  NAND3_X1 pe_1_6_4_U54 ( .A1(pe_1_6_4_n43), .A2(pe_1_6_4_n63), .A3(
        pe_1_6_4_n60), .ZN(pe_1_6_4_n38) );
  NAND3_X1 pe_1_6_4_U53 ( .A1(pe_1_6_4_n61), .A2(pe_1_6_4_n63), .A3(
        pe_1_6_4_n43), .ZN(pe_1_6_4_n37) );
  DFFR_X1 pe_1_6_4_int_q_acc_reg_6_ ( .D(pe_1_6_4_n78), .CK(pe_1_6_4_net3496), 
        .RN(pe_1_6_4_n71), .Q(int_data_res_6__4__6_) );
  DFFR_X1 pe_1_6_4_int_q_acc_reg_5_ ( .D(pe_1_6_4_n79), .CK(pe_1_6_4_net3496), 
        .RN(pe_1_6_4_n71), .Q(int_data_res_6__4__5_) );
  DFFR_X1 pe_1_6_4_int_q_acc_reg_4_ ( .D(pe_1_6_4_n80), .CK(pe_1_6_4_net3496), 
        .RN(pe_1_6_4_n71), .Q(int_data_res_6__4__4_) );
  DFFR_X1 pe_1_6_4_int_q_acc_reg_3_ ( .D(pe_1_6_4_n81), .CK(pe_1_6_4_net3496), 
        .RN(pe_1_6_4_n71), .Q(int_data_res_6__4__3_) );
  DFFR_X1 pe_1_6_4_int_q_acc_reg_2_ ( .D(pe_1_6_4_n82), .CK(pe_1_6_4_net3496), 
        .RN(pe_1_6_4_n71), .Q(int_data_res_6__4__2_) );
  DFFR_X1 pe_1_6_4_int_q_acc_reg_1_ ( .D(pe_1_6_4_n83), .CK(pe_1_6_4_net3496), 
        .RN(pe_1_6_4_n71), .Q(int_data_res_6__4__1_) );
  DFFR_X1 pe_1_6_4_int_q_acc_reg_7_ ( .D(pe_1_6_4_n77), .CK(pe_1_6_4_net3496), 
        .RN(pe_1_6_4_n71), .Q(int_data_res_6__4__7_) );
  CLKGATETST_X1 pe_1_6_4_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_6_4_n88), .SE(1'b0), .GCK(pe_1_6_4_net3435) );
  CLKGATETST_X1 pe_1_6_4_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_6_4_n87), .SE(1'b0), .GCK(pe_1_6_4_net3441) );
  CLKGATETST_X1 pe_1_6_4_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_6_4_n86), .SE(1'b0), .GCK(pe_1_6_4_net3446) );
  CLKGATETST_X1 pe_1_6_4_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_6_4_n85), .SE(1'b0), .GCK(pe_1_6_4_net3451) );
  CLKGATETST_X1 pe_1_6_4_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_6_4_n90), .SE(1'b0), .GCK(pe_1_6_4_net3456) );
  CLKGATETST_X1 pe_1_6_4_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_6_4_n89), .SE(1'b0), .GCK(pe_1_6_4_net3461) );
  CLKGATETST_X1 pe_1_6_4_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_6_4_N64), .SE(1'b0), .GCK(pe_1_6_4_net3466) );
  CLKGATETST_X1 pe_1_6_4_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_6_4_N63), .SE(1'b0), .GCK(pe_1_6_4_net3471) );
  CLKGATETST_X1 pe_1_6_4_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_6_4_N62), .SE(1'b0), .GCK(pe_1_6_4_net3476) );
  CLKGATETST_X1 pe_1_6_4_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_6_4_N61), .SE(1'b0), .GCK(pe_1_6_4_net3481) );
  CLKGATETST_X1 pe_1_6_4_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_6_4_N60), .SE(1'b0), .GCK(pe_1_6_4_net3486) );
  CLKGATETST_X1 pe_1_6_4_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_6_4_N59), .SE(1'b0), .GCK(pe_1_6_4_net3491) );
  CLKGATETST_X1 pe_1_6_4_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_6_4_N90), .SE(1'b0), .GCK(pe_1_6_4_net3496) );
  CLKBUF_X1 pe_1_6_5_U112 ( .A(pe_1_6_5_n72), .Z(pe_1_6_5_n71) );
  INV_X1 pe_1_6_5_U111 ( .A(n77), .ZN(pe_1_6_5_n70) );
  INV_X1 pe_1_6_5_U110 ( .A(n69), .ZN(pe_1_6_5_n69) );
  INV_X1 pe_1_6_5_U109 ( .A(n69), .ZN(pe_1_6_5_n68) );
  INV_X1 pe_1_6_5_U108 ( .A(n69), .ZN(pe_1_6_5_n67) );
  INV_X1 pe_1_6_5_U107 ( .A(pe_1_6_5_n69), .ZN(pe_1_6_5_n66) );
  INV_X1 pe_1_6_5_U106 ( .A(pe_1_6_5_n63), .ZN(pe_1_6_5_n62) );
  INV_X1 pe_1_6_5_U105 ( .A(pe_1_6_5_n61), .ZN(pe_1_6_5_n60) );
  INV_X1 pe_1_6_5_U104 ( .A(n29), .ZN(pe_1_6_5_n59) );
  INV_X1 pe_1_6_5_U103 ( .A(pe_1_6_5_n59), .ZN(pe_1_6_5_n58) );
  INV_X1 pe_1_6_5_U102 ( .A(n21), .ZN(pe_1_6_5_n57) );
  MUX2_X1 pe_1_6_5_U101 ( .A(pe_1_6_5_n54), .B(pe_1_6_5_n51), .S(n53), .Z(
        int_data_x_6__5__3_) );
  MUX2_X1 pe_1_6_5_U100 ( .A(pe_1_6_5_n53), .B(pe_1_6_5_n52), .S(pe_1_6_5_n62), 
        .Z(pe_1_6_5_n54) );
  MUX2_X1 pe_1_6_5_U99 ( .A(pe_1_6_5_int_q_reg_h[23]), .B(
        pe_1_6_5_int_q_reg_h[19]), .S(pe_1_6_5_n56), .Z(pe_1_6_5_n53) );
  MUX2_X1 pe_1_6_5_U98 ( .A(pe_1_6_5_int_q_reg_h[15]), .B(
        pe_1_6_5_int_q_reg_h[11]), .S(pe_1_6_5_n56), .Z(pe_1_6_5_n52) );
  MUX2_X1 pe_1_6_5_U97 ( .A(pe_1_6_5_int_q_reg_h[7]), .B(
        pe_1_6_5_int_q_reg_h[3]), .S(pe_1_6_5_n56), .Z(pe_1_6_5_n51) );
  MUX2_X1 pe_1_6_5_U96 ( .A(pe_1_6_5_n50), .B(pe_1_6_5_n47), .S(n53), .Z(
        int_data_x_6__5__2_) );
  MUX2_X1 pe_1_6_5_U95 ( .A(pe_1_6_5_n49), .B(pe_1_6_5_n48), .S(pe_1_6_5_n62), 
        .Z(pe_1_6_5_n50) );
  MUX2_X1 pe_1_6_5_U94 ( .A(pe_1_6_5_int_q_reg_h[22]), .B(
        pe_1_6_5_int_q_reg_h[18]), .S(pe_1_6_5_n56), .Z(pe_1_6_5_n49) );
  MUX2_X1 pe_1_6_5_U93 ( .A(pe_1_6_5_int_q_reg_h[14]), .B(
        pe_1_6_5_int_q_reg_h[10]), .S(pe_1_6_5_n56), .Z(pe_1_6_5_n48) );
  MUX2_X1 pe_1_6_5_U92 ( .A(pe_1_6_5_int_q_reg_h[6]), .B(
        pe_1_6_5_int_q_reg_h[2]), .S(pe_1_6_5_n56), .Z(pe_1_6_5_n47) );
  MUX2_X1 pe_1_6_5_U91 ( .A(pe_1_6_5_n46), .B(pe_1_6_5_n24), .S(n53), .Z(
        int_data_x_6__5__1_) );
  MUX2_X1 pe_1_6_5_U90 ( .A(pe_1_6_5_n45), .B(pe_1_6_5_n25), .S(pe_1_6_5_n62), 
        .Z(pe_1_6_5_n46) );
  MUX2_X1 pe_1_6_5_U89 ( .A(pe_1_6_5_int_q_reg_h[21]), .B(
        pe_1_6_5_int_q_reg_h[17]), .S(pe_1_6_5_n56), .Z(pe_1_6_5_n45) );
  MUX2_X1 pe_1_6_5_U88 ( .A(pe_1_6_5_int_q_reg_h[13]), .B(
        pe_1_6_5_int_q_reg_h[9]), .S(pe_1_6_5_n56), .Z(pe_1_6_5_n25) );
  MUX2_X1 pe_1_6_5_U87 ( .A(pe_1_6_5_int_q_reg_h[5]), .B(
        pe_1_6_5_int_q_reg_h[1]), .S(pe_1_6_5_n56), .Z(pe_1_6_5_n24) );
  MUX2_X1 pe_1_6_5_U86 ( .A(pe_1_6_5_n23), .B(pe_1_6_5_n20), .S(n53), .Z(
        int_data_x_6__5__0_) );
  MUX2_X1 pe_1_6_5_U85 ( .A(pe_1_6_5_n22), .B(pe_1_6_5_n21), .S(pe_1_6_5_n62), 
        .Z(pe_1_6_5_n23) );
  MUX2_X1 pe_1_6_5_U84 ( .A(pe_1_6_5_int_q_reg_h[20]), .B(
        pe_1_6_5_int_q_reg_h[16]), .S(pe_1_6_5_n56), .Z(pe_1_6_5_n22) );
  MUX2_X1 pe_1_6_5_U83 ( .A(pe_1_6_5_int_q_reg_h[12]), .B(
        pe_1_6_5_int_q_reg_h[8]), .S(pe_1_6_5_n56), .Z(pe_1_6_5_n21) );
  MUX2_X1 pe_1_6_5_U82 ( .A(pe_1_6_5_int_q_reg_h[4]), .B(
        pe_1_6_5_int_q_reg_h[0]), .S(pe_1_6_5_n56), .Z(pe_1_6_5_n20) );
  MUX2_X1 pe_1_6_5_U81 ( .A(pe_1_6_5_n19), .B(pe_1_6_5_n16), .S(n53), .Z(
        int_data_y_6__5__3_) );
  MUX2_X1 pe_1_6_5_U80 ( .A(pe_1_6_5_n18), .B(pe_1_6_5_n17), .S(pe_1_6_5_n62), 
        .Z(pe_1_6_5_n19) );
  MUX2_X1 pe_1_6_5_U79 ( .A(pe_1_6_5_int_q_reg_v[23]), .B(
        pe_1_6_5_int_q_reg_v[19]), .S(pe_1_6_5_n55), .Z(pe_1_6_5_n18) );
  MUX2_X1 pe_1_6_5_U78 ( .A(pe_1_6_5_int_q_reg_v[15]), .B(
        pe_1_6_5_int_q_reg_v[11]), .S(pe_1_6_5_n55), .Z(pe_1_6_5_n17) );
  MUX2_X1 pe_1_6_5_U77 ( .A(pe_1_6_5_int_q_reg_v[7]), .B(
        pe_1_6_5_int_q_reg_v[3]), .S(pe_1_6_5_n55), .Z(pe_1_6_5_n16) );
  MUX2_X1 pe_1_6_5_U76 ( .A(pe_1_6_5_n15), .B(pe_1_6_5_n12), .S(n53), .Z(
        int_data_y_6__5__2_) );
  MUX2_X1 pe_1_6_5_U75 ( .A(pe_1_6_5_n14), .B(pe_1_6_5_n13), .S(pe_1_6_5_n62), 
        .Z(pe_1_6_5_n15) );
  MUX2_X1 pe_1_6_5_U74 ( .A(pe_1_6_5_int_q_reg_v[22]), .B(
        pe_1_6_5_int_q_reg_v[18]), .S(pe_1_6_5_n55), .Z(pe_1_6_5_n14) );
  MUX2_X1 pe_1_6_5_U73 ( .A(pe_1_6_5_int_q_reg_v[14]), .B(
        pe_1_6_5_int_q_reg_v[10]), .S(pe_1_6_5_n55), .Z(pe_1_6_5_n13) );
  MUX2_X1 pe_1_6_5_U72 ( .A(pe_1_6_5_int_q_reg_v[6]), .B(
        pe_1_6_5_int_q_reg_v[2]), .S(pe_1_6_5_n55), .Z(pe_1_6_5_n12) );
  MUX2_X1 pe_1_6_5_U71 ( .A(pe_1_6_5_n11), .B(pe_1_6_5_n8), .S(n53), .Z(
        int_data_y_6__5__1_) );
  MUX2_X1 pe_1_6_5_U70 ( .A(pe_1_6_5_n10), .B(pe_1_6_5_n9), .S(pe_1_6_5_n62), 
        .Z(pe_1_6_5_n11) );
  MUX2_X1 pe_1_6_5_U69 ( .A(pe_1_6_5_int_q_reg_v[21]), .B(
        pe_1_6_5_int_q_reg_v[17]), .S(pe_1_6_5_n55), .Z(pe_1_6_5_n10) );
  MUX2_X1 pe_1_6_5_U68 ( .A(pe_1_6_5_int_q_reg_v[13]), .B(
        pe_1_6_5_int_q_reg_v[9]), .S(pe_1_6_5_n55), .Z(pe_1_6_5_n9) );
  MUX2_X1 pe_1_6_5_U67 ( .A(pe_1_6_5_int_q_reg_v[5]), .B(
        pe_1_6_5_int_q_reg_v[1]), .S(pe_1_6_5_n55), .Z(pe_1_6_5_n8) );
  MUX2_X1 pe_1_6_5_U66 ( .A(pe_1_6_5_n7), .B(pe_1_6_5_n4), .S(n53), .Z(
        int_data_y_6__5__0_) );
  MUX2_X1 pe_1_6_5_U65 ( .A(pe_1_6_5_n6), .B(pe_1_6_5_n5), .S(pe_1_6_5_n62), 
        .Z(pe_1_6_5_n7) );
  MUX2_X1 pe_1_6_5_U64 ( .A(pe_1_6_5_int_q_reg_v[20]), .B(
        pe_1_6_5_int_q_reg_v[16]), .S(pe_1_6_5_n55), .Z(pe_1_6_5_n6) );
  MUX2_X1 pe_1_6_5_U63 ( .A(pe_1_6_5_int_q_reg_v[12]), .B(
        pe_1_6_5_int_q_reg_v[8]), .S(pe_1_6_5_n55), .Z(pe_1_6_5_n5) );
  MUX2_X1 pe_1_6_5_U62 ( .A(pe_1_6_5_int_q_reg_v[4]), .B(
        pe_1_6_5_int_q_reg_v[0]), .S(pe_1_6_5_n55), .Z(pe_1_6_5_n4) );
  AOI222_X1 pe_1_6_5_U61 ( .A1(int_data_res_7__5__2_), .A2(pe_1_6_5_n64), .B1(
        pe_1_6_5_N80), .B2(pe_1_6_5_n27), .C1(pe_1_6_5_N72), .C2(pe_1_6_5_n28), 
        .ZN(pe_1_6_5_n33) );
  INV_X1 pe_1_6_5_U60 ( .A(pe_1_6_5_n33), .ZN(pe_1_6_5_n82) );
  AOI222_X1 pe_1_6_5_U59 ( .A1(int_data_res_7__5__6_), .A2(pe_1_6_5_n64), .B1(
        pe_1_6_5_N84), .B2(pe_1_6_5_n27), .C1(pe_1_6_5_N76), .C2(pe_1_6_5_n28), 
        .ZN(pe_1_6_5_n29) );
  INV_X1 pe_1_6_5_U58 ( .A(pe_1_6_5_n29), .ZN(pe_1_6_5_n78) );
  XNOR2_X1 pe_1_6_5_U57 ( .A(pe_1_6_5_n73), .B(int_data_res_6__5__0_), .ZN(
        pe_1_6_5_N70) );
  AOI222_X1 pe_1_6_5_U52 ( .A1(int_data_res_7__5__0_), .A2(pe_1_6_5_n64), .B1(
        pe_1_6_5_n1), .B2(pe_1_6_5_n27), .C1(pe_1_6_5_N70), .C2(pe_1_6_5_n28), 
        .ZN(pe_1_6_5_n35) );
  INV_X1 pe_1_6_5_U51 ( .A(pe_1_6_5_n35), .ZN(pe_1_6_5_n84) );
  AOI222_X1 pe_1_6_5_U50 ( .A1(int_data_res_7__5__1_), .A2(pe_1_6_5_n64), .B1(
        pe_1_6_5_N79), .B2(pe_1_6_5_n27), .C1(pe_1_6_5_N71), .C2(pe_1_6_5_n28), 
        .ZN(pe_1_6_5_n34) );
  INV_X1 pe_1_6_5_U49 ( .A(pe_1_6_5_n34), .ZN(pe_1_6_5_n83) );
  AOI222_X1 pe_1_6_5_U48 ( .A1(int_data_res_7__5__3_), .A2(pe_1_6_5_n64), .B1(
        pe_1_6_5_N81), .B2(pe_1_6_5_n27), .C1(pe_1_6_5_N73), .C2(pe_1_6_5_n28), 
        .ZN(pe_1_6_5_n32) );
  INV_X1 pe_1_6_5_U47 ( .A(pe_1_6_5_n32), .ZN(pe_1_6_5_n81) );
  AOI222_X1 pe_1_6_5_U46 ( .A1(int_data_res_7__5__4_), .A2(pe_1_6_5_n64), .B1(
        pe_1_6_5_N82), .B2(pe_1_6_5_n27), .C1(pe_1_6_5_N74), .C2(pe_1_6_5_n28), 
        .ZN(pe_1_6_5_n31) );
  INV_X1 pe_1_6_5_U45 ( .A(pe_1_6_5_n31), .ZN(pe_1_6_5_n80) );
  AOI222_X1 pe_1_6_5_U44 ( .A1(int_data_res_7__5__5_), .A2(pe_1_6_5_n64), .B1(
        pe_1_6_5_N83), .B2(pe_1_6_5_n27), .C1(pe_1_6_5_N75), .C2(pe_1_6_5_n28), 
        .ZN(pe_1_6_5_n30) );
  INV_X1 pe_1_6_5_U43 ( .A(pe_1_6_5_n30), .ZN(pe_1_6_5_n79) );
  NAND2_X1 pe_1_6_5_U42 ( .A1(pe_1_6_5_int_data_0_), .A2(pe_1_6_5_n3), .ZN(
        pe_1_6_5_sub_81_carry[1]) );
  INV_X1 pe_1_6_5_U41 ( .A(pe_1_6_5_int_data_1_), .ZN(pe_1_6_5_n74) );
  INV_X1 pe_1_6_5_U40 ( .A(pe_1_6_5_int_data_2_), .ZN(pe_1_6_5_n75) );
  AND2_X1 pe_1_6_5_U39 ( .A1(pe_1_6_5_int_data_0_), .A2(int_data_res_6__5__0_), 
        .ZN(pe_1_6_5_n2) );
  AOI222_X1 pe_1_6_5_U38 ( .A1(pe_1_6_5_n64), .A2(int_data_res_7__5__7_), .B1(
        pe_1_6_5_N85), .B2(pe_1_6_5_n27), .C1(pe_1_6_5_N77), .C2(pe_1_6_5_n28), 
        .ZN(pe_1_6_5_n26) );
  INV_X1 pe_1_6_5_U37 ( .A(pe_1_6_5_n26), .ZN(pe_1_6_5_n77) );
  NOR3_X1 pe_1_6_5_U36 ( .A1(pe_1_6_5_n59), .A2(pe_1_6_5_n65), .A3(int_ckg[10]), .ZN(pe_1_6_5_n36) );
  OR2_X1 pe_1_6_5_U35 ( .A1(pe_1_6_5_n36), .A2(pe_1_6_5_n64), .ZN(pe_1_6_5_N90) );
  INV_X1 pe_1_6_5_U34 ( .A(n41), .ZN(pe_1_6_5_n63) );
  AND2_X1 pe_1_6_5_U33 ( .A1(int_data_x_6__5__2_), .A2(pe_1_6_5_n58), .ZN(
        pe_1_6_5_int_data_2_) );
  AND2_X1 pe_1_6_5_U32 ( .A1(int_data_x_6__5__1_), .A2(pe_1_6_5_n58), .ZN(
        pe_1_6_5_int_data_1_) );
  AND2_X1 pe_1_6_5_U31 ( .A1(int_data_x_6__5__3_), .A2(pe_1_6_5_n58), .ZN(
        pe_1_6_5_int_data_3_) );
  BUF_X1 pe_1_6_5_U30 ( .A(n63), .Z(pe_1_6_5_n64) );
  INV_X1 pe_1_6_5_U29 ( .A(n35), .ZN(pe_1_6_5_n61) );
  AND2_X1 pe_1_6_5_U28 ( .A1(int_data_x_6__5__0_), .A2(pe_1_6_5_n58), .ZN(
        pe_1_6_5_int_data_0_) );
  NAND2_X1 pe_1_6_5_U27 ( .A1(pe_1_6_5_n44), .A2(pe_1_6_5_n61), .ZN(
        pe_1_6_5_n41) );
  AND3_X1 pe_1_6_5_U26 ( .A1(n77), .A2(pe_1_6_5_n63), .A3(n53), .ZN(
        pe_1_6_5_n44) );
  INV_X1 pe_1_6_5_U25 ( .A(pe_1_6_5_int_data_3_), .ZN(pe_1_6_5_n76) );
  NOR2_X1 pe_1_6_5_U24 ( .A1(pe_1_6_5_n70), .A2(n53), .ZN(pe_1_6_5_n43) );
  NOR2_X1 pe_1_6_5_U23 ( .A1(pe_1_6_5_n57), .A2(pe_1_6_5_n64), .ZN(
        pe_1_6_5_n28) );
  NOR2_X1 pe_1_6_5_U22 ( .A1(n21), .A2(pe_1_6_5_n64), .ZN(pe_1_6_5_n27) );
  INV_X1 pe_1_6_5_U21 ( .A(pe_1_6_5_int_data_0_), .ZN(pe_1_6_5_n73) );
  INV_X1 pe_1_6_5_U20 ( .A(pe_1_6_5_n41), .ZN(pe_1_6_5_n90) );
  INV_X1 pe_1_6_5_U19 ( .A(pe_1_6_5_n37), .ZN(pe_1_6_5_n88) );
  INV_X1 pe_1_6_5_U18 ( .A(pe_1_6_5_n38), .ZN(pe_1_6_5_n87) );
  INV_X1 pe_1_6_5_U17 ( .A(pe_1_6_5_n39), .ZN(pe_1_6_5_n86) );
  NOR2_X1 pe_1_6_5_U16 ( .A1(pe_1_6_5_n68), .A2(pe_1_6_5_n42), .ZN(
        pe_1_6_5_N59) );
  NOR2_X1 pe_1_6_5_U15 ( .A1(pe_1_6_5_n68), .A2(pe_1_6_5_n41), .ZN(
        pe_1_6_5_N60) );
  NOR2_X1 pe_1_6_5_U14 ( .A1(pe_1_6_5_n68), .A2(pe_1_6_5_n38), .ZN(
        pe_1_6_5_N63) );
  NOR2_X1 pe_1_6_5_U13 ( .A1(pe_1_6_5_n67), .A2(pe_1_6_5_n40), .ZN(
        pe_1_6_5_N61) );
  NOR2_X1 pe_1_6_5_U12 ( .A1(pe_1_6_5_n67), .A2(pe_1_6_5_n39), .ZN(
        pe_1_6_5_N62) );
  NOR2_X1 pe_1_6_5_U11 ( .A1(pe_1_6_5_n37), .A2(pe_1_6_5_n67), .ZN(
        pe_1_6_5_N64) );
  NAND2_X1 pe_1_6_5_U10 ( .A1(pe_1_6_5_n44), .A2(pe_1_6_5_n60), .ZN(
        pe_1_6_5_n42) );
  BUF_X1 pe_1_6_5_U9 ( .A(pe_1_6_5_n60), .Z(pe_1_6_5_n55) );
  INV_X1 pe_1_6_5_U8 ( .A(pe_1_6_5_n69), .ZN(pe_1_6_5_n65) );
  BUF_X1 pe_1_6_5_U7 ( .A(pe_1_6_5_n60), .Z(pe_1_6_5_n56) );
  INV_X1 pe_1_6_5_U6 ( .A(pe_1_6_5_n42), .ZN(pe_1_6_5_n89) );
  INV_X1 pe_1_6_5_U5 ( .A(pe_1_6_5_n40), .ZN(pe_1_6_5_n85) );
  INV_X2 pe_1_6_5_U4 ( .A(n85), .ZN(pe_1_6_5_n72) );
  XOR2_X1 pe_1_6_5_U3 ( .A(pe_1_6_5_int_data_0_), .B(int_data_res_6__5__0_), 
        .Z(pe_1_6_5_n1) );
  DFFR_X1 pe_1_6_5_int_q_acc_reg_0_ ( .D(pe_1_6_5_n84), .CK(pe_1_6_5_net3418), 
        .RN(pe_1_6_5_n72), .Q(int_data_res_6__5__0_), .QN(pe_1_6_5_n3) );
  DFFR_X1 pe_1_6_5_int_q_reg_v_reg_0__0_ ( .D(int_data_y_7__5__0_), .CK(
        pe_1_6_5_net3388), .RN(pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_v[20]) );
  DFFR_X1 pe_1_6_5_int_q_reg_v_reg_0__1_ ( .D(int_data_y_7__5__1_), .CK(
        pe_1_6_5_net3388), .RN(pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_v[21]) );
  DFFR_X1 pe_1_6_5_int_q_reg_v_reg_0__2_ ( .D(int_data_y_7__5__2_), .CK(
        pe_1_6_5_net3388), .RN(pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_v[22]) );
  DFFR_X1 pe_1_6_5_int_q_reg_v_reg_0__3_ ( .D(int_data_y_7__5__3_), .CK(
        pe_1_6_5_net3388), .RN(pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_v[23]) );
  DFFR_X1 pe_1_6_5_int_q_reg_v_reg_1__0_ ( .D(int_data_y_7__5__0_), .CK(
        pe_1_6_5_net3393), .RN(pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_v[16]) );
  DFFR_X1 pe_1_6_5_int_q_reg_v_reg_1__1_ ( .D(int_data_y_7__5__1_), .CK(
        pe_1_6_5_net3393), .RN(pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_v[17]) );
  DFFR_X1 pe_1_6_5_int_q_reg_v_reg_1__2_ ( .D(int_data_y_7__5__2_), .CK(
        pe_1_6_5_net3393), .RN(pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_v[18]) );
  DFFR_X1 pe_1_6_5_int_q_reg_v_reg_1__3_ ( .D(int_data_y_7__5__3_), .CK(
        pe_1_6_5_net3393), .RN(pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_v[19]) );
  DFFR_X1 pe_1_6_5_int_q_reg_v_reg_2__0_ ( .D(int_data_y_7__5__0_), .CK(
        pe_1_6_5_net3398), .RN(pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_v[12]) );
  DFFR_X1 pe_1_6_5_int_q_reg_v_reg_2__1_ ( .D(int_data_y_7__5__1_), .CK(
        pe_1_6_5_net3398), .RN(pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_v[13]) );
  DFFR_X1 pe_1_6_5_int_q_reg_v_reg_2__2_ ( .D(int_data_y_7__5__2_), .CK(
        pe_1_6_5_net3398), .RN(pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_v[14]) );
  DFFR_X1 pe_1_6_5_int_q_reg_v_reg_2__3_ ( .D(int_data_y_7__5__3_), .CK(
        pe_1_6_5_net3398), .RN(pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_v[15]) );
  DFFR_X1 pe_1_6_5_int_q_reg_v_reg_3__0_ ( .D(int_data_y_7__5__0_), .CK(
        pe_1_6_5_net3403), .RN(pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_v[8]) );
  DFFR_X1 pe_1_6_5_int_q_reg_v_reg_3__1_ ( .D(int_data_y_7__5__1_), .CK(
        pe_1_6_5_net3403), .RN(pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_v[9]) );
  DFFR_X1 pe_1_6_5_int_q_reg_v_reg_3__2_ ( .D(int_data_y_7__5__2_), .CK(
        pe_1_6_5_net3403), .RN(pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_v[10]) );
  DFFR_X1 pe_1_6_5_int_q_reg_v_reg_3__3_ ( .D(int_data_y_7__5__3_), .CK(
        pe_1_6_5_net3403), .RN(pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_v[11]) );
  DFFR_X1 pe_1_6_5_int_q_reg_v_reg_4__0_ ( .D(int_data_y_7__5__0_), .CK(
        pe_1_6_5_net3408), .RN(pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_v[4]) );
  DFFR_X1 pe_1_6_5_int_q_reg_v_reg_4__1_ ( .D(int_data_y_7__5__1_), .CK(
        pe_1_6_5_net3408), .RN(pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_v[5]) );
  DFFR_X1 pe_1_6_5_int_q_reg_v_reg_4__2_ ( .D(int_data_y_7__5__2_), .CK(
        pe_1_6_5_net3408), .RN(pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_v[6]) );
  DFFR_X1 pe_1_6_5_int_q_reg_v_reg_4__3_ ( .D(int_data_y_7__5__3_), .CK(
        pe_1_6_5_net3408), .RN(pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_v[7]) );
  DFFR_X1 pe_1_6_5_int_q_reg_v_reg_5__0_ ( .D(int_data_y_7__5__0_), .CK(
        pe_1_6_5_net3413), .RN(pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_v[0]) );
  DFFR_X1 pe_1_6_5_int_q_reg_v_reg_5__1_ ( .D(int_data_y_7__5__1_), .CK(
        pe_1_6_5_net3413), .RN(pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_v[1]) );
  DFFR_X1 pe_1_6_5_int_q_reg_v_reg_5__2_ ( .D(int_data_y_7__5__2_), .CK(
        pe_1_6_5_net3413), .RN(pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_v[2]) );
  DFFR_X1 pe_1_6_5_int_q_reg_v_reg_5__3_ ( .D(int_data_y_7__5__3_), .CK(
        pe_1_6_5_net3413), .RN(pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_6_5_int_q_reg_h_reg_0__0_ ( .D(int_data_x_6__6__0_), .SI(
        int_data_y_7__5__0_), .SE(pe_1_6_5_n65), .CK(pe_1_6_5_net3357), .RN(
        pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_6_5_int_q_reg_h_reg_0__1_ ( .D(int_data_x_6__6__1_), .SI(
        int_data_y_7__5__1_), .SE(pe_1_6_5_n65), .CK(pe_1_6_5_net3357), .RN(
        pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_6_5_int_q_reg_h_reg_0__2_ ( .D(int_data_x_6__6__2_), .SI(
        int_data_y_7__5__2_), .SE(pe_1_6_5_n65), .CK(pe_1_6_5_net3357), .RN(
        pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_6_5_int_q_reg_h_reg_0__3_ ( .D(int_data_x_6__6__3_), .SI(
        int_data_y_7__5__3_), .SE(pe_1_6_5_n65), .CK(pe_1_6_5_net3357), .RN(
        pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_6_5_int_q_reg_h_reg_1__0_ ( .D(int_data_x_6__6__0_), .SI(
        int_data_y_7__5__0_), .SE(pe_1_6_5_n65), .CK(pe_1_6_5_net3363), .RN(
        pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_6_5_int_q_reg_h_reg_1__1_ ( .D(int_data_x_6__6__1_), .SI(
        int_data_y_7__5__1_), .SE(pe_1_6_5_n65), .CK(pe_1_6_5_net3363), .RN(
        pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_6_5_int_q_reg_h_reg_1__2_ ( .D(int_data_x_6__6__2_), .SI(
        int_data_y_7__5__2_), .SE(pe_1_6_5_n65), .CK(pe_1_6_5_net3363), .RN(
        pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_6_5_int_q_reg_h_reg_1__3_ ( .D(int_data_x_6__6__3_), .SI(
        int_data_y_7__5__3_), .SE(pe_1_6_5_n65), .CK(pe_1_6_5_net3363), .RN(
        pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_6_5_int_q_reg_h_reg_2__0_ ( .D(int_data_x_6__6__0_), .SI(
        int_data_y_7__5__0_), .SE(pe_1_6_5_n65), .CK(pe_1_6_5_net3368), .RN(
        pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_6_5_int_q_reg_h_reg_2__1_ ( .D(int_data_x_6__6__1_), .SI(
        int_data_y_7__5__1_), .SE(pe_1_6_5_n65), .CK(pe_1_6_5_net3368), .RN(
        pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_6_5_int_q_reg_h_reg_2__2_ ( .D(int_data_x_6__6__2_), .SI(
        int_data_y_7__5__2_), .SE(pe_1_6_5_n65), .CK(pe_1_6_5_net3368), .RN(
        pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_6_5_int_q_reg_h_reg_2__3_ ( .D(int_data_x_6__6__3_), .SI(
        int_data_y_7__5__3_), .SE(pe_1_6_5_n65), .CK(pe_1_6_5_net3368), .RN(
        pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_6_5_int_q_reg_h_reg_3__0_ ( .D(int_data_x_6__6__0_), .SI(
        int_data_y_7__5__0_), .SE(pe_1_6_5_n65), .CK(pe_1_6_5_net3373), .RN(
        pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_6_5_int_q_reg_h_reg_3__1_ ( .D(int_data_x_6__6__1_), .SI(
        int_data_y_7__5__1_), .SE(pe_1_6_5_n65), .CK(pe_1_6_5_net3373), .RN(
        pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_6_5_int_q_reg_h_reg_3__2_ ( .D(int_data_x_6__6__2_), .SI(
        int_data_y_7__5__2_), .SE(pe_1_6_5_n65), .CK(pe_1_6_5_net3373), .RN(
        pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_6_5_int_q_reg_h_reg_3__3_ ( .D(int_data_x_6__6__3_), .SI(
        int_data_y_7__5__3_), .SE(pe_1_6_5_n65), .CK(pe_1_6_5_net3373), .RN(
        pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_6_5_int_q_reg_h_reg_4__0_ ( .D(int_data_x_6__6__0_), .SI(
        int_data_y_7__5__0_), .SE(pe_1_6_5_n66), .CK(pe_1_6_5_net3378), .RN(
        pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_6_5_int_q_reg_h_reg_4__1_ ( .D(int_data_x_6__6__1_), .SI(
        int_data_y_7__5__1_), .SE(pe_1_6_5_n66), .CK(pe_1_6_5_net3378), .RN(
        pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_6_5_int_q_reg_h_reg_4__2_ ( .D(int_data_x_6__6__2_), .SI(
        int_data_y_7__5__2_), .SE(pe_1_6_5_n66), .CK(pe_1_6_5_net3378), .RN(
        pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_6_5_int_q_reg_h_reg_4__3_ ( .D(int_data_x_6__6__3_), .SI(
        int_data_y_7__5__3_), .SE(pe_1_6_5_n66), .CK(pe_1_6_5_net3378), .RN(
        pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_6_5_int_q_reg_h_reg_5__0_ ( .D(int_data_x_6__6__0_), .SI(
        int_data_y_7__5__0_), .SE(pe_1_6_5_n66), .CK(pe_1_6_5_net3383), .RN(
        pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_6_5_int_q_reg_h_reg_5__1_ ( .D(int_data_x_6__6__1_), .SI(
        int_data_y_7__5__1_), .SE(pe_1_6_5_n66), .CK(pe_1_6_5_net3383), .RN(
        pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_6_5_int_q_reg_h_reg_5__2_ ( .D(int_data_x_6__6__2_), .SI(
        int_data_y_7__5__2_), .SE(pe_1_6_5_n66), .CK(pe_1_6_5_net3383), .RN(
        pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_6_5_int_q_reg_h_reg_5__3_ ( .D(int_data_x_6__6__3_), .SI(
        int_data_y_7__5__3_), .SE(pe_1_6_5_n66), .CK(pe_1_6_5_net3383), .RN(
        pe_1_6_5_n72), .Q(pe_1_6_5_int_q_reg_h[3]) );
  FA_X1 pe_1_6_5_sub_81_U2_7 ( .A(int_data_res_6__5__7_), .B(pe_1_6_5_n76), 
        .CI(pe_1_6_5_sub_81_carry[7]), .S(pe_1_6_5_N77) );
  FA_X1 pe_1_6_5_sub_81_U2_6 ( .A(int_data_res_6__5__6_), .B(pe_1_6_5_n76), 
        .CI(pe_1_6_5_sub_81_carry[6]), .CO(pe_1_6_5_sub_81_carry[7]), .S(
        pe_1_6_5_N76) );
  FA_X1 pe_1_6_5_sub_81_U2_5 ( .A(int_data_res_6__5__5_), .B(pe_1_6_5_n76), 
        .CI(pe_1_6_5_sub_81_carry[5]), .CO(pe_1_6_5_sub_81_carry[6]), .S(
        pe_1_6_5_N75) );
  FA_X1 pe_1_6_5_sub_81_U2_4 ( .A(int_data_res_6__5__4_), .B(pe_1_6_5_n76), 
        .CI(pe_1_6_5_sub_81_carry[4]), .CO(pe_1_6_5_sub_81_carry[5]), .S(
        pe_1_6_5_N74) );
  FA_X1 pe_1_6_5_sub_81_U2_3 ( .A(int_data_res_6__5__3_), .B(pe_1_6_5_n76), 
        .CI(pe_1_6_5_sub_81_carry[3]), .CO(pe_1_6_5_sub_81_carry[4]), .S(
        pe_1_6_5_N73) );
  FA_X1 pe_1_6_5_sub_81_U2_2 ( .A(int_data_res_6__5__2_), .B(pe_1_6_5_n75), 
        .CI(pe_1_6_5_sub_81_carry[2]), .CO(pe_1_6_5_sub_81_carry[3]), .S(
        pe_1_6_5_N72) );
  FA_X1 pe_1_6_5_sub_81_U2_1 ( .A(int_data_res_6__5__1_), .B(pe_1_6_5_n74), 
        .CI(pe_1_6_5_sub_81_carry[1]), .CO(pe_1_6_5_sub_81_carry[2]), .S(
        pe_1_6_5_N71) );
  FA_X1 pe_1_6_5_add_83_U1_7 ( .A(int_data_res_6__5__7_), .B(
        pe_1_6_5_int_data_3_), .CI(pe_1_6_5_add_83_carry[7]), .S(pe_1_6_5_N85)
         );
  FA_X1 pe_1_6_5_add_83_U1_6 ( .A(int_data_res_6__5__6_), .B(
        pe_1_6_5_int_data_3_), .CI(pe_1_6_5_add_83_carry[6]), .CO(
        pe_1_6_5_add_83_carry[7]), .S(pe_1_6_5_N84) );
  FA_X1 pe_1_6_5_add_83_U1_5 ( .A(int_data_res_6__5__5_), .B(
        pe_1_6_5_int_data_3_), .CI(pe_1_6_5_add_83_carry[5]), .CO(
        pe_1_6_5_add_83_carry[6]), .S(pe_1_6_5_N83) );
  FA_X1 pe_1_6_5_add_83_U1_4 ( .A(int_data_res_6__5__4_), .B(
        pe_1_6_5_int_data_3_), .CI(pe_1_6_5_add_83_carry[4]), .CO(
        pe_1_6_5_add_83_carry[5]), .S(pe_1_6_5_N82) );
  FA_X1 pe_1_6_5_add_83_U1_3 ( .A(int_data_res_6__5__3_), .B(
        pe_1_6_5_int_data_3_), .CI(pe_1_6_5_add_83_carry[3]), .CO(
        pe_1_6_5_add_83_carry[4]), .S(pe_1_6_5_N81) );
  FA_X1 pe_1_6_5_add_83_U1_2 ( .A(int_data_res_6__5__2_), .B(
        pe_1_6_5_int_data_2_), .CI(pe_1_6_5_add_83_carry[2]), .CO(
        pe_1_6_5_add_83_carry[3]), .S(pe_1_6_5_N80) );
  FA_X1 pe_1_6_5_add_83_U1_1 ( .A(int_data_res_6__5__1_), .B(
        pe_1_6_5_int_data_1_), .CI(pe_1_6_5_n2), .CO(pe_1_6_5_add_83_carry[2]), 
        .S(pe_1_6_5_N79) );
  NAND3_X1 pe_1_6_5_U56 ( .A1(pe_1_6_5_n60), .A2(pe_1_6_5_n43), .A3(
        pe_1_6_5_n62), .ZN(pe_1_6_5_n40) );
  NAND3_X1 pe_1_6_5_U55 ( .A1(pe_1_6_5_n43), .A2(pe_1_6_5_n61), .A3(
        pe_1_6_5_n62), .ZN(pe_1_6_5_n39) );
  NAND3_X1 pe_1_6_5_U54 ( .A1(pe_1_6_5_n43), .A2(pe_1_6_5_n63), .A3(
        pe_1_6_5_n60), .ZN(pe_1_6_5_n38) );
  NAND3_X1 pe_1_6_5_U53 ( .A1(pe_1_6_5_n61), .A2(pe_1_6_5_n63), .A3(
        pe_1_6_5_n43), .ZN(pe_1_6_5_n37) );
  DFFR_X1 pe_1_6_5_int_q_acc_reg_6_ ( .D(pe_1_6_5_n78), .CK(pe_1_6_5_net3418), 
        .RN(pe_1_6_5_n71), .Q(int_data_res_6__5__6_) );
  DFFR_X1 pe_1_6_5_int_q_acc_reg_5_ ( .D(pe_1_6_5_n79), .CK(pe_1_6_5_net3418), 
        .RN(pe_1_6_5_n71), .Q(int_data_res_6__5__5_) );
  DFFR_X1 pe_1_6_5_int_q_acc_reg_4_ ( .D(pe_1_6_5_n80), .CK(pe_1_6_5_net3418), 
        .RN(pe_1_6_5_n71), .Q(int_data_res_6__5__4_) );
  DFFR_X1 pe_1_6_5_int_q_acc_reg_3_ ( .D(pe_1_6_5_n81), .CK(pe_1_6_5_net3418), 
        .RN(pe_1_6_5_n71), .Q(int_data_res_6__5__3_) );
  DFFR_X1 pe_1_6_5_int_q_acc_reg_2_ ( .D(pe_1_6_5_n82), .CK(pe_1_6_5_net3418), 
        .RN(pe_1_6_5_n71), .Q(int_data_res_6__5__2_) );
  DFFR_X1 pe_1_6_5_int_q_acc_reg_1_ ( .D(pe_1_6_5_n83), .CK(pe_1_6_5_net3418), 
        .RN(pe_1_6_5_n71), .Q(int_data_res_6__5__1_) );
  DFFR_X1 pe_1_6_5_int_q_acc_reg_7_ ( .D(pe_1_6_5_n77), .CK(pe_1_6_5_net3418), 
        .RN(pe_1_6_5_n71), .Q(int_data_res_6__5__7_) );
  CLKGATETST_X1 pe_1_6_5_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_6_5_n88), .SE(1'b0), .GCK(pe_1_6_5_net3357) );
  CLKGATETST_X1 pe_1_6_5_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_6_5_n87), .SE(1'b0), .GCK(pe_1_6_5_net3363) );
  CLKGATETST_X1 pe_1_6_5_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_6_5_n86), .SE(1'b0), .GCK(pe_1_6_5_net3368) );
  CLKGATETST_X1 pe_1_6_5_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_6_5_n85), .SE(1'b0), .GCK(pe_1_6_5_net3373) );
  CLKGATETST_X1 pe_1_6_5_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_6_5_n90), .SE(1'b0), .GCK(pe_1_6_5_net3378) );
  CLKGATETST_X1 pe_1_6_5_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_6_5_n89), .SE(1'b0), .GCK(pe_1_6_5_net3383) );
  CLKGATETST_X1 pe_1_6_5_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_6_5_N64), .SE(1'b0), .GCK(pe_1_6_5_net3388) );
  CLKGATETST_X1 pe_1_6_5_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_6_5_N63), .SE(1'b0), .GCK(pe_1_6_5_net3393) );
  CLKGATETST_X1 pe_1_6_5_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_6_5_N62), .SE(1'b0), .GCK(pe_1_6_5_net3398) );
  CLKGATETST_X1 pe_1_6_5_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_6_5_N61), .SE(1'b0), .GCK(pe_1_6_5_net3403) );
  CLKGATETST_X1 pe_1_6_5_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_6_5_N60), .SE(1'b0), .GCK(pe_1_6_5_net3408) );
  CLKGATETST_X1 pe_1_6_5_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_6_5_N59), .SE(1'b0), .GCK(pe_1_6_5_net3413) );
  CLKGATETST_X1 pe_1_6_5_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_6_5_N90), .SE(1'b0), .GCK(pe_1_6_5_net3418) );
  CLKBUF_X1 pe_1_6_6_U112 ( .A(pe_1_6_6_n72), .Z(pe_1_6_6_n71) );
  INV_X1 pe_1_6_6_U111 ( .A(n77), .ZN(pe_1_6_6_n70) );
  INV_X1 pe_1_6_6_U110 ( .A(n69), .ZN(pe_1_6_6_n69) );
  INV_X1 pe_1_6_6_U109 ( .A(n69), .ZN(pe_1_6_6_n68) );
  INV_X1 pe_1_6_6_U108 ( .A(n69), .ZN(pe_1_6_6_n67) );
  INV_X1 pe_1_6_6_U107 ( .A(pe_1_6_6_n69), .ZN(pe_1_6_6_n66) );
  INV_X1 pe_1_6_6_U106 ( .A(pe_1_6_6_n63), .ZN(pe_1_6_6_n62) );
  INV_X1 pe_1_6_6_U105 ( .A(pe_1_6_6_n61), .ZN(pe_1_6_6_n60) );
  INV_X1 pe_1_6_6_U104 ( .A(n29), .ZN(pe_1_6_6_n59) );
  INV_X1 pe_1_6_6_U103 ( .A(pe_1_6_6_n59), .ZN(pe_1_6_6_n58) );
  INV_X1 pe_1_6_6_U102 ( .A(n21), .ZN(pe_1_6_6_n57) );
  MUX2_X1 pe_1_6_6_U101 ( .A(pe_1_6_6_n54), .B(pe_1_6_6_n51), .S(n53), .Z(
        int_data_x_6__6__3_) );
  MUX2_X1 pe_1_6_6_U100 ( .A(pe_1_6_6_n53), .B(pe_1_6_6_n52), .S(pe_1_6_6_n62), 
        .Z(pe_1_6_6_n54) );
  MUX2_X1 pe_1_6_6_U99 ( .A(pe_1_6_6_int_q_reg_h[23]), .B(
        pe_1_6_6_int_q_reg_h[19]), .S(pe_1_6_6_n56), .Z(pe_1_6_6_n53) );
  MUX2_X1 pe_1_6_6_U98 ( .A(pe_1_6_6_int_q_reg_h[15]), .B(
        pe_1_6_6_int_q_reg_h[11]), .S(pe_1_6_6_n56), .Z(pe_1_6_6_n52) );
  MUX2_X1 pe_1_6_6_U97 ( .A(pe_1_6_6_int_q_reg_h[7]), .B(
        pe_1_6_6_int_q_reg_h[3]), .S(pe_1_6_6_n56), .Z(pe_1_6_6_n51) );
  MUX2_X1 pe_1_6_6_U96 ( .A(pe_1_6_6_n50), .B(pe_1_6_6_n47), .S(n53), .Z(
        int_data_x_6__6__2_) );
  MUX2_X1 pe_1_6_6_U95 ( .A(pe_1_6_6_n49), .B(pe_1_6_6_n48), .S(pe_1_6_6_n62), 
        .Z(pe_1_6_6_n50) );
  MUX2_X1 pe_1_6_6_U94 ( .A(pe_1_6_6_int_q_reg_h[22]), .B(
        pe_1_6_6_int_q_reg_h[18]), .S(pe_1_6_6_n56), .Z(pe_1_6_6_n49) );
  MUX2_X1 pe_1_6_6_U93 ( .A(pe_1_6_6_int_q_reg_h[14]), .B(
        pe_1_6_6_int_q_reg_h[10]), .S(pe_1_6_6_n56), .Z(pe_1_6_6_n48) );
  MUX2_X1 pe_1_6_6_U92 ( .A(pe_1_6_6_int_q_reg_h[6]), .B(
        pe_1_6_6_int_q_reg_h[2]), .S(pe_1_6_6_n56), .Z(pe_1_6_6_n47) );
  MUX2_X1 pe_1_6_6_U91 ( .A(pe_1_6_6_n46), .B(pe_1_6_6_n24), .S(n53), .Z(
        int_data_x_6__6__1_) );
  MUX2_X1 pe_1_6_6_U90 ( .A(pe_1_6_6_n45), .B(pe_1_6_6_n25), .S(pe_1_6_6_n62), 
        .Z(pe_1_6_6_n46) );
  MUX2_X1 pe_1_6_6_U89 ( .A(pe_1_6_6_int_q_reg_h[21]), .B(
        pe_1_6_6_int_q_reg_h[17]), .S(pe_1_6_6_n56), .Z(pe_1_6_6_n45) );
  MUX2_X1 pe_1_6_6_U88 ( .A(pe_1_6_6_int_q_reg_h[13]), .B(
        pe_1_6_6_int_q_reg_h[9]), .S(pe_1_6_6_n56), .Z(pe_1_6_6_n25) );
  MUX2_X1 pe_1_6_6_U87 ( .A(pe_1_6_6_int_q_reg_h[5]), .B(
        pe_1_6_6_int_q_reg_h[1]), .S(pe_1_6_6_n56), .Z(pe_1_6_6_n24) );
  MUX2_X1 pe_1_6_6_U86 ( .A(pe_1_6_6_n23), .B(pe_1_6_6_n20), .S(n53), .Z(
        int_data_x_6__6__0_) );
  MUX2_X1 pe_1_6_6_U85 ( .A(pe_1_6_6_n22), .B(pe_1_6_6_n21), .S(pe_1_6_6_n62), 
        .Z(pe_1_6_6_n23) );
  MUX2_X1 pe_1_6_6_U84 ( .A(pe_1_6_6_int_q_reg_h[20]), .B(
        pe_1_6_6_int_q_reg_h[16]), .S(pe_1_6_6_n56), .Z(pe_1_6_6_n22) );
  MUX2_X1 pe_1_6_6_U83 ( .A(pe_1_6_6_int_q_reg_h[12]), .B(
        pe_1_6_6_int_q_reg_h[8]), .S(pe_1_6_6_n56), .Z(pe_1_6_6_n21) );
  MUX2_X1 pe_1_6_6_U82 ( .A(pe_1_6_6_int_q_reg_h[4]), .B(
        pe_1_6_6_int_q_reg_h[0]), .S(pe_1_6_6_n56), .Z(pe_1_6_6_n20) );
  MUX2_X1 pe_1_6_6_U81 ( .A(pe_1_6_6_n19), .B(pe_1_6_6_n16), .S(n53), .Z(
        int_data_y_6__6__3_) );
  MUX2_X1 pe_1_6_6_U80 ( .A(pe_1_6_6_n18), .B(pe_1_6_6_n17), .S(pe_1_6_6_n62), 
        .Z(pe_1_6_6_n19) );
  MUX2_X1 pe_1_6_6_U79 ( .A(pe_1_6_6_int_q_reg_v[23]), .B(
        pe_1_6_6_int_q_reg_v[19]), .S(pe_1_6_6_n55), .Z(pe_1_6_6_n18) );
  MUX2_X1 pe_1_6_6_U78 ( .A(pe_1_6_6_int_q_reg_v[15]), .B(
        pe_1_6_6_int_q_reg_v[11]), .S(pe_1_6_6_n55), .Z(pe_1_6_6_n17) );
  MUX2_X1 pe_1_6_6_U77 ( .A(pe_1_6_6_int_q_reg_v[7]), .B(
        pe_1_6_6_int_q_reg_v[3]), .S(pe_1_6_6_n55), .Z(pe_1_6_6_n16) );
  MUX2_X1 pe_1_6_6_U76 ( .A(pe_1_6_6_n15), .B(pe_1_6_6_n12), .S(n53), .Z(
        int_data_y_6__6__2_) );
  MUX2_X1 pe_1_6_6_U75 ( .A(pe_1_6_6_n14), .B(pe_1_6_6_n13), .S(pe_1_6_6_n62), 
        .Z(pe_1_6_6_n15) );
  MUX2_X1 pe_1_6_6_U74 ( .A(pe_1_6_6_int_q_reg_v[22]), .B(
        pe_1_6_6_int_q_reg_v[18]), .S(pe_1_6_6_n55), .Z(pe_1_6_6_n14) );
  MUX2_X1 pe_1_6_6_U73 ( .A(pe_1_6_6_int_q_reg_v[14]), .B(
        pe_1_6_6_int_q_reg_v[10]), .S(pe_1_6_6_n55), .Z(pe_1_6_6_n13) );
  MUX2_X1 pe_1_6_6_U72 ( .A(pe_1_6_6_int_q_reg_v[6]), .B(
        pe_1_6_6_int_q_reg_v[2]), .S(pe_1_6_6_n55), .Z(pe_1_6_6_n12) );
  MUX2_X1 pe_1_6_6_U71 ( .A(pe_1_6_6_n11), .B(pe_1_6_6_n8), .S(n53), .Z(
        int_data_y_6__6__1_) );
  MUX2_X1 pe_1_6_6_U70 ( .A(pe_1_6_6_n10), .B(pe_1_6_6_n9), .S(pe_1_6_6_n62), 
        .Z(pe_1_6_6_n11) );
  MUX2_X1 pe_1_6_6_U69 ( .A(pe_1_6_6_int_q_reg_v[21]), .B(
        pe_1_6_6_int_q_reg_v[17]), .S(pe_1_6_6_n55), .Z(pe_1_6_6_n10) );
  MUX2_X1 pe_1_6_6_U68 ( .A(pe_1_6_6_int_q_reg_v[13]), .B(
        pe_1_6_6_int_q_reg_v[9]), .S(pe_1_6_6_n55), .Z(pe_1_6_6_n9) );
  MUX2_X1 pe_1_6_6_U67 ( .A(pe_1_6_6_int_q_reg_v[5]), .B(
        pe_1_6_6_int_q_reg_v[1]), .S(pe_1_6_6_n55), .Z(pe_1_6_6_n8) );
  MUX2_X1 pe_1_6_6_U66 ( .A(pe_1_6_6_n7), .B(pe_1_6_6_n4), .S(n53), .Z(
        int_data_y_6__6__0_) );
  MUX2_X1 pe_1_6_6_U65 ( .A(pe_1_6_6_n6), .B(pe_1_6_6_n5), .S(pe_1_6_6_n62), 
        .Z(pe_1_6_6_n7) );
  MUX2_X1 pe_1_6_6_U64 ( .A(pe_1_6_6_int_q_reg_v[20]), .B(
        pe_1_6_6_int_q_reg_v[16]), .S(pe_1_6_6_n55), .Z(pe_1_6_6_n6) );
  MUX2_X1 pe_1_6_6_U63 ( .A(pe_1_6_6_int_q_reg_v[12]), .B(
        pe_1_6_6_int_q_reg_v[8]), .S(pe_1_6_6_n55), .Z(pe_1_6_6_n5) );
  MUX2_X1 pe_1_6_6_U62 ( .A(pe_1_6_6_int_q_reg_v[4]), .B(
        pe_1_6_6_int_q_reg_v[0]), .S(pe_1_6_6_n55), .Z(pe_1_6_6_n4) );
  AOI222_X1 pe_1_6_6_U61 ( .A1(int_data_res_7__6__2_), .A2(pe_1_6_6_n64), .B1(
        pe_1_6_6_N80), .B2(pe_1_6_6_n27), .C1(pe_1_6_6_N72), .C2(pe_1_6_6_n28), 
        .ZN(pe_1_6_6_n33) );
  INV_X1 pe_1_6_6_U60 ( .A(pe_1_6_6_n33), .ZN(pe_1_6_6_n82) );
  AOI222_X1 pe_1_6_6_U59 ( .A1(int_data_res_7__6__6_), .A2(pe_1_6_6_n64), .B1(
        pe_1_6_6_N84), .B2(pe_1_6_6_n27), .C1(pe_1_6_6_N76), .C2(pe_1_6_6_n28), 
        .ZN(pe_1_6_6_n29) );
  INV_X1 pe_1_6_6_U58 ( .A(pe_1_6_6_n29), .ZN(pe_1_6_6_n78) );
  XNOR2_X1 pe_1_6_6_U57 ( .A(pe_1_6_6_n73), .B(int_data_res_6__6__0_), .ZN(
        pe_1_6_6_N70) );
  AOI222_X1 pe_1_6_6_U52 ( .A1(int_data_res_7__6__0_), .A2(pe_1_6_6_n64), .B1(
        pe_1_6_6_n1), .B2(pe_1_6_6_n27), .C1(pe_1_6_6_N70), .C2(pe_1_6_6_n28), 
        .ZN(pe_1_6_6_n35) );
  INV_X1 pe_1_6_6_U51 ( .A(pe_1_6_6_n35), .ZN(pe_1_6_6_n84) );
  AOI222_X1 pe_1_6_6_U50 ( .A1(int_data_res_7__6__1_), .A2(pe_1_6_6_n64), .B1(
        pe_1_6_6_N79), .B2(pe_1_6_6_n27), .C1(pe_1_6_6_N71), .C2(pe_1_6_6_n28), 
        .ZN(pe_1_6_6_n34) );
  INV_X1 pe_1_6_6_U49 ( .A(pe_1_6_6_n34), .ZN(pe_1_6_6_n83) );
  AOI222_X1 pe_1_6_6_U48 ( .A1(int_data_res_7__6__3_), .A2(pe_1_6_6_n64), .B1(
        pe_1_6_6_N81), .B2(pe_1_6_6_n27), .C1(pe_1_6_6_N73), .C2(pe_1_6_6_n28), 
        .ZN(pe_1_6_6_n32) );
  INV_X1 pe_1_6_6_U47 ( .A(pe_1_6_6_n32), .ZN(pe_1_6_6_n81) );
  AOI222_X1 pe_1_6_6_U46 ( .A1(int_data_res_7__6__4_), .A2(pe_1_6_6_n64), .B1(
        pe_1_6_6_N82), .B2(pe_1_6_6_n27), .C1(pe_1_6_6_N74), .C2(pe_1_6_6_n28), 
        .ZN(pe_1_6_6_n31) );
  INV_X1 pe_1_6_6_U45 ( .A(pe_1_6_6_n31), .ZN(pe_1_6_6_n80) );
  AOI222_X1 pe_1_6_6_U44 ( .A1(int_data_res_7__6__5_), .A2(pe_1_6_6_n64), .B1(
        pe_1_6_6_N83), .B2(pe_1_6_6_n27), .C1(pe_1_6_6_N75), .C2(pe_1_6_6_n28), 
        .ZN(pe_1_6_6_n30) );
  INV_X1 pe_1_6_6_U43 ( .A(pe_1_6_6_n30), .ZN(pe_1_6_6_n79) );
  NAND2_X1 pe_1_6_6_U42 ( .A1(pe_1_6_6_int_data_0_), .A2(pe_1_6_6_n3), .ZN(
        pe_1_6_6_sub_81_carry[1]) );
  INV_X1 pe_1_6_6_U41 ( .A(pe_1_6_6_int_data_1_), .ZN(pe_1_6_6_n74) );
  INV_X1 pe_1_6_6_U40 ( .A(pe_1_6_6_int_data_2_), .ZN(pe_1_6_6_n75) );
  AND2_X1 pe_1_6_6_U39 ( .A1(pe_1_6_6_int_data_0_), .A2(int_data_res_6__6__0_), 
        .ZN(pe_1_6_6_n2) );
  AOI222_X1 pe_1_6_6_U38 ( .A1(pe_1_6_6_n64), .A2(int_data_res_7__6__7_), .B1(
        pe_1_6_6_N85), .B2(pe_1_6_6_n27), .C1(pe_1_6_6_N77), .C2(pe_1_6_6_n28), 
        .ZN(pe_1_6_6_n26) );
  INV_X1 pe_1_6_6_U37 ( .A(pe_1_6_6_n26), .ZN(pe_1_6_6_n77) );
  NOR3_X1 pe_1_6_6_U36 ( .A1(pe_1_6_6_n59), .A2(pe_1_6_6_n65), .A3(int_ckg[9]), 
        .ZN(pe_1_6_6_n36) );
  OR2_X1 pe_1_6_6_U35 ( .A1(pe_1_6_6_n36), .A2(pe_1_6_6_n64), .ZN(pe_1_6_6_N90) );
  INV_X1 pe_1_6_6_U34 ( .A(n41), .ZN(pe_1_6_6_n63) );
  AND2_X1 pe_1_6_6_U33 ( .A1(int_data_x_6__6__2_), .A2(pe_1_6_6_n58), .ZN(
        pe_1_6_6_int_data_2_) );
  AND2_X1 pe_1_6_6_U32 ( .A1(int_data_x_6__6__1_), .A2(pe_1_6_6_n58), .ZN(
        pe_1_6_6_int_data_1_) );
  AND2_X1 pe_1_6_6_U31 ( .A1(int_data_x_6__6__3_), .A2(pe_1_6_6_n58), .ZN(
        pe_1_6_6_int_data_3_) );
  BUF_X1 pe_1_6_6_U30 ( .A(n63), .Z(pe_1_6_6_n64) );
  INV_X1 pe_1_6_6_U29 ( .A(n35), .ZN(pe_1_6_6_n61) );
  AND2_X1 pe_1_6_6_U28 ( .A1(int_data_x_6__6__0_), .A2(pe_1_6_6_n58), .ZN(
        pe_1_6_6_int_data_0_) );
  NAND2_X1 pe_1_6_6_U27 ( .A1(pe_1_6_6_n44), .A2(pe_1_6_6_n61), .ZN(
        pe_1_6_6_n41) );
  AND3_X1 pe_1_6_6_U26 ( .A1(n77), .A2(pe_1_6_6_n63), .A3(n53), .ZN(
        pe_1_6_6_n44) );
  INV_X1 pe_1_6_6_U25 ( .A(pe_1_6_6_int_data_3_), .ZN(pe_1_6_6_n76) );
  NOR2_X1 pe_1_6_6_U24 ( .A1(pe_1_6_6_n70), .A2(n53), .ZN(pe_1_6_6_n43) );
  NOR2_X1 pe_1_6_6_U23 ( .A1(pe_1_6_6_n57), .A2(pe_1_6_6_n64), .ZN(
        pe_1_6_6_n28) );
  NOR2_X1 pe_1_6_6_U22 ( .A1(n21), .A2(pe_1_6_6_n64), .ZN(pe_1_6_6_n27) );
  INV_X1 pe_1_6_6_U21 ( .A(pe_1_6_6_int_data_0_), .ZN(pe_1_6_6_n73) );
  INV_X1 pe_1_6_6_U20 ( .A(pe_1_6_6_n41), .ZN(pe_1_6_6_n90) );
  INV_X1 pe_1_6_6_U19 ( .A(pe_1_6_6_n37), .ZN(pe_1_6_6_n88) );
  INV_X1 pe_1_6_6_U18 ( .A(pe_1_6_6_n38), .ZN(pe_1_6_6_n87) );
  INV_X1 pe_1_6_6_U17 ( .A(pe_1_6_6_n39), .ZN(pe_1_6_6_n86) );
  NOR2_X1 pe_1_6_6_U16 ( .A1(pe_1_6_6_n68), .A2(pe_1_6_6_n42), .ZN(
        pe_1_6_6_N59) );
  NOR2_X1 pe_1_6_6_U15 ( .A1(pe_1_6_6_n68), .A2(pe_1_6_6_n41), .ZN(
        pe_1_6_6_N60) );
  NOR2_X1 pe_1_6_6_U14 ( .A1(pe_1_6_6_n68), .A2(pe_1_6_6_n38), .ZN(
        pe_1_6_6_N63) );
  NOR2_X1 pe_1_6_6_U13 ( .A1(pe_1_6_6_n67), .A2(pe_1_6_6_n40), .ZN(
        pe_1_6_6_N61) );
  NOR2_X1 pe_1_6_6_U12 ( .A1(pe_1_6_6_n67), .A2(pe_1_6_6_n39), .ZN(
        pe_1_6_6_N62) );
  NOR2_X1 pe_1_6_6_U11 ( .A1(pe_1_6_6_n37), .A2(pe_1_6_6_n67), .ZN(
        pe_1_6_6_N64) );
  NAND2_X1 pe_1_6_6_U10 ( .A1(pe_1_6_6_n44), .A2(pe_1_6_6_n60), .ZN(
        pe_1_6_6_n42) );
  BUF_X1 pe_1_6_6_U9 ( .A(pe_1_6_6_n60), .Z(pe_1_6_6_n55) );
  INV_X1 pe_1_6_6_U8 ( .A(pe_1_6_6_n69), .ZN(pe_1_6_6_n65) );
  BUF_X1 pe_1_6_6_U7 ( .A(pe_1_6_6_n60), .Z(pe_1_6_6_n56) );
  INV_X1 pe_1_6_6_U6 ( .A(pe_1_6_6_n42), .ZN(pe_1_6_6_n89) );
  INV_X1 pe_1_6_6_U5 ( .A(pe_1_6_6_n40), .ZN(pe_1_6_6_n85) );
  INV_X2 pe_1_6_6_U4 ( .A(n85), .ZN(pe_1_6_6_n72) );
  XOR2_X1 pe_1_6_6_U3 ( .A(pe_1_6_6_int_data_0_), .B(int_data_res_6__6__0_), 
        .Z(pe_1_6_6_n1) );
  DFFR_X1 pe_1_6_6_int_q_acc_reg_0_ ( .D(pe_1_6_6_n84), .CK(pe_1_6_6_net3340), 
        .RN(pe_1_6_6_n72), .Q(int_data_res_6__6__0_), .QN(pe_1_6_6_n3) );
  DFFR_X1 pe_1_6_6_int_q_reg_v_reg_0__0_ ( .D(int_data_y_7__6__0_), .CK(
        pe_1_6_6_net3310), .RN(pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_v[20]) );
  DFFR_X1 pe_1_6_6_int_q_reg_v_reg_0__1_ ( .D(int_data_y_7__6__1_), .CK(
        pe_1_6_6_net3310), .RN(pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_v[21]) );
  DFFR_X1 pe_1_6_6_int_q_reg_v_reg_0__2_ ( .D(int_data_y_7__6__2_), .CK(
        pe_1_6_6_net3310), .RN(pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_v[22]) );
  DFFR_X1 pe_1_6_6_int_q_reg_v_reg_0__3_ ( .D(int_data_y_7__6__3_), .CK(
        pe_1_6_6_net3310), .RN(pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_v[23]) );
  DFFR_X1 pe_1_6_6_int_q_reg_v_reg_1__0_ ( .D(int_data_y_7__6__0_), .CK(
        pe_1_6_6_net3315), .RN(pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_v[16]) );
  DFFR_X1 pe_1_6_6_int_q_reg_v_reg_1__1_ ( .D(int_data_y_7__6__1_), .CK(
        pe_1_6_6_net3315), .RN(pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_v[17]) );
  DFFR_X1 pe_1_6_6_int_q_reg_v_reg_1__2_ ( .D(int_data_y_7__6__2_), .CK(
        pe_1_6_6_net3315), .RN(pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_v[18]) );
  DFFR_X1 pe_1_6_6_int_q_reg_v_reg_1__3_ ( .D(int_data_y_7__6__3_), .CK(
        pe_1_6_6_net3315), .RN(pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_v[19]) );
  DFFR_X1 pe_1_6_6_int_q_reg_v_reg_2__0_ ( .D(int_data_y_7__6__0_), .CK(
        pe_1_6_6_net3320), .RN(pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_v[12]) );
  DFFR_X1 pe_1_6_6_int_q_reg_v_reg_2__1_ ( .D(int_data_y_7__6__1_), .CK(
        pe_1_6_6_net3320), .RN(pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_v[13]) );
  DFFR_X1 pe_1_6_6_int_q_reg_v_reg_2__2_ ( .D(int_data_y_7__6__2_), .CK(
        pe_1_6_6_net3320), .RN(pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_v[14]) );
  DFFR_X1 pe_1_6_6_int_q_reg_v_reg_2__3_ ( .D(int_data_y_7__6__3_), .CK(
        pe_1_6_6_net3320), .RN(pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_v[15]) );
  DFFR_X1 pe_1_6_6_int_q_reg_v_reg_3__0_ ( .D(int_data_y_7__6__0_), .CK(
        pe_1_6_6_net3325), .RN(pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_v[8]) );
  DFFR_X1 pe_1_6_6_int_q_reg_v_reg_3__1_ ( .D(int_data_y_7__6__1_), .CK(
        pe_1_6_6_net3325), .RN(pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_v[9]) );
  DFFR_X1 pe_1_6_6_int_q_reg_v_reg_3__2_ ( .D(int_data_y_7__6__2_), .CK(
        pe_1_6_6_net3325), .RN(pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_v[10]) );
  DFFR_X1 pe_1_6_6_int_q_reg_v_reg_3__3_ ( .D(int_data_y_7__6__3_), .CK(
        pe_1_6_6_net3325), .RN(pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_v[11]) );
  DFFR_X1 pe_1_6_6_int_q_reg_v_reg_4__0_ ( .D(int_data_y_7__6__0_), .CK(
        pe_1_6_6_net3330), .RN(pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_v[4]) );
  DFFR_X1 pe_1_6_6_int_q_reg_v_reg_4__1_ ( .D(int_data_y_7__6__1_), .CK(
        pe_1_6_6_net3330), .RN(pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_v[5]) );
  DFFR_X1 pe_1_6_6_int_q_reg_v_reg_4__2_ ( .D(int_data_y_7__6__2_), .CK(
        pe_1_6_6_net3330), .RN(pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_v[6]) );
  DFFR_X1 pe_1_6_6_int_q_reg_v_reg_4__3_ ( .D(int_data_y_7__6__3_), .CK(
        pe_1_6_6_net3330), .RN(pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_v[7]) );
  DFFR_X1 pe_1_6_6_int_q_reg_v_reg_5__0_ ( .D(int_data_y_7__6__0_), .CK(
        pe_1_6_6_net3335), .RN(pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_v[0]) );
  DFFR_X1 pe_1_6_6_int_q_reg_v_reg_5__1_ ( .D(int_data_y_7__6__1_), .CK(
        pe_1_6_6_net3335), .RN(pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_v[1]) );
  DFFR_X1 pe_1_6_6_int_q_reg_v_reg_5__2_ ( .D(int_data_y_7__6__2_), .CK(
        pe_1_6_6_net3335), .RN(pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_v[2]) );
  DFFR_X1 pe_1_6_6_int_q_reg_v_reg_5__3_ ( .D(int_data_y_7__6__3_), .CK(
        pe_1_6_6_net3335), .RN(pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_6_6_int_q_reg_h_reg_0__0_ ( .D(int_data_x_6__7__0_), .SI(
        int_data_y_7__6__0_), .SE(pe_1_6_6_n65), .CK(pe_1_6_6_net3279), .RN(
        pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_6_6_int_q_reg_h_reg_0__1_ ( .D(int_data_x_6__7__1_), .SI(
        int_data_y_7__6__1_), .SE(pe_1_6_6_n65), .CK(pe_1_6_6_net3279), .RN(
        pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_6_6_int_q_reg_h_reg_0__2_ ( .D(int_data_x_6__7__2_), .SI(
        int_data_y_7__6__2_), .SE(pe_1_6_6_n65), .CK(pe_1_6_6_net3279), .RN(
        pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_6_6_int_q_reg_h_reg_0__3_ ( .D(int_data_x_6__7__3_), .SI(
        int_data_y_7__6__3_), .SE(pe_1_6_6_n65), .CK(pe_1_6_6_net3279), .RN(
        pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_6_6_int_q_reg_h_reg_1__0_ ( .D(int_data_x_6__7__0_), .SI(
        int_data_y_7__6__0_), .SE(pe_1_6_6_n65), .CK(pe_1_6_6_net3285), .RN(
        pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_6_6_int_q_reg_h_reg_1__1_ ( .D(int_data_x_6__7__1_), .SI(
        int_data_y_7__6__1_), .SE(pe_1_6_6_n65), .CK(pe_1_6_6_net3285), .RN(
        pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_6_6_int_q_reg_h_reg_1__2_ ( .D(int_data_x_6__7__2_), .SI(
        int_data_y_7__6__2_), .SE(pe_1_6_6_n65), .CK(pe_1_6_6_net3285), .RN(
        pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_6_6_int_q_reg_h_reg_1__3_ ( .D(int_data_x_6__7__3_), .SI(
        int_data_y_7__6__3_), .SE(pe_1_6_6_n65), .CK(pe_1_6_6_net3285), .RN(
        pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_6_6_int_q_reg_h_reg_2__0_ ( .D(int_data_x_6__7__0_), .SI(
        int_data_y_7__6__0_), .SE(pe_1_6_6_n65), .CK(pe_1_6_6_net3290), .RN(
        pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_6_6_int_q_reg_h_reg_2__1_ ( .D(int_data_x_6__7__1_), .SI(
        int_data_y_7__6__1_), .SE(pe_1_6_6_n65), .CK(pe_1_6_6_net3290), .RN(
        pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_6_6_int_q_reg_h_reg_2__2_ ( .D(int_data_x_6__7__2_), .SI(
        int_data_y_7__6__2_), .SE(pe_1_6_6_n65), .CK(pe_1_6_6_net3290), .RN(
        pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_6_6_int_q_reg_h_reg_2__3_ ( .D(int_data_x_6__7__3_), .SI(
        int_data_y_7__6__3_), .SE(pe_1_6_6_n65), .CK(pe_1_6_6_net3290), .RN(
        pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_6_6_int_q_reg_h_reg_3__0_ ( .D(int_data_x_6__7__0_), .SI(
        int_data_y_7__6__0_), .SE(pe_1_6_6_n65), .CK(pe_1_6_6_net3295), .RN(
        pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_6_6_int_q_reg_h_reg_3__1_ ( .D(int_data_x_6__7__1_), .SI(
        int_data_y_7__6__1_), .SE(pe_1_6_6_n65), .CK(pe_1_6_6_net3295), .RN(
        pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_6_6_int_q_reg_h_reg_3__2_ ( .D(int_data_x_6__7__2_), .SI(
        int_data_y_7__6__2_), .SE(pe_1_6_6_n65), .CK(pe_1_6_6_net3295), .RN(
        pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_6_6_int_q_reg_h_reg_3__3_ ( .D(int_data_x_6__7__3_), .SI(
        int_data_y_7__6__3_), .SE(pe_1_6_6_n65), .CK(pe_1_6_6_net3295), .RN(
        pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_6_6_int_q_reg_h_reg_4__0_ ( .D(int_data_x_6__7__0_), .SI(
        int_data_y_7__6__0_), .SE(pe_1_6_6_n66), .CK(pe_1_6_6_net3300), .RN(
        pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_6_6_int_q_reg_h_reg_4__1_ ( .D(int_data_x_6__7__1_), .SI(
        int_data_y_7__6__1_), .SE(pe_1_6_6_n66), .CK(pe_1_6_6_net3300), .RN(
        pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_6_6_int_q_reg_h_reg_4__2_ ( .D(int_data_x_6__7__2_), .SI(
        int_data_y_7__6__2_), .SE(pe_1_6_6_n66), .CK(pe_1_6_6_net3300), .RN(
        pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_6_6_int_q_reg_h_reg_4__3_ ( .D(int_data_x_6__7__3_), .SI(
        int_data_y_7__6__3_), .SE(pe_1_6_6_n66), .CK(pe_1_6_6_net3300), .RN(
        pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_6_6_int_q_reg_h_reg_5__0_ ( .D(int_data_x_6__7__0_), .SI(
        int_data_y_7__6__0_), .SE(pe_1_6_6_n66), .CK(pe_1_6_6_net3305), .RN(
        pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_6_6_int_q_reg_h_reg_5__1_ ( .D(int_data_x_6__7__1_), .SI(
        int_data_y_7__6__1_), .SE(pe_1_6_6_n66), .CK(pe_1_6_6_net3305), .RN(
        pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_6_6_int_q_reg_h_reg_5__2_ ( .D(int_data_x_6__7__2_), .SI(
        int_data_y_7__6__2_), .SE(pe_1_6_6_n66), .CK(pe_1_6_6_net3305), .RN(
        pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_6_6_int_q_reg_h_reg_5__3_ ( .D(int_data_x_6__7__3_), .SI(
        int_data_y_7__6__3_), .SE(pe_1_6_6_n66), .CK(pe_1_6_6_net3305), .RN(
        pe_1_6_6_n72), .Q(pe_1_6_6_int_q_reg_h[3]) );
  FA_X1 pe_1_6_6_sub_81_U2_7 ( .A(int_data_res_6__6__7_), .B(pe_1_6_6_n76), 
        .CI(pe_1_6_6_sub_81_carry[7]), .S(pe_1_6_6_N77) );
  FA_X1 pe_1_6_6_sub_81_U2_6 ( .A(int_data_res_6__6__6_), .B(pe_1_6_6_n76), 
        .CI(pe_1_6_6_sub_81_carry[6]), .CO(pe_1_6_6_sub_81_carry[7]), .S(
        pe_1_6_6_N76) );
  FA_X1 pe_1_6_6_sub_81_U2_5 ( .A(int_data_res_6__6__5_), .B(pe_1_6_6_n76), 
        .CI(pe_1_6_6_sub_81_carry[5]), .CO(pe_1_6_6_sub_81_carry[6]), .S(
        pe_1_6_6_N75) );
  FA_X1 pe_1_6_6_sub_81_U2_4 ( .A(int_data_res_6__6__4_), .B(pe_1_6_6_n76), 
        .CI(pe_1_6_6_sub_81_carry[4]), .CO(pe_1_6_6_sub_81_carry[5]), .S(
        pe_1_6_6_N74) );
  FA_X1 pe_1_6_6_sub_81_U2_3 ( .A(int_data_res_6__6__3_), .B(pe_1_6_6_n76), 
        .CI(pe_1_6_6_sub_81_carry[3]), .CO(pe_1_6_6_sub_81_carry[4]), .S(
        pe_1_6_6_N73) );
  FA_X1 pe_1_6_6_sub_81_U2_2 ( .A(int_data_res_6__6__2_), .B(pe_1_6_6_n75), 
        .CI(pe_1_6_6_sub_81_carry[2]), .CO(pe_1_6_6_sub_81_carry[3]), .S(
        pe_1_6_6_N72) );
  FA_X1 pe_1_6_6_sub_81_U2_1 ( .A(int_data_res_6__6__1_), .B(pe_1_6_6_n74), 
        .CI(pe_1_6_6_sub_81_carry[1]), .CO(pe_1_6_6_sub_81_carry[2]), .S(
        pe_1_6_6_N71) );
  FA_X1 pe_1_6_6_add_83_U1_7 ( .A(int_data_res_6__6__7_), .B(
        pe_1_6_6_int_data_3_), .CI(pe_1_6_6_add_83_carry[7]), .S(pe_1_6_6_N85)
         );
  FA_X1 pe_1_6_6_add_83_U1_6 ( .A(int_data_res_6__6__6_), .B(
        pe_1_6_6_int_data_3_), .CI(pe_1_6_6_add_83_carry[6]), .CO(
        pe_1_6_6_add_83_carry[7]), .S(pe_1_6_6_N84) );
  FA_X1 pe_1_6_6_add_83_U1_5 ( .A(int_data_res_6__6__5_), .B(
        pe_1_6_6_int_data_3_), .CI(pe_1_6_6_add_83_carry[5]), .CO(
        pe_1_6_6_add_83_carry[6]), .S(pe_1_6_6_N83) );
  FA_X1 pe_1_6_6_add_83_U1_4 ( .A(int_data_res_6__6__4_), .B(
        pe_1_6_6_int_data_3_), .CI(pe_1_6_6_add_83_carry[4]), .CO(
        pe_1_6_6_add_83_carry[5]), .S(pe_1_6_6_N82) );
  FA_X1 pe_1_6_6_add_83_U1_3 ( .A(int_data_res_6__6__3_), .B(
        pe_1_6_6_int_data_3_), .CI(pe_1_6_6_add_83_carry[3]), .CO(
        pe_1_6_6_add_83_carry[4]), .S(pe_1_6_6_N81) );
  FA_X1 pe_1_6_6_add_83_U1_2 ( .A(int_data_res_6__6__2_), .B(
        pe_1_6_6_int_data_2_), .CI(pe_1_6_6_add_83_carry[2]), .CO(
        pe_1_6_6_add_83_carry[3]), .S(pe_1_6_6_N80) );
  FA_X1 pe_1_6_6_add_83_U1_1 ( .A(int_data_res_6__6__1_), .B(
        pe_1_6_6_int_data_1_), .CI(pe_1_6_6_n2), .CO(pe_1_6_6_add_83_carry[2]), 
        .S(pe_1_6_6_N79) );
  NAND3_X1 pe_1_6_6_U56 ( .A1(pe_1_6_6_n60), .A2(pe_1_6_6_n43), .A3(
        pe_1_6_6_n62), .ZN(pe_1_6_6_n40) );
  NAND3_X1 pe_1_6_6_U55 ( .A1(pe_1_6_6_n43), .A2(pe_1_6_6_n61), .A3(
        pe_1_6_6_n62), .ZN(pe_1_6_6_n39) );
  NAND3_X1 pe_1_6_6_U54 ( .A1(pe_1_6_6_n43), .A2(pe_1_6_6_n63), .A3(
        pe_1_6_6_n60), .ZN(pe_1_6_6_n38) );
  NAND3_X1 pe_1_6_6_U53 ( .A1(pe_1_6_6_n61), .A2(pe_1_6_6_n63), .A3(
        pe_1_6_6_n43), .ZN(pe_1_6_6_n37) );
  DFFR_X1 pe_1_6_6_int_q_acc_reg_6_ ( .D(pe_1_6_6_n78), .CK(pe_1_6_6_net3340), 
        .RN(pe_1_6_6_n71), .Q(int_data_res_6__6__6_) );
  DFFR_X1 pe_1_6_6_int_q_acc_reg_5_ ( .D(pe_1_6_6_n79), .CK(pe_1_6_6_net3340), 
        .RN(pe_1_6_6_n71), .Q(int_data_res_6__6__5_) );
  DFFR_X1 pe_1_6_6_int_q_acc_reg_4_ ( .D(pe_1_6_6_n80), .CK(pe_1_6_6_net3340), 
        .RN(pe_1_6_6_n71), .Q(int_data_res_6__6__4_) );
  DFFR_X1 pe_1_6_6_int_q_acc_reg_3_ ( .D(pe_1_6_6_n81), .CK(pe_1_6_6_net3340), 
        .RN(pe_1_6_6_n71), .Q(int_data_res_6__6__3_) );
  DFFR_X1 pe_1_6_6_int_q_acc_reg_2_ ( .D(pe_1_6_6_n82), .CK(pe_1_6_6_net3340), 
        .RN(pe_1_6_6_n71), .Q(int_data_res_6__6__2_) );
  DFFR_X1 pe_1_6_6_int_q_acc_reg_1_ ( .D(pe_1_6_6_n83), .CK(pe_1_6_6_net3340), 
        .RN(pe_1_6_6_n71), .Q(int_data_res_6__6__1_) );
  DFFR_X1 pe_1_6_6_int_q_acc_reg_7_ ( .D(pe_1_6_6_n77), .CK(pe_1_6_6_net3340), 
        .RN(pe_1_6_6_n71), .Q(int_data_res_6__6__7_) );
  CLKGATETST_X1 pe_1_6_6_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_6_6_n88), .SE(1'b0), .GCK(pe_1_6_6_net3279) );
  CLKGATETST_X1 pe_1_6_6_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_6_6_n87), .SE(1'b0), .GCK(pe_1_6_6_net3285) );
  CLKGATETST_X1 pe_1_6_6_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_6_6_n86), .SE(1'b0), .GCK(pe_1_6_6_net3290) );
  CLKGATETST_X1 pe_1_6_6_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_6_6_n85), .SE(1'b0), .GCK(pe_1_6_6_net3295) );
  CLKGATETST_X1 pe_1_6_6_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_6_6_n90), .SE(1'b0), .GCK(pe_1_6_6_net3300) );
  CLKGATETST_X1 pe_1_6_6_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_6_6_n89), .SE(1'b0), .GCK(pe_1_6_6_net3305) );
  CLKGATETST_X1 pe_1_6_6_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_6_6_N64), .SE(1'b0), .GCK(pe_1_6_6_net3310) );
  CLKGATETST_X1 pe_1_6_6_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_6_6_N63), .SE(1'b0), .GCK(pe_1_6_6_net3315) );
  CLKGATETST_X1 pe_1_6_6_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_6_6_N62), .SE(1'b0), .GCK(pe_1_6_6_net3320) );
  CLKGATETST_X1 pe_1_6_6_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_6_6_N61), .SE(1'b0), .GCK(pe_1_6_6_net3325) );
  CLKGATETST_X1 pe_1_6_6_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_6_6_N60), .SE(1'b0), .GCK(pe_1_6_6_net3330) );
  CLKGATETST_X1 pe_1_6_6_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_6_6_N59), .SE(1'b0), .GCK(pe_1_6_6_net3335) );
  CLKGATETST_X1 pe_1_6_6_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_6_6_N90), .SE(1'b0), .GCK(pe_1_6_6_net3340) );
  CLKBUF_X1 pe_1_6_7_U112 ( .A(pe_1_6_7_n72), .Z(pe_1_6_7_n71) );
  INV_X1 pe_1_6_7_U111 ( .A(n77), .ZN(pe_1_6_7_n70) );
  INV_X1 pe_1_6_7_U110 ( .A(n69), .ZN(pe_1_6_7_n69) );
  INV_X1 pe_1_6_7_U109 ( .A(n69), .ZN(pe_1_6_7_n68) );
  INV_X1 pe_1_6_7_U108 ( .A(n69), .ZN(pe_1_6_7_n67) );
  INV_X1 pe_1_6_7_U107 ( .A(pe_1_6_7_n69), .ZN(pe_1_6_7_n66) );
  INV_X1 pe_1_6_7_U106 ( .A(pe_1_6_7_n63), .ZN(pe_1_6_7_n62) );
  INV_X1 pe_1_6_7_U105 ( .A(pe_1_6_7_n61), .ZN(pe_1_6_7_n60) );
  INV_X1 pe_1_6_7_U104 ( .A(n29), .ZN(pe_1_6_7_n59) );
  INV_X1 pe_1_6_7_U103 ( .A(pe_1_6_7_n59), .ZN(pe_1_6_7_n58) );
  INV_X1 pe_1_6_7_U102 ( .A(n21), .ZN(pe_1_6_7_n57) );
  MUX2_X1 pe_1_6_7_U101 ( .A(pe_1_6_7_n54), .B(pe_1_6_7_n51), .S(n54), .Z(
        int_data_x_6__7__3_) );
  MUX2_X1 pe_1_6_7_U100 ( .A(pe_1_6_7_n53), .B(pe_1_6_7_n52), .S(pe_1_6_7_n62), 
        .Z(pe_1_6_7_n54) );
  MUX2_X1 pe_1_6_7_U99 ( .A(pe_1_6_7_int_q_reg_h[23]), .B(
        pe_1_6_7_int_q_reg_h[19]), .S(pe_1_6_7_n56), .Z(pe_1_6_7_n53) );
  MUX2_X1 pe_1_6_7_U98 ( .A(pe_1_6_7_int_q_reg_h[15]), .B(
        pe_1_6_7_int_q_reg_h[11]), .S(pe_1_6_7_n56), .Z(pe_1_6_7_n52) );
  MUX2_X1 pe_1_6_7_U97 ( .A(pe_1_6_7_int_q_reg_h[7]), .B(
        pe_1_6_7_int_q_reg_h[3]), .S(pe_1_6_7_n56), .Z(pe_1_6_7_n51) );
  MUX2_X1 pe_1_6_7_U96 ( .A(pe_1_6_7_n50), .B(pe_1_6_7_n47), .S(n54), .Z(
        int_data_x_6__7__2_) );
  MUX2_X1 pe_1_6_7_U95 ( .A(pe_1_6_7_n49), .B(pe_1_6_7_n48), .S(pe_1_6_7_n62), 
        .Z(pe_1_6_7_n50) );
  MUX2_X1 pe_1_6_7_U94 ( .A(pe_1_6_7_int_q_reg_h[22]), .B(
        pe_1_6_7_int_q_reg_h[18]), .S(pe_1_6_7_n56), .Z(pe_1_6_7_n49) );
  MUX2_X1 pe_1_6_7_U93 ( .A(pe_1_6_7_int_q_reg_h[14]), .B(
        pe_1_6_7_int_q_reg_h[10]), .S(pe_1_6_7_n56), .Z(pe_1_6_7_n48) );
  MUX2_X1 pe_1_6_7_U92 ( .A(pe_1_6_7_int_q_reg_h[6]), .B(
        pe_1_6_7_int_q_reg_h[2]), .S(pe_1_6_7_n56), .Z(pe_1_6_7_n47) );
  MUX2_X1 pe_1_6_7_U91 ( .A(pe_1_6_7_n46), .B(pe_1_6_7_n24), .S(n54), .Z(
        int_data_x_6__7__1_) );
  MUX2_X1 pe_1_6_7_U90 ( .A(pe_1_6_7_n45), .B(pe_1_6_7_n25), .S(pe_1_6_7_n62), 
        .Z(pe_1_6_7_n46) );
  MUX2_X1 pe_1_6_7_U89 ( .A(pe_1_6_7_int_q_reg_h[21]), .B(
        pe_1_6_7_int_q_reg_h[17]), .S(pe_1_6_7_n56), .Z(pe_1_6_7_n45) );
  MUX2_X1 pe_1_6_7_U88 ( .A(pe_1_6_7_int_q_reg_h[13]), .B(
        pe_1_6_7_int_q_reg_h[9]), .S(pe_1_6_7_n56), .Z(pe_1_6_7_n25) );
  MUX2_X1 pe_1_6_7_U87 ( .A(pe_1_6_7_int_q_reg_h[5]), .B(
        pe_1_6_7_int_q_reg_h[1]), .S(pe_1_6_7_n56), .Z(pe_1_6_7_n24) );
  MUX2_X1 pe_1_6_7_U86 ( .A(pe_1_6_7_n23), .B(pe_1_6_7_n20), .S(n54), .Z(
        int_data_x_6__7__0_) );
  MUX2_X1 pe_1_6_7_U85 ( .A(pe_1_6_7_n22), .B(pe_1_6_7_n21), .S(pe_1_6_7_n62), 
        .Z(pe_1_6_7_n23) );
  MUX2_X1 pe_1_6_7_U84 ( .A(pe_1_6_7_int_q_reg_h[20]), .B(
        pe_1_6_7_int_q_reg_h[16]), .S(pe_1_6_7_n56), .Z(pe_1_6_7_n22) );
  MUX2_X1 pe_1_6_7_U83 ( .A(pe_1_6_7_int_q_reg_h[12]), .B(
        pe_1_6_7_int_q_reg_h[8]), .S(pe_1_6_7_n56), .Z(pe_1_6_7_n21) );
  MUX2_X1 pe_1_6_7_U82 ( .A(pe_1_6_7_int_q_reg_h[4]), .B(
        pe_1_6_7_int_q_reg_h[0]), .S(pe_1_6_7_n56), .Z(pe_1_6_7_n20) );
  MUX2_X1 pe_1_6_7_U81 ( .A(pe_1_6_7_n19), .B(pe_1_6_7_n16), .S(n54), .Z(
        int_data_y_6__7__3_) );
  MUX2_X1 pe_1_6_7_U80 ( .A(pe_1_6_7_n18), .B(pe_1_6_7_n17), .S(pe_1_6_7_n62), 
        .Z(pe_1_6_7_n19) );
  MUX2_X1 pe_1_6_7_U79 ( .A(pe_1_6_7_int_q_reg_v[23]), .B(
        pe_1_6_7_int_q_reg_v[19]), .S(pe_1_6_7_n55), .Z(pe_1_6_7_n18) );
  MUX2_X1 pe_1_6_7_U78 ( .A(pe_1_6_7_int_q_reg_v[15]), .B(
        pe_1_6_7_int_q_reg_v[11]), .S(pe_1_6_7_n55), .Z(pe_1_6_7_n17) );
  MUX2_X1 pe_1_6_7_U77 ( .A(pe_1_6_7_int_q_reg_v[7]), .B(
        pe_1_6_7_int_q_reg_v[3]), .S(pe_1_6_7_n55), .Z(pe_1_6_7_n16) );
  MUX2_X1 pe_1_6_7_U76 ( .A(pe_1_6_7_n15), .B(pe_1_6_7_n12), .S(n54), .Z(
        int_data_y_6__7__2_) );
  MUX2_X1 pe_1_6_7_U75 ( .A(pe_1_6_7_n14), .B(pe_1_6_7_n13), .S(pe_1_6_7_n62), 
        .Z(pe_1_6_7_n15) );
  MUX2_X1 pe_1_6_7_U74 ( .A(pe_1_6_7_int_q_reg_v[22]), .B(
        pe_1_6_7_int_q_reg_v[18]), .S(pe_1_6_7_n55), .Z(pe_1_6_7_n14) );
  MUX2_X1 pe_1_6_7_U73 ( .A(pe_1_6_7_int_q_reg_v[14]), .B(
        pe_1_6_7_int_q_reg_v[10]), .S(pe_1_6_7_n55), .Z(pe_1_6_7_n13) );
  MUX2_X1 pe_1_6_7_U72 ( .A(pe_1_6_7_int_q_reg_v[6]), .B(
        pe_1_6_7_int_q_reg_v[2]), .S(pe_1_6_7_n55), .Z(pe_1_6_7_n12) );
  MUX2_X1 pe_1_6_7_U71 ( .A(pe_1_6_7_n11), .B(pe_1_6_7_n8), .S(n54), .Z(
        int_data_y_6__7__1_) );
  MUX2_X1 pe_1_6_7_U70 ( .A(pe_1_6_7_n10), .B(pe_1_6_7_n9), .S(pe_1_6_7_n62), 
        .Z(pe_1_6_7_n11) );
  MUX2_X1 pe_1_6_7_U69 ( .A(pe_1_6_7_int_q_reg_v[21]), .B(
        pe_1_6_7_int_q_reg_v[17]), .S(pe_1_6_7_n55), .Z(pe_1_6_7_n10) );
  MUX2_X1 pe_1_6_7_U68 ( .A(pe_1_6_7_int_q_reg_v[13]), .B(
        pe_1_6_7_int_q_reg_v[9]), .S(pe_1_6_7_n55), .Z(pe_1_6_7_n9) );
  MUX2_X1 pe_1_6_7_U67 ( .A(pe_1_6_7_int_q_reg_v[5]), .B(
        pe_1_6_7_int_q_reg_v[1]), .S(pe_1_6_7_n55), .Z(pe_1_6_7_n8) );
  MUX2_X1 pe_1_6_7_U66 ( .A(pe_1_6_7_n7), .B(pe_1_6_7_n4), .S(n54), .Z(
        int_data_y_6__7__0_) );
  MUX2_X1 pe_1_6_7_U65 ( .A(pe_1_6_7_n6), .B(pe_1_6_7_n5), .S(pe_1_6_7_n62), 
        .Z(pe_1_6_7_n7) );
  MUX2_X1 pe_1_6_7_U64 ( .A(pe_1_6_7_int_q_reg_v[20]), .B(
        pe_1_6_7_int_q_reg_v[16]), .S(pe_1_6_7_n55), .Z(pe_1_6_7_n6) );
  MUX2_X1 pe_1_6_7_U63 ( .A(pe_1_6_7_int_q_reg_v[12]), .B(
        pe_1_6_7_int_q_reg_v[8]), .S(pe_1_6_7_n55), .Z(pe_1_6_7_n5) );
  MUX2_X1 pe_1_6_7_U62 ( .A(pe_1_6_7_int_q_reg_v[4]), .B(
        pe_1_6_7_int_q_reg_v[0]), .S(pe_1_6_7_n55), .Z(pe_1_6_7_n4) );
  AOI222_X1 pe_1_6_7_U61 ( .A1(int_data_res_7__7__2_), .A2(pe_1_6_7_n64), .B1(
        pe_1_6_7_N80), .B2(pe_1_6_7_n27), .C1(pe_1_6_7_N72), .C2(pe_1_6_7_n28), 
        .ZN(pe_1_6_7_n33) );
  INV_X1 pe_1_6_7_U60 ( .A(pe_1_6_7_n33), .ZN(pe_1_6_7_n82) );
  AOI222_X1 pe_1_6_7_U59 ( .A1(int_data_res_7__7__6_), .A2(pe_1_6_7_n64), .B1(
        pe_1_6_7_N84), .B2(pe_1_6_7_n27), .C1(pe_1_6_7_N76), .C2(pe_1_6_7_n28), 
        .ZN(pe_1_6_7_n29) );
  INV_X1 pe_1_6_7_U58 ( .A(pe_1_6_7_n29), .ZN(pe_1_6_7_n78) );
  XNOR2_X1 pe_1_6_7_U57 ( .A(pe_1_6_7_n73), .B(int_data_res_6__7__0_), .ZN(
        pe_1_6_7_N70) );
  AOI222_X1 pe_1_6_7_U52 ( .A1(int_data_res_7__7__0_), .A2(pe_1_6_7_n64), .B1(
        pe_1_6_7_n1), .B2(pe_1_6_7_n27), .C1(pe_1_6_7_N70), .C2(pe_1_6_7_n28), 
        .ZN(pe_1_6_7_n35) );
  INV_X1 pe_1_6_7_U51 ( .A(pe_1_6_7_n35), .ZN(pe_1_6_7_n84) );
  AOI222_X1 pe_1_6_7_U50 ( .A1(int_data_res_7__7__1_), .A2(pe_1_6_7_n64), .B1(
        pe_1_6_7_N79), .B2(pe_1_6_7_n27), .C1(pe_1_6_7_N71), .C2(pe_1_6_7_n28), 
        .ZN(pe_1_6_7_n34) );
  INV_X1 pe_1_6_7_U49 ( .A(pe_1_6_7_n34), .ZN(pe_1_6_7_n83) );
  AOI222_X1 pe_1_6_7_U48 ( .A1(int_data_res_7__7__3_), .A2(pe_1_6_7_n64), .B1(
        pe_1_6_7_N81), .B2(pe_1_6_7_n27), .C1(pe_1_6_7_N73), .C2(pe_1_6_7_n28), 
        .ZN(pe_1_6_7_n32) );
  INV_X1 pe_1_6_7_U47 ( .A(pe_1_6_7_n32), .ZN(pe_1_6_7_n81) );
  AOI222_X1 pe_1_6_7_U46 ( .A1(int_data_res_7__7__4_), .A2(pe_1_6_7_n64), .B1(
        pe_1_6_7_N82), .B2(pe_1_6_7_n27), .C1(pe_1_6_7_N74), .C2(pe_1_6_7_n28), 
        .ZN(pe_1_6_7_n31) );
  INV_X1 pe_1_6_7_U45 ( .A(pe_1_6_7_n31), .ZN(pe_1_6_7_n80) );
  AOI222_X1 pe_1_6_7_U44 ( .A1(int_data_res_7__7__5_), .A2(pe_1_6_7_n64), .B1(
        pe_1_6_7_N83), .B2(pe_1_6_7_n27), .C1(pe_1_6_7_N75), .C2(pe_1_6_7_n28), 
        .ZN(pe_1_6_7_n30) );
  INV_X1 pe_1_6_7_U43 ( .A(pe_1_6_7_n30), .ZN(pe_1_6_7_n79) );
  NAND2_X1 pe_1_6_7_U42 ( .A1(pe_1_6_7_int_data_0_), .A2(pe_1_6_7_n3), .ZN(
        pe_1_6_7_sub_81_carry[1]) );
  INV_X1 pe_1_6_7_U41 ( .A(pe_1_6_7_int_data_1_), .ZN(pe_1_6_7_n74) );
  INV_X1 pe_1_6_7_U40 ( .A(pe_1_6_7_int_data_2_), .ZN(pe_1_6_7_n75) );
  AND2_X1 pe_1_6_7_U39 ( .A1(pe_1_6_7_int_data_0_), .A2(int_data_res_6__7__0_), 
        .ZN(pe_1_6_7_n2) );
  AOI222_X1 pe_1_6_7_U38 ( .A1(pe_1_6_7_n64), .A2(int_data_res_7__7__7_), .B1(
        pe_1_6_7_N85), .B2(pe_1_6_7_n27), .C1(pe_1_6_7_N77), .C2(pe_1_6_7_n28), 
        .ZN(pe_1_6_7_n26) );
  INV_X1 pe_1_6_7_U37 ( .A(pe_1_6_7_n26), .ZN(pe_1_6_7_n77) );
  NOR3_X1 pe_1_6_7_U36 ( .A1(pe_1_6_7_n59), .A2(pe_1_6_7_n65), .A3(int_ckg[8]), 
        .ZN(pe_1_6_7_n36) );
  OR2_X1 pe_1_6_7_U35 ( .A1(pe_1_6_7_n36), .A2(pe_1_6_7_n64), .ZN(pe_1_6_7_N90) );
  INV_X1 pe_1_6_7_U34 ( .A(n41), .ZN(pe_1_6_7_n63) );
  AND2_X1 pe_1_6_7_U33 ( .A1(int_data_x_6__7__2_), .A2(pe_1_6_7_n58), .ZN(
        pe_1_6_7_int_data_2_) );
  AND2_X1 pe_1_6_7_U32 ( .A1(int_data_x_6__7__1_), .A2(pe_1_6_7_n58), .ZN(
        pe_1_6_7_int_data_1_) );
  AND2_X1 pe_1_6_7_U31 ( .A1(int_data_x_6__7__3_), .A2(pe_1_6_7_n58), .ZN(
        pe_1_6_7_int_data_3_) );
  BUF_X1 pe_1_6_7_U30 ( .A(n63), .Z(pe_1_6_7_n64) );
  INV_X1 pe_1_6_7_U29 ( .A(n35), .ZN(pe_1_6_7_n61) );
  AND2_X1 pe_1_6_7_U28 ( .A1(int_data_x_6__7__0_), .A2(pe_1_6_7_n58), .ZN(
        pe_1_6_7_int_data_0_) );
  NAND2_X1 pe_1_6_7_U27 ( .A1(pe_1_6_7_n44), .A2(pe_1_6_7_n61), .ZN(
        pe_1_6_7_n41) );
  AND3_X1 pe_1_6_7_U26 ( .A1(n77), .A2(pe_1_6_7_n63), .A3(n54), .ZN(
        pe_1_6_7_n44) );
  INV_X1 pe_1_6_7_U25 ( .A(pe_1_6_7_int_data_3_), .ZN(pe_1_6_7_n76) );
  NOR2_X1 pe_1_6_7_U24 ( .A1(pe_1_6_7_n70), .A2(n54), .ZN(pe_1_6_7_n43) );
  NOR2_X1 pe_1_6_7_U23 ( .A1(pe_1_6_7_n57), .A2(pe_1_6_7_n64), .ZN(
        pe_1_6_7_n28) );
  NOR2_X1 pe_1_6_7_U22 ( .A1(n21), .A2(pe_1_6_7_n64), .ZN(pe_1_6_7_n27) );
  INV_X1 pe_1_6_7_U21 ( .A(pe_1_6_7_int_data_0_), .ZN(pe_1_6_7_n73) );
  INV_X1 pe_1_6_7_U20 ( .A(pe_1_6_7_n41), .ZN(pe_1_6_7_n90) );
  INV_X1 pe_1_6_7_U19 ( .A(pe_1_6_7_n37), .ZN(pe_1_6_7_n88) );
  INV_X1 pe_1_6_7_U18 ( .A(pe_1_6_7_n38), .ZN(pe_1_6_7_n87) );
  INV_X1 pe_1_6_7_U17 ( .A(pe_1_6_7_n39), .ZN(pe_1_6_7_n86) );
  NOR2_X1 pe_1_6_7_U16 ( .A1(pe_1_6_7_n68), .A2(pe_1_6_7_n42), .ZN(
        pe_1_6_7_N59) );
  NOR2_X1 pe_1_6_7_U15 ( .A1(pe_1_6_7_n68), .A2(pe_1_6_7_n41), .ZN(
        pe_1_6_7_N60) );
  NOR2_X1 pe_1_6_7_U14 ( .A1(pe_1_6_7_n68), .A2(pe_1_6_7_n38), .ZN(
        pe_1_6_7_N63) );
  NOR2_X1 pe_1_6_7_U13 ( .A1(pe_1_6_7_n67), .A2(pe_1_6_7_n40), .ZN(
        pe_1_6_7_N61) );
  NOR2_X1 pe_1_6_7_U12 ( .A1(pe_1_6_7_n67), .A2(pe_1_6_7_n39), .ZN(
        pe_1_6_7_N62) );
  NOR2_X1 pe_1_6_7_U11 ( .A1(pe_1_6_7_n37), .A2(pe_1_6_7_n67), .ZN(
        pe_1_6_7_N64) );
  NAND2_X1 pe_1_6_7_U10 ( .A1(pe_1_6_7_n44), .A2(pe_1_6_7_n60), .ZN(
        pe_1_6_7_n42) );
  BUF_X1 pe_1_6_7_U9 ( .A(pe_1_6_7_n60), .Z(pe_1_6_7_n55) );
  INV_X1 pe_1_6_7_U8 ( .A(pe_1_6_7_n69), .ZN(pe_1_6_7_n65) );
  BUF_X1 pe_1_6_7_U7 ( .A(pe_1_6_7_n60), .Z(pe_1_6_7_n56) );
  INV_X1 pe_1_6_7_U6 ( .A(pe_1_6_7_n42), .ZN(pe_1_6_7_n89) );
  INV_X1 pe_1_6_7_U5 ( .A(pe_1_6_7_n40), .ZN(pe_1_6_7_n85) );
  INV_X2 pe_1_6_7_U4 ( .A(n85), .ZN(pe_1_6_7_n72) );
  XOR2_X1 pe_1_6_7_U3 ( .A(pe_1_6_7_int_data_0_), .B(int_data_res_6__7__0_), 
        .Z(pe_1_6_7_n1) );
  DFFR_X1 pe_1_6_7_int_q_acc_reg_0_ ( .D(pe_1_6_7_n84), .CK(pe_1_6_7_net3262), 
        .RN(pe_1_6_7_n72), .Q(int_data_res_6__7__0_), .QN(pe_1_6_7_n3) );
  DFFR_X1 pe_1_6_7_int_q_reg_v_reg_0__0_ ( .D(int_data_y_7__7__0_), .CK(
        pe_1_6_7_net3232), .RN(pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_v[20]) );
  DFFR_X1 pe_1_6_7_int_q_reg_v_reg_0__1_ ( .D(int_data_y_7__7__1_), .CK(
        pe_1_6_7_net3232), .RN(pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_v[21]) );
  DFFR_X1 pe_1_6_7_int_q_reg_v_reg_0__2_ ( .D(int_data_y_7__7__2_), .CK(
        pe_1_6_7_net3232), .RN(pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_v[22]) );
  DFFR_X1 pe_1_6_7_int_q_reg_v_reg_0__3_ ( .D(int_data_y_7__7__3_), .CK(
        pe_1_6_7_net3232), .RN(pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_v[23]) );
  DFFR_X1 pe_1_6_7_int_q_reg_v_reg_1__0_ ( .D(int_data_y_7__7__0_), .CK(
        pe_1_6_7_net3237), .RN(pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_v[16]) );
  DFFR_X1 pe_1_6_7_int_q_reg_v_reg_1__1_ ( .D(int_data_y_7__7__1_), .CK(
        pe_1_6_7_net3237), .RN(pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_v[17]) );
  DFFR_X1 pe_1_6_7_int_q_reg_v_reg_1__2_ ( .D(int_data_y_7__7__2_), .CK(
        pe_1_6_7_net3237), .RN(pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_v[18]) );
  DFFR_X1 pe_1_6_7_int_q_reg_v_reg_1__3_ ( .D(int_data_y_7__7__3_), .CK(
        pe_1_6_7_net3237), .RN(pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_v[19]) );
  DFFR_X1 pe_1_6_7_int_q_reg_v_reg_2__0_ ( .D(int_data_y_7__7__0_), .CK(
        pe_1_6_7_net3242), .RN(pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_v[12]) );
  DFFR_X1 pe_1_6_7_int_q_reg_v_reg_2__1_ ( .D(int_data_y_7__7__1_), .CK(
        pe_1_6_7_net3242), .RN(pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_v[13]) );
  DFFR_X1 pe_1_6_7_int_q_reg_v_reg_2__2_ ( .D(int_data_y_7__7__2_), .CK(
        pe_1_6_7_net3242), .RN(pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_v[14]) );
  DFFR_X1 pe_1_6_7_int_q_reg_v_reg_2__3_ ( .D(int_data_y_7__7__3_), .CK(
        pe_1_6_7_net3242), .RN(pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_v[15]) );
  DFFR_X1 pe_1_6_7_int_q_reg_v_reg_3__0_ ( .D(int_data_y_7__7__0_), .CK(
        pe_1_6_7_net3247), .RN(pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_v[8]) );
  DFFR_X1 pe_1_6_7_int_q_reg_v_reg_3__1_ ( .D(int_data_y_7__7__1_), .CK(
        pe_1_6_7_net3247), .RN(pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_v[9]) );
  DFFR_X1 pe_1_6_7_int_q_reg_v_reg_3__2_ ( .D(int_data_y_7__7__2_), .CK(
        pe_1_6_7_net3247), .RN(pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_v[10]) );
  DFFR_X1 pe_1_6_7_int_q_reg_v_reg_3__3_ ( .D(int_data_y_7__7__3_), .CK(
        pe_1_6_7_net3247), .RN(pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_v[11]) );
  DFFR_X1 pe_1_6_7_int_q_reg_v_reg_4__0_ ( .D(int_data_y_7__7__0_), .CK(
        pe_1_6_7_net3252), .RN(pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_v[4]) );
  DFFR_X1 pe_1_6_7_int_q_reg_v_reg_4__1_ ( .D(int_data_y_7__7__1_), .CK(
        pe_1_6_7_net3252), .RN(pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_v[5]) );
  DFFR_X1 pe_1_6_7_int_q_reg_v_reg_4__2_ ( .D(int_data_y_7__7__2_), .CK(
        pe_1_6_7_net3252), .RN(pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_v[6]) );
  DFFR_X1 pe_1_6_7_int_q_reg_v_reg_4__3_ ( .D(int_data_y_7__7__3_), .CK(
        pe_1_6_7_net3252), .RN(pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_v[7]) );
  DFFR_X1 pe_1_6_7_int_q_reg_v_reg_5__0_ ( .D(int_data_y_7__7__0_), .CK(
        pe_1_6_7_net3257), .RN(pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_v[0]) );
  DFFR_X1 pe_1_6_7_int_q_reg_v_reg_5__1_ ( .D(int_data_y_7__7__1_), .CK(
        pe_1_6_7_net3257), .RN(pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_v[1]) );
  DFFR_X1 pe_1_6_7_int_q_reg_v_reg_5__2_ ( .D(int_data_y_7__7__2_), .CK(
        pe_1_6_7_net3257), .RN(pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_v[2]) );
  DFFR_X1 pe_1_6_7_int_q_reg_v_reg_5__3_ ( .D(int_data_y_7__7__3_), .CK(
        pe_1_6_7_net3257), .RN(pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_6_7_int_q_reg_h_reg_0__0_ ( .D(i_data_conv_h[4]), .SI(
        int_data_y_7__7__0_), .SE(pe_1_6_7_n65), .CK(pe_1_6_7_net3201), .RN(
        pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_6_7_int_q_reg_h_reg_0__1_ ( .D(i_data_conv_h[5]), .SI(
        int_data_y_7__7__1_), .SE(pe_1_6_7_n65), .CK(pe_1_6_7_net3201), .RN(
        pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_6_7_int_q_reg_h_reg_0__2_ ( .D(i_data_conv_h[6]), .SI(
        int_data_y_7__7__2_), .SE(pe_1_6_7_n65), .CK(pe_1_6_7_net3201), .RN(
        pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_6_7_int_q_reg_h_reg_0__3_ ( .D(i_data_conv_h[7]), .SI(
        int_data_y_7__7__3_), .SE(pe_1_6_7_n65), .CK(pe_1_6_7_net3201), .RN(
        pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_6_7_int_q_reg_h_reg_1__0_ ( .D(i_data_conv_h[4]), .SI(
        int_data_y_7__7__0_), .SE(pe_1_6_7_n65), .CK(pe_1_6_7_net3207), .RN(
        pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_6_7_int_q_reg_h_reg_1__1_ ( .D(i_data_conv_h[5]), .SI(
        int_data_y_7__7__1_), .SE(pe_1_6_7_n65), .CK(pe_1_6_7_net3207), .RN(
        pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_6_7_int_q_reg_h_reg_1__2_ ( .D(i_data_conv_h[6]), .SI(
        int_data_y_7__7__2_), .SE(pe_1_6_7_n65), .CK(pe_1_6_7_net3207), .RN(
        pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_6_7_int_q_reg_h_reg_1__3_ ( .D(i_data_conv_h[7]), .SI(
        int_data_y_7__7__3_), .SE(pe_1_6_7_n65), .CK(pe_1_6_7_net3207), .RN(
        pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_6_7_int_q_reg_h_reg_2__0_ ( .D(i_data_conv_h[4]), .SI(
        int_data_y_7__7__0_), .SE(pe_1_6_7_n65), .CK(pe_1_6_7_net3212), .RN(
        pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_6_7_int_q_reg_h_reg_2__1_ ( .D(i_data_conv_h[5]), .SI(
        int_data_y_7__7__1_), .SE(pe_1_6_7_n65), .CK(pe_1_6_7_net3212), .RN(
        pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_6_7_int_q_reg_h_reg_2__2_ ( .D(i_data_conv_h[6]), .SI(
        int_data_y_7__7__2_), .SE(pe_1_6_7_n65), .CK(pe_1_6_7_net3212), .RN(
        pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_6_7_int_q_reg_h_reg_2__3_ ( .D(i_data_conv_h[7]), .SI(
        int_data_y_7__7__3_), .SE(pe_1_6_7_n65), .CK(pe_1_6_7_net3212), .RN(
        pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_6_7_int_q_reg_h_reg_3__0_ ( .D(i_data_conv_h[4]), .SI(
        int_data_y_7__7__0_), .SE(pe_1_6_7_n65), .CK(pe_1_6_7_net3217), .RN(
        pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_6_7_int_q_reg_h_reg_3__1_ ( .D(i_data_conv_h[5]), .SI(
        int_data_y_7__7__1_), .SE(pe_1_6_7_n65), .CK(pe_1_6_7_net3217), .RN(
        pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_6_7_int_q_reg_h_reg_3__2_ ( .D(i_data_conv_h[6]), .SI(
        int_data_y_7__7__2_), .SE(pe_1_6_7_n65), .CK(pe_1_6_7_net3217), .RN(
        pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_6_7_int_q_reg_h_reg_3__3_ ( .D(i_data_conv_h[7]), .SI(
        int_data_y_7__7__3_), .SE(pe_1_6_7_n65), .CK(pe_1_6_7_net3217), .RN(
        pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_6_7_int_q_reg_h_reg_4__0_ ( .D(i_data_conv_h[4]), .SI(
        int_data_y_7__7__0_), .SE(pe_1_6_7_n66), .CK(pe_1_6_7_net3222), .RN(
        pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_6_7_int_q_reg_h_reg_4__1_ ( .D(i_data_conv_h[5]), .SI(
        int_data_y_7__7__1_), .SE(pe_1_6_7_n66), .CK(pe_1_6_7_net3222), .RN(
        pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_6_7_int_q_reg_h_reg_4__2_ ( .D(i_data_conv_h[6]), .SI(
        int_data_y_7__7__2_), .SE(pe_1_6_7_n66), .CK(pe_1_6_7_net3222), .RN(
        pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_6_7_int_q_reg_h_reg_4__3_ ( .D(i_data_conv_h[7]), .SI(
        int_data_y_7__7__3_), .SE(pe_1_6_7_n66), .CK(pe_1_6_7_net3222), .RN(
        pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_6_7_int_q_reg_h_reg_5__0_ ( .D(i_data_conv_h[4]), .SI(
        int_data_y_7__7__0_), .SE(pe_1_6_7_n66), .CK(pe_1_6_7_net3227), .RN(
        pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_6_7_int_q_reg_h_reg_5__1_ ( .D(i_data_conv_h[5]), .SI(
        int_data_y_7__7__1_), .SE(pe_1_6_7_n66), .CK(pe_1_6_7_net3227), .RN(
        pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_6_7_int_q_reg_h_reg_5__2_ ( .D(i_data_conv_h[6]), .SI(
        int_data_y_7__7__2_), .SE(pe_1_6_7_n66), .CK(pe_1_6_7_net3227), .RN(
        pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_6_7_int_q_reg_h_reg_5__3_ ( .D(i_data_conv_h[7]), .SI(
        int_data_y_7__7__3_), .SE(pe_1_6_7_n66), .CK(pe_1_6_7_net3227), .RN(
        pe_1_6_7_n72), .Q(pe_1_6_7_int_q_reg_h[3]) );
  FA_X1 pe_1_6_7_sub_81_U2_7 ( .A(int_data_res_6__7__7_), .B(pe_1_6_7_n76), 
        .CI(pe_1_6_7_sub_81_carry[7]), .S(pe_1_6_7_N77) );
  FA_X1 pe_1_6_7_sub_81_U2_6 ( .A(int_data_res_6__7__6_), .B(pe_1_6_7_n76), 
        .CI(pe_1_6_7_sub_81_carry[6]), .CO(pe_1_6_7_sub_81_carry[7]), .S(
        pe_1_6_7_N76) );
  FA_X1 pe_1_6_7_sub_81_U2_5 ( .A(int_data_res_6__7__5_), .B(pe_1_6_7_n76), 
        .CI(pe_1_6_7_sub_81_carry[5]), .CO(pe_1_6_7_sub_81_carry[6]), .S(
        pe_1_6_7_N75) );
  FA_X1 pe_1_6_7_sub_81_U2_4 ( .A(int_data_res_6__7__4_), .B(pe_1_6_7_n76), 
        .CI(pe_1_6_7_sub_81_carry[4]), .CO(pe_1_6_7_sub_81_carry[5]), .S(
        pe_1_6_7_N74) );
  FA_X1 pe_1_6_7_sub_81_U2_3 ( .A(int_data_res_6__7__3_), .B(pe_1_6_7_n76), 
        .CI(pe_1_6_7_sub_81_carry[3]), .CO(pe_1_6_7_sub_81_carry[4]), .S(
        pe_1_6_7_N73) );
  FA_X1 pe_1_6_7_sub_81_U2_2 ( .A(int_data_res_6__7__2_), .B(pe_1_6_7_n75), 
        .CI(pe_1_6_7_sub_81_carry[2]), .CO(pe_1_6_7_sub_81_carry[3]), .S(
        pe_1_6_7_N72) );
  FA_X1 pe_1_6_7_sub_81_U2_1 ( .A(int_data_res_6__7__1_), .B(pe_1_6_7_n74), 
        .CI(pe_1_6_7_sub_81_carry[1]), .CO(pe_1_6_7_sub_81_carry[2]), .S(
        pe_1_6_7_N71) );
  FA_X1 pe_1_6_7_add_83_U1_7 ( .A(int_data_res_6__7__7_), .B(
        pe_1_6_7_int_data_3_), .CI(pe_1_6_7_add_83_carry[7]), .S(pe_1_6_7_N85)
         );
  FA_X1 pe_1_6_7_add_83_U1_6 ( .A(int_data_res_6__7__6_), .B(
        pe_1_6_7_int_data_3_), .CI(pe_1_6_7_add_83_carry[6]), .CO(
        pe_1_6_7_add_83_carry[7]), .S(pe_1_6_7_N84) );
  FA_X1 pe_1_6_7_add_83_U1_5 ( .A(int_data_res_6__7__5_), .B(
        pe_1_6_7_int_data_3_), .CI(pe_1_6_7_add_83_carry[5]), .CO(
        pe_1_6_7_add_83_carry[6]), .S(pe_1_6_7_N83) );
  FA_X1 pe_1_6_7_add_83_U1_4 ( .A(int_data_res_6__7__4_), .B(
        pe_1_6_7_int_data_3_), .CI(pe_1_6_7_add_83_carry[4]), .CO(
        pe_1_6_7_add_83_carry[5]), .S(pe_1_6_7_N82) );
  FA_X1 pe_1_6_7_add_83_U1_3 ( .A(int_data_res_6__7__3_), .B(
        pe_1_6_7_int_data_3_), .CI(pe_1_6_7_add_83_carry[3]), .CO(
        pe_1_6_7_add_83_carry[4]), .S(pe_1_6_7_N81) );
  FA_X1 pe_1_6_7_add_83_U1_2 ( .A(int_data_res_6__7__2_), .B(
        pe_1_6_7_int_data_2_), .CI(pe_1_6_7_add_83_carry[2]), .CO(
        pe_1_6_7_add_83_carry[3]), .S(pe_1_6_7_N80) );
  FA_X1 pe_1_6_7_add_83_U1_1 ( .A(int_data_res_6__7__1_), .B(
        pe_1_6_7_int_data_1_), .CI(pe_1_6_7_n2), .CO(pe_1_6_7_add_83_carry[2]), 
        .S(pe_1_6_7_N79) );
  NAND3_X1 pe_1_6_7_U56 ( .A1(pe_1_6_7_n60), .A2(pe_1_6_7_n43), .A3(
        pe_1_6_7_n62), .ZN(pe_1_6_7_n40) );
  NAND3_X1 pe_1_6_7_U55 ( .A1(pe_1_6_7_n43), .A2(pe_1_6_7_n61), .A3(
        pe_1_6_7_n62), .ZN(pe_1_6_7_n39) );
  NAND3_X1 pe_1_6_7_U54 ( .A1(pe_1_6_7_n43), .A2(pe_1_6_7_n63), .A3(
        pe_1_6_7_n60), .ZN(pe_1_6_7_n38) );
  NAND3_X1 pe_1_6_7_U53 ( .A1(pe_1_6_7_n61), .A2(pe_1_6_7_n63), .A3(
        pe_1_6_7_n43), .ZN(pe_1_6_7_n37) );
  DFFR_X1 pe_1_6_7_int_q_acc_reg_6_ ( .D(pe_1_6_7_n78), .CK(pe_1_6_7_net3262), 
        .RN(pe_1_6_7_n71), .Q(int_data_res_6__7__6_) );
  DFFR_X1 pe_1_6_7_int_q_acc_reg_5_ ( .D(pe_1_6_7_n79), .CK(pe_1_6_7_net3262), 
        .RN(pe_1_6_7_n71), .Q(int_data_res_6__7__5_) );
  DFFR_X1 pe_1_6_7_int_q_acc_reg_4_ ( .D(pe_1_6_7_n80), .CK(pe_1_6_7_net3262), 
        .RN(pe_1_6_7_n71), .Q(int_data_res_6__7__4_) );
  DFFR_X1 pe_1_6_7_int_q_acc_reg_3_ ( .D(pe_1_6_7_n81), .CK(pe_1_6_7_net3262), 
        .RN(pe_1_6_7_n71), .Q(int_data_res_6__7__3_) );
  DFFR_X1 pe_1_6_7_int_q_acc_reg_2_ ( .D(pe_1_6_7_n82), .CK(pe_1_6_7_net3262), 
        .RN(pe_1_6_7_n71), .Q(int_data_res_6__7__2_) );
  DFFR_X1 pe_1_6_7_int_q_acc_reg_1_ ( .D(pe_1_6_7_n83), .CK(pe_1_6_7_net3262), 
        .RN(pe_1_6_7_n71), .Q(int_data_res_6__7__1_) );
  DFFR_X1 pe_1_6_7_int_q_acc_reg_7_ ( .D(pe_1_6_7_n77), .CK(pe_1_6_7_net3262), 
        .RN(pe_1_6_7_n71), .Q(int_data_res_6__7__7_) );
  CLKGATETST_X1 pe_1_6_7_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_6_7_n88), .SE(1'b0), .GCK(pe_1_6_7_net3201) );
  CLKGATETST_X1 pe_1_6_7_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_6_7_n87), .SE(1'b0), .GCK(pe_1_6_7_net3207) );
  CLKGATETST_X1 pe_1_6_7_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_6_7_n86), .SE(1'b0), .GCK(pe_1_6_7_net3212) );
  CLKGATETST_X1 pe_1_6_7_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_6_7_n85), .SE(1'b0), .GCK(pe_1_6_7_net3217) );
  CLKGATETST_X1 pe_1_6_7_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_6_7_n90), .SE(1'b0), .GCK(pe_1_6_7_net3222) );
  CLKGATETST_X1 pe_1_6_7_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_6_7_n89), .SE(1'b0), .GCK(pe_1_6_7_net3227) );
  CLKGATETST_X1 pe_1_6_7_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_6_7_N64), .SE(1'b0), .GCK(pe_1_6_7_net3232) );
  CLKGATETST_X1 pe_1_6_7_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_6_7_N63), .SE(1'b0), .GCK(pe_1_6_7_net3237) );
  CLKGATETST_X1 pe_1_6_7_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_6_7_N62), .SE(1'b0), .GCK(pe_1_6_7_net3242) );
  CLKGATETST_X1 pe_1_6_7_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_6_7_N61), .SE(1'b0), .GCK(pe_1_6_7_net3247) );
  CLKGATETST_X1 pe_1_6_7_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_6_7_N60), .SE(1'b0), .GCK(pe_1_6_7_net3252) );
  CLKGATETST_X1 pe_1_6_7_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_6_7_N59), .SE(1'b0), .GCK(pe_1_6_7_net3257) );
  CLKGATETST_X1 pe_1_6_7_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_6_7_N90), .SE(1'b0), .GCK(pe_1_6_7_net3262) );
  CLKBUF_X1 pe_1_7_0_U112 ( .A(pe_1_7_0_n72), .Z(pe_1_7_0_n71) );
  INV_X1 pe_1_7_0_U111 ( .A(n77), .ZN(pe_1_7_0_n70) );
  INV_X1 pe_1_7_0_U110 ( .A(n69), .ZN(pe_1_7_0_n69) );
  INV_X1 pe_1_7_0_U109 ( .A(n69), .ZN(pe_1_7_0_n68) );
  INV_X1 pe_1_7_0_U108 ( .A(n69), .ZN(pe_1_7_0_n67) );
  INV_X1 pe_1_7_0_U107 ( .A(pe_1_7_0_n69), .ZN(pe_1_7_0_n66) );
  INV_X1 pe_1_7_0_U106 ( .A(pe_1_7_0_n63), .ZN(pe_1_7_0_n62) );
  INV_X1 pe_1_7_0_U105 ( .A(pe_1_7_0_n61), .ZN(pe_1_7_0_n60) );
  INV_X1 pe_1_7_0_U104 ( .A(n29), .ZN(pe_1_7_0_n59) );
  INV_X1 pe_1_7_0_U103 ( .A(pe_1_7_0_n59), .ZN(pe_1_7_0_n58) );
  INV_X1 pe_1_7_0_U102 ( .A(n21), .ZN(pe_1_7_0_n57) );
  MUX2_X1 pe_1_7_0_U101 ( .A(pe_1_7_0_n54), .B(pe_1_7_0_n51), .S(n54), .Z(
        pe_1_7_0_o_data_h_3_) );
  MUX2_X1 pe_1_7_0_U100 ( .A(pe_1_7_0_n53), .B(pe_1_7_0_n52), .S(pe_1_7_0_n62), 
        .Z(pe_1_7_0_n54) );
  MUX2_X1 pe_1_7_0_U99 ( .A(pe_1_7_0_int_q_reg_h[23]), .B(
        pe_1_7_0_int_q_reg_h[19]), .S(pe_1_7_0_n56), .Z(pe_1_7_0_n53) );
  MUX2_X1 pe_1_7_0_U98 ( .A(pe_1_7_0_int_q_reg_h[15]), .B(
        pe_1_7_0_int_q_reg_h[11]), .S(pe_1_7_0_n56), .Z(pe_1_7_0_n52) );
  MUX2_X1 pe_1_7_0_U97 ( .A(pe_1_7_0_int_q_reg_h[7]), .B(
        pe_1_7_0_int_q_reg_h[3]), .S(pe_1_7_0_n56), .Z(pe_1_7_0_n51) );
  MUX2_X1 pe_1_7_0_U96 ( .A(pe_1_7_0_n50), .B(pe_1_7_0_n47), .S(n54), .Z(
        pe_1_7_0_o_data_h_2_) );
  MUX2_X1 pe_1_7_0_U95 ( .A(pe_1_7_0_n49), .B(pe_1_7_0_n48), .S(pe_1_7_0_n62), 
        .Z(pe_1_7_0_n50) );
  MUX2_X1 pe_1_7_0_U94 ( .A(pe_1_7_0_int_q_reg_h[22]), .B(
        pe_1_7_0_int_q_reg_h[18]), .S(pe_1_7_0_n56), .Z(pe_1_7_0_n49) );
  MUX2_X1 pe_1_7_0_U93 ( .A(pe_1_7_0_int_q_reg_h[14]), .B(
        pe_1_7_0_int_q_reg_h[10]), .S(pe_1_7_0_n56), .Z(pe_1_7_0_n48) );
  MUX2_X1 pe_1_7_0_U92 ( .A(pe_1_7_0_int_q_reg_h[6]), .B(
        pe_1_7_0_int_q_reg_h[2]), .S(pe_1_7_0_n56), .Z(pe_1_7_0_n47) );
  MUX2_X1 pe_1_7_0_U91 ( .A(pe_1_7_0_n46), .B(pe_1_7_0_n24), .S(n54), .Z(
        pe_1_7_0_o_data_h_1_) );
  MUX2_X1 pe_1_7_0_U90 ( .A(pe_1_7_0_n45), .B(pe_1_7_0_n25), .S(pe_1_7_0_n62), 
        .Z(pe_1_7_0_n46) );
  MUX2_X1 pe_1_7_0_U89 ( .A(pe_1_7_0_int_q_reg_h[21]), .B(
        pe_1_7_0_int_q_reg_h[17]), .S(pe_1_7_0_n56), .Z(pe_1_7_0_n45) );
  MUX2_X1 pe_1_7_0_U88 ( .A(pe_1_7_0_int_q_reg_h[13]), .B(
        pe_1_7_0_int_q_reg_h[9]), .S(pe_1_7_0_n56), .Z(pe_1_7_0_n25) );
  MUX2_X1 pe_1_7_0_U87 ( .A(pe_1_7_0_int_q_reg_h[5]), .B(
        pe_1_7_0_int_q_reg_h[1]), .S(pe_1_7_0_n56), .Z(pe_1_7_0_n24) );
  MUX2_X1 pe_1_7_0_U86 ( .A(pe_1_7_0_n23), .B(pe_1_7_0_n20), .S(n54), .Z(
        pe_1_7_0_o_data_h_0_) );
  MUX2_X1 pe_1_7_0_U85 ( .A(pe_1_7_0_n22), .B(pe_1_7_0_n21), .S(pe_1_7_0_n62), 
        .Z(pe_1_7_0_n23) );
  MUX2_X1 pe_1_7_0_U84 ( .A(pe_1_7_0_int_q_reg_h[20]), .B(
        pe_1_7_0_int_q_reg_h[16]), .S(pe_1_7_0_n56), .Z(pe_1_7_0_n22) );
  MUX2_X1 pe_1_7_0_U83 ( .A(pe_1_7_0_int_q_reg_h[12]), .B(
        pe_1_7_0_int_q_reg_h[8]), .S(pe_1_7_0_n56), .Z(pe_1_7_0_n21) );
  MUX2_X1 pe_1_7_0_U82 ( .A(pe_1_7_0_int_q_reg_h[4]), .B(
        pe_1_7_0_int_q_reg_h[0]), .S(pe_1_7_0_n56), .Z(pe_1_7_0_n20) );
  MUX2_X1 pe_1_7_0_U81 ( .A(pe_1_7_0_n19), .B(pe_1_7_0_n16), .S(n54), .Z(
        int_data_y_7__0__3_) );
  MUX2_X1 pe_1_7_0_U80 ( .A(pe_1_7_0_n18), .B(pe_1_7_0_n17), .S(pe_1_7_0_n62), 
        .Z(pe_1_7_0_n19) );
  MUX2_X1 pe_1_7_0_U79 ( .A(pe_1_7_0_int_q_reg_v[23]), .B(
        pe_1_7_0_int_q_reg_v[19]), .S(pe_1_7_0_n55), .Z(pe_1_7_0_n18) );
  MUX2_X1 pe_1_7_0_U78 ( .A(pe_1_7_0_int_q_reg_v[15]), .B(
        pe_1_7_0_int_q_reg_v[11]), .S(pe_1_7_0_n55), .Z(pe_1_7_0_n17) );
  MUX2_X1 pe_1_7_0_U77 ( .A(pe_1_7_0_int_q_reg_v[7]), .B(
        pe_1_7_0_int_q_reg_v[3]), .S(pe_1_7_0_n55), .Z(pe_1_7_0_n16) );
  MUX2_X1 pe_1_7_0_U76 ( .A(pe_1_7_0_n15), .B(pe_1_7_0_n12), .S(n54), .Z(
        int_data_y_7__0__2_) );
  MUX2_X1 pe_1_7_0_U75 ( .A(pe_1_7_0_n14), .B(pe_1_7_0_n13), .S(pe_1_7_0_n62), 
        .Z(pe_1_7_0_n15) );
  MUX2_X1 pe_1_7_0_U74 ( .A(pe_1_7_0_int_q_reg_v[22]), .B(
        pe_1_7_0_int_q_reg_v[18]), .S(pe_1_7_0_n55), .Z(pe_1_7_0_n14) );
  MUX2_X1 pe_1_7_0_U73 ( .A(pe_1_7_0_int_q_reg_v[14]), .B(
        pe_1_7_0_int_q_reg_v[10]), .S(pe_1_7_0_n55), .Z(pe_1_7_0_n13) );
  MUX2_X1 pe_1_7_0_U72 ( .A(pe_1_7_0_int_q_reg_v[6]), .B(
        pe_1_7_0_int_q_reg_v[2]), .S(pe_1_7_0_n55), .Z(pe_1_7_0_n12) );
  MUX2_X1 pe_1_7_0_U71 ( .A(pe_1_7_0_n11), .B(pe_1_7_0_n8), .S(n54), .Z(
        int_data_y_7__0__1_) );
  MUX2_X1 pe_1_7_0_U70 ( .A(pe_1_7_0_n10), .B(pe_1_7_0_n9), .S(pe_1_7_0_n62), 
        .Z(pe_1_7_0_n11) );
  MUX2_X1 pe_1_7_0_U69 ( .A(pe_1_7_0_int_q_reg_v[21]), .B(
        pe_1_7_0_int_q_reg_v[17]), .S(pe_1_7_0_n55), .Z(pe_1_7_0_n10) );
  MUX2_X1 pe_1_7_0_U68 ( .A(pe_1_7_0_int_q_reg_v[13]), .B(
        pe_1_7_0_int_q_reg_v[9]), .S(pe_1_7_0_n55), .Z(pe_1_7_0_n9) );
  MUX2_X1 pe_1_7_0_U67 ( .A(pe_1_7_0_int_q_reg_v[5]), .B(
        pe_1_7_0_int_q_reg_v[1]), .S(pe_1_7_0_n55), .Z(pe_1_7_0_n8) );
  MUX2_X1 pe_1_7_0_U66 ( .A(pe_1_7_0_n7), .B(pe_1_7_0_n4), .S(n54), .Z(
        int_data_y_7__0__0_) );
  MUX2_X1 pe_1_7_0_U65 ( .A(pe_1_7_0_n6), .B(pe_1_7_0_n5), .S(pe_1_7_0_n62), 
        .Z(pe_1_7_0_n7) );
  MUX2_X1 pe_1_7_0_U64 ( .A(pe_1_7_0_int_q_reg_v[20]), .B(
        pe_1_7_0_int_q_reg_v[16]), .S(pe_1_7_0_n55), .Z(pe_1_7_0_n6) );
  MUX2_X1 pe_1_7_0_U63 ( .A(pe_1_7_0_int_q_reg_v[12]), .B(
        pe_1_7_0_int_q_reg_v[8]), .S(pe_1_7_0_n55), .Z(pe_1_7_0_n5) );
  MUX2_X1 pe_1_7_0_U62 ( .A(pe_1_7_0_int_q_reg_v[4]), .B(
        pe_1_7_0_int_q_reg_v[0]), .S(pe_1_7_0_n55), .Z(pe_1_7_0_n4) );
  AND2_X1 pe_1_7_0_U61 ( .A1(pe_1_7_0_o_data_h_3_), .A2(pe_1_7_0_n58), .ZN(
        pe_1_7_0_int_data_3_) );
  NAND2_X1 pe_1_7_0_U60 ( .A1(pe_1_7_0_int_data_0_), .A2(pe_1_7_0_n3), .ZN(
        pe_1_7_0_sub_81_carry[1]) );
  INV_X1 pe_1_7_0_U59 ( .A(pe_1_7_0_int_data_1_), .ZN(pe_1_7_0_n74) );
  AOI222_X1 pe_1_7_0_U58 ( .A1(pe_1_7_0_n64), .A2(i_data_acc[63]), .B1(
        pe_1_7_0_N85), .B2(pe_1_7_0_n27), .C1(pe_1_7_0_N77), .C2(pe_1_7_0_n28), 
        .ZN(pe_1_7_0_n26) );
  INV_X1 pe_1_7_0_U57 ( .A(pe_1_7_0_n26), .ZN(pe_1_7_0_n77) );
  AOI222_X1 pe_1_7_0_U52 ( .A1(i_data_acc[57]), .A2(pe_1_7_0_n64), .B1(
        pe_1_7_0_N79), .B2(pe_1_7_0_n27), .C1(pe_1_7_0_N71), .C2(pe_1_7_0_n28), 
        .ZN(pe_1_7_0_n34) );
  INV_X1 pe_1_7_0_U51 ( .A(pe_1_7_0_n34), .ZN(pe_1_7_0_n83) );
  AOI222_X1 pe_1_7_0_U50 ( .A1(i_data_acc[58]), .A2(pe_1_7_0_n64), .B1(
        pe_1_7_0_N80), .B2(pe_1_7_0_n27), .C1(pe_1_7_0_N72), .C2(pe_1_7_0_n28), 
        .ZN(pe_1_7_0_n33) );
  INV_X1 pe_1_7_0_U49 ( .A(pe_1_7_0_n33), .ZN(pe_1_7_0_n82) );
  AOI222_X1 pe_1_7_0_U48 ( .A1(i_data_acc[62]), .A2(pe_1_7_0_n64), .B1(
        pe_1_7_0_N84), .B2(pe_1_7_0_n27), .C1(pe_1_7_0_N76), .C2(pe_1_7_0_n28), 
        .ZN(pe_1_7_0_n29) );
  INV_X1 pe_1_7_0_U47 ( .A(pe_1_7_0_n29), .ZN(pe_1_7_0_n78) );
  AND2_X1 pe_1_7_0_U46 ( .A1(pe_1_7_0_o_data_h_2_), .A2(pe_1_7_0_n58), .ZN(
        pe_1_7_0_int_data_2_) );
  AND2_X1 pe_1_7_0_U45 ( .A1(pe_1_7_0_o_data_h_1_), .A2(pe_1_7_0_n58), .ZN(
        pe_1_7_0_int_data_1_) );
  INV_X1 pe_1_7_0_U44 ( .A(pe_1_7_0_int_data_2_), .ZN(pe_1_7_0_n75) );
  AND2_X1 pe_1_7_0_U43 ( .A1(pe_1_7_0_int_data_0_), .A2(int_data_res_7__0__0_), 
        .ZN(pe_1_7_0_n2) );
  AND2_X1 pe_1_7_0_U42 ( .A1(pe_1_7_0_o_data_h_0_), .A2(pe_1_7_0_n58), .ZN(
        pe_1_7_0_int_data_0_) );
  XNOR2_X1 pe_1_7_0_U41 ( .A(pe_1_7_0_n73), .B(int_data_res_7__0__0_), .ZN(
        pe_1_7_0_N70) );
  AOI222_X1 pe_1_7_0_U40 ( .A1(i_data_acc[56]), .A2(pe_1_7_0_n64), .B1(
        pe_1_7_0_n1), .B2(pe_1_7_0_n27), .C1(pe_1_7_0_N70), .C2(pe_1_7_0_n28), 
        .ZN(pe_1_7_0_n35) );
  INV_X1 pe_1_7_0_U39 ( .A(pe_1_7_0_n35), .ZN(pe_1_7_0_n84) );
  AOI222_X1 pe_1_7_0_U38 ( .A1(i_data_acc[59]), .A2(pe_1_7_0_n64), .B1(
        pe_1_7_0_N81), .B2(pe_1_7_0_n27), .C1(pe_1_7_0_N73), .C2(pe_1_7_0_n28), 
        .ZN(pe_1_7_0_n32) );
  INV_X1 pe_1_7_0_U37 ( .A(pe_1_7_0_n32), .ZN(pe_1_7_0_n81) );
  AOI222_X1 pe_1_7_0_U36 ( .A1(i_data_acc[60]), .A2(pe_1_7_0_n64), .B1(
        pe_1_7_0_N82), .B2(pe_1_7_0_n27), .C1(pe_1_7_0_N74), .C2(pe_1_7_0_n28), 
        .ZN(pe_1_7_0_n31) );
  INV_X1 pe_1_7_0_U35 ( .A(pe_1_7_0_n31), .ZN(pe_1_7_0_n80) );
  AOI222_X1 pe_1_7_0_U34 ( .A1(i_data_acc[61]), .A2(pe_1_7_0_n64), .B1(
        pe_1_7_0_N83), .B2(pe_1_7_0_n27), .C1(pe_1_7_0_N75), .C2(pe_1_7_0_n28), 
        .ZN(pe_1_7_0_n30) );
  INV_X1 pe_1_7_0_U33 ( .A(pe_1_7_0_n30), .ZN(pe_1_7_0_n79) );
  NOR3_X1 pe_1_7_0_U32 ( .A1(pe_1_7_0_n59), .A2(pe_1_7_0_n65), .A3(int_ckg[7]), 
        .ZN(pe_1_7_0_n36) );
  OR2_X1 pe_1_7_0_U31 ( .A1(pe_1_7_0_n36), .A2(pe_1_7_0_n64), .ZN(pe_1_7_0_N90) );
  INV_X1 pe_1_7_0_U30 ( .A(pe_1_7_0_int_data_0_), .ZN(pe_1_7_0_n73) );
  INV_X1 pe_1_7_0_U29 ( .A(n41), .ZN(pe_1_7_0_n63) );
  INV_X1 pe_1_7_0_U28 ( .A(n35), .ZN(pe_1_7_0_n61) );
  INV_X1 pe_1_7_0_U27 ( .A(pe_1_7_0_int_data_3_), .ZN(pe_1_7_0_n76) );
  BUF_X1 pe_1_7_0_U26 ( .A(n63), .Z(pe_1_7_0_n64) );
  NAND2_X1 pe_1_7_0_U25 ( .A1(pe_1_7_0_n44), .A2(pe_1_7_0_n61), .ZN(
        pe_1_7_0_n41) );
  AND3_X1 pe_1_7_0_U24 ( .A1(n77), .A2(pe_1_7_0_n63), .A3(n54), .ZN(
        pe_1_7_0_n44) );
  NOR2_X1 pe_1_7_0_U23 ( .A1(pe_1_7_0_n70), .A2(n54), .ZN(pe_1_7_0_n43) );
  NOR2_X1 pe_1_7_0_U22 ( .A1(pe_1_7_0_n57), .A2(pe_1_7_0_n64), .ZN(
        pe_1_7_0_n28) );
  NOR2_X1 pe_1_7_0_U21 ( .A1(n21), .A2(pe_1_7_0_n64), .ZN(pe_1_7_0_n27) );
  INV_X1 pe_1_7_0_U20 ( .A(pe_1_7_0_n41), .ZN(pe_1_7_0_n90) );
  INV_X1 pe_1_7_0_U19 ( .A(pe_1_7_0_n37), .ZN(pe_1_7_0_n88) );
  INV_X1 pe_1_7_0_U18 ( .A(pe_1_7_0_n38), .ZN(pe_1_7_0_n87) );
  INV_X1 pe_1_7_0_U17 ( .A(pe_1_7_0_n39), .ZN(pe_1_7_0_n86) );
  NOR2_X1 pe_1_7_0_U16 ( .A1(pe_1_7_0_n68), .A2(pe_1_7_0_n42), .ZN(
        pe_1_7_0_N59) );
  NOR2_X1 pe_1_7_0_U15 ( .A1(pe_1_7_0_n68), .A2(pe_1_7_0_n41), .ZN(
        pe_1_7_0_N60) );
  NOR2_X1 pe_1_7_0_U14 ( .A1(pe_1_7_0_n68), .A2(pe_1_7_0_n38), .ZN(
        pe_1_7_0_N63) );
  NOR2_X1 pe_1_7_0_U13 ( .A1(pe_1_7_0_n67), .A2(pe_1_7_0_n40), .ZN(
        pe_1_7_0_N61) );
  NOR2_X1 pe_1_7_0_U12 ( .A1(pe_1_7_0_n67), .A2(pe_1_7_0_n39), .ZN(
        pe_1_7_0_N62) );
  NOR2_X1 pe_1_7_0_U11 ( .A1(pe_1_7_0_n37), .A2(pe_1_7_0_n67), .ZN(
        pe_1_7_0_N64) );
  NAND2_X1 pe_1_7_0_U10 ( .A1(pe_1_7_0_n44), .A2(pe_1_7_0_n60), .ZN(
        pe_1_7_0_n42) );
  BUF_X1 pe_1_7_0_U9 ( .A(pe_1_7_0_n60), .Z(pe_1_7_0_n55) );
  BUF_X1 pe_1_7_0_U8 ( .A(pe_1_7_0_n60), .Z(pe_1_7_0_n56) );
  INV_X1 pe_1_7_0_U7 ( .A(pe_1_7_0_n69), .ZN(pe_1_7_0_n65) );
  INV_X1 pe_1_7_0_U6 ( .A(pe_1_7_0_n42), .ZN(pe_1_7_0_n89) );
  INV_X1 pe_1_7_0_U5 ( .A(pe_1_7_0_n40), .ZN(pe_1_7_0_n85) );
  INV_X2 pe_1_7_0_U4 ( .A(n85), .ZN(pe_1_7_0_n72) );
  XOR2_X1 pe_1_7_0_U3 ( .A(pe_1_7_0_int_data_0_), .B(int_data_res_7__0__0_), 
        .Z(pe_1_7_0_n1) );
  DFFR_X1 pe_1_7_0_int_q_acc_reg_0_ ( .D(pe_1_7_0_n84), .CK(pe_1_7_0_net3184), 
        .RN(pe_1_7_0_n72), .Q(int_data_res_7__0__0_), .QN(pe_1_7_0_n3) );
  DFFR_X1 pe_1_7_0_int_q_reg_v_reg_0__0_ ( .D(i_data_conv_v[28]), .CK(
        pe_1_7_0_net3154), .RN(pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_v[20]) );
  DFFR_X1 pe_1_7_0_int_q_reg_v_reg_0__1_ ( .D(i_data_conv_v[29]), .CK(
        pe_1_7_0_net3154), .RN(pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_v[21]) );
  DFFR_X1 pe_1_7_0_int_q_reg_v_reg_0__2_ ( .D(i_data_conv_v[30]), .CK(
        pe_1_7_0_net3154), .RN(pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_v[22]) );
  DFFR_X1 pe_1_7_0_int_q_reg_v_reg_0__3_ ( .D(i_data_conv_v[31]), .CK(
        pe_1_7_0_net3154), .RN(pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_v[23]) );
  DFFR_X1 pe_1_7_0_int_q_reg_v_reg_1__0_ ( .D(i_data_conv_v[28]), .CK(
        pe_1_7_0_net3159), .RN(pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_v[16]) );
  DFFR_X1 pe_1_7_0_int_q_reg_v_reg_1__1_ ( .D(i_data_conv_v[29]), .CK(
        pe_1_7_0_net3159), .RN(pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_v[17]) );
  DFFR_X1 pe_1_7_0_int_q_reg_v_reg_1__2_ ( .D(i_data_conv_v[30]), .CK(
        pe_1_7_0_net3159), .RN(pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_v[18]) );
  DFFR_X1 pe_1_7_0_int_q_reg_v_reg_1__3_ ( .D(i_data_conv_v[31]), .CK(
        pe_1_7_0_net3159), .RN(pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_v[19]) );
  DFFR_X1 pe_1_7_0_int_q_reg_v_reg_2__0_ ( .D(i_data_conv_v[28]), .CK(
        pe_1_7_0_net3164), .RN(pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_v[12]) );
  DFFR_X1 pe_1_7_0_int_q_reg_v_reg_2__1_ ( .D(i_data_conv_v[29]), .CK(
        pe_1_7_0_net3164), .RN(pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_v[13]) );
  DFFR_X1 pe_1_7_0_int_q_reg_v_reg_2__2_ ( .D(i_data_conv_v[30]), .CK(
        pe_1_7_0_net3164), .RN(pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_v[14]) );
  DFFR_X1 pe_1_7_0_int_q_reg_v_reg_2__3_ ( .D(i_data_conv_v[31]), .CK(
        pe_1_7_0_net3164), .RN(pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_v[15]) );
  DFFR_X1 pe_1_7_0_int_q_reg_v_reg_3__0_ ( .D(i_data_conv_v[28]), .CK(
        pe_1_7_0_net3169), .RN(pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_v[8]) );
  DFFR_X1 pe_1_7_0_int_q_reg_v_reg_3__1_ ( .D(i_data_conv_v[29]), .CK(
        pe_1_7_0_net3169), .RN(pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_v[9]) );
  DFFR_X1 pe_1_7_0_int_q_reg_v_reg_3__2_ ( .D(i_data_conv_v[30]), .CK(
        pe_1_7_0_net3169), .RN(pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_v[10]) );
  DFFR_X1 pe_1_7_0_int_q_reg_v_reg_3__3_ ( .D(i_data_conv_v[31]), .CK(
        pe_1_7_0_net3169), .RN(pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_v[11]) );
  DFFR_X1 pe_1_7_0_int_q_reg_v_reg_4__0_ ( .D(i_data_conv_v[28]), .CK(
        pe_1_7_0_net3174), .RN(pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_v[4]) );
  DFFR_X1 pe_1_7_0_int_q_reg_v_reg_4__1_ ( .D(i_data_conv_v[29]), .CK(
        pe_1_7_0_net3174), .RN(pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_v[5]) );
  DFFR_X1 pe_1_7_0_int_q_reg_v_reg_4__2_ ( .D(i_data_conv_v[30]), .CK(
        pe_1_7_0_net3174), .RN(pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_v[6]) );
  DFFR_X1 pe_1_7_0_int_q_reg_v_reg_4__3_ ( .D(i_data_conv_v[31]), .CK(
        pe_1_7_0_net3174), .RN(pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_v[7]) );
  DFFR_X1 pe_1_7_0_int_q_reg_v_reg_5__0_ ( .D(i_data_conv_v[28]), .CK(
        pe_1_7_0_net3179), .RN(pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_v[0]) );
  DFFR_X1 pe_1_7_0_int_q_reg_v_reg_5__1_ ( .D(i_data_conv_v[29]), .CK(
        pe_1_7_0_net3179), .RN(pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_v[1]) );
  DFFR_X1 pe_1_7_0_int_q_reg_v_reg_5__2_ ( .D(i_data_conv_v[30]), .CK(
        pe_1_7_0_net3179), .RN(pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_v[2]) );
  DFFR_X1 pe_1_7_0_int_q_reg_v_reg_5__3_ ( .D(i_data_conv_v[31]), .CK(
        pe_1_7_0_net3179), .RN(pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_7_0_int_q_reg_h_reg_0__0_ ( .D(int_data_x_7__1__0_), .SI(
        i_data_conv_v[28]), .SE(pe_1_7_0_n65), .CK(pe_1_7_0_net3123), .RN(
        pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_7_0_int_q_reg_h_reg_0__1_ ( .D(int_data_x_7__1__1_), .SI(
        i_data_conv_v[29]), .SE(pe_1_7_0_n65), .CK(pe_1_7_0_net3123), .RN(
        pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_7_0_int_q_reg_h_reg_0__2_ ( .D(int_data_x_7__1__2_), .SI(
        i_data_conv_v[30]), .SE(pe_1_7_0_n65), .CK(pe_1_7_0_net3123), .RN(
        pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_7_0_int_q_reg_h_reg_0__3_ ( .D(int_data_x_7__1__3_), .SI(
        i_data_conv_v[31]), .SE(pe_1_7_0_n65), .CK(pe_1_7_0_net3123), .RN(
        pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_7_0_int_q_reg_h_reg_1__0_ ( .D(int_data_x_7__1__0_), .SI(
        i_data_conv_v[28]), .SE(pe_1_7_0_n65), .CK(pe_1_7_0_net3129), .RN(
        pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_7_0_int_q_reg_h_reg_1__1_ ( .D(int_data_x_7__1__1_), .SI(
        i_data_conv_v[29]), .SE(pe_1_7_0_n65), .CK(pe_1_7_0_net3129), .RN(
        pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_7_0_int_q_reg_h_reg_1__2_ ( .D(int_data_x_7__1__2_), .SI(
        i_data_conv_v[30]), .SE(pe_1_7_0_n65), .CK(pe_1_7_0_net3129), .RN(
        pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_7_0_int_q_reg_h_reg_1__3_ ( .D(int_data_x_7__1__3_), .SI(
        i_data_conv_v[31]), .SE(pe_1_7_0_n65), .CK(pe_1_7_0_net3129), .RN(
        pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_7_0_int_q_reg_h_reg_2__0_ ( .D(int_data_x_7__1__0_), .SI(
        i_data_conv_v[28]), .SE(pe_1_7_0_n65), .CK(pe_1_7_0_net3134), .RN(
        pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_7_0_int_q_reg_h_reg_2__1_ ( .D(int_data_x_7__1__1_), .SI(
        i_data_conv_v[29]), .SE(pe_1_7_0_n65), .CK(pe_1_7_0_net3134), .RN(
        pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_7_0_int_q_reg_h_reg_2__2_ ( .D(int_data_x_7__1__2_), .SI(
        i_data_conv_v[30]), .SE(pe_1_7_0_n65), .CK(pe_1_7_0_net3134), .RN(
        pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_7_0_int_q_reg_h_reg_2__3_ ( .D(int_data_x_7__1__3_), .SI(
        i_data_conv_v[31]), .SE(pe_1_7_0_n65), .CK(pe_1_7_0_net3134), .RN(
        pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_7_0_int_q_reg_h_reg_3__0_ ( .D(int_data_x_7__1__0_), .SI(
        i_data_conv_v[28]), .SE(pe_1_7_0_n65), .CK(pe_1_7_0_net3139), .RN(
        pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_7_0_int_q_reg_h_reg_3__1_ ( .D(int_data_x_7__1__1_), .SI(
        i_data_conv_v[29]), .SE(pe_1_7_0_n65), .CK(pe_1_7_0_net3139), .RN(
        pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_7_0_int_q_reg_h_reg_3__2_ ( .D(int_data_x_7__1__2_), .SI(
        i_data_conv_v[30]), .SE(pe_1_7_0_n65), .CK(pe_1_7_0_net3139), .RN(
        pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_7_0_int_q_reg_h_reg_3__3_ ( .D(int_data_x_7__1__3_), .SI(
        i_data_conv_v[31]), .SE(pe_1_7_0_n65), .CK(pe_1_7_0_net3139), .RN(
        pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_7_0_int_q_reg_h_reg_4__0_ ( .D(int_data_x_7__1__0_), .SI(
        i_data_conv_v[28]), .SE(pe_1_7_0_n66), .CK(pe_1_7_0_net3144), .RN(
        pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_7_0_int_q_reg_h_reg_4__1_ ( .D(int_data_x_7__1__1_), .SI(
        i_data_conv_v[29]), .SE(pe_1_7_0_n66), .CK(pe_1_7_0_net3144), .RN(
        pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_7_0_int_q_reg_h_reg_4__2_ ( .D(int_data_x_7__1__2_), .SI(
        i_data_conv_v[30]), .SE(pe_1_7_0_n66), .CK(pe_1_7_0_net3144), .RN(
        pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_7_0_int_q_reg_h_reg_4__3_ ( .D(int_data_x_7__1__3_), .SI(
        i_data_conv_v[31]), .SE(pe_1_7_0_n66), .CK(pe_1_7_0_net3144), .RN(
        pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_7_0_int_q_reg_h_reg_5__0_ ( .D(int_data_x_7__1__0_), .SI(
        i_data_conv_v[28]), .SE(pe_1_7_0_n66), .CK(pe_1_7_0_net3149), .RN(
        pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_7_0_int_q_reg_h_reg_5__1_ ( .D(int_data_x_7__1__1_), .SI(
        i_data_conv_v[29]), .SE(pe_1_7_0_n66), .CK(pe_1_7_0_net3149), .RN(
        pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_7_0_int_q_reg_h_reg_5__2_ ( .D(int_data_x_7__1__2_), .SI(
        i_data_conv_v[30]), .SE(pe_1_7_0_n66), .CK(pe_1_7_0_net3149), .RN(
        pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_7_0_int_q_reg_h_reg_5__3_ ( .D(int_data_x_7__1__3_), .SI(
        i_data_conv_v[31]), .SE(pe_1_7_0_n66), .CK(pe_1_7_0_net3149), .RN(
        pe_1_7_0_n72), .Q(pe_1_7_0_int_q_reg_h[3]) );
  FA_X1 pe_1_7_0_sub_81_U2_7 ( .A(int_data_res_7__0__7_), .B(pe_1_7_0_n76), 
        .CI(pe_1_7_0_sub_81_carry[7]), .S(pe_1_7_0_N77) );
  FA_X1 pe_1_7_0_sub_81_U2_6 ( .A(int_data_res_7__0__6_), .B(pe_1_7_0_n76), 
        .CI(pe_1_7_0_sub_81_carry[6]), .CO(pe_1_7_0_sub_81_carry[7]), .S(
        pe_1_7_0_N76) );
  FA_X1 pe_1_7_0_sub_81_U2_5 ( .A(int_data_res_7__0__5_), .B(pe_1_7_0_n76), 
        .CI(pe_1_7_0_sub_81_carry[5]), .CO(pe_1_7_0_sub_81_carry[6]), .S(
        pe_1_7_0_N75) );
  FA_X1 pe_1_7_0_sub_81_U2_4 ( .A(int_data_res_7__0__4_), .B(pe_1_7_0_n76), 
        .CI(pe_1_7_0_sub_81_carry[4]), .CO(pe_1_7_0_sub_81_carry[5]), .S(
        pe_1_7_0_N74) );
  FA_X1 pe_1_7_0_sub_81_U2_3 ( .A(int_data_res_7__0__3_), .B(pe_1_7_0_n76), 
        .CI(pe_1_7_0_sub_81_carry[3]), .CO(pe_1_7_0_sub_81_carry[4]), .S(
        pe_1_7_0_N73) );
  FA_X1 pe_1_7_0_sub_81_U2_2 ( .A(int_data_res_7__0__2_), .B(pe_1_7_0_n75), 
        .CI(pe_1_7_0_sub_81_carry[2]), .CO(pe_1_7_0_sub_81_carry[3]), .S(
        pe_1_7_0_N72) );
  FA_X1 pe_1_7_0_sub_81_U2_1 ( .A(int_data_res_7__0__1_), .B(pe_1_7_0_n74), 
        .CI(pe_1_7_0_sub_81_carry[1]), .CO(pe_1_7_0_sub_81_carry[2]), .S(
        pe_1_7_0_N71) );
  FA_X1 pe_1_7_0_add_83_U1_7 ( .A(int_data_res_7__0__7_), .B(
        pe_1_7_0_int_data_3_), .CI(pe_1_7_0_add_83_carry[7]), .S(pe_1_7_0_N85)
         );
  FA_X1 pe_1_7_0_add_83_U1_6 ( .A(int_data_res_7__0__6_), .B(
        pe_1_7_0_int_data_3_), .CI(pe_1_7_0_add_83_carry[6]), .CO(
        pe_1_7_0_add_83_carry[7]), .S(pe_1_7_0_N84) );
  FA_X1 pe_1_7_0_add_83_U1_5 ( .A(int_data_res_7__0__5_), .B(
        pe_1_7_0_int_data_3_), .CI(pe_1_7_0_add_83_carry[5]), .CO(
        pe_1_7_0_add_83_carry[6]), .S(pe_1_7_0_N83) );
  FA_X1 pe_1_7_0_add_83_U1_4 ( .A(int_data_res_7__0__4_), .B(
        pe_1_7_0_int_data_3_), .CI(pe_1_7_0_add_83_carry[4]), .CO(
        pe_1_7_0_add_83_carry[5]), .S(pe_1_7_0_N82) );
  FA_X1 pe_1_7_0_add_83_U1_3 ( .A(int_data_res_7__0__3_), .B(
        pe_1_7_0_int_data_3_), .CI(pe_1_7_0_add_83_carry[3]), .CO(
        pe_1_7_0_add_83_carry[4]), .S(pe_1_7_0_N81) );
  FA_X1 pe_1_7_0_add_83_U1_2 ( .A(int_data_res_7__0__2_), .B(
        pe_1_7_0_int_data_2_), .CI(pe_1_7_0_add_83_carry[2]), .CO(
        pe_1_7_0_add_83_carry[3]), .S(pe_1_7_0_N80) );
  FA_X1 pe_1_7_0_add_83_U1_1 ( .A(int_data_res_7__0__1_), .B(
        pe_1_7_0_int_data_1_), .CI(pe_1_7_0_n2), .CO(pe_1_7_0_add_83_carry[2]), 
        .S(pe_1_7_0_N79) );
  NAND3_X1 pe_1_7_0_U56 ( .A1(pe_1_7_0_n60), .A2(pe_1_7_0_n43), .A3(
        pe_1_7_0_n62), .ZN(pe_1_7_0_n40) );
  NAND3_X1 pe_1_7_0_U55 ( .A1(pe_1_7_0_n43), .A2(pe_1_7_0_n61), .A3(
        pe_1_7_0_n62), .ZN(pe_1_7_0_n39) );
  NAND3_X1 pe_1_7_0_U54 ( .A1(pe_1_7_0_n43), .A2(pe_1_7_0_n63), .A3(
        pe_1_7_0_n60), .ZN(pe_1_7_0_n38) );
  NAND3_X1 pe_1_7_0_U53 ( .A1(pe_1_7_0_n61), .A2(pe_1_7_0_n63), .A3(
        pe_1_7_0_n43), .ZN(pe_1_7_0_n37) );
  DFFR_X1 pe_1_7_0_int_q_acc_reg_6_ ( .D(pe_1_7_0_n78), .CK(pe_1_7_0_net3184), 
        .RN(pe_1_7_0_n71), .Q(int_data_res_7__0__6_) );
  DFFR_X1 pe_1_7_0_int_q_acc_reg_5_ ( .D(pe_1_7_0_n79), .CK(pe_1_7_0_net3184), 
        .RN(pe_1_7_0_n71), .Q(int_data_res_7__0__5_) );
  DFFR_X1 pe_1_7_0_int_q_acc_reg_4_ ( .D(pe_1_7_0_n80), .CK(pe_1_7_0_net3184), 
        .RN(pe_1_7_0_n71), .Q(int_data_res_7__0__4_) );
  DFFR_X1 pe_1_7_0_int_q_acc_reg_3_ ( .D(pe_1_7_0_n81), .CK(pe_1_7_0_net3184), 
        .RN(pe_1_7_0_n71), .Q(int_data_res_7__0__3_) );
  DFFR_X1 pe_1_7_0_int_q_acc_reg_2_ ( .D(pe_1_7_0_n82), .CK(pe_1_7_0_net3184), 
        .RN(pe_1_7_0_n71), .Q(int_data_res_7__0__2_) );
  DFFR_X1 pe_1_7_0_int_q_acc_reg_1_ ( .D(pe_1_7_0_n83), .CK(pe_1_7_0_net3184), 
        .RN(pe_1_7_0_n71), .Q(int_data_res_7__0__1_) );
  DFFR_X1 pe_1_7_0_int_q_acc_reg_7_ ( .D(pe_1_7_0_n77), .CK(pe_1_7_0_net3184), 
        .RN(pe_1_7_0_n71), .Q(int_data_res_7__0__7_) );
  CLKGATETST_X1 pe_1_7_0_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_7_0_n88), .SE(1'b0), .GCK(pe_1_7_0_net3123) );
  CLKGATETST_X1 pe_1_7_0_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_7_0_n87), .SE(1'b0), .GCK(pe_1_7_0_net3129) );
  CLKGATETST_X1 pe_1_7_0_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_7_0_n86), .SE(1'b0), .GCK(pe_1_7_0_net3134) );
  CLKGATETST_X1 pe_1_7_0_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_7_0_n85), .SE(1'b0), .GCK(pe_1_7_0_net3139) );
  CLKGATETST_X1 pe_1_7_0_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_7_0_n90), .SE(1'b0), .GCK(pe_1_7_0_net3144) );
  CLKGATETST_X1 pe_1_7_0_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_7_0_n89), .SE(1'b0), .GCK(pe_1_7_0_net3149) );
  CLKGATETST_X1 pe_1_7_0_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_7_0_N64), .SE(1'b0), .GCK(pe_1_7_0_net3154) );
  CLKGATETST_X1 pe_1_7_0_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_7_0_N63), .SE(1'b0), .GCK(pe_1_7_0_net3159) );
  CLKGATETST_X1 pe_1_7_0_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_7_0_N62), .SE(1'b0), .GCK(pe_1_7_0_net3164) );
  CLKGATETST_X1 pe_1_7_0_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_7_0_N61), .SE(1'b0), .GCK(pe_1_7_0_net3169) );
  CLKGATETST_X1 pe_1_7_0_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_7_0_N60), .SE(1'b0), .GCK(pe_1_7_0_net3174) );
  CLKGATETST_X1 pe_1_7_0_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_7_0_N59), .SE(1'b0), .GCK(pe_1_7_0_net3179) );
  CLKGATETST_X1 pe_1_7_0_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_7_0_N90), .SE(1'b0), .GCK(pe_1_7_0_net3184) );
  CLKBUF_X1 pe_1_7_1_U112 ( .A(pe_1_7_1_n72), .Z(pe_1_7_1_n71) );
  INV_X1 pe_1_7_1_U111 ( .A(n77), .ZN(pe_1_7_1_n70) );
  INV_X1 pe_1_7_1_U110 ( .A(n69), .ZN(pe_1_7_1_n69) );
  INV_X1 pe_1_7_1_U109 ( .A(n69), .ZN(pe_1_7_1_n68) );
  INV_X1 pe_1_7_1_U108 ( .A(n69), .ZN(pe_1_7_1_n67) );
  INV_X1 pe_1_7_1_U107 ( .A(pe_1_7_1_n69), .ZN(pe_1_7_1_n66) );
  INV_X1 pe_1_7_1_U106 ( .A(pe_1_7_1_n63), .ZN(pe_1_7_1_n62) );
  INV_X1 pe_1_7_1_U105 ( .A(pe_1_7_1_n61), .ZN(pe_1_7_1_n60) );
  INV_X1 pe_1_7_1_U104 ( .A(n29), .ZN(pe_1_7_1_n59) );
  INV_X1 pe_1_7_1_U103 ( .A(pe_1_7_1_n59), .ZN(pe_1_7_1_n58) );
  INV_X1 pe_1_7_1_U102 ( .A(n21), .ZN(pe_1_7_1_n57) );
  MUX2_X1 pe_1_7_1_U101 ( .A(pe_1_7_1_n54), .B(pe_1_7_1_n51), .S(n54), .Z(
        int_data_x_7__1__3_) );
  MUX2_X1 pe_1_7_1_U100 ( .A(pe_1_7_1_n53), .B(pe_1_7_1_n52), .S(pe_1_7_1_n62), 
        .Z(pe_1_7_1_n54) );
  MUX2_X1 pe_1_7_1_U99 ( .A(pe_1_7_1_int_q_reg_h[23]), .B(
        pe_1_7_1_int_q_reg_h[19]), .S(pe_1_7_1_n56), .Z(pe_1_7_1_n53) );
  MUX2_X1 pe_1_7_1_U98 ( .A(pe_1_7_1_int_q_reg_h[15]), .B(
        pe_1_7_1_int_q_reg_h[11]), .S(pe_1_7_1_n56), .Z(pe_1_7_1_n52) );
  MUX2_X1 pe_1_7_1_U97 ( .A(pe_1_7_1_int_q_reg_h[7]), .B(
        pe_1_7_1_int_q_reg_h[3]), .S(pe_1_7_1_n56), .Z(pe_1_7_1_n51) );
  MUX2_X1 pe_1_7_1_U96 ( .A(pe_1_7_1_n50), .B(pe_1_7_1_n47), .S(n54), .Z(
        int_data_x_7__1__2_) );
  MUX2_X1 pe_1_7_1_U95 ( .A(pe_1_7_1_n49), .B(pe_1_7_1_n48), .S(pe_1_7_1_n62), 
        .Z(pe_1_7_1_n50) );
  MUX2_X1 pe_1_7_1_U94 ( .A(pe_1_7_1_int_q_reg_h[22]), .B(
        pe_1_7_1_int_q_reg_h[18]), .S(pe_1_7_1_n56), .Z(pe_1_7_1_n49) );
  MUX2_X1 pe_1_7_1_U93 ( .A(pe_1_7_1_int_q_reg_h[14]), .B(
        pe_1_7_1_int_q_reg_h[10]), .S(pe_1_7_1_n56), .Z(pe_1_7_1_n48) );
  MUX2_X1 pe_1_7_1_U92 ( .A(pe_1_7_1_int_q_reg_h[6]), .B(
        pe_1_7_1_int_q_reg_h[2]), .S(pe_1_7_1_n56), .Z(pe_1_7_1_n47) );
  MUX2_X1 pe_1_7_1_U91 ( .A(pe_1_7_1_n46), .B(pe_1_7_1_n24), .S(n54), .Z(
        int_data_x_7__1__1_) );
  MUX2_X1 pe_1_7_1_U90 ( .A(pe_1_7_1_n45), .B(pe_1_7_1_n25), .S(pe_1_7_1_n62), 
        .Z(pe_1_7_1_n46) );
  MUX2_X1 pe_1_7_1_U89 ( .A(pe_1_7_1_int_q_reg_h[21]), .B(
        pe_1_7_1_int_q_reg_h[17]), .S(pe_1_7_1_n56), .Z(pe_1_7_1_n45) );
  MUX2_X1 pe_1_7_1_U88 ( .A(pe_1_7_1_int_q_reg_h[13]), .B(
        pe_1_7_1_int_q_reg_h[9]), .S(pe_1_7_1_n56), .Z(pe_1_7_1_n25) );
  MUX2_X1 pe_1_7_1_U87 ( .A(pe_1_7_1_int_q_reg_h[5]), .B(
        pe_1_7_1_int_q_reg_h[1]), .S(pe_1_7_1_n56), .Z(pe_1_7_1_n24) );
  MUX2_X1 pe_1_7_1_U86 ( .A(pe_1_7_1_n23), .B(pe_1_7_1_n20), .S(n54), .Z(
        int_data_x_7__1__0_) );
  MUX2_X1 pe_1_7_1_U85 ( .A(pe_1_7_1_n22), .B(pe_1_7_1_n21), .S(pe_1_7_1_n62), 
        .Z(pe_1_7_1_n23) );
  MUX2_X1 pe_1_7_1_U84 ( .A(pe_1_7_1_int_q_reg_h[20]), .B(
        pe_1_7_1_int_q_reg_h[16]), .S(pe_1_7_1_n56), .Z(pe_1_7_1_n22) );
  MUX2_X1 pe_1_7_1_U83 ( .A(pe_1_7_1_int_q_reg_h[12]), .B(
        pe_1_7_1_int_q_reg_h[8]), .S(pe_1_7_1_n56), .Z(pe_1_7_1_n21) );
  MUX2_X1 pe_1_7_1_U82 ( .A(pe_1_7_1_int_q_reg_h[4]), .B(
        pe_1_7_1_int_q_reg_h[0]), .S(pe_1_7_1_n56), .Z(pe_1_7_1_n20) );
  MUX2_X1 pe_1_7_1_U81 ( .A(pe_1_7_1_n19), .B(pe_1_7_1_n16), .S(n54), .Z(
        int_data_y_7__1__3_) );
  MUX2_X1 pe_1_7_1_U80 ( .A(pe_1_7_1_n18), .B(pe_1_7_1_n17), .S(pe_1_7_1_n62), 
        .Z(pe_1_7_1_n19) );
  MUX2_X1 pe_1_7_1_U79 ( .A(pe_1_7_1_int_q_reg_v[23]), .B(
        pe_1_7_1_int_q_reg_v[19]), .S(pe_1_7_1_n55), .Z(pe_1_7_1_n18) );
  MUX2_X1 pe_1_7_1_U78 ( .A(pe_1_7_1_int_q_reg_v[15]), .B(
        pe_1_7_1_int_q_reg_v[11]), .S(pe_1_7_1_n55), .Z(pe_1_7_1_n17) );
  MUX2_X1 pe_1_7_1_U77 ( .A(pe_1_7_1_int_q_reg_v[7]), .B(
        pe_1_7_1_int_q_reg_v[3]), .S(pe_1_7_1_n55), .Z(pe_1_7_1_n16) );
  MUX2_X1 pe_1_7_1_U76 ( .A(pe_1_7_1_n15), .B(pe_1_7_1_n12), .S(n54), .Z(
        int_data_y_7__1__2_) );
  MUX2_X1 pe_1_7_1_U75 ( .A(pe_1_7_1_n14), .B(pe_1_7_1_n13), .S(pe_1_7_1_n62), 
        .Z(pe_1_7_1_n15) );
  MUX2_X1 pe_1_7_1_U74 ( .A(pe_1_7_1_int_q_reg_v[22]), .B(
        pe_1_7_1_int_q_reg_v[18]), .S(pe_1_7_1_n55), .Z(pe_1_7_1_n14) );
  MUX2_X1 pe_1_7_1_U73 ( .A(pe_1_7_1_int_q_reg_v[14]), .B(
        pe_1_7_1_int_q_reg_v[10]), .S(pe_1_7_1_n55), .Z(pe_1_7_1_n13) );
  MUX2_X1 pe_1_7_1_U72 ( .A(pe_1_7_1_int_q_reg_v[6]), .B(
        pe_1_7_1_int_q_reg_v[2]), .S(pe_1_7_1_n55), .Z(pe_1_7_1_n12) );
  MUX2_X1 pe_1_7_1_U71 ( .A(pe_1_7_1_n11), .B(pe_1_7_1_n8), .S(n54), .Z(
        int_data_y_7__1__1_) );
  MUX2_X1 pe_1_7_1_U70 ( .A(pe_1_7_1_n10), .B(pe_1_7_1_n9), .S(pe_1_7_1_n62), 
        .Z(pe_1_7_1_n11) );
  MUX2_X1 pe_1_7_1_U69 ( .A(pe_1_7_1_int_q_reg_v[21]), .B(
        pe_1_7_1_int_q_reg_v[17]), .S(pe_1_7_1_n55), .Z(pe_1_7_1_n10) );
  MUX2_X1 pe_1_7_1_U68 ( .A(pe_1_7_1_int_q_reg_v[13]), .B(
        pe_1_7_1_int_q_reg_v[9]), .S(pe_1_7_1_n55), .Z(pe_1_7_1_n9) );
  MUX2_X1 pe_1_7_1_U67 ( .A(pe_1_7_1_int_q_reg_v[5]), .B(
        pe_1_7_1_int_q_reg_v[1]), .S(pe_1_7_1_n55), .Z(pe_1_7_1_n8) );
  MUX2_X1 pe_1_7_1_U66 ( .A(pe_1_7_1_n7), .B(pe_1_7_1_n4), .S(n54), .Z(
        int_data_y_7__1__0_) );
  MUX2_X1 pe_1_7_1_U65 ( .A(pe_1_7_1_n6), .B(pe_1_7_1_n5), .S(pe_1_7_1_n62), 
        .Z(pe_1_7_1_n7) );
  MUX2_X1 pe_1_7_1_U64 ( .A(pe_1_7_1_int_q_reg_v[20]), .B(
        pe_1_7_1_int_q_reg_v[16]), .S(pe_1_7_1_n55), .Z(pe_1_7_1_n6) );
  MUX2_X1 pe_1_7_1_U63 ( .A(pe_1_7_1_int_q_reg_v[12]), .B(
        pe_1_7_1_int_q_reg_v[8]), .S(pe_1_7_1_n55), .Z(pe_1_7_1_n5) );
  MUX2_X1 pe_1_7_1_U62 ( .A(pe_1_7_1_int_q_reg_v[4]), .B(
        pe_1_7_1_int_q_reg_v[0]), .S(pe_1_7_1_n55), .Z(pe_1_7_1_n4) );
  AOI222_X1 pe_1_7_1_U61 ( .A1(i_data_acc[50]), .A2(pe_1_7_1_n64), .B1(
        pe_1_7_1_N80), .B2(pe_1_7_1_n27), .C1(pe_1_7_1_N72), .C2(pe_1_7_1_n28), 
        .ZN(pe_1_7_1_n33) );
  INV_X1 pe_1_7_1_U60 ( .A(pe_1_7_1_n33), .ZN(pe_1_7_1_n82) );
  AOI222_X1 pe_1_7_1_U59 ( .A1(i_data_acc[54]), .A2(pe_1_7_1_n64), .B1(
        pe_1_7_1_N84), .B2(pe_1_7_1_n27), .C1(pe_1_7_1_N76), .C2(pe_1_7_1_n28), 
        .ZN(pe_1_7_1_n29) );
  INV_X1 pe_1_7_1_U58 ( .A(pe_1_7_1_n29), .ZN(pe_1_7_1_n78) );
  XNOR2_X1 pe_1_7_1_U57 ( .A(pe_1_7_1_n73), .B(int_data_res_7__1__0_), .ZN(
        pe_1_7_1_N70) );
  AOI222_X1 pe_1_7_1_U52 ( .A1(i_data_acc[48]), .A2(pe_1_7_1_n64), .B1(
        pe_1_7_1_n1), .B2(pe_1_7_1_n27), .C1(pe_1_7_1_N70), .C2(pe_1_7_1_n28), 
        .ZN(pe_1_7_1_n35) );
  INV_X1 pe_1_7_1_U51 ( .A(pe_1_7_1_n35), .ZN(pe_1_7_1_n84) );
  AOI222_X1 pe_1_7_1_U50 ( .A1(i_data_acc[49]), .A2(pe_1_7_1_n64), .B1(
        pe_1_7_1_N79), .B2(pe_1_7_1_n27), .C1(pe_1_7_1_N71), .C2(pe_1_7_1_n28), 
        .ZN(pe_1_7_1_n34) );
  INV_X1 pe_1_7_1_U49 ( .A(pe_1_7_1_n34), .ZN(pe_1_7_1_n83) );
  AOI222_X1 pe_1_7_1_U48 ( .A1(i_data_acc[51]), .A2(pe_1_7_1_n64), .B1(
        pe_1_7_1_N81), .B2(pe_1_7_1_n27), .C1(pe_1_7_1_N73), .C2(pe_1_7_1_n28), 
        .ZN(pe_1_7_1_n32) );
  INV_X1 pe_1_7_1_U47 ( .A(pe_1_7_1_n32), .ZN(pe_1_7_1_n81) );
  AOI222_X1 pe_1_7_1_U46 ( .A1(i_data_acc[52]), .A2(pe_1_7_1_n64), .B1(
        pe_1_7_1_N82), .B2(pe_1_7_1_n27), .C1(pe_1_7_1_N74), .C2(pe_1_7_1_n28), 
        .ZN(pe_1_7_1_n31) );
  INV_X1 pe_1_7_1_U45 ( .A(pe_1_7_1_n31), .ZN(pe_1_7_1_n80) );
  AOI222_X1 pe_1_7_1_U44 ( .A1(i_data_acc[53]), .A2(pe_1_7_1_n64), .B1(
        pe_1_7_1_N83), .B2(pe_1_7_1_n27), .C1(pe_1_7_1_N75), .C2(pe_1_7_1_n28), 
        .ZN(pe_1_7_1_n30) );
  INV_X1 pe_1_7_1_U43 ( .A(pe_1_7_1_n30), .ZN(pe_1_7_1_n79) );
  NAND2_X1 pe_1_7_1_U42 ( .A1(pe_1_7_1_int_data_0_), .A2(pe_1_7_1_n3), .ZN(
        pe_1_7_1_sub_81_carry[1]) );
  INV_X1 pe_1_7_1_U41 ( .A(pe_1_7_1_int_data_1_), .ZN(pe_1_7_1_n74) );
  INV_X1 pe_1_7_1_U40 ( .A(pe_1_7_1_int_data_2_), .ZN(pe_1_7_1_n75) );
  AND2_X1 pe_1_7_1_U39 ( .A1(pe_1_7_1_int_data_0_), .A2(int_data_res_7__1__0_), 
        .ZN(pe_1_7_1_n2) );
  AOI222_X1 pe_1_7_1_U38 ( .A1(pe_1_7_1_n64), .A2(i_data_acc[55]), .B1(
        pe_1_7_1_N85), .B2(pe_1_7_1_n27), .C1(pe_1_7_1_N77), .C2(pe_1_7_1_n28), 
        .ZN(pe_1_7_1_n26) );
  INV_X1 pe_1_7_1_U37 ( .A(pe_1_7_1_n26), .ZN(pe_1_7_1_n77) );
  NOR3_X1 pe_1_7_1_U36 ( .A1(pe_1_7_1_n59), .A2(pe_1_7_1_n65), .A3(int_ckg[6]), 
        .ZN(pe_1_7_1_n36) );
  OR2_X1 pe_1_7_1_U35 ( .A1(pe_1_7_1_n36), .A2(pe_1_7_1_n64), .ZN(pe_1_7_1_N90) );
  INV_X1 pe_1_7_1_U34 ( .A(n41), .ZN(pe_1_7_1_n63) );
  AND2_X1 pe_1_7_1_U33 ( .A1(int_data_x_7__1__2_), .A2(pe_1_7_1_n58), .ZN(
        pe_1_7_1_int_data_2_) );
  AND2_X1 pe_1_7_1_U32 ( .A1(int_data_x_7__1__1_), .A2(pe_1_7_1_n58), .ZN(
        pe_1_7_1_int_data_1_) );
  AND2_X1 pe_1_7_1_U31 ( .A1(int_data_x_7__1__3_), .A2(pe_1_7_1_n58), .ZN(
        pe_1_7_1_int_data_3_) );
  BUF_X1 pe_1_7_1_U30 ( .A(n63), .Z(pe_1_7_1_n64) );
  INV_X1 pe_1_7_1_U29 ( .A(n35), .ZN(pe_1_7_1_n61) );
  AND2_X1 pe_1_7_1_U28 ( .A1(int_data_x_7__1__0_), .A2(pe_1_7_1_n58), .ZN(
        pe_1_7_1_int_data_0_) );
  NAND2_X1 pe_1_7_1_U27 ( .A1(pe_1_7_1_n44), .A2(pe_1_7_1_n61), .ZN(
        pe_1_7_1_n41) );
  AND3_X1 pe_1_7_1_U26 ( .A1(n77), .A2(pe_1_7_1_n63), .A3(n54), .ZN(
        pe_1_7_1_n44) );
  INV_X1 pe_1_7_1_U25 ( .A(pe_1_7_1_int_data_3_), .ZN(pe_1_7_1_n76) );
  NOR2_X1 pe_1_7_1_U24 ( .A1(pe_1_7_1_n70), .A2(n54), .ZN(pe_1_7_1_n43) );
  NOR2_X1 pe_1_7_1_U23 ( .A1(pe_1_7_1_n57), .A2(pe_1_7_1_n64), .ZN(
        pe_1_7_1_n28) );
  NOR2_X1 pe_1_7_1_U22 ( .A1(n21), .A2(pe_1_7_1_n64), .ZN(pe_1_7_1_n27) );
  INV_X1 pe_1_7_1_U21 ( .A(pe_1_7_1_int_data_0_), .ZN(pe_1_7_1_n73) );
  INV_X1 pe_1_7_1_U20 ( .A(pe_1_7_1_n41), .ZN(pe_1_7_1_n90) );
  INV_X1 pe_1_7_1_U19 ( .A(pe_1_7_1_n37), .ZN(pe_1_7_1_n88) );
  INV_X1 pe_1_7_1_U18 ( .A(pe_1_7_1_n38), .ZN(pe_1_7_1_n87) );
  INV_X1 pe_1_7_1_U17 ( .A(pe_1_7_1_n39), .ZN(pe_1_7_1_n86) );
  NOR2_X1 pe_1_7_1_U16 ( .A1(pe_1_7_1_n68), .A2(pe_1_7_1_n42), .ZN(
        pe_1_7_1_N59) );
  NOR2_X1 pe_1_7_1_U15 ( .A1(pe_1_7_1_n68), .A2(pe_1_7_1_n41), .ZN(
        pe_1_7_1_N60) );
  NOR2_X1 pe_1_7_1_U14 ( .A1(pe_1_7_1_n68), .A2(pe_1_7_1_n38), .ZN(
        pe_1_7_1_N63) );
  NOR2_X1 pe_1_7_1_U13 ( .A1(pe_1_7_1_n67), .A2(pe_1_7_1_n40), .ZN(
        pe_1_7_1_N61) );
  NOR2_X1 pe_1_7_1_U12 ( .A1(pe_1_7_1_n67), .A2(pe_1_7_1_n39), .ZN(
        pe_1_7_1_N62) );
  NOR2_X1 pe_1_7_1_U11 ( .A1(pe_1_7_1_n37), .A2(pe_1_7_1_n67), .ZN(
        pe_1_7_1_N64) );
  NAND2_X1 pe_1_7_1_U10 ( .A1(pe_1_7_1_n44), .A2(pe_1_7_1_n60), .ZN(
        pe_1_7_1_n42) );
  BUF_X1 pe_1_7_1_U9 ( .A(pe_1_7_1_n60), .Z(pe_1_7_1_n55) );
  INV_X1 pe_1_7_1_U8 ( .A(pe_1_7_1_n69), .ZN(pe_1_7_1_n65) );
  BUF_X1 pe_1_7_1_U7 ( .A(pe_1_7_1_n60), .Z(pe_1_7_1_n56) );
  INV_X1 pe_1_7_1_U6 ( .A(pe_1_7_1_n42), .ZN(pe_1_7_1_n89) );
  INV_X1 pe_1_7_1_U5 ( .A(pe_1_7_1_n40), .ZN(pe_1_7_1_n85) );
  INV_X2 pe_1_7_1_U4 ( .A(n85), .ZN(pe_1_7_1_n72) );
  XOR2_X1 pe_1_7_1_U3 ( .A(pe_1_7_1_int_data_0_), .B(int_data_res_7__1__0_), 
        .Z(pe_1_7_1_n1) );
  DFFR_X1 pe_1_7_1_int_q_acc_reg_0_ ( .D(pe_1_7_1_n84), .CK(pe_1_7_1_net3106), 
        .RN(pe_1_7_1_n72), .Q(int_data_res_7__1__0_), .QN(pe_1_7_1_n3) );
  DFFR_X1 pe_1_7_1_int_q_reg_v_reg_0__0_ ( .D(i_data_conv_v[24]), .CK(
        pe_1_7_1_net3076), .RN(pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_v[20]) );
  DFFR_X1 pe_1_7_1_int_q_reg_v_reg_0__1_ ( .D(i_data_conv_v[25]), .CK(
        pe_1_7_1_net3076), .RN(pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_v[21]) );
  DFFR_X1 pe_1_7_1_int_q_reg_v_reg_0__2_ ( .D(i_data_conv_v[26]), .CK(
        pe_1_7_1_net3076), .RN(pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_v[22]) );
  DFFR_X1 pe_1_7_1_int_q_reg_v_reg_0__3_ ( .D(i_data_conv_v[27]), .CK(
        pe_1_7_1_net3076), .RN(pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_v[23]) );
  DFFR_X1 pe_1_7_1_int_q_reg_v_reg_1__0_ ( .D(i_data_conv_v[24]), .CK(
        pe_1_7_1_net3081), .RN(pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_v[16]) );
  DFFR_X1 pe_1_7_1_int_q_reg_v_reg_1__1_ ( .D(i_data_conv_v[25]), .CK(
        pe_1_7_1_net3081), .RN(pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_v[17]) );
  DFFR_X1 pe_1_7_1_int_q_reg_v_reg_1__2_ ( .D(i_data_conv_v[26]), .CK(
        pe_1_7_1_net3081), .RN(pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_v[18]) );
  DFFR_X1 pe_1_7_1_int_q_reg_v_reg_1__3_ ( .D(i_data_conv_v[27]), .CK(
        pe_1_7_1_net3081), .RN(pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_v[19]) );
  DFFR_X1 pe_1_7_1_int_q_reg_v_reg_2__0_ ( .D(i_data_conv_v[24]), .CK(
        pe_1_7_1_net3086), .RN(pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_v[12]) );
  DFFR_X1 pe_1_7_1_int_q_reg_v_reg_2__1_ ( .D(i_data_conv_v[25]), .CK(
        pe_1_7_1_net3086), .RN(pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_v[13]) );
  DFFR_X1 pe_1_7_1_int_q_reg_v_reg_2__2_ ( .D(i_data_conv_v[26]), .CK(
        pe_1_7_1_net3086), .RN(pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_v[14]) );
  DFFR_X1 pe_1_7_1_int_q_reg_v_reg_2__3_ ( .D(i_data_conv_v[27]), .CK(
        pe_1_7_1_net3086), .RN(pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_v[15]) );
  DFFR_X1 pe_1_7_1_int_q_reg_v_reg_3__0_ ( .D(i_data_conv_v[24]), .CK(
        pe_1_7_1_net3091), .RN(pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_v[8]) );
  DFFR_X1 pe_1_7_1_int_q_reg_v_reg_3__1_ ( .D(i_data_conv_v[25]), .CK(
        pe_1_7_1_net3091), .RN(pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_v[9]) );
  DFFR_X1 pe_1_7_1_int_q_reg_v_reg_3__2_ ( .D(i_data_conv_v[26]), .CK(
        pe_1_7_1_net3091), .RN(pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_v[10]) );
  DFFR_X1 pe_1_7_1_int_q_reg_v_reg_3__3_ ( .D(i_data_conv_v[27]), .CK(
        pe_1_7_1_net3091), .RN(pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_v[11]) );
  DFFR_X1 pe_1_7_1_int_q_reg_v_reg_4__0_ ( .D(i_data_conv_v[24]), .CK(
        pe_1_7_1_net3096), .RN(pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_v[4]) );
  DFFR_X1 pe_1_7_1_int_q_reg_v_reg_4__1_ ( .D(i_data_conv_v[25]), .CK(
        pe_1_7_1_net3096), .RN(pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_v[5]) );
  DFFR_X1 pe_1_7_1_int_q_reg_v_reg_4__2_ ( .D(i_data_conv_v[26]), .CK(
        pe_1_7_1_net3096), .RN(pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_v[6]) );
  DFFR_X1 pe_1_7_1_int_q_reg_v_reg_4__3_ ( .D(i_data_conv_v[27]), .CK(
        pe_1_7_1_net3096), .RN(pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_v[7]) );
  DFFR_X1 pe_1_7_1_int_q_reg_v_reg_5__0_ ( .D(i_data_conv_v[24]), .CK(
        pe_1_7_1_net3101), .RN(pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_v[0]) );
  DFFR_X1 pe_1_7_1_int_q_reg_v_reg_5__1_ ( .D(i_data_conv_v[25]), .CK(
        pe_1_7_1_net3101), .RN(pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_v[1]) );
  DFFR_X1 pe_1_7_1_int_q_reg_v_reg_5__2_ ( .D(i_data_conv_v[26]), .CK(
        pe_1_7_1_net3101), .RN(pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_v[2]) );
  DFFR_X1 pe_1_7_1_int_q_reg_v_reg_5__3_ ( .D(i_data_conv_v[27]), .CK(
        pe_1_7_1_net3101), .RN(pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_7_1_int_q_reg_h_reg_0__0_ ( .D(int_data_x_7__2__0_), .SI(
        i_data_conv_v[24]), .SE(pe_1_7_1_n65), .CK(pe_1_7_1_net3045), .RN(
        pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_7_1_int_q_reg_h_reg_0__1_ ( .D(int_data_x_7__2__1_), .SI(
        i_data_conv_v[25]), .SE(pe_1_7_1_n65), .CK(pe_1_7_1_net3045), .RN(
        pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_7_1_int_q_reg_h_reg_0__2_ ( .D(int_data_x_7__2__2_), .SI(
        i_data_conv_v[26]), .SE(pe_1_7_1_n65), .CK(pe_1_7_1_net3045), .RN(
        pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_7_1_int_q_reg_h_reg_0__3_ ( .D(int_data_x_7__2__3_), .SI(
        i_data_conv_v[27]), .SE(pe_1_7_1_n65), .CK(pe_1_7_1_net3045), .RN(
        pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_7_1_int_q_reg_h_reg_1__0_ ( .D(int_data_x_7__2__0_), .SI(
        i_data_conv_v[24]), .SE(pe_1_7_1_n65), .CK(pe_1_7_1_net3051), .RN(
        pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_7_1_int_q_reg_h_reg_1__1_ ( .D(int_data_x_7__2__1_), .SI(
        i_data_conv_v[25]), .SE(pe_1_7_1_n65), .CK(pe_1_7_1_net3051), .RN(
        pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_7_1_int_q_reg_h_reg_1__2_ ( .D(int_data_x_7__2__2_), .SI(
        i_data_conv_v[26]), .SE(pe_1_7_1_n65), .CK(pe_1_7_1_net3051), .RN(
        pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_7_1_int_q_reg_h_reg_1__3_ ( .D(int_data_x_7__2__3_), .SI(
        i_data_conv_v[27]), .SE(pe_1_7_1_n65), .CK(pe_1_7_1_net3051), .RN(
        pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_7_1_int_q_reg_h_reg_2__0_ ( .D(int_data_x_7__2__0_), .SI(
        i_data_conv_v[24]), .SE(pe_1_7_1_n65), .CK(pe_1_7_1_net3056), .RN(
        pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_7_1_int_q_reg_h_reg_2__1_ ( .D(int_data_x_7__2__1_), .SI(
        i_data_conv_v[25]), .SE(pe_1_7_1_n65), .CK(pe_1_7_1_net3056), .RN(
        pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_7_1_int_q_reg_h_reg_2__2_ ( .D(int_data_x_7__2__2_), .SI(
        i_data_conv_v[26]), .SE(pe_1_7_1_n65), .CK(pe_1_7_1_net3056), .RN(
        pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_7_1_int_q_reg_h_reg_2__3_ ( .D(int_data_x_7__2__3_), .SI(
        i_data_conv_v[27]), .SE(pe_1_7_1_n65), .CK(pe_1_7_1_net3056), .RN(
        pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_7_1_int_q_reg_h_reg_3__0_ ( .D(int_data_x_7__2__0_), .SI(
        i_data_conv_v[24]), .SE(pe_1_7_1_n65), .CK(pe_1_7_1_net3061), .RN(
        pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_7_1_int_q_reg_h_reg_3__1_ ( .D(int_data_x_7__2__1_), .SI(
        i_data_conv_v[25]), .SE(pe_1_7_1_n65), .CK(pe_1_7_1_net3061), .RN(
        pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_7_1_int_q_reg_h_reg_3__2_ ( .D(int_data_x_7__2__2_), .SI(
        i_data_conv_v[26]), .SE(pe_1_7_1_n65), .CK(pe_1_7_1_net3061), .RN(
        pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_7_1_int_q_reg_h_reg_3__3_ ( .D(int_data_x_7__2__3_), .SI(
        i_data_conv_v[27]), .SE(pe_1_7_1_n65), .CK(pe_1_7_1_net3061), .RN(
        pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_7_1_int_q_reg_h_reg_4__0_ ( .D(int_data_x_7__2__0_), .SI(
        i_data_conv_v[24]), .SE(pe_1_7_1_n66), .CK(pe_1_7_1_net3066), .RN(
        pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_7_1_int_q_reg_h_reg_4__1_ ( .D(int_data_x_7__2__1_), .SI(
        i_data_conv_v[25]), .SE(pe_1_7_1_n66), .CK(pe_1_7_1_net3066), .RN(
        pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_7_1_int_q_reg_h_reg_4__2_ ( .D(int_data_x_7__2__2_), .SI(
        i_data_conv_v[26]), .SE(pe_1_7_1_n66), .CK(pe_1_7_1_net3066), .RN(
        pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_7_1_int_q_reg_h_reg_4__3_ ( .D(int_data_x_7__2__3_), .SI(
        i_data_conv_v[27]), .SE(pe_1_7_1_n66), .CK(pe_1_7_1_net3066), .RN(
        pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_7_1_int_q_reg_h_reg_5__0_ ( .D(int_data_x_7__2__0_), .SI(
        i_data_conv_v[24]), .SE(pe_1_7_1_n66), .CK(pe_1_7_1_net3071), .RN(
        pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_7_1_int_q_reg_h_reg_5__1_ ( .D(int_data_x_7__2__1_), .SI(
        i_data_conv_v[25]), .SE(pe_1_7_1_n66), .CK(pe_1_7_1_net3071), .RN(
        pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_7_1_int_q_reg_h_reg_5__2_ ( .D(int_data_x_7__2__2_), .SI(
        i_data_conv_v[26]), .SE(pe_1_7_1_n66), .CK(pe_1_7_1_net3071), .RN(
        pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_7_1_int_q_reg_h_reg_5__3_ ( .D(int_data_x_7__2__3_), .SI(
        i_data_conv_v[27]), .SE(pe_1_7_1_n66), .CK(pe_1_7_1_net3071), .RN(
        pe_1_7_1_n72), .Q(pe_1_7_1_int_q_reg_h[3]) );
  FA_X1 pe_1_7_1_sub_81_U2_7 ( .A(int_data_res_7__1__7_), .B(pe_1_7_1_n76), 
        .CI(pe_1_7_1_sub_81_carry[7]), .S(pe_1_7_1_N77) );
  FA_X1 pe_1_7_1_sub_81_U2_6 ( .A(int_data_res_7__1__6_), .B(pe_1_7_1_n76), 
        .CI(pe_1_7_1_sub_81_carry[6]), .CO(pe_1_7_1_sub_81_carry[7]), .S(
        pe_1_7_1_N76) );
  FA_X1 pe_1_7_1_sub_81_U2_5 ( .A(int_data_res_7__1__5_), .B(pe_1_7_1_n76), 
        .CI(pe_1_7_1_sub_81_carry[5]), .CO(pe_1_7_1_sub_81_carry[6]), .S(
        pe_1_7_1_N75) );
  FA_X1 pe_1_7_1_sub_81_U2_4 ( .A(int_data_res_7__1__4_), .B(pe_1_7_1_n76), 
        .CI(pe_1_7_1_sub_81_carry[4]), .CO(pe_1_7_1_sub_81_carry[5]), .S(
        pe_1_7_1_N74) );
  FA_X1 pe_1_7_1_sub_81_U2_3 ( .A(int_data_res_7__1__3_), .B(pe_1_7_1_n76), 
        .CI(pe_1_7_1_sub_81_carry[3]), .CO(pe_1_7_1_sub_81_carry[4]), .S(
        pe_1_7_1_N73) );
  FA_X1 pe_1_7_1_sub_81_U2_2 ( .A(int_data_res_7__1__2_), .B(pe_1_7_1_n75), 
        .CI(pe_1_7_1_sub_81_carry[2]), .CO(pe_1_7_1_sub_81_carry[3]), .S(
        pe_1_7_1_N72) );
  FA_X1 pe_1_7_1_sub_81_U2_1 ( .A(int_data_res_7__1__1_), .B(pe_1_7_1_n74), 
        .CI(pe_1_7_1_sub_81_carry[1]), .CO(pe_1_7_1_sub_81_carry[2]), .S(
        pe_1_7_1_N71) );
  FA_X1 pe_1_7_1_add_83_U1_7 ( .A(int_data_res_7__1__7_), .B(
        pe_1_7_1_int_data_3_), .CI(pe_1_7_1_add_83_carry[7]), .S(pe_1_7_1_N85)
         );
  FA_X1 pe_1_7_1_add_83_U1_6 ( .A(int_data_res_7__1__6_), .B(
        pe_1_7_1_int_data_3_), .CI(pe_1_7_1_add_83_carry[6]), .CO(
        pe_1_7_1_add_83_carry[7]), .S(pe_1_7_1_N84) );
  FA_X1 pe_1_7_1_add_83_U1_5 ( .A(int_data_res_7__1__5_), .B(
        pe_1_7_1_int_data_3_), .CI(pe_1_7_1_add_83_carry[5]), .CO(
        pe_1_7_1_add_83_carry[6]), .S(pe_1_7_1_N83) );
  FA_X1 pe_1_7_1_add_83_U1_4 ( .A(int_data_res_7__1__4_), .B(
        pe_1_7_1_int_data_3_), .CI(pe_1_7_1_add_83_carry[4]), .CO(
        pe_1_7_1_add_83_carry[5]), .S(pe_1_7_1_N82) );
  FA_X1 pe_1_7_1_add_83_U1_3 ( .A(int_data_res_7__1__3_), .B(
        pe_1_7_1_int_data_3_), .CI(pe_1_7_1_add_83_carry[3]), .CO(
        pe_1_7_1_add_83_carry[4]), .S(pe_1_7_1_N81) );
  FA_X1 pe_1_7_1_add_83_U1_2 ( .A(int_data_res_7__1__2_), .B(
        pe_1_7_1_int_data_2_), .CI(pe_1_7_1_add_83_carry[2]), .CO(
        pe_1_7_1_add_83_carry[3]), .S(pe_1_7_1_N80) );
  FA_X1 pe_1_7_1_add_83_U1_1 ( .A(int_data_res_7__1__1_), .B(
        pe_1_7_1_int_data_1_), .CI(pe_1_7_1_n2), .CO(pe_1_7_1_add_83_carry[2]), 
        .S(pe_1_7_1_N79) );
  NAND3_X1 pe_1_7_1_U56 ( .A1(pe_1_7_1_n60), .A2(pe_1_7_1_n43), .A3(
        pe_1_7_1_n62), .ZN(pe_1_7_1_n40) );
  NAND3_X1 pe_1_7_1_U55 ( .A1(pe_1_7_1_n43), .A2(pe_1_7_1_n61), .A3(
        pe_1_7_1_n62), .ZN(pe_1_7_1_n39) );
  NAND3_X1 pe_1_7_1_U54 ( .A1(pe_1_7_1_n43), .A2(pe_1_7_1_n63), .A3(
        pe_1_7_1_n60), .ZN(pe_1_7_1_n38) );
  NAND3_X1 pe_1_7_1_U53 ( .A1(pe_1_7_1_n61), .A2(pe_1_7_1_n63), .A3(
        pe_1_7_1_n43), .ZN(pe_1_7_1_n37) );
  DFFR_X1 pe_1_7_1_int_q_acc_reg_6_ ( .D(pe_1_7_1_n78), .CK(pe_1_7_1_net3106), 
        .RN(pe_1_7_1_n71), .Q(int_data_res_7__1__6_) );
  DFFR_X1 pe_1_7_1_int_q_acc_reg_5_ ( .D(pe_1_7_1_n79), .CK(pe_1_7_1_net3106), 
        .RN(pe_1_7_1_n71), .Q(int_data_res_7__1__5_) );
  DFFR_X1 pe_1_7_1_int_q_acc_reg_4_ ( .D(pe_1_7_1_n80), .CK(pe_1_7_1_net3106), 
        .RN(pe_1_7_1_n71), .Q(int_data_res_7__1__4_) );
  DFFR_X1 pe_1_7_1_int_q_acc_reg_3_ ( .D(pe_1_7_1_n81), .CK(pe_1_7_1_net3106), 
        .RN(pe_1_7_1_n71), .Q(int_data_res_7__1__3_) );
  DFFR_X1 pe_1_7_1_int_q_acc_reg_2_ ( .D(pe_1_7_1_n82), .CK(pe_1_7_1_net3106), 
        .RN(pe_1_7_1_n71), .Q(int_data_res_7__1__2_) );
  DFFR_X1 pe_1_7_1_int_q_acc_reg_1_ ( .D(pe_1_7_1_n83), .CK(pe_1_7_1_net3106), 
        .RN(pe_1_7_1_n71), .Q(int_data_res_7__1__1_) );
  DFFR_X1 pe_1_7_1_int_q_acc_reg_7_ ( .D(pe_1_7_1_n77), .CK(pe_1_7_1_net3106), 
        .RN(pe_1_7_1_n71), .Q(int_data_res_7__1__7_) );
  CLKGATETST_X1 pe_1_7_1_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_7_1_n88), .SE(1'b0), .GCK(pe_1_7_1_net3045) );
  CLKGATETST_X1 pe_1_7_1_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_7_1_n87), .SE(1'b0), .GCK(pe_1_7_1_net3051) );
  CLKGATETST_X1 pe_1_7_1_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_7_1_n86), .SE(1'b0), .GCK(pe_1_7_1_net3056) );
  CLKGATETST_X1 pe_1_7_1_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_7_1_n85), .SE(1'b0), .GCK(pe_1_7_1_net3061) );
  CLKGATETST_X1 pe_1_7_1_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_7_1_n90), .SE(1'b0), .GCK(pe_1_7_1_net3066) );
  CLKGATETST_X1 pe_1_7_1_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_7_1_n89), .SE(1'b0), .GCK(pe_1_7_1_net3071) );
  CLKGATETST_X1 pe_1_7_1_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_7_1_N64), .SE(1'b0), .GCK(pe_1_7_1_net3076) );
  CLKGATETST_X1 pe_1_7_1_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_7_1_N63), .SE(1'b0), .GCK(pe_1_7_1_net3081) );
  CLKGATETST_X1 pe_1_7_1_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_7_1_N62), .SE(1'b0), .GCK(pe_1_7_1_net3086) );
  CLKGATETST_X1 pe_1_7_1_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_7_1_N61), .SE(1'b0), .GCK(pe_1_7_1_net3091) );
  CLKGATETST_X1 pe_1_7_1_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_7_1_N60), .SE(1'b0), .GCK(pe_1_7_1_net3096) );
  CLKGATETST_X1 pe_1_7_1_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_7_1_N59), .SE(1'b0), .GCK(pe_1_7_1_net3101) );
  CLKGATETST_X1 pe_1_7_1_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_7_1_N90), .SE(1'b0), .GCK(pe_1_7_1_net3106) );
  CLKBUF_X1 pe_1_7_2_U112 ( .A(pe_1_7_2_n72), .Z(pe_1_7_2_n71) );
  INV_X1 pe_1_7_2_U111 ( .A(n77), .ZN(pe_1_7_2_n70) );
  INV_X1 pe_1_7_2_U110 ( .A(n69), .ZN(pe_1_7_2_n69) );
  INV_X1 pe_1_7_2_U109 ( .A(n69), .ZN(pe_1_7_2_n68) );
  INV_X1 pe_1_7_2_U108 ( .A(n69), .ZN(pe_1_7_2_n67) );
  INV_X1 pe_1_7_2_U107 ( .A(pe_1_7_2_n69), .ZN(pe_1_7_2_n66) );
  INV_X1 pe_1_7_2_U106 ( .A(pe_1_7_2_n63), .ZN(pe_1_7_2_n62) );
  INV_X1 pe_1_7_2_U105 ( .A(pe_1_7_2_n61), .ZN(pe_1_7_2_n60) );
  INV_X1 pe_1_7_2_U104 ( .A(n29), .ZN(pe_1_7_2_n59) );
  INV_X1 pe_1_7_2_U103 ( .A(pe_1_7_2_n59), .ZN(pe_1_7_2_n58) );
  INV_X1 pe_1_7_2_U102 ( .A(n21), .ZN(pe_1_7_2_n57) );
  MUX2_X1 pe_1_7_2_U101 ( .A(pe_1_7_2_n54), .B(pe_1_7_2_n51), .S(n54), .Z(
        int_data_x_7__2__3_) );
  MUX2_X1 pe_1_7_2_U100 ( .A(pe_1_7_2_n53), .B(pe_1_7_2_n52), .S(pe_1_7_2_n62), 
        .Z(pe_1_7_2_n54) );
  MUX2_X1 pe_1_7_2_U99 ( .A(pe_1_7_2_int_q_reg_h[23]), .B(
        pe_1_7_2_int_q_reg_h[19]), .S(pe_1_7_2_n56), .Z(pe_1_7_2_n53) );
  MUX2_X1 pe_1_7_2_U98 ( .A(pe_1_7_2_int_q_reg_h[15]), .B(
        pe_1_7_2_int_q_reg_h[11]), .S(pe_1_7_2_n56), .Z(pe_1_7_2_n52) );
  MUX2_X1 pe_1_7_2_U97 ( .A(pe_1_7_2_int_q_reg_h[7]), .B(
        pe_1_7_2_int_q_reg_h[3]), .S(pe_1_7_2_n56), .Z(pe_1_7_2_n51) );
  MUX2_X1 pe_1_7_2_U96 ( .A(pe_1_7_2_n50), .B(pe_1_7_2_n47), .S(n54), .Z(
        int_data_x_7__2__2_) );
  MUX2_X1 pe_1_7_2_U95 ( .A(pe_1_7_2_n49), .B(pe_1_7_2_n48), .S(pe_1_7_2_n62), 
        .Z(pe_1_7_2_n50) );
  MUX2_X1 pe_1_7_2_U94 ( .A(pe_1_7_2_int_q_reg_h[22]), .B(
        pe_1_7_2_int_q_reg_h[18]), .S(pe_1_7_2_n56), .Z(pe_1_7_2_n49) );
  MUX2_X1 pe_1_7_2_U93 ( .A(pe_1_7_2_int_q_reg_h[14]), .B(
        pe_1_7_2_int_q_reg_h[10]), .S(pe_1_7_2_n56), .Z(pe_1_7_2_n48) );
  MUX2_X1 pe_1_7_2_U92 ( .A(pe_1_7_2_int_q_reg_h[6]), .B(
        pe_1_7_2_int_q_reg_h[2]), .S(pe_1_7_2_n56), .Z(pe_1_7_2_n47) );
  MUX2_X1 pe_1_7_2_U91 ( .A(pe_1_7_2_n46), .B(pe_1_7_2_n24), .S(n54), .Z(
        int_data_x_7__2__1_) );
  MUX2_X1 pe_1_7_2_U90 ( .A(pe_1_7_2_n45), .B(pe_1_7_2_n25), .S(pe_1_7_2_n62), 
        .Z(pe_1_7_2_n46) );
  MUX2_X1 pe_1_7_2_U89 ( .A(pe_1_7_2_int_q_reg_h[21]), .B(
        pe_1_7_2_int_q_reg_h[17]), .S(pe_1_7_2_n56), .Z(pe_1_7_2_n45) );
  MUX2_X1 pe_1_7_2_U88 ( .A(pe_1_7_2_int_q_reg_h[13]), .B(
        pe_1_7_2_int_q_reg_h[9]), .S(pe_1_7_2_n56), .Z(pe_1_7_2_n25) );
  MUX2_X1 pe_1_7_2_U87 ( .A(pe_1_7_2_int_q_reg_h[5]), .B(
        pe_1_7_2_int_q_reg_h[1]), .S(pe_1_7_2_n56), .Z(pe_1_7_2_n24) );
  MUX2_X1 pe_1_7_2_U86 ( .A(pe_1_7_2_n23), .B(pe_1_7_2_n20), .S(n54), .Z(
        int_data_x_7__2__0_) );
  MUX2_X1 pe_1_7_2_U85 ( .A(pe_1_7_2_n22), .B(pe_1_7_2_n21), .S(pe_1_7_2_n62), 
        .Z(pe_1_7_2_n23) );
  MUX2_X1 pe_1_7_2_U84 ( .A(pe_1_7_2_int_q_reg_h[20]), .B(
        pe_1_7_2_int_q_reg_h[16]), .S(pe_1_7_2_n56), .Z(pe_1_7_2_n22) );
  MUX2_X1 pe_1_7_2_U83 ( .A(pe_1_7_2_int_q_reg_h[12]), .B(
        pe_1_7_2_int_q_reg_h[8]), .S(pe_1_7_2_n56), .Z(pe_1_7_2_n21) );
  MUX2_X1 pe_1_7_2_U82 ( .A(pe_1_7_2_int_q_reg_h[4]), .B(
        pe_1_7_2_int_q_reg_h[0]), .S(pe_1_7_2_n56), .Z(pe_1_7_2_n20) );
  MUX2_X1 pe_1_7_2_U81 ( .A(pe_1_7_2_n19), .B(pe_1_7_2_n16), .S(n54), .Z(
        int_data_y_7__2__3_) );
  MUX2_X1 pe_1_7_2_U80 ( .A(pe_1_7_2_n18), .B(pe_1_7_2_n17), .S(pe_1_7_2_n62), 
        .Z(pe_1_7_2_n19) );
  MUX2_X1 pe_1_7_2_U79 ( .A(pe_1_7_2_int_q_reg_v[23]), .B(
        pe_1_7_2_int_q_reg_v[19]), .S(pe_1_7_2_n55), .Z(pe_1_7_2_n18) );
  MUX2_X1 pe_1_7_2_U78 ( .A(pe_1_7_2_int_q_reg_v[15]), .B(
        pe_1_7_2_int_q_reg_v[11]), .S(pe_1_7_2_n55), .Z(pe_1_7_2_n17) );
  MUX2_X1 pe_1_7_2_U77 ( .A(pe_1_7_2_int_q_reg_v[7]), .B(
        pe_1_7_2_int_q_reg_v[3]), .S(pe_1_7_2_n55), .Z(pe_1_7_2_n16) );
  MUX2_X1 pe_1_7_2_U76 ( .A(pe_1_7_2_n15), .B(pe_1_7_2_n12), .S(n54), .Z(
        int_data_y_7__2__2_) );
  MUX2_X1 pe_1_7_2_U75 ( .A(pe_1_7_2_n14), .B(pe_1_7_2_n13), .S(pe_1_7_2_n62), 
        .Z(pe_1_7_2_n15) );
  MUX2_X1 pe_1_7_2_U74 ( .A(pe_1_7_2_int_q_reg_v[22]), .B(
        pe_1_7_2_int_q_reg_v[18]), .S(pe_1_7_2_n55), .Z(pe_1_7_2_n14) );
  MUX2_X1 pe_1_7_2_U73 ( .A(pe_1_7_2_int_q_reg_v[14]), .B(
        pe_1_7_2_int_q_reg_v[10]), .S(pe_1_7_2_n55), .Z(pe_1_7_2_n13) );
  MUX2_X1 pe_1_7_2_U72 ( .A(pe_1_7_2_int_q_reg_v[6]), .B(
        pe_1_7_2_int_q_reg_v[2]), .S(pe_1_7_2_n55), .Z(pe_1_7_2_n12) );
  MUX2_X1 pe_1_7_2_U71 ( .A(pe_1_7_2_n11), .B(pe_1_7_2_n8), .S(n54), .Z(
        int_data_y_7__2__1_) );
  MUX2_X1 pe_1_7_2_U70 ( .A(pe_1_7_2_n10), .B(pe_1_7_2_n9), .S(pe_1_7_2_n62), 
        .Z(pe_1_7_2_n11) );
  MUX2_X1 pe_1_7_2_U69 ( .A(pe_1_7_2_int_q_reg_v[21]), .B(
        pe_1_7_2_int_q_reg_v[17]), .S(pe_1_7_2_n55), .Z(pe_1_7_2_n10) );
  MUX2_X1 pe_1_7_2_U68 ( .A(pe_1_7_2_int_q_reg_v[13]), .B(
        pe_1_7_2_int_q_reg_v[9]), .S(pe_1_7_2_n55), .Z(pe_1_7_2_n9) );
  MUX2_X1 pe_1_7_2_U67 ( .A(pe_1_7_2_int_q_reg_v[5]), .B(
        pe_1_7_2_int_q_reg_v[1]), .S(pe_1_7_2_n55), .Z(pe_1_7_2_n8) );
  MUX2_X1 pe_1_7_2_U66 ( .A(pe_1_7_2_n7), .B(pe_1_7_2_n4), .S(n54), .Z(
        int_data_y_7__2__0_) );
  MUX2_X1 pe_1_7_2_U65 ( .A(pe_1_7_2_n6), .B(pe_1_7_2_n5), .S(pe_1_7_2_n62), 
        .Z(pe_1_7_2_n7) );
  MUX2_X1 pe_1_7_2_U64 ( .A(pe_1_7_2_int_q_reg_v[20]), .B(
        pe_1_7_2_int_q_reg_v[16]), .S(pe_1_7_2_n55), .Z(pe_1_7_2_n6) );
  MUX2_X1 pe_1_7_2_U63 ( .A(pe_1_7_2_int_q_reg_v[12]), .B(
        pe_1_7_2_int_q_reg_v[8]), .S(pe_1_7_2_n55), .Z(pe_1_7_2_n5) );
  MUX2_X1 pe_1_7_2_U62 ( .A(pe_1_7_2_int_q_reg_v[4]), .B(
        pe_1_7_2_int_q_reg_v[0]), .S(pe_1_7_2_n55), .Z(pe_1_7_2_n4) );
  AOI222_X1 pe_1_7_2_U61 ( .A1(i_data_acc[42]), .A2(pe_1_7_2_n64), .B1(
        pe_1_7_2_N80), .B2(pe_1_7_2_n27), .C1(pe_1_7_2_N72), .C2(pe_1_7_2_n28), 
        .ZN(pe_1_7_2_n33) );
  INV_X1 pe_1_7_2_U60 ( .A(pe_1_7_2_n33), .ZN(pe_1_7_2_n82) );
  AOI222_X1 pe_1_7_2_U59 ( .A1(i_data_acc[46]), .A2(pe_1_7_2_n64), .B1(
        pe_1_7_2_N84), .B2(pe_1_7_2_n27), .C1(pe_1_7_2_N76), .C2(pe_1_7_2_n28), 
        .ZN(pe_1_7_2_n29) );
  INV_X1 pe_1_7_2_U58 ( .A(pe_1_7_2_n29), .ZN(pe_1_7_2_n78) );
  XNOR2_X1 pe_1_7_2_U57 ( .A(pe_1_7_2_n73), .B(int_data_res_7__2__0_), .ZN(
        pe_1_7_2_N70) );
  AOI222_X1 pe_1_7_2_U52 ( .A1(i_data_acc[40]), .A2(pe_1_7_2_n64), .B1(
        pe_1_7_2_n1), .B2(pe_1_7_2_n27), .C1(pe_1_7_2_N70), .C2(pe_1_7_2_n28), 
        .ZN(pe_1_7_2_n35) );
  INV_X1 pe_1_7_2_U51 ( .A(pe_1_7_2_n35), .ZN(pe_1_7_2_n84) );
  AOI222_X1 pe_1_7_2_U50 ( .A1(i_data_acc[41]), .A2(pe_1_7_2_n64), .B1(
        pe_1_7_2_N79), .B2(pe_1_7_2_n27), .C1(pe_1_7_2_N71), .C2(pe_1_7_2_n28), 
        .ZN(pe_1_7_2_n34) );
  INV_X1 pe_1_7_2_U49 ( .A(pe_1_7_2_n34), .ZN(pe_1_7_2_n83) );
  AOI222_X1 pe_1_7_2_U48 ( .A1(i_data_acc[43]), .A2(pe_1_7_2_n64), .B1(
        pe_1_7_2_N81), .B2(pe_1_7_2_n27), .C1(pe_1_7_2_N73), .C2(pe_1_7_2_n28), 
        .ZN(pe_1_7_2_n32) );
  INV_X1 pe_1_7_2_U47 ( .A(pe_1_7_2_n32), .ZN(pe_1_7_2_n81) );
  AOI222_X1 pe_1_7_2_U46 ( .A1(i_data_acc[44]), .A2(pe_1_7_2_n64), .B1(
        pe_1_7_2_N82), .B2(pe_1_7_2_n27), .C1(pe_1_7_2_N74), .C2(pe_1_7_2_n28), 
        .ZN(pe_1_7_2_n31) );
  INV_X1 pe_1_7_2_U45 ( .A(pe_1_7_2_n31), .ZN(pe_1_7_2_n80) );
  AOI222_X1 pe_1_7_2_U44 ( .A1(i_data_acc[45]), .A2(pe_1_7_2_n64), .B1(
        pe_1_7_2_N83), .B2(pe_1_7_2_n27), .C1(pe_1_7_2_N75), .C2(pe_1_7_2_n28), 
        .ZN(pe_1_7_2_n30) );
  INV_X1 pe_1_7_2_U43 ( .A(pe_1_7_2_n30), .ZN(pe_1_7_2_n79) );
  NAND2_X1 pe_1_7_2_U42 ( .A1(pe_1_7_2_int_data_0_), .A2(pe_1_7_2_n3), .ZN(
        pe_1_7_2_sub_81_carry[1]) );
  INV_X1 pe_1_7_2_U41 ( .A(pe_1_7_2_int_data_1_), .ZN(pe_1_7_2_n74) );
  INV_X1 pe_1_7_2_U40 ( .A(pe_1_7_2_int_data_2_), .ZN(pe_1_7_2_n75) );
  AND2_X1 pe_1_7_2_U39 ( .A1(pe_1_7_2_int_data_0_), .A2(int_data_res_7__2__0_), 
        .ZN(pe_1_7_2_n2) );
  AOI222_X1 pe_1_7_2_U38 ( .A1(pe_1_7_2_n64), .A2(i_data_acc[47]), .B1(
        pe_1_7_2_N85), .B2(pe_1_7_2_n27), .C1(pe_1_7_2_N77), .C2(pe_1_7_2_n28), 
        .ZN(pe_1_7_2_n26) );
  INV_X1 pe_1_7_2_U37 ( .A(pe_1_7_2_n26), .ZN(pe_1_7_2_n77) );
  NOR3_X1 pe_1_7_2_U36 ( .A1(pe_1_7_2_n59), .A2(pe_1_7_2_n65), .A3(int_ckg[5]), 
        .ZN(pe_1_7_2_n36) );
  OR2_X1 pe_1_7_2_U35 ( .A1(pe_1_7_2_n36), .A2(pe_1_7_2_n64), .ZN(pe_1_7_2_N90) );
  INV_X1 pe_1_7_2_U34 ( .A(n41), .ZN(pe_1_7_2_n63) );
  AND2_X1 pe_1_7_2_U33 ( .A1(int_data_x_7__2__2_), .A2(pe_1_7_2_n58), .ZN(
        pe_1_7_2_int_data_2_) );
  AND2_X1 pe_1_7_2_U32 ( .A1(int_data_x_7__2__1_), .A2(pe_1_7_2_n58), .ZN(
        pe_1_7_2_int_data_1_) );
  AND2_X1 pe_1_7_2_U31 ( .A1(int_data_x_7__2__3_), .A2(pe_1_7_2_n58), .ZN(
        pe_1_7_2_int_data_3_) );
  BUF_X1 pe_1_7_2_U30 ( .A(n63), .Z(pe_1_7_2_n64) );
  INV_X1 pe_1_7_2_U29 ( .A(n35), .ZN(pe_1_7_2_n61) );
  AND2_X1 pe_1_7_2_U28 ( .A1(int_data_x_7__2__0_), .A2(pe_1_7_2_n58), .ZN(
        pe_1_7_2_int_data_0_) );
  NAND2_X1 pe_1_7_2_U27 ( .A1(pe_1_7_2_n44), .A2(pe_1_7_2_n61), .ZN(
        pe_1_7_2_n41) );
  AND3_X1 pe_1_7_2_U26 ( .A1(n77), .A2(pe_1_7_2_n63), .A3(n54), .ZN(
        pe_1_7_2_n44) );
  INV_X1 pe_1_7_2_U25 ( .A(pe_1_7_2_int_data_3_), .ZN(pe_1_7_2_n76) );
  NOR2_X1 pe_1_7_2_U24 ( .A1(pe_1_7_2_n70), .A2(n54), .ZN(pe_1_7_2_n43) );
  NOR2_X1 pe_1_7_2_U23 ( .A1(pe_1_7_2_n57), .A2(pe_1_7_2_n64), .ZN(
        pe_1_7_2_n28) );
  NOR2_X1 pe_1_7_2_U22 ( .A1(n21), .A2(pe_1_7_2_n64), .ZN(pe_1_7_2_n27) );
  INV_X1 pe_1_7_2_U21 ( .A(pe_1_7_2_int_data_0_), .ZN(pe_1_7_2_n73) );
  INV_X1 pe_1_7_2_U20 ( .A(pe_1_7_2_n41), .ZN(pe_1_7_2_n90) );
  INV_X1 pe_1_7_2_U19 ( .A(pe_1_7_2_n37), .ZN(pe_1_7_2_n88) );
  INV_X1 pe_1_7_2_U18 ( .A(pe_1_7_2_n38), .ZN(pe_1_7_2_n87) );
  INV_X1 pe_1_7_2_U17 ( .A(pe_1_7_2_n39), .ZN(pe_1_7_2_n86) );
  NOR2_X1 pe_1_7_2_U16 ( .A1(pe_1_7_2_n68), .A2(pe_1_7_2_n42), .ZN(
        pe_1_7_2_N59) );
  NOR2_X1 pe_1_7_2_U15 ( .A1(pe_1_7_2_n68), .A2(pe_1_7_2_n41), .ZN(
        pe_1_7_2_N60) );
  NOR2_X1 pe_1_7_2_U14 ( .A1(pe_1_7_2_n68), .A2(pe_1_7_2_n38), .ZN(
        pe_1_7_2_N63) );
  NOR2_X1 pe_1_7_2_U13 ( .A1(pe_1_7_2_n67), .A2(pe_1_7_2_n40), .ZN(
        pe_1_7_2_N61) );
  NOR2_X1 pe_1_7_2_U12 ( .A1(pe_1_7_2_n67), .A2(pe_1_7_2_n39), .ZN(
        pe_1_7_2_N62) );
  NOR2_X1 pe_1_7_2_U11 ( .A1(pe_1_7_2_n37), .A2(pe_1_7_2_n67), .ZN(
        pe_1_7_2_N64) );
  NAND2_X1 pe_1_7_2_U10 ( .A1(pe_1_7_2_n44), .A2(pe_1_7_2_n60), .ZN(
        pe_1_7_2_n42) );
  BUF_X1 pe_1_7_2_U9 ( .A(pe_1_7_2_n60), .Z(pe_1_7_2_n55) );
  INV_X1 pe_1_7_2_U8 ( .A(pe_1_7_2_n69), .ZN(pe_1_7_2_n65) );
  BUF_X1 pe_1_7_2_U7 ( .A(pe_1_7_2_n60), .Z(pe_1_7_2_n56) );
  INV_X1 pe_1_7_2_U6 ( .A(pe_1_7_2_n42), .ZN(pe_1_7_2_n89) );
  INV_X1 pe_1_7_2_U5 ( .A(pe_1_7_2_n40), .ZN(pe_1_7_2_n85) );
  INV_X2 pe_1_7_2_U4 ( .A(n85), .ZN(pe_1_7_2_n72) );
  XOR2_X1 pe_1_7_2_U3 ( .A(pe_1_7_2_int_data_0_), .B(int_data_res_7__2__0_), 
        .Z(pe_1_7_2_n1) );
  DFFR_X1 pe_1_7_2_int_q_acc_reg_0_ ( .D(pe_1_7_2_n84), .CK(pe_1_7_2_net3028), 
        .RN(pe_1_7_2_n72), .Q(int_data_res_7__2__0_), .QN(pe_1_7_2_n3) );
  DFFR_X1 pe_1_7_2_int_q_reg_v_reg_0__0_ ( .D(i_data_conv_v[20]), .CK(
        pe_1_7_2_net2998), .RN(pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_v[20]) );
  DFFR_X1 pe_1_7_2_int_q_reg_v_reg_0__1_ ( .D(i_data_conv_v[21]), .CK(
        pe_1_7_2_net2998), .RN(pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_v[21]) );
  DFFR_X1 pe_1_7_2_int_q_reg_v_reg_0__2_ ( .D(i_data_conv_v[22]), .CK(
        pe_1_7_2_net2998), .RN(pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_v[22]) );
  DFFR_X1 pe_1_7_2_int_q_reg_v_reg_0__3_ ( .D(i_data_conv_v[23]), .CK(
        pe_1_7_2_net2998), .RN(pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_v[23]) );
  DFFR_X1 pe_1_7_2_int_q_reg_v_reg_1__0_ ( .D(i_data_conv_v[20]), .CK(
        pe_1_7_2_net3003), .RN(pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_v[16]) );
  DFFR_X1 pe_1_7_2_int_q_reg_v_reg_1__1_ ( .D(i_data_conv_v[21]), .CK(
        pe_1_7_2_net3003), .RN(pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_v[17]) );
  DFFR_X1 pe_1_7_2_int_q_reg_v_reg_1__2_ ( .D(i_data_conv_v[22]), .CK(
        pe_1_7_2_net3003), .RN(pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_v[18]) );
  DFFR_X1 pe_1_7_2_int_q_reg_v_reg_1__3_ ( .D(i_data_conv_v[23]), .CK(
        pe_1_7_2_net3003), .RN(pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_v[19]) );
  DFFR_X1 pe_1_7_2_int_q_reg_v_reg_2__0_ ( .D(i_data_conv_v[20]), .CK(
        pe_1_7_2_net3008), .RN(pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_v[12]) );
  DFFR_X1 pe_1_7_2_int_q_reg_v_reg_2__1_ ( .D(i_data_conv_v[21]), .CK(
        pe_1_7_2_net3008), .RN(pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_v[13]) );
  DFFR_X1 pe_1_7_2_int_q_reg_v_reg_2__2_ ( .D(i_data_conv_v[22]), .CK(
        pe_1_7_2_net3008), .RN(pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_v[14]) );
  DFFR_X1 pe_1_7_2_int_q_reg_v_reg_2__3_ ( .D(i_data_conv_v[23]), .CK(
        pe_1_7_2_net3008), .RN(pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_v[15]) );
  DFFR_X1 pe_1_7_2_int_q_reg_v_reg_3__0_ ( .D(i_data_conv_v[20]), .CK(
        pe_1_7_2_net3013), .RN(pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_v[8]) );
  DFFR_X1 pe_1_7_2_int_q_reg_v_reg_3__1_ ( .D(i_data_conv_v[21]), .CK(
        pe_1_7_2_net3013), .RN(pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_v[9]) );
  DFFR_X1 pe_1_7_2_int_q_reg_v_reg_3__2_ ( .D(i_data_conv_v[22]), .CK(
        pe_1_7_2_net3013), .RN(pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_v[10]) );
  DFFR_X1 pe_1_7_2_int_q_reg_v_reg_3__3_ ( .D(i_data_conv_v[23]), .CK(
        pe_1_7_2_net3013), .RN(pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_v[11]) );
  DFFR_X1 pe_1_7_2_int_q_reg_v_reg_4__0_ ( .D(i_data_conv_v[20]), .CK(
        pe_1_7_2_net3018), .RN(pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_v[4]) );
  DFFR_X1 pe_1_7_2_int_q_reg_v_reg_4__1_ ( .D(i_data_conv_v[21]), .CK(
        pe_1_7_2_net3018), .RN(pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_v[5]) );
  DFFR_X1 pe_1_7_2_int_q_reg_v_reg_4__2_ ( .D(i_data_conv_v[22]), .CK(
        pe_1_7_2_net3018), .RN(pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_v[6]) );
  DFFR_X1 pe_1_7_2_int_q_reg_v_reg_4__3_ ( .D(i_data_conv_v[23]), .CK(
        pe_1_7_2_net3018), .RN(pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_v[7]) );
  DFFR_X1 pe_1_7_2_int_q_reg_v_reg_5__0_ ( .D(i_data_conv_v[20]), .CK(
        pe_1_7_2_net3023), .RN(pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_v[0]) );
  DFFR_X1 pe_1_7_2_int_q_reg_v_reg_5__1_ ( .D(i_data_conv_v[21]), .CK(
        pe_1_7_2_net3023), .RN(pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_v[1]) );
  DFFR_X1 pe_1_7_2_int_q_reg_v_reg_5__2_ ( .D(i_data_conv_v[22]), .CK(
        pe_1_7_2_net3023), .RN(pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_v[2]) );
  DFFR_X1 pe_1_7_2_int_q_reg_v_reg_5__3_ ( .D(i_data_conv_v[23]), .CK(
        pe_1_7_2_net3023), .RN(pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_7_2_int_q_reg_h_reg_0__0_ ( .D(int_data_x_7__3__0_), .SI(
        i_data_conv_v[20]), .SE(pe_1_7_2_n65), .CK(pe_1_7_2_net2967), .RN(
        pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_7_2_int_q_reg_h_reg_0__1_ ( .D(int_data_x_7__3__1_), .SI(
        i_data_conv_v[21]), .SE(pe_1_7_2_n65), .CK(pe_1_7_2_net2967), .RN(
        pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_7_2_int_q_reg_h_reg_0__2_ ( .D(int_data_x_7__3__2_), .SI(
        i_data_conv_v[22]), .SE(pe_1_7_2_n65), .CK(pe_1_7_2_net2967), .RN(
        pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_7_2_int_q_reg_h_reg_0__3_ ( .D(int_data_x_7__3__3_), .SI(
        i_data_conv_v[23]), .SE(pe_1_7_2_n65), .CK(pe_1_7_2_net2967), .RN(
        pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_7_2_int_q_reg_h_reg_1__0_ ( .D(int_data_x_7__3__0_), .SI(
        i_data_conv_v[20]), .SE(pe_1_7_2_n65), .CK(pe_1_7_2_net2973), .RN(
        pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_7_2_int_q_reg_h_reg_1__1_ ( .D(int_data_x_7__3__1_), .SI(
        i_data_conv_v[21]), .SE(pe_1_7_2_n65), .CK(pe_1_7_2_net2973), .RN(
        pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_7_2_int_q_reg_h_reg_1__2_ ( .D(int_data_x_7__3__2_), .SI(
        i_data_conv_v[22]), .SE(pe_1_7_2_n65), .CK(pe_1_7_2_net2973), .RN(
        pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_7_2_int_q_reg_h_reg_1__3_ ( .D(int_data_x_7__3__3_), .SI(
        i_data_conv_v[23]), .SE(pe_1_7_2_n65), .CK(pe_1_7_2_net2973), .RN(
        pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_7_2_int_q_reg_h_reg_2__0_ ( .D(int_data_x_7__3__0_), .SI(
        i_data_conv_v[20]), .SE(pe_1_7_2_n65), .CK(pe_1_7_2_net2978), .RN(
        pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_7_2_int_q_reg_h_reg_2__1_ ( .D(int_data_x_7__3__1_), .SI(
        i_data_conv_v[21]), .SE(pe_1_7_2_n65), .CK(pe_1_7_2_net2978), .RN(
        pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_7_2_int_q_reg_h_reg_2__2_ ( .D(int_data_x_7__3__2_), .SI(
        i_data_conv_v[22]), .SE(pe_1_7_2_n65), .CK(pe_1_7_2_net2978), .RN(
        pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_7_2_int_q_reg_h_reg_2__3_ ( .D(int_data_x_7__3__3_), .SI(
        i_data_conv_v[23]), .SE(pe_1_7_2_n65), .CK(pe_1_7_2_net2978), .RN(
        pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_7_2_int_q_reg_h_reg_3__0_ ( .D(int_data_x_7__3__0_), .SI(
        i_data_conv_v[20]), .SE(pe_1_7_2_n65), .CK(pe_1_7_2_net2983), .RN(
        pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_7_2_int_q_reg_h_reg_3__1_ ( .D(int_data_x_7__3__1_), .SI(
        i_data_conv_v[21]), .SE(pe_1_7_2_n65), .CK(pe_1_7_2_net2983), .RN(
        pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_7_2_int_q_reg_h_reg_3__2_ ( .D(int_data_x_7__3__2_), .SI(
        i_data_conv_v[22]), .SE(pe_1_7_2_n65), .CK(pe_1_7_2_net2983), .RN(
        pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_7_2_int_q_reg_h_reg_3__3_ ( .D(int_data_x_7__3__3_), .SI(
        i_data_conv_v[23]), .SE(pe_1_7_2_n65), .CK(pe_1_7_2_net2983), .RN(
        pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_7_2_int_q_reg_h_reg_4__0_ ( .D(int_data_x_7__3__0_), .SI(
        i_data_conv_v[20]), .SE(pe_1_7_2_n66), .CK(pe_1_7_2_net2988), .RN(
        pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_7_2_int_q_reg_h_reg_4__1_ ( .D(int_data_x_7__3__1_), .SI(
        i_data_conv_v[21]), .SE(pe_1_7_2_n66), .CK(pe_1_7_2_net2988), .RN(
        pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_7_2_int_q_reg_h_reg_4__2_ ( .D(int_data_x_7__3__2_), .SI(
        i_data_conv_v[22]), .SE(pe_1_7_2_n66), .CK(pe_1_7_2_net2988), .RN(
        pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_7_2_int_q_reg_h_reg_4__3_ ( .D(int_data_x_7__3__3_), .SI(
        i_data_conv_v[23]), .SE(pe_1_7_2_n66), .CK(pe_1_7_2_net2988), .RN(
        pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_7_2_int_q_reg_h_reg_5__0_ ( .D(int_data_x_7__3__0_), .SI(
        i_data_conv_v[20]), .SE(pe_1_7_2_n66), .CK(pe_1_7_2_net2993), .RN(
        pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_7_2_int_q_reg_h_reg_5__1_ ( .D(int_data_x_7__3__1_), .SI(
        i_data_conv_v[21]), .SE(pe_1_7_2_n66), .CK(pe_1_7_2_net2993), .RN(
        pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_7_2_int_q_reg_h_reg_5__2_ ( .D(int_data_x_7__3__2_), .SI(
        i_data_conv_v[22]), .SE(pe_1_7_2_n66), .CK(pe_1_7_2_net2993), .RN(
        pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_7_2_int_q_reg_h_reg_5__3_ ( .D(int_data_x_7__3__3_), .SI(
        i_data_conv_v[23]), .SE(pe_1_7_2_n66), .CK(pe_1_7_2_net2993), .RN(
        pe_1_7_2_n72), .Q(pe_1_7_2_int_q_reg_h[3]) );
  FA_X1 pe_1_7_2_sub_81_U2_7 ( .A(int_data_res_7__2__7_), .B(pe_1_7_2_n76), 
        .CI(pe_1_7_2_sub_81_carry[7]), .S(pe_1_7_2_N77) );
  FA_X1 pe_1_7_2_sub_81_U2_6 ( .A(int_data_res_7__2__6_), .B(pe_1_7_2_n76), 
        .CI(pe_1_7_2_sub_81_carry[6]), .CO(pe_1_7_2_sub_81_carry[7]), .S(
        pe_1_7_2_N76) );
  FA_X1 pe_1_7_2_sub_81_U2_5 ( .A(int_data_res_7__2__5_), .B(pe_1_7_2_n76), 
        .CI(pe_1_7_2_sub_81_carry[5]), .CO(pe_1_7_2_sub_81_carry[6]), .S(
        pe_1_7_2_N75) );
  FA_X1 pe_1_7_2_sub_81_U2_4 ( .A(int_data_res_7__2__4_), .B(pe_1_7_2_n76), 
        .CI(pe_1_7_2_sub_81_carry[4]), .CO(pe_1_7_2_sub_81_carry[5]), .S(
        pe_1_7_2_N74) );
  FA_X1 pe_1_7_2_sub_81_U2_3 ( .A(int_data_res_7__2__3_), .B(pe_1_7_2_n76), 
        .CI(pe_1_7_2_sub_81_carry[3]), .CO(pe_1_7_2_sub_81_carry[4]), .S(
        pe_1_7_2_N73) );
  FA_X1 pe_1_7_2_sub_81_U2_2 ( .A(int_data_res_7__2__2_), .B(pe_1_7_2_n75), 
        .CI(pe_1_7_2_sub_81_carry[2]), .CO(pe_1_7_2_sub_81_carry[3]), .S(
        pe_1_7_2_N72) );
  FA_X1 pe_1_7_2_sub_81_U2_1 ( .A(int_data_res_7__2__1_), .B(pe_1_7_2_n74), 
        .CI(pe_1_7_2_sub_81_carry[1]), .CO(pe_1_7_2_sub_81_carry[2]), .S(
        pe_1_7_2_N71) );
  FA_X1 pe_1_7_2_add_83_U1_7 ( .A(int_data_res_7__2__7_), .B(
        pe_1_7_2_int_data_3_), .CI(pe_1_7_2_add_83_carry[7]), .S(pe_1_7_2_N85)
         );
  FA_X1 pe_1_7_2_add_83_U1_6 ( .A(int_data_res_7__2__6_), .B(
        pe_1_7_2_int_data_3_), .CI(pe_1_7_2_add_83_carry[6]), .CO(
        pe_1_7_2_add_83_carry[7]), .S(pe_1_7_2_N84) );
  FA_X1 pe_1_7_2_add_83_U1_5 ( .A(int_data_res_7__2__5_), .B(
        pe_1_7_2_int_data_3_), .CI(pe_1_7_2_add_83_carry[5]), .CO(
        pe_1_7_2_add_83_carry[6]), .S(pe_1_7_2_N83) );
  FA_X1 pe_1_7_2_add_83_U1_4 ( .A(int_data_res_7__2__4_), .B(
        pe_1_7_2_int_data_3_), .CI(pe_1_7_2_add_83_carry[4]), .CO(
        pe_1_7_2_add_83_carry[5]), .S(pe_1_7_2_N82) );
  FA_X1 pe_1_7_2_add_83_U1_3 ( .A(int_data_res_7__2__3_), .B(
        pe_1_7_2_int_data_3_), .CI(pe_1_7_2_add_83_carry[3]), .CO(
        pe_1_7_2_add_83_carry[4]), .S(pe_1_7_2_N81) );
  FA_X1 pe_1_7_2_add_83_U1_2 ( .A(int_data_res_7__2__2_), .B(
        pe_1_7_2_int_data_2_), .CI(pe_1_7_2_add_83_carry[2]), .CO(
        pe_1_7_2_add_83_carry[3]), .S(pe_1_7_2_N80) );
  FA_X1 pe_1_7_2_add_83_U1_1 ( .A(int_data_res_7__2__1_), .B(
        pe_1_7_2_int_data_1_), .CI(pe_1_7_2_n2), .CO(pe_1_7_2_add_83_carry[2]), 
        .S(pe_1_7_2_N79) );
  NAND3_X1 pe_1_7_2_U56 ( .A1(pe_1_7_2_n60), .A2(pe_1_7_2_n43), .A3(
        pe_1_7_2_n62), .ZN(pe_1_7_2_n40) );
  NAND3_X1 pe_1_7_2_U55 ( .A1(pe_1_7_2_n43), .A2(pe_1_7_2_n61), .A3(
        pe_1_7_2_n62), .ZN(pe_1_7_2_n39) );
  NAND3_X1 pe_1_7_2_U54 ( .A1(pe_1_7_2_n43), .A2(pe_1_7_2_n63), .A3(
        pe_1_7_2_n60), .ZN(pe_1_7_2_n38) );
  NAND3_X1 pe_1_7_2_U53 ( .A1(pe_1_7_2_n61), .A2(pe_1_7_2_n63), .A3(
        pe_1_7_2_n43), .ZN(pe_1_7_2_n37) );
  DFFR_X1 pe_1_7_2_int_q_acc_reg_6_ ( .D(pe_1_7_2_n78), .CK(pe_1_7_2_net3028), 
        .RN(pe_1_7_2_n71), .Q(int_data_res_7__2__6_) );
  DFFR_X1 pe_1_7_2_int_q_acc_reg_5_ ( .D(pe_1_7_2_n79), .CK(pe_1_7_2_net3028), 
        .RN(pe_1_7_2_n71), .Q(int_data_res_7__2__5_) );
  DFFR_X1 pe_1_7_2_int_q_acc_reg_4_ ( .D(pe_1_7_2_n80), .CK(pe_1_7_2_net3028), 
        .RN(pe_1_7_2_n71), .Q(int_data_res_7__2__4_) );
  DFFR_X1 pe_1_7_2_int_q_acc_reg_3_ ( .D(pe_1_7_2_n81), .CK(pe_1_7_2_net3028), 
        .RN(pe_1_7_2_n71), .Q(int_data_res_7__2__3_) );
  DFFR_X1 pe_1_7_2_int_q_acc_reg_2_ ( .D(pe_1_7_2_n82), .CK(pe_1_7_2_net3028), 
        .RN(pe_1_7_2_n71), .Q(int_data_res_7__2__2_) );
  DFFR_X1 pe_1_7_2_int_q_acc_reg_1_ ( .D(pe_1_7_2_n83), .CK(pe_1_7_2_net3028), 
        .RN(pe_1_7_2_n71), .Q(int_data_res_7__2__1_) );
  DFFR_X1 pe_1_7_2_int_q_acc_reg_7_ ( .D(pe_1_7_2_n77), .CK(pe_1_7_2_net3028), 
        .RN(pe_1_7_2_n71), .Q(int_data_res_7__2__7_) );
  CLKGATETST_X1 pe_1_7_2_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_7_2_n88), .SE(1'b0), .GCK(pe_1_7_2_net2967) );
  CLKGATETST_X1 pe_1_7_2_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_7_2_n87), .SE(1'b0), .GCK(pe_1_7_2_net2973) );
  CLKGATETST_X1 pe_1_7_2_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_7_2_n86), .SE(1'b0), .GCK(pe_1_7_2_net2978) );
  CLKGATETST_X1 pe_1_7_2_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_7_2_n85), .SE(1'b0), .GCK(pe_1_7_2_net2983) );
  CLKGATETST_X1 pe_1_7_2_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_7_2_n90), .SE(1'b0), .GCK(pe_1_7_2_net2988) );
  CLKGATETST_X1 pe_1_7_2_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_7_2_n89), .SE(1'b0), .GCK(pe_1_7_2_net2993) );
  CLKGATETST_X1 pe_1_7_2_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_7_2_N64), .SE(1'b0), .GCK(pe_1_7_2_net2998) );
  CLKGATETST_X1 pe_1_7_2_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_7_2_N63), .SE(1'b0), .GCK(pe_1_7_2_net3003) );
  CLKGATETST_X1 pe_1_7_2_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_7_2_N62), .SE(1'b0), .GCK(pe_1_7_2_net3008) );
  CLKGATETST_X1 pe_1_7_2_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_7_2_N61), .SE(1'b0), .GCK(pe_1_7_2_net3013) );
  CLKGATETST_X1 pe_1_7_2_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_7_2_N60), .SE(1'b0), .GCK(pe_1_7_2_net3018) );
  CLKGATETST_X1 pe_1_7_2_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_7_2_N59), .SE(1'b0), .GCK(pe_1_7_2_net3023) );
  CLKGATETST_X1 pe_1_7_2_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_7_2_N90), .SE(1'b0), .GCK(pe_1_7_2_net3028) );
  CLKBUF_X1 pe_1_7_3_U112 ( .A(pe_1_7_3_n72), .Z(pe_1_7_3_n71) );
  INV_X1 pe_1_7_3_U111 ( .A(n77), .ZN(pe_1_7_3_n70) );
  INV_X1 pe_1_7_3_U110 ( .A(n69), .ZN(pe_1_7_3_n69) );
  INV_X1 pe_1_7_3_U109 ( .A(n69), .ZN(pe_1_7_3_n68) );
  INV_X1 pe_1_7_3_U108 ( .A(n69), .ZN(pe_1_7_3_n67) );
  INV_X1 pe_1_7_3_U107 ( .A(pe_1_7_3_n69), .ZN(pe_1_7_3_n66) );
  INV_X1 pe_1_7_3_U106 ( .A(pe_1_7_3_n63), .ZN(pe_1_7_3_n62) );
  INV_X1 pe_1_7_3_U105 ( .A(pe_1_7_3_n61), .ZN(pe_1_7_3_n60) );
  INV_X1 pe_1_7_3_U104 ( .A(n29), .ZN(pe_1_7_3_n59) );
  INV_X1 pe_1_7_3_U103 ( .A(pe_1_7_3_n59), .ZN(pe_1_7_3_n58) );
  INV_X1 pe_1_7_3_U102 ( .A(n21), .ZN(pe_1_7_3_n57) );
  MUX2_X1 pe_1_7_3_U101 ( .A(pe_1_7_3_n54), .B(pe_1_7_3_n51), .S(n54), .Z(
        int_data_x_7__3__3_) );
  MUX2_X1 pe_1_7_3_U100 ( .A(pe_1_7_3_n53), .B(pe_1_7_3_n52), .S(pe_1_7_3_n62), 
        .Z(pe_1_7_3_n54) );
  MUX2_X1 pe_1_7_3_U99 ( .A(pe_1_7_3_int_q_reg_h[23]), .B(
        pe_1_7_3_int_q_reg_h[19]), .S(pe_1_7_3_n56), .Z(pe_1_7_3_n53) );
  MUX2_X1 pe_1_7_3_U98 ( .A(pe_1_7_3_int_q_reg_h[15]), .B(
        pe_1_7_3_int_q_reg_h[11]), .S(pe_1_7_3_n56), .Z(pe_1_7_3_n52) );
  MUX2_X1 pe_1_7_3_U97 ( .A(pe_1_7_3_int_q_reg_h[7]), .B(
        pe_1_7_3_int_q_reg_h[3]), .S(pe_1_7_3_n56), .Z(pe_1_7_3_n51) );
  MUX2_X1 pe_1_7_3_U96 ( .A(pe_1_7_3_n50), .B(pe_1_7_3_n47), .S(n54), .Z(
        int_data_x_7__3__2_) );
  MUX2_X1 pe_1_7_3_U95 ( .A(pe_1_7_3_n49), .B(pe_1_7_3_n48), .S(pe_1_7_3_n62), 
        .Z(pe_1_7_3_n50) );
  MUX2_X1 pe_1_7_3_U94 ( .A(pe_1_7_3_int_q_reg_h[22]), .B(
        pe_1_7_3_int_q_reg_h[18]), .S(pe_1_7_3_n56), .Z(pe_1_7_3_n49) );
  MUX2_X1 pe_1_7_3_U93 ( .A(pe_1_7_3_int_q_reg_h[14]), .B(
        pe_1_7_3_int_q_reg_h[10]), .S(pe_1_7_3_n56), .Z(pe_1_7_3_n48) );
  MUX2_X1 pe_1_7_3_U92 ( .A(pe_1_7_3_int_q_reg_h[6]), .B(
        pe_1_7_3_int_q_reg_h[2]), .S(pe_1_7_3_n56), .Z(pe_1_7_3_n47) );
  MUX2_X1 pe_1_7_3_U91 ( .A(pe_1_7_3_n46), .B(pe_1_7_3_n24), .S(n54), .Z(
        int_data_x_7__3__1_) );
  MUX2_X1 pe_1_7_3_U90 ( .A(pe_1_7_3_n45), .B(pe_1_7_3_n25), .S(pe_1_7_3_n62), 
        .Z(pe_1_7_3_n46) );
  MUX2_X1 pe_1_7_3_U89 ( .A(pe_1_7_3_int_q_reg_h[21]), .B(
        pe_1_7_3_int_q_reg_h[17]), .S(pe_1_7_3_n56), .Z(pe_1_7_3_n45) );
  MUX2_X1 pe_1_7_3_U88 ( .A(pe_1_7_3_int_q_reg_h[13]), .B(
        pe_1_7_3_int_q_reg_h[9]), .S(pe_1_7_3_n56), .Z(pe_1_7_3_n25) );
  MUX2_X1 pe_1_7_3_U87 ( .A(pe_1_7_3_int_q_reg_h[5]), .B(
        pe_1_7_3_int_q_reg_h[1]), .S(pe_1_7_3_n56), .Z(pe_1_7_3_n24) );
  MUX2_X1 pe_1_7_3_U86 ( .A(pe_1_7_3_n23), .B(pe_1_7_3_n20), .S(n54), .Z(
        int_data_x_7__3__0_) );
  MUX2_X1 pe_1_7_3_U85 ( .A(pe_1_7_3_n22), .B(pe_1_7_3_n21), .S(pe_1_7_3_n62), 
        .Z(pe_1_7_3_n23) );
  MUX2_X1 pe_1_7_3_U84 ( .A(pe_1_7_3_int_q_reg_h[20]), .B(
        pe_1_7_3_int_q_reg_h[16]), .S(pe_1_7_3_n56), .Z(pe_1_7_3_n22) );
  MUX2_X1 pe_1_7_3_U83 ( .A(pe_1_7_3_int_q_reg_h[12]), .B(
        pe_1_7_3_int_q_reg_h[8]), .S(pe_1_7_3_n56), .Z(pe_1_7_3_n21) );
  MUX2_X1 pe_1_7_3_U82 ( .A(pe_1_7_3_int_q_reg_h[4]), .B(
        pe_1_7_3_int_q_reg_h[0]), .S(pe_1_7_3_n56), .Z(pe_1_7_3_n20) );
  MUX2_X1 pe_1_7_3_U81 ( .A(pe_1_7_3_n19), .B(pe_1_7_3_n16), .S(n54), .Z(
        int_data_y_7__3__3_) );
  MUX2_X1 pe_1_7_3_U80 ( .A(pe_1_7_3_n18), .B(pe_1_7_3_n17), .S(pe_1_7_3_n62), 
        .Z(pe_1_7_3_n19) );
  MUX2_X1 pe_1_7_3_U79 ( .A(pe_1_7_3_int_q_reg_v[23]), .B(
        pe_1_7_3_int_q_reg_v[19]), .S(pe_1_7_3_n55), .Z(pe_1_7_3_n18) );
  MUX2_X1 pe_1_7_3_U78 ( .A(pe_1_7_3_int_q_reg_v[15]), .B(
        pe_1_7_3_int_q_reg_v[11]), .S(pe_1_7_3_n55), .Z(pe_1_7_3_n17) );
  MUX2_X1 pe_1_7_3_U77 ( .A(pe_1_7_3_int_q_reg_v[7]), .B(
        pe_1_7_3_int_q_reg_v[3]), .S(pe_1_7_3_n55), .Z(pe_1_7_3_n16) );
  MUX2_X1 pe_1_7_3_U76 ( .A(pe_1_7_3_n15), .B(pe_1_7_3_n12), .S(n54), .Z(
        int_data_y_7__3__2_) );
  MUX2_X1 pe_1_7_3_U75 ( .A(pe_1_7_3_n14), .B(pe_1_7_3_n13), .S(pe_1_7_3_n62), 
        .Z(pe_1_7_3_n15) );
  MUX2_X1 pe_1_7_3_U74 ( .A(pe_1_7_3_int_q_reg_v[22]), .B(
        pe_1_7_3_int_q_reg_v[18]), .S(pe_1_7_3_n55), .Z(pe_1_7_3_n14) );
  MUX2_X1 pe_1_7_3_U73 ( .A(pe_1_7_3_int_q_reg_v[14]), .B(
        pe_1_7_3_int_q_reg_v[10]), .S(pe_1_7_3_n55), .Z(pe_1_7_3_n13) );
  MUX2_X1 pe_1_7_3_U72 ( .A(pe_1_7_3_int_q_reg_v[6]), .B(
        pe_1_7_3_int_q_reg_v[2]), .S(pe_1_7_3_n55), .Z(pe_1_7_3_n12) );
  MUX2_X1 pe_1_7_3_U71 ( .A(pe_1_7_3_n11), .B(pe_1_7_3_n8), .S(n54), .Z(
        int_data_y_7__3__1_) );
  MUX2_X1 pe_1_7_3_U70 ( .A(pe_1_7_3_n10), .B(pe_1_7_3_n9), .S(pe_1_7_3_n62), 
        .Z(pe_1_7_3_n11) );
  MUX2_X1 pe_1_7_3_U69 ( .A(pe_1_7_3_int_q_reg_v[21]), .B(
        pe_1_7_3_int_q_reg_v[17]), .S(pe_1_7_3_n55), .Z(pe_1_7_3_n10) );
  MUX2_X1 pe_1_7_3_U68 ( .A(pe_1_7_3_int_q_reg_v[13]), .B(
        pe_1_7_3_int_q_reg_v[9]), .S(pe_1_7_3_n55), .Z(pe_1_7_3_n9) );
  MUX2_X1 pe_1_7_3_U67 ( .A(pe_1_7_3_int_q_reg_v[5]), .B(
        pe_1_7_3_int_q_reg_v[1]), .S(pe_1_7_3_n55), .Z(pe_1_7_3_n8) );
  MUX2_X1 pe_1_7_3_U66 ( .A(pe_1_7_3_n7), .B(pe_1_7_3_n4), .S(n54), .Z(
        int_data_y_7__3__0_) );
  MUX2_X1 pe_1_7_3_U65 ( .A(pe_1_7_3_n6), .B(pe_1_7_3_n5), .S(pe_1_7_3_n62), 
        .Z(pe_1_7_3_n7) );
  MUX2_X1 pe_1_7_3_U64 ( .A(pe_1_7_3_int_q_reg_v[20]), .B(
        pe_1_7_3_int_q_reg_v[16]), .S(pe_1_7_3_n55), .Z(pe_1_7_3_n6) );
  MUX2_X1 pe_1_7_3_U63 ( .A(pe_1_7_3_int_q_reg_v[12]), .B(
        pe_1_7_3_int_q_reg_v[8]), .S(pe_1_7_3_n55), .Z(pe_1_7_3_n5) );
  MUX2_X1 pe_1_7_3_U62 ( .A(pe_1_7_3_int_q_reg_v[4]), .B(
        pe_1_7_3_int_q_reg_v[0]), .S(pe_1_7_3_n55), .Z(pe_1_7_3_n4) );
  AOI222_X1 pe_1_7_3_U61 ( .A1(i_data_acc[34]), .A2(pe_1_7_3_n64), .B1(
        pe_1_7_3_N80), .B2(pe_1_7_3_n27), .C1(pe_1_7_3_N72), .C2(pe_1_7_3_n28), 
        .ZN(pe_1_7_3_n33) );
  INV_X1 pe_1_7_3_U60 ( .A(pe_1_7_3_n33), .ZN(pe_1_7_3_n82) );
  AOI222_X1 pe_1_7_3_U59 ( .A1(i_data_acc[38]), .A2(pe_1_7_3_n64), .B1(
        pe_1_7_3_N84), .B2(pe_1_7_3_n27), .C1(pe_1_7_3_N76), .C2(pe_1_7_3_n28), 
        .ZN(pe_1_7_3_n29) );
  INV_X1 pe_1_7_3_U58 ( .A(pe_1_7_3_n29), .ZN(pe_1_7_3_n78) );
  XNOR2_X1 pe_1_7_3_U57 ( .A(pe_1_7_3_n73), .B(int_data_res_7__3__0_), .ZN(
        pe_1_7_3_N70) );
  AOI222_X1 pe_1_7_3_U52 ( .A1(i_data_acc[32]), .A2(pe_1_7_3_n64), .B1(
        pe_1_7_3_n1), .B2(pe_1_7_3_n27), .C1(pe_1_7_3_N70), .C2(pe_1_7_3_n28), 
        .ZN(pe_1_7_3_n35) );
  INV_X1 pe_1_7_3_U51 ( .A(pe_1_7_3_n35), .ZN(pe_1_7_3_n84) );
  AOI222_X1 pe_1_7_3_U50 ( .A1(i_data_acc[33]), .A2(pe_1_7_3_n64), .B1(
        pe_1_7_3_N79), .B2(pe_1_7_3_n27), .C1(pe_1_7_3_N71), .C2(pe_1_7_3_n28), 
        .ZN(pe_1_7_3_n34) );
  INV_X1 pe_1_7_3_U49 ( .A(pe_1_7_3_n34), .ZN(pe_1_7_3_n83) );
  AOI222_X1 pe_1_7_3_U48 ( .A1(i_data_acc[35]), .A2(pe_1_7_3_n64), .B1(
        pe_1_7_3_N81), .B2(pe_1_7_3_n27), .C1(pe_1_7_3_N73), .C2(pe_1_7_3_n28), 
        .ZN(pe_1_7_3_n32) );
  INV_X1 pe_1_7_3_U47 ( .A(pe_1_7_3_n32), .ZN(pe_1_7_3_n81) );
  AOI222_X1 pe_1_7_3_U46 ( .A1(i_data_acc[36]), .A2(pe_1_7_3_n64), .B1(
        pe_1_7_3_N82), .B2(pe_1_7_3_n27), .C1(pe_1_7_3_N74), .C2(pe_1_7_3_n28), 
        .ZN(pe_1_7_3_n31) );
  INV_X1 pe_1_7_3_U45 ( .A(pe_1_7_3_n31), .ZN(pe_1_7_3_n80) );
  AOI222_X1 pe_1_7_3_U44 ( .A1(i_data_acc[37]), .A2(pe_1_7_3_n64), .B1(
        pe_1_7_3_N83), .B2(pe_1_7_3_n27), .C1(pe_1_7_3_N75), .C2(pe_1_7_3_n28), 
        .ZN(pe_1_7_3_n30) );
  INV_X1 pe_1_7_3_U43 ( .A(pe_1_7_3_n30), .ZN(pe_1_7_3_n79) );
  NAND2_X1 pe_1_7_3_U42 ( .A1(pe_1_7_3_int_data_0_), .A2(pe_1_7_3_n3), .ZN(
        pe_1_7_3_sub_81_carry[1]) );
  INV_X1 pe_1_7_3_U41 ( .A(pe_1_7_3_int_data_1_), .ZN(pe_1_7_3_n74) );
  INV_X1 pe_1_7_3_U40 ( .A(pe_1_7_3_int_data_2_), .ZN(pe_1_7_3_n75) );
  AND2_X1 pe_1_7_3_U39 ( .A1(pe_1_7_3_int_data_0_), .A2(int_data_res_7__3__0_), 
        .ZN(pe_1_7_3_n2) );
  AOI222_X1 pe_1_7_3_U38 ( .A1(pe_1_7_3_n64), .A2(i_data_acc[39]), .B1(
        pe_1_7_3_N85), .B2(pe_1_7_3_n27), .C1(pe_1_7_3_N77), .C2(pe_1_7_3_n28), 
        .ZN(pe_1_7_3_n26) );
  INV_X1 pe_1_7_3_U37 ( .A(pe_1_7_3_n26), .ZN(pe_1_7_3_n77) );
  NOR3_X1 pe_1_7_3_U36 ( .A1(pe_1_7_3_n59), .A2(pe_1_7_3_n65), .A3(int_ckg[4]), 
        .ZN(pe_1_7_3_n36) );
  OR2_X1 pe_1_7_3_U35 ( .A1(pe_1_7_3_n36), .A2(pe_1_7_3_n64), .ZN(pe_1_7_3_N90) );
  INV_X1 pe_1_7_3_U34 ( .A(n41), .ZN(pe_1_7_3_n63) );
  AND2_X1 pe_1_7_3_U33 ( .A1(int_data_x_7__3__2_), .A2(pe_1_7_3_n58), .ZN(
        pe_1_7_3_int_data_2_) );
  AND2_X1 pe_1_7_3_U32 ( .A1(int_data_x_7__3__1_), .A2(pe_1_7_3_n58), .ZN(
        pe_1_7_3_int_data_1_) );
  AND2_X1 pe_1_7_3_U31 ( .A1(int_data_x_7__3__3_), .A2(pe_1_7_3_n58), .ZN(
        pe_1_7_3_int_data_3_) );
  BUF_X1 pe_1_7_3_U30 ( .A(n63), .Z(pe_1_7_3_n64) );
  INV_X1 pe_1_7_3_U29 ( .A(n35), .ZN(pe_1_7_3_n61) );
  AND2_X1 pe_1_7_3_U28 ( .A1(int_data_x_7__3__0_), .A2(pe_1_7_3_n58), .ZN(
        pe_1_7_3_int_data_0_) );
  NAND2_X1 pe_1_7_3_U27 ( .A1(pe_1_7_3_n44), .A2(pe_1_7_3_n61), .ZN(
        pe_1_7_3_n41) );
  AND3_X1 pe_1_7_3_U26 ( .A1(n77), .A2(pe_1_7_3_n63), .A3(n54), .ZN(
        pe_1_7_3_n44) );
  INV_X1 pe_1_7_3_U25 ( .A(pe_1_7_3_int_data_3_), .ZN(pe_1_7_3_n76) );
  NOR2_X1 pe_1_7_3_U24 ( .A1(pe_1_7_3_n70), .A2(n54), .ZN(pe_1_7_3_n43) );
  NOR2_X1 pe_1_7_3_U23 ( .A1(pe_1_7_3_n57), .A2(pe_1_7_3_n64), .ZN(
        pe_1_7_3_n28) );
  NOR2_X1 pe_1_7_3_U22 ( .A1(n21), .A2(pe_1_7_3_n64), .ZN(pe_1_7_3_n27) );
  INV_X1 pe_1_7_3_U21 ( .A(pe_1_7_3_int_data_0_), .ZN(pe_1_7_3_n73) );
  INV_X1 pe_1_7_3_U20 ( .A(pe_1_7_3_n41), .ZN(pe_1_7_3_n90) );
  INV_X1 pe_1_7_3_U19 ( .A(pe_1_7_3_n37), .ZN(pe_1_7_3_n88) );
  INV_X1 pe_1_7_3_U18 ( .A(pe_1_7_3_n38), .ZN(pe_1_7_3_n87) );
  INV_X1 pe_1_7_3_U17 ( .A(pe_1_7_3_n39), .ZN(pe_1_7_3_n86) );
  NOR2_X1 pe_1_7_3_U16 ( .A1(pe_1_7_3_n68), .A2(pe_1_7_3_n42), .ZN(
        pe_1_7_3_N59) );
  NOR2_X1 pe_1_7_3_U15 ( .A1(pe_1_7_3_n68), .A2(pe_1_7_3_n41), .ZN(
        pe_1_7_3_N60) );
  NOR2_X1 pe_1_7_3_U14 ( .A1(pe_1_7_3_n68), .A2(pe_1_7_3_n38), .ZN(
        pe_1_7_3_N63) );
  NOR2_X1 pe_1_7_3_U13 ( .A1(pe_1_7_3_n67), .A2(pe_1_7_3_n40), .ZN(
        pe_1_7_3_N61) );
  NOR2_X1 pe_1_7_3_U12 ( .A1(pe_1_7_3_n67), .A2(pe_1_7_3_n39), .ZN(
        pe_1_7_3_N62) );
  NOR2_X1 pe_1_7_3_U11 ( .A1(pe_1_7_3_n37), .A2(pe_1_7_3_n67), .ZN(
        pe_1_7_3_N64) );
  NAND2_X1 pe_1_7_3_U10 ( .A1(pe_1_7_3_n44), .A2(pe_1_7_3_n60), .ZN(
        pe_1_7_3_n42) );
  BUF_X1 pe_1_7_3_U9 ( .A(pe_1_7_3_n60), .Z(pe_1_7_3_n55) );
  INV_X1 pe_1_7_3_U8 ( .A(pe_1_7_3_n69), .ZN(pe_1_7_3_n65) );
  BUF_X1 pe_1_7_3_U7 ( .A(pe_1_7_3_n60), .Z(pe_1_7_3_n56) );
  INV_X1 pe_1_7_3_U6 ( .A(pe_1_7_3_n42), .ZN(pe_1_7_3_n89) );
  INV_X1 pe_1_7_3_U5 ( .A(pe_1_7_3_n40), .ZN(pe_1_7_3_n85) );
  INV_X2 pe_1_7_3_U4 ( .A(n85), .ZN(pe_1_7_3_n72) );
  XOR2_X1 pe_1_7_3_U3 ( .A(pe_1_7_3_int_data_0_), .B(int_data_res_7__3__0_), 
        .Z(pe_1_7_3_n1) );
  DFFR_X1 pe_1_7_3_int_q_acc_reg_0_ ( .D(pe_1_7_3_n84), .CK(pe_1_7_3_net2950), 
        .RN(pe_1_7_3_n72), .Q(int_data_res_7__3__0_), .QN(pe_1_7_3_n3) );
  DFFR_X1 pe_1_7_3_int_q_reg_v_reg_0__0_ ( .D(i_data_conv_v[16]), .CK(
        pe_1_7_3_net2920), .RN(pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_v[20]) );
  DFFR_X1 pe_1_7_3_int_q_reg_v_reg_0__1_ ( .D(i_data_conv_v[17]), .CK(
        pe_1_7_3_net2920), .RN(pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_v[21]) );
  DFFR_X1 pe_1_7_3_int_q_reg_v_reg_0__2_ ( .D(i_data_conv_v[18]), .CK(
        pe_1_7_3_net2920), .RN(pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_v[22]) );
  DFFR_X1 pe_1_7_3_int_q_reg_v_reg_0__3_ ( .D(i_data_conv_v[19]), .CK(
        pe_1_7_3_net2920), .RN(pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_v[23]) );
  DFFR_X1 pe_1_7_3_int_q_reg_v_reg_1__0_ ( .D(i_data_conv_v[16]), .CK(
        pe_1_7_3_net2925), .RN(pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_v[16]) );
  DFFR_X1 pe_1_7_3_int_q_reg_v_reg_1__1_ ( .D(i_data_conv_v[17]), .CK(
        pe_1_7_3_net2925), .RN(pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_v[17]) );
  DFFR_X1 pe_1_7_3_int_q_reg_v_reg_1__2_ ( .D(i_data_conv_v[18]), .CK(
        pe_1_7_3_net2925), .RN(pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_v[18]) );
  DFFR_X1 pe_1_7_3_int_q_reg_v_reg_1__3_ ( .D(i_data_conv_v[19]), .CK(
        pe_1_7_3_net2925), .RN(pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_v[19]) );
  DFFR_X1 pe_1_7_3_int_q_reg_v_reg_2__0_ ( .D(i_data_conv_v[16]), .CK(
        pe_1_7_3_net2930), .RN(pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_v[12]) );
  DFFR_X1 pe_1_7_3_int_q_reg_v_reg_2__1_ ( .D(i_data_conv_v[17]), .CK(
        pe_1_7_3_net2930), .RN(pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_v[13]) );
  DFFR_X1 pe_1_7_3_int_q_reg_v_reg_2__2_ ( .D(i_data_conv_v[18]), .CK(
        pe_1_7_3_net2930), .RN(pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_v[14]) );
  DFFR_X1 pe_1_7_3_int_q_reg_v_reg_2__3_ ( .D(i_data_conv_v[19]), .CK(
        pe_1_7_3_net2930), .RN(pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_v[15]) );
  DFFR_X1 pe_1_7_3_int_q_reg_v_reg_3__0_ ( .D(i_data_conv_v[16]), .CK(
        pe_1_7_3_net2935), .RN(pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_v[8]) );
  DFFR_X1 pe_1_7_3_int_q_reg_v_reg_3__1_ ( .D(i_data_conv_v[17]), .CK(
        pe_1_7_3_net2935), .RN(pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_v[9]) );
  DFFR_X1 pe_1_7_3_int_q_reg_v_reg_3__2_ ( .D(i_data_conv_v[18]), .CK(
        pe_1_7_3_net2935), .RN(pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_v[10]) );
  DFFR_X1 pe_1_7_3_int_q_reg_v_reg_3__3_ ( .D(i_data_conv_v[19]), .CK(
        pe_1_7_3_net2935), .RN(pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_v[11]) );
  DFFR_X1 pe_1_7_3_int_q_reg_v_reg_4__0_ ( .D(i_data_conv_v[16]), .CK(
        pe_1_7_3_net2940), .RN(pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_v[4]) );
  DFFR_X1 pe_1_7_3_int_q_reg_v_reg_4__1_ ( .D(i_data_conv_v[17]), .CK(
        pe_1_7_3_net2940), .RN(pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_v[5]) );
  DFFR_X1 pe_1_7_3_int_q_reg_v_reg_4__2_ ( .D(i_data_conv_v[18]), .CK(
        pe_1_7_3_net2940), .RN(pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_v[6]) );
  DFFR_X1 pe_1_7_3_int_q_reg_v_reg_4__3_ ( .D(i_data_conv_v[19]), .CK(
        pe_1_7_3_net2940), .RN(pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_v[7]) );
  DFFR_X1 pe_1_7_3_int_q_reg_v_reg_5__0_ ( .D(i_data_conv_v[16]), .CK(
        pe_1_7_3_net2945), .RN(pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_v[0]) );
  DFFR_X1 pe_1_7_3_int_q_reg_v_reg_5__1_ ( .D(i_data_conv_v[17]), .CK(
        pe_1_7_3_net2945), .RN(pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_v[1]) );
  DFFR_X1 pe_1_7_3_int_q_reg_v_reg_5__2_ ( .D(i_data_conv_v[18]), .CK(
        pe_1_7_3_net2945), .RN(pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_v[2]) );
  DFFR_X1 pe_1_7_3_int_q_reg_v_reg_5__3_ ( .D(i_data_conv_v[19]), .CK(
        pe_1_7_3_net2945), .RN(pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_7_3_int_q_reg_h_reg_0__0_ ( .D(int_data_x_7__4__0_), .SI(
        i_data_conv_v[16]), .SE(pe_1_7_3_n65), .CK(pe_1_7_3_net2889), .RN(
        pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_7_3_int_q_reg_h_reg_0__1_ ( .D(int_data_x_7__4__1_), .SI(
        i_data_conv_v[17]), .SE(pe_1_7_3_n65), .CK(pe_1_7_3_net2889), .RN(
        pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_7_3_int_q_reg_h_reg_0__2_ ( .D(int_data_x_7__4__2_), .SI(
        i_data_conv_v[18]), .SE(pe_1_7_3_n65), .CK(pe_1_7_3_net2889), .RN(
        pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_7_3_int_q_reg_h_reg_0__3_ ( .D(int_data_x_7__4__3_), .SI(
        i_data_conv_v[19]), .SE(pe_1_7_3_n65), .CK(pe_1_7_3_net2889), .RN(
        pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_7_3_int_q_reg_h_reg_1__0_ ( .D(int_data_x_7__4__0_), .SI(
        i_data_conv_v[16]), .SE(pe_1_7_3_n65), .CK(pe_1_7_3_net2895), .RN(
        pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_7_3_int_q_reg_h_reg_1__1_ ( .D(int_data_x_7__4__1_), .SI(
        i_data_conv_v[17]), .SE(pe_1_7_3_n65), .CK(pe_1_7_3_net2895), .RN(
        pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_7_3_int_q_reg_h_reg_1__2_ ( .D(int_data_x_7__4__2_), .SI(
        i_data_conv_v[18]), .SE(pe_1_7_3_n65), .CK(pe_1_7_3_net2895), .RN(
        pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_7_3_int_q_reg_h_reg_1__3_ ( .D(int_data_x_7__4__3_), .SI(
        i_data_conv_v[19]), .SE(pe_1_7_3_n65), .CK(pe_1_7_3_net2895), .RN(
        pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_7_3_int_q_reg_h_reg_2__0_ ( .D(int_data_x_7__4__0_), .SI(
        i_data_conv_v[16]), .SE(pe_1_7_3_n65), .CK(pe_1_7_3_net2900), .RN(
        pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_7_3_int_q_reg_h_reg_2__1_ ( .D(int_data_x_7__4__1_), .SI(
        i_data_conv_v[17]), .SE(pe_1_7_3_n65), .CK(pe_1_7_3_net2900), .RN(
        pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_7_3_int_q_reg_h_reg_2__2_ ( .D(int_data_x_7__4__2_), .SI(
        i_data_conv_v[18]), .SE(pe_1_7_3_n65), .CK(pe_1_7_3_net2900), .RN(
        pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_7_3_int_q_reg_h_reg_2__3_ ( .D(int_data_x_7__4__3_), .SI(
        i_data_conv_v[19]), .SE(pe_1_7_3_n65), .CK(pe_1_7_3_net2900), .RN(
        pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_7_3_int_q_reg_h_reg_3__0_ ( .D(int_data_x_7__4__0_), .SI(
        i_data_conv_v[16]), .SE(pe_1_7_3_n65), .CK(pe_1_7_3_net2905), .RN(
        pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_7_3_int_q_reg_h_reg_3__1_ ( .D(int_data_x_7__4__1_), .SI(
        i_data_conv_v[17]), .SE(pe_1_7_3_n65), .CK(pe_1_7_3_net2905), .RN(
        pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_7_3_int_q_reg_h_reg_3__2_ ( .D(int_data_x_7__4__2_), .SI(
        i_data_conv_v[18]), .SE(pe_1_7_3_n65), .CK(pe_1_7_3_net2905), .RN(
        pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_7_3_int_q_reg_h_reg_3__3_ ( .D(int_data_x_7__4__3_), .SI(
        i_data_conv_v[19]), .SE(pe_1_7_3_n65), .CK(pe_1_7_3_net2905), .RN(
        pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_7_3_int_q_reg_h_reg_4__0_ ( .D(int_data_x_7__4__0_), .SI(
        i_data_conv_v[16]), .SE(pe_1_7_3_n66), .CK(pe_1_7_3_net2910), .RN(
        pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_7_3_int_q_reg_h_reg_4__1_ ( .D(int_data_x_7__4__1_), .SI(
        i_data_conv_v[17]), .SE(pe_1_7_3_n66), .CK(pe_1_7_3_net2910), .RN(
        pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_7_3_int_q_reg_h_reg_4__2_ ( .D(int_data_x_7__4__2_), .SI(
        i_data_conv_v[18]), .SE(pe_1_7_3_n66), .CK(pe_1_7_3_net2910), .RN(
        pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_7_3_int_q_reg_h_reg_4__3_ ( .D(int_data_x_7__4__3_), .SI(
        i_data_conv_v[19]), .SE(pe_1_7_3_n66), .CK(pe_1_7_3_net2910), .RN(
        pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_7_3_int_q_reg_h_reg_5__0_ ( .D(int_data_x_7__4__0_), .SI(
        i_data_conv_v[16]), .SE(pe_1_7_3_n66), .CK(pe_1_7_3_net2915), .RN(
        pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_7_3_int_q_reg_h_reg_5__1_ ( .D(int_data_x_7__4__1_), .SI(
        i_data_conv_v[17]), .SE(pe_1_7_3_n66), .CK(pe_1_7_3_net2915), .RN(
        pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_7_3_int_q_reg_h_reg_5__2_ ( .D(int_data_x_7__4__2_), .SI(
        i_data_conv_v[18]), .SE(pe_1_7_3_n66), .CK(pe_1_7_3_net2915), .RN(
        pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_7_3_int_q_reg_h_reg_5__3_ ( .D(int_data_x_7__4__3_), .SI(
        i_data_conv_v[19]), .SE(pe_1_7_3_n66), .CK(pe_1_7_3_net2915), .RN(
        pe_1_7_3_n72), .Q(pe_1_7_3_int_q_reg_h[3]) );
  FA_X1 pe_1_7_3_sub_81_U2_7 ( .A(int_data_res_7__3__7_), .B(pe_1_7_3_n76), 
        .CI(pe_1_7_3_sub_81_carry[7]), .S(pe_1_7_3_N77) );
  FA_X1 pe_1_7_3_sub_81_U2_6 ( .A(int_data_res_7__3__6_), .B(pe_1_7_3_n76), 
        .CI(pe_1_7_3_sub_81_carry[6]), .CO(pe_1_7_3_sub_81_carry[7]), .S(
        pe_1_7_3_N76) );
  FA_X1 pe_1_7_3_sub_81_U2_5 ( .A(int_data_res_7__3__5_), .B(pe_1_7_3_n76), 
        .CI(pe_1_7_3_sub_81_carry[5]), .CO(pe_1_7_3_sub_81_carry[6]), .S(
        pe_1_7_3_N75) );
  FA_X1 pe_1_7_3_sub_81_U2_4 ( .A(int_data_res_7__3__4_), .B(pe_1_7_3_n76), 
        .CI(pe_1_7_3_sub_81_carry[4]), .CO(pe_1_7_3_sub_81_carry[5]), .S(
        pe_1_7_3_N74) );
  FA_X1 pe_1_7_3_sub_81_U2_3 ( .A(int_data_res_7__3__3_), .B(pe_1_7_3_n76), 
        .CI(pe_1_7_3_sub_81_carry[3]), .CO(pe_1_7_3_sub_81_carry[4]), .S(
        pe_1_7_3_N73) );
  FA_X1 pe_1_7_3_sub_81_U2_2 ( .A(int_data_res_7__3__2_), .B(pe_1_7_3_n75), 
        .CI(pe_1_7_3_sub_81_carry[2]), .CO(pe_1_7_3_sub_81_carry[3]), .S(
        pe_1_7_3_N72) );
  FA_X1 pe_1_7_3_sub_81_U2_1 ( .A(int_data_res_7__3__1_), .B(pe_1_7_3_n74), 
        .CI(pe_1_7_3_sub_81_carry[1]), .CO(pe_1_7_3_sub_81_carry[2]), .S(
        pe_1_7_3_N71) );
  FA_X1 pe_1_7_3_add_83_U1_7 ( .A(int_data_res_7__3__7_), .B(
        pe_1_7_3_int_data_3_), .CI(pe_1_7_3_add_83_carry[7]), .S(pe_1_7_3_N85)
         );
  FA_X1 pe_1_7_3_add_83_U1_6 ( .A(int_data_res_7__3__6_), .B(
        pe_1_7_3_int_data_3_), .CI(pe_1_7_3_add_83_carry[6]), .CO(
        pe_1_7_3_add_83_carry[7]), .S(pe_1_7_3_N84) );
  FA_X1 pe_1_7_3_add_83_U1_5 ( .A(int_data_res_7__3__5_), .B(
        pe_1_7_3_int_data_3_), .CI(pe_1_7_3_add_83_carry[5]), .CO(
        pe_1_7_3_add_83_carry[6]), .S(pe_1_7_3_N83) );
  FA_X1 pe_1_7_3_add_83_U1_4 ( .A(int_data_res_7__3__4_), .B(
        pe_1_7_3_int_data_3_), .CI(pe_1_7_3_add_83_carry[4]), .CO(
        pe_1_7_3_add_83_carry[5]), .S(pe_1_7_3_N82) );
  FA_X1 pe_1_7_3_add_83_U1_3 ( .A(int_data_res_7__3__3_), .B(
        pe_1_7_3_int_data_3_), .CI(pe_1_7_3_add_83_carry[3]), .CO(
        pe_1_7_3_add_83_carry[4]), .S(pe_1_7_3_N81) );
  FA_X1 pe_1_7_3_add_83_U1_2 ( .A(int_data_res_7__3__2_), .B(
        pe_1_7_3_int_data_2_), .CI(pe_1_7_3_add_83_carry[2]), .CO(
        pe_1_7_3_add_83_carry[3]), .S(pe_1_7_3_N80) );
  FA_X1 pe_1_7_3_add_83_U1_1 ( .A(int_data_res_7__3__1_), .B(
        pe_1_7_3_int_data_1_), .CI(pe_1_7_3_n2), .CO(pe_1_7_3_add_83_carry[2]), 
        .S(pe_1_7_3_N79) );
  NAND3_X1 pe_1_7_3_U56 ( .A1(pe_1_7_3_n60), .A2(pe_1_7_3_n43), .A3(
        pe_1_7_3_n62), .ZN(pe_1_7_3_n40) );
  NAND3_X1 pe_1_7_3_U55 ( .A1(pe_1_7_3_n43), .A2(pe_1_7_3_n61), .A3(
        pe_1_7_3_n62), .ZN(pe_1_7_3_n39) );
  NAND3_X1 pe_1_7_3_U54 ( .A1(pe_1_7_3_n43), .A2(pe_1_7_3_n63), .A3(
        pe_1_7_3_n60), .ZN(pe_1_7_3_n38) );
  NAND3_X1 pe_1_7_3_U53 ( .A1(pe_1_7_3_n61), .A2(pe_1_7_3_n63), .A3(
        pe_1_7_3_n43), .ZN(pe_1_7_3_n37) );
  DFFR_X1 pe_1_7_3_int_q_acc_reg_6_ ( .D(pe_1_7_3_n78), .CK(pe_1_7_3_net2950), 
        .RN(pe_1_7_3_n71), .Q(int_data_res_7__3__6_) );
  DFFR_X1 pe_1_7_3_int_q_acc_reg_5_ ( .D(pe_1_7_3_n79), .CK(pe_1_7_3_net2950), 
        .RN(pe_1_7_3_n71), .Q(int_data_res_7__3__5_) );
  DFFR_X1 pe_1_7_3_int_q_acc_reg_4_ ( .D(pe_1_7_3_n80), .CK(pe_1_7_3_net2950), 
        .RN(pe_1_7_3_n71), .Q(int_data_res_7__3__4_) );
  DFFR_X1 pe_1_7_3_int_q_acc_reg_3_ ( .D(pe_1_7_3_n81), .CK(pe_1_7_3_net2950), 
        .RN(pe_1_7_3_n71), .Q(int_data_res_7__3__3_) );
  DFFR_X1 pe_1_7_3_int_q_acc_reg_2_ ( .D(pe_1_7_3_n82), .CK(pe_1_7_3_net2950), 
        .RN(pe_1_7_3_n71), .Q(int_data_res_7__3__2_) );
  DFFR_X1 pe_1_7_3_int_q_acc_reg_1_ ( .D(pe_1_7_3_n83), .CK(pe_1_7_3_net2950), 
        .RN(pe_1_7_3_n71), .Q(int_data_res_7__3__1_) );
  DFFR_X1 pe_1_7_3_int_q_acc_reg_7_ ( .D(pe_1_7_3_n77), .CK(pe_1_7_3_net2950), 
        .RN(pe_1_7_3_n71), .Q(int_data_res_7__3__7_) );
  CLKGATETST_X1 pe_1_7_3_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_7_3_n88), .SE(1'b0), .GCK(pe_1_7_3_net2889) );
  CLKGATETST_X1 pe_1_7_3_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_7_3_n87), .SE(1'b0), .GCK(pe_1_7_3_net2895) );
  CLKGATETST_X1 pe_1_7_3_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_7_3_n86), .SE(1'b0), .GCK(pe_1_7_3_net2900) );
  CLKGATETST_X1 pe_1_7_3_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_7_3_n85), .SE(1'b0), .GCK(pe_1_7_3_net2905) );
  CLKGATETST_X1 pe_1_7_3_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_7_3_n90), .SE(1'b0), .GCK(pe_1_7_3_net2910) );
  CLKGATETST_X1 pe_1_7_3_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_7_3_n89), .SE(1'b0), .GCK(pe_1_7_3_net2915) );
  CLKGATETST_X1 pe_1_7_3_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_7_3_N64), .SE(1'b0), .GCK(pe_1_7_3_net2920) );
  CLKGATETST_X1 pe_1_7_3_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_7_3_N63), .SE(1'b0), .GCK(pe_1_7_3_net2925) );
  CLKGATETST_X1 pe_1_7_3_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_7_3_N62), .SE(1'b0), .GCK(pe_1_7_3_net2930) );
  CLKGATETST_X1 pe_1_7_3_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_7_3_N61), .SE(1'b0), .GCK(pe_1_7_3_net2935) );
  CLKGATETST_X1 pe_1_7_3_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_7_3_N60), .SE(1'b0), .GCK(pe_1_7_3_net2940) );
  CLKGATETST_X1 pe_1_7_3_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_7_3_N59), .SE(1'b0), .GCK(pe_1_7_3_net2945) );
  CLKGATETST_X1 pe_1_7_3_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_7_3_N90), .SE(1'b0), .GCK(pe_1_7_3_net2950) );
  CLKBUF_X1 pe_1_7_4_U106 ( .A(pe_1_7_4_n66), .Z(pe_1_7_4_n65) );
  INV_X1 pe_1_7_4_U105 ( .A(n78), .ZN(pe_1_7_4_n64) );
  INV_X1 pe_1_7_4_U104 ( .A(n70), .ZN(pe_1_7_4_n63) );
  INV_X1 pe_1_7_4_U103 ( .A(n30), .ZN(pe_1_7_4_n58) );
  INV_X1 pe_1_7_4_U102 ( .A(n22), .ZN(pe_1_7_4_n57) );
  MUX2_X1 pe_1_7_4_U101 ( .A(pe_1_7_4_n54), .B(pe_1_7_4_n51), .S(n55), .Z(
        int_data_x_7__4__3_) );
  MUX2_X1 pe_1_7_4_U100 ( .A(pe_1_7_4_n53), .B(pe_1_7_4_n52), .S(n42), .Z(
        pe_1_7_4_n54) );
  MUX2_X1 pe_1_7_4_U99 ( .A(pe_1_7_4_int_q_reg_h[23]), .B(
        pe_1_7_4_int_q_reg_h[19]), .S(pe_1_7_4_n56), .Z(pe_1_7_4_n53) );
  MUX2_X1 pe_1_7_4_U98 ( .A(pe_1_7_4_int_q_reg_h[15]), .B(
        pe_1_7_4_int_q_reg_h[11]), .S(pe_1_7_4_n56), .Z(pe_1_7_4_n52) );
  MUX2_X1 pe_1_7_4_U97 ( .A(pe_1_7_4_int_q_reg_h[7]), .B(
        pe_1_7_4_int_q_reg_h[3]), .S(pe_1_7_4_n56), .Z(pe_1_7_4_n51) );
  MUX2_X1 pe_1_7_4_U96 ( .A(pe_1_7_4_n50), .B(pe_1_7_4_n47), .S(n55), .Z(
        int_data_x_7__4__2_) );
  MUX2_X1 pe_1_7_4_U95 ( .A(pe_1_7_4_n49), .B(pe_1_7_4_n48), .S(n42), .Z(
        pe_1_7_4_n50) );
  MUX2_X1 pe_1_7_4_U94 ( .A(pe_1_7_4_int_q_reg_h[22]), .B(
        pe_1_7_4_int_q_reg_h[18]), .S(pe_1_7_4_n56), .Z(pe_1_7_4_n49) );
  MUX2_X1 pe_1_7_4_U93 ( .A(pe_1_7_4_int_q_reg_h[14]), .B(
        pe_1_7_4_int_q_reg_h[10]), .S(pe_1_7_4_n56), .Z(pe_1_7_4_n48) );
  MUX2_X1 pe_1_7_4_U92 ( .A(pe_1_7_4_int_q_reg_h[6]), .B(
        pe_1_7_4_int_q_reg_h[2]), .S(pe_1_7_4_n56), .Z(pe_1_7_4_n47) );
  MUX2_X1 pe_1_7_4_U91 ( .A(pe_1_7_4_n46), .B(pe_1_7_4_n24), .S(n55), .Z(
        int_data_x_7__4__1_) );
  MUX2_X1 pe_1_7_4_U90 ( .A(pe_1_7_4_n45), .B(pe_1_7_4_n25), .S(n42), .Z(
        pe_1_7_4_n46) );
  MUX2_X1 pe_1_7_4_U89 ( .A(pe_1_7_4_int_q_reg_h[21]), .B(
        pe_1_7_4_int_q_reg_h[17]), .S(pe_1_7_4_n56), .Z(pe_1_7_4_n45) );
  MUX2_X1 pe_1_7_4_U88 ( .A(pe_1_7_4_int_q_reg_h[13]), .B(
        pe_1_7_4_int_q_reg_h[9]), .S(pe_1_7_4_n56), .Z(pe_1_7_4_n25) );
  MUX2_X1 pe_1_7_4_U87 ( .A(pe_1_7_4_int_q_reg_h[5]), .B(
        pe_1_7_4_int_q_reg_h[1]), .S(pe_1_7_4_n56), .Z(pe_1_7_4_n24) );
  MUX2_X1 pe_1_7_4_U86 ( .A(pe_1_7_4_n23), .B(pe_1_7_4_n20), .S(n55), .Z(
        int_data_x_7__4__0_) );
  MUX2_X1 pe_1_7_4_U85 ( .A(pe_1_7_4_n22), .B(pe_1_7_4_n21), .S(n42), .Z(
        pe_1_7_4_n23) );
  MUX2_X1 pe_1_7_4_U84 ( .A(pe_1_7_4_int_q_reg_h[20]), .B(
        pe_1_7_4_int_q_reg_h[16]), .S(pe_1_7_4_n56), .Z(pe_1_7_4_n22) );
  MUX2_X1 pe_1_7_4_U83 ( .A(pe_1_7_4_int_q_reg_h[12]), .B(
        pe_1_7_4_int_q_reg_h[8]), .S(pe_1_7_4_n56), .Z(pe_1_7_4_n21) );
  MUX2_X1 pe_1_7_4_U82 ( .A(pe_1_7_4_int_q_reg_h[4]), .B(
        pe_1_7_4_int_q_reg_h[0]), .S(pe_1_7_4_n56), .Z(pe_1_7_4_n20) );
  MUX2_X1 pe_1_7_4_U81 ( .A(pe_1_7_4_n19), .B(pe_1_7_4_n16), .S(n55), .Z(
        int_data_y_7__4__3_) );
  MUX2_X1 pe_1_7_4_U80 ( .A(pe_1_7_4_n18), .B(pe_1_7_4_n17), .S(n42), .Z(
        pe_1_7_4_n19) );
  MUX2_X1 pe_1_7_4_U79 ( .A(pe_1_7_4_int_q_reg_v[23]), .B(
        pe_1_7_4_int_q_reg_v[19]), .S(pe_1_7_4_n55), .Z(pe_1_7_4_n18) );
  MUX2_X1 pe_1_7_4_U78 ( .A(pe_1_7_4_int_q_reg_v[15]), .B(
        pe_1_7_4_int_q_reg_v[11]), .S(pe_1_7_4_n55), .Z(pe_1_7_4_n17) );
  MUX2_X1 pe_1_7_4_U77 ( .A(pe_1_7_4_int_q_reg_v[7]), .B(
        pe_1_7_4_int_q_reg_v[3]), .S(pe_1_7_4_n55), .Z(pe_1_7_4_n16) );
  MUX2_X1 pe_1_7_4_U76 ( .A(pe_1_7_4_n15), .B(pe_1_7_4_n12), .S(n55), .Z(
        int_data_y_7__4__2_) );
  MUX2_X1 pe_1_7_4_U75 ( .A(pe_1_7_4_n14), .B(pe_1_7_4_n13), .S(n42), .Z(
        pe_1_7_4_n15) );
  MUX2_X1 pe_1_7_4_U74 ( .A(pe_1_7_4_int_q_reg_v[22]), .B(
        pe_1_7_4_int_q_reg_v[18]), .S(pe_1_7_4_n55), .Z(pe_1_7_4_n14) );
  MUX2_X1 pe_1_7_4_U73 ( .A(pe_1_7_4_int_q_reg_v[14]), .B(
        pe_1_7_4_int_q_reg_v[10]), .S(pe_1_7_4_n55), .Z(pe_1_7_4_n13) );
  MUX2_X1 pe_1_7_4_U72 ( .A(pe_1_7_4_int_q_reg_v[6]), .B(
        pe_1_7_4_int_q_reg_v[2]), .S(pe_1_7_4_n55), .Z(pe_1_7_4_n12) );
  MUX2_X1 pe_1_7_4_U71 ( .A(pe_1_7_4_n11), .B(pe_1_7_4_n8), .S(n55), .Z(
        int_data_y_7__4__1_) );
  MUX2_X1 pe_1_7_4_U70 ( .A(pe_1_7_4_n10), .B(pe_1_7_4_n9), .S(n42), .Z(
        pe_1_7_4_n11) );
  MUX2_X1 pe_1_7_4_U69 ( .A(pe_1_7_4_int_q_reg_v[21]), .B(
        pe_1_7_4_int_q_reg_v[17]), .S(pe_1_7_4_n55), .Z(pe_1_7_4_n10) );
  MUX2_X1 pe_1_7_4_U68 ( .A(pe_1_7_4_int_q_reg_v[13]), .B(
        pe_1_7_4_int_q_reg_v[9]), .S(pe_1_7_4_n55), .Z(pe_1_7_4_n9) );
  MUX2_X1 pe_1_7_4_U67 ( .A(pe_1_7_4_int_q_reg_v[5]), .B(
        pe_1_7_4_int_q_reg_v[1]), .S(pe_1_7_4_n55), .Z(pe_1_7_4_n8) );
  MUX2_X1 pe_1_7_4_U66 ( .A(pe_1_7_4_n7), .B(pe_1_7_4_n4), .S(n55), .Z(
        int_data_y_7__4__0_) );
  MUX2_X1 pe_1_7_4_U65 ( .A(pe_1_7_4_n6), .B(pe_1_7_4_n5), .S(n42), .Z(
        pe_1_7_4_n7) );
  MUX2_X1 pe_1_7_4_U64 ( .A(pe_1_7_4_int_q_reg_v[20]), .B(
        pe_1_7_4_int_q_reg_v[16]), .S(pe_1_7_4_n55), .Z(pe_1_7_4_n6) );
  MUX2_X1 pe_1_7_4_U63 ( .A(pe_1_7_4_int_q_reg_v[12]), .B(
        pe_1_7_4_int_q_reg_v[8]), .S(pe_1_7_4_n55), .Z(pe_1_7_4_n5) );
  MUX2_X1 pe_1_7_4_U62 ( .A(pe_1_7_4_int_q_reg_v[4]), .B(
        pe_1_7_4_int_q_reg_v[0]), .S(pe_1_7_4_n55), .Z(pe_1_7_4_n4) );
  AOI222_X1 pe_1_7_4_U61 ( .A1(i_data_acc[25]), .A2(pe_1_7_4_n61), .B1(
        pe_1_7_4_N79), .B2(pe_1_7_4_n27), .C1(pe_1_7_4_N71), .C2(pe_1_7_4_n28), 
        .ZN(pe_1_7_4_n34) );
  INV_X1 pe_1_7_4_U60 ( .A(pe_1_7_4_n34), .ZN(pe_1_7_4_n77) );
  AOI222_X1 pe_1_7_4_U59 ( .A1(i_data_acc[26]), .A2(pe_1_7_4_n61), .B1(
        pe_1_7_4_N80), .B2(pe_1_7_4_n27), .C1(pe_1_7_4_N72), .C2(pe_1_7_4_n28), 
        .ZN(pe_1_7_4_n33) );
  INV_X1 pe_1_7_4_U58 ( .A(pe_1_7_4_n33), .ZN(pe_1_7_4_n76) );
  AOI222_X1 pe_1_7_4_U57 ( .A1(i_data_acc[27]), .A2(pe_1_7_4_n61), .B1(
        pe_1_7_4_N81), .B2(pe_1_7_4_n27), .C1(pe_1_7_4_N73), .C2(pe_1_7_4_n28), 
        .ZN(pe_1_7_4_n32) );
  INV_X1 pe_1_7_4_U52 ( .A(pe_1_7_4_n32), .ZN(pe_1_7_4_n75) );
  AOI222_X1 pe_1_7_4_U51 ( .A1(i_data_acc[28]), .A2(pe_1_7_4_n61), .B1(
        pe_1_7_4_N82), .B2(pe_1_7_4_n27), .C1(pe_1_7_4_N74), .C2(pe_1_7_4_n28), 
        .ZN(pe_1_7_4_n31) );
  INV_X1 pe_1_7_4_U50 ( .A(pe_1_7_4_n31), .ZN(pe_1_7_4_n74) );
  AOI222_X1 pe_1_7_4_U49 ( .A1(i_data_acc[29]), .A2(pe_1_7_4_n61), .B1(
        pe_1_7_4_N83), .B2(pe_1_7_4_n27), .C1(pe_1_7_4_N75), .C2(pe_1_7_4_n28), 
        .ZN(pe_1_7_4_n30) );
  INV_X1 pe_1_7_4_U48 ( .A(pe_1_7_4_n30), .ZN(pe_1_7_4_n73) );
  AOI222_X1 pe_1_7_4_U47 ( .A1(i_data_acc[30]), .A2(pe_1_7_4_n61), .B1(
        pe_1_7_4_N84), .B2(pe_1_7_4_n27), .C1(pe_1_7_4_N76), .C2(pe_1_7_4_n28), 
        .ZN(pe_1_7_4_n29) );
  INV_X1 pe_1_7_4_U46 ( .A(pe_1_7_4_n29), .ZN(pe_1_7_4_n72) );
  XNOR2_X1 pe_1_7_4_U45 ( .A(pe_1_7_4_n67), .B(int_data_res_7__4__0_), .ZN(
        pe_1_7_4_N70) );
  AOI222_X1 pe_1_7_4_U44 ( .A1(i_data_acc[24]), .A2(pe_1_7_4_n61), .B1(
        pe_1_7_4_n1), .B2(pe_1_7_4_n27), .C1(pe_1_7_4_N70), .C2(pe_1_7_4_n28), 
        .ZN(pe_1_7_4_n35) );
  INV_X1 pe_1_7_4_U43 ( .A(pe_1_7_4_n35), .ZN(pe_1_7_4_n78) );
  NAND2_X1 pe_1_7_4_U42 ( .A1(pe_1_7_4_int_data_0_), .A2(pe_1_7_4_n3), .ZN(
        pe_1_7_4_sub_81_carry[1]) );
  INV_X1 pe_1_7_4_U41 ( .A(pe_1_7_4_int_data_1_), .ZN(pe_1_7_4_n68) );
  INV_X1 pe_1_7_4_U40 ( .A(pe_1_7_4_int_data_2_), .ZN(pe_1_7_4_n69) );
  AND2_X1 pe_1_7_4_U39 ( .A1(pe_1_7_4_int_data_0_), .A2(int_data_res_7__4__0_), 
        .ZN(pe_1_7_4_n2) );
  AOI222_X1 pe_1_7_4_U38 ( .A1(pe_1_7_4_n61), .A2(i_data_acc[31]), .B1(
        pe_1_7_4_N85), .B2(pe_1_7_4_n27), .C1(pe_1_7_4_N77), .C2(pe_1_7_4_n28), 
        .ZN(pe_1_7_4_n26) );
  INV_X1 pe_1_7_4_U37 ( .A(pe_1_7_4_n26), .ZN(pe_1_7_4_n71) );
  NOR3_X1 pe_1_7_4_U36 ( .A1(pe_1_7_4_n58), .A2(pe_1_7_4_n62), .A3(int_ckg[3]), 
        .ZN(pe_1_7_4_n36) );
  OR2_X1 pe_1_7_4_U35 ( .A1(pe_1_7_4_n36), .A2(pe_1_7_4_n61), .ZN(pe_1_7_4_N90) );
  AND2_X1 pe_1_7_4_U34 ( .A1(int_data_x_7__4__2_), .A2(n30), .ZN(
        pe_1_7_4_int_data_2_) );
  AND2_X1 pe_1_7_4_U33 ( .A1(int_data_x_7__4__1_), .A2(n30), .ZN(
        pe_1_7_4_int_data_1_) );
  INV_X1 pe_1_7_4_U32 ( .A(n42), .ZN(pe_1_7_4_n60) );
  BUF_X1 pe_1_7_4_U31 ( .A(n64), .Z(pe_1_7_4_n61) );
  AND2_X1 pe_1_7_4_U30 ( .A1(int_data_x_7__4__3_), .A2(n30), .ZN(
        pe_1_7_4_int_data_3_) );
  AND2_X1 pe_1_7_4_U29 ( .A1(int_data_x_7__4__0_), .A2(n30), .ZN(
        pe_1_7_4_int_data_0_) );
  INV_X1 pe_1_7_4_U28 ( .A(n36), .ZN(pe_1_7_4_n59) );
  NAND2_X1 pe_1_7_4_U27 ( .A1(pe_1_7_4_n44), .A2(pe_1_7_4_n59), .ZN(
        pe_1_7_4_n41) );
  AND3_X1 pe_1_7_4_U26 ( .A1(n78), .A2(pe_1_7_4_n60), .A3(n55), .ZN(
        pe_1_7_4_n44) );
  INV_X1 pe_1_7_4_U25 ( .A(pe_1_7_4_int_data_3_), .ZN(pe_1_7_4_n70) );
  NOR2_X1 pe_1_7_4_U24 ( .A1(pe_1_7_4_n64), .A2(n55), .ZN(pe_1_7_4_n43) );
  NOR2_X1 pe_1_7_4_U23 ( .A1(pe_1_7_4_n57), .A2(pe_1_7_4_n61), .ZN(
        pe_1_7_4_n28) );
  NOR2_X1 pe_1_7_4_U22 ( .A1(n22), .A2(pe_1_7_4_n61), .ZN(pe_1_7_4_n27) );
  INV_X1 pe_1_7_4_U21 ( .A(pe_1_7_4_int_data_0_), .ZN(pe_1_7_4_n67) );
  INV_X1 pe_1_7_4_U20 ( .A(pe_1_7_4_n41), .ZN(pe_1_7_4_n84) );
  INV_X1 pe_1_7_4_U19 ( .A(pe_1_7_4_n37), .ZN(pe_1_7_4_n82) );
  INV_X1 pe_1_7_4_U18 ( .A(pe_1_7_4_n38), .ZN(pe_1_7_4_n81) );
  INV_X1 pe_1_7_4_U17 ( .A(pe_1_7_4_n39), .ZN(pe_1_7_4_n80) );
  NOR2_X1 pe_1_7_4_U16 ( .A1(pe_1_7_4_n63), .A2(pe_1_7_4_n42), .ZN(
        pe_1_7_4_N59) );
  NOR2_X1 pe_1_7_4_U15 ( .A1(pe_1_7_4_n63), .A2(pe_1_7_4_n41), .ZN(
        pe_1_7_4_N60) );
  NOR2_X1 pe_1_7_4_U14 ( .A1(pe_1_7_4_n63), .A2(pe_1_7_4_n38), .ZN(
        pe_1_7_4_N63) );
  NOR2_X1 pe_1_7_4_U13 ( .A1(pe_1_7_4_n63), .A2(pe_1_7_4_n40), .ZN(
        pe_1_7_4_N61) );
  NOR2_X1 pe_1_7_4_U12 ( .A1(pe_1_7_4_n63), .A2(pe_1_7_4_n39), .ZN(
        pe_1_7_4_N62) );
  NOR2_X1 pe_1_7_4_U11 ( .A1(pe_1_7_4_n37), .A2(pe_1_7_4_n63), .ZN(
        pe_1_7_4_N64) );
  NAND2_X1 pe_1_7_4_U10 ( .A1(pe_1_7_4_n44), .A2(n36), .ZN(pe_1_7_4_n42) );
  BUF_X1 pe_1_7_4_U9 ( .A(n36), .Z(pe_1_7_4_n55) );
  INV_X1 pe_1_7_4_U8 ( .A(pe_1_7_4_n63), .ZN(pe_1_7_4_n62) );
  BUF_X1 pe_1_7_4_U7 ( .A(n36), .Z(pe_1_7_4_n56) );
  INV_X1 pe_1_7_4_U6 ( .A(pe_1_7_4_n42), .ZN(pe_1_7_4_n83) );
  INV_X1 pe_1_7_4_U5 ( .A(pe_1_7_4_n40), .ZN(pe_1_7_4_n79) );
  INV_X2 pe_1_7_4_U4 ( .A(n86), .ZN(pe_1_7_4_n66) );
  XOR2_X1 pe_1_7_4_U3 ( .A(pe_1_7_4_int_data_0_), .B(int_data_res_7__4__0_), 
        .Z(pe_1_7_4_n1) );
  DFFR_X1 pe_1_7_4_int_q_acc_reg_0_ ( .D(pe_1_7_4_n78), .CK(pe_1_7_4_net2872), 
        .RN(pe_1_7_4_n66), .Q(int_data_res_7__4__0_), .QN(pe_1_7_4_n3) );
  DFFR_X1 pe_1_7_4_int_q_reg_v_reg_0__0_ ( .D(i_data_conv_v[12]), .CK(
        pe_1_7_4_net2842), .RN(pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_v[20]) );
  DFFR_X1 pe_1_7_4_int_q_reg_v_reg_0__1_ ( .D(i_data_conv_v[13]), .CK(
        pe_1_7_4_net2842), .RN(pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_v[21]) );
  DFFR_X1 pe_1_7_4_int_q_reg_v_reg_0__2_ ( .D(i_data_conv_v[14]), .CK(
        pe_1_7_4_net2842), .RN(pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_v[22]) );
  DFFR_X1 pe_1_7_4_int_q_reg_v_reg_0__3_ ( .D(i_data_conv_v[15]), .CK(
        pe_1_7_4_net2842), .RN(pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_v[23]) );
  DFFR_X1 pe_1_7_4_int_q_reg_v_reg_1__0_ ( .D(i_data_conv_v[12]), .CK(
        pe_1_7_4_net2847), .RN(pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_v[16]) );
  DFFR_X1 pe_1_7_4_int_q_reg_v_reg_1__1_ ( .D(i_data_conv_v[13]), .CK(
        pe_1_7_4_net2847), .RN(pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_v[17]) );
  DFFR_X1 pe_1_7_4_int_q_reg_v_reg_1__2_ ( .D(i_data_conv_v[14]), .CK(
        pe_1_7_4_net2847), .RN(pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_v[18]) );
  DFFR_X1 pe_1_7_4_int_q_reg_v_reg_1__3_ ( .D(i_data_conv_v[15]), .CK(
        pe_1_7_4_net2847), .RN(pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_v[19]) );
  DFFR_X1 pe_1_7_4_int_q_reg_v_reg_2__0_ ( .D(i_data_conv_v[12]), .CK(
        pe_1_7_4_net2852), .RN(pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_v[12]) );
  DFFR_X1 pe_1_7_4_int_q_reg_v_reg_2__1_ ( .D(i_data_conv_v[13]), .CK(
        pe_1_7_4_net2852), .RN(pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_v[13]) );
  DFFR_X1 pe_1_7_4_int_q_reg_v_reg_2__2_ ( .D(i_data_conv_v[14]), .CK(
        pe_1_7_4_net2852), .RN(pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_v[14]) );
  DFFR_X1 pe_1_7_4_int_q_reg_v_reg_2__3_ ( .D(i_data_conv_v[15]), .CK(
        pe_1_7_4_net2852), .RN(pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_v[15]) );
  DFFR_X1 pe_1_7_4_int_q_reg_v_reg_3__0_ ( .D(i_data_conv_v[12]), .CK(
        pe_1_7_4_net2857), .RN(pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_v[8]) );
  DFFR_X1 pe_1_7_4_int_q_reg_v_reg_3__1_ ( .D(i_data_conv_v[13]), .CK(
        pe_1_7_4_net2857), .RN(pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_v[9]) );
  DFFR_X1 pe_1_7_4_int_q_reg_v_reg_3__2_ ( .D(i_data_conv_v[14]), .CK(
        pe_1_7_4_net2857), .RN(pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_v[10]) );
  DFFR_X1 pe_1_7_4_int_q_reg_v_reg_3__3_ ( .D(i_data_conv_v[15]), .CK(
        pe_1_7_4_net2857), .RN(pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_v[11]) );
  DFFR_X1 pe_1_7_4_int_q_reg_v_reg_4__0_ ( .D(i_data_conv_v[12]), .CK(
        pe_1_7_4_net2862), .RN(pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_v[4]) );
  DFFR_X1 pe_1_7_4_int_q_reg_v_reg_4__1_ ( .D(i_data_conv_v[13]), .CK(
        pe_1_7_4_net2862), .RN(pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_v[5]) );
  DFFR_X1 pe_1_7_4_int_q_reg_v_reg_4__2_ ( .D(i_data_conv_v[14]), .CK(
        pe_1_7_4_net2862), .RN(pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_v[6]) );
  DFFR_X1 pe_1_7_4_int_q_reg_v_reg_4__3_ ( .D(i_data_conv_v[15]), .CK(
        pe_1_7_4_net2862), .RN(pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_v[7]) );
  DFFR_X1 pe_1_7_4_int_q_reg_v_reg_5__0_ ( .D(i_data_conv_v[12]), .CK(
        pe_1_7_4_net2867), .RN(pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_v[0]) );
  DFFR_X1 pe_1_7_4_int_q_reg_v_reg_5__1_ ( .D(i_data_conv_v[13]), .CK(
        pe_1_7_4_net2867), .RN(pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_v[1]) );
  DFFR_X1 pe_1_7_4_int_q_reg_v_reg_5__2_ ( .D(i_data_conv_v[14]), .CK(
        pe_1_7_4_net2867), .RN(pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_v[2]) );
  DFFR_X1 pe_1_7_4_int_q_reg_v_reg_5__3_ ( .D(i_data_conv_v[15]), .CK(
        pe_1_7_4_net2867), .RN(pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_7_4_int_q_reg_h_reg_0__0_ ( .D(int_data_x_7__5__0_), .SI(
        i_data_conv_v[12]), .SE(pe_1_7_4_n62), .CK(pe_1_7_4_net2811), .RN(
        pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_7_4_int_q_reg_h_reg_0__1_ ( .D(int_data_x_7__5__1_), .SI(
        i_data_conv_v[13]), .SE(pe_1_7_4_n62), .CK(pe_1_7_4_net2811), .RN(
        pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_7_4_int_q_reg_h_reg_0__2_ ( .D(int_data_x_7__5__2_), .SI(
        i_data_conv_v[14]), .SE(pe_1_7_4_n62), .CK(pe_1_7_4_net2811), .RN(
        pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_7_4_int_q_reg_h_reg_0__3_ ( .D(int_data_x_7__5__3_), .SI(
        i_data_conv_v[15]), .SE(pe_1_7_4_n62), .CK(pe_1_7_4_net2811), .RN(
        pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_7_4_int_q_reg_h_reg_1__0_ ( .D(int_data_x_7__5__0_), .SI(
        i_data_conv_v[12]), .SE(pe_1_7_4_n62), .CK(pe_1_7_4_net2817), .RN(
        pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_7_4_int_q_reg_h_reg_1__1_ ( .D(int_data_x_7__5__1_), .SI(
        i_data_conv_v[13]), .SE(pe_1_7_4_n62), .CK(pe_1_7_4_net2817), .RN(
        pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_7_4_int_q_reg_h_reg_1__2_ ( .D(int_data_x_7__5__2_), .SI(
        i_data_conv_v[14]), .SE(pe_1_7_4_n62), .CK(pe_1_7_4_net2817), .RN(
        pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_7_4_int_q_reg_h_reg_1__3_ ( .D(int_data_x_7__5__3_), .SI(
        i_data_conv_v[15]), .SE(pe_1_7_4_n62), .CK(pe_1_7_4_net2817), .RN(
        pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_7_4_int_q_reg_h_reg_2__0_ ( .D(int_data_x_7__5__0_), .SI(
        i_data_conv_v[12]), .SE(pe_1_7_4_n62), .CK(pe_1_7_4_net2822), .RN(
        pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_7_4_int_q_reg_h_reg_2__1_ ( .D(int_data_x_7__5__1_), .SI(
        i_data_conv_v[13]), .SE(pe_1_7_4_n62), .CK(pe_1_7_4_net2822), .RN(
        pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_7_4_int_q_reg_h_reg_2__2_ ( .D(int_data_x_7__5__2_), .SI(
        i_data_conv_v[14]), .SE(pe_1_7_4_n62), .CK(pe_1_7_4_net2822), .RN(
        pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_7_4_int_q_reg_h_reg_2__3_ ( .D(int_data_x_7__5__3_), .SI(
        i_data_conv_v[15]), .SE(pe_1_7_4_n62), .CK(pe_1_7_4_net2822), .RN(
        pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_7_4_int_q_reg_h_reg_3__0_ ( .D(int_data_x_7__5__0_), .SI(
        i_data_conv_v[12]), .SE(pe_1_7_4_n62), .CK(pe_1_7_4_net2827), .RN(
        pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_7_4_int_q_reg_h_reg_3__1_ ( .D(int_data_x_7__5__1_), .SI(
        i_data_conv_v[13]), .SE(pe_1_7_4_n62), .CK(pe_1_7_4_net2827), .RN(
        pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_7_4_int_q_reg_h_reg_3__2_ ( .D(int_data_x_7__5__2_), .SI(
        i_data_conv_v[14]), .SE(pe_1_7_4_n62), .CK(pe_1_7_4_net2827), .RN(
        pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_7_4_int_q_reg_h_reg_3__3_ ( .D(int_data_x_7__5__3_), .SI(
        i_data_conv_v[15]), .SE(pe_1_7_4_n62), .CK(pe_1_7_4_net2827), .RN(
        pe_1_7_4_n66), .Q(pe_1_7_4_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_7_4_int_q_reg_h_reg_4__0_ ( .D(int_data_x_7__5__0_), .SI(
        i_data_conv_v[12]), .SE(n70), .CK(pe_1_7_4_net2832), .RN(pe_1_7_4_n66), 
        .Q(pe_1_7_4_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_7_4_int_q_reg_h_reg_4__1_ ( .D(int_data_x_7__5__1_), .SI(
        i_data_conv_v[13]), .SE(n70), .CK(pe_1_7_4_net2832), .RN(pe_1_7_4_n66), 
        .Q(pe_1_7_4_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_7_4_int_q_reg_h_reg_4__2_ ( .D(int_data_x_7__5__2_), .SI(
        i_data_conv_v[14]), .SE(n70), .CK(pe_1_7_4_net2832), .RN(pe_1_7_4_n66), 
        .Q(pe_1_7_4_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_7_4_int_q_reg_h_reg_4__3_ ( .D(int_data_x_7__5__3_), .SI(
        i_data_conv_v[15]), .SE(n70), .CK(pe_1_7_4_net2832), .RN(pe_1_7_4_n66), 
        .Q(pe_1_7_4_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_7_4_int_q_reg_h_reg_5__0_ ( .D(int_data_x_7__5__0_), .SI(
        i_data_conv_v[12]), .SE(n70), .CK(pe_1_7_4_net2837), .RN(pe_1_7_4_n66), 
        .Q(pe_1_7_4_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_7_4_int_q_reg_h_reg_5__1_ ( .D(int_data_x_7__5__1_), .SI(
        i_data_conv_v[13]), .SE(n70), .CK(pe_1_7_4_net2837), .RN(pe_1_7_4_n66), 
        .Q(pe_1_7_4_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_7_4_int_q_reg_h_reg_5__2_ ( .D(int_data_x_7__5__2_), .SI(
        i_data_conv_v[14]), .SE(n70), .CK(pe_1_7_4_net2837), .RN(pe_1_7_4_n66), 
        .Q(pe_1_7_4_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_7_4_int_q_reg_h_reg_5__3_ ( .D(int_data_x_7__5__3_), .SI(
        i_data_conv_v[15]), .SE(n70), .CK(pe_1_7_4_net2837), .RN(pe_1_7_4_n66), 
        .Q(pe_1_7_4_int_q_reg_h[3]) );
  FA_X1 pe_1_7_4_sub_81_U2_7 ( .A(int_data_res_7__4__7_), .B(pe_1_7_4_n70), 
        .CI(pe_1_7_4_sub_81_carry[7]), .S(pe_1_7_4_N77) );
  FA_X1 pe_1_7_4_sub_81_U2_6 ( .A(int_data_res_7__4__6_), .B(pe_1_7_4_n70), 
        .CI(pe_1_7_4_sub_81_carry[6]), .CO(pe_1_7_4_sub_81_carry[7]), .S(
        pe_1_7_4_N76) );
  FA_X1 pe_1_7_4_sub_81_U2_5 ( .A(int_data_res_7__4__5_), .B(pe_1_7_4_n70), 
        .CI(pe_1_7_4_sub_81_carry[5]), .CO(pe_1_7_4_sub_81_carry[6]), .S(
        pe_1_7_4_N75) );
  FA_X1 pe_1_7_4_sub_81_U2_4 ( .A(int_data_res_7__4__4_), .B(pe_1_7_4_n70), 
        .CI(pe_1_7_4_sub_81_carry[4]), .CO(pe_1_7_4_sub_81_carry[5]), .S(
        pe_1_7_4_N74) );
  FA_X1 pe_1_7_4_sub_81_U2_3 ( .A(int_data_res_7__4__3_), .B(pe_1_7_4_n70), 
        .CI(pe_1_7_4_sub_81_carry[3]), .CO(pe_1_7_4_sub_81_carry[4]), .S(
        pe_1_7_4_N73) );
  FA_X1 pe_1_7_4_sub_81_U2_2 ( .A(int_data_res_7__4__2_), .B(pe_1_7_4_n69), 
        .CI(pe_1_7_4_sub_81_carry[2]), .CO(pe_1_7_4_sub_81_carry[3]), .S(
        pe_1_7_4_N72) );
  FA_X1 pe_1_7_4_sub_81_U2_1 ( .A(int_data_res_7__4__1_), .B(pe_1_7_4_n68), 
        .CI(pe_1_7_4_sub_81_carry[1]), .CO(pe_1_7_4_sub_81_carry[2]), .S(
        pe_1_7_4_N71) );
  FA_X1 pe_1_7_4_add_83_U1_7 ( .A(int_data_res_7__4__7_), .B(
        pe_1_7_4_int_data_3_), .CI(pe_1_7_4_add_83_carry[7]), .S(pe_1_7_4_N85)
         );
  FA_X1 pe_1_7_4_add_83_U1_6 ( .A(int_data_res_7__4__6_), .B(
        pe_1_7_4_int_data_3_), .CI(pe_1_7_4_add_83_carry[6]), .CO(
        pe_1_7_4_add_83_carry[7]), .S(pe_1_7_4_N84) );
  FA_X1 pe_1_7_4_add_83_U1_5 ( .A(int_data_res_7__4__5_), .B(
        pe_1_7_4_int_data_3_), .CI(pe_1_7_4_add_83_carry[5]), .CO(
        pe_1_7_4_add_83_carry[6]), .S(pe_1_7_4_N83) );
  FA_X1 pe_1_7_4_add_83_U1_4 ( .A(int_data_res_7__4__4_), .B(
        pe_1_7_4_int_data_3_), .CI(pe_1_7_4_add_83_carry[4]), .CO(
        pe_1_7_4_add_83_carry[5]), .S(pe_1_7_4_N82) );
  FA_X1 pe_1_7_4_add_83_U1_3 ( .A(int_data_res_7__4__3_), .B(
        pe_1_7_4_int_data_3_), .CI(pe_1_7_4_add_83_carry[3]), .CO(
        pe_1_7_4_add_83_carry[4]), .S(pe_1_7_4_N81) );
  FA_X1 pe_1_7_4_add_83_U1_2 ( .A(int_data_res_7__4__2_), .B(
        pe_1_7_4_int_data_2_), .CI(pe_1_7_4_add_83_carry[2]), .CO(
        pe_1_7_4_add_83_carry[3]), .S(pe_1_7_4_N80) );
  FA_X1 pe_1_7_4_add_83_U1_1 ( .A(int_data_res_7__4__1_), .B(
        pe_1_7_4_int_data_1_), .CI(pe_1_7_4_n2), .CO(pe_1_7_4_add_83_carry[2]), 
        .S(pe_1_7_4_N79) );
  NAND3_X1 pe_1_7_4_U56 ( .A1(n36), .A2(pe_1_7_4_n43), .A3(n42), .ZN(
        pe_1_7_4_n40) );
  NAND3_X1 pe_1_7_4_U55 ( .A1(pe_1_7_4_n43), .A2(pe_1_7_4_n59), .A3(n42), .ZN(
        pe_1_7_4_n39) );
  NAND3_X1 pe_1_7_4_U54 ( .A1(pe_1_7_4_n43), .A2(pe_1_7_4_n60), .A3(n36), .ZN(
        pe_1_7_4_n38) );
  NAND3_X1 pe_1_7_4_U53 ( .A1(pe_1_7_4_n59), .A2(pe_1_7_4_n60), .A3(
        pe_1_7_4_n43), .ZN(pe_1_7_4_n37) );
  DFFR_X1 pe_1_7_4_int_q_acc_reg_6_ ( .D(pe_1_7_4_n72), .CK(pe_1_7_4_net2872), 
        .RN(pe_1_7_4_n65), .Q(int_data_res_7__4__6_) );
  DFFR_X1 pe_1_7_4_int_q_acc_reg_5_ ( .D(pe_1_7_4_n73), .CK(pe_1_7_4_net2872), 
        .RN(pe_1_7_4_n65), .Q(int_data_res_7__4__5_) );
  DFFR_X1 pe_1_7_4_int_q_acc_reg_4_ ( .D(pe_1_7_4_n74), .CK(pe_1_7_4_net2872), 
        .RN(pe_1_7_4_n65), .Q(int_data_res_7__4__4_) );
  DFFR_X1 pe_1_7_4_int_q_acc_reg_3_ ( .D(pe_1_7_4_n75), .CK(pe_1_7_4_net2872), 
        .RN(pe_1_7_4_n65), .Q(int_data_res_7__4__3_) );
  DFFR_X1 pe_1_7_4_int_q_acc_reg_2_ ( .D(pe_1_7_4_n76), .CK(pe_1_7_4_net2872), 
        .RN(pe_1_7_4_n65), .Q(int_data_res_7__4__2_) );
  DFFR_X1 pe_1_7_4_int_q_acc_reg_1_ ( .D(pe_1_7_4_n77), .CK(pe_1_7_4_net2872), 
        .RN(pe_1_7_4_n65), .Q(int_data_res_7__4__1_) );
  DFFR_X1 pe_1_7_4_int_q_acc_reg_7_ ( .D(pe_1_7_4_n71), .CK(pe_1_7_4_net2872), 
        .RN(pe_1_7_4_n65), .Q(int_data_res_7__4__7_) );
  CLKGATETST_X1 pe_1_7_4_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_7_4_n82), .SE(1'b0), .GCK(pe_1_7_4_net2811) );
  CLKGATETST_X1 pe_1_7_4_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_7_4_n81), .SE(1'b0), .GCK(pe_1_7_4_net2817) );
  CLKGATETST_X1 pe_1_7_4_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_7_4_n80), .SE(1'b0), .GCK(pe_1_7_4_net2822) );
  CLKGATETST_X1 pe_1_7_4_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_7_4_n79), .SE(1'b0), .GCK(pe_1_7_4_net2827) );
  CLKGATETST_X1 pe_1_7_4_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_7_4_n84), .SE(1'b0), .GCK(pe_1_7_4_net2832) );
  CLKGATETST_X1 pe_1_7_4_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_7_4_n83), .SE(1'b0), .GCK(pe_1_7_4_net2837) );
  CLKGATETST_X1 pe_1_7_4_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_7_4_N64), .SE(1'b0), .GCK(pe_1_7_4_net2842) );
  CLKGATETST_X1 pe_1_7_4_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_7_4_N63), .SE(1'b0), .GCK(pe_1_7_4_net2847) );
  CLKGATETST_X1 pe_1_7_4_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_7_4_N62), .SE(1'b0), .GCK(pe_1_7_4_net2852) );
  CLKGATETST_X1 pe_1_7_4_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_7_4_N61), .SE(1'b0), .GCK(pe_1_7_4_net2857) );
  CLKGATETST_X1 pe_1_7_4_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_7_4_N60), .SE(1'b0), .GCK(pe_1_7_4_net2862) );
  CLKGATETST_X1 pe_1_7_4_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_7_4_N59), .SE(1'b0), .GCK(pe_1_7_4_net2867) );
  CLKGATETST_X1 pe_1_7_4_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_7_4_N90), .SE(1'b0), .GCK(pe_1_7_4_net2872) );
  CLKBUF_X1 pe_1_7_5_U106 ( .A(pe_1_7_5_n66), .Z(pe_1_7_5_n65) );
  INV_X1 pe_1_7_5_U105 ( .A(n78), .ZN(pe_1_7_5_n64) );
  INV_X1 pe_1_7_5_U104 ( .A(n70), .ZN(pe_1_7_5_n63) );
  INV_X1 pe_1_7_5_U103 ( .A(n30), .ZN(pe_1_7_5_n58) );
  INV_X1 pe_1_7_5_U102 ( .A(n22), .ZN(pe_1_7_5_n57) );
  MUX2_X1 pe_1_7_5_U101 ( .A(pe_1_7_5_n54), .B(pe_1_7_5_n51), .S(n55), .Z(
        int_data_x_7__5__3_) );
  MUX2_X1 pe_1_7_5_U100 ( .A(pe_1_7_5_n53), .B(pe_1_7_5_n52), .S(n42), .Z(
        pe_1_7_5_n54) );
  MUX2_X1 pe_1_7_5_U99 ( .A(pe_1_7_5_int_q_reg_h[23]), .B(
        pe_1_7_5_int_q_reg_h[19]), .S(pe_1_7_5_n56), .Z(pe_1_7_5_n53) );
  MUX2_X1 pe_1_7_5_U98 ( .A(pe_1_7_5_int_q_reg_h[15]), .B(
        pe_1_7_5_int_q_reg_h[11]), .S(pe_1_7_5_n56), .Z(pe_1_7_5_n52) );
  MUX2_X1 pe_1_7_5_U97 ( .A(pe_1_7_5_int_q_reg_h[7]), .B(
        pe_1_7_5_int_q_reg_h[3]), .S(pe_1_7_5_n56), .Z(pe_1_7_5_n51) );
  MUX2_X1 pe_1_7_5_U96 ( .A(pe_1_7_5_n50), .B(pe_1_7_5_n47), .S(n55), .Z(
        int_data_x_7__5__2_) );
  MUX2_X1 pe_1_7_5_U95 ( .A(pe_1_7_5_n49), .B(pe_1_7_5_n48), .S(n42), .Z(
        pe_1_7_5_n50) );
  MUX2_X1 pe_1_7_5_U94 ( .A(pe_1_7_5_int_q_reg_h[22]), .B(
        pe_1_7_5_int_q_reg_h[18]), .S(pe_1_7_5_n56), .Z(pe_1_7_5_n49) );
  MUX2_X1 pe_1_7_5_U93 ( .A(pe_1_7_5_int_q_reg_h[14]), .B(
        pe_1_7_5_int_q_reg_h[10]), .S(pe_1_7_5_n56), .Z(pe_1_7_5_n48) );
  MUX2_X1 pe_1_7_5_U92 ( .A(pe_1_7_5_int_q_reg_h[6]), .B(
        pe_1_7_5_int_q_reg_h[2]), .S(pe_1_7_5_n56), .Z(pe_1_7_5_n47) );
  MUX2_X1 pe_1_7_5_U91 ( .A(pe_1_7_5_n46), .B(pe_1_7_5_n24), .S(n55), .Z(
        int_data_x_7__5__1_) );
  MUX2_X1 pe_1_7_5_U90 ( .A(pe_1_7_5_n45), .B(pe_1_7_5_n25), .S(n42), .Z(
        pe_1_7_5_n46) );
  MUX2_X1 pe_1_7_5_U89 ( .A(pe_1_7_5_int_q_reg_h[21]), .B(
        pe_1_7_5_int_q_reg_h[17]), .S(pe_1_7_5_n56), .Z(pe_1_7_5_n45) );
  MUX2_X1 pe_1_7_5_U88 ( .A(pe_1_7_5_int_q_reg_h[13]), .B(
        pe_1_7_5_int_q_reg_h[9]), .S(pe_1_7_5_n56), .Z(pe_1_7_5_n25) );
  MUX2_X1 pe_1_7_5_U87 ( .A(pe_1_7_5_int_q_reg_h[5]), .B(
        pe_1_7_5_int_q_reg_h[1]), .S(pe_1_7_5_n56), .Z(pe_1_7_5_n24) );
  MUX2_X1 pe_1_7_5_U86 ( .A(pe_1_7_5_n23), .B(pe_1_7_5_n20), .S(n55), .Z(
        int_data_x_7__5__0_) );
  MUX2_X1 pe_1_7_5_U85 ( .A(pe_1_7_5_n22), .B(pe_1_7_5_n21), .S(n42), .Z(
        pe_1_7_5_n23) );
  MUX2_X1 pe_1_7_5_U84 ( .A(pe_1_7_5_int_q_reg_h[20]), .B(
        pe_1_7_5_int_q_reg_h[16]), .S(pe_1_7_5_n56), .Z(pe_1_7_5_n22) );
  MUX2_X1 pe_1_7_5_U83 ( .A(pe_1_7_5_int_q_reg_h[12]), .B(
        pe_1_7_5_int_q_reg_h[8]), .S(pe_1_7_5_n56), .Z(pe_1_7_5_n21) );
  MUX2_X1 pe_1_7_5_U82 ( .A(pe_1_7_5_int_q_reg_h[4]), .B(
        pe_1_7_5_int_q_reg_h[0]), .S(pe_1_7_5_n56), .Z(pe_1_7_5_n20) );
  MUX2_X1 pe_1_7_5_U81 ( .A(pe_1_7_5_n19), .B(pe_1_7_5_n16), .S(n55), .Z(
        int_data_y_7__5__3_) );
  MUX2_X1 pe_1_7_5_U80 ( .A(pe_1_7_5_n18), .B(pe_1_7_5_n17), .S(n42), .Z(
        pe_1_7_5_n19) );
  MUX2_X1 pe_1_7_5_U79 ( .A(pe_1_7_5_int_q_reg_v[23]), .B(
        pe_1_7_5_int_q_reg_v[19]), .S(pe_1_7_5_n55), .Z(pe_1_7_5_n18) );
  MUX2_X1 pe_1_7_5_U78 ( .A(pe_1_7_5_int_q_reg_v[15]), .B(
        pe_1_7_5_int_q_reg_v[11]), .S(pe_1_7_5_n55), .Z(pe_1_7_5_n17) );
  MUX2_X1 pe_1_7_5_U77 ( .A(pe_1_7_5_int_q_reg_v[7]), .B(
        pe_1_7_5_int_q_reg_v[3]), .S(pe_1_7_5_n55), .Z(pe_1_7_5_n16) );
  MUX2_X1 pe_1_7_5_U76 ( .A(pe_1_7_5_n15), .B(pe_1_7_5_n12), .S(n55), .Z(
        int_data_y_7__5__2_) );
  MUX2_X1 pe_1_7_5_U75 ( .A(pe_1_7_5_n14), .B(pe_1_7_5_n13), .S(n42), .Z(
        pe_1_7_5_n15) );
  MUX2_X1 pe_1_7_5_U74 ( .A(pe_1_7_5_int_q_reg_v[22]), .B(
        pe_1_7_5_int_q_reg_v[18]), .S(pe_1_7_5_n55), .Z(pe_1_7_5_n14) );
  MUX2_X1 pe_1_7_5_U73 ( .A(pe_1_7_5_int_q_reg_v[14]), .B(
        pe_1_7_5_int_q_reg_v[10]), .S(pe_1_7_5_n55), .Z(pe_1_7_5_n13) );
  MUX2_X1 pe_1_7_5_U72 ( .A(pe_1_7_5_int_q_reg_v[6]), .B(
        pe_1_7_5_int_q_reg_v[2]), .S(pe_1_7_5_n55), .Z(pe_1_7_5_n12) );
  MUX2_X1 pe_1_7_5_U71 ( .A(pe_1_7_5_n11), .B(pe_1_7_5_n8), .S(n55), .Z(
        int_data_y_7__5__1_) );
  MUX2_X1 pe_1_7_5_U70 ( .A(pe_1_7_5_n10), .B(pe_1_7_5_n9), .S(n42), .Z(
        pe_1_7_5_n11) );
  MUX2_X1 pe_1_7_5_U69 ( .A(pe_1_7_5_int_q_reg_v[21]), .B(
        pe_1_7_5_int_q_reg_v[17]), .S(pe_1_7_5_n55), .Z(pe_1_7_5_n10) );
  MUX2_X1 pe_1_7_5_U68 ( .A(pe_1_7_5_int_q_reg_v[13]), .B(
        pe_1_7_5_int_q_reg_v[9]), .S(pe_1_7_5_n55), .Z(pe_1_7_5_n9) );
  MUX2_X1 pe_1_7_5_U67 ( .A(pe_1_7_5_int_q_reg_v[5]), .B(
        pe_1_7_5_int_q_reg_v[1]), .S(pe_1_7_5_n55), .Z(pe_1_7_5_n8) );
  MUX2_X1 pe_1_7_5_U66 ( .A(pe_1_7_5_n7), .B(pe_1_7_5_n4), .S(n55), .Z(
        int_data_y_7__5__0_) );
  MUX2_X1 pe_1_7_5_U65 ( .A(pe_1_7_5_n6), .B(pe_1_7_5_n5), .S(n42), .Z(
        pe_1_7_5_n7) );
  MUX2_X1 pe_1_7_5_U64 ( .A(pe_1_7_5_int_q_reg_v[20]), .B(
        pe_1_7_5_int_q_reg_v[16]), .S(pe_1_7_5_n55), .Z(pe_1_7_5_n6) );
  MUX2_X1 pe_1_7_5_U63 ( .A(pe_1_7_5_int_q_reg_v[12]), .B(
        pe_1_7_5_int_q_reg_v[8]), .S(pe_1_7_5_n55), .Z(pe_1_7_5_n5) );
  MUX2_X1 pe_1_7_5_U62 ( .A(pe_1_7_5_int_q_reg_v[4]), .B(
        pe_1_7_5_int_q_reg_v[0]), .S(pe_1_7_5_n55), .Z(pe_1_7_5_n4) );
  AOI222_X1 pe_1_7_5_U61 ( .A1(i_data_acc[17]), .A2(pe_1_7_5_n61), .B1(
        pe_1_7_5_N79), .B2(pe_1_7_5_n27), .C1(pe_1_7_5_N71), .C2(pe_1_7_5_n28), 
        .ZN(pe_1_7_5_n34) );
  INV_X1 pe_1_7_5_U60 ( .A(pe_1_7_5_n34), .ZN(pe_1_7_5_n77) );
  AOI222_X1 pe_1_7_5_U59 ( .A1(i_data_acc[18]), .A2(pe_1_7_5_n61), .B1(
        pe_1_7_5_N80), .B2(pe_1_7_5_n27), .C1(pe_1_7_5_N72), .C2(pe_1_7_5_n28), 
        .ZN(pe_1_7_5_n33) );
  INV_X1 pe_1_7_5_U58 ( .A(pe_1_7_5_n33), .ZN(pe_1_7_5_n76) );
  AOI222_X1 pe_1_7_5_U57 ( .A1(i_data_acc[19]), .A2(pe_1_7_5_n61), .B1(
        pe_1_7_5_N81), .B2(pe_1_7_5_n27), .C1(pe_1_7_5_N73), .C2(pe_1_7_5_n28), 
        .ZN(pe_1_7_5_n32) );
  INV_X1 pe_1_7_5_U52 ( .A(pe_1_7_5_n32), .ZN(pe_1_7_5_n75) );
  AOI222_X1 pe_1_7_5_U51 ( .A1(i_data_acc[20]), .A2(pe_1_7_5_n61), .B1(
        pe_1_7_5_N82), .B2(pe_1_7_5_n27), .C1(pe_1_7_5_N74), .C2(pe_1_7_5_n28), 
        .ZN(pe_1_7_5_n31) );
  INV_X1 pe_1_7_5_U50 ( .A(pe_1_7_5_n31), .ZN(pe_1_7_5_n74) );
  AOI222_X1 pe_1_7_5_U49 ( .A1(i_data_acc[21]), .A2(pe_1_7_5_n61), .B1(
        pe_1_7_5_N83), .B2(pe_1_7_5_n27), .C1(pe_1_7_5_N75), .C2(pe_1_7_5_n28), 
        .ZN(pe_1_7_5_n30) );
  INV_X1 pe_1_7_5_U48 ( .A(pe_1_7_5_n30), .ZN(pe_1_7_5_n73) );
  AOI222_X1 pe_1_7_5_U47 ( .A1(i_data_acc[22]), .A2(pe_1_7_5_n61), .B1(
        pe_1_7_5_N84), .B2(pe_1_7_5_n27), .C1(pe_1_7_5_N76), .C2(pe_1_7_5_n28), 
        .ZN(pe_1_7_5_n29) );
  INV_X1 pe_1_7_5_U46 ( .A(pe_1_7_5_n29), .ZN(pe_1_7_5_n72) );
  XNOR2_X1 pe_1_7_5_U45 ( .A(pe_1_7_5_n67), .B(int_data_res_7__5__0_), .ZN(
        pe_1_7_5_N70) );
  AOI222_X1 pe_1_7_5_U44 ( .A1(i_data_acc[16]), .A2(pe_1_7_5_n61), .B1(
        pe_1_7_5_n1), .B2(pe_1_7_5_n27), .C1(pe_1_7_5_N70), .C2(pe_1_7_5_n28), 
        .ZN(pe_1_7_5_n35) );
  INV_X1 pe_1_7_5_U43 ( .A(pe_1_7_5_n35), .ZN(pe_1_7_5_n78) );
  NAND2_X1 pe_1_7_5_U42 ( .A1(pe_1_7_5_int_data_0_), .A2(pe_1_7_5_n3), .ZN(
        pe_1_7_5_sub_81_carry[1]) );
  INV_X1 pe_1_7_5_U41 ( .A(pe_1_7_5_int_data_1_), .ZN(pe_1_7_5_n68) );
  INV_X1 pe_1_7_5_U40 ( .A(pe_1_7_5_int_data_2_), .ZN(pe_1_7_5_n69) );
  AND2_X1 pe_1_7_5_U39 ( .A1(pe_1_7_5_int_data_0_), .A2(int_data_res_7__5__0_), 
        .ZN(pe_1_7_5_n2) );
  AOI222_X1 pe_1_7_5_U38 ( .A1(pe_1_7_5_n61), .A2(i_data_acc[23]), .B1(
        pe_1_7_5_N85), .B2(pe_1_7_5_n27), .C1(pe_1_7_5_N77), .C2(pe_1_7_5_n28), 
        .ZN(pe_1_7_5_n26) );
  INV_X1 pe_1_7_5_U37 ( .A(pe_1_7_5_n26), .ZN(pe_1_7_5_n71) );
  NOR3_X1 pe_1_7_5_U36 ( .A1(pe_1_7_5_n58), .A2(pe_1_7_5_n62), .A3(int_ckg[2]), 
        .ZN(pe_1_7_5_n36) );
  OR2_X1 pe_1_7_5_U35 ( .A1(pe_1_7_5_n36), .A2(pe_1_7_5_n61), .ZN(pe_1_7_5_N90) );
  AND2_X1 pe_1_7_5_U34 ( .A1(int_data_x_7__5__2_), .A2(n30), .ZN(
        pe_1_7_5_int_data_2_) );
  AND2_X1 pe_1_7_5_U33 ( .A1(int_data_x_7__5__1_), .A2(n30), .ZN(
        pe_1_7_5_int_data_1_) );
  INV_X1 pe_1_7_5_U32 ( .A(n42), .ZN(pe_1_7_5_n60) );
  BUF_X1 pe_1_7_5_U31 ( .A(n64), .Z(pe_1_7_5_n61) );
  AND2_X1 pe_1_7_5_U30 ( .A1(int_data_x_7__5__3_), .A2(n30), .ZN(
        pe_1_7_5_int_data_3_) );
  AND2_X1 pe_1_7_5_U29 ( .A1(int_data_x_7__5__0_), .A2(n30), .ZN(
        pe_1_7_5_int_data_0_) );
  INV_X1 pe_1_7_5_U28 ( .A(n36), .ZN(pe_1_7_5_n59) );
  NAND2_X1 pe_1_7_5_U27 ( .A1(pe_1_7_5_n44), .A2(pe_1_7_5_n59), .ZN(
        pe_1_7_5_n41) );
  AND3_X1 pe_1_7_5_U26 ( .A1(n78), .A2(pe_1_7_5_n60), .A3(n55), .ZN(
        pe_1_7_5_n44) );
  INV_X1 pe_1_7_5_U25 ( .A(pe_1_7_5_int_data_3_), .ZN(pe_1_7_5_n70) );
  NOR2_X1 pe_1_7_5_U24 ( .A1(pe_1_7_5_n64), .A2(n55), .ZN(pe_1_7_5_n43) );
  NOR2_X1 pe_1_7_5_U23 ( .A1(pe_1_7_5_n57), .A2(pe_1_7_5_n61), .ZN(
        pe_1_7_5_n28) );
  NOR2_X1 pe_1_7_5_U22 ( .A1(n22), .A2(pe_1_7_5_n61), .ZN(pe_1_7_5_n27) );
  INV_X1 pe_1_7_5_U21 ( .A(pe_1_7_5_int_data_0_), .ZN(pe_1_7_5_n67) );
  INV_X1 pe_1_7_5_U20 ( .A(pe_1_7_5_n41), .ZN(pe_1_7_5_n84) );
  INV_X1 pe_1_7_5_U19 ( .A(pe_1_7_5_n37), .ZN(pe_1_7_5_n82) );
  INV_X1 pe_1_7_5_U18 ( .A(pe_1_7_5_n38), .ZN(pe_1_7_5_n81) );
  INV_X1 pe_1_7_5_U17 ( .A(pe_1_7_5_n39), .ZN(pe_1_7_5_n80) );
  NOR2_X1 pe_1_7_5_U16 ( .A1(pe_1_7_5_n63), .A2(pe_1_7_5_n42), .ZN(
        pe_1_7_5_N59) );
  NOR2_X1 pe_1_7_5_U15 ( .A1(pe_1_7_5_n63), .A2(pe_1_7_5_n41), .ZN(
        pe_1_7_5_N60) );
  NOR2_X1 pe_1_7_5_U14 ( .A1(pe_1_7_5_n63), .A2(pe_1_7_5_n38), .ZN(
        pe_1_7_5_N63) );
  NOR2_X1 pe_1_7_5_U13 ( .A1(pe_1_7_5_n63), .A2(pe_1_7_5_n40), .ZN(
        pe_1_7_5_N61) );
  NOR2_X1 pe_1_7_5_U12 ( .A1(pe_1_7_5_n63), .A2(pe_1_7_5_n39), .ZN(
        pe_1_7_5_N62) );
  NOR2_X1 pe_1_7_5_U11 ( .A1(pe_1_7_5_n37), .A2(pe_1_7_5_n63), .ZN(
        pe_1_7_5_N64) );
  NAND2_X1 pe_1_7_5_U10 ( .A1(pe_1_7_5_n44), .A2(n36), .ZN(pe_1_7_5_n42) );
  BUF_X1 pe_1_7_5_U9 ( .A(n36), .Z(pe_1_7_5_n55) );
  INV_X1 pe_1_7_5_U8 ( .A(pe_1_7_5_n63), .ZN(pe_1_7_5_n62) );
  BUF_X1 pe_1_7_5_U7 ( .A(n36), .Z(pe_1_7_5_n56) );
  INV_X1 pe_1_7_5_U6 ( .A(pe_1_7_5_n42), .ZN(pe_1_7_5_n83) );
  INV_X1 pe_1_7_5_U5 ( .A(pe_1_7_5_n40), .ZN(pe_1_7_5_n79) );
  INV_X2 pe_1_7_5_U4 ( .A(n86), .ZN(pe_1_7_5_n66) );
  XOR2_X1 pe_1_7_5_U3 ( .A(pe_1_7_5_int_data_0_), .B(int_data_res_7__5__0_), 
        .Z(pe_1_7_5_n1) );
  DFFR_X1 pe_1_7_5_int_q_acc_reg_0_ ( .D(pe_1_7_5_n78), .CK(pe_1_7_5_net2794), 
        .RN(pe_1_7_5_n66), .Q(int_data_res_7__5__0_), .QN(pe_1_7_5_n3) );
  DFFR_X1 pe_1_7_5_int_q_reg_v_reg_0__0_ ( .D(i_data_conv_v[8]), .CK(
        pe_1_7_5_net2764), .RN(pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_v[20]) );
  DFFR_X1 pe_1_7_5_int_q_reg_v_reg_0__1_ ( .D(i_data_conv_v[9]), .CK(
        pe_1_7_5_net2764), .RN(pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_v[21]) );
  DFFR_X1 pe_1_7_5_int_q_reg_v_reg_0__2_ ( .D(i_data_conv_v[10]), .CK(
        pe_1_7_5_net2764), .RN(pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_v[22]) );
  DFFR_X1 pe_1_7_5_int_q_reg_v_reg_0__3_ ( .D(i_data_conv_v[11]), .CK(
        pe_1_7_5_net2764), .RN(pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_v[23]) );
  DFFR_X1 pe_1_7_5_int_q_reg_v_reg_1__0_ ( .D(i_data_conv_v[8]), .CK(
        pe_1_7_5_net2769), .RN(pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_v[16]) );
  DFFR_X1 pe_1_7_5_int_q_reg_v_reg_1__1_ ( .D(i_data_conv_v[9]), .CK(
        pe_1_7_5_net2769), .RN(pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_v[17]) );
  DFFR_X1 pe_1_7_5_int_q_reg_v_reg_1__2_ ( .D(i_data_conv_v[10]), .CK(
        pe_1_7_5_net2769), .RN(pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_v[18]) );
  DFFR_X1 pe_1_7_5_int_q_reg_v_reg_1__3_ ( .D(i_data_conv_v[11]), .CK(
        pe_1_7_5_net2769), .RN(pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_v[19]) );
  DFFR_X1 pe_1_7_5_int_q_reg_v_reg_2__0_ ( .D(i_data_conv_v[8]), .CK(
        pe_1_7_5_net2774), .RN(pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_v[12]) );
  DFFR_X1 pe_1_7_5_int_q_reg_v_reg_2__1_ ( .D(i_data_conv_v[9]), .CK(
        pe_1_7_5_net2774), .RN(pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_v[13]) );
  DFFR_X1 pe_1_7_5_int_q_reg_v_reg_2__2_ ( .D(i_data_conv_v[10]), .CK(
        pe_1_7_5_net2774), .RN(pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_v[14]) );
  DFFR_X1 pe_1_7_5_int_q_reg_v_reg_2__3_ ( .D(i_data_conv_v[11]), .CK(
        pe_1_7_5_net2774), .RN(pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_v[15]) );
  DFFR_X1 pe_1_7_5_int_q_reg_v_reg_3__0_ ( .D(i_data_conv_v[8]), .CK(
        pe_1_7_5_net2779), .RN(pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_v[8]) );
  DFFR_X1 pe_1_7_5_int_q_reg_v_reg_3__1_ ( .D(i_data_conv_v[9]), .CK(
        pe_1_7_5_net2779), .RN(pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_v[9]) );
  DFFR_X1 pe_1_7_5_int_q_reg_v_reg_3__2_ ( .D(i_data_conv_v[10]), .CK(
        pe_1_7_5_net2779), .RN(pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_v[10]) );
  DFFR_X1 pe_1_7_5_int_q_reg_v_reg_3__3_ ( .D(i_data_conv_v[11]), .CK(
        pe_1_7_5_net2779), .RN(pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_v[11]) );
  DFFR_X1 pe_1_7_5_int_q_reg_v_reg_4__0_ ( .D(i_data_conv_v[8]), .CK(
        pe_1_7_5_net2784), .RN(pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_v[4]) );
  DFFR_X1 pe_1_7_5_int_q_reg_v_reg_4__1_ ( .D(i_data_conv_v[9]), .CK(
        pe_1_7_5_net2784), .RN(pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_v[5]) );
  DFFR_X1 pe_1_7_5_int_q_reg_v_reg_4__2_ ( .D(i_data_conv_v[10]), .CK(
        pe_1_7_5_net2784), .RN(pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_v[6]) );
  DFFR_X1 pe_1_7_5_int_q_reg_v_reg_4__3_ ( .D(i_data_conv_v[11]), .CK(
        pe_1_7_5_net2784), .RN(pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_v[7]) );
  DFFR_X1 pe_1_7_5_int_q_reg_v_reg_5__0_ ( .D(i_data_conv_v[8]), .CK(
        pe_1_7_5_net2789), .RN(pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_v[0]) );
  DFFR_X1 pe_1_7_5_int_q_reg_v_reg_5__1_ ( .D(i_data_conv_v[9]), .CK(
        pe_1_7_5_net2789), .RN(pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_v[1]) );
  DFFR_X1 pe_1_7_5_int_q_reg_v_reg_5__2_ ( .D(i_data_conv_v[10]), .CK(
        pe_1_7_5_net2789), .RN(pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_v[2]) );
  DFFR_X1 pe_1_7_5_int_q_reg_v_reg_5__3_ ( .D(i_data_conv_v[11]), .CK(
        pe_1_7_5_net2789), .RN(pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_7_5_int_q_reg_h_reg_0__0_ ( .D(int_data_x_7__6__0_), .SI(
        i_data_conv_v[8]), .SE(pe_1_7_5_n62), .CK(pe_1_7_5_net2733), .RN(
        pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_7_5_int_q_reg_h_reg_0__1_ ( .D(int_data_x_7__6__1_), .SI(
        i_data_conv_v[9]), .SE(pe_1_7_5_n62), .CK(pe_1_7_5_net2733), .RN(
        pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_7_5_int_q_reg_h_reg_0__2_ ( .D(int_data_x_7__6__2_), .SI(
        i_data_conv_v[10]), .SE(pe_1_7_5_n62), .CK(pe_1_7_5_net2733), .RN(
        pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_7_5_int_q_reg_h_reg_0__3_ ( .D(int_data_x_7__6__3_), .SI(
        i_data_conv_v[11]), .SE(pe_1_7_5_n62), .CK(pe_1_7_5_net2733), .RN(
        pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_7_5_int_q_reg_h_reg_1__0_ ( .D(int_data_x_7__6__0_), .SI(
        i_data_conv_v[8]), .SE(pe_1_7_5_n62), .CK(pe_1_7_5_net2739), .RN(
        pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_7_5_int_q_reg_h_reg_1__1_ ( .D(int_data_x_7__6__1_), .SI(
        i_data_conv_v[9]), .SE(pe_1_7_5_n62), .CK(pe_1_7_5_net2739), .RN(
        pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_7_5_int_q_reg_h_reg_1__2_ ( .D(int_data_x_7__6__2_), .SI(
        i_data_conv_v[10]), .SE(pe_1_7_5_n62), .CK(pe_1_7_5_net2739), .RN(
        pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_7_5_int_q_reg_h_reg_1__3_ ( .D(int_data_x_7__6__3_), .SI(
        i_data_conv_v[11]), .SE(pe_1_7_5_n62), .CK(pe_1_7_5_net2739), .RN(
        pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_7_5_int_q_reg_h_reg_2__0_ ( .D(int_data_x_7__6__0_), .SI(
        i_data_conv_v[8]), .SE(pe_1_7_5_n62), .CK(pe_1_7_5_net2744), .RN(
        pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_7_5_int_q_reg_h_reg_2__1_ ( .D(int_data_x_7__6__1_), .SI(
        i_data_conv_v[9]), .SE(pe_1_7_5_n62), .CK(pe_1_7_5_net2744), .RN(
        pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_7_5_int_q_reg_h_reg_2__2_ ( .D(int_data_x_7__6__2_), .SI(
        i_data_conv_v[10]), .SE(pe_1_7_5_n62), .CK(pe_1_7_5_net2744), .RN(
        pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_7_5_int_q_reg_h_reg_2__3_ ( .D(int_data_x_7__6__3_), .SI(
        i_data_conv_v[11]), .SE(pe_1_7_5_n62), .CK(pe_1_7_5_net2744), .RN(
        pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_7_5_int_q_reg_h_reg_3__0_ ( .D(int_data_x_7__6__0_), .SI(
        i_data_conv_v[8]), .SE(pe_1_7_5_n62), .CK(pe_1_7_5_net2749), .RN(
        pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_7_5_int_q_reg_h_reg_3__1_ ( .D(int_data_x_7__6__1_), .SI(
        i_data_conv_v[9]), .SE(pe_1_7_5_n62), .CK(pe_1_7_5_net2749), .RN(
        pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_7_5_int_q_reg_h_reg_3__2_ ( .D(int_data_x_7__6__2_), .SI(
        i_data_conv_v[10]), .SE(pe_1_7_5_n62), .CK(pe_1_7_5_net2749), .RN(
        pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_7_5_int_q_reg_h_reg_3__3_ ( .D(int_data_x_7__6__3_), .SI(
        i_data_conv_v[11]), .SE(pe_1_7_5_n62), .CK(pe_1_7_5_net2749), .RN(
        pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_7_5_int_q_reg_h_reg_4__0_ ( .D(int_data_x_7__6__0_), .SI(
        i_data_conv_v[8]), .SE(pe_1_7_5_n62), .CK(pe_1_7_5_net2754), .RN(
        pe_1_7_5_n66), .Q(pe_1_7_5_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_7_5_int_q_reg_h_reg_4__1_ ( .D(int_data_x_7__6__1_), .SI(
        i_data_conv_v[9]), .SE(n70), .CK(pe_1_7_5_net2754), .RN(pe_1_7_5_n66), 
        .Q(pe_1_7_5_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_7_5_int_q_reg_h_reg_4__2_ ( .D(int_data_x_7__6__2_), .SI(
        i_data_conv_v[10]), .SE(n70), .CK(pe_1_7_5_net2754), .RN(pe_1_7_5_n66), 
        .Q(pe_1_7_5_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_7_5_int_q_reg_h_reg_4__3_ ( .D(int_data_x_7__6__3_), .SI(
        i_data_conv_v[11]), .SE(n70), .CK(pe_1_7_5_net2754), .RN(pe_1_7_5_n66), 
        .Q(pe_1_7_5_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_7_5_int_q_reg_h_reg_5__0_ ( .D(int_data_x_7__6__0_), .SI(
        i_data_conv_v[8]), .SE(n70), .CK(pe_1_7_5_net2759), .RN(pe_1_7_5_n66), 
        .Q(pe_1_7_5_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_7_5_int_q_reg_h_reg_5__1_ ( .D(int_data_x_7__6__1_), .SI(
        i_data_conv_v[9]), .SE(n70), .CK(pe_1_7_5_net2759), .RN(pe_1_7_5_n66), 
        .Q(pe_1_7_5_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_7_5_int_q_reg_h_reg_5__2_ ( .D(int_data_x_7__6__2_), .SI(
        i_data_conv_v[10]), .SE(n70), .CK(pe_1_7_5_net2759), .RN(pe_1_7_5_n66), 
        .Q(pe_1_7_5_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_7_5_int_q_reg_h_reg_5__3_ ( .D(int_data_x_7__6__3_), .SI(
        i_data_conv_v[11]), .SE(n70), .CK(pe_1_7_5_net2759), .RN(pe_1_7_5_n66), 
        .Q(pe_1_7_5_int_q_reg_h[3]) );
  FA_X1 pe_1_7_5_sub_81_U2_7 ( .A(int_data_res_7__5__7_), .B(pe_1_7_5_n70), 
        .CI(pe_1_7_5_sub_81_carry[7]), .S(pe_1_7_5_N77) );
  FA_X1 pe_1_7_5_sub_81_U2_6 ( .A(int_data_res_7__5__6_), .B(pe_1_7_5_n70), 
        .CI(pe_1_7_5_sub_81_carry[6]), .CO(pe_1_7_5_sub_81_carry[7]), .S(
        pe_1_7_5_N76) );
  FA_X1 pe_1_7_5_sub_81_U2_5 ( .A(int_data_res_7__5__5_), .B(pe_1_7_5_n70), 
        .CI(pe_1_7_5_sub_81_carry[5]), .CO(pe_1_7_5_sub_81_carry[6]), .S(
        pe_1_7_5_N75) );
  FA_X1 pe_1_7_5_sub_81_U2_4 ( .A(int_data_res_7__5__4_), .B(pe_1_7_5_n70), 
        .CI(pe_1_7_5_sub_81_carry[4]), .CO(pe_1_7_5_sub_81_carry[5]), .S(
        pe_1_7_5_N74) );
  FA_X1 pe_1_7_5_sub_81_U2_3 ( .A(int_data_res_7__5__3_), .B(pe_1_7_5_n70), 
        .CI(pe_1_7_5_sub_81_carry[3]), .CO(pe_1_7_5_sub_81_carry[4]), .S(
        pe_1_7_5_N73) );
  FA_X1 pe_1_7_5_sub_81_U2_2 ( .A(int_data_res_7__5__2_), .B(pe_1_7_5_n69), 
        .CI(pe_1_7_5_sub_81_carry[2]), .CO(pe_1_7_5_sub_81_carry[3]), .S(
        pe_1_7_5_N72) );
  FA_X1 pe_1_7_5_sub_81_U2_1 ( .A(int_data_res_7__5__1_), .B(pe_1_7_5_n68), 
        .CI(pe_1_7_5_sub_81_carry[1]), .CO(pe_1_7_5_sub_81_carry[2]), .S(
        pe_1_7_5_N71) );
  FA_X1 pe_1_7_5_add_83_U1_7 ( .A(int_data_res_7__5__7_), .B(
        pe_1_7_5_int_data_3_), .CI(pe_1_7_5_add_83_carry[7]), .S(pe_1_7_5_N85)
         );
  FA_X1 pe_1_7_5_add_83_U1_6 ( .A(int_data_res_7__5__6_), .B(
        pe_1_7_5_int_data_3_), .CI(pe_1_7_5_add_83_carry[6]), .CO(
        pe_1_7_5_add_83_carry[7]), .S(pe_1_7_5_N84) );
  FA_X1 pe_1_7_5_add_83_U1_5 ( .A(int_data_res_7__5__5_), .B(
        pe_1_7_5_int_data_3_), .CI(pe_1_7_5_add_83_carry[5]), .CO(
        pe_1_7_5_add_83_carry[6]), .S(pe_1_7_5_N83) );
  FA_X1 pe_1_7_5_add_83_U1_4 ( .A(int_data_res_7__5__4_), .B(
        pe_1_7_5_int_data_3_), .CI(pe_1_7_5_add_83_carry[4]), .CO(
        pe_1_7_5_add_83_carry[5]), .S(pe_1_7_5_N82) );
  FA_X1 pe_1_7_5_add_83_U1_3 ( .A(int_data_res_7__5__3_), .B(
        pe_1_7_5_int_data_3_), .CI(pe_1_7_5_add_83_carry[3]), .CO(
        pe_1_7_5_add_83_carry[4]), .S(pe_1_7_5_N81) );
  FA_X1 pe_1_7_5_add_83_U1_2 ( .A(int_data_res_7__5__2_), .B(
        pe_1_7_5_int_data_2_), .CI(pe_1_7_5_add_83_carry[2]), .CO(
        pe_1_7_5_add_83_carry[3]), .S(pe_1_7_5_N80) );
  FA_X1 pe_1_7_5_add_83_U1_1 ( .A(int_data_res_7__5__1_), .B(
        pe_1_7_5_int_data_1_), .CI(pe_1_7_5_n2), .CO(pe_1_7_5_add_83_carry[2]), 
        .S(pe_1_7_5_N79) );
  NAND3_X1 pe_1_7_5_U56 ( .A1(n36), .A2(pe_1_7_5_n43), .A3(n42), .ZN(
        pe_1_7_5_n40) );
  NAND3_X1 pe_1_7_5_U55 ( .A1(pe_1_7_5_n43), .A2(pe_1_7_5_n59), .A3(n42), .ZN(
        pe_1_7_5_n39) );
  NAND3_X1 pe_1_7_5_U54 ( .A1(pe_1_7_5_n43), .A2(pe_1_7_5_n60), .A3(n36), .ZN(
        pe_1_7_5_n38) );
  NAND3_X1 pe_1_7_5_U53 ( .A1(pe_1_7_5_n59), .A2(pe_1_7_5_n60), .A3(
        pe_1_7_5_n43), .ZN(pe_1_7_5_n37) );
  DFFR_X1 pe_1_7_5_int_q_acc_reg_6_ ( .D(pe_1_7_5_n72), .CK(pe_1_7_5_net2794), 
        .RN(pe_1_7_5_n65), .Q(int_data_res_7__5__6_) );
  DFFR_X1 pe_1_7_5_int_q_acc_reg_5_ ( .D(pe_1_7_5_n73), .CK(pe_1_7_5_net2794), 
        .RN(pe_1_7_5_n65), .Q(int_data_res_7__5__5_) );
  DFFR_X1 pe_1_7_5_int_q_acc_reg_4_ ( .D(pe_1_7_5_n74), .CK(pe_1_7_5_net2794), 
        .RN(pe_1_7_5_n65), .Q(int_data_res_7__5__4_) );
  DFFR_X1 pe_1_7_5_int_q_acc_reg_3_ ( .D(pe_1_7_5_n75), .CK(pe_1_7_5_net2794), 
        .RN(pe_1_7_5_n65), .Q(int_data_res_7__5__3_) );
  DFFR_X1 pe_1_7_5_int_q_acc_reg_2_ ( .D(pe_1_7_5_n76), .CK(pe_1_7_5_net2794), 
        .RN(pe_1_7_5_n65), .Q(int_data_res_7__5__2_) );
  DFFR_X1 pe_1_7_5_int_q_acc_reg_1_ ( .D(pe_1_7_5_n77), .CK(pe_1_7_5_net2794), 
        .RN(pe_1_7_5_n65), .Q(int_data_res_7__5__1_) );
  DFFR_X1 pe_1_7_5_int_q_acc_reg_7_ ( .D(pe_1_7_5_n71), .CK(pe_1_7_5_net2794), 
        .RN(pe_1_7_5_n65), .Q(int_data_res_7__5__7_) );
  CLKGATETST_X1 pe_1_7_5_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_7_5_n82), .SE(1'b0), .GCK(pe_1_7_5_net2733) );
  CLKGATETST_X1 pe_1_7_5_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_7_5_n81), .SE(1'b0), .GCK(pe_1_7_5_net2739) );
  CLKGATETST_X1 pe_1_7_5_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_7_5_n80), .SE(1'b0), .GCK(pe_1_7_5_net2744) );
  CLKGATETST_X1 pe_1_7_5_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_7_5_n79), .SE(1'b0), .GCK(pe_1_7_5_net2749) );
  CLKGATETST_X1 pe_1_7_5_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_7_5_n84), .SE(1'b0), .GCK(pe_1_7_5_net2754) );
  CLKGATETST_X1 pe_1_7_5_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_7_5_n83), .SE(1'b0), .GCK(pe_1_7_5_net2759) );
  CLKGATETST_X1 pe_1_7_5_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_7_5_N64), .SE(1'b0), .GCK(pe_1_7_5_net2764) );
  CLKGATETST_X1 pe_1_7_5_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_7_5_N63), .SE(1'b0), .GCK(pe_1_7_5_net2769) );
  CLKGATETST_X1 pe_1_7_5_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_7_5_N62), .SE(1'b0), .GCK(pe_1_7_5_net2774) );
  CLKGATETST_X1 pe_1_7_5_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_7_5_N61), .SE(1'b0), .GCK(pe_1_7_5_net2779) );
  CLKGATETST_X1 pe_1_7_5_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_7_5_N60), .SE(1'b0), .GCK(pe_1_7_5_net2784) );
  CLKGATETST_X1 pe_1_7_5_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_7_5_N59), .SE(1'b0), .GCK(pe_1_7_5_net2789) );
  CLKGATETST_X1 pe_1_7_5_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_7_5_N90), .SE(1'b0), .GCK(pe_1_7_5_net2794) );
  CLKBUF_X1 pe_1_7_6_U107 ( .A(pe_1_7_6_n67), .Z(pe_1_7_6_n66) );
  INV_X1 pe_1_7_6_U106 ( .A(n78), .ZN(pe_1_7_6_n65) );
  INV_X1 pe_1_7_6_U105 ( .A(n70), .ZN(pe_1_7_6_n64) );
  INV_X1 pe_1_7_6_U104 ( .A(pe_1_7_6_n61), .ZN(pe_1_7_6_n60) );
  INV_X1 pe_1_7_6_U103 ( .A(n30), .ZN(pe_1_7_6_n58) );
  INV_X1 pe_1_7_6_U102 ( .A(n22), .ZN(pe_1_7_6_n57) );
  MUX2_X1 pe_1_7_6_U101 ( .A(pe_1_7_6_n54), .B(pe_1_7_6_n51), .S(n55), .Z(
        int_data_x_7__6__3_) );
  MUX2_X1 pe_1_7_6_U100 ( .A(pe_1_7_6_n53), .B(pe_1_7_6_n52), .S(pe_1_7_6_n60), 
        .Z(pe_1_7_6_n54) );
  MUX2_X1 pe_1_7_6_U99 ( .A(pe_1_7_6_int_q_reg_h[23]), .B(
        pe_1_7_6_int_q_reg_h[19]), .S(pe_1_7_6_n56), .Z(pe_1_7_6_n53) );
  MUX2_X1 pe_1_7_6_U98 ( .A(pe_1_7_6_int_q_reg_h[15]), .B(
        pe_1_7_6_int_q_reg_h[11]), .S(pe_1_7_6_n56), .Z(pe_1_7_6_n52) );
  MUX2_X1 pe_1_7_6_U97 ( .A(pe_1_7_6_int_q_reg_h[7]), .B(
        pe_1_7_6_int_q_reg_h[3]), .S(pe_1_7_6_n56), .Z(pe_1_7_6_n51) );
  MUX2_X1 pe_1_7_6_U96 ( .A(pe_1_7_6_n50), .B(pe_1_7_6_n47), .S(n55), .Z(
        int_data_x_7__6__2_) );
  MUX2_X1 pe_1_7_6_U95 ( .A(pe_1_7_6_n49), .B(pe_1_7_6_n48), .S(pe_1_7_6_n60), 
        .Z(pe_1_7_6_n50) );
  MUX2_X1 pe_1_7_6_U94 ( .A(pe_1_7_6_int_q_reg_h[22]), .B(
        pe_1_7_6_int_q_reg_h[18]), .S(pe_1_7_6_n56), .Z(pe_1_7_6_n49) );
  MUX2_X1 pe_1_7_6_U93 ( .A(pe_1_7_6_int_q_reg_h[14]), .B(
        pe_1_7_6_int_q_reg_h[10]), .S(pe_1_7_6_n56), .Z(pe_1_7_6_n48) );
  MUX2_X1 pe_1_7_6_U92 ( .A(pe_1_7_6_int_q_reg_h[6]), .B(
        pe_1_7_6_int_q_reg_h[2]), .S(pe_1_7_6_n56), .Z(pe_1_7_6_n47) );
  MUX2_X1 pe_1_7_6_U91 ( .A(pe_1_7_6_n46), .B(pe_1_7_6_n24), .S(n55), .Z(
        int_data_x_7__6__1_) );
  MUX2_X1 pe_1_7_6_U90 ( .A(pe_1_7_6_n45), .B(pe_1_7_6_n25), .S(pe_1_7_6_n60), 
        .Z(pe_1_7_6_n46) );
  MUX2_X1 pe_1_7_6_U89 ( .A(pe_1_7_6_int_q_reg_h[21]), .B(
        pe_1_7_6_int_q_reg_h[17]), .S(pe_1_7_6_n56), .Z(pe_1_7_6_n45) );
  MUX2_X1 pe_1_7_6_U88 ( .A(pe_1_7_6_int_q_reg_h[13]), .B(
        pe_1_7_6_int_q_reg_h[9]), .S(pe_1_7_6_n56), .Z(pe_1_7_6_n25) );
  MUX2_X1 pe_1_7_6_U87 ( .A(pe_1_7_6_int_q_reg_h[5]), .B(
        pe_1_7_6_int_q_reg_h[1]), .S(pe_1_7_6_n56), .Z(pe_1_7_6_n24) );
  MUX2_X1 pe_1_7_6_U86 ( .A(pe_1_7_6_n23), .B(pe_1_7_6_n20), .S(n55), .Z(
        int_data_x_7__6__0_) );
  MUX2_X1 pe_1_7_6_U85 ( .A(pe_1_7_6_n22), .B(pe_1_7_6_n21), .S(pe_1_7_6_n60), 
        .Z(pe_1_7_6_n23) );
  MUX2_X1 pe_1_7_6_U84 ( .A(pe_1_7_6_int_q_reg_h[20]), .B(
        pe_1_7_6_int_q_reg_h[16]), .S(pe_1_7_6_n56), .Z(pe_1_7_6_n22) );
  MUX2_X1 pe_1_7_6_U83 ( .A(pe_1_7_6_int_q_reg_h[12]), .B(
        pe_1_7_6_int_q_reg_h[8]), .S(pe_1_7_6_n56), .Z(pe_1_7_6_n21) );
  MUX2_X1 pe_1_7_6_U82 ( .A(pe_1_7_6_int_q_reg_h[4]), .B(
        pe_1_7_6_int_q_reg_h[0]), .S(pe_1_7_6_n56), .Z(pe_1_7_6_n20) );
  MUX2_X1 pe_1_7_6_U81 ( .A(pe_1_7_6_n19), .B(pe_1_7_6_n16), .S(n55), .Z(
        int_data_y_7__6__3_) );
  MUX2_X1 pe_1_7_6_U80 ( .A(pe_1_7_6_n18), .B(pe_1_7_6_n17), .S(pe_1_7_6_n60), 
        .Z(pe_1_7_6_n19) );
  MUX2_X1 pe_1_7_6_U79 ( .A(pe_1_7_6_int_q_reg_v[23]), .B(
        pe_1_7_6_int_q_reg_v[19]), .S(pe_1_7_6_n55), .Z(pe_1_7_6_n18) );
  MUX2_X1 pe_1_7_6_U78 ( .A(pe_1_7_6_int_q_reg_v[15]), .B(
        pe_1_7_6_int_q_reg_v[11]), .S(pe_1_7_6_n55), .Z(pe_1_7_6_n17) );
  MUX2_X1 pe_1_7_6_U77 ( .A(pe_1_7_6_int_q_reg_v[7]), .B(
        pe_1_7_6_int_q_reg_v[3]), .S(pe_1_7_6_n55), .Z(pe_1_7_6_n16) );
  MUX2_X1 pe_1_7_6_U76 ( .A(pe_1_7_6_n15), .B(pe_1_7_6_n12), .S(n55), .Z(
        int_data_y_7__6__2_) );
  MUX2_X1 pe_1_7_6_U75 ( .A(pe_1_7_6_n14), .B(pe_1_7_6_n13), .S(pe_1_7_6_n60), 
        .Z(pe_1_7_6_n15) );
  MUX2_X1 pe_1_7_6_U74 ( .A(pe_1_7_6_int_q_reg_v[22]), .B(
        pe_1_7_6_int_q_reg_v[18]), .S(pe_1_7_6_n55), .Z(pe_1_7_6_n14) );
  MUX2_X1 pe_1_7_6_U73 ( .A(pe_1_7_6_int_q_reg_v[14]), .B(
        pe_1_7_6_int_q_reg_v[10]), .S(pe_1_7_6_n55), .Z(pe_1_7_6_n13) );
  MUX2_X1 pe_1_7_6_U72 ( .A(pe_1_7_6_int_q_reg_v[6]), .B(
        pe_1_7_6_int_q_reg_v[2]), .S(pe_1_7_6_n55), .Z(pe_1_7_6_n12) );
  MUX2_X1 pe_1_7_6_U71 ( .A(pe_1_7_6_n11), .B(pe_1_7_6_n8), .S(n55), .Z(
        int_data_y_7__6__1_) );
  MUX2_X1 pe_1_7_6_U70 ( .A(pe_1_7_6_n10), .B(pe_1_7_6_n9), .S(pe_1_7_6_n60), 
        .Z(pe_1_7_6_n11) );
  MUX2_X1 pe_1_7_6_U69 ( .A(pe_1_7_6_int_q_reg_v[21]), .B(
        pe_1_7_6_int_q_reg_v[17]), .S(pe_1_7_6_n55), .Z(pe_1_7_6_n10) );
  MUX2_X1 pe_1_7_6_U68 ( .A(pe_1_7_6_int_q_reg_v[13]), .B(
        pe_1_7_6_int_q_reg_v[9]), .S(pe_1_7_6_n55), .Z(pe_1_7_6_n9) );
  MUX2_X1 pe_1_7_6_U67 ( .A(pe_1_7_6_int_q_reg_v[5]), .B(
        pe_1_7_6_int_q_reg_v[1]), .S(pe_1_7_6_n55), .Z(pe_1_7_6_n8) );
  MUX2_X1 pe_1_7_6_U66 ( .A(pe_1_7_6_n7), .B(pe_1_7_6_n4), .S(n55), .Z(
        int_data_y_7__6__0_) );
  MUX2_X1 pe_1_7_6_U65 ( .A(pe_1_7_6_n6), .B(pe_1_7_6_n5), .S(pe_1_7_6_n60), 
        .Z(pe_1_7_6_n7) );
  MUX2_X1 pe_1_7_6_U64 ( .A(pe_1_7_6_int_q_reg_v[20]), .B(
        pe_1_7_6_int_q_reg_v[16]), .S(pe_1_7_6_n55), .Z(pe_1_7_6_n6) );
  MUX2_X1 pe_1_7_6_U63 ( .A(pe_1_7_6_int_q_reg_v[12]), .B(
        pe_1_7_6_int_q_reg_v[8]), .S(pe_1_7_6_n55), .Z(pe_1_7_6_n5) );
  MUX2_X1 pe_1_7_6_U62 ( .A(pe_1_7_6_int_q_reg_v[4]), .B(
        pe_1_7_6_int_q_reg_v[0]), .S(pe_1_7_6_n55), .Z(pe_1_7_6_n4) );
  AOI222_X1 pe_1_7_6_U61 ( .A1(i_data_acc[9]), .A2(pe_1_7_6_n62), .B1(
        pe_1_7_6_N79), .B2(pe_1_7_6_n27), .C1(pe_1_7_6_N71), .C2(pe_1_7_6_n28), 
        .ZN(pe_1_7_6_n34) );
  INV_X1 pe_1_7_6_U60 ( .A(pe_1_7_6_n34), .ZN(pe_1_7_6_n78) );
  AOI222_X1 pe_1_7_6_U59 ( .A1(i_data_acc[10]), .A2(pe_1_7_6_n62), .B1(
        pe_1_7_6_N80), .B2(pe_1_7_6_n27), .C1(pe_1_7_6_N72), .C2(pe_1_7_6_n28), 
        .ZN(pe_1_7_6_n33) );
  INV_X1 pe_1_7_6_U58 ( .A(pe_1_7_6_n33), .ZN(pe_1_7_6_n77) );
  AOI222_X1 pe_1_7_6_U57 ( .A1(i_data_acc[11]), .A2(pe_1_7_6_n62), .B1(
        pe_1_7_6_N81), .B2(pe_1_7_6_n27), .C1(pe_1_7_6_N73), .C2(pe_1_7_6_n28), 
        .ZN(pe_1_7_6_n32) );
  INV_X1 pe_1_7_6_U52 ( .A(pe_1_7_6_n32), .ZN(pe_1_7_6_n76) );
  AOI222_X1 pe_1_7_6_U51 ( .A1(i_data_acc[12]), .A2(pe_1_7_6_n62), .B1(
        pe_1_7_6_N82), .B2(pe_1_7_6_n27), .C1(pe_1_7_6_N74), .C2(pe_1_7_6_n28), 
        .ZN(pe_1_7_6_n31) );
  INV_X1 pe_1_7_6_U50 ( .A(pe_1_7_6_n31), .ZN(pe_1_7_6_n75) );
  AOI222_X1 pe_1_7_6_U49 ( .A1(i_data_acc[13]), .A2(pe_1_7_6_n62), .B1(
        pe_1_7_6_N83), .B2(pe_1_7_6_n27), .C1(pe_1_7_6_N75), .C2(pe_1_7_6_n28), 
        .ZN(pe_1_7_6_n30) );
  INV_X1 pe_1_7_6_U48 ( .A(pe_1_7_6_n30), .ZN(pe_1_7_6_n74) );
  AOI222_X1 pe_1_7_6_U47 ( .A1(i_data_acc[14]), .A2(pe_1_7_6_n62), .B1(
        pe_1_7_6_N84), .B2(pe_1_7_6_n27), .C1(pe_1_7_6_N76), .C2(pe_1_7_6_n28), 
        .ZN(pe_1_7_6_n29) );
  INV_X1 pe_1_7_6_U46 ( .A(pe_1_7_6_n29), .ZN(pe_1_7_6_n73) );
  XNOR2_X1 pe_1_7_6_U45 ( .A(pe_1_7_6_n68), .B(int_data_res_7__6__0_), .ZN(
        pe_1_7_6_N70) );
  AOI222_X1 pe_1_7_6_U44 ( .A1(i_data_acc[8]), .A2(pe_1_7_6_n62), .B1(
        pe_1_7_6_n1), .B2(pe_1_7_6_n27), .C1(pe_1_7_6_N70), .C2(pe_1_7_6_n28), 
        .ZN(pe_1_7_6_n35) );
  INV_X1 pe_1_7_6_U43 ( .A(pe_1_7_6_n35), .ZN(pe_1_7_6_n79) );
  NAND2_X1 pe_1_7_6_U42 ( .A1(pe_1_7_6_int_data_0_), .A2(pe_1_7_6_n3), .ZN(
        pe_1_7_6_sub_81_carry[1]) );
  INV_X1 pe_1_7_6_U41 ( .A(pe_1_7_6_int_data_1_), .ZN(pe_1_7_6_n69) );
  INV_X1 pe_1_7_6_U40 ( .A(pe_1_7_6_int_data_2_), .ZN(pe_1_7_6_n70) );
  AND2_X1 pe_1_7_6_U39 ( .A1(pe_1_7_6_int_data_0_), .A2(int_data_res_7__6__0_), 
        .ZN(pe_1_7_6_n2) );
  AOI222_X1 pe_1_7_6_U38 ( .A1(pe_1_7_6_n62), .A2(i_data_acc[15]), .B1(
        pe_1_7_6_N85), .B2(pe_1_7_6_n27), .C1(pe_1_7_6_N77), .C2(pe_1_7_6_n28), 
        .ZN(pe_1_7_6_n26) );
  INV_X1 pe_1_7_6_U37 ( .A(pe_1_7_6_n26), .ZN(pe_1_7_6_n72) );
  NOR3_X1 pe_1_7_6_U36 ( .A1(pe_1_7_6_n58), .A2(pe_1_7_6_n63), .A3(int_ckg[1]), 
        .ZN(pe_1_7_6_n36) );
  OR2_X1 pe_1_7_6_U35 ( .A1(pe_1_7_6_n36), .A2(pe_1_7_6_n62), .ZN(pe_1_7_6_N90) );
  AND2_X1 pe_1_7_6_U34 ( .A1(int_data_x_7__6__2_), .A2(n30), .ZN(
        pe_1_7_6_int_data_2_) );
  AND2_X1 pe_1_7_6_U33 ( .A1(int_data_x_7__6__1_), .A2(n30), .ZN(
        pe_1_7_6_int_data_1_) );
  INV_X1 pe_1_7_6_U32 ( .A(n42), .ZN(pe_1_7_6_n61) );
  BUF_X1 pe_1_7_6_U31 ( .A(n64), .Z(pe_1_7_6_n62) );
  AND2_X1 pe_1_7_6_U30 ( .A1(int_data_x_7__6__3_), .A2(n30), .ZN(
        pe_1_7_6_int_data_3_) );
  AND2_X1 pe_1_7_6_U29 ( .A1(int_data_x_7__6__0_), .A2(n30), .ZN(
        pe_1_7_6_int_data_0_) );
  INV_X1 pe_1_7_6_U28 ( .A(n36), .ZN(pe_1_7_6_n59) );
  NAND2_X1 pe_1_7_6_U27 ( .A1(pe_1_7_6_n44), .A2(pe_1_7_6_n59), .ZN(
        pe_1_7_6_n41) );
  AND3_X1 pe_1_7_6_U26 ( .A1(n78), .A2(pe_1_7_6_n61), .A3(n55), .ZN(
        pe_1_7_6_n44) );
  INV_X1 pe_1_7_6_U25 ( .A(pe_1_7_6_int_data_3_), .ZN(pe_1_7_6_n71) );
  NOR2_X1 pe_1_7_6_U24 ( .A1(pe_1_7_6_n65), .A2(n55), .ZN(pe_1_7_6_n43) );
  NOR2_X1 pe_1_7_6_U23 ( .A1(pe_1_7_6_n57), .A2(pe_1_7_6_n62), .ZN(
        pe_1_7_6_n28) );
  NOR2_X1 pe_1_7_6_U22 ( .A1(n22), .A2(pe_1_7_6_n62), .ZN(pe_1_7_6_n27) );
  INV_X1 pe_1_7_6_U21 ( .A(pe_1_7_6_int_data_0_), .ZN(pe_1_7_6_n68) );
  INV_X1 pe_1_7_6_U20 ( .A(pe_1_7_6_n41), .ZN(pe_1_7_6_n85) );
  INV_X1 pe_1_7_6_U19 ( .A(pe_1_7_6_n37), .ZN(pe_1_7_6_n83) );
  INV_X1 pe_1_7_6_U18 ( .A(pe_1_7_6_n38), .ZN(pe_1_7_6_n82) );
  INV_X1 pe_1_7_6_U17 ( .A(pe_1_7_6_n39), .ZN(pe_1_7_6_n81) );
  NOR2_X1 pe_1_7_6_U16 ( .A1(pe_1_7_6_n64), .A2(pe_1_7_6_n42), .ZN(
        pe_1_7_6_N59) );
  NOR2_X1 pe_1_7_6_U15 ( .A1(pe_1_7_6_n64), .A2(pe_1_7_6_n41), .ZN(
        pe_1_7_6_N60) );
  NOR2_X1 pe_1_7_6_U14 ( .A1(pe_1_7_6_n64), .A2(pe_1_7_6_n38), .ZN(
        pe_1_7_6_N63) );
  NOR2_X1 pe_1_7_6_U13 ( .A1(pe_1_7_6_n64), .A2(pe_1_7_6_n40), .ZN(
        pe_1_7_6_N61) );
  NOR2_X1 pe_1_7_6_U12 ( .A1(pe_1_7_6_n64), .A2(pe_1_7_6_n39), .ZN(
        pe_1_7_6_N62) );
  NOR2_X1 pe_1_7_6_U11 ( .A1(pe_1_7_6_n37), .A2(pe_1_7_6_n64), .ZN(
        pe_1_7_6_N64) );
  NAND2_X1 pe_1_7_6_U10 ( .A1(pe_1_7_6_n44), .A2(n36), .ZN(pe_1_7_6_n42) );
  BUF_X1 pe_1_7_6_U9 ( .A(n36), .Z(pe_1_7_6_n55) );
  INV_X1 pe_1_7_6_U8 ( .A(pe_1_7_6_n64), .ZN(pe_1_7_6_n63) );
  BUF_X1 pe_1_7_6_U7 ( .A(n36), .Z(pe_1_7_6_n56) );
  INV_X1 pe_1_7_6_U6 ( .A(pe_1_7_6_n42), .ZN(pe_1_7_6_n84) );
  INV_X1 pe_1_7_6_U5 ( .A(pe_1_7_6_n40), .ZN(pe_1_7_6_n80) );
  INV_X2 pe_1_7_6_U4 ( .A(n86), .ZN(pe_1_7_6_n67) );
  XOR2_X1 pe_1_7_6_U3 ( .A(pe_1_7_6_int_data_0_), .B(int_data_res_7__6__0_), 
        .Z(pe_1_7_6_n1) );
  DFFR_X1 pe_1_7_6_int_q_acc_reg_0_ ( .D(pe_1_7_6_n79), .CK(pe_1_7_6_net2716), 
        .RN(pe_1_7_6_n67), .Q(int_data_res_7__6__0_), .QN(pe_1_7_6_n3) );
  DFFR_X1 pe_1_7_6_int_q_reg_v_reg_0__0_ ( .D(i_data_conv_v[4]), .CK(
        pe_1_7_6_net2686), .RN(pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_v[20]) );
  DFFR_X1 pe_1_7_6_int_q_reg_v_reg_0__1_ ( .D(i_data_conv_v[5]), .CK(
        pe_1_7_6_net2686), .RN(pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_v[21]) );
  DFFR_X1 pe_1_7_6_int_q_reg_v_reg_0__2_ ( .D(i_data_conv_v[6]), .CK(
        pe_1_7_6_net2686), .RN(pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_v[22]) );
  DFFR_X1 pe_1_7_6_int_q_reg_v_reg_0__3_ ( .D(i_data_conv_v[7]), .CK(
        pe_1_7_6_net2686), .RN(pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_v[23]) );
  DFFR_X1 pe_1_7_6_int_q_reg_v_reg_1__0_ ( .D(i_data_conv_v[4]), .CK(
        pe_1_7_6_net2691), .RN(pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_v[16]) );
  DFFR_X1 pe_1_7_6_int_q_reg_v_reg_1__1_ ( .D(i_data_conv_v[5]), .CK(
        pe_1_7_6_net2691), .RN(pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_v[17]) );
  DFFR_X1 pe_1_7_6_int_q_reg_v_reg_1__2_ ( .D(i_data_conv_v[6]), .CK(
        pe_1_7_6_net2691), .RN(pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_v[18]) );
  DFFR_X1 pe_1_7_6_int_q_reg_v_reg_1__3_ ( .D(i_data_conv_v[7]), .CK(
        pe_1_7_6_net2691), .RN(pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_v[19]) );
  DFFR_X1 pe_1_7_6_int_q_reg_v_reg_2__0_ ( .D(i_data_conv_v[4]), .CK(
        pe_1_7_6_net2696), .RN(pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_v[12]) );
  DFFR_X1 pe_1_7_6_int_q_reg_v_reg_2__1_ ( .D(i_data_conv_v[5]), .CK(
        pe_1_7_6_net2696), .RN(pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_v[13]) );
  DFFR_X1 pe_1_7_6_int_q_reg_v_reg_2__2_ ( .D(i_data_conv_v[6]), .CK(
        pe_1_7_6_net2696), .RN(pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_v[14]) );
  DFFR_X1 pe_1_7_6_int_q_reg_v_reg_2__3_ ( .D(i_data_conv_v[7]), .CK(
        pe_1_7_6_net2696), .RN(pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_v[15]) );
  DFFR_X1 pe_1_7_6_int_q_reg_v_reg_3__0_ ( .D(i_data_conv_v[4]), .CK(
        pe_1_7_6_net2701), .RN(pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_v[8]) );
  DFFR_X1 pe_1_7_6_int_q_reg_v_reg_3__1_ ( .D(i_data_conv_v[5]), .CK(
        pe_1_7_6_net2701), .RN(pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_v[9]) );
  DFFR_X1 pe_1_7_6_int_q_reg_v_reg_3__2_ ( .D(i_data_conv_v[6]), .CK(
        pe_1_7_6_net2701), .RN(pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_v[10]) );
  DFFR_X1 pe_1_7_6_int_q_reg_v_reg_3__3_ ( .D(i_data_conv_v[7]), .CK(
        pe_1_7_6_net2701), .RN(pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_v[11]) );
  DFFR_X1 pe_1_7_6_int_q_reg_v_reg_4__0_ ( .D(i_data_conv_v[4]), .CK(
        pe_1_7_6_net2706), .RN(pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_v[4]) );
  DFFR_X1 pe_1_7_6_int_q_reg_v_reg_4__1_ ( .D(i_data_conv_v[5]), .CK(
        pe_1_7_6_net2706), .RN(pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_v[5]) );
  DFFR_X1 pe_1_7_6_int_q_reg_v_reg_4__2_ ( .D(i_data_conv_v[6]), .CK(
        pe_1_7_6_net2706), .RN(pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_v[6]) );
  DFFR_X1 pe_1_7_6_int_q_reg_v_reg_4__3_ ( .D(i_data_conv_v[7]), .CK(
        pe_1_7_6_net2706), .RN(pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_v[7]) );
  DFFR_X1 pe_1_7_6_int_q_reg_v_reg_5__0_ ( .D(i_data_conv_v[4]), .CK(
        pe_1_7_6_net2711), .RN(pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_v[0]) );
  DFFR_X1 pe_1_7_6_int_q_reg_v_reg_5__1_ ( .D(i_data_conv_v[5]), .CK(
        pe_1_7_6_net2711), .RN(pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_v[1]) );
  DFFR_X1 pe_1_7_6_int_q_reg_v_reg_5__2_ ( .D(i_data_conv_v[6]), .CK(
        pe_1_7_6_net2711), .RN(pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_v[2]) );
  DFFR_X1 pe_1_7_6_int_q_reg_v_reg_5__3_ ( .D(i_data_conv_v[7]), .CK(
        pe_1_7_6_net2711), .RN(pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_7_6_int_q_reg_h_reg_0__0_ ( .D(int_data_x_7__7__0_), .SI(
        i_data_conv_v[4]), .SE(pe_1_7_6_n63), .CK(pe_1_7_6_net2655), .RN(
        pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_7_6_int_q_reg_h_reg_0__1_ ( .D(int_data_x_7__7__1_), .SI(
        i_data_conv_v[5]), .SE(pe_1_7_6_n63), .CK(pe_1_7_6_net2655), .RN(
        pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_7_6_int_q_reg_h_reg_0__2_ ( .D(int_data_x_7__7__2_), .SI(
        i_data_conv_v[6]), .SE(pe_1_7_6_n63), .CK(pe_1_7_6_net2655), .RN(
        pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_7_6_int_q_reg_h_reg_0__3_ ( .D(int_data_x_7__7__3_), .SI(
        i_data_conv_v[7]), .SE(pe_1_7_6_n63), .CK(pe_1_7_6_net2655), .RN(
        pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_7_6_int_q_reg_h_reg_1__0_ ( .D(int_data_x_7__7__0_), .SI(
        i_data_conv_v[4]), .SE(pe_1_7_6_n63), .CK(pe_1_7_6_net2661), .RN(
        pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_7_6_int_q_reg_h_reg_1__1_ ( .D(int_data_x_7__7__1_), .SI(
        i_data_conv_v[5]), .SE(pe_1_7_6_n63), .CK(pe_1_7_6_net2661), .RN(
        pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_7_6_int_q_reg_h_reg_1__2_ ( .D(int_data_x_7__7__2_), .SI(
        i_data_conv_v[6]), .SE(pe_1_7_6_n63), .CK(pe_1_7_6_net2661), .RN(
        pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_7_6_int_q_reg_h_reg_1__3_ ( .D(int_data_x_7__7__3_), .SI(
        i_data_conv_v[7]), .SE(pe_1_7_6_n63), .CK(pe_1_7_6_net2661), .RN(
        pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_7_6_int_q_reg_h_reg_2__0_ ( .D(int_data_x_7__7__0_), .SI(
        i_data_conv_v[4]), .SE(pe_1_7_6_n63), .CK(pe_1_7_6_net2666), .RN(
        pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_7_6_int_q_reg_h_reg_2__1_ ( .D(int_data_x_7__7__1_), .SI(
        i_data_conv_v[5]), .SE(pe_1_7_6_n63), .CK(pe_1_7_6_net2666), .RN(
        pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_7_6_int_q_reg_h_reg_2__2_ ( .D(int_data_x_7__7__2_), .SI(
        i_data_conv_v[6]), .SE(pe_1_7_6_n63), .CK(pe_1_7_6_net2666), .RN(
        pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_7_6_int_q_reg_h_reg_2__3_ ( .D(int_data_x_7__7__3_), .SI(
        i_data_conv_v[7]), .SE(pe_1_7_6_n63), .CK(pe_1_7_6_net2666), .RN(
        pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_7_6_int_q_reg_h_reg_3__0_ ( .D(int_data_x_7__7__0_), .SI(
        i_data_conv_v[4]), .SE(pe_1_7_6_n63), .CK(pe_1_7_6_net2671), .RN(
        pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_7_6_int_q_reg_h_reg_3__1_ ( .D(int_data_x_7__7__1_), .SI(
        i_data_conv_v[5]), .SE(pe_1_7_6_n63), .CK(pe_1_7_6_net2671), .RN(
        pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_7_6_int_q_reg_h_reg_3__2_ ( .D(int_data_x_7__7__2_), .SI(
        i_data_conv_v[6]), .SE(pe_1_7_6_n63), .CK(pe_1_7_6_net2671), .RN(
        pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_7_6_int_q_reg_h_reg_3__3_ ( .D(int_data_x_7__7__3_), .SI(
        i_data_conv_v[7]), .SE(pe_1_7_6_n63), .CK(pe_1_7_6_net2671), .RN(
        pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_7_6_int_q_reg_h_reg_4__0_ ( .D(int_data_x_7__7__0_), .SI(
        i_data_conv_v[4]), .SE(n70), .CK(pe_1_7_6_net2676), .RN(pe_1_7_6_n67), 
        .Q(pe_1_7_6_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_7_6_int_q_reg_h_reg_4__1_ ( .D(int_data_x_7__7__1_), .SI(
        i_data_conv_v[5]), .SE(n70), .CK(pe_1_7_6_net2676), .RN(pe_1_7_6_n67), 
        .Q(pe_1_7_6_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_7_6_int_q_reg_h_reg_4__2_ ( .D(int_data_x_7__7__2_), .SI(
        i_data_conv_v[6]), .SE(n70), .CK(pe_1_7_6_net2676), .RN(pe_1_7_6_n67), 
        .Q(pe_1_7_6_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_7_6_int_q_reg_h_reg_4__3_ ( .D(int_data_x_7__7__3_), .SI(
        i_data_conv_v[7]), .SE(n70), .CK(pe_1_7_6_net2676), .RN(pe_1_7_6_n67), 
        .Q(pe_1_7_6_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_7_6_int_q_reg_h_reg_5__0_ ( .D(int_data_x_7__7__0_), .SI(
        i_data_conv_v[4]), .SE(pe_1_7_6_n63), .CK(pe_1_7_6_net2681), .RN(
        pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_7_6_int_q_reg_h_reg_5__1_ ( .D(int_data_x_7__7__1_), .SI(
        i_data_conv_v[5]), .SE(pe_1_7_6_n63), .CK(pe_1_7_6_net2681), .RN(
        pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_7_6_int_q_reg_h_reg_5__2_ ( .D(int_data_x_7__7__2_), .SI(
        i_data_conv_v[6]), .SE(pe_1_7_6_n63), .CK(pe_1_7_6_net2681), .RN(
        pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_7_6_int_q_reg_h_reg_5__3_ ( .D(int_data_x_7__7__3_), .SI(
        i_data_conv_v[7]), .SE(pe_1_7_6_n63), .CK(pe_1_7_6_net2681), .RN(
        pe_1_7_6_n67), .Q(pe_1_7_6_int_q_reg_h[3]) );
  FA_X1 pe_1_7_6_sub_81_U2_7 ( .A(int_data_res_7__6__7_), .B(pe_1_7_6_n71), 
        .CI(pe_1_7_6_sub_81_carry[7]), .S(pe_1_7_6_N77) );
  FA_X1 pe_1_7_6_sub_81_U2_6 ( .A(int_data_res_7__6__6_), .B(pe_1_7_6_n71), 
        .CI(pe_1_7_6_sub_81_carry[6]), .CO(pe_1_7_6_sub_81_carry[7]), .S(
        pe_1_7_6_N76) );
  FA_X1 pe_1_7_6_sub_81_U2_5 ( .A(int_data_res_7__6__5_), .B(pe_1_7_6_n71), 
        .CI(pe_1_7_6_sub_81_carry[5]), .CO(pe_1_7_6_sub_81_carry[6]), .S(
        pe_1_7_6_N75) );
  FA_X1 pe_1_7_6_sub_81_U2_4 ( .A(int_data_res_7__6__4_), .B(pe_1_7_6_n71), 
        .CI(pe_1_7_6_sub_81_carry[4]), .CO(pe_1_7_6_sub_81_carry[5]), .S(
        pe_1_7_6_N74) );
  FA_X1 pe_1_7_6_sub_81_U2_3 ( .A(int_data_res_7__6__3_), .B(pe_1_7_6_n71), 
        .CI(pe_1_7_6_sub_81_carry[3]), .CO(pe_1_7_6_sub_81_carry[4]), .S(
        pe_1_7_6_N73) );
  FA_X1 pe_1_7_6_sub_81_U2_2 ( .A(int_data_res_7__6__2_), .B(pe_1_7_6_n70), 
        .CI(pe_1_7_6_sub_81_carry[2]), .CO(pe_1_7_6_sub_81_carry[3]), .S(
        pe_1_7_6_N72) );
  FA_X1 pe_1_7_6_sub_81_U2_1 ( .A(int_data_res_7__6__1_), .B(pe_1_7_6_n69), 
        .CI(pe_1_7_6_sub_81_carry[1]), .CO(pe_1_7_6_sub_81_carry[2]), .S(
        pe_1_7_6_N71) );
  FA_X1 pe_1_7_6_add_83_U1_7 ( .A(int_data_res_7__6__7_), .B(
        pe_1_7_6_int_data_3_), .CI(pe_1_7_6_add_83_carry[7]), .S(pe_1_7_6_N85)
         );
  FA_X1 pe_1_7_6_add_83_U1_6 ( .A(int_data_res_7__6__6_), .B(
        pe_1_7_6_int_data_3_), .CI(pe_1_7_6_add_83_carry[6]), .CO(
        pe_1_7_6_add_83_carry[7]), .S(pe_1_7_6_N84) );
  FA_X1 pe_1_7_6_add_83_U1_5 ( .A(int_data_res_7__6__5_), .B(
        pe_1_7_6_int_data_3_), .CI(pe_1_7_6_add_83_carry[5]), .CO(
        pe_1_7_6_add_83_carry[6]), .S(pe_1_7_6_N83) );
  FA_X1 pe_1_7_6_add_83_U1_4 ( .A(int_data_res_7__6__4_), .B(
        pe_1_7_6_int_data_3_), .CI(pe_1_7_6_add_83_carry[4]), .CO(
        pe_1_7_6_add_83_carry[5]), .S(pe_1_7_6_N82) );
  FA_X1 pe_1_7_6_add_83_U1_3 ( .A(int_data_res_7__6__3_), .B(
        pe_1_7_6_int_data_3_), .CI(pe_1_7_6_add_83_carry[3]), .CO(
        pe_1_7_6_add_83_carry[4]), .S(pe_1_7_6_N81) );
  FA_X1 pe_1_7_6_add_83_U1_2 ( .A(int_data_res_7__6__2_), .B(
        pe_1_7_6_int_data_2_), .CI(pe_1_7_6_add_83_carry[2]), .CO(
        pe_1_7_6_add_83_carry[3]), .S(pe_1_7_6_N80) );
  FA_X1 pe_1_7_6_add_83_U1_1 ( .A(int_data_res_7__6__1_), .B(
        pe_1_7_6_int_data_1_), .CI(pe_1_7_6_n2), .CO(pe_1_7_6_add_83_carry[2]), 
        .S(pe_1_7_6_N79) );
  NAND3_X1 pe_1_7_6_U56 ( .A1(n36), .A2(pe_1_7_6_n43), .A3(pe_1_7_6_n60), .ZN(
        pe_1_7_6_n40) );
  NAND3_X1 pe_1_7_6_U55 ( .A1(pe_1_7_6_n43), .A2(pe_1_7_6_n59), .A3(
        pe_1_7_6_n60), .ZN(pe_1_7_6_n39) );
  NAND3_X1 pe_1_7_6_U54 ( .A1(pe_1_7_6_n43), .A2(pe_1_7_6_n61), .A3(n36), .ZN(
        pe_1_7_6_n38) );
  NAND3_X1 pe_1_7_6_U53 ( .A1(pe_1_7_6_n59), .A2(pe_1_7_6_n61), .A3(
        pe_1_7_6_n43), .ZN(pe_1_7_6_n37) );
  DFFR_X1 pe_1_7_6_int_q_acc_reg_6_ ( .D(pe_1_7_6_n73), .CK(pe_1_7_6_net2716), 
        .RN(pe_1_7_6_n66), .Q(int_data_res_7__6__6_) );
  DFFR_X1 pe_1_7_6_int_q_acc_reg_5_ ( .D(pe_1_7_6_n74), .CK(pe_1_7_6_net2716), 
        .RN(pe_1_7_6_n66), .Q(int_data_res_7__6__5_) );
  DFFR_X1 pe_1_7_6_int_q_acc_reg_4_ ( .D(pe_1_7_6_n75), .CK(pe_1_7_6_net2716), 
        .RN(pe_1_7_6_n66), .Q(int_data_res_7__6__4_) );
  DFFR_X1 pe_1_7_6_int_q_acc_reg_3_ ( .D(pe_1_7_6_n76), .CK(pe_1_7_6_net2716), 
        .RN(pe_1_7_6_n66), .Q(int_data_res_7__6__3_) );
  DFFR_X1 pe_1_7_6_int_q_acc_reg_2_ ( .D(pe_1_7_6_n77), .CK(pe_1_7_6_net2716), 
        .RN(pe_1_7_6_n66), .Q(int_data_res_7__6__2_) );
  DFFR_X1 pe_1_7_6_int_q_acc_reg_1_ ( .D(pe_1_7_6_n78), .CK(pe_1_7_6_net2716), 
        .RN(pe_1_7_6_n66), .Q(int_data_res_7__6__1_) );
  DFFR_X1 pe_1_7_6_int_q_acc_reg_7_ ( .D(pe_1_7_6_n72), .CK(pe_1_7_6_net2716), 
        .RN(pe_1_7_6_n66), .Q(int_data_res_7__6__7_) );
  CLKGATETST_X1 pe_1_7_6_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_7_6_n83), .SE(1'b0), .GCK(pe_1_7_6_net2655) );
  CLKGATETST_X1 pe_1_7_6_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_7_6_n82), .SE(1'b0), .GCK(pe_1_7_6_net2661) );
  CLKGATETST_X1 pe_1_7_6_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_7_6_n81), .SE(1'b0), .GCK(pe_1_7_6_net2666) );
  CLKGATETST_X1 pe_1_7_6_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_7_6_n80), .SE(1'b0), .GCK(pe_1_7_6_net2671) );
  CLKGATETST_X1 pe_1_7_6_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_7_6_n85), .SE(1'b0), .GCK(pe_1_7_6_net2676) );
  CLKGATETST_X1 pe_1_7_6_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_7_6_n84), .SE(1'b0), .GCK(pe_1_7_6_net2681) );
  CLKGATETST_X1 pe_1_7_6_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_7_6_N64), .SE(1'b0), .GCK(pe_1_7_6_net2686) );
  CLKGATETST_X1 pe_1_7_6_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_7_6_N63), .SE(1'b0), .GCK(pe_1_7_6_net2691) );
  CLKGATETST_X1 pe_1_7_6_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_7_6_N62), .SE(1'b0), .GCK(pe_1_7_6_net2696) );
  CLKGATETST_X1 pe_1_7_6_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_7_6_N61), .SE(1'b0), .GCK(pe_1_7_6_net2701) );
  CLKGATETST_X1 pe_1_7_6_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_7_6_N60), .SE(1'b0), .GCK(pe_1_7_6_net2706) );
  CLKGATETST_X1 pe_1_7_6_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_7_6_N59), .SE(1'b0), .GCK(pe_1_7_6_net2711) );
  CLKGATETST_X1 pe_1_7_6_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_7_6_N90), .SE(1'b0), .GCK(pe_1_7_6_net2716) );
  CLKBUF_X1 pe_1_7_7_U108 ( .A(pe_1_7_7_n68), .Z(pe_1_7_7_n67) );
  INV_X1 pe_1_7_7_U107 ( .A(n78), .ZN(pe_1_7_7_n66) );
  INV_X1 pe_1_7_7_U106 ( .A(n70), .ZN(pe_1_7_7_n65) );
  INV_X1 pe_1_7_7_U105 ( .A(pe_1_7_7_n65), .ZN(pe_1_7_7_n64) );
  INV_X1 pe_1_7_7_U104 ( .A(pe_1_7_7_n61), .ZN(pe_1_7_7_n60) );
  INV_X1 pe_1_7_7_U103 ( .A(n30), .ZN(pe_1_7_7_n58) );
  INV_X1 pe_1_7_7_U102 ( .A(n22), .ZN(pe_1_7_7_n57) );
  MUX2_X1 pe_1_7_7_U101 ( .A(pe_1_7_7_n54), .B(pe_1_7_7_n51), .S(n55), .Z(
        int_data_x_7__7__3_) );
  MUX2_X1 pe_1_7_7_U100 ( .A(pe_1_7_7_n53), .B(pe_1_7_7_n52), .S(pe_1_7_7_n60), 
        .Z(pe_1_7_7_n54) );
  MUX2_X1 pe_1_7_7_U99 ( .A(pe_1_7_7_int_q_reg_h[23]), .B(
        pe_1_7_7_int_q_reg_h[19]), .S(pe_1_7_7_n56), .Z(pe_1_7_7_n53) );
  MUX2_X1 pe_1_7_7_U98 ( .A(pe_1_7_7_int_q_reg_h[15]), .B(
        pe_1_7_7_int_q_reg_h[11]), .S(pe_1_7_7_n56), .Z(pe_1_7_7_n52) );
  MUX2_X1 pe_1_7_7_U97 ( .A(pe_1_7_7_int_q_reg_h[7]), .B(
        pe_1_7_7_int_q_reg_h[3]), .S(pe_1_7_7_n56), .Z(pe_1_7_7_n51) );
  MUX2_X1 pe_1_7_7_U96 ( .A(pe_1_7_7_n50), .B(pe_1_7_7_n47), .S(n55), .Z(
        int_data_x_7__7__2_) );
  MUX2_X1 pe_1_7_7_U95 ( .A(pe_1_7_7_n49), .B(pe_1_7_7_n48), .S(pe_1_7_7_n60), 
        .Z(pe_1_7_7_n50) );
  MUX2_X1 pe_1_7_7_U94 ( .A(pe_1_7_7_int_q_reg_h[22]), .B(
        pe_1_7_7_int_q_reg_h[18]), .S(pe_1_7_7_n56), .Z(pe_1_7_7_n49) );
  MUX2_X1 pe_1_7_7_U93 ( .A(pe_1_7_7_int_q_reg_h[14]), .B(
        pe_1_7_7_int_q_reg_h[10]), .S(pe_1_7_7_n56), .Z(pe_1_7_7_n48) );
  MUX2_X1 pe_1_7_7_U92 ( .A(pe_1_7_7_int_q_reg_h[6]), .B(
        pe_1_7_7_int_q_reg_h[2]), .S(pe_1_7_7_n56), .Z(pe_1_7_7_n47) );
  MUX2_X1 pe_1_7_7_U91 ( .A(pe_1_7_7_n46), .B(pe_1_7_7_n24), .S(n55), .Z(
        int_data_x_7__7__1_) );
  MUX2_X1 pe_1_7_7_U90 ( .A(pe_1_7_7_n45), .B(pe_1_7_7_n25), .S(pe_1_7_7_n60), 
        .Z(pe_1_7_7_n46) );
  MUX2_X1 pe_1_7_7_U89 ( .A(pe_1_7_7_int_q_reg_h[21]), .B(
        pe_1_7_7_int_q_reg_h[17]), .S(pe_1_7_7_n56), .Z(pe_1_7_7_n45) );
  MUX2_X1 pe_1_7_7_U88 ( .A(pe_1_7_7_int_q_reg_h[13]), .B(
        pe_1_7_7_int_q_reg_h[9]), .S(pe_1_7_7_n56), .Z(pe_1_7_7_n25) );
  MUX2_X1 pe_1_7_7_U87 ( .A(pe_1_7_7_int_q_reg_h[5]), .B(
        pe_1_7_7_int_q_reg_h[1]), .S(pe_1_7_7_n56), .Z(pe_1_7_7_n24) );
  MUX2_X1 pe_1_7_7_U86 ( .A(pe_1_7_7_n23), .B(pe_1_7_7_n20), .S(n55), .Z(
        int_data_x_7__7__0_) );
  MUX2_X1 pe_1_7_7_U85 ( .A(pe_1_7_7_n22), .B(pe_1_7_7_n21), .S(pe_1_7_7_n60), 
        .Z(pe_1_7_7_n23) );
  MUX2_X1 pe_1_7_7_U84 ( .A(pe_1_7_7_int_q_reg_h[20]), .B(
        pe_1_7_7_int_q_reg_h[16]), .S(pe_1_7_7_n56), .Z(pe_1_7_7_n22) );
  MUX2_X1 pe_1_7_7_U83 ( .A(pe_1_7_7_int_q_reg_h[12]), .B(
        pe_1_7_7_int_q_reg_h[8]), .S(pe_1_7_7_n56), .Z(pe_1_7_7_n21) );
  MUX2_X1 pe_1_7_7_U82 ( .A(pe_1_7_7_int_q_reg_h[4]), .B(
        pe_1_7_7_int_q_reg_h[0]), .S(pe_1_7_7_n56), .Z(pe_1_7_7_n20) );
  MUX2_X1 pe_1_7_7_U81 ( .A(pe_1_7_7_n19), .B(pe_1_7_7_n16), .S(n55), .Z(
        int_data_y_7__7__3_) );
  MUX2_X1 pe_1_7_7_U80 ( .A(pe_1_7_7_n18), .B(pe_1_7_7_n17), .S(pe_1_7_7_n60), 
        .Z(pe_1_7_7_n19) );
  MUX2_X1 pe_1_7_7_U79 ( .A(pe_1_7_7_int_q_reg_v[23]), .B(
        pe_1_7_7_int_q_reg_v[19]), .S(pe_1_7_7_n55), .Z(pe_1_7_7_n18) );
  MUX2_X1 pe_1_7_7_U78 ( .A(pe_1_7_7_int_q_reg_v[15]), .B(
        pe_1_7_7_int_q_reg_v[11]), .S(pe_1_7_7_n55), .Z(pe_1_7_7_n17) );
  MUX2_X1 pe_1_7_7_U77 ( .A(pe_1_7_7_int_q_reg_v[7]), .B(
        pe_1_7_7_int_q_reg_v[3]), .S(pe_1_7_7_n55), .Z(pe_1_7_7_n16) );
  MUX2_X1 pe_1_7_7_U76 ( .A(pe_1_7_7_n15), .B(pe_1_7_7_n12), .S(n55), .Z(
        int_data_y_7__7__2_) );
  MUX2_X1 pe_1_7_7_U75 ( .A(pe_1_7_7_n14), .B(pe_1_7_7_n13), .S(pe_1_7_7_n60), 
        .Z(pe_1_7_7_n15) );
  MUX2_X1 pe_1_7_7_U74 ( .A(pe_1_7_7_int_q_reg_v[22]), .B(
        pe_1_7_7_int_q_reg_v[18]), .S(pe_1_7_7_n55), .Z(pe_1_7_7_n14) );
  MUX2_X1 pe_1_7_7_U73 ( .A(pe_1_7_7_int_q_reg_v[14]), .B(
        pe_1_7_7_int_q_reg_v[10]), .S(pe_1_7_7_n55), .Z(pe_1_7_7_n13) );
  MUX2_X1 pe_1_7_7_U72 ( .A(pe_1_7_7_int_q_reg_v[6]), .B(
        pe_1_7_7_int_q_reg_v[2]), .S(pe_1_7_7_n55), .Z(pe_1_7_7_n12) );
  MUX2_X1 pe_1_7_7_U71 ( .A(pe_1_7_7_n11), .B(pe_1_7_7_n8), .S(n55), .Z(
        int_data_y_7__7__1_) );
  MUX2_X1 pe_1_7_7_U70 ( .A(pe_1_7_7_n10), .B(pe_1_7_7_n9), .S(pe_1_7_7_n60), 
        .Z(pe_1_7_7_n11) );
  MUX2_X1 pe_1_7_7_U69 ( .A(pe_1_7_7_int_q_reg_v[21]), .B(
        pe_1_7_7_int_q_reg_v[17]), .S(pe_1_7_7_n55), .Z(pe_1_7_7_n10) );
  MUX2_X1 pe_1_7_7_U68 ( .A(pe_1_7_7_int_q_reg_v[13]), .B(
        pe_1_7_7_int_q_reg_v[9]), .S(pe_1_7_7_n55), .Z(pe_1_7_7_n9) );
  MUX2_X1 pe_1_7_7_U67 ( .A(pe_1_7_7_int_q_reg_v[5]), .B(
        pe_1_7_7_int_q_reg_v[1]), .S(pe_1_7_7_n55), .Z(pe_1_7_7_n8) );
  MUX2_X1 pe_1_7_7_U66 ( .A(pe_1_7_7_n7), .B(pe_1_7_7_n4), .S(n55), .Z(
        int_data_y_7__7__0_) );
  MUX2_X1 pe_1_7_7_U65 ( .A(pe_1_7_7_n6), .B(pe_1_7_7_n5), .S(pe_1_7_7_n60), 
        .Z(pe_1_7_7_n7) );
  MUX2_X1 pe_1_7_7_U64 ( .A(pe_1_7_7_int_q_reg_v[20]), .B(
        pe_1_7_7_int_q_reg_v[16]), .S(pe_1_7_7_n55), .Z(pe_1_7_7_n6) );
  MUX2_X1 pe_1_7_7_U63 ( .A(pe_1_7_7_int_q_reg_v[12]), .B(
        pe_1_7_7_int_q_reg_v[8]), .S(pe_1_7_7_n55), .Z(pe_1_7_7_n5) );
  MUX2_X1 pe_1_7_7_U62 ( .A(pe_1_7_7_int_q_reg_v[4]), .B(
        pe_1_7_7_int_q_reg_v[0]), .S(pe_1_7_7_n55), .Z(pe_1_7_7_n4) );
  AOI222_X1 pe_1_7_7_U61 ( .A1(i_data_acc[1]), .A2(pe_1_7_7_n62), .B1(
        pe_1_7_7_N79), .B2(pe_1_7_7_n27), .C1(pe_1_7_7_N71), .C2(pe_1_7_7_n28), 
        .ZN(pe_1_7_7_n34) );
  INV_X1 pe_1_7_7_U60 ( .A(pe_1_7_7_n34), .ZN(pe_1_7_7_n79) );
  AOI222_X1 pe_1_7_7_U59 ( .A1(i_data_acc[2]), .A2(pe_1_7_7_n62), .B1(
        pe_1_7_7_N80), .B2(pe_1_7_7_n27), .C1(pe_1_7_7_N72), .C2(pe_1_7_7_n28), 
        .ZN(pe_1_7_7_n33) );
  INV_X1 pe_1_7_7_U58 ( .A(pe_1_7_7_n33), .ZN(pe_1_7_7_n78) );
  AOI222_X1 pe_1_7_7_U57 ( .A1(i_data_acc[3]), .A2(pe_1_7_7_n62), .B1(
        pe_1_7_7_N81), .B2(pe_1_7_7_n27), .C1(pe_1_7_7_N73), .C2(pe_1_7_7_n28), 
        .ZN(pe_1_7_7_n32) );
  INV_X1 pe_1_7_7_U52 ( .A(pe_1_7_7_n32), .ZN(pe_1_7_7_n77) );
  AOI222_X1 pe_1_7_7_U51 ( .A1(i_data_acc[4]), .A2(pe_1_7_7_n62), .B1(
        pe_1_7_7_N82), .B2(pe_1_7_7_n27), .C1(pe_1_7_7_N74), .C2(pe_1_7_7_n28), 
        .ZN(pe_1_7_7_n31) );
  INV_X1 pe_1_7_7_U50 ( .A(pe_1_7_7_n31), .ZN(pe_1_7_7_n76) );
  AOI222_X1 pe_1_7_7_U49 ( .A1(i_data_acc[5]), .A2(pe_1_7_7_n62), .B1(
        pe_1_7_7_N83), .B2(pe_1_7_7_n27), .C1(pe_1_7_7_N75), .C2(pe_1_7_7_n28), 
        .ZN(pe_1_7_7_n30) );
  INV_X1 pe_1_7_7_U48 ( .A(pe_1_7_7_n30), .ZN(pe_1_7_7_n75) );
  AOI222_X1 pe_1_7_7_U47 ( .A1(i_data_acc[6]), .A2(pe_1_7_7_n62), .B1(
        pe_1_7_7_N84), .B2(pe_1_7_7_n27), .C1(pe_1_7_7_N76), .C2(pe_1_7_7_n28), 
        .ZN(pe_1_7_7_n29) );
  INV_X1 pe_1_7_7_U46 ( .A(pe_1_7_7_n29), .ZN(pe_1_7_7_n74) );
  XNOR2_X1 pe_1_7_7_U45 ( .A(pe_1_7_7_n69), .B(int_data_res_7__7__0_), .ZN(
        pe_1_7_7_N70) );
  AOI222_X1 pe_1_7_7_U44 ( .A1(i_data_acc[0]), .A2(pe_1_7_7_n62), .B1(
        pe_1_7_7_n1), .B2(pe_1_7_7_n27), .C1(pe_1_7_7_N70), .C2(pe_1_7_7_n28), 
        .ZN(pe_1_7_7_n35) );
  INV_X1 pe_1_7_7_U43 ( .A(pe_1_7_7_n35), .ZN(pe_1_7_7_n80) );
  NAND2_X1 pe_1_7_7_U42 ( .A1(pe_1_7_7_int_data_0_), .A2(pe_1_7_7_n3), .ZN(
        pe_1_7_7_sub_81_carry[1]) );
  INV_X1 pe_1_7_7_U41 ( .A(pe_1_7_7_int_data_1_), .ZN(pe_1_7_7_n70) );
  INV_X1 pe_1_7_7_U40 ( .A(pe_1_7_7_int_data_2_), .ZN(pe_1_7_7_n71) );
  AND2_X1 pe_1_7_7_U39 ( .A1(pe_1_7_7_int_data_0_), .A2(int_data_res_7__7__0_), 
        .ZN(pe_1_7_7_n2) );
  AOI222_X1 pe_1_7_7_U38 ( .A1(pe_1_7_7_n62), .A2(i_data_acc[7]), .B1(
        pe_1_7_7_N85), .B2(pe_1_7_7_n27), .C1(pe_1_7_7_N77), .C2(pe_1_7_7_n28), 
        .ZN(pe_1_7_7_n26) );
  INV_X1 pe_1_7_7_U37 ( .A(pe_1_7_7_n26), .ZN(pe_1_7_7_n73) );
  NOR3_X1 pe_1_7_7_U36 ( .A1(pe_1_7_7_n58), .A2(pe_1_7_7_n63), .A3(int_ckg[0]), 
        .ZN(pe_1_7_7_n36) );
  OR2_X1 pe_1_7_7_U35 ( .A1(pe_1_7_7_n36), .A2(pe_1_7_7_n62), .ZN(pe_1_7_7_N90) );
  AND2_X1 pe_1_7_7_U34 ( .A1(int_data_x_7__7__2_), .A2(n30), .ZN(
        pe_1_7_7_int_data_2_) );
  AND2_X1 pe_1_7_7_U33 ( .A1(int_data_x_7__7__1_), .A2(n30), .ZN(
        pe_1_7_7_int_data_1_) );
  INV_X1 pe_1_7_7_U32 ( .A(n42), .ZN(pe_1_7_7_n61) );
  BUF_X1 pe_1_7_7_U31 ( .A(n64), .Z(pe_1_7_7_n62) );
  AND2_X1 pe_1_7_7_U30 ( .A1(int_data_x_7__7__3_), .A2(n30), .ZN(
        pe_1_7_7_int_data_3_) );
  AND2_X1 pe_1_7_7_U29 ( .A1(int_data_x_7__7__0_), .A2(n30), .ZN(
        pe_1_7_7_int_data_0_) );
  INV_X1 pe_1_7_7_U28 ( .A(n36), .ZN(pe_1_7_7_n59) );
  NAND2_X1 pe_1_7_7_U27 ( .A1(pe_1_7_7_n44), .A2(pe_1_7_7_n59), .ZN(
        pe_1_7_7_n41) );
  AND3_X1 pe_1_7_7_U26 ( .A1(n78), .A2(pe_1_7_7_n61), .A3(n55), .ZN(
        pe_1_7_7_n44) );
  INV_X1 pe_1_7_7_U25 ( .A(pe_1_7_7_int_data_3_), .ZN(pe_1_7_7_n72) );
  NOR2_X1 pe_1_7_7_U24 ( .A1(pe_1_7_7_n66), .A2(n55), .ZN(pe_1_7_7_n43) );
  NOR2_X1 pe_1_7_7_U23 ( .A1(pe_1_7_7_n57), .A2(pe_1_7_7_n62), .ZN(
        pe_1_7_7_n28) );
  NOR2_X1 pe_1_7_7_U22 ( .A1(n22), .A2(pe_1_7_7_n62), .ZN(pe_1_7_7_n27) );
  INV_X1 pe_1_7_7_U21 ( .A(pe_1_7_7_int_data_0_), .ZN(pe_1_7_7_n69) );
  INV_X1 pe_1_7_7_U20 ( .A(pe_1_7_7_n41), .ZN(pe_1_7_7_n86) );
  INV_X1 pe_1_7_7_U19 ( .A(pe_1_7_7_n37), .ZN(pe_1_7_7_n84) );
  INV_X1 pe_1_7_7_U18 ( .A(pe_1_7_7_n38), .ZN(pe_1_7_7_n83) );
  INV_X1 pe_1_7_7_U17 ( .A(pe_1_7_7_n39), .ZN(pe_1_7_7_n82) );
  NOR2_X1 pe_1_7_7_U16 ( .A1(pe_1_7_7_n65), .A2(pe_1_7_7_n42), .ZN(
        pe_1_7_7_N59) );
  NOR2_X1 pe_1_7_7_U15 ( .A1(pe_1_7_7_n65), .A2(pe_1_7_7_n41), .ZN(
        pe_1_7_7_N60) );
  NOR2_X1 pe_1_7_7_U14 ( .A1(pe_1_7_7_n65), .A2(pe_1_7_7_n38), .ZN(
        pe_1_7_7_N63) );
  NOR2_X1 pe_1_7_7_U13 ( .A1(pe_1_7_7_n65), .A2(pe_1_7_7_n40), .ZN(
        pe_1_7_7_N61) );
  NOR2_X1 pe_1_7_7_U12 ( .A1(pe_1_7_7_n65), .A2(pe_1_7_7_n39), .ZN(
        pe_1_7_7_N62) );
  NOR2_X1 pe_1_7_7_U11 ( .A1(pe_1_7_7_n37), .A2(pe_1_7_7_n65), .ZN(
        pe_1_7_7_N64) );
  NAND2_X1 pe_1_7_7_U10 ( .A1(pe_1_7_7_n44), .A2(n36), .ZN(pe_1_7_7_n42) );
  BUF_X1 pe_1_7_7_U9 ( .A(n36), .Z(pe_1_7_7_n55) );
  INV_X1 pe_1_7_7_U8 ( .A(pe_1_7_7_n65), .ZN(pe_1_7_7_n63) );
  BUF_X1 pe_1_7_7_U7 ( .A(n36), .Z(pe_1_7_7_n56) );
  INV_X1 pe_1_7_7_U6 ( .A(pe_1_7_7_n42), .ZN(pe_1_7_7_n85) );
  INV_X1 pe_1_7_7_U5 ( .A(pe_1_7_7_n40), .ZN(pe_1_7_7_n81) );
  INV_X2 pe_1_7_7_U4 ( .A(n86), .ZN(pe_1_7_7_n68) );
  XOR2_X1 pe_1_7_7_U3 ( .A(pe_1_7_7_int_data_0_), .B(int_data_res_7__7__0_), 
        .Z(pe_1_7_7_n1) );
  DFFR_X1 pe_1_7_7_int_q_acc_reg_0_ ( .D(pe_1_7_7_n80), .CK(pe_1_7_7_net2638), 
        .RN(pe_1_7_7_n68), .Q(int_data_res_7__7__0_), .QN(pe_1_7_7_n3) );
  DFFR_X1 pe_1_7_7_int_q_reg_v_reg_0__0_ ( .D(i_data_conv_v[0]), .CK(
        pe_1_7_7_net2608), .RN(pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_v[20]) );
  DFFR_X1 pe_1_7_7_int_q_reg_v_reg_0__1_ ( .D(i_data_conv_v[1]), .CK(
        pe_1_7_7_net2608), .RN(pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_v[21]) );
  DFFR_X1 pe_1_7_7_int_q_reg_v_reg_0__2_ ( .D(i_data_conv_v[2]), .CK(
        pe_1_7_7_net2608), .RN(pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_v[22]) );
  DFFR_X1 pe_1_7_7_int_q_reg_v_reg_0__3_ ( .D(i_data_conv_v[3]), .CK(
        pe_1_7_7_net2608), .RN(pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_v[23]) );
  DFFR_X1 pe_1_7_7_int_q_reg_v_reg_1__0_ ( .D(i_data_conv_v[0]), .CK(
        pe_1_7_7_net2613), .RN(pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_v[16]) );
  DFFR_X1 pe_1_7_7_int_q_reg_v_reg_1__1_ ( .D(i_data_conv_v[1]), .CK(
        pe_1_7_7_net2613), .RN(pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_v[17]) );
  DFFR_X1 pe_1_7_7_int_q_reg_v_reg_1__2_ ( .D(i_data_conv_v[2]), .CK(
        pe_1_7_7_net2613), .RN(pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_v[18]) );
  DFFR_X1 pe_1_7_7_int_q_reg_v_reg_1__3_ ( .D(i_data_conv_v[3]), .CK(
        pe_1_7_7_net2613), .RN(pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_v[19]) );
  DFFR_X1 pe_1_7_7_int_q_reg_v_reg_2__0_ ( .D(i_data_conv_v[0]), .CK(
        pe_1_7_7_net2618), .RN(pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_v[12]) );
  DFFR_X1 pe_1_7_7_int_q_reg_v_reg_2__1_ ( .D(i_data_conv_v[1]), .CK(
        pe_1_7_7_net2618), .RN(pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_v[13]) );
  DFFR_X1 pe_1_7_7_int_q_reg_v_reg_2__2_ ( .D(i_data_conv_v[2]), .CK(
        pe_1_7_7_net2618), .RN(pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_v[14]) );
  DFFR_X1 pe_1_7_7_int_q_reg_v_reg_2__3_ ( .D(i_data_conv_v[3]), .CK(
        pe_1_7_7_net2618), .RN(pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_v[15]) );
  DFFR_X1 pe_1_7_7_int_q_reg_v_reg_3__0_ ( .D(i_data_conv_v[0]), .CK(
        pe_1_7_7_net2623), .RN(pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_v[8]) );
  DFFR_X1 pe_1_7_7_int_q_reg_v_reg_3__1_ ( .D(i_data_conv_v[1]), .CK(
        pe_1_7_7_net2623), .RN(pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_v[9]) );
  DFFR_X1 pe_1_7_7_int_q_reg_v_reg_3__2_ ( .D(i_data_conv_v[2]), .CK(
        pe_1_7_7_net2623), .RN(pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_v[10]) );
  DFFR_X1 pe_1_7_7_int_q_reg_v_reg_3__3_ ( .D(i_data_conv_v[3]), .CK(
        pe_1_7_7_net2623), .RN(pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_v[11]) );
  DFFR_X1 pe_1_7_7_int_q_reg_v_reg_4__0_ ( .D(i_data_conv_v[0]), .CK(
        pe_1_7_7_net2628), .RN(pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_v[4]) );
  DFFR_X1 pe_1_7_7_int_q_reg_v_reg_4__1_ ( .D(i_data_conv_v[1]), .CK(
        pe_1_7_7_net2628), .RN(pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_v[5]) );
  DFFR_X1 pe_1_7_7_int_q_reg_v_reg_4__2_ ( .D(i_data_conv_v[2]), .CK(
        pe_1_7_7_net2628), .RN(pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_v[6]) );
  DFFR_X1 pe_1_7_7_int_q_reg_v_reg_4__3_ ( .D(i_data_conv_v[3]), .CK(
        pe_1_7_7_net2628), .RN(pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_v[7]) );
  DFFR_X1 pe_1_7_7_int_q_reg_v_reg_5__0_ ( .D(i_data_conv_v[0]), .CK(
        pe_1_7_7_net2633), .RN(pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_v[0]) );
  DFFR_X1 pe_1_7_7_int_q_reg_v_reg_5__1_ ( .D(i_data_conv_v[1]), .CK(
        pe_1_7_7_net2633), .RN(pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_v[1]) );
  DFFR_X1 pe_1_7_7_int_q_reg_v_reg_5__2_ ( .D(i_data_conv_v[2]), .CK(
        pe_1_7_7_net2633), .RN(pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_v[2]) );
  DFFR_X1 pe_1_7_7_int_q_reg_v_reg_5__3_ ( .D(i_data_conv_v[3]), .CK(
        pe_1_7_7_net2633), .RN(pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_v[3]) );
  SDFFR_X1 pe_1_7_7_int_q_reg_h_reg_0__0_ ( .D(i_data_conv_h[0]), .SI(
        i_data_conv_v[0]), .SE(pe_1_7_7_n63), .CK(pe_1_7_7_net2577), .RN(
        pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_h[20]) );
  SDFFR_X1 pe_1_7_7_int_q_reg_h_reg_0__1_ ( .D(i_data_conv_h[1]), .SI(
        i_data_conv_v[1]), .SE(pe_1_7_7_n63), .CK(pe_1_7_7_net2577), .RN(
        pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_h[21]) );
  SDFFR_X1 pe_1_7_7_int_q_reg_h_reg_0__2_ ( .D(i_data_conv_h[2]), .SI(
        i_data_conv_v[2]), .SE(pe_1_7_7_n63), .CK(pe_1_7_7_net2577), .RN(
        pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_h[22]) );
  SDFFR_X1 pe_1_7_7_int_q_reg_h_reg_0__3_ ( .D(i_data_conv_h[3]), .SI(
        i_data_conv_v[3]), .SE(pe_1_7_7_n63), .CK(pe_1_7_7_net2577), .RN(
        pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_h[23]) );
  SDFFR_X1 pe_1_7_7_int_q_reg_h_reg_1__0_ ( .D(i_data_conv_h[0]), .SI(
        i_data_conv_v[0]), .SE(pe_1_7_7_n63), .CK(pe_1_7_7_net2583), .RN(
        pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_h[16]) );
  SDFFR_X1 pe_1_7_7_int_q_reg_h_reg_1__1_ ( .D(i_data_conv_h[1]), .SI(
        i_data_conv_v[1]), .SE(pe_1_7_7_n63), .CK(pe_1_7_7_net2583), .RN(
        pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_h[17]) );
  SDFFR_X1 pe_1_7_7_int_q_reg_h_reg_1__2_ ( .D(i_data_conv_h[2]), .SI(
        i_data_conv_v[2]), .SE(pe_1_7_7_n63), .CK(pe_1_7_7_net2583), .RN(
        pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_h[18]) );
  SDFFR_X1 pe_1_7_7_int_q_reg_h_reg_1__3_ ( .D(i_data_conv_h[3]), .SI(
        i_data_conv_v[3]), .SE(pe_1_7_7_n63), .CK(pe_1_7_7_net2583), .RN(
        pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_h[19]) );
  SDFFR_X1 pe_1_7_7_int_q_reg_h_reg_2__0_ ( .D(i_data_conv_h[0]), .SI(
        i_data_conv_v[0]), .SE(pe_1_7_7_n63), .CK(pe_1_7_7_net2588), .RN(
        pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_h[12]) );
  SDFFR_X1 pe_1_7_7_int_q_reg_h_reg_2__1_ ( .D(i_data_conv_h[1]), .SI(
        i_data_conv_v[1]), .SE(pe_1_7_7_n63), .CK(pe_1_7_7_net2588), .RN(
        pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_h[13]) );
  SDFFR_X1 pe_1_7_7_int_q_reg_h_reg_2__2_ ( .D(i_data_conv_h[2]), .SI(
        i_data_conv_v[2]), .SE(pe_1_7_7_n63), .CK(pe_1_7_7_net2588), .RN(
        pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_h[14]) );
  SDFFR_X1 pe_1_7_7_int_q_reg_h_reg_2__3_ ( .D(i_data_conv_h[3]), .SI(
        i_data_conv_v[3]), .SE(pe_1_7_7_n63), .CK(pe_1_7_7_net2588), .RN(
        pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_h[15]) );
  SDFFR_X1 pe_1_7_7_int_q_reg_h_reg_3__0_ ( .D(i_data_conv_h[0]), .SI(
        i_data_conv_v[0]), .SE(pe_1_7_7_n63), .CK(pe_1_7_7_net2593), .RN(
        pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_h[8]) );
  SDFFR_X1 pe_1_7_7_int_q_reg_h_reg_3__1_ ( .D(i_data_conv_h[1]), .SI(
        i_data_conv_v[1]), .SE(pe_1_7_7_n63), .CK(pe_1_7_7_net2593), .RN(
        pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_h[9]) );
  SDFFR_X1 pe_1_7_7_int_q_reg_h_reg_3__2_ ( .D(i_data_conv_h[2]), .SI(
        i_data_conv_v[2]), .SE(pe_1_7_7_n63), .CK(pe_1_7_7_net2593), .RN(
        pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_h[10]) );
  SDFFR_X1 pe_1_7_7_int_q_reg_h_reg_3__3_ ( .D(i_data_conv_h[3]), .SI(
        i_data_conv_v[3]), .SE(pe_1_7_7_n63), .CK(pe_1_7_7_net2593), .RN(
        pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_h[11]) );
  SDFFR_X1 pe_1_7_7_int_q_reg_h_reg_4__0_ ( .D(i_data_conv_h[0]), .SI(
        i_data_conv_v[0]), .SE(pe_1_7_7_n64), .CK(pe_1_7_7_net2598), .RN(
        pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_h[4]) );
  SDFFR_X1 pe_1_7_7_int_q_reg_h_reg_4__1_ ( .D(i_data_conv_h[1]), .SI(
        i_data_conv_v[1]), .SE(pe_1_7_7_n64), .CK(pe_1_7_7_net2598), .RN(
        pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_h[5]) );
  SDFFR_X1 pe_1_7_7_int_q_reg_h_reg_4__2_ ( .D(i_data_conv_h[2]), .SI(
        i_data_conv_v[2]), .SE(pe_1_7_7_n64), .CK(pe_1_7_7_net2598), .RN(
        pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_h[6]) );
  SDFFR_X1 pe_1_7_7_int_q_reg_h_reg_4__3_ ( .D(i_data_conv_h[3]), .SI(
        i_data_conv_v[3]), .SE(pe_1_7_7_n64), .CK(pe_1_7_7_net2598), .RN(
        pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_h[7]) );
  SDFFR_X1 pe_1_7_7_int_q_reg_h_reg_5__0_ ( .D(i_data_conv_h[0]), .SI(
        i_data_conv_v[0]), .SE(pe_1_7_7_n64), .CK(pe_1_7_7_net2603), .RN(
        pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_h[0]) );
  SDFFR_X1 pe_1_7_7_int_q_reg_h_reg_5__1_ ( .D(i_data_conv_h[1]), .SI(
        i_data_conv_v[1]), .SE(pe_1_7_7_n64), .CK(pe_1_7_7_net2603), .RN(
        pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_h[1]) );
  SDFFR_X1 pe_1_7_7_int_q_reg_h_reg_5__2_ ( .D(i_data_conv_h[2]), .SI(
        i_data_conv_v[2]), .SE(pe_1_7_7_n64), .CK(pe_1_7_7_net2603), .RN(
        pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_h[2]) );
  SDFFR_X1 pe_1_7_7_int_q_reg_h_reg_5__3_ ( .D(i_data_conv_h[3]), .SI(
        i_data_conv_v[3]), .SE(pe_1_7_7_n64), .CK(pe_1_7_7_net2603), .RN(
        pe_1_7_7_n68), .Q(pe_1_7_7_int_q_reg_h[3]) );
  FA_X1 pe_1_7_7_sub_81_U2_7 ( .A(int_data_res_7__7__7_), .B(pe_1_7_7_n72), 
        .CI(pe_1_7_7_sub_81_carry[7]), .S(pe_1_7_7_N77) );
  FA_X1 pe_1_7_7_sub_81_U2_6 ( .A(int_data_res_7__7__6_), .B(pe_1_7_7_n72), 
        .CI(pe_1_7_7_sub_81_carry[6]), .CO(pe_1_7_7_sub_81_carry[7]), .S(
        pe_1_7_7_N76) );
  FA_X1 pe_1_7_7_sub_81_U2_5 ( .A(int_data_res_7__7__5_), .B(pe_1_7_7_n72), 
        .CI(pe_1_7_7_sub_81_carry[5]), .CO(pe_1_7_7_sub_81_carry[6]), .S(
        pe_1_7_7_N75) );
  FA_X1 pe_1_7_7_sub_81_U2_4 ( .A(int_data_res_7__7__4_), .B(pe_1_7_7_n72), 
        .CI(pe_1_7_7_sub_81_carry[4]), .CO(pe_1_7_7_sub_81_carry[5]), .S(
        pe_1_7_7_N74) );
  FA_X1 pe_1_7_7_sub_81_U2_3 ( .A(int_data_res_7__7__3_), .B(pe_1_7_7_n72), 
        .CI(pe_1_7_7_sub_81_carry[3]), .CO(pe_1_7_7_sub_81_carry[4]), .S(
        pe_1_7_7_N73) );
  FA_X1 pe_1_7_7_sub_81_U2_2 ( .A(int_data_res_7__7__2_), .B(pe_1_7_7_n71), 
        .CI(pe_1_7_7_sub_81_carry[2]), .CO(pe_1_7_7_sub_81_carry[3]), .S(
        pe_1_7_7_N72) );
  FA_X1 pe_1_7_7_sub_81_U2_1 ( .A(int_data_res_7__7__1_), .B(pe_1_7_7_n70), 
        .CI(pe_1_7_7_sub_81_carry[1]), .CO(pe_1_7_7_sub_81_carry[2]), .S(
        pe_1_7_7_N71) );
  FA_X1 pe_1_7_7_add_83_U1_7 ( .A(int_data_res_7__7__7_), .B(
        pe_1_7_7_int_data_3_), .CI(pe_1_7_7_add_83_carry[7]), .S(pe_1_7_7_N85)
         );
  FA_X1 pe_1_7_7_add_83_U1_6 ( .A(int_data_res_7__7__6_), .B(
        pe_1_7_7_int_data_3_), .CI(pe_1_7_7_add_83_carry[6]), .CO(
        pe_1_7_7_add_83_carry[7]), .S(pe_1_7_7_N84) );
  FA_X1 pe_1_7_7_add_83_U1_5 ( .A(int_data_res_7__7__5_), .B(
        pe_1_7_7_int_data_3_), .CI(pe_1_7_7_add_83_carry[5]), .CO(
        pe_1_7_7_add_83_carry[6]), .S(pe_1_7_7_N83) );
  FA_X1 pe_1_7_7_add_83_U1_4 ( .A(int_data_res_7__7__4_), .B(
        pe_1_7_7_int_data_3_), .CI(pe_1_7_7_add_83_carry[4]), .CO(
        pe_1_7_7_add_83_carry[5]), .S(pe_1_7_7_N82) );
  FA_X1 pe_1_7_7_add_83_U1_3 ( .A(int_data_res_7__7__3_), .B(
        pe_1_7_7_int_data_3_), .CI(pe_1_7_7_add_83_carry[3]), .CO(
        pe_1_7_7_add_83_carry[4]), .S(pe_1_7_7_N81) );
  FA_X1 pe_1_7_7_add_83_U1_2 ( .A(int_data_res_7__7__2_), .B(
        pe_1_7_7_int_data_2_), .CI(pe_1_7_7_add_83_carry[2]), .CO(
        pe_1_7_7_add_83_carry[3]), .S(pe_1_7_7_N80) );
  FA_X1 pe_1_7_7_add_83_U1_1 ( .A(int_data_res_7__7__1_), .B(
        pe_1_7_7_int_data_1_), .CI(pe_1_7_7_n2), .CO(pe_1_7_7_add_83_carry[2]), 
        .S(pe_1_7_7_N79) );
  NAND3_X1 pe_1_7_7_U56 ( .A1(n36), .A2(pe_1_7_7_n43), .A3(pe_1_7_7_n60), .ZN(
        pe_1_7_7_n40) );
  NAND3_X1 pe_1_7_7_U55 ( .A1(pe_1_7_7_n43), .A2(pe_1_7_7_n59), .A3(
        pe_1_7_7_n60), .ZN(pe_1_7_7_n39) );
  NAND3_X1 pe_1_7_7_U54 ( .A1(pe_1_7_7_n43), .A2(pe_1_7_7_n61), .A3(n36), .ZN(
        pe_1_7_7_n38) );
  NAND3_X1 pe_1_7_7_U53 ( .A1(pe_1_7_7_n59), .A2(pe_1_7_7_n61), .A3(
        pe_1_7_7_n43), .ZN(pe_1_7_7_n37) );
  DFFR_X1 pe_1_7_7_int_q_acc_reg_6_ ( .D(pe_1_7_7_n74), .CK(pe_1_7_7_net2638), 
        .RN(pe_1_7_7_n67), .Q(int_data_res_7__7__6_) );
  DFFR_X1 pe_1_7_7_int_q_acc_reg_5_ ( .D(pe_1_7_7_n75), .CK(pe_1_7_7_net2638), 
        .RN(pe_1_7_7_n67), .Q(int_data_res_7__7__5_) );
  DFFR_X1 pe_1_7_7_int_q_acc_reg_4_ ( .D(pe_1_7_7_n76), .CK(pe_1_7_7_net2638), 
        .RN(pe_1_7_7_n67), .Q(int_data_res_7__7__4_) );
  DFFR_X1 pe_1_7_7_int_q_acc_reg_3_ ( .D(pe_1_7_7_n77), .CK(pe_1_7_7_net2638), 
        .RN(pe_1_7_7_n67), .Q(int_data_res_7__7__3_) );
  DFFR_X1 pe_1_7_7_int_q_acc_reg_2_ ( .D(pe_1_7_7_n78), .CK(pe_1_7_7_net2638), 
        .RN(pe_1_7_7_n67), .Q(int_data_res_7__7__2_) );
  DFFR_X1 pe_1_7_7_int_q_acc_reg_1_ ( .D(pe_1_7_7_n79), .CK(pe_1_7_7_net2638), 
        .RN(pe_1_7_7_n67), .Q(int_data_res_7__7__1_) );
  DFFR_X1 pe_1_7_7_int_q_acc_reg_7_ ( .D(pe_1_7_7_n73), .CK(pe_1_7_7_net2638), 
        .RN(pe_1_7_7_n67), .Q(int_data_res_7__7__7_) );
  CLKGATETST_X1 pe_1_7_7_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), .E(
        pe_1_7_7_n84), .SE(1'b0), .GCK(pe_1_7_7_net2577) );
  CLKGATETST_X1 pe_1_7_7_clk_gate_int_q_reg_h_reg_1__latch ( .CK(ck), .E(
        pe_1_7_7_n83), .SE(1'b0), .GCK(pe_1_7_7_net2583) );
  CLKGATETST_X1 pe_1_7_7_clk_gate_int_q_reg_h_reg_2__latch ( .CK(ck), .E(
        pe_1_7_7_n82), .SE(1'b0), .GCK(pe_1_7_7_net2588) );
  CLKGATETST_X1 pe_1_7_7_clk_gate_int_q_reg_h_reg_3__latch ( .CK(ck), .E(
        pe_1_7_7_n81), .SE(1'b0), .GCK(pe_1_7_7_net2593) );
  CLKGATETST_X1 pe_1_7_7_clk_gate_int_q_reg_h_reg_4__latch ( .CK(ck), .E(
        pe_1_7_7_n86), .SE(1'b0), .GCK(pe_1_7_7_net2598) );
  CLKGATETST_X1 pe_1_7_7_clk_gate_int_q_reg_h_reg_5__latch ( .CK(ck), .E(
        pe_1_7_7_n85), .SE(1'b0), .GCK(pe_1_7_7_net2603) );
  CLKGATETST_X1 pe_1_7_7_clk_gate_int_q_reg_v_reg_0__latch ( .CK(ck), .E(
        pe_1_7_7_N64), .SE(1'b0), .GCK(pe_1_7_7_net2608) );
  CLKGATETST_X1 pe_1_7_7_clk_gate_int_q_reg_v_reg_1__latch ( .CK(ck), .E(
        pe_1_7_7_N63), .SE(1'b0), .GCK(pe_1_7_7_net2613) );
  CLKGATETST_X1 pe_1_7_7_clk_gate_int_q_reg_v_reg_2__latch ( .CK(ck), .E(
        pe_1_7_7_N62), .SE(1'b0), .GCK(pe_1_7_7_net2618) );
  CLKGATETST_X1 pe_1_7_7_clk_gate_int_q_reg_v_reg_3__latch ( .CK(ck), .E(
        pe_1_7_7_N61), .SE(1'b0), .GCK(pe_1_7_7_net2623) );
  CLKGATETST_X1 pe_1_7_7_clk_gate_int_q_reg_v_reg_4__latch ( .CK(ck), .E(
        pe_1_7_7_N60), .SE(1'b0), .GCK(pe_1_7_7_net2628) );
  CLKGATETST_X1 pe_1_7_7_clk_gate_int_q_reg_v_reg_5__latch ( .CK(ck), .E(
        pe_1_7_7_N59), .SE(1'b0), .GCK(pe_1_7_7_net2633) );
  CLKGATETST_X1 pe_1_7_7_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        pe_1_7_7_N90), .SE(1'b0), .GCK(pe_1_7_7_net2638) );
endmodule

