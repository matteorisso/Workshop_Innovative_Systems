library verilog;
use verilog.vl_types.all;
entity cfg_sv_unit is
end cfg_sv_unit;
