
module dp ( ck, rst, i_acth, i_actv, i_weight, i_gamma, i_beta, arv_npu, 
        arv_ckg, arv_k, arv_tile, arv_ifmaps, arv_ofmaps, ctrl_en_npu, 
        ctrl_ldh_v_n, ctrl_en_hmode, ctrl_en_vmode, ctrl_wr_pipe, s_tc_hmode, 
        s_tc_vmode, s_tc_res, s_tc_npu_ptr, s_tc_tilev, s_tc_tileh, 
        s_tc_ifmaps, s_tc_ofmaps, i_weight_addr, i_data_ev_odd_n, 
        i_data_even_addr, i_data_odd_addr, o_data_ev_odd_n, o_data_even_addr, 
        o_data_odd_addr, o_data );
  input [15:0] i_acth;
  input [15:0] i_actv;
  input [1:0] i_weight;
  input [7:0] i_gamma;
  input [7:0] i_beta;
  input [2:0] arv_npu;
  input [2:0] arv_ckg;
  input [2:0] arv_k;
  input [1:0] arv_tile;
  input [2:0] arv_ifmaps;
  input [3:0] arv_ofmaps;
  output [31:0] i_weight_addr;
  output [9:0] i_data_even_addr;
  output [9:0] i_data_odd_addr;
  output [9:0] o_data_even_addr;
  output [9:0] o_data_odd_addr;
  output [63:0] o_data;
  input ck, rst, ctrl_en_npu, ctrl_ldh_v_n, ctrl_en_hmode, ctrl_en_vmode,
         ctrl_wr_pipe;
  output s_tc_hmode, s_tc_vmode, s_tc_res, s_tc_npu_ptr, s_tc_tilev,
         s_tc_tileh, s_tc_ifmaps, s_tc_ofmaps, i_data_ev_odd_n,
         o_data_ev_odd_n;
  wire   ps_ctrl_en_npu, ps_ctrl_ldh_v_n, ps_ctrl_wr_pipe, ps_int_s_tc_tilev,
         ps_int_s_tc_tileh, int_en_hmode, int_en_vmode, int_en_npu_ptr,
         int_en_tilev_ptr, int_inc_i_data_even, int_inc_i_data_odd,
         int_rst_i_data_addr, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28,
         int_inc_i_w_addr, net2652, net2658, net2663, net2668, n5, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, act_buffer_inst_n196,
         act_buffer_inst_n195, act_buffer_inst_n194, act_buffer_inst_n193,
         act_buffer_inst_n192, act_buffer_inst_n191, act_buffer_inst_n190,
         act_buffer_inst_n189, act_buffer_inst_n188, act_buffer_inst_n187,
         act_buffer_inst_n186, act_buffer_inst_n185, act_buffer_inst_n184,
         act_buffer_inst_n183, act_buffer_inst_n182, act_buffer_inst_n181,
         act_buffer_inst_n180, act_buffer_inst_n179, act_buffer_inst_n178,
         act_buffer_inst_n177, act_buffer_inst_n176, act_buffer_inst_n175,
         act_buffer_inst_n174, act_buffer_inst_n173, act_buffer_inst_n172,
         act_buffer_inst_n171, act_buffer_inst_n170, act_buffer_inst_n169,
         act_buffer_inst_n168, act_buffer_inst_n167, act_buffer_inst_n166,
         act_buffer_inst_n165, act_buffer_inst_n164, act_buffer_inst_n163,
         act_buffer_inst_n162, act_buffer_inst_n161, act_buffer_inst_n160,
         act_buffer_inst_n159, act_buffer_inst_n9, act_buffer_inst_n8,
         act_buffer_inst_n7, act_buffer_inst_n6, act_buffer_inst_n5,
         act_buffer_inst_n4, act_buffer_inst_n3, act_buffer_inst_n2,
         act_buffer_inst_n1, act_buffer_inst_n158, act_buffer_inst_n157,
         act_buffer_inst_n156, act_buffer_inst_n155, act_buffer_inst_n154,
         act_buffer_inst_n153, act_buffer_inst_n152, act_buffer_inst_n151,
         act_buffer_inst_n150, act_buffer_inst_n149, act_buffer_inst_n148,
         act_buffer_inst_n147, act_buffer_inst_n146, act_buffer_inst_n145,
         act_buffer_inst_n144, act_buffer_inst_n143, act_buffer_inst_n142,
         act_buffer_inst_n141, act_buffer_inst_n140, act_buffer_inst_n139,
         act_buffer_inst_n138, act_buffer_inst_n137, act_buffer_inst_n136,
         act_buffer_inst_n135, act_buffer_inst_n134, act_buffer_inst_n133,
         act_buffer_inst_n132, act_buffer_inst_n131, act_buffer_inst_n130,
         act_buffer_inst_n129, act_buffer_inst_n128, act_buffer_inst_n127,
         act_buffer_inst_n126, act_buffer_inst_n125, act_buffer_inst_n124,
         act_buffer_inst_n123, act_buffer_inst_n122, act_buffer_inst_n121,
         act_buffer_inst_n120, act_buffer_inst_n119, act_buffer_inst_n118,
         act_buffer_inst_n117, act_buffer_inst_n116, act_buffer_inst_n115,
         act_buffer_inst_n114, act_buffer_inst_n113, act_buffer_inst_n112,
         act_buffer_inst_n111, act_buffer_inst_n110, act_buffer_inst_n109,
         act_buffer_inst_n108, act_buffer_inst_n107, act_buffer_inst_n106,
         act_buffer_inst_n105, act_buffer_inst_n104, act_buffer_inst_n103,
         act_buffer_inst_n102, act_buffer_inst_n101, act_buffer_inst_n100,
         act_buffer_inst_n99, act_buffer_inst_n98, act_buffer_inst_n97,
         act_buffer_inst_n96, act_buffer_inst_n95, act_buffer_inst_n94,
         act_buffer_inst_n93, act_buffer_inst_n92, act_buffer_inst_n91,
         act_buffer_inst_n90, act_buffer_inst_n89, act_buffer_inst_n88,
         act_buffer_inst_n87, act_buffer_inst_n86, act_buffer_inst_n85,
         act_buffer_inst_n84, act_buffer_inst_n83, act_buffer_inst_n82,
         act_buffer_inst_n81, act_buffer_inst_n80, act_buffer_inst_n79,
         act_buffer_inst_n78, act_buffer_inst_n77, act_buffer_inst_n76,
         act_buffer_inst_n75, act_buffer_inst_n74, act_buffer_inst_n73,
         act_buffer_inst_n72, act_buffer_inst_n71, act_buffer_inst_n70,
         act_buffer_inst_n69, act_buffer_inst_n68, act_buffer_inst_n67,
         act_buffer_inst_n66, act_buffer_inst_n65, act_buffer_inst_n64,
         act_buffer_inst_n63, act_buffer_inst_n62, act_buffer_inst_n61,
         act_buffer_inst_n60, act_buffer_inst_n59, act_buffer_inst_n58,
         act_buffer_inst_n57, act_buffer_inst_n56, act_buffer_inst_n55,
         act_buffer_inst_n54, act_buffer_inst_n53, act_buffer_inst_n52,
         act_buffer_inst_n51, act_buffer_inst_n50, act_buffer_inst_n49,
         act_buffer_inst_n48, act_buffer_inst_n47, act_buffer_inst_n46,
         act_buffer_inst_n45, act_buffer_inst_n44, act_buffer_inst_n43,
         act_buffer_inst_n42, act_buffer_inst_n41, act_buffer_inst_n40,
         act_buffer_inst_n39, act_buffer_inst_n38, act_buffer_inst_n37,
         act_buffer_inst_n36, act_buffer_inst_n35, act_buffer_inst_n34,
         act_buffer_inst_n33, act_buffer_inst_n32, act_buffer_inst_n31,
         act_buffer_inst_n30, act_buffer_inst_n29, act_buffer_inst_n28,
         act_buffer_inst_n27, act_buffer_inst_n26, act_buffer_inst_n25,
         act_buffer_inst_n24, act_buffer_inst_n23, act_buffer_inst_n22,
         act_buffer_inst_n21, act_buffer_inst_n20, act_buffer_inst_n19,
         act_buffer_inst_n18, act_buffer_inst_n17, act_buffer_inst_n16,
         act_buffer_inst_n15, act_buffer_inst_n14, act_buffer_inst_n13,
         act_buffer_inst_n12, act_buffer_inst_n11, act_buffer_inst_n10,
         act_buffer_inst_net4552, act_buffer_inst_net4547,
         act_buffer_inst_net4542, act_buffer_inst_net4537,
         act_buffer_inst_net4532, act_buffer_inst_net4527,
         act_buffer_inst_net4522, act_buffer_inst_net4517,
         act_buffer_inst_net4512, act_buffer_inst_net4507,
         act_buffer_inst_net4502, act_buffer_inst_net4497,
         act_buffer_inst_net4492, act_buffer_inst_net4487,
         act_buffer_inst_net4482, act_buffer_inst_net4477,
         act_buffer_inst_net4472, act_buffer_inst_net4467,
         act_buffer_inst_net4462, act_buffer_inst_net4457,
         act_buffer_inst_net4452, act_buffer_inst_net4447,
         act_buffer_inst_net4442, act_buffer_inst_net4437,
         act_buffer_inst_net4432, act_buffer_inst_net4427,
         act_buffer_inst_net4422, act_buffer_inst_net4417,
         act_buffer_inst_net4412, act_buffer_inst_net4407,
         act_buffer_inst_net4402, act_buffer_inst_net4397,
         act_buffer_inst_net4392, act_buffer_inst_net4387,
         act_buffer_inst_net4382, act_buffer_inst_net4377,
         act_buffer_inst_net4372, act_buffer_inst_net4367,
         act_buffer_inst_net4362, act_buffer_inst_net4357,
         act_buffer_inst_net4352, act_buffer_inst_net4347,
         act_buffer_inst_net4342, act_buffer_inst_net4337,
         act_buffer_inst_net4332, act_buffer_inst_net4327,
         act_buffer_inst_net4322, act_buffer_inst_net4316,
         act_buffer_inst_N162, act_buffer_inst_N161, act_buffer_inst_N160,
         act_buffer_inst_N159, act_buffer_inst_N158, act_buffer_inst_N157,
         act_buffer_inst_N156, act_buffer_inst_N155, act_buffer_inst_N154,
         act_buffer_inst_N153, act_buffer_inst_N152, act_buffer_inst_N151,
         act_buffer_inst_N150, act_buffer_inst_N149, act_buffer_inst_N148,
         act_buffer_inst_N147, act_buffer_inst_N146, act_buffer_inst_N145,
         act_buffer_inst_N144, act_buffer_inst_N143, act_buffer_inst_N142,
         act_buffer_inst_N141, act_buffer_inst_N140, act_buffer_inst_N139,
         act_buffer_inst_N138, act_buffer_inst_N137, act_buffer_inst_N136,
         act_buffer_inst_N135, act_buffer_inst_N134, act_buffer_inst_N133,
         act_buffer_inst_N132, act_buffer_inst_N131, act_buffer_inst_N130,
         act_buffer_inst_N129, act_buffer_inst_N128, act_buffer_inst_N127,
         act_buffer_inst_N126, act_buffer_inst_N125, act_buffer_inst_N124,
         act_buffer_inst_N123, act_buffer_inst_N122, act_buffer_inst_N121,
         act_buffer_inst_N120, act_buffer_inst_N119, act_buffer_inst_N118,
         act_buffer_inst_N117, act_buffer_inst_N116, act_buffer_inst_N115,
         act_if_inst_n312, act_if_inst_n311, act_if_inst_n310,
         act_if_inst_n309, act_if_inst_n308, act_if_inst_n307,
         act_if_inst_n306, act_if_inst_n305, act_if_inst_n304,
         act_if_inst_n303, act_if_inst_n302, act_if_inst_n301,
         act_if_inst_n300, act_if_inst_n299, act_if_inst_n298,
         act_if_inst_n297, act_if_inst_n296, act_if_inst_n295,
         act_if_inst_n294, act_if_inst_n293, act_if_inst_n292,
         act_if_inst_n291, act_if_inst_n290, act_if_inst_n289,
         act_if_inst_n288, act_if_inst_n287, act_if_inst_n286,
         act_if_inst_n285, act_if_inst_n284, act_if_inst_n283,
         act_if_inst_n282, act_if_inst_n281, act_if_inst_n280,
         act_if_inst_n279, act_if_inst_n278, act_if_inst_n277,
         act_if_inst_n276, act_if_inst_n275, act_if_inst_n274,
         act_if_inst_n273, act_if_inst_n272, act_if_inst_n271,
         act_if_inst_n270, act_if_inst_n269, act_if_inst_n268,
         act_if_inst_n267, act_if_inst_n266, act_if_inst_n265,
         act_if_inst_n264, act_if_inst_n263, act_if_inst_n262,
         act_if_inst_n261, act_if_inst_n260, act_if_inst_n259,
         act_if_inst_n258, act_if_inst_n257, act_if_inst_n256,
         act_if_inst_n255, act_if_inst_n254, act_if_inst_n253,
         act_if_inst_n252, act_if_inst_n251, act_if_inst_n250,
         act_if_inst_n249, act_if_inst_n248, act_if_inst_n247,
         act_if_inst_n246, act_if_inst_n245, act_if_inst_n244,
         act_if_inst_n243, act_if_inst_n242, act_if_inst_n241,
         act_if_inst_n240, act_if_inst_n239, act_if_inst_n238,
         act_if_inst_n237, act_if_inst_n236, act_if_inst_n235,
         act_if_inst_n234, act_if_inst_n233, act_if_inst_n232,
         act_if_inst_n231, act_if_inst_n230, act_if_inst_n229,
         act_if_inst_n228, act_if_inst_n227, act_if_inst_n226,
         act_if_inst_n225, act_if_inst_n224, act_if_inst_n223,
         act_if_inst_n222, act_if_inst_n221, act_if_inst_n220,
         act_if_inst_n219, act_if_inst_n218, act_if_inst_n217,
         act_if_inst_n216, act_if_inst_n215, act_if_inst_n214,
         act_if_inst_n213, act_if_inst_n212, act_if_inst_n211,
         act_if_inst_n210, act_if_inst_n209, act_if_inst_n208,
         act_if_inst_n207, act_if_inst_n206, act_if_inst_n205,
         act_if_inst_n204, act_if_inst_n203, act_if_inst_n202,
         act_if_inst_n201, act_if_inst_n200, act_if_inst_n199,
         act_if_inst_n198, act_if_inst_n197, act_if_inst_n196,
         act_if_inst_n195, act_if_inst_n194, act_if_inst_n193,
         act_if_inst_n192, act_if_inst_n191, act_if_inst_n190,
         act_if_inst_n189, act_if_inst_n188, act_if_inst_n187,
         act_if_inst_n186, act_if_inst_n185, act_if_inst_n184,
         act_if_inst_n183, act_if_inst_n182, act_if_inst_n181,
         act_if_inst_n180, act_if_inst_n179, act_if_inst_n178,
         act_if_inst_n177, act_if_inst_n176, act_if_inst_n175,
         act_if_inst_n174, act_if_inst_n173, act_if_inst_n172,
         act_if_inst_n171, act_if_inst_n170, act_if_inst_n169,
         act_if_inst_n168, act_if_inst_n167, act_if_inst_n166,
         act_if_inst_n165, act_if_inst_n164, act_if_inst_n163,
         act_if_inst_n162, act_if_inst_n161, act_if_inst_n160,
         act_if_inst_n159, act_if_inst_n158, act_if_inst_n157,
         act_if_inst_n156, act_if_inst_n155, act_if_inst_n154,
         act_if_inst_n153, act_if_inst_n152, act_if_inst_n151,
         act_if_inst_n150, act_if_inst_n149, act_if_inst_n148,
         act_if_inst_n147, act_if_inst_n146, act_if_inst_n145,
         act_if_inst_n144, act_if_inst_n143, act_if_inst_n142,
         act_if_inst_n141, act_if_inst_n140, act_if_inst_n139,
         act_if_inst_n138, act_if_inst_n137, act_if_inst_n136,
         act_if_inst_n135, act_if_inst_n134, act_if_inst_n133,
         act_if_inst_n132, act_if_inst_n131, act_if_inst_n130,
         act_if_inst_n129, act_if_inst_n128, act_if_inst_n127,
         act_if_inst_n126, act_if_inst_n125, act_if_inst_n124,
         act_if_inst_n123, act_if_inst_n122, act_if_inst_n121,
         act_if_inst_n120, act_if_inst_n119, act_if_inst_n118,
         act_if_inst_n117, act_if_inst_n116, act_if_inst_n115,
         act_if_inst_n114, act_if_inst_n113, act_if_inst_n112,
         act_if_inst_n111, act_if_inst_n110, act_if_inst_n109,
         act_if_inst_n108, act_if_inst_n107, act_if_inst_n106,
         act_if_inst_n105, act_if_inst_n104, act_if_inst_n103,
         act_if_inst_n102, act_if_inst_n101, act_if_inst_n100, act_if_inst_n99,
         act_if_inst_n98, act_if_inst_n97, act_if_inst_n96, act_if_inst_n95,
         act_if_inst_n94, act_if_inst_n93, act_if_inst_n92, act_if_inst_n91,
         act_if_inst_n90, act_if_inst_n89, act_if_inst_n88, act_if_inst_n87,
         act_if_inst_n86, act_if_inst_n85, act_if_inst_n84, act_if_inst_n83,
         act_if_inst_n82, act_if_inst_n81, act_if_inst_n80, act_if_inst_n79,
         act_if_inst_n78, act_if_inst_n77, act_if_inst_n76, act_if_inst_n75,
         act_if_inst_n74, act_if_inst_n73, act_if_inst_n72, act_if_inst_n71,
         act_if_inst_n70, act_if_inst_n69, act_if_inst_n68, act_if_inst_n67,
         act_if_inst_n66, act_if_inst_n65, act_if_inst_n64, act_if_inst_n63,
         act_if_inst_n62, act_if_inst_n61, act_if_inst_n60, act_if_inst_n59,
         act_if_inst_n58, act_if_inst_n57, act_if_inst_n56, act_if_inst_n55,
         act_if_inst_n54, act_if_inst_n53, act_if_inst_n52, act_if_inst_n51,
         act_if_inst_n50, act_if_inst_n49, act_if_inst_n48, act_if_inst_n47,
         act_if_inst_n46, act_if_inst_n45, act_if_inst_n44, act_if_inst_n43,
         act_if_inst_n42, act_if_inst_n41, act_if_inst_n40, act_if_inst_n39,
         act_if_inst_n2, act_if_inst_n1, act_if_inst_n38, act_if_inst_n37,
         act_if_inst_n36, act_if_inst_n35, act_if_inst_n34, act_if_inst_n33,
         act_if_inst_n32, act_if_inst_n31, act_if_inst_n30, act_if_inst_n29,
         act_if_inst_n28, act_if_inst_n27, act_if_inst_n26, act_if_inst_n25,
         act_if_inst_n24, act_if_inst_n23, act_if_inst_n22, act_if_inst_n21,
         act_if_inst_n20, act_if_inst_n19, act_if_inst_n18, act_if_inst_n17,
         act_if_inst_n16, act_if_inst_n15, act_if_inst_n14, act_if_inst_n13,
         act_if_inst_n12, act_if_inst_n11, act_if_inst_n10, act_if_inst_n9,
         act_if_inst_n8, act_if_inst_n7, act_if_inst_n6, act_if_inst_n5,
         act_if_inst_n4, act_if_inst_n3, npu_inst_n143, npu_inst_n142,
         npu_inst_n141, npu_inst_n140, npu_inst_n139, npu_inst_n138,
         npu_inst_n137, npu_inst_n136, npu_inst_n135, npu_inst_n134,
         npu_inst_n133, npu_inst_n132, npu_inst_n131, npu_inst_n130,
         npu_inst_n129, npu_inst_n128, npu_inst_n127, npu_inst_n126,
         npu_inst_n125, npu_inst_n124, npu_inst_n123, npu_inst_n122,
         npu_inst_n121, npu_inst_n120, npu_inst_n119, npu_inst_n118,
         npu_inst_n117, npu_inst_n116, npu_inst_n115, npu_inst_n114,
         npu_inst_n113, npu_inst_n112, npu_inst_n111, npu_inst_n110,
         npu_inst_n109, npu_inst_n108, npu_inst_n107, npu_inst_n106,
         npu_inst_n105, npu_inst_n104, npu_inst_n103, npu_inst_n102,
         npu_inst_n101, npu_inst_n100, npu_inst_n99, npu_inst_n98,
         npu_inst_n97, npu_inst_n96, npu_inst_n95, npu_inst_n94, npu_inst_n93,
         npu_inst_n92, npu_inst_n91, npu_inst_n90, npu_inst_n89, npu_inst_n88,
         npu_inst_n87, npu_inst_n86, npu_inst_n85, npu_inst_n84, npu_inst_n83,
         npu_inst_n82, npu_inst_n81, npu_inst_n80, npu_inst_n79, npu_inst_n78,
         npu_inst_n77, npu_inst_n76, npu_inst_n75, npu_inst_n74, npu_inst_n73,
         npu_inst_n72, npu_inst_n71, npu_inst_n70, npu_inst_n69, npu_inst_n68,
         npu_inst_n67, npu_inst_n66, npu_inst_n65, npu_inst_n64, npu_inst_n63,
         npu_inst_n62, npu_inst_n61, npu_inst_n60, npu_inst_n59, npu_inst_n58,
         npu_inst_n57, npu_inst_n56, npu_inst_n55, npu_inst_n54, npu_inst_n53,
         npu_inst_n52, npu_inst_n51, npu_inst_n50, npu_inst_n49, npu_inst_n48,
         npu_inst_n47, npu_inst_n46, npu_inst_n45, npu_inst_n44, npu_inst_n43,
         npu_inst_n42, npu_inst_n41, npu_inst_n40, npu_inst_n39, npu_inst_n38,
         npu_inst_n37, npu_inst_n36, npu_inst_n35, npu_inst_n34, npu_inst_n33,
         npu_inst_n32, npu_inst_n31, npu_inst_n30, npu_inst_n29, npu_inst_n28,
         npu_inst_n27, npu_inst_n26, npu_inst_n25, npu_inst_n24, npu_inst_n23,
         npu_inst_n22, npu_inst_n21, npu_inst_n20, npu_inst_n19, npu_inst_n18,
         npu_inst_n17, npu_inst_n16, npu_inst_n15, npu_inst_n14, npu_inst_n13,
         npu_inst_n12, npu_inst_n11, npu_inst_n10, npu_inst_n9, npu_inst_n8,
         npu_inst_n7, npu_inst_n6, npu_inst_n5, npu_inst_n4, npu_inst_n3,
         npu_inst_n2, npu_inst_n1, npu_inst_int_data_res_7__7__0_,
         npu_inst_int_data_res_7__7__1_, npu_inst_int_data_res_7__7__2_,
         npu_inst_int_data_res_7__7__3_, npu_inst_int_data_res_7__7__4_,
         npu_inst_int_data_res_7__7__5_, npu_inst_int_data_res_7__7__6_,
         npu_inst_int_data_res_7__7__7_, npu_inst_int_data_res_7__6__0_,
         npu_inst_int_data_res_7__6__1_, npu_inst_int_data_res_7__6__2_,
         npu_inst_int_data_res_7__6__3_, npu_inst_int_data_res_7__6__4_,
         npu_inst_int_data_res_7__6__5_, npu_inst_int_data_res_7__6__6_,
         npu_inst_int_data_res_7__6__7_, npu_inst_int_data_res_7__5__0_,
         npu_inst_int_data_res_7__5__1_, npu_inst_int_data_res_7__5__2_,
         npu_inst_int_data_res_7__5__3_, npu_inst_int_data_res_7__5__4_,
         npu_inst_int_data_res_7__5__5_, npu_inst_int_data_res_7__5__6_,
         npu_inst_int_data_res_7__5__7_, npu_inst_int_data_res_7__4__0_,
         npu_inst_int_data_res_7__4__1_, npu_inst_int_data_res_7__4__2_,
         npu_inst_int_data_res_7__4__3_, npu_inst_int_data_res_7__4__4_,
         npu_inst_int_data_res_7__4__5_, npu_inst_int_data_res_7__4__6_,
         npu_inst_int_data_res_7__4__7_, npu_inst_int_data_res_7__3__0_,
         npu_inst_int_data_res_7__3__1_, npu_inst_int_data_res_7__3__2_,
         npu_inst_int_data_res_7__3__3_, npu_inst_int_data_res_7__3__4_,
         npu_inst_int_data_res_7__3__5_, npu_inst_int_data_res_7__3__6_,
         npu_inst_int_data_res_7__3__7_, npu_inst_int_data_res_7__2__0_,
         npu_inst_int_data_res_7__2__1_, npu_inst_int_data_res_7__2__2_,
         npu_inst_int_data_res_7__2__3_, npu_inst_int_data_res_7__2__4_,
         npu_inst_int_data_res_7__2__5_, npu_inst_int_data_res_7__2__6_,
         npu_inst_int_data_res_7__2__7_, npu_inst_int_data_res_7__1__0_,
         npu_inst_int_data_res_7__1__1_, npu_inst_int_data_res_7__1__2_,
         npu_inst_int_data_res_7__1__3_, npu_inst_int_data_res_7__1__4_,
         npu_inst_int_data_res_7__1__5_, npu_inst_int_data_res_7__1__6_,
         npu_inst_int_data_res_7__1__7_, npu_inst_int_data_res_7__0__0_,
         npu_inst_int_data_res_7__0__1_, npu_inst_int_data_res_7__0__2_,
         npu_inst_int_data_res_7__0__3_, npu_inst_int_data_res_7__0__4_,
         npu_inst_int_data_res_7__0__5_, npu_inst_int_data_res_7__0__6_,
         npu_inst_int_data_res_7__0__7_, npu_inst_int_data_res_6__7__0_,
         npu_inst_int_data_res_6__7__1_, npu_inst_int_data_res_6__7__2_,
         npu_inst_int_data_res_6__7__3_, npu_inst_int_data_res_6__7__4_,
         npu_inst_int_data_res_6__7__5_, npu_inst_int_data_res_6__7__6_,
         npu_inst_int_data_res_6__7__7_, npu_inst_int_data_res_6__6__0_,
         npu_inst_int_data_res_6__6__1_, npu_inst_int_data_res_6__6__2_,
         npu_inst_int_data_res_6__6__3_, npu_inst_int_data_res_6__6__4_,
         npu_inst_int_data_res_6__6__5_, npu_inst_int_data_res_6__6__6_,
         npu_inst_int_data_res_6__6__7_, npu_inst_int_data_res_6__5__0_,
         npu_inst_int_data_res_6__5__1_, npu_inst_int_data_res_6__5__2_,
         npu_inst_int_data_res_6__5__3_, npu_inst_int_data_res_6__5__4_,
         npu_inst_int_data_res_6__5__5_, npu_inst_int_data_res_6__5__6_,
         npu_inst_int_data_res_6__5__7_, npu_inst_int_data_res_6__4__0_,
         npu_inst_int_data_res_6__4__1_, npu_inst_int_data_res_6__4__2_,
         npu_inst_int_data_res_6__4__3_, npu_inst_int_data_res_6__4__4_,
         npu_inst_int_data_res_6__4__5_, npu_inst_int_data_res_6__4__6_,
         npu_inst_int_data_res_6__4__7_, npu_inst_int_data_res_6__3__0_,
         npu_inst_int_data_res_6__3__1_, npu_inst_int_data_res_6__3__2_,
         npu_inst_int_data_res_6__3__3_, npu_inst_int_data_res_6__3__4_,
         npu_inst_int_data_res_6__3__5_, npu_inst_int_data_res_6__3__6_,
         npu_inst_int_data_res_6__3__7_, npu_inst_int_data_res_6__2__0_,
         npu_inst_int_data_res_6__2__1_, npu_inst_int_data_res_6__2__2_,
         npu_inst_int_data_res_6__2__3_, npu_inst_int_data_res_6__2__4_,
         npu_inst_int_data_res_6__2__5_, npu_inst_int_data_res_6__2__6_,
         npu_inst_int_data_res_6__2__7_, npu_inst_int_data_res_6__1__0_,
         npu_inst_int_data_res_6__1__1_, npu_inst_int_data_res_6__1__2_,
         npu_inst_int_data_res_6__1__3_, npu_inst_int_data_res_6__1__4_,
         npu_inst_int_data_res_6__1__5_, npu_inst_int_data_res_6__1__6_,
         npu_inst_int_data_res_6__1__7_, npu_inst_int_data_res_6__0__0_,
         npu_inst_int_data_res_6__0__1_, npu_inst_int_data_res_6__0__2_,
         npu_inst_int_data_res_6__0__3_, npu_inst_int_data_res_6__0__4_,
         npu_inst_int_data_res_6__0__5_, npu_inst_int_data_res_6__0__6_,
         npu_inst_int_data_res_6__0__7_, npu_inst_int_data_res_5__7__0_,
         npu_inst_int_data_res_5__7__1_, npu_inst_int_data_res_5__7__2_,
         npu_inst_int_data_res_5__7__3_, npu_inst_int_data_res_5__7__4_,
         npu_inst_int_data_res_5__7__5_, npu_inst_int_data_res_5__7__6_,
         npu_inst_int_data_res_5__7__7_, npu_inst_int_data_res_5__6__0_,
         npu_inst_int_data_res_5__6__1_, npu_inst_int_data_res_5__6__2_,
         npu_inst_int_data_res_5__6__3_, npu_inst_int_data_res_5__6__4_,
         npu_inst_int_data_res_5__6__5_, npu_inst_int_data_res_5__6__6_,
         npu_inst_int_data_res_5__6__7_, npu_inst_int_data_res_5__5__0_,
         npu_inst_int_data_res_5__5__1_, npu_inst_int_data_res_5__5__2_,
         npu_inst_int_data_res_5__5__3_, npu_inst_int_data_res_5__5__4_,
         npu_inst_int_data_res_5__5__5_, npu_inst_int_data_res_5__5__6_,
         npu_inst_int_data_res_5__5__7_, npu_inst_int_data_res_5__4__0_,
         npu_inst_int_data_res_5__4__1_, npu_inst_int_data_res_5__4__2_,
         npu_inst_int_data_res_5__4__3_, npu_inst_int_data_res_5__4__4_,
         npu_inst_int_data_res_5__4__5_, npu_inst_int_data_res_5__4__6_,
         npu_inst_int_data_res_5__4__7_, npu_inst_int_data_res_5__3__0_,
         npu_inst_int_data_res_5__3__1_, npu_inst_int_data_res_5__3__2_,
         npu_inst_int_data_res_5__3__3_, npu_inst_int_data_res_5__3__4_,
         npu_inst_int_data_res_5__3__5_, npu_inst_int_data_res_5__3__6_,
         npu_inst_int_data_res_5__3__7_, npu_inst_int_data_res_5__2__0_,
         npu_inst_int_data_res_5__2__1_, npu_inst_int_data_res_5__2__2_,
         npu_inst_int_data_res_5__2__3_, npu_inst_int_data_res_5__2__4_,
         npu_inst_int_data_res_5__2__5_, npu_inst_int_data_res_5__2__6_,
         npu_inst_int_data_res_5__2__7_, npu_inst_int_data_res_5__1__0_,
         npu_inst_int_data_res_5__1__1_, npu_inst_int_data_res_5__1__2_,
         npu_inst_int_data_res_5__1__3_, npu_inst_int_data_res_5__1__4_,
         npu_inst_int_data_res_5__1__5_, npu_inst_int_data_res_5__1__6_,
         npu_inst_int_data_res_5__1__7_, npu_inst_int_data_res_5__0__0_,
         npu_inst_int_data_res_5__0__1_, npu_inst_int_data_res_5__0__2_,
         npu_inst_int_data_res_5__0__3_, npu_inst_int_data_res_5__0__4_,
         npu_inst_int_data_res_5__0__5_, npu_inst_int_data_res_5__0__6_,
         npu_inst_int_data_res_5__0__7_, npu_inst_int_data_res_4__7__0_,
         npu_inst_int_data_res_4__7__1_, npu_inst_int_data_res_4__7__2_,
         npu_inst_int_data_res_4__7__3_, npu_inst_int_data_res_4__7__4_,
         npu_inst_int_data_res_4__7__5_, npu_inst_int_data_res_4__7__6_,
         npu_inst_int_data_res_4__7__7_, npu_inst_int_data_res_4__6__0_,
         npu_inst_int_data_res_4__6__1_, npu_inst_int_data_res_4__6__2_,
         npu_inst_int_data_res_4__6__3_, npu_inst_int_data_res_4__6__4_,
         npu_inst_int_data_res_4__6__5_, npu_inst_int_data_res_4__6__6_,
         npu_inst_int_data_res_4__6__7_, npu_inst_int_data_res_4__5__0_,
         npu_inst_int_data_res_4__5__1_, npu_inst_int_data_res_4__5__2_,
         npu_inst_int_data_res_4__5__3_, npu_inst_int_data_res_4__5__4_,
         npu_inst_int_data_res_4__5__5_, npu_inst_int_data_res_4__5__6_,
         npu_inst_int_data_res_4__5__7_, npu_inst_int_data_res_4__4__0_,
         npu_inst_int_data_res_4__4__1_, npu_inst_int_data_res_4__4__2_,
         npu_inst_int_data_res_4__4__3_, npu_inst_int_data_res_4__4__4_,
         npu_inst_int_data_res_4__4__5_, npu_inst_int_data_res_4__4__6_,
         npu_inst_int_data_res_4__4__7_, npu_inst_int_data_res_4__3__0_,
         npu_inst_int_data_res_4__3__1_, npu_inst_int_data_res_4__3__2_,
         npu_inst_int_data_res_4__3__3_, npu_inst_int_data_res_4__3__4_,
         npu_inst_int_data_res_4__3__5_, npu_inst_int_data_res_4__3__6_,
         npu_inst_int_data_res_4__3__7_, npu_inst_int_data_res_4__2__0_,
         npu_inst_int_data_res_4__2__1_, npu_inst_int_data_res_4__2__2_,
         npu_inst_int_data_res_4__2__3_, npu_inst_int_data_res_4__2__4_,
         npu_inst_int_data_res_4__2__5_, npu_inst_int_data_res_4__2__6_,
         npu_inst_int_data_res_4__2__7_, npu_inst_int_data_res_4__1__0_,
         npu_inst_int_data_res_4__1__1_, npu_inst_int_data_res_4__1__2_,
         npu_inst_int_data_res_4__1__3_, npu_inst_int_data_res_4__1__4_,
         npu_inst_int_data_res_4__1__5_, npu_inst_int_data_res_4__1__6_,
         npu_inst_int_data_res_4__1__7_, npu_inst_int_data_res_4__0__0_,
         npu_inst_int_data_res_4__0__1_, npu_inst_int_data_res_4__0__2_,
         npu_inst_int_data_res_4__0__3_, npu_inst_int_data_res_4__0__4_,
         npu_inst_int_data_res_4__0__5_, npu_inst_int_data_res_4__0__6_,
         npu_inst_int_data_res_4__0__7_, npu_inst_int_data_res_3__7__0_,
         npu_inst_int_data_res_3__7__1_, npu_inst_int_data_res_3__7__2_,
         npu_inst_int_data_res_3__7__3_, npu_inst_int_data_res_3__7__4_,
         npu_inst_int_data_res_3__7__5_, npu_inst_int_data_res_3__7__6_,
         npu_inst_int_data_res_3__7__7_, npu_inst_int_data_res_3__6__0_,
         npu_inst_int_data_res_3__6__1_, npu_inst_int_data_res_3__6__2_,
         npu_inst_int_data_res_3__6__3_, npu_inst_int_data_res_3__6__4_,
         npu_inst_int_data_res_3__6__5_, npu_inst_int_data_res_3__6__6_,
         npu_inst_int_data_res_3__6__7_, npu_inst_int_data_res_3__5__0_,
         npu_inst_int_data_res_3__5__1_, npu_inst_int_data_res_3__5__2_,
         npu_inst_int_data_res_3__5__3_, npu_inst_int_data_res_3__5__4_,
         npu_inst_int_data_res_3__5__5_, npu_inst_int_data_res_3__5__6_,
         npu_inst_int_data_res_3__5__7_, npu_inst_int_data_res_3__4__0_,
         npu_inst_int_data_res_3__4__1_, npu_inst_int_data_res_3__4__2_,
         npu_inst_int_data_res_3__4__3_, npu_inst_int_data_res_3__4__4_,
         npu_inst_int_data_res_3__4__5_, npu_inst_int_data_res_3__4__6_,
         npu_inst_int_data_res_3__4__7_, npu_inst_int_data_res_3__3__0_,
         npu_inst_int_data_res_3__3__1_, npu_inst_int_data_res_3__3__2_,
         npu_inst_int_data_res_3__3__3_, npu_inst_int_data_res_3__3__4_,
         npu_inst_int_data_res_3__3__5_, npu_inst_int_data_res_3__3__6_,
         npu_inst_int_data_res_3__3__7_, npu_inst_int_data_res_3__2__0_,
         npu_inst_int_data_res_3__2__1_, npu_inst_int_data_res_3__2__2_,
         npu_inst_int_data_res_3__2__3_, npu_inst_int_data_res_3__2__4_,
         npu_inst_int_data_res_3__2__5_, npu_inst_int_data_res_3__2__6_,
         npu_inst_int_data_res_3__2__7_, npu_inst_int_data_res_3__1__0_,
         npu_inst_int_data_res_3__1__1_, npu_inst_int_data_res_3__1__2_,
         npu_inst_int_data_res_3__1__3_, npu_inst_int_data_res_3__1__4_,
         npu_inst_int_data_res_3__1__5_, npu_inst_int_data_res_3__1__6_,
         npu_inst_int_data_res_3__1__7_, npu_inst_int_data_res_3__0__0_,
         npu_inst_int_data_res_3__0__1_, npu_inst_int_data_res_3__0__2_,
         npu_inst_int_data_res_3__0__3_, npu_inst_int_data_res_3__0__4_,
         npu_inst_int_data_res_3__0__5_, npu_inst_int_data_res_3__0__6_,
         npu_inst_int_data_res_3__0__7_, npu_inst_int_data_res_2__7__0_,
         npu_inst_int_data_res_2__7__1_, npu_inst_int_data_res_2__7__2_,
         npu_inst_int_data_res_2__7__3_, npu_inst_int_data_res_2__7__4_,
         npu_inst_int_data_res_2__7__5_, npu_inst_int_data_res_2__7__6_,
         npu_inst_int_data_res_2__7__7_, npu_inst_int_data_res_2__6__0_,
         npu_inst_int_data_res_2__6__1_, npu_inst_int_data_res_2__6__2_,
         npu_inst_int_data_res_2__6__3_, npu_inst_int_data_res_2__6__4_,
         npu_inst_int_data_res_2__6__5_, npu_inst_int_data_res_2__6__6_,
         npu_inst_int_data_res_2__6__7_, npu_inst_int_data_res_2__5__0_,
         npu_inst_int_data_res_2__5__1_, npu_inst_int_data_res_2__5__2_,
         npu_inst_int_data_res_2__5__3_, npu_inst_int_data_res_2__5__4_,
         npu_inst_int_data_res_2__5__5_, npu_inst_int_data_res_2__5__6_,
         npu_inst_int_data_res_2__5__7_, npu_inst_int_data_res_2__4__0_,
         npu_inst_int_data_res_2__4__1_, npu_inst_int_data_res_2__4__2_,
         npu_inst_int_data_res_2__4__3_, npu_inst_int_data_res_2__4__4_,
         npu_inst_int_data_res_2__4__5_, npu_inst_int_data_res_2__4__6_,
         npu_inst_int_data_res_2__4__7_, npu_inst_int_data_res_2__3__0_,
         npu_inst_int_data_res_2__3__1_, npu_inst_int_data_res_2__3__2_,
         npu_inst_int_data_res_2__3__3_, npu_inst_int_data_res_2__3__4_,
         npu_inst_int_data_res_2__3__5_, npu_inst_int_data_res_2__3__6_,
         npu_inst_int_data_res_2__3__7_, npu_inst_int_data_res_2__2__0_,
         npu_inst_int_data_res_2__2__1_, npu_inst_int_data_res_2__2__2_,
         npu_inst_int_data_res_2__2__3_, npu_inst_int_data_res_2__2__4_,
         npu_inst_int_data_res_2__2__5_, npu_inst_int_data_res_2__2__6_,
         npu_inst_int_data_res_2__2__7_, npu_inst_int_data_res_2__1__0_,
         npu_inst_int_data_res_2__1__1_, npu_inst_int_data_res_2__1__2_,
         npu_inst_int_data_res_2__1__3_, npu_inst_int_data_res_2__1__4_,
         npu_inst_int_data_res_2__1__5_, npu_inst_int_data_res_2__1__6_,
         npu_inst_int_data_res_2__1__7_, npu_inst_int_data_res_2__0__0_,
         npu_inst_int_data_res_2__0__1_, npu_inst_int_data_res_2__0__2_,
         npu_inst_int_data_res_2__0__3_, npu_inst_int_data_res_2__0__4_,
         npu_inst_int_data_res_2__0__5_, npu_inst_int_data_res_2__0__6_,
         npu_inst_int_data_res_2__0__7_, npu_inst_int_data_res_1__7__0_,
         npu_inst_int_data_res_1__7__1_, npu_inst_int_data_res_1__7__2_,
         npu_inst_int_data_res_1__7__3_, npu_inst_int_data_res_1__7__4_,
         npu_inst_int_data_res_1__7__5_, npu_inst_int_data_res_1__7__6_,
         npu_inst_int_data_res_1__7__7_, npu_inst_int_data_res_1__6__0_,
         npu_inst_int_data_res_1__6__1_, npu_inst_int_data_res_1__6__2_,
         npu_inst_int_data_res_1__6__3_, npu_inst_int_data_res_1__6__4_,
         npu_inst_int_data_res_1__6__5_, npu_inst_int_data_res_1__6__6_,
         npu_inst_int_data_res_1__6__7_, npu_inst_int_data_res_1__5__0_,
         npu_inst_int_data_res_1__5__1_, npu_inst_int_data_res_1__5__2_,
         npu_inst_int_data_res_1__5__3_, npu_inst_int_data_res_1__5__4_,
         npu_inst_int_data_res_1__5__5_, npu_inst_int_data_res_1__5__6_,
         npu_inst_int_data_res_1__5__7_, npu_inst_int_data_res_1__4__0_,
         npu_inst_int_data_res_1__4__1_, npu_inst_int_data_res_1__4__2_,
         npu_inst_int_data_res_1__4__3_, npu_inst_int_data_res_1__4__4_,
         npu_inst_int_data_res_1__4__5_, npu_inst_int_data_res_1__4__6_,
         npu_inst_int_data_res_1__4__7_, npu_inst_int_data_res_1__3__0_,
         npu_inst_int_data_res_1__3__1_, npu_inst_int_data_res_1__3__2_,
         npu_inst_int_data_res_1__3__3_, npu_inst_int_data_res_1__3__4_,
         npu_inst_int_data_res_1__3__5_, npu_inst_int_data_res_1__3__6_,
         npu_inst_int_data_res_1__3__7_, npu_inst_int_data_res_1__2__0_,
         npu_inst_int_data_res_1__2__1_, npu_inst_int_data_res_1__2__2_,
         npu_inst_int_data_res_1__2__3_, npu_inst_int_data_res_1__2__4_,
         npu_inst_int_data_res_1__2__5_, npu_inst_int_data_res_1__2__6_,
         npu_inst_int_data_res_1__2__7_, npu_inst_int_data_res_1__1__0_,
         npu_inst_int_data_res_1__1__1_, npu_inst_int_data_res_1__1__2_,
         npu_inst_int_data_res_1__1__3_, npu_inst_int_data_res_1__1__4_,
         npu_inst_int_data_res_1__1__5_, npu_inst_int_data_res_1__1__6_,
         npu_inst_int_data_res_1__1__7_, npu_inst_int_data_res_1__0__0_,
         npu_inst_int_data_res_1__0__1_, npu_inst_int_data_res_1__0__2_,
         npu_inst_int_data_res_1__0__3_, npu_inst_int_data_res_1__0__4_,
         npu_inst_int_data_res_1__0__5_, npu_inst_int_data_res_1__0__6_,
         npu_inst_int_data_res_1__0__7_, npu_inst_int_data_y_7__7__0_,
         npu_inst_int_data_y_7__7__1_, npu_inst_int_data_y_7__6__0_,
         npu_inst_int_data_y_7__6__1_, npu_inst_int_data_y_7__5__0_,
         npu_inst_int_data_y_7__5__1_, npu_inst_int_data_y_7__4__0_,
         npu_inst_int_data_y_7__4__1_, npu_inst_int_data_y_7__3__0_,
         npu_inst_int_data_y_7__3__1_, npu_inst_int_data_y_7__2__0_,
         npu_inst_int_data_y_7__2__1_, npu_inst_int_data_y_7__1__0_,
         npu_inst_int_data_y_7__1__1_, npu_inst_int_data_y_7__0__0_,
         npu_inst_int_data_y_7__0__1_, npu_inst_int_data_y_6__7__0_,
         npu_inst_int_data_y_6__7__1_, npu_inst_int_data_y_6__6__0_,
         npu_inst_int_data_y_6__6__1_, npu_inst_int_data_y_6__5__0_,
         npu_inst_int_data_y_6__5__1_, npu_inst_int_data_y_6__4__0_,
         npu_inst_int_data_y_6__4__1_, npu_inst_int_data_y_6__3__0_,
         npu_inst_int_data_y_6__3__1_, npu_inst_int_data_y_6__2__0_,
         npu_inst_int_data_y_6__2__1_, npu_inst_int_data_y_6__1__0_,
         npu_inst_int_data_y_6__1__1_, npu_inst_int_data_y_6__0__0_,
         npu_inst_int_data_y_6__0__1_, npu_inst_int_data_y_5__7__0_,
         npu_inst_int_data_y_5__7__1_, npu_inst_int_data_y_5__6__0_,
         npu_inst_int_data_y_5__6__1_, npu_inst_int_data_y_5__5__0_,
         npu_inst_int_data_y_5__5__1_, npu_inst_int_data_y_5__4__0_,
         npu_inst_int_data_y_5__4__1_, npu_inst_int_data_y_5__3__0_,
         npu_inst_int_data_y_5__3__1_, npu_inst_int_data_y_5__2__0_,
         npu_inst_int_data_y_5__2__1_, npu_inst_int_data_y_5__1__0_,
         npu_inst_int_data_y_5__1__1_, npu_inst_int_data_y_5__0__0_,
         npu_inst_int_data_y_5__0__1_, npu_inst_int_data_y_4__7__0_,
         npu_inst_int_data_y_4__7__1_, npu_inst_int_data_y_4__6__0_,
         npu_inst_int_data_y_4__6__1_, npu_inst_int_data_y_4__5__0_,
         npu_inst_int_data_y_4__5__1_, npu_inst_int_data_y_4__4__0_,
         npu_inst_int_data_y_4__4__1_, npu_inst_int_data_y_4__3__0_,
         npu_inst_int_data_y_4__3__1_, npu_inst_int_data_y_4__2__0_,
         npu_inst_int_data_y_4__2__1_, npu_inst_int_data_y_4__1__0_,
         npu_inst_int_data_y_4__1__1_, npu_inst_int_data_y_4__0__0_,
         npu_inst_int_data_y_4__0__1_, npu_inst_int_data_y_3__7__0_,
         npu_inst_int_data_y_3__7__1_, npu_inst_int_data_y_3__6__0_,
         npu_inst_int_data_y_3__6__1_, npu_inst_int_data_y_3__5__0_,
         npu_inst_int_data_y_3__5__1_, npu_inst_int_data_y_3__4__0_,
         npu_inst_int_data_y_3__4__1_, npu_inst_int_data_y_3__3__0_,
         npu_inst_int_data_y_3__3__1_, npu_inst_int_data_y_3__2__0_,
         npu_inst_int_data_y_3__2__1_, npu_inst_int_data_y_3__1__0_,
         npu_inst_int_data_y_3__1__1_, npu_inst_int_data_y_3__0__0_,
         npu_inst_int_data_y_3__0__1_, npu_inst_int_data_y_2__7__0_,
         npu_inst_int_data_y_2__7__1_, npu_inst_int_data_y_2__6__0_,
         npu_inst_int_data_y_2__6__1_, npu_inst_int_data_y_2__5__0_,
         npu_inst_int_data_y_2__5__1_, npu_inst_int_data_y_2__4__0_,
         npu_inst_int_data_y_2__4__1_, npu_inst_int_data_y_2__3__0_,
         npu_inst_int_data_y_2__3__1_, npu_inst_int_data_y_2__2__0_,
         npu_inst_int_data_y_2__2__1_, npu_inst_int_data_y_2__1__0_,
         npu_inst_int_data_y_2__1__1_, npu_inst_int_data_y_2__0__0_,
         npu_inst_int_data_y_2__0__1_, npu_inst_int_data_y_1__7__0_,
         npu_inst_int_data_y_1__7__1_, npu_inst_int_data_y_1__6__0_,
         npu_inst_int_data_y_1__6__1_, npu_inst_int_data_y_1__5__0_,
         npu_inst_int_data_y_1__5__1_, npu_inst_int_data_y_1__4__0_,
         npu_inst_int_data_y_1__4__1_, npu_inst_int_data_y_1__3__0_,
         npu_inst_int_data_y_1__3__1_, npu_inst_int_data_y_1__2__0_,
         npu_inst_int_data_y_1__2__1_, npu_inst_int_data_y_1__1__0_,
         npu_inst_int_data_y_1__1__1_, npu_inst_int_data_y_1__0__0_,
         npu_inst_int_data_y_1__0__1_, npu_inst_int_data_x_7__7__0_,
         npu_inst_int_data_x_7__7__1_, npu_inst_int_data_x_7__6__0_,
         npu_inst_int_data_x_7__6__1_, npu_inst_int_data_x_7__5__0_,
         npu_inst_int_data_x_7__5__1_, npu_inst_int_data_x_7__4__0_,
         npu_inst_int_data_x_7__4__1_, npu_inst_int_data_x_7__3__0_,
         npu_inst_int_data_x_7__3__1_, npu_inst_int_data_x_7__2__0_,
         npu_inst_int_data_x_7__2__1_, npu_inst_int_data_x_7__1__0_,
         npu_inst_int_data_x_7__1__1_, npu_inst_int_data_x_6__7__0_,
         npu_inst_int_data_x_6__7__1_, npu_inst_int_data_x_6__6__0_,
         npu_inst_int_data_x_6__6__1_, npu_inst_int_data_x_6__5__0_,
         npu_inst_int_data_x_6__5__1_, npu_inst_int_data_x_6__4__0_,
         npu_inst_int_data_x_6__4__1_, npu_inst_int_data_x_6__3__0_,
         npu_inst_int_data_x_6__3__1_, npu_inst_int_data_x_6__2__0_,
         npu_inst_int_data_x_6__2__1_, npu_inst_int_data_x_6__1__0_,
         npu_inst_int_data_x_6__1__1_, npu_inst_int_data_x_5__7__0_,
         npu_inst_int_data_x_5__7__1_, npu_inst_int_data_x_5__6__0_,
         npu_inst_int_data_x_5__6__1_, npu_inst_int_data_x_5__5__0_,
         npu_inst_int_data_x_5__5__1_, npu_inst_int_data_x_5__4__0_,
         npu_inst_int_data_x_5__4__1_, npu_inst_int_data_x_5__3__0_,
         npu_inst_int_data_x_5__3__1_, npu_inst_int_data_x_5__2__0_,
         npu_inst_int_data_x_5__2__1_, npu_inst_int_data_x_5__1__0_,
         npu_inst_int_data_x_5__1__1_, npu_inst_int_data_x_4__7__0_,
         npu_inst_int_data_x_4__7__1_, npu_inst_int_data_x_4__6__0_,
         npu_inst_int_data_x_4__6__1_, npu_inst_int_data_x_4__5__0_,
         npu_inst_int_data_x_4__5__1_, npu_inst_int_data_x_4__4__0_,
         npu_inst_int_data_x_4__4__1_, npu_inst_int_data_x_4__3__0_,
         npu_inst_int_data_x_4__3__1_, npu_inst_int_data_x_4__2__0_,
         npu_inst_int_data_x_4__2__1_, npu_inst_int_data_x_4__1__0_,
         npu_inst_int_data_x_4__1__1_, npu_inst_int_data_x_3__7__0_,
         npu_inst_int_data_x_3__7__1_, npu_inst_int_data_x_3__6__0_,
         npu_inst_int_data_x_3__6__1_, npu_inst_int_data_x_3__5__0_,
         npu_inst_int_data_x_3__5__1_, npu_inst_int_data_x_3__4__0_,
         npu_inst_int_data_x_3__4__1_, npu_inst_int_data_x_3__3__0_,
         npu_inst_int_data_x_3__3__1_, npu_inst_int_data_x_3__2__0_,
         npu_inst_int_data_x_3__2__1_, npu_inst_int_data_x_3__1__0_,
         npu_inst_int_data_x_3__1__1_, npu_inst_int_data_x_2__7__0_,
         npu_inst_int_data_x_2__7__1_, npu_inst_int_data_x_2__6__0_,
         npu_inst_int_data_x_2__6__1_, npu_inst_int_data_x_2__5__0_,
         npu_inst_int_data_x_2__5__1_, npu_inst_int_data_x_2__4__0_,
         npu_inst_int_data_x_2__4__1_, npu_inst_int_data_x_2__3__0_,
         npu_inst_int_data_x_2__3__1_, npu_inst_int_data_x_2__2__0_,
         npu_inst_int_data_x_2__2__1_, npu_inst_int_data_x_2__1__0_,
         npu_inst_int_data_x_2__1__1_, npu_inst_int_data_x_1__7__0_,
         npu_inst_int_data_x_1__7__1_, npu_inst_int_data_x_1__6__0_,
         npu_inst_int_data_x_1__6__1_, npu_inst_int_data_x_1__5__0_,
         npu_inst_int_data_x_1__5__1_, npu_inst_int_data_x_1__4__0_,
         npu_inst_int_data_x_1__4__1_, npu_inst_int_data_x_1__3__0_,
         npu_inst_int_data_x_1__3__1_, npu_inst_int_data_x_1__2__0_,
         npu_inst_int_data_x_1__2__1_, npu_inst_int_data_x_1__1__0_,
         npu_inst_int_data_x_1__1__1_, npu_inst_int_data_x_0__7__0_,
         npu_inst_int_data_x_0__7__1_, npu_inst_int_data_x_0__6__0_,
         npu_inst_int_data_x_0__6__1_, npu_inst_int_data_x_0__5__0_,
         npu_inst_int_data_x_0__5__1_, npu_inst_int_data_x_0__4__0_,
         npu_inst_int_data_x_0__4__1_, npu_inst_int_data_x_0__3__0_,
         npu_inst_int_data_x_0__3__1_, npu_inst_int_data_x_0__2__0_,
         npu_inst_int_data_x_0__2__1_, npu_inst_int_data_x_0__1__0_,
         npu_inst_int_data_x_0__1__1_, npu_inst_pe_1_0_0_n118,
         npu_inst_pe_1_0_0_n117, npu_inst_pe_1_0_0_n116,
         npu_inst_pe_1_0_0_n115, npu_inst_pe_1_0_0_n114,
         npu_inst_pe_1_0_0_n113, npu_inst_pe_1_0_0_n112,
         npu_inst_pe_1_0_0_n111, npu_inst_pe_1_0_0_n110,
         npu_inst_pe_1_0_0_n109, npu_inst_pe_1_0_0_n108,
         npu_inst_pe_1_0_0_n107, npu_inst_pe_1_0_0_n106,
         npu_inst_pe_1_0_0_n105, npu_inst_pe_1_0_0_n104,
         npu_inst_pe_1_0_0_n103, npu_inst_pe_1_0_0_n102,
         npu_inst_pe_1_0_0_n101, npu_inst_pe_1_0_0_n100, npu_inst_pe_1_0_0_n99,
         npu_inst_pe_1_0_0_n98, npu_inst_pe_1_0_0_n36, npu_inst_pe_1_0_0_n35,
         npu_inst_pe_1_0_0_n34, npu_inst_pe_1_0_0_n33, npu_inst_pe_1_0_0_n32,
         npu_inst_pe_1_0_0_n31, npu_inst_pe_1_0_0_n30, npu_inst_pe_1_0_0_n29,
         npu_inst_pe_1_0_0_n28, npu_inst_pe_1_0_0_n25, npu_inst_pe_1_0_0_n24,
         npu_inst_pe_1_0_0_n23, npu_inst_pe_1_0_0_n22, npu_inst_pe_1_0_0_n21,
         npu_inst_pe_1_0_0_n20, npu_inst_pe_1_0_0_n19, npu_inst_pe_1_0_0_n18,
         npu_inst_pe_1_0_0_n17, npu_inst_pe_1_0_0_n16, npu_inst_pe_1_0_0_n15,
         npu_inst_pe_1_0_0_n14, npu_inst_pe_1_0_0_n13, npu_inst_pe_1_0_0_n12,
         npu_inst_pe_1_0_0_n11, npu_inst_pe_1_0_0_n10, npu_inst_pe_1_0_0_n9,
         npu_inst_pe_1_0_0_n8, npu_inst_pe_1_0_0_n7, npu_inst_pe_1_0_0_n6,
         npu_inst_pe_1_0_0_n5, npu_inst_pe_1_0_0_n4, npu_inst_pe_1_0_0_n3,
         npu_inst_pe_1_0_0_n2, npu_inst_pe_1_0_0_n1,
         npu_inst_pe_1_0_0_sub_77_carry_7_, npu_inst_pe_1_0_0_sub_77_carry_6_,
         npu_inst_pe_1_0_0_sub_77_carry_5_, npu_inst_pe_1_0_0_sub_77_carry_4_,
         npu_inst_pe_1_0_0_sub_77_carry_3_, npu_inst_pe_1_0_0_sub_77_carry_2_,
         npu_inst_pe_1_0_0_sub_77_carry_1_, npu_inst_pe_1_0_0_add_79_carry_7_,
         npu_inst_pe_1_0_0_add_79_carry_6_, npu_inst_pe_1_0_0_add_79_carry_5_,
         npu_inst_pe_1_0_0_add_79_carry_4_, npu_inst_pe_1_0_0_add_79_carry_3_,
         npu_inst_pe_1_0_0_add_79_carry_2_, npu_inst_pe_1_0_0_add_79_carry_1_,
         npu_inst_pe_1_0_0_n97, npu_inst_pe_1_0_0_n96, npu_inst_pe_1_0_0_n95,
         npu_inst_pe_1_0_0_n94, npu_inst_pe_1_0_0_n93, npu_inst_pe_1_0_0_n92,
         npu_inst_pe_1_0_0_n91, npu_inst_pe_1_0_0_n90, npu_inst_pe_1_0_0_n89,
         npu_inst_pe_1_0_0_n88, npu_inst_pe_1_0_0_n87, npu_inst_pe_1_0_0_n86,
         npu_inst_pe_1_0_0_n85, npu_inst_pe_1_0_0_n84, npu_inst_pe_1_0_0_n83,
         npu_inst_pe_1_0_0_n82, npu_inst_pe_1_0_0_n81, npu_inst_pe_1_0_0_n80,
         npu_inst_pe_1_0_0_n79, npu_inst_pe_1_0_0_n78, npu_inst_pe_1_0_0_n77,
         npu_inst_pe_1_0_0_n76, npu_inst_pe_1_0_0_n75, npu_inst_pe_1_0_0_n74,
         npu_inst_pe_1_0_0_n73, npu_inst_pe_1_0_0_n72, npu_inst_pe_1_0_0_n71,
         npu_inst_pe_1_0_0_n70, npu_inst_pe_1_0_0_n69, npu_inst_pe_1_0_0_n68,
         npu_inst_pe_1_0_0_n67, npu_inst_pe_1_0_0_n66, npu_inst_pe_1_0_0_n65,
         npu_inst_pe_1_0_0_n64, npu_inst_pe_1_0_0_n63, npu_inst_pe_1_0_0_n62,
         npu_inst_pe_1_0_0_n61, npu_inst_pe_1_0_0_n60, npu_inst_pe_1_0_0_n59,
         npu_inst_pe_1_0_0_n58, npu_inst_pe_1_0_0_n57, npu_inst_pe_1_0_0_n56,
         npu_inst_pe_1_0_0_n55, npu_inst_pe_1_0_0_n54, npu_inst_pe_1_0_0_n53,
         npu_inst_pe_1_0_0_n52, npu_inst_pe_1_0_0_n51, npu_inst_pe_1_0_0_n50,
         npu_inst_pe_1_0_0_n49, npu_inst_pe_1_0_0_n48, npu_inst_pe_1_0_0_n47,
         npu_inst_pe_1_0_0_n46, npu_inst_pe_1_0_0_n45, npu_inst_pe_1_0_0_n44,
         npu_inst_pe_1_0_0_n43, npu_inst_pe_1_0_0_n42, npu_inst_pe_1_0_0_n41,
         npu_inst_pe_1_0_0_n40, npu_inst_pe_1_0_0_n39, npu_inst_pe_1_0_0_n38,
         npu_inst_pe_1_0_0_n37, npu_inst_pe_1_0_0_n27, npu_inst_pe_1_0_0_n26,
         npu_inst_pe_1_0_0_net4299, npu_inst_pe_1_0_0_net4293,
         npu_inst_pe_1_0_0_N94, npu_inst_pe_1_0_0_N93, npu_inst_pe_1_0_0_N84,
         npu_inst_pe_1_0_0_N80, npu_inst_pe_1_0_0_N79, npu_inst_pe_1_0_0_N78,
         npu_inst_pe_1_0_0_N77, npu_inst_pe_1_0_0_N76, npu_inst_pe_1_0_0_N75,
         npu_inst_pe_1_0_0_N74, npu_inst_pe_1_0_0_N73, npu_inst_pe_1_0_0_N72,
         npu_inst_pe_1_0_0_N71, npu_inst_pe_1_0_0_N70, npu_inst_pe_1_0_0_N69,
         npu_inst_pe_1_0_0_N68, npu_inst_pe_1_0_0_N67, npu_inst_pe_1_0_0_N66,
         npu_inst_pe_1_0_0_N65, npu_inst_pe_1_0_0_int_q_acc_0_,
         npu_inst_pe_1_0_0_int_q_acc_1_, npu_inst_pe_1_0_0_int_q_acc_2_,
         npu_inst_pe_1_0_0_int_q_acc_3_, npu_inst_pe_1_0_0_int_q_acc_4_,
         npu_inst_pe_1_0_0_int_q_acc_5_, npu_inst_pe_1_0_0_int_q_acc_6_,
         npu_inst_pe_1_0_0_int_q_acc_7_, npu_inst_pe_1_0_0_int_data_0_,
         npu_inst_pe_1_0_0_int_data_1_, npu_inst_pe_1_0_0_int_q_weight_0_,
         npu_inst_pe_1_0_0_int_q_weight_1_,
         npu_inst_pe_1_0_0_int_q_reg_v_5__0_,
         npu_inst_pe_1_0_0_int_q_reg_v_5__1_,
         npu_inst_pe_1_0_0_int_q_reg_v_4__0_,
         npu_inst_pe_1_0_0_int_q_reg_v_4__1_,
         npu_inst_pe_1_0_0_int_q_reg_v_3__0_,
         npu_inst_pe_1_0_0_int_q_reg_v_3__1_,
         npu_inst_pe_1_0_0_int_q_reg_v_2__0_,
         npu_inst_pe_1_0_0_int_q_reg_v_2__1_,
         npu_inst_pe_1_0_0_int_q_reg_v_1__0_,
         npu_inst_pe_1_0_0_int_q_reg_v_1__1_,
         npu_inst_pe_1_0_0_int_q_reg_v_0__0_,
         npu_inst_pe_1_0_0_int_q_reg_v_0__1_,
         npu_inst_pe_1_0_0_int_q_reg_h_5__0_,
         npu_inst_pe_1_0_0_int_q_reg_h_5__1_,
         npu_inst_pe_1_0_0_int_q_reg_h_4__0_,
         npu_inst_pe_1_0_0_int_q_reg_h_4__1_,
         npu_inst_pe_1_0_0_int_q_reg_h_3__0_,
         npu_inst_pe_1_0_0_int_q_reg_h_3__1_,
         npu_inst_pe_1_0_0_int_q_reg_h_2__0_,
         npu_inst_pe_1_0_0_int_q_reg_h_2__1_,
         npu_inst_pe_1_0_0_int_q_reg_h_1__0_,
         npu_inst_pe_1_0_0_int_q_reg_h_1__1_,
         npu_inst_pe_1_0_0_int_q_reg_h_0__0_,
         npu_inst_pe_1_0_0_int_q_reg_h_0__1_, npu_inst_pe_1_0_0_o_data_v_0_,
         npu_inst_pe_1_0_0_o_data_v_1_, npu_inst_pe_1_0_0_o_data_h_0_,
         npu_inst_pe_1_0_0_o_data_h_1_, npu_inst_pe_1_0_1_n117,
         npu_inst_pe_1_0_1_n116, npu_inst_pe_1_0_1_n115,
         npu_inst_pe_1_0_1_n114, npu_inst_pe_1_0_1_n113,
         npu_inst_pe_1_0_1_n112, npu_inst_pe_1_0_1_n111,
         npu_inst_pe_1_0_1_n110, npu_inst_pe_1_0_1_n109,
         npu_inst_pe_1_0_1_n108, npu_inst_pe_1_0_1_n107,
         npu_inst_pe_1_0_1_n106, npu_inst_pe_1_0_1_n105,
         npu_inst_pe_1_0_1_n104, npu_inst_pe_1_0_1_n103,
         npu_inst_pe_1_0_1_n102, npu_inst_pe_1_0_1_n101,
         npu_inst_pe_1_0_1_n100, npu_inst_pe_1_0_1_n99, npu_inst_pe_1_0_1_n98,
         npu_inst_pe_1_0_1_n36, npu_inst_pe_1_0_1_n35, npu_inst_pe_1_0_1_n34,
         npu_inst_pe_1_0_1_n33, npu_inst_pe_1_0_1_n32, npu_inst_pe_1_0_1_n31,
         npu_inst_pe_1_0_1_n30, npu_inst_pe_1_0_1_n29, npu_inst_pe_1_0_1_n28,
         npu_inst_pe_1_0_1_n25, npu_inst_pe_1_0_1_n24, npu_inst_pe_1_0_1_n23,
         npu_inst_pe_1_0_1_n22, npu_inst_pe_1_0_1_n21, npu_inst_pe_1_0_1_n20,
         npu_inst_pe_1_0_1_n19, npu_inst_pe_1_0_1_n18, npu_inst_pe_1_0_1_n17,
         npu_inst_pe_1_0_1_n16, npu_inst_pe_1_0_1_n15, npu_inst_pe_1_0_1_n14,
         npu_inst_pe_1_0_1_n13, npu_inst_pe_1_0_1_n12, npu_inst_pe_1_0_1_n11,
         npu_inst_pe_1_0_1_n10, npu_inst_pe_1_0_1_n9, npu_inst_pe_1_0_1_n8,
         npu_inst_pe_1_0_1_n7, npu_inst_pe_1_0_1_n6, npu_inst_pe_1_0_1_n5,
         npu_inst_pe_1_0_1_n4, npu_inst_pe_1_0_1_n3, npu_inst_pe_1_0_1_n2,
         npu_inst_pe_1_0_1_n1, npu_inst_pe_1_0_1_sub_77_carry_7_,
         npu_inst_pe_1_0_1_sub_77_carry_6_, npu_inst_pe_1_0_1_sub_77_carry_5_,
         npu_inst_pe_1_0_1_sub_77_carry_4_, npu_inst_pe_1_0_1_sub_77_carry_3_,
         npu_inst_pe_1_0_1_sub_77_carry_2_, npu_inst_pe_1_0_1_sub_77_carry_1_,
         npu_inst_pe_1_0_1_add_79_carry_7_, npu_inst_pe_1_0_1_add_79_carry_6_,
         npu_inst_pe_1_0_1_add_79_carry_5_, npu_inst_pe_1_0_1_add_79_carry_4_,
         npu_inst_pe_1_0_1_add_79_carry_3_, npu_inst_pe_1_0_1_add_79_carry_2_,
         npu_inst_pe_1_0_1_add_79_carry_1_, npu_inst_pe_1_0_1_n97,
         npu_inst_pe_1_0_1_n96, npu_inst_pe_1_0_1_n95, npu_inst_pe_1_0_1_n94,
         npu_inst_pe_1_0_1_n93, npu_inst_pe_1_0_1_n92, npu_inst_pe_1_0_1_n91,
         npu_inst_pe_1_0_1_n90, npu_inst_pe_1_0_1_n89, npu_inst_pe_1_0_1_n88,
         npu_inst_pe_1_0_1_n87, npu_inst_pe_1_0_1_n86, npu_inst_pe_1_0_1_n85,
         npu_inst_pe_1_0_1_n84, npu_inst_pe_1_0_1_n83, npu_inst_pe_1_0_1_n82,
         npu_inst_pe_1_0_1_n81, npu_inst_pe_1_0_1_n80, npu_inst_pe_1_0_1_n79,
         npu_inst_pe_1_0_1_n78, npu_inst_pe_1_0_1_n77, npu_inst_pe_1_0_1_n76,
         npu_inst_pe_1_0_1_n75, npu_inst_pe_1_0_1_n74, npu_inst_pe_1_0_1_n73,
         npu_inst_pe_1_0_1_n72, npu_inst_pe_1_0_1_n71, npu_inst_pe_1_0_1_n70,
         npu_inst_pe_1_0_1_n69, npu_inst_pe_1_0_1_n68, npu_inst_pe_1_0_1_n67,
         npu_inst_pe_1_0_1_n66, npu_inst_pe_1_0_1_n65, npu_inst_pe_1_0_1_n64,
         npu_inst_pe_1_0_1_n63, npu_inst_pe_1_0_1_n62, npu_inst_pe_1_0_1_n61,
         npu_inst_pe_1_0_1_n60, npu_inst_pe_1_0_1_n59, npu_inst_pe_1_0_1_n58,
         npu_inst_pe_1_0_1_n57, npu_inst_pe_1_0_1_n56, npu_inst_pe_1_0_1_n55,
         npu_inst_pe_1_0_1_n54, npu_inst_pe_1_0_1_n53, npu_inst_pe_1_0_1_n52,
         npu_inst_pe_1_0_1_n51, npu_inst_pe_1_0_1_n50, npu_inst_pe_1_0_1_n49,
         npu_inst_pe_1_0_1_n48, npu_inst_pe_1_0_1_n47, npu_inst_pe_1_0_1_n46,
         npu_inst_pe_1_0_1_n45, npu_inst_pe_1_0_1_n44, npu_inst_pe_1_0_1_n43,
         npu_inst_pe_1_0_1_n42, npu_inst_pe_1_0_1_n41, npu_inst_pe_1_0_1_n40,
         npu_inst_pe_1_0_1_n39, npu_inst_pe_1_0_1_n38, npu_inst_pe_1_0_1_n37,
         npu_inst_pe_1_0_1_n27, npu_inst_pe_1_0_1_n26,
         npu_inst_pe_1_0_1_net4276, npu_inst_pe_1_0_1_net4270,
         npu_inst_pe_1_0_1_N94, npu_inst_pe_1_0_1_N93, npu_inst_pe_1_0_1_N84,
         npu_inst_pe_1_0_1_N80, npu_inst_pe_1_0_1_N79, npu_inst_pe_1_0_1_N78,
         npu_inst_pe_1_0_1_N77, npu_inst_pe_1_0_1_N76, npu_inst_pe_1_0_1_N75,
         npu_inst_pe_1_0_1_N74, npu_inst_pe_1_0_1_N73, npu_inst_pe_1_0_1_N72,
         npu_inst_pe_1_0_1_N71, npu_inst_pe_1_0_1_N70, npu_inst_pe_1_0_1_N69,
         npu_inst_pe_1_0_1_N68, npu_inst_pe_1_0_1_N67, npu_inst_pe_1_0_1_N66,
         npu_inst_pe_1_0_1_N65, npu_inst_pe_1_0_1_int_q_acc_0_,
         npu_inst_pe_1_0_1_int_q_acc_1_, npu_inst_pe_1_0_1_int_q_acc_2_,
         npu_inst_pe_1_0_1_int_q_acc_3_, npu_inst_pe_1_0_1_int_q_acc_4_,
         npu_inst_pe_1_0_1_int_q_acc_5_, npu_inst_pe_1_0_1_int_q_acc_6_,
         npu_inst_pe_1_0_1_int_q_acc_7_, npu_inst_pe_1_0_1_int_data_0_,
         npu_inst_pe_1_0_1_int_data_1_, npu_inst_pe_1_0_1_int_q_weight_0_,
         npu_inst_pe_1_0_1_int_q_weight_1_,
         npu_inst_pe_1_0_1_int_q_reg_v_5__0_,
         npu_inst_pe_1_0_1_int_q_reg_v_5__1_,
         npu_inst_pe_1_0_1_int_q_reg_v_4__0_,
         npu_inst_pe_1_0_1_int_q_reg_v_4__1_,
         npu_inst_pe_1_0_1_int_q_reg_v_3__0_,
         npu_inst_pe_1_0_1_int_q_reg_v_3__1_,
         npu_inst_pe_1_0_1_int_q_reg_v_2__0_,
         npu_inst_pe_1_0_1_int_q_reg_v_2__1_,
         npu_inst_pe_1_0_1_int_q_reg_v_1__0_,
         npu_inst_pe_1_0_1_int_q_reg_v_1__1_,
         npu_inst_pe_1_0_1_int_q_reg_v_0__0_,
         npu_inst_pe_1_0_1_int_q_reg_v_0__1_,
         npu_inst_pe_1_0_1_int_q_reg_h_5__0_,
         npu_inst_pe_1_0_1_int_q_reg_h_5__1_,
         npu_inst_pe_1_0_1_int_q_reg_h_4__0_,
         npu_inst_pe_1_0_1_int_q_reg_h_4__1_,
         npu_inst_pe_1_0_1_int_q_reg_h_3__0_,
         npu_inst_pe_1_0_1_int_q_reg_h_3__1_,
         npu_inst_pe_1_0_1_int_q_reg_h_2__0_,
         npu_inst_pe_1_0_1_int_q_reg_h_2__1_,
         npu_inst_pe_1_0_1_int_q_reg_h_1__0_,
         npu_inst_pe_1_0_1_int_q_reg_h_1__1_,
         npu_inst_pe_1_0_1_int_q_reg_h_0__0_,
         npu_inst_pe_1_0_1_int_q_reg_h_0__1_, npu_inst_pe_1_0_1_o_data_v_0_,
         npu_inst_pe_1_0_1_o_data_v_1_, npu_inst_pe_1_0_2_n118,
         npu_inst_pe_1_0_2_n117, npu_inst_pe_1_0_2_n116,
         npu_inst_pe_1_0_2_n115, npu_inst_pe_1_0_2_n114,
         npu_inst_pe_1_0_2_n113, npu_inst_pe_1_0_2_n112,
         npu_inst_pe_1_0_2_n111, npu_inst_pe_1_0_2_n110,
         npu_inst_pe_1_0_2_n109, npu_inst_pe_1_0_2_n108,
         npu_inst_pe_1_0_2_n107, npu_inst_pe_1_0_2_n106,
         npu_inst_pe_1_0_2_n105, npu_inst_pe_1_0_2_n104,
         npu_inst_pe_1_0_2_n103, npu_inst_pe_1_0_2_n102,
         npu_inst_pe_1_0_2_n101, npu_inst_pe_1_0_2_n100, npu_inst_pe_1_0_2_n99,
         npu_inst_pe_1_0_2_n98, npu_inst_pe_1_0_2_n36, npu_inst_pe_1_0_2_n35,
         npu_inst_pe_1_0_2_n34, npu_inst_pe_1_0_2_n33, npu_inst_pe_1_0_2_n32,
         npu_inst_pe_1_0_2_n31, npu_inst_pe_1_0_2_n30, npu_inst_pe_1_0_2_n29,
         npu_inst_pe_1_0_2_n28, npu_inst_pe_1_0_2_n25, npu_inst_pe_1_0_2_n24,
         npu_inst_pe_1_0_2_n23, npu_inst_pe_1_0_2_n22, npu_inst_pe_1_0_2_n21,
         npu_inst_pe_1_0_2_n20, npu_inst_pe_1_0_2_n19, npu_inst_pe_1_0_2_n18,
         npu_inst_pe_1_0_2_n17, npu_inst_pe_1_0_2_n16, npu_inst_pe_1_0_2_n15,
         npu_inst_pe_1_0_2_n14, npu_inst_pe_1_0_2_n13, npu_inst_pe_1_0_2_n12,
         npu_inst_pe_1_0_2_n11, npu_inst_pe_1_0_2_n10, npu_inst_pe_1_0_2_n9,
         npu_inst_pe_1_0_2_n8, npu_inst_pe_1_0_2_n7, npu_inst_pe_1_0_2_n6,
         npu_inst_pe_1_0_2_n5, npu_inst_pe_1_0_2_n4, npu_inst_pe_1_0_2_n3,
         npu_inst_pe_1_0_2_n2, npu_inst_pe_1_0_2_n1,
         npu_inst_pe_1_0_2_sub_77_carry_7_, npu_inst_pe_1_0_2_sub_77_carry_6_,
         npu_inst_pe_1_0_2_sub_77_carry_5_, npu_inst_pe_1_0_2_sub_77_carry_4_,
         npu_inst_pe_1_0_2_sub_77_carry_3_, npu_inst_pe_1_0_2_sub_77_carry_2_,
         npu_inst_pe_1_0_2_sub_77_carry_1_, npu_inst_pe_1_0_2_add_79_carry_7_,
         npu_inst_pe_1_0_2_add_79_carry_6_, npu_inst_pe_1_0_2_add_79_carry_5_,
         npu_inst_pe_1_0_2_add_79_carry_4_, npu_inst_pe_1_0_2_add_79_carry_3_,
         npu_inst_pe_1_0_2_add_79_carry_2_, npu_inst_pe_1_0_2_add_79_carry_1_,
         npu_inst_pe_1_0_2_n97, npu_inst_pe_1_0_2_n96, npu_inst_pe_1_0_2_n95,
         npu_inst_pe_1_0_2_n94, npu_inst_pe_1_0_2_n93, npu_inst_pe_1_0_2_n92,
         npu_inst_pe_1_0_2_n91, npu_inst_pe_1_0_2_n90, npu_inst_pe_1_0_2_n89,
         npu_inst_pe_1_0_2_n88, npu_inst_pe_1_0_2_n87, npu_inst_pe_1_0_2_n86,
         npu_inst_pe_1_0_2_n85, npu_inst_pe_1_0_2_n84, npu_inst_pe_1_0_2_n83,
         npu_inst_pe_1_0_2_n82, npu_inst_pe_1_0_2_n81, npu_inst_pe_1_0_2_n80,
         npu_inst_pe_1_0_2_n79, npu_inst_pe_1_0_2_n78, npu_inst_pe_1_0_2_n77,
         npu_inst_pe_1_0_2_n76, npu_inst_pe_1_0_2_n75, npu_inst_pe_1_0_2_n74,
         npu_inst_pe_1_0_2_n73, npu_inst_pe_1_0_2_n72, npu_inst_pe_1_0_2_n71,
         npu_inst_pe_1_0_2_n70, npu_inst_pe_1_0_2_n69, npu_inst_pe_1_0_2_n68,
         npu_inst_pe_1_0_2_n67, npu_inst_pe_1_0_2_n66, npu_inst_pe_1_0_2_n65,
         npu_inst_pe_1_0_2_n64, npu_inst_pe_1_0_2_n63, npu_inst_pe_1_0_2_n62,
         npu_inst_pe_1_0_2_n61, npu_inst_pe_1_0_2_n60, npu_inst_pe_1_0_2_n59,
         npu_inst_pe_1_0_2_n58, npu_inst_pe_1_0_2_n57, npu_inst_pe_1_0_2_n56,
         npu_inst_pe_1_0_2_n55, npu_inst_pe_1_0_2_n54, npu_inst_pe_1_0_2_n53,
         npu_inst_pe_1_0_2_n52, npu_inst_pe_1_0_2_n51, npu_inst_pe_1_0_2_n50,
         npu_inst_pe_1_0_2_n49, npu_inst_pe_1_0_2_n48, npu_inst_pe_1_0_2_n47,
         npu_inst_pe_1_0_2_n46, npu_inst_pe_1_0_2_n45, npu_inst_pe_1_0_2_n44,
         npu_inst_pe_1_0_2_n43, npu_inst_pe_1_0_2_n42, npu_inst_pe_1_0_2_n41,
         npu_inst_pe_1_0_2_n40, npu_inst_pe_1_0_2_n39, npu_inst_pe_1_0_2_n38,
         npu_inst_pe_1_0_2_n37, npu_inst_pe_1_0_2_n27, npu_inst_pe_1_0_2_n26,
         npu_inst_pe_1_0_2_net4253, npu_inst_pe_1_0_2_net4247,
         npu_inst_pe_1_0_2_N94, npu_inst_pe_1_0_2_N93, npu_inst_pe_1_0_2_N84,
         npu_inst_pe_1_0_2_N80, npu_inst_pe_1_0_2_N79, npu_inst_pe_1_0_2_N78,
         npu_inst_pe_1_0_2_N77, npu_inst_pe_1_0_2_N76, npu_inst_pe_1_0_2_N75,
         npu_inst_pe_1_0_2_N74, npu_inst_pe_1_0_2_N73, npu_inst_pe_1_0_2_N72,
         npu_inst_pe_1_0_2_N71, npu_inst_pe_1_0_2_N70, npu_inst_pe_1_0_2_N69,
         npu_inst_pe_1_0_2_N68, npu_inst_pe_1_0_2_N67, npu_inst_pe_1_0_2_N66,
         npu_inst_pe_1_0_2_N65, npu_inst_pe_1_0_2_int_q_acc_0_,
         npu_inst_pe_1_0_2_int_q_acc_1_, npu_inst_pe_1_0_2_int_q_acc_2_,
         npu_inst_pe_1_0_2_int_q_acc_3_, npu_inst_pe_1_0_2_int_q_acc_4_,
         npu_inst_pe_1_0_2_int_q_acc_5_, npu_inst_pe_1_0_2_int_q_acc_6_,
         npu_inst_pe_1_0_2_int_q_acc_7_, npu_inst_pe_1_0_2_int_data_0_,
         npu_inst_pe_1_0_2_int_data_1_, npu_inst_pe_1_0_2_int_q_weight_0_,
         npu_inst_pe_1_0_2_int_q_weight_1_,
         npu_inst_pe_1_0_2_int_q_reg_v_5__0_,
         npu_inst_pe_1_0_2_int_q_reg_v_5__1_,
         npu_inst_pe_1_0_2_int_q_reg_v_4__0_,
         npu_inst_pe_1_0_2_int_q_reg_v_4__1_,
         npu_inst_pe_1_0_2_int_q_reg_v_3__0_,
         npu_inst_pe_1_0_2_int_q_reg_v_3__1_,
         npu_inst_pe_1_0_2_int_q_reg_v_2__0_,
         npu_inst_pe_1_0_2_int_q_reg_v_2__1_,
         npu_inst_pe_1_0_2_int_q_reg_v_1__0_,
         npu_inst_pe_1_0_2_int_q_reg_v_1__1_,
         npu_inst_pe_1_0_2_int_q_reg_v_0__0_,
         npu_inst_pe_1_0_2_int_q_reg_v_0__1_,
         npu_inst_pe_1_0_2_int_q_reg_h_5__0_,
         npu_inst_pe_1_0_2_int_q_reg_h_5__1_,
         npu_inst_pe_1_0_2_int_q_reg_h_4__0_,
         npu_inst_pe_1_0_2_int_q_reg_h_4__1_,
         npu_inst_pe_1_0_2_int_q_reg_h_3__0_,
         npu_inst_pe_1_0_2_int_q_reg_h_3__1_,
         npu_inst_pe_1_0_2_int_q_reg_h_2__0_,
         npu_inst_pe_1_0_2_int_q_reg_h_2__1_,
         npu_inst_pe_1_0_2_int_q_reg_h_1__0_,
         npu_inst_pe_1_0_2_int_q_reg_h_1__1_,
         npu_inst_pe_1_0_2_int_q_reg_h_0__0_,
         npu_inst_pe_1_0_2_int_q_reg_h_0__1_, npu_inst_pe_1_0_2_o_data_v_0_,
         npu_inst_pe_1_0_2_o_data_v_1_, npu_inst_pe_1_0_3_n119,
         npu_inst_pe_1_0_3_n118, npu_inst_pe_1_0_3_n117,
         npu_inst_pe_1_0_3_n116, npu_inst_pe_1_0_3_n115,
         npu_inst_pe_1_0_3_n114, npu_inst_pe_1_0_3_n113,
         npu_inst_pe_1_0_3_n112, npu_inst_pe_1_0_3_n111,
         npu_inst_pe_1_0_3_n110, npu_inst_pe_1_0_3_n109,
         npu_inst_pe_1_0_3_n108, npu_inst_pe_1_0_3_n107,
         npu_inst_pe_1_0_3_n106, npu_inst_pe_1_0_3_n105,
         npu_inst_pe_1_0_3_n104, npu_inst_pe_1_0_3_n103,
         npu_inst_pe_1_0_3_n102, npu_inst_pe_1_0_3_n101,
         npu_inst_pe_1_0_3_n100, npu_inst_pe_1_0_3_n99, npu_inst_pe_1_0_3_n98,
         npu_inst_pe_1_0_3_n36, npu_inst_pe_1_0_3_n35, npu_inst_pe_1_0_3_n34,
         npu_inst_pe_1_0_3_n33, npu_inst_pe_1_0_3_n32, npu_inst_pe_1_0_3_n31,
         npu_inst_pe_1_0_3_n30, npu_inst_pe_1_0_3_n29, npu_inst_pe_1_0_3_n28,
         npu_inst_pe_1_0_3_n25, npu_inst_pe_1_0_3_n24, npu_inst_pe_1_0_3_n23,
         npu_inst_pe_1_0_3_n22, npu_inst_pe_1_0_3_n21, npu_inst_pe_1_0_3_n20,
         npu_inst_pe_1_0_3_n19, npu_inst_pe_1_0_3_n18, npu_inst_pe_1_0_3_n17,
         npu_inst_pe_1_0_3_n16, npu_inst_pe_1_0_3_n15, npu_inst_pe_1_0_3_n14,
         npu_inst_pe_1_0_3_n13, npu_inst_pe_1_0_3_n12, npu_inst_pe_1_0_3_n11,
         npu_inst_pe_1_0_3_n10, npu_inst_pe_1_0_3_n9, npu_inst_pe_1_0_3_n8,
         npu_inst_pe_1_0_3_n7, npu_inst_pe_1_0_3_n6, npu_inst_pe_1_0_3_n5,
         npu_inst_pe_1_0_3_n4, npu_inst_pe_1_0_3_n3, npu_inst_pe_1_0_3_n2,
         npu_inst_pe_1_0_3_n1, npu_inst_pe_1_0_3_sub_77_carry_7_,
         npu_inst_pe_1_0_3_sub_77_carry_6_, npu_inst_pe_1_0_3_sub_77_carry_5_,
         npu_inst_pe_1_0_3_sub_77_carry_4_, npu_inst_pe_1_0_3_sub_77_carry_3_,
         npu_inst_pe_1_0_3_sub_77_carry_2_, npu_inst_pe_1_0_3_sub_77_carry_1_,
         npu_inst_pe_1_0_3_add_79_carry_7_, npu_inst_pe_1_0_3_add_79_carry_6_,
         npu_inst_pe_1_0_3_add_79_carry_5_, npu_inst_pe_1_0_3_add_79_carry_4_,
         npu_inst_pe_1_0_3_add_79_carry_3_, npu_inst_pe_1_0_3_add_79_carry_2_,
         npu_inst_pe_1_0_3_add_79_carry_1_, npu_inst_pe_1_0_3_n97,
         npu_inst_pe_1_0_3_n96, npu_inst_pe_1_0_3_n95, npu_inst_pe_1_0_3_n94,
         npu_inst_pe_1_0_3_n93, npu_inst_pe_1_0_3_n92, npu_inst_pe_1_0_3_n91,
         npu_inst_pe_1_0_3_n90, npu_inst_pe_1_0_3_n89, npu_inst_pe_1_0_3_n88,
         npu_inst_pe_1_0_3_n87, npu_inst_pe_1_0_3_n86, npu_inst_pe_1_0_3_n85,
         npu_inst_pe_1_0_3_n84, npu_inst_pe_1_0_3_n83, npu_inst_pe_1_0_3_n82,
         npu_inst_pe_1_0_3_n81, npu_inst_pe_1_0_3_n80, npu_inst_pe_1_0_3_n79,
         npu_inst_pe_1_0_3_n78, npu_inst_pe_1_0_3_n77, npu_inst_pe_1_0_3_n76,
         npu_inst_pe_1_0_3_n75, npu_inst_pe_1_0_3_n74, npu_inst_pe_1_0_3_n73,
         npu_inst_pe_1_0_3_n72, npu_inst_pe_1_0_3_n71, npu_inst_pe_1_0_3_n70,
         npu_inst_pe_1_0_3_n69, npu_inst_pe_1_0_3_n68, npu_inst_pe_1_0_3_n67,
         npu_inst_pe_1_0_3_n66, npu_inst_pe_1_0_3_n65, npu_inst_pe_1_0_3_n64,
         npu_inst_pe_1_0_3_n63, npu_inst_pe_1_0_3_n62, npu_inst_pe_1_0_3_n61,
         npu_inst_pe_1_0_3_n60, npu_inst_pe_1_0_3_n59, npu_inst_pe_1_0_3_n58,
         npu_inst_pe_1_0_3_n57, npu_inst_pe_1_0_3_n56, npu_inst_pe_1_0_3_n55,
         npu_inst_pe_1_0_3_n54, npu_inst_pe_1_0_3_n53, npu_inst_pe_1_0_3_n52,
         npu_inst_pe_1_0_3_n51, npu_inst_pe_1_0_3_n50, npu_inst_pe_1_0_3_n49,
         npu_inst_pe_1_0_3_n48, npu_inst_pe_1_0_3_n47, npu_inst_pe_1_0_3_n46,
         npu_inst_pe_1_0_3_n45, npu_inst_pe_1_0_3_n44, npu_inst_pe_1_0_3_n43,
         npu_inst_pe_1_0_3_n42, npu_inst_pe_1_0_3_n41, npu_inst_pe_1_0_3_n40,
         npu_inst_pe_1_0_3_n39, npu_inst_pe_1_0_3_n38, npu_inst_pe_1_0_3_n37,
         npu_inst_pe_1_0_3_n27, npu_inst_pe_1_0_3_n26,
         npu_inst_pe_1_0_3_net4230, npu_inst_pe_1_0_3_net4224,
         npu_inst_pe_1_0_3_N94, npu_inst_pe_1_0_3_N93, npu_inst_pe_1_0_3_N84,
         npu_inst_pe_1_0_3_N80, npu_inst_pe_1_0_3_N79, npu_inst_pe_1_0_3_N78,
         npu_inst_pe_1_0_3_N77, npu_inst_pe_1_0_3_N76, npu_inst_pe_1_0_3_N75,
         npu_inst_pe_1_0_3_N74, npu_inst_pe_1_0_3_N73, npu_inst_pe_1_0_3_N72,
         npu_inst_pe_1_0_3_N71, npu_inst_pe_1_0_3_N70, npu_inst_pe_1_0_3_N69,
         npu_inst_pe_1_0_3_N68, npu_inst_pe_1_0_3_N67, npu_inst_pe_1_0_3_N66,
         npu_inst_pe_1_0_3_N65, npu_inst_pe_1_0_3_int_q_acc_0_,
         npu_inst_pe_1_0_3_int_q_acc_1_, npu_inst_pe_1_0_3_int_q_acc_2_,
         npu_inst_pe_1_0_3_int_q_acc_3_, npu_inst_pe_1_0_3_int_q_acc_4_,
         npu_inst_pe_1_0_3_int_q_acc_5_, npu_inst_pe_1_0_3_int_q_acc_6_,
         npu_inst_pe_1_0_3_int_q_acc_7_, npu_inst_pe_1_0_3_int_data_0_,
         npu_inst_pe_1_0_3_int_data_1_, npu_inst_pe_1_0_3_int_q_weight_0_,
         npu_inst_pe_1_0_3_int_q_weight_1_,
         npu_inst_pe_1_0_3_int_q_reg_v_5__0_,
         npu_inst_pe_1_0_3_int_q_reg_v_5__1_,
         npu_inst_pe_1_0_3_int_q_reg_v_4__0_,
         npu_inst_pe_1_0_3_int_q_reg_v_4__1_,
         npu_inst_pe_1_0_3_int_q_reg_v_3__0_,
         npu_inst_pe_1_0_3_int_q_reg_v_3__1_,
         npu_inst_pe_1_0_3_int_q_reg_v_2__0_,
         npu_inst_pe_1_0_3_int_q_reg_v_2__1_,
         npu_inst_pe_1_0_3_int_q_reg_v_1__0_,
         npu_inst_pe_1_0_3_int_q_reg_v_1__1_,
         npu_inst_pe_1_0_3_int_q_reg_v_0__0_,
         npu_inst_pe_1_0_3_int_q_reg_v_0__1_,
         npu_inst_pe_1_0_3_int_q_reg_h_5__0_,
         npu_inst_pe_1_0_3_int_q_reg_h_5__1_,
         npu_inst_pe_1_0_3_int_q_reg_h_4__0_,
         npu_inst_pe_1_0_3_int_q_reg_h_4__1_,
         npu_inst_pe_1_0_3_int_q_reg_h_3__0_,
         npu_inst_pe_1_0_3_int_q_reg_h_3__1_,
         npu_inst_pe_1_0_3_int_q_reg_h_2__0_,
         npu_inst_pe_1_0_3_int_q_reg_h_2__1_,
         npu_inst_pe_1_0_3_int_q_reg_h_1__0_,
         npu_inst_pe_1_0_3_int_q_reg_h_1__1_,
         npu_inst_pe_1_0_3_int_q_reg_h_0__0_,
         npu_inst_pe_1_0_3_int_q_reg_h_0__1_, npu_inst_pe_1_0_3_o_data_v_0_,
         npu_inst_pe_1_0_3_o_data_v_1_, npu_inst_pe_1_0_4_n118,
         npu_inst_pe_1_0_4_n117, npu_inst_pe_1_0_4_n116,
         npu_inst_pe_1_0_4_n115, npu_inst_pe_1_0_4_n114,
         npu_inst_pe_1_0_4_n113, npu_inst_pe_1_0_4_n112,
         npu_inst_pe_1_0_4_n111, npu_inst_pe_1_0_4_n110,
         npu_inst_pe_1_0_4_n109, npu_inst_pe_1_0_4_n108,
         npu_inst_pe_1_0_4_n107, npu_inst_pe_1_0_4_n106,
         npu_inst_pe_1_0_4_n105, npu_inst_pe_1_0_4_n104,
         npu_inst_pe_1_0_4_n103, npu_inst_pe_1_0_4_n102,
         npu_inst_pe_1_0_4_n101, npu_inst_pe_1_0_4_n100, npu_inst_pe_1_0_4_n99,
         npu_inst_pe_1_0_4_n98, npu_inst_pe_1_0_4_n36, npu_inst_pe_1_0_4_n35,
         npu_inst_pe_1_0_4_n34, npu_inst_pe_1_0_4_n33, npu_inst_pe_1_0_4_n32,
         npu_inst_pe_1_0_4_n31, npu_inst_pe_1_0_4_n30, npu_inst_pe_1_0_4_n29,
         npu_inst_pe_1_0_4_n28, npu_inst_pe_1_0_4_n25, npu_inst_pe_1_0_4_n24,
         npu_inst_pe_1_0_4_n23, npu_inst_pe_1_0_4_n22, npu_inst_pe_1_0_4_n21,
         npu_inst_pe_1_0_4_n20, npu_inst_pe_1_0_4_n19, npu_inst_pe_1_0_4_n18,
         npu_inst_pe_1_0_4_n17, npu_inst_pe_1_0_4_n16, npu_inst_pe_1_0_4_n15,
         npu_inst_pe_1_0_4_n14, npu_inst_pe_1_0_4_n13, npu_inst_pe_1_0_4_n12,
         npu_inst_pe_1_0_4_n11, npu_inst_pe_1_0_4_n10, npu_inst_pe_1_0_4_n9,
         npu_inst_pe_1_0_4_n8, npu_inst_pe_1_0_4_n7, npu_inst_pe_1_0_4_n6,
         npu_inst_pe_1_0_4_n5, npu_inst_pe_1_0_4_n4, npu_inst_pe_1_0_4_n3,
         npu_inst_pe_1_0_4_n2, npu_inst_pe_1_0_4_n1,
         npu_inst_pe_1_0_4_sub_77_carry_7_, npu_inst_pe_1_0_4_sub_77_carry_6_,
         npu_inst_pe_1_0_4_sub_77_carry_5_, npu_inst_pe_1_0_4_sub_77_carry_4_,
         npu_inst_pe_1_0_4_sub_77_carry_3_, npu_inst_pe_1_0_4_sub_77_carry_2_,
         npu_inst_pe_1_0_4_sub_77_carry_1_, npu_inst_pe_1_0_4_add_79_carry_7_,
         npu_inst_pe_1_0_4_add_79_carry_6_, npu_inst_pe_1_0_4_add_79_carry_5_,
         npu_inst_pe_1_0_4_add_79_carry_4_, npu_inst_pe_1_0_4_add_79_carry_3_,
         npu_inst_pe_1_0_4_add_79_carry_2_, npu_inst_pe_1_0_4_add_79_carry_1_,
         npu_inst_pe_1_0_4_n97, npu_inst_pe_1_0_4_n96, npu_inst_pe_1_0_4_n95,
         npu_inst_pe_1_0_4_n94, npu_inst_pe_1_0_4_n93, npu_inst_pe_1_0_4_n92,
         npu_inst_pe_1_0_4_n91, npu_inst_pe_1_0_4_n90, npu_inst_pe_1_0_4_n89,
         npu_inst_pe_1_0_4_n88, npu_inst_pe_1_0_4_n87, npu_inst_pe_1_0_4_n86,
         npu_inst_pe_1_0_4_n85, npu_inst_pe_1_0_4_n84, npu_inst_pe_1_0_4_n83,
         npu_inst_pe_1_0_4_n82, npu_inst_pe_1_0_4_n81, npu_inst_pe_1_0_4_n80,
         npu_inst_pe_1_0_4_n79, npu_inst_pe_1_0_4_n78, npu_inst_pe_1_0_4_n77,
         npu_inst_pe_1_0_4_n76, npu_inst_pe_1_0_4_n75, npu_inst_pe_1_0_4_n74,
         npu_inst_pe_1_0_4_n73, npu_inst_pe_1_0_4_n72, npu_inst_pe_1_0_4_n71,
         npu_inst_pe_1_0_4_n70, npu_inst_pe_1_0_4_n69, npu_inst_pe_1_0_4_n68,
         npu_inst_pe_1_0_4_n67, npu_inst_pe_1_0_4_n66, npu_inst_pe_1_0_4_n65,
         npu_inst_pe_1_0_4_n64, npu_inst_pe_1_0_4_n63, npu_inst_pe_1_0_4_n62,
         npu_inst_pe_1_0_4_n61, npu_inst_pe_1_0_4_n60, npu_inst_pe_1_0_4_n59,
         npu_inst_pe_1_0_4_n58, npu_inst_pe_1_0_4_n57, npu_inst_pe_1_0_4_n56,
         npu_inst_pe_1_0_4_n55, npu_inst_pe_1_0_4_n54, npu_inst_pe_1_0_4_n53,
         npu_inst_pe_1_0_4_n52, npu_inst_pe_1_0_4_n51, npu_inst_pe_1_0_4_n50,
         npu_inst_pe_1_0_4_n49, npu_inst_pe_1_0_4_n48, npu_inst_pe_1_0_4_n47,
         npu_inst_pe_1_0_4_n46, npu_inst_pe_1_0_4_n45, npu_inst_pe_1_0_4_n44,
         npu_inst_pe_1_0_4_n43, npu_inst_pe_1_0_4_n42, npu_inst_pe_1_0_4_n41,
         npu_inst_pe_1_0_4_n40, npu_inst_pe_1_0_4_n39, npu_inst_pe_1_0_4_n38,
         npu_inst_pe_1_0_4_n37, npu_inst_pe_1_0_4_n27, npu_inst_pe_1_0_4_n26,
         npu_inst_pe_1_0_4_net4207, npu_inst_pe_1_0_4_net4201,
         npu_inst_pe_1_0_4_N94, npu_inst_pe_1_0_4_N93, npu_inst_pe_1_0_4_N84,
         npu_inst_pe_1_0_4_N80, npu_inst_pe_1_0_4_N79, npu_inst_pe_1_0_4_N78,
         npu_inst_pe_1_0_4_N77, npu_inst_pe_1_0_4_N76, npu_inst_pe_1_0_4_N75,
         npu_inst_pe_1_0_4_N74, npu_inst_pe_1_0_4_N73, npu_inst_pe_1_0_4_N72,
         npu_inst_pe_1_0_4_N71, npu_inst_pe_1_0_4_N70, npu_inst_pe_1_0_4_N69,
         npu_inst_pe_1_0_4_N68, npu_inst_pe_1_0_4_N67, npu_inst_pe_1_0_4_N66,
         npu_inst_pe_1_0_4_N65, npu_inst_pe_1_0_4_int_q_acc_0_,
         npu_inst_pe_1_0_4_int_q_acc_1_, npu_inst_pe_1_0_4_int_q_acc_2_,
         npu_inst_pe_1_0_4_int_q_acc_3_, npu_inst_pe_1_0_4_int_q_acc_4_,
         npu_inst_pe_1_0_4_int_q_acc_5_, npu_inst_pe_1_0_4_int_q_acc_6_,
         npu_inst_pe_1_0_4_int_q_acc_7_, npu_inst_pe_1_0_4_int_data_0_,
         npu_inst_pe_1_0_4_int_data_1_, npu_inst_pe_1_0_4_int_q_weight_0_,
         npu_inst_pe_1_0_4_int_q_weight_1_,
         npu_inst_pe_1_0_4_int_q_reg_v_5__0_,
         npu_inst_pe_1_0_4_int_q_reg_v_5__1_,
         npu_inst_pe_1_0_4_int_q_reg_v_4__0_,
         npu_inst_pe_1_0_4_int_q_reg_v_4__1_,
         npu_inst_pe_1_0_4_int_q_reg_v_3__0_,
         npu_inst_pe_1_0_4_int_q_reg_v_3__1_,
         npu_inst_pe_1_0_4_int_q_reg_v_2__0_,
         npu_inst_pe_1_0_4_int_q_reg_v_2__1_,
         npu_inst_pe_1_0_4_int_q_reg_v_1__0_,
         npu_inst_pe_1_0_4_int_q_reg_v_1__1_,
         npu_inst_pe_1_0_4_int_q_reg_v_0__0_,
         npu_inst_pe_1_0_4_int_q_reg_v_0__1_,
         npu_inst_pe_1_0_4_int_q_reg_h_5__0_,
         npu_inst_pe_1_0_4_int_q_reg_h_5__1_,
         npu_inst_pe_1_0_4_int_q_reg_h_4__0_,
         npu_inst_pe_1_0_4_int_q_reg_h_4__1_,
         npu_inst_pe_1_0_4_int_q_reg_h_3__0_,
         npu_inst_pe_1_0_4_int_q_reg_h_3__1_,
         npu_inst_pe_1_0_4_int_q_reg_h_2__0_,
         npu_inst_pe_1_0_4_int_q_reg_h_2__1_,
         npu_inst_pe_1_0_4_int_q_reg_h_1__0_,
         npu_inst_pe_1_0_4_int_q_reg_h_1__1_,
         npu_inst_pe_1_0_4_int_q_reg_h_0__0_,
         npu_inst_pe_1_0_4_int_q_reg_h_0__1_, npu_inst_pe_1_0_4_o_data_v_0_,
         npu_inst_pe_1_0_4_o_data_v_1_, npu_inst_pe_1_0_5_n119,
         npu_inst_pe_1_0_5_n118, npu_inst_pe_1_0_5_n117,
         npu_inst_pe_1_0_5_n116, npu_inst_pe_1_0_5_n115,
         npu_inst_pe_1_0_5_n114, npu_inst_pe_1_0_5_n113,
         npu_inst_pe_1_0_5_n112, npu_inst_pe_1_0_5_n111,
         npu_inst_pe_1_0_5_n110, npu_inst_pe_1_0_5_n109,
         npu_inst_pe_1_0_5_n108, npu_inst_pe_1_0_5_n107,
         npu_inst_pe_1_0_5_n106, npu_inst_pe_1_0_5_n105,
         npu_inst_pe_1_0_5_n104, npu_inst_pe_1_0_5_n103,
         npu_inst_pe_1_0_5_n102, npu_inst_pe_1_0_5_n101,
         npu_inst_pe_1_0_5_n100, npu_inst_pe_1_0_5_n99, npu_inst_pe_1_0_5_n98,
         npu_inst_pe_1_0_5_n36, npu_inst_pe_1_0_5_n35, npu_inst_pe_1_0_5_n34,
         npu_inst_pe_1_0_5_n33, npu_inst_pe_1_0_5_n32, npu_inst_pe_1_0_5_n31,
         npu_inst_pe_1_0_5_n30, npu_inst_pe_1_0_5_n29, npu_inst_pe_1_0_5_n28,
         npu_inst_pe_1_0_5_n25, npu_inst_pe_1_0_5_n24, npu_inst_pe_1_0_5_n23,
         npu_inst_pe_1_0_5_n22, npu_inst_pe_1_0_5_n21, npu_inst_pe_1_0_5_n20,
         npu_inst_pe_1_0_5_n19, npu_inst_pe_1_0_5_n18, npu_inst_pe_1_0_5_n17,
         npu_inst_pe_1_0_5_n16, npu_inst_pe_1_0_5_n15, npu_inst_pe_1_0_5_n14,
         npu_inst_pe_1_0_5_n13, npu_inst_pe_1_0_5_n12, npu_inst_pe_1_0_5_n11,
         npu_inst_pe_1_0_5_n10, npu_inst_pe_1_0_5_n9, npu_inst_pe_1_0_5_n8,
         npu_inst_pe_1_0_5_n7, npu_inst_pe_1_0_5_n6, npu_inst_pe_1_0_5_n5,
         npu_inst_pe_1_0_5_n4, npu_inst_pe_1_0_5_n3, npu_inst_pe_1_0_5_n2,
         npu_inst_pe_1_0_5_n1, npu_inst_pe_1_0_5_sub_77_carry_7_,
         npu_inst_pe_1_0_5_sub_77_carry_6_, npu_inst_pe_1_0_5_sub_77_carry_5_,
         npu_inst_pe_1_0_5_sub_77_carry_4_, npu_inst_pe_1_0_5_sub_77_carry_3_,
         npu_inst_pe_1_0_5_sub_77_carry_2_, npu_inst_pe_1_0_5_sub_77_carry_1_,
         npu_inst_pe_1_0_5_add_79_carry_7_, npu_inst_pe_1_0_5_add_79_carry_6_,
         npu_inst_pe_1_0_5_add_79_carry_5_, npu_inst_pe_1_0_5_add_79_carry_4_,
         npu_inst_pe_1_0_5_add_79_carry_3_, npu_inst_pe_1_0_5_add_79_carry_2_,
         npu_inst_pe_1_0_5_add_79_carry_1_, npu_inst_pe_1_0_5_n97,
         npu_inst_pe_1_0_5_n96, npu_inst_pe_1_0_5_n95, npu_inst_pe_1_0_5_n94,
         npu_inst_pe_1_0_5_n93, npu_inst_pe_1_0_5_n92, npu_inst_pe_1_0_5_n91,
         npu_inst_pe_1_0_5_n90, npu_inst_pe_1_0_5_n89, npu_inst_pe_1_0_5_n88,
         npu_inst_pe_1_0_5_n87, npu_inst_pe_1_0_5_n86, npu_inst_pe_1_0_5_n85,
         npu_inst_pe_1_0_5_n84, npu_inst_pe_1_0_5_n83, npu_inst_pe_1_0_5_n82,
         npu_inst_pe_1_0_5_n81, npu_inst_pe_1_0_5_n80, npu_inst_pe_1_0_5_n79,
         npu_inst_pe_1_0_5_n78, npu_inst_pe_1_0_5_n77, npu_inst_pe_1_0_5_n76,
         npu_inst_pe_1_0_5_n75, npu_inst_pe_1_0_5_n74, npu_inst_pe_1_0_5_n73,
         npu_inst_pe_1_0_5_n72, npu_inst_pe_1_0_5_n71, npu_inst_pe_1_0_5_n70,
         npu_inst_pe_1_0_5_n69, npu_inst_pe_1_0_5_n68, npu_inst_pe_1_0_5_n67,
         npu_inst_pe_1_0_5_n66, npu_inst_pe_1_0_5_n65, npu_inst_pe_1_0_5_n64,
         npu_inst_pe_1_0_5_n63, npu_inst_pe_1_0_5_n62, npu_inst_pe_1_0_5_n61,
         npu_inst_pe_1_0_5_n60, npu_inst_pe_1_0_5_n59, npu_inst_pe_1_0_5_n58,
         npu_inst_pe_1_0_5_n57, npu_inst_pe_1_0_5_n56, npu_inst_pe_1_0_5_n55,
         npu_inst_pe_1_0_5_n54, npu_inst_pe_1_0_5_n53, npu_inst_pe_1_0_5_n52,
         npu_inst_pe_1_0_5_n51, npu_inst_pe_1_0_5_n50, npu_inst_pe_1_0_5_n49,
         npu_inst_pe_1_0_5_n48, npu_inst_pe_1_0_5_n47, npu_inst_pe_1_0_5_n46,
         npu_inst_pe_1_0_5_n45, npu_inst_pe_1_0_5_n44, npu_inst_pe_1_0_5_n43,
         npu_inst_pe_1_0_5_n42, npu_inst_pe_1_0_5_n41, npu_inst_pe_1_0_5_n40,
         npu_inst_pe_1_0_5_n39, npu_inst_pe_1_0_5_n38, npu_inst_pe_1_0_5_n37,
         npu_inst_pe_1_0_5_n27, npu_inst_pe_1_0_5_n26,
         npu_inst_pe_1_0_5_net4184, npu_inst_pe_1_0_5_net4178,
         npu_inst_pe_1_0_5_N94, npu_inst_pe_1_0_5_N93, npu_inst_pe_1_0_5_N84,
         npu_inst_pe_1_0_5_N80, npu_inst_pe_1_0_5_N79, npu_inst_pe_1_0_5_N78,
         npu_inst_pe_1_0_5_N77, npu_inst_pe_1_0_5_N76, npu_inst_pe_1_0_5_N75,
         npu_inst_pe_1_0_5_N74, npu_inst_pe_1_0_5_N73, npu_inst_pe_1_0_5_N72,
         npu_inst_pe_1_0_5_N71, npu_inst_pe_1_0_5_N70, npu_inst_pe_1_0_5_N69,
         npu_inst_pe_1_0_5_N68, npu_inst_pe_1_0_5_N67, npu_inst_pe_1_0_5_N66,
         npu_inst_pe_1_0_5_N65, npu_inst_pe_1_0_5_int_q_acc_0_,
         npu_inst_pe_1_0_5_int_q_acc_1_, npu_inst_pe_1_0_5_int_q_acc_2_,
         npu_inst_pe_1_0_5_int_q_acc_3_, npu_inst_pe_1_0_5_int_q_acc_4_,
         npu_inst_pe_1_0_5_int_q_acc_5_, npu_inst_pe_1_0_5_int_q_acc_6_,
         npu_inst_pe_1_0_5_int_q_acc_7_, npu_inst_pe_1_0_5_int_data_0_,
         npu_inst_pe_1_0_5_int_data_1_, npu_inst_pe_1_0_5_int_q_weight_0_,
         npu_inst_pe_1_0_5_int_q_weight_1_,
         npu_inst_pe_1_0_5_int_q_reg_v_5__0_,
         npu_inst_pe_1_0_5_int_q_reg_v_5__1_,
         npu_inst_pe_1_0_5_int_q_reg_v_4__0_,
         npu_inst_pe_1_0_5_int_q_reg_v_4__1_,
         npu_inst_pe_1_0_5_int_q_reg_v_3__0_,
         npu_inst_pe_1_0_5_int_q_reg_v_3__1_,
         npu_inst_pe_1_0_5_int_q_reg_v_2__0_,
         npu_inst_pe_1_0_5_int_q_reg_v_2__1_,
         npu_inst_pe_1_0_5_int_q_reg_v_1__0_,
         npu_inst_pe_1_0_5_int_q_reg_v_1__1_,
         npu_inst_pe_1_0_5_int_q_reg_v_0__0_,
         npu_inst_pe_1_0_5_int_q_reg_v_0__1_,
         npu_inst_pe_1_0_5_int_q_reg_h_5__0_,
         npu_inst_pe_1_0_5_int_q_reg_h_5__1_,
         npu_inst_pe_1_0_5_int_q_reg_h_4__0_,
         npu_inst_pe_1_0_5_int_q_reg_h_4__1_,
         npu_inst_pe_1_0_5_int_q_reg_h_3__0_,
         npu_inst_pe_1_0_5_int_q_reg_h_3__1_,
         npu_inst_pe_1_0_5_int_q_reg_h_2__0_,
         npu_inst_pe_1_0_5_int_q_reg_h_2__1_,
         npu_inst_pe_1_0_5_int_q_reg_h_1__0_,
         npu_inst_pe_1_0_5_int_q_reg_h_1__1_,
         npu_inst_pe_1_0_5_int_q_reg_h_0__0_,
         npu_inst_pe_1_0_5_int_q_reg_h_0__1_, npu_inst_pe_1_0_5_o_data_v_0_,
         npu_inst_pe_1_0_5_o_data_v_1_, npu_inst_pe_1_0_6_n119,
         npu_inst_pe_1_0_6_n118, npu_inst_pe_1_0_6_n117,
         npu_inst_pe_1_0_6_n116, npu_inst_pe_1_0_6_n115,
         npu_inst_pe_1_0_6_n114, npu_inst_pe_1_0_6_n113,
         npu_inst_pe_1_0_6_n112, npu_inst_pe_1_0_6_n111,
         npu_inst_pe_1_0_6_n110, npu_inst_pe_1_0_6_n109,
         npu_inst_pe_1_0_6_n108, npu_inst_pe_1_0_6_n107,
         npu_inst_pe_1_0_6_n106, npu_inst_pe_1_0_6_n105,
         npu_inst_pe_1_0_6_n104, npu_inst_pe_1_0_6_n103,
         npu_inst_pe_1_0_6_n102, npu_inst_pe_1_0_6_n101,
         npu_inst_pe_1_0_6_n100, npu_inst_pe_1_0_6_n99, npu_inst_pe_1_0_6_n98,
         npu_inst_pe_1_0_6_n36, npu_inst_pe_1_0_6_n35, npu_inst_pe_1_0_6_n34,
         npu_inst_pe_1_0_6_n33, npu_inst_pe_1_0_6_n32, npu_inst_pe_1_0_6_n31,
         npu_inst_pe_1_0_6_n30, npu_inst_pe_1_0_6_n29, npu_inst_pe_1_0_6_n28,
         npu_inst_pe_1_0_6_n25, npu_inst_pe_1_0_6_n24, npu_inst_pe_1_0_6_n23,
         npu_inst_pe_1_0_6_n22, npu_inst_pe_1_0_6_n21, npu_inst_pe_1_0_6_n20,
         npu_inst_pe_1_0_6_n19, npu_inst_pe_1_0_6_n18, npu_inst_pe_1_0_6_n17,
         npu_inst_pe_1_0_6_n16, npu_inst_pe_1_0_6_n15, npu_inst_pe_1_0_6_n14,
         npu_inst_pe_1_0_6_n13, npu_inst_pe_1_0_6_n12, npu_inst_pe_1_0_6_n11,
         npu_inst_pe_1_0_6_n10, npu_inst_pe_1_0_6_n9, npu_inst_pe_1_0_6_n8,
         npu_inst_pe_1_0_6_n7, npu_inst_pe_1_0_6_n6, npu_inst_pe_1_0_6_n5,
         npu_inst_pe_1_0_6_n4, npu_inst_pe_1_0_6_n3, npu_inst_pe_1_0_6_n2,
         npu_inst_pe_1_0_6_n1, npu_inst_pe_1_0_6_sub_77_carry_7_,
         npu_inst_pe_1_0_6_sub_77_carry_6_, npu_inst_pe_1_0_6_sub_77_carry_5_,
         npu_inst_pe_1_0_6_sub_77_carry_4_, npu_inst_pe_1_0_6_sub_77_carry_3_,
         npu_inst_pe_1_0_6_sub_77_carry_2_, npu_inst_pe_1_0_6_sub_77_carry_1_,
         npu_inst_pe_1_0_6_add_79_carry_7_, npu_inst_pe_1_0_6_add_79_carry_6_,
         npu_inst_pe_1_0_6_add_79_carry_5_, npu_inst_pe_1_0_6_add_79_carry_4_,
         npu_inst_pe_1_0_6_add_79_carry_3_, npu_inst_pe_1_0_6_add_79_carry_2_,
         npu_inst_pe_1_0_6_add_79_carry_1_, npu_inst_pe_1_0_6_n97,
         npu_inst_pe_1_0_6_n96, npu_inst_pe_1_0_6_n95, npu_inst_pe_1_0_6_n94,
         npu_inst_pe_1_0_6_n93, npu_inst_pe_1_0_6_n92, npu_inst_pe_1_0_6_n91,
         npu_inst_pe_1_0_6_n90, npu_inst_pe_1_0_6_n89, npu_inst_pe_1_0_6_n88,
         npu_inst_pe_1_0_6_n87, npu_inst_pe_1_0_6_n86, npu_inst_pe_1_0_6_n85,
         npu_inst_pe_1_0_6_n84, npu_inst_pe_1_0_6_n83, npu_inst_pe_1_0_6_n82,
         npu_inst_pe_1_0_6_n81, npu_inst_pe_1_0_6_n80, npu_inst_pe_1_0_6_n79,
         npu_inst_pe_1_0_6_n78, npu_inst_pe_1_0_6_n77, npu_inst_pe_1_0_6_n76,
         npu_inst_pe_1_0_6_n75, npu_inst_pe_1_0_6_n74, npu_inst_pe_1_0_6_n73,
         npu_inst_pe_1_0_6_n72, npu_inst_pe_1_0_6_n71, npu_inst_pe_1_0_6_n70,
         npu_inst_pe_1_0_6_n69, npu_inst_pe_1_0_6_n68, npu_inst_pe_1_0_6_n67,
         npu_inst_pe_1_0_6_n66, npu_inst_pe_1_0_6_n65, npu_inst_pe_1_0_6_n64,
         npu_inst_pe_1_0_6_n63, npu_inst_pe_1_0_6_n62, npu_inst_pe_1_0_6_n61,
         npu_inst_pe_1_0_6_n60, npu_inst_pe_1_0_6_n59, npu_inst_pe_1_0_6_n58,
         npu_inst_pe_1_0_6_n57, npu_inst_pe_1_0_6_n56, npu_inst_pe_1_0_6_n55,
         npu_inst_pe_1_0_6_n54, npu_inst_pe_1_0_6_n53, npu_inst_pe_1_0_6_n52,
         npu_inst_pe_1_0_6_n51, npu_inst_pe_1_0_6_n50, npu_inst_pe_1_0_6_n49,
         npu_inst_pe_1_0_6_n48, npu_inst_pe_1_0_6_n47, npu_inst_pe_1_0_6_n46,
         npu_inst_pe_1_0_6_n45, npu_inst_pe_1_0_6_n44, npu_inst_pe_1_0_6_n43,
         npu_inst_pe_1_0_6_n42, npu_inst_pe_1_0_6_n41, npu_inst_pe_1_0_6_n40,
         npu_inst_pe_1_0_6_n39, npu_inst_pe_1_0_6_n38, npu_inst_pe_1_0_6_n37,
         npu_inst_pe_1_0_6_n27, npu_inst_pe_1_0_6_n26,
         npu_inst_pe_1_0_6_net4161, npu_inst_pe_1_0_6_net4155,
         npu_inst_pe_1_0_6_N94, npu_inst_pe_1_0_6_N93, npu_inst_pe_1_0_6_N84,
         npu_inst_pe_1_0_6_N80, npu_inst_pe_1_0_6_N79, npu_inst_pe_1_0_6_N78,
         npu_inst_pe_1_0_6_N77, npu_inst_pe_1_0_6_N76, npu_inst_pe_1_0_6_N75,
         npu_inst_pe_1_0_6_N74, npu_inst_pe_1_0_6_N73, npu_inst_pe_1_0_6_N72,
         npu_inst_pe_1_0_6_N71, npu_inst_pe_1_0_6_N70, npu_inst_pe_1_0_6_N69,
         npu_inst_pe_1_0_6_N68, npu_inst_pe_1_0_6_N67, npu_inst_pe_1_0_6_N66,
         npu_inst_pe_1_0_6_N65, npu_inst_pe_1_0_6_int_q_acc_0_,
         npu_inst_pe_1_0_6_int_q_acc_1_, npu_inst_pe_1_0_6_int_q_acc_2_,
         npu_inst_pe_1_0_6_int_q_acc_3_, npu_inst_pe_1_0_6_int_q_acc_4_,
         npu_inst_pe_1_0_6_int_q_acc_5_, npu_inst_pe_1_0_6_int_q_acc_6_,
         npu_inst_pe_1_0_6_int_q_acc_7_, npu_inst_pe_1_0_6_int_data_0_,
         npu_inst_pe_1_0_6_int_data_1_, npu_inst_pe_1_0_6_int_q_weight_0_,
         npu_inst_pe_1_0_6_int_q_weight_1_,
         npu_inst_pe_1_0_6_int_q_reg_v_5__0_,
         npu_inst_pe_1_0_6_int_q_reg_v_5__1_,
         npu_inst_pe_1_0_6_int_q_reg_v_4__0_,
         npu_inst_pe_1_0_6_int_q_reg_v_4__1_,
         npu_inst_pe_1_0_6_int_q_reg_v_3__0_,
         npu_inst_pe_1_0_6_int_q_reg_v_3__1_,
         npu_inst_pe_1_0_6_int_q_reg_v_2__0_,
         npu_inst_pe_1_0_6_int_q_reg_v_2__1_,
         npu_inst_pe_1_0_6_int_q_reg_v_1__0_,
         npu_inst_pe_1_0_6_int_q_reg_v_1__1_,
         npu_inst_pe_1_0_6_int_q_reg_v_0__0_,
         npu_inst_pe_1_0_6_int_q_reg_v_0__1_,
         npu_inst_pe_1_0_6_int_q_reg_h_5__0_,
         npu_inst_pe_1_0_6_int_q_reg_h_5__1_,
         npu_inst_pe_1_0_6_int_q_reg_h_4__0_,
         npu_inst_pe_1_0_6_int_q_reg_h_4__1_,
         npu_inst_pe_1_0_6_int_q_reg_h_3__0_,
         npu_inst_pe_1_0_6_int_q_reg_h_3__1_,
         npu_inst_pe_1_0_6_int_q_reg_h_2__0_,
         npu_inst_pe_1_0_6_int_q_reg_h_2__1_,
         npu_inst_pe_1_0_6_int_q_reg_h_1__0_,
         npu_inst_pe_1_0_6_int_q_reg_h_1__1_,
         npu_inst_pe_1_0_6_int_q_reg_h_0__0_,
         npu_inst_pe_1_0_6_int_q_reg_h_0__1_, npu_inst_pe_1_0_6_o_data_v_0_,
         npu_inst_pe_1_0_6_o_data_v_1_, npu_inst_pe_1_0_7_n119,
         npu_inst_pe_1_0_7_n118, npu_inst_pe_1_0_7_n117,
         npu_inst_pe_1_0_7_n116, npu_inst_pe_1_0_7_n115,
         npu_inst_pe_1_0_7_n114, npu_inst_pe_1_0_7_n113,
         npu_inst_pe_1_0_7_n112, npu_inst_pe_1_0_7_n111,
         npu_inst_pe_1_0_7_n110, npu_inst_pe_1_0_7_n109,
         npu_inst_pe_1_0_7_n108, npu_inst_pe_1_0_7_n107,
         npu_inst_pe_1_0_7_n106, npu_inst_pe_1_0_7_n105,
         npu_inst_pe_1_0_7_n104, npu_inst_pe_1_0_7_n103,
         npu_inst_pe_1_0_7_n102, npu_inst_pe_1_0_7_n101,
         npu_inst_pe_1_0_7_n100, npu_inst_pe_1_0_7_n99, npu_inst_pe_1_0_7_n98,
         npu_inst_pe_1_0_7_n36, npu_inst_pe_1_0_7_n35, npu_inst_pe_1_0_7_n34,
         npu_inst_pe_1_0_7_n33, npu_inst_pe_1_0_7_n32, npu_inst_pe_1_0_7_n31,
         npu_inst_pe_1_0_7_n30, npu_inst_pe_1_0_7_n29, npu_inst_pe_1_0_7_n28,
         npu_inst_pe_1_0_7_n25, npu_inst_pe_1_0_7_n24, npu_inst_pe_1_0_7_n23,
         npu_inst_pe_1_0_7_n22, npu_inst_pe_1_0_7_n21, npu_inst_pe_1_0_7_n20,
         npu_inst_pe_1_0_7_n19, npu_inst_pe_1_0_7_n18, npu_inst_pe_1_0_7_n17,
         npu_inst_pe_1_0_7_n16, npu_inst_pe_1_0_7_n15, npu_inst_pe_1_0_7_n14,
         npu_inst_pe_1_0_7_n13, npu_inst_pe_1_0_7_n12, npu_inst_pe_1_0_7_n11,
         npu_inst_pe_1_0_7_n10, npu_inst_pe_1_0_7_n9, npu_inst_pe_1_0_7_n8,
         npu_inst_pe_1_0_7_n7, npu_inst_pe_1_0_7_n6, npu_inst_pe_1_0_7_n5,
         npu_inst_pe_1_0_7_n4, npu_inst_pe_1_0_7_n3, npu_inst_pe_1_0_7_n2,
         npu_inst_pe_1_0_7_n1, npu_inst_pe_1_0_7_sub_77_carry_7_,
         npu_inst_pe_1_0_7_sub_77_carry_6_, npu_inst_pe_1_0_7_sub_77_carry_5_,
         npu_inst_pe_1_0_7_sub_77_carry_4_, npu_inst_pe_1_0_7_sub_77_carry_3_,
         npu_inst_pe_1_0_7_sub_77_carry_2_, npu_inst_pe_1_0_7_sub_77_carry_1_,
         npu_inst_pe_1_0_7_add_79_carry_7_, npu_inst_pe_1_0_7_add_79_carry_6_,
         npu_inst_pe_1_0_7_add_79_carry_5_, npu_inst_pe_1_0_7_add_79_carry_4_,
         npu_inst_pe_1_0_7_add_79_carry_3_, npu_inst_pe_1_0_7_add_79_carry_2_,
         npu_inst_pe_1_0_7_add_79_carry_1_, npu_inst_pe_1_0_7_n97,
         npu_inst_pe_1_0_7_n96, npu_inst_pe_1_0_7_n95, npu_inst_pe_1_0_7_n94,
         npu_inst_pe_1_0_7_n93, npu_inst_pe_1_0_7_n92, npu_inst_pe_1_0_7_n91,
         npu_inst_pe_1_0_7_n90, npu_inst_pe_1_0_7_n89, npu_inst_pe_1_0_7_n88,
         npu_inst_pe_1_0_7_n87, npu_inst_pe_1_0_7_n86, npu_inst_pe_1_0_7_n85,
         npu_inst_pe_1_0_7_n84, npu_inst_pe_1_0_7_n83, npu_inst_pe_1_0_7_n82,
         npu_inst_pe_1_0_7_n81, npu_inst_pe_1_0_7_n80, npu_inst_pe_1_0_7_n79,
         npu_inst_pe_1_0_7_n78, npu_inst_pe_1_0_7_n77, npu_inst_pe_1_0_7_n76,
         npu_inst_pe_1_0_7_n75, npu_inst_pe_1_0_7_n74, npu_inst_pe_1_0_7_n73,
         npu_inst_pe_1_0_7_n72, npu_inst_pe_1_0_7_n71, npu_inst_pe_1_0_7_n70,
         npu_inst_pe_1_0_7_n69, npu_inst_pe_1_0_7_n68, npu_inst_pe_1_0_7_n67,
         npu_inst_pe_1_0_7_n66, npu_inst_pe_1_0_7_n65, npu_inst_pe_1_0_7_n64,
         npu_inst_pe_1_0_7_n63, npu_inst_pe_1_0_7_n62, npu_inst_pe_1_0_7_n61,
         npu_inst_pe_1_0_7_n60, npu_inst_pe_1_0_7_n59, npu_inst_pe_1_0_7_n58,
         npu_inst_pe_1_0_7_n57, npu_inst_pe_1_0_7_n56, npu_inst_pe_1_0_7_n55,
         npu_inst_pe_1_0_7_n54, npu_inst_pe_1_0_7_n53, npu_inst_pe_1_0_7_n52,
         npu_inst_pe_1_0_7_n51, npu_inst_pe_1_0_7_n50, npu_inst_pe_1_0_7_n49,
         npu_inst_pe_1_0_7_n48, npu_inst_pe_1_0_7_n47, npu_inst_pe_1_0_7_n46,
         npu_inst_pe_1_0_7_n45, npu_inst_pe_1_0_7_n44, npu_inst_pe_1_0_7_n43,
         npu_inst_pe_1_0_7_n42, npu_inst_pe_1_0_7_n41, npu_inst_pe_1_0_7_n40,
         npu_inst_pe_1_0_7_n39, npu_inst_pe_1_0_7_n38, npu_inst_pe_1_0_7_n37,
         npu_inst_pe_1_0_7_n27, npu_inst_pe_1_0_7_n26,
         npu_inst_pe_1_0_7_net4138, npu_inst_pe_1_0_7_net4132,
         npu_inst_pe_1_0_7_N94, npu_inst_pe_1_0_7_N93, npu_inst_pe_1_0_7_N84,
         npu_inst_pe_1_0_7_N80, npu_inst_pe_1_0_7_N79, npu_inst_pe_1_0_7_N78,
         npu_inst_pe_1_0_7_N77, npu_inst_pe_1_0_7_N76, npu_inst_pe_1_0_7_N75,
         npu_inst_pe_1_0_7_N74, npu_inst_pe_1_0_7_N73, npu_inst_pe_1_0_7_N72,
         npu_inst_pe_1_0_7_N71, npu_inst_pe_1_0_7_N70, npu_inst_pe_1_0_7_N69,
         npu_inst_pe_1_0_7_N68, npu_inst_pe_1_0_7_N67, npu_inst_pe_1_0_7_N66,
         npu_inst_pe_1_0_7_N65, npu_inst_pe_1_0_7_int_q_acc_0_,
         npu_inst_pe_1_0_7_int_q_acc_1_, npu_inst_pe_1_0_7_int_q_acc_2_,
         npu_inst_pe_1_0_7_int_q_acc_3_, npu_inst_pe_1_0_7_int_q_acc_4_,
         npu_inst_pe_1_0_7_int_q_acc_5_, npu_inst_pe_1_0_7_int_q_acc_6_,
         npu_inst_pe_1_0_7_int_q_acc_7_, npu_inst_pe_1_0_7_int_data_0_,
         npu_inst_pe_1_0_7_int_data_1_, npu_inst_pe_1_0_7_int_q_weight_0_,
         npu_inst_pe_1_0_7_int_q_weight_1_,
         npu_inst_pe_1_0_7_int_q_reg_v_5__0_,
         npu_inst_pe_1_0_7_int_q_reg_v_5__1_,
         npu_inst_pe_1_0_7_int_q_reg_v_4__0_,
         npu_inst_pe_1_0_7_int_q_reg_v_4__1_,
         npu_inst_pe_1_0_7_int_q_reg_v_3__0_,
         npu_inst_pe_1_0_7_int_q_reg_v_3__1_,
         npu_inst_pe_1_0_7_int_q_reg_v_2__0_,
         npu_inst_pe_1_0_7_int_q_reg_v_2__1_,
         npu_inst_pe_1_0_7_int_q_reg_v_1__0_,
         npu_inst_pe_1_0_7_int_q_reg_v_1__1_,
         npu_inst_pe_1_0_7_int_q_reg_v_0__0_,
         npu_inst_pe_1_0_7_int_q_reg_v_0__1_,
         npu_inst_pe_1_0_7_int_q_reg_h_5__0_,
         npu_inst_pe_1_0_7_int_q_reg_h_5__1_,
         npu_inst_pe_1_0_7_int_q_reg_h_4__0_,
         npu_inst_pe_1_0_7_int_q_reg_h_4__1_,
         npu_inst_pe_1_0_7_int_q_reg_h_3__0_,
         npu_inst_pe_1_0_7_int_q_reg_h_3__1_,
         npu_inst_pe_1_0_7_int_q_reg_h_2__0_,
         npu_inst_pe_1_0_7_int_q_reg_h_2__1_,
         npu_inst_pe_1_0_7_int_q_reg_h_1__0_,
         npu_inst_pe_1_0_7_int_q_reg_h_1__1_,
         npu_inst_pe_1_0_7_int_q_reg_h_0__0_,
         npu_inst_pe_1_0_7_int_q_reg_h_0__1_, npu_inst_pe_1_0_7_o_data_v_0_,
         npu_inst_pe_1_0_7_o_data_v_1_, npu_inst_pe_1_1_0_n119,
         npu_inst_pe_1_1_0_n118, npu_inst_pe_1_1_0_n117,
         npu_inst_pe_1_1_0_n116, npu_inst_pe_1_1_0_n115,
         npu_inst_pe_1_1_0_n114, npu_inst_pe_1_1_0_n113,
         npu_inst_pe_1_1_0_n112, npu_inst_pe_1_1_0_n111,
         npu_inst_pe_1_1_0_n110, npu_inst_pe_1_1_0_n109,
         npu_inst_pe_1_1_0_n108, npu_inst_pe_1_1_0_n107,
         npu_inst_pe_1_1_0_n106, npu_inst_pe_1_1_0_n105,
         npu_inst_pe_1_1_0_n104, npu_inst_pe_1_1_0_n103,
         npu_inst_pe_1_1_0_n102, npu_inst_pe_1_1_0_n101,
         npu_inst_pe_1_1_0_n100, npu_inst_pe_1_1_0_n99, npu_inst_pe_1_1_0_n98,
         npu_inst_pe_1_1_0_n36, npu_inst_pe_1_1_0_n35, npu_inst_pe_1_1_0_n34,
         npu_inst_pe_1_1_0_n33, npu_inst_pe_1_1_0_n32, npu_inst_pe_1_1_0_n31,
         npu_inst_pe_1_1_0_n30, npu_inst_pe_1_1_0_n29, npu_inst_pe_1_1_0_n28,
         npu_inst_pe_1_1_0_n25, npu_inst_pe_1_1_0_n24, npu_inst_pe_1_1_0_n23,
         npu_inst_pe_1_1_0_n22, npu_inst_pe_1_1_0_n21, npu_inst_pe_1_1_0_n20,
         npu_inst_pe_1_1_0_n19, npu_inst_pe_1_1_0_n18, npu_inst_pe_1_1_0_n17,
         npu_inst_pe_1_1_0_n16, npu_inst_pe_1_1_0_n15, npu_inst_pe_1_1_0_n14,
         npu_inst_pe_1_1_0_n13, npu_inst_pe_1_1_0_n12, npu_inst_pe_1_1_0_n11,
         npu_inst_pe_1_1_0_n10, npu_inst_pe_1_1_0_n9, npu_inst_pe_1_1_0_n8,
         npu_inst_pe_1_1_0_n7, npu_inst_pe_1_1_0_n6, npu_inst_pe_1_1_0_n5,
         npu_inst_pe_1_1_0_n4, npu_inst_pe_1_1_0_n3, npu_inst_pe_1_1_0_n2,
         npu_inst_pe_1_1_0_n1, npu_inst_pe_1_1_0_sub_77_carry_7_,
         npu_inst_pe_1_1_0_sub_77_carry_6_, npu_inst_pe_1_1_0_sub_77_carry_5_,
         npu_inst_pe_1_1_0_sub_77_carry_4_, npu_inst_pe_1_1_0_sub_77_carry_3_,
         npu_inst_pe_1_1_0_sub_77_carry_2_, npu_inst_pe_1_1_0_sub_77_carry_1_,
         npu_inst_pe_1_1_0_add_79_carry_7_, npu_inst_pe_1_1_0_add_79_carry_6_,
         npu_inst_pe_1_1_0_add_79_carry_5_, npu_inst_pe_1_1_0_add_79_carry_4_,
         npu_inst_pe_1_1_0_add_79_carry_3_, npu_inst_pe_1_1_0_add_79_carry_2_,
         npu_inst_pe_1_1_0_add_79_carry_1_, npu_inst_pe_1_1_0_n97,
         npu_inst_pe_1_1_0_n96, npu_inst_pe_1_1_0_n95, npu_inst_pe_1_1_0_n94,
         npu_inst_pe_1_1_0_n93, npu_inst_pe_1_1_0_n92, npu_inst_pe_1_1_0_n91,
         npu_inst_pe_1_1_0_n90, npu_inst_pe_1_1_0_n89, npu_inst_pe_1_1_0_n88,
         npu_inst_pe_1_1_0_n87, npu_inst_pe_1_1_0_n86, npu_inst_pe_1_1_0_n85,
         npu_inst_pe_1_1_0_n84, npu_inst_pe_1_1_0_n83, npu_inst_pe_1_1_0_n82,
         npu_inst_pe_1_1_0_n81, npu_inst_pe_1_1_0_n80, npu_inst_pe_1_1_0_n79,
         npu_inst_pe_1_1_0_n78, npu_inst_pe_1_1_0_n77, npu_inst_pe_1_1_0_n76,
         npu_inst_pe_1_1_0_n75, npu_inst_pe_1_1_0_n74, npu_inst_pe_1_1_0_n73,
         npu_inst_pe_1_1_0_n72, npu_inst_pe_1_1_0_n71, npu_inst_pe_1_1_0_n70,
         npu_inst_pe_1_1_0_n69, npu_inst_pe_1_1_0_n68, npu_inst_pe_1_1_0_n67,
         npu_inst_pe_1_1_0_n66, npu_inst_pe_1_1_0_n65, npu_inst_pe_1_1_0_n64,
         npu_inst_pe_1_1_0_n63, npu_inst_pe_1_1_0_n62, npu_inst_pe_1_1_0_n61,
         npu_inst_pe_1_1_0_n60, npu_inst_pe_1_1_0_n59, npu_inst_pe_1_1_0_n58,
         npu_inst_pe_1_1_0_n57, npu_inst_pe_1_1_0_n56, npu_inst_pe_1_1_0_n55,
         npu_inst_pe_1_1_0_n54, npu_inst_pe_1_1_0_n53, npu_inst_pe_1_1_0_n52,
         npu_inst_pe_1_1_0_n51, npu_inst_pe_1_1_0_n50, npu_inst_pe_1_1_0_n49,
         npu_inst_pe_1_1_0_n48, npu_inst_pe_1_1_0_n47, npu_inst_pe_1_1_0_n46,
         npu_inst_pe_1_1_0_n45, npu_inst_pe_1_1_0_n44, npu_inst_pe_1_1_0_n43,
         npu_inst_pe_1_1_0_n42, npu_inst_pe_1_1_0_n41, npu_inst_pe_1_1_0_n40,
         npu_inst_pe_1_1_0_n39, npu_inst_pe_1_1_0_n38, npu_inst_pe_1_1_0_n37,
         npu_inst_pe_1_1_0_n27, npu_inst_pe_1_1_0_n26,
         npu_inst_pe_1_1_0_net4115, npu_inst_pe_1_1_0_net4109,
         npu_inst_pe_1_1_0_N94, npu_inst_pe_1_1_0_N93, npu_inst_pe_1_1_0_N84,
         npu_inst_pe_1_1_0_N80, npu_inst_pe_1_1_0_N79, npu_inst_pe_1_1_0_N78,
         npu_inst_pe_1_1_0_N77, npu_inst_pe_1_1_0_N76, npu_inst_pe_1_1_0_N75,
         npu_inst_pe_1_1_0_N74, npu_inst_pe_1_1_0_N73, npu_inst_pe_1_1_0_N72,
         npu_inst_pe_1_1_0_N71, npu_inst_pe_1_1_0_N70, npu_inst_pe_1_1_0_N69,
         npu_inst_pe_1_1_0_N68, npu_inst_pe_1_1_0_N67, npu_inst_pe_1_1_0_N66,
         npu_inst_pe_1_1_0_N65, npu_inst_pe_1_1_0_int_q_acc_0_,
         npu_inst_pe_1_1_0_int_q_acc_1_, npu_inst_pe_1_1_0_int_q_acc_2_,
         npu_inst_pe_1_1_0_int_q_acc_3_, npu_inst_pe_1_1_0_int_q_acc_4_,
         npu_inst_pe_1_1_0_int_q_acc_5_, npu_inst_pe_1_1_0_int_q_acc_6_,
         npu_inst_pe_1_1_0_int_q_acc_7_, npu_inst_pe_1_1_0_int_data_0_,
         npu_inst_pe_1_1_0_int_data_1_, npu_inst_pe_1_1_0_int_q_weight_0_,
         npu_inst_pe_1_1_0_int_q_weight_1_,
         npu_inst_pe_1_1_0_int_q_reg_v_5__0_,
         npu_inst_pe_1_1_0_int_q_reg_v_5__1_,
         npu_inst_pe_1_1_0_int_q_reg_v_4__0_,
         npu_inst_pe_1_1_0_int_q_reg_v_4__1_,
         npu_inst_pe_1_1_0_int_q_reg_v_3__0_,
         npu_inst_pe_1_1_0_int_q_reg_v_3__1_,
         npu_inst_pe_1_1_0_int_q_reg_v_2__0_,
         npu_inst_pe_1_1_0_int_q_reg_v_2__1_,
         npu_inst_pe_1_1_0_int_q_reg_v_1__0_,
         npu_inst_pe_1_1_0_int_q_reg_v_1__1_,
         npu_inst_pe_1_1_0_int_q_reg_v_0__0_,
         npu_inst_pe_1_1_0_int_q_reg_v_0__1_,
         npu_inst_pe_1_1_0_int_q_reg_h_5__0_,
         npu_inst_pe_1_1_0_int_q_reg_h_5__1_,
         npu_inst_pe_1_1_0_int_q_reg_h_4__0_,
         npu_inst_pe_1_1_0_int_q_reg_h_4__1_,
         npu_inst_pe_1_1_0_int_q_reg_h_3__0_,
         npu_inst_pe_1_1_0_int_q_reg_h_3__1_,
         npu_inst_pe_1_1_0_int_q_reg_h_2__0_,
         npu_inst_pe_1_1_0_int_q_reg_h_2__1_,
         npu_inst_pe_1_1_0_int_q_reg_h_1__0_,
         npu_inst_pe_1_1_0_int_q_reg_h_1__1_,
         npu_inst_pe_1_1_0_int_q_reg_h_0__0_,
         npu_inst_pe_1_1_0_int_q_reg_h_0__1_, npu_inst_pe_1_1_0_o_data_h_0_,
         npu_inst_pe_1_1_0_o_data_h_1_, npu_inst_pe_1_1_1_n119,
         npu_inst_pe_1_1_1_n118, npu_inst_pe_1_1_1_n117,
         npu_inst_pe_1_1_1_n116, npu_inst_pe_1_1_1_n115,
         npu_inst_pe_1_1_1_n114, npu_inst_pe_1_1_1_n113,
         npu_inst_pe_1_1_1_n112, npu_inst_pe_1_1_1_n111,
         npu_inst_pe_1_1_1_n110, npu_inst_pe_1_1_1_n109,
         npu_inst_pe_1_1_1_n108, npu_inst_pe_1_1_1_n107,
         npu_inst_pe_1_1_1_n106, npu_inst_pe_1_1_1_n105,
         npu_inst_pe_1_1_1_n104, npu_inst_pe_1_1_1_n103,
         npu_inst_pe_1_1_1_n102, npu_inst_pe_1_1_1_n101,
         npu_inst_pe_1_1_1_n100, npu_inst_pe_1_1_1_n99, npu_inst_pe_1_1_1_n98,
         npu_inst_pe_1_1_1_n36, npu_inst_pe_1_1_1_n35, npu_inst_pe_1_1_1_n34,
         npu_inst_pe_1_1_1_n33, npu_inst_pe_1_1_1_n32, npu_inst_pe_1_1_1_n31,
         npu_inst_pe_1_1_1_n30, npu_inst_pe_1_1_1_n29, npu_inst_pe_1_1_1_n28,
         npu_inst_pe_1_1_1_n25, npu_inst_pe_1_1_1_n24, npu_inst_pe_1_1_1_n23,
         npu_inst_pe_1_1_1_n22, npu_inst_pe_1_1_1_n21, npu_inst_pe_1_1_1_n20,
         npu_inst_pe_1_1_1_n19, npu_inst_pe_1_1_1_n18, npu_inst_pe_1_1_1_n17,
         npu_inst_pe_1_1_1_n16, npu_inst_pe_1_1_1_n15, npu_inst_pe_1_1_1_n14,
         npu_inst_pe_1_1_1_n13, npu_inst_pe_1_1_1_n12, npu_inst_pe_1_1_1_n11,
         npu_inst_pe_1_1_1_n10, npu_inst_pe_1_1_1_n9, npu_inst_pe_1_1_1_n8,
         npu_inst_pe_1_1_1_n7, npu_inst_pe_1_1_1_n6, npu_inst_pe_1_1_1_n5,
         npu_inst_pe_1_1_1_n4, npu_inst_pe_1_1_1_n3, npu_inst_pe_1_1_1_n2,
         npu_inst_pe_1_1_1_n1, npu_inst_pe_1_1_1_sub_77_carry_7_,
         npu_inst_pe_1_1_1_sub_77_carry_6_, npu_inst_pe_1_1_1_sub_77_carry_5_,
         npu_inst_pe_1_1_1_sub_77_carry_4_, npu_inst_pe_1_1_1_sub_77_carry_3_,
         npu_inst_pe_1_1_1_sub_77_carry_2_, npu_inst_pe_1_1_1_sub_77_carry_1_,
         npu_inst_pe_1_1_1_add_79_carry_7_, npu_inst_pe_1_1_1_add_79_carry_6_,
         npu_inst_pe_1_1_1_add_79_carry_5_, npu_inst_pe_1_1_1_add_79_carry_4_,
         npu_inst_pe_1_1_1_add_79_carry_3_, npu_inst_pe_1_1_1_add_79_carry_2_,
         npu_inst_pe_1_1_1_add_79_carry_1_, npu_inst_pe_1_1_1_n97,
         npu_inst_pe_1_1_1_n96, npu_inst_pe_1_1_1_n95, npu_inst_pe_1_1_1_n94,
         npu_inst_pe_1_1_1_n93, npu_inst_pe_1_1_1_n92, npu_inst_pe_1_1_1_n91,
         npu_inst_pe_1_1_1_n90, npu_inst_pe_1_1_1_n89, npu_inst_pe_1_1_1_n88,
         npu_inst_pe_1_1_1_n87, npu_inst_pe_1_1_1_n86, npu_inst_pe_1_1_1_n85,
         npu_inst_pe_1_1_1_n84, npu_inst_pe_1_1_1_n83, npu_inst_pe_1_1_1_n82,
         npu_inst_pe_1_1_1_n81, npu_inst_pe_1_1_1_n80, npu_inst_pe_1_1_1_n79,
         npu_inst_pe_1_1_1_n78, npu_inst_pe_1_1_1_n77, npu_inst_pe_1_1_1_n76,
         npu_inst_pe_1_1_1_n75, npu_inst_pe_1_1_1_n74, npu_inst_pe_1_1_1_n73,
         npu_inst_pe_1_1_1_n72, npu_inst_pe_1_1_1_n71, npu_inst_pe_1_1_1_n70,
         npu_inst_pe_1_1_1_n69, npu_inst_pe_1_1_1_n68, npu_inst_pe_1_1_1_n67,
         npu_inst_pe_1_1_1_n66, npu_inst_pe_1_1_1_n65, npu_inst_pe_1_1_1_n64,
         npu_inst_pe_1_1_1_n63, npu_inst_pe_1_1_1_n62, npu_inst_pe_1_1_1_n61,
         npu_inst_pe_1_1_1_n60, npu_inst_pe_1_1_1_n59, npu_inst_pe_1_1_1_n58,
         npu_inst_pe_1_1_1_n57, npu_inst_pe_1_1_1_n56, npu_inst_pe_1_1_1_n55,
         npu_inst_pe_1_1_1_n54, npu_inst_pe_1_1_1_n53, npu_inst_pe_1_1_1_n52,
         npu_inst_pe_1_1_1_n51, npu_inst_pe_1_1_1_n50, npu_inst_pe_1_1_1_n49,
         npu_inst_pe_1_1_1_n48, npu_inst_pe_1_1_1_n47, npu_inst_pe_1_1_1_n46,
         npu_inst_pe_1_1_1_n45, npu_inst_pe_1_1_1_n44, npu_inst_pe_1_1_1_n43,
         npu_inst_pe_1_1_1_n42, npu_inst_pe_1_1_1_n41, npu_inst_pe_1_1_1_n40,
         npu_inst_pe_1_1_1_n39, npu_inst_pe_1_1_1_n38, npu_inst_pe_1_1_1_n37,
         npu_inst_pe_1_1_1_n27, npu_inst_pe_1_1_1_n26,
         npu_inst_pe_1_1_1_net4092, npu_inst_pe_1_1_1_net4086,
         npu_inst_pe_1_1_1_N94, npu_inst_pe_1_1_1_N93, npu_inst_pe_1_1_1_N84,
         npu_inst_pe_1_1_1_N80, npu_inst_pe_1_1_1_N79, npu_inst_pe_1_1_1_N78,
         npu_inst_pe_1_1_1_N77, npu_inst_pe_1_1_1_N76, npu_inst_pe_1_1_1_N75,
         npu_inst_pe_1_1_1_N74, npu_inst_pe_1_1_1_N73, npu_inst_pe_1_1_1_N72,
         npu_inst_pe_1_1_1_N71, npu_inst_pe_1_1_1_N70, npu_inst_pe_1_1_1_N69,
         npu_inst_pe_1_1_1_N68, npu_inst_pe_1_1_1_N67, npu_inst_pe_1_1_1_N66,
         npu_inst_pe_1_1_1_N65, npu_inst_pe_1_1_1_int_q_acc_0_,
         npu_inst_pe_1_1_1_int_q_acc_1_, npu_inst_pe_1_1_1_int_q_acc_2_,
         npu_inst_pe_1_1_1_int_q_acc_3_, npu_inst_pe_1_1_1_int_q_acc_4_,
         npu_inst_pe_1_1_1_int_q_acc_5_, npu_inst_pe_1_1_1_int_q_acc_6_,
         npu_inst_pe_1_1_1_int_q_acc_7_, npu_inst_pe_1_1_1_int_data_0_,
         npu_inst_pe_1_1_1_int_data_1_, npu_inst_pe_1_1_1_int_q_weight_0_,
         npu_inst_pe_1_1_1_int_q_weight_1_,
         npu_inst_pe_1_1_1_int_q_reg_v_5__0_,
         npu_inst_pe_1_1_1_int_q_reg_v_5__1_,
         npu_inst_pe_1_1_1_int_q_reg_v_4__0_,
         npu_inst_pe_1_1_1_int_q_reg_v_4__1_,
         npu_inst_pe_1_1_1_int_q_reg_v_3__0_,
         npu_inst_pe_1_1_1_int_q_reg_v_3__1_,
         npu_inst_pe_1_1_1_int_q_reg_v_2__0_,
         npu_inst_pe_1_1_1_int_q_reg_v_2__1_,
         npu_inst_pe_1_1_1_int_q_reg_v_1__0_,
         npu_inst_pe_1_1_1_int_q_reg_v_1__1_,
         npu_inst_pe_1_1_1_int_q_reg_v_0__0_,
         npu_inst_pe_1_1_1_int_q_reg_v_0__1_,
         npu_inst_pe_1_1_1_int_q_reg_h_5__0_,
         npu_inst_pe_1_1_1_int_q_reg_h_5__1_,
         npu_inst_pe_1_1_1_int_q_reg_h_4__0_,
         npu_inst_pe_1_1_1_int_q_reg_h_4__1_,
         npu_inst_pe_1_1_1_int_q_reg_h_3__0_,
         npu_inst_pe_1_1_1_int_q_reg_h_3__1_,
         npu_inst_pe_1_1_1_int_q_reg_h_2__0_,
         npu_inst_pe_1_1_1_int_q_reg_h_2__1_,
         npu_inst_pe_1_1_1_int_q_reg_h_1__0_,
         npu_inst_pe_1_1_1_int_q_reg_h_1__1_,
         npu_inst_pe_1_1_1_int_q_reg_h_0__0_,
         npu_inst_pe_1_1_1_int_q_reg_h_0__1_, npu_inst_pe_1_1_2_n119,
         npu_inst_pe_1_1_2_n118, npu_inst_pe_1_1_2_n117,
         npu_inst_pe_1_1_2_n116, npu_inst_pe_1_1_2_n115,
         npu_inst_pe_1_1_2_n114, npu_inst_pe_1_1_2_n113,
         npu_inst_pe_1_1_2_n112, npu_inst_pe_1_1_2_n111,
         npu_inst_pe_1_1_2_n110, npu_inst_pe_1_1_2_n109,
         npu_inst_pe_1_1_2_n108, npu_inst_pe_1_1_2_n107,
         npu_inst_pe_1_1_2_n106, npu_inst_pe_1_1_2_n105,
         npu_inst_pe_1_1_2_n104, npu_inst_pe_1_1_2_n103,
         npu_inst_pe_1_1_2_n102, npu_inst_pe_1_1_2_n101,
         npu_inst_pe_1_1_2_n100, npu_inst_pe_1_1_2_n99, npu_inst_pe_1_1_2_n98,
         npu_inst_pe_1_1_2_n36, npu_inst_pe_1_1_2_n35, npu_inst_pe_1_1_2_n34,
         npu_inst_pe_1_1_2_n33, npu_inst_pe_1_1_2_n32, npu_inst_pe_1_1_2_n31,
         npu_inst_pe_1_1_2_n30, npu_inst_pe_1_1_2_n29, npu_inst_pe_1_1_2_n28,
         npu_inst_pe_1_1_2_n25, npu_inst_pe_1_1_2_n24, npu_inst_pe_1_1_2_n23,
         npu_inst_pe_1_1_2_n22, npu_inst_pe_1_1_2_n21, npu_inst_pe_1_1_2_n20,
         npu_inst_pe_1_1_2_n19, npu_inst_pe_1_1_2_n18, npu_inst_pe_1_1_2_n17,
         npu_inst_pe_1_1_2_n16, npu_inst_pe_1_1_2_n15, npu_inst_pe_1_1_2_n14,
         npu_inst_pe_1_1_2_n13, npu_inst_pe_1_1_2_n12, npu_inst_pe_1_1_2_n11,
         npu_inst_pe_1_1_2_n10, npu_inst_pe_1_1_2_n9, npu_inst_pe_1_1_2_n8,
         npu_inst_pe_1_1_2_n7, npu_inst_pe_1_1_2_n6, npu_inst_pe_1_1_2_n5,
         npu_inst_pe_1_1_2_n4, npu_inst_pe_1_1_2_n3, npu_inst_pe_1_1_2_n2,
         npu_inst_pe_1_1_2_n1, npu_inst_pe_1_1_2_sub_77_carry_7_,
         npu_inst_pe_1_1_2_sub_77_carry_6_, npu_inst_pe_1_1_2_sub_77_carry_5_,
         npu_inst_pe_1_1_2_sub_77_carry_4_, npu_inst_pe_1_1_2_sub_77_carry_3_,
         npu_inst_pe_1_1_2_sub_77_carry_2_, npu_inst_pe_1_1_2_sub_77_carry_1_,
         npu_inst_pe_1_1_2_add_79_carry_7_, npu_inst_pe_1_1_2_add_79_carry_6_,
         npu_inst_pe_1_1_2_add_79_carry_5_, npu_inst_pe_1_1_2_add_79_carry_4_,
         npu_inst_pe_1_1_2_add_79_carry_3_, npu_inst_pe_1_1_2_add_79_carry_2_,
         npu_inst_pe_1_1_2_add_79_carry_1_, npu_inst_pe_1_1_2_n97,
         npu_inst_pe_1_1_2_n96, npu_inst_pe_1_1_2_n95, npu_inst_pe_1_1_2_n94,
         npu_inst_pe_1_1_2_n93, npu_inst_pe_1_1_2_n92, npu_inst_pe_1_1_2_n91,
         npu_inst_pe_1_1_2_n90, npu_inst_pe_1_1_2_n89, npu_inst_pe_1_1_2_n88,
         npu_inst_pe_1_1_2_n87, npu_inst_pe_1_1_2_n86, npu_inst_pe_1_1_2_n85,
         npu_inst_pe_1_1_2_n84, npu_inst_pe_1_1_2_n83, npu_inst_pe_1_1_2_n82,
         npu_inst_pe_1_1_2_n81, npu_inst_pe_1_1_2_n80, npu_inst_pe_1_1_2_n79,
         npu_inst_pe_1_1_2_n78, npu_inst_pe_1_1_2_n77, npu_inst_pe_1_1_2_n76,
         npu_inst_pe_1_1_2_n75, npu_inst_pe_1_1_2_n74, npu_inst_pe_1_1_2_n73,
         npu_inst_pe_1_1_2_n72, npu_inst_pe_1_1_2_n71, npu_inst_pe_1_1_2_n70,
         npu_inst_pe_1_1_2_n69, npu_inst_pe_1_1_2_n68, npu_inst_pe_1_1_2_n67,
         npu_inst_pe_1_1_2_n66, npu_inst_pe_1_1_2_n65, npu_inst_pe_1_1_2_n64,
         npu_inst_pe_1_1_2_n63, npu_inst_pe_1_1_2_n62, npu_inst_pe_1_1_2_n61,
         npu_inst_pe_1_1_2_n60, npu_inst_pe_1_1_2_n59, npu_inst_pe_1_1_2_n58,
         npu_inst_pe_1_1_2_n57, npu_inst_pe_1_1_2_n56, npu_inst_pe_1_1_2_n55,
         npu_inst_pe_1_1_2_n54, npu_inst_pe_1_1_2_n53, npu_inst_pe_1_1_2_n52,
         npu_inst_pe_1_1_2_n51, npu_inst_pe_1_1_2_n50, npu_inst_pe_1_1_2_n49,
         npu_inst_pe_1_1_2_n48, npu_inst_pe_1_1_2_n47, npu_inst_pe_1_1_2_n46,
         npu_inst_pe_1_1_2_n45, npu_inst_pe_1_1_2_n44, npu_inst_pe_1_1_2_n43,
         npu_inst_pe_1_1_2_n42, npu_inst_pe_1_1_2_n41, npu_inst_pe_1_1_2_n40,
         npu_inst_pe_1_1_2_n39, npu_inst_pe_1_1_2_n38, npu_inst_pe_1_1_2_n37,
         npu_inst_pe_1_1_2_n27, npu_inst_pe_1_1_2_n26,
         npu_inst_pe_1_1_2_net4069, npu_inst_pe_1_1_2_net4063,
         npu_inst_pe_1_1_2_N94, npu_inst_pe_1_1_2_N93, npu_inst_pe_1_1_2_N84,
         npu_inst_pe_1_1_2_N80, npu_inst_pe_1_1_2_N79, npu_inst_pe_1_1_2_N78,
         npu_inst_pe_1_1_2_N77, npu_inst_pe_1_1_2_N76, npu_inst_pe_1_1_2_N75,
         npu_inst_pe_1_1_2_N74, npu_inst_pe_1_1_2_N73, npu_inst_pe_1_1_2_N72,
         npu_inst_pe_1_1_2_N71, npu_inst_pe_1_1_2_N70, npu_inst_pe_1_1_2_N69,
         npu_inst_pe_1_1_2_N68, npu_inst_pe_1_1_2_N67, npu_inst_pe_1_1_2_N66,
         npu_inst_pe_1_1_2_N65, npu_inst_pe_1_1_2_int_q_acc_0_,
         npu_inst_pe_1_1_2_int_q_acc_1_, npu_inst_pe_1_1_2_int_q_acc_2_,
         npu_inst_pe_1_1_2_int_q_acc_3_, npu_inst_pe_1_1_2_int_q_acc_4_,
         npu_inst_pe_1_1_2_int_q_acc_5_, npu_inst_pe_1_1_2_int_q_acc_6_,
         npu_inst_pe_1_1_2_int_q_acc_7_, npu_inst_pe_1_1_2_int_data_0_,
         npu_inst_pe_1_1_2_int_data_1_, npu_inst_pe_1_1_2_int_q_weight_0_,
         npu_inst_pe_1_1_2_int_q_weight_1_,
         npu_inst_pe_1_1_2_int_q_reg_v_5__0_,
         npu_inst_pe_1_1_2_int_q_reg_v_5__1_,
         npu_inst_pe_1_1_2_int_q_reg_v_4__0_,
         npu_inst_pe_1_1_2_int_q_reg_v_4__1_,
         npu_inst_pe_1_1_2_int_q_reg_v_3__0_,
         npu_inst_pe_1_1_2_int_q_reg_v_3__1_,
         npu_inst_pe_1_1_2_int_q_reg_v_2__0_,
         npu_inst_pe_1_1_2_int_q_reg_v_2__1_,
         npu_inst_pe_1_1_2_int_q_reg_v_1__0_,
         npu_inst_pe_1_1_2_int_q_reg_v_1__1_,
         npu_inst_pe_1_1_2_int_q_reg_v_0__0_,
         npu_inst_pe_1_1_2_int_q_reg_v_0__1_,
         npu_inst_pe_1_1_2_int_q_reg_h_5__0_,
         npu_inst_pe_1_1_2_int_q_reg_h_5__1_,
         npu_inst_pe_1_1_2_int_q_reg_h_4__0_,
         npu_inst_pe_1_1_2_int_q_reg_h_4__1_,
         npu_inst_pe_1_1_2_int_q_reg_h_3__0_,
         npu_inst_pe_1_1_2_int_q_reg_h_3__1_,
         npu_inst_pe_1_1_2_int_q_reg_h_2__0_,
         npu_inst_pe_1_1_2_int_q_reg_h_2__1_,
         npu_inst_pe_1_1_2_int_q_reg_h_1__0_,
         npu_inst_pe_1_1_2_int_q_reg_h_1__1_,
         npu_inst_pe_1_1_2_int_q_reg_h_0__0_,
         npu_inst_pe_1_1_2_int_q_reg_h_0__1_, npu_inst_pe_1_1_3_n119,
         npu_inst_pe_1_1_3_n118, npu_inst_pe_1_1_3_n117,
         npu_inst_pe_1_1_3_n116, npu_inst_pe_1_1_3_n115,
         npu_inst_pe_1_1_3_n114, npu_inst_pe_1_1_3_n113,
         npu_inst_pe_1_1_3_n112, npu_inst_pe_1_1_3_n111,
         npu_inst_pe_1_1_3_n110, npu_inst_pe_1_1_3_n109,
         npu_inst_pe_1_1_3_n108, npu_inst_pe_1_1_3_n107,
         npu_inst_pe_1_1_3_n106, npu_inst_pe_1_1_3_n105,
         npu_inst_pe_1_1_3_n104, npu_inst_pe_1_1_3_n103,
         npu_inst_pe_1_1_3_n102, npu_inst_pe_1_1_3_n101,
         npu_inst_pe_1_1_3_n100, npu_inst_pe_1_1_3_n99, npu_inst_pe_1_1_3_n98,
         npu_inst_pe_1_1_3_n36, npu_inst_pe_1_1_3_n35, npu_inst_pe_1_1_3_n34,
         npu_inst_pe_1_1_3_n33, npu_inst_pe_1_1_3_n32, npu_inst_pe_1_1_3_n31,
         npu_inst_pe_1_1_3_n30, npu_inst_pe_1_1_3_n29, npu_inst_pe_1_1_3_n28,
         npu_inst_pe_1_1_3_n25, npu_inst_pe_1_1_3_n24, npu_inst_pe_1_1_3_n23,
         npu_inst_pe_1_1_3_n22, npu_inst_pe_1_1_3_n21, npu_inst_pe_1_1_3_n20,
         npu_inst_pe_1_1_3_n19, npu_inst_pe_1_1_3_n18, npu_inst_pe_1_1_3_n17,
         npu_inst_pe_1_1_3_n16, npu_inst_pe_1_1_3_n15, npu_inst_pe_1_1_3_n14,
         npu_inst_pe_1_1_3_n13, npu_inst_pe_1_1_3_n12, npu_inst_pe_1_1_3_n11,
         npu_inst_pe_1_1_3_n10, npu_inst_pe_1_1_3_n9, npu_inst_pe_1_1_3_n8,
         npu_inst_pe_1_1_3_n7, npu_inst_pe_1_1_3_n6, npu_inst_pe_1_1_3_n5,
         npu_inst_pe_1_1_3_n4, npu_inst_pe_1_1_3_n3, npu_inst_pe_1_1_3_n2,
         npu_inst_pe_1_1_3_n1, npu_inst_pe_1_1_3_sub_77_carry_7_,
         npu_inst_pe_1_1_3_sub_77_carry_6_, npu_inst_pe_1_1_3_sub_77_carry_5_,
         npu_inst_pe_1_1_3_sub_77_carry_4_, npu_inst_pe_1_1_3_sub_77_carry_3_,
         npu_inst_pe_1_1_3_sub_77_carry_2_, npu_inst_pe_1_1_3_sub_77_carry_1_,
         npu_inst_pe_1_1_3_add_79_carry_7_, npu_inst_pe_1_1_3_add_79_carry_6_,
         npu_inst_pe_1_1_3_add_79_carry_5_, npu_inst_pe_1_1_3_add_79_carry_4_,
         npu_inst_pe_1_1_3_add_79_carry_3_, npu_inst_pe_1_1_3_add_79_carry_2_,
         npu_inst_pe_1_1_3_add_79_carry_1_, npu_inst_pe_1_1_3_n97,
         npu_inst_pe_1_1_3_n96, npu_inst_pe_1_1_3_n95, npu_inst_pe_1_1_3_n94,
         npu_inst_pe_1_1_3_n93, npu_inst_pe_1_1_3_n92, npu_inst_pe_1_1_3_n91,
         npu_inst_pe_1_1_3_n90, npu_inst_pe_1_1_3_n89, npu_inst_pe_1_1_3_n88,
         npu_inst_pe_1_1_3_n87, npu_inst_pe_1_1_3_n86, npu_inst_pe_1_1_3_n85,
         npu_inst_pe_1_1_3_n84, npu_inst_pe_1_1_3_n83, npu_inst_pe_1_1_3_n82,
         npu_inst_pe_1_1_3_n81, npu_inst_pe_1_1_3_n80, npu_inst_pe_1_1_3_n79,
         npu_inst_pe_1_1_3_n78, npu_inst_pe_1_1_3_n77, npu_inst_pe_1_1_3_n76,
         npu_inst_pe_1_1_3_n75, npu_inst_pe_1_1_3_n74, npu_inst_pe_1_1_3_n73,
         npu_inst_pe_1_1_3_n72, npu_inst_pe_1_1_3_n71, npu_inst_pe_1_1_3_n70,
         npu_inst_pe_1_1_3_n69, npu_inst_pe_1_1_3_n68, npu_inst_pe_1_1_3_n67,
         npu_inst_pe_1_1_3_n66, npu_inst_pe_1_1_3_n65, npu_inst_pe_1_1_3_n64,
         npu_inst_pe_1_1_3_n63, npu_inst_pe_1_1_3_n62, npu_inst_pe_1_1_3_n61,
         npu_inst_pe_1_1_3_n60, npu_inst_pe_1_1_3_n59, npu_inst_pe_1_1_3_n58,
         npu_inst_pe_1_1_3_n57, npu_inst_pe_1_1_3_n56, npu_inst_pe_1_1_3_n55,
         npu_inst_pe_1_1_3_n54, npu_inst_pe_1_1_3_n53, npu_inst_pe_1_1_3_n52,
         npu_inst_pe_1_1_3_n51, npu_inst_pe_1_1_3_n50, npu_inst_pe_1_1_3_n49,
         npu_inst_pe_1_1_3_n48, npu_inst_pe_1_1_3_n47, npu_inst_pe_1_1_3_n46,
         npu_inst_pe_1_1_3_n45, npu_inst_pe_1_1_3_n44, npu_inst_pe_1_1_3_n43,
         npu_inst_pe_1_1_3_n42, npu_inst_pe_1_1_3_n41, npu_inst_pe_1_1_3_n40,
         npu_inst_pe_1_1_3_n39, npu_inst_pe_1_1_3_n38, npu_inst_pe_1_1_3_n37,
         npu_inst_pe_1_1_3_n27, npu_inst_pe_1_1_3_n26,
         npu_inst_pe_1_1_3_net4046, npu_inst_pe_1_1_3_net4040,
         npu_inst_pe_1_1_3_N94, npu_inst_pe_1_1_3_N93, npu_inst_pe_1_1_3_N84,
         npu_inst_pe_1_1_3_N80, npu_inst_pe_1_1_3_N79, npu_inst_pe_1_1_3_N78,
         npu_inst_pe_1_1_3_N77, npu_inst_pe_1_1_3_N76, npu_inst_pe_1_1_3_N75,
         npu_inst_pe_1_1_3_N74, npu_inst_pe_1_1_3_N73, npu_inst_pe_1_1_3_N72,
         npu_inst_pe_1_1_3_N71, npu_inst_pe_1_1_3_N70, npu_inst_pe_1_1_3_N69,
         npu_inst_pe_1_1_3_N68, npu_inst_pe_1_1_3_N67, npu_inst_pe_1_1_3_N66,
         npu_inst_pe_1_1_3_N65, npu_inst_pe_1_1_3_int_q_acc_0_,
         npu_inst_pe_1_1_3_int_q_acc_1_, npu_inst_pe_1_1_3_int_q_acc_2_,
         npu_inst_pe_1_1_3_int_q_acc_3_, npu_inst_pe_1_1_3_int_q_acc_4_,
         npu_inst_pe_1_1_3_int_q_acc_5_, npu_inst_pe_1_1_3_int_q_acc_6_,
         npu_inst_pe_1_1_3_int_q_acc_7_, npu_inst_pe_1_1_3_int_data_0_,
         npu_inst_pe_1_1_3_int_data_1_, npu_inst_pe_1_1_3_int_q_weight_0_,
         npu_inst_pe_1_1_3_int_q_weight_1_,
         npu_inst_pe_1_1_3_int_q_reg_v_5__0_,
         npu_inst_pe_1_1_3_int_q_reg_v_5__1_,
         npu_inst_pe_1_1_3_int_q_reg_v_4__0_,
         npu_inst_pe_1_1_3_int_q_reg_v_4__1_,
         npu_inst_pe_1_1_3_int_q_reg_v_3__0_,
         npu_inst_pe_1_1_3_int_q_reg_v_3__1_,
         npu_inst_pe_1_1_3_int_q_reg_v_2__0_,
         npu_inst_pe_1_1_3_int_q_reg_v_2__1_,
         npu_inst_pe_1_1_3_int_q_reg_v_1__0_,
         npu_inst_pe_1_1_3_int_q_reg_v_1__1_,
         npu_inst_pe_1_1_3_int_q_reg_v_0__0_,
         npu_inst_pe_1_1_3_int_q_reg_v_0__1_,
         npu_inst_pe_1_1_3_int_q_reg_h_5__0_,
         npu_inst_pe_1_1_3_int_q_reg_h_5__1_,
         npu_inst_pe_1_1_3_int_q_reg_h_4__0_,
         npu_inst_pe_1_1_3_int_q_reg_h_4__1_,
         npu_inst_pe_1_1_3_int_q_reg_h_3__0_,
         npu_inst_pe_1_1_3_int_q_reg_h_3__1_,
         npu_inst_pe_1_1_3_int_q_reg_h_2__0_,
         npu_inst_pe_1_1_3_int_q_reg_h_2__1_,
         npu_inst_pe_1_1_3_int_q_reg_h_1__0_,
         npu_inst_pe_1_1_3_int_q_reg_h_1__1_,
         npu_inst_pe_1_1_3_int_q_reg_h_0__0_,
         npu_inst_pe_1_1_3_int_q_reg_h_0__1_, npu_inst_pe_1_1_4_n119,
         npu_inst_pe_1_1_4_n118, npu_inst_pe_1_1_4_n117,
         npu_inst_pe_1_1_4_n116, npu_inst_pe_1_1_4_n115,
         npu_inst_pe_1_1_4_n114, npu_inst_pe_1_1_4_n113,
         npu_inst_pe_1_1_4_n112, npu_inst_pe_1_1_4_n111,
         npu_inst_pe_1_1_4_n110, npu_inst_pe_1_1_4_n109,
         npu_inst_pe_1_1_4_n108, npu_inst_pe_1_1_4_n107,
         npu_inst_pe_1_1_4_n106, npu_inst_pe_1_1_4_n105,
         npu_inst_pe_1_1_4_n104, npu_inst_pe_1_1_4_n103,
         npu_inst_pe_1_1_4_n102, npu_inst_pe_1_1_4_n101,
         npu_inst_pe_1_1_4_n100, npu_inst_pe_1_1_4_n99, npu_inst_pe_1_1_4_n98,
         npu_inst_pe_1_1_4_n36, npu_inst_pe_1_1_4_n35, npu_inst_pe_1_1_4_n34,
         npu_inst_pe_1_1_4_n33, npu_inst_pe_1_1_4_n32, npu_inst_pe_1_1_4_n31,
         npu_inst_pe_1_1_4_n30, npu_inst_pe_1_1_4_n29, npu_inst_pe_1_1_4_n28,
         npu_inst_pe_1_1_4_n25, npu_inst_pe_1_1_4_n24, npu_inst_pe_1_1_4_n23,
         npu_inst_pe_1_1_4_n22, npu_inst_pe_1_1_4_n21, npu_inst_pe_1_1_4_n20,
         npu_inst_pe_1_1_4_n19, npu_inst_pe_1_1_4_n18, npu_inst_pe_1_1_4_n17,
         npu_inst_pe_1_1_4_n16, npu_inst_pe_1_1_4_n15, npu_inst_pe_1_1_4_n14,
         npu_inst_pe_1_1_4_n13, npu_inst_pe_1_1_4_n12, npu_inst_pe_1_1_4_n11,
         npu_inst_pe_1_1_4_n10, npu_inst_pe_1_1_4_n9, npu_inst_pe_1_1_4_n8,
         npu_inst_pe_1_1_4_n7, npu_inst_pe_1_1_4_n6, npu_inst_pe_1_1_4_n5,
         npu_inst_pe_1_1_4_n4, npu_inst_pe_1_1_4_n3, npu_inst_pe_1_1_4_n2,
         npu_inst_pe_1_1_4_n1, npu_inst_pe_1_1_4_sub_77_carry_7_,
         npu_inst_pe_1_1_4_sub_77_carry_6_, npu_inst_pe_1_1_4_sub_77_carry_5_,
         npu_inst_pe_1_1_4_sub_77_carry_4_, npu_inst_pe_1_1_4_sub_77_carry_3_,
         npu_inst_pe_1_1_4_sub_77_carry_2_, npu_inst_pe_1_1_4_sub_77_carry_1_,
         npu_inst_pe_1_1_4_add_79_carry_7_, npu_inst_pe_1_1_4_add_79_carry_6_,
         npu_inst_pe_1_1_4_add_79_carry_5_, npu_inst_pe_1_1_4_add_79_carry_4_,
         npu_inst_pe_1_1_4_add_79_carry_3_, npu_inst_pe_1_1_4_add_79_carry_2_,
         npu_inst_pe_1_1_4_add_79_carry_1_, npu_inst_pe_1_1_4_n97,
         npu_inst_pe_1_1_4_n96, npu_inst_pe_1_1_4_n95, npu_inst_pe_1_1_4_n94,
         npu_inst_pe_1_1_4_n93, npu_inst_pe_1_1_4_n92, npu_inst_pe_1_1_4_n91,
         npu_inst_pe_1_1_4_n90, npu_inst_pe_1_1_4_n89, npu_inst_pe_1_1_4_n88,
         npu_inst_pe_1_1_4_n87, npu_inst_pe_1_1_4_n86, npu_inst_pe_1_1_4_n85,
         npu_inst_pe_1_1_4_n84, npu_inst_pe_1_1_4_n83, npu_inst_pe_1_1_4_n82,
         npu_inst_pe_1_1_4_n81, npu_inst_pe_1_1_4_n80, npu_inst_pe_1_1_4_n79,
         npu_inst_pe_1_1_4_n78, npu_inst_pe_1_1_4_n77, npu_inst_pe_1_1_4_n76,
         npu_inst_pe_1_1_4_n75, npu_inst_pe_1_1_4_n74, npu_inst_pe_1_1_4_n73,
         npu_inst_pe_1_1_4_n72, npu_inst_pe_1_1_4_n71, npu_inst_pe_1_1_4_n70,
         npu_inst_pe_1_1_4_n69, npu_inst_pe_1_1_4_n68, npu_inst_pe_1_1_4_n67,
         npu_inst_pe_1_1_4_n66, npu_inst_pe_1_1_4_n65, npu_inst_pe_1_1_4_n64,
         npu_inst_pe_1_1_4_n63, npu_inst_pe_1_1_4_n62, npu_inst_pe_1_1_4_n61,
         npu_inst_pe_1_1_4_n60, npu_inst_pe_1_1_4_n59, npu_inst_pe_1_1_4_n58,
         npu_inst_pe_1_1_4_n57, npu_inst_pe_1_1_4_n56, npu_inst_pe_1_1_4_n55,
         npu_inst_pe_1_1_4_n54, npu_inst_pe_1_1_4_n53, npu_inst_pe_1_1_4_n52,
         npu_inst_pe_1_1_4_n51, npu_inst_pe_1_1_4_n50, npu_inst_pe_1_1_4_n49,
         npu_inst_pe_1_1_4_n48, npu_inst_pe_1_1_4_n47, npu_inst_pe_1_1_4_n46,
         npu_inst_pe_1_1_4_n45, npu_inst_pe_1_1_4_n44, npu_inst_pe_1_1_4_n43,
         npu_inst_pe_1_1_4_n42, npu_inst_pe_1_1_4_n41, npu_inst_pe_1_1_4_n40,
         npu_inst_pe_1_1_4_n39, npu_inst_pe_1_1_4_n38, npu_inst_pe_1_1_4_n37,
         npu_inst_pe_1_1_4_n27, npu_inst_pe_1_1_4_n26,
         npu_inst_pe_1_1_4_net4023, npu_inst_pe_1_1_4_net4017,
         npu_inst_pe_1_1_4_N94, npu_inst_pe_1_1_4_N93, npu_inst_pe_1_1_4_N84,
         npu_inst_pe_1_1_4_N80, npu_inst_pe_1_1_4_N79, npu_inst_pe_1_1_4_N78,
         npu_inst_pe_1_1_4_N77, npu_inst_pe_1_1_4_N76, npu_inst_pe_1_1_4_N75,
         npu_inst_pe_1_1_4_N74, npu_inst_pe_1_1_4_N73, npu_inst_pe_1_1_4_N72,
         npu_inst_pe_1_1_4_N71, npu_inst_pe_1_1_4_N70, npu_inst_pe_1_1_4_N69,
         npu_inst_pe_1_1_4_N68, npu_inst_pe_1_1_4_N67, npu_inst_pe_1_1_4_N66,
         npu_inst_pe_1_1_4_N65, npu_inst_pe_1_1_4_int_q_acc_0_,
         npu_inst_pe_1_1_4_int_q_acc_1_, npu_inst_pe_1_1_4_int_q_acc_2_,
         npu_inst_pe_1_1_4_int_q_acc_3_, npu_inst_pe_1_1_4_int_q_acc_4_,
         npu_inst_pe_1_1_4_int_q_acc_5_, npu_inst_pe_1_1_4_int_q_acc_6_,
         npu_inst_pe_1_1_4_int_q_acc_7_, npu_inst_pe_1_1_4_int_data_0_,
         npu_inst_pe_1_1_4_int_data_1_, npu_inst_pe_1_1_4_int_q_weight_0_,
         npu_inst_pe_1_1_4_int_q_weight_1_,
         npu_inst_pe_1_1_4_int_q_reg_v_5__0_,
         npu_inst_pe_1_1_4_int_q_reg_v_5__1_,
         npu_inst_pe_1_1_4_int_q_reg_v_4__0_,
         npu_inst_pe_1_1_4_int_q_reg_v_4__1_,
         npu_inst_pe_1_1_4_int_q_reg_v_3__0_,
         npu_inst_pe_1_1_4_int_q_reg_v_3__1_,
         npu_inst_pe_1_1_4_int_q_reg_v_2__0_,
         npu_inst_pe_1_1_4_int_q_reg_v_2__1_,
         npu_inst_pe_1_1_4_int_q_reg_v_1__0_,
         npu_inst_pe_1_1_4_int_q_reg_v_1__1_,
         npu_inst_pe_1_1_4_int_q_reg_v_0__0_,
         npu_inst_pe_1_1_4_int_q_reg_v_0__1_,
         npu_inst_pe_1_1_4_int_q_reg_h_5__0_,
         npu_inst_pe_1_1_4_int_q_reg_h_5__1_,
         npu_inst_pe_1_1_4_int_q_reg_h_4__0_,
         npu_inst_pe_1_1_4_int_q_reg_h_4__1_,
         npu_inst_pe_1_1_4_int_q_reg_h_3__0_,
         npu_inst_pe_1_1_4_int_q_reg_h_3__1_,
         npu_inst_pe_1_1_4_int_q_reg_h_2__0_,
         npu_inst_pe_1_1_4_int_q_reg_h_2__1_,
         npu_inst_pe_1_1_4_int_q_reg_h_1__0_,
         npu_inst_pe_1_1_4_int_q_reg_h_1__1_,
         npu_inst_pe_1_1_4_int_q_reg_h_0__0_,
         npu_inst_pe_1_1_4_int_q_reg_h_0__1_, npu_inst_pe_1_1_5_n119,
         npu_inst_pe_1_1_5_n118, npu_inst_pe_1_1_5_n117,
         npu_inst_pe_1_1_5_n116, npu_inst_pe_1_1_5_n115,
         npu_inst_pe_1_1_5_n114, npu_inst_pe_1_1_5_n113,
         npu_inst_pe_1_1_5_n112, npu_inst_pe_1_1_5_n111,
         npu_inst_pe_1_1_5_n110, npu_inst_pe_1_1_5_n109,
         npu_inst_pe_1_1_5_n108, npu_inst_pe_1_1_5_n107,
         npu_inst_pe_1_1_5_n106, npu_inst_pe_1_1_5_n105,
         npu_inst_pe_1_1_5_n104, npu_inst_pe_1_1_5_n103,
         npu_inst_pe_1_1_5_n102, npu_inst_pe_1_1_5_n101,
         npu_inst_pe_1_1_5_n100, npu_inst_pe_1_1_5_n99, npu_inst_pe_1_1_5_n98,
         npu_inst_pe_1_1_5_n36, npu_inst_pe_1_1_5_n35, npu_inst_pe_1_1_5_n34,
         npu_inst_pe_1_1_5_n33, npu_inst_pe_1_1_5_n32, npu_inst_pe_1_1_5_n31,
         npu_inst_pe_1_1_5_n30, npu_inst_pe_1_1_5_n29, npu_inst_pe_1_1_5_n28,
         npu_inst_pe_1_1_5_n25, npu_inst_pe_1_1_5_n24, npu_inst_pe_1_1_5_n23,
         npu_inst_pe_1_1_5_n22, npu_inst_pe_1_1_5_n21, npu_inst_pe_1_1_5_n20,
         npu_inst_pe_1_1_5_n19, npu_inst_pe_1_1_5_n18, npu_inst_pe_1_1_5_n17,
         npu_inst_pe_1_1_5_n16, npu_inst_pe_1_1_5_n15, npu_inst_pe_1_1_5_n14,
         npu_inst_pe_1_1_5_n13, npu_inst_pe_1_1_5_n12, npu_inst_pe_1_1_5_n11,
         npu_inst_pe_1_1_5_n10, npu_inst_pe_1_1_5_n9, npu_inst_pe_1_1_5_n8,
         npu_inst_pe_1_1_5_n7, npu_inst_pe_1_1_5_n6, npu_inst_pe_1_1_5_n5,
         npu_inst_pe_1_1_5_n4, npu_inst_pe_1_1_5_n3, npu_inst_pe_1_1_5_n2,
         npu_inst_pe_1_1_5_n1, npu_inst_pe_1_1_5_sub_77_carry_7_,
         npu_inst_pe_1_1_5_sub_77_carry_6_, npu_inst_pe_1_1_5_sub_77_carry_5_,
         npu_inst_pe_1_1_5_sub_77_carry_4_, npu_inst_pe_1_1_5_sub_77_carry_3_,
         npu_inst_pe_1_1_5_sub_77_carry_2_, npu_inst_pe_1_1_5_sub_77_carry_1_,
         npu_inst_pe_1_1_5_add_79_carry_7_, npu_inst_pe_1_1_5_add_79_carry_6_,
         npu_inst_pe_1_1_5_add_79_carry_5_, npu_inst_pe_1_1_5_add_79_carry_4_,
         npu_inst_pe_1_1_5_add_79_carry_3_, npu_inst_pe_1_1_5_add_79_carry_2_,
         npu_inst_pe_1_1_5_add_79_carry_1_, npu_inst_pe_1_1_5_n97,
         npu_inst_pe_1_1_5_n96, npu_inst_pe_1_1_5_n95, npu_inst_pe_1_1_5_n94,
         npu_inst_pe_1_1_5_n93, npu_inst_pe_1_1_5_n92, npu_inst_pe_1_1_5_n91,
         npu_inst_pe_1_1_5_n90, npu_inst_pe_1_1_5_n89, npu_inst_pe_1_1_5_n88,
         npu_inst_pe_1_1_5_n87, npu_inst_pe_1_1_5_n86, npu_inst_pe_1_1_5_n85,
         npu_inst_pe_1_1_5_n84, npu_inst_pe_1_1_5_n83, npu_inst_pe_1_1_5_n82,
         npu_inst_pe_1_1_5_n81, npu_inst_pe_1_1_5_n80, npu_inst_pe_1_1_5_n79,
         npu_inst_pe_1_1_5_n78, npu_inst_pe_1_1_5_n77, npu_inst_pe_1_1_5_n76,
         npu_inst_pe_1_1_5_n75, npu_inst_pe_1_1_5_n74, npu_inst_pe_1_1_5_n73,
         npu_inst_pe_1_1_5_n72, npu_inst_pe_1_1_5_n71, npu_inst_pe_1_1_5_n70,
         npu_inst_pe_1_1_5_n69, npu_inst_pe_1_1_5_n68, npu_inst_pe_1_1_5_n67,
         npu_inst_pe_1_1_5_n66, npu_inst_pe_1_1_5_n65, npu_inst_pe_1_1_5_n64,
         npu_inst_pe_1_1_5_n63, npu_inst_pe_1_1_5_n62, npu_inst_pe_1_1_5_n61,
         npu_inst_pe_1_1_5_n60, npu_inst_pe_1_1_5_n59, npu_inst_pe_1_1_5_n58,
         npu_inst_pe_1_1_5_n57, npu_inst_pe_1_1_5_n56, npu_inst_pe_1_1_5_n55,
         npu_inst_pe_1_1_5_n54, npu_inst_pe_1_1_5_n53, npu_inst_pe_1_1_5_n52,
         npu_inst_pe_1_1_5_n51, npu_inst_pe_1_1_5_n50, npu_inst_pe_1_1_5_n49,
         npu_inst_pe_1_1_5_n48, npu_inst_pe_1_1_5_n47, npu_inst_pe_1_1_5_n46,
         npu_inst_pe_1_1_5_n45, npu_inst_pe_1_1_5_n44, npu_inst_pe_1_1_5_n43,
         npu_inst_pe_1_1_5_n42, npu_inst_pe_1_1_5_n41, npu_inst_pe_1_1_5_n40,
         npu_inst_pe_1_1_5_n39, npu_inst_pe_1_1_5_n38, npu_inst_pe_1_1_5_n37,
         npu_inst_pe_1_1_5_n27, npu_inst_pe_1_1_5_n26,
         npu_inst_pe_1_1_5_net4000, npu_inst_pe_1_1_5_net3994,
         npu_inst_pe_1_1_5_N94, npu_inst_pe_1_1_5_N93, npu_inst_pe_1_1_5_N84,
         npu_inst_pe_1_1_5_N80, npu_inst_pe_1_1_5_N79, npu_inst_pe_1_1_5_N78,
         npu_inst_pe_1_1_5_N77, npu_inst_pe_1_1_5_N76, npu_inst_pe_1_1_5_N75,
         npu_inst_pe_1_1_5_N74, npu_inst_pe_1_1_5_N73, npu_inst_pe_1_1_5_N72,
         npu_inst_pe_1_1_5_N71, npu_inst_pe_1_1_5_N70, npu_inst_pe_1_1_5_N69,
         npu_inst_pe_1_1_5_N68, npu_inst_pe_1_1_5_N67, npu_inst_pe_1_1_5_N66,
         npu_inst_pe_1_1_5_N65, npu_inst_pe_1_1_5_int_q_acc_0_,
         npu_inst_pe_1_1_5_int_q_acc_1_, npu_inst_pe_1_1_5_int_q_acc_2_,
         npu_inst_pe_1_1_5_int_q_acc_3_, npu_inst_pe_1_1_5_int_q_acc_4_,
         npu_inst_pe_1_1_5_int_q_acc_5_, npu_inst_pe_1_1_5_int_q_acc_6_,
         npu_inst_pe_1_1_5_int_q_acc_7_, npu_inst_pe_1_1_5_int_data_0_,
         npu_inst_pe_1_1_5_int_data_1_, npu_inst_pe_1_1_5_int_q_weight_0_,
         npu_inst_pe_1_1_5_int_q_weight_1_,
         npu_inst_pe_1_1_5_int_q_reg_v_5__0_,
         npu_inst_pe_1_1_5_int_q_reg_v_5__1_,
         npu_inst_pe_1_1_5_int_q_reg_v_4__0_,
         npu_inst_pe_1_1_5_int_q_reg_v_4__1_,
         npu_inst_pe_1_1_5_int_q_reg_v_3__0_,
         npu_inst_pe_1_1_5_int_q_reg_v_3__1_,
         npu_inst_pe_1_1_5_int_q_reg_v_2__0_,
         npu_inst_pe_1_1_5_int_q_reg_v_2__1_,
         npu_inst_pe_1_1_5_int_q_reg_v_1__0_,
         npu_inst_pe_1_1_5_int_q_reg_v_1__1_,
         npu_inst_pe_1_1_5_int_q_reg_v_0__0_,
         npu_inst_pe_1_1_5_int_q_reg_v_0__1_,
         npu_inst_pe_1_1_5_int_q_reg_h_5__0_,
         npu_inst_pe_1_1_5_int_q_reg_h_5__1_,
         npu_inst_pe_1_1_5_int_q_reg_h_4__0_,
         npu_inst_pe_1_1_5_int_q_reg_h_4__1_,
         npu_inst_pe_1_1_5_int_q_reg_h_3__0_,
         npu_inst_pe_1_1_5_int_q_reg_h_3__1_,
         npu_inst_pe_1_1_5_int_q_reg_h_2__0_,
         npu_inst_pe_1_1_5_int_q_reg_h_2__1_,
         npu_inst_pe_1_1_5_int_q_reg_h_1__0_,
         npu_inst_pe_1_1_5_int_q_reg_h_1__1_,
         npu_inst_pe_1_1_5_int_q_reg_h_0__0_,
         npu_inst_pe_1_1_5_int_q_reg_h_0__1_, npu_inst_pe_1_1_6_n119,
         npu_inst_pe_1_1_6_n118, npu_inst_pe_1_1_6_n117,
         npu_inst_pe_1_1_6_n116, npu_inst_pe_1_1_6_n115,
         npu_inst_pe_1_1_6_n114, npu_inst_pe_1_1_6_n113,
         npu_inst_pe_1_1_6_n112, npu_inst_pe_1_1_6_n111,
         npu_inst_pe_1_1_6_n110, npu_inst_pe_1_1_6_n109,
         npu_inst_pe_1_1_6_n108, npu_inst_pe_1_1_6_n107,
         npu_inst_pe_1_1_6_n106, npu_inst_pe_1_1_6_n105,
         npu_inst_pe_1_1_6_n104, npu_inst_pe_1_1_6_n103,
         npu_inst_pe_1_1_6_n102, npu_inst_pe_1_1_6_n101,
         npu_inst_pe_1_1_6_n100, npu_inst_pe_1_1_6_n99, npu_inst_pe_1_1_6_n98,
         npu_inst_pe_1_1_6_n36, npu_inst_pe_1_1_6_n35, npu_inst_pe_1_1_6_n34,
         npu_inst_pe_1_1_6_n33, npu_inst_pe_1_1_6_n32, npu_inst_pe_1_1_6_n31,
         npu_inst_pe_1_1_6_n30, npu_inst_pe_1_1_6_n29, npu_inst_pe_1_1_6_n28,
         npu_inst_pe_1_1_6_n25, npu_inst_pe_1_1_6_n24, npu_inst_pe_1_1_6_n23,
         npu_inst_pe_1_1_6_n22, npu_inst_pe_1_1_6_n21, npu_inst_pe_1_1_6_n20,
         npu_inst_pe_1_1_6_n19, npu_inst_pe_1_1_6_n18, npu_inst_pe_1_1_6_n17,
         npu_inst_pe_1_1_6_n16, npu_inst_pe_1_1_6_n15, npu_inst_pe_1_1_6_n14,
         npu_inst_pe_1_1_6_n13, npu_inst_pe_1_1_6_n12, npu_inst_pe_1_1_6_n11,
         npu_inst_pe_1_1_6_n10, npu_inst_pe_1_1_6_n9, npu_inst_pe_1_1_6_n8,
         npu_inst_pe_1_1_6_n7, npu_inst_pe_1_1_6_n6, npu_inst_pe_1_1_6_n5,
         npu_inst_pe_1_1_6_n4, npu_inst_pe_1_1_6_n3, npu_inst_pe_1_1_6_n2,
         npu_inst_pe_1_1_6_n1, npu_inst_pe_1_1_6_sub_77_carry_7_,
         npu_inst_pe_1_1_6_sub_77_carry_6_, npu_inst_pe_1_1_6_sub_77_carry_5_,
         npu_inst_pe_1_1_6_sub_77_carry_4_, npu_inst_pe_1_1_6_sub_77_carry_3_,
         npu_inst_pe_1_1_6_sub_77_carry_2_, npu_inst_pe_1_1_6_sub_77_carry_1_,
         npu_inst_pe_1_1_6_add_79_carry_7_, npu_inst_pe_1_1_6_add_79_carry_6_,
         npu_inst_pe_1_1_6_add_79_carry_5_, npu_inst_pe_1_1_6_add_79_carry_4_,
         npu_inst_pe_1_1_6_add_79_carry_3_, npu_inst_pe_1_1_6_add_79_carry_2_,
         npu_inst_pe_1_1_6_add_79_carry_1_, npu_inst_pe_1_1_6_n97,
         npu_inst_pe_1_1_6_n96, npu_inst_pe_1_1_6_n95, npu_inst_pe_1_1_6_n94,
         npu_inst_pe_1_1_6_n93, npu_inst_pe_1_1_6_n92, npu_inst_pe_1_1_6_n91,
         npu_inst_pe_1_1_6_n90, npu_inst_pe_1_1_6_n89, npu_inst_pe_1_1_6_n88,
         npu_inst_pe_1_1_6_n87, npu_inst_pe_1_1_6_n86, npu_inst_pe_1_1_6_n85,
         npu_inst_pe_1_1_6_n84, npu_inst_pe_1_1_6_n83, npu_inst_pe_1_1_6_n82,
         npu_inst_pe_1_1_6_n81, npu_inst_pe_1_1_6_n80, npu_inst_pe_1_1_6_n79,
         npu_inst_pe_1_1_6_n78, npu_inst_pe_1_1_6_n77, npu_inst_pe_1_1_6_n76,
         npu_inst_pe_1_1_6_n75, npu_inst_pe_1_1_6_n74, npu_inst_pe_1_1_6_n73,
         npu_inst_pe_1_1_6_n72, npu_inst_pe_1_1_6_n71, npu_inst_pe_1_1_6_n70,
         npu_inst_pe_1_1_6_n69, npu_inst_pe_1_1_6_n68, npu_inst_pe_1_1_6_n67,
         npu_inst_pe_1_1_6_n66, npu_inst_pe_1_1_6_n65, npu_inst_pe_1_1_6_n64,
         npu_inst_pe_1_1_6_n63, npu_inst_pe_1_1_6_n62, npu_inst_pe_1_1_6_n61,
         npu_inst_pe_1_1_6_n60, npu_inst_pe_1_1_6_n59, npu_inst_pe_1_1_6_n58,
         npu_inst_pe_1_1_6_n57, npu_inst_pe_1_1_6_n56, npu_inst_pe_1_1_6_n55,
         npu_inst_pe_1_1_6_n54, npu_inst_pe_1_1_6_n53, npu_inst_pe_1_1_6_n52,
         npu_inst_pe_1_1_6_n51, npu_inst_pe_1_1_6_n50, npu_inst_pe_1_1_6_n49,
         npu_inst_pe_1_1_6_n48, npu_inst_pe_1_1_6_n47, npu_inst_pe_1_1_6_n46,
         npu_inst_pe_1_1_6_n45, npu_inst_pe_1_1_6_n44, npu_inst_pe_1_1_6_n43,
         npu_inst_pe_1_1_6_n42, npu_inst_pe_1_1_6_n41, npu_inst_pe_1_1_6_n40,
         npu_inst_pe_1_1_6_n39, npu_inst_pe_1_1_6_n38, npu_inst_pe_1_1_6_n37,
         npu_inst_pe_1_1_6_n27, npu_inst_pe_1_1_6_n26,
         npu_inst_pe_1_1_6_net3977, npu_inst_pe_1_1_6_net3971,
         npu_inst_pe_1_1_6_N94, npu_inst_pe_1_1_6_N93, npu_inst_pe_1_1_6_N84,
         npu_inst_pe_1_1_6_N80, npu_inst_pe_1_1_6_N79, npu_inst_pe_1_1_6_N78,
         npu_inst_pe_1_1_6_N77, npu_inst_pe_1_1_6_N76, npu_inst_pe_1_1_6_N75,
         npu_inst_pe_1_1_6_N74, npu_inst_pe_1_1_6_N73, npu_inst_pe_1_1_6_N72,
         npu_inst_pe_1_1_6_N71, npu_inst_pe_1_1_6_N70, npu_inst_pe_1_1_6_N69,
         npu_inst_pe_1_1_6_N68, npu_inst_pe_1_1_6_N67, npu_inst_pe_1_1_6_N66,
         npu_inst_pe_1_1_6_N65, npu_inst_pe_1_1_6_int_q_acc_0_,
         npu_inst_pe_1_1_6_int_q_acc_1_, npu_inst_pe_1_1_6_int_q_acc_2_,
         npu_inst_pe_1_1_6_int_q_acc_3_, npu_inst_pe_1_1_6_int_q_acc_4_,
         npu_inst_pe_1_1_6_int_q_acc_5_, npu_inst_pe_1_1_6_int_q_acc_6_,
         npu_inst_pe_1_1_6_int_q_acc_7_, npu_inst_pe_1_1_6_int_data_0_,
         npu_inst_pe_1_1_6_int_data_1_, npu_inst_pe_1_1_6_int_q_weight_0_,
         npu_inst_pe_1_1_6_int_q_weight_1_,
         npu_inst_pe_1_1_6_int_q_reg_v_5__0_,
         npu_inst_pe_1_1_6_int_q_reg_v_5__1_,
         npu_inst_pe_1_1_6_int_q_reg_v_4__0_,
         npu_inst_pe_1_1_6_int_q_reg_v_4__1_,
         npu_inst_pe_1_1_6_int_q_reg_v_3__0_,
         npu_inst_pe_1_1_6_int_q_reg_v_3__1_,
         npu_inst_pe_1_1_6_int_q_reg_v_2__0_,
         npu_inst_pe_1_1_6_int_q_reg_v_2__1_,
         npu_inst_pe_1_1_6_int_q_reg_v_1__0_,
         npu_inst_pe_1_1_6_int_q_reg_v_1__1_,
         npu_inst_pe_1_1_6_int_q_reg_v_0__0_,
         npu_inst_pe_1_1_6_int_q_reg_v_0__1_,
         npu_inst_pe_1_1_6_int_q_reg_h_5__0_,
         npu_inst_pe_1_1_6_int_q_reg_h_5__1_,
         npu_inst_pe_1_1_6_int_q_reg_h_4__0_,
         npu_inst_pe_1_1_6_int_q_reg_h_4__1_,
         npu_inst_pe_1_1_6_int_q_reg_h_3__0_,
         npu_inst_pe_1_1_6_int_q_reg_h_3__1_,
         npu_inst_pe_1_1_6_int_q_reg_h_2__0_,
         npu_inst_pe_1_1_6_int_q_reg_h_2__1_,
         npu_inst_pe_1_1_6_int_q_reg_h_1__0_,
         npu_inst_pe_1_1_6_int_q_reg_h_1__1_,
         npu_inst_pe_1_1_6_int_q_reg_h_0__0_,
         npu_inst_pe_1_1_6_int_q_reg_h_0__1_, npu_inst_pe_1_1_7_n119,
         npu_inst_pe_1_1_7_n118, npu_inst_pe_1_1_7_n117,
         npu_inst_pe_1_1_7_n116, npu_inst_pe_1_1_7_n115,
         npu_inst_pe_1_1_7_n114, npu_inst_pe_1_1_7_n113,
         npu_inst_pe_1_1_7_n112, npu_inst_pe_1_1_7_n111,
         npu_inst_pe_1_1_7_n110, npu_inst_pe_1_1_7_n109,
         npu_inst_pe_1_1_7_n108, npu_inst_pe_1_1_7_n107,
         npu_inst_pe_1_1_7_n106, npu_inst_pe_1_1_7_n105,
         npu_inst_pe_1_1_7_n104, npu_inst_pe_1_1_7_n103,
         npu_inst_pe_1_1_7_n102, npu_inst_pe_1_1_7_n101,
         npu_inst_pe_1_1_7_n100, npu_inst_pe_1_1_7_n99, npu_inst_pe_1_1_7_n98,
         npu_inst_pe_1_1_7_n36, npu_inst_pe_1_1_7_n35, npu_inst_pe_1_1_7_n34,
         npu_inst_pe_1_1_7_n33, npu_inst_pe_1_1_7_n32, npu_inst_pe_1_1_7_n31,
         npu_inst_pe_1_1_7_n30, npu_inst_pe_1_1_7_n29, npu_inst_pe_1_1_7_n28,
         npu_inst_pe_1_1_7_n25, npu_inst_pe_1_1_7_n24, npu_inst_pe_1_1_7_n23,
         npu_inst_pe_1_1_7_n22, npu_inst_pe_1_1_7_n21, npu_inst_pe_1_1_7_n20,
         npu_inst_pe_1_1_7_n19, npu_inst_pe_1_1_7_n18, npu_inst_pe_1_1_7_n17,
         npu_inst_pe_1_1_7_n16, npu_inst_pe_1_1_7_n15, npu_inst_pe_1_1_7_n14,
         npu_inst_pe_1_1_7_n13, npu_inst_pe_1_1_7_n12, npu_inst_pe_1_1_7_n11,
         npu_inst_pe_1_1_7_n10, npu_inst_pe_1_1_7_n9, npu_inst_pe_1_1_7_n8,
         npu_inst_pe_1_1_7_n7, npu_inst_pe_1_1_7_n6, npu_inst_pe_1_1_7_n5,
         npu_inst_pe_1_1_7_n4, npu_inst_pe_1_1_7_n3, npu_inst_pe_1_1_7_n2,
         npu_inst_pe_1_1_7_n1, npu_inst_pe_1_1_7_sub_77_carry_7_,
         npu_inst_pe_1_1_7_sub_77_carry_6_, npu_inst_pe_1_1_7_sub_77_carry_5_,
         npu_inst_pe_1_1_7_sub_77_carry_4_, npu_inst_pe_1_1_7_sub_77_carry_3_,
         npu_inst_pe_1_1_7_sub_77_carry_2_, npu_inst_pe_1_1_7_sub_77_carry_1_,
         npu_inst_pe_1_1_7_add_79_carry_7_, npu_inst_pe_1_1_7_add_79_carry_6_,
         npu_inst_pe_1_1_7_add_79_carry_5_, npu_inst_pe_1_1_7_add_79_carry_4_,
         npu_inst_pe_1_1_7_add_79_carry_3_, npu_inst_pe_1_1_7_add_79_carry_2_,
         npu_inst_pe_1_1_7_add_79_carry_1_, npu_inst_pe_1_1_7_n97,
         npu_inst_pe_1_1_7_n96, npu_inst_pe_1_1_7_n95, npu_inst_pe_1_1_7_n94,
         npu_inst_pe_1_1_7_n93, npu_inst_pe_1_1_7_n92, npu_inst_pe_1_1_7_n91,
         npu_inst_pe_1_1_7_n90, npu_inst_pe_1_1_7_n89, npu_inst_pe_1_1_7_n88,
         npu_inst_pe_1_1_7_n87, npu_inst_pe_1_1_7_n86, npu_inst_pe_1_1_7_n85,
         npu_inst_pe_1_1_7_n84, npu_inst_pe_1_1_7_n83, npu_inst_pe_1_1_7_n82,
         npu_inst_pe_1_1_7_n81, npu_inst_pe_1_1_7_n80, npu_inst_pe_1_1_7_n79,
         npu_inst_pe_1_1_7_n78, npu_inst_pe_1_1_7_n77, npu_inst_pe_1_1_7_n76,
         npu_inst_pe_1_1_7_n75, npu_inst_pe_1_1_7_n74, npu_inst_pe_1_1_7_n73,
         npu_inst_pe_1_1_7_n72, npu_inst_pe_1_1_7_n71, npu_inst_pe_1_1_7_n70,
         npu_inst_pe_1_1_7_n69, npu_inst_pe_1_1_7_n68, npu_inst_pe_1_1_7_n67,
         npu_inst_pe_1_1_7_n66, npu_inst_pe_1_1_7_n65, npu_inst_pe_1_1_7_n64,
         npu_inst_pe_1_1_7_n63, npu_inst_pe_1_1_7_n62, npu_inst_pe_1_1_7_n61,
         npu_inst_pe_1_1_7_n60, npu_inst_pe_1_1_7_n59, npu_inst_pe_1_1_7_n58,
         npu_inst_pe_1_1_7_n57, npu_inst_pe_1_1_7_n56, npu_inst_pe_1_1_7_n55,
         npu_inst_pe_1_1_7_n54, npu_inst_pe_1_1_7_n53, npu_inst_pe_1_1_7_n52,
         npu_inst_pe_1_1_7_n51, npu_inst_pe_1_1_7_n50, npu_inst_pe_1_1_7_n49,
         npu_inst_pe_1_1_7_n48, npu_inst_pe_1_1_7_n47, npu_inst_pe_1_1_7_n46,
         npu_inst_pe_1_1_7_n45, npu_inst_pe_1_1_7_n44, npu_inst_pe_1_1_7_n43,
         npu_inst_pe_1_1_7_n42, npu_inst_pe_1_1_7_n41, npu_inst_pe_1_1_7_n40,
         npu_inst_pe_1_1_7_n39, npu_inst_pe_1_1_7_n38, npu_inst_pe_1_1_7_n37,
         npu_inst_pe_1_1_7_n27, npu_inst_pe_1_1_7_n26,
         npu_inst_pe_1_1_7_net3954, npu_inst_pe_1_1_7_net3948,
         npu_inst_pe_1_1_7_N94, npu_inst_pe_1_1_7_N93, npu_inst_pe_1_1_7_N84,
         npu_inst_pe_1_1_7_N80, npu_inst_pe_1_1_7_N79, npu_inst_pe_1_1_7_N78,
         npu_inst_pe_1_1_7_N77, npu_inst_pe_1_1_7_N76, npu_inst_pe_1_1_7_N75,
         npu_inst_pe_1_1_7_N74, npu_inst_pe_1_1_7_N73, npu_inst_pe_1_1_7_N72,
         npu_inst_pe_1_1_7_N71, npu_inst_pe_1_1_7_N70, npu_inst_pe_1_1_7_N69,
         npu_inst_pe_1_1_7_N68, npu_inst_pe_1_1_7_N67, npu_inst_pe_1_1_7_N66,
         npu_inst_pe_1_1_7_N65, npu_inst_pe_1_1_7_int_q_acc_0_,
         npu_inst_pe_1_1_7_int_q_acc_1_, npu_inst_pe_1_1_7_int_q_acc_2_,
         npu_inst_pe_1_1_7_int_q_acc_3_, npu_inst_pe_1_1_7_int_q_acc_4_,
         npu_inst_pe_1_1_7_int_q_acc_5_, npu_inst_pe_1_1_7_int_q_acc_6_,
         npu_inst_pe_1_1_7_int_q_acc_7_, npu_inst_pe_1_1_7_int_data_0_,
         npu_inst_pe_1_1_7_int_data_1_, npu_inst_pe_1_1_7_int_q_weight_0_,
         npu_inst_pe_1_1_7_int_q_weight_1_,
         npu_inst_pe_1_1_7_int_q_reg_v_5__0_,
         npu_inst_pe_1_1_7_int_q_reg_v_5__1_,
         npu_inst_pe_1_1_7_int_q_reg_v_4__0_,
         npu_inst_pe_1_1_7_int_q_reg_v_4__1_,
         npu_inst_pe_1_1_7_int_q_reg_v_3__0_,
         npu_inst_pe_1_1_7_int_q_reg_v_3__1_,
         npu_inst_pe_1_1_7_int_q_reg_v_2__0_,
         npu_inst_pe_1_1_7_int_q_reg_v_2__1_,
         npu_inst_pe_1_1_7_int_q_reg_v_1__0_,
         npu_inst_pe_1_1_7_int_q_reg_v_1__1_,
         npu_inst_pe_1_1_7_int_q_reg_v_0__0_,
         npu_inst_pe_1_1_7_int_q_reg_v_0__1_,
         npu_inst_pe_1_1_7_int_q_reg_h_5__0_,
         npu_inst_pe_1_1_7_int_q_reg_h_5__1_,
         npu_inst_pe_1_1_7_int_q_reg_h_4__0_,
         npu_inst_pe_1_1_7_int_q_reg_h_4__1_,
         npu_inst_pe_1_1_7_int_q_reg_h_3__0_,
         npu_inst_pe_1_1_7_int_q_reg_h_3__1_,
         npu_inst_pe_1_1_7_int_q_reg_h_2__0_,
         npu_inst_pe_1_1_7_int_q_reg_h_2__1_,
         npu_inst_pe_1_1_7_int_q_reg_h_1__0_,
         npu_inst_pe_1_1_7_int_q_reg_h_1__1_,
         npu_inst_pe_1_1_7_int_q_reg_h_0__0_,
         npu_inst_pe_1_1_7_int_q_reg_h_0__1_, npu_inst_pe_1_2_0_n118,
         npu_inst_pe_1_2_0_n117, npu_inst_pe_1_2_0_n116,
         npu_inst_pe_1_2_0_n115, npu_inst_pe_1_2_0_n114,
         npu_inst_pe_1_2_0_n113, npu_inst_pe_1_2_0_n112,
         npu_inst_pe_1_2_0_n111, npu_inst_pe_1_2_0_n110,
         npu_inst_pe_1_2_0_n109, npu_inst_pe_1_2_0_n108,
         npu_inst_pe_1_2_0_n107, npu_inst_pe_1_2_0_n106,
         npu_inst_pe_1_2_0_n105, npu_inst_pe_1_2_0_n104,
         npu_inst_pe_1_2_0_n103, npu_inst_pe_1_2_0_n102,
         npu_inst_pe_1_2_0_n101, npu_inst_pe_1_2_0_n100, npu_inst_pe_1_2_0_n99,
         npu_inst_pe_1_2_0_n98, npu_inst_pe_1_2_0_n36, npu_inst_pe_1_2_0_n35,
         npu_inst_pe_1_2_0_n34, npu_inst_pe_1_2_0_n33, npu_inst_pe_1_2_0_n32,
         npu_inst_pe_1_2_0_n31, npu_inst_pe_1_2_0_n30, npu_inst_pe_1_2_0_n29,
         npu_inst_pe_1_2_0_n28, npu_inst_pe_1_2_0_n25, npu_inst_pe_1_2_0_n24,
         npu_inst_pe_1_2_0_n23, npu_inst_pe_1_2_0_n22, npu_inst_pe_1_2_0_n21,
         npu_inst_pe_1_2_0_n20, npu_inst_pe_1_2_0_n19, npu_inst_pe_1_2_0_n18,
         npu_inst_pe_1_2_0_n17, npu_inst_pe_1_2_0_n16, npu_inst_pe_1_2_0_n15,
         npu_inst_pe_1_2_0_n14, npu_inst_pe_1_2_0_n13, npu_inst_pe_1_2_0_n12,
         npu_inst_pe_1_2_0_n11, npu_inst_pe_1_2_0_n10, npu_inst_pe_1_2_0_n9,
         npu_inst_pe_1_2_0_n8, npu_inst_pe_1_2_0_n7, npu_inst_pe_1_2_0_n6,
         npu_inst_pe_1_2_0_n5, npu_inst_pe_1_2_0_n4, npu_inst_pe_1_2_0_n3,
         npu_inst_pe_1_2_0_n2, npu_inst_pe_1_2_0_n1,
         npu_inst_pe_1_2_0_sub_77_carry_7_, npu_inst_pe_1_2_0_sub_77_carry_6_,
         npu_inst_pe_1_2_0_sub_77_carry_5_, npu_inst_pe_1_2_0_sub_77_carry_4_,
         npu_inst_pe_1_2_0_sub_77_carry_3_, npu_inst_pe_1_2_0_sub_77_carry_2_,
         npu_inst_pe_1_2_0_sub_77_carry_1_, npu_inst_pe_1_2_0_add_79_carry_7_,
         npu_inst_pe_1_2_0_add_79_carry_6_, npu_inst_pe_1_2_0_add_79_carry_5_,
         npu_inst_pe_1_2_0_add_79_carry_4_, npu_inst_pe_1_2_0_add_79_carry_3_,
         npu_inst_pe_1_2_0_add_79_carry_2_, npu_inst_pe_1_2_0_add_79_carry_1_,
         npu_inst_pe_1_2_0_n97, npu_inst_pe_1_2_0_n96, npu_inst_pe_1_2_0_n95,
         npu_inst_pe_1_2_0_n94, npu_inst_pe_1_2_0_n93, npu_inst_pe_1_2_0_n92,
         npu_inst_pe_1_2_0_n91, npu_inst_pe_1_2_0_n90, npu_inst_pe_1_2_0_n89,
         npu_inst_pe_1_2_0_n88, npu_inst_pe_1_2_0_n87, npu_inst_pe_1_2_0_n86,
         npu_inst_pe_1_2_0_n85, npu_inst_pe_1_2_0_n84, npu_inst_pe_1_2_0_n83,
         npu_inst_pe_1_2_0_n82, npu_inst_pe_1_2_0_n81, npu_inst_pe_1_2_0_n80,
         npu_inst_pe_1_2_0_n79, npu_inst_pe_1_2_0_n78, npu_inst_pe_1_2_0_n77,
         npu_inst_pe_1_2_0_n76, npu_inst_pe_1_2_0_n75, npu_inst_pe_1_2_0_n74,
         npu_inst_pe_1_2_0_n73, npu_inst_pe_1_2_0_n72, npu_inst_pe_1_2_0_n71,
         npu_inst_pe_1_2_0_n70, npu_inst_pe_1_2_0_n69, npu_inst_pe_1_2_0_n68,
         npu_inst_pe_1_2_0_n67, npu_inst_pe_1_2_0_n66, npu_inst_pe_1_2_0_n65,
         npu_inst_pe_1_2_0_n64, npu_inst_pe_1_2_0_n63, npu_inst_pe_1_2_0_n62,
         npu_inst_pe_1_2_0_n61, npu_inst_pe_1_2_0_n60, npu_inst_pe_1_2_0_n59,
         npu_inst_pe_1_2_0_n58, npu_inst_pe_1_2_0_n57, npu_inst_pe_1_2_0_n56,
         npu_inst_pe_1_2_0_n55, npu_inst_pe_1_2_0_n54, npu_inst_pe_1_2_0_n53,
         npu_inst_pe_1_2_0_n52, npu_inst_pe_1_2_0_n51, npu_inst_pe_1_2_0_n50,
         npu_inst_pe_1_2_0_n49, npu_inst_pe_1_2_0_n48, npu_inst_pe_1_2_0_n47,
         npu_inst_pe_1_2_0_n46, npu_inst_pe_1_2_0_n45, npu_inst_pe_1_2_0_n44,
         npu_inst_pe_1_2_0_n43, npu_inst_pe_1_2_0_n42, npu_inst_pe_1_2_0_n41,
         npu_inst_pe_1_2_0_n40, npu_inst_pe_1_2_0_n39, npu_inst_pe_1_2_0_n38,
         npu_inst_pe_1_2_0_n37, npu_inst_pe_1_2_0_n27, npu_inst_pe_1_2_0_n26,
         npu_inst_pe_1_2_0_net3931, npu_inst_pe_1_2_0_net3925,
         npu_inst_pe_1_2_0_N94, npu_inst_pe_1_2_0_N93, npu_inst_pe_1_2_0_N84,
         npu_inst_pe_1_2_0_N80, npu_inst_pe_1_2_0_N79, npu_inst_pe_1_2_0_N78,
         npu_inst_pe_1_2_0_N77, npu_inst_pe_1_2_0_N76, npu_inst_pe_1_2_0_N75,
         npu_inst_pe_1_2_0_N74, npu_inst_pe_1_2_0_N73, npu_inst_pe_1_2_0_N72,
         npu_inst_pe_1_2_0_N71, npu_inst_pe_1_2_0_N70, npu_inst_pe_1_2_0_N69,
         npu_inst_pe_1_2_0_N68, npu_inst_pe_1_2_0_N67, npu_inst_pe_1_2_0_N66,
         npu_inst_pe_1_2_0_N65, npu_inst_pe_1_2_0_int_q_acc_0_,
         npu_inst_pe_1_2_0_int_q_acc_1_, npu_inst_pe_1_2_0_int_q_acc_2_,
         npu_inst_pe_1_2_0_int_q_acc_3_, npu_inst_pe_1_2_0_int_q_acc_4_,
         npu_inst_pe_1_2_0_int_q_acc_5_, npu_inst_pe_1_2_0_int_q_acc_6_,
         npu_inst_pe_1_2_0_int_q_acc_7_, npu_inst_pe_1_2_0_int_data_0_,
         npu_inst_pe_1_2_0_int_data_1_, npu_inst_pe_1_2_0_int_q_weight_0_,
         npu_inst_pe_1_2_0_int_q_weight_1_,
         npu_inst_pe_1_2_0_int_q_reg_v_5__0_,
         npu_inst_pe_1_2_0_int_q_reg_v_5__1_,
         npu_inst_pe_1_2_0_int_q_reg_v_4__0_,
         npu_inst_pe_1_2_0_int_q_reg_v_4__1_,
         npu_inst_pe_1_2_0_int_q_reg_v_3__0_,
         npu_inst_pe_1_2_0_int_q_reg_v_3__1_,
         npu_inst_pe_1_2_0_int_q_reg_v_2__0_,
         npu_inst_pe_1_2_0_int_q_reg_v_2__1_,
         npu_inst_pe_1_2_0_int_q_reg_v_1__0_,
         npu_inst_pe_1_2_0_int_q_reg_v_1__1_,
         npu_inst_pe_1_2_0_int_q_reg_v_0__0_,
         npu_inst_pe_1_2_0_int_q_reg_v_0__1_,
         npu_inst_pe_1_2_0_int_q_reg_h_5__0_,
         npu_inst_pe_1_2_0_int_q_reg_h_5__1_,
         npu_inst_pe_1_2_0_int_q_reg_h_4__0_,
         npu_inst_pe_1_2_0_int_q_reg_h_4__1_,
         npu_inst_pe_1_2_0_int_q_reg_h_3__0_,
         npu_inst_pe_1_2_0_int_q_reg_h_3__1_,
         npu_inst_pe_1_2_0_int_q_reg_h_2__0_,
         npu_inst_pe_1_2_0_int_q_reg_h_2__1_,
         npu_inst_pe_1_2_0_int_q_reg_h_1__0_,
         npu_inst_pe_1_2_0_int_q_reg_h_1__1_,
         npu_inst_pe_1_2_0_int_q_reg_h_0__0_,
         npu_inst_pe_1_2_0_int_q_reg_h_0__1_, npu_inst_pe_1_2_0_o_data_h_0_,
         npu_inst_pe_1_2_0_o_data_h_1_, npu_inst_pe_1_2_1_n119,
         npu_inst_pe_1_2_1_n118, npu_inst_pe_1_2_1_n117,
         npu_inst_pe_1_2_1_n116, npu_inst_pe_1_2_1_n115,
         npu_inst_pe_1_2_1_n114, npu_inst_pe_1_2_1_n113,
         npu_inst_pe_1_2_1_n112, npu_inst_pe_1_2_1_n111,
         npu_inst_pe_1_2_1_n110, npu_inst_pe_1_2_1_n109,
         npu_inst_pe_1_2_1_n108, npu_inst_pe_1_2_1_n107,
         npu_inst_pe_1_2_1_n106, npu_inst_pe_1_2_1_n105,
         npu_inst_pe_1_2_1_n104, npu_inst_pe_1_2_1_n103,
         npu_inst_pe_1_2_1_n102, npu_inst_pe_1_2_1_n101,
         npu_inst_pe_1_2_1_n100, npu_inst_pe_1_2_1_n99, npu_inst_pe_1_2_1_n98,
         npu_inst_pe_1_2_1_n36, npu_inst_pe_1_2_1_n35, npu_inst_pe_1_2_1_n34,
         npu_inst_pe_1_2_1_n33, npu_inst_pe_1_2_1_n32, npu_inst_pe_1_2_1_n31,
         npu_inst_pe_1_2_1_n30, npu_inst_pe_1_2_1_n29, npu_inst_pe_1_2_1_n28,
         npu_inst_pe_1_2_1_n25, npu_inst_pe_1_2_1_n24, npu_inst_pe_1_2_1_n23,
         npu_inst_pe_1_2_1_n22, npu_inst_pe_1_2_1_n21, npu_inst_pe_1_2_1_n20,
         npu_inst_pe_1_2_1_n19, npu_inst_pe_1_2_1_n18, npu_inst_pe_1_2_1_n17,
         npu_inst_pe_1_2_1_n16, npu_inst_pe_1_2_1_n15, npu_inst_pe_1_2_1_n14,
         npu_inst_pe_1_2_1_n13, npu_inst_pe_1_2_1_n12, npu_inst_pe_1_2_1_n11,
         npu_inst_pe_1_2_1_n10, npu_inst_pe_1_2_1_n9, npu_inst_pe_1_2_1_n8,
         npu_inst_pe_1_2_1_n7, npu_inst_pe_1_2_1_n6, npu_inst_pe_1_2_1_n5,
         npu_inst_pe_1_2_1_n4, npu_inst_pe_1_2_1_n3, npu_inst_pe_1_2_1_n2,
         npu_inst_pe_1_2_1_n1, npu_inst_pe_1_2_1_sub_77_carry_7_,
         npu_inst_pe_1_2_1_sub_77_carry_6_, npu_inst_pe_1_2_1_sub_77_carry_5_,
         npu_inst_pe_1_2_1_sub_77_carry_4_, npu_inst_pe_1_2_1_sub_77_carry_3_,
         npu_inst_pe_1_2_1_sub_77_carry_2_, npu_inst_pe_1_2_1_sub_77_carry_1_,
         npu_inst_pe_1_2_1_add_79_carry_7_, npu_inst_pe_1_2_1_add_79_carry_6_,
         npu_inst_pe_1_2_1_add_79_carry_5_, npu_inst_pe_1_2_1_add_79_carry_4_,
         npu_inst_pe_1_2_1_add_79_carry_3_, npu_inst_pe_1_2_1_add_79_carry_2_,
         npu_inst_pe_1_2_1_add_79_carry_1_, npu_inst_pe_1_2_1_n97,
         npu_inst_pe_1_2_1_n96, npu_inst_pe_1_2_1_n95, npu_inst_pe_1_2_1_n94,
         npu_inst_pe_1_2_1_n93, npu_inst_pe_1_2_1_n92, npu_inst_pe_1_2_1_n91,
         npu_inst_pe_1_2_1_n90, npu_inst_pe_1_2_1_n89, npu_inst_pe_1_2_1_n88,
         npu_inst_pe_1_2_1_n87, npu_inst_pe_1_2_1_n86, npu_inst_pe_1_2_1_n85,
         npu_inst_pe_1_2_1_n84, npu_inst_pe_1_2_1_n83, npu_inst_pe_1_2_1_n82,
         npu_inst_pe_1_2_1_n81, npu_inst_pe_1_2_1_n80, npu_inst_pe_1_2_1_n79,
         npu_inst_pe_1_2_1_n78, npu_inst_pe_1_2_1_n77, npu_inst_pe_1_2_1_n76,
         npu_inst_pe_1_2_1_n75, npu_inst_pe_1_2_1_n74, npu_inst_pe_1_2_1_n73,
         npu_inst_pe_1_2_1_n72, npu_inst_pe_1_2_1_n71, npu_inst_pe_1_2_1_n70,
         npu_inst_pe_1_2_1_n69, npu_inst_pe_1_2_1_n68, npu_inst_pe_1_2_1_n67,
         npu_inst_pe_1_2_1_n66, npu_inst_pe_1_2_1_n65, npu_inst_pe_1_2_1_n64,
         npu_inst_pe_1_2_1_n63, npu_inst_pe_1_2_1_n62, npu_inst_pe_1_2_1_n61,
         npu_inst_pe_1_2_1_n60, npu_inst_pe_1_2_1_n59, npu_inst_pe_1_2_1_n58,
         npu_inst_pe_1_2_1_n57, npu_inst_pe_1_2_1_n56, npu_inst_pe_1_2_1_n55,
         npu_inst_pe_1_2_1_n54, npu_inst_pe_1_2_1_n53, npu_inst_pe_1_2_1_n52,
         npu_inst_pe_1_2_1_n51, npu_inst_pe_1_2_1_n50, npu_inst_pe_1_2_1_n49,
         npu_inst_pe_1_2_1_n48, npu_inst_pe_1_2_1_n47, npu_inst_pe_1_2_1_n46,
         npu_inst_pe_1_2_1_n45, npu_inst_pe_1_2_1_n44, npu_inst_pe_1_2_1_n43,
         npu_inst_pe_1_2_1_n42, npu_inst_pe_1_2_1_n41, npu_inst_pe_1_2_1_n40,
         npu_inst_pe_1_2_1_n39, npu_inst_pe_1_2_1_n38, npu_inst_pe_1_2_1_n37,
         npu_inst_pe_1_2_1_n27, npu_inst_pe_1_2_1_n26,
         npu_inst_pe_1_2_1_net3908, npu_inst_pe_1_2_1_net3902,
         npu_inst_pe_1_2_1_N94, npu_inst_pe_1_2_1_N93, npu_inst_pe_1_2_1_N84,
         npu_inst_pe_1_2_1_N80, npu_inst_pe_1_2_1_N79, npu_inst_pe_1_2_1_N78,
         npu_inst_pe_1_2_1_N77, npu_inst_pe_1_2_1_N76, npu_inst_pe_1_2_1_N75,
         npu_inst_pe_1_2_1_N74, npu_inst_pe_1_2_1_N73, npu_inst_pe_1_2_1_N72,
         npu_inst_pe_1_2_1_N71, npu_inst_pe_1_2_1_N70, npu_inst_pe_1_2_1_N69,
         npu_inst_pe_1_2_1_N68, npu_inst_pe_1_2_1_N67, npu_inst_pe_1_2_1_N66,
         npu_inst_pe_1_2_1_N65, npu_inst_pe_1_2_1_int_q_acc_0_,
         npu_inst_pe_1_2_1_int_q_acc_1_, npu_inst_pe_1_2_1_int_q_acc_2_,
         npu_inst_pe_1_2_1_int_q_acc_3_, npu_inst_pe_1_2_1_int_q_acc_4_,
         npu_inst_pe_1_2_1_int_q_acc_5_, npu_inst_pe_1_2_1_int_q_acc_6_,
         npu_inst_pe_1_2_1_int_q_acc_7_, npu_inst_pe_1_2_1_int_data_0_,
         npu_inst_pe_1_2_1_int_data_1_, npu_inst_pe_1_2_1_int_q_weight_0_,
         npu_inst_pe_1_2_1_int_q_weight_1_,
         npu_inst_pe_1_2_1_int_q_reg_v_5__0_,
         npu_inst_pe_1_2_1_int_q_reg_v_5__1_,
         npu_inst_pe_1_2_1_int_q_reg_v_4__0_,
         npu_inst_pe_1_2_1_int_q_reg_v_4__1_,
         npu_inst_pe_1_2_1_int_q_reg_v_3__0_,
         npu_inst_pe_1_2_1_int_q_reg_v_3__1_,
         npu_inst_pe_1_2_1_int_q_reg_v_2__0_,
         npu_inst_pe_1_2_1_int_q_reg_v_2__1_,
         npu_inst_pe_1_2_1_int_q_reg_v_1__0_,
         npu_inst_pe_1_2_1_int_q_reg_v_1__1_,
         npu_inst_pe_1_2_1_int_q_reg_v_0__0_,
         npu_inst_pe_1_2_1_int_q_reg_v_0__1_,
         npu_inst_pe_1_2_1_int_q_reg_h_5__0_,
         npu_inst_pe_1_2_1_int_q_reg_h_5__1_,
         npu_inst_pe_1_2_1_int_q_reg_h_4__0_,
         npu_inst_pe_1_2_1_int_q_reg_h_4__1_,
         npu_inst_pe_1_2_1_int_q_reg_h_3__0_,
         npu_inst_pe_1_2_1_int_q_reg_h_3__1_,
         npu_inst_pe_1_2_1_int_q_reg_h_2__0_,
         npu_inst_pe_1_2_1_int_q_reg_h_2__1_,
         npu_inst_pe_1_2_1_int_q_reg_h_1__0_,
         npu_inst_pe_1_2_1_int_q_reg_h_1__1_,
         npu_inst_pe_1_2_1_int_q_reg_h_0__0_,
         npu_inst_pe_1_2_1_int_q_reg_h_0__1_, npu_inst_pe_1_2_2_n119,
         npu_inst_pe_1_2_2_n118, npu_inst_pe_1_2_2_n117,
         npu_inst_pe_1_2_2_n116, npu_inst_pe_1_2_2_n115,
         npu_inst_pe_1_2_2_n114, npu_inst_pe_1_2_2_n113,
         npu_inst_pe_1_2_2_n112, npu_inst_pe_1_2_2_n111,
         npu_inst_pe_1_2_2_n110, npu_inst_pe_1_2_2_n109,
         npu_inst_pe_1_2_2_n108, npu_inst_pe_1_2_2_n107,
         npu_inst_pe_1_2_2_n106, npu_inst_pe_1_2_2_n105,
         npu_inst_pe_1_2_2_n104, npu_inst_pe_1_2_2_n103,
         npu_inst_pe_1_2_2_n102, npu_inst_pe_1_2_2_n101,
         npu_inst_pe_1_2_2_n100, npu_inst_pe_1_2_2_n99, npu_inst_pe_1_2_2_n98,
         npu_inst_pe_1_2_2_n36, npu_inst_pe_1_2_2_n35, npu_inst_pe_1_2_2_n34,
         npu_inst_pe_1_2_2_n33, npu_inst_pe_1_2_2_n32, npu_inst_pe_1_2_2_n31,
         npu_inst_pe_1_2_2_n30, npu_inst_pe_1_2_2_n29, npu_inst_pe_1_2_2_n28,
         npu_inst_pe_1_2_2_n25, npu_inst_pe_1_2_2_n24, npu_inst_pe_1_2_2_n23,
         npu_inst_pe_1_2_2_n22, npu_inst_pe_1_2_2_n21, npu_inst_pe_1_2_2_n20,
         npu_inst_pe_1_2_2_n19, npu_inst_pe_1_2_2_n18, npu_inst_pe_1_2_2_n17,
         npu_inst_pe_1_2_2_n16, npu_inst_pe_1_2_2_n15, npu_inst_pe_1_2_2_n14,
         npu_inst_pe_1_2_2_n13, npu_inst_pe_1_2_2_n12, npu_inst_pe_1_2_2_n11,
         npu_inst_pe_1_2_2_n10, npu_inst_pe_1_2_2_n9, npu_inst_pe_1_2_2_n8,
         npu_inst_pe_1_2_2_n7, npu_inst_pe_1_2_2_n6, npu_inst_pe_1_2_2_n5,
         npu_inst_pe_1_2_2_n4, npu_inst_pe_1_2_2_n3, npu_inst_pe_1_2_2_n2,
         npu_inst_pe_1_2_2_n1, npu_inst_pe_1_2_2_sub_77_carry_7_,
         npu_inst_pe_1_2_2_sub_77_carry_6_, npu_inst_pe_1_2_2_sub_77_carry_5_,
         npu_inst_pe_1_2_2_sub_77_carry_4_, npu_inst_pe_1_2_2_sub_77_carry_3_,
         npu_inst_pe_1_2_2_sub_77_carry_2_, npu_inst_pe_1_2_2_sub_77_carry_1_,
         npu_inst_pe_1_2_2_add_79_carry_7_, npu_inst_pe_1_2_2_add_79_carry_6_,
         npu_inst_pe_1_2_2_add_79_carry_5_, npu_inst_pe_1_2_2_add_79_carry_4_,
         npu_inst_pe_1_2_2_add_79_carry_3_, npu_inst_pe_1_2_2_add_79_carry_2_,
         npu_inst_pe_1_2_2_add_79_carry_1_, npu_inst_pe_1_2_2_n97,
         npu_inst_pe_1_2_2_n96, npu_inst_pe_1_2_2_n95, npu_inst_pe_1_2_2_n94,
         npu_inst_pe_1_2_2_n93, npu_inst_pe_1_2_2_n92, npu_inst_pe_1_2_2_n91,
         npu_inst_pe_1_2_2_n90, npu_inst_pe_1_2_2_n89, npu_inst_pe_1_2_2_n88,
         npu_inst_pe_1_2_2_n87, npu_inst_pe_1_2_2_n86, npu_inst_pe_1_2_2_n85,
         npu_inst_pe_1_2_2_n84, npu_inst_pe_1_2_2_n83, npu_inst_pe_1_2_2_n82,
         npu_inst_pe_1_2_2_n81, npu_inst_pe_1_2_2_n80, npu_inst_pe_1_2_2_n79,
         npu_inst_pe_1_2_2_n78, npu_inst_pe_1_2_2_n77, npu_inst_pe_1_2_2_n76,
         npu_inst_pe_1_2_2_n75, npu_inst_pe_1_2_2_n74, npu_inst_pe_1_2_2_n73,
         npu_inst_pe_1_2_2_n72, npu_inst_pe_1_2_2_n71, npu_inst_pe_1_2_2_n70,
         npu_inst_pe_1_2_2_n69, npu_inst_pe_1_2_2_n68, npu_inst_pe_1_2_2_n67,
         npu_inst_pe_1_2_2_n66, npu_inst_pe_1_2_2_n65, npu_inst_pe_1_2_2_n64,
         npu_inst_pe_1_2_2_n63, npu_inst_pe_1_2_2_n62, npu_inst_pe_1_2_2_n61,
         npu_inst_pe_1_2_2_n60, npu_inst_pe_1_2_2_n59, npu_inst_pe_1_2_2_n58,
         npu_inst_pe_1_2_2_n57, npu_inst_pe_1_2_2_n56, npu_inst_pe_1_2_2_n55,
         npu_inst_pe_1_2_2_n54, npu_inst_pe_1_2_2_n53, npu_inst_pe_1_2_2_n52,
         npu_inst_pe_1_2_2_n51, npu_inst_pe_1_2_2_n50, npu_inst_pe_1_2_2_n49,
         npu_inst_pe_1_2_2_n48, npu_inst_pe_1_2_2_n47, npu_inst_pe_1_2_2_n46,
         npu_inst_pe_1_2_2_n45, npu_inst_pe_1_2_2_n44, npu_inst_pe_1_2_2_n43,
         npu_inst_pe_1_2_2_n42, npu_inst_pe_1_2_2_n41, npu_inst_pe_1_2_2_n40,
         npu_inst_pe_1_2_2_n39, npu_inst_pe_1_2_2_n38, npu_inst_pe_1_2_2_n37,
         npu_inst_pe_1_2_2_n27, npu_inst_pe_1_2_2_n26,
         npu_inst_pe_1_2_2_net3885, npu_inst_pe_1_2_2_net3879,
         npu_inst_pe_1_2_2_N94, npu_inst_pe_1_2_2_N93, npu_inst_pe_1_2_2_N84,
         npu_inst_pe_1_2_2_N80, npu_inst_pe_1_2_2_N79, npu_inst_pe_1_2_2_N78,
         npu_inst_pe_1_2_2_N77, npu_inst_pe_1_2_2_N76, npu_inst_pe_1_2_2_N75,
         npu_inst_pe_1_2_2_N74, npu_inst_pe_1_2_2_N73, npu_inst_pe_1_2_2_N72,
         npu_inst_pe_1_2_2_N71, npu_inst_pe_1_2_2_N70, npu_inst_pe_1_2_2_N69,
         npu_inst_pe_1_2_2_N68, npu_inst_pe_1_2_2_N67, npu_inst_pe_1_2_2_N66,
         npu_inst_pe_1_2_2_N65, npu_inst_pe_1_2_2_int_q_acc_0_,
         npu_inst_pe_1_2_2_int_q_acc_1_, npu_inst_pe_1_2_2_int_q_acc_2_,
         npu_inst_pe_1_2_2_int_q_acc_3_, npu_inst_pe_1_2_2_int_q_acc_4_,
         npu_inst_pe_1_2_2_int_q_acc_5_, npu_inst_pe_1_2_2_int_q_acc_6_,
         npu_inst_pe_1_2_2_int_q_acc_7_, npu_inst_pe_1_2_2_int_data_0_,
         npu_inst_pe_1_2_2_int_data_1_, npu_inst_pe_1_2_2_int_q_weight_0_,
         npu_inst_pe_1_2_2_int_q_weight_1_,
         npu_inst_pe_1_2_2_int_q_reg_v_5__0_,
         npu_inst_pe_1_2_2_int_q_reg_v_5__1_,
         npu_inst_pe_1_2_2_int_q_reg_v_4__0_,
         npu_inst_pe_1_2_2_int_q_reg_v_4__1_,
         npu_inst_pe_1_2_2_int_q_reg_v_3__0_,
         npu_inst_pe_1_2_2_int_q_reg_v_3__1_,
         npu_inst_pe_1_2_2_int_q_reg_v_2__0_,
         npu_inst_pe_1_2_2_int_q_reg_v_2__1_,
         npu_inst_pe_1_2_2_int_q_reg_v_1__0_,
         npu_inst_pe_1_2_2_int_q_reg_v_1__1_,
         npu_inst_pe_1_2_2_int_q_reg_v_0__0_,
         npu_inst_pe_1_2_2_int_q_reg_v_0__1_,
         npu_inst_pe_1_2_2_int_q_reg_h_5__0_,
         npu_inst_pe_1_2_2_int_q_reg_h_5__1_,
         npu_inst_pe_1_2_2_int_q_reg_h_4__0_,
         npu_inst_pe_1_2_2_int_q_reg_h_4__1_,
         npu_inst_pe_1_2_2_int_q_reg_h_3__0_,
         npu_inst_pe_1_2_2_int_q_reg_h_3__1_,
         npu_inst_pe_1_2_2_int_q_reg_h_2__0_,
         npu_inst_pe_1_2_2_int_q_reg_h_2__1_,
         npu_inst_pe_1_2_2_int_q_reg_h_1__0_,
         npu_inst_pe_1_2_2_int_q_reg_h_1__1_,
         npu_inst_pe_1_2_2_int_q_reg_h_0__0_,
         npu_inst_pe_1_2_2_int_q_reg_h_0__1_, npu_inst_pe_1_2_3_n119,
         npu_inst_pe_1_2_3_n118, npu_inst_pe_1_2_3_n117,
         npu_inst_pe_1_2_3_n116, npu_inst_pe_1_2_3_n115,
         npu_inst_pe_1_2_3_n114, npu_inst_pe_1_2_3_n113,
         npu_inst_pe_1_2_3_n112, npu_inst_pe_1_2_3_n111,
         npu_inst_pe_1_2_3_n110, npu_inst_pe_1_2_3_n109,
         npu_inst_pe_1_2_3_n108, npu_inst_pe_1_2_3_n107,
         npu_inst_pe_1_2_3_n106, npu_inst_pe_1_2_3_n105,
         npu_inst_pe_1_2_3_n104, npu_inst_pe_1_2_3_n103,
         npu_inst_pe_1_2_3_n102, npu_inst_pe_1_2_3_n101,
         npu_inst_pe_1_2_3_n100, npu_inst_pe_1_2_3_n99, npu_inst_pe_1_2_3_n98,
         npu_inst_pe_1_2_3_n36, npu_inst_pe_1_2_3_n35, npu_inst_pe_1_2_3_n34,
         npu_inst_pe_1_2_3_n33, npu_inst_pe_1_2_3_n32, npu_inst_pe_1_2_3_n31,
         npu_inst_pe_1_2_3_n30, npu_inst_pe_1_2_3_n29, npu_inst_pe_1_2_3_n28,
         npu_inst_pe_1_2_3_n25, npu_inst_pe_1_2_3_n24, npu_inst_pe_1_2_3_n23,
         npu_inst_pe_1_2_3_n22, npu_inst_pe_1_2_3_n21, npu_inst_pe_1_2_3_n20,
         npu_inst_pe_1_2_3_n19, npu_inst_pe_1_2_3_n18, npu_inst_pe_1_2_3_n17,
         npu_inst_pe_1_2_3_n16, npu_inst_pe_1_2_3_n15, npu_inst_pe_1_2_3_n14,
         npu_inst_pe_1_2_3_n13, npu_inst_pe_1_2_3_n12, npu_inst_pe_1_2_3_n11,
         npu_inst_pe_1_2_3_n10, npu_inst_pe_1_2_3_n9, npu_inst_pe_1_2_3_n8,
         npu_inst_pe_1_2_3_n7, npu_inst_pe_1_2_3_n6, npu_inst_pe_1_2_3_n5,
         npu_inst_pe_1_2_3_n4, npu_inst_pe_1_2_3_n3, npu_inst_pe_1_2_3_n2,
         npu_inst_pe_1_2_3_n1, npu_inst_pe_1_2_3_sub_77_carry_7_,
         npu_inst_pe_1_2_3_sub_77_carry_6_, npu_inst_pe_1_2_3_sub_77_carry_5_,
         npu_inst_pe_1_2_3_sub_77_carry_4_, npu_inst_pe_1_2_3_sub_77_carry_3_,
         npu_inst_pe_1_2_3_sub_77_carry_2_, npu_inst_pe_1_2_3_sub_77_carry_1_,
         npu_inst_pe_1_2_3_add_79_carry_7_, npu_inst_pe_1_2_3_add_79_carry_6_,
         npu_inst_pe_1_2_3_add_79_carry_5_, npu_inst_pe_1_2_3_add_79_carry_4_,
         npu_inst_pe_1_2_3_add_79_carry_3_, npu_inst_pe_1_2_3_add_79_carry_2_,
         npu_inst_pe_1_2_3_add_79_carry_1_, npu_inst_pe_1_2_3_n97,
         npu_inst_pe_1_2_3_n96, npu_inst_pe_1_2_3_n95, npu_inst_pe_1_2_3_n94,
         npu_inst_pe_1_2_3_n93, npu_inst_pe_1_2_3_n92, npu_inst_pe_1_2_3_n91,
         npu_inst_pe_1_2_3_n90, npu_inst_pe_1_2_3_n89, npu_inst_pe_1_2_3_n88,
         npu_inst_pe_1_2_3_n87, npu_inst_pe_1_2_3_n86, npu_inst_pe_1_2_3_n85,
         npu_inst_pe_1_2_3_n84, npu_inst_pe_1_2_3_n83, npu_inst_pe_1_2_3_n82,
         npu_inst_pe_1_2_3_n81, npu_inst_pe_1_2_3_n80, npu_inst_pe_1_2_3_n79,
         npu_inst_pe_1_2_3_n78, npu_inst_pe_1_2_3_n77, npu_inst_pe_1_2_3_n76,
         npu_inst_pe_1_2_3_n75, npu_inst_pe_1_2_3_n74, npu_inst_pe_1_2_3_n73,
         npu_inst_pe_1_2_3_n72, npu_inst_pe_1_2_3_n71, npu_inst_pe_1_2_3_n70,
         npu_inst_pe_1_2_3_n69, npu_inst_pe_1_2_3_n68, npu_inst_pe_1_2_3_n67,
         npu_inst_pe_1_2_3_n66, npu_inst_pe_1_2_3_n65, npu_inst_pe_1_2_3_n64,
         npu_inst_pe_1_2_3_n63, npu_inst_pe_1_2_3_n62, npu_inst_pe_1_2_3_n61,
         npu_inst_pe_1_2_3_n60, npu_inst_pe_1_2_3_n59, npu_inst_pe_1_2_3_n58,
         npu_inst_pe_1_2_3_n57, npu_inst_pe_1_2_3_n56, npu_inst_pe_1_2_3_n55,
         npu_inst_pe_1_2_3_n54, npu_inst_pe_1_2_3_n53, npu_inst_pe_1_2_3_n52,
         npu_inst_pe_1_2_3_n51, npu_inst_pe_1_2_3_n50, npu_inst_pe_1_2_3_n49,
         npu_inst_pe_1_2_3_n48, npu_inst_pe_1_2_3_n47, npu_inst_pe_1_2_3_n46,
         npu_inst_pe_1_2_3_n45, npu_inst_pe_1_2_3_n44, npu_inst_pe_1_2_3_n43,
         npu_inst_pe_1_2_3_n42, npu_inst_pe_1_2_3_n41, npu_inst_pe_1_2_3_n40,
         npu_inst_pe_1_2_3_n39, npu_inst_pe_1_2_3_n38, npu_inst_pe_1_2_3_n37,
         npu_inst_pe_1_2_3_n27, npu_inst_pe_1_2_3_n26,
         npu_inst_pe_1_2_3_net3862, npu_inst_pe_1_2_3_net3856,
         npu_inst_pe_1_2_3_N94, npu_inst_pe_1_2_3_N93, npu_inst_pe_1_2_3_N84,
         npu_inst_pe_1_2_3_N80, npu_inst_pe_1_2_3_N79, npu_inst_pe_1_2_3_N78,
         npu_inst_pe_1_2_3_N77, npu_inst_pe_1_2_3_N76, npu_inst_pe_1_2_3_N75,
         npu_inst_pe_1_2_3_N74, npu_inst_pe_1_2_3_N73, npu_inst_pe_1_2_3_N72,
         npu_inst_pe_1_2_3_N71, npu_inst_pe_1_2_3_N70, npu_inst_pe_1_2_3_N69,
         npu_inst_pe_1_2_3_N68, npu_inst_pe_1_2_3_N67, npu_inst_pe_1_2_3_N66,
         npu_inst_pe_1_2_3_N65, npu_inst_pe_1_2_3_int_q_acc_0_,
         npu_inst_pe_1_2_3_int_q_acc_1_, npu_inst_pe_1_2_3_int_q_acc_2_,
         npu_inst_pe_1_2_3_int_q_acc_3_, npu_inst_pe_1_2_3_int_q_acc_4_,
         npu_inst_pe_1_2_3_int_q_acc_5_, npu_inst_pe_1_2_3_int_q_acc_6_,
         npu_inst_pe_1_2_3_int_q_acc_7_, npu_inst_pe_1_2_3_int_data_0_,
         npu_inst_pe_1_2_3_int_data_1_, npu_inst_pe_1_2_3_int_q_weight_0_,
         npu_inst_pe_1_2_3_int_q_weight_1_,
         npu_inst_pe_1_2_3_int_q_reg_v_5__0_,
         npu_inst_pe_1_2_3_int_q_reg_v_5__1_,
         npu_inst_pe_1_2_3_int_q_reg_v_4__0_,
         npu_inst_pe_1_2_3_int_q_reg_v_4__1_,
         npu_inst_pe_1_2_3_int_q_reg_v_3__0_,
         npu_inst_pe_1_2_3_int_q_reg_v_3__1_,
         npu_inst_pe_1_2_3_int_q_reg_v_2__0_,
         npu_inst_pe_1_2_3_int_q_reg_v_2__1_,
         npu_inst_pe_1_2_3_int_q_reg_v_1__0_,
         npu_inst_pe_1_2_3_int_q_reg_v_1__1_,
         npu_inst_pe_1_2_3_int_q_reg_v_0__0_,
         npu_inst_pe_1_2_3_int_q_reg_v_0__1_,
         npu_inst_pe_1_2_3_int_q_reg_h_5__0_,
         npu_inst_pe_1_2_3_int_q_reg_h_5__1_,
         npu_inst_pe_1_2_3_int_q_reg_h_4__0_,
         npu_inst_pe_1_2_3_int_q_reg_h_4__1_,
         npu_inst_pe_1_2_3_int_q_reg_h_3__0_,
         npu_inst_pe_1_2_3_int_q_reg_h_3__1_,
         npu_inst_pe_1_2_3_int_q_reg_h_2__0_,
         npu_inst_pe_1_2_3_int_q_reg_h_2__1_,
         npu_inst_pe_1_2_3_int_q_reg_h_1__0_,
         npu_inst_pe_1_2_3_int_q_reg_h_1__1_,
         npu_inst_pe_1_2_3_int_q_reg_h_0__0_,
         npu_inst_pe_1_2_3_int_q_reg_h_0__1_, npu_inst_pe_1_2_4_n119,
         npu_inst_pe_1_2_4_n118, npu_inst_pe_1_2_4_n117,
         npu_inst_pe_1_2_4_n116, npu_inst_pe_1_2_4_n115,
         npu_inst_pe_1_2_4_n114, npu_inst_pe_1_2_4_n113,
         npu_inst_pe_1_2_4_n112, npu_inst_pe_1_2_4_n111,
         npu_inst_pe_1_2_4_n110, npu_inst_pe_1_2_4_n109,
         npu_inst_pe_1_2_4_n108, npu_inst_pe_1_2_4_n107,
         npu_inst_pe_1_2_4_n106, npu_inst_pe_1_2_4_n105,
         npu_inst_pe_1_2_4_n104, npu_inst_pe_1_2_4_n103,
         npu_inst_pe_1_2_4_n102, npu_inst_pe_1_2_4_n101,
         npu_inst_pe_1_2_4_n100, npu_inst_pe_1_2_4_n99, npu_inst_pe_1_2_4_n98,
         npu_inst_pe_1_2_4_n36, npu_inst_pe_1_2_4_n35, npu_inst_pe_1_2_4_n34,
         npu_inst_pe_1_2_4_n33, npu_inst_pe_1_2_4_n32, npu_inst_pe_1_2_4_n31,
         npu_inst_pe_1_2_4_n30, npu_inst_pe_1_2_4_n29, npu_inst_pe_1_2_4_n28,
         npu_inst_pe_1_2_4_n25, npu_inst_pe_1_2_4_n24, npu_inst_pe_1_2_4_n23,
         npu_inst_pe_1_2_4_n22, npu_inst_pe_1_2_4_n21, npu_inst_pe_1_2_4_n20,
         npu_inst_pe_1_2_4_n19, npu_inst_pe_1_2_4_n18, npu_inst_pe_1_2_4_n17,
         npu_inst_pe_1_2_4_n16, npu_inst_pe_1_2_4_n15, npu_inst_pe_1_2_4_n14,
         npu_inst_pe_1_2_4_n13, npu_inst_pe_1_2_4_n12, npu_inst_pe_1_2_4_n11,
         npu_inst_pe_1_2_4_n10, npu_inst_pe_1_2_4_n9, npu_inst_pe_1_2_4_n8,
         npu_inst_pe_1_2_4_n7, npu_inst_pe_1_2_4_n6, npu_inst_pe_1_2_4_n5,
         npu_inst_pe_1_2_4_n4, npu_inst_pe_1_2_4_n3, npu_inst_pe_1_2_4_n2,
         npu_inst_pe_1_2_4_n1, npu_inst_pe_1_2_4_sub_77_carry_7_,
         npu_inst_pe_1_2_4_sub_77_carry_6_, npu_inst_pe_1_2_4_sub_77_carry_5_,
         npu_inst_pe_1_2_4_sub_77_carry_4_, npu_inst_pe_1_2_4_sub_77_carry_3_,
         npu_inst_pe_1_2_4_sub_77_carry_2_, npu_inst_pe_1_2_4_sub_77_carry_1_,
         npu_inst_pe_1_2_4_add_79_carry_7_, npu_inst_pe_1_2_4_add_79_carry_6_,
         npu_inst_pe_1_2_4_add_79_carry_5_, npu_inst_pe_1_2_4_add_79_carry_4_,
         npu_inst_pe_1_2_4_add_79_carry_3_, npu_inst_pe_1_2_4_add_79_carry_2_,
         npu_inst_pe_1_2_4_add_79_carry_1_, npu_inst_pe_1_2_4_n97,
         npu_inst_pe_1_2_4_n96, npu_inst_pe_1_2_4_n95, npu_inst_pe_1_2_4_n94,
         npu_inst_pe_1_2_4_n93, npu_inst_pe_1_2_4_n92, npu_inst_pe_1_2_4_n91,
         npu_inst_pe_1_2_4_n90, npu_inst_pe_1_2_4_n89, npu_inst_pe_1_2_4_n88,
         npu_inst_pe_1_2_4_n87, npu_inst_pe_1_2_4_n86, npu_inst_pe_1_2_4_n85,
         npu_inst_pe_1_2_4_n84, npu_inst_pe_1_2_4_n83, npu_inst_pe_1_2_4_n82,
         npu_inst_pe_1_2_4_n81, npu_inst_pe_1_2_4_n80, npu_inst_pe_1_2_4_n79,
         npu_inst_pe_1_2_4_n78, npu_inst_pe_1_2_4_n77, npu_inst_pe_1_2_4_n76,
         npu_inst_pe_1_2_4_n75, npu_inst_pe_1_2_4_n74, npu_inst_pe_1_2_4_n73,
         npu_inst_pe_1_2_4_n72, npu_inst_pe_1_2_4_n71, npu_inst_pe_1_2_4_n70,
         npu_inst_pe_1_2_4_n69, npu_inst_pe_1_2_4_n68, npu_inst_pe_1_2_4_n67,
         npu_inst_pe_1_2_4_n66, npu_inst_pe_1_2_4_n65, npu_inst_pe_1_2_4_n64,
         npu_inst_pe_1_2_4_n63, npu_inst_pe_1_2_4_n62, npu_inst_pe_1_2_4_n61,
         npu_inst_pe_1_2_4_n60, npu_inst_pe_1_2_4_n59, npu_inst_pe_1_2_4_n58,
         npu_inst_pe_1_2_4_n57, npu_inst_pe_1_2_4_n56, npu_inst_pe_1_2_4_n55,
         npu_inst_pe_1_2_4_n54, npu_inst_pe_1_2_4_n53, npu_inst_pe_1_2_4_n52,
         npu_inst_pe_1_2_4_n51, npu_inst_pe_1_2_4_n50, npu_inst_pe_1_2_4_n49,
         npu_inst_pe_1_2_4_n48, npu_inst_pe_1_2_4_n47, npu_inst_pe_1_2_4_n46,
         npu_inst_pe_1_2_4_n45, npu_inst_pe_1_2_4_n44, npu_inst_pe_1_2_4_n43,
         npu_inst_pe_1_2_4_n42, npu_inst_pe_1_2_4_n41, npu_inst_pe_1_2_4_n40,
         npu_inst_pe_1_2_4_n39, npu_inst_pe_1_2_4_n38, npu_inst_pe_1_2_4_n37,
         npu_inst_pe_1_2_4_n27, npu_inst_pe_1_2_4_n26,
         npu_inst_pe_1_2_4_net3839, npu_inst_pe_1_2_4_net3833,
         npu_inst_pe_1_2_4_N94, npu_inst_pe_1_2_4_N93, npu_inst_pe_1_2_4_N84,
         npu_inst_pe_1_2_4_N80, npu_inst_pe_1_2_4_N79, npu_inst_pe_1_2_4_N78,
         npu_inst_pe_1_2_4_N77, npu_inst_pe_1_2_4_N76, npu_inst_pe_1_2_4_N75,
         npu_inst_pe_1_2_4_N74, npu_inst_pe_1_2_4_N73, npu_inst_pe_1_2_4_N72,
         npu_inst_pe_1_2_4_N71, npu_inst_pe_1_2_4_N70, npu_inst_pe_1_2_4_N69,
         npu_inst_pe_1_2_4_N68, npu_inst_pe_1_2_4_N67, npu_inst_pe_1_2_4_N66,
         npu_inst_pe_1_2_4_N65, npu_inst_pe_1_2_4_int_q_acc_0_,
         npu_inst_pe_1_2_4_int_q_acc_1_, npu_inst_pe_1_2_4_int_q_acc_2_,
         npu_inst_pe_1_2_4_int_q_acc_3_, npu_inst_pe_1_2_4_int_q_acc_4_,
         npu_inst_pe_1_2_4_int_q_acc_5_, npu_inst_pe_1_2_4_int_q_acc_6_,
         npu_inst_pe_1_2_4_int_q_acc_7_, npu_inst_pe_1_2_4_int_data_0_,
         npu_inst_pe_1_2_4_int_data_1_, npu_inst_pe_1_2_4_int_q_weight_0_,
         npu_inst_pe_1_2_4_int_q_weight_1_,
         npu_inst_pe_1_2_4_int_q_reg_v_5__0_,
         npu_inst_pe_1_2_4_int_q_reg_v_5__1_,
         npu_inst_pe_1_2_4_int_q_reg_v_4__0_,
         npu_inst_pe_1_2_4_int_q_reg_v_4__1_,
         npu_inst_pe_1_2_4_int_q_reg_v_3__0_,
         npu_inst_pe_1_2_4_int_q_reg_v_3__1_,
         npu_inst_pe_1_2_4_int_q_reg_v_2__0_,
         npu_inst_pe_1_2_4_int_q_reg_v_2__1_,
         npu_inst_pe_1_2_4_int_q_reg_v_1__0_,
         npu_inst_pe_1_2_4_int_q_reg_v_1__1_,
         npu_inst_pe_1_2_4_int_q_reg_v_0__0_,
         npu_inst_pe_1_2_4_int_q_reg_v_0__1_,
         npu_inst_pe_1_2_4_int_q_reg_h_5__0_,
         npu_inst_pe_1_2_4_int_q_reg_h_5__1_,
         npu_inst_pe_1_2_4_int_q_reg_h_4__0_,
         npu_inst_pe_1_2_4_int_q_reg_h_4__1_,
         npu_inst_pe_1_2_4_int_q_reg_h_3__0_,
         npu_inst_pe_1_2_4_int_q_reg_h_3__1_,
         npu_inst_pe_1_2_4_int_q_reg_h_2__0_,
         npu_inst_pe_1_2_4_int_q_reg_h_2__1_,
         npu_inst_pe_1_2_4_int_q_reg_h_1__0_,
         npu_inst_pe_1_2_4_int_q_reg_h_1__1_,
         npu_inst_pe_1_2_4_int_q_reg_h_0__0_,
         npu_inst_pe_1_2_4_int_q_reg_h_0__1_, npu_inst_pe_1_2_5_n119,
         npu_inst_pe_1_2_5_n118, npu_inst_pe_1_2_5_n117,
         npu_inst_pe_1_2_5_n116, npu_inst_pe_1_2_5_n115,
         npu_inst_pe_1_2_5_n114, npu_inst_pe_1_2_5_n113,
         npu_inst_pe_1_2_5_n112, npu_inst_pe_1_2_5_n111,
         npu_inst_pe_1_2_5_n110, npu_inst_pe_1_2_5_n109,
         npu_inst_pe_1_2_5_n108, npu_inst_pe_1_2_5_n107,
         npu_inst_pe_1_2_5_n106, npu_inst_pe_1_2_5_n105,
         npu_inst_pe_1_2_5_n104, npu_inst_pe_1_2_5_n103,
         npu_inst_pe_1_2_5_n102, npu_inst_pe_1_2_5_n101,
         npu_inst_pe_1_2_5_n100, npu_inst_pe_1_2_5_n99, npu_inst_pe_1_2_5_n98,
         npu_inst_pe_1_2_5_n36, npu_inst_pe_1_2_5_n35, npu_inst_pe_1_2_5_n34,
         npu_inst_pe_1_2_5_n33, npu_inst_pe_1_2_5_n32, npu_inst_pe_1_2_5_n31,
         npu_inst_pe_1_2_5_n30, npu_inst_pe_1_2_5_n29, npu_inst_pe_1_2_5_n28,
         npu_inst_pe_1_2_5_n25, npu_inst_pe_1_2_5_n24, npu_inst_pe_1_2_5_n23,
         npu_inst_pe_1_2_5_n22, npu_inst_pe_1_2_5_n21, npu_inst_pe_1_2_5_n20,
         npu_inst_pe_1_2_5_n19, npu_inst_pe_1_2_5_n18, npu_inst_pe_1_2_5_n17,
         npu_inst_pe_1_2_5_n16, npu_inst_pe_1_2_5_n15, npu_inst_pe_1_2_5_n14,
         npu_inst_pe_1_2_5_n13, npu_inst_pe_1_2_5_n12, npu_inst_pe_1_2_5_n11,
         npu_inst_pe_1_2_5_n10, npu_inst_pe_1_2_5_n9, npu_inst_pe_1_2_5_n8,
         npu_inst_pe_1_2_5_n7, npu_inst_pe_1_2_5_n6, npu_inst_pe_1_2_5_n5,
         npu_inst_pe_1_2_5_n4, npu_inst_pe_1_2_5_n3, npu_inst_pe_1_2_5_n2,
         npu_inst_pe_1_2_5_n1, npu_inst_pe_1_2_5_sub_77_carry_7_,
         npu_inst_pe_1_2_5_sub_77_carry_6_, npu_inst_pe_1_2_5_sub_77_carry_5_,
         npu_inst_pe_1_2_5_sub_77_carry_4_, npu_inst_pe_1_2_5_sub_77_carry_3_,
         npu_inst_pe_1_2_5_sub_77_carry_2_, npu_inst_pe_1_2_5_sub_77_carry_1_,
         npu_inst_pe_1_2_5_add_79_carry_7_, npu_inst_pe_1_2_5_add_79_carry_6_,
         npu_inst_pe_1_2_5_add_79_carry_5_, npu_inst_pe_1_2_5_add_79_carry_4_,
         npu_inst_pe_1_2_5_add_79_carry_3_, npu_inst_pe_1_2_5_add_79_carry_2_,
         npu_inst_pe_1_2_5_add_79_carry_1_, npu_inst_pe_1_2_5_n97,
         npu_inst_pe_1_2_5_n96, npu_inst_pe_1_2_5_n95, npu_inst_pe_1_2_5_n94,
         npu_inst_pe_1_2_5_n93, npu_inst_pe_1_2_5_n92, npu_inst_pe_1_2_5_n91,
         npu_inst_pe_1_2_5_n90, npu_inst_pe_1_2_5_n89, npu_inst_pe_1_2_5_n88,
         npu_inst_pe_1_2_5_n87, npu_inst_pe_1_2_5_n86, npu_inst_pe_1_2_5_n85,
         npu_inst_pe_1_2_5_n84, npu_inst_pe_1_2_5_n83, npu_inst_pe_1_2_5_n82,
         npu_inst_pe_1_2_5_n81, npu_inst_pe_1_2_5_n80, npu_inst_pe_1_2_5_n79,
         npu_inst_pe_1_2_5_n78, npu_inst_pe_1_2_5_n77, npu_inst_pe_1_2_5_n76,
         npu_inst_pe_1_2_5_n75, npu_inst_pe_1_2_5_n74, npu_inst_pe_1_2_5_n73,
         npu_inst_pe_1_2_5_n72, npu_inst_pe_1_2_5_n71, npu_inst_pe_1_2_5_n70,
         npu_inst_pe_1_2_5_n69, npu_inst_pe_1_2_5_n68, npu_inst_pe_1_2_5_n67,
         npu_inst_pe_1_2_5_n66, npu_inst_pe_1_2_5_n65, npu_inst_pe_1_2_5_n64,
         npu_inst_pe_1_2_5_n63, npu_inst_pe_1_2_5_n62, npu_inst_pe_1_2_5_n61,
         npu_inst_pe_1_2_5_n60, npu_inst_pe_1_2_5_n59, npu_inst_pe_1_2_5_n58,
         npu_inst_pe_1_2_5_n57, npu_inst_pe_1_2_5_n56, npu_inst_pe_1_2_5_n55,
         npu_inst_pe_1_2_5_n54, npu_inst_pe_1_2_5_n53, npu_inst_pe_1_2_5_n52,
         npu_inst_pe_1_2_5_n51, npu_inst_pe_1_2_5_n50, npu_inst_pe_1_2_5_n49,
         npu_inst_pe_1_2_5_n48, npu_inst_pe_1_2_5_n47, npu_inst_pe_1_2_5_n46,
         npu_inst_pe_1_2_5_n45, npu_inst_pe_1_2_5_n44, npu_inst_pe_1_2_5_n43,
         npu_inst_pe_1_2_5_n42, npu_inst_pe_1_2_5_n41, npu_inst_pe_1_2_5_n40,
         npu_inst_pe_1_2_5_n39, npu_inst_pe_1_2_5_n38, npu_inst_pe_1_2_5_n37,
         npu_inst_pe_1_2_5_n27, npu_inst_pe_1_2_5_n26,
         npu_inst_pe_1_2_5_net3816, npu_inst_pe_1_2_5_net3810,
         npu_inst_pe_1_2_5_N94, npu_inst_pe_1_2_5_N93, npu_inst_pe_1_2_5_N84,
         npu_inst_pe_1_2_5_N80, npu_inst_pe_1_2_5_N79, npu_inst_pe_1_2_5_N78,
         npu_inst_pe_1_2_5_N77, npu_inst_pe_1_2_5_N76, npu_inst_pe_1_2_5_N75,
         npu_inst_pe_1_2_5_N74, npu_inst_pe_1_2_5_N73, npu_inst_pe_1_2_5_N72,
         npu_inst_pe_1_2_5_N71, npu_inst_pe_1_2_5_N70, npu_inst_pe_1_2_5_N69,
         npu_inst_pe_1_2_5_N68, npu_inst_pe_1_2_5_N67, npu_inst_pe_1_2_5_N66,
         npu_inst_pe_1_2_5_N65, npu_inst_pe_1_2_5_int_q_acc_0_,
         npu_inst_pe_1_2_5_int_q_acc_1_, npu_inst_pe_1_2_5_int_q_acc_2_,
         npu_inst_pe_1_2_5_int_q_acc_3_, npu_inst_pe_1_2_5_int_q_acc_4_,
         npu_inst_pe_1_2_5_int_q_acc_5_, npu_inst_pe_1_2_5_int_q_acc_6_,
         npu_inst_pe_1_2_5_int_q_acc_7_, npu_inst_pe_1_2_5_int_data_0_,
         npu_inst_pe_1_2_5_int_data_1_, npu_inst_pe_1_2_5_int_q_weight_0_,
         npu_inst_pe_1_2_5_int_q_weight_1_,
         npu_inst_pe_1_2_5_int_q_reg_v_5__0_,
         npu_inst_pe_1_2_5_int_q_reg_v_5__1_,
         npu_inst_pe_1_2_5_int_q_reg_v_4__0_,
         npu_inst_pe_1_2_5_int_q_reg_v_4__1_,
         npu_inst_pe_1_2_5_int_q_reg_v_3__0_,
         npu_inst_pe_1_2_5_int_q_reg_v_3__1_,
         npu_inst_pe_1_2_5_int_q_reg_v_2__0_,
         npu_inst_pe_1_2_5_int_q_reg_v_2__1_,
         npu_inst_pe_1_2_5_int_q_reg_v_1__0_,
         npu_inst_pe_1_2_5_int_q_reg_v_1__1_,
         npu_inst_pe_1_2_5_int_q_reg_v_0__0_,
         npu_inst_pe_1_2_5_int_q_reg_v_0__1_,
         npu_inst_pe_1_2_5_int_q_reg_h_5__0_,
         npu_inst_pe_1_2_5_int_q_reg_h_5__1_,
         npu_inst_pe_1_2_5_int_q_reg_h_4__0_,
         npu_inst_pe_1_2_5_int_q_reg_h_4__1_,
         npu_inst_pe_1_2_5_int_q_reg_h_3__0_,
         npu_inst_pe_1_2_5_int_q_reg_h_3__1_,
         npu_inst_pe_1_2_5_int_q_reg_h_2__0_,
         npu_inst_pe_1_2_5_int_q_reg_h_2__1_,
         npu_inst_pe_1_2_5_int_q_reg_h_1__0_,
         npu_inst_pe_1_2_5_int_q_reg_h_1__1_,
         npu_inst_pe_1_2_5_int_q_reg_h_0__0_,
         npu_inst_pe_1_2_5_int_q_reg_h_0__1_, npu_inst_pe_1_2_6_n119,
         npu_inst_pe_1_2_6_n118, npu_inst_pe_1_2_6_n117,
         npu_inst_pe_1_2_6_n116, npu_inst_pe_1_2_6_n115,
         npu_inst_pe_1_2_6_n114, npu_inst_pe_1_2_6_n113,
         npu_inst_pe_1_2_6_n112, npu_inst_pe_1_2_6_n111,
         npu_inst_pe_1_2_6_n110, npu_inst_pe_1_2_6_n109,
         npu_inst_pe_1_2_6_n108, npu_inst_pe_1_2_6_n107,
         npu_inst_pe_1_2_6_n106, npu_inst_pe_1_2_6_n105,
         npu_inst_pe_1_2_6_n104, npu_inst_pe_1_2_6_n103,
         npu_inst_pe_1_2_6_n102, npu_inst_pe_1_2_6_n101,
         npu_inst_pe_1_2_6_n100, npu_inst_pe_1_2_6_n99, npu_inst_pe_1_2_6_n98,
         npu_inst_pe_1_2_6_n36, npu_inst_pe_1_2_6_n35, npu_inst_pe_1_2_6_n34,
         npu_inst_pe_1_2_6_n33, npu_inst_pe_1_2_6_n32, npu_inst_pe_1_2_6_n31,
         npu_inst_pe_1_2_6_n30, npu_inst_pe_1_2_6_n29, npu_inst_pe_1_2_6_n28,
         npu_inst_pe_1_2_6_n25, npu_inst_pe_1_2_6_n24, npu_inst_pe_1_2_6_n23,
         npu_inst_pe_1_2_6_n22, npu_inst_pe_1_2_6_n21, npu_inst_pe_1_2_6_n20,
         npu_inst_pe_1_2_6_n19, npu_inst_pe_1_2_6_n18, npu_inst_pe_1_2_6_n17,
         npu_inst_pe_1_2_6_n16, npu_inst_pe_1_2_6_n15, npu_inst_pe_1_2_6_n14,
         npu_inst_pe_1_2_6_n13, npu_inst_pe_1_2_6_n12, npu_inst_pe_1_2_6_n11,
         npu_inst_pe_1_2_6_n10, npu_inst_pe_1_2_6_n9, npu_inst_pe_1_2_6_n8,
         npu_inst_pe_1_2_6_n7, npu_inst_pe_1_2_6_n6, npu_inst_pe_1_2_6_n5,
         npu_inst_pe_1_2_6_n4, npu_inst_pe_1_2_6_n3, npu_inst_pe_1_2_6_n2,
         npu_inst_pe_1_2_6_n1, npu_inst_pe_1_2_6_sub_77_carry_7_,
         npu_inst_pe_1_2_6_sub_77_carry_6_, npu_inst_pe_1_2_6_sub_77_carry_5_,
         npu_inst_pe_1_2_6_sub_77_carry_4_, npu_inst_pe_1_2_6_sub_77_carry_3_,
         npu_inst_pe_1_2_6_sub_77_carry_2_, npu_inst_pe_1_2_6_sub_77_carry_1_,
         npu_inst_pe_1_2_6_add_79_carry_7_, npu_inst_pe_1_2_6_add_79_carry_6_,
         npu_inst_pe_1_2_6_add_79_carry_5_, npu_inst_pe_1_2_6_add_79_carry_4_,
         npu_inst_pe_1_2_6_add_79_carry_3_, npu_inst_pe_1_2_6_add_79_carry_2_,
         npu_inst_pe_1_2_6_add_79_carry_1_, npu_inst_pe_1_2_6_n97,
         npu_inst_pe_1_2_6_n96, npu_inst_pe_1_2_6_n95, npu_inst_pe_1_2_6_n94,
         npu_inst_pe_1_2_6_n93, npu_inst_pe_1_2_6_n92, npu_inst_pe_1_2_6_n91,
         npu_inst_pe_1_2_6_n90, npu_inst_pe_1_2_6_n89, npu_inst_pe_1_2_6_n88,
         npu_inst_pe_1_2_6_n87, npu_inst_pe_1_2_6_n86, npu_inst_pe_1_2_6_n85,
         npu_inst_pe_1_2_6_n84, npu_inst_pe_1_2_6_n83, npu_inst_pe_1_2_6_n82,
         npu_inst_pe_1_2_6_n81, npu_inst_pe_1_2_6_n80, npu_inst_pe_1_2_6_n79,
         npu_inst_pe_1_2_6_n78, npu_inst_pe_1_2_6_n77, npu_inst_pe_1_2_6_n76,
         npu_inst_pe_1_2_6_n75, npu_inst_pe_1_2_6_n74, npu_inst_pe_1_2_6_n73,
         npu_inst_pe_1_2_6_n72, npu_inst_pe_1_2_6_n71, npu_inst_pe_1_2_6_n70,
         npu_inst_pe_1_2_6_n69, npu_inst_pe_1_2_6_n68, npu_inst_pe_1_2_6_n67,
         npu_inst_pe_1_2_6_n66, npu_inst_pe_1_2_6_n65, npu_inst_pe_1_2_6_n64,
         npu_inst_pe_1_2_6_n63, npu_inst_pe_1_2_6_n62, npu_inst_pe_1_2_6_n61,
         npu_inst_pe_1_2_6_n60, npu_inst_pe_1_2_6_n59, npu_inst_pe_1_2_6_n58,
         npu_inst_pe_1_2_6_n57, npu_inst_pe_1_2_6_n56, npu_inst_pe_1_2_6_n55,
         npu_inst_pe_1_2_6_n54, npu_inst_pe_1_2_6_n53, npu_inst_pe_1_2_6_n52,
         npu_inst_pe_1_2_6_n51, npu_inst_pe_1_2_6_n50, npu_inst_pe_1_2_6_n49,
         npu_inst_pe_1_2_6_n48, npu_inst_pe_1_2_6_n47, npu_inst_pe_1_2_6_n46,
         npu_inst_pe_1_2_6_n45, npu_inst_pe_1_2_6_n44, npu_inst_pe_1_2_6_n43,
         npu_inst_pe_1_2_6_n42, npu_inst_pe_1_2_6_n41, npu_inst_pe_1_2_6_n40,
         npu_inst_pe_1_2_6_n39, npu_inst_pe_1_2_6_n38, npu_inst_pe_1_2_6_n37,
         npu_inst_pe_1_2_6_n27, npu_inst_pe_1_2_6_n26,
         npu_inst_pe_1_2_6_net3793, npu_inst_pe_1_2_6_net3787,
         npu_inst_pe_1_2_6_N94, npu_inst_pe_1_2_6_N93, npu_inst_pe_1_2_6_N84,
         npu_inst_pe_1_2_6_N80, npu_inst_pe_1_2_6_N79, npu_inst_pe_1_2_6_N78,
         npu_inst_pe_1_2_6_N77, npu_inst_pe_1_2_6_N76, npu_inst_pe_1_2_6_N75,
         npu_inst_pe_1_2_6_N74, npu_inst_pe_1_2_6_N73, npu_inst_pe_1_2_6_N72,
         npu_inst_pe_1_2_6_N71, npu_inst_pe_1_2_6_N70, npu_inst_pe_1_2_6_N69,
         npu_inst_pe_1_2_6_N68, npu_inst_pe_1_2_6_N67, npu_inst_pe_1_2_6_N66,
         npu_inst_pe_1_2_6_N65, npu_inst_pe_1_2_6_int_q_acc_0_,
         npu_inst_pe_1_2_6_int_q_acc_1_, npu_inst_pe_1_2_6_int_q_acc_2_,
         npu_inst_pe_1_2_6_int_q_acc_3_, npu_inst_pe_1_2_6_int_q_acc_4_,
         npu_inst_pe_1_2_6_int_q_acc_5_, npu_inst_pe_1_2_6_int_q_acc_6_,
         npu_inst_pe_1_2_6_int_q_acc_7_, npu_inst_pe_1_2_6_int_data_0_,
         npu_inst_pe_1_2_6_int_data_1_, npu_inst_pe_1_2_6_int_q_weight_0_,
         npu_inst_pe_1_2_6_int_q_weight_1_,
         npu_inst_pe_1_2_6_int_q_reg_v_5__0_,
         npu_inst_pe_1_2_6_int_q_reg_v_5__1_,
         npu_inst_pe_1_2_6_int_q_reg_v_4__0_,
         npu_inst_pe_1_2_6_int_q_reg_v_4__1_,
         npu_inst_pe_1_2_6_int_q_reg_v_3__0_,
         npu_inst_pe_1_2_6_int_q_reg_v_3__1_,
         npu_inst_pe_1_2_6_int_q_reg_v_2__0_,
         npu_inst_pe_1_2_6_int_q_reg_v_2__1_,
         npu_inst_pe_1_2_6_int_q_reg_v_1__0_,
         npu_inst_pe_1_2_6_int_q_reg_v_1__1_,
         npu_inst_pe_1_2_6_int_q_reg_v_0__0_,
         npu_inst_pe_1_2_6_int_q_reg_v_0__1_,
         npu_inst_pe_1_2_6_int_q_reg_h_5__0_,
         npu_inst_pe_1_2_6_int_q_reg_h_5__1_,
         npu_inst_pe_1_2_6_int_q_reg_h_4__0_,
         npu_inst_pe_1_2_6_int_q_reg_h_4__1_,
         npu_inst_pe_1_2_6_int_q_reg_h_3__0_,
         npu_inst_pe_1_2_6_int_q_reg_h_3__1_,
         npu_inst_pe_1_2_6_int_q_reg_h_2__0_,
         npu_inst_pe_1_2_6_int_q_reg_h_2__1_,
         npu_inst_pe_1_2_6_int_q_reg_h_1__0_,
         npu_inst_pe_1_2_6_int_q_reg_h_1__1_,
         npu_inst_pe_1_2_6_int_q_reg_h_0__0_,
         npu_inst_pe_1_2_6_int_q_reg_h_0__1_, npu_inst_pe_1_2_7_n119,
         npu_inst_pe_1_2_7_n118, npu_inst_pe_1_2_7_n117,
         npu_inst_pe_1_2_7_n116, npu_inst_pe_1_2_7_n115,
         npu_inst_pe_1_2_7_n114, npu_inst_pe_1_2_7_n113,
         npu_inst_pe_1_2_7_n112, npu_inst_pe_1_2_7_n111,
         npu_inst_pe_1_2_7_n110, npu_inst_pe_1_2_7_n109,
         npu_inst_pe_1_2_7_n108, npu_inst_pe_1_2_7_n107,
         npu_inst_pe_1_2_7_n106, npu_inst_pe_1_2_7_n105,
         npu_inst_pe_1_2_7_n104, npu_inst_pe_1_2_7_n103,
         npu_inst_pe_1_2_7_n102, npu_inst_pe_1_2_7_n101,
         npu_inst_pe_1_2_7_n100, npu_inst_pe_1_2_7_n99, npu_inst_pe_1_2_7_n98,
         npu_inst_pe_1_2_7_n36, npu_inst_pe_1_2_7_n35, npu_inst_pe_1_2_7_n34,
         npu_inst_pe_1_2_7_n33, npu_inst_pe_1_2_7_n32, npu_inst_pe_1_2_7_n31,
         npu_inst_pe_1_2_7_n30, npu_inst_pe_1_2_7_n29, npu_inst_pe_1_2_7_n28,
         npu_inst_pe_1_2_7_n25, npu_inst_pe_1_2_7_n24, npu_inst_pe_1_2_7_n23,
         npu_inst_pe_1_2_7_n22, npu_inst_pe_1_2_7_n21, npu_inst_pe_1_2_7_n20,
         npu_inst_pe_1_2_7_n19, npu_inst_pe_1_2_7_n18, npu_inst_pe_1_2_7_n17,
         npu_inst_pe_1_2_7_n16, npu_inst_pe_1_2_7_n15, npu_inst_pe_1_2_7_n14,
         npu_inst_pe_1_2_7_n13, npu_inst_pe_1_2_7_n12, npu_inst_pe_1_2_7_n11,
         npu_inst_pe_1_2_7_n10, npu_inst_pe_1_2_7_n9, npu_inst_pe_1_2_7_n8,
         npu_inst_pe_1_2_7_n7, npu_inst_pe_1_2_7_n6, npu_inst_pe_1_2_7_n5,
         npu_inst_pe_1_2_7_n4, npu_inst_pe_1_2_7_n3, npu_inst_pe_1_2_7_n2,
         npu_inst_pe_1_2_7_n1, npu_inst_pe_1_2_7_sub_77_carry_7_,
         npu_inst_pe_1_2_7_sub_77_carry_6_, npu_inst_pe_1_2_7_sub_77_carry_5_,
         npu_inst_pe_1_2_7_sub_77_carry_4_, npu_inst_pe_1_2_7_sub_77_carry_3_,
         npu_inst_pe_1_2_7_sub_77_carry_2_, npu_inst_pe_1_2_7_sub_77_carry_1_,
         npu_inst_pe_1_2_7_add_79_carry_7_, npu_inst_pe_1_2_7_add_79_carry_6_,
         npu_inst_pe_1_2_7_add_79_carry_5_, npu_inst_pe_1_2_7_add_79_carry_4_,
         npu_inst_pe_1_2_7_add_79_carry_3_, npu_inst_pe_1_2_7_add_79_carry_2_,
         npu_inst_pe_1_2_7_add_79_carry_1_, npu_inst_pe_1_2_7_n97,
         npu_inst_pe_1_2_7_n96, npu_inst_pe_1_2_7_n95, npu_inst_pe_1_2_7_n94,
         npu_inst_pe_1_2_7_n93, npu_inst_pe_1_2_7_n92, npu_inst_pe_1_2_7_n91,
         npu_inst_pe_1_2_7_n90, npu_inst_pe_1_2_7_n89, npu_inst_pe_1_2_7_n88,
         npu_inst_pe_1_2_7_n87, npu_inst_pe_1_2_7_n86, npu_inst_pe_1_2_7_n85,
         npu_inst_pe_1_2_7_n84, npu_inst_pe_1_2_7_n83, npu_inst_pe_1_2_7_n82,
         npu_inst_pe_1_2_7_n81, npu_inst_pe_1_2_7_n80, npu_inst_pe_1_2_7_n79,
         npu_inst_pe_1_2_7_n78, npu_inst_pe_1_2_7_n77, npu_inst_pe_1_2_7_n76,
         npu_inst_pe_1_2_7_n75, npu_inst_pe_1_2_7_n74, npu_inst_pe_1_2_7_n73,
         npu_inst_pe_1_2_7_n72, npu_inst_pe_1_2_7_n71, npu_inst_pe_1_2_7_n70,
         npu_inst_pe_1_2_7_n69, npu_inst_pe_1_2_7_n68, npu_inst_pe_1_2_7_n67,
         npu_inst_pe_1_2_7_n66, npu_inst_pe_1_2_7_n65, npu_inst_pe_1_2_7_n64,
         npu_inst_pe_1_2_7_n63, npu_inst_pe_1_2_7_n62, npu_inst_pe_1_2_7_n61,
         npu_inst_pe_1_2_7_n60, npu_inst_pe_1_2_7_n59, npu_inst_pe_1_2_7_n58,
         npu_inst_pe_1_2_7_n57, npu_inst_pe_1_2_7_n56, npu_inst_pe_1_2_7_n55,
         npu_inst_pe_1_2_7_n54, npu_inst_pe_1_2_7_n53, npu_inst_pe_1_2_7_n52,
         npu_inst_pe_1_2_7_n51, npu_inst_pe_1_2_7_n50, npu_inst_pe_1_2_7_n49,
         npu_inst_pe_1_2_7_n48, npu_inst_pe_1_2_7_n47, npu_inst_pe_1_2_7_n46,
         npu_inst_pe_1_2_7_n45, npu_inst_pe_1_2_7_n44, npu_inst_pe_1_2_7_n43,
         npu_inst_pe_1_2_7_n42, npu_inst_pe_1_2_7_n41, npu_inst_pe_1_2_7_n40,
         npu_inst_pe_1_2_7_n39, npu_inst_pe_1_2_7_n38, npu_inst_pe_1_2_7_n37,
         npu_inst_pe_1_2_7_n27, npu_inst_pe_1_2_7_n26,
         npu_inst_pe_1_2_7_net3770, npu_inst_pe_1_2_7_net3764,
         npu_inst_pe_1_2_7_N94, npu_inst_pe_1_2_7_N93, npu_inst_pe_1_2_7_N84,
         npu_inst_pe_1_2_7_N80, npu_inst_pe_1_2_7_N79, npu_inst_pe_1_2_7_N78,
         npu_inst_pe_1_2_7_N77, npu_inst_pe_1_2_7_N76, npu_inst_pe_1_2_7_N75,
         npu_inst_pe_1_2_7_N74, npu_inst_pe_1_2_7_N73, npu_inst_pe_1_2_7_N72,
         npu_inst_pe_1_2_7_N71, npu_inst_pe_1_2_7_N70, npu_inst_pe_1_2_7_N69,
         npu_inst_pe_1_2_7_N68, npu_inst_pe_1_2_7_N67, npu_inst_pe_1_2_7_N66,
         npu_inst_pe_1_2_7_N65, npu_inst_pe_1_2_7_int_q_acc_0_,
         npu_inst_pe_1_2_7_int_q_acc_1_, npu_inst_pe_1_2_7_int_q_acc_2_,
         npu_inst_pe_1_2_7_int_q_acc_3_, npu_inst_pe_1_2_7_int_q_acc_4_,
         npu_inst_pe_1_2_7_int_q_acc_5_, npu_inst_pe_1_2_7_int_q_acc_6_,
         npu_inst_pe_1_2_7_int_q_acc_7_, npu_inst_pe_1_2_7_int_data_0_,
         npu_inst_pe_1_2_7_int_data_1_, npu_inst_pe_1_2_7_int_q_weight_0_,
         npu_inst_pe_1_2_7_int_q_weight_1_,
         npu_inst_pe_1_2_7_int_q_reg_v_5__0_,
         npu_inst_pe_1_2_7_int_q_reg_v_5__1_,
         npu_inst_pe_1_2_7_int_q_reg_v_4__0_,
         npu_inst_pe_1_2_7_int_q_reg_v_4__1_,
         npu_inst_pe_1_2_7_int_q_reg_v_3__0_,
         npu_inst_pe_1_2_7_int_q_reg_v_3__1_,
         npu_inst_pe_1_2_7_int_q_reg_v_2__0_,
         npu_inst_pe_1_2_7_int_q_reg_v_2__1_,
         npu_inst_pe_1_2_7_int_q_reg_v_1__0_,
         npu_inst_pe_1_2_7_int_q_reg_v_1__1_,
         npu_inst_pe_1_2_7_int_q_reg_v_0__0_,
         npu_inst_pe_1_2_7_int_q_reg_v_0__1_,
         npu_inst_pe_1_2_7_int_q_reg_h_5__0_,
         npu_inst_pe_1_2_7_int_q_reg_h_5__1_,
         npu_inst_pe_1_2_7_int_q_reg_h_4__0_,
         npu_inst_pe_1_2_7_int_q_reg_h_4__1_,
         npu_inst_pe_1_2_7_int_q_reg_h_3__0_,
         npu_inst_pe_1_2_7_int_q_reg_h_3__1_,
         npu_inst_pe_1_2_7_int_q_reg_h_2__0_,
         npu_inst_pe_1_2_7_int_q_reg_h_2__1_,
         npu_inst_pe_1_2_7_int_q_reg_h_1__0_,
         npu_inst_pe_1_2_7_int_q_reg_h_1__1_,
         npu_inst_pe_1_2_7_int_q_reg_h_0__0_,
         npu_inst_pe_1_2_7_int_q_reg_h_0__1_, npu_inst_pe_1_3_0_n119,
         npu_inst_pe_1_3_0_n118, npu_inst_pe_1_3_0_n117,
         npu_inst_pe_1_3_0_n116, npu_inst_pe_1_3_0_n115,
         npu_inst_pe_1_3_0_n114, npu_inst_pe_1_3_0_n113,
         npu_inst_pe_1_3_0_n112, npu_inst_pe_1_3_0_n111,
         npu_inst_pe_1_3_0_n110, npu_inst_pe_1_3_0_n109,
         npu_inst_pe_1_3_0_n108, npu_inst_pe_1_3_0_n107,
         npu_inst_pe_1_3_0_n106, npu_inst_pe_1_3_0_n105,
         npu_inst_pe_1_3_0_n104, npu_inst_pe_1_3_0_n103,
         npu_inst_pe_1_3_0_n102, npu_inst_pe_1_3_0_n101,
         npu_inst_pe_1_3_0_n100, npu_inst_pe_1_3_0_n99, npu_inst_pe_1_3_0_n98,
         npu_inst_pe_1_3_0_n36, npu_inst_pe_1_3_0_n35, npu_inst_pe_1_3_0_n34,
         npu_inst_pe_1_3_0_n33, npu_inst_pe_1_3_0_n32, npu_inst_pe_1_3_0_n31,
         npu_inst_pe_1_3_0_n30, npu_inst_pe_1_3_0_n29, npu_inst_pe_1_3_0_n28,
         npu_inst_pe_1_3_0_n25, npu_inst_pe_1_3_0_n24, npu_inst_pe_1_3_0_n23,
         npu_inst_pe_1_3_0_n22, npu_inst_pe_1_3_0_n21, npu_inst_pe_1_3_0_n20,
         npu_inst_pe_1_3_0_n19, npu_inst_pe_1_3_0_n18, npu_inst_pe_1_3_0_n17,
         npu_inst_pe_1_3_0_n16, npu_inst_pe_1_3_0_n15, npu_inst_pe_1_3_0_n14,
         npu_inst_pe_1_3_0_n13, npu_inst_pe_1_3_0_n12, npu_inst_pe_1_3_0_n11,
         npu_inst_pe_1_3_0_n10, npu_inst_pe_1_3_0_n9, npu_inst_pe_1_3_0_n8,
         npu_inst_pe_1_3_0_n7, npu_inst_pe_1_3_0_n6, npu_inst_pe_1_3_0_n5,
         npu_inst_pe_1_3_0_n4, npu_inst_pe_1_3_0_n3, npu_inst_pe_1_3_0_n2,
         npu_inst_pe_1_3_0_n1, npu_inst_pe_1_3_0_sub_77_carry_7_,
         npu_inst_pe_1_3_0_sub_77_carry_6_, npu_inst_pe_1_3_0_sub_77_carry_5_,
         npu_inst_pe_1_3_0_sub_77_carry_4_, npu_inst_pe_1_3_0_sub_77_carry_3_,
         npu_inst_pe_1_3_0_sub_77_carry_2_, npu_inst_pe_1_3_0_sub_77_carry_1_,
         npu_inst_pe_1_3_0_add_79_carry_7_, npu_inst_pe_1_3_0_add_79_carry_6_,
         npu_inst_pe_1_3_0_add_79_carry_5_, npu_inst_pe_1_3_0_add_79_carry_4_,
         npu_inst_pe_1_3_0_add_79_carry_3_, npu_inst_pe_1_3_0_add_79_carry_2_,
         npu_inst_pe_1_3_0_add_79_carry_1_, npu_inst_pe_1_3_0_n97,
         npu_inst_pe_1_3_0_n96, npu_inst_pe_1_3_0_n95, npu_inst_pe_1_3_0_n94,
         npu_inst_pe_1_3_0_n93, npu_inst_pe_1_3_0_n92, npu_inst_pe_1_3_0_n91,
         npu_inst_pe_1_3_0_n90, npu_inst_pe_1_3_0_n89, npu_inst_pe_1_3_0_n88,
         npu_inst_pe_1_3_0_n87, npu_inst_pe_1_3_0_n86, npu_inst_pe_1_3_0_n85,
         npu_inst_pe_1_3_0_n84, npu_inst_pe_1_3_0_n83, npu_inst_pe_1_3_0_n82,
         npu_inst_pe_1_3_0_n81, npu_inst_pe_1_3_0_n80, npu_inst_pe_1_3_0_n79,
         npu_inst_pe_1_3_0_n78, npu_inst_pe_1_3_0_n77, npu_inst_pe_1_3_0_n76,
         npu_inst_pe_1_3_0_n75, npu_inst_pe_1_3_0_n74, npu_inst_pe_1_3_0_n73,
         npu_inst_pe_1_3_0_n72, npu_inst_pe_1_3_0_n71, npu_inst_pe_1_3_0_n70,
         npu_inst_pe_1_3_0_n69, npu_inst_pe_1_3_0_n68, npu_inst_pe_1_3_0_n67,
         npu_inst_pe_1_3_0_n66, npu_inst_pe_1_3_0_n65, npu_inst_pe_1_3_0_n64,
         npu_inst_pe_1_3_0_n63, npu_inst_pe_1_3_0_n62, npu_inst_pe_1_3_0_n61,
         npu_inst_pe_1_3_0_n60, npu_inst_pe_1_3_0_n59, npu_inst_pe_1_3_0_n58,
         npu_inst_pe_1_3_0_n57, npu_inst_pe_1_3_0_n56, npu_inst_pe_1_3_0_n55,
         npu_inst_pe_1_3_0_n54, npu_inst_pe_1_3_0_n53, npu_inst_pe_1_3_0_n52,
         npu_inst_pe_1_3_0_n51, npu_inst_pe_1_3_0_n50, npu_inst_pe_1_3_0_n49,
         npu_inst_pe_1_3_0_n48, npu_inst_pe_1_3_0_n47, npu_inst_pe_1_3_0_n46,
         npu_inst_pe_1_3_0_n45, npu_inst_pe_1_3_0_n44, npu_inst_pe_1_3_0_n43,
         npu_inst_pe_1_3_0_n42, npu_inst_pe_1_3_0_n41, npu_inst_pe_1_3_0_n40,
         npu_inst_pe_1_3_0_n39, npu_inst_pe_1_3_0_n38, npu_inst_pe_1_3_0_n37,
         npu_inst_pe_1_3_0_n27, npu_inst_pe_1_3_0_n26,
         npu_inst_pe_1_3_0_net3747, npu_inst_pe_1_3_0_net3741,
         npu_inst_pe_1_3_0_N94, npu_inst_pe_1_3_0_N93, npu_inst_pe_1_3_0_N84,
         npu_inst_pe_1_3_0_N80, npu_inst_pe_1_3_0_N79, npu_inst_pe_1_3_0_N78,
         npu_inst_pe_1_3_0_N77, npu_inst_pe_1_3_0_N76, npu_inst_pe_1_3_0_N75,
         npu_inst_pe_1_3_0_N74, npu_inst_pe_1_3_0_N73, npu_inst_pe_1_3_0_N72,
         npu_inst_pe_1_3_0_N71, npu_inst_pe_1_3_0_N70, npu_inst_pe_1_3_0_N69,
         npu_inst_pe_1_3_0_N68, npu_inst_pe_1_3_0_N67, npu_inst_pe_1_3_0_N66,
         npu_inst_pe_1_3_0_N65, npu_inst_pe_1_3_0_int_q_acc_0_,
         npu_inst_pe_1_3_0_int_q_acc_1_, npu_inst_pe_1_3_0_int_q_acc_2_,
         npu_inst_pe_1_3_0_int_q_acc_3_, npu_inst_pe_1_3_0_int_q_acc_4_,
         npu_inst_pe_1_3_0_int_q_acc_5_, npu_inst_pe_1_3_0_int_q_acc_6_,
         npu_inst_pe_1_3_0_int_q_acc_7_, npu_inst_pe_1_3_0_int_data_0_,
         npu_inst_pe_1_3_0_int_data_1_, npu_inst_pe_1_3_0_int_q_weight_0_,
         npu_inst_pe_1_3_0_int_q_weight_1_,
         npu_inst_pe_1_3_0_int_q_reg_v_5__0_,
         npu_inst_pe_1_3_0_int_q_reg_v_5__1_,
         npu_inst_pe_1_3_0_int_q_reg_v_4__0_,
         npu_inst_pe_1_3_0_int_q_reg_v_4__1_,
         npu_inst_pe_1_3_0_int_q_reg_v_3__0_,
         npu_inst_pe_1_3_0_int_q_reg_v_3__1_,
         npu_inst_pe_1_3_0_int_q_reg_v_2__0_,
         npu_inst_pe_1_3_0_int_q_reg_v_2__1_,
         npu_inst_pe_1_3_0_int_q_reg_v_1__0_,
         npu_inst_pe_1_3_0_int_q_reg_v_1__1_,
         npu_inst_pe_1_3_0_int_q_reg_v_0__0_,
         npu_inst_pe_1_3_0_int_q_reg_v_0__1_,
         npu_inst_pe_1_3_0_int_q_reg_h_5__0_,
         npu_inst_pe_1_3_0_int_q_reg_h_5__1_,
         npu_inst_pe_1_3_0_int_q_reg_h_4__0_,
         npu_inst_pe_1_3_0_int_q_reg_h_4__1_,
         npu_inst_pe_1_3_0_int_q_reg_h_3__0_,
         npu_inst_pe_1_3_0_int_q_reg_h_3__1_,
         npu_inst_pe_1_3_0_int_q_reg_h_2__0_,
         npu_inst_pe_1_3_0_int_q_reg_h_2__1_,
         npu_inst_pe_1_3_0_int_q_reg_h_1__0_,
         npu_inst_pe_1_3_0_int_q_reg_h_1__1_,
         npu_inst_pe_1_3_0_int_q_reg_h_0__0_,
         npu_inst_pe_1_3_0_int_q_reg_h_0__1_, npu_inst_pe_1_3_0_o_data_h_0_,
         npu_inst_pe_1_3_0_o_data_h_1_, npu_inst_pe_1_3_1_n119,
         npu_inst_pe_1_3_1_n118, npu_inst_pe_1_3_1_n117,
         npu_inst_pe_1_3_1_n116, npu_inst_pe_1_3_1_n115,
         npu_inst_pe_1_3_1_n114, npu_inst_pe_1_3_1_n113,
         npu_inst_pe_1_3_1_n112, npu_inst_pe_1_3_1_n111,
         npu_inst_pe_1_3_1_n110, npu_inst_pe_1_3_1_n109,
         npu_inst_pe_1_3_1_n108, npu_inst_pe_1_3_1_n107,
         npu_inst_pe_1_3_1_n106, npu_inst_pe_1_3_1_n105,
         npu_inst_pe_1_3_1_n104, npu_inst_pe_1_3_1_n103,
         npu_inst_pe_1_3_1_n102, npu_inst_pe_1_3_1_n101,
         npu_inst_pe_1_3_1_n100, npu_inst_pe_1_3_1_n99, npu_inst_pe_1_3_1_n98,
         npu_inst_pe_1_3_1_n36, npu_inst_pe_1_3_1_n35, npu_inst_pe_1_3_1_n34,
         npu_inst_pe_1_3_1_n33, npu_inst_pe_1_3_1_n32, npu_inst_pe_1_3_1_n31,
         npu_inst_pe_1_3_1_n30, npu_inst_pe_1_3_1_n29, npu_inst_pe_1_3_1_n28,
         npu_inst_pe_1_3_1_n25, npu_inst_pe_1_3_1_n24, npu_inst_pe_1_3_1_n23,
         npu_inst_pe_1_3_1_n22, npu_inst_pe_1_3_1_n21, npu_inst_pe_1_3_1_n20,
         npu_inst_pe_1_3_1_n19, npu_inst_pe_1_3_1_n18, npu_inst_pe_1_3_1_n17,
         npu_inst_pe_1_3_1_n16, npu_inst_pe_1_3_1_n15, npu_inst_pe_1_3_1_n14,
         npu_inst_pe_1_3_1_n13, npu_inst_pe_1_3_1_n12, npu_inst_pe_1_3_1_n11,
         npu_inst_pe_1_3_1_n10, npu_inst_pe_1_3_1_n9, npu_inst_pe_1_3_1_n8,
         npu_inst_pe_1_3_1_n7, npu_inst_pe_1_3_1_n6, npu_inst_pe_1_3_1_n5,
         npu_inst_pe_1_3_1_n4, npu_inst_pe_1_3_1_n3, npu_inst_pe_1_3_1_n2,
         npu_inst_pe_1_3_1_n1, npu_inst_pe_1_3_1_sub_77_carry_7_,
         npu_inst_pe_1_3_1_sub_77_carry_6_, npu_inst_pe_1_3_1_sub_77_carry_5_,
         npu_inst_pe_1_3_1_sub_77_carry_4_, npu_inst_pe_1_3_1_sub_77_carry_3_,
         npu_inst_pe_1_3_1_sub_77_carry_2_, npu_inst_pe_1_3_1_sub_77_carry_1_,
         npu_inst_pe_1_3_1_add_79_carry_7_, npu_inst_pe_1_3_1_add_79_carry_6_,
         npu_inst_pe_1_3_1_add_79_carry_5_, npu_inst_pe_1_3_1_add_79_carry_4_,
         npu_inst_pe_1_3_1_add_79_carry_3_, npu_inst_pe_1_3_1_add_79_carry_2_,
         npu_inst_pe_1_3_1_add_79_carry_1_, npu_inst_pe_1_3_1_n97,
         npu_inst_pe_1_3_1_n96, npu_inst_pe_1_3_1_n95, npu_inst_pe_1_3_1_n94,
         npu_inst_pe_1_3_1_n93, npu_inst_pe_1_3_1_n92, npu_inst_pe_1_3_1_n91,
         npu_inst_pe_1_3_1_n90, npu_inst_pe_1_3_1_n89, npu_inst_pe_1_3_1_n88,
         npu_inst_pe_1_3_1_n87, npu_inst_pe_1_3_1_n86, npu_inst_pe_1_3_1_n85,
         npu_inst_pe_1_3_1_n84, npu_inst_pe_1_3_1_n83, npu_inst_pe_1_3_1_n82,
         npu_inst_pe_1_3_1_n81, npu_inst_pe_1_3_1_n80, npu_inst_pe_1_3_1_n79,
         npu_inst_pe_1_3_1_n78, npu_inst_pe_1_3_1_n77, npu_inst_pe_1_3_1_n76,
         npu_inst_pe_1_3_1_n75, npu_inst_pe_1_3_1_n74, npu_inst_pe_1_3_1_n73,
         npu_inst_pe_1_3_1_n72, npu_inst_pe_1_3_1_n71, npu_inst_pe_1_3_1_n70,
         npu_inst_pe_1_3_1_n69, npu_inst_pe_1_3_1_n68, npu_inst_pe_1_3_1_n67,
         npu_inst_pe_1_3_1_n66, npu_inst_pe_1_3_1_n65, npu_inst_pe_1_3_1_n64,
         npu_inst_pe_1_3_1_n63, npu_inst_pe_1_3_1_n62, npu_inst_pe_1_3_1_n61,
         npu_inst_pe_1_3_1_n60, npu_inst_pe_1_3_1_n59, npu_inst_pe_1_3_1_n58,
         npu_inst_pe_1_3_1_n57, npu_inst_pe_1_3_1_n56, npu_inst_pe_1_3_1_n55,
         npu_inst_pe_1_3_1_n54, npu_inst_pe_1_3_1_n53, npu_inst_pe_1_3_1_n52,
         npu_inst_pe_1_3_1_n51, npu_inst_pe_1_3_1_n50, npu_inst_pe_1_3_1_n49,
         npu_inst_pe_1_3_1_n48, npu_inst_pe_1_3_1_n47, npu_inst_pe_1_3_1_n46,
         npu_inst_pe_1_3_1_n45, npu_inst_pe_1_3_1_n44, npu_inst_pe_1_3_1_n43,
         npu_inst_pe_1_3_1_n42, npu_inst_pe_1_3_1_n41, npu_inst_pe_1_3_1_n40,
         npu_inst_pe_1_3_1_n39, npu_inst_pe_1_3_1_n38, npu_inst_pe_1_3_1_n37,
         npu_inst_pe_1_3_1_n27, npu_inst_pe_1_3_1_n26,
         npu_inst_pe_1_3_1_net3724, npu_inst_pe_1_3_1_net3718,
         npu_inst_pe_1_3_1_N94, npu_inst_pe_1_3_1_N93, npu_inst_pe_1_3_1_N84,
         npu_inst_pe_1_3_1_N80, npu_inst_pe_1_3_1_N79, npu_inst_pe_1_3_1_N78,
         npu_inst_pe_1_3_1_N77, npu_inst_pe_1_3_1_N76, npu_inst_pe_1_3_1_N75,
         npu_inst_pe_1_3_1_N74, npu_inst_pe_1_3_1_N73, npu_inst_pe_1_3_1_N72,
         npu_inst_pe_1_3_1_N71, npu_inst_pe_1_3_1_N70, npu_inst_pe_1_3_1_N69,
         npu_inst_pe_1_3_1_N68, npu_inst_pe_1_3_1_N67, npu_inst_pe_1_3_1_N66,
         npu_inst_pe_1_3_1_N65, npu_inst_pe_1_3_1_int_q_acc_0_,
         npu_inst_pe_1_3_1_int_q_acc_1_, npu_inst_pe_1_3_1_int_q_acc_2_,
         npu_inst_pe_1_3_1_int_q_acc_3_, npu_inst_pe_1_3_1_int_q_acc_4_,
         npu_inst_pe_1_3_1_int_q_acc_5_, npu_inst_pe_1_3_1_int_q_acc_6_,
         npu_inst_pe_1_3_1_int_q_acc_7_, npu_inst_pe_1_3_1_int_data_0_,
         npu_inst_pe_1_3_1_int_data_1_, npu_inst_pe_1_3_1_int_q_weight_0_,
         npu_inst_pe_1_3_1_int_q_weight_1_,
         npu_inst_pe_1_3_1_int_q_reg_v_5__0_,
         npu_inst_pe_1_3_1_int_q_reg_v_5__1_,
         npu_inst_pe_1_3_1_int_q_reg_v_4__0_,
         npu_inst_pe_1_3_1_int_q_reg_v_4__1_,
         npu_inst_pe_1_3_1_int_q_reg_v_3__0_,
         npu_inst_pe_1_3_1_int_q_reg_v_3__1_,
         npu_inst_pe_1_3_1_int_q_reg_v_2__0_,
         npu_inst_pe_1_3_1_int_q_reg_v_2__1_,
         npu_inst_pe_1_3_1_int_q_reg_v_1__0_,
         npu_inst_pe_1_3_1_int_q_reg_v_1__1_,
         npu_inst_pe_1_3_1_int_q_reg_v_0__0_,
         npu_inst_pe_1_3_1_int_q_reg_v_0__1_,
         npu_inst_pe_1_3_1_int_q_reg_h_5__0_,
         npu_inst_pe_1_3_1_int_q_reg_h_5__1_,
         npu_inst_pe_1_3_1_int_q_reg_h_4__0_,
         npu_inst_pe_1_3_1_int_q_reg_h_4__1_,
         npu_inst_pe_1_3_1_int_q_reg_h_3__0_,
         npu_inst_pe_1_3_1_int_q_reg_h_3__1_,
         npu_inst_pe_1_3_1_int_q_reg_h_2__0_,
         npu_inst_pe_1_3_1_int_q_reg_h_2__1_,
         npu_inst_pe_1_3_1_int_q_reg_h_1__0_,
         npu_inst_pe_1_3_1_int_q_reg_h_1__1_,
         npu_inst_pe_1_3_1_int_q_reg_h_0__0_,
         npu_inst_pe_1_3_1_int_q_reg_h_0__1_, npu_inst_pe_1_3_2_n119,
         npu_inst_pe_1_3_2_n118, npu_inst_pe_1_3_2_n117,
         npu_inst_pe_1_3_2_n116, npu_inst_pe_1_3_2_n115,
         npu_inst_pe_1_3_2_n114, npu_inst_pe_1_3_2_n113,
         npu_inst_pe_1_3_2_n112, npu_inst_pe_1_3_2_n111,
         npu_inst_pe_1_3_2_n110, npu_inst_pe_1_3_2_n109,
         npu_inst_pe_1_3_2_n108, npu_inst_pe_1_3_2_n107,
         npu_inst_pe_1_3_2_n106, npu_inst_pe_1_3_2_n105,
         npu_inst_pe_1_3_2_n104, npu_inst_pe_1_3_2_n103,
         npu_inst_pe_1_3_2_n102, npu_inst_pe_1_3_2_n101,
         npu_inst_pe_1_3_2_n100, npu_inst_pe_1_3_2_n99, npu_inst_pe_1_3_2_n98,
         npu_inst_pe_1_3_2_n36, npu_inst_pe_1_3_2_n35, npu_inst_pe_1_3_2_n34,
         npu_inst_pe_1_3_2_n33, npu_inst_pe_1_3_2_n32, npu_inst_pe_1_3_2_n31,
         npu_inst_pe_1_3_2_n30, npu_inst_pe_1_3_2_n29, npu_inst_pe_1_3_2_n28,
         npu_inst_pe_1_3_2_n25, npu_inst_pe_1_3_2_n24, npu_inst_pe_1_3_2_n23,
         npu_inst_pe_1_3_2_n22, npu_inst_pe_1_3_2_n21, npu_inst_pe_1_3_2_n20,
         npu_inst_pe_1_3_2_n19, npu_inst_pe_1_3_2_n18, npu_inst_pe_1_3_2_n17,
         npu_inst_pe_1_3_2_n16, npu_inst_pe_1_3_2_n15, npu_inst_pe_1_3_2_n14,
         npu_inst_pe_1_3_2_n13, npu_inst_pe_1_3_2_n12, npu_inst_pe_1_3_2_n11,
         npu_inst_pe_1_3_2_n10, npu_inst_pe_1_3_2_n9, npu_inst_pe_1_3_2_n8,
         npu_inst_pe_1_3_2_n7, npu_inst_pe_1_3_2_n6, npu_inst_pe_1_3_2_n5,
         npu_inst_pe_1_3_2_n4, npu_inst_pe_1_3_2_n3, npu_inst_pe_1_3_2_n2,
         npu_inst_pe_1_3_2_n1, npu_inst_pe_1_3_2_sub_77_carry_7_,
         npu_inst_pe_1_3_2_sub_77_carry_6_, npu_inst_pe_1_3_2_sub_77_carry_5_,
         npu_inst_pe_1_3_2_sub_77_carry_4_, npu_inst_pe_1_3_2_sub_77_carry_3_,
         npu_inst_pe_1_3_2_sub_77_carry_2_, npu_inst_pe_1_3_2_sub_77_carry_1_,
         npu_inst_pe_1_3_2_add_79_carry_7_, npu_inst_pe_1_3_2_add_79_carry_6_,
         npu_inst_pe_1_3_2_add_79_carry_5_, npu_inst_pe_1_3_2_add_79_carry_4_,
         npu_inst_pe_1_3_2_add_79_carry_3_, npu_inst_pe_1_3_2_add_79_carry_2_,
         npu_inst_pe_1_3_2_add_79_carry_1_, npu_inst_pe_1_3_2_n97,
         npu_inst_pe_1_3_2_n96, npu_inst_pe_1_3_2_n95, npu_inst_pe_1_3_2_n94,
         npu_inst_pe_1_3_2_n93, npu_inst_pe_1_3_2_n92, npu_inst_pe_1_3_2_n91,
         npu_inst_pe_1_3_2_n90, npu_inst_pe_1_3_2_n89, npu_inst_pe_1_3_2_n88,
         npu_inst_pe_1_3_2_n87, npu_inst_pe_1_3_2_n86, npu_inst_pe_1_3_2_n85,
         npu_inst_pe_1_3_2_n84, npu_inst_pe_1_3_2_n83, npu_inst_pe_1_3_2_n82,
         npu_inst_pe_1_3_2_n81, npu_inst_pe_1_3_2_n80, npu_inst_pe_1_3_2_n79,
         npu_inst_pe_1_3_2_n78, npu_inst_pe_1_3_2_n77, npu_inst_pe_1_3_2_n76,
         npu_inst_pe_1_3_2_n75, npu_inst_pe_1_3_2_n74, npu_inst_pe_1_3_2_n73,
         npu_inst_pe_1_3_2_n72, npu_inst_pe_1_3_2_n71, npu_inst_pe_1_3_2_n70,
         npu_inst_pe_1_3_2_n69, npu_inst_pe_1_3_2_n68, npu_inst_pe_1_3_2_n67,
         npu_inst_pe_1_3_2_n66, npu_inst_pe_1_3_2_n65, npu_inst_pe_1_3_2_n64,
         npu_inst_pe_1_3_2_n63, npu_inst_pe_1_3_2_n62, npu_inst_pe_1_3_2_n61,
         npu_inst_pe_1_3_2_n60, npu_inst_pe_1_3_2_n59, npu_inst_pe_1_3_2_n58,
         npu_inst_pe_1_3_2_n57, npu_inst_pe_1_3_2_n56, npu_inst_pe_1_3_2_n55,
         npu_inst_pe_1_3_2_n54, npu_inst_pe_1_3_2_n53, npu_inst_pe_1_3_2_n52,
         npu_inst_pe_1_3_2_n51, npu_inst_pe_1_3_2_n50, npu_inst_pe_1_3_2_n49,
         npu_inst_pe_1_3_2_n48, npu_inst_pe_1_3_2_n47, npu_inst_pe_1_3_2_n46,
         npu_inst_pe_1_3_2_n45, npu_inst_pe_1_3_2_n44, npu_inst_pe_1_3_2_n43,
         npu_inst_pe_1_3_2_n42, npu_inst_pe_1_3_2_n41, npu_inst_pe_1_3_2_n40,
         npu_inst_pe_1_3_2_n39, npu_inst_pe_1_3_2_n38, npu_inst_pe_1_3_2_n37,
         npu_inst_pe_1_3_2_n27, npu_inst_pe_1_3_2_n26,
         npu_inst_pe_1_3_2_net3701, npu_inst_pe_1_3_2_net3695,
         npu_inst_pe_1_3_2_N94, npu_inst_pe_1_3_2_N93, npu_inst_pe_1_3_2_N84,
         npu_inst_pe_1_3_2_N80, npu_inst_pe_1_3_2_N79, npu_inst_pe_1_3_2_N78,
         npu_inst_pe_1_3_2_N77, npu_inst_pe_1_3_2_N76, npu_inst_pe_1_3_2_N75,
         npu_inst_pe_1_3_2_N74, npu_inst_pe_1_3_2_N73, npu_inst_pe_1_3_2_N72,
         npu_inst_pe_1_3_2_N71, npu_inst_pe_1_3_2_N70, npu_inst_pe_1_3_2_N69,
         npu_inst_pe_1_3_2_N68, npu_inst_pe_1_3_2_N67, npu_inst_pe_1_3_2_N66,
         npu_inst_pe_1_3_2_N65, npu_inst_pe_1_3_2_int_q_acc_0_,
         npu_inst_pe_1_3_2_int_q_acc_1_, npu_inst_pe_1_3_2_int_q_acc_2_,
         npu_inst_pe_1_3_2_int_q_acc_3_, npu_inst_pe_1_3_2_int_q_acc_4_,
         npu_inst_pe_1_3_2_int_q_acc_5_, npu_inst_pe_1_3_2_int_q_acc_6_,
         npu_inst_pe_1_3_2_int_q_acc_7_, npu_inst_pe_1_3_2_int_data_0_,
         npu_inst_pe_1_3_2_int_data_1_, npu_inst_pe_1_3_2_int_q_weight_0_,
         npu_inst_pe_1_3_2_int_q_weight_1_,
         npu_inst_pe_1_3_2_int_q_reg_v_5__0_,
         npu_inst_pe_1_3_2_int_q_reg_v_5__1_,
         npu_inst_pe_1_3_2_int_q_reg_v_4__0_,
         npu_inst_pe_1_3_2_int_q_reg_v_4__1_,
         npu_inst_pe_1_3_2_int_q_reg_v_3__0_,
         npu_inst_pe_1_3_2_int_q_reg_v_3__1_,
         npu_inst_pe_1_3_2_int_q_reg_v_2__0_,
         npu_inst_pe_1_3_2_int_q_reg_v_2__1_,
         npu_inst_pe_1_3_2_int_q_reg_v_1__0_,
         npu_inst_pe_1_3_2_int_q_reg_v_1__1_,
         npu_inst_pe_1_3_2_int_q_reg_v_0__0_,
         npu_inst_pe_1_3_2_int_q_reg_v_0__1_,
         npu_inst_pe_1_3_2_int_q_reg_h_5__0_,
         npu_inst_pe_1_3_2_int_q_reg_h_5__1_,
         npu_inst_pe_1_3_2_int_q_reg_h_4__0_,
         npu_inst_pe_1_3_2_int_q_reg_h_4__1_,
         npu_inst_pe_1_3_2_int_q_reg_h_3__0_,
         npu_inst_pe_1_3_2_int_q_reg_h_3__1_,
         npu_inst_pe_1_3_2_int_q_reg_h_2__0_,
         npu_inst_pe_1_3_2_int_q_reg_h_2__1_,
         npu_inst_pe_1_3_2_int_q_reg_h_1__0_,
         npu_inst_pe_1_3_2_int_q_reg_h_1__1_,
         npu_inst_pe_1_3_2_int_q_reg_h_0__0_,
         npu_inst_pe_1_3_2_int_q_reg_h_0__1_, npu_inst_pe_1_3_3_n119,
         npu_inst_pe_1_3_3_n118, npu_inst_pe_1_3_3_n117,
         npu_inst_pe_1_3_3_n116, npu_inst_pe_1_3_3_n115,
         npu_inst_pe_1_3_3_n114, npu_inst_pe_1_3_3_n113,
         npu_inst_pe_1_3_3_n112, npu_inst_pe_1_3_3_n111,
         npu_inst_pe_1_3_3_n110, npu_inst_pe_1_3_3_n109,
         npu_inst_pe_1_3_3_n108, npu_inst_pe_1_3_3_n107,
         npu_inst_pe_1_3_3_n106, npu_inst_pe_1_3_3_n105,
         npu_inst_pe_1_3_3_n104, npu_inst_pe_1_3_3_n103,
         npu_inst_pe_1_3_3_n102, npu_inst_pe_1_3_3_n101,
         npu_inst_pe_1_3_3_n100, npu_inst_pe_1_3_3_n99, npu_inst_pe_1_3_3_n98,
         npu_inst_pe_1_3_3_n36, npu_inst_pe_1_3_3_n35, npu_inst_pe_1_3_3_n34,
         npu_inst_pe_1_3_3_n33, npu_inst_pe_1_3_3_n32, npu_inst_pe_1_3_3_n31,
         npu_inst_pe_1_3_3_n30, npu_inst_pe_1_3_3_n29, npu_inst_pe_1_3_3_n28,
         npu_inst_pe_1_3_3_n25, npu_inst_pe_1_3_3_n24, npu_inst_pe_1_3_3_n23,
         npu_inst_pe_1_3_3_n22, npu_inst_pe_1_3_3_n21, npu_inst_pe_1_3_3_n20,
         npu_inst_pe_1_3_3_n19, npu_inst_pe_1_3_3_n18, npu_inst_pe_1_3_3_n17,
         npu_inst_pe_1_3_3_n16, npu_inst_pe_1_3_3_n15, npu_inst_pe_1_3_3_n14,
         npu_inst_pe_1_3_3_n13, npu_inst_pe_1_3_3_n12, npu_inst_pe_1_3_3_n11,
         npu_inst_pe_1_3_3_n10, npu_inst_pe_1_3_3_n9, npu_inst_pe_1_3_3_n8,
         npu_inst_pe_1_3_3_n7, npu_inst_pe_1_3_3_n6, npu_inst_pe_1_3_3_n5,
         npu_inst_pe_1_3_3_n4, npu_inst_pe_1_3_3_n3, npu_inst_pe_1_3_3_n2,
         npu_inst_pe_1_3_3_n1, npu_inst_pe_1_3_3_sub_77_carry_7_,
         npu_inst_pe_1_3_3_sub_77_carry_6_, npu_inst_pe_1_3_3_sub_77_carry_5_,
         npu_inst_pe_1_3_3_sub_77_carry_4_, npu_inst_pe_1_3_3_sub_77_carry_3_,
         npu_inst_pe_1_3_3_sub_77_carry_2_, npu_inst_pe_1_3_3_sub_77_carry_1_,
         npu_inst_pe_1_3_3_add_79_carry_7_, npu_inst_pe_1_3_3_add_79_carry_6_,
         npu_inst_pe_1_3_3_add_79_carry_5_, npu_inst_pe_1_3_3_add_79_carry_4_,
         npu_inst_pe_1_3_3_add_79_carry_3_, npu_inst_pe_1_3_3_add_79_carry_2_,
         npu_inst_pe_1_3_3_add_79_carry_1_, npu_inst_pe_1_3_3_n97,
         npu_inst_pe_1_3_3_n96, npu_inst_pe_1_3_3_n95, npu_inst_pe_1_3_3_n94,
         npu_inst_pe_1_3_3_n93, npu_inst_pe_1_3_3_n92, npu_inst_pe_1_3_3_n91,
         npu_inst_pe_1_3_3_n90, npu_inst_pe_1_3_3_n89, npu_inst_pe_1_3_3_n88,
         npu_inst_pe_1_3_3_n87, npu_inst_pe_1_3_3_n86, npu_inst_pe_1_3_3_n85,
         npu_inst_pe_1_3_3_n84, npu_inst_pe_1_3_3_n83, npu_inst_pe_1_3_3_n82,
         npu_inst_pe_1_3_3_n81, npu_inst_pe_1_3_3_n80, npu_inst_pe_1_3_3_n79,
         npu_inst_pe_1_3_3_n78, npu_inst_pe_1_3_3_n77, npu_inst_pe_1_3_3_n76,
         npu_inst_pe_1_3_3_n75, npu_inst_pe_1_3_3_n74, npu_inst_pe_1_3_3_n73,
         npu_inst_pe_1_3_3_n72, npu_inst_pe_1_3_3_n71, npu_inst_pe_1_3_3_n70,
         npu_inst_pe_1_3_3_n69, npu_inst_pe_1_3_3_n68, npu_inst_pe_1_3_3_n67,
         npu_inst_pe_1_3_3_n66, npu_inst_pe_1_3_3_n65, npu_inst_pe_1_3_3_n64,
         npu_inst_pe_1_3_3_n63, npu_inst_pe_1_3_3_n62, npu_inst_pe_1_3_3_n61,
         npu_inst_pe_1_3_3_n60, npu_inst_pe_1_3_3_n59, npu_inst_pe_1_3_3_n58,
         npu_inst_pe_1_3_3_n57, npu_inst_pe_1_3_3_n56, npu_inst_pe_1_3_3_n55,
         npu_inst_pe_1_3_3_n54, npu_inst_pe_1_3_3_n53, npu_inst_pe_1_3_3_n52,
         npu_inst_pe_1_3_3_n51, npu_inst_pe_1_3_3_n50, npu_inst_pe_1_3_3_n49,
         npu_inst_pe_1_3_3_n48, npu_inst_pe_1_3_3_n47, npu_inst_pe_1_3_3_n46,
         npu_inst_pe_1_3_3_n45, npu_inst_pe_1_3_3_n44, npu_inst_pe_1_3_3_n43,
         npu_inst_pe_1_3_3_n42, npu_inst_pe_1_3_3_n41, npu_inst_pe_1_3_3_n40,
         npu_inst_pe_1_3_3_n39, npu_inst_pe_1_3_3_n38, npu_inst_pe_1_3_3_n37,
         npu_inst_pe_1_3_3_n27, npu_inst_pe_1_3_3_n26,
         npu_inst_pe_1_3_3_net3678, npu_inst_pe_1_3_3_net3672,
         npu_inst_pe_1_3_3_N94, npu_inst_pe_1_3_3_N93, npu_inst_pe_1_3_3_N84,
         npu_inst_pe_1_3_3_N80, npu_inst_pe_1_3_3_N79, npu_inst_pe_1_3_3_N78,
         npu_inst_pe_1_3_3_N77, npu_inst_pe_1_3_3_N76, npu_inst_pe_1_3_3_N75,
         npu_inst_pe_1_3_3_N74, npu_inst_pe_1_3_3_N73, npu_inst_pe_1_3_3_N72,
         npu_inst_pe_1_3_3_N71, npu_inst_pe_1_3_3_N70, npu_inst_pe_1_3_3_N69,
         npu_inst_pe_1_3_3_N68, npu_inst_pe_1_3_3_N67, npu_inst_pe_1_3_3_N66,
         npu_inst_pe_1_3_3_N65, npu_inst_pe_1_3_3_int_q_acc_0_,
         npu_inst_pe_1_3_3_int_q_acc_1_, npu_inst_pe_1_3_3_int_q_acc_2_,
         npu_inst_pe_1_3_3_int_q_acc_3_, npu_inst_pe_1_3_3_int_q_acc_4_,
         npu_inst_pe_1_3_3_int_q_acc_5_, npu_inst_pe_1_3_3_int_q_acc_6_,
         npu_inst_pe_1_3_3_int_q_acc_7_, npu_inst_pe_1_3_3_int_data_0_,
         npu_inst_pe_1_3_3_int_data_1_, npu_inst_pe_1_3_3_int_q_weight_0_,
         npu_inst_pe_1_3_3_int_q_weight_1_,
         npu_inst_pe_1_3_3_int_q_reg_v_5__0_,
         npu_inst_pe_1_3_3_int_q_reg_v_5__1_,
         npu_inst_pe_1_3_3_int_q_reg_v_4__0_,
         npu_inst_pe_1_3_3_int_q_reg_v_4__1_,
         npu_inst_pe_1_3_3_int_q_reg_v_3__0_,
         npu_inst_pe_1_3_3_int_q_reg_v_3__1_,
         npu_inst_pe_1_3_3_int_q_reg_v_2__0_,
         npu_inst_pe_1_3_3_int_q_reg_v_2__1_,
         npu_inst_pe_1_3_3_int_q_reg_v_1__0_,
         npu_inst_pe_1_3_3_int_q_reg_v_1__1_,
         npu_inst_pe_1_3_3_int_q_reg_v_0__0_,
         npu_inst_pe_1_3_3_int_q_reg_v_0__1_,
         npu_inst_pe_1_3_3_int_q_reg_h_5__0_,
         npu_inst_pe_1_3_3_int_q_reg_h_5__1_,
         npu_inst_pe_1_3_3_int_q_reg_h_4__0_,
         npu_inst_pe_1_3_3_int_q_reg_h_4__1_,
         npu_inst_pe_1_3_3_int_q_reg_h_3__0_,
         npu_inst_pe_1_3_3_int_q_reg_h_3__1_,
         npu_inst_pe_1_3_3_int_q_reg_h_2__0_,
         npu_inst_pe_1_3_3_int_q_reg_h_2__1_,
         npu_inst_pe_1_3_3_int_q_reg_h_1__0_,
         npu_inst_pe_1_3_3_int_q_reg_h_1__1_,
         npu_inst_pe_1_3_3_int_q_reg_h_0__0_,
         npu_inst_pe_1_3_3_int_q_reg_h_0__1_, npu_inst_pe_1_3_4_n118,
         npu_inst_pe_1_3_4_n117, npu_inst_pe_1_3_4_n116,
         npu_inst_pe_1_3_4_n115, npu_inst_pe_1_3_4_n114,
         npu_inst_pe_1_3_4_n113, npu_inst_pe_1_3_4_n112,
         npu_inst_pe_1_3_4_n111, npu_inst_pe_1_3_4_n110,
         npu_inst_pe_1_3_4_n109, npu_inst_pe_1_3_4_n108,
         npu_inst_pe_1_3_4_n107, npu_inst_pe_1_3_4_n106,
         npu_inst_pe_1_3_4_n105, npu_inst_pe_1_3_4_n104,
         npu_inst_pe_1_3_4_n103, npu_inst_pe_1_3_4_n102,
         npu_inst_pe_1_3_4_n101, npu_inst_pe_1_3_4_n100, npu_inst_pe_1_3_4_n99,
         npu_inst_pe_1_3_4_n98, npu_inst_pe_1_3_4_n36, npu_inst_pe_1_3_4_n35,
         npu_inst_pe_1_3_4_n34, npu_inst_pe_1_3_4_n33, npu_inst_pe_1_3_4_n32,
         npu_inst_pe_1_3_4_n31, npu_inst_pe_1_3_4_n30, npu_inst_pe_1_3_4_n29,
         npu_inst_pe_1_3_4_n28, npu_inst_pe_1_3_4_n25, npu_inst_pe_1_3_4_n24,
         npu_inst_pe_1_3_4_n23, npu_inst_pe_1_3_4_n22, npu_inst_pe_1_3_4_n21,
         npu_inst_pe_1_3_4_n20, npu_inst_pe_1_3_4_n19, npu_inst_pe_1_3_4_n18,
         npu_inst_pe_1_3_4_n17, npu_inst_pe_1_3_4_n16, npu_inst_pe_1_3_4_n15,
         npu_inst_pe_1_3_4_n14, npu_inst_pe_1_3_4_n13, npu_inst_pe_1_3_4_n12,
         npu_inst_pe_1_3_4_n11, npu_inst_pe_1_3_4_n10, npu_inst_pe_1_3_4_n9,
         npu_inst_pe_1_3_4_n8, npu_inst_pe_1_3_4_n7, npu_inst_pe_1_3_4_n6,
         npu_inst_pe_1_3_4_n5, npu_inst_pe_1_3_4_n4, npu_inst_pe_1_3_4_n3,
         npu_inst_pe_1_3_4_n2, npu_inst_pe_1_3_4_n1,
         npu_inst_pe_1_3_4_sub_77_carry_7_, npu_inst_pe_1_3_4_sub_77_carry_6_,
         npu_inst_pe_1_3_4_sub_77_carry_5_, npu_inst_pe_1_3_4_sub_77_carry_4_,
         npu_inst_pe_1_3_4_sub_77_carry_3_, npu_inst_pe_1_3_4_sub_77_carry_2_,
         npu_inst_pe_1_3_4_sub_77_carry_1_, npu_inst_pe_1_3_4_add_79_carry_7_,
         npu_inst_pe_1_3_4_add_79_carry_6_, npu_inst_pe_1_3_4_add_79_carry_5_,
         npu_inst_pe_1_3_4_add_79_carry_4_, npu_inst_pe_1_3_4_add_79_carry_3_,
         npu_inst_pe_1_3_4_add_79_carry_2_, npu_inst_pe_1_3_4_add_79_carry_1_,
         npu_inst_pe_1_3_4_n97, npu_inst_pe_1_3_4_n96, npu_inst_pe_1_3_4_n95,
         npu_inst_pe_1_3_4_n94, npu_inst_pe_1_3_4_n93, npu_inst_pe_1_3_4_n92,
         npu_inst_pe_1_3_4_n91, npu_inst_pe_1_3_4_n90, npu_inst_pe_1_3_4_n89,
         npu_inst_pe_1_3_4_n88, npu_inst_pe_1_3_4_n87, npu_inst_pe_1_3_4_n86,
         npu_inst_pe_1_3_4_n85, npu_inst_pe_1_3_4_n84, npu_inst_pe_1_3_4_n83,
         npu_inst_pe_1_3_4_n82, npu_inst_pe_1_3_4_n81, npu_inst_pe_1_3_4_n80,
         npu_inst_pe_1_3_4_n79, npu_inst_pe_1_3_4_n78, npu_inst_pe_1_3_4_n77,
         npu_inst_pe_1_3_4_n76, npu_inst_pe_1_3_4_n75, npu_inst_pe_1_3_4_n74,
         npu_inst_pe_1_3_4_n73, npu_inst_pe_1_3_4_n72, npu_inst_pe_1_3_4_n71,
         npu_inst_pe_1_3_4_n70, npu_inst_pe_1_3_4_n69, npu_inst_pe_1_3_4_n68,
         npu_inst_pe_1_3_4_n67, npu_inst_pe_1_3_4_n66, npu_inst_pe_1_3_4_n65,
         npu_inst_pe_1_3_4_n64, npu_inst_pe_1_3_4_n63, npu_inst_pe_1_3_4_n62,
         npu_inst_pe_1_3_4_n61, npu_inst_pe_1_3_4_n60, npu_inst_pe_1_3_4_n59,
         npu_inst_pe_1_3_4_n58, npu_inst_pe_1_3_4_n57, npu_inst_pe_1_3_4_n56,
         npu_inst_pe_1_3_4_n55, npu_inst_pe_1_3_4_n54, npu_inst_pe_1_3_4_n53,
         npu_inst_pe_1_3_4_n52, npu_inst_pe_1_3_4_n51, npu_inst_pe_1_3_4_n50,
         npu_inst_pe_1_3_4_n49, npu_inst_pe_1_3_4_n48, npu_inst_pe_1_3_4_n47,
         npu_inst_pe_1_3_4_n46, npu_inst_pe_1_3_4_n45, npu_inst_pe_1_3_4_n44,
         npu_inst_pe_1_3_4_n43, npu_inst_pe_1_3_4_n42, npu_inst_pe_1_3_4_n41,
         npu_inst_pe_1_3_4_n40, npu_inst_pe_1_3_4_n39, npu_inst_pe_1_3_4_n38,
         npu_inst_pe_1_3_4_n37, npu_inst_pe_1_3_4_n27, npu_inst_pe_1_3_4_n26,
         npu_inst_pe_1_3_4_net3655, npu_inst_pe_1_3_4_net3649,
         npu_inst_pe_1_3_4_N94, npu_inst_pe_1_3_4_N93, npu_inst_pe_1_3_4_N84,
         npu_inst_pe_1_3_4_N80, npu_inst_pe_1_3_4_N79, npu_inst_pe_1_3_4_N78,
         npu_inst_pe_1_3_4_N77, npu_inst_pe_1_3_4_N76, npu_inst_pe_1_3_4_N75,
         npu_inst_pe_1_3_4_N74, npu_inst_pe_1_3_4_N73, npu_inst_pe_1_3_4_N72,
         npu_inst_pe_1_3_4_N71, npu_inst_pe_1_3_4_N70, npu_inst_pe_1_3_4_N69,
         npu_inst_pe_1_3_4_N68, npu_inst_pe_1_3_4_N67, npu_inst_pe_1_3_4_N66,
         npu_inst_pe_1_3_4_N65, npu_inst_pe_1_3_4_int_q_acc_0_,
         npu_inst_pe_1_3_4_int_q_acc_1_, npu_inst_pe_1_3_4_int_q_acc_2_,
         npu_inst_pe_1_3_4_int_q_acc_3_, npu_inst_pe_1_3_4_int_q_acc_4_,
         npu_inst_pe_1_3_4_int_q_acc_5_, npu_inst_pe_1_3_4_int_q_acc_6_,
         npu_inst_pe_1_3_4_int_q_acc_7_, npu_inst_pe_1_3_4_int_data_0_,
         npu_inst_pe_1_3_4_int_data_1_, npu_inst_pe_1_3_4_int_q_weight_0_,
         npu_inst_pe_1_3_4_int_q_weight_1_,
         npu_inst_pe_1_3_4_int_q_reg_v_5__0_,
         npu_inst_pe_1_3_4_int_q_reg_v_5__1_,
         npu_inst_pe_1_3_4_int_q_reg_v_4__0_,
         npu_inst_pe_1_3_4_int_q_reg_v_4__1_,
         npu_inst_pe_1_3_4_int_q_reg_v_3__0_,
         npu_inst_pe_1_3_4_int_q_reg_v_3__1_,
         npu_inst_pe_1_3_4_int_q_reg_v_2__0_,
         npu_inst_pe_1_3_4_int_q_reg_v_2__1_,
         npu_inst_pe_1_3_4_int_q_reg_v_1__0_,
         npu_inst_pe_1_3_4_int_q_reg_v_1__1_,
         npu_inst_pe_1_3_4_int_q_reg_v_0__0_,
         npu_inst_pe_1_3_4_int_q_reg_v_0__1_,
         npu_inst_pe_1_3_4_int_q_reg_h_5__0_,
         npu_inst_pe_1_3_4_int_q_reg_h_5__1_,
         npu_inst_pe_1_3_4_int_q_reg_h_4__0_,
         npu_inst_pe_1_3_4_int_q_reg_h_4__1_,
         npu_inst_pe_1_3_4_int_q_reg_h_3__0_,
         npu_inst_pe_1_3_4_int_q_reg_h_3__1_,
         npu_inst_pe_1_3_4_int_q_reg_h_2__0_,
         npu_inst_pe_1_3_4_int_q_reg_h_2__1_,
         npu_inst_pe_1_3_4_int_q_reg_h_1__0_,
         npu_inst_pe_1_3_4_int_q_reg_h_1__1_,
         npu_inst_pe_1_3_4_int_q_reg_h_0__0_,
         npu_inst_pe_1_3_4_int_q_reg_h_0__1_, npu_inst_pe_1_3_5_n119,
         npu_inst_pe_1_3_5_n118, npu_inst_pe_1_3_5_n117,
         npu_inst_pe_1_3_5_n116, npu_inst_pe_1_3_5_n115,
         npu_inst_pe_1_3_5_n114, npu_inst_pe_1_3_5_n113,
         npu_inst_pe_1_3_5_n112, npu_inst_pe_1_3_5_n111,
         npu_inst_pe_1_3_5_n110, npu_inst_pe_1_3_5_n109,
         npu_inst_pe_1_3_5_n108, npu_inst_pe_1_3_5_n107,
         npu_inst_pe_1_3_5_n106, npu_inst_pe_1_3_5_n105,
         npu_inst_pe_1_3_5_n104, npu_inst_pe_1_3_5_n103,
         npu_inst_pe_1_3_5_n102, npu_inst_pe_1_3_5_n101,
         npu_inst_pe_1_3_5_n100, npu_inst_pe_1_3_5_n99, npu_inst_pe_1_3_5_n98,
         npu_inst_pe_1_3_5_n36, npu_inst_pe_1_3_5_n35, npu_inst_pe_1_3_5_n34,
         npu_inst_pe_1_3_5_n33, npu_inst_pe_1_3_5_n32, npu_inst_pe_1_3_5_n31,
         npu_inst_pe_1_3_5_n30, npu_inst_pe_1_3_5_n29, npu_inst_pe_1_3_5_n28,
         npu_inst_pe_1_3_5_n25, npu_inst_pe_1_3_5_n24, npu_inst_pe_1_3_5_n23,
         npu_inst_pe_1_3_5_n22, npu_inst_pe_1_3_5_n21, npu_inst_pe_1_3_5_n20,
         npu_inst_pe_1_3_5_n19, npu_inst_pe_1_3_5_n18, npu_inst_pe_1_3_5_n17,
         npu_inst_pe_1_3_5_n16, npu_inst_pe_1_3_5_n15, npu_inst_pe_1_3_5_n14,
         npu_inst_pe_1_3_5_n13, npu_inst_pe_1_3_5_n12, npu_inst_pe_1_3_5_n11,
         npu_inst_pe_1_3_5_n10, npu_inst_pe_1_3_5_n9, npu_inst_pe_1_3_5_n8,
         npu_inst_pe_1_3_5_n7, npu_inst_pe_1_3_5_n6, npu_inst_pe_1_3_5_n5,
         npu_inst_pe_1_3_5_n4, npu_inst_pe_1_3_5_n3, npu_inst_pe_1_3_5_n2,
         npu_inst_pe_1_3_5_n1, npu_inst_pe_1_3_5_sub_77_carry_7_,
         npu_inst_pe_1_3_5_sub_77_carry_6_, npu_inst_pe_1_3_5_sub_77_carry_5_,
         npu_inst_pe_1_3_5_sub_77_carry_4_, npu_inst_pe_1_3_5_sub_77_carry_3_,
         npu_inst_pe_1_3_5_sub_77_carry_2_, npu_inst_pe_1_3_5_sub_77_carry_1_,
         npu_inst_pe_1_3_5_add_79_carry_7_, npu_inst_pe_1_3_5_add_79_carry_6_,
         npu_inst_pe_1_3_5_add_79_carry_5_, npu_inst_pe_1_3_5_add_79_carry_4_,
         npu_inst_pe_1_3_5_add_79_carry_3_, npu_inst_pe_1_3_5_add_79_carry_2_,
         npu_inst_pe_1_3_5_add_79_carry_1_, npu_inst_pe_1_3_5_n97,
         npu_inst_pe_1_3_5_n96, npu_inst_pe_1_3_5_n95, npu_inst_pe_1_3_5_n94,
         npu_inst_pe_1_3_5_n93, npu_inst_pe_1_3_5_n92, npu_inst_pe_1_3_5_n91,
         npu_inst_pe_1_3_5_n90, npu_inst_pe_1_3_5_n89, npu_inst_pe_1_3_5_n88,
         npu_inst_pe_1_3_5_n87, npu_inst_pe_1_3_5_n86, npu_inst_pe_1_3_5_n85,
         npu_inst_pe_1_3_5_n84, npu_inst_pe_1_3_5_n83, npu_inst_pe_1_3_5_n82,
         npu_inst_pe_1_3_5_n81, npu_inst_pe_1_3_5_n80, npu_inst_pe_1_3_5_n79,
         npu_inst_pe_1_3_5_n78, npu_inst_pe_1_3_5_n77, npu_inst_pe_1_3_5_n76,
         npu_inst_pe_1_3_5_n75, npu_inst_pe_1_3_5_n74, npu_inst_pe_1_3_5_n73,
         npu_inst_pe_1_3_5_n72, npu_inst_pe_1_3_5_n71, npu_inst_pe_1_3_5_n70,
         npu_inst_pe_1_3_5_n69, npu_inst_pe_1_3_5_n68, npu_inst_pe_1_3_5_n67,
         npu_inst_pe_1_3_5_n66, npu_inst_pe_1_3_5_n65, npu_inst_pe_1_3_5_n64,
         npu_inst_pe_1_3_5_n63, npu_inst_pe_1_3_5_n62, npu_inst_pe_1_3_5_n61,
         npu_inst_pe_1_3_5_n60, npu_inst_pe_1_3_5_n59, npu_inst_pe_1_3_5_n58,
         npu_inst_pe_1_3_5_n57, npu_inst_pe_1_3_5_n56, npu_inst_pe_1_3_5_n55,
         npu_inst_pe_1_3_5_n54, npu_inst_pe_1_3_5_n53, npu_inst_pe_1_3_5_n52,
         npu_inst_pe_1_3_5_n51, npu_inst_pe_1_3_5_n50, npu_inst_pe_1_3_5_n49,
         npu_inst_pe_1_3_5_n48, npu_inst_pe_1_3_5_n47, npu_inst_pe_1_3_5_n46,
         npu_inst_pe_1_3_5_n45, npu_inst_pe_1_3_5_n44, npu_inst_pe_1_3_5_n43,
         npu_inst_pe_1_3_5_n42, npu_inst_pe_1_3_5_n41, npu_inst_pe_1_3_5_n40,
         npu_inst_pe_1_3_5_n39, npu_inst_pe_1_3_5_n38, npu_inst_pe_1_3_5_n37,
         npu_inst_pe_1_3_5_n27, npu_inst_pe_1_3_5_n26,
         npu_inst_pe_1_3_5_net3632, npu_inst_pe_1_3_5_net3626,
         npu_inst_pe_1_3_5_N94, npu_inst_pe_1_3_5_N93, npu_inst_pe_1_3_5_N84,
         npu_inst_pe_1_3_5_N80, npu_inst_pe_1_3_5_N79, npu_inst_pe_1_3_5_N78,
         npu_inst_pe_1_3_5_N77, npu_inst_pe_1_3_5_N76, npu_inst_pe_1_3_5_N75,
         npu_inst_pe_1_3_5_N74, npu_inst_pe_1_3_5_N73, npu_inst_pe_1_3_5_N72,
         npu_inst_pe_1_3_5_N71, npu_inst_pe_1_3_5_N70, npu_inst_pe_1_3_5_N69,
         npu_inst_pe_1_3_5_N68, npu_inst_pe_1_3_5_N67, npu_inst_pe_1_3_5_N66,
         npu_inst_pe_1_3_5_N65, npu_inst_pe_1_3_5_int_q_acc_0_,
         npu_inst_pe_1_3_5_int_q_acc_1_, npu_inst_pe_1_3_5_int_q_acc_2_,
         npu_inst_pe_1_3_5_int_q_acc_3_, npu_inst_pe_1_3_5_int_q_acc_4_,
         npu_inst_pe_1_3_5_int_q_acc_5_, npu_inst_pe_1_3_5_int_q_acc_6_,
         npu_inst_pe_1_3_5_int_q_acc_7_, npu_inst_pe_1_3_5_int_data_0_,
         npu_inst_pe_1_3_5_int_data_1_, npu_inst_pe_1_3_5_int_q_weight_0_,
         npu_inst_pe_1_3_5_int_q_weight_1_,
         npu_inst_pe_1_3_5_int_q_reg_v_5__0_,
         npu_inst_pe_1_3_5_int_q_reg_v_5__1_,
         npu_inst_pe_1_3_5_int_q_reg_v_4__0_,
         npu_inst_pe_1_3_5_int_q_reg_v_4__1_,
         npu_inst_pe_1_3_5_int_q_reg_v_3__0_,
         npu_inst_pe_1_3_5_int_q_reg_v_3__1_,
         npu_inst_pe_1_3_5_int_q_reg_v_2__0_,
         npu_inst_pe_1_3_5_int_q_reg_v_2__1_,
         npu_inst_pe_1_3_5_int_q_reg_v_1__0_,
         npu_inst_pe_1_3_5_int_q_reg_v_1__1_,
         npu_inst_pe_1_3_5_int_q_reg_v_0__0_,
         npu_inst_pe_1_3_5_int_q_reg_v_0__1_,
         npu_inst_pe_1_3_5_int_q_reg_h_5__0_,
         npu_inst_pe_1_3_5_int_q_reg_h_5__1_,
         npu_inst_pe_1_3_5_int_q_reg_h_4__0_,
         npu_inst_pe_1_3_5_int_q_reg_h_4__1_,
         npu_inst_pe_1_3_5_int_q_reg_h_3__0_,
         npu_inst_pe_1_3_5_int_q_reg_h_3__1_,
         npu_inst_pe_1_3_5_int_q_reg_h_2__0_,
         npu_inst_pe_1_3_5_int_q_reg_h_2__1_,
         npu_inst_pe_1_3_5_int_q_reg_h_1__0_,
         npu_inst_pe_1_3_5_int_q_reg_h_1__1_,
         npu_inst_pe_1_3_5_int_q_reg_h_0__0_,
         npu_inst_pe_1_3_5_int_q_reg_h_0__1_, npu_inst_pe_1_3_6_n119,
         npu_inst_pe_1_3_6_n118, npu_inst_pe_1_3_6_n117,
         npu_inst_pe_1_3_6_n116, npu_inst_pe_1_3_6_n115,
         npu_inst_pe_1_3_6_n114, npu_inst_pe_1_3_6_n113,
         npu_inst_pe_1_3_6_n112, npu_inst_pe_1_3_6_n111,
         npu_inst_pe_1_3_6_n110, npu_inst_pe_1_3_6_n109,
         npu_inst_pe_1_3_6_n108, npu_inst_pe_1_3_6_n107,
         npu_inst_pe_1_3_6_n106, npu_inst_pe_1_3_6_n105,
         npu_inst_pe_1_3_6_n104, npu_inst_pe_1_3_6_n103,
         npu_inst_pe_1_3_6_n102, npu_inst_pe_1_3_6_n101,
         npu_inst_pe_1_3_6_n100, npu_inst_pe_1_3_6_n99, npu_inst_pe_1_3_6_n98,
         npu_inst_pe_1_3_6_n36, npu_inst_pe_1_3_6_n35, npu_inst_pe_1_3_6_n34,
         npu_inst_pe_1_3_6_n33, npu_inst_pe_1_3_6_n32, npu_inst_pe_1_3_6_n31,
         npu_inst_pe_1_3_6_n30, npu_inst_pe_1_3_6_n29, npu_inst_pe_1_3_6_n28,
         npu_inst_pe_1_3_6_n25, npu_inst_pe_1_3_6_n24, npu_inst_pe_1_3_6_n23,
         npu_inst_pe_1_3_6_n22, npu_inst_pe_1_3_6_n21, npu_inst_pe_1_3_6_n20,
         npu_inst_pe_1_3_6_n19, npu_inst_pe_1_3_6_n18, npu_inst_pe_1_3_6_n17,
         npu_inst_pe_1_3_6_n16, npu_inst_pe_1_3_6_n15, npu_inst_pe_1_3_6_n14,
         npu_inst_pe_1_3_6_n13, npu_inst_pe_1_3_6_n12, npu_inst_pe_1_3_6_n11,
         npu_inst_pe_1_3_6_n10, npu_inst_pe_1_3_6_n9, npu_inst_pe_1_3_6_n8,
         npu_inst_pe_1_3_6_n7, npu_inst_pe_1_3_6_n6, npu_inst_pe_1_3_6_n5,
         npu_inst_pe_1_3_6_n4, npu_inst_pe_1_3_6_n3, npu_inst_pe_1_3_6_n2,
         npu_inst_pe_1_3_6_n1, npu_inst_pe_1_3_6_sub_77_carry_7_,
         npu_inst_pe_1_3_6_sub_77_carry_6_, npu_inst_pe_1_3_6_sub_77_carry_5_,
         npu_inst_pe_1_3_6_sub_77_carry_4_, npu_inst_pe_1_3_6_sub_77_carry_3_,
         npu_inst_pe_1_3_6_sub_77_carry_2_, npu_inst_pe_1_3_6_sub_77_carry_1_,
         npu_inst_pe_1_3_6_add_79_carry_7_, npu_inst_pe_1_3_6_add_79_carry_6_,
         npu_inst_pe_1_3_6_add_79_carry_5_, npu_inst_pe_1_3_6_add_79_carry_4_,
         npu_inst_pe_1_3_6_add_79_carry_3_, npu_inst_pe_1_3_6_add_79_carry_2_,
         npu_inst_pe_1_3_6_add_79_carry_1_, npu_inst_pe_1_3_6_n97,
         npu_inst_pe_1_3_6_n96, npu_inst_pe_1_3_6_n95, npu_inst_pe_1_3_6_n94,
         npu_inst_pe_1_3_6_n93, npu_inst_pe_1_3_6_n92, npu_inst_pe_1_3_6_n91,
         npu_inst_pe_1_3_6_n90, npu_inst_pe_1_3_6_n89, npu_inst_pe_1_3_6_n88,
         npu_inst_pe_1_3_6_n87, npu_inst_pe_1_3_6_n86, npu_inst_pe_1_3_6_n85,
         npu_inst_pe_1_3_6_n84, npu_inst_pe_1_3_6_n83, npu_inst_pe_1_3_6_n82,
         npu_inst_pe_1_3_6_n81, npu_inst_pe_1_3_6_n80, npu_inst_pe_1_3_6_n79,
         npu_inst_pe_1_3_6_n78, npu_inst_pe_1_3_6_n77, npu_inst_pe_1_3_6_n76,
         npu_inst_pe_1_3_6_n75, npu_inst_pe_1_3_6_n74, npu_inst_pe_1_3_6_n73,
         npu_inst_pe_1_3_6_n72, npu_inst_pe_1_3_6_n71, npu_inst_pe_1_3_6_n70,
         npu_inst_pe_1_3_6_n69, npu_inst_pe_1_3_6_n68, npu_inst_pe_1_3_6_n67,
         npu_inst_pe_1_3_6_n66, npu_inst_pe_1_3_6_n65, npu_inst_pe_1_3_6_n64,
         npu_inst_pe_1_3_6_n63, npu_inst_pe_1_3_6_n62, npu_inst_pe_1_3_6_n61,
         npu_inst_pe_1_3_6_n60, npu_inst_pe_1_3_6_n59, npu_inst_pe_1_3_6_n58,
         npu_inst_pe_1_3_6_n57, npu_inst_pe_1_3_6_n56, npu_inst_pe_1_3_6_n55,
         npu_inst_pe_1_3_6_n54, npu_inst_pe_1_3_6_n53, npu_inst_pe_1_3_6_n52,
         npu_inst_pe_1_3_6_n51, npu_inst_pe_1_3_6_n50, npu_inst_pe_1_3_6_n49,
         npu_inst_pe_1_3_6_n48, npu_inst_pe_1_3_6_n47, npu_inst_pe_1_3_6_n46,
         npu_inst_pe_1_3_6_n45, npu_inst_pe_1_3_6_n44, npu_inst_pe_1_3_6_n43,
         npu_inst_pe_1_3_6_n42, npu_inst_pe_1_3_6_n41, npu_inst_pe_1_3_6_n40,
         npu_inst_pe_1_3_6_n39, npu_inst_pe_1_3_6_n38, npu_inst_pe_1_3_6_n37,
         npu_inst_pe_1_3_6_n27, npu_inst_pe_1_3_6_n26,
         npu_inst_pe_1_3_6_net3609, npu_inst_pe_1_3_6_net3603,
         npu_inst_pe_1_3_6_N94, npu_inst_pe_1_3_6_N93, npu_inst_pe_1_3_6_N84,
         npu_inst_pe_1_3_6_N80, npu_inst_pe_1_3_6_N79, npu_inst_pe_1_3_6_N78,
         npu_inst_pe_1_3_6_N77, npu_inst_pe_1_3_6_N76, npu_inst_pe_1_3_6_N75,
         npu_inst_pe_1_3_6_N74, npu_inst_pe_1_3_6_N73, npu_inst_pe_1_3_6_N72,
         npu_inst_pe_1_3_6_N71, npu_inst_pe_1_3_6_N70, npu_inst_pe_1_3_6_N69,
         npu_inst_pe_1_3_6_N68, npu_inst_pe_1_3_6_N67, npu_inst_pe_1_3_6_N66,
         npu_inst_pe_1_3_6_N65, npu_inst_pe_1_3_6_int_q_acc_0_,
         npu_inst_pe_1_3_6_int_q_acc_1_, npu_inst_pe_1_3_6_int_q_acc_2_,
         npu_inst_pe_1_3_6_int_q_acc_3_, npu_inst_pe_1_3_6_int_q_acc_4_,
         npu_inst_pe_1_3_6_int_q_acc_5_, npu_inst_pe_1_3_6_int_q_acc_6_,
         npu_inst_pe_1_3_6_int_q_acc_7_, npu_inst_pe_1_3_6_int_data_0_,
         npu_inst_pe_1_3_6_int_data_1_, npu_inst_pe_1_3_6_int_q_weight_0_,
         npu_inst_pe_1_3_6_int_q_weight_1_,
         npu_inst_pe_1_3_6_int_q_reg_v_5__0_,
         npu_inst_pe_1_3_6_int_q_reg_v_5__1_,
         npu_inst_pe_1_3_6_int_q_reg_v_4__0_,
         npu_inst_pe_1_3_6_int_q_reg_v_4__1_,
         npu_inst_pe_1_3_6_int_q_reg_v_3__0_,
         npu_inst_pe_1_3_6_int_q_reg_v_3__1_,
         npu_inst_pe_1_3_6_int_q_reg_v_2__0_,
         npu_inst_pe_1_3_6_int_q_reg_v_2__1_,
         npu_inst_pe_1_3_6_int_q_reg_v_1__0_,
         npu_inst_pe_1_3_6_int_q_reg_v_1__1_,
         npu_inst_pe_1_3_6_int_q_reg_v_0__0_,
         npu_inst_pe_1_3_6_int_q_reg_v_0__1_,
         npu_inst_pe_1_3_6_int_q_reg_h_5__0_,
         npu_inst_pe_1_3_6_int_q_reg_h_5__1_,
         npu_inst_pe_1_3_6_int_q_reg_h_4__0_,
         npu_inst_pe_1_3_6_int_q_reg_h_4__1_,
         npu_inst_pe_1_3_6_int_q_reg_h_3__0_,
         npu_inst_pe_1_3_6_int_q_reg_h_3__1_,
         npu_inst_pe_1_3_6_int_q_reg_h_2__0_,
         npu_inst_pe_1_3_6_int_q_reg_h_2__1_,
         npu_inst_pe_1_3_6_int_q_reg_h_1__0_,
         npu_inst_pe_1_3_6_int_q_reg_h_1__1_,
         npu_inst_pe_1_3_6_int_q_reg_h_0__0_,
         npu_inst_pe_1_3_6_int_q_reg_h_0__1_, npu_inst_pe_1_3_7_n119,
         npu_inst_pe_1_3_7_n118, npu_inst_pe_1_3_7_n117,
         npu_inst_pe_1_3_7_n116, npu_inst_pe_1_3_7_n115,
         npu_inst_pe_1_3_7_n114, npu_inst_pe_1_3_7_n113,
         npu_inst_pe_1_3_7_n112, npu_inst_pe_1_3_7_n111,
         npu_inst_pe_1_3_7_n110, npu_inst_pe_1_3_7_n109,
         npu_inst_pe_1_3_7_n108, npu_inst_pe_1_3_7_n107,
         npu_inst_pe_1_3_7_n106, npu_inst_pe_1_3_7_n105,
         npu_inst_pe_1_3_7_n104, npu_inst_pe_1_3_7_n103,
         npu_inst_pe_1_3_7_n102, npu_inst_pe_1_3_7_n101,
         npu_inst_pe_1_3_7_n100, npu_inst_pe_1_3_7_n99, npu_inst_pe_1_3_7_n98,
         npu_inst_pe_1_3_7_n36, npu_inst_pe_1_3_7_n35, npu_inst_pe_1_3_7_n34,
         npu_inst_pe_1_3_7_n33, npu_inst_pe_1_3_7_n32, npu_inst_pe_1_3_7_n31,
         npu_inst_pe_1_3_7_n30, npu_inst_pe_1_3_7_n29, npu_inst_pe_1_3_7_n28,
         npu_inst_pe_1_3_7_n25, npu_inst_pe_1_3_7_n24, npu_inst_pe_1_3_7_n23,
         npu_inst_pe_1_3_7_n22, npu_inst_pe_1_3_7_n21, npu_inst_pe_1_3_7_n20,
         npu_inst_pe_1_3_7_n19, npu_inst_pe_1_3_7_n18, npu_inst_pe_1_3_7_n17,
         npu_inst_pe_1_3_7_n16, npu_inst_pe_1_3_7_n15, npu_inst_pe_1_3_7_n14,
         npu_inst_pe_1_3_7_n13, npu_inst_pe_1_3_7_n12, npu_inst_pe_1_3_7_n11,
         npu_inst_pe_1_3_7_n10, npu_inst_pe_1_3_7_n9, npu_inst_pe_1_3_7_n8,
         npu_inst_pe_1_3_7_n7, npu_inst_pe_1_3_7_n6, npu_inst_pe_1_3_7_n5,
         npu_inst_pe_1_3_7_n4, npu_inst_pe_1_3_7_n3, npu_inst_pe_1_3_7_n2,
         npu_inst_pe_1_3_7_n1, npu_inst_pe_1_3_7_sub_77_carry_7_,
         npu_inst_pe_1_3_7_sub_77_carry_6_, npu_inst_pe_1_3_7_sub_77_carry_5_,
         npu_inst_pe_1_3_7_sub_77_carry_4_, npu_inst_pe_1_3_7_sub_77_carry_3_,
         npu_inst_pe_1_3_7_sub_77_carry_2_, npu_inst_pe_1_3_7_sub_77_carry_1_,
         npu_inst_pe_1_3_7_add_79_carry_7_, npu_inst_pe_1_3_7_add_79_carry_6_,
         npu_inst_pe_1_3_7_add_79_carry_5_, npu_inst_pe_1_3_7_add_79_carry_4_,
         npu_inst_pe_1_3_7_add_79_carry_3_, npu_inst_pe_1_3_7_add_79_carry_2_,
         npu_inst_pe_1_3_7_add_79_carry_1_, npu_inst_pe_1_3_7_n97,
         npu_inst_pe_1_3_7_n96, npu_inst_pe_1_3_7_n95, npu_inst_pe_1_3_7_n94,
         npu_inst_pe_1_3_7_n93, npu_inst_pe_1_3_7_n92, npu_inst_pe_1_3_7_n91,
         npu_inst_pe_1_3_7_n90, npu_inst_pe_1_3_7_n89, npu_inst_pe_1_3_7_n88,
         npu_inst_pe_1_3_7_n87, npu_inst_pe_1_3_7_n86, npu_inst_pe_1_3_7_n85,
         npu_inst_pe_1_3_7_n84, npu_inst_pe_1_3_7_n83, npu_inst_pe_1_3_7_n82,
         npu_inst_pe_1_3_7_n81, npu_inst_pe_1_3_7_n80, npu_inst_pe_1_3_7_n79,
         npu_inst_pe_1_3_7_n78, npu_inst_pe_1_3_7_n77, npu_inst_pe_1_3_7_n76,
         npu_inst_pe_1_3_7_n75, npu_inst_pe_1_3_7_n74, npu_inst_pe_1_3_7_n73,
         npu_inst_pe_1_3_7_n72, npu_inst_pe_1_3_7_n71, npu_inst_pe_1_3_7_n70,
         npu_inst_pe_1_3_7_n69, npu_inst_pe_1_3_7_n68, npu_inst_pe_1_3_7_n67,
         npu_inst_pe_1_3_7_n66, npu_inst_pe_1_3_7_n65, npu_inst_pe_1_3_7_n64,
         npu_inst_pe_1_3_7_n63, npu_inst_pe_1_3_7_n62, npu_inst_pe_1_3_7_n61,
         npu_inst_pe_1_3_7_n60, npu_inst_pe_1_3_7_n59, npu_inst_pe_1_3_7_n58,
         npu_inst_pe_1_3_7_n57, npu_inst_pe_1_3_7_n56, npu_inst_pe_1_3_7_n55,
         npu_inst_pe_1_3_7_n54, npu_inst_pe_1_3_7_n53, npu_inst_pe_1_3_7_n52,
         npu_inst_pe_1_3_7_n51, npu_inst_pe_1_3_7_n50, npu_inst_pe_1_3_7_n49,
         npu_inst_pe_1_3_7_n48, npu_inst_pe_1_3_7_n47, npu_inst_pe_1_3_7_n46,
         npu_inst_pe_1_3_7_n45, npu_inst_pe_1_3_7_n44, npu_inst_pe_1_3_7_n43,
         npu_inst_pe_1_3_7_n42, npu_inst_pe_1_3_7_n41, npu_inst_pe_1_3_7_n40,
         npu_inst_pe_1_3_7_n39, npu_inst_pe_1_3_7_n38, npu_inst_pe_1_3_7_n37,
         npu_inst_pe_1_3_7_n27, npu_inst_pe_1_3_7_n26,
         npu_inst_pe_1_3_7_net3586, npu_inst_pe_1_3_7_net3580,
         npu_inst_pe_1_3_7_N94, npu_inst_pe_1_3_7_N93, npu_inst_pe_1_3_7_N84,
         npu_inst_pe_1_3_7_N80, npu_inst_pe_1_3_7_N79, npu_inst_pe_1_3_7_N78,
         npu_inst_pe_1_3_7_N77, npu_inst_pe_1_3_7_N76, npu_inst_pe_1_3_7_N75,
         npu_inst_pe_1_3_7_N74, npu_inst_pe_1_3_7_N73, npu_inst_pe_1_3_7_N72,
         npu_inst_pe_1_3_7_N71, npu_inst_pe_1_3_7_N70, npu_inst_pe_1_3_7_N69,
         npu_inst_pe_1_3_7_N68, npu_inst_pe_1_3_7_N67, npu_inst_pe_1_3_7_N66,
         npu_inst_pe_1_3_7_N65, npu_inst_pe_1_3_7_int_q_acc_0_,
         npu_inst_pe_1_3_7_int_q_acc_1_, npu_inst_pe_1_3_7_int_q_acc_2_,
         npu_inst_pe_1_3_7_int_q_acc_3_, npu_inst_pe_1_3_7_int_q_acc_4_,
         npu_inst_pe_1_3_7_int_q_acc_5_, npu_inst_pe_1_3_7_int_q_acc_6_,
         npu_inst_pe_1_3_7_int_q_acc_7_, npu_inst_pe_1_3_7_int_data_0_,
         npu_inst_pe_1_3_7_int_data_1_, npu_inst_pe_1_3_7_int_q_weight_0_,
         npu_inst_pe_1_3_7_int_q_weight_1_,
         npu_inst_pe_1_3_7_int_q_reg_v_5__0_,
         npu_inst_pe_1_3_7_int_q_reg_v_5__1_,
         npu_inst_pe_1_3_7_int_q_reg_v_4__0_,
         npu_inst_pe_1_3_7_int_q_reg_v_4__1_,
         npu_inst_pe_1_3_7_int_q_reg_v_3__0_,
         npu_inst_pe_1_3_7_int_q_reg_v_3__1_,
         npu_inst_pe_1_3_7_int_q_reg_v_2__0_,
         npu_inst_pe_1_3_7_int_q_reg_v_2__1_,
         npu_inst_pe_1_3_7_int_q_reg_v_1__0_,
         npu_inst_pe_1_3_7_int_q_reg_v_1__1_,
         npu_inst_pe_1_3_7_int_q_reg_v_0__0_,
         npu_inst_pe_1_3_7_int_q_reg_v_0__1_,
         npu_inst_pe_1_3_7_int_q_reg_h_5__0_,
         npu_inst_pe_1_3_7_int_q_reg_h_5__1_,
         npu_inst_pe_1_3_7_int_q_reg_h_4__0_,
         npu_inst_pe_1_3_7_int_q_reg_h_4__1_,
         npu_inst_pe_1_3_7_int_q_reg_h_3__0_,
         npu_inst_pe_1_3_7_int_q_reg_h_3__1_,
         npu_inst_pe_1_3_7_int_q_reg_h_2__0_,
         npu_inst_pe_1_3_7_int_q_reg_h_2__1_,
         npu_inst_pe_1_3_7_int_q_reg_h_1__0_,
         npu_inst_pe_1_3_7_int_q_reg_h_1__1_,
         npu_inst_pe_1_3_7_int_q_reg_h_0__0_,
         npu_inst_pe_1_3_7_int_q_reg_h_0__1_, npu_inst_pe_1_4_0_n119,
         npu_inst_pe_1_4_0_n118, npu_inst_pe_1_4_0_n117,
         npu_inst_pe_1_4_0_n116, npu_inst_pe_1_4_0_n115,
         npu_inst_pe_1_4_0_n114, npu_inst_pe_1_4_0_n113,
         npu_inst_pe_1_4_0_n112, npu_inst_pe_1_4_0_n111,
         npu_inst_pe_1_4_0_n110, npu_inst_pe_1_4_0_n109,
         npu_inst_pe_1_4_0_n108, npu_inst_pe_1_4_0_n107,
         npu_inst_pe_1_4_0_n106, npu_inst_pe_1_4_0_n105,
         npu_inst_pe_1_4_0_n104, npu_inst_pe_1_4_0_n103,
         npu_inst_pe_1_4_0_n102, npu_inst_pe_1_4_0_n101,
         npu_inst_pe_1_4_0_n100, npu_inst_pe_1_4_0_n99, npu_inst_pe_1_4_0_n98,
         npu_inst_pe_1_4_0_n36, npu_inst_pe_1_4_0_n35, npu_inst_pe_1_4_0_n34,
         npu_inst_pe_1_4_0_n33, npu_inst_pe_1_4_0_n32, npu_inst_pe_1_4_0_n31,
         npu_inst_pe_1_4_0_n30, npu_inst_pe_1_4_0_n29, npu_inst_pe_1_4_0_n28,
         npu_inst_pe_1_4_0_n25, npu_inst_pe_1_4_0_n24, npu_inst_pe_1_4_0_n23,
         npu_inst_pe_1_4_0_n22, npu_inst_pe_1_4_0_n21, npu_inst_pe_1_4_0_n20,
         npu_inst_pe_1_4_0_n19, npu_inst_pe_1_4_0_n18, npu_inst_pe_1_4_0_n17,
         npu_inst_pe_1_4_0_n16, npu_inst_pe_1_4_0_n15, npu_inst_pe_1_4_0_n14,
         npu_inst_pe_1_4_0_n13, npu_inst_pe_1_4_0_n12, npu_inst_pe_1_4_0_n11,
         npu_inst_pe_1_4_0_n10, npu_inst_pe_1_4_0_n9, npu_inst_pe_1_4_0_n8,
         npu_inst_pe_1_4_0_n7, npu_inst_pe_1_4_0_n6, npu_inst_pe_1_4_0_n5,
         npu_inst_pe_1_4_0_n4, npu_inst_pe_1_4_0_n3, npu_inst_pe_1_4_0_n2,
         npu_inst_pe_1_4_0_n1, npu_inst_pe_1_4_0_sub_77_carry_7_,
         npu_inst_pe_1_4_0_sub_77_carry_6_, npu_inst_pe_1_4_0_sub_77_carry_5_,
         npu_inst_pe_1_4_0_sub_77_carry_4_, npu_inst_pe_1_4_0_sub_77_carry_3_,
         npu_inst_pe_1_4_0_sub_77_carry_2_, npu_inst_pe_1_4_0_sub_77_carry_1_,
         npu_inst_pe_1_4_0_add_79_carry_7_, npu_inst_pe_1_4_0_add_79_carry_6_,
         npu_inst_pe_1_4_0_add_79_carry_5_, npu_inst_pe_1_4_0_add_79_carry_4_,
         npu_inst_pe_1_4_0_add_79_carry_3_, npu_inst_pe_1_4_0_add_79_carry_2_,
         npu_inst_pe_1_4_0_add_79_carry_1_, npu_inst_pe_1_4_0_n97,
         npu_inst_pe_1_4_0_n96, npu_inst_pe_1_4_0_n95, npu_inst_pe_1_4_0_n94,
         npu_inst_pe_1_4_0_n93, npu_inst_pe_1_4_0_n92, npu_inst_pe_1_4_0_n91,
         npu_inst_pe_1_4_0_n90, npu_inst_pe_1_4_0_n89, npu_inst_pe_1_4_0_n88,
         npu_inst_pe_1_4_0_n87, npu_inst_pe_1_4_0_n86, npu_inst_pe_1_4_0_n85,
         npu_inst_pe_1_4_0_n84, npu_inst_pe_1_4_0_n83, npu_inst_pe_1_4_0_n82,
         npu_inst_pe_1_4_0_n81, npu_inst_pe_1_4_0_n80, npu_inst_pe_1_4_0_n79,
         npu_inst_pe_1_4_0_n78, npu_inst_pe_1_4_0_n77, npu_inst_pe_1_4_0_n76,
         npu_inst_pe_1_4_0_n75, npu_inst_pe_1_4_0_n74, npu_inst_pe_1_4_0_n73,
         npu_inst_pe_1_4_0_n72, npu_inst_pe_1_4_0_n71, npu_inst_pe_1_4_0_n70,
         npu_inst_pe_1_4_0_n69, npu_inst_pe_1_4_0_n68, npu_inst_pe_1_4_0_n67,
         npu_inst_pe_1_4_0_n66, npu_inst_pe_1_4_0_n65, npu_inst_pe_1_4_0_n64,
         npu_inst_pe_1_4_0_n63, npu_inst_pe_1_4_0_n62, npu_inst_pe_1_4_0_n61,
         npu_inst_pe_1_4_0_n60, npu_inst_pe_1_4_0_n59, npu_inst_pe_1_4_0_n58,
         npu_inst_pe_1_4_0_n57, npu_inst_pe_1_4_0_n56, npu_inst_pe_1_4_0_n55,
         npu_inst_pe_1_4_0_n54, npu_inst_pe_1_4_0_n53, npu_inst_pe_1_4_0_n52,
         npu_inst_pe_1_4_0_n51, npu_inst_pe_1_4_0_n50, npu_inst_pe_1_4_0_n49,
         npu_inst_pe_1_4_0_n48, npu_inst_pe_1_4_0_n47, npu_inst_pe_1_4_0_n46,
         npu_inst_pe_1_4_0_n45, npu_inst_pe_1_4_0_n44, npu_inst_pe_1_4_0_n43,
         npu_inst_pe_1_4_0_n42, npu_inst_pe_1_4_0_n41, npu_inst_pe_1_4_0_n40,
         npu_inst_pe_1_4_0_n39, npu_inst_pe_1_4_0_n38, npu_inst_pe_1_4_0_n37,
         npu_inst_pe_1_4_0_n27, npu_inst_pe_1_4_0_n26,
         npu_inst_pe_1_4_0_net3563, npu_inst_pe_1_4_0_net3557,
         npu_inst_pe_1_4_0_N94, npu_inst_pe_1_4_0_N93, npu_inst_pe_1_4_0_N84,
         npu_inst_pe_1_4_0_N80, npu_inst_pe_1_4_0_N79, npu_inst_pe_1_4_0_N78,
         npu_inst_pe_1_4_0_N77, npu_inst_pe_1_4_0_N76, npu_inst_pe_1_4_0_N75,
         npu_inst_pe_1_4_0_N74, npu_inst_pe_1_4_0_N73, npu_inst_pe_1_4_0_N72,
         npu_inst_pe_1_4_0_N71, npu_inst_pe_1_4_0_N70, npu_inst_pe_1_4_0_N69,
         npu_inst_pe_1_4_0_N68, npu_inst_pe_1_4_0_N67, npu_inst_pe_1_4_0_N66,
         npu_inst_pe_1_4_0_N65, npu_inst_pe_1_4_0_int_q_acc_0_,
         npu_inst_pe_1_4_0_int_q_acc_1_, npu_inst_pe_1_4_0_int_q_acc_2_,
         npu_inst_pe_1_4_0_int_q_acc_3_, npu_inst_pe_1_4_0_int_q_acc_4_,
         npu_inst_pe_1_4_0_int_q_acc_5_, npu_inst_pe_1_4_0_int_q_acc_6_,
         npu_inst_pe_1_4_0_int_q_acc_7_, npu_inst_pe_1_4_0_int_data_0_,
         npu_inst_pe_1_4_0_int_data_1_, npu_inst_pe_1_4_0_int_q_weight_0_,
         npu_inst_pe_1_4_0_int_q_weight_1_,
         npu_inst_pe_1_4_0_int_q_reg_v_5__0_,
         npu_inst_pe_1_4_0_int_q_reg_v_5__1_,
         npu_inst_pe_1_4_0_int_q_reg_v_4__0_,
         npu_inst_pe_1_4_0_int_q_reg_v_4__1_,
         npu_inst_pe_1_4_0_int_q_reg_v_3__0_,
         npu_inst_pe_1_4_0_int_q_reg_v_3__1_,
         npu_inst_pe_1_4_0_int_q_reg_v_2__0_,
         npu_inst_pe_1_4_0_int_q_reg_v_2__1_,
         npu_inst_pe_1_4_0_int_q_reg_v_1__0_,
         npu_inst_pe_1_4_0_int_q_reg_v_1__1_,
         npu_inst_pe_1_4_0_int_q_reg_v_0__0_,
         npu_inst_pe_1_4_0_int_q_reg_v_0__1_,
         npu_inst_pe_1_4_0_int_q_reg_h_5__0_,
         npu_inst_pe_1_4_0_int_q_reg_h_5__1_,
         npu_inst_pe_1_4_0_int_q_reg_h_4__0_,
         npu_inst_pe_1_4_0_int_q_reg_h_4__1_,
         npu_inst_pe_1_4_0_int_q_reg_h_3__0_,
         npu_inst_pe_1_4_0_int_q_reg_h_3__1_,
         npu_inst_pe_1_4_0_int_q_reg_h_2__0_,
         npu_inst_pe_1_4_0_int_q_reg_h_2__1_,
         npu_inst_pe_1_4_0_int_q_reg_h_1__0_,
         npu_inst_pe_1_4_0_int_q_reg_h_1__1_,
         npu_inst_pe_1_4_0_int_q_reg_h_0__0_,
         npu_inst_pe_1_4_0_int_q_reg_h_0__1_, npu_inst_pe_1_4_0_o_data_h_0_,
         npu_inst_pe_1_4_0_o_data_h_1_, npu_inst_pe_1_4_1_n119,
         npu_inst_pe_1_4_1_n118, npu_inst_pe_1_4_1_n117,
         npu_inst_pe_1_4_1_n116, npu_inst_pe_1_4_1_n115,
         npu_inst_pe_1_4_1_n114, npu_inst_pe_1_4_1_n113,
         npu_inst_pe_1_4_1_n112, npu_inst_pe_1_4_1_n111,
         npu_inst_pe_1_4_1_n110, npu_inst_pe_1_4_1_n109,
         npu_inst_pe_1_4_1_n108, npu_inst_pe_1_4_1_n107,
         npu_inst_pe_1_4_1_n106, npu_inst_pe_1_4_1_n105,
         npu_inst_pe_1_4_1_n104, npu_inst_pe_1_4_1_n103,
         npu_inst_pe_1_4_1_n102, npu_inst_pe_1_4_1_n101,
         npu_inst_pe_1_4_1_n100, npu_inst_pe_1_4_1_n99, npu_inst_pe_1_4_1_n98,
         npu_inst_pe_1_4_1_n36, npu_inst_pe_1_4_1_n35, npu_inst_pe_1_4_1_n34,
         npu_inst_pe_1_4_1_n33, npu_inst_pe_1_4_1_n32, npu_inst_pe_1_4_1_n31,
         npu_inst_pe_1_4_1_n30, npu_inst_pe_1_4_1_n29, npu_inst_pe_1_4_1_n28,
         npu_inst_pe_1_4_1_n25, npu_inst_pe_1_4_1_n24, npu_inst_pe_1_4_1_n23,
         npu_inst_pe_1_4_1_n22, npu_inst_pe_1_4_1_n21, npu_inst_pe_1_4_1_n20,
         npu_inst_pe_1_4_1_n19, npu_inst_pe_1_4_1_n18, npu_inst_pe_1_4_1_n17,
         npu_inst_pe_1_4_1_n16, npu_inst_pe_1_4_1_n15, npu_inst_pe_1_4_1_n14,
         npu_inst_pe_1_4_1_n13, npu_inst_pe_1_4_1_n12, npu_inst_pe_1_4_1_n11,
         npu_inst_pe_1_4_1_n10, npu_inst_pe_1_4_1_n9, npu_inst_pe_1_4_1_n8,
         npu_inst_pe_1_4_1_n7, npu_inst_pe_1_4_1_n6, npu_inst_pe_1_4_1_n5,
         npu_inst_pe_1_4_1_n4, npu_inst_pe_1_4_1_n3, npu_inst_pe_1_4_1_n2,
         npu_inst_pe_1_4_1_n1, npu_inst_pe_1_4_1_sub_77_carry_7_,
         npu_inst_pe_1_4_1_sub_77_carry_6_, npu_inst_pe_1_4_1_sub_77_carry_5_,
         npu_inst_pe_1_4_1_sub_77_carry_4_, npu_inst_pe_1_4_1_sub_77_carry_3_,
         npu_inst_pe_1_4_1_sub_77_carry_2_, npu_inst_pe_1_4_1_sub_77_carry_1_,
         npu_inst_pe_1_4_1_add_79_carry_7_, npu_inst_pe_1_4_1_add_79_carry_6_,
         npu_inst_pe_1_4_1_add_79_carry_5_, npu_inst_pe_1_4_1_add_79_carry_4_,
         npu_inst_pe_1_4_1_add_79_carry_3_, npu_inst_pe_1_4_1_add_79_carry_2_,
         npu_inst_pe_1_4_1_add_79_carry_1_, npu_inst_pe_1_4_1_n97,
         npu_inst_pe_1_4_1_n96, npu_inst_pe_1_4_1_n95, npu_inst_pe_1_4_1_n94,
         npu_inst_pe_1_4_1_n93, npu_inst_pe_1_4_1_n92, npu_inst_pe_1_4_1_n91,
         npu_inst_pe_1_4_1_n90, npu_inst_pe_1_4_1_n89, npu_inst_pe_1_4_1_n88,
         npu_inst_pe_1_4_1_n87, npu_inst_pe_1_4_1_n86, npu_inst_pe_1_4_1_n85,
         npu_inst_pe_1_4_1_n84, npu_inst_pe_1_4_1_n83, npu_inst_pe_1_4_1_n82,
         npu_inst_pe_1_4_1_n81, npu_inst_pe_1_4_1_n80, npu_inst_pe_1_4_1_n79,
         npu_inst_pe_1_4_1_n78, npu_inst_pe_1_4_1_n77, npu_inst_pe_1_4_1_n76,
         npu_inst_pe_1_4_1_n75, npu_inst_pe_1_4_1_n74, npu_inst_pe_1_4_1_n73,
         npu_inst_pe_1_4_1_n72, npu_inst_pe_1_4_1_n71, npu_inst_pe_1_4_1_n70,
         npu_inst_pe_1_4_1_n69, npu_inst_pe_1_4_1_n68, npu_inst_pe_1_4_1_n67,
         npu_inst_pe_1_4_1_n66, npu_inst_pe_1_4_1_n65, npu_inst_pe_1_4_1_n64,
         npu_inst_pe_1_4_1_n63, npu_inst_pe_1_4_1_n62, npu_inst_pe_1_4_1_n61,
         npu_inst_pe_1_4_1_n60, npu_inst_pe_1_4_1_n59, npu_inst_pe_1_4_1_n58,
         npu_inst_pe_1_4_1_n57, npu_inst_pe_1_4_1_n56, npu_inst_pe_1_4_1_n55,
         npu_inst_pe_1_4_1_n54, npu_inst_pe_1_4_1_n53, npu_inst_pe_1_4_1_n52,
         npu_inst_pe_1_4_1_n51, npu_inst_pe_1_4_1_n50, npu_inst_pe_1_4_1_n49,
         npu_inst_pe_1_4_1_n48, npu_inst_pe_1_4_1_n47, npu_inst_pe_1_4_1_n46,
         npu_inst_pe_1_4_1_n45, npu_inst_pe_1_4_1_n44, npu_inst_pe_1_4_1_n43,
         npu_inst_pe_1_4_1_n42, npu_inst_pe_1_4_1_n41, npu_inst_pe_1_4_1_n40,
         npu_inst_pe_1_4_1_n39, npu_inst_pe_1_4_1_n38, npu_inst_pe_1_4_1_n37,
         npu_inst_pe_1_4_1_n27, npu_inst_pe_1_4_1_n26,
         npu_inst_pe_1_4_1_net3540, npu_inst_pe_1_4_1_net3534,
         npu_inst_pe_1_4_1_N94, npu_inst_pe_1_4_1_N93, npu_inst_pe_1_4_1_N84,
         npu_inst_pe_1_4_1_N80, npu_inst_pe_1_4_1_N79, npu_inst_pe_1_4_1_N78,
         npu_inst_pe_1_4_1_N77, npu_inst_pe_1_4_1_N76, npu_inst_pe_1_4_1_N75,
         npu_inst_pe_1_4_1_N74, npu_inst_pe_1_4_1_N73, npu_inst_pe_1_4_1_N72,
         npu_inst_pe_1_4_1_N71, npu_inst_pe_1_4_1_N70, npu_inst_pe_1_4_1_N69,
         npu_inst_pe_1_4_1_N68, npu_inst_pe_1_4_1_N67, npu_inst_pe_1_4_1_N66,
         npu_inst_pe_1_4_1_N65, npu_inst_pe_1_4_1_int_q_acc_0_,
         npu_inst_pe_1_4_1_int_q_acc_1_, npu_inst_pe_1_4_1_int_q_acc_2_,
         npu_inst_pe_1_4_1_int_q_acc_3_, npu_inst_pe_1_4_1_int_q_acc_4_,
         npu_inst_pe_1_4_1_int_q_acc_5_, npu_inst_pe_1_4_1_int_q_acc_6_,
         npu_inst_pe_1_4_1_int_q_acc_7_, npu_inst_pe_1_4_1_int_data_0_,
         npu_inst_pe_1_4_1_int_data_1_, npu_inst_pe_1_4_1_int_q_weight_0_,
         npu_inst_pe_1_4_1_int_q_weight_1_,
         npu_inst_pe_1_4_1_int_q_reg_v_5__0_,
         npu_inst_pe_1_4_1_int_q_reg_v_5__1_,
         npu_inst_pe_1_4_1_int_q_reg_v_4__0_,
         npu_inst_pe_1_4_1_int_q_reg_v_4__1_,
         npu_inst_pe_1_4_1_int_q_reg_v_3__0_,
         npu_inst_pe_1_4_1_int_q_reg_v_3__1_,
         npu_inst_pe_1_4_1_int_q_reg_v_2__0_,
         npu_inst_pe_1_4_1_int_q_reg_v_2__1_,
         npu_inst_pe_1_4_1_int_q_reg_v_1__0_,
         npu_inst_pe_1_4_1_int_q_reg_v_1__1_,
         npu_inst_pe_1_4_1_int_q_reg_v_0__0_,
         npu_inst_pe_1_4_1_int_q_reg_v_0__1_,
         npu_inst_pe_1_4_1_int_q_reg_h_5__0_,
         npu_inst_pe_1_4_1_int_q_reg_h_5__1_,
         npu_inst_pe_1_4_1_int_q_reg_h_4__0_,
         npu_inst_pe_1_4_1_int_q_reg_h_4__1_,
         npu_inst_pe_1_4_1_int_q_reg_h_3__0_,
         npu_inst_pe_1_4_1_int_q_reg_h_3__1_,
         npu_inst_pe_1_4_1_int_q_reg_h_2__0_,
         npu_inst_pe_1_4_1_int_q_reg_h_2__1_,
         npu_inst_pe_1_4_1_int_q_reg_h_1__0_,
         npu_inst_pe_1_4_1_int_q_reg_h_1__1_,
         npu_inst_pe_1_4_1_int_q_reg_h_0__0_,
         npu_inst_pe_1_4_1_int_q_reg_h_0__1_, npu_inst_pe_1_4_2_n119,
         npu_inst_pe_1_4_2_n118, npu_inst_pe_1_4_2_n117,
         npu_inst_pe_1_4_2_n116, npu_inst_pe_1_4_2_n115,
         npu_inst_pe_1_4_2_n114, npu_inst_pe_1_4_2_n113,
         npu_inst_pe_1_4_2_n112, npu_inst_pe_1_4_2_n111,
         npu_inst_pe_1_4_2_n110, npu_inst_pe_1_4_2_n109,
         npu_inst_pe_1_4_2_n108, npu_inst_pe_1_4_2_n107,
         npu_inst_pe_1_4_2_n106, npu_inst_pe_1_4_2_n105,
         npu_inst_pe_1_4_2_n104, npu_inst_pe_1_4_2_n103,
         npu_inst_pe_1_4_2_n102, npu_inst_pe_1_4_2_n101,
         npu_inst_pe_1_4_2_n100, npu_inst_pe_1_4_2_n99, npu_inst_pe_1_4_2_n98,
         npu_inst_pe_1_4_2_n36, npu_inst_pe_1_4_2_n35, npu_inst_pe_1_4_2_n34,
         npu_inst_pe_1_4_2_n33, npu_inst_pe_1_4_2_n32, npu_inst_pe_1_4_2_n31,
         npu_inst_pe_1_4_2_n30, npu_inst_pe_1_4_2_n29, npu_inst_pe_1_4_2_n28,
         npu_inst_pe_1_4_2_n25, npu_inst_pe_1_4_2_n24, npu_inst_pe_1_4_2_n23,
         npu_inst_pe_1_4_2_n22, npu_inst_pe_1_4_2_n21, npu_inst_pe_1_4_2_n20,
         npu_inst_pe_1_4_2_n19, npu_inst_pe_1_4_2_n18, npu_inst_pe_1_4_2_n17,
         npu_inst_pe_1_4_2_n16, npu_inst_pe_1_4_2_n15, npu_inst_pe_1_4_2_n14,
         npu_inst_pe_1_4_2_n13, npu_inst_pe_1_4_2_n12, npu_inst_pe_1_4_2_n11,
         npu_inst_pe_1_4_2_n10, npu_inst_pe_1_4_2_n9, npu_inst_pe_1_4_2_n8,
         npu_inst_pe_1_4_2_n7, npu_inst_pe_1_4_2_n6, npu_inst_pe_1_4_2_n5,
         npu_inst_pe_1_4_2_n4, npu_inst_pe_1_4_2_n3, npu_inst_pe_1_4_2_n2,
         npu_inst_pe_1_4_2_n1, npu_inst_pe_1_4_2_sub_77_carry_7_,
         npu_inst_pe_1_4_2_sub_77_carry_6_, npu_inst_pe_1_4_2_sub_77_carry_5_,
         npu_inst_pe_1_4_2_sub_77_carry_4_, npu_inst_pe_1_4_2_sub_77_carry_3_,
         npu_inst_pe_1_4_2_sub_77_carry_2_, npu_inst_pe_1_4_2_sub_77_carry_1_,
         npu_inst_pe_1_4_2_add_79_carry_7_, npu_inst_pe_1_4_2_add_79_carry_6_,
         npu_inst_pe_1_4_2_add_79_carry_5_, npu_inst_pe_1_4_2_add_79_carry_4_,
         npu_inst_pe_1_4_2_add_79_carry_3_, npu_inst_pe_1_4_2_add_79_carry_2_,
         npu_inst_pe_1_4_2_add_79_carry_1_, npu_inst_pe_1_4_2_n97,
         npu_inst_pe_1_4_2_n96, npu_inst_pe_1_4_2_n95, npu_inst_pe_1_4_2_n94,
         npu_inst_pe_1_4_2_n93, npu_inst_pe_1_4_2_n92, npu_inst_pe_1_4_2_n91,
         npu_inst_pe_1_4_2_n90, npu_inst_pe_1_4_2_n89, npu_inst_pe_1_4_2_n88,
         npu_inst_pe_1_4_2_n87, npu_inst_pe_1_4_2_n86, npu_inst_pe_1_4_2_n85,
         npu_inst_pe_1_4_2_n84, npu_inst_pe_1_4_2_n83, npu_inst_pe_1_4_2_n82,
         npu_inst_pe_1_4_2_n81, npu_inst_pe_1_4_2_n80, npu_inst_pe_1_4_2_n79,
         npu_inst_pe_1_4_2_n78, npu_inst_pe_1_4_2_n77, npu_inst_pe_1_4_2_n76,
         npu_inst_pe_1_4_2_n75, npu_inst_pe_1_4_2_n74, npu_inst_pe_1_4_2_n73,
         npu_inst_pe_1_4_2_n72, npu_inst_pe_1_4_2_n71, npu_inst_pe_1_4_2_n70,
         npu_inst_pe_1_4_2_n69, npu_inst_pe_1_4_2_n68, npu_inst_pe_1_4_2_n67,
         npu_inst_pe_1_4_2_n66, npu_inst_pe_1_4_2_n65, npu_inst_pe_1_4_2_n64,
         npu_inst_pe_1_4_2_n63, npu_inst_pe_1_4_2_n62, npu_inst_pe_1_4_2_n61,
         npu_inst_pe_1_4_2_n60, npu_inst_pe_1_4_2_n59, npu_inst_pe_1_4_2_n58,
         npu_inst_pe_1_4_2_n57, npu_inst_pe_1_4_2_n56, npu_inst_pe_1_4_2_n55,
         npu_inst_pe_1_4_2_n54, npu_inst_pe_1_4_2_n53, npu_inst_pe_1_4_2_n52,
         npu_inst_pe_1_4_2_n51, npu_inst_pe_1_4_2_n50, npu_inst_pe_1_4_2_n49,
         npu_inst_pe_1_4_2_n48, npu_inst_pe_1_4_2_n47, npu_inst_pe_1_4_2_n46,
         npu_inst_pe_1_4_2_n45, npu_inst_pe_1_4_2_n44, npu_inst_pe_1_4_2_n43,
         npu_inst_pe_1_4_2_n42, npu_inst_pe_1_4_2_n41, npu_inst_pe_1_4_2_n40,
         npu_inst_pe_1_4_2_n39, npu_inst_pe_1_4_2_n38, npu_inst_pe_1_4_2_n37,
         npu_inst_pe_1_4_2_n27, npu_inst_pe_1_4_2_n26,
         npu_inst_pe_1_4_2_net3517, npu_inst_pe_1_4_2_net3511,
         npu_inst_pe_1_4_2_N94, npu_inst_pe_1_4_2_N93, npu_inst_pe_1_4_2_N84,
         npu_inst_pe_1_4_2_N80, npu_inst_pe_1_4_2_N79, npu_inst_pe_1_4_2_N78,
         npu_inst_pe_1_4_2_N77, npu_inst_pe_1_4_2_N76, npu_inst_pe_1_4_2_N75,
         npu_inst_pe_1_4_2_N74, npu_inst_pe_1_4_2_N73, npu_inst_pe_1_4_2_N72,
         npu_inst_pe_1_4_2_N71, npu_inst_pe_1_4_2_N70, npu_inst_pe_1_4_2_N69,
         npu_inst_pe_1_4_2_N68, npu_inst_pe_1_4_2_N67, npu_inst_pe_1_4_2_N66,
         npu_inst_pe_1_4_2_N65, npu_inst_pe_1_4_2_int_q_acc_0_,
         npu_inst_pe_1_4_2_int_q_acc_1_, npu_inst_pe_1_4_2_int_q_acc_2_,
         npu_inst_pe_1_4_2_int_q_acc_3_, npu_inst_pe_1_4_2_int_q_acc_4_,
         npu_inst_pe_1_4_2_int_q_acc_5_, npu_inst_pe_1_4_2_int_q_acc_6_,
         npu_inst_pe_1_4_2_int_q_acc_7_, npu_inst_pe_1_4_2_int_data_0_,
         npu_inst_pe_1_4_2_int_data_1_, npu_inst_pe_1_4_2_int_q_weight_0_,
         npu_inst_pe_1_4_2_int_q_weight_1_,
         npu_inst_pe_1_4_2_int_q_reg_v_5__0_,
         npu_inst_pe_1_4_2_int_q_reg_v_5__1_,
         npu_inst_pe_1_4_2_int_q_reg_v_4__0_,
         npu_inst_pe_1_4_2_int_q_reg_v_4__1_,
         npu_inst_pe_1_4_2_int_q_reg_v_3__0_,
         npu_inst_pe_1_4_2_int_q_reg_v_3__1_,
         npu_inst_pe_1_4_2_int_q_reg_v_2__0_,
         npu_inst_pe_1_4_2_int_q_reg_v_2__1_,
         npu_inst_pe_1_4_2_int_q_reg_v_1__0_,
         npu_inst_pe_1_4_2_int_q_reg_v_1__1_,
         npu_inst_pe_1_4_2_int_q_reg_v_0__0_,
         npu_inst_pe_1_4_2_int_q_reg_v_0__1_,
         npu_inst_pe_1_4_2_int_q_reg_h_5__0_,
         npu_inst_pe_1_4_2_int_q_reg_h_5__1_,
         npu_inst_pe_1_4_2_int_q_reg_h_4__0_,
         npu_inst_pe_1_4_2_int_q_reg_h_4__1_,
         npu_inst_pe_1_4_2_int_q_reg_h_3__0_,
         npu_inst_pe_1_4_2_int_q_reg_h_3__1_,
         npu_inst_pe_1_4_2_int_q_reg_h_2__0_,
         npu_inst_pe_1_4_2_int_q_reg_h_2__1_,
         npu_inst_pe_1_4_2_int_q_reg_h_1__0_,
         npu_inst_pe_1_4_2_int_q_reg_h_1__1_,
         npu_inst_pe_1_4_2_int_q_reg_h_0__0_,
         npu_inst_pe_1_4_2_int_q_reg_h_0__1_, npu_inst_pe_1_4_3_n119,
         npu_inst_pe_1_4_3_n118, npu_inst_pe_1_4_3_n117,
         npu_inst_pe_1_4_3_n116, npu_inst_pe_1_4_3_n115,
         npu_inst_pe_1_4_3_n114, npu_inst_pe_1_4_3_n113,
         npu_inst_pe_1_4_3_n112, npu_inst_pe_1_4_3_n111,
         npu_inst_pe_1_4_3_n110, npu_inst_pe_1_4_3_n109,
         npu_inst_pe_1_4_3_n108, npu_inst_pe_1_4_3_n107,
         npu_inst_pe_1_4_3_n106, npu_inst_pe_1_4_3_n105,
         npu_inst_pe_1_4_3_n104, npu_inst_pe_1_4_3_n103,
         npu_inst_pe_1_4_3_n102, npu_inst_pe_1_4_3_n101,
         npu_inst_pe_1_4_3_n100, npu_inst_pe_1_4_3_n99, npu_inst_pe_1_4_3_n98,
         npu_inst_pe_1_4_3_n36, npu_inst_pe_1_4_3_n35, npu_inst_pe_1_4_3_n34,
         npu_inst_pe_1_4_3_n33, npu_inst_pe_1_4_3_n32, npu_inst_pe_1_4_3_n31,
         npu_inst_pe_1_4_3_n30, npu_inst_pe_1_4_3_n29, npu_inst_pe_1_4_3_n28,
         npu_inst_pe_1_4_3_n25, npu_inst_pe_1_4_3_n24, npu_inst_pe_1_4_3_n23,
         npu_inst_pe_1_4_3_n22, npu_inst_pe_1_4_3_n21, npu_inst_pe_1_4_3_n20,
         npu_inst_pe_1_4_3_n19, npu_inst_pe_1_4_3_n18, npu_inst_pe_1_4_3_n17,
         npu_inst_pe_1_4_3_n16, npu_inst_pe_1_4_3_n15, npu_inst_pe_1_4_3_n14,
         npu_inst_pe_1_4_3_n13, npu_inst_pe_1_4_3_n12, npu_inst_pe_1_4_3_n11,
         npu_inst_pe_1_4_3_n10, npu_inst_pe_1_4_3_n9, npu_inst_pe_1_4_3_n8,
         npu_inst_pe_1_4_3_n7, npu_inst_pe_1_4_3_n6, npu_inst_pe_1_4_3_n5,
         npu_inst_pe_1_4_3_n4, npu_inst_pe_1_4_3_n3, npu_inst_pe_1_4_3_n2,
         npu_inst_pe_1_4_3_n1, npu_inst_pe_1_4_3_sub_77_carry_7_,
         npu_inst_pe_1_4_3_sub_77_carry_6_, npu_inst_pe_1_4_3_sub_77_carry_5_,
         npu_inst_pe_1_4_3_sub_77_carry_4_, npu_inst_pe_1_4_3_sub_77_carry_3_,
         npu_inst_pe_1_4_3_sub_77_carry_2_, npu_inst_pe_1_4_3_sub_77_carry_1_,
         npu_inst_pe_1_4_3_add_79_carry_7_, npu_inst_pe_1_4_3_add_79_carry_6_,
         npu_inst_pe_1_4_3_add_79_carry_5_, npu_inst_pe_1_4_3_add_79_carry_4_,
         npu_inst_pe_1_4_3_add_79_carry_3_, npu_inst_pe_1_4_3_add_79_carry_2_,
         npu_inst_pe_1_4_3_add_79_carry_1_, npu_inst_pe_1_4_3_n97,
         npu_inst_pe_1_4_3_n96, npu_inst_pe_1_4_3_n95, npu_inst_pe_1_4_3_n94,
         npu_inst_pe_1_4_3_n93, npu_inst_pe_1_4_3_n92, npu_inst_pe_1_4_3_n91,
         npu_inst_pe_1_4_3_n90, npu_inst_pe_1_4_3_n89, npu_inst_pe_1_4_3_n88,
         npu_inst_pe_1_4_3_n87, npu_inst_pe_1_4_3_n86, npu_inst_pe_1_4_3_n85,
         npu_inst_pe_1_4_3_n84, npu_inst_pe_1_4_3_n83, npu_inst_pe_1_4_3_n82,
         npu_inst_pe_1_4_3_n81, npu_inst_pe_1_4_3_n80, npu_inst_pe_1_4_3_n79,
         npu_inst_pe_1_4_3_n78, npu_inst_pe_1_4_3_n77, npu_inst_pe_1_4_3_n76,
         npu_inst_pe_1_4_3_n75, npu_inst_pe_1_4_3_n74, npu_inst_pe_1_4_3_n73,
         npu_inst_pe_1_4_3_n72, npu_inst_pe_1_4_3_n71, npu_inst_pe_1_4_3_n70,
         npu_inst_pe_1_4_3_n69, npu_inst_pe_1_4_3_n68, npu_inst_pe_1_4_3_n67,
         npu_inst_pe_1_4_3_n66, npu_inst_pe_1_4_3_n65, npu_inst_pe_1_4_3_n64,
         npu_inst_pe_1_4_3_n63, npu_inst_pe_1_4_3_n62, npu_inst_pe_1_4_3_n61,
         npu_inst_pe_1_4_3_n60, npu_inst_pe_1_4_3_n59, npu_inst_pe_1_4_3_n58,
         npu_inst_pe_1_4_3_n57, npu_inst_pe_1_4_3_n56, npu_inst_pe_1_4_3_n55,
         npu_inst_pe_1_4_3_n54, npu_inst_pe_1_4_3_n53, npu_inst_pe_1_4_3_n52,
         npu_inst_pe_1_4_3_n51, npu_inst_pe_1_4_3_n50, npu_inst_pe_1_4_3_n49,
         npu_inst_pe_1_4_3_n48, npu_inst_pe_1_4_3_n47, npu_inst_pe_1_4_3_n46,
         npu_inst_pe_1_4_3_n45, npu_inst_pe_1_4_3_n44, npu_inst_pe_1_4_3_n43,
         npu_inst_pe_1_4_3_n42, npu_inst_pe_1_4_3_n41, npu_inst_pe_1_4_3_n40,
         npu_inst_pe_1_4_3_n39, npu_inst_pe_1_4_3_n38, npu_inst_pe_1_4_3_n37,
         npu_inst_pe_1_4_3_n27, npu_inst_pe_1_4_3_n26,
         npu_inst_pe_1_4_3_net3494, npu_inst_pe_1_4_3_net3488,
         npu_inst_pe_1_4_3_N94, npu_inst_pe_1_4_3_N93, npu_inst_pe_1_4_3_N84,
         npu_inst_pe_1_4_3_N80, npu_inst_pe_1_4_3_N79, npu_inst_pe_1_4_3_N78,
         npu_inst_pe_1_4_3_N77, npu_inst_pe_1_4_3_N76, npu_inst_pe_1_4_3_N75,
         npu_inst_pe_1_4_3_N74, npu_inst_pe_1_4_3_N73, npu_inst_pe_1_4_3_N72,
         npu_inst_pe_1_4_3_N71, npu_inst_pe_1_4_3_N70, npu_inst_pe_1_4_3_N69,
         npu_inst_pe_1_4_3_N68, npu_inst_pe_1_4_3_N67, npu_inst_pe_1_4_3_N66,
         npu_inst_pe_1_4_3_N65, npu_inst_pe_1_4_3_int_q_acc_0_,
         npu_inst_pe_1_4_3_int_q_acc_1_, npu_inst_pe_1_4_3_int_q_acc_2_,
         npu_inst_pe_1_4_3_int_q_acc_3_, npu_inst_pe_1_4_3_int_q_acc_4_,
         npu_inst_pe_1_4_3_int_q_acc_5_, npu_inst_pe_1_4_3_int_q_acc_6_,
         npu_inst_pe_1_4_3_int_q_acc_7_, npu_inst_pe_1_4_3_int_data_0_,
         npu_inst_pe_1_4_3_int_data_1_, npu_inst_pe_1_4_3_int_q_weight_0_,
         npu_inst_pe_1_4_3_int_q_weight_1_,
         npu_inst_pe_1_4_3_int_q_reg_v_5__0_,
         npu_inst_pe_1_4_3_int_q_reg_v_5__1_,
         npu_inst_pe_1_4_3_int_q_reg_v_4__0_,
         npu_inst_pe_1_4_3_int_q_reg_v_4__1_,
         npu_inst_pe_1_4_3_int_q_reg_v_3__0_,
         npu_inst_pe_1_4_3_int_q_reg_v_3__1_,
         npu_inst_pe_1_4_3_int_q_reg_v_2__0_,
         npu_inst_pe_1_4_3_int_q_reg_v_2__1_,
         npu_inst_pe_1_4_3_int_q_reg_v_1__0_,
         npu_inst_pe_1_4_3_int_q_reg_v_1__1_,
         npu_inst_pe_1_4_3_int_q_reg_v_0__0_,
         npu_inst_pe_1_4_3_int_q_reg_v_0__1_,
         npu_inst_pe_1_4_3_int_q_reg_h_5__0_,
         npu_inst_pe_1_4_3_int_q_reg_h_5__1_,
         npu_inst_pe_1_4_3_int_q_reg_h_4__0_,
         npu_inst_pe_1_4_3_int_q_reg_h_4__1_,
         npu_inst_pe_1_4_3_int_q_reg_h_3__0_,
         npu_inst_pe_1_4_3_int_q_reg_h_3__1_,
         npu_inst_pe_1_4_3_int_q_reg_h_2__0_,
         npu_inst_pe_1_4_3_int_q_reg_h_2__1_,
         npu_inst_pe_1_4_3_int_q_reg_h_1__0_,
         npu_inst_pe_1_4_3_int_q_reg_h_1__1_,
         npu_inst_pe_1_4_3_int_q_reg_h_0__0_,
         npu_inst_pe_1_4_3_int_q_reg_h_0__1_, npu_inst_pe_1_4_4_n119,
         npu_inst_pe_1_4_4_n118, npu_inst_pe_1_4_4_n117,
         npu_inst_pe_1_4_4_n116, npu_inst_pe_1_4_4_n115,
         npu_inst_pe_1_4_4_n114, npu_inst_pe_1_4_4_n113,
         npu_inst_pe_1_4_4_n112, npu_inst_pe_1_4_4_n111,
         npu_inst_pe_1_4_4_n110, npu_inst_pe_1_4_4_n109,
         npu_inst_pe_1_4_4_n108, npu_inst_pe_1_4_4_n107,
         npu_inst_pe_1_4_4_n106, npu_inst_pe_1_4_4_n105,
         npu_inst_pe_1_4_4_n104, npu_inst_pe_1_4_4_n103,
         npu_inst_pe_1_4_4_n102, npu_inst_pe_1_4_4_n101,
         npu_inst_pe_1_4_4_n100, npu_inst_pe_1_4_4_n99, npu_inst_pe_1_4_4_n98,
         npu_inst_pe_1_4_4_n36, npu_inst_pe_1_4_4_n35, npu_inst_pe_1_4_4_n34,
         npu_inst_pe_1_4_4_n33, npu_inst_pe_1_4_4_n32, npu_inst_pe_1_4_4_n31,
         npu_inst_pe_1_4_4_n30, npu_inst_pe_1_4_4_n29, npu_inst_pe_1_4_4_n28,
         npu_inst_pe_1_4_4_n25, npu_inst_pe_1_4_4_n24, npu_inst_pe_1_4_4_n23,
         npu_inst_pe_1_4_4_n22, npu_inst_pe_1_4_4_n21, npu_inst_pe_1_4_4_n20,
         npu_inst_pe_1_4_4_n19, npu_inst_pe_1_4_4_n18, npu_inst_pe_1_4_4_n17,
         npu_inst_pe_1_4_4_n16, npu_inst_pe_1_4_4_n15, npu_inst_pe_1_4_4_n14,
         npu_inst_pe_1_4_4_n13, npu_inst_pe_1_4_4_n12, npu_inst_pe_1_4_4_n11,
         npu_inst_pe_1_4_4_n10, npu_inst_pe_1_4_4_n9, npu_inst_pe_1_4_4_n8,
         npu_inst_pe_1_4_4_n7, npu_inst_pe_1_4_4_n6, npu_inst_pe_1_4_4_n5,
         npu_inst_pe_1_4_4_n4, npu_inst_pe_1_4_4_n3, npu_inst_pe_1_4_4_n2,
         npu_inst_pe_1_4_4_n1, npu_inst_pe_1_4_4_sub_77_carry_7_,
         npu_inst_pe_1_4_4_sub_77_carry_6_, npu_inst_pe_1_4_4_sub_77_carry_5_,
         npu_inst_pe_1_4_4_sub_77_carry_4_, npu_inst_pe_1_4_4_sub_77_carry_3_,
         npu_inst_pe_1_4_4_sub_77_carry_2_, npu_inst_pe_1_4_4_sub_77_carry_1_,
         npu_inst_pe_1_4_4_add_79_carry_7_, npu_inst_pe_1_4_4_add_79_carry_6_,
         npu_inst_pe_1_4_4_add_79_carry_5_, npu_inst_pe_1_4_4_add_79_carry_4_,
         npu_inst_pe_1_4_4_add_79_carry_3_, npu_inst_pe_1_4_4_add_79_carry_2_,
         npu_inst_pe_1_4_4_add_79_carry_1_, npu_inst_pe_1_4_4_n97,
         npu_inst_pe_1_4_4_n96, npu_inst_pe_1_4_4_n95, npu_inst_pe_1_4_4_n94,
         npu_inst_pe_1_4_4_n93, npu_inst_pe_1_4_4_n92, npu_inst_pe_1_4_4_n91,
         npu_inst_pe_1_4_4_n90, npu_inst_pe_1_4_4_n89, npu_inst_pe_1_4_4_n88,
         npu_inst_pe_1_4_4_n87, npu_inst_pe_1_4_4_n86, npu_inst_pe_1_4_4_n85,
         npu_inst_pe_1_4_4_n84, npu_inst_pe_1_4_4_n83, npu_inst_pe_1_4_4_n82,
         npu_inst_pe_1_4_4_n81, npu_inst_pe_1_4_4_n80, npu_inst_pe_1_4_4_n79,
         npu_inst_pe_1_4_4_n78, npu_inst_pe_1_4_4_n77, npu_inst_pe_1_4_4_n76,
         npu_inst_pe_1_4_4_n75, npu_inst_pe_1_4_4_n74, npu_inst_pe_1_4_4_n73,
         npu_inst_pe_1_4_4_n72, npu_inst_pe_1_4_4_n71, npu_inst_pe_1_4_4_n70,
         npu_inst_pe_1_4_4_n69, npu_inst_pe_1_4_4_n68, npu_inst_pe_1_4_4_n67,
         npu_inst_pe_1_4_4_n66, npu_inst_pe_1_4_4_n65, npu_inst_pe_1_4_4_n64,
         npu_inst_pe_1_4_4_n63, npu_inst_pe_1_4_4_n62, npu_inst_pe_1_4_4_n61,
         npu_inst_pe_1_4_4_n60, npu_inst_pe_1_4_4_n59, npu_inst_pe_1_4_4_n58,
         npu_inst_pe_1_4_4_n57, npu_inst_pe_1_4_4_n56, npu_inst_pe_1_4_4_n55,
         npu_inst_pe_1_4_4_n54, npu_inst_pe_1_4_4_n53, npu_inst_pe_1_4_4_n52,
         npu_inst_pe_1_4_4_n51, npu_inst_pe_1_4_4_n50, npu_inst_pe_1_4_4_n49,
         npu_inst_pe_1_4_4_n48, npu_inst_pe_1_4_4_n47, npu_inst_pe_1_4_4_n46,
         npu_inst_pe_1_4_4_n45, npu_inst_pe_1_4_4_n44, npu_inst_pe_1_4_4_n43,
         npu_inst_pe_1_4_4_n42, npu_inst_pe_1_4_4_n41, npu_inst_pe_1_4_4_n40,
         npu_inst_pe_1_4_4_n39, npu_inst_pe_1_4_4_n38, npu_inst_pe_1_4_4_n37,
         npu_inst_pe_1_4_4_n27, npu_inst_pe_1_4_4_n26,
         npu_inst_pe_1_4_4_net3471, npu_inst_pe_1_4_4_net3465,
         npu_inst_pe_1_4_4_N94, npu_inst_pe_1_4_4_N93, npu_inst_pe_1_4_4_N84,
         npu_inst_pe_1_4_4_N80, npu_inst_pe_1_4_4_N79, npu_inst_pe_1_4_4_N78,
         npu_inst_pe_1_4_4_N77, npu_inst_pe_1_4_4_N76, npu_inst_pe_1_4_4_N75,
         npu_inst_pe_1_4_4_N74, npu_inst_pe_1_4_4_N73, npu_inst_pe_1_4_4_N72,
         npu_inst_pe_1_4_4_N71, npu_inst_pe_1_4_4_N70, npu_inst_pe_1_4_4_N69,
         npu_inst_pe_1_4_4_N68, npu_inst_pe_1_4_4_N67, npu_inst_pe_1_4_4_N66,
         npu_inst_pe_1_4_4_N65, npu_inst_pe_1_4_4_int_q_acc_0_,
         npu_inst_pe_1_4_4_int_q_acc_1_, npu_inst_pe_1_4_4_int_q_acc_2_,
         npu_inst_pe_1_4_4_int_q_acc_3_, npu_inst_pe_1_4_4_int_q_acc_4_,
         npu_inst_pe_1_4_4_int_q_acc_5_, npu_inst_pe_1_4_4_int_q_acc_6_,
         npu_inst_pe_1_4_4_int_q_acc_7_, npu_inst_pe_1_4_4_int_data_0_,
         npu_inst_pe_1_4_4_int_data_1_, npu_inst_pe_1_4_4_int_q_weight_0_,
         npu_inst_pe_1_4_4_int_q_weight_1_,
         npu_inst_pe_1_4_4_int_q_reg_v_5__0_,
         npu_inst_pe_1_4_4_int_q_reg_v_5__1_,
         npu_inst_pe_1_4_4_int_q_reg_v_4__0_,
         npu_inst_pe_1_4_4_int_q_reg_v_4__1_,
         npu_inst_pe_1_4_4_int_q_reg_v_3__0_,
         npu_inst_pe_1_4_4_int_q_reg_v_3__1_,
         npu_inst_pe_1_4_4_int_q_reg_v_2__0_,
         npu_inst_pe_1_4_4_int_q_reg_v_2__1_,
         npu_inst_pe_1_4_4_int_q_reg_v_1__0_,
         npu_inst_pe_1_4_4_int_q_reg_v_1__1_,
         npu_inst_pe_1_4_4_int_q_reg_v_0__0_,
         npu_inst_pe_1_4_4_int_q_reg_v_0__1_,
         npu_inst_pe_1_4_4_int_q_reg_h_5__0_,
         npu_inst_pe_1_4_4_int_q_reg_h_5__1_,
         npu_inst_pe_1_4_4_int_q_reg_h_4__0_,
         npu_inst_pe_1_4_4_int_q_reg_h_4__1_,
         npu_inst_pe_1_4_4_int_q_reg_h_3__0_,
         npu_inst_pe_1_4_4_int_q_reg_h_3__1_,
         npu_inst_pe_1_4_4_int_q_reg_h_2__0_,
         npu_inst_pe_1_4_4_int_q_reg_h_2__1_,
         npu_inst_pe_1_4_4_int_q_reg_h_1__0_,
         npu_inst_pe_1_4_4_int_q_reg_h_1__1_,
         npu_inst_pe_1_4_4_int_q_reg_h_0__0_,
         npu_inst_pe_1_4_4_int_q_reg_h_0__1_, npu_inst_pe_1_4_5_n119,
         npu_inst_pe_1_4_5_n118, npu_inst_pe_1_4_5_n117,
         npu_inst_pe_1_4_5_n116, npu_inst_pe_1_4_5_n115,
         npu_inst_pe_1_4_5_n114, npu_inst_pe_1_4_5_n113,
         npu_inst_pe_1_4_5_n112, npu_inst_pe_1_4_5_n111,
         npu_inst_pe_1_4_5_n110, npu_inst_pe_1_4_5_n109,
         npu_inst_pe_1_4_5_n108, npu_inst_pe_1_4_5_n107,
         npu_inst_pe_1_4_5_n106, npu_inst_pe_1_4_5_n105,
         npu_inst_pe_1_4_5_n104, npu_inst_pe_1_4_5_n103,
         npu_inst_pe_1_4_5_n102, npu_inst_pe_1_4_5_n101,
         npu_inst_pe_1_4_5_n100, npu_inst_pe_1_4_5_n99, npu_inst_pe_1_4_5_n98,
         npu_inst_pe_1_4_5_n36, npu_inst_pe_1_4_5_n35, npu_inst_pe_1_4_5_n34,
         npu_inst_pe_1_4_5_n33, npu_inst_pe_1_4_5_n32, npu_inst_pe_1_4_5_n31,
         npu_inst_pe_1_4_5_n30, npu_inst_pe_1_4_5_n29, npu_inst_pe_1_4_5_n28,
         npu_inst_pe_1_4_5_n25, npu_inst_pe_1_4_5_n24, npu_inst_pe_1_4_5_n23,
         npu_inst_pe_1_4_5_n22, npu_inst_pe_1_4_5_n21, npu_inst_pe_1_4_5_n20,
         npu_inst_pe_1_4_5_n19, npu_inst_pe_1_4_5_n18, npu_inst_pe_1_4_5_n17,
         npu_inst_pe_1_4_5_n16, npu_inst_pe_1_4_5_n15, npu_inst_pe_1_4_5_n14,
         npu_inst_pe_1_4_5_n13, npu_inst_pe_1_4_5_n12, npu_inst_pe_1_4_5_n11,
         npu_inst_pe_1_4_5_n10, npu_inst_pe_1_4_5_n9, npu_inst_pe_1_4_5_n8,
         npu_inst_pe_1_4_5_n7, npu_inst_pe_1_4_5_n6, npu_inst_pe_1_4_5_n5,
         npu_inst_pe_1_4_5_n4, npu_inst_pe_1_4_5_n3, npu_inst_pe_1_4_5_n2,
         npu_inst_pe_1_4_5_n1, npu_inst_pe_1_4_5_sub_77_carry_7_,
         npu_inst_pe_1_4_5_sub_77_carry_6_, npu_inst_pe_1_4_5_sub_77_carry_5_,
         npu_inst_pe_1_4_5_sub_77_carry_4_, npu_inst_pe_1_4_5_sub_77_carry_3_,
         npu_inst_pe_1_4_5_sub_77_carry_2_, npu_inst_pe_1_4_5_sub_77_carry_1_,
         npu_inst_pe_1_4_5_add_79_carry_7_, npu_inst_pe_1_4_5_add_79_carry_6_,
         npu_inst_pe_1_4_5_add_79_carry_5_, npu_inst_pe_1_4_5_add_79_carry_4_,
         npu_inst_pe_1_4_5_add_79_carry_3_, npu_inst_pe_1_4_5_add_79_carry_2_,
         npu_inst_pe_1_4_5_add_79_carry_1_, npu_inst_pe_1_4_5_n97,
         npu_inst_pe_1_4_5_n96, npu_inst_pe_1_4_5_n95, npu_inst_pe_1_4_5_n94,
         npu_inst_pe_1_4_5_n93, npu_inst_pe_1_4_5_n92, npu_inst_pe_1_4_5_n91,
         npu_inst_pe_1_4_5_n90, npu_inst_pe_1_4_5_n89, npu_inst_pe_1_4_5_n88,
         npu_inst_pe_1_4_5_n87, npu_inst_pe_1_4_5_n86, npu_inst_pe_1_4_5_n85,
         npu_inst_pe_1_4_5_n84, npu_inst_pe_1_4_5_n83, npu_inst_pe_1_4_5_n82,
         npu_inst_pe_1_4_5_n81, npu_inst_pe_1_4_5_n80, npu_inst_pe_1_4_5_n79,
         npu_inst_pe_1_4_5_n78, npu_inst_pe_1_4_5_n77, npu_inst_pe_1_4_5_n76,
         npu_inst_pe_1_4_5_n75, npu_inst_pe_1_4_5_n74, npu_inst_pe_1_4_5_n73,
         npu_inst_pe_1_4_5_n72, npu_inst_pe_1_4_5_n71, npu_inst_pe_1_4_5_n70,
         npu_inst_pe_1_4_5_n69, npu_inst_pe_1_4_5_n68, npu_inst_pe_1_4_5_n67,
         npu_inst_pe_1_4_5_n66, npu_inst_pe_1_4_5_n65, npu_inst_pe_1_4_5_n64,
         npu_inst_pe_1_4_5_n63, npu_inst_pe_1_4_5_n62, npu_inst_pe_1_4_5_n61,
         npu_inst_pe_1_4_5_n60, npu_inst_pe_1_4_5_n59, npu_inst_pe_1_4_5_n58,
         npu_inst_pe_1_4_5_n57, npu_inst_pe_1_4_5_n56, npu_inst_pe_1_4_5_n55,
         npu_inst_pe_1_4_5_n54, npu_inst_pe_1_4_5_n53, npu_inst_pe_1_4_5_n52,
         npu_inst_pe_1_4_5_n51, npu_inst_pe_1_4_5_n50, npu_inst_pe_1_4_5_n49,
         npu_inst_pe_1_4_5_n48, npu_inst_pe_1_4_5_n47, npu_inst_pe_1_4_5_n46,
         npu_inst_pe_1_4_5_n45, npu_inst_pe_1_4_5_n44, npu_inst_pe_1_4_5_n43,
         npu_inst_pe_1_4_5_n42, npu_inst_pe_1_4_5_n41, npu_inst_pe_1_4_5_n40,
         npu_inst_pe_1_4_5_n39, npu_inst_pe_1_4_5_n38, npu_inst_pe_1_4_5_n37,
         npu_inst_pe_1_4_5_n27, npu_inst_pe_1_4_5_n26,
         npu_inst_pe_1_4_5_net3448, npu_inst_pe_1_4_5_net3442,
         npu_inst_pe_1_4_5_N94, npu_inst_pe_1_4_5_N93, npu_inst_pe_1_4_5_N84,
         npu_inst_pe_1_4_5_N80, npu_inst_pe_1_4_5_N79, npu_inst_pe_1_4_5_N78,
         npu_inst_pe_1_4_5_N77, npu_inst_pe_1_4_5_N76, npu_inst_pe_1_4_5_N75,
         npu_inst_pe_1_4_5_N74, npu_inst_pe_1_4_5_N73, npu_inst_pe_1_4_5_N72,
         npu_inst_pe_1_4_5_N71, npu_inst_pe_1_4_5_N70, npu_inst_pe_1_4_5_N69,
         npu_inst_pe_1_4_5_N68, npu_inst_pe_1_4_5_N67, npu_inst_pe_1_4_5_N66,
         npu_inst_pe_1_4_5_N65, npu_inst_pe_1_4_5_int_q_acc_0_,
         npu_inst_pe_1_4_5_int_q_acc_1_, npu_inst_pe_1_4_5_int_q_acc_2_,
         npu_inst_pe_1_4_5_int_q_acc_3_, npu_inst_pe_1_4_5_int_q_acc_4_,
         npu_inst_pe_1_4_5_int_q_acc_5_, npu_inst_pe_1_4_5_int_q_acc_6_,
         npu_inst_pe_1_4_5_int_q_acc_7_, npu_inst_pe_1_4_5_int_data_0_,
         npu_inst_pe_1_4_5_int_data_1_, npu_inst_pe_1_4_5_int_q_weight_0_,
         npu_inst_pe_1_4_5_int_q_weight_1_,
         npu_inst_pe_1_4_5_int_q_reg_v_5__0_,
         npu_inst_pe_1_4_5_int_q_reg_v_5__1_,
         npu_inst_pe_1_4_5_int_q_reg_v_4__0_,
         npu_inst_pe_1_4_5_int_q_reg_v_4__1_,
         npu_inst_pe_1_4_5_int_q_reg_v_3__0_,
         npu_inst_pe_1_4_5_int_q_reg_v_3__1_,
         npu_inst_pe_1_4_5_int_q_reg_v_2__0_,
         npu_inst_pe_1_4_5_int_q_reg_v_2__1_,
         npu_inst_pe_1_4_5_int_q_reg_v_1__0_,
         npu_inst_pe_1_4_5_int_q_reg_v_1__1_,
         npu_inst_pe_1_4_5_int_q_reg_v_0__0_,
         npu_inst_pe_1_4_5_int_q_reg_v_0__1_,
         npu_inst_pe_1_4_5_int_q_reg_h_5__0_,
         npu_inst_pe_1_4_5_int_q_reg_h_5__1_,
         npu_inst_pe_1_4_5_int_q_reg_h_4__0_,
         npu_inst_pe_1_4_5_int_q_reg_h_4__1_,
         npu_inst_pe_1_4_5_int_q_reg_h_3__0_,
         npu_inst_pe_1_4_5_int_q_reg_h_3__1_,
         npu_inst_pe_1_4_5_int_q_reg_h_2__0_,
         npu_inst_pe_1_4_5_int_q_reg_h_2__1_,
         npu_inst_pe_1_4_5_int_q_reg_h_1__0_,
         npu_inst_pe_1_4_5_int_q_reg_h_1__1_,
         npu_inst_pe_1_4_5_int_q_reg_h_0__0_,
         npu_inst_pe_1_4_5_int_q_reg_h_0__1_, npu_inst_pe_1_4_6_n119,
         npu_inst_pe_1_4_6_n118, npu_inst_pe_1_4_6_n117,
         npu_inst_pe_1_4_6_n116, npu_inst_pe_1_4_6_n115,
         npu_inst_pe_1_4_6_n114, npu_inst_pe_1_4_6_n113,
         npu_inst_pe_1_4_6_n112, npu_inst_pe_1_4_6_n111,
         npu_inst_pe_1_4_6_n110, npu_inst_pe_1_4_6_n109,
         npu_inst_pe_1_4_6_n108, npu_inst_pe_1_4_6_n107,
         npu_inst_pe_1_4_6_n106, npu_inst_pe_1_4_6_n105,
         npu_inst_pe_1_4_6_n104, npu_inst_pe_1_4_6_n103,
         npu_inst_pe_1_4_6_n102, npu_inst_pe_1_4_6_n101,
         npu_inst_pe_1_4_6_n100, npu_inst_pe_1_4_6_n99, npu_inst_pe_1_4_6_n98,
         npu_inst_pe_1_4_6_n36, npu_inst_pe_1_4_6_n35, npu_inst_pe_1_4_6_n34,
         npu_inst_pe_1_4_6_n33, npu_inst_pe_1_4_6_n32, npu_inst_pe_1_4_6_n31,
         npu_inst_pe_1_4_6_n30, npu_inst_pe_1_4_6_n29, npu_inst_pe_1_4_6_n28,
         npu_inst_pe_1_4_6_n25, npu_inst_pe_1_4_6_n24, npu_inst_pe_1_4_6_n23,
         npu_inst_pe_1_4_6_n22, npu_inst_pe_1_4_6_n21, npu_inst_pe_1_4_6_n20,
         npu_inst_pe_1_4_6_n19, npu_inst_pe_1_4_6_n18, npu_inst_pe_1_4_6_n17,
         npu_inst_pe_1_4_6_n16, npu_inst_pe_1_4_6_n15, npu_inst_pe_1_4_6_n14,
         npu_inst_pe_1_4_6_n13, npu_inst_pe_1_4_6_n12, npu_inst_pe_1_4_6_n11,
         npu_inst_pe_1_4_6_n10, npu_inst_pe_1_4_6_n9, npu_inst_pe_1_4_6_n8,
         npu_inst_pe_1_4_6_n7, npu_inst_pe_1_4_6_n6, npu_inst_pe_1_4_6_n5,
         npu_inst_pe_1_4_6_n4, npu_inst_pe_1_4_6_n3, npu_inst_pe_1_4_6_n2,
         npu_inst_pe_1_4_6_n1, npu_inst_pe_1_4_6_sub_77_carry_7_,
         npu_inst_pe_1_4_6_sub_77_carry_6_, npu_inst_pe_1_4_6_sub_77_carry_5_,
         npu_inst_pe_1_4_6_sub_77_carry_4_, npu_inst_pe_1_4_6_sub_77_carry_3_,
         npu_inst_pe_1_4_6_sub_77_carry_2_, npu_inst_pe_1_4_6_sub_77_carry_1_,
         npu_inst_pe_1_4_6_add_79_carry_7_, npu_inst_pe_1_4_6_add_79_carry_6_,
         npu_inst_pe_1_4_6_add_79_carry_5_, npu_inst_pe_1_4_6_add_79_carry_4_,
         npu_inst_pe_1_4_6_add_79_carry_3_, npu_inst_pe_1_4_6_add_79_carry_2_,
         npu_inst_pe_1_4_6_add_79_carry_1_, npu_inst_pe_1_4_6_n97,
         npu_inst_pe_1_4_6_n96, npu_inst_pe_1_4_6_n95, npu_inst_pe_1_4_6_n94,
         npu_inst_pe_1_4_6_n93, npu_inst_pe_1_4_6_n92, npu_inst_pe_1_4_6_n91,
         npu_inst_pe_1_4_6_n90, npu_inst_pe_1_4_6_n89, npu_inst_pe_1_4_6_n88,
         npu_inst_pe_1_4_6_n87, npu_inst_pe_1_4_6_n86, npu_inst_pe_1_4_6_n85,
         npu_inst_pe_1_4_6_n84, npu_inst_pe_1_4_6_n83, npu_inst_pe_1_4_6_n82,
         npu_inst_pe_1_4_6_n81, npu_inst_pe_1_4_6_n80, npu_inst_pe_1_4_6_n79,
         npu_inst_pe_1_4_6_n78, npu_inst_pe_1_4_6_n77, npu_inst_pe_1_4_6_n76,
         npu_inst_pe_1_4_6_n75, npu_inst_pe_1_4_6_n74, npu_inst_pe_1_4_6_n73,
         npu_inst_pe_1_4_6_n72, npu_inst_pe_1_4_6_n71, npu_inst_pe_1_4_6_n70,
         npu_inst_pe_1_4_6_n69, npu_inst_pe_1_4_6_n68, npu_inst_pe_1_4_6_n67,
         npu_inst_pe_1_4_6_n66, npu_inst_pe_1_4_6_n65, npu_inst_pe_1_4_6_n64,
         npu_inst_pe_1_4_6_n63, npu_inst_pe_1_4_6_n62, npu_inst_pe_1_4_6_n61,
         npu_inst_pe_1_4_6_n60, npu_inst_pe_1_4_6_n59, npu_inst_pe_1_4_6_n58,
         npu_inst_pe_1_4_6_n57, npu_inst_pe_1_4_6_n56, npu_inst_pe_1_4_6_n55,
         npu_inst_pe_1_4_6_n54, npu_inst_pe_1_4_6_n53, npu_inst_pe_1_4_6_n52,
         npu_inst_pe_1_4_6_n51, npu_inst_pe_1_4_6_n50, npu_inst_pe_1_4_6_n49,
         npu_inst_pe_1_4_6_n48, npu_inst_pe_1_4_6_n47, npu_inst_pe_1_4_6_n46,
         npu_inst_pe_1_4_6_n45, npu_inst_pe_1_4_6_n44, npu_inst_pe_1_4_6_n43,
         npu_inst_pe_1_4_6_n42, npu_inst_pe_1_4_6_n41, npu_inst_pe_1_4_6_n40,
         npu_inst_pe_1_4_6_n39, npu_inst_pe_1_4_6_n38, npu_inst_pe_1_4_6_n37,
         npu_inst_pe_1_4_6_n27, npu_inst_pe_1_4_6_n26,
         npu_inst_pe_1_4_6_net3425, npu_inst_pe_1_4_6_net3419,
         npu_inst_pe_1_4_6_N94, npu_inst_pe_1_4_6_N93, npu_inst_pe_1_4_6_N84,
         npu_inst_pe_1_4_6_N80, npu_inst_pe_1_4_6_N79, npu_inst_pe_1_4_6_N78,
         npu_inst_pe_1_4_6_N77, npu_inst_pe_1_4_6_N76, npu_inst_pe_1_4_6_N75,
         npu_inst_pe_1_4_6_N74, npu_inst_pe_1_4_6_N73, npu_inst_pe_1_4_6_N72,
         npu_inst_pe_1_4_6_N71, npu_inst_pe_1_4_6_N70, npu_inst_pe_1_4_6_N69,
         npu_inst_pe_1_4_6_N68, npu_inst_pe_1_4_6_N67, npu_inst_pe_1_4_6_N66,
         npu_inst_pe_1_4_6_N65, npu_inst_pe_1_4_6_int_q_acc_0_,
         npu_inst_pe_1_4_6_int_q_acc_1_, npu_inst_pe_1_4_6_int_q_acc_2_,
         npu_inst_pe_1_4_6_int_q_acc_3_, npu_inst_pe_1_4_6_int_q_acc_4_,
         npu_inst_pe_1_4_6_int_q_acc_5_, npu_inst_pe_1_4_6_int_q_acc_6_,
         npu_inst_pe_1_4_6_int_q_acc_7_, npu_inst_pe_1_4_6_int_data_0_,
         npu_inst_pe_1_4_6_int_data_1_, npu_inst_pe_1_4_6_int_q_weight_0_,
         npu_inst_pe_1_4_6_int_q_weight_1_,
         npu_inst_pe_1_4_6_int_q_reg_v_5__0_,
         npu_inst_pe_1_4_6_int_q_reg_v_5__1_,
         npu_inst_pe_1_4_6_int_q_reg_v_4__0_,
         npu_inst_pe_1_4_6_int_q_reg_v_4__1_,
         npu_inst_pe_1_4_6_int_q_reg_v_3__0_,
         npu_inst_pe_1_4_6_int_q_reg_v_3__1_,
         npu_inst_pe_1_4_6_int_q_reg_v_2__0_,
         npu_inst_pe_1_4_6_int_q_reg_v_2__1_,
         npu_inst_pe_1_4_6_int_q_reg_v_1__0_,
         npu_inst_pe_1_4_6_int_q_reg_v_1__1_,
         npu_inst_pe_1_4_6_int_q_reg_v_0__0_,
         npu_inst_pe_1_4_6_int_q_reg_v_0__1_,
         npu_inst_pe_1_4_6_int_q_reg_h_5__0_,
         npu_inst_pe_1_4_6_int_q_reg_h_5__1_,
         npu_inst_pe_1_4_6_int_q_reg_h_4__0_,
         npu_inst_pe_1_4_6_int_q_reg_h_4__1_,
         npu_inst_pe_1_4_6_int_q_reg_h_3__0_,
         npu_inst_pe_1_4_6_int_q_reg_h_3__1_,
         npu_inst_pe_1_4_6_int_q_reg_h_2__0_,
         npu_inst_pe_1_4_6_int_q_reg_h_2__1_,
         npu_inst_pe_1_4_6_int_q_reg_h_1__0_,
         npu_inst_pe_1_4_6_int_q_reg_h_1__1_,
         npu_inst_pe_1_4_6_int_q_reg_h_0__0_,
         npu_inst_pe_1_4_6_int_q_reg_h_0__1_, npu_inst_pe_1_4_7_n119,
         npu_inst_pe_1_4_7_n118, npu_inst_pe_1_4_7_n117,
         npu_inst_pe_1_4_7_n116, npu_inst_pe_1_4_7_n115,
         npu_inst_pe_1_4_7_n114, npu_inst_pe_1_4_7_n113,
         npu_inst_pe_1_4_7_n112, npu_inst_pe_1_4_7_n111,
         npu_inst_pe_1_4_7_n110, npu_inst_pe_1_4_7_n109,
         npu_inst_pe_1_4_7_n108, npu_inst_pe_1_4_7_n107,
         npu_inst_pe_1_4_7_n106, npu_inst_pe_1_4_7_n105,
         npu_inst_pe_1_4_7_n104, npu_inst_pe_1_4_7_n103,
         npu_inst_pe_1_4_7_n102, npu_inst_pe_1_4_7_n101,
         npu_inst_pe_1_4_7_n100, npu_inst_pe_1_4_7_n99, npu_inst_pe_1_4_7_n98,
         npu_inst_pe_1_4_7_n36, npu_inst_pe_1_4_7_n35, npu_inst_pe_1_4_7_n34,
         npu_inst_pe_1_4_7_n33, npu_inst_pe_1_4_7_n32, npu_inst_pe_1_4_7_n31,
         npu_inst_pe_1_4_7_n30, npu_inst_pe_1_4_7_n29, npu_inst_pe_1_4_7_n28,
         npu_inst_pe_1_4_7_n25, npu_inst_pe_1_4_7_n24, npu_inst_pe_1_4_7_n23,
         npu_inst_pe_1_4_7_n22, npu_inst_pe_1_4_7_n21, npu_inst_pe_1_4_7_n20,
         npu_inst_pe_1_4_7_n19, npu_inst_pe_1_4_7_n18, npu_inst_pe_1_4_7_n17,
         npu_inst_pe_1_4_7_n16, npu_inst_pe_1_4_7_n15, npu_inst_pe_1_4_7_n14,
         npu_inst_pe_1_4_7_n13, npu_inst_pe_1_4_7_n12, npu_inst_pe_1_4_7_n11,
         npu_inst_pe_1_4_7_n10, npu_inst_pe_1_4_7_n9, npu_inst_pe_1_4_7_n8,
         npu_inst_pe_1_4_7_n7, npu_inst_pe_1_4_7_n6, npu_inst_pe_1_4_7_n5,
         npu_inst_pe_1_4_7_n4, npu_inst_pe_1_4_7_n3, npu_inst_pe_1_4_7_n2,
         npu_inst_pe_1_4_7_n1, npu_inst_pe_1_4_7_sub_77_carry_7_,
         npu_inst_pe_1_4_7_sub_77_carry_6_, npu_inst_pe_1_4_7_sub_77_carry_5_,
         npu_inst_pe_1_4_7_sub_77_carry_4_, npu_inst_pe_1_4_7_sub_77_carry_3_,
         npu_inst_pe_1_4_7_sub_77_carry_2_, npu_inst_pe_1_4_7_sub_77_carry_1_,
         npu_inst_pe_1_4_7_add_79_carry_7_, npu_inst_pe_1_4_7_add_79_carry_6_,
         npu_inst_pe_1_4_7_add_79_carry_5_, npu_inst_pe_1_4_7_add_79_carry_4_,
         npu_inst_pe_1_4_7_add_79_carry_3_, npu_inst_pe_1_4_7_add_79_carry_2_,
         npu_inst_pe_1_4_7_add_79_carry_1_, npu_inst_pe_1_4_7_n97,
         npu_inst_pe_1_4_7_n96, npu_inst_pe_1_4_7_n95, npu_inst_pe_1_4_7_n94,
         npu_inst_pe_1_4_7_n93, npu_inst_pe_1_4_7_n92, npu_inst_pe_1_4_7_n91,
         npu_inst_pe_1_4_7_n90, npu_inst_pe_1_4_7_n89, npu_inst_pe_1_4_7_n88,
         npu_inst_pe_1_4_7_n87, npu_inst_pe_1_4_7_n86, npu_inst_pe_1_4_7_n85,
         npu_inst_pe_1_4_7_n84, npu_inst_pe_1_4_7_n83, npu_inst_pe_1_4_7_n82,
         npu_inst_pe_1_4_7_n81, npu_inst_pe_1_4_7_n80, npu_inst_pe_1_4_7_n79,
         npu_inst_pe_1_4_7_n78, npu_inst_pe_1_4_7_n77, npu_inst_pe_1_4_7_n76,
         npu_inst_pe_1_4_7_n75, npu_inst_pe_1_4_7_n74, npu_inst_pe_1_4_7_n73,
         npu_inst_pe_1_4_7_n72, npu_inst_pe_1_4_7_n71, npu_inst_pe_1_4_7_n70,
         npu_inst_pe_1_4_7_n69, npu_inst_pe_1_4_7_n68, npu_inst_pe_1_4_7_n67,
         npu_inst_pe_1_4_7_n66, npu_inst_pe_1_4_7_n65, npu_inst_pe_1_4_7_n64,
         npu_inst_pe_1_4_7_n63, npu_inst_pe_1_4_7_n62, npu_inst_pe_1_4_7_n61,
         npu_inst_pe_1_4_7_n60, npu_inst_pe_1_4_7_n59, npu_inst_pe_1_4_7_n58,
         npu_inst_pe_1_4_7_n57, npu_inst_pe_1_4_7_n56, npu_inst_pe_1_4_7_n55,
         npu_inst_pe_1_4_7_n54, npu_inst_pe_1_4_7_n53, npu_inst_pe_1_4_7_n52,
         npu_inst_pe_1_4_7_n51, npu_inst_pe_1_4_7_n50, npu_inst_pe_1_4_7_n49,
         npu_inst_pe_1_4_7_n48, npu_inst_pe_1_4_7_n47, npu_inst_pe_1_4_7_n46,
         npu_inst_pe_1_4_7_n45, npu_inst_pe_1_4_7_n44, npu_inst_pe_1_4_7_n43,
         npu_inst_pe_1_4_7_n42, npu_inst_pe_1_4_7_n41, npu_inst_pe_1_4_7_n40,
         npu_inst_pe_1_4_7_n39, npu_inst_pe_1_4_7_n38, npu_inst_pe_1_4_7_n37,
         npu_inst_pe_1_4_7_n27, npu_inst_pe_1_4_7_n26,
         npu_inst_pe_1_4_7_net3402, npu_inst_pe_1_4_7_net3396,
         npu_inst_pe_1_4_7_N94, npu_inst_pe_1_4_7_N93, npu_inst_pe_1_4_7_N84,
         npu_inst_pe_1_4_7_N80, npu_inst_pe_1_4_7_N79, npu_inst_pe_1_4_7_N78,
         npu_inst_pe_1_4_7_N77, npu_inst_pe_1_4_7_N76, npu_inst_pe_1_4_7_N75,
         npu_inst_pe_1_4_7_N74, npu_inst_pe_1_4_7_N73, npu_inst_pe_1_4_7_N72,
         npu_inst_pe_1_4_7_N71, npu_inst_pe_1_4_7_N70, npu_inst_pe_1_4_7_N69,
         npu_inst_pe_1_4_7_N68, npu_inst_pe_1_4_7_N67, npu_inst_pe_1_4_7_N66,
         npu_inst_pe_1_4_7_N65, npu_inst_pe_1_4_7_int_q_acc_0_,
         npu_inst_pe_1_4_7_int_q_acc_1_, npu_inst_pe_1_4_7_int_q_acc_2_,
         npu_inst_pe_1_4_7_int_q_acc_3_, npu_inst_pe_1_4_7_int_q_acc_4_,
         npu_inst_pe_1_4_7_int_q_acc_5_, npu_inst_pe_1_4_7_int_q_acc_6_,
         npu_inst_pe_1_4_7_int_q_acc_7_, npu_inst_pe_1_4_7_int_data_0_,
         npu_inst_pe_1_4_7_int_data_1_, npu_inst_pe_1_4_7_int_q_weight_0_,
         npu_inst_pe_1_4_7_int_q_weight_1_,
         npu_inst_pe_1_4_7_int_q_reg_v_5__0_,
         npu_inst_pe_1_4_7_int_q_reg_v_5__1_,
         npu_inst_pe_1_4_7_int_q_reg_v_4__0_,
         npu_inst_pe_1_4_7_int_q_reg_v_4__1_,
         npu_inst_pe_1_4_7_int_q_reg_v_3__0_,
         npu_inst_pe_1_4_7_int_q_reg_v_3__1_,
         npu_inst_pe_1_4_7_int_q_reg_v_2__0_,
         npu_inst_pe_1_4_7_int_q_reg_v_2__1_,
         npu_inst_pe_1_4_7_int_q_reg_v_1__0_,
         npu_inst_pe_1_4_7_int_q_reg_v_1__1_,
         npu_inst_pe_1_4_7_int_q_reg_v_0__0_,
         npu_inst_pe_1_4_7_int_q_reg_v_0__1_,
         npu_inst_pe_1_4_7_int_q_reg_h_5__0_,
         npu_inst_pe_1_4_7_int_q_reg_h_5__1_,
         npu_inst_pe_1_4_7_int_q_reg_h_4__0_,
         npu_inst_pe_1_4_7_int_q_reg_h_4__1_,
         npu_inst_pe_1_4_7_int_q_reg_h_3__0_,
         npu_inst_pe_1_4_7_int_q_reg_h_3__1_,
         npu_inst_pe_1_4_7_int_q_reg_h_2__0_,
         npu_inst_pe_1_4_7_int_q_reg_h_2__1_,
         npu_inst_pe_1_4_7_int_q_reg_h_1__0_,
         npu_inst_pe_1_4_7_int_q_reg_h_1__1_,
         npu_inst_pe_1_4_7_int_q_reg_h_0__0_,
         npu_inst_pe_1_4_7_int_q_reg_h_0__1_, npu_inst_pe_1_5_0_n118,
         npu_inst_pe_1_5_0_n117, npu_inst_pe_1_5_0_n116,
         npu_inst_pe_1_5_0_n115, npu_inst_pe_1_5_0_n114,
         npu_inst_pe_1_5_0_n113, npu_inst_pe_1_5_0_n112,
         npu_inst_pe_1_5_0_n111, npu_inst_pe_1_5_0_n110,
         npu_inst_pe_1_5_0_n109, npu_inst_pe_1_5_0_n108,
         npu_inst_pe_1_5_0_n107, npu_inst_pe_1_5_0_n106,
         npu_inst_pe_1_5_0_n105, npu_inst_pe_1_5_0_n104,
         npu_inst_pe_1_5_0_n103, npu_inst_pe_1_5_0_n102,
         npu_inst_pe_1_5_0_n101, npu_inst_pe_1_5_0_n100, npu_inst_pe_1_5_0_n99,
         npu_inst_pe_1_5_0_n98, npu_inst_pe_1_5_0_n36, npu_inst_pe_1_5_0_n35,
         npu_inst_pe_1_5_0_n34, npu_inst_pe_1_5_0_n33, npu_inst_pe_1_5_0_n32,
         npu_inst_pe_1_5_0_n31, npu_inst_pe_1_5_0_n30, npu_inst_pe_1_5_0_n29,
         npu_inst_pe_1_5_0_n28, npu_inst_pe_1_5_0_n25, npu_inst_pe_1_5_0_n24,
         npu_inst_pe_1_5_0_n23, npu_inst_pe_1_5_0_n22, npu_inst_pe_1_5_0_n21,
         npu_inst_pe_1_5_0_n20, npu_inst_pe_1_5_0_n19, npu_inst_pe_1_5_0_n18,
         npu_inst_pe_1_5_0_n17, npu_inst_pe_1_5_0_n16, npu_inst_pe_1_5_0_n15,
         npu_inst_pe_1_5_0_n14, npu_inst_pe_1_5_0_n13, npu_inst_pe_1_5_0_n12,
         npu_inst_pe_1_5_0_n11, npu_inst_pe_1_5_0_n10, npu_inst_pe_1_5_0_n9,
         npu_inst_pe_1_5_0_n8, npu_inst_pe_1_5_0_n7, npu_inst_pe_1_5_0_n6,
         npu_inst_pe_1_5_0_n5, npu_inst_pe_1_5_0_n4, npu_inst_pe_1_5_0_n3,
         npu_inst_pe_1_5_0_n2, npu_inst_pe_1_5_0_n1,
         npu_inst_pe_1_5_0_sub_77_carry_7_, npu_inst_pe_1_5_0_sub_77_carry_6_,
         npu_inst_pe_1_5_0_sub_77_carry_5_, npu_inst_pe_1_5_0_sub_77_carry_4_,
         npu_inst_pe_1_5_0_sub_77_carry_3_, npu_inst_pe_1_5_0_sub_77_carry_2_,
         npu_inst_pe_1_5_0_sub_77_carry_1_, npu_inst_pe_1_5_0_add_79_carry_7_,
         npu_inst_pe_1_5_0_add_79_carry_6_, npu_inst_pe_1_5_0_add_79_carry_5_,
         npu_inst_pe_1_5_0_add_79_carry_4_, npu_inst_pe_1_5_0_add_79_carry_3_,
         npu_inst_pe_1_5_0_add_79_carry_2_, npu_inst_pe_1_5_0_add_79_carry_1_,
         npu_inst_pe_1_5_0_n97, npu_inst_pe_1_5_0_n96, npu_inst_pe_1_5_0_n95,
         npu_inst_pe_1_5_0_n94, npu_inst_pe_1_5_0_n93, npu_inst_pe_1_5_0_n92,
         npu_inst_pe_1_5_0_n91, npu_inst_pe_1_5_0_n90, npu_inst_pe_1_5_0_n89,
         npu_inst_pe_1_5_0_n88, npu_inst_pe_1_5_0_n87, npu_inst_pe_1_5_0_n86,
         npu_inst_pe_1_5_0_n85, npu_inst_pe_1_5_0_n84, npu_inst_pe_1_5_0_n83,
         npu_inst_pe_1_5_0_n82, npu_inst_pe_1_5_0_n81, npu_inst_pe_1_5_0_n80,
         npu_inst_pe_1_5_0_n79, npu_inst_pe_1_5_0_n78, npu_inst_pe_1_5_0_n77,
         npu_inst_pe_1_5_0_n76, npu_inst_pe_1_5_0_n75, npu_inst_pe_1_5_0_n74,
         npu_inst_pe_1_5_0_n73, npu_inst_pe_1_5_0_n72, npu_inst_pe_1_5_0_n71,
         npu_inst_pe_1_5_0_n70, npu_inst_pe_1_5_0_n69, npu_inst_pe_1_5_0_n68,
         npu_inst_pe_1_5_0_n67, npu_inst_pe_1_5_0_n66, npu_inst_pe_1_5_0_n65,
         npu_inst_pe_1_5_0_n64, npu_inst_pe_1_5_0_n63, npu_inst_pe_1_5_0_n62,
         npu_inst_pe_1_5_0_n61, npu_inst_pe_1_5_0_n60, npu_inst_pe_1_5_0_n59,
         npu_inst_pe_1_5_0_n58, npu_inst_pe_1_5_0_n57, npu_inst_pe_1_5_0_n56,
         npu_inst_pe_1_5_0_n55, npu_inst_pe_1_5_0_n54, npu_inst_pe_1_5_0_n53,
         npu_inst_pe_1_5_0_n52, npu_inst_pe_1_5_0_n51, npu_inst_pe_1_5_0_n50,
         npu_inst_pe_1_5_0_n49, npu_inst_pe_1_5_0_n48, npu_inst_pe_1_5_0_n47,
         npu_inst_pe_1_5_0_n46, npu_inst_pe_1_5_0_n45, npu_inst_pe_1_5_0_n44,
         npu_inst_pe_1_5_0_n43, npu_inst_pe_1_5_0_n42, npu_inst_pe_1_5_0_n41,
         npu_inst_pe_1_5_0_n40, npu_inst_pe_1_5_0_n39, npu_inst_pe_1_5_0_n38,
         npu_inst_pe_1_5_0_n37, npu_inst_pe_1_5_0_n27, npu_inst_pe_1_5_0_n26,
         npu_inst_pe_1_5_0_net3379, npu_inst_pe_1_5_0_net3373,
         npu_inst_pe_1_5_0_N94, npu_inst_pe_1_5_0_N93, npu_inst_pe_1_5_0_N84,
         npu_inst_pe_1_5_0_N80, npu_inst_pe_1_5_0_N79, npu_inst_pe_1_5_0_N78,
         npu_inst_pe_1_5_0_N77, npu_inst_pe_1_5_0_N76, npu_inst_pe_1_5_0_N75,
         npu_inst_pe_1_5_0_N74, npu_inst_pe_1_5_0_N73, npu_inst_pe_1_5_0_N72,
         npu_inst_pe_1_5_0_N71, npu_inst_pe_1_5_0_N70, npu_inst_pe_1_5_0_N69,
         npu_inst_pe_1_5_0_N68, npu_inst_pe_1_5_0_N67, npu_inst_pe_1_5_0_N66,
         npu_inst_pe_1_5_0_N65, npu_inst_pe_1_5_0_int_q_acc_0_,
         npu_inst_pe_1_5_0_int_q_acc_1_, npu_inst_pe_1_5_0_int_q_acc_2_,
         npu_inst_pe_1_5_0_int_q_acc_3_, npu_inst_pe_1_5_0_int_q_acc_4_,
         npu_inst_pe_1_5_0_int_q_acc_5_, npu_inst_pe_1_5_0_int_q_acc_6_,
         npu_inst_pe_1_5_0_int_q_acc_7_, npu_inst_pe_1_5_0_int_data_0_,
         npu_inst_pe_1_5_0_int_data_1_, npu_inst_pe_1_5_0_int_q_weight_0_,
         npu_inst_pe_1_5_0_int_q_weight_1_,
         npu_inst_pe_1_5_0_int_q_reg_v_5__0_,
         npu_inst_pe_1_5_0_int_q_reg_v_5__1_,
         npu_inst_pe_1_5_0_int_q_reg_v_4__0_,
         npu_inst_pe_1_5_0_int_q_reg_v_4__1_,
         npu_inst_pe_1_5_0_int_q_reg_v_3__0_,
         npu_inst_pe_1_5_0_int_q_reg_v_3__1_,
         npu_inst_pe_1_5_0_int_q_reg_v_2__0_,
         npu_inst_pe_1_5_0_int_q_reg_v_2__1_,
         npu_inst_pe_1_5_0_int_q_reg_v_1__0_,
         npu_inst_pe_1_5_0_int_q_reg_v_1__1_,
         npu_inst_pe_1_5_0_int_q_reg_v_0__0_,
         npu_inst_pe_1_5_0_int_q_reg_v_0__1_,
         npu_inst_pe_1_5_0_int_q_reg_h_5__0_,
         npu_inst_pe_1_5_0_int_q_reg_h_5__1_,
         npu_inst_pe_1_5_0_int_q_reg_h_4__0_,
         npu_inst_pe_1_5_0_int_q_reg_h_4__1_,
         npu_inst_pe_1_5_0_int_q_reg_h_3__0_,
         npu_inst_pe_1_5_0_int_q_reg_h_3__1_,
         npu_inst_pe_1_5_0_int_q_reg_h_2__0_,
         npu_inst_pe_1_5_0_int_q_reg_h_2__1_,
         npu_inst_pe_1_5_0_int_q_reg_h_1__0_,
         npu_inst_pe_1_5_0_int_q_reg_h_1__1_,
         npu_inst_pe_1_5_0_int_q_reg_h_0__0_,
         npu_inst_pe_1_5_0_int_q_reg_h_0__1_, npu_inst_pe_1_5_0_o_data_h_0_,
         npu_inst_pe_1_5_0_o_data_h_1_, npu_inst_pe_1_5_1_n119,
         npu_inst_pe_1_5_1_n118, npu_inst_pe_1_5_1_n117,
         npu_inst_pe_1_5_1_n116, npu_inst_pe_1_5_1_n115,
         npu_inst_pe_1_5_1_n114, npu_inst_pe_1_5_1_n113,
         npu_inst_pe_1_5_1_n112, npu_inst_pe_1_5_1_n111,
         npu_inst_pe_1_5_1_n110, npu_inst_pe_1_5_1_n109,
         npu_inst_pe_1_5_1_n108, npu_inst_pe_1_5_1_n107,
         npu_inst_pe_1_5_1_n106, npu_inst_pe_1_5_1_n105,
         npu_inst_pe_1_5_1_n104, npu_inst_pe_1_5_1_n103,
         npu_inst_pe_1_5_1_n102, npu_inst_pe_1_5_1_n101,
         npu_inst_pe_1_5_1_n100, npu_inst_pe_1_5_1_n99, npu_inst_pe_1_5_1_n98,
         npu_inst_pe_1_5_1_n36, npu_inst_pe_1_5_1_n35, npu_inst_pe_1_5_1_n34,
         npu_inst_pe_1_5_1_n33, npu_inst_pe_1_5_1_n32, npu_inst_pe_1_5_1_n31,
         npu_inst_pe_1_5_1_n30, npu_inst_pe_1_5_1_n29, npu_inst_pe_1_5_1_n28,
         npu_inst_pe_1_5_1_n25, npu_inst_pe_1_5_1_n24, npu_inst_pe_1_5_1_n23,
         npu_inst_pe_1_5_1_n22, npu_inst_pe_1_5_1_n21, npu_inst_pe_1_5_1_n20,
         npu_inst_pe_1_5_1_n19, npu_inst_pe_1_5_1_n18, npu_inst_pe_1_5_1_n17,
         npu_inst_pe_1_5_1_n16, npu_inst_pe_1_5_1_n15, npu_inst_pe_1_5_1_n14,
         npu_inst_pe_1_5_1_n13, npu_inst_pe_1_5_1_n12, npu_inst_pe_1_5_1_n11,
         npu_inst_pe_1_5_1_n10, npu_inst_pe_1_5_1_n9, npu_inst_pe_1_5_1_n8,
         npu_inst_pe_1_5_1_n7, npu_inst_pe_1_5_1_n6, npu_inst_pe_1_5_1_n5,
         npu_inst_pe_1_5_1_n4, npu_inst_pe_1_5_1_n3, npu_inst_pe_1_5_1_n2,
         npu_inst_pe_1_5_1_n1, npu_inst_pe_1_5_1_sub_77_carry_7_,
         npu_inst_pe_1_5_1_sub_77_carry_6_, npu_inst_pe_1_5_1_sub_77_carry_5_,
         npu_inst_pe_1_5_1_sub_77_carry_4_, npu_inst_pe_1_5_1_sub_77_carry_3_,
         npu_inst_pe_1_5_1_sub_77_carry_2_, npu_inst_pe_1_5_1_sub_77_carry_1_,
         npu_inst_pe_1_5_1_add_79_carry_7_, npu_inst_pe_1_5_1_add_79_carry_6_,
         npu_inst_pe_1_5_1_add_79_carry_5_, npu_inst_pe_1_5_1_add_79_carry_4_,
         npu_inst_pe_1_5_1_add_79_carry_3_, npu_inst_pe_1_5_1_add_79_carry_2_,
         npu_inst_pe_1_5_1_add_79_carry_1_, npu_inst_pe_1_5_1_n97,
         npu_inst_pe_1_5_1_n96, npu_inst_pe_1_5_1_n95, npu_inst_pe_1_5_1_n94,
         npu_inst_pe_1_5_1_n93, npu_inst_pe_1_5_1_n92, npu_inst_pe_1_5_1_n91,
         npu_inst_pe_1_5_1_n90, npu_inst_pe_1_5_1_n89, npu_inst_pe_1_5_1_n88,
         npu_inst_pe_1_5_1_n87, npu_inst_pe_1_5_1_n86, npu_inst_pe_1_5_1_n85,
         npu_inst_pe_1_5_1_n84, npu_inst_pe_1_5_1_n83, npu_inst_pe_1_5_1_n82,
         npu_inst_pe_1_5_1_n81, npu_inst_pe_1_5_1_n80, npu_inst_pe_1_5_1_n79,
         npu_inst_pe_1_5_1_n78, npu_inst_pe_1_5_1_n77, npu_inst_pe_1_5_1_n76,
         npu_inst_pe_1_5_1_n75, npu_inst_pe_1_5_1_n74, npu_inst_pe_1_5_1_n73,
         npu_inst_pe_1_5_1_n72, npu_inst_pe_1_5_1_n71, npu_inst_pe_1_5_1_n70,
         npu_inst_pe_1_5_1_n69, npu_inst_pe_1_5_1_n68, npu_inst_pe_1_5_1_n67,
         npu_inst_pe_1_5_1_n66, npu_inst_pe_1_5_1_n65, npu_inst_pe_1_5_1_n64,
         npu_inst_pe_1_5_1_n63, npu_inst_pe_1_5_1_n62, npu_inst_pe_1_5_1_n61,
         npu_inst_pe_1_5_1_n60, npu_inst_pe_1_5_1_n59, npu_inst_pe_1_5_1_n58,
         npu_inst_pe_1_5_1_n57, npu_inst_pe_1_5_1_n56, npu_inst_pe_1_5_1_n55,
         npu_inst_pe_1_5_1_n54, npu_inst_pe_1_5_1_n53, npu_inst_pe_1_5_1_n52,
         npu_inst_pe_1_5_1_n51, npu_inst_pe_1_5_1_n50, npu_inst_pe_1_5_1_n49,
         npu_inst_pe_1_5_1_n48, npu_inst_pe_1_5_1_n47, npu_inst_pe_1_5_1_n46,
         npu_inst_pe_1_5_1_n45, npu_inst_pe_1_5_1_n44, npu_inst_pe_1_5_1_n43,
         npu_inst_pe_1_5_1_n42, npu_inst_pe_1_5_1_n41, npu_inst_pe_1_5_1_n40,
         npu_inst_pe_1_5_1_n39, npu_inst_pe_1_5_1_n38, npu_inst_pe_1_5_1_n37,
         npu_inst_pe_1_5_1_n27, npu_inst_pe_1_5_1_n26,
         npu_inst_pe_1_5_1_net3356, npu_inst_pe_1_5_1_net3350,
         npu_inst_pe_1_5_1_N94, npu_inst_pe_1_5_1_N93, npu_inst_pe_1_5_1_N84,
         npu_inst_pe_1_5_1_N80, npu_inst_pe_1_5_1_N79, npu_inst_pe_1_5_1_N78,
         npu_inst_pe_1_5_1_N77, npu_inst_pe_1_5_1_N76, npu_inst_pe_1_5_1_N75,
         npu_inst_pe_1_5_1_N74, npu_inst_pe_1_5_1_N73, npu_inst_pe_1_5_1_N72,
         npu_inst_pe_1_5_1_N71, npu_inst_pe_1_5_1_N70, npu_inst_pe_1_5_1_N69,
         npu_inst_pe_1_5_1_N68, npu_inst_pe_1_5_1_N67, npu_inst_pe_1_5_1_N66,
         npu_inst_pe_1_5_1_N65, npu_inst_pe_1_5_1_int_q_acc_0_,
         npu_inst_pe_1_5_1_int_q_acc_1_, npu_inst_pe_1_5_1_int_q_acc_2_,
         npu_inst_pe_1_5_1_int_q_acc_3_, npu_inst_pe_1_5_1_int_q_acc_4_,
         npu_inst_pe_1_5_1_int_q_acc_5_, npu_inst_pe_1_5_1_int_q_acc_6_,
         npu_inst_pe_1_5_1_int_q_acc_7_, npu_inst_pe_1_5_1_int_data_0_,
         npu_inst_pe_1_5_1_int_data_1_, npu_inst_pe_1_5_1_int_q_weight_0_,
         npu_inst_pe_1_5_1_int_q_weight_1_,
         npu_inst_pe_1_5_1_int_q_reg_v_5__0_,
         npu_inst_pe_1_5_1_int_q_reg_v_5__1_,
         npu_inst_pe_1_5_1_int_q_reg_v_4__0_,
         npu_inst_pe_1_5_1_int_q_reg_v_4__1_,
         npu_inst_pe_1_5_1_int_q_reg_v_3__0_,
         npu_inst_pe_1_5_1_int_q_reg_v_3__1_,
         npu_inst_pe_1_5_1_int_q_reg_v_2__0_,
         npu_inst_pe_1_5_1_int_q_reg_v_2__1_,
         npu_inst_pe_1_5_1_int_q_reg_v_1__0_,
         npu_inst_pe_1_5_1_int_q_reg_v_1__1_,
         npu_inst_pe_1_5_1_int_q_reg_v_0__0_,
         npu_inst_pe_1_5_1_int_q_reg_v_0__1_,
         npu_inst_pe_1_5_1_int_q_reg_h_5__0_,
         npu_inst_pe_1_5_1_int_q_reg_h_5__1_,
         npu_inst_pe_1_5_1_int_q_reg_h_4__0_,
         npu_inst_pe_1_5_1_int_q_reg_h_4__1_,
         npu_inst_pe_1_5_1_int_q_reg_h_3__0_,
         npu_inst_pe_1_5_1_int_q_reg_h_3__1_,
         npu_inst_pe_1_5_1_int_q_reg_h_2__0_,
         npu_inst_pe_1_5_1_int_q_reg_h_2__1_,
         npu_inst_pe_1_5_1_int_q_reg_h_1__0_,
         npu_inst_pe_1_5_1_int_q_reg_h_1__1_,
         npu_inst_pe_1_5_1_int_q_reg_h_0__0_,
         npu_inst_pe_1_5_1_int_q_reg_h_0__1_, npu_inst_pe_1_5_2_n119,
         npu_inst_pe_1_5_2_n118, npu_inst_pe_1_5_2_n117,
         npu_inst_pe_1_5_2_n116, npu_inst_pe_1_5_2_n115,
         npu_inst_pe_1_5_2_n114, npu_inst_pe_1_5_2_n113,
         npu_inst_pe_1_5_2_n112, npu_inst_pe_1_5_2_n111,
         npu_inst_pe_1_5_2_n110, npu_inst_pe_1_5_2_n109,
         npu_inst_pe_1_5_2_n108, npu_inst_pe_1_5_2_n107,
         npu_inst_pe_1_5_2_n106, npu_inst_pe_1_5_2_n105,
         npu_inst_pe_1_5_2_n104, npu_inst_pe_1_5_2_n103,
         npu_inst_pe_1_5_2_n102, npu_inst_pe_1_5_2_n101,
         npu_inst_pe_1_5_2_n100, npu_inst_pe_1_5_2_n99, npu_inst_pe_1_5_2_n98,
         npu_inst_pe_1_5_2_n36, npu_inst_pe_1_5_2_n35, npu_inst_pe_1_5_2_n34,
         npu_inst_pe_1_5_2_n33, npu_inst_pe_1_5_2_n32, npu_inst_pe_1_5_2_n31,
         npu_inst_pe_1_5_2_n30, npu_inst_pe_1_5_2_n29, npu_inst_pe_1_5_2_n28,
         npu_inst_pe_1_5_2_n25, npu_inst_pe_1_5_2_n24, npu_inst_pe_1_5_2_n23,
         npu_inst_pe_1_5_2_n22, npu_inst_pe_1_5_2_n21, npu_inst_pe_1_5_2_n20,
         npu_inst_pe_1_5_2_n19, npu_inst_pe_1_5_2_n18, npu_inst_pe_1_5_2_n17,
         npu_inst_pe_1_5_2_n16, npu_inst_pe_1_5_2_n15, npu_inst_pe_1_5_2_n14,
         npu_inst_pe_1_5_2_n13, npu_inst_pe_1_5_2_n12, npu_inst_pe_1_5_2_n11,
         npu_inst_pe_1_5_2_n10, npu_inst_pe_1_5_2_n9, npu_inst_pe_1_5_2_n8,
         npu_inst_pe_1_5_2_n7, npu_inst_pe_1_5_2_n6, npu_inst_pe_1_5_2_n5,
         npu_inst_pe_1_5_2_n4, npu_inst_pe_1_5_2_n3, npu_inst_pe_1_5_2_n2,
         npu_inst_pe_1_5_2_n1, npu_inst_pe_1_5_2_sub_77_carry_7_,
         npu_inst_pe_1_5_2_sub_77_carry_6_, npu_inst_pe_1_5_2_sub_77_carry_5_,
         npu_inst_pe_1_5_2_sub_77_carry_4_, npu_inst_pe_1_5_2_sub_77_carry_3_,
         npu_inst_pe_1_5_2_sub_77_carry_2_, npu_inst_pe_1_5_2_sub_77_carry_1_,
         npu_inst_pe_1_5_2_add_79_carry_7_, npu_inst_pe_1_5_2_add_79_carry_6_,
         npu_inst_pe_1_5_2_add_79_carry_5_, npu_inst_pe_1_5_2_add_79_carry_4_,
         npu_inst_pe_1_5_2_add_79_carry_3_, npu_inst_pe_1_5_2_add_79_carry_2_,
         npu_inst_pe_1_5_2_add_79_carry_1_, npu_inst_pe_1_5_2_n97,
         npu_inst_pe_1_5_2_n96, npu_inst_pe_1_5_2_n95, npu_inst_pe_1_5_2_n94,
         npu_inst_pe_1_5_2_n93, npu_inst_pe_1_5_2_n92, npu_inst_pe_1_5_2_n91,
         npu_inst_pe_1_5_2_n90, npu_inst_pe_1_5_2_n89, npu_inst_pe_1_5_2_n88,
         npu_inst_pe_1_5_2_n87, npu_inst_pe_1_5_2_n86, npu_inst_pe_1_5_2_n85,
         npu_inst_pe_1_5_2_n84, npu_inst_pe_1_5_2_n83, npu_inst_pe_1_5_2_n82,
         npu_inst_pe_1_5_2_n81, npu_inst_pe_1_5_2_n80, npu_inst_pe_1_5_2_n79,
         npu_inst_pe_1_5_2_n78, npu_inst_pe_1_5_2_n77, npu_inst_pe_1_5_2_n76,
         npu_inst_pe_1_5_2_n75, npu_inst_pe_1_5_2_n74, npu_inst_pe_1_5_2_n73,
         npu_inst_pe_1_5_2_n72, npu_inst_pe_1_5_2_n71, npu_inst_pe_1_5_2_n70,
         npu_inst_pe_1_5_2_n69, npu_inst_pe_1_5_2_n68, npu_inst_pe_1_5_2_n67,
         npu_inst_pe_1_5_2_n66, npu_inst_pe_1_5_2_n65, npu_inst_pe_1_5_2_n64,
         npu_inst_pe_1_5_2_n63, npu_inst_pe_1_5_2_n62, npu_inst_pe_1_5_2_n61,
         npu_inst_pe_1_5_2_n60, npu_inst_pe_1_5_2_n59, npu_inst_pe_1_5_2_n58,
         npu_inst_pe_1_5_2_n57, npu_inst_pe_1_5_2_n56, npu_inst_pe_1_5_2_n55,
         npu_inst_pe_1_5_2_n54, npu_inst_pe_1_5_2_n53, npu_inst_pe_1_5_2_n52,
         npu_inst_pe_1_5_2_n51, npu_inst_pe_1_5_2_n50, npu_inst_pe_1_5_2_n49,
         npu_inst_pe_1_5_2_n48, npu_inst_pe_1_5_2_n47, npu_inst_pe_1_5_2_n46,
         npu_inst_pe_1_5_2_n45, npu_inst_pe_1_5_2_n44, npu_inst_pe_1_5_2_n43,
         npu_inst_pe_1_5_2_n42, npu_inst_pe_1_5_2_n41, npu_inst_pe_1_5_2_n40,
         npu_inst_pe_1_5_2_n39, npu_inst_pe_1_5_2_n38, npu_inst_pe_1_5_2_n37,
         npu_inst_pe_1_5_2_n27, npu_inst_pe_1_5_2_n26,
         npu_inst_pe_1_5_2_net3333, npu_inst_pe_1_5_2_net3327,
         npu_inst_pe_1_5_2_N94, npu_inst_pe_1_5_2_N93, npu_inst_pe_1_5_2_N84,
         npu_inst_pe_1_5_2_N80, npu_inst_pe_1_5_2_N79, npu_inst_pe_1_5_2_N78,
         npu_inst_pe_1_5_2_N77, npu_inst_pe_1_5_2_N76, npu_inst_pe_1_5_2_N75,
         npu_inst_pe_1_5_2_N74, npu_inst_pe_1_5_2_N73, npu_inst_pe_1_5_2_N72,
         npu_inst_pe_1_5_2_N71, npu_inst_pe_1_5_2_N70, npu_inst_pe_1_5_2_N69,
         npu_inst_pe_1_5_2_N68, npu_inst_pe_1_5_2_N67, npu_inst_pe_1_5_2_N66,
         npu_inst_pe_1_5_2_N65, npu_inst_pe_1_5_2_int_q_acc_0_,
         npu_inst_pe_1_5_2_int_q_acc_1_, npu_inst_pe_1_5_2_int_q_acc_2_,
         npu_inst_pe_1_5_2_int_q_acc_3_, npu_inst_pe_1_5_2_int_q_acc_4_,
         npu_inst_pe_1_5_2_int_q_acc_5_, npu_inst_pe_1_5_2_int_q_acc_6_,
         npu_inst_pe_1_5_2_int_q_acc_7_, npu_inst_pe_1_5_2_int_data_0_,
         npu_inst_pe_1_5_2_int_data_1_, npu_inst_pe_1_5_2_int_q_weight_0_,
         npu_inst_pe_1_5_2_int_q_weight_1_,
         npu_inst_pe_1_5_2_int_q_reg_v_5__0_,
         npu_inst_pe_1_5_2_int_q_reg_v_5__1_,
         npu_inst_pe_1_5_2_int_q_reg_v_4__0_,
         npu_inst_pe_1_5_2_int_q_reg_v_4__1_,
         npu_inst_pe_1_5_2_int_q_reg_v_3__0_,
         npu_inst_pe_1_5_2_int_q_reg_v_3__1_,
         npu_inst_pe_1_5_2_int_q_reg_v_2__0_,
         npu_inst_pe_1_5_2_int_q_reg_v_2__1_,
         npu_inst_pe_1_5_2_int_q_reg_v_1__0_,
         npu_inst_pe_1_5_2_int_q_reg_v_1__1_,
         npu_inst_pe_1_5_2_int_q_reg_v_0__0_,
         npu_inst_pe_1_5_2_int_q_reg_v_0__1_,
         npu_inst_pe_1_5_2_int_q_reg_h_5__0_,
         npu_inst_pe_1_5_2_int_q_reg_h_5__1_,
         npu_inst_pe_1_5_2_int_q_reg_h_4__0_,
         npu_inst_pe_1_5_2_int_q_reg_h_4__1_,
         npu_inst_pe_1_5_2_int_q_reg_h_3__0_,
         npu_inst_pe_1_5_2_int_q_reg_h_3__1_,
         npu_inst_pe_1_5_2_int_q_reg_h_2__0_,
         npu_inst_pe_1_5_2_int_q_reg_h_2__1_,
         npu_inst_pe_1_5_2_int_q_reg_h_1__0_,
         npu_inst_pe_1_5_2_int_q_reg_h_1__1_,
         npu_inst_pe_1_5_2_int_q_reg_h_0__0_,
         npu_inst_pe_1_5_2_int_q_reg_h_0__1_, npu_inst_pe_1_5_3_n119,
         npu_inst_pe_1_5_3_n118, npu_inst_pe_1_5_3_n117,
         npu_inst_pe_1_5_3_n116, npu_inst_pe_1_5_3_n115,
         npu_inst_pe_1_5_3_n114, npu_inst_pe_1_5_3_n113,
         npu_inst_pe_1_5_3_n112, npu_inst_pe_1_5_3_n111,
         npu_inst_pe_1_5_3_n110, npu_inst_pe_1_5_3_n109,
         npu_inst_pe_1_5_3_n108, npu_inst_pe_1_5_3_n107,
         npu_inst_pe_1_5_3_n106, npu_inst_pe_1_5_3_n105,
         npu_inst_pe_1_5_3_n104, npu_inst_pe_1_5_3_n103,
         npu_inst_pe_1_5_3_n102, npu_inst_pe_1_5_3_n101,
         npu_inst_pe_1_5_3_n100, npu_inst_pe_1_5_3_n99, npu_inst_pe_1_5_3_n98,
         npu_inst_pe_1_5_3_n36, npu_inst_pe_1_5_3_n35, npu_inst_pe_1_5_3_n34,
         npu_inst_pe_1_5_3_n33, npu_inst_pe_1_5_3_n32, npu_inst_pe_1_5_3_n31,
         npu_inst_pe_1_5_3_n30, npu_inst_pe_1_5_3_n29, npu_inst_pe_1_5_3_n28,
         npu_inst_pe_1_5_3_n25, npu_inst_pe_1_5_3_n24, npu_inst_pe_1_5_3_n23,
         npu_inst_pe_1_5_3_n22, npu_inst_pe_1_5_3_n21, npu_inst_pe_1_5_3_n20,
         npu_inst_pe_1_5_3_n19, npu_inst_pe_1_5_3_n18, npu_inst_pe_1_5_3_n17,
         npu_inst_pe_1_5_3_n16, npu_inst_pe_1_5_3_n15, npu_inst_pe_1_5_3_n14,
         npu_inst_pe_1_5_3_n13, npu_inst_pe_1_5_3_n12, npu_inst_pe_1_5_3_n11,
         npu_inst_pe_1_5_3_n10, npu_inst_pe_1_5_3_n9, npu_inst_pe_1_5_3_n8,
         npu_inst_pe_1_5_3_n7, npu_inst_pe_1_5_3_n6, npu_inst_pe_1_5_3_n5,
         npu_inst_pe_1_5_3_n4, npu_inst_pe_1_5_3_n3, npu_inst_pe_1_5_3_n2,
         npu_inst_pe_1_5_3_n1, npu_inst_pe_1_5_3_sub_77_carry_7_,
         npu_inst_pe_1_5_3_sub_77_carry_6_, npu_inst_pe_1_5_3_sub_77_carry_5_,
         npu_inst_pe_1_5_3_sub_77_carry_4_, npu_inst_pe_1_5_3_sub_77_carry_3_,
         npu_inst_pe_1_5_3_sub_77_carry_2_, npu_inst_pe_1_5_3_sub_77_carry_1_,
         npu_inst_pe_1_5_3_add_79_carry_7_, npu_inst_pe_1_5_3_add_79_carry_6_,
         npu_inst_pe_1_5_3_add_79_carry_5_, npu_inst_pe_1_5_3_add_79_carry_4_,
         npu_inst_pe_1_5_3_add_79_carry_3_, npu_inst_pe_1_5_3_add_79_carry_2_,
         npu_inst_pe_1_5_3_add_79_carry_1_, npu_inst_pe_1_5_3_n97,
         npu_inst_pe_1_5_3_n96, npu_inst_pe_1_5_3_n95, npu_inst_pe_1_5_3_n94,
         npu_inst_pe_1_5_3_n93, npu_inst_pe_1_5_3_n92, npu_inst_pe_1_5_3_n91,
         npu_inst_pe_1_5_3_n90, npu_inst_pe_1_5_3_n89, npu_inst_pe_1_5_3_n88,
         npu_inst_pe_1_5_3_n87, npu_inst_pe_1_5_3_n86, npu_inst_pe_1_5_3_n85,
         npu_inst_pe_1_5_3_n84, npu_inst_pe_1_5_3_n83, npu_inst_pe_1_5_3_n82,
         npu_inst_pe_1_5_3_n81, npu_inst_pe_1_5_3_n80, npu_inst_pe_1_5_3_n79,
         npu_inst_pe_1_5_3_n78, npu_inst_pe_1_5_3_n77, npu_inst_pe_1_5_3_n76,
         npu_inst_pe_1_5_3_n75, npu_inst_pe_1_5_3_n74, npu_inst_pe_1_5_3_n73,
         npu_inst_pe_1_5_3_n72, npu_inst_pe_1_5_3_n71, npu_inst_pe_1_5_3_n70,
         npu_inst_pe_1_5_3_n69, npu_inst_pe_1_5_3_n68, npu_inst_pe_1_5_3_n67,
         npu_inst_pe_1_5_3_n66, npu_inst_pe_1_5_3_n65, npu_inst_pe_1_5_3_n64,
         npu_inst_pe_1_5_3_n63, npu_inst_pe_1_5_3_n62, npu_inst_pe_1_5_3_n61,
         npu_inst_pe_1_5_3_n60, npu_inst_pe_1_5_3_n59, npu_inst_pe_1_5_3_n58,
         npu_inst_pe_1_5_3_n57, npu_inst_pe_1_5_3_n56, npu_inst_pe_1_5_3_n55,
         npu_inst_pe_1_5_3_n54, npu_inst_pe_1_5_3_n53, npu_inst_pe_1_5_3_n52,
         npu_inst_pe_1_5_3_n51, npu_inst_pe_1_5_3_n50, npu_inst_pe_1_5_3_n49,
         npu_inst_pe_1_5_3_n48, npu_inst_pe_1_5_3_n47, npu_inst_pe_1_5_3_n46,
         npu_inst_pe_1_5_3_n45, npu_inst_pe_1_5_3_n44, npu_inst_pe_1_5_3_n43,
         npu_inst_pe_1_5_3_n42, npu_inst_pe_1_5_3_n41, npu_inst_pe_1_5_3_n40,
         npu_inst_pe_1_5_3_n39, npu_inst_pe_1_5_3_n38, npu_inst_pe_1_5_3_n37,
         npu_inst_pe_1_5_3_n27, npu_inst_pe_1_5_3_n26,
         npu_inst_pe_1_5_3_net3310, npu_inst_pe_1_5_3_net3304,
         npu_inst_pe_1_5_3_N94, npu_inst_pe_1_5_3_N93, npu_inst_pe_1_5_3_N84,
         npu_inst_pe_1_5_3_N80, npu_inst_pe_1_5_3_N79, npu_inst_pe_1_5_3_N78,
         npu_inst_pe_1_5_3_N77, npu_inst_pe_1_5_3_N76, npu_inst_pe_1_5_3_N75,
         npu_inst_pe_1_5_3_N74, npu_inst_pe_1_5_3_N73, npu_inst_pe_1_5_3_N72,
         npu_inst_pe_1_5_3_N71, npu_inst_pe_1_5_3_N70, npu_inst_pe_1_5_3_N69,
         npu_inst_pe_1_5_3_N68, npu_inst_pe_1_5_3_N67, npu_inst_pe_1_5_3_N66,
         npu_inst_pe_1_5_3_N65, npu_inst_pe_1_5_3_int_q_acc_0_,
         npu_inst_pe_1_5_3_int_q_acc_1_, npu_inst_pe_1_5_3_int_q_acc_2_,
         npu_inst_pe_1_5_3_int_q_acc_3_, npu_inst_pe_1_5_3_int_q_acc_4_,
         npu_inst_pe_1_5_3_int_q_acc_5_, npu_inst_pe_1_5_3_int_q_acc_6_,
         npu_inst_pe_1_5_3_int_q_acc_7_, npu_inst_pe_1_5_3_int_data_0_,
         npu_inst_pe_1_5_3_int_data_1_, npu_inst_pe_1_5_3_int_q_weight_0_,
         npu_inst_pe_1_5_3_int_q_weight_1_,
         npu_inst_pe_1_5_3_int_q_reg_v_5__0_,
         npu_inst_pe_1_5_3_int_q_reg_v_5__1_,
         npu_inst_pe_1_5_3_int_q_reg_v_4__0_,
         npu_inst_pe_1_5_3_int_q_reg_v_4__1_,
         npu_inst_pe_1_5_3_int_q_reg_v_3__0_,
         npu_inst_pe_1_5_3_int_q_reg_v_3__1_,
         npu_inst_pe_1_5_3_int_q_reg_v_2__0_,
         npu_inst_pe_1_5_3_int_q_reg_v_2__1_,
         npu_inst_pe_1_5_3_int_q_reg_v_1__0_,
         npu_inst_pe_1_5_3_int_q_reg_v_1__1_,
         npu_inst_pe_1_5_3_int_q_reg_v_0__0_,
         npu_inst_pe_1_5_3_int_q_reg_v_0__1_,
         npu_inst_pe_1_5_3_int_q_reg_h_5__0_,
         npu_inst_pe_1_5_3_int_q_reg_h_5__1_,
         npu_inst_pe_1_5_3_int_q_reg_h_4__0_,
         npu_inst_pe_1_5_3_int_q_reg_h_4__1_,
         npu_inst_pe_1_5_3_int_q_reg_h_3__0_,
         npu_inst_pe_1_5_3_int_q_reg_h_3__1_,
         npu_inst_pe_1_5_3_int_q_reg_h_2__0_,
         npu_inst_pe_1_5_3_int_q_reg_h_2__1_,
         npu_inst_pe_1_5_3_int_q_reg_h_1__0_,
         npu_inst_pe_1_5_3_int_q_reg_h_1__1_,
         npu_inst_pe_1_5_3_int_q_reg_h_0__0_,
         npu_inst_pe_1_5_3_int_q_reg_h_0__1_, npu_inst_pe_1_5_4_n119,
         npu_inst_pe_1_5_4_n118, npu_inst_pe_1_5_4_n117,
         npu_inst_pe_1_5_4_n116, npu_inst_pe_1_5_4_n115,
         npu_inst_pe_1_5_4_n114, npu_inst_pe_1_5_4_n113,
         npu_inst_pe_1_5_4_n112, npu_inst_pe_1_5_4_n111,
         npu_inst_pe_1_5_4_n110, npu_inst_pe_1_5_4_n109,
         npu_inst_pe_1_5_4_n108, npu_inst_pe_1_5_4_n107,
         npu_inst_pe_1_5_4_n106, npu_inst_pe_1_5_4_n105,
         npu_inst_pe_1_5_4_n104, npu_inst_pe_1_5_4_n103,
         npu_inst_pe_1_5_4_n102, npu_inst_pe_1_5_4_n101,
         npu_inst_pe_1_5_4_n100, npu_inst_pe_1_5_4_n99, npu_inst_pe_1_5_4_n98,
         npu_inst_pe_1_5_4_n36, npu_inst_pe_1_5_4_n35, npu_inst_pe_1_5_4_n34,
         npu_inst_pe_1_5_4_n33, npu_inst_pe_1_5_4_n32, npu_inst_pe_1_5_4_n31,
         npu_inst_pe_1_5_4_n30, npu_inst_pe_1_5_4_n29, npu_inst_pe_1_5_4_n28,
         npu_inst_pe_1_5_4_n25, npu_inst_pe_1_5_4_n24, npu_inst_pe_1_5_4_n23,
         npu_inst_pe_1_5_4_n22, npu_inst_pe_1_5_4_n21, npu_inst_pe_1_5_4_n20,
         npu_inst_pe_1_5_4_n19, npu_inst_pe_1_5_4_n18, npu_inst_pe_1_5_4_n17,
         npu_inst_pe_1_5_4_n16, npu_inst_pe_1_5_4_n15, npu_inst_pe_1_5_4_n14,
         npu_inst_pe_1_5_4_n13, npu_inst_pe_1_5_4_n12, npu_inst_pe_1_5_4_n11,
         npu_inst_pe_1_5_4_n10, npu_inst_pe_1_5_4_n9, npu_inst_pe_1_5_4_n8,
         npu_inst_pe_1_5_4_n7, npu_inst_pe_1_5_4_n6, npu_inst_pe_1_5_4_n5,
         npu_inst_pe_1_5_4_n4, npu_inst_pe_1_5_4_n3, npu_inst_pe_1_5_4_n2,
         npu_inst_pe_1_5_4_n1, npu_inst_pe_1_5_4_sub_77_carry_7_,
         npu_inst_pe_1_5_4_sub_77_carry_6_, npu_inst_pe_1_5_4_sub_77_carry_5_,
         npu_inst_pe_1_5_4_sub_77_carry_4_, npu_inst_pe_1_5_4_sub_77_carry_3_,
         npu_inst_pe_1_5_4_sub_77_carry_2_, npu_inst_pe_1_5_4_sub_77_carry_1_,
         npu_inst_pe_1_5_4_add_79_carry_7_, npu_inst_pe_1_5_4_add_79_carry_6_,
         npu_inst_pe_1_5_4_add_79_carry_5_, npu_inst_pe_1_5_4_add_79_carry_4_,
         npu_inst_pe_1_5_4_add_79_carry_3_, npu_inst_pe_1_5_4_add_79_carry_2_,
         npu_inst_pe_1_5_4_add_79_carry_1_, npu_inst_pe_1_5_4_n97,
         npu_inst_pe_1_5_4_n96, npu_inst_pe_1_5_4_n95, npu_inst_pe_1_5_4_n94,
         npu_inst_pe_1_5_4_n93, npu_inst_pe_1_5_4_n92, npu_inst_pe_1_5_4_n91,
         npu_inst_pe_1_5_4_n90, npu_inst_pe_1_5_4_n89, npu_inst_pe_1_5_4_n88,
         npu_inst_pe_1_5_4_n87, npu_inst_pe_1_5_4_n86, npu_inst_pe_1_5_4_n85,
         npu_inst_pe_1_5_4_n84, npu_inst_pe_1_5_4_n83, npu_inst_pe_1_5_4_n82,
         npu_inst_pe_1_5_4_n81, npu_inst_pe_1_5_4_n80, npu_inst_pe_1_5_4_n79,
         npu_inst_pe_1_5_4_n78, npu_inst_pe_1_5_4_n77, npu_inst_pe_1_5_4_n76,
         npu_inst_pe_1_5_4_n75, npu_inst_pe_1_5_4_n74, npu_inst_pe_1_5_4_n73,
         npu_inst_pe_1_5_4_n72, npu_inst_pe_1_5_4_n71, npu_inst_pe_1_5_4_n70,
         npu_inst_pe_1_5_4_n69, npu_inst_pe_1_5_4_n68, npu_inst_pe_1_5_4_n67,
         npu_inst_pe_1_5_4_n66, npu_inst_pe_1_5_4_n65, npu_inst_pe_1_5_4_n64,
         npu_inst_pe_1_5_4_n63, npu_inst_pe_1_5_4_n62, npu_inst_pe_1_5_4_n61,
         npu_inst_pe_1_5_4_n60, npu_inst_pe_1_5_4_n59, npu_inst_pe_1_5_4_n58,
         npu_inst_pe_1_5_4_n57, npu_inst_pe_1_5_4_n56, npu_inst_pe_1_5_4_n55,
         npu_inst_pe_1_5_4_n54, npu_inst_pe_1_5_4_n53, npu_inst_pe_1_5_4_n52,
         npu_inst_pe_1_5_4_n51, npu_inst_pe_1_5_4_n50, npu_inst_pe_1_5_4_n49,
         npu_inst_pe_1_5_4_n48, npu_inst_pe_1_5_4_n47, npu_inst_pe_1_5_4_n46,
         npu_inst_pe_1_5_4_n45, npu_inst_pe_1_5_4_n44, npu_inst_pe_1_5_4_n43,
         npu_inst_pe_1_5_4_n42, npu_inst_pe_1_5_4_n41, npu_inst_pe_1_5_4_n40,
         npu_inst_pe_1_5_4_n39, npu_inst_pe_1_5_4_n38, npu_inst_pe_1_5_4_n37,
         npu_inst_pe_1_5_4_n27, npu_inst_pe_1_5_4_n26,
         npu_inst_pe_1_5_4_net3287, npu_inst_pe_1_5_4_net3281,
         npu_inst_pe_1_5_4_N94, npu_inst_pe_1_5_4_N93, npu_inst_pe_1_5_4_N84,
         npu_inst_pe_1_5_4_N80, npu_inst_pe_1_5_4_N79, npu_inst_pe_1_5_4_N78,
         npu_inst_pe_1_5_4_N77, npu_inst_pe_1_5_4_N76, npu_inst_pe_1_5_4_N75,
         npu_inst_pe_1_5_4_N74, npu_inst_pe_1_5_4_N73, npu_inst_pe_1_5_4_N72,
         npu_inst_pe_1_5_4_N71, npu_inst_pe_1_5_4_N70, npu_inst_pe_1_5_4_N69,
         npu_inst_pe_1_5_4_N68, npu_inst_pe_1_5_4_N67, npu_inst_pe_1_5_4_N66,
         npu_inst_pe_1_5_4_N65, npu_inst_pe_1_5_4_int_q_acc_0_,
         npu_inst_pe_1_5_4_int_q_acc_1_, npu_inst_pe_1_5_4_int_q_acc_2_,
         npu_inst_pe_1_5_4_int_q_acc_3_, npu_inst_pe_1_5_4_int_q_acc_4_,
         npu_inst_pe_1_5_4_int_q_acc_5_, npu_inst_pe_1_5_4_int_q_acc_6_,
         npu_inst_pe_1_5_4_int_q_acc_7_, npu_inst_pe_1_5_4_int_data_0_,
         npu_inst_pe_1_5_4_int_data_1_, npu_inst_pe_1_5_4_int_q_weight_0_,
         npu_inst_pe_1_5_4_int_q_weight_1_,
         npu_inst_pe_1_5_4_int_q_reg_v_5__0_,
         npu_inst_pe_1_5_4_int_q_reg_v_5__1_,
         npu_inst_pe_1_5_4_int_q_reg_v_4__0_,
         npu_inst_pe_1_5_4_int_q_reg_v_4__1_,
         npu_inst_pe_1_5_4_int_q_reg_v_3__0_,
         npu_inst_pe_1_5_4_int_q_reg_v_3__1_,
         npu_inst_pe_1_5_4_int_q_reg_v_2__0_,
         npu_inst_pe_1_5_4_int_q_reg_v_2__1_,
         npu_inst_pe_1_5_4_int_q_reg_v_1__0_,
         npu_inst_pe_1_5_4_int_q_reg_v_1__1_,
         npu_inst_pe_1_5_4_int_q_reg_v_0__0_,
         npu_inst_pe_1_5_4_int_q_reg_v_0__1_,
         npu_inst_pe_1_5_4_int_q_reg_h_5__0_,
         npu_inst_pe_1_5_4_int_q_reg_h_5__1_,
         npu_inst_pe_1_5_4_int_q_reg_h_4__0_,
         npu_inst_pe_1_5_4_int_q_reg_h_4__1_,
         npu_inst_pe_1_5_4_int_q_reg_h_3__0_,
         npu_inst_pe_1_5_4_int_q_reg_h_3__1_,
         npu_inst_pe_1_5_4_int_q_reg_h_2__0_,
         npu_inst_pe_1_5_4_int_q_reg_h_2__1_,
         npu_inst_pe_1_5_4_int_q_reg_h_1__0_,
         npu_inst_pe_1_5_4_int_q_reg_h_1__1_,
         npu_inst_pe_1_5_4_int_q_reg_h_0__0_,
         npu_inst_pe_1_5_4_int_q_reg_h_0__1_, npu_inst_pe_1_5_5_n119,
         npu_inst_pe_1_5_5_n118, npu_inst_pe_1_5_5_n117,
         npu_inst_pe_1_5_5_n116, npu_inst_pe_1_5_5_n115,
         npu_inst_pe_1_5_5_n114, npu_inst_pe_1_5_5_n113,
         npu_inst_pe_1_5_5_n112, npu_inst_pe_1_5_5_n111,
         npu_inst_pe_1_5_5_n110, npu_inst_pe_1_5_5_n109,
         npu_inst_pe_1_5_5_n108, npu_inst_pe_1_5_5_n107,
         npu_inst_pe_1_5_5_n106, npu_inst_pe_1_5_5_n105,
         npu_inst_pe_1_5_5_n104, npu_inst_pe_1_5_5_n103,
         npu_inst_pe_1_5_5_n102, npu_inst_pe_1_5_5_n101,
         npu_inst_pe_1_5_5_n100, npu_inst_pe_1_5_5_n99, npu_inst_pe_1_5_5_n98,
         npu_inst_pe_1_5_5_n36, npu_inst_pe_1_5_5_n35, npu_inst_pe_1_5_5_n34,
         npu_inst_pe_1_5_5_n33, npu_inst_pe_1_5_5_n32, npu_inst_pe_1_5_5_n31,
         npu_inst_pe_1_5_5_n30, npu_inst_pe_1_5_5_n29, npu_inst_pe_1_5_5_n28,
         npu_inst_pe_1_5_5_n25, npu_inst_pe_1_5_5_n24, npu_inst_pe_1_5_5_n23,
         npu_inst_pe_1_5_5_n22, npu_inst_pe_1_5_5_n21, npu_inst_pe_1_5_5_n20,
         npu_inst_pe_1_5_5_n19, npu_inst_pe_1_5_5_n18, npu_inst_pe_1_5_5_n17,
         npu_inst_pe_1_5_5_n16, npu_inst_pe_1_5_5_n15, npu_inst_pe_1_5_5_n14,
         npu_inst_pe_1_5_5_n13, npu_inst_pe_1_5_5_n12, npu_inst_pe_1_5_5_n11,
         npu_inst_pe_1_5_5_n10, npu_inst_pe_1_5_5_n9, npu_inst_pe_1_5_5_n8,
         npu_inst_pe_1_5_5_n7, npu_inst_pe_1_5_5_n6, npu_inst_pe_1_5_5_n5,
         npu_inst_pe_1_5_5_n4, npu_inst_pe_1_5_5_n3, npu_inst_pe_1_5_5_n2,
         npu_inst_pe_1_5_5_n1, npu_inst_pe_1_5_5_sub_77_carry_7_,
         npu_inst_pe_1_5_5_sub_77_carry_6_, npu_inst_pe_1_5_5_sub_77_carry_5_,
         npu_inst_pe_1_5_5_sub_77_carry_4_, npu_inst_pe_1_5_5_sub_77_carry_3_,
         npu_inst_pe_1_5_5_sub_77_carry_2_, npu_inst_pe_1_5_5_sub_77_carry_1_,
         npu_inst_pe_1_5_5_add_79_carry_7_, npu_inst_pe_1_5_5_add_79_carry_6_,
         npu_inst_pe_1_5_5_add_79_carry_5_, npu_inst_pe_1_5_5_add_79_carry_4_,
         npu_inst_pe_1_5_5_add_79_carry_3_, npu_inst_pe_1_5_5_add_79_carry_2_,
         npu_inst_pe_1_5_5_add_79_carry_1_, npu_inst_pe_1_5_5_n97,
         npu_inst_pe_1_5_5_n96, npu_inst_pe_1_5_5_n95, npu_inst_pe_1_5_5_n94,
         npu_inst_pe_1_5_5_n93, npu_inst_pe_1_5_5_n92, npu_inst_pe_1_5_5_n91,
         npu_inst_pe_1_5_5_n90, npu_inst_pe_1_5_5_n89, npu_inst_pe_1_5_5_n88,
         npu_inst_pe_1_5_5_n87, npu_inst_pe_1_5_5_n86, npu_inst_pe_1_5_5_n85,
         npu_inst_pe_1_5_5_n84, npu_inst_pe_1_5_5_n83, npu_inst_pe_1_5_5_n82,
         npu_inst_pe_1_5_5_n81, npu_inst_pe_1_5_5_n80, npu_inst_pe_1_5_5_n79,
         npu_inst_pe_1_5_5_n78, npu_inst_pe_1_5_5_n77, npu_inst_pe_1_5_5_n76,
         npu_inst_pe_1_5_5_n75, npu_inst_pe_1_5_5_n74, npu_inst_pe_1_5_5_n73,
         npu_inst_pe_1_5_5_n72, npu_inst_pe_1_5_5_n71, npu_inst_pe_1_5_5_n70,
         npu_inst_pe_1_5_5_n69, npu_inst_pe_1_5_5_n68, npu_inst_pe_1_5_5_n67,
         npu_inst_pe_1_5_5_n66, npu_inst_pe_1_5_5_n65, npu_inst_pe_1_5_5_n64,
         npu_inst_pe_1_5_5_n63, npu_inst_pe_1_5_5_n62, npu_inst_pe_1_5_5_n61,
         npu_inst_pe_1_5_5_n60, npu_inst_pe_1_5_5_n59, npu_inst_pe_1_5_5_n58,
         npu_inst_pe_1_5_5_n57, npu_inst_pe_1_5_5_n56, npu_inst_pe_1_5_5_n55,
         npu_inst_pe_1_5_5_n54, npu_inst_pe_1_5_5_n53, npu_inst_pe_1_5_5_n52,
         npu_inst_pe_1_5_5_n51, npu_inst_pe_1_5_5_n50, npu_inst_pe_1_5_5_n49,
         npu_inst_pe_1_5_5_n48, npu_inst_pe_1_5_5_n47, npu_inst_pe_1_5_5_n46,
         npu_inst_pe_1_5_5_n45, npu_inst_pe_1_5_5_n44, npu_inst_pe_1_5_5_n43,
         npu_inst_pe_1_5_5_n42, npu_inst_pe_1_5_5_n41, npu_inst_pe_1_5_5_n40,
         npu_inst_pe_1_5_5_n39, npu_inst_pe_1_5_5_n38, npu_inst_pe_1_5_5_n37,
         npu_inst_pe_1_5_5_n27, npu_inst_pe_1_5_5_n26,
         npu_inst_pe_1_5_5_net3264, npu_inst_pe_1_5_5_net3258,
         npu_inst_pe_1_5_5_N94, npu_inst_pe_1_5_5_N93, npu_inst_pe_1_5_5_N84,
         npu_inst_pe_1_5_5_N80, npu_inst_pe_1_5_5_N79, npu_inst_pe_1_5_5_N78,
         npu_inst_pe_1_5_5_N77, npu_inst_pe_1_5_5_N76, npu_inst_pe_1_5_5_N75,
         npu_inst_pe_1_5_5_N74, npu_inst_pe_1_5_5_N73, npu_inst_pe_1_5_5_N72,
         npu_inst_pe_1_5_5_N71, npu_inst_pe_1_5_5_N70, npu_inst_pe_1_5_5_N69,
         npu_inst_pe_1_5_5_N68, npu_inst_pe_1_5_5_N67, npu_inst_pe_1_5_5_N66,
         npu_inst_pe_1_5_5_N65, npu_inst_pe_1_5_5_int_q_acc_0_,
         npu_inst_pe_1_5_5_int_q_acc_1_, npu_inst_pe_1_5_5_int_q_acc_2_,
         npu_inst_pe_1_5_5_int_q_acc_3_, npu_inst_pe_1_5_5_int_q_acc_4_,
         npu_inst_pe_1_5_5_int_q_acc_5_, npu_inst_pe_1_5_5_int_q_acc_6_,
         npu_inst_pe_1_5_5_int_q_acc_7_, npu_inst_pe_1_5_5_int_data_0_,
         npu_inst_pe_1_5_5_int_data_1_, npu_inst_pe_1_5_5_int_q_weight_0_,
         npu_inst_pe_1_5_5_int_q_weight_1_,
         npu_inst_pe_1_5_5_int_q_reg_v_5__0_,
         npu_inst_pe_1_5_5_int_q_reg_v_5__1_,
         npu_inst_pe_1_5_5_int_q_reg_v_4__0_,
         npu_inst_pe_1_5_5_int_q_reg_v_4__1_,
         npu_inst_pe_1_5_5_int_q_reg_v_3__0_,
         npu_inst_pe_1_5_5_int_q_reg_v_3__1_,
         npu_inst_pe_1_5_5_int_q_reg_v_2__0_,
         npu_inst_pe_1_5_5_int_q_reg_v_2__1_,
         npu_inst_pe_1_5_5_int_q_reg_v_1__0_,
         npu_inst_pe_1_5_5_int_q_reg_v_1__1_,
         npu_inst_pe_1_5_5_int_q_reg_v_0__0_,
         npu_inst_pe_1_5_5_int_q_reg_v_0__1_,
         npu_inst_pe_1_5_5_int_q_reg_h_5__0_,
         npu_inst_pe_1_5_5_int_q_reg_h_5__1_,
         npu_inst_pe_1_5_5_int_q_reg_h_4__0_,
         npu_inst_pe_1_5_5_int_q_reg_h_4__1_,
         npu_inst_pe_1_5_5_int_q_reg_h_3__0_,
         npu_inst_pe_1_5_5_int_q_reg_h_3__1_,
         npu_inst_pe_1_5_5_int_q_reg_h_2__0_,
         npu_inst_pe_1_5_5_int_q_reg_h_2__1_,
         npu_inst_pe_1_5_5_int_q_reg_h_1__0_,
         npu_inst_pe_1_5_5_int_q_reg_h_1__1_,
         npu_inst_pe_1_5_5_int_q_reg_h_0__0_,
         npu_inst_pe_1_5_5_int_q_reg_h_0__1_, npu_inst_pe_1_5_6_n119,
         npu_inst_pe_1_5_6_n118, npu_inst_pe_1_5_6_n117,
         npu_inst_pe_1_5_6_n116, npu_inst_pe_1_5_6_n115,
         npu_inst_pe_1_5_6_n114, npu_inst_pe_1_5_6_n113,
         npu_inst_pe_1_5_6_n112, npu_inst_pe_1_5_6_n111,
         npu_inst_pe_1_5_6_n110, npu_inst_pe_1_5_6_n109,
         npu_inst_pe_1_5_6_n108, npu_inst_pe_1_5_6_n107,
         npu_inst_pe_1_5_6_n106, npu_inst_pe_1_5_6_n105,
         npu_inst_pe_1_5_6_n104, npu_inst_pe_1_5_6_n103,
         npu_inst_pe_1_5_6_n102, npu_inst_pe_1_5_6_n101,
         npu_inst_pe_1_5_6_n100, npu_inst_pe_1_5_6_n99, npu_inst_pe_1_5_6_n98,
         npu_inst_pe_1_5_6_n36, npu_inst_pe_1_5_6_n35, npu_inst_pe_1_5_6_n34,
         npu_inst_pe_1_5_6_n33, npu_inst_pe_1_5_6_n32, npu_inst_pe_1_5_6_n31,
         npu_inst_pe_1_5_6_n30, npu_inst_pe_1_5_6_n29, npu_inst_pe_1_5_6_n28,
         npu_inst_pe_1_5_6_n25, npu_inst_pe_1_5_6_n24, npu_inst_pe_1_5_6_n23,
         npu_inst_pe_1_5_6_n22, npu_inst_pe_1_5_6_n21, npu_inst_pe_1_5_6_n20,
         npu_inst_pe_1_5_6_n19, npu_inst_pe_1_5_6_n18, npu_inst_pe_1_5_6_n17,
         npu_inst_pe_1_5_6_n16, npu_inst_pe_1_5_6_n15, npu_inst_pe_1_5_6_n14,
         npu_inst_pe_1_5_6_n13, npu_inst_pe_1_5_6_n12, npu_inst_pe_1_5_6_n11,
         npu_inst_pe_1_5_6_n10, npu_inst_pe_1_5_6_n9, npu_inst_pe_1_5_6_n8,
         npu_inst_pe_1_5_6_n7, npu_inst_pe_1_5_6_n6, npu_inst_pe_1_5_6_n5,
         npu_inst_pe_1_5_6_n4, npu_inst_pe_1_5_6_n3, npu_inst_pe_1_5_6_n2,
         npu_inst_pe_1_5_6_n1, npu_inst_pe_1_5_6_sub_77_carry_7_,
         npu_inst_pe_1_5_6_sub_77_carry_6_, npu_inst_pe_1_5_6_sub_77_carry_5_,
         npu_inst_pe_1_5_6_sub_77_carry_4_, npu_inst_pe_1_5_6_sub_77_carry_3_,
         npu_inst_pe_1_5_6_sub_77_carry_2_, npu_inst_pe_1_5_6_sub_77_carry_1_,
         npu_inst_pe_1_5_6_add_79_carry_7_, npu_inst_pe_1_5_6_add_79_carry_6_,
         npu_inst_pe_1_5_6_add_79_carry_5_, npu_inst_pe_1_5_6_add_79_carry_4_,
         npu_inst_pe_1_5_6_add_79_carry_3_, npu_inst_pe_1_5_6_add_79_carry_2_,
         npu_inst_pe_1_5_6_add_79_carry_1_, npu_inst_pe_1_5_6_n97,
         npu_inst_pe_1_5_6_n96, npu_inst_pe_1_5_6_n95, npu_inst_pe_1_5_6_n94,
         npu_inst_pe_1_5_6_n93, npu_inst_pe_1_5_6_n92, npu_inst_pe_1_5_6_n91,
         npu_inst_pe_1_5_6_n90, npu_inst_pe_1_5_6_n89, npu_inst_pe_1_5_6_n88,
         npu_inst_pe_1_5_6_n87, npu_inst_pe_1_5_6_n86, npu_inst_pe_1_5_6_n85,
         npu_inst_pe_1_5_6_n84, npu_inst_pe_1_5_6_n83, npu_inst_pe_1_5_6_n82,
         npu_inst_pe_1_5_6_n81, npu_inst_pe_1_5_6_n80, npu_inst_pe_1_5_6_n79,
         npu_inst_pe_1_5_6_n78, npu_inst_pe_1_5_6_n77, npu_inst_pe_1_5_6_n76,
         npu_inst_pe_1_5_6_n75, npu_inst_pe_1_5_6_n74, npu_inst_pe_1_5_6_n73,
         npu_inst_pe_1_5_6_n72, npu_inst_pe_1_5_6_n71, npu_inst_pe_1_5_6_n70,
         npu_inst_pe_1_5_6_n69, npu_inst_pe_1_5_6_n68, npu_inst_pe_1_5_6_n67,
         npu_inst_pe_1_5_6_n66, npu_inst_pe_1_5_6_n65, npu_inst_pe_1_5_6_n64,
         npu_inst_pe_1_5_6_n63, npu_inst_pe_1_5_6_n62, npu_inst_pe_1_5_6_n61,
         npu_inst_pe_1_5_6_n60, npu_inst_pe_1_5_6_n59, npu_inst_pe_1_5_6_n58,
         npu_inst_pe_1_5_6_n57, npu_inst_pe_1_5_6_n56, npu_inst_pe_1_5_6_n55,
         npu_inst_pe_1_5_6_n54, npu_inst_pe_1_5_6_n53, npu_inst_pe_1_5_6_n52,
         npu_inst_pe_1_5_6_n51, npu_inst_pe_1_5_6_n50, npu_inst_pe_1_5_6_n49,
         npu_inst_pe_1_5_6_n48, npu_inst_pe_1_5_6_n47, npu_inst_pe_1_5_6_n46,
         npu_inst_pe_1_5_6_n45, npu_inst_pe_1_5_6_n44, npu_inst_pe_1_5_6_n43,
         npu_inst_pe_1_5_6_n42, npu_inst_pe_1_5_6_n41, npu_inst_pe_1_5_6_n40,
         npu_inst_pe_1_5_6_n39, npu_inst_pe_1_5_6_n38, npu_inst_pe_1_5_6_n37,
         npu_inst_pe_1_5_6_n27, npu_inst_pe_1_5_6_n26,
         npu_inst_pe_1_5_6_net3241, npu_inst_pe_1_5_6_net3235,
         npu_inst_pe_1_5_6_N94, npu_inst_pe_1_5_6_N93, npu_inst_pe_1_5_6_N84,
         npu_inst_pe_1_5_6_N80, npu_inst_pe_1_5_6_N79, npu_inst_pe_1_5_6_N78,
         npu_inst_pe_1_5_6_N77, npu_inst_pe_1_5_6_N76, npu_inst_pe_1_5_6_N75,
         npu_inst_pe_1_5_6_N74, npu_inst_pe_1_5_6_N73, npu_inst_pe_1_5_6_N72,
         npu_inst_pe_1_5_6_N71, npu_inst_pe_1_5_6_N70, npu_inst_pe_1_5_6_N69,
         npu_inst_pe_1_5_6_N68, npu_inst_pe_1_5_6_N67, npu_inst_pe_1_5_6_N66,
         npu_inst_pe_1_5_6_N65, npu_inst_pe_1_5_6_int_q_acc_0_,
         npu_inst_pe_1_5_6_int_q_acc_1_, npu_inst_pe_1_5_6_int_q_acc_2_,
         npu_inst_pe_1_5_6_int_q_acc_3_, npu_inst_pe_1_5_6_int_q_acc_4_,
         npu_inst_pe_1_5_6_int_q_acc_5_, npu_inst_pe_1_5_6_int_q_acc_6_,
         npu_inst_pe_1_5_6_int_q_acc_7_, npu_inst_pe_1_5_6_int_data_0_,
         npu_inst_pe_1_5_6_int_data_1_, npu_inst_pe_1_5_6_int_q_weight_0_,
         npu_inst_pe_1_5_6_int_q_weight_1_,
         npu_inst_pe_1_5_6_int_q_reg_v_5__0_,
         npu_inst_pe_1_5_6_int_q_reg_v_5__1_,
         npu_inst_pe_1_5_6_int_q_reg_v_4__0_,
         npu_inst_pe_1_5_6_int_q_reg_v_4__1_,
         npu_inst_pe_1_5_6_int_q_reg_v_3__0_,
         npu_inst_pe_1_5_6_int_q_reg_v_3__1_,
         npu_inst_pe_1_5_6_int_q_reg_v_2__0_,
         npu_inst_pe_1_5_6_int_q_reg_v_2__1_,
         npu_inst_pe_1_5_6_int_q_reg_v_1__0_,
         npu_inst_pe_1_5_6_int_q_reg_v_1__1_,
         npu_inst_pe_1_5_6_int_q_reg_v_0__0_,
         npu_inst_pe_1_5_6_int_q_reg_v_0__1_,
         npu_inst_pe_1_5_6_int_q_reg_h_5__0_,
         npu_inst_pe_1_5_6_int_q_reg_h_5__1_,
         npu_inst_pe_1_5_6_int_q_reg_h_4__0_,
         npu_inst_pe_1_5_6_int_q_reg_h_4__1_,
         npu_inst_pe_1_5_6_int_q_reg_h_3__0_,
         npu_inst_pe_1_5_6_int_q_reg_h_3__1_,
         npu_inst_pe_1_5_6_int_q_reg_h_2__0_,
         npu_inst_pe_1_5_6_int_q_reg_h_2__1_,
         npu_inst_pe_1_5_6_int_q_reg_h_1__0_,
         npu_inst_pe_1_5_6_int_q_reg_h_1__1_,
         npu_inst_pe_1_5_6_int_q_reg_h_0__0_,
         npu_inst_pe_1_5_6_int_q_reg_h_0__1_, npu_inst_pe_1_5_7_n119,
         npu_inst_pe_1_5_7_n118, npu_inst_pe_1_5_7_n117,
         npu_inst_pe_1_5_7_n116, npu_inst_pe_1_5_7_n115,
         npu_inst_pe_1_5_7_n114, npu_inst_pe_1_5_7_n113,
         npu_inst_pe_1_5_7_n112, npu_inst_pe_1_5_7_n111,
         npu_inst_pe_1_5_7_n110, npu_inst_pe_1_5_7_n109,
         npu_inst_pe_1_5_7_n108, npu_inst_pe_1_5_7_n107,
         npu_inst_pe_1_5_7_n106, npu_inst_pe_1_5_7_n105,
         npu_inst_pe_1_5_7_n104, npu_inst_pe_1_5_7_n103,
         npu_inst_pe_1_5_7_n102, npu_inst_pe_1_5_7_n101,
         npu_inst_pe_1_5_7_n100, npu_inst_pe_1_5_7_n99, npu_inst_pe_1_5_7_n98,
         npu_inst_pe_1_5_7_n36, npu_inst_pe_1_5_7_n35, npu_inst_pe_1_5_7_n34,
         npu_inst_pe_1_5_7_n33, npu_inst_pe_1_5_7_n32, npu_inst_pe_1_5_7_n31,
         npu_inst_pe_1_5_7_n30, npu_inst_pe_1_5_7_n29, npu_inst_pe_1_5_7_n28,
         npu_inst_pe_1_5_7_n25, npu_inst_pe_1_5_7_n24, npu_inst_pe_1_5_7_n23,
         npu_inst_pe_1_5_7_n22, npu_inst_pe_1_5_7_n21, npu_inst_pe_1_5_7_n20,
         npu_inst_pe_1_5_7_n19, npu_inst_pe_1_5_7_n18, npu_inst_pe_1_5_7_n17,
         npu_inst_pe_1_5_7_n16, npu_inst_pe_1_5_7_n15, npu_inst_pe_1_5_7_n14,
         npu_inst_pe_1_5_7_n13, npu_inst_pe_1_5_7_n12, npu_inst_pe_1_5_7_n11,
         npu_inst_pe_1_5_7_n10, npu_inst_pe_1_5_7_n9, npu_inst_pe_1_5_7_n8,
         npu_inst_pe_1_5_7_n7, npu_inst_pe_1_5_7_n6, npu_inst_pe_1_5_7_n5,
         npu_inst_pe_1_5_7_n4, npu_inst_pe_1_5_7_n3, npu_inst_pe_1_5_7_n2,
         npu_inst_pe_1_5_7_n1, npu_inst_pe_1_5_7_sub_77_carry_7_,
         npu_inst_pe_1_5_7_sub_77_carry_6_, npu_inst_pe_1_5_7_sub_77_carry_5_,
         npu_inst_pe_1_5_7_sub_77_carry_4_, npu_inst_pe_1_5_7_sub_77_carry_3_,
         npu_inst_pe_1_5_7_sub_77_carry_2_, npu_inst_pe_1_5_7_sub_77_carry_1_,
         npu_inst_pe_1_5_7_add_79_carry_7_, npu_inst_pe_1_5_7_add_79_carry_6_,
         npu_inst_pe_1_5_7_add_79_carry_5_, npu_inst_pe_1_5_7_add_79_carry_4_,
         npu_inst_pe_1_5_7_add_79_carry_3_, npu_inst_pe_1_5_7_add_79_carry_2_,
         npu_inst_pe_1_5_7_add_79_carry_1_, npu_inst_pe_1_5_7_n97,
         npu_inst_pe_1_5_7_n96, npu_inst_pe_1_5_7_n95, npu_inst_pe_1_5_7_n94,
         npu_inst_pe_1_5_7_n93, npu_inst_pe_1_5_7_n92, npu_inst_pe_1_5_7_n91,
         npu_inst_pe_1_5_7_n90, npu_inst_pe_1_5_7_n89, npu_inst_pe_1_5_7_n88,
         npu_inst_pe_1_5_7_n87, npu_inst_pe_1_5_7_n86, npu_inst_pe_1_5_7_n85,
         npu_inst_pe_1_5_7_n84, npu_inst_pe_1_5_7_n83, npu_inst_pe_1_5_7_n82,
         npu_inst_pe_1_5_7_n81, npu_inst_pe_1_5_7_n80, npu_inst_pe_1_5_7_n79,
         npu_inst_pe_1_5_7_n78, npu_inst_pe_1_5_7_n77, npu_inst_pe_1_5_7_n76,
         npu_inst_pe_1_5_7_n75, npu_inst_pe_1_5_7_n74, npu_inst_pe_1_5_7_n73,
         npu_inst_pe_1_5_7_n72, npu_inst_pe_1_5_7_n71, npu_inst_pe_1_5_7_n70,
         npu_inst_pe_1_5_7_n69, npu_inst_pe_1_5_7_n68, npu_inst_pe_1_5_7_n67,
         npu_inst_pe_1_5_7_n66, npu_inst_pe_1_5_7_n65, npu_inst_pe_1_5_7_n64,
         npu_inst_pe_1_5_7_n63, npu_inst_pe_1_5_7_n62, npu_inst_pe_1_5_7_n61,
         npu_inst_pe_1_5_7_n60, npu_inst_pe_1_5_7_n59, npu_inst_pe_1_5_7_n58,
         npu_inst_pe_1_5_7_n57, npu_inst_pe_1_5_7_n56, npu_inst_pe_1_5_7_n55,
         npu_inst_pe_1_5_7_n54, npu_inst_pe_1_5_7_n53, npu_inst_pe_1_5_7_n52,
         npu_inst_pe_1_5_7_n51, npu_inst_pe_1_5_7_n50, npu_inst_pe_1_5_7_n49,
         npu_inst_pe_1_5_7_n48, npu_inst_pe_1_5_7_n47, npu_inst_pe_1_5_7_n46,
         npu_inst_pe_1_5_7_n45, npu_inst_pe_1_5_7_n44, npu_inst_pe_1_5_7_n43,
         npu_inst_pe_1_5_7_n42, npu_inst_pe_1_5_7_n41, npu_inst_pe_1_5_7_n40,
         npu_inst_pe_1_5_7_n39, npu_inst_pe_1_5_7_n38, npu_inst_pe_1_5_7_n37,
         npu_inst_pe_1_5_7_n27, npu_inst_pe_1_5_7_n26,
         npu_inst_pe_1_5_7_net3218, npu_inst_pe_1_5_7_net3212,
         npu_inst_pe_1_5_7_N94, npu_inst_pe_1_5_7_N93, npu_inst_pe_1_5_7_N84,
         npu_inst_pe_1_5_7_N80, npu_inst_pe_1_5_7_N79, npu_inst_pe_1_5_7_N78,
         npu_inst_pe_1_5_7_N77, npu_inst_pe_1_5_7_N76, npu_inst_pe_1_5_7_N75,
         npu_inst_pe_1_5_7_N74, npu_inst_pe_1_5_7_N73, npu_inst_pe_1_5_7_N72,
         npu_inst_pe_1_5_7_N71, npu_inst_pe_1_5_7_N70, npu_inst_pe_1_5_7_N69,
         npu_inst_pe_1_5_7_N68, npu_inst_pe_1_5_7_N67, npu_inst_pe_1_5_7_N66,
         npu_inst_pe_1_5_7_N65, npu_inst_pe_1_5_7_int_q_acc_0_,
         npu_inst_pe_1_5_7_int_q_acc_1_, npu_inst_pe_1_5_7_int_q_acc_2_,
         npu_inst_pe_1_5_7_int_q_acc_3_, npu_inst_pe_1_5_7_int_q_acc_4_,
         npu_inst_pe_1_5_7_int_q_acc_5_, npu_inst_pe_1_5_7_int_q_acc_6_,
         npu_inst_pe_1_5_7_int_q_acc_7_, npu_inst_pe_1_5_7_int_data_0_,
         npu_inst_pe_1_5_7_int_data_1_, npu_inst_pe_1_5_7_int_q_weight_0_,
         npu_inst_pe_1_5_7_int_q_weight_1_,
         npu_inst_pe_1_5_7_int_q_reg_v_5__0_,
         npu_inst_pe_1_5_7_int_q_reg_v_5__1_,
         npu_inst_pe_1_5_7_int_q_reg_v_4__0_,
         npu_inst_pe_1_5_7_int_q_reg_v_4__1_,
         npu_inst_pe_1_5_7_int_q_reg_v_3__0_,
         npu_inst_pe_1_5_7_int_q_reg_v_3__1_,
         npu_inst_pe_1_5_7_int_q_reg_v_2__0_,
         npu_inst_pe_1_5_7_int_q_reg_v_2__1_,
         npu_inst_pe_1_5_7_int_q_reg_v_1__0_,
         npu_inst_pe_1_5_7_int_q_reg_v_1__1_,
         npu_inst_pe_1_5_7_int_q_reg_v_0__0_,
         npu_inst_pe_1_5_7_int_q_reg_v_0__1_,
         npu_inst_pe_1_5_7_int_q_reg_h_5__0_,
         npu_inst_pe_1_5_7_int_q_reg_h_5__1_,
         npu_inst_pe_1_5_7_int_q_reg_h_4__0_,
         npu_inst_pe_1_5_7_int_q_reg_h_4__1_,
         npu_inst_pe_1_5_7_int_q_reg_h_3__0_,
         npu_inst_pe_1_5_7_int_q_reg_h_3__1_,
         npu_inst_pe_1_5_7_int_q_reg_h_2__0_,
         npu_inst_pe_1_5_7_int_q_reg_h_2__1_,
         npu_inst_pe_1_5_7_int_q_reg_h_1__0_,
         npu_inst_pe_1_5_7_int_q_reg_h_1__1_,
         npu_inst_pe_1_5_7_int_q_reg_h_0__0_,
         npu_inst_pe_1_5_7_int_q_reg_h_0__1_, npu_inst_pe_1_6_0_n119,
         npu_inst_pe_1_6_0_n118, npu_inst_pe_1_6_0_n117,
         npu_inst_pe_1_6_0_n116, npu_inst_pe_1_6_0_n115,
         npu_inst_pe_1_6_0_n114, npu_inst_pe_1_6_0_n113,
         npu_inst_pe_1_6_0_n112, npu_inst_pe_1_6_0_n111,
         npu_inst_pe_1_6_0_n110, npu_inst_pe_1_6_0_n109,
         npu_inst_pe_1_6_0_n108, npu_inst_pe_1_6_0_n107,
         npu_inst_pe_1_6_0_n106, npu_inst_pe_1_6_0_n105,
         npu_inst_pe_1_6_0_n104, npu_inst_pe_1_6_0_n103,
         npu_inst_pe_1_6_0_n102, npu_inst_pe_1_6_0_n101,
         npu_inst_pe_1_6_0_n100, npu_inst_pe_1_6_0_n99, npu_inst_pe_1_6_0_n98,
         npu_inst_pe_1_6_0_n36, npu_inst_pe_1_6_0_n35, npu_inst_pe_1_6_0_n34,
         npu_inst_pe_1_6_0_n33, npu_inst_pe_1_6_0_n32, npu_inst_pe_1_6_0_n31,
         npu_inst_pe_1_6_0_n30, npu_inst_pe_1_6_0_n29, npu_inst_pe_1_6_0_n28,
         npu_inst_pe_1_6_0_n25, npu_inst_pe_1_6_0_n24, npu_inst_pe_1_6_0_n23,
         npu_inst_pe_1_6_0_n22, npu_inst_pe_1_6_0_n21, npu_inst_pe_1_6_0_n20,
         npu_inst_pe_1_6_0_n19, npu_inst_pe_1_6_0_n18, npu_inst_pe_1_6_0_n17,
         npu_inst_pe_1_6_0_n16, npu_inst_pe_1_6_0_n15, npu_inst_pe_1_6_0_n14,
         npu_inst_pe_1_6_0_n13, npu_inst_pe_1_6_0_n12, npu_inst_pe_1_6_0_n11,
         npu_inst_pe_1_6_0_n10, npu_inst_pe_1_6_0_n9, npu_inst_pe_1_6_0_n8,
         npu_inst_pe_1_6_0_n7, npu_inst_pe_1_6_0_n6, npu_inst_pe_1_6_0_n5,
         npu_inst_pe_1_6_0_n4, npu_inst_pe_1_6_0_n3, npu_inst_pe_1_6_0_n2,
         npu_inst_pe_1_6_0_n1, npu_inst_pe_1_6_0_sub_77_carry_7_,
         npu_inst_pe_1_6_0_sub_77_carry_6_, npu_inst_pe_1_6_0_sub_77_carry_5_,
         npu_inst_pe_1_6_0_sub_77_carry_4_, npu_inst_pe_1_6_0_sub_77_carry_3_,
         npu_inst_pe_1_6_0_sub_77_carry_2_, npu_inst_pe_1_6_0_sub_77_carry_1_,
         npu_inst_pe_1_6_0_add_79_carry_7_, npu_inst_pe_1_6_0_add_79_carry_6_,
         npu_inst_pe_1_6_0_add_79_carry_5_, npu_inst_pe_1_6_0_add_79_carry_4_,
         npu_inst_pe_1_6_0_add_79_carry_3_, npu_inst_pe_1_6_0_add_79_carry_2_,
         npu_inst_pe_1_6_0_add_79_carry_1_, npu_inst_pe_1_6_0_n97,
         npu_inst_pe_1_6_0_n96, npu_inst_pe_1_6_0_n95, npu_inst_pe_1_6_0_n94,
         npu_inst_pe_1_6_0_n93, npu_inst_pe_1_6_0_n92, npu_inst_pe_1_6_0_n91,
         npu_inst_pe_1_6_0_n90, npu_inst_pe_1_6_0_n89, npu_inst_pe_1_6_0_n88,
         npu_inst_pe_1_6_0_n87, npu_inst_pe_1_6_0_n86, npu_inst_pe_1_6_0_n85,
         npu_inst_pe_1_6_0_n84, npu_inst_pe_1_6_0_n83, npu_inst_pe_1_6_0_n82,
         npu_inst_pe_1_6_0_n81, npu_inst_pe_1_6_0_n80, npu_inst_pe_1_6_0_n79,
         npu_inst_pe_1_6_0_n78, npu_inst_pe_1_6_0_n77, npu_inst_pe_1_6_0_n76,
         npu_inst_pe_1_6_0_n75, npu_inst_pe_1_6_0_n74, npu_inst_pe_1_6_0_n73,
         npu_inst_pe_1_6_0_n72, npu_inst_pe_1_6_0_n71, npu_inst_pe_1_6_0_n70,
         npu_inst_pe_1_6_0_n69, npu_inst_pe_1_6_0_n68, npu_inst_pe_1_6_0_n67,
         npu_inst_pe_1_6_0_n66, npu_inst_pe_1_6_0_n65, npu_inst_pe_1_6_0_n64,
         npu_inst_pe_1_6_0_n63, npu_inst_pe_1_6_0_n62, npu_inst_pe_1_6_0_n61,
         npu_inst_pe_1_6_0_n60, npu_inst_pe_1_6_0_n59, npu_inst_pe_1_6_0_n58,
         npu_inst_pe_1_6_0_n57, npu_inst_pe_1_6_0_n56, npu_inst_pe_1_6_0_n55,
         npu_inst_pe_1_6_0_n54, npu_inst_pe_1_6_0_n53, npu_inst_pe_1_6_0_n52,
         npu_inst_pe_1_6_0_n51, npu_inst_pe_1_6_0_n50, npu_inst_pe_1_6_0_n49,
         npu_inst_pe_1_6_0_n48, npu_inst_pe_1_6_0_n47, npu_inst_pe_1_6_0_n46,
         npu_inst_pe_1_6_0_n45, npu_inst_pe_1_6_0_n44, npu_inst_pe_1_6_0_n43,
         npu_inst_pe_1_6_0_n42, npu_inst_pe_1_6_0_n41, npu_inst_pe_1_6_0_n40,
         npu_inst_pe_1_6_0_n39, npu_inst_pe_1_6_0_n38, npu_inst_pe_1_6_0_n37,
         npu_inst_pe_1_6_0_n27, npu_inst_pe_1_6_0_n26,
         npu_inst_pe_1_6_0_net3195, npu_inst_pe_1_6_0_net3189,
         npu_inst_pe_1_6_0_N94, npu_inst_pe_1_6_0_N93, npu_inst_pe_1_6_0_N84,
         npu_inst_pe_1_6_0_N80, npu_inst_pe_1_6_0_N79, npu_inst_pe_1_6_0_N78,
         npu_inst_pe_1_6_0_N77, npu_inst_pe_1_6_0_N76, npu_inst_pe_1_6_0_N75,
         npu_inst_pe_1_6_0_N74, npu_inst_pe_1_6_0_N73, npu_inst_pe_1_6_0_N72,
         npu_inst_pe_1_6_0_N71, npu_inst_pe_1_6_0_N70, npu_inst_pe_1_6_0_N69,
         npu_inst_pe_1_6_0_N68, npu_inst_pe_1_6_0_N67, npu_inst_pe_1_6_0_N66,
         npu_inst_pe_1_6_0_N65, npu_inst_pe_1_6_0_int_q_acc_0_,
         npu_inst_pe_1_6_0_int_q_acc_1_, npu_inst_pe_1_6_0_int_q_acc_2_,
         npu_inst_pe_1_6_0_int_q_acc_3_, npu_inst_pe_1_6_0_int_q_acc_4_,
         npu_inst_pe_1_6_0_int_q_acc_5_, npu_inst_pe_1_6_0_int_q_acc_6_,
         npu_inst_pe_1_6_0_int_q_acc_7_, npu_inst_pe_1_6_0_int_data_0_,
         npu_inst_pe_1_6_0_int_data_1_, npu_inst_pe_1_6_0_int_q_weight_0_,
         npu_inst_pe_1_6_0_int_q_weight_1_,
         npu_inst_pe_1_6_0_int_q_reg_v_5__0_,
         npu_inst_pe_1_6_0_int_q_reg_v_5__1_,
         npu_inst_pe_1_6_0_int_q_reg_v_4__0_,
         npu_inst_pe_1_6_0_int_q_reg_v_4__1_,
         npu_inst_pe_1_6_0_int_q_reg_v_3__0_,
         npu_inst_pe_1_6_0_int_q_reg_v_3__1_,
         npu_inst_pe_1_6_0_int_q_reg_v_2__0_,
         npu_inst_pe_1_6_0_int_q_reg_v_2__1_,
         npu_inst_pe_1_6_0_int_q_reg_v_1__0_,
         npu_inst_pe_1_6_0_int_q_reg_v_1__1_,
         npu_inst_pe_1_6_0_int_q_reg_v_0__0_,
         npu_inst_pe_1_6_0_int_q_reg_v_0__1_,
         npu_inst_pe_1_6_0_int_q_reg_h_5__0_,
         npu_inst_pe_1_6_0_int_q_reg_h_5__1_,
         npu_inst_pe_1_6_0_int_q_reg_h_4__0_,
         npu_inst_pe_1_6_0_int_q_reg_h_4__1_,
         npu_inst_pe_1_6_0_int_q_reg_h_3__0_,
         npu_inst_pe_1_6_0_int_q_reg_h_3__1_,
         npu_inst_pe_1_6_0_int_q_reg_h_2__0_,
         npu_inst_pe_1_6_0_int_q_reg_h_2__1_,
         npu_inst_pe_1_6_0_int_q_reg_h_1__0_,
         npu_inst_pe_1_6_0_int_q_reg_h_1__1_,
         npu_inst_pe_1_6_0_int_q_reg_h_0__0_,
         npu_inst_pe_1_6_0_int_q_reg_h_0__1_, npu_inst_pe_1_6_0_o_data_h_0_,
         npu_inst_pe_1_6_0_o_data_h_1_, npu_inst_pe_1_6_1_n119,
         npu_inst_pe_1_6_1_n118, npu_inst_pe_1_6_1_n117,
         npu_inst_pe_1_6_1_n116, npu_inst_pe_1_6_1_n115,
         npu_inst_pe_1_6_1_n114, npu_inst_pe_1_6_1_n113,
         npu_inst_pe_1_6_1_n112, npu_inst_pe_1_6_1_n111,
         npu_inst_pe_1_6_1_n110, npu_inst_pe_1_6_1_n109,
         npu_inst_pe_1_6_1_n108, npu_inst_pe_1_6_1_n107,
         npu_inst_pe_1_6_1_n106, npu_inst_pe_1_6_1_n105,
         npu_inst_pe_1_6_1_n104, npu_inst_pe_1_6_1_n103,
         npu_inst_pe_1_6_1_n102, npu_inst_pe_1_6_1_n101,
         npu_inst_pe_1_6_1_n100, npu_inst_pe_1_6_1_n99, npu_inst_pe_1_6_1_n98,
         npu_inst_pe_1_6_1_n36, npu_inst_pe_1_6_1_n35, npu_inst_pe_1_6_1_n34,
         npu_inst_pe_1_6_1_n33, npu_inst_pe_1_6_1_n32, npu_inst_pe_1_6_1_n31,
         npu_inst_pe_1_6_1_n30, npu_inst_pe_1_6_1_n29, npu_inst_pe_1_6_1_n28,
         npu_inst_pe_1_6_1_n25, npu_inst_pe_1_6_1_n24, npu_inst_pe_1_6_1_n23,
         npu_inst_pe_1_6_1_n22, npu_inst_pe_1_6_1_n21, npu_inst_pe_1_6_1_n20,
         npu_inst_pe_1_6_1_n19, npu_inst_pe_1_6_1_n18, npu_inst_pe_1_6_1_n17,
         npu_inst_pe_1_6_1_n16, npu_inst_pe_1_6_1_n15, npu_inst_pe_1_6_1_n14,
         npu_inst_pe_1_6_1_n13, npu_inst_pe_1_6_1_n12, npu_inst_pe_1_6_1_n11,
         npu_inst_pe_1_6_1_n10, npu_inst_pe_1_6_1_n9, npu_inst_pe_1_6_1_n8,
         npu_inst_pe_1_6_1_n7, npu_inst_pe_1_6_1_n6, npu_inst_pe_1_6_1_n5,
         npu_inst_pe_1_6_1_n4, npu_inst_pe_1_6_1_n3, npu_inst_pe_1_6_1_n2,
         npu_inst_pe_1_6_1_n1, npu_inst_pe_1_6_1_sub_77_carry_7_,
         npu_inst_pe_1_6_1_sub_77_carry_6_, npu_inst_pe_1_6_1_sub_77_carry_5_,
         npu_inst_pe_1_6_1_sub_77_carry_4_, npu_inst_pe_1_6_1_sub_77_carry_3_,
         npu_inst_pe_1_6_1_sub_77_carry_2_, npu_inst_pe_1_6_1_sub_77_carry_1_,
         npu_inst_pe_1_6_1_add_79_carry_7_, npu_inst_pe_1_6_1_add_79_carry_6_,
         npu_inst_pe_1_6_1_add_79_carry_5_, npu_inst_pe_1_6_1_add_79_carry_4_,
         npu_inst_pe_1_6_1_add_79_carry_3_, npu_inst_pe_1_6_1_add_79_carry_2_,
         npu_inst_pe_1_6_1_add_79_carry_1_, npu_inst_pe_1_6_1_n97,
         npu_inst_pe_1_6_1_n96, npu_inst_pe_1_6_1_n95, npu_inst_pe_1_6_1_n94,
         npu_inst_pe_1_6_1_n93, npu_inst_pe_1_6_1_n92, npu_inst_pe_1_6_1_n91,
         npu_inst_pe_1_6_1_n90, npu_inst_pe_1_6_1_n89, npu_inst_pe_1_6_1_n88,
         npu_inst_pe_1_6_1_n87, npu_inst_pe_1_6_1_n86, npu_inst_pe_1_6_1_n85,
         npu_inst_pe_1_6_1_n84, npu_inst_pe_1_6_1_n83, npu_inst_pe_1_6_1_n82,
         npu_inst_pe_1_6_1_n81, npu_inst_pe_1_6_1_n80, npu_inst_pe_1_6_1_n79,
         npu_inst_pe_1_6_1_n78, npu_inst_pe_1_6_1_n77, npu_inst_pe_1_6_1_n76,
         npu_inst_pe_1_6_1_n75, npu_inst_pe_1_6_1_n74, npu_inst_pe_1_6_1_n73,
         npu_inst_pe_1_6_1_n72, npu_inst_pe_1_6_1_n71, npu_inst_pe_1_6_1_n70,
         npu_inst_pe_1_6_1_n69, npu_inst_pe_1_6_1_n68, npu_inst_pe_1_6_1_n67,
         npu_inst_pe_1_6_1_n66, npu_inst_pe_1_6_1_n65, npu_inst_pe_1_6_1_n64,
         npu_inst_pe_1_6_1_n63, npu_inst_pe_1_6_1_n62, npu_inst_pe_1_6_1_n61,
         npu_inst_pe_1_6_1_n60, npu_inst_pe_1_6_1_n59, npu_inst_pe_1_6_1_n58,
         npu_inst_pe_1_6_1_n57, npu_inst_pe_1_6_1_n56, npu_inst_pe_1_6_1_n55,
         npu_inst_pe_1_6_1_n54, npu_inst_pe_1_6_1_n53, npu_inst_pe_1_6_1_n52,
         npu_inst_pe_1_6_1_n51, npu_inst_pe_1_6_1_n50, npu_inst_pe_1_6_1_n49,
         npu_inst_pe_1_6_1_n48, npu_inst_pe_1_6_1_n47, npu_inst_pe_1_6_1_n46,
         npu_inst_pe_1_6_1_n45, npu_inst_pe_1_6_1_n44, npu_inst_pe_1_6_1_n43,
         npu_inst_pe_1_6_1_n42, npu_inst_pe_1_6_1_n41, npu_inst_pe_1_6_1_n40,
         npu_inst_pe_1_6_1_n39, npu_inst_pe_1_6_1_n38, npu_inst_pe_1_6_1_n37,
         npu_inst_pe_1_6_1_n27, npu_inst_pe_1_6_1_n26,
         npu_inst_pe_1_6_1_net3172, npu_inst_pe_1_6_1_net3166,
         npu_inst_pe_1_6_1_N94, npu_inst_pe_1_6_1_N93, npu_inst_pe_1_6_1_N84,
         npu_inst_pe_1_6_1_N80, npu_inst_pe_1_6_1_N79, npu_inst_pe_1_6_1_N78,
         npu_inst_pe_1_6_1_N77, npu_inst_pe_1_6_1_N76, npu_inst_pe_1_6_1_N75,
         npu_inst_pe_1_6_1_N74, npu_inst_pe_1_6_1_N73, npu_inst_pe_1_6_1_N72,
         npu_inst_pe_1_6_1_N71, npu_inst_pe_1_6_1_N70, npu_inst_pe_1_6_1_N69,
         npu_inst_pe_1_6_1_N68, npu_inst_pe_1_6_1_N67, npu_inst_pe_1_6_1_N66,
         npu_inst_pe_1_6_1_N65, npu_inst_pe_1_6_1_int_q_acc_0_,
         npu_inst_pe_1_6_1_int_q_acc_1_, npu_inst_pe_1_6_1_int_q_acc_2_,
         npu_inst_pe_1_6_1_int_q_acc_3_, npu_inst_pe_1_6_1_int_q_acc_4_,
         npu_inst_pe_1_6_1_int_q_acc_5_, npu_inst_pe_1_6_1_int_q_acc_6_,
         npu_inst_pe_1_6_1_int_q_acc_7_, npu_inst_pe_1_6_1_int_data_0_,
         npu_inst_pe_1_6_1_int_data_1_, npu_inst_pe_1_6_1_int_q_weight_0_,
         npu_inst_pe_1_6_1_int_q_weight_1_,
         npu_inst_pe_1_6_1_int_q_reg_v_5__0_,
         npu_inst_pe_1_6_1_int_q_reg_v_5__1_,
         npu_inst_pe_1_6_1_int_q_reg_v_4__0_,
         npu_inst_pe_1_6_1_int_q_reg_v_4__1_,
         npu_inst_pe_1_6_1_int_q_reg_v_3__0_,
         npu_inst_pe_1_6_1_int_q_reg_v_3__1_,
         npu_inst_pe_1_6_1_int_q_reg_v_2__0_,
         npu_inst_pe_1_6_1_int_q_reg_v_2__1_,
         npu_inst_pe_1_6_1_int_q_reg_v_1__0_,
         npu_inst_pe_1_6_1_int_q_reg_v_1__1_,
         npu_inst_pe_1_6_1_int_q_reg_v_0__0_,
         npu_inst_pe_1_6_1_int_q_reg_v_0__1_,
         npu_inst_pe_1_6_1_int_q_reg_h_5__0_,
         npu_inst_pe_1_6_1_int_q_reg_h_5__1_,
         npu_inst_pe_1_6_1_int_q_reg_h_4__0_,
         npu_inst_pe_1_6_1_int_q_reg_h_4__1_,
         npu_inst_pe_1_6_1_int_q_reg_h_3__0_,
         npu_inst_pe_1_6_1_int_q_reg_h_3__1_,
         npu_inst_pe_1_6_1_int_q_reg_h_2__0_,
         npu_inst_pe_1_6_1_int_q_reg_h_2__1_,
         npu_inst_pe_1_6_1_int_q_reg_h_1__0_,
         npu_inst_pe_1_6_1_int_q_reg_h_1__1_,
         npu_inst_pe_1_6_1_int_q_reg_h_0__0_,
         npu_inst_pe_1_6_1_int_q_reg_h_0__1_, npu_inst_pe_1_6_2_n119,
         npu_inst_pe_1_6_2_n118, npu_inst_pe_1_6_2_n117,
         npu_inst_pe_1_6_2_n116, npu_inst_pe_1_6_2_n115,
         npu_inst_pe_1_6_2_n114, npu_inst_pe_1_6_2_n113,
         npu_inst_pe_1_6_2_n112, npu_inst_pe_1_6_2_n111,
         npu_inst_pe_1_6_2_n110, npu_inst_pe_1_6_2_n109,
         npu_inst_pe_1_6_2_n108, npu_inst_pe_1_6_2_n107,
         npu_inst_pe_1_6_2_n106, npu_inst_pe_1_6_2_n105,
         npu_inst_pe_1_6_2_n104, npu_inst_pe_1_6_2_n103,
         npu_inst_pe_1_6_2_n102, npu_inst_pe_1_6_2_n101,
         npu_inst_pe_1_6_2_n100, npu_inst_pe_1_6_2_n99, npu_inst_pe_1_6_2_n98,
         npu_inst_pe_1_6_2_n36, npu_inst_pe_1_6_2_n35, npu_inst_pe_1_6_2_n34,
         npu_inst_pe_1_6_2_n33, npu_inst_pe_1_6_2_n32, npu_inst_pe_1_6_2_n31,
         npu_inst_pe_1_6_2_n30, npu_inst_pe_1_6_2_n29, npu_inst_pe_1_6_2_n28,
         npu_inst_pe_1_6_2_n25, npu_inst_pe_1_6_2_n24, npu_inst_pe_1_6_2_n23,
         npu_inst_pe_1_6_2_n22, npu_inst_pe_1_6_2_n21, npu_inst_pe_1_6_2_n20,
         npu_inst_pe_1_6_2_n19, npu_inst_pe_1_6_2_n18, npu_inst_pe_1_6_2_n17,
         npu_inst_pe_1_6_2_n16, npu_inst_pe_1_6_2_n15, npu_inst_pe_1_6_2_n14,
         npu_inst_pe_1_6_2_n13, npu_inst_pe_1_6_2_n12, npu_inst_pe_1_6_2_n11,
         npu_inst_pe_1_6_2_n10, npu_inst_pe_1_6_2_n9, npu_inst_pe_1_6_2_n8,
         npu_inst_pe_1_6_2_n7, npu_inst_pe_1_6_2_n6, npu_inst_pe_1_6_2_n5,
         npu_inst_pe_1_6_2_n4, npu_inst_pe_1_6_2_n3, npu_inst_pe_1_6_2_n2,
         npu_inst_pe_1_6_2_n1, npu_inst_pe_1_6_2_sub_77_carry_7_,
         npu_inst_pe_1_6_2_sub_77_carry_6_, npu_inst_pe_1_6_2_sub_77_carry_5_,
         npu_inst_pe_1_6_2_sub_77_carry_4_, npu_inst_pe_1_6_2_sub_77_carry_3_,
         npu_inst_pe_1_6_2_sub_77_carry_2_, npu_inst_pe_1_6_2_sub_77_carry_1_,
         npu_inst_pe_1_6_2_add_79_carry_7_, npu_inst_pe_1_6_2_add_79_carry_6_,
         npu_inst_pe_1_6_2_add_79_carry_5_, npu_inst_pe_1_6_2_add_79_carry_4_,
         npu_inst_pe_1_6_2_add_79_carry_3_, npu_inst_pe_1_6_2_add_79_carry_2_,
         npu_inst_pe_1_6_2_add_79_carry_1_, npu_inst_pe_1_6_2_n97,
         npu_inst_pe_1_6_2_n96, npu_inst_pe_1_6_2_n95, npu_inst_pe_1_6_2_n94,
         npu_inst_pe_1_6_2_n93, npu_inst_pe_1_6_2_n92, npu_inst_pe_1_6_2_n91,
         npu_inst_pe_1_6_2_n90, npu_inst_pe_1_6_2_n89, npu_inst_pe_1_6_2_n88,
         npu_inst_pe_1_6_2_n87, npu_inst_pe_1_6_2_n86, npu_inst_pe_1_6_2_n85,
         npu_inst_pe_1_6_2_n84, npu_inst_pe_1_6_2_n83, npu_inst_pe_1_6_2_n82,
         npu_inst_pe_1_6_2_n81, npu_inst_pe_1_6_2_n80, npu_inst_pe_1_6_2_n79,
         npu_inst_pe_1_6_2_n78, npu_inst_pe_1_6_2_n77, npu_inst_pe_1_6_2_n76,
         npu_inst_pe_1_6_2_n75, npu_inst_pe_1_6_2_n74, npu_inst_pe_1_6_2_n73,
         npu_inst_pe_1_6_2_n72, npu_inst_pe_1_6_2_n71, npu_inst_pe_1_6_2_n70,
         npu_inst_pe_1_6_2_n69, npu_inst_pe_1_6_2_n68, npu_inst_pe_1_6_2_n67,
         npu_inst_pe_1_6_2_n66, npu_inst_pe_1_6_2_n65, npu_inst_pe_1_6_2_n64,
         npu_inst_pe_1_6_2_n63, npu_inst_pe_1_6_2_n62, npu_inst_pe_1_6_2_n61,
         npu_inst_pe_1_6_2_n60, npu_inst_pe_1_6_2_n59, npu_inst_pe_1_6_2_n58,
         npu_inst_pe_1_6_2_n57, npu_inst_pe_1_6_2_n56, npu_inst_pe_1_6_2_n55,
         npu_inst_pe_1_6_2_n54, npu_inst_pe_1_6_2_n53, npu_inst_pe_1_6_2_n52,
         npu_inst_pe_1_6_2_n51, npu_inst_pe_1_6_2_n50, npu_inst_pe_1_6_2_n49,
         npu_inst_pe_1_6_2_n48, npu_inst_pe_1_6_2_n47, npu_inst_pe_1_6_2_n46,
         npu_inst_pe_1_6_2_n45, npu_inst_pe_1_6_2_n44, npu_inst_pe_1_6_2_n43,
         npu_inst_pe_1_6_2_n42, npu_inst_pe_1_6_2_n41, npu_inst_pe_1_6_2_n40,
         npu_inst_pe_1_6_2_n39, npu_inst_pe_1_6_2_n38, npu_inst_pe_1_6_2_n37,
         npu_inst_pe_1_6_2_n27, npu_inst_pe_1_6_2_n26,
         npu_inst_pe_1_6_2_net3149, npu_inst_pe_1_6_2_net3143,
         npu_inst_pe_1_6_2_N94, npu_inst_pe_1_6_2_N93, npu_inst_pe_1_6_2_N84,
         npu_inst_pe_1_6_2_N80, npu_inst_pe_1_6_2_N79, npu_inst_pe_1_6_2_N78,
         npu_inst_pe_1_6_2_N77, npu_inst_pe_1_6_2_N76, npu_inst_pe_1_6_2_N75,
         npu_inst_pe_1_6_2_N74, npu_inst_pe_1_6_2_N73, npu_inst_pe_1_6_2_N72,
         npu_inst_pe_1_6_2_N71, npu_inst_pe_1_6_2_N70, npu_inst_pe_1_6_2_N69,
         npu_inst_pe_1_6_2_N68, npu_inst_pe_1_6_2_N67, npu_inst_pe_1_6_2_N66,
         npu_inst_pe_1_6_2_N65, npu_inst_pe_1_6_2_int_q_acc_0_,
         npu_inst_pe_1_6_2_int_q_acc_1_, npu_inst_pe_1_6_2_int_q_acc_2_,
         npu_inst_pe_1_6_2_int_q_acc_3_, npu_inst_pe_1_6_2_int_q_acc_4_,
         npu_inst_pe_1_6_2_int_q_acc_5_, npu_inst_pe_1_6_2_int_q_acc_6_,
         npu_inst_pe_1_6_2_int_q_acc_7_, npu_inst_pe_1_6_2_int_data_0_,
         npu_inst_pe_1_6_2_int_data_1_, npu_inst_pe_1_6_2_int_q_weight_0_,
         npu_inst_pe_1_6_2_int_q_weight_1_,
         npu_inst_pe_1_6_2_int_q_reg_v_5__0_,
         npu_inst_pe_1_6_2_int_q_reg_v_5__1_,
         npu_inst_pe_1_6_2_int_q_reg_v_4__0_,
         npu_inst_pe_1_6_2_int_q_reg_v_4__1_,
         npu_inst_pe_1_6_2_int_q_reg_v_3__0_,
         npu_inst_pe_1_6_2_int_q_reg_v_3__1_,
         npu_inst_pe_1_6_2_int_q_reg_v_2__0_,
         npu_inst_pe_1_6_2_int_q_reg_v_2__1_,
         npu_inst_pe_1_6_2_int_q_reg_v_1__0_,
         npu_inst_pe_1_6_2_int_q_reg_v_1__1_,
         npu_inst_pe_1_6_2_int_q_reg_v_0__0_,
         npu_inst_pe_1_6_2_int_q_reg_v_0__1_,
         npu_inst_pe_1_6_2_int_q_reg_h_5__0_,
         npu_inst_pe_1_6_2_int_q_reg_h_5__1_,
         npu_inst_pe_1_6_2_int_q_reg_h_4__0_,
         npu_inst_pe_1_6_2_int_q_reg_h_4__1_,
         npu_inst_pe_1_6_2_int_q_reg_h_3__0_,
         npu_inst_pe_1_6_2_int_q_reg_h_3__1_,
         npu_inst_pe_1_6_2_int_q_reg_h_2__0_,
         npu_inst_pe_1_6_2_int_q_reg_h_2__1_,
         npu_inst_pe_1_6_2_int_q_reg_h_1__0_,
         npu_inst_pe_1_6_2_int_q_reg_h_1__1_,
         npu_inst_pe_1_6_2_int_q_reg_h_0__0_,
         npu_inst_pe_1_6_2_int_q_reg_h_0__1_, npu_inst_pe_1_6_3_n119,
         npu_inst_pe_1_6_3_n118, npu_inst_pe_1_6_3_n117,
         npu_inst_pe_1_6_3_n116, npu_inst_pe_1_6_3_n115,
         npu_inst_pe_1_6_3_n114, npu_inst_pe_1_6_3_n113,
         npu_inst_pe_1_6_3_n112, npu_inst_pe_1_6_3_n111,
         npu_inst_pe_1_6_3_n110, npu_inst_pe_1_6_3_n109,
         npu_inst_pe_1_6_3_n108, npu_inst_pe_1_6_3_n107,
         npu_inst_pe_1_6_3_n106, npu_inst_pe_1_6_3_n105,
         npu_inst_pe_1_6_3_n104, npu_inst_pe_1_6_3_n103,
         npu_inst_pe_1_6_3_n102, npu_inst_pe_1_6_3_n101,
         npu_inst_pe_1_6_3_n100, npu_inst_pe_1_6_3_n99, npu_inst_pe_1_6_3_n98,
         npu_inst_pe_1_6_3_n36, npu_inst_pe_1_6_3_n35, npu_inst_pe_1_6_3_n34,
         npu_inst_pe_1_6_3_n33, npu_inst_pe_1_6_3_n32, npu_inst_pe_1_6_3_n31,
         npu_inst_pe_1_6_3_n30, npu_inst_pe_1_6_3_n29, npu_inst_pe_1_6_3_n28,
         npu_inst_pe_1_6_3_n25, npu_inst_pe_1_6_3_n24, npu_inst_pe_1_6_3_n23,
         npu_inst_pe_1_6_3_n22, npu_inst_pe_1_6_3_n21, npu_inst_pe_1_6_3_n20,
         npu_inst_pe_1_6_3_n19, npu_inst_pe_1_6_3_n18, npu_inst_pe_1_6_3_n17,
         npu_inst_pe_1_6_3_n16, npu_inst_pe_1_6_3_n15, npu_inst_pe_1_6_3_n14,
         npu_inst_pe_1_6_3_n13, npu_inst_pe_1_6_3_n12, npu_inst_pe_1_6_3_n11,
         npu_inst_pe_1_6_3_n10, npu_inst_pe_1_6_3_n9, npu_inst_pe_1_6_3_n8,
         npu_inst_pe_1_6_3_n7, npu_inst_pe_1_6_3_n6, npu_inst_pe_1_6_3_n5,
         npu_inst_pe_1_6_3_n4, npu_inst_pe_1_6_3_n3, npu_inst_pe_1_6_3_n2,
         npu_inst_pe_1_6_3_n1, npu_inst_pe_1_6_3_sub_77_carry_7_,
         npu_inst_pe_1_6_3_sub_77_carry_6_, npu_inst_pe_1_6_3_sub_77_carry_5_,
         npu_inst_pe_1_6_3_sub_77_carry_4_, npu_inst_pe_1_6_3_sub_77_carry_3_,
         npu_inst_pe_1_6_3_sub_77_carry_2_, npu_inst_pe_1_6_3_sub_77_carry_1_,
         npu_inst_pe_1_6_3_add_79_carry_7_, npu_inst_pe_1_6_3_add_79_carry_6_,
         npu_inst_pe_1_6_3_add_79_carry_5_, npu_inst_pe_1_6_3_add_79_carry_4_,
         npu_inst_pe_1_6_3_add_79_carry_3_, npu_inst_pe_1_6_3_add_79_carry_2_,
         npu_inst_pe_1_6_3_add_79_carry_1_, npu_inst_pe_1_6_3_n97,
         npu_inst_pe_1_6_3_n96, npu_inst_pe_1_6_3_n95, npu_inst_pe_1_6_3_n94,
         npu_inst_pe_1_6_3_n93, npu_inst_pe_1_6_3_n92, npu_inst_pe_1_6_3_n91,
         npu_inst_pe_1_6_3_n90, npu_inst_pe_1_6_3_n89, npu_inst_pe_1_6_3_n88,
         npu_inst_pe_1_6_3_n87, npu_inst_pe_1_6_3_n86, npu_inst_pe_1_6_3_n85,
         npu_inst_pe_1_6_3_n84, npu_inst_pe_1_6_3_n83, npu_inst_pe_1_6_3_n82,
         npu_inst_pe_1_6_3_n81, npu_inst_pe_1_6_3_n80, npu_inst_pe_1_6_3_n79,
         npu_inst_pe_1_6_3_n78, npu_inst_pe_1_6_3_n77, npu_inst_pe_1_6_3_n76,
         npu_inst_pe_1_6_3_n75, npu_inst_pe_1_6_3_n74, npu_inst_pe_1_6_3_n73,
         npu_inst_pe_1_6_3_n72, npu_inst_pe_1_6_3_n71, npu_inst_pe_1_6_3_n70,
         npu_inst_pe_1_6_3_n69, npu_inst_pe_1_6_3_n68, npu_inst_pe_1_6_3_n67,
         npu_inst_pe_1_6_3_n66, npu_inst_pe_1_6_3_n65, npu_inst_pe_1_6_3_n64,
         npu_inst_pe_1_6_3_n63, npu_inst_pe_1_6_3_n62, npu_inst_pe_1_6_3_n61,
         npu_inst_pe_1_6_3_n60, npu_inst_pe_1_6_3_n59, npu_inst_pe_1_6_3_n58,
         npu_inst_pe_1_6_3_n57, npu_inst_pe_1_6_3_n56, npu_inst_pe_1_6_3_n55,
         npu_inst_pe_1_6_3_n54, npu_inst_pe_1_6_3_n53, npu_inst_pe_1_6_3_n52,
         npu_inst_pe_1_6_3_n51, npu_inst_pe_1_6_3_n50, npu_inst_pe_1_6_3_n49,
         npu_inst_pe_1_6_3_n48, npu_inst_pe_1_6_3_n47, npu_inst_pe_1_6_3_n46,
         npu_inst_pe_1_6_3_n45, npu_inst_pe_1_6_3_n44, npu_inst_pe_1_6_3_n43,
         npu_inst_pe_1_6_3_n42, npu_inst_pe_1_6_3_n41, npu_inst_pe_1_6_3_n40,
         npu_inst_pe_1_6_3_n39, npu_inst_pe_1_6_3_n38, npu_inst_pe_1_6_3_n37,
         npu_inst_pe_1_6_3_n27, npu_inst_pe_1_6_3_n26,
         npu_inst_pe_1_6_3_net3126, npu_inst_pe_1_6_3_net3120,
         npu_inst_pe_1_6_3_N94, npu_inst_pe_1_6_3_N93, npu_inst_pe_1_6_3_N84,
         npu_inst_pe_1_6_3_N80, npu_inst_pe_1_6_3_N79, npu_inst_pe_1_6_3_N78,
         npu_inst_pe_1_6_3_N77, npu_inst_pe_1_6_3_N76, npu_inst_pe_1_6_3_N75,
         npu_inst_pe_1_6_3_N74, npu_inst_pe_1_6_3_N73, npu_inst_pe_1_6_3_N72,
         npu_inst_pe_1_6_3_N71, npu_inst_pe_1_6_3_N70, npu_inst_pe_1_6_3_N69,
         npu_inst_pe_1_6_3_N68, npu_inst_pe_1_6_3_N67, npu_inst_pe_1_6_3_N66,
         npu_inst_pe_1_6_3_N65, npu_inst_pe_1_6_3_int_q_acc_0_,
         npu_inst_pe_1_6_3_int_q_acc_1_, npu_inst_pe_1_6_3_int_q_acc_2_,
         npu_inst_pe_1_6_3_int_q_acc_3_, npu_inst_pe_1_6_3_int_q_acc_4_,
         npu_inst_pe_1_6_3_int_q_acc_5_, npu_inst_pe_1_6_3_int_q_acc_6_,
         npu_inst_pe_1_6_3_int_q_acc_7_, npu_inst_pe_1_6_3_int_data_0_,
         npu_inst_pe_1_6_3_int_data_1_, npu_inst_pe_1_6_3_int_q_weight_0_,
         npu_inst_pe_1_6_3_int_q_weight_1_,
         npu_inst_pe_1_6_3_int_q_reg_v_5__0_,
         npu_inst_pe_1_6_3_int_q_reg_v_5__1_,
         npu_inst_pe_1_6_3_int_q_reg_v_4__0_,
         npu_inst_pe_1_6_3_int_q_reg_v_4__1_,
         npu_inst_pe_1_6_3_int_q_reg_v_3__0_,
         npu_inst_pe_1_6_3_int_q_reg_v_3__1_,
         npu_inst_pe_1_6_3_int_q_reg_v_2__0_,
         npu_inst_pe_1_6_3_int_q_reg_v_2__1_,
         npu_inst_pe_1_6_3_int_q_reg_v_1__0_,
         npu_inst_pe_1_6_3_int_q_reg_v_1__1_,
         npu_inst_pe_1_6_3_int_q_reg_v_0__0_,
         npu_inst_pe_1_6_3_int_q_reg_v_0__1_,
         npu_inst_pe_1_6_3_int_q_reg_h_5__0_,
         npu_inst_pe_1_6_3_int_q_reg_h_5__1_,
         npu_inst_pe_1_6_3_int_q_reg_h_4__0_,
         npu_inst_pe_1_6_3_int_q_reg_h_4__1_,
         npu_inst_pe_1_6_3_int_q_reg_h_3__0_,
         npu_inst_pe_1_6_3_int_q_reg_h_3__1_,
         npu_inst_pe_1_6_3_int_q_reg_h_2__0_,
         npu_inst_pe_1_6_3_int_q_reg_h_2__1_,
         npu_inst_pe_1_6_3_int_q_reg_h_1__0_,
         npu_inst_pe_1_6_3_int_q_reg_h_1__1_,
         npu_inst_pe_1_6_3_int_q_reg_h_0__0_,
         npu_inst_pe_1_6_3_int_q_reg_h_0__1_, npu_inst_pe_1_6_4_n118,
         npu_inst_pe_1_6_4_n117, npu_inst_pe_1_6_4_n116,
         npu_inst_pe_1_6_4_n115, npu_inst_pe_1_6_4_n114,
         npu_inst_pe_1_6_4_n113, npu_inst_pe_1_6_4_n112,
         npu_inst_pe_1_6_4_n111, npu_inst_pe_1_6_4_n110,
         npu_inst_pe_1_6_4_n109, npu_inst_pe_1_6_4_n108,
         npu_inst_pe_1_6_4_n107, npu_inst_pe_1_6_4_n106,
         npu_inst_pe_1_6_4_n105, npu_inst_pe_1_6_4_n104,
         npu_inst_pe_1_6_4_n103, npu_inst_pe_1_6_4_n102,
         npu_inst_pe_1_6_4_n101, npu_inst_pe_1_6_4_n100, npu_inst_pe_1_6_4_n99,
         npu_inst_pe_1_6_4_n98, npu_inst_pe_1_6_4_n36, npu_inst_pe_1_6_4_n35,
         npu_inst_pe_1_6_4_n34, npu_inst_pe_1_6_4_n33, npu_inst_pe_1_6_4_n32,
         npu_inst_pe_1_6_4_n31, npu_inst_pe_1_6_4_n30, npu_inst_pe_1_6_4_n29,
         npu_inst_pe_1_6_4_n28, npu_inst_pe_1_6_4_n25, npu_inst_pe_1_6_4_n24,
         npu_inst_pe_1_6_4_n23, npu_inst_pe_1_6_4_n22, npu_inst_pe_1_6_4_n21,
         npu_inst_pe_1_6_4_n20, npu_inst_pe_1_6_4_n19, npu_inst_pe_1_6_4_n18,
         npu_inst_pe_1_6_4_n17, npu_inst_pe_1_6_4_n16, npu_inst_pe_1_6_4_n15,
         npu_inst_pe_1_6_4_n14, npu_inst_pe_1_6_4_n13, npu_inst_pe_1_6_4_n12,
         npu_inst_pe_1_6_4_n11, npu_inst_pe_1_6_4_n10, npu_inst_pe_1_6_4_n9,
         npu_inst_pe_1_6_4_n8, npu_inst_pe_1_6_4_n7, npu_inst_pe_1_6_4_n6,
         npu_inst_pe_1_6_4_n5, npu_inst_pe_1_6_4_n4, npu_inst_pe_1_6_4_n3,
         npu_inst_pe_1_6_4_n2, npu_inst_pe_1_6_4_n1,
         npu_inst_pe_1_6_4_sub_77_carry_7_, npu_inst_pe_1_6_4_sub_77_carry_6_,
         npu_inst_pe_1_6_4_sub_77_carry_5_, npu_inst_pe_1_6_4_sub_77_carry_4_,
         npu_inst_pe_1_6_4_sub_77_carry_3_, npu_inst_pe_1_6_4_sub_77_carry_2_,
         npu_inst_pe_1_6_4_sub_77_carry_1_, npu_inst_pe_1_6_4_add_79_carry_7_,
         npu_inst_pe_1_6_4_add_79_carry_6_, npu_inst_pe_1_6_4_add_79_carry_5_,
         npu_inst_pe_1_6_4_add_79_carry_4_, npu_inst_pe_1_6_4_add_79_carry_3_,
         npu_inst_pe_1_6_4_add_79_carry_2_, npu_inst_pe_1_6_4_add_79_carry_1_,
         npu_inst_pe_1_6_4_n97, npu_inst_pe_1_6_4_n96, npu_inst_pe_1_6_4_n95,
         npu_inst_pe_1_6_4_n94, npu_inst_pe_1_6_4_n93, npu_inst_pe_1_6_4_n92,
         npu_inst_pe_1_6_4_n91, npu_inst_pe_1_6_4_n90, npu_inst_pe_1_6_4_n89,
         npu_inst_pe_1_6_4_n88, npu_inst_pe_1_6_4_n87, npu_inst_pe_1_6_4_n86,
         npu_inst_pe_1_6_4_n85, npu_inst_pe_1_6_4_n84, npu_inst_pe_1_6_4_n83,
         npu_inst_pe_1_6_4_n82, npu_inst_pe_1_6_4_n81, npu_inst_pe_1_6_4_n80,
         npu_inst_pe_1_6_4_n79, npu_inst_pe_1_6_4_n78, npu_inst_pe_1_6_4_n77,
         npu_inst_pe_1_6_4_n76, npu_inst_pe_1_6_4_n75, npu_inst_pe_1_6_4_n74,
         npu_inst_pe_1_6_4_n73, npu_inst_pe_1_6_4_n72, npu_inst_pe_1_6_4_n71,
         npu_inst_pe_1_6_4_n70, npu_inst_pe_1_6_4_n69, npu_inst_pe_1_6_4_n68,
         npu_inst_pe_1_6_4_n67, npu_inst_pe_1_6_4_n66, npu_inst_pe_1_6_4_n65,
         npu_inst_pe_1_6_4_n64, npu_inst_pe_1_6_4_n63, npu_inst_pe_1_6_4_n62,
         npu_inst_pe_1_6_4_n61, npu_inst_pe_1_6_4_n60, npu_inst_pe_1_6_4_n59,
         npu_inst_pe_1_6_4_n58, npu_inst_pe_1_6_4_n57, npu_inst_pe_1_6_4_n56,
         npu_inst_pe_1_6_4_n55, npu_inst_pe_1_6_4_n54, npu_inst_pe_1_6_4_n53,
         npu_inst_pe_1_6_4_n52, npu_inst_pe_1_6_4_n51, npu_inst_pe_1_6_4_n50,
         npu_inst_pe_1_6_4_n49, npu_inst_pe_1_6_4_n48, npu_inst_pe_1_6_4_n47,
         npu_inst_pe_1_6_4_n46, npu_inst_pe_1_6_4_n45, npu_inst_pe_1_6_4_n44,
         npu_inst_pe_1_6_4_n43, npu_inst_pe_1_6_4_n42, npu_inst_pe_1_6_4_n41,
         npu_inst_pe_1_6_4_n40, npu_inst_pe_1_6_4_n39, npu_inst_pe_1_6_4_n38,
         npu_inst_pe_1_6_4_n37, npu_inst_pe_1_6_4_n27, npu_inst_pe_1_6_4_n26,
         npu_inst_pe_1_6_4_net3103, npu_inst_pe_1_6_4_net3097,
         npu_inst_pe_1_6_4_N94, npu_inst_pe_1_6_4_N93, npu_inst_pe_1_6_4_N84,
         npu_inst_pe_1_6_4_N80, npu_inst_pe_1_6_4_N79, npu_inst_pe_1_6_4_N78,
         npu_inst_pe_1_6_4_N77, npu_inst_pe_1_6_4_N76, npu_inst_pe_1_6_4_N75,
         npu_inst_pe_1_6_4_N74, npu_inst_pe_1_6_4_N73, npu_inst_pe_1_6_4_N72,
         npu_inst_pe_1_6_4_N71, npu_inst_pe_1_6_4_N70, npu_inst_pe_1_6_4_N69,
         npu_inst_pe_1_6_4_N68, npu_inst_pe_1_6_4_N67, npu_inst_pe_1_6_4_N66,
         npu_inst_pe_1_6_4_N65, npu_inst_pe_1_6_4_int_q_acc_0_,
         npu_inst_pe_1_6_4_int_q_acc_1_, npu_inst_pe_1_6_4_int_q_acc_2_,
         npu_inst_pe_1_6_4_int_q_acc_3_, npu_inst_pe_1_6_4_int_q_acc_4_,
         npu_inst_pe_1_6_4_int_q_acc_5_, npu_inst_pe_1_6_4_int_q_acc_6_,
         npu_inst_pe_1_6_4_int_q_acc_7_, npu_inst_pe_1_6_4_int_data_0_,
         npu_inst_pe_1_6_4_int_data_1_, npu_inst_pe_1_6_4_int_q_weight_0_,
         npu_inst_pe_1_6_4_int_q_weight_1_,
         npu_inst_pe_1_6_4_int_q_reg_v_5__0_,
         npu_inst_pe_1_6_4_int_q_reg_v_5__1_,
         npu_inst_pe_1_6_4_int_q_reg_v_4__0_,
         npu_inst_pe_1_6_4_int_q_reg_v_4__1_,
         npu_inst_pe_1_6_4_int_q_reg_v_3__0_,
         npu_inst_pe_1_6_4_int_q_reg_v_3__1_,
         npu_inst_pe_1_6_4_int_q_reg_v_2__0_,
         npu_inst_pe_1_6_4_int_q_reg_v_2__1_,
         npu_inst_pe_1_6_4_int_q_reg_v_1__0_,
         npu_inst_pe_1_6_4_int_q_reg_v_1__1_,
         npu_inst_pe_1_6_4_int_q_reg_v_0__0_,
         npu_inst_pe_1_6_4_int_q_reg_v_0__1_,
         npu_inst_pe_1_6_4_int_q_reg_h_5__0_,
         npu_inst_pe_1_6_4_int_q_reg_h_5__1_,
         npu_inst_pe_1_6_4_int_q_reg_h_4__0_,
         npu_inst_pe_1_6_4_int_q_reg_h_4__1_,
         npu_inst_pe_1_6_4_int_q_reg_h_3__0_,
         npu_inst_pe_1_6_4_int_q_reg_h_3__1_,
         npu_inst_pe_1_6_4_int_q_reg_h_2__0_,
         npu_inst_pe_1_6_4_int_q_reg_h_2__1_,
         npu_inst_pe_1_6_4_int_q_reg_h_1__0_,
         npu_inst_pe_1_6_4_int_q_reg_h_1__1_,
         npu_inst_pe_1_6_4_int_q_reg_h_0__0_,
         npu_inst_pe_1_6_4_int_q_reg_h_0__1_, npu_inst_pe_1_6_5_n119,
         npu_inst_pe_1_6_5_n118, npu_inst_pe_1_6_5_n117,
         npu_inst_pe_1_6_5_n116, npu_inst_pe_1_6_5_n115,
         npu_inst_pe_1_6_5_n114, npu_inst_pe_1_6_5_n113,
         npu_inst_pe_1_6_5_n112, npu_inst_pe_1_6_5_n111,
         npu_inst_pe_1_6_5_n110, npu_inst_pe_1_6_5_n109,
         npu_inst_pe_1_6_5_n108, npu_inst_pe_1_6_5_n107,
         npu_inst_pe_1_6_5_n106, npu_inst_pe_1_6_5_n105,
         npu_inst_pe_1_6_5_n104, npu_inst_pe_1_6_5_n103,
         npu_inst_pe_1_6_5_n102, npu_inst_pe_1_6_5_n101,
         npu_inst_pe_1_6_5_n100, npu_inst_pe_1_6_5_n99, npu_inst_pe_1_6_5_n98,
         npu_inst_pe_1_6_5_n36, npu_inst_pe_1_6_5_n35, npu_inst_pe_1_6_5_n34,
         npu_inst_pe_1_6_5_n33, npu_inst_pe_1_6_5_n32, npu_inst_pe_1_6_5_n31,
         npu_inst_pe_1_6_5_n30, npu_inst_pe_1_6_5_n29, npu_inst_pe_1_6_5_n28,
         npu_inst_pe_1_6_5_n25, npu_inst_pe_1_6_5_n24, npu_inst_pe_1_6_5_n23,
         npu_inst_pe_1_6_5_n22, npu_inst_pe_1_6_5_n21, npu_inst_pe_1_6_5_n20,
         npu_inst_pe_1_6_5_n19, npu_inst_pe_1_6_5_n18, npu_inst_pe_1_6_5_n17,
         npu_inst_pe_1_6_5_n16, npu_inst_pe_1_6_5_n15, npu_inst_pe_1_6_5_n14,
         npu_inst_pe_1_6_5_n13, npu_inst_pe_1_6_5_n12, npu_inst_pe_1_6_5_n11,
         npu_inst_pe_1_6_5_n10, npu_inst_pe_1_6_5_n9, npu_inst_pe_1_6_5_n8,
         npu_inst_pe_1_6_5_n7, npu_inst_pe_1_6_5_n6, npu_inst_pe_1_6_5_n5,
         npu_inst_pe_1_6_5_n4, npu_inst_pe_1_6_5_n3, npu_inst_pe_1_6_5_n2,
         npu_inst_pe_1_6_5_n1, npu_inst_pe_1_6_5_sub_77_carry_7_,
         npu_inst_pe_1_6_5_sub_77_carry_6_, npu_inst_pe_1_6_5_sub_77_carry_5_,
         npu_inst_pe_1_6_5_sub_77_carry_4_, npu_inst_pe_1_6_5_sub_77_carry_3_,
         npu_inst_pe_1_6_5_sub_77_carry_2_, npu_inst_pe_1_6_5_sub_77_carry_1_,
         npu_inst_pe_1_6_5_add_79_carry_7_, npu_inst_pe_1_6_5_add_79_carry_6_,
         npu_inst_pe_1_6_5_add_79_carry_5_, npu_inst_pe_1_6_5_add_79_carry_4_,
         npu_inst_pe_1_6_5_add_79_carry_3_, npu_inst_pe_1_6_5_add_79_carry_2_,
         npu_inst_pe_1_6_5_add_79_carry_1_, npu_inst_pe_1_6_5_n97,
         npu_inst_pe_1_6_5_n96, npu_inst_pe_1_6_5_n95, npu_inst_pe_1_6_5_n94,
         npu_inst_pe_1_6_5_n93, npu_inst_pe_1_6_5_n92, npu_inst_pe_1_6_5_n91,
         npu_inst_pe_1_6_5_n90, npu_inst_pe_1_6_5_n89, npu_inst_pe_1_6_5_n88,
         npu_inst_pe_1_6_5_n87, npu_inst_pe_1_6_5_n86, npu_inst_pe_1_6_5_n85,
         npu_inst_pe_1_6_5_n84, npu_inst_pe_1_6_5_n83, npu_inst_pe_1_6_5_n82,
         npu_inst_pe_1_6_5_n81, npu_inst_pe_1_6_5_n80, npu_inst_pe_1_6_5_n79,
         npu_inst_pe_1_6_5_n78, npu_inst_pe_1_6_5_n77, npu_inst_pe_1_6_5_n76,
         npu_inst_pe_1_6_5_n75, npu_inst_pe_1_6_5_n74, npu_inst_pe_1_6_5_n73,
         npu_inst_pe_1_6_5_n72, npu_inst_pe_1_6_5_n71, npu_inst_pe_1_6_5_n70,
         npu_inst_pe_1_6_5_n69, npu_inst_pe_1_6_5_n68, npu_inst_pe_1_6_5_n67,
         npu_inst_pe_1_6_5_n66, npu_inst_pe_1_6_5_n65, npu_inst_pe_1_6_5_n64,
         npu_inst_pe_1_6_5_n63, npu_inst_pe_1_6_5_n62, npu_inst_pe_1_6_5_n61,
         npu_inst_pe_1_6_5_n60, npu_inst_pe_1_6_5_n59, npu_inst_pe_1_6_5_n58,
         npu_inst_pe_1_6_5_n57, npu_inst_pe_1_6_5_n56, npu_inst_pe_1_6_5_n55,
         npu_inst_pe_1_6_5_n54, npu_inst_pe_1_6_5_n53, npu_inst_pe_1_6_5_n52,
         npu_inst_pe_1_6_5_n51, npu_inst_pe_1_6_5_n50, npu_inst_pe_1_6_5_n49,
         npu_inst_pe_1_6_5_n48, npu_inst_pe_1_6_5_n47, npu_inst_pe_1_6_5_n46,
         npu_inst_pe_1_6_5_n45, npu_inst_pe_1_6_5_n44, npu_inst_pe_1_6_5_n43,
         npu_inst_pe_1_6_5_n42, npu_inst_pe_1_6_5_n41, npu_inst_pe_1_6_5_n40,
         npu_inst_pe_1_6_5_n39, npu_inst_pe_1_6_5_n38, npu_inst_pe_1_6_5_n37,
         npu_inst_pe_1_6_5_n27, npu_inst_pe_1_6_5_n26,
         npu_inst_pe_1_6_5_net3080, npu_inst_pe_1_6_5_net3074,
         npu_inst_pe_1_6_5_N94, npu_inst_pe_1_6_5_N93, npu_inst_pe_1_6_5_N84,
         npu_inst_pe_1_6_5_N80, npu_inst_pe_1_6_5_N79, npu_inst_pe_1_6_5_N78,
         npu_inst_pe_1_6_5_N77, npu_inst_pe_1_6_5_N76, npu_inst_pe_1_6_5_N75,
         npu_inst_pe_1_6_5_N74, npu_inst_pe_1_6_5_N73, npu_inst_pe_1_6_5_N72,
         npu_inst_pe_1_6_5_N71, npu_inst_pe_1_6_5_N70, npu_inst_pe_1_6_5_N69,
         npu_inst_pe_1_6_5_N68, npu_inst_pe_1_6_5_N67, npu_inst_pe_1_6_5_N66,
         npu_inst_pe_1_6_5_N65, npu_inst_pe_1_6_5_int_q_acc_0_,
         npu_inst_pe_1_6_5_int_q_acc_1_, npu_inst_pe_1_6_5_int_q_acc_2_,
         npu_inst_pe_1_6_5_int_q_acc_3_, npu_inst_pe_1_6_5_int_q_acc_4_,
         npu_inst_pe_1_6_5_int_q_acc_5_, npu_inst_pe_1_6_5_int_q_acc_6_,
         npu_inst_pe_1_6_5_int_q_acc_7_, npu_inst_pe_1_6_5_int_data_0_,
         npu_inst_pe_1_6_5_int_data_1_, npu_inst_pe_1_6_5_int_q_weight_0_,
         npu_inst_pe_1_6_5_int_q_weight_1_,
         npu_inst_pe_1_6_5_int_q_reg_v_5__0_,
         npu_inst_pe_1_6_5_int_q_reg_v_5__1_,
         npu_inst_pe_1_6_5_int_q_reg_v_4__0_,
         npu_inst_pe_1_6_5_int_q_reg_v_4__1_,
         npu_inst_pe_1_6_5_int_q_reg_v_3__0_,
         npu_inst_pe_1_6_5_int_q_reg_v_3__1_,
         npu_inst_pe_1_6_5_int_q_reg_v_2__0_,
         npu_inst_pe_1_6_5_int_q_reg_v_2__1_,
         npu_inst_pe_1_6_5_int_q_reg_v_1__0_,
         npu_inst_pe_1_6_5_int_q_reg_v_1__1_,
         npu_inst_pe_1_6_5_int_q_reg_v_0__0_,
         npu_inst_pe_1_6_5_int_q_reg_v_0__1_,
         npu_inst_pe_1_6_5_int_q_reg_h_5__0_,
         npu_inst_pe_1_6_5_int_q_reg_h_5__1_,
         npu_inst_pe_1_6_5_int_q_reg_h_4__0_,
         npu_inst_pe_1_6_5_int_q_reg_h_4__1_,
         npu_inst_pe_1_6_5_int_q_reg_h_3__0_,
         npu_inst_pe_1_6_5_int_q_reg_h_3__1_,
         npu_inst_pe_1_6_5_int_q_reg_h_2__0_,
         npu_inst_pe_1_6_5_int_q_reg_h_2__1_,
         npu_inst_pe_1_6_5_int_q_reg_h_1__0_,
         npu_inst_pe_1_6_5_int_q_reg_h_1__1_,
         npu_inst_pe_1_6_5_int_q_reg_h_0__0_,
         npu_inst_pe_1_6_5_int_q_reg_h_0__1_, npu_inst_pe_1_6_6_n119,
         npu_inst_pe_1_6_6_n118, npu_inst_pe_1_6_6_n117,
         npu_inst_pe_1_6_6_n116, npu_inst_pe_1_6_6_n115,
         npu_inst_pe_1_6_6_n114, npu_inst_pe_1_6_6_n113,
         npu_inst_pe_1_6_6_n112, npu_inst_pe_1_6_6_n111,
         npu_inst_pe_1_6_6_n110, npu_inst_pe_1_6_6_n109,
         npu_inst_pe_1_6_6_n108, npu_inst_pe_1_6_6_n107,
         npu_inst_pe_1_6_6_n106, npu_inst_pe_1_6_6_n105,
         npu_inst_pe_1_6_6_n104, npu_inst_pe_1_6_6_n103,
         npu_inst_pe_1_6_6_n102, npu_inst_pe_1_6_6_n101,
         npu_inst_pe_1_6_6_n100, npu_inst_pe_1_6_6_n99, npu_inst_pe_1_6_6_n98,
         npu_inst_pe_1_6_6_n36, npu_inst_pe_1_6_6_n35, npu_inst_pe_1_6_6_n34,
         npu_inst_pe_1_6_6_n33, npu_inst_pe_1_6_6_n32, npu_inst_pe_1_6_6_n31,
         npu_inst_pe_1_6_6_n30, npu_inst_pe_1_6_6_n29, npu_inst_pe_1_6_6_n28,
         npu_inst_pe_1_6_6_n25, npu_inst_pe_1_6_6_n24, npu_inst_pe_1_6_6_n23,
         npu_inst_pe_1_6_6_n22, npu_inst_pe_1_6_6_n21, npu_inst_pe_1_6_6_n20,
         npu_inst_pe_1_6_6_n19, npu_inst_pe_1_6_6_n18, npu_inst_pe_1_6_6_n17,
         npu_inst_pe_1_6_6_n16, npu_inst_pe_1_6_6_n15, npu_inst_pe_1_6_6_n14,
         npu_inst_pe_1_6_6_n13, npu_inst_pe_1_6_6_n12, npu_inst_pe_1_6_6_n11,
         npu_inst_pe_1_6_6_n10, npu_inst_pe_1_6_6_n9, npu_inst_pe_1_6_6_n8,
         npu_inst_pe_1_6_6_n7, npu_inst_pe_1_6_6_n6, npu_inst_pe_1_6_6_n5,
         npu_inst_pe_1_6_6_n4, npu_inst_pe_1_6_6_n3, npu_inst_pe_1_6_6_n2,
         npu_inst_pe_1_6_6_n1, npu_inst_pe_1_6_6_sub_77_carry_7_,
         npu_inst_pe_1_6_6_sub_77_carry_6_, npu_inst_pe_1_6_6_sub_77_carry_5_,
         npu_inst_pe_1_6_6_sub_77_carry_4_, npu_inst_pe_1_6_6_sub_77_carry_3_,
         npu_inst_pe_1_6_6_sub_77_carry_2_, npu_inst_pe_1_6_6_sub_77_carry_1_,
         npu_inst_pe_1_6_6_add_79_carry_7_, npu_inst_pe_1_6_6_add_79_carry_6_,
         npu_inst_pe_1_6_6_add_79_carry_5_, npu_inst_pe_1_6_6_add_79_carry_4_,
         npu_inst_pe_1_6_6_add_79_carry_3_, npu_inst_pe_1_6_6_add_79_carry_2_,
         npu_inst_pe_1_6_6_add_79_carry_1_, npu_inst_pe_1_6_6_n97,
         npu_inst_pe_1_6_6_n96, npu_inst_pe_1_6_6_n95, npu_inst_pe_1_6_6_n94,
         npu_inst_pe_1_6_6_n93, npu_inst_pe_1_6_6_n92, npu_inst_pe_1_6_6_n91,
         npu_inst_pe_1_6_6_n90, npu_inst_pe_1_6_6_n89, npu_inst_pe_1_6_6_n88,
         npu_inst_pe_1_6_6_n87, npu_inst_pe_1_6_6_n86, npu_inst_pe_1_6_6_n85,
         npu_inst_pe_1_6_6_n84, npu_inst_pe_1_6_6_n83, npu_inst_pe_1_6_6_n82,
         npu_inst_pe_1_6_6_n81, npu_inst_pe_1_6_6_n80, npu_inst_pe_1_6_6_n79,
         npu_inst_pe_1_6_6_n78, npu_inst_pe_1_6_6_n77, npu_inst_pe_1_6_6_n76,
         npu_inst_pe_1_6_6_n75, npu_inst_pe_1_6_6_n74, npu_inst_pe_1_6_6_n73,
         npu_inst_pe_1_6_6_n72, npu_inst_pe_1_6_6_n71, npu_inst_pe_1_6_6_n70,
         npu_inst_pe_1_6_6_n69, npu_inst_pe_1_6_6_n68, npu_inst_pe_1_6_6_n67,
         npu_inst_pe_1_6_6_n66, npu_inst_pe_1_6_6_n65, npu_inst_pe_1_6_6_n64,
         npu_inst_pe_1_6_6_n63, npu_inst_pe_1_6_6_n62, npu_inst_pe_1_6_6_n61,
         npu_inst_pe_1_6_6_n60, npu_inst_pe_1_6_6_n59, npu_inst_pe_1_6_6_n58,
         npu_inst_pe_1_6_6_n57, npu_inst_pe_1_6_6_n56, npu_inst_pe_1_6_6_n55,
         npu_inst_pe_1_6_6_n54, npu_inst_pe_1_6_6_n53, npu_inst_pe_1_6_6_n52,
         npu_inst_pe_1_6_6_n51, npu_inst_pe_1_6_6_n50, npu_inst_pe_1_6_6_n49,
         npu_inst_pe_1_6_6_n48, npu_inst_pe_1_6_6_n47, npu_inst_pe_1_6_6_n46,
         npu_inst_pe_1_6_6_n45, npu_inst_pe_1_6_6_n44, npu_inst_pe_1_6_6_n43,
         npu_inst_pe_1_6_6_n42, npu_inst_pe_1_6_6_n41, npu_inst_pe_1_6_6_n40,
         npu_inst_pe_1_6_6_n39, npu_inst_pe_1_6_6_n38, npu_inst_pe_1_6_6_n37,
         npu_inst_pe_1_6_6_n27, npu_inst_pe_1_6_6_n26,
         npu_inst_pe_1_6_6_net3057, npu_inst_pe_1_6_6_net3051,
         npu_inst_pe_1_6_6_N94, npu_inst_pe_1_6_6_N93, npu_inst_pe_1_6_6_N84,
         npu_inst_pe_1_6_6_N80, npu_inst_pe_1_6_6_N79, npu_inst_pe_1_6_6_N78,
         npu_inst_pe_1_6_6_N77, npu_inst_pe_1_6_6_N76, npu_inst_pe_1_6_6_N75,
         npu_inst_pe_1_6_6_N74, npu_inst_pe_1_6_6_N73, npu_inst_pe_1_6_6_N72,
         npu_inst_pe_1_6_6_N71, npu_inst_pe_1_6_6_N70, npu_inst_pe_1_6_6_N69,
         npu_inst_pe_1_6_6_N68, npu_inst_pe_1_6_6_N67, npu_inst_pe_1_6_6_N66,
         npu_inst_pe_1_6_6_N65, npu_inst_pe_1_6_6_int_q_acc_0_,
         npu_inst_pe_1_6_6_int_q_acc_1_, npu_inst_pe_1_6_6_int_q_acc_2_,
         npu_inst_pe_1_6_6_int_q_acc_3_, npu_inst_pe_1_6_6_int_q_acc_4_,
         npu_inst_pe_1_6_6_int_q_acc_5_, npu_inst_pe_1_6_6_int_q_acc_6_,
         npu_inst_pe_1_6_6_int_q_acc_7_, npu_inst_pe_1_6_6_int_data_0_,
         npu_inst_pe_1_6_6_int_data_1_, npu_inst_pe_1_6_6_int_q_weight_0_,
         npu_inst_pe_1_6_6_int_q_weight_1_,
         npu_inst_pe_1_6_6_int_q_reg_v_5__0_,
         npu_inst_pe_1_6_6_int_q_reg_v_5__1_,
         npu_inst_pe_1_6_6_int_q_reg_v_4__0_,
         npu_inst_pe_1_6_6_int_q_reg_v_4__1_,
         npu_inst_pe_1_6_6_int_q_reg_v_3__0_,
         npu_inst_pe_1_6_6_int_q_reg_v_3__1_,
         npu_inst_pe_1_6_6_int_q_reg_v_2__0_,
         npu_inst_pe_1_6_6_int_q_reg_v_2__1_,
         npu_inst_pe_1_6_6_int_q_reg_v_1__0_,
         npu_inst_pe_1_6_6_int_q_reg_v_1__1_,
         npu_inst_pe_1_6_6_int_q_reg_v_0__0_,
         npu_inst_pe_1_6_6_int_q_reg_v_0__1_,
         npu_inst_pe_1_6_6_int_q_reg_h_5__0_,
         npu_inst_pe_1_6_6_int_q_reg_h_5__1_,
         npu_inst_pe_1_6_6_int_q_reg_h_4__0_,
         npu_inst_pe_1_6_6_int_q_reg_h_4__1_,
         npu_inst_pe_1_6_6_int_q_reg_h_3__0_,
         npu_inst_pe_1_6_6_int_q_reg_h_3__1_,
         npu_inst_pe_1_6_6_int_q_reg_h_2__0_,
         npu_inst_pe_1_6_6_int_q_reg_h_2__1_,
         npu_inst_pe_1_6_6_int_q_reg_h_1__0_,
         npu_inst_pe_1_6_6_int_q_reg_h_1__1_,
         npu_inst_pe_1_6_6_int_q_reg_h_0__0_,
         npu_inst_pe_1_6_6_int_q_reg_h_0__1_, npu_inst_pe_1_6_7_n119,
         npu_inst_pe_1_6_7_n118, npu_inst_pe_1_6_7_n117,
         npu_inst_pe_1_6_7_n116, npu_inst_pe_1_6_7_n115,
         npu_inst_pe_1_6_7_n114, npu_inst_pe_1_6_7_n113,
         npu_inst_pe_1_6_7_n112, npu_inst_pe_1_6_7_n111,
         npu_inst_pe_1_6_7_n110, npu_inst_pe_1_6_7_n109,
         npu_inst_pe_1_6_7_n108, npu_inst_pe_1_6_7_n107,
         npu_inst_pe_1_6_7_n106, npu_inst_pe_1_6_7_n105,
         npu_inst_pe_1_6_7_n104, npu_inst_pe_1_6_7_n103,
         npu_inst_pe_1_6_7_n102, npu_inst_pe_1_6_7_n101,
         npu_inst_pe_1_6_7_n100, npu_inst_pe_1_6_7_n99, npu_inst_pe_1_6_7_n98,
         npu_inst_pe_1_6_7_n36, npu_inst_pe_1_6_7_n35, npu_inst_pe_1_6_7_n34,
         npu_inst_pe_1_6_7_n33, npu_inst_pe_1_6_7_n32, npu_inst_pe_1_6_7_n31,
         npu_inst_pe_1_6_7_n30, npu_inst_pe_1_6_7_n29, npu_inst_pe_1_6_7_n28,
         npu_inst_pe_1_6_7_n25, npu_inst_pe_1_6_7_n24, npu_inst_pe_1_6_7_n23,
         npu_inst_pe_1_6_7_n22, npu_inst_pe_1_6_7_n21, npu_inst_pe_1_6_7_n20,
         npu_inst_pe_1_6_7_n19, npu_inst_pe_1_6_7_n18, npu_inst_pe_1_6_7_n17,
         npu_inst_pe_1_6_7_n16, npu_inst_pe_1_6_7_n15, npu_inst_pe_1_6_7_n14,
         npu_inst_pe_1_6_7_n13, npu_inst_pe_1_6_7_n12, npu_inst_pe_1_6_7_n11,
         npu_inst_pe_1_6_7_n10, npu_inst_pe_1_6_7_n9, npu_inst_pe_1_6_7_n8,
         npu_inst_pe_1_6_7_n7, npu_inst_pe_1_6_7_n6, npu_inst_pe_1_6_7_n5,
         npu_inst_pe_1_6_7_n4, npu_inst_pe_1_6_7_n3, npu_inst_pe_1_6_7_n2,
         npu_inst_pe_1_6_7_n1, npu_inst_pe_1_6_7_sub_77_carry_7_,
         npu_inst_pe_1_6_7_sub_77_carry_6_, npu_inst_pe_1_6_7_sub_77_carry_5_,
         npu_inst_pe_1_6_7_sub_77_carry_4_, npu_inst_pe_1_6_7_sub_77_carry_3_,
         npu_inst_pe_1_6_7_sub_77_carry_2_, npu_inst_pe_1_6_7_sub_77_carry_1_,
         npu_inst_pe_1_6_7_add_79_carry_7_, npu_inst_pe_1_6_7_add_79_carry_6_,
         npu_inst_pe_1_6_7_add_79_carry_5_, npu_inst_pe_1_6_7_add_79_carry_4_,
         npu_inst_pe_1_6_7_add_79_carry_3_, npu_inst_pe_1_6_7_add_79_carry_2_,
         npu_inst_pe_1_6_7_add_79_carry_1_, npu_inst_pe_1_6_7_n97,
         npu_inst_pe_1_6_7_n96, npu_inst_pe_1_6_7_n95, npu_inst_pe_1_6_7_n94,
         npu_inst_pe_1_6_7_n93, npu_inst_pe_1_6_7_n92, npu_inst_pe_1_6_7_n91,
         npu_inst_pe_1_6_7_n90, npu_inst_pe_1_6_7_n89, npu_inst_pe_1_6_7_n88,
         npu_inst_pe_1_6_7_n87, npu_inst_pe_1_6_7_n86, npu_inst_pe_1_6_7_n85,
         npu_inst_pe_1_6_7_n84, npu_inst_pe_1_6_7_n83, npu_inst_pe_1_6_7_n82,
         npu_inst_pe_1_6_7_n81, npu_inst_pe_1_6_7_n80, npu_inst_pe_1_6_7_n79,
         npu_inst_pe_1_6_7_n78, npu_inst_pe_1_6_7_n77, npu_inst_pe_1_6_7_n76,
         npu_inst_pe_1_6_7_n75, npu_inst_pe_1_6_7_n74, npu_inst_pe_1_6_7_n73,
         npu_inst_pe_1_6_7_n72, npu_inst_pe_1_6_7_n71, npu_inst_pe_1_6_7_n70,
         npu_inst_pe_1_6_7_n69, npu_inst_pe_1_6_7_n68, npu_inst_pe_1_6_7_n67,
         npu_inst_pe_1_6_7_n66, npu_inst_pe_1_6_7_n65, npu_inst_pe_1_6_7_n64,
         npu_inst_pe_1_6_7_n63, npu_inst_pe_1_6_7_n62, npu_inst_pe_1_6_7_n61,
         npu_inst_pe_1_6_7_n60, npu_inst_pe_1_6_7_n59, npu_inst_pe_1_6_7_n58,
         npu_inst_pe_1_6_7_n57, npu_inst_pe_1_6_7_n56, npu_inst_pe_1_6_7_n55,
         npu_inst_pe_1_6_7_n54, npu_inst_pe_1_6_7_n53, npu_inst_pe_1_6_7_n52,
         npu_inst_pe_1_6_7_n51, npu_inst_pe_1_6_7_n50, npu_inst_pe_1_6_7_n49,
         npu_inst_pe_1_6_7_n48, npu_inst_pe_1_6_7_n47, npu_inst_pe_1_6_7_n46,
         npu_inst_pe_1_6_7_n45, npu_inst_pe_1_6_7_n44, npu_inst_pe_1_6_7_n43,
         npu_inst_pe_1_6_7_n42, npu_inst_pe_1_6_7_n41, npu_inst_pe_1_6_7_n40,
         npu_inst_pe_1_6_7_n39, npu_inst_pe_1_6_7_n38, npu_inst_pe_1_6_7_n37,
         npu_inst_pe_1_6_7_n27, npu_inst_pe_1_6_7_n26,
         npu_inst_pe_1_6_7_net3034, npu_inst_pe_1_6_7_net3028,
         npu_inst_pe_1_6_7_N94, npu_inst_pe_1_6_7_N93, npu_inst_pe_1_6_7_N84,
         npu_inst_pe_1_6_7_N80, npu_inst_pe_1_6_7_N79, npu_inst_pe_1_6_7_N78,
         npu_inst_pe_1_6_7_N77, npu_inst_pe_1_6_7_N76, npu_inst_pe_1_6_7_N75,
         npu_inst_pe_1_6_7_N74, npu_inst_pe_1_6_7_N73, npu_inst_pe_1_6_7_N72,
         npu_inst_pe_1_6_7_N71, npu_inst_pe_1_6_7_N70, npu_inst_pe_1_6_7_N69,
         npu_inst_pe_1_6_7_N68, npu_inst_pe_1_6_7_N67, npu_inst_pe_1_6_7_N66,
         npu_inst_pe_1_6_7_N65, npu_inst_pe_1_6_7_int_q_acc_0_,
         npu_inst_pe_1_6_7_int_q_acc_1_, npu_inst_pe_1_6_7_int_q_acc_2_,
         npu_inst_pe_1_6_7_int_q_acc_3_, npu_inst_pe_1_6_7_int_q_acc_4_,
         npu_inst_pe_1_6_7_int_q_acc_5_, npu_inst_pe_1_6_7_int_q_acc_6_,
         npu_inst_pe_1_6_7_int_q_acc_7_, npu_inst_pe_1_6_7_int_data_0_,
         npu_inst_pe_1_6_7_int_data_1_, npu_inst_pe_1_6_7_int_q_weight_0_,
         npu_inst_pe_1_6_7_int_q_weight_1_,
         npu_inst_pe_1_6_7_int_q_reg_v_5__0_,
         npu_inst_pe_1_6_7_int_q_reg_v_5__1_,
         npu_inst_pe_1_6_7_int_q_reg_v_4__0_,
         npu_inst_pe_1_6_7_int_q_reg_v_4__1_,
         npu_inst_pe_1_6_7_int_q_reg_v_3__0_,
         npu_inst_pe_1_6_7_int_q_reg_v_3__1_,
         npu_inst_pe_1_6_7_int_q_reg_v_2__0_,
         npu_inst_pe_1_6_7_int_q_reg_v_2__1_,
         npu_inst_pe_1_6_7_int_q_reg_v_1__0_,
         npu_inst_pe_1_6_7_int_q_reg_v_1__1_,
         npu_inst_pe_1_6_7_int_q_reg_v_0__0_,
         npu_inst_pe_1_6_7_int_q_reg_v_0__1_,
         npu_inst_pe_1_6_7_int_q_reg_h_5__0_,
         npu_inst_pe_1_6_7_int_q_reg_h_5__1_,
         npu_inst_pe_1_6_7_int_q_reg_h_4__0_,
         npu_inst_pe_1_6_7_int_q_reg_h_4__1_,
         npu_inst_pe_1_6_7_int_q_reg_h_3__0_,
         npu_inst_pe_1_6_7_int_q_reg_h_3__1_,
         npu_inst_pe_1_6_7_int_q_reg_h_2__0_,
         npu_inst_pe_1_6_7_int_q_reg_h_2__1_,
         npu_inst_pe_1_6_7_int_q_reg_h_1__0_,
         npu_inst_pe_1_6_7_int_q_reg_h_1__1_,
         npu_inst_pe_1_6_7_int_q_reg_h_0__0_,
         npu_inst_pe_1_6_7_int_q_reg_h_0__1_, npu_inst_pe_1_7_0_n119,
         npu_inst_pe_1_7_0_n118, npu_inst_pe_1_7_0_n117,
         npu_inst_pe_1_7_0_n116, npu_inst_pe_1_7_0_n115,
         npu_inst_pe_1_7_0_n114, npu_inst_pe_1_7_0_n113,
         npu_inst_pe_1_7_0_n112, npu_inst_pe_1_7_0_n111,
         npu_inst_pe_1_7_0_n110, npu_inst_pe_1_7_0_n109,
         npu_inst_pe_1_7_0_n108, npu_inst_pe_1_7_0_n107,
         npu_inst_pe_1_7_0_n106, npu_inst_pe_1_7_0_n105,
         npu_inst_pe_1_7_0_n104, npu_inst_pe_1_7_0_n103,
         npu_inst_pe_1_7_0_n102, npu_inst_pe_1_7_0_n101,
         npu_inst_pe_1_7_0_n100, npu_inst_pe_1_7_0_n99, npu_inst_pe_1_7_0_n98,
         npu_inst_pe_1_7_0_n36, npu_inst_pe_1_7_0_n35, npu_inst_pe_1_7_0_n34,
         npu_inst_pe_1_7_0_n33, npu_inst_pe_1_7_0_n32, npu_inst_pe_1_7_0_n31,
         npu_inst_pe_1_7_0_n30, npu_inst_pe_1_7_0_n29, npu_inst_pe_1_7_0_n28,
         npu_inst_pe_1_7_0_n25, npu_inst_pe_1_7_0_n24, npu_inst_pe_1_7_0_n23,
         npu_inst_pe_1_7_0_n22, npu_inst_pe_1_7_0_n21, npu_inst_pe_1_7_0_n20,
         npu_inst_pe_1_7_0_n19, npu_inst_pe_1_7_0_n18, npu_inst_pe_1_7_0_n17,
         npu_inst_pe_1_7_0_n16, npu_inst_pe_1_7_0_n15, npu_inst_pe_1_7_0_n14,
         npu_inst_pe_1_7_0_n13, npu_inst_pe_1_7_0_n12, npu_inst_pe_1_7_0_n11,
         npu_inst_pe_1_7_0_n10, npu_inst_pe_1_7_0_n9, npu_inst_pe_1_7_0_n8,
         npu_inst_pe_1_7_0_n7, npu_inst_pe_1_7_0_n6, npu_inst_pe_1_7_0_n5,
         npu_inst_pe_1_7_0_n4, npu_inst_pe_1_7_0_n3, npu_inst_pe_1_7_0_n2,
         npu_inst_pe_1_7_0_n1, npu_inst_pe_1_7_0_sub_77_carry_7_,
         npu_inst_pe_1_7_0_sub_77_carry_6_, npu_inst_pe_1_7_0_sub_77_carry_5_,
         npu_inst_pe_1_7_0_sub_77_carry_4_, npu_inst_pe_1_7_0_sub_77_carry_3_,
         npu_inst_pe_1_7_0_sub_77_carry_2_, npu_inst_pe_1_7_0_sub_77_carry_1_,
         npu_inst_pe_1_7_0_add_79_carry_7_, npu_inst_pe_1_7_0_add_79_carry_6_,
         npu_inst_pe_1_7_0_add_79_carry_5_, npu_inst_pe_1_7_0_add_79_carry_4_,
         npu_inst_pe_1_7_0_add_79_carry_3_, npu_inst_pe_1_7_0_add_79_carry_2_,
         npu_inst_pe_1_7_0_add_79_carry_1_, npu_inst_pe_1_7_0_n97,
         npu_inst_pe_1_7_0_n96, npu_inst_pe_1_7_0_n95, npu_inst_pe_1_7_0_n94,
         npu_inst_pe_1_7_0_n93, npu_inst_pe_1_7_0_n92, npu_inst_pe_1_7_0_n91,
         npu_inst_pe_1_7_0_n90, npu_inst_pe_1_7_0_n89, npu_inst_pe_1_7_0_n88,
         npu_inst_pe_1_7_0_n87, npu_inst_pe_1_7_0_n86, npu_inst_pe_1_7_0_n85,
         npu_inst_pe_1_7_0_n84, npu_inst_pe_1_7_0_n83, npu_inst_pe_1_7_0_n82,
         npu_inst_pe_1_7_0_n81, npu_inst_pe_1_7_0_n80, npu_inst_pe_1_7_0_n79,
         npu_inst_pe_1_7_0_n78, npu_inst_pe_1_7_0_n77, npu_inst_pe_1_7_0_n76,
         npu_inst_pe_1_7_0_n75, npu_inst_pe_1_7_0_n74, npu_inst_pe_1_7_0_n73,
         npu_inst_pe_1_7_0_n72, npu_inst_pe_1_7_0_n71, npu_inst_pe_1_7_0_n70,
         npu_inst_pe_1_7_0_n69, npu_inst_pe_1_7_0_n68, npu_inst_pe_1_7_0_n67,
         npu_inst_pe_1_7_0_n66, npu_inst_pe_1_7_0_n65, npu_inst_pe_1_7_0_n64,
         npu_inst_pe_1_7_0_n63, npu_inst_pe_1_7_0_n62, npu_inst_pe_1_7_0_n61,
         npu_inst_pe_1_7_0_n60, npu_inst_pe_1_7_0_n59, npu_inst_pe_1_7_0_n58,
         npu_inst_pe_1_7_0_n57, npu_inst_pe_1_7_0_n56, npu_inst_pe_1_7_0_n55,
         npu_inst_pe_1_7_0_n54, npu_inst_pe_1_7_0_n53, npu_inst_pe_1_7_0_n52,
         npu_inst_pe_1_7_0_n51, npu_inst_pe_1_7_0_n50, npu_inst_pe_1_7_0_n49,
         npu_inst_pe_1_7_0_n48, npu_inst_pe_1_7_0_n47, npu_inst_pe_1_7_0_n46,
         npu_inst_pe_1_7_0_n45, npu_inst_pe_1_7_0_n44, npu_inst_pe_1_7_0_n43,
         npu_inst_pe_1_7_0_n42, npu_inst_pe_1_7_0_n41, npu_inst_pe_1_7_0_n40,
         npu_inst_pe_1_7_0_n39, npu_inst_pe_1_7_0_n38, npu_inst_pe_1_7_0_n37,
         npu_inst_pe_1_7_0_n27, npu_inst_pe_1_7_0_n26,
         npu_inst_pe_1_7_0_net3011, npu_inst_pe_1_7_0_net3005,
         npu_inst_pe_1_7_0_N94, npu_inst_pe_1_7_0_N93, npu_inst_pe_1_7_0_N84,
         npu_inst_pe_1_7_0_N80, npu_inst_pe_1_7_0_N79, npu_inst_pe_1_7_0_N78,
         npu_inst_pe_1_7_0_N77, npu_inst_pe_1_7_0_N76, npu_inst_pe_1_7_0_N75,
         npu_inst_pe_1_7_0_N74, npu_inst_pe_1_7_0_N73, npu_inst_pe_1_7_0_N72,
         npu_inst_pe_1_7_0_N71, npu_inst_pe_1_7_0_N70, npu_inst_pe_1_7_0_N69,
         npu_inst_pe_1_7_0_N68, npu_inst_pe_1_7_0_N67, npu_inst_pe_1_7_0_N66,
         npu_inst_pe_1_7_0_N65, npu_inst_pe_1_7_0_int_q_acc_0_,
         npu_inst_pe_1_7_0_int_q_acc_1_, npu_inst_pe_1_7_0_int_q_acc_2_,
         npu_inst_pe_1_7_0_int_q_acc_3_, npu_inst_pe_1_7_0_int_q_acc_4_,
         npu_inst_pe_1_7_0_int_q_acc_5_, npu_inst_pe_1_7_0_int_q_acc_6_,
         npu_inst_pe_1_7_0_int_q_acc_7_, npu_inst_pe_1_7_0_int_data_0_,
         npu_inst_pe_1_7_0_int_data_1_, npu_inst_pe_1_7_0_int_q_weight_0_,
         npu_inst_pe_1_7_0_int_q_weight_1_,
         npu_inst_pe_1_7_0_int_q_reg_v_5__0_,
         npu_inst_pe_1_7_0_int_q_reg_v_5__1_,
         npu_inst_pe_1_7_0_int_q_reg_v_4__0_,
         npu_inst_pe_1_7_0_int_q_reg_v_4__1_,
         npu_inst_pe_1_7_0_int_q_reg_v_3__0_,
         npu_inst_pe_1_7_0_int_q_reg_v_3__1_,
         npu_inst_pe_1_7_0_int_q_reg_v_2__0_,
         npu_inst_pe_1_7_0_int_q_reg_v_2__1_,
         npu_inst_pe_1_7_0_int_q_reg_v_1__0_,
         npu_inst_pe_1_7_0_int_q_reg_v_1__1_,
         npu_inst_pe_1_7_0_int_q_reg_v_0__0_,
         npu_inst_pe_1_7_0_int_q_reg_v_0__1_,
         npu_inst_pe_1_7_0_int_q_reg_h_5__0_,
         npu_inst_pe_1_7_0_int_q_reg_h_5__1_,
         npu_inst_pe_1_7_0_int_q_reg_h_4__0_,
         npu_inst_pe_1_7_0_int_q_reg_h_4__1_,
         npu_inst_pe_1_7_0_int_q_reg_h_3__0_,
         npu_inst_pe_1_7_0_int_q_reg_h_3__1_,
         npu_inst_pe_1_7_0_int_q_reg_h_2__0_,
         npu_inst_pe_1_7_0_int_q_reg_h_2__1_,
         npu_inst_pe_1_7_0_int_q_reg_h_1__0_,
         npu_inst_pe_1_7_0_int_q_reg_h_1__1_,
         npu_inst_pe_1_7_0_int_q_reg_h_0__0_,
         npu_inst_pe_1_7_0_int_q_reg_h_0__1_, npu_inst_pe_1_7_0_o_data_h_0_,
         npu_inst_pe_1_7_0_o_data_h_1_, npu_inst_pe_1_7_1_n119,
         npu_inst_pe_1_7_1_n118, npu_inst_pe_1_7_1_n117,
         npu_inst_pe_1_7_1_n116, npu_inst_pe_1_7_1_n115,
         npu_inst_pe_1_7_1_n114, npu_inst_pe_1_7_1_n113,
         npu_inst_pe_1_7_1_n112, npu_inst_pe_1_7_1_n111,
         npu_inst_pe_1_7_1_n110, npu_inst_pe_1_7_1_n109,
         npu_inst_pe_1_7_1_n108, npu_inst_pe_1_7_1_n107,
         npu_inst_pe_1_7_1_n106, npu_inst_pe_1_7_1_n105,
         npu_inst_pe_1_7_1_n104, npu_inst_pe_1_7_1_n103,
         npu_inst_pe_1_7_1_n102, npu_inst_pe_1_7_1_n101,
         npu_inst_pe_1_7_1_n100, npu_inst_pe_1_7_1_n99, npu_inst_pe_1_7_1_n98,
         npu_inst_pe_1_7_1_n36, npu_inst_pe_1_7_1_n35, npu_inst_pe_1_7_1_n34,
         npu_inst_pe_1_7_1_n33, npu_inst_pe_1_7_1_n32, npu_inst_pe_1_7_1_n31,
         npu_inst_pe_1_7_1_n30, npu_inst_pe_1_7_1_n29, npu_inst_pe_1_7_1_n28,
         npu_inst_pe_1_7_1_n25, npu_inst_pe_1_7_1_n24, npu_inst_pe_1_7_1_n23,
         npu_inst_pe_1_7_1_n22, npu_inst_pe_1_7_1_n21, npu_inst_pe_1_7_1_n20,
         npu_inst_pe_1_7_1_n19, npu_inst_pe_1_7_1_n18, npu_inst_pe_1_7_1_n17,
         npu_inst_pe_1_7_1_n16, npu_inst_pe_1_7_1_n15, npu_inst_pe_1_7_1_n14,
         npu_inst_pe_1_7_1_n13, npu_inst_pe_1_7_1_n12, npu_inst_pe_1_7_1_n11,
         npu_inst_pe_1_7_1_n10, npu_inst_pe_1_7_1_n9, npu_inst_pe_1_7_1_n8,
         npu_inst_pe_1_7_1_n7, npu_inst_pe_1_7_1_n6, npu_inst_pe_1_7_1_n5,
         npu_inst_pe_1_7_1_n4, npu_inst_pe_1_7_1_n3, npu_inst_pe_1_7_1_n2,
         npu_inst_pe_1_7_1_n1, npu_inst_pe_1_7_1_sub_77_carry_7_,
         npu_inst_pe_1_7_1_sub_77_carry_6_, npu_inst_pe_1_7_1_sub_77_carry_5_,
         npu_inst_pe_1_7_1_sub_77_carry_4_, npu_inst_pe_1_7_1_sub_77_carry_3_,
         npu_inst_pe_1_7_1_sub_77_carry_2_, npu_inst_pe_1_7_1_sub_77_carry_1_,
         npu_inst_pe_1_7_1_add_79_carry_7_, npu_inst_pe_1_7_1_add_79_carry_6_,
         npu_inst_pe_1_7_1_add_79_carry_5_, npu_inst_pe_1_7_1_add_79_carry_4_,
         npu_inst_pe_1_7_1_add_79_carry_3_, npu_inst_pe_1_7_1_add_79_carry_2_,
         npu_inst_pe_1_7_1_add_79_carry_1_, npu_inst_pe_1_7_1_n97,
         npu_inst_pe_1_7_1_n96, npu_inst_pe_1_7_1_n95, npu_inst_pe_1_7_1_n94,
         npu_inst_pe_1_7_1_n93, npu_inst_pe_1_7_1_n92, npu_inst_pe_1_7_1_n91,
         npu_inst_pe_1_7_1_n90, npu_inst_pe_1_7_1_n89, npu_inst_pe_1_7_1_n88,
         npu_inst_pe_1_7_1_n87, npu_inst_pe_1_7_1_n86, npu_inst_pe_1_7_1_n85,
         npu_inst_pe_1_7_1_n84, npu_inst_pe_1_7_1_n83, npu_inst_pe_1_7_1_n82,
         npu_inst_pe_1_7_1_n81, npu_inst_pe_1_7_1_n80, npu_inst_pe_1_7_1_n79,
         npu_inst_pe_1_7_1_n78, npu_inst_pe_1_7_1_n77, npu_inst_pe_1_7_1_n76,
         npu_inst_pe_1_7_1_n75, npu_inst_pe_1_7_1_n74, npu_inst_pe_1_7_1_n73,
         npu_inst_pe_1_7_1_n72, npu_inst_pe_1_7_1_n71, npu_inst_pe_1_7_1_n70,
         npu_inst_pe_1_7_1_n69, npu_inst_pe_1_7_1_n68, npu_inst_pe_1_7_1_n67,
         npu_inst_pe_1_7_1_n66, npu_inst_pe_1_7_1_n65, npu_inst_pe_1_7_1_n64,
         npu_inst_pe_1_7_1_n63, npu_inst_pe_1_7_1_n62, npu_inst_pe_1_7_1_n61,
         npu_inst_pe_1_7_1_n60, npu_inst_pe_1_7_1_n59, npu_inst_pe_1_7_1_n58,
         npu_inst_pe_1_7_1_n57, npu_inst_pe_1_7_1_n56, npu_inst_pe_1_7_1_n55,
         npu_inst_pe_1_7_1_n54, npu_inst_pe_1_7_1_n53, npu_inst_pe_1_7_1_n52,
         npu_inst_pe_1_7_1_n51, npu_inst_pe_1_7_1_n50, npu_inst_pe_1_7_1_n49,
         npu_inst_pe_1_7_1_n48, npu_inst_pe_1_7_1_n47, npu_inst_pe_1_7_1_n46,
         npu_inst_pe_1_7_1_n45, npu_inst_pe_1_7_1_n44, npu_inst_pe_1_7_1_n43,
         npu_inst_pe_1_7_1_n42, npu_inst_pe_1_7_1_n41, npu_inst_pe_1_7_1_n40,
         npu_inst_pe_1_7_1_n39, npu_inst_pe_1_7_1_n38, npu_inst_pe_1_7_1_n37,
         npu_inst_pe_1_7_1_n27, npu_inst_pe_1_7_1_n26,
         npu_inst_pe_1_7_1_net2988, npu_inst_pe_1_7_1_net2982,
         npu_inst_pe_1_7_1_N94, npu_inst_pe_1_7_1_N93, npu_inst_pe_1_7_1_N84,
         npu_inst_pe_1_7_1_N80, npu_inst_pe_1_7_1_N79, npu_inst_pe_1_7_1_N78,
         npu_inst_pe_1_7_1_N77, npu_inst_pe_1_7_1_N76, npu_inst_pe_1_7_1_N75,
         npu_inst_pe_1_7_1_N74, npu_inst_pe_1_7_1_N73, npu_inst_pe_1_7_1_N72,
         npu_inst_pe_1_7_1_N71, npu_inst_pe_1_7_1_N70, npu_inst_pe_1_7_1_N69,
         npu_inst_pe_1_7_1_N68, npu_inst_pe_1_7_1_N67, npu_inst_pe_1_7_1_N66,
         npu_inst_pe_1_7_1_N65, npu_inst_pe_1_7_1_int_q_acc_0_,
         npu_inst_pe_1_7_1_int_q_acc_1_, npu_inst_pe_1_7_1_int_q_acc_2_,
         npu_inst_pe_1_7_1_int_q_acc_3_, npu_inst_pe_1_7_1_int_q_acc_4_,
         npu_inst_pe_1_7_1_int_q_acc_5_, npu_inst_pe_1_7_1_int_q_acc_6_,
         npu_inst_pe_1_7_1_int_q_acc_7_, npu_inst_pe_1_7_1_int_data_0_,
         npu_inst_pe_1_7_1_int_data_1_, npu_inst_pe_1_7_1_int_q_weight_0_,
         npu_inst_pe_1_7_1_int_q_weight_1_,
         npu_inst_pe_1_7_1_int_q_reg_v_5__0_,
         npu_inst_pe_1_7_1_int_q_reg_v_5__1_,
         npu_inst_pe_1_7_1_int_q_reg_v_4__0_,
         npu_inst_pe_1_7_1_int_q_reg_v_4__1_,
         npu_inst_pe_1_7_1_int_q_reg_v_3__0_,
         npu_inst_pe_1_7_1_int_q_reg_v_3__1_,
         npu_inst_pe_1_7_1_int_q_reg_v_2__0_,
         npu_inst_pe_1_7_1_int_q_reg_v_2__1_,
         npu_inst_pe_1_7_1_int_q_reg_v_1__0_,
         npu_inst_pe_1_7_1_int_q_reg_v_1__1_,
         npu_inst_pe_1_7_1_int_q_reg_v_0__0_,
         npu_inst_pe_1_7_1_int_q_reg_v_0__1_,
         npu_inst_pe_1_7_1_int_q_reg_h_5__0_,
         npu_inst_pe_1_7_1_int_q_reg_h_5__1_,
         npu_inst_pe_1_7_1_int_q_reg_h_4__0_,
         npu_inst_pe_1_7_1_int_q_reg_h_4__1_,
         npu_inst_pe_1_7_1_int_q_reg_h_3__0_,
         npu_inst_pe_1_7_1_int_q_reg_h_3__1_,
         npu_inst_pe_1_7_1_int_q_reg_h_2__0_,
         npu_inst_pe_1_7_1_int_q_reg_h_2__1_,
         npu_inst_pe_1_7_1_int_q_reg_h_1__0_,
         npu_inst_pe_1_7_1_int_q_reg_h_1__1_,
         npu_inst_pe_1_7_1_int_q_reg_h_0__0_,
         npu_inst_pe_1_7_1_int_q_reg_h_0__1_, npu_inst_pe_1_7_2_n119,
         npu_inst_pe_1_7_2_n118, npu_inst_pe_1_7_2_n117,
         npu_inst_pe_1_7_2_n116, npu_inst_pe_1_7_2_n115,
         npu_inst_pe_1_7_2_n114, npu_inst_pe_1_7_2_n113,
         npu_inst_pe_1_7_2_n112, npu_inst_pe_1_7_2_n111,
         npu_inst_pe_1_7_2_n110, npu_inst_pe_1_7_2_n109,
         npu_inst_pe_1_7_2_n108, npu_inst_pe_1_7_2_n107,
         npu_inst_pe_1_7_2_n106, npu_inst_pe_1_7_2_n105,
         npu_inst_pe_1_7_2_n104, npu_inst_pe_1_7_2_n103,
         npu_inst_pe_1_7_2_n102, npu_inst_pe_1_7_2_n101,
         npu_inst_pe_1_7_2_n100, npu_inst_pe_1_7_2_n99, npu_inst_pe_1_7_2_n98,
         npu_inst_pe_1_7_2_n36, npu_inst_pe_1_7_2_n35, npu_inst_pe_1_7_2_n34,
         npu_inst_pe_1_7_2_n33, npu_inst_pe_1_7_2_n32, npu_inst_pe_1_7_2_n31,
         npu_inst_pe_1_7_2_n30, npu_inst_pe_1_7_2_n29, npu_inst_pe_1_7_2_n28,
         npu_inst_pe_1_7_2_n25, npu_inst_pe_1_7_2_n24, npu_inst_pe_1_7_2_n23,
         npu_inst_pe_1_7_2_n22, npu_inst_pe_1_7_2_n21, npu_inst_pe_1_7_2_n20,
         npu_inst_pe_1_7_2_n19, npu_inst_pe_1_7_2_n18, npu_inst_pe_1_7_2_n17,
         npu_inst_pe_1_7_2_n16, npu_inst_pe_1_7_2_n15, npu_inst_pe_1_7_2_n14,
         npu_inst_pe_1_7_2_n13, npu_inst_pe_1_7_2_n12, npu_inst_pe_1_7_2_n11,
         npu_inst_pe_1_7_2_n10, npu_inst_pe_1_7_2_n9, npu_inst_pe_1_7_2_n8,
         npu_inst_pe_1_7_2_n7, npu_inst_pe_1_7_2_n6, npu_inst_pe_1_7_2_n5,
         npu_inst_pe_1_7_2_n4, npu_inst_pe_1_7_2_n3, npu_inst_pe_1_7_2_n2,
         npu_inst_pe_1_7_2_n1, npu_inst_pe_1_7_2_sub_77_carry_7_,
         npu_inst_pe_1_7_2_sub_77_carry_6_, npu_inst_pe_1_7_2_sub_77_carry_5_,
         npu_inst_pe_1_7_2_sub_77_carry_4_, npu_inst_pe_1_7_2_sub_77_carry_3_,
         npu_inst_pe_1_7_2_sub_77_carry_2_, npu_inst_pe_1_7_2_sub_77_carry_1_,
         npu_inst_pe_1_7_2_add_79_carry_7_, npu_inst_pe_1_7_2_add_79_carry_6_,
         npu_inst_pe_1_7_2_add_79_carry_5_, npu_inst_pe_1_7_2_add_79_carry_4_,
         npu_inst_pe_1_7_2_add_79_carry_3_, npu_inst_pe_1_7_2_add_79_carry_2_,
         npu_inst_pe_1_7_2_add_79_carry_1_, npu_inst_pe_1_7_2_n97,
         npu_inst_pe_1_7_2_n96, npu_inst_pe_1_7_2_n95, npu_inst_pe_1_7_2_n94,
         npu_inst_pe_1_7_2_n93, npu_inst_pe_1_7_2_n92, npu_inst_pe_1_7_2_n91,
         npu_inst_pe_1_7_2_n90, npu_inst_pe_1_7_2_n89, npu_inst_pe_1_7_2_n88,
         npu_inst_pe_1_7_2_n87, npu_inst_pe_1_7_2_n86, npu_inst_pe_1_7_2_n85,
         npu_inst_pe_1_7_2_n84, npu_inst_pe_1_7_2_n83, npu_inst_pe_1_7_2_n82,
         npu_inst_pe_1_7_2_n81, npu_inst_pe_1_7_2_n80, npu_inst_pe_1_7_2_n79,
         npu_inst_pe_1_7_2_n78, npu_inst_pe_1_7_2_n77, npu_inst_pe_1_7_2_n76,
         npu_inst_pe_1_7_2_n75, npu_inst_pe_1_7_2_n74, npu_inst_pe_1_7_2_n73,
         npu_inst_pe_1_7_2_n72, npu_inst_pe_1_7_2_n71, npu_inst_pe_1_7_2_n70,
         npu_inst_pe_1_7_2_n69, npu_inst_pe_1_7_2_n68, npu_inst_pe_1_7_2_n67,
         npu_inst_pe_1_7_2_n66, npu_inst_pe_1_7_2_n65, npu_inst_pe_1_7_2_n64,
         npu_inst_pe_1_7_2_n63, npu_inst_pe_1_7_2_n62, npu_inst_pe_1_7_2_n61,
         npu_inst_pe_1_7_2_n60, npu_inst_pe_1_7_2_n59, npu_inst_pe_1_7_2_n58,
         npu_inst_pe_1_7_2_n57, npu_inst_pe_1_7_2_n56, npu_inst_pe_1_7_2_n55,
         npu_inst_pe_1_7_2_n54, npu_inst_pe_1_7_2_n53, npu_inst_pe_1_7_2_n52,
         npu_inst_pe_1_7_2_n51, npu_inst_pe_1_7_2_n50, npu_inst_pe_1_7_2_n49,
         npu_inst_pe_1_7_2_n48, npu_inst_pe_1_7_2_n47, npu_inst_pe_1_7_2_n46,
         npu_inst_pe_1_7_2_n45, npu_inst_pe_1_7_2_n44, npu_inst_pe_1_7_2_n43,
         npu_inst_pe_1_7_2_n42, npu_inst_pe_1_7_2_n41, npu_inst_pe_1_7_2_n40,
         npu_inst_pe_1_7_2_n39, npu_inst_pe_1_7_2_n38, npu_inst_pe_1_7_2_n37,
         npu_inst_pe_1_7_2_n27, npu_inst_pe_1_7_2_n26,
         npu_inst_pe_1_7_2_net2965, npu_inst_pe_1_7_2_net2959,
         npu_inst_pe_1_7_2_N94, npu_inst_pe_1_7_2_N93, npu_inst_pe_1_7_2_N84,
         npu_inst_pe_1_7_2_N80, npu_inst_pe_1_7_2_N79, npu_inst_pe_1_7_2_N78,
         npu_inst_pe_1_7_2_N77, npu_inst_pe_1_7_2_N76, npu_inst_pe_1_7_2_N75,
         npu_inst_pe_1_7_2_N74, npu_inst_pe_1_7_2_N73, npu_inst_pe_1_7_2_N72,
         npu_inst_pe_1_7_2_N71, npu_inst_pe_1_7_2_N70, npu_inst_pe_1_7_2_N69,
         npu_inst_pe_1_7_2_N68, npu_inst_pe_1_7_2_N67, npu_inst_pe_1_7_2_N66,
         npu_inst_pe_1_7_2_N65, npu_inst_pe_1_7_2_int_q_acc_0_,
         npu_inst_pe_1_7_2_int_q_acc_1_, npu_inst_pe_1_7_2_int_q_acc_2_,
         npu_inst_pe_1_7_2_int_q_acc_3_, npu_inst_pe_1_7_2_int_q_acc_4_,
         npu_inst_pe_1_7_2_int_q_acc_5_, npu_inst_pe_1_7_2_int_q_acc_6_,
         npu_inst_pe_1_7_2_int_q_acc_7_, npu_inst_pe_1_7_2_int_data_0_,
         npu_inst_pe_1_7_2_int_data_1_, npu_inst_pe_1_7_2_int_q_weight_0_,
         npu_inst_pe_1_7_2_int_q_weight_1_,
         npu_inst_pe_1_7_2_int_q_reg_v_5__0_,
         npu_inst_pe_1_7_2_int_q_reg_v_5__1_,
         npu_inst_pe_1_7_2_int_q_reg_v_4__0_,
         npu_inst_pe_1_7_2_int_q_reg_v_4__1_,
         npu_inst_pe_1_7_2_int_q_reg_v_3__0_,
         npu_inst_pe_1_7_2_int_q_reg_v_3__1_,
         npu_inst_pe_1_7_2_int_q_reg_v_2__0_,
         npu_inst_pe_1_7_2_int_q_reg_v_2__1_,
         npu_inst_pe_1_7_2_int_q_reg_v_1__0_,
         npu_inst_pe_1_7_2_int_q_reg_v_1__1_,
         npu_inst_pe_1_7_2_int_q_reg_v_0__0_,
         npu_inst_pe_1_7_2_int_q_reg_v_0__1_,
         npu_inst_pe_1_7_2_int_q_reg_h_5__0_,
         npu_inst_pe_1_7_2_int_q_reg_h_5__1_,
         npu_inst_pe_1_7_2_int_q_reg_h_4__0_,
         npu_inst_pe_1_7_2_int_q_reg_h_4__1_,
         npu_inst_pe_1_7_2_int_q_reg_h_3__0_,
         npu_inst_pe_1_7_2_int_q_reg_h_3__1_,
         npu_inst_pe_1_7_2_int_q_reg_h_2__0_,
         npu_inst_pe_1_7_2_int_q_reg_h_2__1_,
         npu_inst_pe_1_7_2_int_q_reg_h_1__0_,
         npu_inst_pe_1_7_2_int_q_reg_h_1__1_,
         npu_inst_pe_1_7_2_int_q_reg_h_0__0_,
         npu_inst_pe_1_7_2_int_q_reg_h_0__1_, npu_inst_pe_1_7_3_n119,
         npu_inst_pe_1_7_3_n118, npu_inst_pe_1_7_3_n117,
         npu_inst_pe_1_7_3_n116, npu_inst_pe_1_7_3_n115,
         npu_inst_pe_1_7_3_n114, npu_inst_pe_1_7_3_n113,
         npu_inst_pe_1_7_3_n112, npu_inst_pe_1_7_3_n111,
         npu_inst_pe_1_7_3_n110, npu_inst_pe_1_7_3_n109,
         npu_inst_pe_1_7_3_n108, npu_inst_pe_1_7_3_n107,
         npu_inst_pe_1_7_3_n106, npu_inst_pe_1_7_3_n105,
         npu_inst_pe_1_7_3_n104, npu_inst_pe_1_7_3_n103,
         npu_inst_pe_1_7_3_n102, npu_inst_pe_1_7_3_n101,
         npu_inst_pe_1_7_3_n100, npu_inst_pe_1_7_3_n99, npu_inst_pe_1_7_3_n98,
         npu_inst_pe_1_7_3_n36, npu_inst_pe_1_7_3_n35, npu_inst_pe_1_7_3_n34,
         npu_inst_pe_1_7_3_n33, npu_inst_pe_1_7_3_n32, npu_inst_pe_1_7_3_n31,
         npu_inst_pe_1_7_3_n30, npu_inst_pe_1_7_3_n29, npu_inst_pe_1_7_3_n28,
         npu_inst_pe_1_7_3_n25, npu_inst_pe_1_7_3_n24, npu_inst_pe_1_7_3_n23,
         npu_inst_pe_1_7_3_n22, npu_inst_pe_1_7_3_n21, npu_inst_pe_1_7_3_n20,
         npu_inst_pe_1_7_3_n19, npu_inst_pe_1_7_3_n18, npu_inst_pe_1_7_3_n17,
         npu_inst_pe_1_7_3_n16, npu_inst_pe_1_7_3_n15, npu_inst_pe_1_7_3_n14,
         npu_inst_pe_1_7_3_n13, npu_inst_pe_1_7_3_n12, npu_inst_pe_1_7_3_n11,
         npu_inst_pe_1_7_3_n10, npu_inst_pe_1_7_3_n9, npu_inst_pe_1_7_3_n8,
         npu_inst_pe_1_7_3_n7, npu_inst_pe_1_7_3_n6, npu_inst_pe_1_7_3_n5,
         npu_inst_pe_1_7_3_n4, npu_inst_pe_1_7_3_n3, npu_inst_pe_1_7_3_n2,
         npu_inst_pe_1_7_3_n1, npu_inst_pe_1_7_3_sub_77_carry_7_,
         npu_inst_pe_1_7_3_sub_77_carry_6_, npu_inst_pe_1_7_3_sub_77_carry_5_,
         npu_inst_pe_1_7_3_sub_77_carry_4_, npu_inst_pe_1_7_3_sub_77_carry_3_,
         npu_inst_pe_1_7_3_sub_77_carry_2_, npu_inst_pe_1_7_3_sub_77_carry_1_,
         npu_inst_pe_1_7_3_add_79_carry_7_, npu_inst_pe_1_7_3_add_79_carry_6_,
         npu_inst_pe_1_7_3_add_79_carry_5_, npu_inst_pe_1_7_3_add_79_carry_4_,
         npu_inst_pe_1_7_3_add_79_carry_3_, npu_inst_pe_1_7_3_add_79_carry_2_,
         npu_inst_pe_1_7_3_add_79_carry_1_, npu_inst_pe_1_7_3_n97,
         npu_inst_pe_1_7_3_n96, npu_inst_pe_1_7_3_n95, npu_inst_pe_1_7_3_n94,
         npu_inst_pe_1_7_3_n93, npu_inst_pe_1_7_3_n92, npu_inst_pe_1_7_3_n91,
         npu_inst_pe_1_7_3_n90, npu_inst_pe_1_7_3_n89, npu_inst_pe_1_7_3_n88,
         npu_inst_pe_1_7_3_n87, npu_inst_pe_1_7_3_n86, npu_inst_pe_1_7_3_n85,
         npu_inst_pe_1_7_3_n84, npu_inst_pe_1_7_3_n83, npu_inst_pe_1_7_3_n82,
         npu_inst_pe_1_7_3_n81, npu_inst_pe_1_7_3_n80, npu_inst_pe_1_7_3_n79,
         npu_inst_pe_1_7_3_n78, npu_inst_pe_1_7_3_n77, npu_inst_pe_1_7_3_n76,
         npu_inst_pe_1_7_3_n75, npu_inst_pe_1_7_3_n74, npu_inst_pe_1_7_3_n73,
         npu_inst_pe_1_7_3_n72, npu_inst_pe_1_7_3_n71, npu_inst_pe_1_7_3_n70,
         npu_inst_pe_1_7_3_n69, npu_inst_pe_1_7_3_n68, npu_inst_pe_1_7_3_n67,
         npu_inst_pe_1_7_3_n66, npu_inst_pe_1_7_3_n65, npu_inst_pe_1_7_3_n64,
         npu_inst_pe_1_7_3_n63, npu_inst_pe_1_7_3_n62, npu_inst_pe_1_7_3_n61,
         npu_inst_pe_1_7_3_n60, npu_inst_pe_1_7_3_n59, npu_inst_pe_1_7_3_n58,
         npu_inst_pe_1_7_3_n57, npu_inst_pe_1_7_3_n56, npu_inst_pe_1_7_3_n55,
         npu_inst_pe_1_7_3_n54, npu_inst_pe_1_7_3_n53, npu_inst_pe_1_7_3_n52,
         npu_inst_pe_1_7_3_n51, npu_inst_pe_1_7_3_n50, npu_inst_pe_1_7_3_n49,
         npu_inst_pe_1_7_3_n48, npu_inst_pe_1_7_3_n47, npu_inst_pe_1_7_3_n46,
         npu_inst_pe_1_7_3_n45, npu_inst_pe_1_7_3_n44, npu_inst_pe_1_7_3_n43,
         npu_inst_pe_1_7_3_n42, npu_inst_pe_1_7_3_n41, npu_inst_pe_1_7_3_n40,
         npu_inst_pe_1_7_3_n39, npu_inst_pe_1_7_3_n38, npu_inst_pe_1_7_3_n37,
         npu_inst_pe_1_7_3_n27, npu_inst_pe_1_7_3_n26,
         npu_inst_pe_1_7_3_net2942, npu_inst_pe_1_7_3_net2936,
         npu_inst_pe_1_7_3_N94, npu_inst_pe_1_7_3_N93, npu_inst_pe_1_7_3_N84,
         npu_inst_pe_1_7_3_N80, npu_inst_pe_1_7_3_N79, npu_inst_pe_1_7_3_N78,
         npu_inst_pe_1_7_3_N77, npu_inst_pe_1_7_3_N76, npu_inst_pe_1_7_3_N75,
         npu_inst_pe_1_7_3_N74, npu_inst_pe_1_7_3_N73, npu_inst_pe_1_7_3_N72,
         npu_inst_pe_1_7_3_N71, npu_inst_pe_1_7_3_N70, npu_inst_pe_1_7_3_N69,
         npu_inst_pe_1_7_3_N68, npu_inst_pe_1_7_3_N67, npu_inst_pe_1_7_3_N66,
         npu_inst_pe_1_7_3_N65, npu_inst_pe_1_7_3_int_q_acc_0_,
         npu_inst_pe_1_7_3_int_q_acc_1_, npu_inst_pe_1_7_3_int_q_acc_2_,
         npu_inst_pe_1_7_3_int_q_acc_3_, npu_inst_pe_1_7_3_int_q_acc_4_,
         npu_inst_pe_1_7_3_int_q_acc_5_, npu_inst_pe_1_7_3_int_q_acc_6_,
         npu_inst_pe_1_7_3_int_q_acc_7_, npu_inst_pe_1_7_3_int_data_0_,
         npu_inst_pe_1_7_3_int_data_1_, npu_inst_pe_1_7_3_int_q_weight_0_,
         npu_inst_pe_1_7_3_int_q_weight_1_,
         npu_inst_pe_1_7_3_int_q_reg_v_5__0_,
         npu_inst_pe_1_7_3_int_q_reg_v_5__1_,
         npu_inst_pe_1_7_3_int_q_reg_v_4__0_,
         npu_inst_pe_1_7_3_int_q_reg_v_4__1_,
         npu_inst_pe_1_7_3_int_q_reg_v_3__0_,
         npu_inst_pe_1_7_3_int_q_reg_v_3__1_,
         npu_inst_pe_1_7_3_int_q_reg_v_2__0_,
         npu_inst_pe_1_7_3_int_q_reg_v_2__1_,
         npu_inst_pe_1_7_3_int_q_reg_v_1__0_,
         npu_inst_pe_1_7_3_int_q_reg_v_1__1_,
         npu_inst_pe_1_7_3_int_q_reg_v_0__0_,
         npu_inst_pe_1_7_3_int_q_reg_v_0__1_,
         npu_inst_pe_1_7_3_int_q_reg_h_5__0_,
         npu_inst_pe_1_7_3_int_q_reg_h_5__1_,
         npu_inst_pe_1_7_3_int_q_reg_h_4__0_,
         npu_inst_pe_1_7_3_int_q_reg_h_4__1_,
         npu_inst_pe_1_7_3_int_q_reg_h_3__0_,
         npu_inst_pe_1_7_3_int_q_reg_h_3__1_,
         npu_inst_pe_1_7_3_int_q_reg_h_2__0_,
         npu_inst_pe_1_7_3_int_q_reg_h_2__1_,
         npu_inst_pe_1_7_3_int_q_reg_h_1__0_,
         npu_inst_pe_1_7_3_int_q_reg_h_1__1_,
         npu_inst_pe_1_7_3_int_q_reg_h_0__0_,
         npu_inst_pe_1_7_3_int_q_reg_h_0__1_, npu_inst_pe_1_7_4_n119,
         npu_inst_pe_1_7_4_n118, npu_inst_pe_1_7_4_n117,
         npu_inst_pe_1_7_4_n116, npu_inst_pe_1_7_4_n115,
         npu_inst_pe_1_7_4_n114, npu_inst_pe_1_7_4_n113,
         npu_inst_pe_1_7_4_n112, npu_inst_pe_1_7_4_n111,
         npu_inst_pe_1_7_4_n110, npu_inst_pe_1_7_4_n109,
         npu_inst_pe_1_7_4_n108, npu_inst_pe_1_7_4_n107,
         npu_inst_pe_1_7_4_n106, npu_inst_pe_1_7_4_n105,
         npu_inst_pe_1_7_4_n104, npu_inst_pe_1_7_4_n103,
         npu_inst_pe_1_7_4_n102, npu_inst_pe_1_7_4_n101,
         npu_inst_pe_1_7_4_n100, npu_inst_pe_1_7_4_n99, npu_inst_pe_1_7_4_n98,
         npu_inst_pe_1_7_4_n36, npu_inst_pe_1_7_4_n35, npu_inst_pe_1_7_4_n34,
         npu_inst_pe_1_7_4_n33, npu_inst_pe_1_7_4_n32, npu_inst_pe_1_7_4_n31,
         npu_inst_pe_1_7_4_n30, npu_inst_pe_1_7_4_n29, npu_inst_pe_1_7_4_n28,
         npu_inst_pe_1_7_4_n25, npu_inst_pe_1_7_4_n24, npu_inst_pe_1_7_4_n23,
         npu_inst_pe_1_7_4_n22, npu_inst_pe_1_7_4_n21, npu_inst_pe_1_7_4_n20,
         npu_inst_pe_1_7_4_n19, npu_inst_pe_1_7_4_n18, npu_inst_pe_1_7_4_n17,
         npu_inst_pe_1_7_4_n16, npu_inst_pe_1_7_4_n15, npu_inst_pe_1_7_4_n14,
         npu_inst_pe_1_7_4_n13, npu_inst_pe_1_7_4_n12, npu_inst_pe_1_7_4_n11,
         npu_inst_pe_1_7_4_n10, npu_inst_pe_1_7_4_n9, npu_inst_pe_1_7_4_n8,
         npu_inst_pe_1_7_4_n7, npu_inst_pe_1_7_4_n6, npu_inst_pe_1_7_4_n5,
         npu_inst_pe_1_7_4_n4, npu_inst_pe_1_7_4_n3, npu_inst_pe_1_7_4_n2,
         npu_inst_pe_1_7_4_n1, npu_inst_pe_1_7_4_sub_77_carry_7_,
         npu_inst_pe_1_7_4_sub_77_carry_6_, npu_inst_pe_1_7_4_sub_77_carry_5_,
         npu_inst_pe_1_7_4_sub_77_carry_4_, npu_inst_pe_1_7_4_sub_77_carry_3_,
         npu_inst_pe_1_7_4_sub_77_carry_2_, npu_inst_pe_1_7_4_sub_77_carry_1_,
         npu_inst_pe_1_7_4_add_79_carry_7_, npu_inst_pe_1_7_4_add_79_carry_6_,
         npu_inst_pe_1_7_4_add_79_carry_5_, npu_inst_pe_1_7_4_add_79_carry_4_,
         npu_inst_pe_1_7_4_add_79_carry_3_, npu_inst_pe_1_7_4_add_79_carry_2_,
         npu_inst_pe_1_7_4_add_79_carry_1_, npu_inst_pe_1_7_4_n97,
         npu_inst_pe_1_7_4_n96, npu_inst_pe_1_7_4_n95, npu_inst_pe_1_7_4_n94,
         npu_inst_pe_1_7_4_n93, npu_inst_pe_1_7_4_n92, npu_inst_pe_1_7_4_n91,
         npu_inst_pe_1_7_4_n90, npu_inst_pe_1_7_4_n89, npu_inst_pe_1_7_4_n88,
         npu_inst_pe_1_7_4_n87, npu_inst_pe_1_7_4_n86, npu_inst_pe_1_7_4_n85,
         npu_inst_pe_1_7_4_n84, npu_inst_pe_1_7_4_n83, npu_inst_pe_1_7_4_n82,
         npu_inst_pe_1_7_4_n81, npu_inst_pe_1_7_4_n80, npu_inst_pe_1_7_4_n79,
         npu_inst_pe_1_7_4_n78, npu_inst_pe_1_7_4_n77, npu_inst_pe_1_7_4_n76,
         npu_inst_pe_1_7_4_n75, npu_inst_pe_1_7_4_n74, npu_inst_pe_1_7_4_n73,
         npu_inst_pe_1_7_4_n72, npu_inst_pe_1_7_4_n71, npu_inst_pe_1_7_4_n70,
         npu_inst_pe_1_7_4_n69, npu_inst_pe_1_7_4_n68, npu_inst_pe_1_7_4_n67,
         npu_inst_pe_1_7_4_n66, npu_inst_pe_1_7_4_n65, npu_inst_pe_1_7_4_n64,
         npu_inst_pe_1_7_4_n63, npu_inst_pe_1_7_4_n62, npu_inst_pe_1_7_4_n61,
         npu_inst_pe_1_7_4_n60, npu_inst_pe_1_7_4_n59, npu_inst_pe_1_7_4_n58,
         npu_inst_pe_1_7_4_n57, npu_inst_pe_1_7_4_n56, npu_inst_pe_1_7_4_n55,
         npu_inst_pe_1_7_4_n54, npu_inst_pe_1_7_4_n53, npu_inst_pe_1_7_4_n52,
         npu_inst_pe_1_7_4_n51, npu_inst_pe_1_7_4_n50, npu_inst_pe_1_7_4_n49,
         npu_inst_pe_1_7_4_n48, npu_inst_pe_1_7_4_n47, npu_inst_pe_1_7_4_n46,
         npu_inst_pe_1_7_4_n45, npu_inst_pe_1_7_4_n44, npu_inst_pe_1_7_4_n43,
         npu_inst_pe_1_7_4_n42, npu_inst_pe_1_7_4_n41, npu_inst_pe_1_7_4_n40,
         npu_inst_pe_1_7_4_n39, npu_inst_pe_1_7_4_n38, npu_inst_pe_1_7_4_n37,
         npu_inst_pe_1_7_4_n27, npu_inst_pe_1_7_4_n26,
         npu_inst_pe_1_7_4_net2919, npu_inst_pe_1_7_4_net2913,
         npu_inst_pe_1_7_4_N94, npu_inst_pe_1_7_4_N93, npu_inst_pe_1_7_4_N84,
         npu_inst_pe_1_7_4_N80, npu_inst_pe_1_7_4_N79, npu_inst_pe_1_7_4_N78,
         npu_inst_pe_1_7_4_N77, npu_inst_pe_1_7_4_N76, npu_inst_pe_1_7_4_N75,
         npu_inst_pe_1_7_4_N74, npu_inst_pe_1_7_4_N73, npu_inst_pe_1_7_4_N72,
         npu_inst_pe_1_7_4_N71, npu_inst_pe_1_7_4_N70, npu_inst_pe_1_7_4_N69,
         npu_inst_pe_1_7_4_N68, npu_inst_pe_1_7_4_N67, npu_inst_pe_1_7_4_N66,
         npu_inst_pe_1_7_4_N65, npu_inst_pe_1_7_4_int_q_acc_0_,
         npu_inst_pe_1_7_4_int_q_acc_1_, npu_inst_pe_1_7_4_int_q_acc_2_,
         npu_inst_pe_1_7_4_int_q_acc_3_, npu_inst_pe_1_7_4_int_q_acc_4_,
         npu_inst_pe_1_7_4_int_q_acc_5_, npu_inst_pe_1_7_4_int_q_acc_6_,
         npu_inst_pe_1_7_4_int_q_acc_7_, npu_inst_pe_1_7_4_int_data_0_,
         npu_inst_pe_1_7_4_int_data_1_, npu_inst_pe_1_7_4_int_q_weight_0_,
         npu_inst_pe_1_7_4_int_q_weight_1_,
         npu_inst_pe_1_7_4_int_q_reg_v_5__0_,
         npu_inst_pe_1_7_4_int_q_reg_v_5__1_,
         npu_inst_pe_1_7_4_int_q_reg_v_4__0_,
         npu_inst_pe_1_7_4_int_q_reg_v_4__1_,
         npu_inst_pe_1_7_4_int_q_reg_v_3__0_,
         npu_inst_pe_1_7_4_int_q_reg_v_3__1_,
         npu_inst_pe_1_7_4_int_q_reg_v_2__0_,
         npu_inst_pe_1_7_4_int_q_reg_v_2__1_,
         npu_inst_pe_1_7_4_int_q_reg_v_1__0_,
         npu_inst_pe_1_7_4_int_q_reg_v_1__1_,
         npu_inst_pe_1_7_4_int_q_reg_v_0__0_,
         npu_inst_pe_1_7_4_int_q_reg_v_0__1_,
         npu_inst_pe_1_7_4_int_q_reg_h_5__0_,
         npu_inst_pe_1_7_4_int_q_reg_h_5__1_,
         npu_inst_pe_1_7_4_int_q_reg_h_4__0_,
         npu_inst_pe_1_7_4_int_q_reg_h_4__1_,
         npu_inst_pe_1_7_4_int_q_reg_h_3__0_,
         npu_inst_pe_1_7_4_int_q_reg_h_3__1_,
         npu_inst_pe_1_7_4_int_q_reg_h_2__0_,
         npu_inst_pe_1_7_4_int_q_reg_h_2__1_,
         npu_inst_pe_1_7_4_int_q_reg_h_1__0_,
         npu_inst_pe_1_7_4_int_q_reg_h_1__1_,
         npu_inst_pe_1_7_4_int_q_reg_h_0__0_,
         npu_inst_pe_1_7_4_int_q_reg_h_0__1_, npu_inst_pe_1_7_5_n119,
         npu_inst_pe_1_7_5_n118, npu_inst_pe_1_7_5_n117,
         npu_inst_pe_1_7_5_n116, npu_inst_pe_1_7_5_n115,
         npu_inst_pe_1_7_5_n114, npu_inst_pe_1_7_5_n113,
         npu_inst_pe_1_7_5_n112, npu_inst_pe_1_7_5_n111,
         npu_inst_pe_1_7_5_n110, npu_inst_pe_1_7_5_n109,
         npu_inst_pe_1_7_5_n108, npu_inst_pe_1_7_5_n107,
         npu_inst_pe_1_7_5_n106, npu_inst_pe_1_7_5_n105,
         npu_inst_pe_1_7_5_n104, npu_inst_pe_1_7_5_n103,
         npu_inst_pe_1_7_5_n102, npu_inst_pe_1_7_5_n101,
         npu_inst_pe_1_7_5_n100, npu_inst_pe_1_7_5_n99, npu_inst_pe_1_7_5_n98,
         npu_inst_pe_1_7_5_n36, npu_inst_pe_1_7_5_n35, npu_inst_pe_1_7_5_n34,
         npu_inst_pe_1_7_5_n33, npu_inst_pe_1_7_5_n32, npu_inst_pe_1_7_5_n31,
         npu_inst_pe_1_7_5_n30, npu_inst_pe_1_7_5_n29, npu_inst_pe_1_7_5_n28,
         npu_inst_pe_1_7_5_n25, npu_inst_pe_1_7_5_n24, npu_inst_pe_1_7_5_n23,
         npu_inst_pe_1_7_5_n22, npu_inst_pe_1_7_5_n21, npu_inst_pe_1_7_5_n20,
         npu_inst_pe_1_7_5_n19, npu_inst_pe_1_7_5_n18, npu_inst_pe_1_7_5_n17,
         npu_inst_pe_1_7_5_n16, npu_inst_pe_1_7_5_n15, npu_inst_pe_1_7_5_n14,
         npu_inst_pe_1_7_5_n13, npu_inst_pe_1_7_5_n12, npu_inst_pe_1_7_5_n11,
         npu_inst_pe_1_7_5_n10, npu_inst_pe_1_7_5_n9, npu_inst_pe_1_7_5_n8,
         npu_inst_pe_1_7_5_n7, npu_inst_pe_1_7_5_n6, npu_inst_pe_1_7_5_n5,
         npu_inst_pe_1_7_5_n4, npu_inst_pe_1_7_5_n3, npu_inst_pe_1_7_5_n2,
         npu_inst_pe_1_7_5_n1, npu_inst_pe_1_7_5_sub_77_carry_7_,
         npu_inst_pe_1_7_5_sub_77_carry_6_, npu_inst_pe_1_7_5_sub_77_carry_5_,
         npu_inst_pe_1_7_5_sub_77_carry_4_, npu_inst_pe_1_7_5_sub_77_carry_3_,
         npu_inst_pe_1_7_5_sub_77_carry_2_, npu_inst_pe_1_7_5_sub_77_carry_1_,
         npu_inst_pe_1_7_5_add_79_carry_7_, npu_inst_pe_1_7_5_add_79_carry_6_,
         npu_inst_pe_1_7_5_add_79_carry_5_, npu_inst_pe_1_7_5_add_79_carry_4_,
         npu_inst_pe_1_7_5_add_79_carry_3_, npu_inst_pe_1_7_5_add_79_carry_2_,
         npu_inst_pe_1_7_5_add_79_carry_1_, npu_inst_pe_1_7_5_n97,
         npu_inst_pe_1_7_5_n96, npu_inst_pe_1_7_5_n95, npu_inst_pe_1_7_5_n94,
         npu_inst_pe_1_7_5_n93, npu_inst_pe_1_7_5_n92, npu_inst_pe_1_7_5_n91,
         npu_inst_pe_1_7_5_n90, npu_inst_pe_1_7_5_n89, npu_inst_pe_1_7_5_n88,
         npu_inst_pe_1_7_5_n87, npu_inst_pe_1_7_5_n86, npu_inst_pe_1_7_5_n85,
         npu_inst_pe_1_7_5_n84, npu_inst_pe_1_7_5_n83, npu_inst_pe_1_7_5_n82,
         npu_inst_pe_1_7_5_n81, npu_inst_pe_1_7_5_n80, npu_inst_pe_1_7_5_n79,
         npu_inst_pe_1_7_5_n78, npu_inst_pe_1_7_5_n77, npu_inst_pe_1_7_5_n76,
         npu_inst_pe_1_7_5_n75, npu_inst_pe_1_7_5_n74, npu_inst_pe_1_7_5_n73,
         npu_inst_pe_1_7_5_n72, npu_inst_pe_1_7_5_n71, npu_inst_pe_1_7_5_n70,
         npu_inst_pe_1_7_5_n69, npu_inst_pe_1_7_5_n68, npu_inst_pe_1_7_5_n67,
         npu_inst_pe_1_7_5_n66, npu_inst_pe_1_7_5_n65, npu_inst_pe_1_7_5_n64,
         npu_inst_pe_1_7_5_n63, npu_inst_pe_1_7_5_n62, npu_inst_pe_1_7_5_n61,
         npu_inst_pe_1_7_5_n60, npu_inst_pe_1_7_5_n59, npu_inst_pe_1_7_5_n58,
         npu_inst_pe_1_7_5_n57, npu_inst_pe_1_7_5_n56, npu_inst_pe_1_7_5_n55,
         npu_inst_pe_1_7_5_n54, npu_inst_pe_1_7_5_n53, npu_inst_pe_1_7_5_n52,
         npu_inst_pe_1_7_5_n51, npu_inst_pe_1_7_5_n50, npu_inst_pe_1_7_5_n49,
         npu_inst_pe_1_7_5_n48, npu_inst_pe_1_7_5_n47, npu_inst_pe_1_7_5_n46,
         npu_inst_pe_1_7_5_n45, npu_inst_pe_1_7_5_n44, npu_inst_pe_1_7_5_n43,
         npu_inst_pe_1_7_5_n42, npu_inst_pe_1_7_5_n41, npu_inst_pe_1_7_5_n40,
         npu_inst_pe_1_7_5_n39, npu_inst_pe_1_7_5_n38, npu_inst_pe_1_7_5_n37,
         npu_inst_pe_1_7_5_n27, npu_inst_pe_1_7_5_n26,
         npu_inst_pe_1_7_5_net2896, npu_inst_pe_1_7_5_net2890,
         npu_inst_pe_1_7_5_N94, npu_inst_pe_1_7_5_N93, npu_inst_pe_1_7_5_N84,
         npu_inst_pe_1_7_5_N80, npu_inst_pe_1_7_5_N79, npu_inst_pe_1_7_5_N78,
         npu_inst_pe_1_7_5_N77, npu_inst_pe_1_7_5_N76, npu_inst_pe_1_7_5_N75,
         npu_inst_pe_1_7_5_N74, npu_inst_pe_1_7_5_N73, npu_inst_pe_1_7_5_N72,
         npu_inst_pe_1_7_5_N71, npu_inst_pe_1_7_5_N70, npu_inst_pe_1_7_5_N69,
         npu_inst_pe_1_7_5_N68, npu_inst_pe_1_7_5_N67, npu_inst_pe_1_7_5_N66,
         npu_inst_pe_1_7_5_N65, npu_inst_pe_1_7_5_int_q_acc_0_,
         npu_inst_pe_1_7_5_int_q_acc_1_, npu_inst_pe_1_7_5_int_q_acc_2_,
         npu_inst_pe_1_7_5_int_q_acc_3_, npu_inst_pe_1_7_5_int_q_acc_4_,
         npu_inst_pe_1_7_5_int_q_acc_5_, npu_inst_pe_1_7_5_int_q_acc_6_,
         npu_inst_pe_1_7_5_int_q_acc_7_, npu_inst_pe_1_7_5_int_data_0_,
         npu_inst_pe_1_7_5_int_data_1_, npu_inst_pe_1_7_5_int_q_weight_0_,
         npu_inst_pe_1_7_5_int_q_weight_1_,
         npu_inst_pe_1_7_5_int_q_reg_v_5__0_,
         npu_inst_pe_1_7_5_int_q_reg_v_5__1_,
         npu_inst_pe_1_7_5_int_q_reg_v_4__0_,
         npu_inst_pe_1_7_5_int_q_reg_v_4__1_,
         npu_inst_pe_1_7_5_int_q_reg_v_3__0_,
         npu_inst_pe_1_7_5_int_q_reg_v_3__1_,
         npu_inst_pe_1_7_5_int_q_reg_v_2__0_,
         npu_inst_pe_1_7_5_int_q_reg_v_2__1_,
         npu_inst_pe_1_7_5_int_q_reg_v_1__0_,
         npu_inst_pe_1_7_5_int_q_reg_v_1__1_,
         npu_inst_pe_1_7_5_int_q_reg_v_0__0_,
         npu_inst_pe_1_7_5_int_q_reg_v_0__1_,
         npu_inst_pe_1_7_5_int_q_reg_h_5__0_,
         npu_inst_pe_1_7_5_int_q_reg_h_5__1_,
         npu_inst_pe_1_7_5_int_q_reg_h_4__0_,
         npu_inst_pe_1_7_5_int_q_reg_h_4__1_,
         npu_inst_pe_1_7_5_int_q_reg_h_3__0_,
         npu_inst_pe_1_7_5_int_q_reg_h_3__1_,
         npu_inst_pe_1_7_5_int_q_reg_h_2__0_,
         npu_inst_pe_1_7_5_int_q_reg_h_2__1_,
         npu_inst_pe_1_7_5_int_q_reg_h_1__0_,
         npu_inst_pe_1_7_5_int_q_reg_h_1__1_,
         npu_inst_pe_1_7_5_int_q_reg_h_0__0_,
         npu_inst_pe_1_7_5_int_q_reg_h_0__1_, npu_inst_pe_1_7_6_n119,
         npu_inst_pe_1_7_6_n118, npu_inst_pe_1_7_6_n117,
         npu_inst_pe_1_7_6_n116, npu_inst_pe_1_7_6_n115,
         npu_inst_pe_1_7_6_n114, npu_inst_pe_1_7_6_n113,
         npu_inst_pe_1_7_6_n112, npu_inst_pe_1_7_6_n111,
         npu_inst_pe_1_7_6_n110, npu_inst_pe_1_7_6_n109,
         npu_inst_pe_1_7_6_n108, npu_inst_pe_1_7_6_n107,
         npu_inst_pe_1_7_6_n106, npu_inst_pe_1_7_6_n105,
         npu_inst_pe_1_7_6_n104, npu_inst_pe_1_7_6_n103,
         npu_inst_pe_1_7_6_n102, npu_inst_pe_1_7_6_n101,
         npu_inst_pe_1_7_6_n100, npu_inst_pe_1_7_6_n99, npu_inst_pe_1_7_6_n98,
         npu_inst_pe_1_7_6_n36, npu_inst_pe_1_7_6_n35, npu_inst_pe_1_7_6_n34,
         npu_inst_pe_1_7_6_n33, npu_inst_pe_1_7_6_n32, npu_inst_pe_1_7_6_n31,
         npu_inst_pe_1_7_6_n30, npu_inst_pe_1_7_6_n29, npu_inst_pe_1_7_6_n28,
         npu_inst_pe_1_7_6_n25, npu_inst_pe_1_7_6_n24, npu_inst_pe_1_7_6_n23,
         npu_inst_pe_1_7_6_n22, npu_inst_pe_1_7_6_n21, npu_inst_pe_1_7_6_n20,
         npu_inst_pe_1_7_6_n19, npu_inst_pe_1_7_6_n18, npu_inst_pe_1_7_6_n17,
         npu_inst_pe_1_7_6_n16, npu_inst_pe_1_7_6_n15, npu_inst_pe_1_7_6_n14,
         npu_inst_pe_1_7_6_n13, npu_inst_pe_1_7_6_n12, npu_inst_pe_1_7_6_n11,
         npu_inst_pe_1_7_6_n10, npu_inst_pe_1_7_6_n9, npu_inst_pe_1_7_6_n8,
         npu_inst_pe_1_7_6_n7, npu_inst_pe_1_7_6_n6, npu_inst_pe_1_7_6_n5,
         npu_inst_pe_1_7_6_n4, npu_inst_pe_1_7_6_n3, npu_inst_pe_1_7_6_n2,
         npu_inst_pe_1_7_6_n1, npu_inst_pe_1_7_6_sub_77_carry_7_,
         npu_inst_pe_1_7_6_sub_77_carry_6_, npu_inst_pe_1_7_6_sub_77_carry_5_,
         npu_inst_pe_1_7_6_sub_77_carry_4_, npu_inst_pe_1_7_6_sub_77_carry_3_,
         npu_inst_pe_1_7_6_sub_77_carry_2_, npu_inst_pe_1_7_6_sub_77_carry_1_,
         npu_inst_pe_1_7_6_add_79_carry_7_, npu_inst_pe_1_7_6_add_79_carry_6_,
         npu_inst_pe_1_7_6_add_79_carry_5_, npu_inst_pe_1_7_6_add_79_carry_4_,
         npu_inst_pe_1_7_6_add_79_carry_3_, npu_inst_pe_1_7_6_add_79_carry_2_,
         npu_inst_pe_1_7_6_add_79_carry_1_, npu_inst_pe_1_7_6_n97,
         npu_inst_pe_1_7_6_n96, npu_inst_pe_1_7_6_n95, npu_inst_pe_1_7_6_n94,
         npu_inst_pe_1_7_6_n93, npu_inst_pe_1_7_6_n92, npu_inst_pe_1_7_6_n91,
         npu_inst_pe_1_7_6_n90, npu_inst_pe_1_7_6_n89, npu_inst_pe_1_7_6_n88,
         npu_inst_pe_1_7_6_n87, npu_inst_pe_1_7_6_n86, npu_inst_pe_1_7_6_n85,
         npu_inst_pe_1_7_6_n84, npu_inst_pe_1_7_6_n83, npu_inst_pe_1_7_6_n82,
         npu_inst_pe_1_7_6_n81, npu_inst_pe_1_7_6_n80, npu_inst_pe_1_7_6_n79,
         npu_inst_pe_1_7_6_n78, npu_inst_pe_1_7_6_n77, npu_inst_pe_1_7_6_n76,
         npu_inst_pe_1_7_6_n75, npu_inst_pe_1_7_6_n74, npu_inst_pe_1_7_6_n73,
         npu_inst_pe_1_7_6_n72, npu_inst_pe_1_7_6_n71, npu_inst_pe_1_7_6_n70,
         npu_inst_pe_1_7_6_n69, npu_inst_pe_1_7_6_n68, npu_inst_pe_1_7_6_n67,
         npu_inst_pe_1_7_6_n66, npu_inst_pe_1_7_6_n65, npu_inst_pe_1_7_6_n64,
         npu_inst_pe_1_7_6_n63, npu_inst_pe_1_7_6_n62, npu_inst_pe_1_7_6_n61,
         npu_inst_pe_1_7_6_n60, npu_inst_pe_1_7_6_n59, npu_inst_pe_1_7_6_n58,
         npu_inst_pe_1_7_6_n57, npu_inst_pe_1_7_6_n56, npu_inst_pe_1_7_6_n55,
         npu_inst_pe_1_7_6_n54, npu_inst_pe_1_7_6_n53, npu_inst_pe_1_7_6_n52,
         npu_inst_pe_1_7_6_n51, npu_inst_pe_1_7_6_n50, npu_inst_pe_1_7_6_n49,
         npu_inst_pe_1_7_6_n48, npu_inst_pe_1_7_6_n47, npu_inst_pe_1_7_6_n46,
         npu_inst_pe_1_7_6_n45, npu_inst_pe_1_7_6_n44, npu_inst_pe_1_7_6_n43,
         npu_inst_pe_1_7_6_n42, npu_inst_pe_1_7_6_n41, npu_inst_pe_1_7_6_n40,
         npu_inst_pe_1_7_6_n39, npu_inst_pe_1_7_6_n38, npu_inst_pe_1_7_6_n37,
         npu_inst_pe_1_7_6_n27, npu_inst_pe_1_7_6_n26,
         npu_inst_pe_1_7_6_net2873, npu_inst_pe_1_7_6_net2867,
         npu_inst_pe_1_7_6_N94, npu_inst_pe_1_7_6_N93, npu_inst_pe_1_7_6_N84,
         npu_inst_pe_1_7_6_N80, npu_inst_pe_1_7_6_N79, npu_inst_pe_1_7_6_N78,
         npu_inst_pe_1_7_6_N77, npu_inst_pe_1_7_6_N76, npu_inst_pe_1_7_6_N75,
         npu_inst_pe_1_7_6_N74, npu_inst_pe_1_7_6_N73, npu_inst_pe_1_7_6_N72,
         npu_inst_pe_1_7_6_N71, npu_inst_pe_1_7_6_N70, npu_inst_pe_1_7_6_N69,
         npu_inst_pe_1_7_6_N68, npu_inst_pe_1_7_6_N67, npu_inst_pe_1_7_6_N66,
         npu_inst_pe_1_7_6_N65, npu_inst_pe_1_7_6_int_q_acc_0_,
         npu_inst_pe_1_7_6_int_q_acc_1_, npu_inst_pe_1_7_6_int_q_acc_2_,
         npu_inst_pe_1_7_6_int_q_acc_3_, npu_inst_pe_1_7_6_int_q_acc_4_,
         npu_inst_pe_1_7_6_int_q_acc_5_, npu_inst_pe_1_7_6_int_q_acc_6_,
         npu_inst_pe_1_7_6_int_q_acc_7_, npu_inst_pe_1_7_6_int_data_0_,
         npu_inst_pe_1_7_6_int_data_1_, npu_inst_pe_1_7_6_int_q_weight_0_,
         npu_inst_pe_1_7_6_int_q_weight_1_,
         npu_inst_pe_1_7_6_int_q_reg_v_5__0_,
         npu_inst_pe_1_7_6_int_q_reg_v_5__1_,
         npu_inst_pe_1_7_6_int_q_reg_v_4__0_,
         npu_inst_pe_1_7_6_int_q_reg_v_4__1_,
         npu_inst_pe_1_7_6_int_q_reg_v_3__0_,
         npu_inst_pe_1_7_6_int_q_reg_v_3__1_,
         npu_inst_pe_1_7_6_int_q_reg_v_2__0_,
         npu_inst_pe_1_7_6_int_q_reg_v_2__1_,
         npu_inst_pe_1_7_6_int_q_reg_v_1__0_,
         npu_inst_pe_1_7_6_int_q_reg_v_1__1_,
         npu_inst_pe_1_7_6_int_q_reg_v_0__0_,
         npu_inst_pe_1_7_6_int_q_reg_v_0__1_,
         npu_inst_pe_1_7_6_int_q_reg_h_5__0_,
         npu_inst_pe_1_7_6_int_q_reg_h_5__1_,
         npu_inst_pe_1_7_6_int_q_reg_h_4__0_,
         npu_inst_pe_1_7_6_int_q_reg_h_4__1_,
         npu_inst_pe_1_7_6_int_q_reg_h_3__0_,
         npu_inst_pe_1_7_6_int_q_reg_h_3__1_,
         npu_inst_pe_1_7_6_int_q_reg_h_2__0_,
         npu_inst_pe_1_7_6_int_q_reg_h_2__1_,
         npu_inst_pe_1_7_6_int_q_reg_h_1__0_,
         npu_inst_pe_1_7_6_int_q_reg_h_1__1_,
         npu_inst_pe_1_7_6_int_q_reg_h_0__0_,
         npu_inst_pe_1_7_6_int_q_reg_h_0__1_, npu_inst_pe_1_7_7_n119,
         npu_inst_pe_1_7_7_n118, npu_inst_pe_1_7_7_n117,
         npu_inst_pe_1_7_7_n116, npu_inst_pe_1_7_7_n115,
         npu_inst_pe_1_7_7_n114, npu_inst_pe_1_7_7_n113,
         npu_inst_pe_1_7_7_n112, npu_inst_pe_1_7_7_n111,
         npu_inst_pe_1_7_7_n110, npu_inst_pe_1_7_7_n109,
         npu_inst_pe_1_7_7_n108, npu_inst_pe_1_7_7_n107,
         npu_inst_pe_1_7_7_n106, npu_inst_pe_1_7_7_n105,
         npu_inst_pe_1_7_7_n104, npu_inst_pe_1_7_7_n103,
         npu_inst_pe_1_7_7_n102, npu_inst_pe_1_7_7_n101,
         npu_inst_pe_1_7_7_n100, npu_inst_pe_1_7_7_n99, npu_inst_pe_1_7_7_n98,
         npu_inst_pe_1_7_7_n36, npu_inst_pe_1_7_7_n35, npu_inst_pe_1_7_7_n34,
         npu_inst_pe_1_7_7_n33, npu_inst_pe_1_7_7_n32, npu_inst_pe_1_7_7_n31,
         npu_inst_pe_1_7_7_n30, npu_inst_pe_1_7_7_n29, npu_inst_pe_1_7_7_n28,
         npu_inst_pe_1_7_7_n25, npu_inst_pe_1_7_7_n24, npu_inst_pe_1_7_7_n23,
         npu_inst_pe_1_7_7_n22, npu_inst_pe_1_7_7_n21, npu_inst_pe_1_7_7_n20,
         npu_inst_pe_1_7_7_n19, npu_inst_pe_1_7_7_n18, npu_inst_pe_1_7_7_n17,
         npu_inst_pe_1_7_7_n16, npu_inst_pe_1_7_7_n15, npu_inst_pe_1_7_7_n14,
         npu_inst_pe_1_7_7_n13, npu_inst_pe_1_7_7_n12, npu_inst_pe_1_7_7_n11,
         npu_inst_pe_1_7_7_n10, npu_inst_pe_1_7_7_n9, npu_inst_pe_1_7_7_n8,
         npu_inst_pe_1_7_7_n7, npu_inst_pe_1_7_7_n6, npu_inst_pe_1_7_7_n5,
         npu_inst_pe_1_7_7_n4, npu_inst_pe_1_7_7_n3, npu_inst_pe_1_7_7_n2,
         npu_inst_pe_1_7_7_n1, npu_inst_pe_1_7_7_sub_77_carry_7_,
         npu_inst_pe_1_7_7_sub_77_carry_6_, npu_inst_pe_1_7_7_sub_77_carry_5_,
         npu_inst_pe_1_7_7_sub_77_carry_4_, npu_inst_pe_1_7_7_sub_77_carry_3_,
         npu_inst_pe_1_7_7_sub_77_carry_2_, npu_inst_pe_1_7_7_sub_77_carry_1_,
         npu_inst_pe_1_7_7_add_79_carry_7_, npu_inst_pe_1_7_7_add_79_carry_6_,
         npu_inst_pe_1_7_7_add_79_carry_5_, npu_inst_pe_1_7_7_add_79_carry_4_,
         npu_inst_pe_1_7_7_add_79_carry_3_, npu_inst_pe_1_7_7_add_79_carry_2_,
         npu_inst_pe_1_7_7_add_79_carry_1_, npu_inst_pe_1_7_7_n97,
         npu_inst_pe_1_7_7_n96, npu_inst_pe_1_7_7_n95, npu_inst_pe_1_7_7_n94,
         npu_inst_pe_1_7_7_n93, npu_inst_pe_1_7_7_n92, npu_inst_pe_1_7_7_n91,
         npu_inst_pe_1_7_7_n90, npu_inst_pe_1_7_7_n89, npu_inst_pe_1_7_7_n88,
         npu_inst_pe_1_7_7_n87, npu_inst_pe_1_7_7_n86, npu_inst_pe_1_7_7_n85,
         npu_inst_pe_1_7_7_n84, npu_inst_pe_1_7_7_n83, npu_inst_pe_1_7_7_n82,
         npu_inst_pe_1_7_7_n81, npu_inst_pe_1_7_7_n80, npu_inst_pe_1_7_7_n79,
         npu_inst_pe_1_7_7_n78, npu_inst_pe_1_7_7_n77, npu_inst_pe_1_7_7_n76,
         npu_inst_pe_1_7_7_n75, npu_inst_pe_1_7_7_n74, npu_inst_pe_1_7_7_n73,
         npu_inst_pe_1_7_7_n72, npu_inst_pe_1_7_7_n71, npu_inst_pe_1_7_7_n70,
         npu_inst_pe_1_7_7_n69, npu_inst_pe_1_7_7_n68, npu_inst_pe_1_7_7_n67,
         npu_inst_pe_1_7_7_n66, npu_inst_pe_1_7_7_n65, npu_inst_pe_1_7_7_n64,
         npu_inst_pe_1_7_7_n63, npu_inst_pe_1_7_7_n62, npu_inst_pe_1_7_7_n61,
         npu_inst_pe_1_7_7_n60, npu_inst_pe_1_7_7_n59, npu_inst_pe_1_7_7_n58,
         npu_inst_pe_1_7_7_n57, npu_inst_pe_1_7_7_n56, npu_inst_pe_1_7_7_n55,
         npu_inst_pe_1_7_7_n54, npu_inst_pe_1_7_7_n53, npu_inst_pe_1_7_7_n52,
         npu_inst_pe_1_7_7_n51, npu_inst_pe_1_7_7_n50, npu_inst_pe_1_7_7_n49,
         npu_inst_pe_1_7_7_n48, npu_inst_pe_1_7_7_n47, npu_inst_pe_1_7_7_n46,
         npu_inst_pe_1_7_7_n45, npu_inst_pe_1_7_7_n44, npu_inst_pe_1_7_7_n43,
         npu_inst_pe_1_7_7_n42, npu_inst_pe_1_7_7_n41, npu_inst_pe_1_7_7_n40,
         npu_inst_pe_1_7_7_n39, npu_inst_pe_1_7_7_n38, npu_inst_pe_1_7_7_n37,
         npu_inst_pe_1_7_7_n27, npu_inst_pe_1_7_7_n26,
         npu_inst_pe_1_7_7_net2850, npu_inst_pe_1_7_7_net2844,
         npu_inst_pe_1_7_7_N94, npu_inst_pe_1_7_7_N93, npu_inst_pe_1_7_7_N84,
         npu_inst_pe_1_7_7_N80, npu_inst_pe_1_7_7_N79, npu_inst_pe_1_7_7_N78,
         npu_inst_pe_1_7_7_N77, npu_inst_pe_1_7_7_N76, npu_inst_pe_1_7_7_N75,
         npu_inst_pe_1_7_7_N74, npu_inst_pe_1_7_7_N73, npu_inst_pe_1_7_7_N72,
         npu_inst_pe_1_7_7_N71, npu_inst_pe_1_7_7_N70, npu_inst_pe_1_7_7_N69,
         npu_inst_pe_1_7_7_N68, npu_inst_pe_1_7_7_N67, npu_inst_pe_1_7_7_N66,
         npu_inst_pe_1_7_7_N65, npu_inst_pe_1_7_7_int_q_acc_0_,
         npu_inst_pe_1_7_7_int_q_acc_1_, npu_inst_pe_1_7_7_int_q_acc_2_,
         npu_inst_pe_1_7_7_int_q_acc_3_, npu_inst_pe_1_7_7_int_q_acc_4_,
         npu_inst_pe_1_7_7_int_q_acc_5_, npu_inst_pe_1_7_7_int_q_acc_6_,
         npu_inst_pe_1_7_7_int_q_acc_7_, npu_inst_pe_1_7_7_int_data_0_,
         npu_inst_pe_1_7_7_int_data_1_, npu_inst_pe_1_7_7_int_q_weight_0_,
         npu_inst_pe_1_7_7_int_q_weight_1_,
         npu_inst_pe_1_7_7_int_q_reg_v_5__0_,
         npu_inst_pe_1_7_7_int_q_reg_v_5__1_,
         npu_inst_pe_1_7_7_int_q_reg_v_4__0_,
         npu_inst_pe_1_7_7_int_q_reg_v_4__1_,
         npu_inst_pe_1_7_7_int_q_reg_v_3__0_,
         npu_inst_pe_1_7_7_int_q_reg_v_3__1_,
         npu_inst_pe_1_7_7_int_q_reg_v_2__0_,
         npu_inst_pe_1_7_7_int_q_reg_v_2__1_,
         npu_inst_pe_1_7_7_int_q_reg_v_1__0_,
         npu_inst_pe_1_7_7_int_q_reg_v_1__1_,
         npu_inst_pe_1_7_7_int_q_reg_v_0__0_,
         npu_inst_pe_1_7_7_int_q_reg_v_0__1_,
         npu_inst_pe_1_7_7_int_q_reg_h_5__0_,
         npu_inst_pe_1_7_7_int_q_reg_h_5__1_,
         npu_inst_pe_1_7_7_int_q_reg_h_4__0_,
         npu_inst_pe_1_7_7_int_q_reg_h_4__1_,
         npu_inst_pe_1_7_7_int_q_reg_h_3__0_,
         npu_inst_pe_1_7_7_int_q_reg_h_3__1_,
         npu_inst_pe_1_7_7_int_q_reg_h_2__0_,
         npu_inst_pe_1_7_7_int_q_reg_h_2__1_,
         npu_inst_pe_1_7_7_int_q_reg_h_1__0_,
         npu_inst_pe_1_7_7_int_q_reg_h_1__1_,
         npu_inst_pe_1_7_7_int_q_reg_h_0__0_,
         npu_inst_pe_1_7_7_int_q_reg_h_0__1_, ckg_ctrl8b_inst_n11,
         ckg_ctrl8b_inst_n10, ckg_ctrl8b_inst_n9, ckg_ctrl8b_inst_n8,
         ckg_ctrl8b_inst_n5, ckg_ctrl8b_inst_n4, ckg_ctrl8b_inst_n3,
         ckg_ctrl8b_inst_n2, ckg_ctrl8b_inst_n1, ckg_ctrl8b_inst_n20,
         ckg_ctrl8b_inst_n19, ckg_ctrl8b_inst_n18, ckg_ctrl8b_inst_n17,
         ckg_ctrl8b_inst_n16, ckg_ctrl8b_inst_n15, ckg_ctrl8b_inst_n14,
         ckg_ctrl8b_inst_n13, ckg_ctrl8b_inst_n12, hmode_cnt_inst_n12,
         hmode_cnt_inst_n6, hmode_cnt_inst_n4, hmode_cnt_inst_n2,
         hmode_cnt_inst_n1, hmode_cnt_inst_n11, hmode_cnt_inst_n10,
         hmode_cnt_inst_n9, hmode_cnt_inst_n8, hmode_cnt_inst_n7,
         hmode_cnt_inst_n5, hmode_cnt_inst_net2826, hmode_cnt_inst_N12,
         hmode_cnt_inst_N10, hmode_cnt_inst_q_2_, vmode_cnt_inst_n12,
         vmode_cnt_inst_n6, vmode_cnt_inst_n4, vmode_cnt_inst_n2,
         vmode_cnt_inst_n1, vmode_cnt_inst_n11, vmode_cnt_inst_n10,
         vmode_cnt_inst_n9, vmode_cnt_inst_n8, vmode_cnt_inst_n7,
         vmode_cnt_inst_n5, vmode_cnt_inst_net2808, vmode_cnt_inst_N12,
         vmode_cnt_inst_N10, vmode_cnt_inst_q_0_, vmode_cnt_inst_q_1_,
         vmode_cnt_inst_q_2_, res_cnt_inst_n2, res_cnt_inst_n1,
         res_cnt_inst_n14, res_cnt_inst_n13, res_cnt_inst_n12,
         res_cnt_inst_n11, res_cnt_inst_n10, res_cnt_inst_n9, res_cnt_inst_n8,
         res_cnt_inst_n7, res_cnt_inst_n5, res_cnt_inst_net2790,
         res_cnt_inst_N12, res_cnt_inst_N10, res_cnt_inst_q_0_,
         res_cnt_inst_q_1_, res_cnt_inst_q_2_, ifmaps_cnt_inst_n12,
         ifmaps_cnt_inst_n6, ifmaps_cnt_inst_n4, ifmaps_cnt_inst_n2,
         ifmaps_cnt_inst_n1, ifmaps_cnt_inst_n11, ifmaps_cnt_inst_n10,
         ifmaps_cnt_inst_n9, ifmaps_cnt_inst_n8, ifmaps_cnt_inst_n7,
         ifmaps_cnt_inst_n5, ifmaps_cnt_inst_net2772, ifmaps_cnt_inst_N12,
         ifmaps_cnt_inst_N10, npu_cnt_inst_n12, npu_cnt_inst_n6,
         npu_cnt_inst_n4, npu_cnt_inst_n2, npu_cnt_inst_n1, npu_cnt_inst_n11,
         npu_cnt_inst_n10, npu_cnt_inst_n9, npu_cnt_inst_n8, npu_cnt_inst_n7,
         npu_cnt_inst_n5, npu_cnt_inst_net2754, npu_cnt_inst_N12,
         npu_cnt_inst_N10, tilev_cnt_inst_n8, tilev_cnt_inst_n6,
         tilev_cnt_inst_n3, tilev_cnt_inst_n2, tilev_cnt_inst_n1,
         tilev_cnt_inst_n17, tilev_cnt_inst_n15, tilev_cnt_inst_n14,
         tilev_cnt_inst_n13, tilev_cnt_inst_n12, tilev_cnt_inst_n11,
         tilev_cnt_inst_n9, tilev_cnt_inst_n7, tilev_cnt_inst_n5,
         tilev_cnt_inst_n4, tilev_cnt_inst_q_0_, tilev_cnt_inst_q_1_,
         tileh_cnt_inst_n24, tileh_cnt_inst_n23, tileh_cnt_inst_n22,
         tileh_cnt_inst_n21, tileh_cnt_inst_n20, tileh_cnt_inst_n19,
         tileh_cnt_inst_n18, tileh_cnt_inst_n17, tileh_cnt_inst_n16,
         tileh_cnt_inst_n10, tileh_cnt_inst_n8, tileh_cnt_inst_n6,
         tileh_cnt_inst_n3, tileh_cnt_inst_n2, tileh_cnt_inst_n1,
         tileh_cnt_inst_q_1_, ofmaps_cnt_inst_n4, ofmaps_cnt_inst_n2,
         ofmaps_cnt_inst_n1, ofmaps_cnt_inst_n19, ofmaps_cnt_inst_n18,
         ofmaps_cnt_inst_n17, ofmaps_cnt_inst_n16, ofmaps_cnt_inst_n15,
         ofmaps_cnt_inst_n14, ofmaps_cnt_inst_n13, ofmaps_cnt_inst_n12,
         ofmaps_cnt_inst_n11, ofmaps_cnt_inst_n10, ofmaps_cnt_inst_n9,
         ofmaps_cnt_inst_n8, ofmaps_cnt_inst_n5, ofmaps_cnt_inst_net2736,
         ofmaps_cnt_inst_N14, ofmaps_cnt_inst_N13, ofmaps_cnt_inst_N11,
         ofmaps_cnt_inst_q_0_, ofmaps_cnt_inst_q_1_, ofmaps_cnt_inst_q_2_,
         ofmaps_cnt_inst_q_3_, i_data_addr_gen_inst_n27,
         i_data_addr_gen_inst_n26, i_data_addr_gen_inst_n25,
         i_data_addr_gen_inst_n24, i_data_addr_gen_inst_n23,
         i_data_addr_gen_inst_n31, i_data_addr_gen_inst_n30,
         i_data_addr_gen_inst_n29, i_data_addr_gen_inst_net2719,
         i_data_addr_gen_inst_net2714, i_data_addr_gen_inst_net2708,
         i_data_addr_gen_inst_N77, i_data_addr_gen_inst_N76,
         i_data_addr_gen_inst_N75, i_data_addr_gen_inst_N74,
         i_data_addr_gen_inst_N73, i_data_addr_gen_inst_N72,
         i_data_addr_gen_inst_N71, i_data_addr_gen_inst_N70,
         i_data_addr_gen_inst_N69, i_data_addr_gen_inst_N68,
         i_data_addr_gen_inst_N67, i_data_addr_gen_inst_N66,
         i_data_addr_gen_inst_N65, i_data_addr_gen_inst_N64,
         i_data_addr_gen_inst_N63, i_data_addr_gen_inst_N62,
         i_data_addr_gen_inst_N61, i_data_addr_gen_inst_N60,
         i_data_addr_gen_inst_N59, i_data_addr_gen_inst_N58,
         i_data_addr_gen_inst_N39, i_data_addr_gen_inst_N38,
         i_data_addr_gen_inst_N37, i_data_addr_gen_inst_N36,
         i_data_addr_gen_inst_N35, i_data_addr_gen_inst_N34,
         i_data_addr_gen_inst_N33, i_data_addr_gen_inst_N32,
         i_data_addr_gen_inst_N31, i_data_addr_gen_inst_N30,
         i_data_addr_gen_inst_N17, i_data_addr_gen_inst_N16,
         i_data_addr_gen_inst_N15, i_data_addr_gen_inst_N14,
         i_data_addr_gen_inst_N13, i_data_addr_gen_inst_N12,
         i_data_addr_gen_inst_N11, i_data_addr_gen_inst_N10,
         i_data_addr_gen_inst_N9, i_data_addr_gen_inst_N8,
         i_data_addr_gen_inst_int_data_offs_addr_0_,
         i_data_addr_gen_inst_int_data_offs_addr_1_,
         i_data_addr_gen_inst_int_data_offs_addr_2_,
         i_data_addr_gen_inst_int_data_offs_addr_3_,
         i_data_addr_gen_inst_int_data_offs_addr_4_,
         i_data_addr_gen_inst_int_data_offs_addr_5_,
         i_data_addr_gen_inst_int_data_offs_addr_6_,
         i_data_addr_gen_inst_int_data_offs_addr_7_,
         i_data_addr_gen_inst_int_data_offs_addr_8_,
         i_data_addr_gen_inst_int_data_offs_addr_9_,
         i_data_addr_gen_inst_add_33_n1, i_data_addr_gen_inst_add_32_n1,
         i_weight_addr_gen_inst_n38, i_weight_addr_gen_inst_n37,
         i_weight_addr_gen_inst_n36, i_weight_addr_gen_inst_n35,
         i_weight_addr_gen_inst_n34, i_weight_addr_gen_inst_net2691,
         i_weight_addr_gen_inst_net2685, i_weight_addr_gen_inst_N38,
         i_weight_addr_gen_inst_N37, i_weight_addr_gen_inst_N36,
         i_weight_addr_gen_inst_N35, i_weight_addr_gen_inst_N34,
         i_weight_addr_gen_inst_N33, i_weight_addr_gen_inst_N32,
         i_weight_addr_gen_inst_N31, i_weight_addr_gen_inst_N30,
         i_weight_addr_gen_inst_N29, i_weight_addr_gen_inst_N28,
         i_weight_addr_gen_inst_N27, i_weight_addr_gen_inst_N26,
         i_weight_addr_gen_inst_N25, i_weight_addr_gen_inst_N24,
         i_weight_addr_gen_inst_N23, i_weight_addr_gen_inst_N22,
         i_weight_addr_gen_inst_N21, i_weight_addr_gen_inst_N20,
         i_weight_addr_gen_inst_N19, i_weight_addr_gen_inst_N18,
         i_weight_addr_gen_inst_N17, i_weight_addr_gen_inst_N16,
         i_weight_addr_gen_inst_N15, i_weight_addr_gen_inst_N14,
         i_weight_addr_gen_inst_N13, i_weight_addr_gen_inst_N12,
         i_weight_addr_gen_inst_N11, i_weight_addr_gen_inst_N10,
         i_weight_addr_gen_inst_N9, i_weight_addr_gen_inst_N8,
         i_weight_addr_gen_inst_N7, i_weight_addr_gen_inst_N6,
         i_weight_addr_gen_inst_int_offs_addr_0_,
         i_weight_addr_gen_inst_int_offs_addr_1_,
         i_weight_addr_gen_inst_int_offs_addr_2_,
         i_weight_addr_gen_inst_int_offs_addr_3_,
         i_weight_addr_gen_inst_int_offs_addr_4_,
         i_weight_addr_gen_inst_int_offs_addr_5_,
         i_weight_addr_gen_inst_int_offs_addr_6_,
         i_weight_addr_gen_inst_int_offs_addr_7_,
         i_weight_addr_gen_inst_int_offs_addr_8_,
         i_weight_addr_gen_inst_int_offs_addr_9_,
         i_weight_addr_gen_inst_int_offs_addr_10_,
         i_weight_addr_gen_inst_int_offs_addr_11_,
         i_weight_addr_gen_inst_int_offs_addr_12_,
         i_weight_addr_gen_inst_int_offs_addr_13_,
         i_weight_addr_gen_inst_int_offs_addr_14_,
         i_weight_addr_gen_inst_int_offs_addr_15_,
         i_weight_addr_gen_inst_int_offs_addr_16_,
         i_weight_addr_gen_inst_int_offs_addr_17_,
         i_weight_addr_gen_inst_int_offs_addr_18_,
         i_weight_addr_gen_inst_int_offs_addr_19_,
         i_weight_addr_gen_inst_int_offs_addr_20_,
         i_weight_addr_gen_inst_int_offs_addr_21_,
         i_weight_addr_gen_inst_int_offs_addr_22_,
         i_weight_addr_gen_inst_int_offs_addr_23_,
         i_weight_addr_gen_inst_int_offs_addr_24_,
         i_weight_addr_gen_inst_int_offs_addr_25_,
         i_weight_addr_gen_inst_int_offs_addr_26_,
         i_weight_addr_gen_inst_int_offs_addr_27_,
         i_weight_addr_gen_inst_int_offs_addr_28_,
         i_weight_addr_gen_inst_int_offs_addr_29_,
         i_weight_addr_gen_inst_int_offs_addr_30_,
         i_weight_addr_gen_inst_int_offs_addr_31_,
         i_weight_addr_gen_inst_add_26_n1;
  wire   [2:0] int_npu_ptr;
  wire   [2:0] int_ifmaps_ptr;
  wire   [2:0] ps_int_ifmaps_ptr;
  wire   [7:0] int_i_data_if1;
  wire   [7:0] int_i_data_if2;
  wire   [7:0] int_i_data_if3;
  wire   [7:0] int_i_data_if4;
  wire   [7:0] int_i_data_if5;
  wire   [7:0] int_i_data_if6;
  wire   [7:0] int_i_data_if7;
  wire   [7:0] int_i_data_if8;
  wire   [1:0] ps_int_hmode_cnt;
  wire   [1:0] int_hmode_cnt;
  wire   [1:0] int_i_data_h_npu1;
  wire   [1:0] int_i_data_h_npu2;
  wire   [1:0] int_i_data_h_npu3;
  wire   [1:0] int_i_data_h_npu4;
  wire   [1:0] int_i_data_h_npu5;
  wire   [1:0] int_i_data_h_npu6;
  wire   [1:0] int_i_data_h_npu7;
  wire   [1:0] int_i_data_h_npu8;
  wire   [15:0] int_i_data_v_npu;
  wire   [0:7] int_ckg_rmask;
  wire   [0:7] int_ckg_cmask;
  wire   [2:0] int_arv_res;
  wire   [2:0] int_d_tc;
  wire   [47:0] act_buffer_inst_int_data8;
  wire   [47:0] act_buffer_inst_int_data7;
  wire   [47:0] act_buffer_inst_int_data6;
  wire   [47:0] act_buffer_inst_int_data5;
  wire   [47:0] act_buffer_inst_int_data4;
  wire   [47:0] act_buffer_inst_int_data3;
  wire   [47:0] act_buffer_inst_int_data2;
  wire   [47:0] act_buffer_inst_int_data1;
  wire   [7:0] act_if_inst_int_data8;
  wire   [7:0] act_if_inst_int_data7;
  wire   [7:0] act_if_inst_int_data6;
  wire   [7:0] act_if_inst_int_data5;
  wire   [7:0] act_if_inst_int_data4;
  wire   [7:0] act_if_inst_int_data3;
  wire   [7:0] act_if_inst_int_data2;
  wire   [7:0] act_if_inst_int_data1;
  wire   [63:0] npu_inst_int_ckg;
  wire   [9:0] i_data_addr_gen_inst_int_data_odd_base_addr;
  wire   [9:0] i_data_addr_gen_inst_int_data_even_base_addr;
  wire   [9:2] i_data_addr_gen_inst_add_78_carry;
  wire   [9:2] i_data_addr_gen_inst_add_62_carry;
  wire   [9:2] i_data_addr_gen_inst_add_46_carry;
  wire   [9:2] i_data_addr_gen_inst_add_33_carry;
  wire   [9:2] i_data_addr_gen_inst_add_32_carry;
  wire   [31:0] i_weight_addr_gen_inst_int_base_addr;
  wire   [31:2] i_weight_addr_gen_inst_add_49_carry;
  wire   [31:2] i_weight_addr_gen_inst_add_26_carry;
  wire   [9:2] add_428_carry;
  wire   [9:2] add_426_carry;

  DFFR_X1 int_q_tc_reg_2_ ( .D(int_d_tc[2]), .CK(net2658), .RN(n13), .Q(
        s_tc_tilev) );
  DFFR_X1 int_q_tc_reg_0_ ( .D(int_d_tc[0]), .CK(net2658), .RN(n13), .Q(
        s_tc_ofmaps) );
  DFFR_X1 int_o_data_ev_odd_n_reg ( .D(i_data_ev_odd_n), .CK(net2658), .RN(n13), .Q(o_data_ev_odd_n), .QN(n8) );
  DFFR_X1 int_o_data_odd_addr_reg_8_ ( .D(N15), .CK(net2663), .RN(n12), .Q(
        o_data_odd_addr[8]) );
  DFFR_X1 int_o_data_odd_addr_reg_9_ ( .D(N16), .CK(net2663), .RN(n12), .Q(
        o_data_odd_addr[9]) );
  DFFR_X1 int_o_data_even_addr_reg_8_ ( .D(N25), .CK(net2668), .RN(n12), .Q(
        o_data_even_addr[8]) );
  DFFR_X1 int_o_data_even_addr_reg_9_ ( .D(N26), .CK(net2668), .RN(n12), .Q(
        o_data_even_addr[9]) );
  DFFR_X1 ps_int_hmode_cnt_reg_1_ ( .D(int_hmode_cnt[1]), .CK(ck), .RN(n14), 
        .Q(ps_int_hmode_cnt[1]) );
  DFFR_X1 ps_int_s_tc_tileh_reg ( .D(s_tc_tileh), .CK(ck), .RN(n14), .Q(
        ps_int_s_tc_tileh) );
  DFFR_X1 ps_int_s_tc_tilev_reg ( .D(s_tc_tilev), .CK(ck), .RN(n14), .Q(
        ps_int_s_tc_tilev) );
  DFFR_X1 ps_int_ifmaps_ptr_reg_1_ ( .D(int_ifmaps_ptr[1]), .CK(ck), .RN(n14), 
        .Q(ps_int_ifmaps_ptr[1]) );
  DFFR_X1 ps_int_hmode_cnt_reg_0_ ( .D(int_hmode_cnt[0]), .CK(ck), .RN(n14), 
        .Q(ps_int_hmode_cnt[0]) );
  DFFR_X1 ps_int_ifmaps_ptr_reg_2_ ( .D(int_ifmaps_ptr[2]), .CK(ck), .RN(n14), 
        .Q(ps_int_ifmaps_ptr[2]) );
  DFFR_X1 int_o_data_odd_addr_reg_0_ ( .D(N7), .CK(net2663), .RN(n14), .Q(
        o_data_odd_addr[0]) );
  DFFR_X1 int_o_data_even_addr_reg_0_ ( .D(N17), .CK(net2668), .RN(n14), .Q(
        o_data_even_addr[0]) );
  DFFR_X1 ps_int_ifmaps_ptr_reg_0_ ( .D(int_ifmaps_ptr[0]), .CK(ck), .RN(n14), 
        .Q(ps_int_ifmaps_ptr[0]) );
  DFFR_X1 int_o_data_odd_addr_reg_1_ ( .D(N8), .CK(net2663), .RN(n14), .Q(
        o_data_odd_addr[1]) );
  DFFR_X1 int_o_data_even_addr_reg_1_ ( .D(N18), .CK(net2668), .RN(n14), .Q(
        o_data_even_addr[1]) );
  DFFR_X1 int_o_data_odd_addr_reg_2_ ( .D(N9), .CK(net2663), .RN(n14), .Q(
        o_data_odd_addr[2]) );
  DFFR_X1 int_o_data_even_addr_reg_2_ ( .D(N19), .CK(net2668), .RN(n14), .Q(
        o_data_even_addr[2]) );
  DFFR_X1 int_o_data_odd_addr_reg_3_ ( .D(N10), .CK(net2663), .RN(n14), .Q(
        o_data_odd_addr[3]) );
  DFFR_X1 int_o_data_even_addr_reg_3_ ( .D(N20), .CK(net2668), .RN(n14), .Q(
        o_data_even_addr[3]) );
  DFFR_X1 int_o_data_odd_addr_reg_4_ ( .D(N11), .CK(net2663), .RN(n14), .Q(
        o_data_odd_addr[4]) );
  DFFR_X1 int_o_data_even_addr_reg_4_ ( .D(N21), .CK(net2668), .RN(n14), .Q(
        o_data_even_addr[4]) );
  DFFR_X1 int_o_data_odd_addr_reg_5_ ( .D(N12), .CK(net2663), .RN(n14), .Q(
        o_data_odd_addr[5]) );
  DFFR_X1 int_o_data_even_addr_reg_5_ ( .D(N22), .CK(net2668), .RN(n14), .Q(
        o_data_even_addr[5]) );
  DFFR_X1 int_i_data_v_npu_reg_15_ ( .D(i_actv[15]), .CK(net2652), .RN(n13), 
        .Q(int_i_data_v_npu[15]) );
  DFFR_X1 int_i_data_v_npu_reg_14_ ( .D(i_actv[14]), .CK(net2652), .RN(n12), 
        .Q(int_i_data_v_npu[14]) );
  DFFR_X1 int_i_data_v_npu_reg_13_ ( .D(i_actv[13]), .CK(net2652), .RN(n13), 
        .Q(int_i_data_v_npu[13]) );
  DFFR_X1 int_i_data_v_npu_reg_12_ ( .D(i_actv[12]), .CK(net2652), .RN(n12), 
        .Q(int_i_data_v_npu[12]) );
  DFFR_X1 int_i_data_v_npu_reg_11_ ( .D(i_actv[11]), .CK(net2652), .RN(n13), 
        .Q(int_i_data_v_npu[11]) );
  DFFR_X1 int_i_data_v_npu_reg_10_ ( .D(i_actv[10]), .CK(net2652), .RN(n12), 
        .Q(int_i_data_v_npu[10]) );
  DFFR_X1 int_i_data_v_npu_reg_9_ ( .D(i_actv[9]), .CK(net2652), .RN(n13), .Q(
        int_i_data_v_npu[9]) );
  DFFR_X1 int_i_data_v_npu_reg_8_ ( .D(i_actv[8]), .CK(net2652), .RN(n12), .Q(
        int_i_data_v_npu[8]) );
  DFFR_X1 int_i_data_v_npu_reg_7_ ( .D(i_actv[7]), .CK(net2652), .RN(n13), .Q(
        int_i_data_v_npu[7]) );
  DFFR_X1 int_i_data_v_npu_reg_6_ ( .D(i_actv[6]), .CK(net2652), .RN(n12), .Q(
        int_i_data_v_npu[6]) );
  DFFR_X1 int_i_data_v_npu_reg_5_ ( .D(i_actv[5]), .CK(net2652), .RN(n13), .Q(
        int_i_data_v_npu[5]) );
  DFFR_X1 int_i_data_v_npu_reg_4_ ( .D(i_actv[4]), .CK(net2652), .RN(n12), .Q(
        int_i_data_v_npu[4]) );
  DFFR_X1 int_i_data_v_npu_reg_3_ ( .D(i_actv[3]), .CK(net2652), .RN(n13), .Q(
        int_i_data_v_npu[3]) );
  DFFR_X1 int_i_data_v_npu_reg_2_ ( .D(i_actv[2]), .CK(net2652), .RN(n12), .Q(
        int_i_data_v_npu[2]) );
  DFFR_X1 int_i_data_v_npu_reg_1_ ( .D(i_actv[1]), .CK(net2652), .RN(n14), .Q(
        int_i_data_v_npu[1]) );
  DFFR_X1 int_i_data_v_npu_reg_0_ ( .D(i_actv[0]), .CK(net2652), .RN(n14), .Q(
        int_i_data_v_npu[0]) );
  DFFR_X1 int_o_data_odd_addr_reg_6_ ( .D(N13), .CK(net2663), .RN(n14), .Q(
        o_data_odd_addr[6]) );
  DFFR_X1 int_o_data_even_addr_reg_6_ ( .D(N23), .CK(net2668), .RN(n14), .Q(
        o_data_even_addr[6]) );
  DFFR_X1 ps_ctrl_en_npu_reg ( .D(ctrl_en_npu), .CK(ck), .RN(n14), .Q(
        ps_ctrl_en_npu) );
  DFFR_X1 ps_ctrl_wr_pipe_reg ( .D(ctrl_wr_pipe), .CK(ck), .RN(n14), .Q(
        ps_ctrl_wr_pipe) );
  DFFR_X1 ps_ctrl_ldh_v_n_reg ( .D(ctrl_ldh_v_n), .CK(ck), .RN(n14), .Q(
        ps_ctrl_ldh_v_n) );
  DFFR_X1 int_o_data_odd_addr_reg_7_ ( .D(N14), .CK(net2663), .RN(n14), .Q(
        o_data_odd_addr[7]) );
  DFFR_X1 int_o_data_even_addr_reg_7_ ( .D(N24), .CK(net2668), .RN(n14), .Q(
        o_data_even_addr[7]) );
  DFFR_X1 int_q_tc_reg_1_ ( .D(int_d_tc[1]), .CK(net2658), .RN(n14), .Q(
        s_tc_tileh) );
  INV_X2 U19 ( .A(n10), .ZN(n14) );
  CLKBUF_X1 U20 ( .A(rst), .Z(n9) );
  INV_X1 U21 ( .A(n5), .ZN(n15) );
  AND2_X1 U22 ( .A1(s_tc_npu_ptr), .A2(int_en_npu_ptr), .ZN(int_en_tilev_ptr)
         );
  AND2_X1 U23 ( .A1(int_d_tc[1]), .A2(n15), .ZN(int_rst_i_data_addr) );
  NAND2_X1 U24 ( .A1(int_d_tc[2]), .A2(int_en_tilev_ptr), .ZN(n5) );
  NOR2_X1 U25 ( .A1(i_data_ev_odd_n), .A2(n5), .ZN(int_inc_i_data_even) );
  AND2_X1 U26 ( .A1(n15), .A2(i_data_ev_odd_n), .ZN(int_inc_i_data_odd) );
  AND2_X1 U27 ( .A1(s_tc_ifmaps), .A2(ctrl_ldh_v_n), .ZN(int_en_npu_ptr) );
  OR2_X1 U28 ( .A1(s_tc_res), .A2(n7), .ZN(int_en_vmode) );
  AND2_X1 U29 ( .A1(ctrl_en_vmode), .A2(s_tc_ifmaps), .ZN(n7) );
  AND2_X1 U30 ( .A1(n8), .A2(ctrl_wr_pipe), .ZN(N27) );
  AND3_X1 U31 ( .A1(s_tc_tileh), .A2(s_tc_res), .A3(s_tc_tilev), .ZN(
        int_inc_i_w_addr) );
  AND2_X1 U32 ( .A1(ctrl_wr_pipe), .A2(o_data_ev_odd_n), .ZN(N28) );
  AND2_X1 U33 ( .A1(ctrl_en_hmode), .A2(s_tc_ifmaps), .ZN(int_en_hmode) );
  BUF_X1 U34 ( .A(rst), .Z(n10) );
  BUF_X1 U35 ( .A(rst), .Z(n11) );
  INV_X1 U36 ( .A(n11), .ZN(n12) );
  INV_X1 U37 ( .A(n11), .ZN(n13) );
  INV_X1 act_buffer_inst_U309 ( .A(ps_int_ifmaps_ptr[0]), .ZN(
        act_buffer_inst_n189) );
  CLKBUF_X1 act_buffer_inst_U308 ( .A(act_buffer_inst_n12), .Z(
        act_buffer_inst_n188) );
  CLKBUF_X1 act_buffer_inst_U307 ( .A(act_buffer_inst_n13), .Z(
        act_buffer_inst_n182) );
  CLKBUF_X1 act_buffer_inst_U306 ( .A(act_buffer_inst_n14), .Z(
        act_buffer_inst_n176) );
  CLKBUF_X1 act_buffer_inst_U305 ( .A(act_buffer_inst_n15), .Z(
        act_buffer_inst_n170) );
  CLKBUF_X1 act_buffer_inst_U304 ( .A(act_buffer_inst_n16), .Z(
        act_buffer_inst_n164) );
  CLKBUF_X1 act_buffer_inst_U303 ( .A(act_buffer_inst_n17), .Z(
        act_buffer_inst_n9) );
  INV_X1 act_buffer_inst_U302 ( .A(int_npu_ptr[2]), .ZN(act_buffer_inst_n193)
         );
  INV_X1 act_buffer_inst_U301 ( .A(int_npu_ptr[1]), .ZN(act_buffer_inst_n192)
         );
  INV_X1 act_buffer_inst_U300 ( .A(int_npu_ptr[0]), .ZN(act_buffer_inst_n191)
         );
  INV_X1 act_buffer_inst_U299 ( .A(int_ifmaps_ptr[0]), .ZN(
        act_buffer_inst_n194) );
  INV_X1 act_buffer_inst_U298 ( .A(int_ifmaps_ptr[2]), .ZN(
        act_buffer_inst_n196) );
  INV_X1 act_buffer_inst_U297 ( .A(int_ifmaps_ptr[1]), .ZN(
        act_buffer_inst_n195) );
  NAND4_X1 act_buffer_inst_U296 ( .A1(ctrl_ldh_v_n), .A2(act_buffer_inst_n194), 
        .A3(act_buffer_inst_n195), .A4(act_buffer_inst_n196), .ZN(
        act_buffer_inst_n145) );
  NAND4_X1 act_buffer_inst_U295 ( .A1(int_ifmaps_ptr[2]), .A2(ctrl_ldh_v_n), 
        .A3(act_buffer_inst_n194), .A4(act_buffer_inst_n195), .ZN(
        act_buffer_inst_n149) );
  NAND4_X1 act_buffer_inst_U294 ( .A1(int_ifmaps_ptr[1]), .A2(ctrl_ldh_v_n), 
        .A3(act_buffer_inst_n194), .A4(act_buffer_inst_n196), .ZN(
        act_buffer_inst_n147) );
  NAND4_X1 act_buffer_inst_U293 ( .A1(int_ifmaps_ptr[2]), .A2(
        int_ifmaps_ptr[0]), .A3(ctrl_ldh_v_n), .A4(act_buffer_inst_n195), .ZN(
        act_buffer_inst_n150) );
  NAND4_X1 act_buffer_inst_U292 ( .A1(int_ifmaps_ptr[1]), .A2(
        int_ifmaps_ptr[0]), .A3(ctrl_ldh_v_n), .A4(act_buffer_inst_n196), .ZN(
        act_buffer_inst_n148) );
  NAND4_X1 act_buffer_inst_U291 ( .A1(int_ifmaps_ptr[0]), .A2(ctrl_ldh_v_n), 
        .A3(act_buffer_inst_n195), .A4(act_buffer_inst_n196), .ZN(
        act_buffer_inst_n146) );
  AOI222_X1 act_buffer_inst_U290 ( .A1(act_buffer_inst_int_data1[43]), .A2(
        act_buffer_inst_n165), .B1(act_buffer_inst_int_data1[27]), .B2(
        act_buffer_inst_n159), .C1(act_buffer_inst_int_data1[35]), .C2(
        act_buffer_inst_n4), .ZN(act_buffer_inst_n136) );
  AOI222_X1 act_buffer_inst_U289 ( .A1(act_buffer_inst_int_data1[19]), .A2(
        act_buffer_inst_n183), .B1(act_buffer_inst_int_data1[3]), .B2(
        act_buffer_inst_n177), .C1(act_buffer_inst_int_data1[11]), .C2(
        act_buffer_inst_n171), .ZN(act_buffer_inst_n137) );
  NAND2_X1 act_buffer_inst_U288 ( .A1(act_buffer_inst_n136), .A2(
        act_buffer_inst_n137), .ZN(int_i_data_if1[3]) );
  AOI222_X1 act_buffer_inst_U287 ( .A1(act_buffer_inst_int_data2[43]), .A2(
        act_buffer_inst_n165), .B1(act_buffer_inst_int_data2[27]), .B2(
        act_buffer_inst_n159), .C1(act_buffer_inst_int_data2[35]), .C2(
        act_buffer_inst_n4), .ZN(act_buffer_inst_n120) );
  AOI222_X1 act_buffer_inst_U286 ( .A1(act_buffer_inst_int_data2[19]), .A2(
        act_buffer_inst_n183), .B1(act_buffer_inst_int_data2[3]), .B2(
        act_buffer_inst_n177), .C1(act_buffer_inst_int_data2[11]), .C2(
        act_buffer_inst_n171), .ZN(act_buffer_inst_n121) );
  NAND2_X1 act_buffer_inst_U285 ( .A1(act_buffer_inst_n120), .A2(
        act_buffer_inst_n121), .ZN(int_i_data_if2[3]) );
  AOI222_X1 act_buffer_inst_U284 ( .A1(act_buffer_inst_int_data5[19]), .A2(
        act_buffer_inst_n185), .B1(act_buffer_inst_int_data5[3]), .B2(
        act_buffer_inst_n179), .C1(act_buffer_inst_int_data5[11]), .C2(
        act_buffer_inst_n173), .ZN(act_buffer_inst_n73) );
  AOI222_X1 act_buffer_inst_U283 ( .A1(act_buffer_inst_int_data5[43]), .A2(
        act_buffer_inst_n167), .B1(act_buffer_inst_int_data5[27]), .B2(
        act_buffer_inst_n161), .C1(act_buffer_inst_int_data5[35]), .C2(
        act_buffer_inst_n6), .ZN(act_buffer_inst_n72) );
  NAND2_X1 act_buffer_inst_U282 ( .A1(act_buffer_inst_n72), .A2(
        act_buffer_inst_n73), .ZN(int_i_data_if5[3]) );
  AOI222_X1 act_buffer_inst_U281 ( .A1(act_buffer_inst_int_data3[19]), .A2(
        act_buffer_inst_n184), .B1(act_buffer_inst_int_data3[3]), .B2(
        act_buffer_inst_n178), .C1(act_buffer_inst_int_data3[11]), .C2(
        act_buffer_inst_n172), .ZN(act_buffer_inst_n105) );
  AOI222_X1 act_buffer_inst_U280 ( .A1(act_buffer_inst_int_data3[43]), .A2(
        act_buffer_inst_n166), .B1(act_buffer_inst_int_data3[27]), .B2(
        act_buffer_inst_n160), .C1(act_buffer_inst_int_data3[35]), .C2(
        act_buffer_inst_n5), .ZN(act_buffer_inst_n104) );
  NAND2_X1 act_buffer_inst_U279 ( .A1(act_buffer_inst_n104), .A2(
        act_buffer_inst_n105), .ZN(int_i_data_if3[3]) );
  AOI222_X1 act_buffer_inst_U278 ( .A1(act_buffer_inst_int_data4[19]), .A2(
        act_buffer_inst_n185), .B1(act_buffer_inst_int_data4[3]), .B2(
        act_buffer_inst_n179), .C1(act_buffer_inst_int_data4[11]), .C2(
        act_buffer_inst_n173), .ZN(act_buffer_inst_n89) );
  AOI222_X1 act_buffer_inst_U277 ( .A1(act_buffer_inst_int_data4[43]), .A2(
        act_buffer_inst_n167), .B1(act_buffer_inst_int_data4[27]), .B2(
        act_buffer_inst_n161), .C1(act_buffer_inst_int_data4[35]), .C2(
        act_buffer_inst_n6), .ZN(act_buffer_inst_n88) );
  NAND2_X1 act_buffer_inst_U276 ( .A1(act_buffer_inst_n88), .A2(
        act_buffer_inst_n89), .ZN(int_i_data_if4[3]) );
  AOI222_X1 act_buffer_inst_U275 ( .A1(act_buffer_inst_int_data1[45]), .A2(
        act_buffer_inst_n165), .B1(act_buffer_inst_int_data1[29]), .B2(
        act_buffer_inst_n159), .C1(act_buffer_inst_int_data1[37]), .C2(
        act_buffer_inst_n4), .ZN(act_buffer_inst_n132) );
  AOI222_X1 act_buffer_inst_U274 ( .A1(act_buffer_inst_int_data1[21]), .A2(
        act_buffer_inst_n183), .B1(act_buffer_inst_int_data1[5]), .B2(
        act_buffer_inst_n177), .C1(act_buffer_inst_int_data1[13]), .C2(
        act_buffer_inst_n171), .ZN(act_buffer_inst_n133) );
  NAND2_X1 act_buffer_inst_U273 ( .A1(act_buffer_inst_n132), .A2(
        act_buffer_inst_n133), .ZN(int_i_data_if1[5]) );
  AOI222_X1 act_buffer_inst_U272 ( .A1(act_buffer_inst_int_data2[21]), .A2(
        act_buffer_inst_n184), .B1(act_buffer_inst_int_data2[5]), .B2(
        act_buffer_inst_n178), .C1(act_buffer_inst_int_data2[13]), .C2(
        act_buffer_inst_n172), .ZN(act_buffer_inst_n117) );
  AOI222_X1 act_buffer_inst_U264 ( .A1(act_buffer_inst_int_data2[45]), .A2(
        act_buffer_inst_n166), .B1(act_buffer_inst_int_data2[29]), .B2(
        act_buffer_inst_n160), .C1(act_buffer_inst_int_data2[37]), .C2(
        act_buffer_inst_n5), .ZN(act_buffer_inst_n116) );
  NAND2_X1 act_buffer_inst_U263 ( .A1(act_buffer_inst_n116), .A2(
        act_buffer_inst_n117), .ZN(int_i_data_if2[5]) );
  AOI222_X1 act_buffer_inst_U262 ( .A1(act_buffer_inst_int_data3[21]), .A2(
        act_buffer_inst_n184), .B1(act_buffer_inst_int_data3[5]), .B2(
        act_buffer_inst_n178), .C1(act_buffer_inst_int_data3[13]), .C2(
        act_buffer_inst_n172), .ZN(act_buffer_inst_n101) );
  AOI222_X1 act_buffer_inst_U261 ( .A1(act_buffer_inst_int_data3[45]), .A2(
        act_buffer_inst_n166), .B1(act_buffer_inst_int_data3[29]), .B2(
        act_buffer_inst_n160), .C1(act_buffer_inst_int_data3[37]), .C2(
        act_buffer_inst_n5), .ZN(act_buffer_inst_n100) );
  NAND2_X1 act_buffer_inst_U260 ( .A1(act_buffer_inst_n100), .A2(
        act_buffer_inst_n101), .ZN(int_i_data_if3[5]) );
  AOI222_X1 act_buffer_inst_U259 ( .A1(act_buffer_inst_int_data4[21]), .A2(
        act_buffer_inst_n185), .B1(act_buffer_inst_int_data4[5]), .B2(
        act_buffer_inst_n179), .C1(act_buffer_inst_int_data4[13]), .C2(
        act_buffer_inst_n173), .ZN(act_buffer_inst_n85) );
  AOI222_X1 act_buffer_inst_U258 ( .A1(act_buffer_inst_int_data4[45]), .A2(
        act_buffer_inst_n167), .B1(act_buffer_inst_int_data4[29]), .B2(
        act_buffer_inst_n161), .C1(act_buffer_inst_int_data4[37]), .C2(
        act_buffer_inst_n6), .ZN(act_buffer_inst_n84) );
  NAND2_X1 act_buffer_inst_U257 ( .A1(act_buffer_inst_n84), .A2(
        act_buffer_inst_n85), .ZN(int_i_data_if4[5]) );
  AOI222_X1 act_buffer_inst_U256 ( .A1(act_buffer_inst_int_data1[47]), .A2(
        act_buffer_inst_n165), .B1(act_buffer_inst_int_data1[31]), .B2(
        act_buffer_inst_n159), .C1(act_buffer_inst_int_data1[39]), .C2(
        act_buffer_inst_n4), .ZN(act_buffer_inst_n128) );
  AOI222_X1 act_buffer_inst_U255 ( .A1(act_buffer_inst_int_data1[23]), .A2(
        act_buffer_inst_n183), .B1(act_buffer_inst_int_data1[7]), .B2(
        act_buffer_inst_n177), .C1(act_buffer_inst_int_data1[15]), .C2(
        act_buffer_inst_n171), .ZN(act_buffer_inst_n129) );
  NAND2_X1 act_buffer_inst_U254 ( .A1(act_buffer_inst_n128), .A2(
        act_buffer_inst_n129), .ZN(int_i_data_if1[7]) );
  AOI222_X1 act_buffer_inst_U253 ( .A1(act_buffer_inst_int_data2[23]), .A2(
        act_buffer_inst_n184), .B1(act_buffer_inst_int_data2[7]), .B2(
        act_buffer_inst_n178), .C1(act_buffer_inst_int_data2[15]), .C2(
        act_buffer_inst_n172), .ZN(act_buffer_inst_n113) );
  AOI222_X1 act_buffer_inst_U252 ( .A1(act_buffer_inst_int_data2[47]), .A2(
        act_buffer_inst_n166), .B1(act_buffer_inst_int_data2[31]), .B2(
        act_buffer_inst_n160), .C1(act_buffer_inst_int_data2[39]), .C2(
        act_buffer_inst_n5), .ZN(act_buffer_inst_n112) );
  NAND2_X1 act_buffer_inst_U251 ( .A1(act_buffer_inst_n112), .A2(
        act_buffer_inst_n113), .ZN(int_i_data_if2[7]) );
  AOI222_X1 act_buffer_inst_U250 ( .A1(act_buffer_inst_int_data3[23]), .A2(
        act_buffer_inst_n184), .B1(act_buffer_inst_int_data3[7]), .B2(
        act_buffer_inst_n178), .C1(act_buffer_inst_int_data3[15]), .C2(
        act_buffer_inst_n172), .ZN(act_buffer_inst_n97) );
  AOI222_X1 act_buffer_inst_U249 ( .A1(act_buffer_inst_int_data3[47]), .A2(
        act_buffer_inst_n166), .B1(act_buffer_inst_int_data3[31]), .B2(
        act_buffer_inst_n160), .C1(act_buffer_inst_int_data3[39]), .C2(
        act_buffer_inst_n5), .ZN(act_buffer_inst_n96) );
  NAND2_X1 act_buffer_inst_U248 ( .A1(act_buffer_inst_n96), .A2(
        act_buffer_inst_n97), .ZN(int_i_data_if3[7]) );
  AOI222_X1 act_buffer_inst_U247 ( .A1(act_buffer_inst_int_data4[23]), .A2(
        act_buffer_inst_n185), .B1(act_buffer_inst_int_data4[7]), .B2(
        act_buffer_inst_n179), .C1(act_buffer_inst_int_data4[15]), .C2(
        act_buffer_inst_n173), .ZN(act_buffer_inst_n81) );
  AOI222_X1 act_buffer_inst_U246 ( .A1(act_buffer_inst_int_data4[47]), .A2(
        act_buffer_inst_n167), .B1(act_buffer_inst_int_data4[31]), .B2(
        act_buffer_inst_n161), .C1(act_buffer_inst_int_data4[39]), .C2(
        act_buffer_inst_n6), .ZN(act_buffer_inst_n80) );
  NAND2_X1 act_buffer_inst_U245 ( .A1(act_buffer_inst_n80), .A2(
        act_buffer_inst_n81), .ZN(int_i_data_if4[7]) );
  AOI222_X1 act_buffer_inst_U244 ( .A1(act_buffer_inst_int_data1[41]), .A2(
        act_buffer_inst_n165), .B1(act_buffer_inst_int_data1[25]), .B2(
        act_buffer_inst_n159), .C1(act_buffer_inst_int_data1[33]), .C2(
        act_buffer_inst_n4), .ZN(act_buffer_inst_n140) );
  AOI222_X1 act_buffer_inst_U243 ( .A1(act_buffer_inst_int_data1[17]), .A2(
        act_buffer_inst_n183), .B1(act_buffer_inst_int_data1[1]), .B2(
        act_buffer_inst_n177), .C1(act_buffer_inst_int_data1[9]), .C2(
        act_buffer_inst_n171), .ZN(act_buffer_inst_n141) );
  NAND2_X1 act_buffer_inst_U242 ( .A1(act_buffer_inst_n140), .A2(
        act_buffer_inst_n141), .ZN(int_i_data_if1[1]) );
  AOI222_X1 act_buffer_inst_U241 ( .A1(act_buffer_inst_int_data2[41]), .A2(
        act_buffer_inst_n165), .B1(act_buffer_inst_int_data2[25]), .B2(
        act_buffer_inst_n159), .C1(act_buffer_inst_int_data2[33]), .C2(
        act_buffer_inst_n4), .ZN(act_buffer_inst_n124) );
  AOI222_X1 act_buffer_inst_U240 ( .A1(act_buffer_inst_int_data2[17]), .A2(
        act_buffer_inst_n183), .B1(act_buffer_inst_int_data2[1]), .B2(
        act_buffer_inst_n177), .C1(act_buffer_inst_int_data2[9]), .C2(
        act_buffer_inst_n171), .ZN(act_buffer_inst_n125) );
  NAND2_X1 act_buffer_inst_U239 ( .A1(act_buffer_inst_n124), .A2(
        act_buffer_inst_n125), .ZN(int_i_data_if2[1]) );
  AOI222_X1 act_buffer_inst_U238 ( .A1(act_buffer_inst_int_data5[17]), .A2(
        act_buffer_inst_n185), .B1(act_buffer_inst_int_data5[1]), .B2(
        act_buffer_inst_n179), .C1(act_buffer_inst_int_data5[9]), .C2(
        act_buffer_inst_n173), .ZN(act_buffer_inst_n77) );
  AOI222_X1 act_buffer_inst_U237 ( .A1(act_buffer_inst_int_data5[41]), .A2(
        act_buffer_inst_n167), .B1(act_buffer_inst_int_data5[25]), .B2(
        act_buffer_inst_n161), .C1(act_buffer_inst_int_data5[33]), .C2(
        act_buffer_inst_n6), .ZN(act_buffer_inst_n76) );
  NAND2_X1 act_buffer_inst_U236 ( .A1(act_buffer_inst_n76), .A2(
        act_buffer_inst_n77), .ZN(int_i_data_if5[1]) );
  AOI222_X1 act_buffer_inst_U235 ( .A1(act_buffer_inst_int_data3[17]), .A2(
        act_buffer_inst_n184), .B1(act_buffer_inst_int_data3[1]), .B2(
        act_buffer_inst_n178), .C1(act_buffer_inst_int_data3[9]), .C2(
        act_buffer_inst_n172), .ZN(act_buffer_inst_n109) );
  AOI222_X1 act_buffer_inst_U234 ( .A1(act_buffer_inst_int_data3[41]), .A2(
        act_buffer_inst_n166), .B1(act_buffer_inst_int_data3[25]), .B2(
        act_buffer_inst_n160), .C1(act_buffer_inst_int_data3[33]), .C2(
        act_buffer_inst_n5), .ZN(act_buffer_inst_n108) );
  NAND2_X1 act_buffer_inst_U233 ( .A1(act_buffer_inst_n108), .A2(
        act_buffer_inst_n109), .ZN(int_i_data_if3[1]) );
  AOI222_X1 act_buffer_inst_U232 ( .A1(act_buffer_inst_int_data4[17]), .A2(
        act_buffer_inst_n185), .B1(act_buffer_inst_int_data4[1]), .B2(
        act_buffer_inst_n179), .C1(act_buffer_inst_int_data4[9]), .C2(
        act_buffer_inst_n173), .ZN(act_buffer_inst_n93) );
  AOI222_X1 act_buffer_inst_U231 ( .A1(act_buffer_inst_int_data4[41]), .A2(
        act_buffer_inst_n167), .B1(act_buffer_inst_int_data4[25]), .B2(
        act_buffer_inst_n161), .C1(act_buffer_inst_int_data4[33]), .C2(
        act_buffer_inst_n6), .ZN(act_buffer_inst_n92) );
  NAND2_X1 act_buffer_inst_U230 ( .A1(act_buffer_inst_n92), .A2(
        act_buffer_inst_n93), .ZN(int_i_data_if4[1]) );
  AOI222_X1 act_buffer_inst_U229 ( .A1(act_buffer_inst_int_data1[42]), .A2(
        act_buffer_inst_n165), .B1(act_buffer_inst_int_data1[26]), .B2(
        act_buffer_inst_n159), .C1(act_buffer_inst_int_data1[34]), .C2(
        act_buffer_inst_n4), .ZN(act_buffer_inst_n138) );
  AOI222_X1 act_buffer_inst_U228 ( .A1(act_buffer_inst_int_data1[18]), .A2(
        act_buffer_inst_n183), .B1(act_buffer_inst_int_data1[2]), .B2(
        act_buffer_inst_n177), .C1(act_buffer_inst_int_data1[10]), .C2(
        act_buffer_inst_n171), .ZN(act_buffer_inst_n139) );
  NAND2_X1 act_buffer_inst_U227 ( .A1(act_buffer_inst_n138), .A2(
        act_buffer_inst_n139), .ZN(int_i_data_if1[2]) );
  AOI222_X1 act_buffer_inst_U226 ( .A1(act_buffer_inst_int_data2[42]), .A2(
        act_buffer_inst_n165), .B1(act_buffer_inst_int_data2[26]), .B2(
        act_buffer_inst_n159), .C1(act_buffer_inst_int_data2[34]), .C2(
        act_buffer_inst_n4), .ZN(act_buffer_inst_n122) );
  AOI222_X1 act_buffer_inst_U225 ( .A1(act_buffer_inst_int_data2[18]), .A2(
        act_buffer_inst_n183), .B1(act_buffer_inst_int_data2[2]), .B2(
        act_buffer_inst_n177), .C1(act_buffer_inst_int_data2[10]), .C2(
        act_buffer_inst_n171), .ZN(act_buffer_inst_n123) );
  NAND2_X1 act_buffer_inst_U224 ( .A1(act_buffer_inst_n122), .A2(
        act_buffer_inst_n123), .ZN(int_i_data_if2[2]) );
  AOI222_X1 act_buffer_inst_U223 ( .A1(act_buffer_inst_int_data5[18]), .A2(
        act_buffer_inst_n185), .B1(act_buffer_inst_int_data5[2]), .B2(
        act_buffer_inst_n179), .C1(act_buffer_inst_int_data5[10]), .C2(
        act_buffer_inst_n173), .ZN(act_buffer_inst_n75) );
  AOI222_X1 act_buffer_inst_U222 ( .A1(act_buffer_inst_int_data5[42]), .A2(
        act_buffer_inst_n167), .B1(act_buffer_inst_int_data5[26]), .B2(
        act_buffer_inst_n161), .C1(act_buffer_inst_int_data5[34]), .C2(
        act_buffer_inst_n6), .ZN(act_buffer_inst_n74) );
  NAND2_X1 act_buffer_inst_U221 ( .A1(act_buffer_inst_n74), .A2(
        act_buffer_inst_n75), .ZN(int_i_data_if5[2]) );
  AOI222_X1 act_buffer_inst_U220 ( .A1(act_buffer_inst_int_data3[18]), .A2(
        act_buffer_inst_n184), .B1(act_buffer_inst_int_data3[2]), .B2(
        act_buffer_inst_n178), .C1(act_buffer_inst_int_data3[10]), .C2(
        act_buffer_inst_n172), .ZN(act_buffer_inst_n107) );
  AOI222_X1 act_buffer_inst_U219 ( .A1(act_buffer_inst_int_data3[42]), .A2(
        act_buffer_inst_n166), .B1(act_buffer_inst_int_data3[26]), .B2(
        act_buffer_inst_n160), .C1(act_buffer_inst_int_data3[34]), .C2(
        act_buffer_inst_n5), .ZN(act_buffer_inst_n106) );
  NAND2_X1 act_buffer_inst_U218 ( .A1(act_buffer_inst_n106), .A2(
        act_buffer_inst_n107), .ZN(int_i_data_if3[2]) );
  AOI222_X1 act_buffer_inst_U217 ( .A1(act_buffer_inst_int_data4[18]), .A2(
        act_buffer_inst_n185), .B1(act_buffer_inst_int_data4[2]), .B2(
        act_buffer_inst_n179), .C1(act_buffer_inst_int_data4[10]), .C2(
        act_buffer_inst_n173), .ZN(act_buffer_inst_n91) );
  AOI222_X1 act_buffer_inst_U216 ( .A1(act_buffer_inst_int_data4[42]), .A2(
        act_buffer_inst_n167), .B1(act_buffer_inst_int_data4[26]), .B2(
        act_buffer_inst_n161), .C1(act_buffer_inst_int_data4[34]), .C2(
        act_buffer_inst_n6), .ZN(act_buffer_inst_n90) );
  NAND2_X1 act_buffer_inst_U215 ( .A1(act_buffer_inst_n90), .A2(
        act_buffer_inst_n91), .ZN(int_i_data_if4[2]) );
  AOI222_X1 act_buffer_inst_U214 ( .A1(act_buffer_inst_int_data1[20]), .A2(
        act_buffer_inst_n183), .B1(act_buffer_inst_int_data1[4]), .B2(
        act_buffer_inst_n177), .C1(act_buffer_inst_int_data1[12]), .C2(
        act_buffer_inst_n171), .ZN(act_buffer_inst_n135) );
  AOI222_X1 act_buffer_inst_U213 ( .A1(act_buffer_inst_int_data1[44]), .A2(
        act_buffer_inst_n165), .B1(act_buffer_inst_int_data1[28]), .B2(
        act_buffer_inst_n159), .C1(act_buffer_inst_int_data1[36]), .C2(
        act_buffer_inst_n4), .ZN(act_buffer_inst_n134) );
  NAND2_X1 act_buffer_inst_U212 ( .A1(act_buffer_inst_n134), .A2(
        act_buffer_inst_n135), .ZN(int_i_data_if1[4]) );
  AOI222_X1 act_buffer_inst_U211 ( .A1(act_buffer_inst_int_data2[20]), .A2(
        act_buffer_inst_n184), .B1(act_buffer_inst_int_data2[4]), .B2(
        act_buffer_inst_n178), .C1(act_buffer_inst_int_data2[12]), .C2(
        act_buffer_inst_n172), .ZN(act_buffer_inst_n119) );
  AOI222_X1 act_buffer_inst_U210 ( .A1(act_buffer_inst_int_data2[44]), .A2(
        act_buffer_inst_n166), .B1(act_buffer_inst_int_data2[28]), .B2(
        act_buffer_inst_n160), .C1(act_buffer_inst_int_data2[36]), .C2(
        act_buffer_inst_n5), .ZN(act_buffer_inst_n118) );
  NAND2_X1 act_buffer_inst_U209 ( .A1(act_buffer_inst_n118), .A2(
        act_buffer_inst_n119), .ZN(int_i_data_if2[4]) );
  AOI222_X1 act_buffer_inst_U208 ( .A1(act_buffer_inst_int_data3[20]), .A2(
        act_buffer_inst_n184), .B1(act_buffer_inst_int_data3[4]), .B2(
        act_buffer_inst_n178), .C1(act_buffer_inst_int_data3[12]), .C2(
        act_buffer_inst_n172), .ZN(act_buffer_inst_n103) );
  AOI222_X1 act_buffer_inst_U207 ( .A1(act_buffer_inst_int_data3[44]), .A2(
        act_buffer_inst_n166), .B1(act_buffer_inst_int_data3[28]), .B2(
        act_buffer_inst_n160), .C1(act_buffer_inst_int_data3[36]), .C2(
        act_buffer_inst_n5), .ZN(act_buffer_inst_n102) );
  NAND2_X1 act_buffer_inst_U206 ( .A1(act_buffer_inst_n102), .A2(
        act_buffer_inst_n103), .ZN(int_i_data_if3[4]) );
  AOI222_X1 act_buffer_inst_U205 ( .A1(act_buffer_inst_int_data4[20]), .A2(
        act_buffer_inst_n185), .B1(act_buffer_inst_int_data4[4]), .B2(
        act_buffer_inst_n179), .C1(act_buffer_inst_int_data4[12]), .C2(
        act_buffer_inst_n173), .ZN(act_buffer_inst_n87) );
  AOI222_X1 act_buffer_inst_U204 ( .A1(act_buffer_inst_int_data4[44]), .A2(
        act_buffer_inst_n167), .B1(act_buffer_inst_int_data4[28]), .B2(
        act_buffer_inst_n161), .C1(act_buffer_inst_int_data4[36]), .C2(
        act_buffer_inst_n6), .ZN(act_buffer_inst_n86) );
  NAND2_X1 act_buffer_inst_U203 ( .A1(act_buffer_inst_n86), .A2(
        act_buffer_inst_n87), .ZN(int_i_data_if4[4]) );
  AOI222_X1 act_buffer_inst_U202 ( .A1(act_buffer_inst_int_data1[46]), .A2(
        act_buffer_inst_n165), .B1(act_buffer_inst_int_data1[30]), .B2(
        act_buffer_inst_n159), .C1(act_buffer_inst_int_data1[38]), .C2(
        act_buffer_inst_n4), .ZN(act_buffer_inst_n130) );
  AOI222_X1 act_buffer_inst_U201 ( .A1(act_buffer_inst_int_data1[22]), .A2(
        act_buffer_inst_n183), .B1(act_buffer_inst_int_data1[6]), .B2(
        act_buffer_inst_n177), .C1(act_buffer_inst_int_data1[14]), .C2(
        act_buffer_inst_n171), .ZN(act_buffer_inst_n131) );
  NAND2_X1 act_buffer_inst_U200 ( .A1(act_buffer_inst_n130), .A2(
        act_buffer_inst_n131), .ZN(int_i_data_if1[6]) );
  AOI222_X1 act_buffer_inst_U199 ( .A1(act_buffer_inst_int_data2[22]), .A2(
        act_buffer_inst_n184), .B1(act_buffer_inst_int_data2[6]), .B2(
        act_buffer_inst_n178), .C1(act_buffer_inst_int_data2[14]), .C2(
        act_buffer_inst_n172), .ZN(act_buffer_inst_n115) );
  AOI222_X1 act_buffer_inst_U198 ( .A1(act_buffer_inst_int_data2[46]), .A2(
        act_buffer_inst_n166), .B1(act_buffer_inst_int_data2[30]), .B2(
        act_buffer_inst_n160), .C1(act_buffer_inst_int_data2[38]), .C2(
        act_buffer_inst_n5), .ZN(act_buffer_inst_n114) );
  NAND2_X1 act_buffer_inst_U197 ( .A1(act_buffer_inst_n114), .A2(
        act_buffer_inst_n115), .ZN(int_i_data_if2[6]) );
  AOI222_X1 act_buffer_inst_U196 ( .A1(act_buffer_inst_int_data3[22]), .A2(
        act_buffer_inst_n184), .B1(act_buffer_inst_int_data3[6]), .B2(
        act_buffer_inst_n178), .C1(act_buffer_inst_int_data3[14]), .C2(
        act_buffer_inst_n172), .ZN(act_buffer_inst_n99) );
  AOI222_X1 act_buffer_inst_U195 ( .A1(act_buffer_inst_int_data3[46]), .A2(
        act_buffer_inst_n166), .B1(act_buffer_inst_int_data3[30]), .B2(
        act_buffer_inst_n160), .C1(act_buffer_inst_int_data3[38]), .C2(
        act_buffer_inst_n5), .ZN(act_buffer_inst_n98) );
  NAND2_X1 act_buffer_inst_U194 ( .A1(act_buffer_inst_n98), .A2(
        act_buffer_inst_n99), .ZN(int_i_data_if3[6]) );
  AOI222_X1 act_buffer_inst_U193 ( .A1(act_buffer_inst_int_data4[22]), .A2(
        act_buffer_inst_n185), .B1(act_buffer_inst_int_data4[6]), .B2(
        act_buffer_inst_n179), .C1(act_buffer_inst_int_data4[14]), .C2(
        act_buffer_inst_n173), .ZN(act_buffer_inst_n83) );
  AOI222_X1 act_buffer_inst_U192 ( .A1(act_buffer_inst_int_data4[46]), .A2(
        act_buffer_inst_n167), .B1(act_buffer_inst_int_data4[30]), .B2(
        act_buffer_inst_n161), .C1(act_buffer_inst_int_data4[38]), .C2(
        act_buffer_inst_n6), .ZN(act_buffer_inst_n82) );
  NAND2_X1 act_buffer_inst_U191 ( .A1(act_buffer_inst_n82), .A2(
        act_buffer_inst_n83), .ZN(int_i_data_if4[6]) );
  AOI222_X1 act_buffer_inst_U190 ( .A1(act_buffer_inst_int_data1[40]), .A2(
        act_buffer_inst_n165), .B1(act_buffer_inst_int_data1[24]), .B2(
        act_buffer_inst_n159), .C1(act_buffer_inst_int_data1[32]), .C2(
        act_buffer_inst_n4), .ZN(act_buffer_inst_n142) );
  AOI222_X1 act_buffer_inst_U189 ( .A1(act_buffer_inst_int_data1[16]), .A2(
        act_buffer_inst_n183), .B1(act_buffer_inst_int_data1[0]), .B2(
        act_buffer_inst_n177), .C1(act_buffer_inst_int_data1[8]), .C2(
        act_buffer_inst_n171), .ZN(act_buffer_inst_n143) );
  NAND2_X1 act_buffer_inst_U188 ( .A1(act_buffer_inst_n142), .A2(
        act_buffer_inst_n143), .ZN(int_i_data_if1[0]) );
  AOI222_X1 act_buffer_inst_U187 ( .A1(act_buffer_inst_int_data2[40]), .A2(
        act_buffer_inst_n165), .B1(act_buffer_inst_int_data2[24]), .B2(
        act_buffer_inst_n159), .C1(act_buffer_inst_int_data2[32]), .C2(
        act_buffer_inst_n4), .ZN(act_buffer_inst_n126) );
  AOI222_X1 act_buffer_inst_U186 ( .A1(act_buffer_inst_int_data2[16]), .A2(
        act_buffer_inst_n183), .B1(act_buffer_inst_int_data2[0]), .B2(
        act_buffer_inst_n177), .C1(act_buffer_inst_int_data2[8]), .C2(
        act_buffer_inst_n171), .ZN(act_buffer_inst_n127) );
  NAND2_X1 act_buffer_inst_U185 ( .A1(act_buffer_inst_n126), .A2(
        act_buffer_inst_n127), .ZN(int_i_data_if2[0]) );
  AOI222_X1 act_buffer_inst_U184 ( .A1(act_buffer_inst_int_data5[16]), .A2(
        act_buffer_inst_n185), .B1(act_buffer_inst_int_data5[0]), .B2(
        act_buffer_inst_n179), .C1(act_buffer_inst_int_data5[8]), .C2(
        act_buffer_inst_n173), .ZN(act_buffer_inst_n79) );
  AOI222_X1 act_buffer_inst_U183 ( .A1(act_buffer_inst_int_data5[40]), .A2(
        act_buffer_inst_n167), .B1(act_buffer_inst_int_data5[24]), .B2(
        act_buffer_inst_n161), .C1(act_buffer_inst_int_data5[32]), .C2(
        act_buffer_inst_n6), .ZN(act_buffer_inst_n78) );
  NAND2_X1 act_buffer_inst_U182 ( .A1(act_buffer_inst_n78), .A2(
        act_buffer_inst_n79), .ZN(int_i_data_if5[0]) );
  AOI222_X1 act_buffer_inst_U181 ( .A1(act_buffer_inst_int_data4[16]), .A2(
        act_buffer_inst_n185), .B1(act_buffer_inst_int_data4[0]), .B2(
        act_buffer_inst_n179), .C1(act_buffer_inst_int_data4[8]), .C2(
        act_buffer_inst_n173), .ZN(act_buffer_inst_n95) );
  AOI222_X1 act_buffer_inst_U180 ( .A1(act_buffer_inst_int_data4[40]), .A2(
        act_buffer_inst_n167), .B1(act_buffer_inst_int_data4[24]), .B2(
        act_buffer_inst_n161), .C1(act_buffer_inst_int_data4[32]), .C2(
        act_buffer_inst_n6), .ZN(act_buffer_inst_n94) );
  NAND2_X1 act_buffer_inst_U179 ( .A1(act_buffer_inst_n94), .A2(
        act_buffer_inst_n95), .ZN(int_i_data_if4[0]) );
  AOI222_X1 act_buffer_inst_U178 ( .A1(act_buffer_inst_int_data3[16]), .A2(
        act_buffer_inst_n184), .B1(act_buffer_inst_int_data3[0]), .B2(
        act_buffer_inst_n178), .C1(act_buffer_inst_int_data3[8]), .C2(
        act_buffer_inst_n172), .ZN(act_buffer_inst_n111) );
  AOI222_X1 act_buffer_inst_U177 ( .A1(act_buffer_inst_int_data3[40]), .A2(
        act_buffer_inst_n166), .B1(act_buffer_inst_int_data3[24]), .B2(
        act_buffer_inst_n160), .C1(act_buffer_inst_int_data3[32]), .C2(
        act_buffer_inst_n5), .ZN(act_buffer_inst_n110) );
  NAND2_X1 act_buffer_inst_U176 ( .A1(act_buffer_inst_n110), .A2(
        act_buffer_inst_n111), .ZN(int_i_data_if3[0]) );
  AOI222_X1 act_buffer_inst_U175 ( .A1(act_buffer_inst_int_data6[19]), .A2(
        act_buffer_inst_n186), .B1(act_buffer_inst_int_data6[3]), .B2(
        act_buffer_inst_n180), .C1(act_buffer_inst_int_data6[11]), .C2(
        act_buffer_inst_n174), .ZN(act_buffer_inst_n57) );
  AOI222_X1 act_buffer_inst_U174 ( .A1(act_buffer_inst_int_data6[43]), .A2(
        act_buffer_inst_n168), .B1(act_buffer_inst_int_data6[27]), .B2(
        act_buffer_inst_n162), .C1(act_buffer_inst_int_data6[35]), .C2(
        act_buffer_inst_n7), .ZN(act_buffer_inst_n56) );
  NAND2_X1 act_buffer_inst_U173 ( .A1(act_buffer_inst_n56), .A2(
        act_buffer_inst_n57), .ZN(int_i_data_if6[3]) );
  AOI222_X1 act_buffer_inst_U172 ( .A1(act_buffer_inst_int_data7[19]), .A2(
        act_buffer_inst_n187), .B1(act_buffer_inst_int_data7[3]), .B2(
        act_buffer_inst_n181), .C1(act_buffer_inst_int_data7[11]), .C2(
        act_buffer_inst_n175), .ZN(act_buffer_inst_n41) );
  AOI222_X1 act_buffer_inst_U171 ( .A1(act_buffer_inst_int_data7[43]), .A2(
        act_buffer_inst_n169), .B1(act_buffer_inst_int_data7[27]), .B2(
        act_buffer_inst_n163), .C1(act_buffer_inst_int_data7[35]), .C2(
        act_buffer_inst_n8), .ZN(act_buffer_inst_n40) );
  NAND2_X1 act_buffer_inst_U170 ( .A1(act_buffer_inst_n40), .A2(
        act_buffer_inst_n41), .ZN(int_i_data_if7[3]) );
  AOI222_X1 act_buffer_inst_U169 ( .A1(act_buffer_inst_int_data8[19]), .A2(
        act_buffer_inst_n187), .B1(act_buffer_inst_int_data8[3]), .B2(
        act_buffer_inst_n181), .C1(act_buffer_inst_int_data8[11]), .C2(
        act_buffer_inst_n175), .ZN(act_buffer_inst_n25) );
  AOI222_X1 act_buffer_inst_U168 ( .A1(act_buffer_inst_int_data8[43]), .A2(
        act_buffer_inst_n169), .B1(act_buffer_inst_int_data8[27]), .B2(
        act_buffer_inst_n163), .C1(act_buffer_inst_int_data8[35]), .C2(
        act_buffer_inst_n8), .ZN(act_buffer_inst_n24) );
  NAND2_X1 act_buffer_inst_U167 ( .A1(act_buffer_inst_n24), .A2(
        act_buffer_inst_n25), .ZN(int_i_data_if8[3]) );
  AOI222_X1 act_buffer_inst_U166 ( .A1(act_buffer_inst_int_data5[21]), .A2(
        act_buffer_inst_n186), .B1(act_buffer_inst_int_data5[5]), .B2(
        act_buffer_inst_n180), .C1(act_buffer_inst_int_data5[13]), .C2(
        act_buffer_inst_n174), .ZN(act_buffer_inst_n69) );
  AOI222_X1 act_buffer_inst_U165 ( .A1(act_buffer_inst_int_data5[45]), .A2(
        act_buffer_inst_n168), .B1(act_buffer_inst_int_data5[29]), .B2(
        act_buffer_inst_n162), .C1(act_buffer_inst_int_data5[37]), .C2(
        act_buffer_inst_n7), .ZN(act_buffer_inst_n68) );
  NAND2_X1 act_buffer_inst_U164 ( .A1(act_buffer_inst_n68), .A2(
        act_buffer_inst_n69), .ZN(int_i_data_if5[5]) );
  AOI222_X1 act_buffer_inst_U163 ( .A1(act_buffer_inst_int_data6[21]), .A2(
        act_buffer_inst_n186), .B1(act_buffer_inst_int_data6[5]), .B2(
        act_buffer_inst_n180), .C1(act_buffer_inst_int_data6[13]), .C2(
        act_buffer_inst_n174), .ZN(act_buffer_inst_n53) );
  AOI222_X1 act_buffer_inst_U162 ( .A1(act_buffer_inst_int_data6[45]), .A2(
        act_buffer_inst_n168), .B1(act_buffer_inst_int_data6[29]), .B2(
        act_buffer_inst_n162), .C1(act_buffer_inst_int_data6[37]), .C2(
        act_buffer_inst_n7), .ZN(act_buffer_inst_n52) );
  NAND2_X1 act_buffer_inst_U161 ( .A1(act_buffer_inst_n52), .A2(
        act_buffer_inst_n53), .ZN(int_i_data_if6[5]) );
  AOI222_X1 act_buffer_inst_U160 ( .A1(act_buffer_inst_int_data8[21]), .A2(
        act_buffer_inst_n188), .B1(act_buffer_inst_int_data8[5]), .B2(
        act_buffer_inst_n182), .C1(act_buffer_inst_int_data8[13]), .C2(
        act_buffer_inst_n176), .ZN(act_buffer_inst_n21) );
  AOI222_X1 act_buffer_inst_U159 ( .A1(act_buffer_inst_int_data8[45]), .A2(
        act_buffer_inst_n170), .B1(act_buffer_inst_int_data8[29]), .B2(
        act_buffer_inst_n164), .C1(act_buffer_inst_int_data8[37]), .C2(
        act_buffer_inst_n9), .ZN(act_buffer_inst_n20) );
  NAND2_X1 act_buffer_inst_U158 ( .A1(act_buffer_inst_n20), .A2(
        act_buffer_inst_n21), .ZN(int_i_data_if8[5]) );
  AOI222_X1 act_buffer_inst_U157 ( .A1(act_buffer_inst_int_data7[21]), .A2(
        act_buffer_inst_n187), .B1(act_buffer_inst_int_data7[5]), .B2(
        act_buffer_inst_n181), .C1(act_buffer_inst_int_data7[13]), .C2(
        act_buffer_inst_n175), .ZN(act_buffer_inst_n37) );
  AOI222_X1 act_buffer_inst_U156 ( .A1(act_buffer_inst_int_data7[45]), .A2(
        act_buffer_inst_n169), .B1(act_buffer_inst_int_data7[29]), .B2(
        act_buffer_inst_n163), .C1(act_buffer_inst_int_data7[37]), .C2(
        act_buffer_inst_n8), .ZN(act_buffer_inst_n36) );
  NAND2_X1 act_buffer_inst_U155 ( .A1(act_buffer_inst_n36), .A2(
        act_buffer_inst_n37), .ZN(int_i_data_if7[5]) );
  AOI222_X1 act_buffer_inst_U154 ( .A1(act_buffer_inst_int_data5[23]), .A2(
        act_buffer_inst_n186), .B1(act_buffer_inst_int_data5[7]), .B2(
        act_buffer_inst_n180), .C1(act_buffer_inst_int_data5[15]), .C2(
        act_buffer_inst_n174), .ZN(act_buffer_inst_n65) );
  AOI222_X1 act_buffer_inst_U153 ( .A1(act_buffer_inst_int_data5[47]), .A2(
        act_buffer_inst_n168), .B1(act_buffer_inst_int_data5[31]), .B2(
        act_buffer_inst_n162), .C1(act_buffer_inst_int_data5[39]), .C2(
        act_buffer_inst_n7), .ZN(act_buffer_inst_n64) );
  NAND2_X1 act_buffer_inst_U152 ( .A1(act_buffer_inst_n64), .A2(
        act_buffer_inst_n65), .ZN(int_i_data_if5[7]) );
  AOI222_X1 act_buffer_inst_U151 ( .A1(act_buffer_inst_int_data6[23]), .A2(
        act_buffer_inst_n186), .B1(act_buffer_inst_int_data6[7]), .B2(
        act_buffer_inst_n180), .C1(act_buffer_inst_int_data6[15]), .C2(
        act_buffer_inst_n174), .ZN(act_buffer_inst_n49) );
  AOI222_X1 act_buffer_inst_U150 ( .A1(act_buffer_inst_int_data6[47]), .A2(
        act_buffer_inst_n168), .B1(act_buffer_inst_int_data6[31]), .B2(
        act_buffer_inst_n162), .C1(act_buffer_inst_int_data6[39]), .C2(
        act_buffer_inst_n7), .ZN(act_buffer_inst_n48) );
  NAND2_X1 act_buffer_inst_U149 ( .A1(act_buffer_inst_n48), .A2(
        act_buffer_inst_n49), .ZN(int_i_data_if6[7]) );
  AOI222_X1 act_buffer_inst_U148 ( .A1(act_buffer_inst_int_data8[47]), .A2(
        act_buffer_inst_n170), .B1(act_buffer_inst_int_data8[31]), .B2(
        act_buffer_inst_n164), .C1(act_buffer_inst_int_data8[39]), .C2(
        act_buffer_inst_n9), .ZN(act_buffer_inst_n10) );
  AOI222_X1 act_buffer_inst_U147 ( .A1(act_buffer_inst_int_data8[23]), .A2(
        act_buffer_inst_n188), .B1(act_buffer_inst_int_data8[7]), .B2(
        act_buffer_inst_n182), .C1(act_buffer_inst_int_data8[15]), .C2(
        act_buffer_inst_n176), .ZN(act_buffer_inst_n11) );
  NAND2_X1 act_buffer_inst_U146 ( .A1(act_buffer_inst_n10), .A2(
        act_buffer_inst_n11), .ZN(int_i_data_if8[7]) );
  AOI222_X1 act_buffer_inst_U145 ( .A1(act_buffer_inst_int_data7[23]), .A2(
        act_buffer_inst_n187), .B1(act_buffer_inst_int_data7[7]), .B2(
        act_buffer_inst_n181), .C1(act_buffer_inst_int_data7[15]), .C2(
        act_buffer_inst_n175), .ZN(act_buffer_inst_n33) );
  AOI222_X1 act_buffer_inst_U144 ( .A1(act_buffer_inst_int_data7[47]), .A2(
        act_buffer_inst_n169), .B1(act_buffer_inst_int_data7[31]), .B2(
        act_buffer_inst_n163), .C1(act_buffer_inst_int_data7[39]), .C2(
        act_buffer_inst_n8), .ZN(act_buffer_inst_n32) );
  NAND2_X1 act_buffer_inst_U143 ( .A1(act_buffer_inst_n32), .A2(
        act_buffer_inst_n33), .ZN(int_i_data_if7[7]) );
  AOI222_X1 act_buffer_inst_U142 ( .A1(act_buffer_inst_int_data6[17]), .A2(
        act_buffer_inst_n186), .B1(act_buffer_inst_int_data6[1]), .B2(
        act_buffer_inst_n180), .C1(act_buffer_inst_int_data6[9]), .C2(
        act_buffer_inst_n174), .ZN(act_buffer_inst_n61) );
  AOI222_X1 act_buffer_inst_U141 ( .A1(act_buffer_inst_int_data6[41]), .A2(
        act_buffer_inst_n168), .B1(act_buffer_inst_int_data6[25]), .B2(
        act_buffer_inst_n162), .C1(act_buffer_inst_int_data6[33]), .C2(
        act_buffer_inst_n7), .ZN(act_buffer_inst_n60) );
  NAND2_X1 act_buffer_inst_U140 ( .A1(act_buffer_inst_n60), .A2(
        act_buffer_inst_n61), .ZN(int_i_data_if6[1]) );
  AOI222_X1 act_buffer_inst_U139 ( .A1(act_buffer_inst_int_data7[17]), .A2(
        act_buffer_inst_n187), .B1(act_buffer_inst_int_data7[1]), .B2(
        act_buffer_inst_n181), .C1(act_buffer_inst_int_data7[9]), .C2(
        act_buffer_inst_n175), .ZN(act_buffer_inst_n45) );
  AOI222_X1 act_buffer_inst_U138 ( .A1(act_buffer_inst_int_data7[41]), .A2(
        act_buffer_inst_n169), .B1(act_buffer_inst_int_data7[25]), .B2(
        act_buffer_inst_n163), .C1(act_buffer_inst_int_data7[33]), .C2(
        act_buffer_inst_n8), .ZN(act_buffer_inst_n44) );
  NAND2_X1 act_buffer_inst_U137 ( .A1(act_buffer_inst_n44), .A2(
        act_buffer_inst_n45), .ZN(int_i_data_if7[1]) );
  AOI222_X1 act_buffer_inst_U136 ( .A1(act_buffer_inst_int_data8[17]), .A2(
        act_buffer_inst_n187), .B1(act_buffer_inst_int_data8[1]), .B2(
        act_buffer_inst_n181), .C1(act_buffer_inst_int_data8[9]), .C2(
        act_buffer_inst_n175), .ZN(act_buffer_inst_n29) );
  AOI222_X1 act_buffer_inst_U135 ( .A1(act_buffer_inst_int_data8[41]), .A2(
        act_buffer_inst_n169), .B1(act_buffer_inst_int_data8[25]), .B2(
        act_buffer_inst_n163), .C1(act_buffer_inst_int_data8[33]), .C2(
        act_buffer_inst_n8), .ZN(act_buffer_inst_n28) );
  NAND2_X1 act_buffer_inst_U134 ( .A1(act_buffer_inst_n28), .A2(
        act_buffer_inst_n29), .ZN(int_i_data_if8[1]) );
  AOI222_X1 act_buffer_inst_U133 ( .A1(act_buffer_inst_int_data6[18]), .A2(
        act_buffer_inst_n186), .B1(act_buffer_inst_int_data6[2]), .B2(
        act_buffer_inst_n180), .C1(act_buffer_inst_int_data6[10]), .C2(
        act_buffer_inst_n174), .ZN(act_buffer_inst_n59) );
  AOI222_X1 act_buffer_inst_U132 ( .A1(act_buffer_inst_int_data6[42]), .A2(
        act_buffer_inst_n168), .B1(act_buffer_inst_int_data6[26]), .B2(
        act_buffer_inst_n162), .C1(act_buffer_inst_int_data6[34]), .C2(
        act_buffer_inst_n7), .ZN(act_buffer_inst_n58) );
  NAND2_X1 act_buffer_inst_U131 ( .A1(act_buffer_inst_n58), .A2(
        act_buffer_inst_n59), .ZN(int_i_data_if6[2]) );
  AOI222_X1 act_buffer_inst_U130 ( .A1(act_buffer_inst_int_data7[18]), .A2(
        act_buffer_inst_n187), .B1(act_buffer_inst_int_data7[2]), .B2(
        act_buffer_inst_n181), .C1(act_buffer_inst_int_data7[10]), .C2(
        act_buffer_inst_n175), .ZN(act_buffer_inst_n43) );
  AOI222_X1 act_buffer_inst_U129 ( .A1(act_buffer_inst_int_data7[42]), .A2(
        act_buffer_inst_n169), .B1(act_buffer_inst_int_data7[26]), .B2(
        act_buffer_inst_n163), .C1(act_buffer_inst_int_data7[34]), .C2(
        act_buffer_inst_n8), .ZN(act_buffer_inst_n42) );
  NAND2_X1 act_buffer_inst_U128 ( .A1(act_buffer_inst_n42), .A2(
        act_buffer_inst_n43), .ZN(int_i_data_if7[2]) );
  AOI222_X1 act_buffer_inst_U127 ( .A1(act_buffer_inst_int_data8[18]), .A2(
        act_buffer_inst_n187), .B1(act_buffer_inst_int_data8[2]), .B2(
        act_buffer_inst_n181), .C1(act_buffer_inst_int_data8[10]), .C2(
        act_buffer_inst_n175), .ZN(act_buffer_inst_n27) );
  AOI222_X1 act_buffer_inst_U126 ( .A1(act_buffer_inst_int_data8[42]), .A2(
        act_buffer_inst_n169), .B1(act_buffer_inst_int_data8[26]), .B2(
        act_buffer_inst_n163), .C1(act_buffer_inst_int_data8[34]), .C2(
        act_buffer_inst_n8), .ZN(act_buffer_inst_n26) );
  NAND2_X1 act_buffer_inst_U125 ( .A1(act_buffer_inst_n26), .A2(
        act_buffer_inst_n27), .ZN(int_i_data_if8[2]) );
  AOI222_X1 act_buffer_inst_U124 ( .A1(act_buffer_inst_int_data6[20]), .A2(
        act_buffer_inst_n186), .B1(act_buffer_inst_int_data6[4]), .B2(
        act_buffer_inst_n180), .C1(act_buffer_inst_int_data6[12]), .C2(
        act_buffer_inst_n174), .ZN(act_buffer_inst_n55) );
  AOI222_X1 act_buffer_inst_U123 ( .A1(act_buffer_inst_int_data6[44]), .A2(
        act_buffer_inst_n168), .B1(act_buffer_inst_int_data6[28]), .B2(
        act_buffer_inst_n162), .C1(act_buffer_inst_int_data6[36]), .C2(
        act_buffer_inst_n7), .ZN(act_buffer_inst_n54) );
  NAND2_X1 act_buffer_inst_U122 ( .A1(act_buffer_inst_n54), .A2(
        act_buffer_inst_n55), .ZN(int_i_data_if6[4]) );
  AOI222_X1 act_buffer_inst_U121 ( .A1(act_buffer_inst_int_data5[20]), .A2(
        act_buffer_inst_n186), .B1(act_buffer_inst_int_data5[4]), .B2(
        act_buffer_inst_n180), .C1(act_buffer_inst_int_data5[12]), .C2(
        act_buffer_inst_n174), .ZN(act_buffer_inst_n71) );
  AOI222_X1 act_buffer_inst_U120 ( .A1(act_buffer_inst_int_data5[44]), .A2(
        act_buffer_inst_n168), .B1(act_buffer_inst_int_data5[28]), .B2(
        act_buffer_inst_n162), .C1(act_buffer_inst_int_data5[36]), .C2(
        act_buffer_inst_n7), .ZN(act_buffer_inst_n70) );
  NAND2_X1 act_buffer_inst_U119 ( .A1(act_buffer_inst_n70), .A2(
        act_buffer_inst_n71), .ZN(int_i_data_if5[4]) );
  AOI222_X1 act_buffer_inst_U118 ( .A1(act_buffer_inst_int_data8[20]), .A2(
        act_buffer_inst_n188), .B1(act_buffer_inst_int_data8[4]), .B2(
        act_buffer_inst_n182), .C1(act_buffer_inst_int_data8[12]), .C2(
        act_buffer_inst_n176), .ZN(act_buffer_inst_n23) );
  AOI222_X1 act_buffer_inst_U117 ( .A1(act_buffer_inst_int_data8[44]), .A2(
        act_buffer_inst_n170), .B1(act_buffer_inst_int_data8[28]), .B2(
        act_buffer_inst_n164), .C1(act_buffer_inst_int_data8[36]), .C2(
        act_buffer_inst_n9), .ZN(act_buffer_inst_n22) );
  NAND2_X1 act_buffer_inst_U116 ( .A1(act_buffer_inst_n22), .A2(
        act_buffer_inst_n23), .ZN(int_i_data_if8[4]) );
  AOI222_X1 act_buffer_inst_U115 ( .A1(act_buffer_inst_int_data7[20]), .A2(
        act_buffer_inst_n187), .B1(act_buffer_inst_int_data7[4]), .B2(
        act_buffer_inst_n181), .C1(act_buffer_inst_int_data7[12]), .C2(
        act_buffer_inst_n175), .ZN(act_buffer_inst_n39) );
  AOI222_X1 act_buffer_inst_U114 ( .A1(act_buffer_inst_int_data7[44]), .A2(
        act_buffer_inst_n169), .B1(act_buffer_inst_int_data7[28]), .B2(
        act_buffer_inst_n163), .C1(act_buffer_inst_int_data7[36]), .C2(
        act_buffer_inst_n8), .ZN(act_buffer_inst_n38) );
  NAND2_X1 act_buffer_inst_U113 ( .A1(act_buffer_inst_n38), .A2(
        act_buffer_inst_n39), .ZN(int_i_data_if7[4]) );
  AOI222_X1 act_buffer_inst_U112 ( .A1(act_buffer_inst_int_data5[22]), .A2(
        act_buffer_inst_n186), .B1(act_buffer_inst_int_data5[6]), .B2(
        act_buffer_inst_n180), .C1(act_buffer_inst_int_data5[14]), .C2(
        act_buffer_inst_n174), .ZN(act_buffer_inst_n67) );
  AOI222_X1 act_buffer_inst_U111 ( .A1(act_buffer_inst_int_data5[46]), .A2(
        act_buffer_inst_n168), .B1(act_buffer_inst_int_data5[30]), .B2(
        act_buffer_inst_n162), .C1(act_buffer_inst_int_data5[38]), .C2(
        act_buffer_inst_n7), .ZN(act_buffer_inst_n66) );
  NAND2_X1 act_buffer_inst_U110 ( .A1(act_buffer_inst_n66), .A2(
        act_buffer_inst_n67), .ZN(int_i_data_if5[6]) );
  AOI222_X1 act_buffer_inst_U109 ( .A1(act_buffer_inst_int_data6[22]), .A2(
        act_buffer_inst_n186), .B1(act_buffer_inst_int_data6[6]), .B2(
        act_buffer_inst_n180), .C1(act_buffer_inst_int_data6[14]), .C2(
        act_buffer_inst_n174), .ZN(act_buffer_inst_n51) );
  AOI222_X1 act_buffer_inst_U108 ( .A1(act_buffer_inst_int_data6[46]), .A2(
        act_buffer_inst_n168), .B1(act_buffer_inst_int_data6[30]), .B2(
        act_buffer_inst_n162), .C1(act_buffer_inst_int_data6[38]), .C2(
        act_buffer_inst_n7), .ZN(act_buffer_inst_n50) );
  NAND2_X1 act_buffer_inst_U107 ( .A1(act_buffer_inst_n50), .A2(
        act_buffer_inst_n51), .ZN(int_i_data_if6[6]) );
  AOI222_X1 act_buffer_inst_U106 ( .A1(act_buffer_inst_int_data8[46]), .A2(
        act_buffer_inst_n170), .B1(act_buffer_inst_int_data8[30]), .B2(
        act_buffer_inst_n164), .C1(act_buffer_inst_int_data8[38]), .C2(
        act_buffer_inst_n9), .ZN(act_buffer_inst_n18) );
  AOI222_X1 act_buffer_inst_U105 ( .A1(act_buffer_inst_int_data8[22]), .A2(
        act_buffer_inst_n188), .B1(act_buffer_inst_int_data8[6]), .B2(
        act_buffer_inst_n182), .C1(act_buffer_inst_int_data8[14]), .C2(
        act_buffer_inst_n176), .ZN(act_buffer_inst_n19) );
  NAND2_X1 act_buffer_inst_U104 ( .A1(act_buffer_inst_n18), .A2(
        act_buffer_inst_n19), .ZN(int_i_data_if8[6]) );
  AOI222_X1 act_buffer_inst_U103 ( .A1(act_buffer_inst_int_data7[22]), .A2(
        act_buffer_inst_n187), .B1(act_buffer_inst_int_data7[6]), .B2(
        act_buffer_inst_n181), .C1(act_buffer_inst_int_data7[14]), .C2(
        act_buffer_inst_n175), .ZN(act_buffer_inst_n35) );
  AOI222_X1 act_buffer_inst_U102 ( .A1(act_buffer_inst_int_data7[46]), .A2(
        act_buffer_inst_n169), .B1(act_buffer_inst_int_data7[30]), .B2(
        act_buffer_inst_n163), .C1(act_buffer_inst_int_data7[38]), .C2(
        act_buffer_inst_n8), .ZN(act_buffer_inst_n34) );
  NAND2_X1 act_buffer_inst_U101 ( .A1(act_buffer_inst_n34), .A2(
        act_buffer_inst_n35), .ZN(int_i_data_if7[6]) );
  AOI222_X1 act_buffer_inst_U100 ( .A1(act_buffer_inst_int_data6[16]), .A2(
        act_buffer_inst_n186), .B1(act_buffer_inst_int_data6[0]), .B2(
        act_buffer_inst_n180), .C1(act_buffer_inst_int_data6[8]), .C2(
        act_buffer_inst_n174), .ZN(act_buffer_inst_n63) );
  AOI222_X1 act_buffer_inst_U99 ( .A1(act_buffer_inst_int_data6[40]), .A2(
        act_buffer_inst_n168), .B1(act_buffer_inst_int_data6[24]), .B2(
        act_buffer_inst_n162), .C1(act_buffer_inst_int_data6[32]), .C2(
        act_buffer_inst_n7), .ZN(act_buffer_inst_n62) );
  NAND2_X1 act_buffer_inst_U98 ( .A1(act_buffer_inst_n62), .A2(
        act_buffer_inst_n63), .ZN(int_i_data_if6[0]) );
  AOI222_X1 act_buffer_inst_U97 ( .A1(act_buffer_inst_int_data8[16]), .A2(
        act_buffer_inst_n187), .B1(act_buffer_inst_int_data8[0]), .B2(
        act_buffer_inst_n181), .C1(act_buffer_inst_int_data8[8]), .C2(
        act_buffer_inst_n175), .ZN(act_buffer_inst_n31) );
  AOI222_X1 act_buffer_inst_U96 ( .A1(act_buffer_inst_int_data8[40]), .A2(
        act_buffer_inst_n169), .B1(act_buffer_inst_int_data8[24]), .B2(
        act_buffer_inst_n163), .C1(act_buffer_inst_int_data8[32]), .C2(
        act_buffer_inst_n8), .ZN(act_buffer_inst_n30) );
  NAND2_X1 act_buffer_inst_U95 ( .A1(act_buffer_inst_n30), .A2(
        act_buffer_inst_n31), .ZN(int_i_data_if8[0]) );
  AOI222_X1 act_buffer_inst_U94 ( .A1(act_buffer_inst_int_data7[16]), .A2(
        act_buffer_inst_n187), .B1(act_buffer_inst_int_data7[0]), .B2(
        act_buffer_inst_n181), .C1(act_buffer_inst_int_data7[8]), .C2(
        act_buffer_inst_n175), .ZN(act_buffer_inst_n47) );
  AOI222_X1 act_buffer_inst_U93 ( .A1(act_buffer_inst_int_data7[40]), .A2(
        act_buffer_inst_n169), .B1(act_buffer_inst_int_data7[24]), .B2(
        act_buffer_inst_n163), .C1(act_buffer_inst_int_data7[32]), .C2(
        act_buffer_inst_n8), .ZN(act_buffer_inst_n46) );
  NAND2_X1 act_buffer_inst_U92 ( .A1(act_buffer_inst_n46), .A2(
        act_buffer_inst_n47), .ZN(int_i_data_if7[0]) );
  INV_X1 act_buffer_inst_U91 ( .A(ps_int_ifmaps_ptr[1]), .ZN(
        act_buffer_inst_n190) );
  AND2_X1 act_buffer_inst_U90 ( .A1(ps_int_ifmaps_ptr[2]), .A2(
        act_buffer_inst_n189), .ZN(act_buffer_inst_n14) );
  AND2_X1 act_buffer_inst_U89 ( .A1(ps_int_ifmaps_ptr[2]), .A2(
        ps_int_ifmaps_ptr[0]), .ZN(act_buffer_inst_n13) );
  NOR2_X1 act_buffer_inst_U88 ( .A1(act_buffer_inst_n190), .A2(
        ps_int_ifmaps_ptr[0]), .ZN(act_buffer_inst_n16) );
  NOR2_X1 act_buffer_inst_U87 ( .A1(act_buffer_inst_n145), .A2(
        act_buffer_inst_n157), .ZN(act_buffer_inst_N120) );
  NOR2_X1 act_buffer_inst_U86 ( .A1(act_buffer_inst_n149), .A2(
        act_buffer_inst_n151), .ZN(act_buffer_inst_N152) );
  NOR2_X1 act_buffer_inst_U85 ( .A1(act_buffer_inst_n145), .A2(
        act_buffer_inst_n151), .ZN(act_buffer_inst_N156) );
  NOR2_X1 act_buffer_inst_U84 ( .A1(act_buffer_inst_n149), .A2(
        act_buffer_inst_n152), .ZN(act_buffer_inst_N146) );
  NOR2_X1 act_buffer_inst_U83 ( .A1(act_buffer_inst_n145), .A2(
        act_buffer_inst_n152), .ZN(act_buffer_inst_N150) );
  NOR2_X1 act_buffer_inst_U82 ( .A1(act_buffer_inst_n149), .A2(
        act_buffer_inst_n153), .ZN(act_buffer_inst_N140) );
  NOR2_X1 act_buffer_inst_U81 ( .A1(act_buffer_inst_n145), .A2(
        act_buffer_inst_n153), .ZN(act_buffer_inst_N144) );
  NOR2_X1 act_buffer_inst_U80 ( .A1(act_buffer_inst_n149), .A2(
        act_buffer_inst_n154), .ZN(act_buffer_inst_N134) );
  NOR2_X1 act_buffer_inst_U79 ( .A1(act_buffer_inst_n145), .A2(
        act_buffer_inst_n154), .ZN(act_buffer_inst_N138) );
  NOR2_X1 act_buffer_inst_U78 ( .A1(act_buffer_inst_n149), .A2(
        act_buffer_inst_n155), .ZN(act_buffer_inst_N128) );
  NOR2_X1 act_buffer_inst_U77 ( .A1(act_buffer_inst_n145), .A2(
        act_buffer_inst_n155), .ZN(act_buffer_inst_N132) );
  NOR2_X1 act_buffer_inst_U76 ( .A1(act_buffer_inst_n149), .A2(
        act_buffer_inst_n156), .ZN(act_buffer_inst_N122) );
  NOR2_X1 act_buffer_inst_U75 ( .A1(act_buffer_inst_n145), .A2(
        act_buffer_inst_n156), .ZN(act_buffer_inst_N126) );
  NOR2_X1 act_buffer_inst_U74 ( .A1(act_buffer_inst_n149), .A2(
        act_buffer_inst_n157), .ZN(act_buffer_inst_N116) );
  NOR2_X1 act_buffer_inst_U73 ( .A1(act_buffer_inst_n147), .A2(
        act_buffer_inst_n151), .ZN(act_buffer_inst_N154) );
  NOR2_X1 act_buffer_inst_U72 ( .A1(act_buffer_inst_n147), .A2(
        act_buffer_inst_n152), .ZN(act_buffer_inst_N148) );
  NOR2_X1 act_buffer_inst_U71 ( .A1(act_buffer_inst_n147), .A2(
        act_buffer_inst_n153), .ZN(act_buffer_inst_N142) );
  NOR2_X1 act_buffer_inst_U70 ( .A1(act_buffer_inst_n147), .A2(
        act_buffer_inst_n154), .ZN(act_buffer_inst_N136) );
  NOR2_X1 act_buffer_inst_U69 ( .A1(act_buffer_inst_n147), .A2(
        act_buffer_inst_n155), .ZN(act_buffer_inst_N130) );
  NOR2_X1 act_buffer_inst_U68 ( .A1(act_buffer_inst_n147), .A2(
        act_buffer_inst_n156), .ZN(act_buffer_inst_N124) );
  NOR2_X1 act_buffer_inst_U67 ( .A1(act_buffer_inst_n147), .A2(
        act_buffer_inst_n157), .ZN(act_buffer_inst_N118) );
  NOR2_X1 act_buffer_inst_U66 ( .A1(act_buffer_inst_n150), .A2(
        act_buffer_inst_n151), .ZN(act_buffer_inst_N151) );
  NOR2_X1 act_buffer_inst_U65 ( .A1(act_buffer_inst_n148), .A2(
        act_buffer_inst_n151), .ZN(act_buffer_inst_N153) );
  NOR2_X1 act_buffer_inst_U64 ( .A1(act_buffer_inst_n150), .A2(
        act_buffer_inst_n152), .ZN(act_buffer_inst_N145) );
  NOR2_X1 act_buffer_inst_U63 ( .A1(act_buffer_inst_n148), .A2(
        act_buffer_inst_n152), .ZN(act_buffer_inst_N147) );
  NOR2_X1 act_buffer_inst_U62 ( .A1(act_buffer_inst_n150), .A2(
        act_buffer_inst_n153), .ZN(act_buffer_inst_N139) );
  NOR2_X1 act_buffer_inst_U61 ( .A1(act_buffer_inst_n148), .A2(
        act_buffer_inst_n153), .ZN(act_buffer_inst_N141) );
  NOR2_X1 act_buffer_inst_U60 ( .A1(act_buffer_inst_n150), .A2(
        act_buffer_inst_n154), .ZN(act_buffer_inst_N133) );
  NOR2_X1 act_buffer_inst_U59 ( .A1(act_buffer_inst_n148), .A2(
        act_buffer_inst_n154), .ZN(act_buffer_inst_N135) );
  NOR2_X1 act_buffer_inst_U58 ( .A1(act_buffer_inst_n150), .A2(
        act_buffer_inst_n155), .ZN(act_buffer_inst_N127) );
  NOR2_X1 act_buffer_inst_U57 ( .A1(act_buffer_inst_n148), .A2(
        act_buffer_inst_n155), .ZN(act_buffer_inst_N129) );
  NOR2_X1 act_buffer_inst_U56 ( .A1(act_buffer_inst_n150), .A2(
        act_buffer_inst_n156), .ZN(act_buffer_inst_N121) );
  NOR2_X1 act_buffer_inst_U55 ( .A1(act_buffer_inst_n148), .A2(
        act_buffer_inst_n156), .ZN(act_buffer_inst_N123) );
  NOR2_X1 act_buffer_inst_U54 ( .A1(act_buffer_inst_n150), .A2(
        act_buffer_inst_n157), .ZN(act_buffer_inst_N115) );
  NOR2_X1 act_buffer_inst_U53 ( .A1(act_buffer_inst_n148), .A2(
        act_buffer_inst_n157), .ZN(act_buffer_inst_N117) );
  NOR2_X1 act_buffer_inst_U52 ( .A1(act_buffer_inst_n146), .A2(
        act_buffer_inst_n151), .ZN(act_buffer_inst_N155) );
  NOR2_X1 act_buffer_inst_U51 ( .A1(act_buffer_inst_n146), .A2(
        act_buffer_inst_n152), .ZN(act_buffer_inst_N149) );
  NOR2_X1 act_buffer_inst_U50 ( .A1(act_buffer_inst_n146), .A2(
        act_buffer_inst_n153), .ZN(act_buffer_inst_N143) );
  NOR2_X1 act_buffer_inst_U49 ( .A1(act_buffer_inst_n146), .A2(
        act_buffer_inst_n154), .ZN(act_buffer_inst_N137) );
  NOR2_X1 act_buffer_inst_U48 ( .A1(act_buffer_inst_n146), .A2(
        act_buffer_inst_n155), .ZN(act_buffer_inst_N131) );
  NOR2_X1 act_buffer_inst_U47 ( .A1(act_buffer_inst_n146), .A2(
        act_buffer_inst_n156), .ZN(act_buffer_inst_N125) );
  NOR2_X1 act_buffer_inst_U46 ( .A1(act_buffer_inst_n146), .A2(
        act_buffer_inst_n157), .ZN(act_buffer_inst_N119) );
  NOR2_X1 act_buffer_inst_U45 ( .A1(act_buffer_inst_n144), .A2(
        act_buffer_inst_n150), .ZN(act_buffer_inst_N157) );
  NOR2_X1 act_buffer_inst_U44 ( .A1(act_buffer_inst_n144), .A2(
        act_buffer_inst_n149), .ZN(act_buffer_inst_N158) );
  NOR2_X1 act_buffer_inst_U43 ( .A1(act_buffer_inst_n144), .A2(
        act_buffer_inst_n148), .ZN(act_buffer_inst_N159) );
  NOR2_X1 act_buffer_inst_U42 ( .A1(act_buffer_inst_n144), .A2(
        act_buffer_inst_n147), .ZN(act_buffer_inst_N160) );
  NOR2_X1 act_buffer_inst_U41 ( .A1(act_buffer_inst_n144), .A2(
        act_buffer_inst_n146), .ZN(act_buffer_inst_N161) );
  NOR2_X1 act_buffer_inst_U40 ( .A1(act_buffer_inst_n144), .A2(
        act_buffer_inst_n145), .ZN(act_buffer_inst_N162) );
  BUF_X1 act_buffer_inst_U39 ( .A(act_buffer_inst_n15), .Z(
        act_buffer_inst_n165) );
  BUF_X1 act_buffer_inst_U38 ( .A(act_buffer_inst_n15), .Z(
        act_buffer_inst_n168) );
  BUF_X1 act_buffer_inst_U37 ( .A(act_buffer_inst_n15), .Z(
        act_buffer_inst_n167) );
  BUF_X1 act_buffer_inst_U36 ( .A(act_buffer_inst_n15), .Z(
        act_buffer_inst_n166) );
  BUF_X1 act_buffer_inst_U35 ( .A(act_buffer_inst_n14), .Z(
        act_buffer_inst_n171) );
  BUF_X1 act_buffer_inst_U34 ( .A(act_buffer_inst_n17), .Z(act_buffer_inst_n4)
         );
  BUF_X1 act_buffer_inst_U33 ( .A(act_buffer_inst_n17), .Z(act_buffer_inst_n7)
         );
  BUF_X1 act_buffer_inst_U32 ( .A(act_buffer_inst_n17), .Z(act_buffer_inst_n6)
         );
  BUF_X1 act_buffer_inst_U31 ( .A(act_buffer_inst_n17), .Z(act_buffer_inst_n8)
         );
  BUF_X1 act_buffer_inst_U30 ( .A(act_buffer_inst_n17), .Z(act_buffer_inst_n5)
         );
  BUF_X1 act_buffer_inst_U29 ( .A(act_buffer_inst_n13), .Z(
        act_buffer_inst_n177) );
  BUF_X1 act_buffer_inst_U28 ( .A(act_buffer_inst_n13), .Z(
        act_buffer_inst_n179) );
  BUF_X1 act_buffer_inst_U27 ( .A(act_buffer_inst_n13), .Z(
        act_buffer_inst_n178) );
  BUF_X1 act_buffer_inst_U26 ( .A(act_buffer_inst_n16), .Z(
        act_buffer_inst_n159) );
  BUF_X1 act_buffer_inst_U25 ( .A(act_buffer_inst_n16), .Z(
        act_buffer_inst_n161) );
  BUF_X1 act_buffer_inst_U24 ( .A(act_buffer_inst_n16), .Z(
        act_buffer_inst_n160) );
  NOR2_X1 act_buffer_inst_U23 ( .A1(act_buffer_inst_n190), .A2(
        act_buffer_inst_n189), .ZN(act_buffer_inst_n12) );
  BUF_X1 act_buffer_inst_U22 ( .A(act_buffer_inst_n15), .Z(
        act_buffer_inst_n169) );
  BUF_X1 act_buffer_inst_U21 ( .A(act_buffer_inst_n14), .Z(
        act_buffer_inst_n174) );
  BUF_X1 act_buffer_inst_U20 ( .A(act_buffer_inst_n14), .Z(
        act_buffer_inst_n173) );
  BUF_X1 act_buffer_inst_U19 ( .A(act_buffer_inst_n14), .Z(
        act_buffer_inst_n175) );
  BUF_X1 act_buffer_inst_U18 ( .A(act_buffer_inst_n14), .Z(
        act_buffer_inst_n172) );
  BUF_X1 act_buffer_inst_U17 ( .A(act_buffer_inst_n13), .Z(
        act_buffer_inst_n180) );
  BUF_X1 act_buffer_inst_U16 ( .A(act_buffer_inst_n13), .Z(
        act_buffer_inst_n181) );
  BUF_X1 act_buffer_inst_U15 ( .A(act_buffer_inst_n16), .Z(
        act_buffer_inst_n162) );
  BUF_X1 act_buffer_inst_U14 ( .A(act_buffer_inst_n16), .Z(
        act_buffer_inst_n163) );
  AND4_X1 act_buffer_inst_U13 ( .A1(act_buffer_inst_n144), .A2(
        act_buffer_inst_n151), .A3(act_buffer_inst_n152), .A4(
        act_buffer_inst_n153), .ZN(act_buffer_inst_n158) );
  NAND4_X1 act_buffer_inst_U12 ( .A1(act_buffer_inst_n155), .A2(
        act_buffer_inst_n154), .A3(act_buffer_inst_n156), .A4(
        act_buffer_inst_n158), .ZN(act_buffer_inst_n157) );
  BUF_X1 act_buffer_inst_U11 ( .A(act_buffer_inst_n12), .Z(
        act_buffer_inst_n183) );
  BUF_X1 act_buffer_inst_U10 ( .A(act_buffer_inst_n12), .Z(
        act_buffer_inst_n186) );
  BUF_X1 act_buffer_inst_U9 ( .A(act_buffer_inst_n12), .Z(act_buffer_inst_n185) );
  BUF_X1 act_buffer_inst_U8 ( .A(act_buffer_inst_n12), .Z(act_buffer_inst_n187) );
  BUF_X1 act_buffer_inst_U7 ( .A(act_buffer_inst_n12), .Z(act_buffer_inst_n184) );
  INV_X8 act_buffer_inst_U6 ( .A(n9), .ZN(act_buffer_inst_n3) );
  INV_X8 act_buffer_inst_U5 ( .A(n9), .ZN(act_buffer_inst_n2) );
  INV_X8 act_buffer_inst_U4 ( .A(n9), .ZN(act_buffer_inst_n1) );
  NOR3_X1 act_buffer_inst_U3 ( .A1(ps_int_ifmaps_ptr[1]), .A2(
        ps_int_ifmaps_ptr[2]), .A3(ps_int_ifmaps_ptr[0]), .ZN(
        act_buffer_inst_n15) );
  NOR3_X1 act_buffer_inst_U2 ( .A1(ps_int_ifmaps_ptr[1]), .A2(
        ps_int_ifmaps_ptr[2]), .A3(act_buffer_inst_n189), .ZN(
        act_buffer_inst_n17) );
  DFFR_X1 act_buffer_inst_int_data1_reg_4__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4337), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data1[8]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_4__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4337), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data1[9]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_4__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4337), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data1[10]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_4__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4337), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data1[11]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_4__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4337), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data1[12]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_4__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4337), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data1[13]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_4__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4337), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data1[14]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_4__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4337), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data1[15]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_5__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4342), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data1[0]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_5__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4342), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data1[1]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_5__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4342), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data1[2]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_5__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4342), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data1[3]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_5__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4342), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data1[4]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_5__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4342), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data1[5]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_5__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4342), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data1[6]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_5__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4342), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data1[7]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_0__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4347), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data2[40]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_0__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4347), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data2[41]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_0__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4347), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data2[42]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_0__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4347), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data2[43]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_0__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4347), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data2[44]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_0__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4347), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data2[45]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_0__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4347), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data2[46]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_0__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4347), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data2[47]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_1__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4352), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data2[32]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_1__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4352), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data2[33]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_1__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4352), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data2[34]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_1__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4352), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data2[35]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_1__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4352), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data2[36]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_1__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4352), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data2[37]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_1__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4352), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data2[38]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_1__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4352), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data2[39]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_2__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4357), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data2[24]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_2__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4357), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data2[25]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_2__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4357), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data2[26]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_2__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4357), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data2[27]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_2__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4357), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data2[28]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_2__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4357), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data2[29]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_2__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4357), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data2[30]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_2__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4357), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data2[31]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_3__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4362), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data2[16]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_3__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4362), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data2[17]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_3__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4362), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data2[18]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_3__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4362), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data2[19]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_3__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4362), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data2[20]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_3__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4362), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data2[21]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_3__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4362), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data2[22]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_3__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4362), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data2[23]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_4__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4367), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data2[8]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_4__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4367), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data2[9]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_4__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4367), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data2[10]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_4__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4367), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data2[11]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_4__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4367), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data2[12]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_4__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4367), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data2[13]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_4__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4367), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data2[14]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_4__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4367), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data2[15]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_5__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4372), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data2[0]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_5__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4372), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data2[1]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_5__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4372), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data2[2]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_5__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4372), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data2[3]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_5__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4372), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data2[4]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_5__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4372), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data2[5]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_5__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4372), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data2[6]) );
  DFFR_X1 act_buffer_inst_int_data2_reg_5__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4372), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data2[7]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_0__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4377), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data3[40]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_0__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4377), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data3[41]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_0__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4377), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data3[42]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_0__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4377), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data3[43]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_0__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4377), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data3[44]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_0__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4377), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data3[45]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_0__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4377), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data3[46]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_0__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4377), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data3[47]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_1__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4382), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data3[32]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_1__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4382), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data3[33]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_1__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4382), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data3[34]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_1__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4382), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data3[35]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_1__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4382), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data3[36]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_1__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4382), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data3[37]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_1__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4382), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data3[38]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_1__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4382), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data3[39]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_2__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4387), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data3[24]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_2__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4387), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data3[25]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_2__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4387), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data3[26]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_2__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4387), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data3[27]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_2__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4387), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data3[28]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_2__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4387), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data3[29]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_2__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4387), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data3[30]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_2__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4387), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data3[31]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_3__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4392), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data3[16]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_3__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4392), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data3[17]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_3__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4392), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data3[18]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_3__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4392), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data3[19]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_3__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4392), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data3[20]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_3__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4392), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data3[21]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_3__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4392), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data3[22]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_3__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4392), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data3[23]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_4__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4397), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data3[8]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_4__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4397), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data3[9]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_4__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4397), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data3[10]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_4__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4397), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data3[11]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_4__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4397), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data3[12]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_4__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4397), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data3[13]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_4__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4397), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data3[14]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_4__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4397), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data3[15]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_5__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4402), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data3[0]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_5__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4402), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data3[1]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_5__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4402), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data3[2]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_5__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4402), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data3[3]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_5__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4402), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data3[4]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_5__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4402), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data3[5]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_5__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4402), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data3[6]) );
  DFFR_X1 act_buffer_inst_int_data3_reg_5__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4402), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data3[7]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_0__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4407), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data4[40]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_0__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4407), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data4[41]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_0__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4407), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data4[42]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_0__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4407), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data4[43]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_0__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4407), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data4[44]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_0__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4407), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data4[45]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_0__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4407), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data4[46]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_0__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4407), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data4[47]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_1__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4412), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data4[32]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_1__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4412), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data4[33]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_1__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4412), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data4[34]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_1__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4412), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data4[35]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_1__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4412), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data4[36]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_1__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4412), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data4[37]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_1__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4412), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data4[38]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_1__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4412), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data4[39]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_2__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4417), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data4[24]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_2__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4417), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data4[25]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_2__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4417), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data4[26]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_2__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4417), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data4[27]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_2__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4417), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data4[28]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_2__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4417), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data4[29]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_2__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4417), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data4[30]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_2__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4417), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data4[31]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_3__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4422), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data4[16]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_3__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4422), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data4[17]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_3__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4422), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data4[18]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_3__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4422), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data4[19]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_3__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4422), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data4[20]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_3__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4422), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data4[21]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_3__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4422), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data4[22]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_3__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4422), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data4[23]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_4__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4427), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data4[8]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_4__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4427), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data4[9]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_4__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4427), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data4[10]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_4__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4427), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data4[11]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_4__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4427), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data4[12]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_4__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4427), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data4[13]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_4__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4427), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data4[14]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_4__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4427), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data4[15]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_5__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4432), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data4[0]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_5__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4432), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data4[1]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_5__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4432), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data4[2]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_5__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4432), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data4[3]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_5__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4432), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data4[4]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_5__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4432), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data4[5]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_5__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4432), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data4[6]) );
  DFFR_X1 act_buffer_inst_int_data4_reg_5__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4432), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data4[7]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_0__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4437), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data5[40]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_0__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4437), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data5[41]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_0__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4437), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data5[42]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_0__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4437), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data5[43]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_0__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4437), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data5[44]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_0__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4437), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data5[45]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_0__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4437), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data5[46]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_0__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4437), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data5[47]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_1__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4442), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data5[32]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_1__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4442), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data5[33]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_1__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4442), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data5[34]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_1__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4442), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data5[35]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_1__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4442), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data5[36]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_1__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4442), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data5[37]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_1__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4442), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data5[38]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_1__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4442), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data5[39]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_2__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4447), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data5[24]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_2__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4447), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data5[25]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_2__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4447), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data5[26]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_2__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4447), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data5[27]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_2__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4447), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data5[28]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_2__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4447), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data5[29]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_2__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4447), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data5[30]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_2__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4447), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data5[31]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_3__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4452), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data5[16]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_3__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4452), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data5[17]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_3__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4452), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data5[18]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_3__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4452), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data5[19]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_3__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4452), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data5[20]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_3__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4452), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data5[21]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_3__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4452), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data5[22]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_3__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4452), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data5[23]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_4__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4457), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data5[8]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_4__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4457), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data5[9]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_4__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4457), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data5[10]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_4__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4457), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data5[11]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_4__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4457), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data5[12]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_4__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4457), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data5[13]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_4__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4457), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data5[14]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_4__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4457), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data5[15]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_5__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4462), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data5[0]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_5__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4462), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data5[1]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_5__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4462), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data5[2]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_5__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4462), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data5[3]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_5__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4462), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data5[4]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_5__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4462), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data5[5]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_5__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4462), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data5[6]) );
  DFFR_X1 act_buffer_inst_int_data5_reg_5__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4462), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data5[7]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_0__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4467), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data6[40]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_0__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4467), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data6[41]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_0__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4467), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data6[42]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_0__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4467), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data6[43]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_0__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4467), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data6[44]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_0__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4467), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data6[45]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_0__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4467), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data6[46]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_0__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4467), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data6[47]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_1__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4472), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data6[32]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_1__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4472), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data6[33]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_1__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4472), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data6[34]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_1__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4472), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data6[35]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_1__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4472), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data6[36]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_1__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4472), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data6[37]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_1__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4472), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data6[38]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_1__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4472), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data6[39]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_2__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4477), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data6[24]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_2__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4477), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data6[25]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_2__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4477), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data6[26]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_2__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4477), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data6[27]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_2__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4477), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data6[28]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_2__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4477), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data6[29]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_2__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4477), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data6[30]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_2__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4477), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data6[31]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_3__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4482), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data6[16]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_3__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4482), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data6[17]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_3__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4482), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data6[18]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_3__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4482), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data6[19]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_3__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4482), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data6[20]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_3__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4482), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data6[21]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_3__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4482), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data6[22]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_3__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4482), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data6[23]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_4__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4487), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data6[8]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_4__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4487), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data6[9]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_4__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4487), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data6[10]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_4__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4487), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data6[11]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_4__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4487), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data6[12]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_4__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4487), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data6[13]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_4__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4487), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data6[14]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_4__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4487), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data6[15]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_5__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4492), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data6[0]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_5__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4492), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data6[1]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_5__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4492), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data6[2]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_5__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4492), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data6[3]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_5__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4492), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data6[4]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_5__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4492), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data6[5]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_5__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4492), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data6[6]) );
  DFFR_X1 act_buffer_inst_int_data6_reg_5__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4492), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data6[7]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_0__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4497), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data7[40]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_0__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4497), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data7[41]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_0__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4497), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data7[42]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_0__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4497), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data7[43]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_0__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4497), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data7[44]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_0__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4497), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data7[45]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_0__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4497), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data7[46]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_0__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4497), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data7[47]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_1__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4502), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data7[32]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_1__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4502), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data7[33]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_1__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4502), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data7[34]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_1__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4502), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data7[35]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_1__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4502), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data7[36]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_1__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4502), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data7[37]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_1__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4502), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data7[38]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_1__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4502), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data7[39]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_2__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4507), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data7[24]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_2__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4507), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data7[25]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_2__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4507), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data7[26]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_2__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4507), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data7[27]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_2__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4507), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data7[28]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_2__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4507), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data7[29]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_2__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4507), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data7[30]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_2__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4507), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data7[31]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_3__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4512), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data7[16]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_3__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4512), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data7[17]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_3__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4512), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data7[18]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_3__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4512), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data7[19]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_3__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4512), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data7[20]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_3__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4512), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data7[21]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_3__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4512), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data7[22]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_3__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4512), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data7[23]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_4__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4517), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data7[8]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_4__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4517), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data7[9]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_4__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4517), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data7[10]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_4__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4517), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data7[11]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_4__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4517), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data7[12]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_4__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4517), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data7[13]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_4__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4517), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data7[14]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_4__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4517), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data7[15]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_5__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4522), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data7[0]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_5__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4522), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data7[1]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_5__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4522), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data7[2]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_5__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4522), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data7[3]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_5__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4522), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data7[4]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_5__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4522), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data7[5]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_5__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4522), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data7[6]) );
  DFFR_X1 act_buffer_inst_int_data7_reg_5__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4522), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data7[7]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_0__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4527), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data8[40]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_0__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4527), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data8[41]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_0__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4527), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data8[42]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_0__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4527), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data8[43]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_0__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4527), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data8[44]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_0__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4527), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data8[45]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_0__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4527), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data8[46]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_0__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4527), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data8[47]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_1__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4532), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data8[32]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_1__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4532), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data8[33]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_1__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4532), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data8[34]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_1__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4532), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data8[35]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_1__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4532), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data8[36]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_1__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4532), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data8[37]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_1__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4532), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data8[38]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_1__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4532), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data8[39]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_2__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4537), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data8[24]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_2__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4537), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data8[25]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_2__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4537), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data8[26]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_2__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4537), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data8[27]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_2__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4537), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data8[28]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_2__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4537), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data8[29]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_2__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4537), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data8[30]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_2__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4537), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data8[31]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_3__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4542), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data8[16]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_3__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4542), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data8[17]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_3__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4542), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data8[18]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_3__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4542), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data8[19]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_3__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4542), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data8[20]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_3__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4542), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data8[21]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_3__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4542), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data8[22]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_3__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4542), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data8[23]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_4__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4547), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data8[8]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_4__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4547), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data8[9]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_4__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4547), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data8[10]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_4__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4547), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data8[11]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_4__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4547), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data8[12]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_4__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4547), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data8[13]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_4__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4547), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data8[14]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_4__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4547), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data8[15]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_5__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4552), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data8[0]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_5__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4552), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data8[1]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_5__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4552), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data8[2]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_5__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4552), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data8[3]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_5__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4552), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data8[4]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_5__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4552), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data8[5]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_5__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4552), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data8[6]) );
  DFFR_X1 act_buffer_inst_int_data8_reg_5__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4552), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data8[7]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_0__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4316), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data1[40]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_0__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4316), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data1[41]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_0__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4316), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data1[42]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_0__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4316), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data1[43]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_0__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4316), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data1[44]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_0__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4316), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data1[45]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_0__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4316), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data1[46]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_0__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4316), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data1[47]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_1__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4322), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data1[32]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_1__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4322), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data1[33]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_1__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4322), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data1[34]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_1__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4322), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data1[35]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_1__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4322), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data1[36]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_1__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4322), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data1[37]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_1__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4322), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data1[38]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_1__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4322), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data1[39]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_2__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4327), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data1[24]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_2__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4327), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data1[25]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_2__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4327), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data1[26]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_2__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4327), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data1[27]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_2__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4327), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data1[28]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_2__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4327), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data1[29]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_2__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4327), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data1[30]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_2__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4327), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data1[31]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_3__0_ ( .D(i_acth[8]), .CK(
        act_buffer_inst_net4332), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data1[16]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_3__1_ ( .D(i_acth[9]), .CK(
        act_buffer_inst_net4332), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data1[17]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_3__2_ ( .D(i_acth[10]), .CK(
        act_buffer_inst_net4332), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data1[18]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_3__3_ ( .D(i_acth[11]), .CK(
        act_buffer_inst_net4332), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data1[19]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_3__4_ ( .D(i_acth[12]), .CK(
        act_buffer_inst_net4332), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data1[20]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_3__5_ ( .D(i_acth[13]), .CK(
        act_buffer_inst_net4332), .RN(act_buffer_inst_n1), .Q(
        act_buffer_inst_int_data1[21]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_3__6_ ( .D(i_acth[14]), .CK(
        act_buffer_inst_net4332), .RN(act_buffer_inst_n2), .Q(
        act_buffer_inst_int_data1[22]) );
  DFFR_X1 act_buffer_inst_int_data1_reg_3__7_ ( .D(i_acth[15]), .CK(
        act_buffer_inst_net4332), .RN(act_buffer_inst_n3), .Q(
        act_buffer_inst_int_data1[23]) );
  NAND3_X1 act_buffer_inst_U271 ( .A1(act_buffer_inst_n191), .A2(
        act_buffer_inst_n193), .A3(int_npu_ptr[1]), .ZN(act_buffer_inst_n155)
         );
  NAND3_X1 act_buffer_inst_U270 ( .A1(int_npu_ptr[0]), .A2(
        act_buffer_inst_n193), .A3(int_npu_ptr[1]), .ZN(act_buffer_inst_n154)
         );
  NAND3_X1 act_buffer_inst_U269 ( .A1(act_buffer_inst_n192), .A2(
        act_buffer_inst_n193), .A3(int_npu_ptr[0]), .ZN(act_buffer_inst_n156)
         );
  NAND3_X1 act_buffer_inst_U268 ( .A1(int_npu_ptr[1]), .A2(int_npu_ptr[0]), 
        .A3(int_npu_ptr[2]), .ZN(act_buffer_inst_n144) );
  NAND3_X1 act_buffer_inst_U267 ( .A1(int_npu_ptr[1]), .A2(
        act_buffer_inst_n191), .A3(int_npu_ptr[2]), .ZN(act_buffer_inst_n151)
         );
  NAND3_X1 act_buffer_inst_U266 ( .A1(int_npu_ptr[0]), .A2(
        act_buffer_inst_n192), .A3(int_npu_ptr[2]), .ZN(act_buffer_inst_n152)
         );
  NAND3_X1 act_buffer_inst_U265 ( .A1(act_buffer_inst_n191), .A2(
        act_buffer_inst_n192), .A3(int_npu_ptr[2]), .ZN(act_buffer_inst_n153)
         );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data1_reg_0__latch ( .CK(ck), .E(
        act_buffer_inst_N120), .SE(1'b0), .GCK(act_buffer_inst_net4316) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data1_reg_1__latch ( .CK(ck), .E(
        act_buffer_inst_N119), .SE(1'b0), .GCK(act_buffer_inst_net4322) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data1_reg_2__latch ( .CK(ck), .E(
        act_buffer_inst_N118), .SE(1'b0), .GCK(act_buffer_inst_net4327) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data1_reg_3__latch ( .CK(ck), .E(
        act_buffer_inst_N117), .SE(1'b0), .GCK(act_buffer_inst_net4332) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data1_reg_4__latch ( .CK(ck), .E(
        act_buffer_inst_N116), .SE(1'b0), .GCK(act_buffer_inst_net4337) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data1_reg_5__latch ( .CK(ck), .E(
        act_buffer_inst_N115), .SE(1'b0), .GCK(act_buffer_inst_net4342) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data2_reg_0__latch ( .CK(ck), .E(
        act_buffer_inst_N126), .SE(1'b0), .GCK(act_buffer_inst_net4347) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data2_reg_1__latch ( .CK(ck), .E(
        act_buffer_inst_N125), .SE(1'b0), .GCK(act_buffer_inst_net4352) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data2_reg_2__latch ( .CK(ck), .E(
        act_buffer_inst_N124), .SE(1'b0), .GCK(act_buffer_inst_net4357) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data2_reg_3__latch ( .CK(ck), .E(
        act_buffer_inst_N123), .SE(1'b0), .GCK(act_buffer_inst_net4362) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data2_reg_4__latch ( .CK(ck), .E(
        act_buffer_inst_N122), .SE(1'b0), .GCK(act_buffer_inst_net4367) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data2_reg_5__latch ( .CK(ck), .E(
        act_buffer_inst_N121), .SE(1'b0), .GCK(act_buffer_inst_net4372) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data3_reg_0__latch ( .CK(ck), .E(
        act_buffer_inst_N132), .SE(1'b0), .GCK(act_buffer_inst_net4377) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data3_reg_1__latch ( .CK(ck), .E(
        act_buffer_inst_N131), .SE(1'b0), .GCK(act_buffer_inst_net4382) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data3_reg_2__latch ( .CK(ck), .E(
        act_buffer_inst_N130), .SE(1'b0), .GCK(act_buffer_inst_net4387) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data3_reg_3__latch ( .CK(ck), .E(
        act_buffer_inst_N129), .SE(1'b0), .GCK(act_buffer_inst_net4392) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data3_reg_4__latch ( .CK(ck), .E(
        act_buffer_inst_N128), .SE(1'b0), .GCK(act_buffer_inst_net4397) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data3_reg_5__latch ( .CK(ck), .E(
        act_buffer_inst_N127), .SE(1'b0), .GCK(act_buffer_inst_net4402) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data4_reg_0__latch ( .CK(ck), .E(
        act_buffer_inst_N138), .SE(1'b0), .GCK(act_buffer_inst_net4407) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data4_reg_1__latch ( .CK(ck), .E(
        act_buffer_inst_N137), .SE(1'b0), .GCK(act_buffer_inst_net4412) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data4_reg_2__latch ( .CK(ck), .E(
        act_buffer_inst_N136), .SE(1'b0), .GCK(act_buffer_inst_net4417) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data4_reg_3__latch ( .CK(ck), .E(
        act_buffer_inst_N135), .SE(1'b0), .GCK(act_buffer_inst_net4422) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data4_reg_4__latch ( .CK(ck), .E(
        act_buffer_inst_N134), .SE(1'b0), .GCK(act_buffer_inst_net4427) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data4_reg_5__latch ( .CK(ck), .E(
        act_buffer_inst_N133), .SE(1'b0), .GCK(act_buffer_inst_net4432) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data5_reg_0__latch ( .CK(ck), .E(
        act_buffer_inst_N144), .SE(1'b0), .GCK(act_buffer_inst_net4437) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data5_reg_1__latch ( .CK(ck), .E(
        act_buffer_inst_N143), .SE(1'b0), .GCK(act_buffer_inst_net4442) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data5_reg_2__latch ( .CK(ck), .E(
        act_buffer_inst_N142), .SE(1'b0), .GCK(act_buffer_inst_net4447) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data5_reg_3__latch ( .CK(ck), .E(
        act_buffer_inst_N141), .SE(1'b0), .GCK(act_buffer_inst_net4452) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data5_reg_4__latch ( .CK(ck), .E(
        act_buffer_inst_N140), .SE(1'b0), .GCK(act_buffer_inst_net4457) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data5_reg_5__latch ( .CK(ck), .E(
        act_buffer_inst_N139), .SE(1'b0), .GCK(act_buffer_inst_net4462) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data6_reg_0__latch ( .CK(ck), .E(
        act_buffer_inst_N150), .SE(1'b0), .GCK(act_buffer_inst_net4467) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data6_reg_1__latch ( .CK(ck), .E(
        act_buffer_inst_N149), .SE(1'b0), .GCK(act_buffer_inst_net4472) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data6_reg_2__latch ( .CK(ck), .E(
        act_buffer_inst_N148), .SE(1'b0), .GCK(act_buffer_inst_net4477) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data6_reg_3__latch ( .CK(ck), .E(
        act_buffer_inst_N147), .SE(1'b0), .GCK(act_buffer_inst_net4482) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data6_reg_4__latch ( .CK(ck), .E(
        act_buffer_inst_N146), .SE(1'b0), .GCK(act_buffer_inst_net4487) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data6_reg_5__latch ( .CK(ck), .E(
        act_buffer_inst_N145), .SE(1'b0), .GCK(act_buffer_inst_net4492) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data7_reg_0__latch ( .CK(ck), .E(
        act_buffer_inst_N156), .SE(1'b0), .GCK(act_buffer_inst_net4497) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data7_reg_1__latch ( .CK(ck), .E(
        act_buffer_inst_N155), .SE(1'b0), .GCK(act_buffer_inst_net4502) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data7_reg_2__latch ( .CK(ck), .E(
        act_buffer_inst_N154), .SE(1'b0), .GCK(act_buffer_inst_net4507) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data7_reg_3__latch ( .CK(ck), .E(
        act_buffer_inst_N153), .SE(1'b0), .GCK(act_buffer_inst_net4512) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data7_reg_4__latch ( .CK(ck), .E(
        act_buffer_inst_N152), .SE(1'b0), .GCK(act_buffer_inst_net4517) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data7_reg_5__latch ( .CK(ck), .E(
        act_buffer_inst_N151), .SE(1'b0), .GCK(act_buffer_inst_net4522) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data8_reg_0__latch ( .CK(ck), .E(
        act_buffer_inst_N162), .SE(1'b0), .GCK(act_buffer_inst_net4527) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data8_reg_1__latch ( .CK(ck), .E(
        act_buffer_inst_N161), .SE(1'b0), .GCK(act_buffer_inst_net4532) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data8_reg_2__latch ( .CK(ck), .E(
        act_buffer_inst_N160), .SE(1'b0), .GCK(act_buffer_inst_net4537) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data8_reg_3__latch ( .CK(ck), .E(
        act_buffer_inst_N159), .SE(1'b0), .GCK(act_buffer_inst_net4542) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data8_reg_4__latch ( .CK(ck), .E(
        act_buffer_inst_N158), .SE(1'b0), .GCK(act_buffer_inst_net4547) );
  CLKGATETST_X1 act_buffer_inst_clk_gate_int_data8_reg_5__latch ( .CK(ck), .E(
        act_buffer_inst_N157), .SE(1'b0), .GCK(act_buffer_inst_net4552) );
  NOR3_X4 act_if_inst_U392 ( .A1(ps_int_hmode_cnt[0]), .A2(1'b0), .A3(
        act_if_inst_n312), .ZN(act_if_inst_n7) );
  CLKBUF_X1 act_if_inst_U391 ( .A(int_npu_ptr[0]), .Z(act_if_inst_n305) );
  CLKBUF_X1 act_if_inst_U390 ( .A(int_npu_ptr[1]), .Z(act_if_inst_n299) );
  CLKBUF_X1 act_if_inst_U389 ( .A(int_npu_ptr[2]), .Z(act_if_inst_n293) );
  MUX2_X1 act_if_inst_U388 ( .A(act_if_inst_n130), .B(act_if_inst_n131), .S(
        act_if_inst_n298), .Z(act_if_inst_n164) );
  MUX2_X1 act_if_inst_U387 ( .A(act_if_inst_n124), .B(act_if_inst_n125), .S(
        act_if_inst_n298), .Z(act_if_inst_n163) );
  MUX2_X1 act_if_inst_U386 ( .A(act_if_inst_n118), .B(act_if_inst_n119), .S(
        act_if_inst_n298), .Z(act_if_inst_n162) );
  MUX2_X1 act_if_inst_U385 ( .A(act_if_inst_n112), .B(act_if_inst_n113), .S(
        act_if_inst_n298), .Z(act_if_inst_n161) );
  MUX2_X1 act_if_inst_U384 ( .A(act_if_inst_n106), .B(act_if_inst_n107), .S(
        act_if_inst_n298), .Z(act_if_inst_n160) );
  MUX2_X1 act_if_inst_U383 ( .A(act_if_inst_n100), .B(act_if_inst_n101), .S(
        act_if_inst_n298), .Z(act_if_inst_n159) );
  MUX2_X1 act_if_inst_U382 ( .A(act_if_inst_n94), .B(act_if_inst_n95), .S(
        act_if_inst_n298), .Z(act_if_inst_n158) );
  MUX2_X1 act_if_inst_U381 ( .A(act_if_inst_n88), .B(act_if_inst_n89), .S(
        act_if_inst_n298), .Z(act_if_inst_n157) );
  MUX2_X1 act_if_inst_U380 ( .A(act_if_inst_n82), .B(act_if_inst_n83), .S(
        act_if_inst_n298), .Z(act_if_inst_n156) );
  MUX2_X1 act_if_inst_U379 ( .A(act_if_inst_n76), .B(act_if_inst_n77), .S(
        act_if_inst_n298), .Z(act_if_inst_n155) );
  MUX2_X1 act_if_inst_U378 ( .A(act_if_inst_n70), .B(act_if_inst_n71), .S(
        act_if_inst_n298), .Z(act_if_inst_n154) );
  MUX2_X1 act_if_inst_U377 ( .A(act_if_inst_n64), .B(act_if_inst_n65), .S(
        act_if_inst_n298), .Z(act_if_inst_n153) );
  MUX2_X1 act_if_inst_U376 ( .A(act_if_inst_n58), .B(act_if_inst_n59), .S(
        act_if_inst_n297), .Z(act_if_inst_n152) );
  MUX2_X1 act_if_inst_U375 ( .A(act_if_inst_n52), .B(act_if_inst_n53), .S(
        act_if_inst_n297), .Z(act_if_inst_n151) );
  MUX2_X1 act_if_inst_U374 ( .A(act_if_inst_n46), .B(act_if_inst_n47), .S(
        act_if_inst_n297), .Z(act_if_inst_n150) );
  MUX2_X1 act_if_inst_U373 ( .A(act_if_inst_n40), .B(act_if_inst_n41), .S(
        act_if_inst_n297), .Z(act_if_inst_n149) );
  MUX2_X1 act_if_inst_U372 ( .A(act_if_inst_n127), .B(act_if_inst_n128), .S(
        act_if_inst_n297), .Z(act_if_inst_n148) );
  MUX2_X1 act_if_inst_U371 ( .A(act_if_inst_n121), .B(act_if_inst_n122), .S(
        act_if_inst_n297), .Z(act_if_inst_n147) );
  MUX2_X1 act_if_inst_U370 ( .A(act_if_inst_n115), .B(act_if_inst_n116), .S(
        act_if_inst_n297), .Z(act_if_inst_n146) );
  MUX2_X1 act_if_inst_U369 ( .A(act_if_inst_n109), .B(act_if_inst_n110), .S(
        act_if_inst_n297), .Z(act_if_inst_n145) );
  MUX2_X1 act_if_inst_U368 ( .A(act_if_inst_n103), .B(act_if_inst_n104), .S(
        act_if_inst_n297), .Z(act_if_inst_n144) );
  MUX2_X1 act_if_inst_U367 ( .A(act_if_inst_n97), .B(act_if_inst_n98), .S(
        act_if_inst_n297), .Z(act_if_inst_n143) );
  MUX2_X1 act_if_inst_U366 ( .A(act_if_inst_n91), .B(act_if_inst_n92), .S(
        act_if_inst_n297), .Z(act_if_inst_n142) );
  MUX2_X1 act_if_inst_U365 ( .A(act_if_inst_n85), .B(act_if_inst_n86), .S(
        act_if_inst_n297), .Z(act_if_inst_n141) );
  MUX2_X1 act_if_inst_U364 ( .A(act_if_inst_n79), .B(act_if_inst_n80), .S(
        act_if_inst_n296), .Z(act_if_inst_n140) );
  MUX2_X1 act_if_inst_U363 ( .A(act_if_inst_n73), .B(act_if_inst_n74), .S(
        act_if_inst_n296), .Z(act_if_inst_n139) );
  MUX2_X1 act_if_inst_U362 ( .A(act_if_inst_n67), .B(act_if_inst_n68), .S(
        act_if_inst_n296), .Z(act_if_inst_n138) );
  MUX2_X1 act_if_inst_U361 ( .A(act_if_inst_n61), .B(act_if_inst_n62), .S(
        act_if_inst_n296), .Z(act_if_inst_n137) );
  MUX2_X1 act_if_inst_U360 ( .A(act_if_inst_n55), .B(act_if_inst_n56), .S(
        act_if_inst_n296), .Z(act_if_inst_n136) );
  MUX2_X1 act_if_inst_U359 ( .A(act_if_inst_n49), .B(act_if_inst_n50), .S(
        act_if_inst_n296), .Z(act_if_inst_n135) );
  MUX2_X1 act_if_inst_U358 ( .A(act_if_inst_n43), .B(act_if_inst_n44), .S(
        act_if_inst_n296), .Z(act_if_inst_n134) );
  MUX2_X1 act_if_inst_U357 ( .A(act_if_inst_n1), .B(act_if_inst_n2), .S(
        act_if_inst_n296), .Z(act_if_inst_n133) );
  MUX2_X1 act_if_inst_U356 ( .A(act_if_inst_n131), .B(act_if_inst_n130), .S(
        act_if_inst_n296), .Z(act_if_inst_n132) );
  MUX2_X1 act_if_inst_U355 ( .A(act_if_inst_n180), .B(act_if_inst_n172), .S(
        act_if_inst_n310), .Z(act_if_inst_n131) );
  MUX2_X1 act_if_inst_U354 ( .A(act_if_inst_n212), .B(act_if_inst_n204), .S(
        act_if_inst_n310), .Z(act_if_inst_n130) );
  MUX2_X1 act_if_inst_U353 ( .A(act_if_inst_n128), .B(act_if_inst_n127), .S(
        act_if_inst_n296), .Z(act_if_inst_n129) );
  MUX2_X1 act_if_inst_U352 ( .A(act_if_inst_n228), .B(act_if_inst_n220), .S(
        act_if_inst_n310), .Z(act_if_inst_n128) );
  MUX2_X1 act_if_inst_U351 ( .A(act_if_inst_n196), .B(act_if_inst_n188), .S(
        act_if_inst_n310), .Z(act_if_inst_n127) );
  MUX2_X1 act_if_inst_U350 ( .A(act_if_inst_n125), .B(act_if_inst_n124), .S(
        act_if_inst_n296), .Z(act_if_inst_n126) );
  MUX2_X1 act_if_inst_U349 ( .A(act_if_inst_n179), .B(act_if_inst_n171), .S(
        act_if_inst_n310), .Z(act_if_inst_n125) );
  MUX2_X1 act_if_inst_U348 ( .A(act_if_inst_n211), .B(act_if_inst_n203), .S(
        act_if_inst_n310), .Z(act_if_inst_n124) );
  MUX2_X1 act_if_inst_U347 ( .A(act_if_inst_n122), .B(act_if_inst_n121), .S(
        act_if_inst_n296), .Z(act_if_inst_n123) );
  MUX2_X1 act_if_inst_U346 ( .A(act_if_inst_n227), .B(act_if_inst_n219), .S(
        act_if_inst_n310), .Z(act_if_inst_n122) );
  MUX2_X1 act_if_inst_U345 ( .A(act_if_inst_n195), .B(act_if_inst_n187), .S(
        act_if_inst_n310), .Z(act_if_inst_n121) );
  MUX2_X1 act_if_inst_U344 ( .A(act_if_inst_n119), .B(act_if_inst_n118), .S(
        act_if_inst_n295), .Z(act_if_inst_n120) );
  MUX2_X1 act_if_inst_U343 ( .A(act_if_inst_n178), .B(act_if_inst_n170), .S(
        act_if_inst_n310), .Z(act_if_inst_n119) );
  MUX2_X1 act_if_inst_U342 ( .A(act_if_inst_n210), .B(act_if_inst_n202), .S(
        act_if_inst_n310), .Z(act_if_inst_n118) );
  MUX2_X1 act_if_inst_U341 ( .A(act_if_inst_n116), .B(act_if_inst_n115), .S(
        act_if_inst_n295), .Z(act_if_inst_n117) );
  MUX2_X1 act_if_inst_U340 ( .A(act_if_inst_n226), .B(act_if_inst_n218), .S(
        act_if_inst_n310), .Z(act_if_inst_n116) );
  MUX2_X1 act_if_inst_U339 ( .A(act_if_inst_n194), .B(act_if_inst_n186), .S(
        act_if_inst_n310), .Z(act_if_inst_n115) );
  MUX2_X1 act_if_inst_U338 ( .A(act_if_inst_n113), .B(act_if_inst_n112), .S(
        act_if_inst_n295), .Z(act_if_inst_n114) );
  MUX2_X1 act_if_inst_U337 ( .A(act_if_inst_n177), .B(act_if_inst_n169), .S(
        act_if_inst_n309), .Z(act_if_inst_n113) );
  MUX2_X1 act_if_inst_U336 ( .A(act_if_inst_n209), .B(act_if_inst_n201), .S(
        act_if_inst_n309), .Z(act_if_inst_n112) );
  MUX2_X1 act_if_inst_U335 ( .A(act_if_inst_n110), .B(act_if_inst_n109), .S(
        act_if_inst_n295), .Z(act_if_inst_n111) );
  MUX2_X1 act_if_inst_U334 ( .A(act_if_inst_n225), .B(act_if_inst_n217), .S(
        act_if_inst_n309), .Z(act_if_inst_n110) );
  MUX2_X1 act_if_inst_U333 ( .A(act_if_inst_n193), .B(act_if_inst_n185), .S(
        act_if_inst_n309), .Z(act_if_inst_n109) );
  MUX2_X1 act_if_inst_U332 ( .A(act_if_inst_n107), .B(act_if_inst_n106), .S(
        act_if_inst_n295), .Z(act_if_inst_n108) );
  MUX2_X1 act_if_inst_U331 ( .A(act_if_inst_n176), .B(act_if_inst_n168), .S(
        act_if_inst_n309), .Z(act_if_inst_n107) );
  MUX2_X1 act_if_inst_U330 ( .A(act_if_inst_n208), .B(act_if_inst_n200), .S(
        act_if_inst_n309), .Z(act_if_inst_n106) );
  MUX2_X1 act_if_inst_U329 ( .A(act_if_inst_n104), .B(act_if_inst_n103), .S(
        act_if_inst_n295), .Z(act_if_inst_n105) );
  MUX2_X1 act_if_inst_U328 ( .A(act_if_inst_n224), .B(act_if_inst_n216), .S(
        act_if_inst_n309), .Z(act_if_inst_n104) );
  MUX2_X1 act_if_inst_U327 ( .A(act_if_inst_n192), .B(act_if_inst_n184), .S(
        act_if_inst_n309), .Z(act_if_inst_n103) );
  MUX2_X1 act_if_inst_U326 ( .A(act_if_inst_n101), .B(act_if_inst_n100), .S(
        act_if_inst_n295), .Z(act_if_inst_n102) );
  MUX2_X1 act_if_inst_U325 ( .A(act_if_inst_n175), .B(act_if_inst_n167), .S(
        act_if_inst_n309), .Z(act_if_inst_n101) );
  MUX2_X1 act_if_inst_U324 ( .A(act_if_inst_n207), .B(act_if_inst_n199), .S(
        act_if_inst_n309), .Z(act_if_inst_n100) );
  MUX2_X1 act_if_inst_U323 ( .A(act_if_inst_n98), .B(act_if_inst_n97), .S(
        act_if_inst_n295), .Z(act_if_inst_n99) );
  MUX2_X1 act_if_inst_U322 ( .A(act_if_inst_n223), .B(act_if_inst_n215), .S(
        act_if_inst_n309), .Z(act_if_inst_n98) );
  MUX2_X1 act_if_inst_U321 ( .A(act_if_inst_n191), .B(act_if_inst_n183), .S(
        act_if_inst_n309), .Z(act_if_inst_n97) );
  MUX2_X1 act_if_inst_U320 ( .A(act_if_inst_n95), .B(act_if_inst_n94), .S(
        act_if_inst_n295), .Z(act_if_inst_n96) );
  MUX2_X1 act_if_inst_U319 ( .A(act_if_inst_n174), .B(act_if_inst_n166), .S(
        act_if_inst_n308), .Z(act_if_inst_n95) );
  MUX2_X1 act_if_inst_U318 ( .A(act_if_inst_n206), .B(act_if_inst_n198), .S(
        act_if_inst_n308), .Z(act_if_inst_n94) );
  MUX2_X1 act_if_inst_U317 ( .A(act_if_inst_n92), .B(act_if_inst_n91), .S(
        act_if_inst_n295), .Z(act_if_inst_n93) );
  MUX2_X1 act_if_inst_U316 ( .A(act_if_inst_n222), .B(act_if_inst_n214), .S(
        act_if_inst_n308), .Z(act_if_inst_n92) );
  MUX2_X1 act_if_inst_U315 ( .A(act_if_inst_n190), .B(act_if_inst_n182), .S(
        act_if_inst_n308), .Z(act_if_inst_n91) );
  MUX2_X1 act_if_inst_U314 ( .A(act_if_inst_n89), .B(act_if_inst_n88), .S(
        act_if_inst_n295), .Z(act_if_inst_n90) );
  MUX2_X1 act_if_inst_U313 ( .A(act_if_inst_n173), .B(act_if_inst_n165), .S(
        act_if_inst_n308), .Z(act_if_inst_n89) );
  MUX2_X1 act_if_inst_U312 ( .A(act_if_inst_n205), .B(act_if_inst_n197), .S(
        act_if_inst_n308), .Z(act_if_inst_n88) );
  MUX2_X1 act_if_inst_U311 ( .A(act_if_inst_n86), .B(act_if_inst_n85), .S(
        act_if_inst_n295), .Z(act_if_inst_n87) );
  MUX2_X1 act_if_inst_U310 ( .A(act_if_inst_n221), .B(act_if_inst_n213), .S(
        act_if_inst_n308), .Z(act_if_inst_n86) );
  MUX2_X1 act_if_inst_U309 ( .A(act_if_inst_n189), .B(act_if_inst_n181), .S(
        act_if_inst_n308), .Z(act_if_inst_n85) );
  MUX2_X1 act_if_inst_U308 ( .A(act_if_inst_n83), .B(act_if_inst_n82), .S(
        act_if_inst_n294), .Z(act_if_inst_n84) );
  MUX2_X1 act_if_inst_U307 ( .A(act_if_inst_n172), .B(act_if_inst_n228), .S(
        act_if_inst_n308), .Z(act_if_inst_n83) );
  MUX2_X1 act_if_inst_U306 ( .A(act_if_inst_n204), .B(act_if_inst_n196), .S(
        act_if_inst_n308), .Z(act_if_inst_n82) );
  MUX2_X1 act_if_inst_U305 ( .A(act_if_inst_n80), .B(act_if_inst_n79), .S(
        act_if_inst_n294), .Z(act_if_inst_n81) );
  MUX2_X1 act_if_inst_U304 ( .A(act_if_inst_n220), .B(act_if_inst_n212), .S(
        act_if_inst_n308), .Z(act_if_inst_n80) );
  MUX2_X1 act_if_inst_U303 ( .A(act_if_inst_n188), .B(act_if_inst_n180), .S(
        act_if_inst_n308), .Z(act_if_inst_n79) );
  MUX2_X1 act_if_inst_U302 ( .A(act_if_inst_n77), .B(act_if_inst_n76), .S(
        act_if_inst_n294), .Z(act_if_inst_n78) );
  MUX2_X1 act_if_inst_U301 ( .A(act_if_inst_n171), .B(act_if_inst_n227), .S(
        act_if_inst_n307), .Z(act_if_inst_n77) );
  MUX2_X1 act_if_inst_U300 ( .A(act_if_inst_n203), .B(act_if_inst_n195), .S(
        act_if_inst_n307), .Z(act_if_inst_n76) );
  MUX2_X1 act_if_inst_U299 ( .A(act_if_inst_n74), .B(act_if_inst_n73), .S(
        act_if_inst_n294), .Z(act_if_inst_n75) );
  MUX2_X1 act_if_inst_U298 ( .A(act_if_inst_n219), .B(act_if_inst_n211), .S(
        act_if_inst_n307), .Z(act_if_inst_n74) );
  MUX2_X1 act_if_inst_U297 ( .A(act_if_inst_n187), .B(act_if_inst_n179), .S(
        act_if_inst_n307), .Z(act_if_inst_n73) );
  MUX2_X1 act_if_inst_U296 ( .A(act_if_inst_n71), .B(act_if_inst_n70), .S(
        act_if_inst_n294), .Z(act_if_inst_n72) );
  MUX2_X1 act_if_inst_U295 ( .A(act_if_inst_n170), .B(act_if_inst_n226), .S(
        act_if_inst_n307), .Z(act_if_inst_n71) );
  MUX2_X1 act_if_inst_U294 ( .A(act_if_inst_n202), .B(act_if_inst_n194), .S(
        act_if_inst_n307), .Z(act_if_inst_n70) );
  MUX2_X1 act_if_inst_U293 ( .A(act_if_inst_n68), .B(act_if_inst_n67), .S(
        act_if_inst_n294), .Z(act_if_inst_n69) );
  MUX2_X1 act_if_inst_U292 ( .A(act_if_inst_n218), .B(act_if_inst_n210), .S(
        act_if_inst_n307), .Z(act_if_inst_n68) );
  MUX2_X1 act_if_inst_U291 ( .A(act_if_inst_n186), .B(act_if_inst_n178), .S(
        act_if_inst_n307), .Z(act_if_inst_n67) );
  MUX2_X1 act_if_inst_U290 ( .A(act_if_inst_n65), .B(act_if_inst_n64), .S(
        act_if_inst_n294), .Z(act_if_inst_n66) );
  MUX2_X1 act_if_inst_U289 ( .A(act_if_inst_n169), .B(act_if_inst_n225), .S(
        act_if_inst_n307), .Z(act_if_inst_n65) );
  MUX2_X1 act_if_inst_U288 ( .A(act_if_inst_n201), .B(act_if_inst_n193), .S(
        act_if_inst_n307), .Z(act_if_inst_n64) );
  MUX2_X1 act_if_inst_U287 ( .A(act_if_inst_n62), .B(act_if_inst_n61), .S(
        act_if_inst_n294), .Z(act_if_inst_n63) );
  MUX2_X1 act_if_inst_U286 ( .A(act_if_inst_n217), .B(act_if_inst_n209), .S(
        act_if_inst_n307), .Z(act_if_inst_n62) );
  MUX2_X1 act_if_inst_U285 ( .A(act_if_inst_n185), .B(act_if_inst_n177), .S(
        act_if_inst_n307), .Z(act_if_inst_n61) );
  MUX2_X1 act_if_inst_U284 ( .A(act_if_inst_n59), .B(act_if_inst_n58), .S(
        act_if_inst_n294), .Z(act_if_inst_n60) );
  MUX2_X1 act_if_inst_U283 ( .A(act_if_inst_n168), .B(act_if_inst_n224), .S(
        act_if_inst_n306), .Z(act_if_inst_n59) );
  MUX2_X1 act_if_inst_U282 ( .A(act_if_inst_n200), .B(act_if_inst_n192), .S(
        act_if_inst_n306), .Z(act_if_inst_n58) );
  MUX2_X1 act_if_inst_U281 ( .A(act_if_inst_n56), .B(act_if_inst_n55), .S(
        act_if_inst_n294), .Z(act_if_inst_n57) );
  MUX2_X1 act_if_inst_U280 ( .A(act_if_inst_n216), .B(act_if_inst_n208), .S(
        act_if_inst_n306), .Z(act_if_inst_n56) );
  MUX2_X1 act_if_inst_U279 ( .A(act_if_inst_n184), .B(act_if_inst_n176), .S(
        act_if_inst_n306), .Z(act_if_inst_n55) );
  MUX2_X1 act_if_inst_U278 ( .A(act_if_inst_n53), .B(act_if_inst_n52), .S(
        act_if_inst_n294), .Z(act_if_inst_n54) );
  MUX2_X1 act_if_inst_U277 ( .A(act_if_inst_n167), .B(act_if_inst_n223), .S(
        act_if_inst_n306), .Z(act_if_inst_n53) );
  MUX2_X1 act_if_inst_U276 ( .A(act_if_inst_n199), .B(act_if_inst_n191), .S(
        act_if_inst_n306), .Z(act_if_inst_n52) );
  MUX2_X1 act_if_inst_U275 ( .A(act_if_inst_n50), .B(act_if_inst_n49), .S(
        act_if_inst_n294), .Z(act_if_inst_n51) );
  MUX2_X1 act_if_inst_U274 ( .A(act_if_inst_n215), .B(act_if_inst_n207), .S(
        act_if_inst_n306), .Z(act_if_inst_n50) );
  MUX2_X1 act_if_inst_U273 ( .A(act_if_inst_n183), .B(act_if_inst_n175), .S(
        act_if_inst_n306), .Z(act_if_inst_n49) );
  MUX2_X1 act_if_inst_U272 ( .A(act_if_inst_n47), .B(act_if_inst_n46), .S(
        act_if_inst_n293), .Z(act_if_inst_n48) );
  MUX2_X1 act_if_inst_U271 ( .A(act_if_inst_n166), .B(act_if_inst_n222), .S(
        act_if_inst_n306), .Z(act_if_inst_n47) );
  MUX2_X1 act_if_inst_U270 ( .A(act_if_inst_n198), .B(act_if_inst_n190), .S(
        act_if_inst_n306), .Z(act_if_inst_n46) );
  MUX2_X1 act_if_inst_U269 ( .A(act_if_inst_n44), .B(act_if_inst_n43), .S(
        act_if_inst_n293), .Z(act_if_inst_n45) );
  MUX2_X1 act_if_inst_U268 ( .A(act_if_inst_n214), .B(act_if_inst_n206), .S(
        act_if_inst_n306), .Z(act_if_inst_n44) );
  MUX2_X1 act_if_inst_U267 ( .A(act_if_inst_n182), .B(act_if_inst_n174), .S(
        act_if_inst_n306), .Z(act_if_inst_n43) );
  MUX2_X1 act_if_inst_U266 ( .A(act_if_inst_n41), .B(act_if_inst_n40), .S(
        act_if_inst_n293), .Z(act_if_inst_n42) );
  MUX2_X1 act_if_inst_U265 ( .A(act_if_inst_n165), .B(act_if_inst_n221), .S(
        act_if_inst_n305), .Z(act_if_inst_n41) );
  MUX2_X1 act_if_inst_U264 ( .A(act_if_inst_n197), .B(act_if_inst_n189), .S(
        act_if_inst_n305), .Z(act_if_inst_n40) );
  MUX2_X1 act_if_inst_U263 ( .A(act_if_inst_n2), .B(act_if_inst_n1), .S(
        act_if_inst_n293), .Z(act_if_inst_n39) );
  MUX2_X1 act_if_inst_U262 ( .A(act_if_inst_n213), .B(act_if_inst_n205), .S(
        act_if_inst_n305), .Z(act_if_inst_n2) );
  MUX2_X1 act_if_inst_U261 ( .A(act_if_inst_n181), .B(act_if_inst_n173), .S(
        act_if_inst_n305), .Z(act_if_inst_n1) );
  MUX2_X1 act_if_inst_U260 ( .A(act_if_inst_n289), .B(act_if_inst_n292), .S(
        act_if_inst_n304), .Z(act_if_inst_int_data1[7]) );
  MUX2_X1 act_if_inst_U259 ( .A(act_if_inst_n285), .B(act_if_inst_n288), .S(
        act_if_inst_n304), .Z(act_if_inst_int_data1[6]) );
  MUX2_X1 act_if_inst_U258 ( .A(act_if_inst_n281), .B(act_if_inst_n284), .S(
        act_if_inst_n304), .Z(act_if_inst_int_data1[5]) );
  MUX2_X1 act_if_inst_U257 ( .A(act_if_inst_n277), .B(act_if_inst_n280), .S(
        act_if_inst_n304), .Z(act_if_inst_int_data1[4]) );
  MUX2_X1 act_if_inst_U256 ( .A(act_if_inst_n273), .B(act_if_inst_n276), .S(
        act_if_inst_n304), .Z(act_if_inst_int_data1[3]) );
  MUX2_X1 act_if_inst_U255 ( .A(act_if_inst_n269), .B(act_if_inst_n272), .S(
        act_if_inst_n304), .Z(act_if_inst_int_data1[2]) );
  MUX2_X1 act_if_inst_U254 ( .A(act_if_inst_n265), .B(act_if_inst_n268), .S(
        act_if_inst_n304), .Z(act_if_inst_int_data1[1]) );
  MUX2_X1 act_if_inst_U253 ( .A(act_if_inst_n261), .B(act_if_inst_n264), .S(
        act_if_inst_n304), .Z(act_if_inst_int_data1[0]) );
  MUX2_X1 act_if_inst_U252 ( .A(act_if_inst_n257), .B(act_if_inst_n260), .S(
        act_if_inst_n304), .Z(act_if_inst_int_data2[7]) );
  MUX2_X1 act_if_inst_U251 ( .A(act_if_inst_n253), .B(act_if_inst_n256), .S(
        act_if_inst_n304), .Z(act_if_inst_int_data2[6]) );
  MUX2_X1 act_if_inst_U250 ( .A(act_if_inst_n249), .B(act_if_inst_n252), .S(
        act_if_inst_n304), .Z(act_if_inst_int_data2[5]) );
  MUX2_X1 act_if_inst_U249 ( .A(act_if_inst_n245), .B(act_if_inst_n248), .S(
        act_if_inst_n304), .Z(act_if_inst_int_data2[4]) );
  MUX2_X1 act_if_inst_U248 ( .A(act_if_inst_n241), .B(act_if_inst_n244), .S(
        act_if_inst_n303), .Z(act_if_inst_int_data2[3]) );
  MUX2_X1 act_if_inst_U247 ( .A(act_if_inst_n237), .B(act_if_inst_n240), .S(
        act_if_inst_n303), .Z(act_if_inst_int_data2[2]) );
  MUX2_X1 act_if_inst_U246 ( .A(act_if_inst_n233), .B(act_if_inst_n236), .S(
        act_if_inst_n303), .Z(act_if_inst_int_data2[1]) );
  MUX2_X1 act_if_inst_U245 ( .A(act_if_inst_n229), .B(act_if_inst_n232), .S(
        act_if_inst_n303), .Z(act_if_inst_int_data2[0]) );
  MUX2_X1 act_if_inst_U244 ( .A(act_if_inst_n292), .B(act_if_inst_n290), .S(
        act_if_inst_n303), .Z(act_if_inst_int_data3[7]) );
  MUX2_X1 act_if_inst_U243 ( .A(act_if_inst_n288), .B(act_if_inst_n286), .S(
        act_if_inst_n303), .Z(act_if_inst_int_data3[6]) );
  MUX2_X1 act_if_inst_U242 ( .A(act_if_inst_n284), .B(act_if_inst_n282), .S(
        act_if_inst_n303), .Z(act_if_inst_int_data3[5]) );
  MUX2_X1 act_if_inst_U241 ( .A(act_if_inst_n280), .B(act_if_inst_n278), .S(
        act_if_inst_n303), .Z(act_if_inst_int_data3[4]) );
  MUX2_X1 act_if_inst_U240 ( .A(act_if_inst_n276), .B(act_if_inst_n274), .S(
        act_if_inst_n303), .Z(act_if_inst_int_data3[3]) );
  MUX2_X1 act_if_inst_U239 ( .A(act_if_inst_n272), .B(act_if_inst_n270), .S(
        act_if_inst_n303), .Z(act_if_inst_int_data3[2]) );
  MUX2_X1 act_if_inst_U238 ( .A(act_if_inst_n268), .B(act_if_inst_n266), .S(
        act_if_inst_n303), .Z(act_if_inst_int_data3[1]) );
  MUX2_X1 act_if_inst_U237 ( .A(act_if_inst_n264), .B(act_if_inst_n262), .S(
        act_if_inst_n303), .Z(act_if_inst_int_data3[0]) );
  MUX2_X1 act_if_inst_U236 ( .A(act_if_inst_n260), .B(act_if_inst_n258), .S(
        act_if_inst_n302), .Z(act_if_inst_int_data4[7]) );
  MUX2_X1 act_if_inst_U235 ( .A(act_if_inst_n256), .B(act_if_inst_n254), .S(
        act_if_inst_n302), .Z(act_if_inst_int_data4[6]) );
  MUX2_X1 act_if_inst_U234 ( .A(act_if_inst_n252), .B(act_if_inst_n250), .S(
        act_if_inst_n302), .Z(act_if_inst_int_data4[5]) );
  MUX2_X1 act_if_inst_U233 ( .A(act_if_inst_n248), .B(act_if_inst_n246), .S(
        act_if_inst_n302), .Z(act_if_inst_int_data4[4]) );
  MUX2_X1 act_if_inst_U232 ( .A(act_if_inst_n244), .B(act_if_inst_n242), .S(
        act_if_inst_n302), .Z(act_if_inst_int_data4[3]) );
  MUX2_X1 act_if_inst_U231 ( .A(act_if_inst_n240), .B(act_if_inst_n238), .S(
        act_if_inst_n302), .Z(act_if_inst_int_data4[2]) );
  MUX2_X1 act_if_inst_U230 ( .A(act_if_inst_n236), .B(act_if_inst_n234), .S(
        act_if_inst_n302), .Z(act_if_inst_int_data4[1]) );
  MUX2_X1 act_if_inst_U229 ( .A(act_if_inst_n232), .B(act_if_inst_n230), .S(
        act_if_inst_n302), .Z(act_if_inst_int_data4[0]) );
  MUX2_X1 act_if_inst_U228 ( .A(act_if_inst_n290), .B(act_if_inst_n291), .S(
        act_if_inst_n302), .Z(act_if_inst_int_data5[7]) );
  MUX2_X1 act_if_inst_U227 ( .A(act_if_inst_n286), .B(act_if_inst_n287), .S(
        act_if_inst_n302), .Z(act_if_inst_int_data5[6]) );
  MUX2_X1 act_if_inst_U226 ( .A(act_if_inst_n282), .B(act_if_inst_n283), .S(
        act_if_inst_n302), .Z(act_if_inst_int_data5[5]) );
  MUX2_X1 act_if_inst_U225 ( .A(act_if_inst_n278), .B(act_if_inst_n279), .S(
        act_if_inst_n302), .Z(act_if_inst_int_data5[4]) );
  MUX2_X1 act_if_inst_U224 ( .A(act_if_inst_n274), .B(act_if_inst_n275), .S(
        act_if_inst_n301), .Z(act_if_inst_int_data5[3]) );
  MUX2_X1 act_if_inst_U223 ( .A(act_if_inst_n270), .B(act_if_inst_n271), .S(
        act_if_inst_n301), .Z(act_if_inst_int_data5[2]) );
  MUX2_X1 act_if_inst_U222 ( .A(act_if_inst_n266), .B(act_if_inst_n267), .S(
        act_if_inst_n301), .Z(act_if_inst_int_data5[1]) );
  MUX2_X1 act_if_inst_U221 ( .A(act_if_inst_n262), .B(act_if_inst_n263), .S(
        act_if_inst_n301), .Z(act_if_inst_int_data5[0]) );
  MUX2_X1 act_if_inst_U220 ( .A(act_if_inst_n258), .B(act_if_inst_n259), .S(
        act_if_inst_n301), .Z(act_if_inst_int_data6[7]) );
  MUX2_X1 act_if_inst_U219 ( .A(act_if_inst_n254), .B(act_if_inst_n255), .S(
        act_if_inst_n301), .Z(act_if_inst_int_data6[6]) );
  MUX2_X1 act_if_inst_U218 ( .A(act_if_inst_n250), .B(act_if_inst_n251), .S(
        act_if_inst_n301), .Z(act_if_inst_int_data6[5]) );
  MUX2_X1 act_if_inst_U217 ( .A(act_if_inst_n246), .B(act_if_inst_n247), .S(
        act_if_inst_n301), .Z(act_if_inst_int_data6[4]) );
  MUX2_X1 act_if_inst_U216 ( .A(act_if_inst_n242), .B(act_if_inst_n243), .S(
        act_if_inst_n301), .Z(act_if_inst_int_data6[3]) );
  MUX2_X1 act_if_inst_U215 ( .A(act_if_inst_n238), .B(act_if_inst_n239), .S(
        act_if_inst_n301), .Z(act_if_inst_int_data6[2]) );
  MUX2_X1 act_if_inst_U214 ( .A(act_if_inst_n234), .B(act_if_inst_n235), .S(
        act_if_inst_n301), .Z(act_if_inst_int_data6[1]) );
  MUX2_X1 act_if_inst_U213 ( .A(act_if_inst_n230), .B(act_if_inst_n231), .S(
        act_if_inst_n301), .Z(act_if_inst_int_data6[0]) );
  MUX2_X1 act_if_inst_U212 ( .A(act_if_inst_n291), .B(act_if_inst_n289), .S(
        act_if_inst_n300), .Z(act_if_inst_int_data7[7]) );
  MUX2_X1 act_if_inst_U211 ( .A(act_if_inst_n287), .B(act_if_inst_n285), .S(
        act_if_inst_n300), .Z(act_if_inst_int_data7[6]) );
  MUX2_X1 act_if_inst_U210 ( .A(act_if_inst_n283), .B(act_if_inst_n281), .S(
        act_if_inst_n300), .Z(act_if_inst_int_data7[5]) );
  MUX2_X1 act_if_inst_U209 ( .A(act_if_inst_n279), .B(act_if_inst_n277), .S(
        act_if_inst_n300), .Z(act_if_inst_int_data7[4]) );
  MUX2_X1 act_if_inst_U208 ( .A(act_if_inst_n275), .B(act_if_inst_n273), .S(
        act_if_inst_n300), .Z(act_if_inst_int_data7[3]) );
  MUX2_X1 act_if_inst_U207 ( .A(act_if_inst_n271), .B(act_if_inst_n269), .S(
        act_if_inst_n300), .Z(act_if_inst_int_data7[2]) );
  MUX2_X1 act_if_inst_U206 ( .A(act_if_inst_n267), .B(act_if_inst_n265), .S(
        act_if_inst_n300), .Z(act_if_inst_int_data7[1]) );
  MUX2_X1 act_if_inst_U205 ( .A(act_if_inst_n263), .B(act_if_inst_n261), .S(
        act_if_inst_n300), .Z(act_if_inst_int_data7[0]) );
  MUX2_X1 act_if_inst_U204 ( .A(act_if_inst_n259), .B(act_if_inst_n257), .S(
        act_if_inst_n300), .Z(act_if_inst_int_data8[7]) );
  MUX2_X1 act_if_inst_U203 ( .A(act_if_inst_n255), .B(act_if_inst_n253), .S(
        act_if_inst_n300), .Z(act_if_inst_int_data8[6]) );
  MUX2_X1 act_if_inst_U202 ( .A(act_if_inst_n251), .B(act_if_inst_n249), .S(
        act_if_inst_n300), .Z(act_if_inst_int_data8[5]) );
  MUX2_X1 act_if_inst_U201 ( .A(act_if_inst_n247), .B(act_if_inst_n245), .S(
        act_if_inst_n300), .Z(act_if_inst_int_data8[4]) );
  MUX2_X1 act_if_inst_U200 ( .A(act_if_inst_n243), .B(act_if_inst_n241), .S(
        act_if_inst_n299), .Z(act_if_inst_int_data8[3]) );
  MUX2_X1 act_if_inst_U199 ( .A(act_if_inst_n239), .B(act_if_inst_n237), .S(
        act_if_inst_n299), .Z(act_if_inst_int_data8[2]) );
  MUX2_X1 act_if_inst_U198 ( .A(act_if_inst_n235), .B(act_if_inst_n233), .S(
        act_if_inst_n299), .Z(act_if_inst_int_data8[1]) );
  MUX2_X1 act_if_inst_U197 ( .A(act_if_inst_n231), .B(act_if_inst_n229), .S(
        act_if_inst_n299), .Z(act_if_inst_int_data8[0]) );
  INV_X1 act_if_inst_U196 ( .A(1'b0), .ZN(act_if_inst_n311) );
  INV_X1 act_if_inst_U195 ( .A(ps_int_hmode_cnt[1]), .ZN(act_if_inst_n312) );
  BUF_X1 act_if_inst_U194 ( .A(int_npu_ptr[0]), .Z(act_if_inst_n310) );
  BUF_X1 act_if_inst_U193 ( .A(int_npu_ptr[2]), .Z(act_if_inst_n295) );
  BUF_X1 act_if_inst_U192 ( .A(int_npu_ptr[2]), .Z(act_if_inst_n296) );
  BUF_X1 act_if_inst_U191 ( .A(int_npu_ptr[2]), .Z(act_if_inst_n294) );
  BUF_X1 act_if_inst_U190 ( .A(int_npu_ptr[2]), .Z(act_if_inst_n298) );
  BUF_X1 act_if_inst_U189 ( .A(int_npu_ptr[2]), .Z(act_if_inst_n297) );
  BUF_X1 act_if_inst_U188 ( .A(int_npu_ptr[1]), .Z(act_if_inst_n304) );
  BUF_X1 act_if_inst_U187 ( .A(int_npu_ptr[1]), .Z(act_if_inst_n303) );
  BUF_X1 act_if_inst_U186 ( .A(int_npu_ptr[1]), .Z(act_if_inst_n302) );
  BUF_X1 act_if_inst_U185 ( .A(int_npu_ptr[1]), .Z(act_if_inst_n301) );
  BUF_X1 act_if_inst_U184 ( .A(int_npu_ptr[1]), .Z(act_if_inst_n300) );
  BUF_X1 act_if_inst_U183 ( .A(int_npu_ptr[0]), .Z(act_if_inst_n309) );
  BUF_X1 act_if_inst_U182 ( .A(int_npu_ptr[0]), .Z(act_if_inst_n308) );
  BUF_X1 act_if_inst_U181 ( .A(int_npu_ptr[0]), .Z(act_if_inst_n306) );
  BUF_X1 act_if_inst_U180 ( .A(int_npu_ptr[0]), .Z(act_if_inst_n307) );
  INV_X1 act_if_inst_U179 ( .A(int_i_data_if1[3]), .ZN(act_if_inst_n224) );
  INV_X1 act_if_inst_U178 ( .A(int_i_data_if2[3]), .ZN(act_if_inst_n216) );
  INV_X1 act_if_inst_U177 ( .A(int_i_data_if5[3]), .ZN(act_if_inst_n192) );
  INV_X1 act_if_inst_U176 ( .A(int_i_data_if3[3]), .ZN(act_if_inst_n208) );
  INV_X1 act_if_inst_U175 ( .A(int_i_data_if4[3]), .ZN(act_if_inst_n200) );
  INV_X1 act_if_inst_U174 ( .A(int_i_data_if1[5]), .ZN(act_if_inst_n226) );
  INV_X1 act_if_inst_U173 ( .A(int_i_data_if2[5]), .ZN(act_if_inst_n218) );
  INV_X1 act_if_inst_U172 ( .A(int_i_data_if3[5]), .ZN(act_if_inst_n210) );
  INV_X1 act_if_inst_U171 ( .A(int_i_data_if4[5]), .ZN(act_if_inst_n202) );
  INV_X1 act_if_inst_U170 ( .A(int_i_data_if1[7]), .ZN(act_if_inst_n228) );
  INV_X1 act_if_inst_U169 ( .A(int_i_data_if2[7]), .ZN(act_if_inst_n220) );
  INV_X1 act_if_inst_U168 ( .A(int_i_data_if3[7]), .ZN(act_if_inst_n212) );
  INV_X1 act_if_inst_U167 ( .A(int_i_data_if4[7]), .ZN(act_if_inst_n204) );
  INV_X1 act_if_inst_U166 ( .A(int_i_data_if1[1]), .ZN(act_if_inst_n222) );
  INV_X1 act_if_inst_U165 ( .A(int_i_data_if2[1]), .ZN(act_if_inst_n214) );
  INV_X1 act_if_inst_U164 ( .A(int_i_data_if5[1]), .ZN(act_if_inst_n190) );
  INV_X1 act_if_inst_U163 ( .A(int_i_data_if3[1]), .ZN(act_if_inst_n206) );
  INV_X1 act_if_inst_U162 ( .A(int_i_data_if4[1]), .ZN(act_if_inst_n198) );
  INV_X1 act_if_inst_U161 ( .A(int_i_data_if1[2]), .ZN(act_if_inst_n223) );
  INV_X1 act_if_inst_U160 ( .A(int_i_data_if2[2]), .ZN(act_if_inst_n215) );
  INV_X1 act_if_inst_U159 ( .A(int_i_data_if5[2]), .ZN(act_if_inst_n191) );
  INV_X1 act_if_inst_U158 ( .A(int_i_data_if3[2]), .ZN(act_if_inst_n207) );
  INV_X1 act_if_inst_U157 ( .A(int_i_data_if4[2]), .ZN(act_if_inst_n199) );
  INV_X1 act_if_inst_U156 ( .A(int_i_data_if1[4]), .ZN(act_if_inst_n225) );
  INV_X1 act_if_inst_U155 ( .A(int_i_data_if2[4]), .ZN(act_if_inst_n217) );
  INV_X1 act_if_inst_U154 ( .A(int_i_data_if3[4]), .ZN(act_if_inst_n209) );
  INV_X1 act_if_inst_U153 ( .A(int_i_data_if4[4]), .ZN(act_if_inst_n201) );
  INV_X1 act_if_inst_U152 ( .A(int_i_data_if1[6]), .ZN(act_if_inst_n227) );
  INV_X1 act_if_inst_U151 ( .A(int_i_data_if2[6]), .ZN(act_if_inst_n219) );
  INV_X1 act_if_inst_U150 ( .A(int_i_data_if3[6]), .ZN(act_if_inst_n211) );
  INV_X1 act_if_inst_U149 ( .A(int_i_data_if4[6]), .ZN(act_if_inst_n203) );
  INV_X1 act_if_inst_U148 ( .A(int_i_data_if1[0]), .ZN(act_if_inst_n221) );
  INV_X1 act_if_inst_U147 ( .A(int_i_data_if2[0]), .ZN(act_if_inst_n213) );
  INV_X1 act_if_inst_U146 ( .A(int_i_data_if5[0]), .ZN(act_if_inst_n189) );
  INV_X1 act_if_inst_U145 ( .A(int_i_data_if4[0]), .ZN(act_if_inst_n197) );
  INV_X1 act_if_inst_U144 ( .A(int_i_data_if3[0]), .ZN(act_if_inst_n205) );
  INV_X1 act_if_inst_U143 ( .A(int_i_data_if6[3]), .ZN(act_if_inst_n184) );
  INV_X1 act_if_inst_U142 ( .A(int_i_data_if7[3]), .ZN(act_if_inst_n176) );
  INV_X1 act_if_inst_U141 ( .A(int_i_data_if8[3]), .ZN(act_if_inst_n168) );
  INV_X1 act_if_inst_U140 ( .A(int_i_data_if5[5]), .ZN(act_if_inst_n194) );
  INV_X1 act_if_inst_U139 ( .A(int_i_data_if6[5]), .ZN(act_if_inst_n186) );
  INV_X1 act_if_inst_U138 ( .A(int_i_data_if8[5]), .ZN(act_if_inst_n170) );
  INV_X1 act_if_inst_U137 ( .A(int_i_data_if7[5]), .ZN(act_if_inst_n178) );
  INV_X1 act_if_inst_U136 ( .A(int_i_data_if5[7]), .ZN(act_if_inst_n196) );
  INV_X1 act_if_inst_U135 ( .A(int_i_data_if6[7]), .ZN(act_if_inst_n188) );
  INV_X1 act_if_inst_U134 ( .A(int_i_data_if8[7]), .ZN(act_if_inst_n172) );
  INV_X1 act_if_inst_U133 ( .A(int_i_data_if7[7]), .ZN(act_if_inst_n180) );
  INV_X1 act_if_inst_U132 ( .A(int_i_data_if6[1]), .ZN(act_if_inst_n182) );
  INV_X1 act_if_inst_U131 ( .A(int_i_data_if7[1]), .ZN(act_if_inst_n174) );
  INV_X1 act_if_inst_U130 ( .A(int_i_data_if8[1]), .ZN(act_if_inst_n166) );
  INV_X1 act_if_inst_U129 ( .A(int_i_data_if6[2]), .ZN(act_if_inst_n183) );
  INV_X1 act_if_inst_U128 ( .A(int_i_data_if7[2]), .ZN(act_if_inst_n175) );
  INV_X1 act_if_inst_U127 ( .A(int_i_data_if8[2]), .ZN(act_if_inst_n167) );
  INV_X1 act_if_inst_U126 ( .A(int_i_data_if6[4]), .ZN(act_if_inst_n185) );
  INV_X1 act_if_inst_U125 ( .A(int_i_data_if5[4]), .ZN(act_if_inst_n193) );
  INV_X1 act_if_inst_U124 ( .A(int_i_data_if8[4]), .ZN(act_if_inst_n169) );
  INV_X1 act_if_inst_U123 ( .A(int_i_data_if7[4]), .ZN(act_if_inst_n177) );
  INV_X1 act_if_inst_U122 ( .A(int_i_data_if5[6]), .ZN(act_if_inst_n195) );
  INV_X1 act_if_inst_U121 ( .A(int_i_data_if6[6]), .ZN(act_if_inst_n187) );
  INV_X1 act_if_inst_U120 ( .A(int_i_data_if8[6]), .ZN(act_if_inst_n171) );
  INV_X1 act_if_inst_U119 ( .A(int_i_data_if7[6]), .ZN(act_if_inst_n179) );
  INV_X1 act_if_inst_U118 ( .A(int_i_data_if6[0]), .ZN(act_if_inst_n181) );
  INV_X1 act_if_inst_U117 ( .A(int_i_data_if8[0]), .ZN(act_if_inst_n165) );
  INV_X1 act_if_inst_U116 ( .A(int_i_data_if7[0]), .ZN(act_if_inst_n173) );
  AOI22_X1 act_if_inst_U115 ( .A1(act_if_inst_int_data8[7]), .A2(
        act_if_inst_n5), .B1(act_if_inst_int_data8[1]), .B2(act_if_inst_n6), 
        .ZN(act_if_inst_n4) );
  AOI22_X1 act_if_inst_U114 ( .A1(act_if_inst_int_data8[3]), .A2(
        act_if_inst_n7), .B1(act_if_inst_int_data8[5]), .B2(act_if_inst_n8), 
        .ZN(act_if_inst_n3) );
  NAND2_X1 act_if_inst_U113 ( .A1(act_if_inst_n3), .A2(act_if_inst_n4), .ZN(
        int_i_data_h_npu8[1]) );
  AOI22_X1 act_if_inst_U112 ( .A1(act_if_inst_int_data8[6]), .A2(
        act_if_inst_n5), .B1(act_if_inst_int_data8[0]), .B2(act_if_inst_n6), 
        .ZN(act_if_inst_n10) );
  AOI22_X1 act_if_inst_U111 ( .A1(act_if_inst_int_data8[2]), .A2(
        act_if_inst_n7), .B1(act_if_inst_int_data8[4]), .B2(act_if_inst_n8), 
        .ZN(act_if_inst_n9) );
  NAND2_X1 act_if_inst_U110 ( .A1(act_if_inst_n9), .A2(act_if_inst_n10), .ZN(
        int_i_data_h_npu8[0]) );
  INV_X1 act_if_inst_U109 ( .A(act_if_inst_n105), .ZN(act_if_inst_n273) );
  INV_X1 act_if_inst_U108 ( .A(act_if_inst_n160), .ZN(act_if_inst_n276) );
  INV_X1 act_if_inst_U107 ( .A(act_if_inst_n117), .ZN(act_if_inst_n281) );
  INV_X1 act_if_inst_U106 ( .A(act_if_inst_n162), .ZN(act_if_inst_n284) );
  INV_X1 act_if_inst_U105 ( .A(act_if_inst_n129), .ZN(act_if_inst_n289) );
  INV_X1 act_if_inst_U104 ( .A(act_if_inst_n164), .ZN(act_if_inst_n292) );
  INV_X1 act_if_inst_U103 ( .A(act_if_inst_n93), .ZN(act_if_inst_n265) );
  INV_X1 act_if_inst_U102 ( .A(act_if_inst_n158), .ZN(act_if_inst_n268) );
  INV_X1 act_if_inst_U101 ( .A(act_if_inst_n99), .ZN(act_if_inst_n269) );
  INV_X1 act_if_inst_U100 ( .A(act_if_inst_n159), .ZN(act_if_inst_n272) );
  INV_X1 act_if_inst_U99 ( .A(act_if_inst_n111), .ZN(act_if_inst_n277) );
  INV_X1 act_if_inst_U98 ( .A(act_if_inst_n161), .ZN(act_if_inst_n280) );
  INV_X1 act_if_inst_U97 ( .A(act_if_inst_n123), .ZN(act_if_inst_n285) );
  INV_X1 act_if_inst_U96 ( .A(act_if_inst_n163), .ZN(act_if_inst_n288) );
  INV_X1 act_if_inst_U95 ( .A(act_if_inst_n87), .ZN(act_if_inst_n261) );
  INV_X1 act_if_inst_U94 ( .A(act_if_inst_n157), .ZN(act_if_inst_n264) );
  INV_X1 act_if_inst_U93 ( .A(act_if_inst_n57), .ZN(act_if_inst_n241) );
  INV_X1 act_if_inst_U92 ( .A(act_if_inst_n152), .ZN(act_if_inst_n244) );
  INV_X1 act_if_inst_U91 ( .A(act_if_inst_n69), .ZN(act_if_inst_n249) );
  INV_X1 act_if_inst_U90 ( .A(act_if_inst_n154), .ZN(act_if_inst_n252) );
  INV_X1 act_if_inst_U89 ( .A(act_if_inst_n81), .ZN(act_if_inst_n257) );
  INV_X1 act_if_inst_U88 ( .A(act_if_inst_n156), .ZN(act_if_inst_n260) );
  INV_X1 act_if_inst_U87 ( .A(act_if_inst_n45), .ZN(act_if_inst_n233) );
  INV_X1 act_if_inst_U86 ( .A(act_if_inst_n150), .ZN(act_if_inst_n236) );
  INV_X1 act_if_inst_U85 ( .A(act_if_inst_n51), .ZN(act_if_inst_n237) );
  INV_X1 act_if_inst_U84 ( .A(act_if_inst_n151), .ZN(act_if_inst_n240) );
  INV_X1 act_if_inst_U83 ( .A(act_if_inst_n63), .ZN(act_if_inst_n245) );
  INV_X1 act_if_inst_U82 ( .A(act_if_inst_n153), .ZN(act_if_inst_n248) );
  INV_X1 act_if_inst_U81 ( .A(act_if_inst_n75), .ZN(act_if_inst_n253) );
  INV_X1 act_if_inst_U80 ( .A(act_if_inst_n155), .ZN(act_if_inst_n256) );
  INV_X1 act_if_inst_U79 ( .A(act_if_inst_n39), .ZN(act_if_inst_n229) );
  INV_X1 act_if_inst_U78 ( .A(act_if_inst_n149), .ZN(act_if_inst_n232) );
  INV_X1 act_if_inst_U77 ( .A(act_if_inst_n144), .ZN(act_if_inst_n274) );
  INV_X1 act_if_inst_U76 ( .A(act_if_inst_n146), .ZN(act_if_inst_n282) );
  INV_X1 act_if_inst_U75 ( .A(act_if_inst_n148), .ZN(act_if_inst_n290) );
  INV_X1 act_if_inst_U74 ( .A(act_if_inst_n142), .ZN(act_if_inst_n266) );
  INV_X1 act_if_inst_U73 ( .A(act_if_inst_n143), .ZN(act_if_inst_n270) );
  INV_X1 act_if_inst_U72 ( .A(act_if_inst_n145), .ZN(act_if_inst_n278) );
  INV_X1 act_if_inst_U71 ( .A(act_if_inst_n147), .ZN(act_if_inst_n286) );
  INV_X1 act_if_inst_U70 ( .A(act_if_inst_n141), .ZN(act_if_inst_n262) );
  INV_X1 act_if_inst_U69 ( .A(act_if_inst_n136), .ZN(act_if_inst_n242) );
  INV_X1 act_if_inst_U68 ( .A(act_if_inst_n138), .ZN(act_if_inst_n250) );
  INV_X1 act_if_inst_U67 ( .A(act_if_inst_n140), .ZN(act_if_inst_n258) );
  INV_X1 act_if_inst_U66 ( .A(act_if_inst_n134), .ZN(act_if_inst_n234) );
  INV_X1 act_if_inst_U65 ( .A(act_if_inst_n135), .ZN(act_if_inst_n238) );
  INV_X1 act_if_inst_U64 ( .A(act_if_inst_n137), .ZN(act_if_inst_n246) );
  INV_X1 act_if_inst_U63 ( .A(act_if_inst_n139), .ZN(act_if_inst_n254) );
  INV_X1 act_if_inst_U62 ( .A(act_if_inst_n133), .ZN(act_if_inst_n230) );
  INV_X1 act_if_inst_U61 ( .A(act_if_inst_n108), .ZN(act_if_inst_n275) );
  INV_X1 act_if_inst_U60 ( .A(act_if_inst_n120), .ZN(act_if_inst_n283) );
  INV_X1 act_if_inst_U59 ( .A(act_if_inst_n132), .ZN(act_if_inst_n291) );
  INV_X1 act_if_inst_U58 ( .A(act_if_inst_n96), .ZN(act_if_inst_n267) );
  INV_X1 act_if_inst_U57 ( .A(act_if_inst_n102), .ZN(act_if_inst_n271) );
  INV_X1 act_if_inst_U56 ( .A(act_if_inst_n114), .ZN(act_if_inst_n279) );
  INV_X1 act_if_inst_U55 ( .A(act_if_inst_n126), .ZN(act_if_inst_n287) );
  INV_X1 act_if_inst_U54 ( .A(act_if_inst_n90), .ZN(act_if_inst_n263) );
  INV_X1 act_if_inst_U53 ( .A(act_if_inst_n60), .ZN(act_if_inst_n243) );
  INV_X1 act_if_inst_U52 ( .A(act_if_inst_n72), .ZN(act_if_inst_n251) );
  INV_X1 act_if_inst_U51 ( .A(act_if_inst_n84), .ZN(act_if_inst_n259) );
  INV_X1 act_if_inst_U50 ( .A(act_if_inst_n48), .ZN(act_if_inst_n235) );
  INV_X1 act_if_inst_U49 ( .A(act_if_inst_n54), .ZN(act_if_inst_n239) );
  INV_X1 act_if_inst_U48 ( .A(act_if_inst_n66), .ZN(act_if_inst_n247) );
  INV_X1 act_if_inst_U47 ( .A(act_if_inst_n78), .ZN(act_if_inst_n255) );
  INV_X1 act_if_inst_U46 ( .A(act_if_inst_n42), .ZN(act_if_inst_n231) );
  AOI22_X1 act_if_inst_U45 ( .A1(act_if_inst_int_data1[7]), .A2(act_if_inst_n5), .B1(act_if_inst_int_data1[1]), .B2(act_if_inst_n6), .ZN(act_if_inst_n36) );
  AOI22_X1 act_if_inst_U44 ( .A1(act_if_inst_int_data1[3]), .A2(act_if_inst_n7), .B1(act_if_inst_int_data1[5]), .B2(act_if_inst_n8), .ZN(act_if_inst_n35) );
  NAND2_X1 act_if_inst_U43 ( .A1(act_if_inst_n35), .A2(act_if_inst_n36), .ZN(
        int_i_data_h_npu1[1]) );
  AOI22_X1 act_if_inst_U42 ( .A1(act_if_inst_int_data1[6]), .A2(act_if_inst_n5), .B1(act_if_inst_int_data1[0]), .B2(act_if_inst_n6), .ZN(act_if_inst_n38) );
  AOI22_X1 act_if_inst_U41 ( .A1(act_if_inst_int_data1[2]), .A2(act_if_inst_n7), .B1(act_if_inst_int_data1[4]), .B2(act_if_inst_n8), .ZN(act_if_inst_n37) );
  NAND2_X1 act_if_inst_U40 ( .A1(act_if_inst_n37), .A2(act_if_inst_n38), .ZN(
        int_i_data_h_npu1[0]) );
  AOI22_X1 act_if_inst_U39 ( .A1(act_if_inst_int_data2[7]), .A2(act_if_inst_n5), .B1(act_if_inst_int_data2[1]), .B2(act_if_inst_n6), .ZN(act_if_inst_n32) );
  AOI22_X1 act_if_inst_U38 ( .A1(act_if_inst_int_data2[3]), .A2(act_if_inst_n7), .B1(act_if_inst_int_data2[5]), .B2(act_if_inst_n8), .ZN(act_if_inst_n31) );
  NAND2_X1 act_if_inst_U37 ( .A1(act_if_inst_n31), .A2(act_if_inst_n32), .ZN(
        int_i_data_h_npu2[1]) );
  AOI22_X1 act_if_inst_U36 ( .A1(act_if_inst_int_data3[7]), .A2(act_if_inst_n5), .B1(act_if_inst_int_data3[1]), .B2(act_if_inst_n6), .ZN(act_if_inst_n28) );
  AOI22_X1 act_if_inst_U35 ( .A1(act_if_inst_int_data3[3]), .A2(act_if_inst_n7), .B1(act_if_inst_int_data3[5]), .B2(act_if_inst_n8), .ZN(act_if_inst_n27) );
  NAND2_X1 act_if_inst_U34 ( .A1(act_if_inst_n27), .A2(act_if_inst_n28), .ZN(
        int_i_data_h_npu3[1]) );
  AOI22_X1 act_if_inst_U33 ( .A1(act_if_inst_int_data3[6]), .A2(act_if_inst_n5), .B1(act_if_inst_int_data3[0]), .B2(act_if_inst_n6), .ZN(act_if_inst_n30) );
  AOI22_X1 act_if_inst_U32 ( .A1(act_if_inst_int_data3[2]), .A2(act_if_inst_n7), .B1(act_if_inst_int_data3[4]), .B2(act_if_inst_n8), .ZN(act_if_inst_n29) );
  NAND2_X1 act_if_inst_U31 ( .A1(act_if_inst_n29), .A2(act_if_inst_n30), .ZN(
        int_i_data_h_npu3[0]) );
  AOI22_X1 act_if_inst_U30 ( .A1(act_if_inst_int_data2[6]), .A2(act_if_inst_n5), .B1(act_if_inst_int_data2[0]), .B2(act_if_inst_n6), .ZN(act_if_inst_n34) );
  AOI22_X1 act_if_inst_U29 ( .A1(act_if_inst_int_data2[2]), .A2(act_if_inst_n7), .B1(act_if_inst_int_data2[4]), .B2(act_if_inst_n8), .ZN(act_if_inst_n33) );
  NAND2_X1 act_if_inst_U28 ( .A1(act_if_inst_n33), .A2(act_if_inst_n34), .ZN(
        int_i_data_h_npu2[0]) );
  AOI22_X1 act_if_inst_U27 ( .A1(act_if_inst_int_data4[7]), .A2(act_if_inst_n5), .B1(act_if_inst_int_data4[1]), .B2(act_if_inst_n6), .ZN(act_if_inst_n24) );
  AOI22_X1 act_if_inst_U26 ( .A1(act_if_inst_int_data4[3]), .A2(act_if_inst_n7), .B1(act_if_inst_int_data4[5]), .B2(act_if_inst_n8), .ZN(act_if_inst_n23) );
  NAND2_X1 act_if_inst_U25 ( .A1(act_if_inst_n23), .A2(act_if_inst_n24), .ZN(
        int_i_data_h_npu4[1]) );
  AOI22_X1 act_if_inst_U24 ( .A1(act_if_inst_int_data4[6]), .A2(act_if_inst_n5), .B1(act_if_inst_int_data4[0]), .B2(act_if_inst_n6), .ZN(act_if_inst_n26) );
  AOI22_X1 act_if_inst_U23 ( .A1(act_if_inst_int_data4[2]), .A2(act_if_inst_n7), .B1(act_if_inst_int_data4[4]), .B2(act_if_inst_n8), .ZN(act_if_inst_n25) );
  NAND2_X1 act_if_inst_U22 ( .A1(act_if_inst_n25), .A2(act_if_inst_n26), .ZN(
        int_i_data_h_npu4[0]) );
  AOI22_X1 act_if_inst_U21 ( .A1(act_if_inst_int_data5[7]), .A2(act_if_inst_n5), .B1(act_if_inst_int_data5[1]), .B2(act_if_inst_n6), .ZN(act_if_inst_n20) );
  AOI22_X1 act_if_inst_U20 ( .A1(act_if_inst_int_data5[3]), .A2(act_if_inst_n7), .B1(act_if_inst_int_data5[5]), .B2(act_if_inst_n8), .ZN(act_if_inst_n19) );
  NAND2_X1 act_if_inst_U19 ( .A1(act_if_inst_n19), .A2(act_if_inst_n20), .ZN(
        int_i_data_h_npu5[1]) );
  AOI22_X1 act_if_inst_U18 ( .A1(act_if_inst_int_data5[6]), .A2(act_if_inst_n5), .B1(act_if_inst_int_data5[0]), .B2(act_if_inst_n6), .ZN(act_if_inst_n22) );
  AOI22_X1 act_if_inst_U17 ( .A1(act_if_inst_int_data5[2]), .A2(act_if_inst_n7), .B1(act_if_inst_int_data5[4]), .B2(act_if_inst_n8), .ZN(act_if_inst_n21) );
  NAND2_X1 act_if_inst_U16 ( .A1(act_if_inst_n21), .A2(act_if_inst_n22), .ZN(
        int_i_data_h_npu5[0]) );
  AOI22_X1 act_if_inst_U15 ( .A1(act_if_inst_int_data6[7]), .A2(act_if_inst_n5), .B1(act_if_inst_int_data6[1]), .B2(act_if_inst_n6), .ZN(act_if_inst_n16) );
  AOI22_X1 act_if_inst_U14 ( .A1(act_if_inst_int_data6[3]), .A2(act_if_inst_n7), .B1(act_if_inst_int_data6[5]), .B2(act_if_inst_n8), .ZN(act_if_inst_n15) );
  NAND2_X1 act_if_inst_U13 ( .A1(act_if_inst_n15), .A2(act_if_inst_n16), .ZN(
        int_i_data_h_npu6[1]) );
  AOI22_X1 act_if_inst_U12 ( .A1(act_if_inst_int_data6[6]), .A2(act_if_inst_n5), .B1(act_if_inst_int_data6[0]), .B2(act_if_inst_n6), .ZN(act_if_inst_n18) );
  AOI22_X1 act_if_inst_U11 ( .A1(act_if_inst_int_data6[2]), .A2(act_if_inst_n7), .B1(act_if_inst_int_data6[4]), .B2(act_if_inst_n8), .ZN(act_if_inst_n17) );
  NAND2_X1 act_if_inst_U10 ( .A1(act_if_inst_n17), .A2(act_if_inst_n18), .ZN(
        int_i_data_h_npu6[0]) );
  AOI22_X1 act_if_inst_U9 ( .A1(act_if_inst_int_data7[7]), .A2(act_if_inst_n5), 
        .B1(act_if_inst_int_data7[1]), .B2(act_if_inst_n6), .ZN(
        act_if_inst_n12) );
  AOI22_X1 act_if_inst_U8 ( .A1(act_if_inst_int_data7[3]), .A2(act_if_inst_n7), 
        .B1(act_if_inst_int_data7[5]), .B2(act_if_inst_n8), .ZN(
        act_if_inst_n11) );
  NAND2_X1 act_if_inst_U7 ( .A1(act_if_inst_n11), .A2(act_if_inst_n12), .ZN(
        int_i_data_h_npu7[1]) );
  AOI22_X1 act_if_inst_U6 ( .A1(act_if_inst_int_data7[6]), .A2(act_if_inst_n5), 
        .B1(act_if_inst_int_data7[0]), .B2(act_if_inst_n6), .ZN(
        act_if_inst_n14) );
  AOI22_X1 act_if_inst_U5 ( .A1(act_if_inst_int_data7[2]), .A2(act_if_inst_n7), 
        .B1(act_if_inst_int_data7[4]), .B2(act_if_inst_n8), .ZN(
        act_if_inst_n13) );
  NAND2_X1 act_if_inst_U4 ( .A1(act_if_inst_n13), .A2(act_if_inst_n14), .ZN(
        int_i_data_h_npu7[0]) );
  AND3_X1 act_if_inst_U3 ( .A1(act_if_inst_n312), .A2(act_if_inst_n311), .A3(
        ps_int_hmode_cnt[0]), .ZN(act_if_inst_n8) );
  AND3_X1 act_if_inst_U2 ( .A1(ps_int_hmode_cnt[0]), .A2(act_if_inst_n311), 
        .A3(ps_int_hmode_cnt[1]), .ZN(act_if_inst_n6) );
  NOR3_X4 act_if_inst_U1 ( .A1(act_if_inst_n7), .A2(act_if_inst_n8), .A3(
        act_if_inst_n6), .ZN(act_if_inst_n5) );
  CLKBUF_X1 npu_inst_U207 ( .A(i_weight[1]), .Z(npu_inst_n119) );
  CLKBUF_X1 npu_inst_U206 ( .A(i_weight[0]), .Z(npu_inst_n113) );
  CLKBUF_X1 npu_inst_U205 ( .A(ps_int_ifmaps_ptr[0]), .Z(npu_inst_n72) );
  INV_X1 npu_inst_U204 ( .A(1'b0), .ZN(npu_inst_n129) );
  INV_X1 npu_inst_U203 ( .A(1'b0), .ZN(npu_inst_n128) );
  NAND2_X1 npu_inst_U202 ( .A1(npu_inst_n129), .A2(npu_inst_n128), .ZN(
        npu_inst_int_ckg[63]) );
  NAND2_X1 npu_inst_U201 ( .A1(npu_inst_n143), .A2(npu_inst_n128), .ZN(
        npu_inst_int_ckg[31]) );
  NAND2_X1 npu_inst_U200 ( .A1(npu_inst_n143), .A2(npu_inst_n138), .ZN(
        npu_inst_int_ckg[27]) );
  BUF_X1 npu_inst_U199 ( .A(ps_ctrl_wr_pipe), .Z(npu_inst_n5) );
  BUF_X1 npu_inst_U198 ( .A(ps_ctrl_ldh_v_n), .Z(npu_inst_n51) );
  BUF_X1 npu_inst_U197 ( .A(ps_ctrl_ldh_v_n), .Z(npu_inst_n50) );
  NAND2_X1 npu_inst_U196 ( .A1(npu_inst_n129), .A2(npu_inst_n138), .ZN(
        npu_inst_int_ckg[59]) );
  BUF_X1 npu_inst_U195 ( .A(ps_ctrl_en_npu), .Z(npu_inst_n66) );
  BUF_X1 npu_inst_U194 ( .A(ps_ctrl_en_npu), .Z(npu_inst_n61) );
  BUF_X1 npu_inst_U193 ( .A(ps_ctrl_en_npu), .Z(npu_inst_n62) );
  BUF_X1 npu_inst_U192 ( .A(ps_ctrl_en_npu), .Z(npu_inst_n63) );
  BUF_X1 npu_inst_U191 ( .A(ps_ctrl_en_npu), .Z(npu_inst_n64) );
  BUF_X1 npu_inst_U190 ( .A(ps_ctrl_en_npu), .Z(npu_inst_n65) );
  BUF_X1 npu_inst_U189 ( .A(i_weight[1]), .Z(npu_inst_n118) );
  BUF_X1 npu_inst_U188 ( .A(i_weight[0]), .Z(npu_inst_n112) );
  BUF_X1 npu_inst_U187 ( .A(i_weight[1]), .Z(npu_inst_n117) );
  BUF_X1 npu_inst_U186 ( .A(i_weight[0]), .Z(npu_inst_n111) );
  BUF_X1 npu_inst_U185 ( .A(i_weight[1]), .Z(npu_inst_n116) );
  BUF_X1 npu_inst_U184 ( .A(i_weight[0]), .Z(npu_inst_n110) );
  BUF_X1 npu_inst_U183 ( .A(i_weight[1]), .Z(npu_inst_n115) );
  BUF_X1 npu_inst_U182 ( .A(i_weight[0]), .Z(npu_inst_n109) );
  BUF_X1 npu_inst_U181 ( .A(i_weight[1]), .Z(npu_inst_n114) );
  BUF_X1 npu_inst_U180 ( .A(i_weight[0]), .Z(npu_inst_n108) );
  INV_X1 npu_inst_U179 ( .A(int_ckg_rmask[4]), .ZN(npu_inst_n143) );
  INV_X1 npu_inst_U178 ( .A(int_ckg_cmask[4]), .ZN(npu_inst_n138) );
  NAND2_X1 npu_inst_U177 ( .A1(npu_inst_n129), .A2(npu_inst_n130), .ZN(
        npu_inst_int_ckg[62]) );
  NAND2_X1 npu_inst_U176 ( .A1(npu_inst_n129), .A2(npu_inst_n136), .ZN(
        npu_inst_int_ckg[61]) );
  NAND2_X1 npu_inst_U175 ( .A1(npu_inst_n129), .A2(npu_inst_n134), .ZN(
        npu_inst_int_ckg[60]) );
  NAND2_X1 npu_inst_U174 ( .A1(npu_inst_n129), .A2(npu_inst_n139), .ZN(
        npu_inst_int_ckg[58]) );
  NAND2_X1 npu_inst_U173 ( .A1(npu_inst_n129), .A2(npu_inst_n140), .ZN(
        npu_inst_int_ckg[57]) );
  NAND2_X1 npu_inst_U172 ( .A1(npu_inst_n129), .A2(npu_inst_n131), .ZN(
        npu_inst_int_ckg[56]) );
  NAND2_X1 npu_inst_U171 ( .A1(npu_inst_n133), .A2(npu_inst_n128), .ZN(
        npu_inst_int_ckg[55]) );
  NAND2_X1 npu_inst_U170 ( .A1(npu_inst_n133), .A2(npu_inst_n130), .ZN(
        npu_inst_int_ckg[54]) );
  NAND2_X1 npu_inst_U169 ( .A1(npu_inst_n133), .A2(npu_inst_n136), .ZN(
        npu_inst_int_ckg[53]) );
  NAND2_X1 npu_inst_U168 ( .A1(npu_inst_n133), .A2(npu_inst_n134), .ZN(
        npu_inst_int_ckg[52]) );
  NAND2_X1 npu_inst_U167 ( .A1(npu_inst_n133), .A2(npu_inst_n138), .ZN(
        npu_inst_int_ckg[51]) );
  NAND2_X1 npu_inst_U166 ( .A1(npu_inst_n133), .A2(npu_inst_n139), .ZN(
        npu_inst_int_ckg[50]) );
  NAND2_X1 npu_inst_U165 ( .A1(npu_inst_n133), .A2(npu_inst_n140), .ZN(
        npu_inst_int_ckg[49]) );
  NAND2_X1 npu_inst_U164 ( .A1(npu_inst_n133), .A2(npu_inst_n131), .ZN(
        npu_inst_int_ckg[48]) );
  NAND2_X1 npu_inst_U163 ( .A1(npu_inst_n137), .A2(npu_inst_n128), .ZN(
        npu_inst_int_ckg[47]) );
  NAND2_X1 npu_inst_U162 ( .A1(npu_inst_n137), .A2(npu_inst_n130), .ZN(
        npu_inst_int_ckg[46]) );
  NAND2_X1 npu_inst_U161 ( .A1(npu_inst_n137), .A2(npu_inst_n136), .ZN(
        npu_inst_int_ckg[45]) );
  NAND2_X1 npu_inst_U160 ( .A1(npu_inst_n137), .A2(npu_inst_n134), .ZN(
        npu_inst_int_ckg[44]) );
  NAND2_X1 npu_inst_U159 ( .A1(npu_inst_n137), .A2(npu_inst_n138), .ZN(
        npu_inst_int_ckg[43]) );
  NAND2_X1 npu_inst_U158 ( .A1(npu_inst_n137), .A2(npu_inst_n139), .ZN(
        npu_inst_int_ckg[42]) );
  NAND2_X1 npu_inst_U157 ( .A1(npu_inst_n137), .A2(npu_inst_n140), .ZN(
        npu_inst_int_ckg[41]) );
  NAND2_X1 npu_inst_U156 ( .A1(npu_inst_n137), .A2(npu_inst_n131), .ZN(
        npu_inst_int_ckg[40]) );
  NAND2_X1 npu_inst_U155 ( .A1(npu_inst_n135), .A2(npu_inst_n128), .ZN(
        npu_inst_int_ckg[39]) );
  NAND2_X1 npu_inst_U154 ( .A1(npu_inst_n135), .A2(npu_inst_n130), .ZN(
        npu_inst_int_ckg[38]) );
  NAND2_X1 npu_inst_U153 ( .A1(npu_inst_n135), .A2(npu_inst_n136), .ZN(
        npu_inst_int_ckg[37]) );
  NAND2_X1 npu_inst_U152 ( .A1(npu_inst_n135), .A2(npu_inst_n134), .ZN(
        npu_inst_int_ckg[36]) );
  NAND2_X1 npu_inst_U151 ( .A1(npu_inst_n135), .A2(npu_inst_n138), .ZN(
        npu_inst_int_ckg[35]) );
  NAND2_X1 npu_inst_U150 ( .A1(npu_inst_n135), .A2(npu_inst_n139), .ZN(
        npu_inst_int_ckg[34]) );
  NAND2_X1 npu_inst_U149 ( .A1(npu_inst_n135), .A2(npu_inst_n140), .ZN(
        npu_inst_int_ckg[33]) );
  NAND2_X1 npu_inst_U148 ( .A1(npu_inst_n135), .A2(npu_inst_n131), .ZN(
        npu_inst_int_ckg[32]) );
  NAND2_X1 npu_inst_U147 ( .A1(npu_inst_n143), .A2(npu_inst_n130), .ZN(
        npu_inst_int_ckg[30]) );
  NAND2_X1 npu_inst_U146 ( .A1(npu_inst_n143), .A2(npu_inst_n136), .ZN(
        npu_inst_int_ckg[29]) );
  NAND2_X1 npu_inst_U145 ( .A1(npu_inst_n143), .A2(npu_inst_n134), .ZN(
        npu_inst_int_ckg[28]) );
  NAND2_X1 npu_inst_U144 ( .A1(npu_inst_n143), .A2(npu_inst_n139), .ZN(
        npu_inst_int_ckg[26]) );
  NAND2_X1 npu_inst_U143 ( .A1(npu_inst_n143), .A2(npu_inst_n140), .ZN(
        npu_inst_int_ckg[25]) );
  NAND2_X1 npu_inst_U142 ( .A1(npu_inst_n143), .A2(npu_inst_n131), .ZN(
        npu_inst_int_ckg[24]) );
  NAND2_X1 npu_inst_U141 ( .A1(npu_inst_n141), .A2(npu_inst_n128), .ZN(
        npu_inst_int_ckg[23]) );
  NAND2_X1 npu_inst_U140 ( .A1(npu_inst_n141), .A2(npu_inst_n130), .ZN(
        npu_inst_int_ckg[22]) );
  NAND2_X1 npu_inst_U139 ( .A1(npu_inst_n141), .A2(npu_inst_n136), .ZN(
        npu_inst_int_ckg[21]) );
  NAND2_X1 npu_inst_U138 ( .A1(npu_inst_n141), .A2(npu_inst_n134), .ZN(
        npu_inst_int_ckg[20]) );
  NAND2_X1 npu_inst_U137 ( .A1(npu_inst_n141), .A2(npu_inst_n138), .ZN(
        npu_inst_int_ckg[19]) );
  NAND2_X1 npu_inst_U136 ( .A1(npu_inst_n141), .A2(npu_inst_n139), .ZN(
        npu_inst_int_ckg[18]) );
  NAND2_X1 npu_inst_U135 ( .A1(npu_inst_n141), .A2(npu_inst_n140), .ZN(
        npu_inst_int_ckg[17]) );
  NAND2_X1 npu_inst_U134 ( .A1(npu_inst_n141), .A2(npu_inst_n131), .ZN(
        npu_inst_int_ckg[16]) );
  NAND2_X1 npu_inst_U133 ( .A1(npu_inst_n142), .A2(npu_inst_n128), .ZN(
        npu_inst_int_ckg[15]) );
  NAND2_X1 npu_inst_U132 ( .A1(npu_inst_n142), .A2(npu_inst_n130), .ZN(
        npu_inst_int_ckg[14]) );
  NAND2_X1 npu_inst_U131 ( .A1(npu_inst_n142), .A2(npu_inst_n136), .ZN(
        npu_inst_int_ckg[13]) );
  NAND2_X1 npu_inst_U130 ( .A1(npu_inst_n142), .A2(npu_inst_n134), .ZN(
        npu_inst_int_ckg[12]) );
  NAND2_X1 npu_inst_U129 ( .A1(npu_inst_n142), .A2(npu_inst_n138), .ZN(
        npu_inst_int_ckg[11]) );
  NAND2_X1 npu_inst_U128 ( .A1(npu_inst_n142), .A2(npu_inst_n139), .ZN(
        npu_inst_int_ckg[10]) );
  NAND2_X1 npu_inst_U127 ( .A1(npu_inst_n142), .A2(npu_inst_n140), .ZN(
        npu_inst_int_ckg[9]) );
  NAND2_X1 npu_inst_U126 ( .A1(npu_inst_n142), .A2(npu_inst_n131), .ZN(
        npu_inst_int_ckg[8]) );
  NAND2_X1 npu_inst_U125 ( .A1(npu_inst_n132), .A2(npu_inst_n128), .ZN(
        npu_inst_int_ckg[7]) );
  NAND2_X1 npu_inst_U124 ( .A1(npu_inst_n132), .A2(npu_inst_n130), .ZN(
        npu_inst_int_ckg[6]) );
  NAND2_X1 npu_inst_U123 ( .A1(npu_inst_n132), .A2(npu_inst_n136), .ZN(
        npu_inst_int_ckg[5]) );
  NAND2_X1 npu_inst_U122 ( .A1(npu_inst_n132), .A2(npu_inst_n134), .ZN(
        npu_inst_int_ckg[4]) );
  NAND2_X1 npu_inst_U121 ( .A1(npu_inst_n132), .A2(npu_inst_n138), .ZN(
        npu_inst_int_ckg[3]) );
  NAND2_X1 npu_inst_U120 ( .A1(npu_inst_n132), .A2(npu_inst_n139), .ZN(
        npu_inst_int_ckg[2]) );
  NAND2_X1 npu_inst_U119 ( .A1(npu_inst_n132), .A2(npu_inst_n140), .ZN(
        npu_inst_int_ckg[1]) );
  NAND2_X1 npu_inst_U118 ( .A1(npu_inst_n132), .A2(npu_inst_n131), .ZN(
        npu_inst_int_ckg[0]) );
  BUF_X1 npu_inst_U117 ( .A(ps_ctrl_wr_pipe), .Z(npu_inst_n6) );
  BUF_X1 npu_inst_U116 ( .A(ps_int_ifmaps_ptr[2]), .Z(npu_inst_n91) );
  BUF_X1 npu_inst_U115 ( .A(ps_int_ifmaps_ptr[2]), .Z(npu_inst_n89) );
  BUF_X1 npu_inst_U114 ( .A(ps_int_ifmaps_ptr[2]), .Z(npu_inst_n90) );
  BUF_X1 npu_inst_U113 ( .A(ps_int_ifmaps_ptr[1]), .Z(npu_inst_n74) );
  BUF_X1 npu_inst_U112 ( .A(ps_int_ifmaps_ptr[1]), .Z(npu_inst_n73) );
  BUF_X1 npu_inst_U111 ( .A(ps_int_ifmaps_ptr[0]), .Z(npu_inst_n71) );
  BUF_X1 npu_inst_U110 ( .A(ps_int_ifmaps_ptr[0]), .Z(npu_inst_n70) );
  BUF_X1 npu_inst_U109 ( .A(ps_int_ifmaps_ptr[0]), .Z(npu_inst_n69) );
  BUF_X1 npu_inst_U108 ( .A(ps_int_ifmaps_ptr[0]), .Z(npu_inst_n68) );
  BUF_X1 npu_inst_U107 ( .A(ps_int_ifmaps_ptr[0]), .Z(npu_inst_n67) );
  INV_X1 npu_inst_U106 ( .A(int_ckg_rmask[6]), .ZN(npu_inst_n142) );
  INV_X1 npu_inst_U105 ( .A(int_ckg_cmask[6]), .ZN(npu_inst_n140) );
  BUF_X1 npu_inst_U104 ( .A(n9), .Z(npu_inst_n121) );
  BUF_X1 npu_inst_U103 ( .A(n9), .Z(npu_inst_n120) );
  BUF_X1 npu_inst_U102 ( .A(npu_inst_n5), .Z(npu_inst_n4) );
  BUF_X1 npu_inst_U101 ( .A(npu_inst_n6), .Z(npu_inst_n2) );
  BUF_X1 npu_inst_U100 ( .A(npu_inst_n5), .Z(npu_inst_n3) );
  BUF_X2 npu_inst_U99 ( .A(npu_inst_n51), .Z(npu_inst_n60) );
  BUF_X2 npu_inst_U98 ( .A(npu_inst_n51), .Z(npu_inst_n59) );
  BUF_X2 npu_inst_U97 ( .A(npu_inst_n51), .Z(npu_inst_n58) );
  BUF_X2 npu_inst_U96 ( .A(npu_inst_n51), .Z(npu_inst_n57) );
  BUF_X2 npu_inst_U95 ( .A(npu_inst_n50), .Z(npu_inst_n56) );
  BUF_X2 npu_inst_U94 ( .A(npu_inst_n50), .Z(npu_inst_n55) );
  BUF_X2 npu_inst_U93 ( .A(npu_inst_n50), .Z(npu_inst_n54) );
  BUF_X2 npu_inst_U92 ( .A(npu_inst_n50), .Z(npu_inst_n53) );
  BUF_X2 npu_inst_U91 ( .A(npu_inst_n50), .Z(npu_inst_n52) );
  BUF_X1 npu_inst_U90 ( .A(npu_inst_n91), .Z(npu_inst_n82) );
  BUF_X1 npu_inst_U89 ( .A(npu_inst_n91), .Z(npu_inst_n81) );
  BUF_X1 npu_inst_U88 ( .A(npu_inst_n89), .Z(npu_inst_n88) );
  BUF_X1 npu_inst_U87 ( .A(npu_inst_n89), .Z(npu_inst_n87) );
  BUF_X1 npu_inst_U86 ( .A(npu_inst_n89), .Z(npu_inst_n86) );
  BUF_X1 npu_inst_U85 ( .A(npu_inst_n90), .Z(npu_inst_n85) );
  BUF_X1 npu_inst_U84 ( .A(npu_inst_n90), .Z(npu_inst_n84) );
  BUF_X1 npu_inst_U83 ( .A(npu_inst_n90), .Z(npu_inst_n83) );
  BUF_X1 npu_inst_U82 ( .A(npu_inst_n6), .Z(npu_inst_n1) );
  BUF_X1 npu_inst_U81 ( .A(npu_inst_n74), .Z(npu_inst_n80) );
  INV_X1 npu_inst_U80 ( .A(int_ckg_rmask[1]), .ZN(npu_inst_n133) );
  INV_X1 npu_inst_U79 ( .A(int_ckg_rmask[2]), .ZN(npu_inst_n137) );
  INV_X1 npu_inst_U78 ( .A(int_ckg_rmask[3]), .ZN(npu_inst_n135) );
  INV_X1 npu_inst_U77 ( .A(int_ckg_rmask[7]), .ZN(npu_inst_n132) );
  INV_X1 npu_inst_U76 ( .A(int_ckg_rmask[5]), .ZN(npu_inst_n141) );
  BUF_X1 npu_inst_U75 ( .A(npu_inst_n74), .Z(npu_inst_n79) );
  BUF_X1 npu_inst_U74 ( .A(npu_inst_n74), .Z(npu_inst_n78) );
  BUF_X1 npu_inst_U73 ( .A(npu_inst_n73), .Z(npu_inst_n77) );
  BUF_X1 npu_inst_U72 ( .A(npu_inst_n73), .Z(npu_inst_n76) );
  BUF_X1 npu_inst_U71 ( .A(npu_inst_n73), .Z(npu_inst_n75) );
  INV_X1 npu_inst_U70 ( .A(int_ckg_cmask[1]), .ZN(npu_inst_n130) );
  INV_X1 npu_inst_U69 ( .A(int_ckg_cmask[2]), .ZN(npu_inst_n136) );
  INV_X1 npu_inst_U68 ( .A(int_ckg_cmask[3]), .ZN(npu_inst_n134) );
  INV_X1 npu_inst_U67 ( .A(int_ckg_cmask[7]), .ZN(npu_inst_n131) );
  INV_X1 npu_inst_U66 ( .A(int_ckg_cmask[5]), .ZN(npu_inst_n139) );
  BUF_X1 npu_inst_U65 ( .A(npu_inst_n121), .Z(npu_inst_n127) );
  BUF_X1 npu_inst_U64 ( .A(npu_inst_n4), .Z(npu_inst_n49) );
  BUF_X1 npu_inst_U63 ( .A(npu_inst_n4), .Z(npu_inst_n48) );
  BUF_X1 npu_inst_U62 ( .A(npu_inst_n1), .Z(npu_inst_n41) );
  BUF_X1 npu_inst_U61 ( .A(npu_inst_n2), .Z(npu_inst_n42) );
  BUF_X1 npu_inst_U60 ( .A(npu_inst_n2), .Z(npu_inst_n43) );
  BUF_X1 npu_inst_U59 ( .A(npu_inst_n2), .Z(npu_inst_n44) );
  BUF_X1 npu_inst_U58 ( .A(npu_inst_n3), .Z(npu_inst_n45) );
  BUF_X1 npu_inst_U57 ( .A(npu_inst_n3), .Z(npu_inst_n46) );
  BUF_X1 npu_inst_U56 ( .A(npu_inst_n3), .Z(npu_inst_n47) );
  BUF_X1 npu_inst_U55 ( .A(npu_inst_n1), .Z(npu_inst_n39) );
  BUF_X1 npu_inst_U54 ( .A(npu_inst_n1), .Z(npu_inst_n40) );
  BUF_X1 npu_inst_U53 ( .A(npu_inst_n88), .Z(npu_inst_n107) );
  BUF_X1 npu_inst_U52 ( .A(npu_inst_n88), .Z(npu_inst_n106) );
  BUF_X1 npu_inst_U51 ( .A(npu_inst_n87), .Z(npu_inst_n105) );
  BUF_X1 npu_inst_U50 ( .A(npu_inst_n87), .Z(npu_inst_n104) );
  BUF_X1 npu_inst_U49 ( .A(npu_inst_n86), .Z(npu_inst_n103) );
  BUF_X1 npu_inst_U48 ( .A(npu_inst_n86), .Z(npu_inst_n102) );
  BUF_X1 npu_inst_U47 ( .A(npu_inst_n85), .Z(npu_inst_n101) );
  BUF_X1 npu_inst_U46 ( .A(npu_inst_n85), .Z(npu_inst_n100) );
  BUF_X1 npu_inst_U45 ( .A(npu_inst_n84), .Z(npu_inst_n99) );
  BUF_X1 npu_inst_U44 ( .A(npu_inst_n84), .Z(npu_inst_n98) );
  BUF_X1 npu_inst_U43 ( .A(npu_inst_n83), .Z(npu_inst_n97) );
  BUF_X1 npu_inst_U42 ( .A(npu_inst_n83), .Z(npu_inst_n96) );
  BUF_X1 npu_inst_U41 ( .A(npu_inst_n82), .Z(npu_inst_n95) );
  BUF_X1 npu_inst_U40 ( .A(npu_inst_n82), .Z(npu_inst_n94) );
  BUF_X1 npu_inst_U39 ( .A(npu_inst_n81), .Z(npu_inst_n93) );
  BUF_X1 npu_inst_U38 ( .A(npu_inst_n81), .Z(npu_inst_n92) );
  BUF_X1 npu_inst_U37 ( .A(npu_inst_n49), .Z(npu_inst_n8) );
  BUF_X1 npu_inst_U36 ( .A(npu_inst_n49), .Z(npu_inst_n7) );
  BUF_X1 npu_inst_U35 ( .A(npu_inst_n40), .Z(npu_inst_n34) );
  BUF_X1 npu_inst_U34 ( .A(npu_inst_n40), .Z(npu_inst_n33) );
  BUF_X1 npu_inst_U33 ( .A(npu_inst_n41), .Z(npu_inst_n32) );
  BUF_X1 npu_inst_U32 ( .A(npu_inst_n41), .Z(npu_inst_n31) );
  BUF_X1 npu_inst_U31 ( .A(npu_inst_n41), .Z(npu_inst_n30) );
  BUF_X1 npu_inst_U30 ( .A(npu_inst_n42), .Z(npu_inst_n29) );
  BUF_X1 npu_inst_U29 ( .A(npu_inst_n42), .Z(npu_inst_n28) );
  BUF_X1 npu_inst_U28 ( .A(npu_inst_n42), .Z(npu_inst_n27) );
  BUF_X1 npu_inst_U27 ( .A(npu_inst_n43), .Z(npu_inst_n26) );
  BUF_X1 npu_inst_U26 ( .A(npu_inst_n43), .Z(npu_inst_n25) );
  BUF_X1 npu_inst_U25 ( .A(npu_inst_n43), .Z(npu_inst_n24) );
  BUF_X1 npu_inst_U24 ( .A(npu_inst_n44), .Z(npu_inst_n23) );
  BUF_X1 npu_inst_U23 ( .A(npu_inst_n44), .Z(npu_inst_n22) );
  BUF_X1 npu_inst_U22 ( .A(npu_inst_n44), .Z(npu_inst_n21) );
  BUF_X1 npu_inst_U21 ( .A(npu_inst_n45), .Z(npu_inst_n20) );
  BUF_X1 npu_inst_U20 ( .A(npu_inst_n45), .Z(npu_inst_n19) );
  BUF_X1 npu_inst_U19 ( .A(npu_inst_n45), .Z(npu_inst_n18) );
  BUF_X1 npu_inst_U18 ( .A(npu_inst_n46), .Z(npu_inst_n17) );
  BUF_X1 npu_inst_U17 ( .A(npu_inst_n46), .Z(npu_inst_n16) );
  BUF_X1 npu_inst_U16 ( .A(npu_inst_n46), .Z(npu_inst_n15) );
  BUF_X1 npu_inst_U15 ( .A(npu_inst_n47), .Z(npu_inst_n14) );
  BUF_X1 npu_inst_U14 ( .A(npu_inst_n47), .Z(npu_inst_n13) );
  BUF_X1 npu_inst_U13 ( .A(npu_inst_n47), .Z(npu_inst_n12) );
  BUF_X1 npu_inst_U12 ( .A(npu_inst_n48), .Z(npu_inst_n11) );
  BUF_X1 npu_inst_U11 ( .A(npu_inst_n48), .Z(npu_inst_n10) );
  BUF_X1 npu_inst_U10 ( .A(npu_inst_n48), .Z(npu_inst_n9) );
  BUF_X1 npu_inst_U9 ( .A(npu_inst_n39), .Z(npu_inst_n38) );
  BUF_X1 npu_inst_U8 ( .A(npu_inst_n39), .Z(npu_inst_n37) );
  BUF_X1 npu_inst_U7 ( .A(npu_inst_n39), .Z(npu_inst_n36) );
  BUF_X1 npu_inst_U6 ( .A(npu_inst_n40), .Z(npu_inst_n35) );
  BUF_X1 npu_inst_U5 ( .A(npu_inst_n121), .Z(npu_inst_n126) );
  BUF_X1 npu_inst_U4 ( .A(npu_inst_n121), .Z(npu_inst_n125) );
  BUF_X1 npu_inst_U3 ( .A(npu_inst_n120), .Z(npu_inst_n124) );
  BUF_X1 npu_inst_U2 ( .A(npu_inst_n120), .Z(npu_inst_n123) );
  BUF_X1 npu_inst_U1 ( .A(npu_inst_n120), .Z(npu_inst_n122) );
  MUX2_X1 npu_inst_pe_1_0_0_U161 ( .A(npu_inst_pe_1_0_0_n31), .B(
        npu_inst_pe_1_0_0_n28), .S(npu_inst_pe_1_0_0_n7), .Z(
        npu_inst_pe_1_0_0_N93) );
  MUX2_X1 npu_inst_pe_1_0_0_U160 ( .A(npu_inst_pe_1_0_0_n30), .B(
        npu_inst_pe_1_0_0_n29), .S(npu_inst_n80), .Z(npu_inst_pe_1_0_0_n31) );
  MUX2_X1 npu_inst_pe_1_0_0_U159 ( .A(npu_inst_pe_1_0_0_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_0_0_int_q_reg_v_1__0_), .S(npu_inst_pe_1_0_0_n4), .Z(
        npu_inst_pe_1_0_0_n30) );
  MUX2_X1 npu_inst_pe_1_0_0_U158 ( .A(npu_inst_pe_1_0_0_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_0_0_int_q_reg_v_3__0_), .S(npu_inst_pe_1_0_0_n4), .Z(
        npu_inst_pe_1_0_0_n29) );
  MUX2_X1 npu_inst_pe_1_0_0_U157 ( .A(npu_inst_pe_1_0_0_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_0_0_int_q_reg_v_5__0_), .S(npu_inst_pe_1_0_0_n4), .Z(
        npu_inst_pe_1_0_0_n28) );
  MUX2_X1 npu_inst_pe_1_0_0_U156 ( .A(npu_inst_pe_1_0_0_n25), .B(
        npu_inst_pe_1_0_0_n22), .S(npu_inst_pe_1_0_0_n7), .Z(
        npu_inst_pe_1_0_0_N94) );
  MUX2_X1 npu_inst_pe_1_0_0_U155 ( .A(npu_inst_pe_1_0_0_n24), .B(
        npu_inst_pe_1_0_0_n23), .S(npu_inst_n80), .Z(npu_inst_pe_1_0_0_n25) );
  MUX2_X1 npu_inst_pe_1_0_0_U154 ( .A(npu_inst_pe_1_0_0_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_0_0_int_q_reg_v_1__1_), .S(npu_inst_pe_1_0_0_n4), .Z(
        npu_inst_pe_1_0_0_n24) );
  MUX2_X1 npu_inst_pe_1_0_0_U153 ( .A(npu_inst_pe_1_0_0_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_0_0_int_q_reg_v_3__1_), .S(npu_inst_pe_1_0_0_n4), .Z(
        npu_inst_pe_1_0_0_n23) );
  MUX2_X1 npu_inst_pe_1_0_0_U152 ( .A(npu_inst_pe_1_0_0_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_0_0_int_q_reg_v_5__1_), .S(npu_inst_pe_1_0_0_n4), .Z(
        npu_inst_pe_1_0_0_n22) );
  MUX2_X1 npu_inst_pe_1_0_0_U151 ( .A(npu_inst_pe_1_0_0_n21), .B(
        npu_inst_pe_1_0_0_n18), .S(npu_inst_pe_1_0_0_n7), .Z(
        npu_inst_pe_1_0_0_o_data_h_1_) );
  MUX2_X1 npu_inst_pe_1_0_0_U150 ( .A(npu_inst_pe_1_0_0_n20), .B(
        npu_inst_pe_1_0_0_n19), .S(npu_inst_n80), .Z(npu_inst_pe_1_0_0_n21) );
  MUX2_X1 npu_inst_pe_1_0_0_U149 ( .A(npu_inst_pe_1_0_0_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_0_0_int_q_reg_h_1__1_), .S(npu_inst_pe_1_0_0_n4), .Z(
        npu_inst_pe_1_0_0_n20) );
  MUX2_X1 npu_inst_pe_1_0_0_U148 ( .A(npu_inst_pe_1_0_0_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_0_0_int_q_reg_h_3__1_), .S(npu_inst_pe_1_0_0_n4), .Z(
        npu_inst_pe_1_0_0_n19) );
  MUX2_X1 npu_inst_pe_1_0_0_U147 ( .A(npu_inst_pe_1_0_0_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_0_0_int_q_reg_h_5__1_), .S(npu_inst_pe_1_0_0_n4), .Z(
        npu_inst_pe_1_0_0_n18) );
  MUX2_X1 npu_inst_pe_1_0_0_U146 ( .A(npu_inst_pe_1_0_0_n17), .B(
        npu_inst_pe_1_0_0_n14), .S(npu_inst_pe_1_0_0_n7), .Z(
        npu_inst_pe_1_0_0_o_data_h_0_) );
  MUX2_X1 npu_inst_pe_1_0_0_U145 ( .A(npu_inst_pe_1_0_0_n16), .B(
        npu_inst_pe_1_0_0_n15), .S(npu_inst_n80), .Z(npu_inst_pe_1_0_0_n17) );
  MUX2_X1 npu_inst_pe_1_0_0_U144 ( .A(npu_inst_pe_1_0_0_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_0_0_int_q_reg_h_1__0_), .S(npu_inst_pe_1_0_0_n4), .Z(
        npu_inst_pe_1_0_0_n16) );
  MUX2_X1 npu_inst_pe_1_0_0_U143 ( .A(npu_inst_pe_1_0_0_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_0_0_int_q_reg_h_3__0_), .S(npu_inst_pe_1_0_0_n4), .Z(
        npu_inst_pe_1_0_0_n15) );
  MUX2_X1 npu_inst_pe_1_0_0_U142 ( .A(npu_inst_pe_1_0_0_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_0_0_int_q_reg_h_5__0_), .S(npu_inst_pe_1_0_0_n4), .Z(
        npu_inst_pe_1_0_0_n14) );
  XOR2_X1 npu_inst_pe_1_0_0_U141 ( .A(npu_inst_pe_1_0_0_int_data_0_), .B(
        npu_inst_pe_1_0_0_int_q_acc_0_), .Z(npu_inst_pe_1_0_0_N73) );
  AND2_X1 npu_inst_pe_1_0_0_U140 ( .A1(npu_inst_pe_1_0_0_int_q_acc_0_), .A2(
        npu_inst_pe_1_0_0_int_data_0_), .ZN(npu_inst_pe_1_0_0_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_0_0_U139 ( .A(npu_inst_pe_1_0_0_int_q_acc_0_), .B(
        npu_inst_pe_1_0_0_n12), .ZN(npu_inst_pe_1_0_0_N65) );
  OR2_X1 npu_inst_pe_1_0_0_U138 ( .A1(npu_inst_pe_1_0_0_n12), .A2(
        npu_inst_pe_1_0_0_int_q_acc_0_), .ZN(npu_inst_pe_1_0_0_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_0_0_U137 ( .A(npu_inst_pe_1_0_0_int_q_acc_2_), .B(
        npu_inst_pe_1_0_0_add_79_carry_2_), .Z(npu_inst_pe_1_0_0_N75) );
  AND2_X1 npu_inst_pe_1_0_0_U136 ( .A1(npu_inst_pe_1_0_0_add_79_carry_2_), 
        .A2(npu_inst_pe_1_0_0_int_q_acc_2_), .ZN(
        npu_inst_pe_1_0_0_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_0_0_U135 ( .A(npu_inst_pe_1_0_0_int_q_acc_3_), .B(
        npu_inst_pe_1_0_0_add_79_carry_3_), .Z(npu_inst_pe_1_0_0_N76) );
  AND2_X1 npu_inst_pe_1_0_0_U134 ( .A1(npu_inst_pe_1_0_0_add_79_carry_3_), 
        .A2(npu_inst_pe_1_0_0_int_q_acc_3_), .ZN(
        npu_inst_pe_1_0_0_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_0_0_U133 ( .A(npu_inst_pe_1_0_0_int_q_acc_4_), .B(
        npu_inst_pe_1_0_0_add_79_carry_4_), .Z(npu_inst_pe_1_0_0_N77) );
  AND2_X1 npu_inst_pe_1_0_0_U132 ( .A1(npu_inst_pe_1_0_0_add_79_carry_4_), 
        .A2(npu_inst_pe_1_0_0_int_q_acc_4_), .ZN(
        npu_inst_pe_1_0_0_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_0_0_U131 ( .A(npu_inst_pe_1_0_0_int_q_acc_5_), .B(
        npu_inst_pe_1_0_0_add_79_carry_5_), .Z(npu_inst_pe_1_0_0_N78) );
  AND2_X1 npu_inst_pe_1_0_0_U130 ( .A1(npu_inst_pe_1_0_0_add_79_carry_5_), 
        .A2(npu_inst_pe_1_0_0_int_q_acc_5_), .ZN(
        npu_inst_pe_1_0_0_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_0_0_U129 ( .A(npu_inst_pe_1_0_0_int_q_acc_6_), .B(
        npu_inst_pe_1_0_0_add_79_carry_6_), .Z(npu_inst_pe_1_0_0_N79) );
  AND2_X1 npu_inst_pe_1_0_0_U128 ( .A1(npu_inst_pe_1_0_0_add_79_carry_6_), 
        .A2(npu_inst_pe_1_0_0_int_q_acc_6_), .ZN(
        npu_inst_pe_1_0_0_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_0_0_U127 ( .A(npu_inst_pe_1_0_0_int_q_acc_7_), .B(
        npu_inst_pe_1_0_0_add_79_carry_7_), .Z(npu_inst_pe_1_0_0_N80) );
  XNOR2_X1 npu_inst_pe_1_0_0_U126 ( .A(npu_inst_pe_1_0_0_sub_77_carry_2_), .B(
        npu_inst_pe_1_0_0_int_q_acc_2_), .ZN(npu_inst_pe_1_0_0_N67) );
  OR2_X1 npu_inst_pe_1_0_0_U125 ( .A1(npu_inst_pe_1_0_0_int_q_acc_2_), .A2(
        npu_inst_pe_1_0_0_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_0_0_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_0_0_U124 ( .A(npu_inst_pe_1_0_0_sub_77_carry_3_), .B(
        npu_inst_pe_1_0_0_int_q_acc_3_), .ZN(npu_inst_pe_1_0_0_N68) );
  OR2_X1 npu_inst_pe_1_0_0_U123 ( .A1(npu_inst_pe_1_0_0_int_q_acc_3_), .A2(
        npu_inst_pe_1_0_0_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_0_0_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_0_0_U122 ( .A(npu_inst_pe_1_0_0_sub_77_carry_4_), .B(
        npu_inst_pe_1_0_0_int_q_acc_4_), .ZN(npu_inst_pe_1_0_0_N69) );
  OR2_X1 npu_inst_pe_1_0_0_U121 ( .A1(npu_inst_pe_1_0_0_int_q_acc_4_), .A2(
        npu_inst_pe_1_0_0_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_0_0_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_0_0_U120 ( .A(npu_inst_pe_1_0_0_sub_77_carry_5_), .B(
        npu_inst_pe_1_0_0_int_q_acc_5_), .ZN(npu_inst_pe_1_0_0_N70) );
  OR2_X1 npu_inst_pe_1_0_0_U119 ( .A1(npu_inst_pe_1_0_0_int_q_acc_5_), .A2(
        npu_inst_pe_1_0_0_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_0_0_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_0_0_U118 ( .A(npu_inst_pe_1_0_0_sub_77_carry_6_), .B(
        npu_inst_pe_1_0_0_int_q_acc_6_), .ZN(npu_inst_pe_1_0_0_N71) );
  OR2_X1 npu_inst_pe_1_0_0_U117 ( .A1(npu_inst_pe_1_0_0_int_q_acc_6_), .A2(
        npu_inst_pe_1_0_0_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_0_0_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_0_0_U116 ( .A(npu_inst_pe_1_0_0_int_q_acc_7_), .B(
        npu_inst_pe_1_0_0_sub_77_carry_7_), .ZN(npu_inst_pe_1_0_0_N72) );
  INV_X1 npu_inst_pe_1_0_0_U115 ( .A(npu_inst_n80), .ZN(npu_inst_pe_1_0_0_n6)
         );
  INV_X1 npu_inst_pe_1_0_0_U114 ( .A(npu_inst_n57), .ZN(npu_inst_pe_1_0_0_n3)
         );
  AOI22_X1 npu_inst_pe_1_0_0_U113 ( .A1(npu_inst_int_data_y_1__0__0_), .A2(
        npu_inst_pe_1_0_0_n58), .B1(npu_inst_pe_1_0_0_n113), .B2(
        npu_inst_pe_1_0_0_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_0_0_n57) );
  INV_X1 npu_inst_pe_1_0_0_U112 ( .A(npu_inst_pe_1_0_0_n57), .ZN(
        npu_inst_pe_1_0_0_n107) );
  AOI22_X1 npu_inst_pe_1_0_0_U111 ( .A1(npu_inst_int_data_y_1__0__0_), .A2(
        npu_inst_pe_1_0_0_n54), .B1(npu_inst_pe_1_0_0_n114), .B2(
        npu_inst_pe_1_0_0_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_0_0_n53) );
  INV_X1 npu_inst_pe_1_0_0_U110 ( .A(npu_inst_pe_1_0_0_n53), .ZN(
        npu_inst_pe_1_0_0_n108) );
  AOI22_X1 npu_inst_pe_1_0_0_U107 ( .A1(npu_inst_int_data_y_1__0__0_), .A2(
        npu_inst_pe_1_0_0_n50), .B1(npu_inst_pe_1_0_0_n115), .B2(
        npu_inst_pe_1_0_0_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_0_0_n49) );
  INV_X1 npu_inst_pe_1_0_0_U106 ( .A(npu_inst_pe_1_0_0_n49), .ZN(
        npu_inst_pe_1_0_0_n109) );
  AOI22_X1 npu_inst_pe_1_0_0_U105 ( .A1(npu_inst_int_data_y_1__0__0_), .A2(
        npu_inst_pe_1_0_0_n46), .B1(npu_inst_pe_1_0_0_n116), .B2(
        npu_inst_pe_1_0_0_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_0_0_n45) );
  INV_X1 npu_inst_pe_1_0_0_U104 ( .A(npu_inst_pe_1_0_0_n45), .ZN(
        npu_inst_pe_1_0_0_n110) );
  AOI22_X1 npu_inst_pe_1_0_0_U103 ( .A1(npu_inst_int_data_y_1__0__0_), .A2(
        npu_inst_pe_1_0_0_n42), .B1(npu_inst_pe_1_0_0_n118), .B2(
        npu_inst_pe_1_0_0_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_0_0_n41) );
  INV_X1 npu_inst_pe_1_0_0_U102 ( .A(npu_inst_pe_1_0_0_n41), .ZN(
        npu_inst_pe_1_0_0_n111) );
  AOI22_X1 npu_inst_pe_1_0_0_U101 ( .A1(npu_inst_int_data_y_1__0__1_), .A2(
        npu_inst_pe_1_0_0_n58), .B1(npu_inst_pe_1_0_0_n113), .B2(
        npu_inst_pe_1_0_0_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_0_0_n59) );
  INV_X1 npu_inst_pe_1_0_0_U100 ( .A(npu_inst_pe_1_0_0_n59), .ZN(
        npu_inst_pe_1_0_0_n101) );
  AOI22_X1 npu_inst_pe_1_0_0_U99 ( .A1(npu_inst_int_data_y_1__0__1_), .A2(
        npu_inst_pe_1_0_0_n54), .B1(npu_inst_pe_1_0_0_n114), .B2(
        npu_inst_pe_1_0_0_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_0_0_n55) );
  INV_X1 npu_inst_pe_1_0_0_U98 ( .A(npu_inst_pe_1_0_0_n55), .ZN(
        npu_inst_pe_1_0_0_n102) );
  AOI22_X1 npu_inst_pe_1_0_0_U97 ( .A1(npu_inst_int_data_y_1__0__1_), .A2(
        npu_inst_pe_1_0_0_n50), .B1(npu_inst_pe_1_0_0_n115), .B2(
        npu_inst_pe_1_0_0_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_0_0_n51) );
  INV_X1 npu_inst_pe_1_0_0_U96 ( .A(npu_inst_pe_1_0_0_n51), .ZN(
        npu_inst_pe_1_0_0_n103) );
  AOI22_X1 npu_inst_pe_1_0_0_U95 ( .A1(npu_inst_int_data_y_1__0__1_), .A2(
        npu_inst_pe_1_0_0_n46), .B1(npu_inst_pe_1_0_0_n116), .B2(
        npu_inst_pe_1_0_0_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_0_0_n47) );
  INV_X1 npu_inst_pe_1_0_0_U94 ( .A(npu_inst_pe_1_0_0_n47), .ZN(
        npu_inst_pe_1_0_0_n104) );
  AOI22_X1 npu_inst_pe_1_0_0_U93 ( .A1(npu_inst_int_data_y_1__0__1_), .A2(
        npu_inst_pe_1_0_0_n42), .B1(npu_inst_pe_1_0_0_n118), .B2(
        npu_inst_pe_1_0_0_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_0_0_n43) );
  INV_X1 npu_inst_pe_1_0_0_U92 ( .A(npu_inst_pe_1_0_0_n43), .ZN(
        npu_inst_pe_1_0_0_n105) );
  AOI22_X1 npu_inst_pe_1_0_0_U91 ( .A1(npu_inst_pe_1_0_0_n38), .A2(
        npu_inst_int_data_y_1__0__1_), .B1(npu_inst_pe_1_0_0_n117), .B2(
        npu_inst_pe_1_0_0_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_0_0_n39) );
  INV_X1 npu_inst_pe_1_0_0_U90 ( .A(npu_inst_pe_1_0_0_n39), .ZN(
        npu_inst_pe_1_0_0_n106) );
  AOI22_X1 npu_inst_pe_1_0_0_U89 ( .A1(npu_inst_pe_1_0_0_n38), .A2(
        npu_inst_int_data_y_1__0__0_), .B1(npu_inst_pe_1_0_0_n117), .B2(
        npu_inst_pe_1_0_0_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_0_0_n37) );
  INV_X1 npu_inst_pe_1_0_0_U88 ( .A(npu_inst_pe_1_0_0_n37), .ZN(
        npu_inst_pe_1_0_0_n112) );
  NOR3_X1 npu_inst_pe_1_0_0_U87 ( .A1(npu_inst_pe_1_0_0_n26), .A2(npu_inst_n57), .A3(npu_inst_int_ckg[63]), .ZN(npu_inst_pe_1_0_0_n85) );
  OR2_X1 npu_inst_pe_1_0_0_U86 ( .A1(npu_inst_pe_1_0_0_n85), .A2(
        npu_inst_pe_1_0_0_n2), .ZN(npu_inst_pe_1_0_0_N84) );
  AND2_X1 npu_inst_pe_1_0_0_U85 ( .A1(npu_inst_pe_1_0_0_n2), .A2(
        npu_inst_pe_1_0_0_int_q_acc_7_), .ZN(o_data[63]) );
  AND2_X1 npu_inst_pe_1_0_0_U84 ( .A1(npu_inst_pe_1_0_0_int_q_acc_6_), .A2(
        npu_inst_pe_1_0_0_n2), .ZN(o_data[62]) );
  AND2_X1 npu_inst_pe_1_0_0_U83 ( .A1(npu_inst_pe_1_0_0_int_q_acc_5_), .A2(
        npu_inst_pe_1_0_0_n2), .ZN(o_data[61]) );
  AND2_X1 npu_inst_pe_1_0_0_U82 ( .A1(npu_inst_pe_1_0_0_int_q_acc_4_), .A2(
        npu_inst_pe_1_0_0_n2), .ZN(o_data[60]) );
  AND2_X1 npu_inst_pe_1_0_0_U81 ( .A1(npu_inst_pe_1_0_0_int_q_acc_3_), .A2(
        npu_inst_pe_1_0_0_n2), .ZN(o_data[59]) );
  NAND2_X1 npu_inst_pe_1_0_0_U80 ( .A1(npu_inst_pe_1_0_0_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_0_0_n60), .ZN(npu_inst_pe_1_0_0_n74) );
  OAI21_X1 npu_inst_pe_1_0_0_U79 ( .B1(npu_inst_pe_1_0_0_n63), .B2(
        npu_inst_pe_1_0_0_n60), .A(npu_inst_pe_1_0_0_n74), .ZN(
        npu_inst_pe_1_0_0_n97) );
  NAND2_X1 npu_inst_pe_1_0_0_U78 ( .A1(npu_inst_pe_1_0_0_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_0_0_n60), .ZN(npu_inst_pe_1_0_0_n73) );
  OAI21_X1 npu_inst_pe_1_0_0_U77 ( .B1(npu_inst_pe_1_0_0_n61), .B2(
        npu_inst_pe_1_0_0_n60), .A(npu_inst_pe_1_0_0_n73), .ZN(
        npu_inst_pe_1_0_0_n96) );
  NAND2_X1 npu_inst_pe_1_0_0_U76 ( .A1(npu_inst_pe_1_0_0_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_0_0_n56), .ZN(npu_inst_pe_1_0_0_n72) );
  OAI21_X1 npu_inst_pe_1_0_0_U75 ( .B1(npu_inst_pe_1_0_0_n63), .B2(
        npu_inst_pe_1_0_0_n56), .A(npu_inst_pe_1_0_0_n72), .ZN(
        npu_inst_pe_1_0_0_n95) );
  NAND2_X1 npu_inst_pe_1_0_0_U74 ( .A1(npu_inst_pe_1_0_0_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_0_0_n56), .ZN(npu_inst_pe_1_0_0_n71) );
  OAI21_X1 npu_inst_pe_1_0_0_U73 ( .B1(npu_inst_pe_1_0_0_n61), .B2(
        npu_inst_pe_1_0_0_n56), .A(npu_inst_pe_1_0_0_n71), .ZN(
        npu_inst_pe_1_0_0_n94) );
  NAND2_X1 npu_inst_pe_1_0_0_U72 ( .A1(npu_inst_pe_1_0_0_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_0_0_n52), .ZN(npu_inst_pe_1_0_0_n70) );
  OAI21_X1 npu_inst_pe_1_0_0_U71 ( .B1(npu_inst_pe_1_0_0_n63), .B2(
        npu_inst_pe_1_0_0_n52), .A(npu_inst_pe_1_0_0_n70), .ZN(
        npu_inst_pe_1_0_0_n93) );
  NAND2_X1 npu_inst_pe_1_0_0_U70 ( .A1(npu_inst_pe_1_0_0_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_0_0_n52), .ZN(npu_inst_pe_1_0_0_n69) );
  OAI21_X1 npu_inst_pe_1_0_0_U69 ( .B1(npu_inst_pe_1_0_0_n61), .B2(
        npu_inst_pe_1_0_0_n52), .A(npu_inst_pe_1_0_0_n69), .ZN(
        npu_inst_pe_1_0_0_n92) );
  NAND2_X1 npu_inst_pe_1_0_0_U68 ( .A1(npu_inst_pe_1_0_0_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_0_0_n48), .ZN(npu_inst_pe_1_0_0_n68) );
  OAI21_X1 npu_inst_pe_1_0_0_U67 ( .B1(npu_inst_pe_1_0_0_n63), .B2(
        npu_inst_pe_1_0_0_n48), .A(npu_inst_pe_1_0_0_n68), .ZN(
        npu_inst_pe_1_0_0_n91) );
  NAND2_X1 npu_inst_pe_1_0_0_U66 ( .A1(npu_inst_pe_1_0_0_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_0_0_n48), .ZN(npu_inst_pe_1_0_0_n67) );
  OAI21_X1 npu_inst_pe_1_0_0_U65 ( .B1(npu_inst_pe_1_0_0_n61), .B2(
        npu_inst_pe_1_0_0_n48), .A(npu_inst_pe_1_0_0_n67), .ZN(
        npu_inst_pe_1_0_0_n90) );
  NAND2_X1 npu_inst_pe_1_0_0_U64 ( .A1(npu_inst_pe_1_0_0_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_0_0_n44), .ZN(npu_inst_pe_1_0_0_n66) );
  OAI21_X1 npu_inst_pe_1_0_0_U63 ( .B1(npu_inst_pe_1_0_0_n63), .B2(
        npu_inst_pe_1_0_0_n44), .A(npu_inst_pe_1_0_0_n66), .ZN(
        npu_inst_pe_1_0_0_n89) );
  NAND2_X1 npu_inst_pe_1_0_0_U62 ( .A1(npu_inst_pe_1_0_0_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_0_0_n44), .ZN(npu_inst_pe_1_0_0_n65) );
  OAI21_X1 npu_inst_pe_1_0_0_U61 ( .B1(npu_inst_pe_1_0_0_n61), .B2(
        npu_inst_pe_1_0_0_n44), .A(npu_inst_pe_1_0_0_n65), .ZN(
        npu_inst_pe_1_0_0_n88) );
  NAND2_X1 npu_inst_pe_1_0_0_U60 ( .A1(npu_inst_pe_1_0_0_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_0_0_n40), .ZN(npu_inst_pe_1_0_0_n64) );
  OAI21_X1 npu_inst_pe_1_0_0_U59 ( .B1(npu_inst_pe_1_0_0_n63), .B2(
        npu_inst_pe_1_0_0_n40), .A(npu_inst_pe_1_0_0_n64), .ZN(
        npu_inst_pe_1_0_0_n87) );
  NAND2_X1 npu_inst_pe_1_0_0_U58 ( .A1(npu_inst_pe_1_0_0_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_0_0_n40), .ZN(npu_inst_pe_1_0_0_n62) );
  OAI21_X1 npu_inst_pe_1_0_0_U57 ( .B1(npu_inst_pe_1_0_0_n61), .B2(
        npu_inst_pe_1_0_0_n40), .A(npu_inst_pe_1_0_0_n62), .ZN(
        npu_inst_pe_1_0_0_n86) );
  AND2_X1 npu_inst_pe_1_0_0_U56 ( .A1(npu_inst_pe_1_0_0_int_q_acc_0_), .A2(
        npu_inst_pe_1_0_0_n1), .ZN(o_data[56]) );
  AND2_X1 npu_inst_pe_1_0_0_U55 ( .A1(npu_inst_pe_1_0_0_int_q_acc_1_), .A2(
        npu_inst_pe_1_0_0_n1), .ZN(o_data[57]) );
  AND2_X1 npu_inst_pe_1_0_0_U54 ( .A1(npu_inst_pe_1_0_0_int_q_acc_2_), .A2(
        npu_inst_pe_1_0_0_n1), .ZN(o_data[58]) );
  AOI222_X1 npu_inst_pe_1_0_0_U53 ( .A1(npu_inst_int_data_res_1__0__0_), .A2(
        npu_inst_pe_1_0_0_n1), .B1(npu_inst_pe_1_0_0_N73), .B2(
        npu_inst_pe_1_0_0_n76), .C1(npu_inst_pe_1_0_0_N65), .C2(
        npu_inst_pe_1_0_0_n77), .ZN(npu_inst_pe_1_0_0_n84) );
  INV_X1 npu_inst_pe_1_0_0_U52 ( .A(npu_inst_pe_1_0_0_n84), .ZN(
        npu_inst_pe_1_0_0_n100) );
  AOI222_X1 npu_inst_pe_1_0_0_U51 ( .A1(npu_inst_int_data_res_1__0__7_), .A2(
        npu_inst_pe_1_0_0_n1), .B1(npu_inst_pe_1_0_0_N80), .B2(
        npu_inst_pe_1_0_0_n76), .C1(npu_inst_pe_1_0_0_N72), .C2(
        npu_inst_pe_1_0_0_n77), .ZN(npu_inst_pe_1_0_0_n75) );
  INV_X1 npu_inst_pe_1_0_0_U50 ( .A(npu_inst_pe_1_0_0_n75), .ZN(
        npu_inst_pe_1_0_0_n32) );
  AOI222_X1 npu_inst_pe_1_0_0_U49 ( .A1(npu_inst_int_data_res_1__0__1_), .A2(
        npu_inst_pe_1_0_0_n1), .B1(npu_inst_pe_1_0_0_N74), .B2(
        npu_inst_pe_1_0_0_n76), .C1(npu_inst_pe_1_0_0_N66), .C2(
        npu_inst_pe_1_0_0_n77), .ZN(npu_inst_pe_1_0_0_n83) );
  INV_X1 npu_inst_pe_1_0_0_U48 ( .A(npu_inst_pe_1_0_0_n83), .ZN(
        npu_inst_pe_1_0_0_n99) );
  AOI222_X1 npu_inst_pe_1_0_0_U47 ( .A1(npu_inst_int_data_res_1__0__2_), .A2(
        npu_inst_pe_1_0_0_n1), .B1(npu_inst_pe_1_0_0_N75), .B2(
        npu_inst_pe_1_0_0_n76), .C1(npu_inst_pe_1_0_0_N67), .C2(
        npu_inst_pe_1_0_0_n77), .ZN(npu_inst_pe_1_0_0_n82) );
  INV_X1 npu_inst_pe_1_0_0_U46 ( .A(npu_inst_pe_1_0_0_n82), .ZN(
        npu_inst_pe_1_0_0_n98) );
  AOI222_X1 npu_inst_pe_1_0_0_U45 ( .A1(npu_inst_int_data_res_1__0__3_), .A2(
        npu_inst_pe_1_0_0_n1), .B1(npu_inst_pe_1_0_0_N76), .B2(
        npu_inst_pe_1_0_0_n76), .C1(npu_inst_pe_1_0_0_N68), .C2(
        npu_inst_pe_1_0_0_n77), .ZN(npu_inst_pe_1_0_0_n81) );
  INV_X1 npu_inst_pe_1_0_0_U44 ( .A(npu_inst_pe_1_0_0_n81), .ZN(
        npu_inst_pe_1_0_0_n36) );
  AOI222_X1 npu_inst_pe_1_0_0_U43 ( .A1(npu_inst_int_data_res_1__0__4_), .A2(
        npu_inst_pe_1_0_0_n1), .B1(npu_inst_pe_1_0_0_N77), .B2(
        npu_inst_pe_1_0_0_n76), .C1(npu_inst_pe_1_0_0_N69), .C2(
        npu_inst_pe_1_0_0_n77), .ZN(npu_inst_pe_1_0_0_n80) );
  INV_X1 npu_inst_pe_1_0_0_U42 ( .A(npu_inst_pe_1_0_0_n80), .ZN(
        npu_inst_pe_1_0_0_n35) );
  AOI222_X1 npu_inst_pe_1_0_0_U41 ( .A1(npu_inst_int_data_res_1__0__5_), .A2(
        npu_inst_pe_1_0_0_n1), .B1(npu_inst_pe_1_0_0_N78), .B2(
        npu_inst_pe_1_0_0_n76), .C1(npu_inst_pe_1_0_0_N70), .C2(
        npu_inst_pe_1_0_0_n77), .ZN(npu_inst_pe_1_0_0_n79) );
  INV_X1 npu_inst_pe_1_0_0_U40 ( .A(npu_inst_pe_1_0_0_n79), .ZN(
        npu_inst_pe_1_0_0_n34) );
  AOI222_X1 npu_inst_pe_1_0_0_U39 ( .A1(npu_inst_int_data_res_1__0__6_), .A2(
        npu_inst_pe_1_0_0_n1), .B1(npu_inst_pe_1_0_0_N79), .B2(
        npu_inst_pe_1_0_0_n76), .C1(npu_inst_pe_1_0_0_N71), .C2(
        npu_inst_pe_1_0_0_n77), .ZN(npu_inst_pe_1_0_0_n78) );
  INV_X1 npu_inst_pe_1_0_0_U38 ( .A(npu_inst_pe_1_0_0_n78), .ZN(
        npu_inst_pe_1_0_0_n33) );
  AND2_X1 npu_inst_pe_1_0_0_U37 ( .A1(npu_inst_pe_1_0_0_o_data_h_1_), .A2(
        npu_inst_pe_1_0_0_int_q_weight_1_), .ZN(npu_inst_pe_1_0_0_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_0_0_U36 ( .A1(npu_inst_pe_1_0_0_o_data_h_0_), .A2(
        npu_inst_pe_1_0_0_int_q_weight_1_), .ZN(npu_inst_pe_1_0_0_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_0_0_U35 ( .A(npu_inst_pe_1_0_0_int_data_1_), .ZN(
        npu_inst_pe_1_0_0_n13) );
  AND2_X1 npu_inst_pe_1_0_0_U34 ( .A1(npu_inst_pe_1_0_0_N93), .A2(npu_inst_n57), .ZN(npu_inst_pe_1_0_0_o_data_v_0_) );
  AND2_X1 npu_inst_pe_1_0_0_U33 ( .A1(npu_inst_n57), .A2(npu_inst_pe_1_0_0_N94), .ZN(npu_inst_pe_1_0_0_o_data_v_1_) );
  AOI22_X1 npu_inst_pe_1_0_0_U32 ( .A1(npu_inst_n57), .A2(
        npu_inst_int_data_y_1__0__1_), .B1(npu_inst_pe_1_0_0_n3), .B2(
        npu_inst_int_data_x_0__1__1_), .ZN(npu_inst_pe_1_0_0_n63) );
  AOI22_X1 npu_inst_pe_1_0_0_U31 ( .A1(npu_inst_n57), .A2(
        npu_inst_int_data_y_1__0__0_), .B1(npu_inst_pe_1_0_0_n3), .B2(
        npu_inst_int_data_x_0__1__0_), .ZN(npu_inst_pe_1_0_0_n61) );
  INV_X1 npu_inst_pe_1_0_0_U30 ( .A(npu_inst_pe_1_0_0_int_data_0_), .ZN(
        npu_inst_pe_1_0_0_n12) );
  INV_X1 npu_inst_pe_1_0_0_U29 ( .A(npu_inst_n72), .ZN(npu_inst_pe_1_0_0_n5)
         );
  OR3_X1 npu_inst_pe_1_0_0_U28 ( .A1(npu_inst_n80), .A2(npu_inst_pe_1_0_0_n7), 
        .A3(npu_inst_pe_1_0_0_n5), .ZN(npu_inst_pe_1_0_0_n56) );
  OR3_X1 npu_inst_pe_1_0_0_U27 ( .A1(npu_inst_pe_1_0_0_n5), .A2(
        npu_inst_pe_1_0_0_n7), .A3(npu_inst_pe_1_0_0_n6), .ZN(
        npu_inst_pe_1_0_0_n48) );
  INV_X1 npu_inst_pe_1_0_0_U26 ( .A(npu_inst_pe_1_0_0_n5), .ZN(
        npu_inst_pe_1_0_0_n4) );
  INV_X1 npu_inst_pe_1_0_0_U25 ( .A(npu_inst_n127), .ZN(npu_inst_pe_1_0_0_n11)
         );
  OR3_X1 npu_inst_pe_1_0_0_U24 ( .A1(npu_inst_pe_1_0_0_n4), .A2(
        npu_inst_pe_1_0_0_n7), .A3(npu_inst_pe_1_0_0_n6), .ZN(
        npu_inst_pe_1_0_0_n52) );
  OR3_X1 npu_inst_pe_1_0_0_U23 ( .A1(npu_inst_n80), .A2(npu_inst_pe_1_0_0_n7), 
        .A3(npu_inst_pe_1_0_0_n4), .ZN(npu_inst_pe_1_0_0_n60) );
  NOR2_X1 npu_inst_pe_1_0_0_U22 ( .A1(npu_inst_pe_1_0_0_n60), .A2(
        npu_inst_pe_1_0_0_n3), .ZN(npu_inst_pe_1_0_0_n58) );
  NOR2_X1 npu_inst_pe_1_0_0_U21 ( .A1(npu_inst_pe_1_0_0_n56), .A2(
        npu_inst_pe_1_0_0_n3), .ZN(npu_inst_pe_1_0_0_n54) );
  NOR2_X1 npu_inst_pe_1_0_0_U20 ( .A1(npu_inst_pe_1_0_0_n52), .A2(
        npu_inst_pe_1_0_0_n3), .ZN(npu_inst_pe_1_0_0_n50) );
  NOR2_X1 npu_inst_pe_1_0_0_U19 ( .A1(npu_inst_pe_1_0_0_n48), .A2(
        npu_inst_pe_1_0_0_n3), .ZN(npu_inst_pe_1_0_0_n46) );
  NOR2_X1 npu_inst_pe_1_0_0_U18 ( .A1(npu_inst_pe_1_0_0_n40), .A2(
        npu_inst_pe_1_0_0_n3), .ZN(npu_inst_pe_1_0_0_n38) );
  NOR2_X1 npu_inst_pe_1_0_0_U17 ( .A1(npu_inst_pe_1_0_0_n44), .A2(
        npu_inst_pe_1_0_0_n3), .ZN(npu_inst_pe_1_0_0_n42) );
  BUF_X1 npu_inst_pe_1_0_0_U16 ( .A(npu_inst_n107), .Z(npu_inst_pe_1_0_0_n7)
         );
  BUF_X1 npu_inst_pe_1_0_0_U15 ( .A(npu_inst_pe_1_0_0_n11), .Z(
        npu_inst_pe_1_0_0_n10) );
  BUF_X1 npu_inst_pe_1_0_0_U14 ( .A(npu_inst_pe_1_0_0_n11), .Z(
        npu_inst_pe_1_0_0_n9) );
  BUF_X1 npu_inst_pe_1_0_0_U13 ( .A(npu_inst_pe_1_0_0_n11), .Z(
        npu_inst_pe_1_0_0_n8) );
  INV_X1 npu_inst_pe_1_0_0_U12 ( .A(npu_inst_pe_1_0_0_n38), .ZN(
        npu_inst_pe_1_0_0_n117) );
  INV_X1 npu_inst_pe_1_0_0_U11 ( .A(npu_inst_pe_1_0_0_n58), .ZN(
        npu_inst_pe_1_0_0_n113) );
  INV_X1 npu_inst_pe_1_0_0_U10 ( .A(npu_inst_pe_1_0_0_n54), .ZN(
        npu_inst_pe_1_0_0_n114) );
  INV_X1 npu_inst_pe_1_0_0_U9 ( .A(npu_inst_pe_1_0_0_n50), .ZN(
        npu_inst_pe_1_0_0_n115) );
  INV_X1 npu_inst_pe_1_0_0_U8 ( .A(npu_inst_pe_1_0_0_n46), .ZN(
        npu_inst_pe_1_0_0_n116) );
  INV_X1 npu_inst_pe_1_0_0_U7 ( .A(npu_inst_pe_1_0_0_n42), .ZN(
        npu_inst_pe_1_0_0_n118) );
  BUF_X1 npu_inst_pe_1_0_0_U6 ( .A(npu_inst_n38), .Z(npu_inst_pe_1_0_0_n2) );
  BUF_X1 npu_inst_pe_1_0_0_U5 ( .A(npu_inst_n38), .Z(npu_inst_pe_1_0_0_n1) );
  NOR2_X1 npu_inst_pe_1_0_0_U4 ( .A1(npu_inst_pe_1_0_0_int_q_weight_0_), .A2(
        npu_inst_pe_1_0_0_n1), .ZN(npu_inst_pe_1_0_0_n76) );
  NOR2_X1 npu_inst_pe_1_0_0_U3 ( .A1(npu_inst_pe_1_0_0_n27), .A2(
        npu_inst_pe_1_0_0_n1), .ZN(npu_inst_pe_1_0_0_n77) );
  FA_X1 npu_inst_pe_1_0_0_sub_77_U2_1 ( .A(npu_inst_pe_1_0_0_int_q_acc_1_), 
        .B(npu_inst_pe_1_0_0_n13), .CI(npu_inst_pe_1_0_0_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_0_0_sub_77_carry_2_), .S(npu_inst_pe_1_0_0_N66) );
  FA_X1 npu_inst_pe_1_0_0_add_79_U1_1 ( .A(npu_inst_pe_1_0_0_int_q_acc_1_), 
        .B(npu_inst_pe_1_0_0_int_data_1_), .CI(
        npu_inst_pe_1_0_0_add_79_carry_1_), .CO(
        npu_inst_pe_1_0_0_add_79_carry_2_), .S(npu_inst_pe_1_0_0_N74) );
  NAND3_X1 npu_inst_pe_1_0_0_U109 ( .A1(npu_inst_pe_1_0_0_n5), .A2(
        npu_inst_pe_1_0_0_n6), .A3(npu_inst_pe_1_0_0_n7), .ZN(
        npu_inst_pe_1_0_0_n44) );
  NAND3_X1 npu_inst_pe_1_0_0_U108 ( .A1(npu_inst_pe_1_0_0_n4), .A2(
        npu_inst_pe_1_0_0_n6), .A3(npu_inst_pe_1_0_0_n7), .ZN(
        npu_inst_pe_1_0_0_n40) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_0_0_n33), .CK(
        npu_inst_pe_1_0_0_net4293), .RN(npu_inst_pe_1_0_0_n8), .Q(
        npu_inst_pe_1_0_0_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_0_0_n34), .CK(
        npu_inst_pe_1_0_0_net4293), .RN(npu_inst_pe_1_0_0_n8), .Q(
        npu_inst_pe_1_0_0_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_0_0_n35), .CK(
        npu_inst_pe_1_0_0_net4293), .RN(npu_inst_pe_1_0_0_n8), .Q(
        npu_inst_pe_1_0_0_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_0_0_n36), .CK(
        npu_inst_pe_1_0_0_net4293), .RN(npu_inst_pe_1_0_0_n8), .Q(
        npu_inst_pe_1_0_0_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_0_0_n98), .CK(
        npu_inst_pe_1_0_0_net4293), .RN(npu_inst_pe_1_0_0_n8), .Q(
        npu_inst_pe_1_0_0_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_0_0_n99), .CK(
        npu_inst_pe_1_0_0_net4293), .RN(npu_inst_pe_1_0_0_n8), .Q(
        npu_inst_pe_1_0_0_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_0_0_n32), .CK(
        npu_inst_pe_1_0_0_net4293), .RN(npu_inst_pe_1_0_0_n8), .Q(
        npu_inst_pe_1_0_0_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_0_0_n100), 
        .CK(npu_inst_pe_1_0_0_net4293), .RN(npu_inst_pe_1_0_0_n8), .Q(
        npu_inst_pe_1_0_0_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_weight_reg_0_ ( .D(npu_inst_n113), .CK(
        npu_inst_pe_1_0_0_net4299), .RN(npu_inst_pe_1_0_0_n8), .Q(
        npu_inst_pe_1_0_0_int_q_weight_0_), .QN(npu_inst_pe_1_0_0_n27) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_weight_reg_1_ ( .D(npu_inst_n119), .CK(
        npu_inst_pe_1_0_0_net4299), .RN(npu_inst_pe_1_0_0_n8), .Q(
        npu_inst_pe_1_0_0_int_q_weight_1_), .QN(npu_inst_pe_1_0_0_n26) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_0_0_n112), 
        .CK(npu_inst_pe_1_0_0_net4299), .RN(npu_inst_pe_1_0_0_n8), .Q(
        npu_inst_pe_1_0_0_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_0_0_n106), 
        .CK(npu_inst_pe_1_0_0_net4299), .RN(npu_inst_pe_1_0_0_n8), .Q(
        npu_inst_pe_1_0_0_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_0_0_n111), 
        .CK(npu_inst_pe_1_0_0_net4299), .RN(npu_inst_pe_1_0_0_n9), .Q(
        npu_inst_pe_1_0_0_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_0_0_n105), 
        .CK(npu_inst_pe_1_0_0_net4299), .RN(npu_inst_pe_1_0_0_n9), .Q(
        npu_inst_pe_1_0_0_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_0_0_n110), 
        .CK(npu_inst_pe_1_0_0_net4299), .RN(npu_inst_pe_1_0_0_n9), .Q(
        npu_inst_pe_1_0_0_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_0_0_n104), 
        .CK(npu_inst_pe_1_0_0_net4299), .RN(npu_inst_pe_1_0_0_n9), .Q(
        npu_inst_pe_1_0_0_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_0_0_n109), 
        .CK(npu_inst_pe_1_0_0_net4299), .RN(npu_inst_pe_1_0_0_n9), .Q(
        npu_inst_pe_1_0_0_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_0_0_n103), 
        .CK(npu_inst_pe_1_0_0_net4299), .RN(npu_inst_pe_1_0_0_n9), .Q(
        npu_inst_pe_1_0_0_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_0_0_n108), 
        .CK(npu_inst_pe_1_0_0_net4299), .RN(npu_inst_pe_1_0_0_n9), .Q(
        npu_inst_pe_1_0_0_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_0_0_n102), 
        .CK(npu_inst_pe_1_0_0_net4299), .RN(npu_inst_pe_1_0_0_n9), .Q(
        npu_inst_pe_1_0_0_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_0_0_n107), 
        .CK(npu_inst_pe_1_0_0_net4299), .RN(npu_inst_pe_1_0_0_n9), .Q(
        npu_inst_pe_1_0_0_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_0_0_n101), 
        .CK(npu_inst_pe_1_0_0_net4299), .RN(npu_inst_pe_1_0_0_n9), .Q(
        npu_inst_pe_1_0_0_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_0_0_n86), 
        .CK(npu_inst_pe_1_0_0_net4299), .RN(npu_inst_pe_1_0_0_n9), .Q(
        npu_inst_pe_1_0_0_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_0_0_n87), 
        .CK(npu_inst_pe_1_0_0_net4299), .RN(npu_inst_pe_1_0_0_n9), .Q(
        npu_inst_pe_1_0_0_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_0_0_n88), 
        .CK(npu_inst_pe_1_0_0_net4299), .RN(npu_inst_pe_1_0_0_n10), .Q(
        npu_inst_pe_1_0_0_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_0_0_n89), 
        .CK(npu_inst_pe_1_0_0_net4299), .RN(npu_inst_pe_1_0_0_n10), .Q(
        npu_inst_pe_1_0_0_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_0_0_n90), 
        .CK(npu_inst_pe_1_0_0_net4299), .RN(npu_inst_pe_1_0_0_n10), .Q(
        npu_inst_pe_1_0_0_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_0_0_n91), 
        .CK(npu_inst_pe_1_0_0_net4299), .RN(npu_inst_pe_1_0_0_n10), .Q(
        npu_inst_pe_1_0_0_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_0_0_n92), 
        .CK(npu_inst_pe_1_0_0_net4299), .RN(npu_inst_pe_1_0_0_n10), .Q(
        npu_inst_pe_1_0_0_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_0_0_n93), 
        .CK(npu_inst_pe_1_0_0_net4299), .RN(npu_inst_pe_1_0_0_n10), .Q(
        npu_inst_pe_1_0_0_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_0_0_n94), 
        .CK(npu_inst_pe_1_0_0_net4299), .RN(npu_inst_pe_1_0_0_n10), .Q(
        npu_inst_pe_1_0_0_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_0_0_n95), 
        .CK(npu_inst_pe_1_0_0_net4299), .RN(npu_inst_pe_1_0_0_n10), .Q(
        npu_inst_pe_1_0_0_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_0_0_n96), 
        .CK(npu_inst_pe_1_0_0_net4299), .RN(npu_inst_pe_1_0_0_n10), .Q(
        npu_inst_pe_1_0_0_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_0_0_n97), 
        .CK(npu_inst_pe_1_0_0_net4299), .RN(npu_inst_pe_1_0_0_n10), .Q(
        npu_inst_pe_1_0_0_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_0_0_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_0_0_N84), .SE(1'b0), .GCK(npu_inst_pe_1_0_0_net4293) );
  CLKGATETST_X1 npu_inst_pe_1_0_0_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n66), .SE(1'b0), .GCK(npu_inst_pe_1_0_0_net4299) );
  MUX2_X1 npu_inst_pe_1_0_1_U160 ( .A(npu_inst_pe_1_0_1_n30), .B(
        npu_inst_pe_1_0_1_n25), .S(npu_inst_pe_1_0_1_n6), .Z(
        npu_inst_pe_1_0_1_N93) );
  MUX2_X1 npu_inst_pe_1_0_1_U159 ( .A(npu_inst_pe_1_0_1_n29), .B(
        npu_inst_pe_1_0_1_n28), .S(npu_inst_n80), .Z(npu_inst_pe_1_0_1_n30) );
  MUX2_X1 npu_inst_pe_1_0_1_U158 ( .A(npu_inst_pe_1_0_1_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_0_1_int_q_reg_v_1__0_), .S(npu_inst_n72), .Z(
        npu_inst_pe_1_0_1_n29) );
  MUX2_X1 npu_inst_pe_1_0_1_U157 ( .A(npu_inst_pe_1_0_1_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_0_1_int_q_reg_v_3__0_), .S(npu_inst_n72), .Z(
        npu_inst_pe_1_0_1_n28) );
  MUX2_X1 npu_inst_pe_1_0_1_U156 ( .A(npu_inst_pe_1_0_1_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_0_1_int_q_reg_v_5__0_), .S(npu_inst_n72), .Z(
        npu_inst_pe_1_0_1_n25) );
  MUX2_X1 npu_inst_pe_1_0_1_U155 ( .A(npu_inst_pe_1_0_1_n24), .B(
        npu_inst_pe_1_0_1_n21), .S(npu_inst_pe_1_0_1_n6), .Z(
        npu_inst_pe_1_0_1_N94) );
  MUX2_X1 npu_inst_pe_1_0_1_U154 ( .A(npu_inst_pe_1_0_1_n23), .B(
        npu_inst_pe_1_0_1_n22), .S(npu_inst_n80), .Z(npu_inst_pe_1_0_1_n24) );
  MUX2_X1 npu_inst_pe_1_0_1_U153 ( .A(npu_inst_pe_1_0_1_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_0_1_int_q_reg_v_1__1_), .S(npu_inst_n72), .Z(
        npu_inst_pe_1_0_1_n23) );
  MUX2_X1 npu_inst_pe_1_0_1_U152 ( .A(npu_inst_pe_1_0_1_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_0_1_int_q_reg_v_3__1_), .S(npu_inst_n72), .Z(
        npu_inst_pe_1_0_1_n22) );
  MUX2_X1 npu_inst_pe_1_0_1_U151 ( .A(npu_inst_pe_1_0_1_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_0_1_int_q_reg_v_5__1_), .S(npu_inst_n72), .Z(
        npu_inst_pe_1_0_1_n21) );
  MUX2_X1 npu_inst_pe_1_0_1_U150 ( .A(npu_inst_pe_1_0_1_n20), .B(
        npu_inst_pe_1_0_1_n17), .S(npu_inst_pe_1_0_1_n6), .Z(
        npu_inst_int_data_x_0__1__1_) );
  MUX2_X1 npu_inst_pe_1_0_1_U149 ( .A(npu_inst_pe_1_0_1_n19), .B(
        npu_inst_pe_1_0_1_n18), .S(npu_inst_n80), .Z(npu_inst_pe_1_0_1_n20) );
  MUX2_X1 npu_inst_pe_1_0_1_U148 ( .A(npu_inst_pe_1_0_1_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_0_1_int_q_reg_h_1__1_), .S(npu_inst_n72), .Z(
        npu_inst_pe_1_0_1_n19) );
  MUX2_X1 npu_inst_pe_1_0_1_U147 ( .A(npu_inst_pe_1_0_1_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_0_1_int_q_reg_h_3__1_), .S(npu_inst_n72), .Z(
        npu_inst_pe_1_0_1_n18) );
  MUX2_X1 npu_inst_pe_1_0_1_U146 ( .A(npu_inst_pe_1_0_1_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_0_1_int_q_reg_h_5__1_), .S(npu_inst_n72), .Z(
        npu_inst_pe_1_0_1_n17) );
  MUX2_X1 npu_inst_pe_1_0_1_U145 ( .A(npu_inst_pe_1_0_1_n16), .B(
        npu_inst_pe_1_0_1_n13), .S(npu_inst_pe_1_0_1_n6), .Z(
        npu_inst_int_data_x_0__1__0_) );
  MUX2_X1 npu_inst_pe_1_0_1_U144 ( .A(npu_inst_pe_1_0_1_n15), .B(
        npu_inst_pe_1_0_1_n14), .S(npu_inst_n80), .Z(npu_inst_pe_1_0_1_n16) );
  MUX2_X1 npu_inst_pe_1_0_1_U143 ( .A(npu_inst_pe_1_0_1_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_0_1_int_q_reg_h_1__0_), .S(npu_inst_n72), .Z(
        npu_inst_pe_1_0_1_n15) );
  MUX2_X1 npu_inst_pe_1_0_1_U142 ( .A(npu_inst_pe_1_0_1_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_0_1_int_q_reg_h_3__0_), .S(npu_inst_n72), .Z(
        npu_inst_pe_1_0_1_n14) );
  MUX2_X1 npu_inst_pe_1_0_1_U141 ( .A(npu_inst_pe_1_0_1_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_0_1_int_q_reg_h_5__0_), .S(npu_inst_n72), .Z(
        npu_inst_pe_1_0_1_n13) );
  XOR2_X1 npu_inst_pe_1_0_1_U140 ( .A(npu_inst_pe_1_0_1_int_data_0_), .B(
        npu_inst_pe_1_0_1_int_q_acc_0_), .Z(npu_inst_pe_1_0_1_N73) );
  AND2_X1 npu_inst_pe_1_0_1_U139 ( .A1(npu_inst_pe_1_0_1_int_q_acc_0_), .A2(
        npu_inst_pe_1_0_1_int_data_0_), .ZN(npu_inst_pe_1_0_1_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_0_1_U138 ( .A(npu_inst_pe_1_0_1_int_q_acc_0_), .B(
        npu_inst_pe_1_0_1_n11), .ZN(npu_inst_pe_1_0_1_N65) );
  OR2_X1 npu_inst_pe_1_0_1_U137 ( .A1(npu_inst_pe_1_0_1_n11), .A2(
        npu_inst_pe_1_0_1_int_q_acc_0_), .ZN(npu_inst_pe_1_0_1_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_0_1_U136 ( .A(npu_inst_pe_1_0_1_int_q_acc_2_), .B(
        npu_inst_pe_1_0_1_add_79_carry_2_), .Z(npu_inst_pe_1_0_1_N75) );
  AND2_X1 npu_inst_pe_1_0_1_U135 ( .A1(npu_inst_pe_1_0_1_add_79_carry_2_), 
        .A2(npu_inst_pe_1_0_1_int_q_acc_2_), .ZN(
        npu_inst_pe_1_0_1_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_0_1_U134 ( .A(npu_inst_pe_1_0_1_int_q_acc_3_), .B(
        npu_inst_pe_1_0_1_add_79_carry_3_), .Z(npu_inst_pe_1_0_1_N76) );
  AND2_X1 npu_inst_pe_1_0_1_U133 ( .A1(npu_inst_pe_1_0_1_add_79_carry_3_), 
        .A2(npu_inst_pe_1_0_1_int_q_acc_3_), .ZN(
        npu_inst_pe_1_0_1_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_0_1_U132 ( .A(npu_inst_pe_1_0_1_int_q_acc_4_), .B(
        npu_inst_pe_1_0_1_add_79_carry_4_), .Z(npu_inst_pe_1_0_1_N77) );
  AND2_X1 npu_inst_pe_1_0_1_U131 ( .A1(npu_inst_pe_1_0_1_add_79_carry_4_), 
        .A2(npu_inst_pe_1_0_1_int_q_acc_4_), .ZN(
        npu_inst_pe_1_0_1_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_0_1_U130 ( .A(npu_inst_pe_1_0_1_int_q_acc_5_), .B(
        npu_inst_pe_1_0_1_add_79_carry_5_), .Z(npu_inst_pe_1_0_1_N78) );
  AND2_X1 npu_inst_pe_1_0_1_U129 ( .A1(npu_inst_pe_1_0_1_add_79_carry_5_), 
        .A2(npu_inst_pe_1_0_1_int_q_acc_5_), .ZN(
        npu_inst_pe_1_0_1_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_0_1_U128 ( .A(npu_inst_pe_1_0_1_int_q_acc_6_), .B(
        npu_inst_pe_1_0_1_add_79_carry_6_), .Z(npu_inst_pe_1_0_1_N79) );
  AND2_X1 npu_inst_pe_1_0_1_U127 ( .A1(npu_inst_pe_1_0_1_add_79_carry_6_), 
        .A2(npu_inst_pe_1_0_1_int_q_acc_6_), .ZN(
        npu_inst_pe_1_0_1_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_0_1_U126 ( .A(npu_inst_pe_1_0_1_int_q_acc_7_), .B(
        npu_inst_pe_1_0_1_add_79_carry_7_), .Z(npu_inst_pe_1_0_1_N80) );
  XNOR2_X1 npu_inst_pe_1_0_1_U125 ( .A(npu_inst_pe_1_0_1_sub_77_carry_2_), .B(
        npu_inst_pe_1_0_1_int_q_acc_2_), .ZN(npu_inst_pe_1_0_1_N67) );
  OR2_X1 npu_inst_pe_1_0_1_U124 ( .A1(npu_inst_pe_1_0_1_int_q_acc_2_), .A2(
        npu_inst_pe_1_0_1_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_0_1_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_0_1_U123 ( .A(npu_inst_pe_1_0_1_sub_77_carry_3_), .B(
        npu_inst_pe_1_0_1_int_q_acc_3_), .ZN(npu_inst_pe_1_0_1_N68) );
  OR2_X1 npu_inst_pe_1_0_1_U122 ( .A1(npu_inst_pe_1_0_1_int_q_acc_3_), .A2(
        npu_inst_pe_1_0_1_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_0_1_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_0_1_U121 ( .A(npu_inst_pe_1_0_1_sub_77_carry_4_), .B(
        npu_inst_pe_1_0_1_int_q_acc_4_), .ZN(npu_inst_pe_1_0_1_N69) );
  OR2_X1 npu_inst_pe_1_0_1_U120 ( .A1(npu_inst_pe_1_0_1_int_q_acc_4_), .A2(
        npu_inst_pe_1_0_1_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_0_1_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_0_1_U119 ( .A(npu_inst_pe_1_0_1_sub_77_carry_5_), .B(
        npu_inst_pe_1_0_1_int_q_acc_5_), .ZN(npu_inst_pe_1_0_1_N70) );
  OR2_X1 npu_inst_pe_1_0_1_U118 ( .A1(npu_inst_pe_1_0_1_int_q_acc_5_), .A2(
        npu_inst_pe_1_0_1_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_0_1_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_0_1_U117 ( .A(npu_inst_pe_1_0_1_sub_77_carry_6_), .B(
        npu_inst_pe_1_0_1_int_q_acc_6_), .ZN(npu_inst_pe_1_0_1_N71) );
  OR2_X1 npu_inst_pe_1_0_1_U116 ( .A1(npu_inst_pe_1_0_1_int_q_acc_6_), .A2(
        npu_inst_pe_1_0_1_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_0_1_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_0_1_U115 ( .A(npu_inst_pe_1_0_1_int_q_acc_7_), .B(
        npu_inst_pe_1_0_1_sub_77_carry_7_), .ZN(npu_inst_pe_1_0_1_N72) );
  INV_X1 npu_inst_pe_1_0_1_U114 ( .A(npu_inst_n80), .ZN(npu_inst_pe_1_0_1_n5)
         );
  INV_X1 npu_inst_pe_1_0_1_U113 ( .A(npu_inst_n60), .ZN(npu_inst_pe_1_0_1_n3)
         );
  AOI22_X1 npu_inst_pe_1_0_1_U112 ( .A1(npu_inst_int_data_y_1__1__0_), .A2(
        npu_inst_pe_1_0_1_n58), .B1(npu_inst_pe_1_0_1_n112), .B2(
        npu_inst_pe_1_0_1_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_0_1_n57) );
  INV_X1 npu_inst_pe_1_0_1_U111 ( .A(npu_inst_pe_1_0_1_n57), .ZN(
        npu_inst_pe_1_0_1_n106) );
  AOI22_X1 npu_inst_pe_1_0_1_U110 ( .A1(npu_inst_int_data_y_1__1__0_), .A2(
        npu_inst_pe_1_0_1_n54), .B1(npu_inst_pe_1_0_1_n113), .B2(
        npu_inst_pe_1_0_1_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_0_1_n53) );
  INV_X1 npu_inst_pe_1_0_1_U107 ( .A(npu_inst_pe_1_0_1_n53), .ZN(
        npu_inst_pe_1_0_1_n107) );
  AOI22_X1 npu_inst_pe_1_0_1_U106 ( .A1(npu_inst_int_data_y_1__1__0_), .A2(
        npu_inst_pe_1_0_1_n50), .B1(npu_inst_pe_1_0_1_n114), .B2(
        npu_inst_pe_1_0_1_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_0_1_n49) );
  INV_X1 npu_inst_pe_1_0_1_U105 ( .A(npu_inst_pe_1_0_1_n49), .ZN(
        npu_inst_pe_1_0_1_n108) );
  AOI22_X1 npu_inst_pe_1_0_1_U104 ( .A1(npu_inst_int_data_y_1__1__0_), .A2(
        npu_inst_pe_1_0_1_n46), .B1(npu_inst_pe_1_0_1_n115), .B2(
        npu_inst_pe_1_0_1_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_0_1_n45) );
  INV_X1 npu_inst_pe_1_0_1_U103 ( .A(npu_inst_pe_1_0_1_n45), .ZN(
        npu_inst_pe_1_0_1_n109) );
  AOI22_X1 npu_inst_pe_1_0_1_U102 ( .A1(npu_inst_int_data_y_1__1__0_), .A2(
        npu_inst_pe_1_0_1_n42), .B1(npu_inst_pe_1_0_1_n117), .B2(
        npu_inst_pe_1_0_1_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_0_1_n41) );
  INV_X1 npu_inst_pe_1_0_1_U101 ( .A(npu_inst_pe_1_0_1_n41), .ZN(
        npu_inst_pe_1_0_1_n110) );
  AOI22_X1 npu_inst_pe_1_0_1_U100 ( .A1(npu_inst_int_data_y_1__1__1_), .A2(
        npu_inst_pe_1_0_1_n58), .B1(npu_inst_pe_1_0_1_n112), .B2(
        npu_inst_pe_1_0_1_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_0_1_n59) );
  INV_X1 npu_inst_pe_1_0_1_U99 ( .A(npu_inst_pe_1_0_1_n59), .ZN(
        npu_inst_pe_1_0_1_n100) );
  AOI22_X1 npu_inst_pe_1_0_1_U98 ( .A1(npu_inst_int_data_y_1__1__1_), .A2(
        npu_inst_pe_1_0_1_n54), .B1(npu_inst_pe_1_0_1_n113), .B2(
        npu_inst_pe_1_0_1_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_0_1_n55) );
  INV_X1 npu_inst_pe_1_0_1_U97 ( .A(npu_inst_pe_1_0_1_n55), .ZN(
        npu_inst_pe_1_0_1_n101) );
  AOI22_X1 npu_inst_pe_1_0_1_U96 ( .A1(npu_inst_int_data_y_1__1__1_), .A2(
        npu_inst_pe_1_0_1_n50), .B1(npu_inst_pe_1_0_1_n114), .B2(
        npu_inst_pe_1_0_1_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_0_1_n51) );
  INV_X1 npu_inst_pe_1_0_1_U95 ( .A(npu_inst_pe_1_0_1_n51), .ZN(
        npu_inst_pe_1_0_1_n102) );
  AOI22_X1 npu_inst_pe_1_0_1_U94 ( .A1(npu_inst_int_data_y_1__1__1_), .A2(
        npu_inst_pe_1_0_1_n46), .B1(npu_inst_pe_1_0_1_n115), .B2(
        npu_inst_pe_1_0_1_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_0_1_n47) );
  INV_X1 npu_inst_pe_1_0_1_U93 ( .A(npu_inst_pe_1_0_1_n47), .ZN(
        npu_inst_pe_1_0_1_n103) );
  AOI22_X1 npu_inst_pe_1_0_1_U92 ( .A1(npu_inst_int_data_y_1__1__1_), .A2(
        npu_inst_pe_1_0_1_n42), .B1(npu_inst_pe_1_0_1_n117), .B2(
        npu_inst_pe_1_0_1_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_0_1_n43) );
  INV_X1 npu_inst_pe_1_0_1_U91 ( .A(npu_inst_pe_1_0_1_n43), .ZN(
        npu_inst_pe_1_0_1_n104) );
  AOI22_X1 npu_inst_pe_1_0_1_U90 ( .A1(npu_inst_pe_1_0_1_n38), .A2(
        npu_inst_int_data_y_1__1__1_), .B1(npu_inst_pe_1_0_1_n116), .B2(
        npu_inst_pe_1_0_1_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_0_1_n39) );
  INV_X1 npu_inst_pe_1_0_1_U89 ( .A(npu_inst_pe_1_0_1_n39), .ZN(
        npu_inst_pe_1_0_1_n105) );
  AOI22_X1 npu_inst_pe_1_0_1_U88 ( .A1(npu_inst_pe_1_0_1_n38), .A2(
        npu_inst_int_data_y_1__1__0_), .B1(npu_inst_pe_1_0_1_n116), .B2(
        npu_inst_pe_1_0_1_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_0_1_n37) );
  INV_X1 npu_inst_pe_1_0_1_U87 ( .A(npu_inst_pe_1_0_1_n37), .ZN(
        npu_inst_pe_1_0_1_n111) );
  AND2_X1 npu_inst_pe_1_0_1_U86 ( .A1(npu_inst_pe_1_0_1_n2), .A2(
        npu_inst_pe_1_0_1_int_q_acc_7_), .ZN(o_data[55]) );
  AND2_X1 npu_inst_pe_1_0_1_U85 ( .A1(npu_inst_pe_1_0_1_int_q_acc_6_), .A2(
        npu_inst_pe_1_0_1_n2), .ZN(o_data[54]) );
  AND2_X1 npu_inst_pe_1_0_1_U84 ( .A1(npu_inst_pe_1_0_1_int_q_acc_5_), .A2(
        npu_inst_pe_1_0_1_n2), .ZN(o_data[53]) );
  AND2_X1 npu_inst_pe_1_0_1_U83 ( .A1(npu_inst_pe_1_0_1_int_q_acc_4_), .A2(
        npu_inst_pe_1_0_1_n2), .ZN(o_data[52]) );
  AND2_X1 npu_inst_pe_1_0_1_U82 ( .A1(npu_inst_pe_1_0_1_int_q_acc_3_), .A2(
        npu_inst_pe_1_0_1_n2), .ZN(o_data[51]) );
  NAND2_X1 npu_inst_pe_1_0_1_U81 ( .A1(npu_inst_pe_1_0_1_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_0_1_n60), .ZN(npu_inst_pe_1_0_1_n74) );
  OAI21_X1 npu_inst_pe_1_0_1_U80 ( .B1(npu_inst_pe_1_0_1_n63), .B2(
        npu_inst_pe_1_0_1_n60), .A(npu_inst_pe_1_0_1_n74), .ZN(
        npu_inst_pe_1_0_1_n97) );
  NAND2_X1 npu_inst_pe_1_0_1_U79 ( .A1(npu_inst_pe_1_0_1_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_0_1_n60), .ZN(npu_inst_pe_1_0_1_n73) );
  OAI21_X1 npu_inst_pe_1_0_1_U78 ( .B1(npu_inst_pe_1_0_1_n61), .B2(
        npu_inst_pe_1_0_1_n60), .A(npu_inst_pe_1_0_1_n73), .ZN(
        npu_inst_pe_1_0_1_n96) );
  NAND2_X1 npu_inst_pe_1_0_1_U77 ( .A1(npu_inst_pe_1_0_1_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_0_1_n56), .ZN(npu_inst_pe_1_0_1_n72) );
  OAI21_X1 npu_inst_pe_1_0_1_U76 ( .B1(npu_inst_pe_1_0_1_n63), .B2(
        npu_inst_pe_1_0_1_n56), .A(npu_inst_pe_1_0_1_n72), .ZN(
        npu_inst_pe_1_0_1_n95) );
  NAND2_X1 npu_inst_pe_1_0_1_U75 ( .A1(npu_inst_pe_1_0_1_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_0_1_n56), .ZN(npu_inst_pe_1_0_1_n71) );
  OAI21_X1 npu_inst_pe_1_0_1_U74 ( .B1(npu_inst_pe_1_0_1_n61), .B2(
        npu_inst_pe_1_0_1_n56), .A(npu_inst_pe_1_0_1_n71), .ZN(
        npu_inst_pe_1_0_1_n94) );
  NAND2_X1 npu_inst_pe_1_0_1_U73 ( .A1(npu_inst_pe_1_0_1_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_0_1_n52), .ZN(npu_inst_pe_1_0_1_n70) );
  OAI21_X1 npu_inst_pe_1_0_1_U72 ( .B1(npu_inst_pe_1_0_1_n63), .B2(
        npu_inst_pe_1_0_1_n52), .A(npu_inst_pe_1_0_1_n70), .ZN(
        npu_inst_pe_1_0_1_n93) );
  NAND2_X1 npu_inst_pe_1_0_1_U71 ( .A1(npu_inst_pe_1_0_1_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_0_1_n52), .ZN(npu_inst_pe_1_0_1_n69) );
  OAI21_X1 npu_inst_pe_1_0_1_U70 ( .B1(npu_inst_pe_1_0_1_n61), .B2(
        npu_inst_pe_1_0_1_n52), .A(npu_inst_pe_1_0_1_n69), .ZN(
        npu_inst_pe_1_0_1_n92) );
  NAND2_X1 npu_inst_pe_1_0_1_U69 ( .A1(npu_inst_pe_1_0_1_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_0_1_n48), .ZN(npu_inst_pe_1_0_1_n68) );
  OAI21_X1 npu_inst_pe_1_0_1_U68 ( .B1(npu_inst_pe_1_0_1_n63), .B2(
        npu_inst_pe_1_0_1_n48), .A(npu_inst_pe_1_0_1_n68), .ZN(
        npu_inst_pe_1_0_1_n91) );
  NAND2_X1 npu_inst_pe_1_0_1_U67 ( .A1(npu_inst_pe_1_0_1_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_0_1_n48), .ZN(npu_inst_pe_1_0_1_n67) );
  OAI21_X1 npu_inst_pe_1_0_1_U66 ( .B1(npu_inst_pe_1_0_1_n61), .B2(
        npu_inst_pe_1_0_1_n48), .A(npu_inst_pe_1_0_1_n67), .ZN(
        npu_inst_pe_1_0_1_n90) );
  NAND2_X1 npu_inst_pe_1_0_1_U65 ( .A1(npu_inst_pe_1_0_1_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_0_1_n44), .ZN(npu_inst_pe_1_0_1_n66) );
  OAI21_X1 npu_inst_pe_1_0_1_U64 ( .B1(npu_inst_pe_1_0_1_n63), .B2(
        npu_inst_pe_1_0_1_n44), .A(npu_inst_pe_1_0_1_n66), .ZN(
        npu_inst_pe_1_0_1_n89) );
  NAND2_X1 npu_inst_pe_1_0_1_U63 ( .A1(npu_inst_pe_1_0_1_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_0_1_n44), .ZN(npu_inst_pe_1_0_1_n65) );
  OAI21_X1 npu_inst_pe_1_0_1_U62 ( .B1(npu_inst_pe_1_0_1_n61), .B2(
        npu_inst_pe_1_0_1_n44), .A(npu_inst_pe_1_0_1_n65), .ZN(
        npu_inst_pe_1_0_1_n88) );
  NAND2_X1 npu_inst_pe_1_0_1_U61 ( .A1(npu_inst_pe_1_0_1_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_0_1_n40), .ZN(npu_inst_pe_1_0_1_n64) );
  OAI21_X1 npu_inst_pe_1_0_1_U60 ( .B1(npu_inst_pe_1_0_1_n63), .B2(
        npu_inst_pe_1_0_1_n40), .A(npu_inst_pe_1_0_1_n64), .ZN(
        npu_inst_pe_1_0_1_n87) );
  NAND2_X1 npu_inst_pe_1_0_1_U59 ( .A1(npu_inst_pe_1_0_1_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_0_1_n40), .ZN(npu_inst_pe_1_0_1_n62) );
  OAI21_X1 npu_inst_pe_1_0_1_U58 ( .B1(npu_inst_pe_1_0_1_n61), .B2(
        npu_inst_pe_1_0_1_n40), .A(npu_inst_pe_1_0_1_n62), .ZN(
        npu_inst_pe_1_0_1_n86) );
  NOR3_X1 npu_inst_pe_1_0_1_U57 ( .A1(npu_inst_pe_1_0_1_n26), .A2(npu_inst_n60), .A3(npu_inst_int_ckg[62]), .ZN(npu_inst_pe_1_0_1_n85) );
  OR2_X1 npu_inst_pe_1_0_1_U56 ( .A1(npu_inst_pe_1_0_1_n85), .A2(
        npu_inst_pe_1_0_1_n2), .ZN(npu_inst_pe_1_0_1_N84) );
  AND2_X1 npu_inst_pe_1_0_1_U55 ( .A1(npu_inst_pe_1_0_1_int_q_acc_0_), .A2(
        npu_inst_pe_1_0_1_n1), .ZN(o_data[48]) );
  AND2_X1 npu_inst_pe_1_0_1_U54 ( .A1(npu_inst_pe_1_0_1_int_q_acc_1_), .A2(
        npu_inst_pe_1_0_1_n1), .ZN(o_data[49]) );
  AND2_X1 npu_inst_pe_1_0_1_U53 ( .A1(npu_inst_pe_1_0_1_int_q_acc_2_), .A2(
        npu_inst_pe_1_0_1_n1), .ZN(o_data[50]) );
  AOI222_X1 npu_inst_pe_1_0_1_U52 ( .A1(npu_inst_int_data_res_1__1__0_), .A2(
        npu_inst_pe_1_0_1_n1), .B1(npu_inst_pe_1_0_1_N73), .B2(
        npu_inst_pe_1_0_1_n76), .C1(npu_inst_pe_1_0_1_N65), .C2(
        npu_inst_pe_1_0_1_n77), .ZN(npu_inst_pe_1_0_1_n84) );
  INV_X1 npu_inst_pe_1_0_1_U51 ( .A(npu_inst_pe_1_0_1_n84), .ZN(
        npu_inst_pe_1_0_1_n99) );
  AOI222_X1 npu_inst_pe_1_0_1_U50 ( .A1(npu_inst_int_data_res_1__1__7_), .A2(
        npu_inst_pe_1_0_1_n1), .B1(npu_inst_pe_1_0_1_N80), .B2(
        npu_inst_pe_1_0_1_n76), .C1(npu_inst_pe_1_0_1_N72), .C2(
        npu_inst_pe_1_0_1_n77), .ZN(npu_inst_pe_1_0_1_n75) );
  INV_X1 npu_inst_pe_1_0_1_U49 ( .A(npu_inst_pe_1_0_1_n75), .ZN(
        npu_inst_pe_1_0_1_n31) );
  AOI222_X1 npu_inst_pe_1_0_1_U48 ( .A1(npu_inst_int_data_res_1__1__1_), .A2(
        npu_inst_pe_1_0_1_n1), .B1(npu_inst_pe_1_0_1_N74), .B2(
        npu_inst_pe_1_0_1_n76), .C1(npu_inst_pe_1_0_1_N66), .C2(
        npu_inst_pe_1_0_1_n77), .ZN(npu_inst_pe_1_0_1_n83) );
  INV_X1 npu_inst_pe_1_0_1_U47 ( .A(npu_inst_pe_1_0_1_n83), .ZN(
        npu_inst_pe_1_0_1_n98) );
  AOI222_X1 npu_inst_pe_1_0_1_U46 ( .A1(npu_inst_int_data_res_1__1__2_), .A2(
        npu_inst_pe_1_0_1_n1), .B1(npu_inst_pe_1_0_1_N75), .B2(
        npu_inst_pe_1_0_1_n76), .C1(npu_inst_pe_1_0_1_N67), .C2(
        npu_inst_pe_1_0_1_n77), .ZN(npu_inst_pe_1_0_1_n82) );
  INV_X1 npu_inst_pe_1_0_1_U45 ( .A(npu_inst_pe_1_0_1_n82), .ZN(
        npu_inst_pe_1_0_1_n36) );
  AOI222_X1 npu_inst_pe_1_0_1_U44 ( .A1(npu_inst_int_data_res_1__1__3_), .A2(
        npu_inst_pe_1_0_1_n1), .B1(npu_inst_pe_1_0_1_N76), .B2(
        npu_inst_pe_1_0_1_n76), .C1(npu_inst_pe_1_0_1_N68), .C2(
        npu_inst_pe_1_0_1_n77), .ZN(npu_inst_pe_1_0_1_n81) );
  INV_X1 npu_inst_pe_1_0_1_U43 ( .A(npu_inst_pe_1_0_1_n81), .ZN(
        npu_inst_pe_1_0_1_n35) );
  AOI222_X1 npu_inst_pe_1_0_1_U42 ( .A1(npu_inst_int_data_res_1__1__4_), .A2(
        npu_inst_pe_1_0_1_n1), .B1(npu_inst_pe_1_0_1_N77), .B2(
        npu_inst_pe_1_0_1_n76), .C1(npu_inst_pe_1_0_1_N69), .C2(
        npu_inst_pe_1_0_1_n77), .ZN(npu_inst_pe_1_0_1_n80) );
  INV_X1 npu_inst_pe_1_0_1_U41 ( .A(npu_inst_pe_1_0_1_n80), .ZN(
        npu_inst_pe_1_0_1_n34) );
  AOI222_X1 npu_inst_pe_1_0_1_U40 ( .A1(npu_inst_int_data_res_1__1__5_), .A2(
        npu_inst_pe_1_0_1_n1), .B1(npu_inst_pe_1_0_1_N78), .B2(
        npu_inst_pe_1_0_1_n76), .C1(npu_inst_pe_1_0_1_N70), .C2(
        npu_inst_pe_1_0_1_n77), .ZN(npu_inst_pe_1_0_1_n79) );
  INV_X1 npu_inst_pe_1_0_1_U39 ( .A(npu_inst_pe_1_0_1_n79), .ZN(
        npu_inst_pe_1_0_1_n33) );
  AOI222_X1 npu_inst_pe_1_0_1_U38 ( .A1(npu_inst_int_data_res_1__1__6_), .A2(
        npu_inst_pe_1_0_1_n1), .B1(npu_inst_pe_1_0_1_N79), .B2(
        npu_inst_pe_1_0_1_n76), .C1(npu_inst_pe_1_0_1_N71), .C2(
        npu_inst_pe_1_0_1_n77), .ZN(npu_inst_pe_1_0_1_n78) );
  INV_X1 npu_inst_pe_1_0_1_U37 ( .A(npu_inst_pe_1_0_1_n78), .ZN(
        npu_inst_pe_1_0_1_n32) );
  INV_X1 npu_inst_pe_1_0_1_U36 ( .A(npu_inst_pe_1_0_1_int_data_1_), .ZN(
        npu_inst_pe_1_0_1_n12) );
  AND2_X1 npu_inst_pe_1_0_1_U35 ( .A1(npu_inst_int_data_x_0__1__1_), .A2(
        npu_inst_pe_1_0_1_int_q_weight_1_), .ZN(npu_inst_pe_1_0_1_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_0_1_U34 ( .A1(npu_inst_int_data_x_0__1__0_), .A2(
        npu_inst_pe_1_0_1_int_q_weight_1_), .ZN(npu_inst_pe_1_0_1_int_data_0_)
         );
  AND2_X1 npu_inst_pe_1_0_1_U33 ( .A1(npu_inst_pe_1_0_1_N93), .A2(npu_inst_n60), .ZN(npu_inst_pe_1_0_1_o_data_v_0_) );
  AND2_X1 npu_inst_pe_1_0_1_U32 ( .A1(npu_inst_n60), .A2(npu_inst_pe_1_0_1_N94), .ZN(npu_inst_pe_1_0_1_o_data_v_1_) );
  AOI22_X1 npu_inst_pe_1_0_1_U31 ( .A1(npu_inst_n60), .A2(
        npu_inst_int_data_y_1__1__1_), .B1(npu_inst_pe_1_0_1_n3), .B2(
        npu_inst_int_data_x_0__2__1_), .ZN(npu_inst_pe_1_0_1_n63) );
  AOI22_X1 npu_inst_pe_1_0_1_U30 ( .A1(npu_inst_n60), .A2(
        npu_inst_int_data_y_1__1__0_), .B1(npu_inst_pe_1_0_1_n3), .B2(
        npu_inst_int_data_x_0__2__0_), .ZN(npu_inst_pe_1_0_1_n61) );
  INV_X1 npu_inst_pe_1_0_1_U29 ( .A(npu_inst_pe_1_0_1_int_data_0_), .ZN(
        npu_inst_pe_1_0_1_n11) );
  INV_X1 npu_inst_pe_1_0_1_U28 ( .A(npu_inst_n72), .ZN(npu_inst_pe_1_0_1_n4)
         );
  OR3_X1 npu_inst_pe_1_0_1_U27 ( .A1(npu_inst_n80), .A2(npu_inst_pe_1_0_1_n6), 
        .A3(npu_inst_pe_1_0_1_n4), .ZN(npu_inst_pe_1_0_1_n56) );
  OR3_X1 npu_inst_pe_1_0_1_U26 ( .A1(npu_inst_pe_1_0_1_n4), .A2(
        npu_inst_pe_1_0_1_n6), .A3(npu_inst_pe_1_0_1_n5), .ZN(
        npu_inst_pe_1_0_1_n48) );
  INV_X1 npu_inst_pe_1_0_1_U25 ( .A(npu_inst_n127), .ZN(npu_inst_pe_1_0_1_n10)
         );
  OR3_X1 npu_inst_pe_1_0_1_U24 ( .A1(npu_inst_n72), .A2(npu_inst_pe_1_0_1_n6), 
        .A3(npu_inst_pe_1_0_1_n5), .ZN(npu_inst_pe_1_0_1_n52) );
  OR3_X1 npu_inst_pe_1_0_1_U23 ( .A1(npu_inst_n80), .A2(npu_inst_pe_1_0_1_n6), 
        .A3(npu_inst_n72), .ZN(npu_inst_pe_1_0_1_n60) );
  NOR2_X1 npu_inst_pe_1_0_1_U22 ( .A1(npu_inst_pe_1_0_1_n60), .A2(
        npu_inst_pe_1_0_1_n3), .ZN(npu_inst_pe_1_0_1_n58) );
  NOR2_X1 npu_inst_pe_1_0_1_U21 ( .A1(npu_inst_pe_1_0_1_n56), .A2(
        npu_inst_pe_1_0_1_n3), .ZN(npu_inst_pe_1_0_1_n54) );
  NOR2_X1 npu_inst_pe_1_0_1_U20 ( .A1(npu_inst_pe_1_0_1_n52), .A2(
        npu_inst_pe_1_0_1_n3), .ZN(npu_inst_pe_1_0_1_n50) );
  NOR2_X1 npu_inst_pe_1_0_1_U19 ( .A1(npu_inst_pe_1_0_1_n48), .A2(
        npu_inst_pe_1_0_1_n3), .ZN(npu_inst_pe_1_0_1_n46) );
  NOR2_X1 npu_inst_pe_1_0_1_U18 ( .A1(npu_inst_pe_1_0_1_n40), .A2(
        npu_inst_pe_1_0_1_n3), .ZN(npu_inst_pe_1_0_1_n38) );
  NOR2_X1 npu_inst_pe_1_0_1_U17 ( .A1(npu_inst_pe_1_0_1_n44), .A2(
        npu_inst_pe_1_0_1_n3), .ZN(npu_inst_pe_1_0_1_n42) );
  BUF_X1 npu_inst_pe_1_0_1_U16 ( .A(npu_inst_n107), .Z(npu_inst_pe_1_0_1_n6)
         );
  BUF_X1 npu_inst_pe_1_0_1_U15 ( .A(npu_inst_pe_1_0_1_n10), .Z(
        npu_inst_pe_1_0_1_n9) );
  BUF_X1 npu_inst_pe_1_0_1_U14 ( .A(npu_inst_pe_1_0_1_n10), .Z(
        npu_inst_pe_1_0_1_n8) );
  BUF_X1 npu_inst_pe_1_0_1_U13 ( .A(npu_inst_pe_1_0_1_n10), .Z(
        npu_inst_pe_1_0_1_n7) );
  INV_X1 npu_inst_pe_1_0_1_U12 ( .A(npu_inst_pe_1_0_1_n38), .ZN(
        npu_inst_pe_1_0_1_n116) );
  INV_X1 npu_inst_pe_1_0_1_U11 ( .A(npu_inst_pe_1_0_1_n58), .ZN(
        npu_inst_pe_1_0_1_n112) );
  INV_X1 npu_inst_pe_1_0_1_U10 ( .A(npu_inst_pe_1_0_1_n54), .ZN(
        npu_inst_pe_1_0_1_n113) );
  INV_X1 npu_inst_pe_1_0_1_U9 ( .A(npu_inst_pe_1_0_1_n50), .ZN(
        npu_inst_pe_1_0_1_n114) );
  INV_X1 npu_inst_pe_1_0_1_U8 ( .A(npu_inst_pe_1_0_1_n46), .ZN(
        npu_inst_pe_1_0_1_n115) );
  INV_X1 npu_inst_pe_1_0_1_U7 ( .A(npu_inst_pe_1_0_1_n42), .ZN(
        npu_inst_pe_1_0_1_n117) );
  BUF_X1 npu_inst_pe_1_0_1_U6 ( .A(npu_inst_n38), .Z(npu_inst_pe_1_0_1_n2) );
  BUF_X1 npu_inst_pe_1_0_1_U5 ( .A(npu_inst_n38), .Z(npu_inst_pe_1_0_1_n1) );
  NOR2_X1 npu_inst_pe_1_0_1_U4 ( .A1(npu_inst_pe_1_0_1_int_q_weight_0_), .A2(
        npu_inst_pe_1_0_1_n1), .ZN(npu_inst_pe_1_0_1_n76) );
  NOR2_X1 npu_inst_pe_1_0_1_U3 ( .A1(npu_inst_pe_1_0_1_n27), .A2(
        npu_inst_pe_1_0_1_n1), .ZN(npu_inst_pe_1_0_1_n77) );
  FA_X1 npu_inst_pe_1_0_1_sub_77_U2_1 ( .A(npu_inst_pe_1_0_1_int_q_acc_1_), 
        .B(npu_inst_pe_1_0_1_n12), .CI(npu_inst_pe_1_0_1_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_0_1_sub_77_carry_2_), .S(npu_inst_pe_1_0_1_N66) );
  FA_X1 npu_inst_pe_1_0_1_add_79_U1_1 ( .A(npu_inst_pe_1_0_1_int_q_acc_1_), 
        .B(npu_inst_pe_1_0_1_int_data_1_), .CI(
        npu_inst_pe_1_0_1_add_79_carry_1_), .CO(
        npu_inst_pe_1_0_1_add_79_carry_2_), .S(npu_inst_pe_1_0_1_N74) );
  NAND3_X1 npu_inst_pe_1_0_1_U109 ( .A1(npu_inst_pe_1_0_1_n4), .A2(
        npu_inst_pe_1_0_1_n5), .A3(npu_inst_pe_1_0_1_n6), .ZN(
        npu_inst_pe_1_0_1_n44) );
  NAND3_X1 npu_inst_pe_1_0_1_U108 ( .A1(npu_inst_n72), .A2(
        npu_inst_pe_1_0_1_n5), .A3(npu_inst_pe_1_0_1_n6), .ZN(
        npu_inst_pe_1_0_1_n40) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_0_1_n32), .CK(
        npu_inst_pe_1_0_1_net4270), .RN(npu_inst_pe_1_0_1_n7), .Q(
        npu_inst_pe_1_0_1_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_0_1_n33), .CK(
        npu_inst_pe_1_0_1_net4270), .RN(npu_inst_pe_1_0_1_n7), .Q(
        npu_inst_pe_1_0_1_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_0_1_n34), .CK(
        npu_inst_pe_1_0_1_net4270), .RN(npu_inst_pe_1_0_1_n7), .Q(
        npu_inst_pe_1_0_1_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_0_1_n35), .CK(
        npu_inst_pe_1_0_1_net4270), .RN(npu_inst_pe_1_0_1_n7), .Q(
        npu_inst_pe_1_0_1_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_0_1_n36), .CK(
        npu_inst_pe_1_0_1_net4270), .RN(npu_inst_pe_1_0_1_n7), .Q(
        npu_inst_pe_1_0_1_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_0_1_n98), .CK(
        npu_inst_pe_1_0_1_net4270), .RN(npu_inst_pe_1_0_1_n7), .Q(
        npu_inst_pe_1_0_1_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_0_1_n31), .CK(
        npu_inst_pe_1_0_1_net4270), .RN(npu_inst_pe_1_0_1_n7), .Q(
        npu_inst_pe_1_0_1_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_0_1_n99), .CK(
        npu_inst_pe_1_0_1_net4270), .RN(npu_inst_pe_1_0_1_n7), .Q(
        npu_inst_pe_1_0_1_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_weight_reg_0_ ( .D(npu_inst_n113), .CK(
        npu_inst_pe_1_0_1_net4276), .RN(npu_inst_pe_1_0_1_n7), .Q(
        npu_inst_pe_1_0_1_int_q_weight_0_), .QN(npu_inst_pe_1_0_1_n27) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_weight_reg_1_ ( .D(npu_inst_n119), .CK(
        npu_inst_pe_1_0_1_net4276), .RN(npu_inst_pe_1_0_1_n7), .Q(
        npu_inst_pe_1_0_1_int_q_weight_1_), .QN(npu_inst_pe_1_0_1_n26) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_0_1_n111), 
        .CK(npu_inst_pe_1_0_1_net4276), .RN(npu_inst_pe_1_0_1_n7), .Q(
        npu_inst_pe_1_0_1_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_0_1_n105), 
        .CK(npu_inst_pe_1_0_1_net4276), .RN(npu_inst_pe_1_0_1_n7), .Q(
        npu_inst_pe_1_0_1_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_0_1_n110), 
        .CK(npu_inst_pe_1_0_1_net4276), .RN(npu_inst_pe_1_0_1_n8), .Q(
        npu_inst_pe_1_0_1_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_0_1_n104), 
        .CK(npu_inst_pe_1_0_1_net4276), .RN(npu_inst_pe_1_0_1_n8), .Q(
        npu_inst_pe_1_0_1_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_0_1_n109), 
        .CK(npu_inst_pe_1_0_1_net4276), .RN(npu_inst_pe_1_0_1_n8), .Q(
        npu_inst_pe_1_0_1_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_0_1_n103), 
        .CK(npu_inst_pe_1_0_1_net4276), .RN(npu_inst_pe_1_0_1_n8), .Q(
        npu_inst_pe_1_0_1_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_0_1_n108), 
        .CK(npu_inst_pe_1_0_1_net4276), .RN(npu_inst_pe_1_0_1_n8), .Q(
        npu_inst_pe_1_0_1_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_0_1_n102), 
        .CK(npu_inst_pe_1_0_1_net4276), .RN(npu_inst_pe_1_0_1_n8), .Q(
        npu_inst_pe_1_0_1_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_0_1_n107), 
        .CK(npu_inst_pe_1_0_1_net4276), .RN(npu_inst_pe_1_0_1_n8), .Q(
        npu_inst_pe_1_0_1_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_0_1_n101), 
        .CK(npu_inst_pe_1_0_1_net4276), .RN(npu_inst_pe_1_0_1_n8), .Q(
        npu_inst_pe_1_0_1_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_0_1_n106), 
        .CK(npu_inst_pe_1_0_1_net4276), .RN(npu_inst_pe_1_0_1_n8), .Q(
        npu_inst_pe_1_0_1_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_0_1_n100), 
        .CK(npu_inst_pe_1_0_1_net4276), .RN(npu_inst_pe_1_0_1_n8), .Q(
        npu_inst_pe_1_0_1_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_0_1_n86), 
        .CK(npu_inst_pe_1_0_1_net4276), .RN(npu_inst_pe_1_0_1_n8), .Q(
        npu_inst_pe_1_0_1_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_0_1_n87), 
        .CK(npu_inst_pe_1_0_1_net4276), .RN(npu_inst_pe_1_0_1_n8), .Q(
        npu_inst_pe_1_0_1_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_0_1_n88), 
        .CK(npu_inst_pe_1_0_1_net4276), .RN(npu_inst_pe_1_0_1_n9), .Q(
        npu_inst_pe_1_0_1_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_0_1_n89), 
        .CK(npu_inst_pe_1_0_1_net4276), .RN(npu_inst_pe_1_0_1_n9), .Q(
        npu_inst_pe_1_0_1_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_0_1_n90), 
        .CK(npu_inst_pe_1_0_1_net4276), .RN(npu_inst_pe_1_0_1_n9), .Q(
        npu_inst_pe_1_0_1_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_0_1_n91), 
        .CK(npu_inst_pe_1_0_1_net4276), .RN(npu_inst_pe_1_0_1_n9), .Q(
        npu_inst_pe_1_0_1_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_0_1_n92), 
        .CK(npu_inst_pe_1_0_1_net4276), .RN(npu_inst_pe_1_0_1_n9), .Q(
        npu_inst_pe_1_0_1_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_0_1_n93), 
        .CK(npu_inst_pe_1_0_1_net4276), .RN(npu_inst_pe_1_0_1_n9), .Q(
        npu_inst_pe_1_0_1_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_0_1_n94), 
        .CK(npu_inst_pe_1_0_1_net4276), .RN(npu_inst_pe_1_0_1_n9), .Q(
        npu_inst_pe_1_0_1_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_0_1_n95), 
        .CK(npu_inst_pe_1_0_1_net4276), .RN(npu_inst_pe_1_0_1_n9), .Q(
        npu_inst_pe_1_0_1_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_0_1_n96), 
        .CK(npu_inst_pe_1_0_1_net4276), .RN(npu_inst_pe_1_0_1_n9), .Q(
        npu_inst_pe_1_0_1_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_0_1_n97), 
        .CK(npu_inst_pe_1_0_1_net4276), .RN(npu_inst_pe_1_0_1_n9), .Q(
        npu_inst_pe_1_0_1_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_0_1_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_0_1_N84), .SE(1'b0), .GCK(npu_inst_pe_1_0_1_net4270) );
  CLKGATETST_X1 npu_inst_pe_1_0_1_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n66), .SE(1'b0), .GCK(npu_inst_pe_1_0_1_net4276) );
  MUX2_X1 npu_inst_pe_1_0_2_U161 ( .A(npu_inst_pe_1_0_2_n31), .B(
        npu_inst_pe_1_0_2_n28), .S(npu_inst_pe_1_0_2_n7), .Z(
        npu_inst_pe_1_0_2_N93) );
  MUX2_X1 npu_inst_pe_1_0_2_U160 ( .A(npu_inst_pe_1_0_2_n30), .B(
        npu_inst_pe_1_0_2_n29), .S(npu_inst_n80), .Z(npu_inst_pe_1_0_2_n31) );
  MUX2_X1 npu_inst_pe_1_0_2_U159 ( .A(npu_inst_pe_1_0_2_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_0_2_int_q_reg_v_1__0_), .S(npu_inst_pe_1_0_2_n4), .Z(
        npu_inst_pe_1_0_2_n30) );
  MUX2_X1 npu_inst_pe_1_0_2_U158 ( .A(npu_inst_pe_1_0_2_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_0_2_int_q_reg_v_3__0_), .S(npu_inst_pe_1_0_2_n4), .Z(
        npu_inst_pe_1_0_2_n29) );
  MUX2_X1 npu_inst_pe_1_0_2_U157 ( .A(npu_inst_pe_1_0_2_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_0_2_int_q_reg_v_5__0_), .S(npu_inst_pe_1_0_2_n4), .Z(
        npu_inst_pe_1_0_2_n28) );
  MUX2_X1 npu_inst_pe_1_0_2_U156 ( .A(npu_inst_pe_1_0_2_n25), .B(
        npu_inst_pe_1_0_2_n22), .S(npu_inst_pe_1_0_2_n7), .Z(
        npu_inst_pe_1_0_2_N94) );
  MUX2_X1 npu_inst_pe_1_0_2_U155 ( .A(npu_inst_pe_1_0_2_n24), .B(
        npu_inst_pe_1_0_2_n23), .S(npu_inst_n80), .Z(npu_inst_pe_1_0_2_n25) );
  MUX2_X1 npu_inst_pe_1_0_2_U154 ( .A(npu_inst_pe_1_0_2_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_0_2_int_q_reg_v_1__1_), .S(npu_inst_pe_1_0_2_n4), .Z(
        npu_inst_pe_1_0_2_n24) );
  MUX2_X1 npu_inst_pe_1_0_2_U153 ( .A(npu_inst_pe_1_0_2_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_0_2_int_q_reg_v_3__1_), .S(npu_inst_pe_1_0_2_n4), .Z(
        npu_inst_pe_1_0_2_n23) );
  MUX2_X1 npu_inst_pe_1_0_2_U152 ( .A(npu_inst_pe_1_0_2_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_0_2_int_q_reg_v_5__1_), .S(npu_inst_pe_1_0_2_n4), .Z(
        npu_inst_pe_1_0_2_n22) );
  MUX2_X1 npu_inst_pe_1_0_2_U151 ( .A(npu_inst_pe_1_0_2_n21), .B(
        npu_inst_pe_1_0_2_n18), .S(npu_inst_pe_1_0_2_n7), .Z(
        npu_inst_int_data_x_0__2__1_) );
  MUX2_X1 npu_inst_pe_1_0_2_U150 ( .A(npu_inst_pe_1_0_2_n20), .B(
        npu_inst_pe_1_0_2_n19), .S(npu_inst_n80), .Z(npu_inst_pe_1_0_2_n21) );
  MUX2_X1 npu_inst_pe_1_0_2_U149 ( .A(npu_inst_pe_1_0_2_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_0_2_int_q_reg_h_1__1_), .S(npu_inst_pe_1_0_2_n4), .Z(
        npu_inst_pe_1_0_2_n20) );
  MUX2_X1 npu_inst_pe_1_0_2_U148 ( .A(npu_inst_pe_1_0_2_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_0_2_int_q_reg_h_3__1_), .S(npu_inst_pe_1_0_2_n4), .Z(
        npu_inst_pe_1_0_2_n19) );
  MUX2_X1 npu_inst_pe_1_0_2_U147 ( .A(npu_inst_pe_1_0_2_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_0_2_int_q_reg_h_5__1_), .S(npu_inst_pe_1_0_2_n4), .Z(
        npu_inst_pe_1_0_2_n18) );
  MUX2_X1 npu_inst_pe_1_0_2_U146 ( .A(npu_inst_pe_1_0_2_n17), .B(
        npu_inst_pe_1_0_2_n14), .S(npu_inst_pe_1_0_2_n7), .Z(
        npu_inst_int_data_x_0__2__0_) );
  MUX2_X1 npu_inst_pe_1_0_2_U145 ( .A(npu_inst_pe_1_0_2_n16), .B(
        npu_inst_pe_1_0_2_n15), .S(npu_inst_n80), .Z(npu_inst_pe_1_0_2_n17) );
  MUX2_X1 npu_inst_pe_1_0_2_U144 ( .A(npu_inst_pe_1_0_2_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_0_2_int_q_reg_h_1__0_), .S(npu_inst_pe_1_0_2_n4), .Z(
        npu_inst_pe_1_0_2_n16) );
  MUX2_X1 npu_inst_pe_1_0_2_U143 ( .A(npu_inst_pe_1_0_2_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_0_2_int_q_reg_h_3__0_), .S(npu_inst_pe_1_0_2_n4), .Z(
        npu_inst_pe_1_0_2_n15) );
  MUX2_X1 npu_inst_pe_1_0_2_U142 ( .A(npu_inst_pe_1_0_2_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_0_2_int_q_reg_h_5__0_), .S(npu_inst_pe_1_0_2_n4), .Z(
        npu_inst_pe_1_0_2_n14) );
  XOR2_X1 npu_inst_pe_1_0_2_U141 ( .A(npu_inst_pe_1_0_2_int_data_0_), .B(
        npu_inst_pe_1_0_2_int_q_acc_0_), .Z(npu_inst_pe_1_0_2_N73) );
  AND2_X1 npu_inst_pe_1_0_2_U140 ( .A1(npu_inst_pe_1_0_2_int_q_acc_0_), .A2(
        npu_inst_pe_1_0_2_int_data_0_), .ZN(npu_inst_pe_1_0_2_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_0_2_U139 ( .A(npu_inst_pe_1_0_2_int_q_acc_0_), .B(
        npu_inst_pe_1_0_2_n12), .ZN(npu_inst_pe_1_0_2_N65) );
  OR2_X1 npu_inst_pe_1_0_2_U138 ( .A1(npu_inst_pe_1_0_2_n12), .A2(
        npu_inst_pe_1_0_2_int_q_acc_0_), .ZN(npu_inst_pe_1_0_2_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_0_2_U137 ( .A(npu_inst_pe_1_0_2_int_q_acc_2_), .B(
        npu_inst_pe_1_0_2_add_79_carry_2_), .Z(npu_inst_pe_1_0_2_N75) );
  AND2_X1 npu_inst_pe_1_0_2_U136 ( .A1(npu_inst_pe_1_0_2_add_79_carry_2_), 
        .A2(npu_inst_pe_1_0_2_int_q_acc_2_), .ZN(
        npu_inst_pe_1_0_2_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_0_2_U135 ( .A(npu_inst_pe_1_0_2_int_q_acc_3_), .B(
        npu_inst_pe_1_0_2_add_79_carry_3_), .Z(npu_inst_pe_1_0_2_N76) );
  AND2_X1 npu_inst_pe_1_0_2_U134 ( .A1(npu_inst_pe_1_0_2_add_79_carry_3_), 
        .A2(npu_inst_pe_1_0_2_int_q_acc_3_), .ZN(
        npu_inst_pe_1_0_2_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_0_2_U133 ( .A(npu_inst_pe_1_0_2_int_q_acc_4_), .B(
        npu_inst_pe_1_0_2_add_79_carry_4_), .Z(npu_inst_pe_1_0_2_N77) );
  AND2_X1 npu_inst_pe_1_0_2_U132 ( .A1(npu_inst_pe_1_0_2_add_79_carry_4_), 
        .A2(npu_inst_pe_1_0_2_int_q_acc_4_), .ZN(
        npu_inst_pe_1_0_2_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_0_2_U131 ( .A(npu_inst_pe_1_0_2_int_q_acc_5_), .B(
        npu_inst_pe_1_0_2_add_79_carry_5_), .Z(npu_inst_pe_1_0_2_N78) );
  AND2_X1 npu_inst_pe_1_0_2_U130 ( .A1(npu_inst_pe_1_0_2_add_79_carry_5_), 
        .A2(npu_inst_pe_1_0_2_int_q_acc_5_), .ZN(
        npu_inst_pe_1_0_2_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_0_2_U129 ( .A(npu_inst_pe_1_0_2_int_q_acc_6_), .B(
        npu_inst_pe_1_0_2_add_79_carry_6_), .Z(npu_inst_pe_1_0_2_N79) );
  AND2_X1 npu_inst_pe_1_0_2_U128 ( .A1(npu_inst_pe_1_0_2_add_79_carry_6_), 
        .A2(npu_inst_pe_1_0_2_int_q_acc_6_), .ZN(
        npu_inst_pe_1_0_2_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_0_2_U127 ( .A(npu_inst_pe_1_0_2_int_q_acc_7_), .B(
        npu_inst_pe_1_0_2_add_79_carry_7_), .Z(npu_inst_pe_1_0_2_N80) );
  XNOR2_X1 npu_inst_pe_1_0_2_U126 ( .A(npu_inst_pe_1_0_2_sub_77_carry_2_), .B(
        npu_inst_pe_1_0_2_int_q_acc_2_), .ZN(npu_inst_pe_1_0_2_N67) );
  OR2_X1 npu_inst_pe_1_0_2_U125 ( .A1(npu_inst_pe_1_0_2_int_q_acc_2_), .A2(
        npu_inst_pe_1_0_2_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_0_2_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_0_2_U124 ( .A(npu_inst_pe_1_0_2_sub_77_carry_3_), .B(
        npu_inst_pe_1_0_2_int_q_acc_3_), .ZN(npu_inst_pe_1_0_2_N68) );
  OR2_X1 npu_inst_pe_1_0_2_U123 ( .A1(npu_inst_pe_1_0_2_int_q_acc_3_), .A2(
        npu_inst_pe_1_0_2_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_0_2_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_0_2_U122 ( .A(npu_inst_pe_1_0_2_sub_77_carry_4_), .B(
        npu_inst_pe_1_0_2_int_q_acc_4_), .ZN(npu_inst_pe_1_0_2_N69) );
  OR2_X1 npu_inst_pe_1_0_2_U121 ( .A1(npu_inst_pe_1_0_2_int_q_acc_4_), .A2(
        npu_inst_pe_1_0_2_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_0_2_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_0_2_U120 ( .A(npu_inst_pe_1_0_2_sub_77_carry_5_), .B(
        npu_inst_pe_1_0_2_int_q_acc_5_), .ZN(npu_inst_pe_1_0_2_N70) );
  OR2_X1 npu_inst_pe_1_0_2_U119 ( .A1(npu_inst_pe_1_0_2_int_q_acc_5_), .A2(
        npu_inst_pe_1_0_2_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_0_2_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_0_2_U118 ( .A(npu_inst_pe_1_0_2_sub_77_carry_6_), .B(
        npu_inst_pe_1_0_2_int_q_acc_6_), .ZN(npu_inst_pe_1_0_2_N71) );
  OR2_X1 npu_inst_pe_1_0_2_U117 ( .A1(npu_inst_pe_1_0_2_int_q_acc_6_), .A2(
        npu_inst_pe_1_0_2_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_0_2_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_0_2_U116 ( .A(npu_inst_pe_1_0_2_int_q_acc_7_), .B(
        npu_inst_pe_1_0_2_sub_77_carry_7_), .ZN(npu_inst_pe_1_0_2_N72) );
  INV_X1 npu_inst_pe_1_0_2_U115 ( .A(npu_inst_n80), .ZN(npu_inst_pe_1_0_2_n6)
         );
  INV_X1 npu_inst_pe_1_0_2_U114 ( .A(npu_inst_n60), .ZN(npu_inst_pe_1_0_2_n3)
         );
  AOI22_X1 npu_inst_pe_1_0_2_U113 ( .A1(npu_inst_int_data_y_1__2__0_), .A2(
        npu_inst_pe_1_0_2_n58), .B1(npu_inst_pe_1_0_2_n113), .B2(
        npu_inst_pe_1_0_2_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_0_2_n57) );
  INV_X1 npu_inst_pe_1_0_2_U112 ( .A(npu_inst_pe_1_0_2_n57), .ZN(
        npu_inst_pe_1_0_2_n107) );
  AOI22_X1 npu_inst_pe_1_0_2_U111 ( .A1(npu_inst_int_data_y_1__2__0_), .A2(
        npu_inst_pe_1_0_2_n54), .B1(npu_inst_pe_1_0_2_n114), .B2(
        npu_inst_pe_1_0_2_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_0_2_n53) );
  INV_X1 npu_inst_pe_1_0_2_U110 ( .A(npu_inst_pe_1_0_2_n53), .ZN(
        npu_inst_pe_1_0_2_n108) );
  AOI22_X1 npu_inst_pe_1_0_2_U107 ( .A1(npu_inst_int_data_y_1__2__0_), .A2(
        npu_inst_pe_1_0_2_n50), .B1(npu_inst_pe_1_0_2_n115), .B2(
        npu_inst_pe_1_0_2_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_0_2_n49) );
  INV_X1 npu_inst_pe_1_0_2_U106 ( .A(npu_inst_pe_1_0_2_n49), .ZN(
        npu_inst_pe_1_0_2_n109) );
  AOI22_X1 npu_inst_pe_1_0_2_U105 ( .A1(npu_inst_int_data_y_1__2__0_), .A2(
        npu_inst_pe_1_0_2_n46), .B1(npu_inst_pe_1_0_2_n116), .B2(
        npu_inst_pe_1_0_2_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_0_2_n45) );
  INV_X1 npu_inst_pe_1_0_2_U104 ( .A(npu_inst_pe_1_0_2_n45), .ZN(
        npu_inst_pe_1_0_2_n110) );
  AOI22_X1 npu_inst_pe_1_0_2_U103 ( .A1(npu_inst_int_data_y_1__2__0_), .A2(
        npu_inst_pe_1_0_2_n42), .B1(npu_inst_pe_1_0_2_n118), .B2(
        npu_inst_pe_1_0_2_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_0_2_n41) );
  INV_X1 npu_inst_pe_1_0_2_U102 ( .A(npu_inst_pe_1_0_2_n41), .ZN(
        npu_inst_pe_1_0_2_n111) );
  AOI22_X1 npu_inst_pe_1_0_2_U101 ( .A1(npu_inst_int_data_y_1__2__1_), .A2(
        npu_inst_pe_1_0_2_n58), .B1(npu_inst_pe_1_0_2_n113), .B2(
        npu_inst_pe_1_0_2_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_0_2_n59) );
  INV_X1 npu_inst_pe_1_0_2_U100 ( .A(npu_inst_pe_1_0_2_n59), .ZN(
        npu_inst_pe_1_0_2_n101) );
  AOI22_X1 npu_inst_pe_1_0_2_U99 ( .A1(npu_inst_int_data_y_1__2__1_), .A2(
        npu_inst_pe_1_0_2_n54), .B1(npu_inst_pe_1_0_2_n114), .B2(
        npu_inst_pe_1_0_2_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_0_2_n55) );
  INV_X1 npu_inst_pe_1_0_2_U98 ( .A(npu_inst_pe_1_0_2_n55), .ZN(
        npu_inst_pe_1_0_2_n102) );
  AOI22_X1 npu_inst_pe_1_0_2_U97 ( .A1(npu_inst_int_data_y_1__2__1_), .A2(
        npu_inst_pe_1_0_2_n50), .B1(npu_inst_pe_1_0_2_n115), .B2(
        npu_inst_pe_1_0_2_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_0_2_n51) );
  INV_X1 npu_inst_pe_1_0_2_U96 ( .A(npu_inst_pe_1_0_2_n51), .ZN(
        npu_inst_pe_1_0_2_n103) );
  AOI22_X1 npu_inst_pe_1_0_2_U95 ( .A1(npu_inst_int_data_y_1__2__1_), .A2(
        npu_inst_pe_1_0_2_n46), .B1(npu_inst_pe_1_0_2_n116), .B2(
        npu_inst_pe_1_0_2_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_0_2_n47) );
  INV_X1 npu_inst_pe_1_0_2_U94 ( .A(npu_inst_pe_1_0_2_n47), .ZN(
        npu_inst_pe_1_0_2_n104) );
  AOI22_X1 npu_inst_pe_1_0_2_U93 ( .A1(npu_inst_int_data_y_1__2__1_), .A2(
        npu_inst_pe_1_0_2_n42), .B1(npu_inst_pe_1_0_2_n118), .B2(
        npu_inst_pe_1_0_2_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_0_2_n43) );
  INV_X1 npu_inst_pe_1_0_2_U92 ( .A(npu_inst_pe_1_0_2_n43), .ZN(
        npu_inst_pe_1_0_2_n105) );
  AOI22_X1 npu_inst_pe_1_0_2_U91 ( .A1(npu_inst_pe_1_0_2_n38), .A2(
        npu_inst_int_data_y_1__2__1_), .B1(npu_inst_pe_1_0_2_n117), .B2(
        npu_inst_pe_1_0_2_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_0_2_n39) );
  INV_X1 npu_inst_pe_1_0_2_U90 ( .A(npu_inst_pe_1_0_2_n39), .ZN(
        npu_inst_pe_1_0_2_n106) );
  AOI22_X1 npu_inst_pe_1_0_2_U89 ( .A1(npu_inst_pe_1_0_2_n38), .A2(
        npu_inst_int_data_y_1__2__0_), .B1(npu_inst_pe_1_0_2_n117), .B2(
        npu_inst_pe_1_0_2_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_0_2_n37) );
  INV_X1 npu_inst_pe_1_0_2_U88 ( .A(npu_inst_pe_1_0_2_n37), .ZN(
        npu_inst_pe_1_0_2_n112) );
  AND2_X1 npu_inst_pe_1_0_2_U87 ( .A1(npu_inst_pe_1_0_2_n2), .A2(
        npu_inst_pe_1_0_2_int_q_acc_7_), .ZN(o_data[47]) );
  AND2_X1 npu_inst_pe_1_0_2_U86 ( .A1(npu_inst_pe_1_0_2_int_q_acc_6_), .A2(
        npu_inst_pe_1_0_2_n2), .ZN(o_data[46]) );
  AND2_X1 npu_inst_pe_1_0_2_U85 ( .A1(npu_inst_pe_1_0_2_int_q_acc_5_), .A2(
        npu_inst_pe_1_0_2_n2), .ZN(o_data[45]) );
  AND2_X1 npu_inst_pe_1_0_2_U84 ( .A1(npu_inst_pe_1_0_2_int_q_acc_4_), .A2(
        npu_inst_pe_1_0_2_n2), .ZN(o_data[44]) );
  AND2_X1 npu_inst_pe_1_0_2_U83 ( .A1(npu_inst_pe_1_0_2_int_q_acc_3_), .A2(
        npu_inst_pe_1_0_2_n2), .ZN(o_data[43]) );
  NAND2_X1 npu_inst_pe_1_0_2_U82 ( .A1(npu_inst_pe_1_0_2_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_0_2_n60), .ZN(npu_inst_pe_1_0_2_n74) );
  OAI21_X1 npu_inst_pe_1_0_2_U81 ( .B1(npu_inst_pe_1_0_2_n63), .B2(
        npu_inst_pe_1_0_2_n60), .A(npu_inst_pe_1_0_2_n74), .ZN(
        npu_inst_pe_1_0_2_n97) );
  NAND2_X1 npu_inst_pe_1_0_2_U80 ( .A1(npu_inst_pe_1_0_2_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_0_2_n60), .ZN(npu_inst_pe_1_0_2_n73) );
  OAI21_X1 npu_inst_pe_1_0_2_U79 ( .B1(npu_inst_pe_1_0_2_n61), .B2(
        npu_inst_pe_1_0_2_n60), .A(npu_inst_pe_1_0_2_n73), .ZN(
        npu_inst_pe_1_0_2_n96) );
  NAND2_X1 npu_inst_pe_1_0_2_U78 ( .A1(npu_inst_pe_1_0_2_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_0_2_n56), .ZN(npu_inst_pe_1_0_2_n72) );
  OAI21_X1 npu_inst_pe_1_0_2_U77 ( .B1(npu_inst_pe_1_0_2_n63), .B2(
        npu_inst_pe_1_0_2_n56), .A(npu_inst_pe_1_0_2_n72), .ZN(
        npu_inst_pe_1_0_2_n95) );
  NAND2_X1 npu_inst_pe_1_0_2_U76 ( .A1(npu_inst_pe_1_0_2_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_0_2_n56), .ZN(npu_inst_pe_1_0_2_n71) );
  OAI21_X1 npu_inst_pe_1_0_2_U75 ( .B1(npu_inst_pe_1_0_2_n61), .B2(
        npu_inst_pe_1_0_2_n56), .A(npu_inst_pe_1_0_2_n71), .ZN(
        npu_inst_pe_1_0_2_n94) );
  NAND2_X1 npu_inst_pe_1_0_2_U74 ( .A1(npu_inst_pe_1_0_2_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_0_2_n52), .ZN(npu_inst_pe_1_0_2_n70) );
  OAI21_X1 npu_inst_pe_1_0_2_U73 ( .B1(npu_inst_pe_1_0_2_n63), .B2(
        npu_inst_pe_1_0_2_n52), .A(npu_inst_pe_1_0_2_n70), .ZN(
        npu_inst_pe_1_0_2_n93) );
  NAND2_X1 npu_inst_pe_1_0_2_U72 ( .A1(npu_inst_pe_1_0_2_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_0_2_n52), .ZN(npu_inst_pe_1_0_2_n69) );
  OAI21_X1 npu_inst_pe_1_0_2_U71 ( .B1(npu_inst_pe_1_0_2_n61), .B2(
        npu_inst_pe_1_0_2_n52), .A(npu_inst_pe_1_0_2_n69), .ZN(
        npu_inst_pe_1_0_2_n92) );
  NAND2_X1 npu_inst_pe_1_0_2_U70 ( .A1(npu_inst_pe_1_0_2_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_0_2_n48), .ZN(npu_inst_pe_1_0_2_n68) );
  OAI21_X1 npu_inst_pe_1_0_2_U69 ( .B1(npu_inst_pe_1_0_2_n63), .B2(
        npu_inst_pe_1_0_2_n48), .A(npu_inst_pe_1_0_2_n68), .ZN(
        npu_inst_pe_1_0_2_n91) );
  NAND2_X1 npu_inst_pe_1_0_2_U68 ( .A1(npu_inst_pe_1_0_2_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_0_2_n48), .ZN(npu_inst_pe_1_0_2_n67) );
  OAI21_X1 npu_inst_pe_1_0_2_U67 ( .B1(npu_inst_pe_1_0_2_n61), .B2(
        npu_inst_pe_1_0_2_n48), .A(npu_inst_pe_1_0_2_n67), .ZN(
        npu_inst_pe_1_0_2_n90) );
  NAND2_X1 npu_inst_pe_1_0_2_U66 ( .A1(npu_inst_pe_1_0_2_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_0_2_n44), .ZN(npu_inst_pe_1_0_2_n66) );
  OAI21_X1 npu_inst_pe_1_0_2_U65 ( .B1(npu_inst_pe_1_0_2_n63), .B2(
        npu_inst_pe_1_0_2_n44), .A(npu_inst_pe_1_0_2_n66), .ZN(
        npu_inst_pe_1_0_2_n89) );
  NAND2_X1 npu_inst_pe_1_0_2_U64 ( .A1(npu_inst_pe_1_0_2_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_0_2_n44), .ZN(npu_inst_pe_1_0_2_n65) );
  OAI21_X1 npu_inst_pe_1_0_2_U63 ( .B1(npu_inst_pe_1_0_2_n61), .B2(
        npu_inst_pe_1_0_2_n44), .A(npu_inst_pe_1_0_2_n65), .ZN(
        npu_inst_pe_1_0_2_n88) );
  NAND2_X1 npu_inst_pe_1_0_2_U62 ( .A1(npu_inst_pe_1_0_2_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_0_2_n40), .ZN(npu_inst_pe_1_0_2_n64) );
  OAI21_X1 npu_inst_pe_1_0_2_U61 ( .B1(npu_inst_pe_1_0_2_n63), .B2(
        npu_inst_pe_1_0_2_n40), .A(npu_inst_pe_1_0_2_n64), .ZN(
        npu_inst_pe_1_0_2_n87) );
  NAND2_X1 npu_inst_pe_1_0_2_U60 ( .A1(npu_inst_pe_1_0_2_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_0_2_n40), .ZN(npu_inst_pe_1_0_2_n62) );
  OAI21_X1 npu_inst_pe_1_0_2_U59 ( .B1(npu_inst_pe_1_0_2_n61), .B2(
        npu_inst_pe_1_0_2_n40), .A(npu_inst_pe_1_0_2_n62), .ZN(
        npu_inst_pe_1_0_2_n86) );
  NOR3_X1 npu_inst_pe_1_0_2_U58 ( .A1(npu_inst_pe_1_0_2_n26), .A2(npu_inst_n60), .A3(npu_inst_int_ckg[61]), .ZN(npu_inst_pe_1_0_2_n85) );
  OR2_X1 npu_inst_pe_1_0_2_U57 ( .A1(npu_inst_pe_1_0_2_n85), .A2(
        npu_inst_pe_1_0_2_n2), .ZN(npu_inst_pe_1_0_2_N84) );
  AND2_X1 npu_inst_pe_1_0_2_U56 ( .A1(npu_inst_pe_1_0_2_int_q_acc_0_), .A2(
        npu_inst_pe_1_0_2_n1), .ZN(o_data[40]) );
  AND2_X1 npu_inst_pe_1_0_2_U55 ( .A1(npu_inst_pe_1_0_2_int_q_acc_1_), .A2(
        npu_inst_pe_1_0_2_n1), .ZN(o_data[41]) );
  AND2_X1 npu_inst_pe_1_0_2_U54 ( .A1(npu_inst_pe_1_0_2_int_q_acc_2_), .A2(
        npu_inst_pe_1_0_2_n1), .ZN(o_data[42]) );
  AOI222_X1 npu_inst_pe_1_0_2_U53 ( .A1(npu_inst_int_data_res_1__2__0_), .A2(
        npu_inst_pe_1_0_2_n1), .B1(npu_inst_pe_1_0_2_N73), .B2(
        npu_inst_pe_1_0_2_n76), .C1(npu_inst_pe_1_0_2_N65), .C2(
        npu_inst_pe_1_0_2_n77), .ZN(npu_inst_pe_1_0_2_n84) );
  INV_X1 npu_inst_pe_1_0_2_U52 ( .A(npu_inst_pe_1_0_2_n84), .ZN(
        npu_inst_pe_1_0_2_n100) );
  AOI222_X1 npu_inst_pe_1_0_2_U51 ( .A1(npu_inst_int_data_res_1__2__7_), .A2(
        npu_inst_pe_1_0_2_n1), .B1(npu_inst_pe_1_0_2_N80), .B2(
        npu_inst_pe_1_0_2_n76), .C1(npu_inst_pe_1_0_2_N72), .C2(
        npu_inst_pe_1_0_2_n77), .ZN(npu_inst_pe_1_0_2_n75) );
  INV_X1 npu_inst_pe_1_0_2_U50 ( .A(npu_inst_pe_1_0_2_n75), .ZN(
        npu_inst_pe_1_0_2_n32) );
  AOI222_X1 npu_inst_pe_1_0_2_U49 ( .A1(npu_inst_int_data_res_1__2__1_), .A2(
        npu_inst_pe_1_0_2_n1), .B1(npu_inst_pe_1_0_2_N74), .B2(
        npu_inst_pe_1_0_2_n76), .C1(npu_inst_pe_1_0_2_N66), .C2(
        npu_inst_pe_1_0_2_n77), .ZN(npu_inst_pe_1_0_2_n83) );
  INV_X1 npu_inst_pe_1_0_2_U48 ( .A(npu_inst_pe_1_0_2_n83), .ZN(
        npu_inst_pe_1_0_2_n99) );
  AOI222_X1 npu_inst_pe_1_0_2_U47 ( .A1(npu_inst_int_data_res_1__2__2_), .A2(
        npu_inst_pe_1_0_2_n1), .B1(npu_inst_pe_1_0_2_N75), .B2(
        npu_inst_pe_1_0_2_n76), .C1(npu_inst_pe_1_0_2_N67), .C2(
        npu_inst_pe_1_0_2_n77), .ZN(npu_inst_pe_1_0_2_n82) );
  INV_X1 npu_inst_pe_1_0_2_U46 ( .A(npu_inst_pe_1_0_2_n82), .ZN(
        npu_inst_pe_1_0_2_n98) );
  AOI222_X1 npu_inst_pe_1_0_2_U45 ( .A1(npu_inst_int_data_res_1__2__3_), .A2(
        npu_inst_pe_1_0_2_n1), .B1(npu_inst_pe_1_0_2_N76), .B2(
        npu_inst_pe_1_0_2_n76), .C1(npu_inst_pe_1_0_2_N68), .C2(
        npu_inst_pe_1_0_2_n77), .ZN(npu_inst_pe_1_0_2_n81) );
  INV_X1 npu_inst_pe_1_0_2_U44 ( .A(npu_inst_pe_1_0_2_n81), .ZN(
        npu_inst_pe_1_0_2_n36) );
  AOI222_X1 npu_inst_pe_1_0_2_U43 ( .A1(npu_inst_int_data_res_1__2__4_), .A2(
        npu_inst_pe_1_0_2_n1), .B1(npu_inst_pe_1_0_2_N77), .B2(
        npu_inst_pe_1_0_2_n76), .C1(npu_inst_pe_1_0_2_N69), .C2(
        npu_inst_pe_1_0_2_n77), .ZN(npu_inst_pe_1_0_2_n80) );
  INV_X1 npu_inst_pe_1_0_2_U42 ( .A(npu_inst_pe_1_0_2_n80), .ZN(
        npu_inst_pe_1_0_2_n35) );
  AOI222_X1 npu_inst_pe_1_0_2_U41 ( .A1(npu_inst_int_data_res_1__2__5_), .A2(
        npu_inst_pe_1_0_2_n1), .B1(npu_inst_pe_1_0_2_N78), .B2(
        npu_inst_pe_1_0_2_n76), .C1(npu_inst_pe_1_0_2_N70), .C2(
        npu_inst_pe_1_0_2_n77), .ZN(npu_inst_pe_1_0_2_n79) );
  INV_X1 npu_inst_pe_1_0_2_U40 ( .A(npu_inst_pe_1_0_2_n79), .ZN(
        npu_inst_pe_1_0_2_n34) );
  AOI222_X1 npu_inst_pe_1_0_2_U39 ( .A1(npu_inst_int_data_res_1__2__6_), .A2(
        npu_inst_pe_1_0_2_n1), .B1(npu_inst_pe_1_0_2_N79), .B2(
        npu_inst_pe_1_0_2_n76), .C1(npu_inst_pe_1_0_2_N71), .C2(
        npu_inst_pe_1_0_2_n77), .ZN(npu_inst_pe_1_0_2_n78) );
  INV_X1 npu_inst_pe_1_0_2_U38 ( .A(npu_inst_pe_1_0_2_n78), .ZN(
        npu_inst_pe_1_0_2_n33) );
  INV_X1 npu_inst_pe_1_0_2_U37 ( .A(npu_inst_pe_1_0_2_int_data_1_), .ZN(
        npu_inst_pe_1_0_2_n13) );
  AND2_X1 npu_inst_pe_1_0_2_U36 ( .A1(npu_inst_int_data_x_0__2__1_), .A2(
        npu_inst_pe_1_0_2_int_q_weight_1_), .ZN(npu_inst_pe_1_0_2_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_0_2_U35 ( .A1(npu_inst_int_data_x_0__2__0_), .A2(
        npu_inst_pe_1_0_2_int_q_weight_1_), .ZN(npu_inst_pe_1_0_2_int_data_0_)
         );
  AND2_X1 npu_inst_pe_1_0_2_U34 ( .A1(npu_inst_pe_1_0_2_N93), .A2(npu_inst_n60), .ZN(npu_inst_pe_1_0_2_o_data_v_0_) );
  AND2_X1 npu_inst_pe_1_0_2_U33 ( .A1(npu_inst_n60), .A2(npu_inst_pe_1_0_2_N94), .ZN(npu_inst_pe_1_0_2_o_data_v_1_) );
  AOI22_X1 npu_inst_pe_1_0_2_U32 ( .A1(npu_inst_n60), .A2(
        npu_inst_int_data_y_1__2__1_), .B1(npu_inst_pe_1_0_2_n3), .B2(
        npu_inst_int_data_x_0__3__1_), .ZN(npu_inst_pe_1_0_2_n63) );
  AOI22_X1 npu_inst_pe_1_0_2_U31 ( .A1(npu_inst_n60), .A2(
        npu_inst_int_data_y_1__2__0_), .B1(npu_inst_pe_1_0_2_n3), .B2(
        npu_inst_int_data_x_0__3__0_), .ZN(npu_inst_pe_1_0_2_n61) );
  INV_X1 npu_inst_pe_1_0_2_U30 ( .A(npu_inst_pe_1_0_2_int_data_0_), .ZN(
        npu_inst_pe_1_0_2_n12) );
  INV_X1 npu_inst_pe_1_0_2_U29 ( .A(npu_inst_n72), .ZN(npu_inst_pe_1_0_2_n5)
         );
  OR3_X1 npu_inst_pe_1_0_2_U28 ( .A1(npu_inst_n80), .A2(npu_inst_pe_1_0_2_n7), 
        .A3(npu_inst_pe_1_0_2_n5), .ZN(npu_inst_pe_1_0_2_n56) );
  OR3_X1 npu_inst_pe_1_0_2_U27 ( .A1(npu_inst_pe_1_0_2_n5), .A2(
        npu_inst_pe_1_0_2_n7), .A3(npu_inst_pe_1_0_2_n6), .ZN(
        npu_inst_pe_1_0_2_n48) );
  INV_X1 npu_inst_pe_1_0_2_U26 ( .A(npu_inst_pe_1_0_2_n5), .ZN(
        npu_inst_pe_1_0_2_n4) );
  INV_X1 npu_inst_pe_1_0_2_U25 ( .A(npu_inst_n127), .ZN(npu_inst_pe_1_0_2_n11)
         );
  OR3_X1 npu_inst_pe_1_0_2_U24 ( .A1(npu_inst_pe_1_0_2_n4), .A2(
        npu_inst_pe_1_0_2_n7), .A3(npu_inst_pe_1_0_2_n6), .ZN(
        npu_inst_pe_1_0_2_n52) );
  OR3_X1 npu_inst_pe_1_0_2_U23 ( .A1(npu_inst_n80), .A2(npu_inst_pe_1_0_2_n7), 
        .A3(npu_inst_pe_1_0_2_n4), .ZN(npu_inst_pe_1_0_2_n60) );
  NOR2_X1 npu_inst_pe_1_0_2_U22 ( .A1(npu_inst_pe_1_0_2_n60), .A2(
        npu_inst_pe_1_0_2_n3), .ZN(npu_inst_pe_1_0_2_n58) );
  NOR2_X1 npu_inst_pe_1_0_2_U21 ( .A1(npu_inst_pe_1_0_2_n56), .A2(
        npu_inst_pe_1_0_2_n3), .ZN(npu_inst_pe_1_0_2_n54) );
  NOR2_X1 npu_inst_pe_1_0_2_U20 ( .A1(npu_inst_pe_1_0_2_n52), .A2(
        npu_inst_pe_1_0_2_n3), .ZN(npu_inst_pe_1_0_2_n50) );
  NOR2_X1 npu_inst_pe_1_0_2_U19 ( .A1(npu_inst_pe_1_0_2_n48), .A2(
        npu_inst_pe_1_0_2_n3), .ZN(npu_inst_pe_1_0_2_n46) );
  NOR2_X1 npu_inst_pe_1_0_2_U18 ( .A1(npu_inst_pe_1_0_2_n40), .A2(
        npu_inst_pe_1_0_2_n3), .ZN(npu_inst_pe_1_0_2_n38) );
  NOR2_X1 npu_inst_pe_1_0_2_U17 ( .A1(npu_inst_pe_1_0_2_n44), .A2(
        npu_inst_pe_1_0_2_n3), .ZN(npu_inst_pe_1_0_2_n42) );
  BUF_X1 npu_inst_pe_1_0_2_U16 ( .A(npu_inst_n107), .Z(npu_inst_pe_1_0_2_n7)
         );
  BUF_X1 npu_inst_pe_1_0_2_U15 ( .A(npu_inst_pe_1_0_2_n11), .Z(
        npu_inst_pe_1_0_2_n10) );
  BUF_X1 npu_inst_pe_1_0_2_U14 ( .A(npu_inst_pe_1_0_2_n11), .Z(
        npu_inst_pe_1_0_2_n9) );
  BUF_X1 npu_inst_pe_1_0_2_U13 ( .A(npu_inst_pe_1_0_2_n11), .Z(
        npu_inst_pe_1_0_2_n8) );
  INV_X1 npu_inst_pe_1_0_2_U12 ( .A(npu_inst_pe_1_0_2_n38), .ZN(
        npu_inst_pe_1_0_2_n117) );
  INV_X1 npu_inst_pe_1_0_2_U11 ( .A(npu_inst_pe_1_0_2_n58), .ZN(
        npu_inst_pe_1_0_2_n113) );
  INV_X1 npu_inst_pe_1_0_2_U10 ( .A(npu_inst_pe_1_0_2_n54), .ZN(
        npu_inst_pe_1_0_2_n114) );
  INV_X1 npu_inst_pe_1_0_2_U9 ( .A(npu_inst_pe_1_0_2_n50), .ZN(
        npu_inst_pe_1_0_2_n115) );
  INV_X1 npu_inst_pe_1_0_2_U8 ( .A(npu_inst_pe_1_0_2_n46), .ZN(
        npu_inst_pe_1_0_2_n116) );
  INV_X1 npu_inst_pe_1_0_2_U7 ( .A(npu_inst_pe_1_0_2_n42), .ZN(
        npu_inst_pe_1_0_2_n118) );
  BUF_X1 npu_inst_pe_1_0_2_U6 ( .A(npu_inst_n37), .Z(npu_inst_pe_1_0_2_n2) );
  BUF_X1 npu_inst_pe_1_0_2_U5 ( .A(npu_inst_n37), .Z(npu_inst_pe_1_0_2_n1) );
  NOR2_X1 npu_inst_pe_1_0_2_U4 ( .A1(npu_inst_pe_1_0_2_int_q_weight_0_), .A2(
        npu_inst_pe_1_0_2_n1), .ZN(npu_inst_pe_1_0_2_n76) );
  NOR2_X1 npu_inst_pe_1_0_2_U3 ( .A1(npu_inst_pe_1_0_2_n27), .A2(
        npu_inst_pe_1_0_2_n1), .ZN(npu_inst_pe_1_0_2_n77) );
  FA_X1 npu_inst_pe_1_0_2_sub_77_U2_1 ( .A(npu_inst_pe_1_0_2_int_q_acc_1_), 
        .B(npu_inst_pe_1_0_2_n13), .CI(npu_inst_pe_1_0_2_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_0_2_sub_77_carry_2_), .S(npu_inst_pe_1_0_2_N66) );
  FA_X1 npu_inst_pe_1_0_2_add_79_U1_1 ( .A(npu_inst_pe_1_0_2_int_q_acc_1_), 
        .B(npu_inst_pe_1_0_2_int_data_1_), .CI(
        npu_inst_pe_1_0_2_add_79_carry_1_), .CO(
        npu_inst_pe_1_0_2_add_79_carry_2_), .S(npu_inst_pe_1_0_2_N74) );
  NAND3_X1 npu_inst_pe_1_0_2_U109 ( .A1(npu_inst_pe_1_0_2_n5), .A2(
        npu_inst_pe_1_0_2_n6), .A3(npu_inst_pe_1_0_2_n7), .ZN(
        npu_inst_pe_1_0_2_n44) );
  NAND3_X1 npu_inst_pe_1_0_2_U108 ( .A1(npu_inst_pe_1_0_2_n4), .A2(
        npu_inst_pe_1_0_2_n6), .A3(npu_inst_pe_1_0_2_n7), .ZN(
        npu_inst_pe_1_0_2_n40) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_0_2_n33), .CK(
        npu_inst_pe_1_0_2_net4247), .RN(npu_inst_pe_1_0_2_n8), .Q(
        npu_inst_pe_1_0_2_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_0_2_n34), .CK(
        npu_inst_pe_1_0_2_net4247), .RN(npu_inst_pe_1_0_2_n8), .Q(
        npu_inst_pe_1_0_2_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_0_2_n35), .CK(
        npu_inst_pe_1_0_2_net4247), .RN(npu_inst_pe_1_0_2_n8), .Q(
        npu_inst_pe_1_0_2_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_0_2_n36), .CK(
        npu_inst_pe_1_0_2_net4247), .RN(npu_inst_pe_1_0_2_n8), .Q(
        npu_inst_pe_1_0_2_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_0_2_n98), .CK(
        npu_inst_pe_1_0_2_net4247), .RN(npu_inst_pe_1_0_2_n8), .Q(
        npu_inst_pe_1_0_2_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_0_2_n99), .CK(
        npu_inst_pe_1_0_2_net4247), .RN(npu_inst_pe_1_0_2_n8), .Q(
        npu_inst_pe_1_0_2_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_0_2_n32), .CK(
        npu_inst_pe_1_0_2_net4247), .RN(npu_inst_pe_1_0_2_n8), .Q(
        npu_inst_pe_1_0_2_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_0_2_n100), 
        .CK(npu_inst_pe_1_0_2_net4247), .RN(npu_inst_pe_1_0_2_n8), .Q(
        npu_inst_pe_1_0_2_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_weight_reg_0_ ( .D(npu_inst_n113), .CK(
        npu_inst_pe_1_0_2_net4253), .RN(npu_inst_pe_1_0_2_n8), .Q(
        npu_inst_pe_1_0_2_int_q_weight_0_), .QN(npu_inst_pe_1_0_2_n27) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_weight_reg_1_ ( .D(npu_inst_n119), .CK(
        npu_inst_pe_1_0_2_net4253), .RN(npu_inst_pe_1_0_2_n8), .Q(
        npu_inst_pe_1_0_2_int_q_weight_1_), .QN(npu_inst_pe_1_0_2_n26) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_0_2_n112), 
        .CK(npu_inst_pe_1_0_2_net4253), .RN(npu_inst_pe_1_0_2_n8), .Q(
        npu_inst_pe_1_0_2_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_0_2_n106), 
        .CK(npu_inst_pe_1_0_2_net4253), .RN(npu_inst_pe_1_0_2_n8), .Q(
        npu_inst_pe_1_0_2_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_0_2_n111), 
        .CK(npu_inst_pe_1_0_2_net4253), .RN(npu_inst_pe_1_0_2_n9), .Q(
        npu_inst_pe_1_0_2_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_0_2_n105), 
        .CK(npu_inst_pe_1_0_2_net4253), .RN(npu_inst_pe_1_0_2_n9), .Q(
        npu_inst_pe_1_0_2_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_0_2_n110), 
        .CK(npu_inst_pe_1_0_2_net4253), .RN(npu_inst_pe_1_0_2_n9), .Q(
        npu_inst_pe_1_0_2_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_0_2_n104), 
        .CK(npu_inst_pe_1_0_2_net4253), .RN(npu_inst_pe_1_0_2_n9), .Q(
        npu_inst_pe_1_0_2_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_0_2_n109), 
        .CK(npu_inst_pe_1_0_2_net4253), .RN(npu_inst_pe_1_0_2_n9), .Q(
        npu_inst_pe_1_0_2_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_0_2_n103), 
        .CK(npu_inst_pe_1_0_2_net4253), .RN(npu_inst_pe_1_0_2_n9), .Q(
        npu_inst_pe_1_0_2_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_0_2_n108), 
        .CK(npu_inst_pe_1_0_2_net4253), .RN(npu_inst_pe_1_0_2_n9), .Q(
        npu_inst_pe_1_0_2_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_0_2_n102), 
        .CK(npu_inst_pe_1_0_2_net4253), .RN(npu_inst_pe_1_0_2_n9), .Q(
        npu_inst_pe_1_0_2_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_0_2_n107), 
        .CK(npu_inst_pe_1_0_2_net4253), .RN(npu_inst_pe_1_0_2_n9), .Q(
        npu_inst_pe_1_0_2_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_0_2_n101), 
        .CK(npu_inst_pe_1_0_2_net4253), .RN(npu_inst_pe_1_0_2_n9), .Q(
        npu_inst_pe_1_0_2_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_0_2_n86), 
        .CK(npu_inst_pe_1_0_2_net4253), .RN(npu_inst_pe_1_0_2_n9), .Q(
        npu_inst_pe_1_0_2_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_0_2_n87), 
        .CK(npu_inst_pe_1_0_2_net4253), .RN(npu_inst_pe_1_0_2_n9), .Q(
        npu_inst_pe_1_0_2_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_0_2_n88), 
        .CK(npu_inst_pe_1_0_2_net4253), .RN(npu_inst_pe_1_0_2_n10), .Q(
        npu_inst_pe_1_0_2_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_0_2_n89), 
        .CK(npu_inst_pe_1_0_2_net4253), .RN(npu_inst_pe_1_0_2_n10), .Q(
        npu_inst_pe_1_0_2_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_0_2_n90), 
        .CK(npu_inst_pe_1_0_2_net4253), .RN(npu_inst_pe_1_0_2_n10), .Q(
        npu_inst_pe_1_0_2_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_0_2_n91), 
        .CK(npu_inst_pe_1_0_2_net4253), .RN(npu_inst_pe_1_0_2_n10), .Q(
        npu_inst_pe_1_0_2_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_0_2_n92), 
        .CK(npu_inst_pe_1_0_2_net4253), .RN(npu_inst_pe_1_0_2_n10), .Q(
        npu_inst_pe_1_0_2_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_0_2_n93), 
        .CK(npu_inst_pe_1_0_2_net4253), .RN(npu_inst_pe_1_0_2_n10), .Q(
        npu_inst_pe_1_0_2_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_0_2_n94), 
        .CK(npu_inst_pe_1_0_2_net4253), .RN(npu_inst_pe_1_0_2_n10), .Q(
        npu_inst_pe_1_0_2_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_0_2_n95), 
        .CK(npu_inst_pe_1_0_2_net4253), .RN(npu_inst_pe_1_0_2_n10), .Q(
        npu_inst_pe_1_0_2_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_0_2_n96), 
        .CK(npu_inst_pe_1_0_2_net4253), .RN(npu_inst_pe_1_0_2_n10), .Q(
        npu_inst_pe_1_0_2_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_0_2_n97), 
        .CK(npu_inst_pe_1_0_2_net4253), .RN(npu_inst_pe_1_0_2_n10), .Q(
        npu_inst_pe_1_0_2_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_0_2_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_0_2_N84), .SE(1'b0), .GCK(npu_inst_pe_1_0_2_net4247) );
  CLKGATETST_X1 npu_inst_pe_1_0_2_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n66), .SE(1'b0), .GCK(npu_inst_pe_1_0_2_net4253) );
  MUX2_X1 npu_inst_pe_1_0_3_U162 ( .A(npu_inst_pe_1_0_3_n32), .B(
        npu_inst_pe_1_0_3_n29), .S(npu_inst_pe_1_0_3_n8), .Z(
        npu_inst_pe_1_0_3_N93) );
  MUX2_X1 npu_inst_pe_1_0_3_U161 ( .A(npu_inst_pe_1_0_3_n31), .B(
        npu_inst_pe_1_0_3_n30), .S(npu_inst_pe_1_0_3_n6), .Z(
        npu_inst_pe_1_0_3_n32) );
  MUX2_X1 npu_inst_pe_1_0_3_U160 ( .A(npu_inst_pe_1_0_3_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_0_3_int_q_reg_v_1__0_), .S(npu_inst_pe_1_0_3_n4), .Z(
        npu_inst_pe_1_0_3_n31) );
  MUX2_X1 npu_inst_pe_1_0_3_U159 ( .A(npu_inst_pe_1_0_3_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_0_3_int_q_reg_v_3__0_), .S(npu_inst_pe_1_0_3_n4), .Z(
        npu_inst_pe_1_0_3_n30) );
  MUX2_X1 npu_inst_pe_1_0_3_U158 ( .A(npu_inst_pe_1_0_3_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_0_3_int_q_reg_v_5__0_), .S(npu_inst_pe_1_0_3_n4), .Z(
        npu_inst_pe_1_0_3_n29) );
  MUX2_X1 npu_inst_pe_1_0_3_U157 ( .A(npu_inst_pe_1_0_3_n28), .B(
        npu_inst_pe_1_0_3_n23), .S(npu_inst_pe_1_0_3_n8), .Z(
        npu_inst_pe_1_0_3_N94) );
  MUX2_X1 npu_inst_pe_1_0_3_U156 ( .A(npu_inst_pe_1_0_3_n25), .B(
        npu_inst_pe_1_0_3_n24), .S(npu_inst_pe_1_0_3_n6), .Z(
        npu_inst_pe_1_0_3_n28) );
  MUX2_X1 npu_inst_pe_1_0_3_U155 ( .A(npu_inst_pe_1_0_3_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_0_3_int_q_reg_v_1__1_), .S(npu_inst_pe_1_0_3_n4), .Z(
        npu_inst_pe_1_0_3_n25) );
  MUX2_X1 npu_inst_pe_1_0_3_U154 ( .A(npu_inst_pe_1_0_3_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_0_3_int_q_reg_v_3__1_), .S(npu_inst_pe_1_0_3_n4), .Z(
        npu_inst_pe_1_0_3_n24) );
  MUX2_X1 npu_inst_pe_1_0_3_U153 ( .A(npu_inst_pe_1_0_3_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_0_3_int_q_reg_v_5__1_), .S(npu_inst_pe_1_0_3_n4), .Z(
        npu_inst_pe_1_0_3_n23) );
  MUX2_X1 npu_inst_pe_1_0_3_U152 ( .A(npu_inst_pe_1_0_3_n22), .B(
        npu_inst_pe_1_0_3_n19), .S(npu_inst_pe_1_0_3_n8), .Z(
        npu_inst_int_data_x_0__3__1_) );
  MUX2_X1 npu_inst_pe_1_0_3_U151 ( .A(npu_inst_pe_1_0_3_n21), .B(
        npu_inst_pe_1_0_3_n20), .S(npu_inst_pe_1_0_3_n6), .Z(
        npu_inst_pe_1_0_3_n22) );
  MUX2_X1 npu_inst_pe_1_0_3_U150 ( .A(npu_inst_pe_1_0_3_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_0_3_int_q_reg_h_1__1_), .S(npu_inst_pe_1_0_3_n4), .Z(
        npu_inst_pe_1_0_3_n21) );
  MUX2_X1 npu_inst_pe_1_0_3_U149 ( .A(npu_inst_pe_1_0_3_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_0_3_int_q_reg_h_3__1_), .S(npu_inst_pe_1_0_3_n4), .Z(
        npu_inst_pe_1_0_3_n20) );
  MUX2_X1 npu_inst_pe_1_0_3_U148 ( .A(npu_inst_pe_1_0_3_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_0_3_int_q_reg_h_5__1_), .S(npu_inst_pe_1_0_3_n4), .Z(
        npu_inst_pe_1_0_3_n19) );
  MUX2_X1 npu_inst_pe_1_0_3_U147 ( .A(npu_inst_pe_1_0_3_n18), .B(
        npu_inst_pe_1_0_3_n15), .S(npu_inst_pe_1_0_3_n8), .Z(
        npu_inst_int_data_x_0__3__0_) );
  MUX2_X1 npu_inst_pe_1_0_3_U146 ( .A(npu_inst_pe_1_0_3_n17), .B(
        npu_inst_pe_1_0_3_n16), .S(npu_inst_pe_1_0_3_n6), .Z(
        npu_inst_pe_1_0_3_n18) );
  MUX2_X1 npu_inst_pe_1_0_3_U145 ( .A(npu_inst_pe_1_0_3_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_0_3_int_q_reg_h_1__0_), .S(npu_inst_pe_1_0_3_n4), .Z(
        npu_inst_pe_1_0_3_n17) );
  MUX2_X1 npu_inst_pe_1_0_3_U144 ( .A(npu_inst_pe_1_0_3_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_0_3_int_q_reg_h_3__0_), .S(npu_inst_pe_1_0_3_n4), .Z(
        npu_inst_pe_1_0_3_n16) );
  MUX2_X1 npu_inst_pe_1_0_3_U143 ( .A(npu_inst_pe_1_0_3_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_0_3_int_q_reg_h_5__0_), .S(npu_inst_pe_1_0_3_n4), .Z(
        npu_inst_pe_1_0_3_n15) );
  XOR2_X1 npu_inst_pe_1_0_3_U142 ( .A(npu_inst_pe_1_0_3_int_data_0_), .B(
        npu_inst_pe_1_0_3_int_q_acc_0_), .Z(npu_inst_pe_1_0_3_N73) );
  AND2_X1 npu_inst_pe_1_0_3_U141 ( .A1(npu_inst_pe_1_0_3_int_q_acc_0_), .A2(
        npu_inst_pe_1_0_3_int_data_0_), .ZN(npu_inst_pe_1_0_3_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_0_3_U140 ( .A(npu_inst_pe_1_0_3_int_q_acc_0_), .B(
        npu_inst_pe_1_0_3_n13), .ZN(npu_inst_pe_1_0_3_N65) );
  OR2_X1 npu_inst_pe_1_0_3_U139 ( .A1(npu_inst_pe_1_0_3_n13), .A2(
        npu_inst_pe_1_0_3_int_q_acc_0_), .ZN(npu_inst_pe_1_0_3_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_0_3_U138 ( .A(npu_inst_pe_1_0_3_int_q_acc_2_), .B(
        npu_inst_pe_1_0_3_add_79_carry_2_), .Z(npu_inst_pe_1_0_3_N75) );
  AND2_X1 npu_inst_pe_1_0_3_U137 ( .A1(npu_inst_pe_1_0_3_add_79_carry_2_), 
        .A2(npu_inst_pe_1_0_3_int_q_acc_2_), .ZN(
        npu_inst_pe_1_0_3_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_0_3_U136 ( .A(npu_inst_pe_1_0_3_int_q_acc_3_), .B(
        npu_inst_pe_1_0_3_add_79_carry_3_), .Z(npu_inst_pe_1_0_3_N76) );
  AND2_X1 npu_inst_pe_1_0_3_U135 ( .A1(npu_inst_pe_1_0_3_add_79_carry_3_), 
        .A2(npu_inst_pe_1_0_3_int_q_acc_3_), .ZN(
        npu_inst_pe_1_0_3_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_0_3_U134 ( .A(npu_inst_pe_1_0_3_int_q_acc_4_), .B(
        npu_inst_pe_1_0_3_add_79_carry_4_), .Z(npu_inst_pe_1_0_3_N77) );
  AND2_X1 npu_inst_pe_1_0_3_U133 ( .A1(npu_inst_pe_1_0_3_add_79_carry_4_), 
        .A2(npu_inst_pe_1_0_3_int_q_acc_4_), .ZN(
        npu_inst_pe_1_0_3_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_0_3_U132 ( .A(npu_inst_pe_1_0_3_int_q_acc_5_), .B(
        npu_inst_pe_1_0_3_add_79_carry_5_), .Z(npu_inst_pe_1_0_3_N78) );
  AND2_X1 npu_inst_pe_1_0_3_U131 ( .A1(npu_inst_pe_1_0_3_add_79_carry_5_), 
        .A2(npu_inst_pe_1_0_3_int_q_acc_5_), .ZN(
        npu_inst_pe_1_0_3_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_0_3_U130 ( .A(npu_inst_pe_1_0_3_int_q_acc_6_), .B(
        npu_inst_pe_1_0_3_add_79_carry_6_), .Z(npu_inst_pe_1_0_3_N79) );
  AND2_X1 npu_inst_pe_1_0_3_U129 ( .A1(npu_inst_pe_1_0_3_add_79_carry_6_), 
        .A2(npu_inst_pe_1_0_3_int_q_acc_6_), .ZN(
        npu_inst_pe_1_0_3_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_0_3_U128 ( .A(npu_inst_pe_1_0_3_int_q_acc_7_), .B(
        npu_inst_pe_1_0_3_add_79_carry_7_), .Z(npu_inst_pe_1_0_3_N80) );
  XNOR2_X1 npu_inst_pe_1_0_3_U127 ( .A(npu_inst_pe_1_0_3_sub_77_carry_2_), .B(
        npu_inst_pe_1_0_3_int_q_acc_2_), .ZN(npu_inst_pe_1_0_3_N67) );
  OR2_X1 npu_inst_pe_1_0_3_U126 ( .A1(npu_inst_pe_1_0_3_int_q_acc_2_), .A2(
        npu_inst_pe_1_0_3_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_0_3_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_0_3_U125 ( .A(npu_inst_pe_1_0_3_sub_77_carry_3_), .B(
        npu_inst_pe_1_0_3_int_q_acc_3_), .ZN(npu_inst_pe_1_0_3_N68) );
  OR2_X1 npu_inst_pe_1_0_3_U124 ( .A1(npu_inst_pe_1_0_3_int_q_acc_3_), .A2(
        npu_inst_pe_1_0_3_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_0_3_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_0_3_U123 ( .A(npu_inst_pe_1_0_3_sub_77_carry_4_), .B(
        npu_inst_pe_1_0_3_int_q_acc_4_), .ZN(npu_inst_pe_1_0_3_N69) );
  OR2_X1 npu_inst_pe_1_0_3_U122 ( .A1(npu_inst_pe_1_0_3_int_q_acc_4_), .A2(
        npu_inst_pe_1_0_3_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_0_3_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_0_3_U121 ( .A(npu_inst_pe_1_0_3_sub_77_carry_5_), .B(
        npu_inst_pe_1_0_3_int_q_acc_5_), .ZN(npu_inst_pe_1_0_3_N70) );
  OR2_X1 npu_inst_pe_1_0_3_U120 ( .A1(npu_inst_pe_1_0_3_int_q_acc_5_), .A2(
        npu_inst_pe_1_0_3_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_0_3_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_0_3_U119 ( .A(npu_inst_pe_1_0_3_sub_77_carry_6_), .B(
        npu_inst_pe_1_0_3_int_q_acc_6_), .ZN(npu_inst_pe_1_0_3_N71) );
  OR2_X1 npu_inst_pe_1_0_3_U118 ( .A1(npu_inst_pe_1_0_3_int_q_acc_6_), .A2(
        npu_inst_pe_1_0_3_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_0_3_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_0_3_U117 ( .A(npu_inst_pe_1_0_3_int_q_acc_7_), .B(
        npu_inst_pe_1_0_3_sub_77_carry_7_), .ZN(npu_inst_pe_1_0_3_N72) );
  INV_X1 npu_inst_pe_1_0_3_U116 ( .A(npu_inst_n80), .ZN(npu_inst_pe_1_0_3_n7)
         );
  INV_X1 npu_inst_pe_1_0_3_U115 ( .A(npu_inst_pe_1_0_3_n7), .ZN(
        npu_inst_pe_1_0_3_n6) );
  INV_X1 npu_inst_pe_1_0_3_U114 ( .A(npu_inst_n60), .ZN(npu_inst_pe_1_0_3_n3)
         );
  AOI22_X1 npu_inst_pe_1_0_3_U113 ( .A1(npu_inst_int_data_y_1__3__0_), .A2(
        npu_inst_pe_1_0_3_n58), .B1(npu_inst_pe_1_0_3_n114), .B2(
        npu_inst_pe_1_0_3_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_0_3_n57) );
  INV_X1 npu_inst_pe_1_0_3_U112 ( .A(npu_inst_pe_1_0_3_n57), .ZN(
        npu_inst_pe_1_0_3_n108) );
  AOI22_X1 npu_inst_pe_1_0_3_U111 ( .A1(npu_inst_int_data_y_1__3__0_), .A2(
        npu_inst_pe_1_0_3_n54), .B1(npu_inst_pe_1_0_3_n115), .B2(
        npu_inst_pe_1_0_3_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_0_3_n53) );
  INV_X1 npu_inst_pe_1_0_3_U110 ( .A(npu_inst_pe_1_0_3_n53), .ZN(
        npu_inst_pe_1_0_3_n109) );
  AOI22_X1 npu_inst_pe_1_0_3_U107 ( .A1(npu_inst_int_data_y_1__3__0_), .A2(
        npu_inst_pe_1_0_3_n50), .B1(npu_inst_pe_1_0_3_n116), .B2(
        npu_inst_pe_1_0_3_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_0_3_n49) );
  INV_X1 npu_inst_pe_1_0_3_U106 ( .A(npu_inst_pe_1_0_3_n49), .ZN(
        npu_inst_pe_1_0_3_n110) );
  AOI22_X1 npu_inst_pe_1_0_3_U105 ( .A1(npu_inst_int_data_y_1__3__0_), .A2(
        npu_inst_pe_1_0_3_n46), .B1(npu_inst_pe_1_0_3_n117), .B2(
        npu_inst_pe_1_0_3_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_0_3_n45) );
  INV_X1 npu_inst_pe_1_0_3_U104 ( .A(npu_inst_pe_1_0_3_n45), .ZN(
        npu_inst_pe_1_0_3_n111) );
  AOI22_X1 npu_inst_pe_1_0_3_U103 ( .A1(npu_inst_int_data_y_1__3__0_), .A2(
        npu_inst_pe_1_0_3_n42), .B1(npu_inst_pe_1_0_3_n119), .B2(
        npu_inst_pe_1_0_3_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_0_3_n41) );
  INV_X1 npu_inst_pe_1_0_3_U102 ( .A(npu_inst_pe_1_0_3_n41), .ZN(
        npu_inst_pe_1_0_3_n112) );
  AOI22_X1 npu_inst_pe_1_0_3_U101 ( .A1(npu_inst_int_data_y_1__3__1_), .A2(
        npu_inst_pe_1_0_3_n58), .B1(npu_inst_pe_1_0_3_n114), .B2(
        npu_inst_pe_1_0_3_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_0_3_n59) );
  INV_X1 npu_inst_pe_1_0_3_U100 ( .A(npu_inst_pe_1_0_3_n59), .ZN(
        npu_inst_pe_1_0_3_n102) );
  AOI22_X1 npu_inst_pe_1_0_3_U99 ( .A1(npu_inst_int_data_y_1__3__1_), .A2(
        npu_inst_pe_1_0_3_n54), .B1(npu_inst_pe_1_0_3_n115), .B2(
        npu_inst_pe_1_0_3_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_0_3_n55) );
  INV_X1 npu_inst_pe_1_0_3_U98 ( .A(npu_inst_pe_1_0_3_n55), .ZN(
        npu_inst_pe_1_0_3_n103) );
  AOI22_X1 npu_inst_pe_1_0_3_U97 ( .A1(npu_inst_int_data_y_1__3__1_), .A2(
        npu_inst_pe_1_0_3_n50), .B1(npu_inst_pe_1_0_3_n116), .B2(
        npu_inst_pe_1_0_3_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_0_3_n51) );
  INV_X1 npu_inst_pe_1_0_3_U96 ( .A(npu_inst_pe_1_0_3_n51), .ZN(
        npu_inst_pe_1_0_3_n104) );
  AOI22_X1 npu_inst_pe_1_0_3_U95 ( .A1(npu_inst_int_data_y_1__3__1_), .A2(
        npu_inst_pe_1_0_3_n46), .B1(npu_inst_pe_1_0_3_n117), .B2(
        npu_inst_pe_1_0_3_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_0_3_n47) );
  INV_X1 npu_inst_pe_1_0_3_U94 ( .A(npu_inst_pe_1_0_3_n47), .ZN(
        npu_inst_pe_1_0_3_n105) );
  AOI22_X1 npu_inst_pe_1_0_3_U93 ( .A1(npu_inst_int_data_y_1__3__1_), .A2(
        npu_inst_pe_1_0_3_n42), .B1(npu_inst_pe_1_0_3_n119), .B2(
        npu_inst_pe_1_0_3_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_0_3_n43) );
  INV_X1 npu_inst_pe_1_0_3_U92 ( .A(npu_inst_pe_1_0_3_n43), .ZN(
        npu_inst_pe_1_0_3_n106) );
  AOI22_X1 npu_inst_pe_1_0_3_U91 ( .A1(npu_inst_pe_1_0_3_n38), .A2(
        npu_inst_int_data_y_1__3__1_), .B1(npu_inst_pe_1_0_3_n118), .B2(
        npu_inst_pe_1_0_3_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_0_3_n39) );
  INV_X1 npu_inst_pe_1_0_3_U90 ( .A(npu_inst_pe_1_0_3_n39), .ZN(
        npu_inst_pe_1_0_3_n107) );
  AOI22_X1 npu_inst_pe_1_0_3_U89 ( .A1(npu_inst_pe_1_0_3_n38), .A2(
        npu_inst_int_data_y_1__3__0_), .B1(npu_inst_pe_1_0_3_n118), .B2(
        npu_inst_pe_1_0_3_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_0_3_n37) );
  INV_X1 npu_inst_pe_1_0_3_U88 ( .A(npu_inst_pe_1_0_3_n37), .ZN(
        npu_inst_pe_1_0_3_n113) );
  AND2_X1 npu_inst_pe_1_0_3_U87 ( .A1(npu_inst_pe_1_0_3_n2), .A2(
        npu_inst_pe_1_0_3_int_q_acc_7_), .ZN(o_data[39]) );
  AND2_X1 npu_inst_pe_1_0_3_U86 ( .A1(npu_inst_pe_1_0_3_int_q_acc_6_), .A2(
        npu_inst_pe_1_0_3_n2), .ZN(o_data[38]) );
  AND2_X1 npu_inst_pe_1_0_3_U85 ( .A1(npu_inst_pe_1_0_3_int_q_acc_5_), .A2(
        npu_inst_pe_1_0_3_n2), .ZN(o_data[37]) );
  AND2_X1 npu_inst_pe_1_0_3_U84 ( .A1(npu_inst_pe_1_0_3_int_q_acc_4_), .A2(
        npu_inst_pe_1_0_3_n2), .ZN(o_data[36]) );
  AND2_X1 npu_inst_pe_1_0_3_U83 ( .A1(npu_inst_pe_1_0_3_int_q_acc_3_), .A2(
        npu_inst_pe_1_0_3_n2), .ZN(o_data[35]) );
  NAND2_X1 npu_inst_pe_1_0_3_U82 ( .A1(npu_inst_pe_1_0_3_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_0_3_n60), .ZN(npu_inst_pe_1_0_3_n74) );
  OAI21_X1 npu_inst_pe_1_0_3_U81 ( .B1(npu_inst_pe_1_0_3_n63), .B2(
        npu_inst_pe_1_0_3_n60), .A(npu_inst_pe_1_0_3_n74), .ZN(
        npu_inst_pe_1_0_3_n97) );
  NAND2_X1 npu_inst_pe_1_0_3_U80 ( .A1(npu_inst_pe_1_0_3_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_0_3_n60), .ZN(npu_inst_pe_1_0_3_n73) );
  OAI21_X1 npu_inst_pe_1_0_3_U79 ( .B1(npu_inst_pe_1_0_3_n61), .B2(
        npu_inst_pe_1_0_3_n60), .A(npu_inst_pe_1_0_3_n73), .ZN(
        npu_inst_pe_1_0_3_n96) );
  NAND2_X1 npu_inst_pe_1_0_3_U78 ( .A1(npu_inst_pe_1_0_3_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_0_3_n56), .ZN(npu_inst_pe_1_0_3_n72) );
  OAI21_X1 npu_inst_pe_1_0_3_U77 ( .B1(npu_inst_pe_1_0_3_n63), .B2(
        npu_inst_pe_1_0_3_n56), .A(npu_inst_pe_1_0_3_n72), .ZN(
        npu_inst_pe_1_0_3_n95) );
  NAND2_X1 npu_inst_pe_1_0_3_U76 ( .A1(npu_inst_pe_1_0_3_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_0_3_n56), .ZN(npu_inst_pe_1_0_3_n71) );
  OAI21_X1 npu_inst_pe_1_0_3_U75 ( .B1(npu_inst_pe_1_0_3_n61), .B2(
        npu_inst_pe_1_0_3_n56), .A(npu_inst_pe_1_0_3_n71), .ZN(
        npu_inst_pe_1_0_3_n94) );
  NAND2_X1 npu_inst_pe_1_0_3_U74 ( .A1(npu_inst_pe_1_0_3_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_0_3_n52), .ZN(npu_inst_pe_1_0_3_n70) );
  OAI21_X1 npu_inst_pe_1_0_3_U73 ( .B1(npu_inst_pe_1_0_3_n63), .B2(
        npu_inst_pe_1_0_3_n52), .A(npu_inst_pe_1_0_3_n70), .ZN(
        npu_inst_pe_1_0_3_n93) );
  NAND2_X1 npu_inst_pe_1_0_3_U72 ( .A1(npu_inst_pe_1_0_3_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_0_3_n52), .ZN(npu_inst_pe_1_0_3_n69) );
  OAI21_X1 npu_inst_pe_1_0_3_U71 ( .B1(npu_inst_pe_1_0_3_n61), .B2(
        npu_inst_pe_1_0_3_n52), .A(npu_inst_pe_1_0_3_n69), .ZN(
        npu_inst_pe_1_0_3_n92) );
  NAND2_X1 npu_inst_pe_1_0_3_U70 ( .A1(npu_inst_pe_1_0_3_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_0_3_n48), .ZN(npu_inst_pe_1_0_3_n68) );
  OAI21_X1 npu_inst_pe_1_0_3_U69 ( .B1(npu_inst_pe_1_0_3_n63), .B2(
        npu_inst_pe_1_0_3_n48), .A(npu_inst_pe_1_0_3_n68), .ZN(
        npu_inst_pe_1_0_3_n91) );
  NAND2_X1 npu_inst_pe_1_0_3_U68 ( .A1(npu_inst_pe_1_0_3_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_0_3_n48), .ZN(npu_inst_pe_1_0_3_n67) );
  OAI21_X1 npu_inst_pe_1_0_3_U67 ( .B1(npu_inst_pe_1_0_3_n61), .B2(
        npu_inst_pe_1_0_3_n48), .A(npu_inst_pe_1_0_3_n67), .ZN(
        npu_inst_pe_1_0_3_n90) );
  NAND2_X1 npu_inst_pe_1_0_3_U66 ( .A1(npu_inst_pe_1_0_3_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_0_3_n44), .ZN(npu_inst_pe_1_0_3_n66) );
  OAI21_X1 npu_inst_pe_1_0_3_U65 ( .B1(npu_inst_pe_1_0_3_n63), .B2(
        npu_inst_pe_1_0_3_n44), .A(npu_inst_pe_1_0_3_n66), .ZN(
        npu_inst_pe_1_0_3_n89) );
  NAND2_X1 npu_inst_pe_1_0_3_U64 ( .A1(npu_inst_pe_1_0_3_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_0_3_n44), .ZN(npu_inst_pe_1_0_3_n65) );
  OAI21_X1 npu_inst_pe_1_0_3_U63 ( .B1(npu_inst_pe_1_0_3_n61), .B2(
        npu_inst_pe_1_0_3_n44), .A(npu_inst_pe_1_0_3_n65), .ZN(
        npu_inst_pe_1_0_3_n88) );
  NAND2_X1 npu_inst_pe_1_0_3_U62 ( .A1(npu_inst_pe_1_0_3_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_0_3_n40), .ZN(npu_inst_pe_1_0_3_n64) );
  OAI21_X1 npu_inst_pe_1_0_3_U61 ( .B1(npu_inst_pe_1_0_3_n63), .B2(
        npu_inst_pe_1_0_3_n40), .A(npu_inst_pe_1_0_3_n64), .ZN(
        npu_inst_pe_1_0_3_n87) );
  NAND2_X1 npu_inst_pe_1_0_3_U60 ( .A1(npu_inst_pe_1_0_3_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_0_3_n40), .ZN(npu_inst_pe_1_0_3_n62) );
  OAI21_X1 npu_inst_pe_1_0_3_U59 ( .B1(npu_inst_pe_1_0_3_n61), .B2(
        npu_inst_pe_1_0_3_n40), .A(npu_inst_pe_1_0_3_n62), .ZN(
        npu_inst_pe_1_0_3_n86) );
  NOR3_X1 npu_inst_pe_1_0_3_U58 ( .A1(npu_inst_pe_1_0_3_n26), .A2(npu_inst_n60), .A3(npu_inst_int_ckg[60]), .ZN(npu_inst_pe_1_0_3_n85) );
  OR2_X1 npu_inst_pe_1_0_3_U57 ( .A1(npu_inst_pe_1_0_3_n85), .A2(
        npu_inst_pe_1_0_3_n2), .ZN(npu_inst_pe_1_0_3_N84) );
  AND2_X1 npu_inst_pe_1_0_3_U56 ( .A1(npu_inst_pe_1_0_3_int_q_acc_0_), .A2(
        npu_inst_pe_1_0_3_n1), .ZN(o_data[32]) );
  AND2_X1 npu_inst_pe_1_0_3_U55 ( .A1(npu_inst_pe_1_0_3_int_q_acc_1_), .A2(
        npu_inst_pe_1_0_3_n1), .ZN(o_data[33]) );
  AND2_X1 npu_inst_pe_1_0_3_U54 ( .A1(npu_inst_pe_1_0_3_int_q_acc_2_), .A2(
        npu_inst_pe_1_0_3_n1), .ZN(o_data[34]) );
  AOI222_X1 npu_inst_pe_1_0_3_U53 ( .A1(npu_inst_int_data_res_1__3__0_), .A2(
        npu_inst_pe_1_0_3_n1), .B1(npu_inst_pe_1_0_3_N73), .B2(
        npu_inst_pe_1_0_3_n76), .C1(npu_inst_pe_1_0_3_N65), .C2(
        npu_inst_pe_1_0_3_n77), .ZN(npu_inst_pe_1_0_3_n84) );
  INV_X1 npu_inst_pe_1_0_3_U52 ( .A(npu_inst_pe_1_0_3_n84), .ZN(
        npu_inst_pe_1_0_3_n101) );
  AOI222_X1 npu_inst_pe_1_0_3_U51 ( .A1(npu_inst_int_data_res_1__3__7_), .A2(
        npu_inst_pe_1_0_3_n1), .B1(npu_inst_pe_1_0_3_N80), .B2(
        npu_inst_pe_1_0_3_n76), .C1(npu_inst_pe_1_0_3_N72), .C2(
        npu_inst_pe_1_0_3_n77), .ZN(npu_inst_pe_1_0_3_n75) );
  INV_X1 npu_inst_pe_1_0_3_U50 ( .A(npu_inst_pe_1_0_3_n75), .ZN(
        npu_inst_pe_1_0_3_n33) );
  AOI222_X1 npu_inst_pe_1_0_3_U49 ( .A1(npu_inst_int_data_res_1__3__1_), .A2(
        npu_inst_pe_1_0_3_n1), .B1(npu_inst_pe_1_0_3_N74), .B2(
        npu_inst_pe_1_0_3_n76), .C1(npu_inst_pe_1_0_3_N66), .C2(
        npu_inst_pe_1_0_3_n77), .ZN(npu_inst_pe_1_0_3_n83) );
  INV_X1 npu_inst_pe_1_0_3_U48 ( .A(npu_inst_pe_1_0_3_n83), .ZN(
        npu_inst_pe_1_0_3_n100) );
  AOI222_X1 npu_inst_pe_1_0_3_U47 ( .A1(npu_inst_int_data_res_1__3__2_), .A2(
        npu_inst_pe_1_0_3_n1), .B1(npu_inst_pe_1_0_3_N75), .B2(
        npu_inst_pe_1_0_3_n76), .C1(npu_inst_pe_1_0_3_N67), .C2(
        npu_inst_pe_1_0_3_n77), .ZN(npu_inst_pe_1_0_3_n82) );
  INV_X1 npu_inst_pe_1_0_3_U46 ( .A(npu_inst_pe_1_0_3_n82), .ZN(
        npu_inst_pe_1_0_3_n99) );
  AOI222_X1 npu_inst_pe_1_0_3_U45 ( .A1(npu_inst_int_data_res_1__3__3_), .A2(
        npu_inst_pe_1_0_3_n1), .B1(npu_inst_pe_1_0_3_N76), .B2(
        npu_inst_pe_1_0_3_n76), .C1(npu_inst_pe_1_0_3_N68), .C2(
        npu_inst_pe_1_0_3_n77), .ZN(npu_inst_pe_1_0_3_n81) );
  INV_X1 npu_inst_pe_1_0_3_U44 ( .A(npu_inst_pe_1_0_3_n81), .ZN(
        npu_inst_pe_1_0_3_n98) );
  AOI222_X1 npu_inst_pe_1_0_3_U43 ( .A1(npu_inst_int_data_res_1__3__4_), .A2(
        npu_inst_pe_1_0_3_n1), .B1(npu_inst_pe_1_0_3_N77), .B2(
        npu_inst_pe_1_0_3_n76), .C1(npu_inst_pe_1_0_3_N69), .C2(
        npu_inst_pe_1_0_3_n77), .ZN(npu_inst_pe_1_0_3_n80) );
  INV_X1 npu_inst_pe_1_0_3_U42 ( .A(npu_inst_pe_1_0_3_n80), .ZN(
        npu_inst_pe_1_0_3_n36) );
  AOI222_X1 npu_inst_pe_1_0_3_U41 ( .A1(npu_inst_int_data_res_1__3__5_), .A2(
        npu_inst_pe_1_0_3_n1), .B1(npu_inst_pe_1_0_3_N78), .B2(
        npu_inst_pe_1_0_3_n76), .C1(npu_inst_pe_1_0_3_N70), .C2(
        npu_inst_pe_1_0_3_n77), .ZN(npu_inst_pe_1_0_3_n79) );
  INV_X1 npu_inst_pe_1_0_3_U40 ( .A(npu_inst_pe_1_0_3_n79), .ZN(
        npu_inst_pe_1_0_3_n35) );
  AOI222_X1 npu_inst_pe_1_0_3_U39 ( .A1(npu_inst_int_data_res_1__3__6_), .A2(
        npu_inst_pe_1_0_3_n1), .B1(npu_inst_pe_1_0_3_N79), .B2(
        npu_inst_pe_1_0_3_n76), .C1(npu_inst_pe_1_0_3_N71), .C2(
        npu_inst_pe_1_0_3_n77), .ZN(npu_inst_pe_1_0_3_n78) );
  INV_X1 npu_inst_pe_1_0_3_U38 ( .A(npu_inst_pe_1_0_3_n78), .ZN(
        npu_inst_pe_1_0_3_n34) );
  INV_X1 npu_inst_pe_1_0_3_U37 ( .A(npu_inst_pe_1_0_3_int_data_1_), .ZN(
        npu_inst_pe_1_0_3_n14) );
  AND2_X1 npu_inst_pe_1_0_3_U36 ( .A1(npu_inst_int_data_x_0__3__1_), .A2(
        npu_inst_pe_1_0_3_int_q_weight_1_), .ZN(npu_inst_pe_1_0_3_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_0_3_U35 ( .A1(npu_inst_int_data_x_0__3__0_), .A2(
        npu_inst_pe_1_0_3_int_q_weight_1_), .ZN(npu_inst_pe_1_0_3_int_data_0_)
         );
  AND2_X1 npu_inst_pe_1_0_3_U34 ( .A1(npu_inst_pe_1_0_3_N93), .A2(npu_inst_n60), .ZN(npu_inst_pe_1_0_3_o_data_v_0_) );
  AND2_X1 npu_inst_pe_1_0_3_U33 ( .A1(npu_inst_n60), .A2(npu_inst_pe_1_0_3_N94), .ZN(npu_inst_pe_1_0_3_o_data_v_1_) );
  AOI22_X1 npu_inst_pe_1_0_3_U32 ( .A1(npu_inst_n60), .A2(
        npu_inst_int_data_y_1__3__1_), .B1(npu_inst_pe_1_0_3_n3), .B2(
        npu_inst_int_data_x_0__4__1_), .ZN(npu_inst_pe_1_0_3_n63) );
  AOI22_X1 npu_inst_pe_1_0_3_U31 ( .A1(npu_inst_n60), .A2(
        npu_inst_int_data_y_1__3__0_), .B1(npu_inst_pe_1_0_3_n3), .B2(
        npu_inst_int_data_x_0__4__0_), .ZN(npu_inst_pe_1_0_3_n61) );
  INV_X1 npu_inst_pe_1_0_3_U30 ( .A(npu_inst_pe_1_0_3_int_data_0_), .ZN(
        npu_inst_pe_1_0_3_n13) );
  INV_X1 npu_inst_pe_1_0_3_U29 ( .A(npu_inst_n72), .ZN(npu_inst_pe_1_0_3_n5)
         );
  OR3_X1 npu_inst_pe_1_0_3_U28 ( .A1(npu_inst_pe_1_0_3_n6), .A2(
        npu_inst_pe_1_0_3_n8), .A3(npu_inst_pe_1_0_3_n5), .ZN(
        npu_inst_pe_1_0_3_n56) );
  OR3_X1 npu_inst_pe_1_0_3_U27 ( .A1(npu_inst_pe_1_0_3_n5), .A2(
        npu_inst_pe_1_0_3_n8), .A3(npu_inst_pe_1_0_3_n7), .ZN(
        npu_inst_pe_1_0_3_n48) );
  INV_X1 npu_inst_pe_1_0_3_U26 ( .A(npu_inst_pe_1_0_3_n5), .ZN(
        npu_inst_pe_1_0_3_n4) );
  INV_X1 npu_inst_pe_1_0_3_U25 ( .A(npu_inst_n127), .ZN(npu_inst_pe_1_0_3_n12)
         );
  OR3_X1 npu_inst_pe_1_0_3_U24 ( .A1(npu_inst_pe_1_0_3_n4), .A2(
        npu_inst_pe_1_0_3_n8), .A3(npu_inst_pe_1_0_3_n7), .ZN(
        npu_inst_pe_1_0_3_n52) );
  OR3_X1 npu_inst_pe_1_0_3_U23 ( .A1(npu_inst_pe_1_0_3_n6), .A2(
        npu_inst_pe_1_0_3_n8), .A3(npu_inst_pe_1_0_3_n4), .ZN(
        npu_inst_pe_1_0_3_n60) );
  NOR2_X1 npu_inst_pe_1_0_3_U22 ( .A1(npu_inst_pe_1_0_3_n60), .A2(
        npu_inst_pe_1_0_3_n3), .ZN(npu_inst_pe_1_0_3_n58) );
  NOR2_X1 npu_inst_pe_1_0_3_U21 ( .A1(npu_inst_pe_1_0_3_n56), .A2(
        npu_inst_pe_1_0_3_n3), .ZN(npu_inst_pe_1_0_3_n54) );
  NOR2_X1 npu_inst_pe_1_0_3_U20 ( .A1(npu_inst_pe_1_0_3_n52), .A2(
        npu_inst_pe_1_0_3_n3), .ZN(npu_inst_pe_1_0_3_n50) );
  NOR2_X1 npu_inst_pe_1_0_3_U19 ( .A1(npu_inst_pe_1_0_3_n48), .A2(
        npu_inst_pe_1_0_3_n3), .ZN(npu_inst_pe_1_0_3_n46) );
  NOR2_X1 npu_inst_pe_1_0_3_U18 ( .A1(npu_inst_pe_1_0_3_n40), .A2(
        npu_inst_pe_1_0_3_n3), .ZN(npu_inst_pe_1_0_3_n38) );
  NOR2_X1 npu_inst_pe_1_0_3_U17 ( .A1(npu_inst_pe_1_0_3_n44), .A2(
        npu_inst_pe_1_0_3_n3), .ZN(npu_inst_pe_1_0_3_n42) );
  BUF_X1 npu_inst_pe_1_0_3_U16 ( .A(npu_inst_n107), .Z(npu_inst_pe_1_0_3_n8)
         );
  BUF_X1 npu_inst_pe_1_0_3_U15 ( .A(npu_inst_pe_1_0_3_n12), .Z(
        npu_inst_pe_1_0_3_n11) );
  BUF_X1 npu_inst_pe_1_0_3_U14 ( .A(npu_inst_pe_1_0_3_n12), .Z(
        npu_inst_pe_1_0_3_n10) );
  BUF_X1 npu_inst_pe_1_0_3_U13 ( .A(npu_inst_pe_1_0_3_n12), .Z(
        npu_inst_pe_1_0_3_n9) );
  INV_X1 npu_inst_pe_1_0_3_U12 ( .A(npu_inst_pe_1_0_3_n38), .ZN(
        npu_inst_pe_1_0_3_n118) );
  INV_X1 npu_inst_pe_1_0_3_U11 ( .A(npu_inst_pe_1_0_3_n58), .ZN(
        npu_inst_pe_1_0_3_n114) );
  INV_X1 npu_inst_pe_1_0_3_U10 ( .A(npu_inst_pe_1_0_3_n54), .ZN(
        npu_inst_pe_1_0_3_n115) );
  INV_X1 npu_inst_pe_1_0_3_U9 ( .A(npu_inst_pe_1_0_3_n50), .ZN(
        npu_inst_pe_1_0_3_n116) );
  INV_X1 npu_inst_pe_1_0_3_U8 ( .A(npu_inst_pe_1_0_3_n46), .ZN(
        npu_inst_pe_1_0_3_n117) );
  INV_X1 npu_inst_pe_1_0_3_U7 ( .A(npu_inst_pe_1_0_3_n42), .ZN(
        npu_inst_pe_1_0_3_n119) );
  BUF_X1 npu_inst_pe_1_0_3_U6 ( .A(npu_inst_n37), .Z(npu_inst_pe_1_0_3_n2) );
  BUF_X1 npu_inst_pe_1_0_3_U5 ( .A(npu_inst_n37), .Z(npu_inst_pe_1_0_3_n1) );
  NOR2_X1 npu_inst_pe_1_0_3_U4 ( .A1(npu_inst_pe_1_0_3_int_q_weight_0_), .A2(
        npu_inst_pe_1_0_3_n1), .ZN(npu_inst_pe_1_0_3_n76) );
  NOR2_X1 npu_inst_pe_1_0_3_U3 ( .A1(npu_inst_pe_1_0_3_n27), .A2(
        npu_inst_pe_1_0_3_n1), .ZN(npu_inst_pe_1_0_3_n77) );
  FA_X1 npu_inst_pe_1_0_3_sub_77_U2_1 ( .A(npu_inst_pe_1_0_3_int_q_acc_1_), 
        .B(npu_inst_pe_1_0_3_n14), .CI(npu_inst_pe_1_0_3_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_0_3_sub_77_carry_2_), .S(npu_inst_pe_1_0_3_N66) );
  FA_X1 npu_inst_pe_1_0_3_add_79_U1_1 ( .A(npu_inst_pe_1_0_3_int_q_acc_1_), 
        .B(npu_inst_pe_1_0_3_int_data_1_), .CI(
        npu_inst_pe_1_0_3_add_79_carry_1_), .CO(
        npu_inst_pe_1_0_3_add_79_carry_2_), .S(npu_inst_pe_1_0_3_N74) );
  NAND3_X1 npu_inst_pe_1_0_3_U109 ( .A1(npu_inst_pe_1_0_3_n5), .A2(
        npu_inst_pe_1_0_3_n7), .A3(npu_inst_pe_1_0_3_n8), .ZN(
        npu_inst_pe_1_0_3_n44) );
  NAND3_X1 npu_inst_pe_1_0_3_U108 ( .A1(npu_inst_pe_1_0_3_n4), .A2(
        npu_inst_pe_1_0_3_n7), .A3(npu_inst_pe_1_0_3_n8), .ZN(
        npu_inst_pe_1_0_3_n40) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_0_3_n34), .CK(
        npu_inst_pe_1_0_3_net4224), .RN(npu_inst_pe_1_0_3_n9), .Q(
        npu_inst_pe_1_0_3_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_0_3_n35), .CK(
        npu_inst_pe_1_0_3_net4224), .RN(npu_inst_pe_1_0_3_n9), .Q(
        npu_inst_pe_1_0_3_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_0_3_n36), .CK(
        npu_inst_pe_1_0_3_net4224), .RN(npu_inst_pe_1_0_3_n9), .Q(
        npu_inst_pe_1_0_3_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_0_3_n98), .CK(
        npu_inst_pe_1_0_3_net4224), .RN(npu_inst_pe_1_0_3_n9), .Q(
        npu_inst_pe_1_0_3_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_0_3_n99), .CK(
        npu_inst_pe_1_0_3_net4224), .RN(npu_inst_pe_1_0_3_n9), .Q(
        npu_inst_pe_1_0_3_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_0_3_n100), 
        .CK(npu_inst_pe_1_0_3_net4224), .RN(npu_inst_pe_1_0_3_n9), .Q(
        npu_inst_pe_1_0_3_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_0_3_n33), .CK(
        npu_inst_pe_1_0_3_net4224), .RN(npu_inst_pe_1_0_3_n9), .Q(
        npu_inst_pe_1_0_3_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_0_3_n101), 
        .CK(npu_inst_pe_1_0_3_net4224), .RN(npu_inst_pe_1_0_3_n9), .Q(
        npu_inst_pe_1_0_3_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_weight_reg_0_ ( .D(npu_inst_n113), .CK(
        npu_inst_pe_1_0_3_net4230), .RN(npu_inst_pe_1_0_3_n9), .Q(
        npu_inst_pe_1_0_3_int_q_weight_0_), .QN(npu_inst_pe_1_0_3_n27) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_weight_reg_1_ ( .D(npu_inst_n119), .CK(
        npu_inst_pe_1_0_3_net4230), .RN(npu_inst_pe_1_0_3_n9), .Q(
        npu_inst_pe_1_0_3_int_q_weight_1_), .QN(npu_inst_pe_1_0_3_n26) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_0_3_n113), 
        .CK(npu_inst_pe_1_0_3_net4230), .RN(npu_inst_pe_1_0_3_n9), .Q(
        npu_inst_pe_1_0_3_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_0_3_n107), 
        .CK(npu_inst_pe_1_0_3_net4230), .RN(npu_inst_pe_1_0_3_n9), .Q(
        npu_inst_pe_1_0_3_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_0_3_n112), 
        .CK(npu_inst_pe_1_0_3_net4230), .RN(npu_inst_pe_1_0_3_n10), .Q(
        npu_inst_pe_1_0_3_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_0_3_n106), 
        .CK(npu_inst_pe_1_0_3_net4230), .RN(npu_inst_pe_1_0_3_n10), .Q(
        npu_inst_pe_1_0_3_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_0_3_n111), 
        .CK(npu_inst_pe_1_0_3_net4230), .RN(npu_inst_pe_1_0_3_n10), .Q(
        npu_inst_pe_1_0_3_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_0_3_n105), 
        .CK(npu_inst_pe_1_0_3_net4230), .RN(npu_inst_pe_1_0_3_n10), .Q(
        npu_inst_pe_1_0_3_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_0_3_n110), 
        .CK(npu_inst_pe_1_0_3_net4230), .RN(npu_inst_pe_1_0_3_n10), .Q(
        npu_inst_pe_1_0_3_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_0_3_n104), 
        .CK(npu_inst_pe_1_0_3_net4230), .RN(npu_inst_pe_1_0_3_n10), .Q(
        npu_inst_pe_1_0_3_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_0_3_n109), 
        .CK(npu_inst_pe_1_0_3_net4230), .RN(npu_inst_pe_1_0_3_n10), .Q(
        npu_inst_pe_1_0_3_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_0_3_n103), 
        .CK(npu_inst_pe_1_0_3_net4230), .RN(npu_inst_pe_1_0_3_n10), .Q(
        npu_inst_pe_1_0_3_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_0_3_n108), 
        .CK(npu_inst_pe_1_0_3_net4230), .RN(npu_inst_pe_1_0_3_n10), .Q(
        npu_inst_pe_1_0_3_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_0_3_n102), 
        .CK(npu_inst_pe_1_0_3_net4230), .RN(npu_inst_pe_1_0_3_n10), .Q(
        npu_inst_pe_1_0_3_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_0_3_n86), 
        .CK(npu_inst_pe_1_0_3_net4230), .RN(npu_inst_pe_1_0_3_n10), .Q(
        npu_inst_pe_1_0_3_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_0_3_n87), 
        .CK(npu_inst_pe_1_0_3_net4230), .RN(npu_inst_pe_1_0_3_n10), .Q(
        npu_inst_pe_1_0_3_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_0_3_n88), 
        .CK(npu_inst_pe_1_0_3_net4230), .RN(npu_inst_pe_1_0_3_n11), .Q(
        npu_inst_pe_1_0_3_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_0_3_n89), 
        .CK(npu_inst_pe_1_0_3_net4230), .RN(npu_inst_pe_1_0_3_n11), .Q(
        npu_inst_pe_1_0_3_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_0_3_n90), 
        .CK(npu_inst_pe_1_0_3_net4230), .RN(npu_inst_pe_1_0_3_n11), .Q(
        npu_inst_pe_1_0_3_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_0_3_n91), 
        .CK(npu_inst_pe_1_0_3_net4230), .RN(npu_inst_pe_1_0_3_n11), .Q(
        npu_inst_pe_1_0_3_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_0_3_n92), 
        .CK(npu_inst_pe_1_0_3_net4230), .RN(npu_inst_pe_1_0_3_n11), .Q(
        npu_inst_pe_1_0_3_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_0_3_n93), 
        .CK(npu_inst_pe_1_0_3_net4230), .RN(npu_inst_pe_1_0_3_n11), .Q(
        npu_inst_pe_1_0_3_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_0_3_n94), 
        .CK(npu_inst_pe_1_0_3_net4230), .RN(npu_inst_pe_1_0_3_n11), .Q(
        npu_inst_pe_1_0_3_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_0_3_n95), 
        .CK(npu_inst_pe_1_0_3_net4230), .RN(npu_inst_pe_1_0_3_n11), .Q(
        npu_inst_pe_1_0_3_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_0_3_n96), 
        .CK(npu_inst_pe_1_0_3_net4230), .RN(npu_inst_pe_1_0_3_n11), .Q(
        npu_inst_pe_1_0_3_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_0_3_n97), 
        .CK(npu_inst_pe_1_0_3_net4230), .RN(npu_inst_pe_1_0_3_n11), .Q(
        npu_inst_pe_1_0_3_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_0_3_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_0_3_N84), .SE(1'b0), .GCK(npu_inst_pe_1_0_3_net4224) );
  CLKGATETST_X1 npu_inst_pe_1_0_3_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n66), .SE(1'b0), .GCK(npu_inst_pe_1_0_3_net4230) );
  MUX2_X1 npu_inst_pe_1_0_4_U161 ( .A(npu_inst_pe_1_0_4_n31), .B(
        npu_inst_pe_1_0_4_n28), .S(npu_inst_pe_1_0_4_n7), .Z(
        npu_inst_pe_1_0_4_N93) );
  MUX2_X1 npu_inst_pe_1_0_4_U160 ( .A(npu_inst_pe_1_0_4_n30), .B(
        npu_inst_pe_1_0_4_n29), .S(npu_inst_n79), .Z(npu_inst_pe_1_0_4_n31) );
  MUX2_X1 npu_inst_pe_1_0_4_U159 ( .A(npu_inst_pe_1_0_4_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_0_4_int_q_reg_v_1__0_), .S(npu_inst_pe_1_0_4_n4), .Z(
        npu_inst_pe_1_0_4_n30) );
  MUX2_X1 npu_inst_pe_1_0_4_U158 ( .A(npu_inst_pe_1_0_4_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_0_4_int_q_reg_v_3__0_), .S(npu_inst_pe_1_0_4_n4), .Z(
        npu_inst_pe_1_0_4_n29) );
  MUX2_X1 npu_inst_pe_1_0_4_U157 ( .A(npu_inst_pe_1_0_4_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_0_4_int_q_reg_v_5__0_), .S(npu_inst_pe_1_0_4_n4), .Z(
        npu_inst_pe_1_0_4_n28) );
  MUX2_X1 npu_inst_pe_1_0_4_U156 ( .A(npu_inst_pe_1_0_4_n25), .B(
        npu_inst_pe_1_0_4_n22), .S(npu_inst_pe_1_0_4_n7), .Z(
        npu_inst_pe_1_0_4_N94) );
  MUX2_X1 npu_inst_pe_1_0_4_U155 ( .A(npu_inst_pe_1_0_4_n24), .B(
        npu_inst_pe_1_0_4_n23), .S(npu_inst_n79), .Z(npu_inst_pe_1_0_4_n25) );
  MUX2_X1 npu_inst_pe_1_0_4_U154 ( .A(npu_inst_pe_1_0_4_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_0_4_int_q_reg_v_1__1_), .S(npu_inst_pe_1_0_4_n4), .Z(
        npu_inst_pe_1_0_4_n24) );
  MUX2_X1 npu_inst_pe_1_0_4_U153 ( .A(npu_inst_pe_1_0_4_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_0_4_int_q_reg_v_3__1_), .S(npu_inst_pe_1_0_4_n4), .Z(
        npu_inst_pe_1_0_4_n23) );
  MUX2_X1 npu_inst_pe_1_0_4_U152 ( .A(npu_inst_pe_1_0_4_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_0_4_int_q_reg_v_5__1_), .S(npu_inst_pe_1_0_4_n4), .Z(
        npu_inst_pe_1_0_4_n22) );
  MUX2_X1 npu_inst_pe_1_0_4_U151 ( .A(npu_inst_pe_1_0_4_n21), .B(
        npu_inst_pe_1_0_4_n18), .S(npu_inst_pe_1_0_4_n7), .Z(
        npu_inst_int_data_x_0__4__1_) );
  MUX2_X1 npu_inst_pe_1_0_4_U150 ( .A(npu_inst_pe_1_0_4_n20), .B(
        npu_inst_pe_1_0_4_n19), .S(npu_inst_n79), .Z(npu_inst_pe_1_0_4_n21) );
  MUX2_X1 npu_inst_pe_1_0_4_U149 ( .A(npu_inst_pe_1_0_4_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_0_4_int_q_reg_h_1__1_), .S(npu_inst_pe_1_0_4_n4), .Z(
        npu_inst_pe_1_0_4_n20) );
  MUX2_X1 npu_inst_pe_1_0_4_U148 ( .A(npu_inst_pe_1_0_4_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_0_4_int_q_reg_h_3__1_), .S(npu_inst_pe_1_0_4_n4), .Z(
        npu_inst_pe_1_0_4_n19) );
  MUX2_X1 npu_inst_pe_1_0_4_U147 ( .A(npu_inst_pe_1_0_4_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_0_4_int_q_reg_h_5__1_), .S(npu_inst_pe_1_0_4_n4), .Z(
        npu_inst_pe_1_0_4_n18) );
  MUX2_X1 npu_inst_pe_1_0_4_U146 ( .A(npu_inst_pe_1_0_4_n17), .B(
        npu_inst_pe_1_0_4_n14), .S(npu_inst_pe_1_0_4_n7), .Z(
        npu_inst_int_data_x_0__4__0_) );
  MUX2_X1 npu_inst_pe_1_0_4_U145 ( .A(npu_inst_pe_1_0_4_n16), .B(
        npu_inst_pe_1_0_4_n15), .S(npu_inst_n79), .Z(npu_inst_pe_1_0_4_n17) );
  MUX2_X1 npu_inst_pe_1_0_4_U144 ( .A(npu_inst_pe_1_0_4_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_0_4_int_q_reg_h_1__0_), .S(npu_inst_pe_1_0_4_n4), .Z(
        npu_inst_pe_1_0_4_n16) );
  MUX2_X1 npu_inst_pe_1_0_4_U143 ( .A(npu_inst_pe_1_0_4_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_0_4_int_q_reg_h_3__0_), .S(npu_inst_pe_1_0_4_n4), .Z(
        npu_inst_pe_1_0_4_n15) );
  MUX2_X1 npu_inst_pe_1_0_4_U142 ( .A(npu_inst_pe_1_0_4_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_0_4_int_q_reg_h_5__0_), .S(npu_inst_pe_1_0_4_n4), .Z(
        npu_inst_pe_1_0_4_n14) );
  XOR2_X1 npu_inst_pe_1_0_4_U141 ( .A(npu_inst_pe_1_0_4_int_data_0_), .B(
        npu_inst_pe_1_0_4_int_q_acc_0_), .Z(npu_inst_pe_1_0_4_N73) );
  AND2_X1 npu_inst_pe_1_0_4_U140 ( .A1(npu_inst_pe_1_0_4_int_q_acc_0_), .A2(
        npu_inst_pe_1_0_4_int_data_0_), .ZN(npu_inst_pe_1_0_4_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_0_4_U139 ( .A(npu_inst_pe_1_0_4_int_q_acc_0_), .B(
        npu_inst_pe_1_0_4_n12), .ZN(npu_inst_pe_1_0_4_N65) );
  OR2_X1 npu_inst_pe_1_0_4_U138 ( .A1(npu_inst_pe_1_0_4_n12), .A2(
        npu_inst_pe_1_0_4_int_q_acc_0_), .ZN(npu_inst_pe_1_0_4_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_0_4_U137 ( .A(npu_inst_pe_1_0_4_int_q_acc_2_), .B(
        npu_inst_pe_1_0_4_add_79_carry_2_), .Z(npu_inst_pe_1_0_4_N75) );
  AND2_X1 npu_inst_pe_1_0_4_U136 ( .A1(npu_inst_pe_1_0_4_add_79_carry_2_), 
        .A2(npu_inst_pe_1_0_4_int_q_acc_2_), .ZN(
        npu_inst_pe_1_0_4_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_0_4_U135 ( .A(npu_inst_pe_1_0_4_int_q_acc_3_), .B(
        npu_inst_pe_1_0_4_add_79_carry_3_), .Z(npu_inst_pe_1_0_4_N76) );
  AND2_X1 npu_inst_pe_1_0_4_U134 ( .A1(npu_inst_pe_1_0_4_add_79_carry_3_), 
        .A2(npu_inst_pe_1_0_4_int_q_acc_3_), .ZN(
        npu_inst_pe_1_0_4_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_0_4_U133 ( .A(npu_inst_pe_1_0_4_int_q_acc_4_), .B(
        npu_inst_pe_1_0_4_add_79_carry_4_), .Z(npu_inst_pe_1_0_4_N77) );
  AND2_X1 npu_inst_pe_1_0_4_U132 ( .A1(npu_inst_pe_1_0_4_add_79_carry_4_), 
        .A2(npu_inst_pe_1_0_4_int_q_acc_4_), .ZN(
        npu_inst_pe_1_0_4_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_0_4_U131 ( .A(npu_inst_pe_1_0_4_int_q_acc_5_), .B(
        npu_inst_pe_1_0_4_add_79_carry_5_), .Z(npu_inst_pe_1_0_4_N78) );
  AND2_X1 npu_inst_pe_1_0_4_U130 ( .A1(npu_inst_pe_1_0_4_add_79_carry_5_), 
        .A2(npu_inst_pe_1_0_4_int_q_acc_5_), .ZN(
        npu_inst_pe_1_0_4_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_0_4_U129 ( .A(npu_inst_pe_1_0_4_int_q_acc_6_), .B(
        npu_inst_pe_1_0_4_add_79_carry_6_), .Z(npu_inst_pe_1_0_4_N79) );
  AND2_X1 npu_inst_pe_1_0_4_U128 ( .A1(npu_inst_pe_1_0_4_add_79_carry_6_), 
        .A2(npu_inst_pe_1_0_4_int_q_acc_6_), .ZN(
        npu_inst_pe_1_0_4_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_0_4_U127 ( .A(npu_inst_pe_1_0_4_int_q_acc_7_), .B(
        npu_inst_pe_1_0_4_add_79_carry_7_), .Z(npu_inst_pe_1_0_4_N80) );
  XNOR2_X1 npu_inst_pe_1_0_4_U126 ( .A(npu_inst_pe_1_0_4_sub_77_carry_2_), .B(
        npu_inst_pe_1_0_4_int_q_acc_2_), .ZN(npu_inst_pe_1_0_4_N67) );
  OR2_X1 npu_inst_pe_1_0_4_U125 ( .A1(npu_inst_pe_1_0_4_int_q_acc_2_), .A2(
        npu_inst_pe_1_0_4_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_0_4_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_0_4_U124 ( .A(npu_inst_pe_1_0_4_sub_77_carry_3_), .B(
        npu_inst_pe_1_0_4_int_q_acc_3_), .ZN(npu_inst_pe_1_0_4_N68) );
  OR2_X1 npu_inst_pe_1_0_4_U123 ( .A1(npu_inst_pe_1_0_4_int_q_acc_3_), .A2(
        npu_inst_pe_1_0_4_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_0_4_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_0_4_U122 ( .A(npu_inst_pe_1_0_4_sub_77_carry_4_), .B(
        npu_inst_pe_1_0_4_int_q_acc_4_), .ZN(npu_inst_pe_1_0_4_N69) );
  OR2_X1 npu_inst_pe_1_0_4_U121 ( .A1(npu_inst_pe_1_0_4_int_q_acc_4_), .A2(
        npu_inst_pe_1_0_4_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_0_4_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_0_4_U120 ( .A(npu_inst_pe_1_0_4_sub_77_carry_5_), .B(
        npu_inst_pe_1_0_4_int_q_acc_5_), .ZN(npu_inst_pe_1_0_4_N70) );
  OR2_X1 npu_inst_pe_1_0_4_U119 ( .A1(npu_inst_pe_1_0_4_int_q_acc_5_), .A2(
        npu_inst_pe_1_0_4_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_0_4_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_0_4_U118 ( .A(npu_inst_pe_1_0_4_sub_77_carry_6_), .B(
        npu_inst_pe_1_0_4_int_q_acc_6_), .ZN(npu_inst_pe_1_0_4_N71) );
  OR2_X1 npu_inst_pe_1_0_4_U117 ( .A1(npu_inst_pe_1_0_4_int_q_acc_6_), .A2(
        npu_inst_pe_1_0_4_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_0_4_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_0_4_U116 ( .A(npu_inst_pe_1_0_4_int_q_acc_7_), .B(
        npu_inst_pe_1_0_4_sub_77_carry_7_), .ZN(npu_inst_pe_1_0_4_N72) );
  INV_X1 npu_inst_pe_1_0_4_U115 ( .A(npu_inst_n79), .ZN(npu_inst_pe_1_0_4_n6)
         );
  INV_X1 npu_inst_pe_1_0_4_U114 ( .A(npu_inst_n60), .ZN(npu_inst_pe_1_0_4_n3)
         );
  AOI22_X1 npu_inst_pe_1_0_4_U113 ( .A1(npu_inst_int_data_y_1__4__0_), .A2(
        npu_inst_pe_1_0_4_n58), .B1(npu_inst_pe_1_0_4_n113), .B2(
        npu_inst_pe_1_0_4_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_0_4_n57) );
  INV_X1 npu_inst_pe_1_0_4_U112 ( .A(npu_inst_pe_1_0_4_n57), .ZN(
        npu_inst_pe_1_0_4_n107) );
  AOI22_X1 npu_inst_pe_1_0_4_U111 ( .A1(npu_inst_int_data_y_1__4__0_), .A2(
        npu_inst_pe_1_0_4_n54), .B1(npu_inst_pe_1_0_4_n114), .B2(
        npu_inst_pe_1_0_4_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_0_4_n53) );
  INV_X1 npu_inst_pe_1_0_4_U110 ( .A(npu_inst_pe_1_0_4_n53), .ZN(
        npu_inst_pe_1_0_4_n108) );
  AOI22_X1 npu_inst_pe_1_0_4_U107 ( .A1(npu_inst_int_data_y_1__4__0_), .A2(
        npu_inst_pe_1_0_4_n50), .B1(npu_inst_pe_1_0_4_n115), .B2(
        npu_inst_pe_1_0_4_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_0_4_n49) );
  INV_X1 npu_inst_pe_1_0_4_U106 ( .A(npu_inst_pe_1_0_4_n49), .ZN(
        npu_inst_pe_1_0_4_n109) );
  AOI22_X1 npu_inst_pe_1_0_4_U105 ( .A1(npu_inst_int_data_y_1__4__0_), .A2(
        npu_inst_pe_1_0_4_n46), .B1(npu_inst_pe_1_0_4_n116), .B2(
        npu_inst_pe_1_0_4_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_0_4_n45) );
  INV_X1 npu_inst_pe_1_0_4_U104 ( .A(npu_inst_pe_1_0_4_n45), .ZN(
        npu_inst_pe_1_0_4_n110) );
  AOI22_X1 npu_inst_pe_1_0_4_U103 ( .A1(npu_inst_int_data_y_1__4__0_), .A2(
        npu_inst_pe_1_0_4_n42), .B1(npu_inst_pe_1_0_4_n118), .B2(
        npu_inst_pe_1_0_4_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_0_4_n41) );
  INV_X1 npu_inst_pe_1_0_4_U102 ( .A(npu_inst_pe_1_0_4_n41), .ZN(
        npu_inst_pe_1_0_4_n111) );
  AOI22_X1 npu_inst_pe_1_0_4_U101 ( .A1(npu_inst_int_data_y_1__4__1_), .A2(
        npu_inst_pe_1_0_4_n58), .B1(npu_inst_pe_1_0_4_n113), .B2(
        npu_inst_pe_1_0_4_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_0_4_n59) );
  INV_X1 npu_inst_pe_1_0_4_U100 ( .A(npu_inst_pe_1_0_4_n59), .ZN(
        npu_inst_pe_1_0_4_n101) );
  AOI22_X1 npu_inst_pe_1_0_4_U99 ( .A1(npu_inst_int_data_y_1__4__1_), .A2(
        npu_inst_pe_1_0_4_n54), .B1(npu_inst_pe_1_0_4_n114), .B2(
        npu_inst_pe_1_0_4_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_0_4_n55) );
  INV_X1 npu_inst_pe_1_0_4_U98 ( .A(npu_inst_pe_1_0_4_n55), .ZN(
        npu_inst_pe_1_0_4_n102) );
  AOI22_X1 npu_inst_pe_1_0_4_U97 ( .A1(npu_inst_int_data_y_1__4__1_), .A2(
        npu_inst_pe_1_0_4_n50), .B1(npu_inst_pe_1_0_4_n115), .B2(
        npu_inst_pe_1_0_4_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_0_4_n51) );
  INV_X1 npu_inst_pe_1_0_4_U96 ( .A(npu_inst_pe_1_0_4_n51), .ZN(
        npu_inst_pe_1_0_4_n103) );
  AOI22_X1 npu_inst_pe_1_0_4_U95 ( .A1(npu_inst_int_data_y_1__4__1_), .A2(
        npu_inst_pe_1_0_4_n46), .B1(npu_inst_pe_1_0_4_n116), .B2(
        npu_inst_pe_1_0_4_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_0_4_n47) );
  INV_X1 npu_inst_pe_1_0_4_U94 ( .A(npu_inst_pe_1_0_4_n47), .ZN(
        npu_inst_pe_1_0_4_n104) );
  AOI22_X1 npu_inst_pe_1_0_4_U93 ( .A1(npu_inst_int_data_y_1__4__1_), .A2(
        npu_inst_pe_1_0_4_n42), .B1(npu_inst_pe_1_0_4_n118), .B2(
        npu_inst_pe_1_0_4_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_0_4_n43) );
  INV_X1 npu_inst_pe_1_0_4_U92 ( .A(npu_inst_pe_1_0_4_n43), .ZN(
        npu_inst_pe_1_0_4_n105) );
  AOI22_X1 npu_inst_pe_1_0_4_U91 ( .A1(npu_inst_pe_1_0_4_n38), .A2(
        npu_inst_int_data_y_1__4__1_), .B1(npu_inst_pe_1_0_4_n117), .B2(
        npu_inst_pe_1_0_4_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_0_4_n39) );
  INV_X1 npu_inst_pe_1_0_4_U90 ( .A(npu_inst_pe_1_0_4_n39), .ZN(
        npu_inst_pe_1_0_4_n106) );
  AOI22_X1 npu_inst_pe_1_0_4_U89 ( .A1(npu_inst_pe_1_0_4_n38), .A2(
        npu_inst_int_data_y_1__4__0_), .B1(npu_inst_pe_1_0_4_n117), .B2(
        npu_inst_pe_1_0_4_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_0_4_n37) );
  INV_X1 npu_inst_pe_1_0_4_U88 ( .A(npu_inst_pe_1_0_4_n37), .ZN(
        npu_inst_pe_1_0_4_n112) );
  AND2_X1 npu_inst_pe_1_0_4_U87 ( .A1(npu_inst_pe_1_0_4_n2), .A2(
        npu_inst_pe_1_0_4_int_q_acc_7_), .ZN(o_data[31]) );
  AND2_X1 npu_inst_pe_1_0_4_U86 ( .A1(npu_inst_pe_1_0_4_int_q_acc_6_), .A2(
        npu_inst_pe_1_0_4_n2), .ZN(o_data[30]) );
  AND2_X1 npu_inst_pe_1_0_4_U85 ( .A1(npu_inst_pe_1_0_4_int_q_acc_5_), .A2(
        npu_inst_pe_1_0_4_n2), .ZN(o_data[29]) );
  AND2_X1 npu_inst_pe_1_0_4_U84 ( .A1(npu_inst_pe_1_0_4_int_q_acc_4_), .A2(
        npu_inst_pe_1_0_4_n2), .ZN(o_data[28]) );
  AND2_X1 npu_inst_pe_1_0_4_U83 ( .A1(npu_inst_pe_1_0_4_int_q_acc_3_), .A2(
        npu_inst_pe_1_0_4_n2), .ZN(o_data[27]) );
  NOR3_X1 npu_inst_pe_1_0_4_U82 ( .A1(npu_inst_pe_1_0_4_n26), .A2(npu_inst_n60), .A3(npu_inst_int_ckg[59]), .ZN(npu_inst_pe_1_0_4_n85) );
  OR2_X1 npu_inst_pe_1_0_4_U81 ( .A1(npu_inst_pe_1_0_4_n85), .A2(
        npu_inst_pe_1_0_4_n2), .ZN(npu_inst_pe_1_0_4_N84) );
  NAND2_X1 npu_inst_pe_1_0_4_U80 ( .A1(npu_inst_pe_1_0_4_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_0_4_n60), .ZN(npu_inst_pe_1_0_4_n74) );
  OAI21_X1 npu_inst_pe_1_0_4_U79 ( .B1(npu_inst_pe_1_0_4_n63), .B2(
        npu_inst_pe_1_0_4_n60), .A(npu_inst_pe_1_0_4_n74), .ZN(
        npu_inst_pe_1_0_4_n97) );
  NAND2_X1 npu_inst_pe_1_0_4_U78 ( .A1(npu_inst_pe_1_0_4_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_0_4_n60), .ZN(npu_inst_pe_1_0_4_n73) );
  OAI21_X1 npu_inst_pe_1_0_4_U77 ( .B1(npu_inst_pe_1_0_4_n61), .B2(
        npu_inst_pe_1_0_4_n60), .A(npu_inst_pe_1_0_4_n73), .ZN(
        npu_inst_pe_1_0_4_n96) );
  NAND2_X1 npu_inst_pe_1_0_4_U76 ( .A1(npu_inst_pe_1_0_4_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_0_4_n56), .ZN(npu_inst_pe_1_0_4_n72) );
  OAI21_X1 npu_inst_pe_1_0_4_U75 ( .B1(npu_inst_pe_1_0_4_n63), .B2(
        npu_inst_pe_1_0_4_n56), .A(npu_inst_pe_1_0_4_n72), .ZN(
        npu_inst_pe_1_0_4_n95) );
  NAND2_X1 npu_inst_pe_1_0_4_U74 ( .A1(npu_inst_pe_1_0_4_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_0_4_n56), .ZN(npu_inst_pe_1_0_4_n71) );
  OAI21_X1 npu_inst_pe_1_0_4_U73 ( .B1(npu_inst_pe_1_0_4_n61), .B2(
        npu_inst_pe_1_0_4_n56), .A(npu_inst_pe_1_0_4_n71), .ZN(
        npu_inst_pe_1_0_4_n94) );
  NAND2_X1 npu_inst_pe_1_0_4_U72 ( .A1(npu_inst_pe_1_0_4_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_0_4_n52), .ZN(npu_inst_pe_1_0_4_n70) );
  OAI21_X1 npu_inst_pe_1_0_4_U71 ( .B1(npu_inst_pe_1_0_4_n63), .B2(
        npu_inst_pe_1_0_4_n52), .A(npu_inst_pe_1_0_4_n70), .ZN(
        npu_inst_pe_1_0_4_n93) );
  NAND2_X1 npu_inst_pe_1_0_4_U70 ( .A1(npu_inst_pe_1_0_4_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_0_4_n52), .ZN(npu_inst_pe_1_0_4_n69) );
  OAI21_X1 npu_inst_pe_1_0_4_U69 ( .B1(npu_inst_pe_1_0_4_n61), .B2(
        npu_inst_pe_1_0_4_n52), .A(npu_inst_pe_1_0_4_n69), .ZN(
        npu_inst_pe_1_0_4_n92) );
  NAND2_X1 npu_inst_pe_1_0_4_U68 ( .A1(npu_inst_pe_1_0_4_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_0_4_n48), .ZN(npu_inst_pe_1_0_4_n68) );
  OAI21_X1 npu_inst_pe_1_0_4_U67 ( .B1(npu_inst_pe_1_0_4_n63), .B2(
        npu_inst_pe_1_0_4_n48), .A(npu_inst_pe_1_0_4_n68), .ZN(
        npu_inst_pe_1_0_4_n91) );
  NAND2_X1 npu_inst_pe_1_0_4_U66 ( .A1(npu_inst_pe_1_0_4_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_0_4_n48), .ZN(npu_inst_pe_1_0_4_n67) );
  OAI21_X1 npu_inst_pe_1_0_4_U65 ( .B1(npu_inst_pe_1_0_4_n61), .B2(
        npu_inst_pe_1_0_4_n48), .A(npu_inst_pe_1_0_4_n67), .ZN(
        npu_inst_pe_1_0_4_n90) );
  NAND2_X1 npu_inst_pe_1_0_4_U64 ( .A1(npu_inst_pe_1_0_4_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_0_4_n44), .ZN(npu_inst_pe_1_0_4_n66) );
  OAI21_X1 npu_inst_pe_1_0_4_U63 ( .B1(npu_inst_pe_1_0_4_n63), .B2(
        npu_inst_pe_1_0_4_n44), .A(npu_inst_pe_1_0_4_n66), .ZN(
        npu_inst_pe_1_0_4_n89) );
  NAND2_X1 npu_inst_pe_1_0_4_U62 ( .A1(npu_inst_pe_1_0_4_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_0_4_n44), .ZN(npu_inst_pe_1_0_4_n65) );
  OAI21_X1 npu_inst_pe_1_0_4_U61 ( .B1(npu_inst_pe_1_0_4_n61), .B2(
        npu_inst_pe_1_0_4_n44), .A(npu_inst_pe_1_0_4_n65), .ZN(
        npu_inst_pe_1_0_4_n88) );
  NAND2_X1 npu_inst_pe_1_0_4_U60 ( .A1(npu_inst_pe_1_0_4_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_0_4_n40), .ZN(npu_inst_pe_1_0_4_n64) );
  OAI21_X1 npu_inst_pe_1_0_4_U59 ( .B1(npu_inst_pe_1_0_4_n63), .B2(
        npu_inst_pe_1_0_4_n40), .A(npu_inst_pe_1_0_4_n64), .ZN(
        npu_inst_pe_1_0_4_n87) );
  NAND2_X1 npu_inst_pe_1_0_4_U58 ( .A1(npu_inst_pe_1_0_4_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_0_4_n40), .ZN(npu_inst_pe_1_0_4_n62) );
  OAI21_X1 npu_inst_pe_1_0_4_U57 ( .B1(npu_inst_pe_1_0_4_n61), .B2(
        npu_inst_pe_1_0_4_n40), .A(npu_inst_pe_1_0_4_n62), .ZN(
        npu_inst_pe_1_0_4_n86) );
  AND2_X1 npu_inst_pe_1_0_4_U56 ( .A1(npu_inst_pe_1_0_4_int_q_acc_0_), .A2(
        npu_inst_pe_1_0_4_n1), .ZN(o_data[24]) );
  AND2_X1 npu_inst_pe_1_0_4_U55 ( .A1(npu_inst_pe_1_0_4_int_q_acc_1_), .A2(
        npu_inst_pe_1_0_4_n1), .ZN(o_data[25]) );
  AND2_X1 npu_inst_pe_1_0_4_U54 ( .A1(npu_inst_pe_1_0_4_int_q_acc_2_), .A2(
        npu_inst_pe_1_0_4_n1), .ZN(o_data[26]) );
  AOI222_X1 npu_inst_pe_1_0_4_U53 ( .A1(npu_inst_int_data_res_1__4__0_), .A2(
        npu_inst_pe_1_0_4_n1), .B1(npu_inst_pe_1_0_4_N73), .B2(
        npu_inst_pe_1_0_4_n76), .C1(npu_inst_pe_1_0_4_N65), .C2(
        npu_inst_pe_1_0_4_n77), .ZN(npu_inst_pe_1_0_4_n84) );
  INV_X1 npu_inst_pe_1_0_4_U52 ( .A(npu_inst_pe_1_0_4_n84), .ZN(
        npu_inst_pe_1_0_4_n100) );
  AOI222_X1 npu_inst_pe_1_0_4_U51 ( .A1(npu_inst_int_data_res_1__4__7_), .A2(
        npu_inst_pe_1_0_4_n1), .B1(npu_inst_pe_1_0_4_N80), .B2(
        npu_inst_pe_1_0_4_n76), .C1(npu_inst_pe_1_0_4_N72), .C2(
        npu_inst_pe_1_0_4_n77), .ZN(npu_inst_pe_1_0_4_n75) );
  INV_X1 npu_inst_pe_1_0_4_U50 ( .A(npu_inst_pe_1_0_4_n75), .ZN(
        npu_inst_pe_1_0_4_n32) );
  AOI222_X1 npu_inst_pe_1_0_4_U49 ( .A1(npu_inst_int_data_res_1__4__1_), .A2(
        npu_inst_pe_1_0_4_n1), .B1(npu_inst_pe_1_0_4_N74), .B2(
        npu_inst_pe_1_0_4_n76), .C1(npu_inst_pe_1_0_4_N66), .C2(
        npu_inst_pe_1_0_4_n77), .ZN(npu_inst_pe_1_0_4_n83) );
  INV_X1 npu_inst_pe_1_0_4_U48 ( .A(npu_inst_pe_1_0_4_n83), .ZN(
        npu_inst_pe_1_0_4_n99) );
  AOI222_X1 npu_inst_pe_1_0_4_U47 ( .A1(npu_inst_int_data_res_1__4__2_), .A2(
        npu_inst_pe_1_0_4_n1), .B1(npu_inst_pe_1_0_4_N75), .B2(
        npu_inst_pe_1_0_4_n76), .C1(npu_inst_pe_1_0_4_N67), .C2(
        npu_inst_pe_1_0_4_n77), .ZN(npu_inst_pe_1_0_4_n82) );
  INV_X1 npu_inst_pe_1_0_4_U46 ( .A(npu_inst_pe_1_0_4_n82), .ZN(
        npu_inst_pe_1_0_4_n98) );
  AOI222_X1 npu_inst_pe_1_0_4_U45 ( .A1(npu_inst_int_data_res_1__4__3_), .A2(
        npu_inst_pe_1_0_4_n1), .B1(npu_inst_pe_1_0_4_N76), .B2(
        npu_inst_pe_1_0_4_n76), .C1(npu_inst_pe_1_0_4_N68), .C2(
        npu_inst_pe_1_0_4_n77), .ZN(npu_inst_pe_1_0_4_n81) );
  INV_X1 npu_inst_pe_1_0_4_U44 ( .A(npu_inst_pe_1_0_4_n81), .ZN(
        npu_inst_pe_1_0_4_n36) );
  AOI222_X1 npu_inst_pe_1_0_4_U43 ( .A1(npu_inst_int_data_res_1__4__4_), .A2(
        npu_inst_pe_1_0_4_n1), .B1(npu_inst_pe_1_0_4_N77), .B2(
        npu_inst_pe_1_0_4_n76), .C1(npu_inst_pe_1_0_4_N69), .C2(
        npu_inst_pe_1_0_4_n77), .ZN(npu_inst_pe_1_0_4_n80) );
  INV_X1 npu_inst_pe_1_0_4_U42 ( .A(npu_inst_pe_1_0_4_n80), .ZN(
        npu_inst_pe_1_0_4_n35) );
  AOI222_X1 npu_inst_pe_1_0_4_U41 ( .A1(npu_inst_int_data_res_1__4__5_), .A2(
        npu_inst_pe_1_0_4_n1), .B1(npu_inst_pe_1_0_4_N78), .B2(
        npu_inst_pe_1_0_4_n76), .C1(npu_inst_pe_1_0_4_N70), .C2(
        npu_inst_pe_1_0_4_n77), .ZN(npu_inst_pe_1_0_4_n79) );
  INV_X1 npu_inst_pe_1_0_4_U40 ( .A(npu_inst_pe_1_0_4_n79), .ZN(
        npu_inst_pe_1_0_4_n34) );
  AOI222_X1 npu_inst_pe_1_0_4_U39 ( .A1(npu_inst_int_data_res_1__4__6_), .A2(
        npu_inst_pe_1_0_4_n1), .B1(npu_inst_pe_1_0_4_N79), .B2(
        npu_inst_pe_1_0_4_n76), .C1(npu_inst_pe_1_0_4_N71), .C2(
        npu_inst_pe_1_0_4_n77), .ZN(npu_inst_pe_1_0_4_n78) );
  INV_X1 npu_inst_pe_1_0_4_U38 ( .A(npu_inst_pe_1_0_4_n78), .ZN(
        npu_inst_pe_1_0_4_n33) );
  INV_X1 npu_inst_pe_1_0_4_U37 ( .A(npu_inst_pe_1_0_4_int_data_1_), .ZN(
        npu_inst_pe_1_0_4_n13) );
  AND2_X1 npu_inst_pe_1_0_4_U36 ( .A1(npu_inst_int_data_x_0__4__1_), .A2(
        npu_inst_pe_1_0_4_int_q_weight_1_), .ZN(npu_inst_pe_1_0_4_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_0_4_U35 ( .A1(npu_inst_int_data_x_0__4__0_), .A2(
        npu_inst_pe_1_0_4_int_q_weight_1_), .ZN(npu_inst_pe_1_0_4_int_data_0_)
         );
  AND2_X1 npu_inst_pe_1_0_4_U34 ( .A1(npu_inst_pe_1_0_4_N93), .A2(npu_inst_n60), .ZN(npu_inst_pe_1_0_4_o_data_v_0_) );
  AND2_X1 npu_inst_pe_1_0_4_U33 ( .A1(npu_inst_n60), .A2(npu_inst_pe_1_0_4_N94), .ZN(npu_inst_pe_1_0_4_o_data_v_1_) );
  AOI22_X1 npu_inst_pe_1_0_4_U32 ( .A1(npu_inst_n60), .A2(
        npu_inst_int_data_y_1__4__1_), .B1(npu_inst_pe_1_0_4_n3), .B2(
        npu_inst_int_data_x_0__5__1_), .ZN(npu_inst_pe_1_0_4_n63) );
  AOI22_X1 npu_inst_pe_1_0_4_U31 ( .A1(npu_inst_n60), .A2(
        npu_inst_int_data_y_1__4__0_), .B1(npu_inst_pe_1_0_4_n3), .B2(
        npu_inst_int_data_x_0__5__0_), .ZN(npu_inst_pe_1_0_4_n61) );
  INV_X1 npu_inst_pe_1_0_4_U30 ( .A(npu_inst_pe_1_0_4_int_data_0_), .ZN(
        npu_inst_pe_1_0_4_n12) );
  INV_X1 npu_inst_pe_1_0_4_U29 ( .A(npu_inst_n71), .ZN(npu_inst_pe_1_0_4_n5)
         );
  OR3_X1 npu_inst_pe_1_0_4_U28 ( .A1(npu_inst_n79), .A2(npu_inst_pe_1_0_4_n7), 
        .A3(npu_inst_pe_1_0_4_n5), .ZN(npu_inst_pe_1_0_4_n56) );
  OR3_X1 npu_inst_pe_1_0_4_U27 ( .A1(npu_inst_pe_1_0_4_n5), .A2(
        npu_inst_pe_1_0_4_n7), .A3(npu_inst_pe_1_0_4_n6), .ZN(
        npu_inst_pe_1_0_4_n48) );
  INV_X1 npu_inst_pe_1_0_4_U26 ( .A(npu_inst_pe_1_0_4_n5), .ZN(
        npu_inst_pe_1_0_4_n4) );
  INV_X1 npu_inst_pe_1_0_4_U25 ( .A(npu_inst_n126), .ZN(npu_inst_pe_1_0_4_n11)
         );
  OR3_X1 npu_inst_pe_1_0_4_U24 ( .A1(npu_inst_pe_1_0_4_n4), .A2(
        npu_inst_pe_1_0_4_n7), .A3(npu_inst_pe_1_0_4_n6), .ZN(
        npu_inst_pe_1_0_4_n52) );
  OR3_X1 npu_inst_pe_1_0_4_U23 ( .A1(npu_inst_n79), .A2(npu_inst_pe_1_0_4_n7), 
        .A3(npu_inst_pe_1_0_4_n4), .ZN(npu_inst_pe_1_0_4_n60) );
  NOR2_X1 npu_inst_pe_1_0_4_U22 ( .A1(npu_inst_pe_1_0_4_n60), .A2(
        npu_inst_pe_1_0_4_n3), .ZN(npu_inst_pe_1_0_4_n58) );
  NOR2_X1 npu_inst_pe_1_0_4_U21 ( .A1(npu_inst_pe_1_0_4_n56), .A2(
        npu_inst_pe_1_0_4_n3), .ZN(npu_inst_pe_1_0_4_n54) );
  NOR2_X1 npu_inst_pe_1_0_4_U20 ( .A1(npu_inst_pe_1_0_4_n52), .A2(
        npu_inst_pe_1_0_4_n3), .ZN(npu_inst_pe_1_0_4_n50) );
  NOR2_X1 npu_inst_pe_1_0_4_U19 ( .A1(npu_inst_pe_1_0_4_n48), .A2(
        npu_inst_pe_1_0_4_n3), .ZN(npu_inst_pe_1_0_4_n46) );
  NOR2_X1 npu_inst_pe_1_0_4_U18 ( .A1(npu_inst_pe_1_0_4_n40), .A2(
        npu_inst_pe_1_0_4_n3), .ZN(npu_inst_pe_1_0_4_n38) );
  NOR2_X1 npu_inst_pe_1_0_4_U17 ( .A1(npu_inst_pe_1_0_4_n44), .A2(
        npu_inst_pe_1_0_4_n3), .ZN(npu_inst_pe_1_0_4_n42) );
  BUF_X1 npu_inst_pe_1_0_4_U16 ( .A(npu_inst_n106), .Z(npu_inst_pe_1_0_4_n7)
         );
  BUF_X1 npu_inst_pe_1_0_4_U15 ( .A(npu_inst_pe_1_0_4_n11), .Z(
        npu_inst_pe_1_0_4_n10) );
  BUF_X1 npu_inst_pe_1_0_4_U14 ( .A(npu_inst_pe_1_0_4_n11), .Z(
        npu_inst_pe_1_0_4_n9) );
  BUF_X1 npu_inst_pe_1_0_4_U13 ( .A(npu_inst_pe_1_0_4_n11), .Z(
        npu_inst_pe_1_0_4_n8) );
  INV_X1 npu_inst_pe_1_0_4_U12 ( .A(npu_inst_pe_1_0_4_n38), .ZN(
        npu_inst_pe_1_0_4_n117) );
  INV_X1 npu_inst_pe_1_0_4_U11 ( .A(npu_inst_pe_1_0_4_n58), .ZN(
        npu_inst_pe_1_0_4_n113) );
  INV_X1 npu_inst_pe_1_0_4_U10 ( .A(npu_inst_pe_1_0_4_n54), .ZN(
        npu_inst_pe_1_0_4_n114) );
  INV_X1 npu_inst_pe_1_0_4_U9 ( .A(npu_inst_pe_1_0_4_n50), .ZN(
        npu_inst_pe_1_0_4_n115) );
  INV_X1 npu_inst_pe_1_0_4_U8 ( .A(npu_inst_pe_1_0_4_n46), .ZN(
        npu_inst_pe_1_0_4_n116) );
  INV_X1 npu_inst_pe_1_0_4_U7 ( .A(npu_inst_pe_1_0_4_n42), .ZN(
        npu_inst_pe_1_0_4_n118) );
  BUF_X1 npu_inst_pe_1_0_4_U6 ( .A(npu_inst_n36), .Z(npu_inst_pe_1_0_4_n2) );
  BUF_X1 npu_inst_pe_1_0_4_U5 ( .A(npu_inst_n36), .Z(npu_inst_pe_1_0_4_n1) );
  NOR2_X1 npu_inst_pe_1_0_4_U4 ( .A1(npu_inst_pe_1_0_4_int_q_weight_0_), .A2(
        npu_inst_pe_1_0_4_n1), .ZN(npu_inst_pe_1_0_4_n76) );
  NOR2_X1 npu_inst_pe_1_0_4_U3 ( .A1(npu_inst_pe_1_0_4_n27), .A2(
        npu_inst_pe_1_0_4_n1), .ZN(npu_inst_pe_1_0_4_n77) );
  FA_X1 npu_inst_pe_1_0_4_sub_77_U2_1 ( .A(npu_inst_pe_1_0_4_int_q_acc_1_), 
        .B(npu_inst_pe_1_0_4_n13), .CI(npu_inst_pe_1_0_4_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_0_4_sub_77_carry_2_), .S(npu_inst_pe_1_0_4_N66) );
  FA_X1 npu_inst_pe_1_0_4_add_79_U1_1 ( .A(npu_inst_pe_1_0_4_int_q_acc_1_), 
        .B(npu_inst_pe_1_0_4_int_data_1_), .CI(
        npu_inst_pe_1_0_4_add_79_carry_1_), .CO(
        npu_inst_pe_1_0_4_add_79_carry_2_), .S(npu_inst_pe_1_0_4_N74) );
  NAND3_X1 npu_inst_pe_1_0_4_U109 ( .A1(npu_inst_pe_1_0_4_n5), .A2(
        npu_inst_pe_1_0_4_n6), .A3(npu_inst_pe_1_0_4_n7), .ZN(
        npu_inst_pe_1_0_4_n44) );
  NAND3_X1 npu_inst_pe_1_0_4_U108 ( .A1(npu_inst_pe_1_0_4_n4), .A2(
        npu_inst_pe_1_0_4_n6), .A3(npu_inst_pe_1_0_4_n7), .ZN(
        npu_inst_pe_1_0_4_n40) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_0_4_n33), .CK(
        npu_inst_pe_1_0_4_net4201), .RN(npu_inst_pe_1_0_4_n8), .Q(
        npu_inst_pe_1_0_4_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_0_4_n34), .CK(
        npu_inst_pe_1_0_4_net4201), .RN(npu_inst_pe_1_0_4_n8), .Q(
        npu_inst_pe_1_0_4_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_0_4_n35), .CK(
        npu_inst_pe_1_0_4_net4201), .RN(npu_inst_pe_1_0_4_n8), .Q(
        npu_inst_pe_1_0_4_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_0_4_n36), .CK(
        npu_inst_pe_1_0_4_net4201), .RN(npu_inst_pe_1_0_4_n8), .Q(
        npu_inst_pe_1_0_4_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_0_4_n98), .CK(
        npu_inst_pe_1_0_4_net4201), .RN(npu_inst_pe_1_0_4_n8), .Q(
        npu_inst_pe_1_0_4_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_0_4_n99), .CK(
        npu_inst_pe_1_0_4_net4201), .RN(npu_inst_pe_1_0_4_n8), .Q(
        npu_inst_pe_1_0_4_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_0_4_n32), .CK(
        npu_inst_pe_1_0_4_net4201), .RN(npu_inst_pe_1_0_4_n8), .Q(
        npu_inst_pe_1_0_4_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_0_4_n100), 
        .CK(npu_inst_pe_1_0_4_net4201), .RN(npu_inst_pe_1_0_4_n8), .Q(
        npu_inst_pe_1_0_4_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_weight_reg_0_ ( .D(npu_inst_n112), .CK(
        npu_inst_pe_1_0_4_net4207), .RN(npu_inst_pe_1_0_4_n8), .Q(
        npu_inst_pe_1_0_4_int_q_weight_0_), .QN(npu_inst_pe_1_0_4_n27) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_weight_reg_1_ ( .D(npu_inst_n118), .CK(
        npu_inst_pe_1_0_4_net4207), .RN(npu_inst_pe_1_0_4_n8), .Q(
        npu_inst_pe_1_0_4_int_q_weight_1_), .QN(npu_inst_pe_1_0_4_n26) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_0_4_n112), 
        .CK(npu_inst_pe_1_0_4_net4207), .RN(npu_inst_pe_1_0_4_n8), .Q(
        npu_inst_pe_1_0_4_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_0_4_n106), 
        .CK(npu_inst_pe_1_0_4_net4207), .RN(npu_inst_pe_1_0_4_n8), .Q(
        npu_inst_pe_1_0_4_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_0_4_n111), 
        .CK(npu_inst_pe_1_0_4_net4207), .RN(npu_inst_pe_1_0_4_n9), .Q(
        npu_inst_pe_1_0_4_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_0_4_n105), 
        .CK(npu_inst_pe_1_0_4_net4207), .RN(npu_inst_pe_1_0_4_n9), .Q(
        npu_inst_pe_1_0_4_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_0_4_n110), 
        .CK(npu_inst_pe_1_0_4_net4207), .RN(npu_inst_pe_1_0_4_n9), .Q(
        npu_inst_pe_1_0_4_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_0_4_n104), 
        .CK(npu_inst_pe_1_0_4_net4207), .RN(npu_inst_pe_1_0_4_n9), .Q(
        npu_inst_pe_1_0_4_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_0_4_n109), 
        .CK(npu_inst_pe_1_0_4_net4207), .RN(npu_inst_pe_1_0_4_n9), .Q(
        npu_inst_pe_1_0_4_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_0_4_n103), 
        .CK(npu_inst_pe_1_0_4_net4207), .RN(npu_inst_pe_1_0_4_n9), .Q(
        npu_inst_pe_1_0_4_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_0_4_n108), 
        .CK(npu_inst_pe_1_0_4_net4207), .RN(npu_inst_pe_1_0_4_n9), .Q(
        npu_inst_pe_1_0_4_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_0_4_n102), 
        .CK(npu_inst_pe_1_0_4_net4207), .RN(npu_inst_pe_1_0_4_n9), .Q(
        npu_inst_pe_1_0_4_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_0_4_n107), 
        .CK(npu_inst_pe_1_0_4_net4207), .RN(npu_inst_pe_1_0_4_n9), .Q(
        npu_inst_pe_1_0_4_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_0_4_n101), 
        .CK(npu_inst_pe_1_0_4_net4207), .RN(npu_inst_pe_1_0_4_n9), .Q(
        npu_inst_pe_1_0_4_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_0_4_n86), 
        .CK(npu_inst_pe_1_0_4_net4207), .RN(npu_inst_pe_1_0_4_n9), .Q(
        npu_inst_pe_1_0_4_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_0_4_n87), 
        .CK(npu_inst_pe_1_0_4_net4207), .RN(npu_inst_pe_1_0_4_n9), .Q(
        npu_inst_pe_1_0_4_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_0_4_n88), 
        .CK(npu_inst_pe_1_0_4_net4207), .RN(npu_inst_pe_1_0_4_n10), .Q(
        npu_inst_pe_1_0_4_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_0_4_n89), 
        .CK(npu_inst_pe_1_0_4_net4207), .RN(npu_inst_pe_1_0_4_n10), .Q(
        npu_inst_pe_1_0_4_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_0_4_n90), 
        .CK(npu_inst_pe_1_0_4_net4207), .RN(npu_inst_pe_1_0_4_n10), .Q(
        npu_inst_pe_1_0_4_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_0_4_n91), 
        .CK(npu_inst_pe_1_0_4_net4207), .RN(npu_inst_pe_1_0_4_n10), .Q(
        npu_inst_pe_1_0_4_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_0_4_n92), 
        .CK(npu_inst_pe_1_0_4_net4207), .RN(npu_inst_pe_1_0_4_n10), .Q(
        npu_inst_pe_1_0_4_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_0_4_n93), 
        .CK(npu_inst_pe_1_0_4_net4207), .RN(npu_inst_pe_1_0_4_n10), .Q(
        npu_inst_pe_1_0_4_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_0_4_n94), 
        .CK(npu_inst_pe_1_0_4_net4207), .RN(npu_inst_pe_1_0_4_n10), .Q(
        npu_inst_pe_1_0_4_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_0_4_n95), 
        .CK(npu_inst_pe_1_0_4_net4207), .RN(npu_inst_pe_1_0_4_n10), .Q(
        npu_inst_pe_1_0_4_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_0_4_n96), 
        .CK(npu_inst_pe_1_0_4_net4207), .RN(npu_inst_pe_1_0_4_n10), .Q(
        npu_inst_pe_1_0_4_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_0_4_n97), 
        .CK(npu_inst_pe_1_0_4_net4207), .RN(npu_inst_pe_1_0_4_n10), .Q(
        npu_inst_pe_1_0_4_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_0_4_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_0_4_N84), .SE(1'b0), .GCK(npu_inst_pe_1_0_4_net4201) );
  CLKGATETST_X1 npu_inst_pe_1_0_4_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n66), .SE(1'b0), .GCK(npu_inst_pe_1_0_4_net4207) );
  MUX2_X1 npu_inst_pe_1_0_5_U162 ( .A(npu_inst_pe_1_0_5_n32), .B(
        npu_inst_pe_1_0_5_n29), .S(npu_inst_pe_1_0_5_n8), .Z(
        npu_inst_pe_1_0_5_N93) );
  MUX2_X1 npu_inst_pe_1_0_5_U161 ( .A(npu_inst_pe_1_0_5_n31), .B(
        npu_inst_pe_1_0_5_n30), .S(npu_inst_pe_1_0_5_n6), .Z(
        npu_inst_pe_1_0_5_n32) );
  MUX2_X1 npu_inst_pe_1_0_5_U160 ( .A(npu_inst_pe_1_0_5_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_0_5_int_q_reg_v_1__0_), .S(npu_inst_pe_1_0_5_n4), .Z(
        npu_inst_pe_1_0_5_n31) );
  MUX2_X1 npu_inst_pe_1_0_5_U159 ( .A(npu_inst_pe_1_0_5_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_0_5_int_q_reg_v_3__0_), .S(npu_inst_pe_1_0_5_n4), .Z(
        npu_inst_pe_1_0_5_n30) );
  MUX2_X1 npu_inst_pe_1_0_5_U158 ( .A(npu_inst_pe_1_0_5_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_0_5_int_q_reg_v_5__0_), .S(npu_inst_pe_1_0_5_n4), .Z(
        npu_inst_pe_1_0_5_n29) );
  MUX2_X1 npu_inst_pe_1_0_5_U157 ( .A(npu_inst_pe_1_0_5_n28), .B(
        npu_inst_pe_1_0_5_n23), .S(npu_inst_pe_1_0_5_n8), .Z(
        npu_inst_pe_1_0_5_N94) );
  MUX2_X1 npu_inst_pe_1_0_5_U156 ( .A(npu_inst_pe_1_0_5_n25), .B(
        npu_inst_pe_1_0_5_n24), .S(npu_inst_pe_1_0_5_n6), .Z(
        npu_inst_pe_1_0_5_n28) );
  MUX2_X1 npu_inst_pe_1_0_5_U155 ( .A(npu_inst_pe_1_0_5_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_0_5_int_q_reg_v_1__1_), .S(npu_inst_pe_1_0_5_n4), .Z(
        npu_inst_pe_1_0_5_n25) );
  MUX2_X1 npu_inst_pe_1_0_5_U154 ( .A(npu_inst_pe_1_0_5_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_0_5_int_q_reg_v_3__1_), .S(npu_inst_pe_1_0_5_n4), .Z(
        npu_inst_pe_1_0_5_n24) );
  MUX2_X1 npu_inst_pe_1_0_5_U153 ( .A(npu_inst_pe_1_0_5_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_0_5_int_q_reg_v_5__1_), .S(npu_inst_pe_1_0_5_n4), .Z(
        npu_inst_pe_1_0_5_n23) );
  MUX2_X1 npu_inst_pe_1_0_5_U152 ( .A(npu_inst_pe_1_0_5_n22), .B(
        npu_inst_pe_1_0_5_n19), .S(npu_inst_pe_1_0_5_n8), .Z(
        npu_inst_int_data_x_0__5__1_) );
  MUX2_X1 npu_inst_pe_1_0_5_U151 ( .A(npu_inst_pe_1_0_5_n21), .B(
        npu_inst_pe_1_0_5_n20), .S(npu_inst_pe_1_0_5_n6), .Z(
        npu_inst_pe_1_0_5_n22) );
  MUX2_X1 npu_inst_pe_1_0_5_U150 ( .A(npu_inst_pe_1_0_5_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_0_5_int_q_reg_h_1__1_), .S(npu_inst_pe_1_0_5_n4), .Z(
        npu_inst_pe_1_0_5_n21) );
  MUX2_X1 npu_inst_pe_1_0_5_U149 ( .A(npu_inst_pe_1_0_5_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_0_5_int_q_reg_h_3__1_), .S(npu_inst_pe_1_0_5_n4), .Z(
        npu_inst_pe_1_0_5_n20) );
  MUX2_X1 npu_inst_pe_1_0_5_U148 ( .A(npu_inst_pe_1_0_5_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_0_5_int_q_reg_h_5__1_), .S(npu_inst_pe_1_0_5_n4), .Z(
        npu_inst_pe_1_0_5_n19) );
  MUX2_X1 npu_inst_pe_1_0_5_U147 ( .A(npu_inst_pe_1_0_5_n18), .B(
        npu_inst_pe_1_0_5_n15), .S(npu_inst_pe_1_0_5_n8), .Z(
        npu_inst_int_data_x_0__5__0_) );
  MUX2_X1 npu_inst_pe_1_0_5_U146 ( .A(npu_inst_pe_1_0_5_n17), .B(
        npu_inst_pe_1_0_5_n16), .S(npu_inst_pe_1_0_5_n6), .Z(
        npu_inst_pe_1_0_5_n18) );
  MUX2_X1 npu_inst_pe_1_0_5_U145 ( .A(npu_inst_pe_1_0_5_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_0_5_int_q_reg_h_1__0_), .S(npu_inst_pe_1_0_5_n4), .Z(
        npu_inst_pe_1_0_5_n17) );
  MUX2_X1 npu_inst_pe_1_0_5_U144 ( .A(npu_inst_pe_1_0_5_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_0_5_int_q_reg_h_3__0_), .S(npu_inst_pe_1_0_5_n4), .Z(
        npu_inst_pe_1_0_5_n16) );
  MUX2_X1 npu_inst_pe_1_0_5_U143 ( .A(npu_inst_pe_1_0_5_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_0_5_int_q_reg_h_5__0_), .S(npu_inst_pe_1_0_5_n4), .Z(
        npu_inst_pe_1_0_5_n15) );
  XOR2_X1 npu_inst_pe_1_0_5_U142 ( .A(npu_inst_pe_1_0_5_int_data_0_), .B(
        npu_inst_pe_1_0_5_int_q_acc_0_), .Z(npu_inst_pe_1_0_5_N73) );
  AND2_X1 npu_inst_pe_1_0_5_U141 ( .A1(npu_inst_pe_1_0_5_int_q_acc_0_), .A2(
        npu_inst_pe_1_0_5_int_data_0_), .ZN(npu_inst_pe_1_0_5_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_0_5_U140 ( .A(npu_inst_pe_1_0_5_int_q_acc_0_), .B(
        npu_inst_pe_1_0_5_n13), .ZN(npu_inst_pe_1_0_5_N65) );
  OR2_X1 npu_inst_pe_1_0_5_U139 ( .A1(npu_inst_pe_1_0_5_n13), .A2(
        npu_inst_pe_1_0_5_int_q_acc_0_), .ZN(npu_inst_pe_1_0_5_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_0_5_U138 ( .A(npu_inst_pe_1_0_5_int_q_acc_2_), .B(
        npu_inst_pe_1_0_5_add_79_carry_2_), .Z(npu_inst_pe_1_0_5_N75) );
  AND2_X1 npu_inst_pe_1_0_5_U137 ( .A1(npu_inst_pe_1_0_5_add_79_carry_2_), 
        .A2(npu_inst_pe_1_0_5_int_q_acc_2_), .ZN(
        npu_inst_pe_1_0_5_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_0_5_U136 ( .A(npu_inst_pe_1_0_5_int_q_acc_3_), .B(
        npu_inst_pe_1_0_5_add_79_carry_3_), .Z(npu_inst_pe_1_0_5_N76) );
  AND2_X1 npu_inst_pe_1_0_5_U135 ( .A1(npu_inst_pe_1_0_5_add_79_carry_3_), 
        .A2(npu_inst_pe_1_0_5_int_q_acc_3_), .ZN(
        npu_inst_pe_1_0_5_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_0_5_U134 ( .A(npu_inst_pe_1_0_5_int_q_acc_4_), .B(
        npu_inst_pe_1_0_5_add_79_carry_4_), .Z(npu_inst_pe_1_0_5_N77) );
  AND2_X1 npu_inst_pe_1_0_5_U133 ( .A1(npu_inst_pe_1_0_5_add_79_carry_4_), 
        .A2(npu_inst_pe_1_0_5_int_q_acc_4_), .ZN(
        npu_inst_pe_1_0_5_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_0_5_U132 ( .A(npu_inst_pe_1_0_5_int_q_acc_5_), .B(
        npu_inst_pe_1_0_5_add_79_carry_5_), .Z(npu_inst_pe_1_0_5_N78) );
  AND2_X1 npu_inst_pe_1_0_5_U131 ( .A1(npu_inst_pe_1_0_5_add_79_carry_5_), 
        .A2(npu_inst_pe_1_0_5_int_q_acc_5_), .ZN(
        npu_inst_pe_1_0_5_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_0_5_U130 ( .A(npu_inst_pe_1_0_5_int_q_acc_6_), .B(
        npu_inst_pe_1_0_5_add_79_carry_6_), .Z(npu_inst_pe_1_0_5_N79) );
  AND2_X1 npu_inst_pe_1_0_5_U129 ( .A1(npu_inst_pe_1_0_5_add_79_carry_6_), 
        .A2(npu_inst_pe_1_0_5_int_q_acc_6_), .ZN(
        npu_inst_pe_1_0_5_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_0_5_U128 ( .A(npu_inst_pe_1_0_5_int_q_acc_7_), .B(
        npu_inst_pe_1_0_5_add_79_carry_7_), .Z(npu_inst_pe_1_0_5_N80) );
  XNOR2_X1 npu_inst_pe_1_0_5_U127 ( .A(npu_inst_pe_1_0_5_sub_77_carry_2_), .B(
        npu_inst_pe_1_0_5_int_q_acc_2_), .ZN(npu_inst_pe_1_0_5_N67) );
  OR2_X1 npu_inst_pe_1_0_5_U126 ( .A1(npu_inst_pe_1_0_5_int_q_acc_2_), .A2(
        npu_inst_pe_1_0_5_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_0_5_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_0_5_U125 ( .A(npu_inst_pe_1_0_5_sub_77_carry_3_), .B(
        npu_inst_pe_1_0_5_int_q_acc_3_), .ZN(npu_inst_pe_1_0_5_N68) );
  OR2_X1 npu_inst_pe_1_0_5_U124 ( .A1(npu_inst_pe_1_0_5_int_q_acc_3_), .A2(
        npu_inst_pe_1_0_5_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_0_5_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_0_5_U123 ( .A(npu_inst_pe_1_0_5_sub_77_carry_4_), .B(
        npu_inst_pe_1_0_5_int_q_acc_4_), .ZN(npu_inst_pe_1_0_5_N69) );
  OR2_X1 npu_inst_pe_1_0_5_U122 ( .A1(npu_inst_pe_1_0_5_int_q_acc_4_), .A2(
        npu_inst_pe_1_0_5_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_0_5_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_0_5_U121 ( .A(npu_inst_pe_1_0_5_sub_77_carry_5_), .B(
        npu_inst_pe_1_0_5_int_q_acc_5_), .ZN(npu_inst_pe_1_0_5_N70) );
  OR2_X1 npu_inst_pe_1_0_5_U120 ( .A1(npu_inst_pe_1_0_5_int_q_acc_5_), .A2(
        npu_inst_pe_1_0_5_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_0_5_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_0_5_U119 ( .A(npu_inst_pe_1_0_5_sub_77_carry_6_), .B(
        npu_inst_pe_1_0_5_int_q_acc_6_), .ZN(npu_inst_pe_1_0_5_N71) );
  OR2_X1 npu_inst_pe_1_0_5_U118 ( .A1(npu_inst_pe_1_0_5_int_q_acc_6_), .A2(
        npu_inst_pe_1_0_5_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_0_5_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_0_5_U117 ( .A(npu_inst_pe_1_0_5_int_q_acc_7_), .B(
        npu_inst_pe_1_0_5_sub_77_carry_7_), .ZN(npu_inst_pe_1_0_5_N72) );
  INV_X1 npu_inst_pe_1_0_5_U116 ( .A(npu_inst_n79), .ZN(npu_inst_pe_1_0_5_n7)
         );
  INV_X1 npu_inst_pe_1_0_5_U115 ( .A(npu_inst_pe_1_0_5_n7), .ZN(
        npu_inst_pe_1_0_5_n6) );
  INV_X1 npu_inst_pe_1_0_5_U114 ( .A(npu_inst_n60), .ZN(npu_inst_pe_1_0_5_n3)
         );
  AOI22_X1 npu_inst_pe_1_0_5_U113 ( .A1(npu_inst_int_data_y_1__5__0_), .A2(
        npu_inst_pe_1_0_5_n58), .B1(npu_inst_pe_1_0_5_n114), .B2(
        npu_inst_pe_1_0_5_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_0_5_n57) );
  INV_X1 npu_inst_pe_1_0_5_U112 ( .A(npu_inst_pe_1_0_5_n57), .ZN(
        npu_inst_pe_1_0_5_n108) );
  AOI22_X1 npu_inst_pe_1_0_5_U111 ( .A1(npu_inst_int_data_y_1__5__0_), .A2(
        npu_inst_pe_1_0_5_n54), .B1(npu_inst_pe_1_0_5_n115), .B2(
        npu_inst_pe_1_0_5_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_0_5_n53) );
  INV_X1 npu_inst_pe_1_0_5_U110 ( .A(npu_inst_pe_1_0_5_n53), .ZN(
        npu_inst_pe_1_0_5_n109) );
  AOI22_X1 npu_inst_pe_1_0_5_U107 ( .A1(npu_inst_int_data_y_1__5__0_), .A2(
        npu_inst_pe_1_0_5_n50), .B1(npu_inst_pe_1_0_5_n116), .B2(
        npu_inst_pe_1_0_5_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_0_5_n49) );
  INV_X1 npu_inst_pe_1_0_5_U106 ( .A(npu_inst_pe_1_0_5_n49), .ZN(
        npu_inst_pe_1_0_5_n110) );
  AOI22_X1 npu_inst_pe_1_0_5_U105 ( .A1(npu_inst_int_data_y_1__5__0_), .A2(
        npu_inst_pe_1_0_5_n46), .B1(npu_inst_pe_1_0_5_n117), .B2(
        npu_inst_pe_1_0_5_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_0_5_n45) );
  INV_X1 npu_inst_pe_1_0_5_U104 ( .A(npu_inst_pe_1_0_5_n45), .ZN(
        npu_inst_pe_1_0_5_n111) );
  AOI22_X1 npu_inst_pe_1_0_5_U103 ( .A1(npu_inst_int_data_y_1__5__0_), .A2(
        npu_inst_pe_1_0_5_n42), .B1(npu_inst_pe_1_0_5_n119), .B2(
        npu_inst_pe_1_0_5_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_0_5_n41) );
  INV_X1 npu_inst_pe_1_0_5_U102 ( .A(npu_inst_pe_1_0_5_n41), .ZN(
        npu_inst_pe_1_0_5_n112) );
  AOI22_X1 npu_inst_pe_1_0_5_U101 ( .A1(npu_inst_int_data_y_1__5__1_), .A2(
        npu_inst_pe_1_0_5_n58), .B1(npu_inst_pe_1_0_5_n114), .B2(
        npu_inst_pe_1_0_5_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_0_5_n59) );
  INV_X1 npu_inst_pe_1_0_5_U100 ( .A(npu_inst_pe_1_0_5_n59), .ZN(
        npu_inst_pe_1_0_5_n102) );
  AOI22_X1 npu_inst_pe_1_0_5_U99 ( .A1(npu_inst_int_data_y_1__5__1_), .A2(
        npu_inst_pe_1_0_5_n54), .B1(npu_inst_pe_1_0_5_n115), .B2(
        npu_inst_pe_1_0_5_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_0_5_n55) );
  INV_X1 npu_inst_pe_1_0_5_U98 ( .A(npu_inst_pe_1_0_5_n55), .ZN(
        npu_inst_pe_1_0_5_n103) );
  AOI22_X1 npu_inst_pe_1_0_5_U97 ( .A1(npu_inst_int_data_y_1__5__1_), .A2(
        npu_inst_pe_1_0_5_n50), .B1(npu_inst_pe_1_0_5_n116), .B2(
        npu_inst_pe_1_0_5_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_0_5_n51) );
  INV_X1 npu_inst_pe_1_0_5_U96 ( .A(npu_inst_pe_1_0_5_n51), .ZN(
        npu_inst_pe_1_0_5_n104) );
  AOI22_X1 npu_inst_pe_1_0_5_U95 ( .A1(npu_inst_int_data_y_1__5__1_), .A2(
        npu_inst_pe_1_0_5_n46), .B1(npu_inst_pe_1_0_5_n117), .B2(
        npu_inst_pe_1_0_5_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_0_5_n47) );
  INV_X1 npu_inst_pe_1_0_5_U94 ( .A(npu_inst_pe_1_0_5_n47), .ZN(
        npu_inst_pe_1_0_5_n105) );
  AOI22_X1 npu_inst_pe_1_0_5_U93 ( .A1(npu_inst_int_data_y_1__5__1_), .A2(
        npu_inst_pe_1_0_5_n42), .B1(npu_inst_pe_1_0_5_n119), .B2(
        npu_inst_pe_1_0_5_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_0_5_n43) );
  INV_X1 npu_inst_pe_1_0_5_U92 ( .A(npu_inst_pe_1_0_5_n43), .ZN(
        npu_inst_pe_1_0_5_n106) );
  AOI22_X1 npu_inst_pe_1_0_5_U91 ( .A1(npu_inst_pe_1_0_5_n38), .A2(
        npu_inst_int_data_y_1__5__1_), .B1(npu_inst_pe_1_0_5_n118), .B2(
        npu_inst_pe_1_0_5_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_0_5_n39) );
  INV_X1 npu_inst_pe_1_0_5_U90 ( .A(npu_inst_pe_1_0_5_n39), .ZN(
        npu_inst_pe_1_0_5_n107) );
  AOI22_X1 npu_inst_pe_1_0_5_U89 ( .A1(npu_inst_pe_1_0_5_n38), .A2(
        npu_inst_int_data_y_1__5__0_), .B1(npu_inst_pe_1_0_5_n118), .B2(
        npu_inst_pe_1_0_5_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_0_5_n37) );
  INV_X1 npu_inst_pe_1_0_5_U88 ( .A(npu_inst_pe_1_0_5_n37), .ZN(
        npu_inst_pe_1_0_5_n113) );
  AND2_X1 npu_inst_pe_1_0_5_U87 ( .A1(npu_inst_pe_1_0_5_n2), .A2(
        npu_inst_pe_1_0_5_int_q_acc_7_), .ZN(o_data[23]) );
  AND2_X1 npu_inst_pe_1_0_5_U86 ( .A1(npu_inst_pe_1_0_5_int_q_acc_6_), .A2(
        npu_inst_pe_1_0_5_n2), .ZN(o_data[22]) );
  AND2_X1 npu_inst_pe_1_0_5_U85 ( .A1(npu_inst_pe_1_0_5_int_q_acc_5_), .A2(
        npu_inst_pe_1_0_5_n2), .ZN(o_data[21]) );
  AND2_X1 npu_inst_pe_1_0_5_U84 ( .A1(npu_inst_pe_1_0_5_int_q_acc_4_), .A2(
        npu_inst_pe_1_0_5_n2), .ZN(o_data[20]) );
  AND2_X1 npu_inst_pe_1_0_5_U83 ( .A1(npu_inst_pe_1_0_5_int_q_acc_3_), .A2(
        npu_inst_pe_1_0_5_n2), .ZN(o_data[19]) );
  NAND2_X1 npu_inst_pe_1_0_5_U82 ( .A1(npu_inst_pe_1_0_5_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_0_5_n60), .ZN(npu_inst_pe_1_0_5_n74) );
  OAI21_X1 npu_inst_pe_1_0_5_U81 ( .B1(npu_inst_pe_1_0_5_n63), .B2(
        npu_inst_pe_1_0_5_n60), .A(npu_inst_pe_1_0_5_n74), .ZN(
        npu_inst_pe_1_0_5_n97) );
  NAND2_X1 npu_inst_pe_1_0_5_U80 ( .A1(npu_inst_pe_1_0_5_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_0_5_n60), .ZN(npu_inst_pe_1_0_5_n73) );
  OAI21_X1 npu_inst_pe_1_0_5_U79 ( .B1(npu_inst_pe_1_0_5_n61), .B2(
        npu_inst_pe_1_0_5_n60), .A(npu_inst_pe_1_0_5_n73), .ZN(
        npu_inst_pe_1_0_5_n96) );
  NAND2_X1 npu_inst_pe_1_0_5_U78 ( .A1(npu_inst_pe_1_0_5_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_0_5_n56), .ZN(npu_inst_pe_1_0_5_n72) );
  OAI21_X1 npu_inst_pe_1_0_5_U77 ( .B1(npu_inst_pe_1_0_5_n63), .B2(
        npu_inst_pe_1_0_5_n56), .A(npu_inst_pe_1_0_5_n72), .ZN(
        npu_inst_pe_1_0_5_n95) );
  NAND2_X1 npu_inst_pe_1_0_5_U76 ( .A1(npu_inst_pe_1_0_5_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_0_5_n56), .ZN(npu_inst_pe_1_0_5_n71) );
  OAI21_X1 npu_inst_pe_1_0_5_U75 ( .B1(npu_inst_pe_1_0_5_n61), .B2(
        npu_inst_pe_1_0_5_n56), .A(npu_inst_pe_1_0_5_n71), .ZN(
        npu_inst_pe_1_0_5_n94) );
  NAND2_X1 npu_inst_pe_1_0_5_U74 ( .A1(npu_inst_pe_1_0_5_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_0_5_n52), .ZN(npu_inst_pe_1_0_5_n70) );
  OAI21_X1 npu_inst_pe_1_0_5_U73 ( .B1(npu_inst_pe_1_0_5_n63), .B2(
        npu_inst_pe_1_0_5_n52), .A(npu_inst_pe_1_0_5_n70), .ZN(
        npu_inst_pe_1_0_5_n93) );
  NAND2_X1 npu_inst_pe_1_0_5_U72 ( .A1(npu_inst_pe_1_0_5_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_0_5_n52), .ZN(npu_inst_pe_1_0_5_n69) );
  OAI21_X1 npu_inst_pe_1_0_5_U71 ( .B1(npu_inst_pe_1_0_5_n61), .B2(
        npu_inst_pe_1_0_5_n52), .A(npu_inst_pe_1_0_5_n69), .ZN(
        npu_inst_pe_1_0_5_n92) );
  NAND2_X1 npu_inst_pe_1_0_5_U70 ( .A1(npu_inst_pe_1_0_5_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_0_5_n48), .ZN(npu_inst_pe_1_0_5_n68) );
  OAI21_X1 npu_inst_pe_1_0_5_U69 ( .B1(npu_inst_pe_1_0_5_n63), .B2(
        npu_inst_pe_1_0_5_n48), .A(npu_inst_pe_1_0_5_n68), .ZN(
        npu_inst_pe_1_0_5_n91) );
  NAND2_X1 npu_inst_pe_1_0_5_U68 ( .A1(npu_inst_pe_1_0_5_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_0_5_n48), .ZN(npu_inst_pe_1_0_5_n67) );
  OAI21_X1 npu_inst_pe_1_0_5_U67 ( .B1(npu_inst_pe_1_0_5_n61), .B2(
        npu_inst_pe_1_0_5_n48), .A(npu_inst_pe_1_0_5_n67), .ZN(
        npu_inst_pe_1_0_5_n90) );
  NAND2_X1 npu_inst_pe_1_0_5_U66 ( .A1(npu_inst_pe_1_0_5_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_0_5_n44), .ZN(npu_inst_pe_1_0_5_n66) );
  OAI21_X1 npu_inst_pe_1_0_5_U65 ( .B1(npu_inst_pe_1_0_5_n63), .B2(
        npu_inst_pe_1_0_5_n44), .A(npu_inst_pe_1_0_5_n66), .ZN(
        npu_inst_pe_1_0_5_n89) );
  NAND2_X1 npu_inst_pe_1_0_5_U64 ( .A1(npu_inst_pe_1_0_5_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_0_5_n44), .ZN(npu_inst_pe_1_0_5_n65) );
  OAI21_X1 npu_inst_pe_1_0_5_U63 ( .B1(npu_inst_pe_1_0_5_n61), .B2(
        npu_inst_pe_1_0_5_n44), .A(npu_inst_pe_1_0_5_n65), .ZN(
        npu_inst_pe_1_0_5_n88) );
  NAND2_X1 npu_inst_pe_1_0_5_U62 ( .A1(npu_inst_pe_1_0_5_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_0_5_n40), .ZN(npu_inst_pe_1_0_5_n64) );
  OAI21_X1 npu_inst_pe_1_0_5_U61 ( .B1(npu_inst_pe_1_0_5_n63), .B2(
        npu_inst_pe_1_0_5_n40), .A(npu_inst_pe_1_0_5_n64), .ZN(
        npu_inst_pe_1_0_5_n87) );
  NAND2_X1 npu_inst_pe_1_0_5_U60 ( .A1(npu_inst_pe_1_0_5_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_0_5_n40), .ZN(npu_inst_pe_1_0_5_n62) );
  OAI21_X1 npu_inst_pe_1_0_5_U59 ( .B1(npu_inst_pe_1_0_5_n61), .B2(
        npu_inst_pe_1_0_5_n40), .A(npu_inst_pe_1_0_5_n62), .ZN(
        npu_inst_pe_1_0_5_n86) );
  NOR3_X1 npu_inst_pe_1_0_5_U58 ( .A1(npu_inst_pe_1_0_5_n26), .A2(npu_inst_n60), .A3(npu_inst_int_ckg[58]), .ZN(npu_inst_pe_1_0_5_n85) );
  OR2_X1 npu_inst_pe_1_0_5_U57 ( .A1(npu_inst_pe_1_0_5_n85), .A2(
        npu_inst_pe_1_0_5_n2), .ZN(npu_inst_pe_1_0_5_N84) );
  AND2_X1 npu_inst_pe_1_0_5_U56 ( .A1(npu_inst_pe_1_0_5_int_q_acc_0_), .A2(
        npu_inst_pe_1_0_5_n1), .ZN(o_data[16]) );
  AND2_X1 npu_inst_pe_1_0_5_U55 ( .A1(npu_inst_pe_1_0_5_int_q_acc_1_), .A2(
        npu_inst_pe_1_0_5_n1), .ZN(o_data[17]) );
  AND2_X1 npu_inst_pe_1_0_5_U54 ( .A1(npu_inst_pe_1_0_5_int_q_acc_2_), .A2(
        npu_inst_pe_1_0_5_n1), .ZN(o_data[18]) );
  AOI222_X1 npu_inst_pe_1_0_5_U53 ( .A1(npu_inst_int_data_res_1__5__0_), .A2(
        npu_inst_pe_1_0_5_n1), .B1(npu_inst_pe_1_0_5_N73), .B2(
        npu_inst_pe_1_0_5_n76), .C1(npu_inst_pe_1_0_5_N65), .C2(
        npu_inst_pe_1_0_5_n77), .ZN(npu_inst_pe_1_0_5_n84) );
  INV_X1 npu_inst_pe_1_0_5_U52 ( .A(npu_inst_pe_1_0_5_n84), .ZN(
        npu_inst_pe_1_0_5_n101) );
  AOI222_X1 npu_inst_pe_1_0_5_U51 ( .A1(npu_inst_int_data_res_1__5__7_), .A2(
        npu_inst_pe_1_0_5_n1), .B1(npu_inst_pe_1_0_5_N80), .B2(
        npu_inst_pe_1_0_5_n76), .C1(npu_inst_pe_1_0_5_N72), .C2(
        npu_inst_pe_1_0_5_n77), .ZN(npu_inst_pe_1_0_5_n75) );
  INV_X1 npu_inst_pe_1_0_5_U50 ( .A(npu_inst_pe_1_0_5_n75), .ZN(
        npu_inst_pe_1_0_5_n33) );
  AOI222_X1 npu_inst_pe_1_0_5_U49 ( .A1(npu_inst_int_data_res_1__5__1_), .A2(
        npu_inst_pe_1_0_5_n1), .B1(npu_inst_pe_1_0_5_N74), .B2(
        npu_inst_pe_1_0_5_n76), .C1(npu_inst_pe_1_0_5_N66), .C2(
        npu_inst_pe_1_0_5_n77), .ZN(npu_inst_pe_1_0_5_n83) );
  INV_X1 npu_inst_pe_1_0_5_U48 ( .A(npu_inst_pe_1_0_5_n83), .ZN(
        npu_inst_pe_1_0_5_n100) );
  AOI222_X1 npu_inst_pe_1_0_5_U47 ( .A1(npu_inst_int_data_res_1__5__2_), .A2(
        npu_inst_pe_1_0_5_n1), .B1(npu_inst_pe_1_0_5_N75), .B2(
        npu_inst_pe_1_0_5_n76), .C1(npu_inst_pe_1_0_5_N67), .C2(
        npu_inst_pe_1_0_5_n77), .ZN(npu_inst_pe_1_0_5_n82) );
  INV_X1 npu_inst_pe_1_0_5_U46 ( .A(npu_inst_pe_1_0_5_n82), .ZN(
        npu_inst_pe_1_0_5_n99) );
  AOI222_X1 npu_inst_pe_1_0_5_U45 ( .A1(npu_inst_int_data_res_1__5__3_), .A2(
        npu_inst_pe_1_0_5_n1), .B1(npu_inst_pe_1_0_5_N76), .B2(
        npu_inst_pe_1_0_5_n76), .C1(npu_inst_pe_1_0_5_N68), .C2(
        npu_inst_pe_1_0_5_n77), .ZN(npu_inst_pe_1_0_5_n81) );
  INV_X1 npu_inst_pe_1_0_5_U44 ( .A(npu_inst_pe_1_0_5_n81), .ZN(
        npu_inst_pe_1_0_5_n98) );
  AOI222_X1 npu_inst_pe_1_0_5_U43 ( .A1(npu_inst_int_data_res_1__5__4_), .A2(
        npu_inst_pe_1_0_5_n1), .B1(npu_inst_pe_1_0_5_N77), .B2(
        npu_inst_pe_1_0_5_n76), .C1(npu_inst_pe_1_0_5_N69), .C2(
        npu_inst_pe_1_0_5_n77), .ZN(npu_inst_pe_1_0_5_n80) );
  INV_X1 npu_inst_pe_1_0_5_U42 ( .A(npu_inst_pe_1_0_5_n80), .ZN(
        npu_inst_pe_1_0_5_n36) );
  AOI222_X1 npu_inst_pe_1_0_5_U41 ( .A1(npu_inst_int_data_res_1__5__5_), .A2(
        npu_inst_pe_1_0_5_n1), .B1(npu_inst_pe_1_0_5_N78), .B2(
        npu_inst_pe_1_0_5_n76), .C1(npu_inst_pe_1_0_5_N70), .C2(
        npu_inst_pe_1_0_5_n77), .ZN(npu_inst_pe_1_0_5_n79) );
  INV_X1 npu_inst_pe_1_0_5_U40 ( .A(npu_inst_pe_1_0_5_n79), .ZN(
        npu_inst_pe_1_0_5_n35) );
  AOI222_X1 npu_inst_pe_1_0_5_U39 ( .A1(npu_inst_int_data_res_1__5__6_), .A2(
        npu_inst_pe_1_0_5_n1), .B1(npu_inst_pe_1_0_5_N79), .B2(
        npu_inst_pe_1_0_5_n76), .C1(npu_inst_pe_1_0_5_N71), .C2(
        npu_inst_pe_1_0_5_n77), .ZN(npu_inst_pe_1_0_5_n78) );
  INV_X1 npu_inst_pe_1_0_5_U38 ( .A(npu_inst_pe_1_0_5_n78), .ZN(
        npu_inst_pe_1_0_5_n34) );
  INV_X1 npu_inst_pe_1_0_5_U37 ( .A(npu_inst_pe_1_0_5_int_data_1_), .ZN(
        npu_inst_pe_1_0_5_n14) );
  AND2_X1 npu_inst_pe_1_0_5_U36 ( .A1(npu_inst_int_data_x_0__5__1_), .A2(
        npu_inst_pe_1_0_5_int_q_weight_1_), .ZN(npu_inst_pe_1_0_5_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_0_5_U35 ( .A1(npu_inst_int_data_x_0__5__0_), .A2(
        npu_inst_pe_1_0_5_int_q_weight_1_), .ZN(npu_inst_pe_1_0_5_int_data_0_)
         );
  AND2_X1 npu_inst_pe_1_0_5_U34 ( .A1(npu_inst_pe_1_0_5_N93), .A2(npu_inst_n60), .ZN(npu_inst_pe_1_0_5_o_data_v_0_) );
  AND2_X1 npu_inst_pe_1_0_5_U33 ( .A1(npu_inst_n60), .A2(npu_inst_pe_1_0_5_N94), .ZN(npu_inst_pe_1_0_5_o_data_v_1_) );
  AOI22_X1 npu_inst_pe_1_0_5_U32 ( .A1(npu_inst_n60), .A2(
        npu_inst_int_data_y_1__5__1_), .B1(npu_inst_pe_1_0_5_n3), .B2(
        npu_inst_int_data_x_0__6__1_), .ZN(npu_inst_pe_1_0_5_n63) );
  AOI22_X1 npu_inst_pe_1_0_5_U31 ( .A1(npu_inst_n60), .A2(
        npu_inst_int_data_y_1__5__0_), .B1(npu_inst_pe_1_0_5_n3), .B2(
        npu_inst_int_data_x_0__6__0_), .ZN(npu_inst_pe_1_0_5_n61) );
  INV_X1 npu_inst_pe_1_0_5_U30 ( .A(npu_inst_pe_1_0_5_int_data_0_), .ZN(
        npu_inst_pe_1_0_5_n13) );
  INV_X1 npu_inst_pe_1_0_5_U29 ( .A(npu_inst_n71), .ZN(npu_inst_pe_1_0_5_n5)
         );
  OR3_X1 npu_inst_pe_1_0_5_U28 ( .A1(npu_inst_pe_1_0_5_n6), .A2(
        npu_inst_pe_1_0_5_n8), .A3(npu_inst_pe_1_0_5_n5), .ZN(
        npu_inst_pe_1_0_5_n56) );
  OR3_X1 npu_inst_pe_1_0_5_U27 ( .A1(npu_inst_pe_1_0_5_n5), .A2(
        npu_inst_pe_1_0_5_n8), .A3(npu_inst_pe_1_0_5_n7), .ZN(
        npu_inst_pe_1_0_5_n48) );
  INV_X1 npu_inst_pe_1_0_5_U26 ( .A(npu_inst_pe_1_0_5_n5), .ZN(
        npu_inst_pe_1_0_5_n4) );
  INV_X1 npu_inst_pe_1_0_5_U25 ( .A(npu_inst_n126), .ZN(npu_inst_pe_1_0_5_n12)
         );
  OR3_X1 npu_inst_pe_1_0_5_U24 ( .A1(npu_inst_pe_1_0_5_n4), .A2(
        npu_inst_pe_1_0_5_n8), .A3(npu_inst_pe_1_0_5_n7), .ZN(
        npu_inst_pe_1_0_5_n52) );
  OR3_X1 npu_inst_pe_1_0_5_U23 ( .A1(npu_inst_pe_1_0_5_n6), .A2(
        npu_inst_pe_1_0_5_n8), .A3(npu_inst_pe_1_0_5_n4), .ZN(
        npu_inst_pe_1_0_5_n60) );
  NOR2_X1 npu_inst_pe_1_0_5_U22 ( .A1(npu_inst_pe_1_0_5_n60), .A2(
        npu_inst_pe_1_0_5_n3), .ZN(npu_inst_pe_1_0_5_n58) );
  NOR2_X1 npu_inst_pe_1_0_5_U21 ( .A1(npu_inst_pe_1_0_5_n56), .A2(
        npu_inst_pe_1_0_5_n3), .ZN(npu_inst_pe_1_0_5_n54) );
  NOR2_X1 npu_inst_pe_1_0_5_U20 ( .A1(npu_inst_pe_1_0_5_n52), .A2(
        npu_inst_pe_1_0_5_n3), .ZN(npu_inst_pe_1_0_5_n50) );
  NOR2_X1 npu_inst_pe_1_0_5_U19 ( .A1(npu_inst_pe_1_0_5_n48), .A2(
        npu_inst_pe_1_0_5_n3), .ZN(npu_inst_pe_1_0_5_n46) );
  NOR2_X1 npu_inst_pe_1_0_5_U18 ( .A1(npu_inst_pe_1_0_5_n40), .A2(
        npu_inst_pe_1_0_5_n3), .ZN(npu_inst_pe_1_0_5_n38) );
  NOR2_X1 npu_inst_pe_1_0_5_U17 ( .A1(npu_inst_pe_1_0_5_n44), .A2(
        npu_inst_pe_1_0_5_n3), .ZN(npu_inst_pe_1_0_5_n42) );
  BUF_X1 npu_inst_pe_1_0_5_U16 ( .A(npu_inst_n106), .Z(npu_inst_pe_1_0_5_n8)
         );
  BUF_X1 npu_inst_pe_1_0_5_U15 ( .A(npu_inst_pe_1_0_5_n12), .Z(
        npu_inst_pe_1_0_5_n11) );
  BUF_X1 npu_inst_pe_1_0_5_U14 ( .A(npu_inst_pe_1_0_5_n12), .Z(
        npu_inst_pe_1_0_5_n10) );
  BUF_X1 npu_inst_pe_1_0_5_U13 ( .A(npu_inst_pe_1_0_5_n12), .Z(
        npu_inst_pe_1_0_5_n9) );
  INV_X1 npu_inst_pe_1_0_5_U12 ( .A(npu_inst_pe_1_0_5_n38), .ZN(
        npu_inst_pe_1_0_5_n118) );
  INV_X1 npu_inst_pe_1_0_5_U11 ( .A(npu_inst_pe_1_0_5_n58), .ZN(
        npu_inst_pe_1_0_5_n114) );
  INV_X1 npu_inst_pe_1_0_5_U10 ( .A(npu_inst_pe_1_0_5_n54), .ZN(
        npu_inst_pe_1_0_5_n115) );
  INV_X1 npu_inst_pe_1_0_5_U9 ( .A(npu_inst_pe_1_0_5_n50), .ZN(
        npu_inst_pe_1_0_5_n116) );
  INV_X1 npu_inst_pe_1_0_5_U8 ( .A(npu_inst_pe_1_0_5_n46), .ZN(
        npu_inst_pe_1_0_5_n117) );
  INV_X1 npu_inst_pe_1_0_5_U7 ( .A(npu_inst_pe_1_0_5_n42), .ZN(
        npu_inst_pe_1_0_5_n119) );
  BUF_X1 npu_inst_pe_1_0_5_U6 ( .A(npu_inst_n36), .Z(npu_inst_pe_1_0_5_n2) );
  BUF_X1 npu_inst_pe_1_0_5_U5 ( .A(npu_inst_n36), .Z(npu_inst_pe_1_0_5_n1) );
  NOR2_X1 npu_inst_pe_1_0_5_U4 ( .A1(npu_inst_pe_1_0_5_int_q_weight_0_), .A2(
        npu_inst_pe_1_0_5_n1), .ZN(npu_inst_pe_1_0_5_n76) );
  NOR2_X1 npu_inst_pe_1_0_5_U3 ( .A1(npu_inst_pe_1_0_5_n27), .A2(
        npu_inst_pe_1_0_5_n1), .ZN(npu_inst_pe_1_0_5_n77) );
  FA_X1 npu_inst_pe_1_0_5_sub_77_U2_1 ( .A(npu_inst_pe_1_0_5_int_q_acc_1_), 
        .B(npu_inst_pe_1_0_5_n14), .CI(npu_inst_pe_1_0_5_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_0_5_sub_77_carry_2_), .S(npu_inst_pe_1_0_5_N66) );
  FA_X1 npu_inst_pe_1_0_5_add_79_U1_1 ( .A(npu_inst_pe_1_0_5_int_q_acc_1_), 
        .B(npu_inst_pe_1_0_5_int_data_1_), .CI(
        npu_inst_pe_1_0_5_add_79_carry_1_), .CO(
        npu_inst_pe_1_0_5_add_79_carry_2_), .S(npu_inst_pe_1_0_5_N74) );
  NAND3_X1 npu_inst_pe_1_0_5_U109 ( .A1(npu_inst_pe_1_0_5_n5), .A2(
        npu_inst_pe_1_0_5_n7), .A3(npu_inst_pe_1_0_5_n8), .ZN(
        npu_inst_pe_1_0_5_n44) );
  NAND3_X1 npu_inst_pe_1_0_5_U108 ( .A1(npu_inst_pe_1_0_5_n4), .A2(
        npu_inst_pe_1_0_5_n7), .A3(npu_inst_pe_1_0_5_n8), .ZN(
        npu_inst_pe_1_0_5_n40) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_0_5_n34), .CK(
        npu_inst_pe_1_0_5_net4178), .RN(npu_inst_pe_1_0_5_n9), .Q(
        npu_inst_pe_1_0_5_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_0_5_n35), .CK(
        npu_inst_pe_1_0_5_net4178), .RN(npu_inst_pe_1_0_5_n9), .Q(
        npu_inst_pe_1_0_5_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_0_5_n36), .CK(
        npu_inst_pe_1_0_5_net4178), .RN(npu_inst_pe_1_0_5_n9), .Q(
        npu_inst_pe_1_0_5_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_0_5_n98), .CK(
        npu_inst_pe_1_0_5_net4178), .RN(npu_inst_pe_1_0_5_n9), .Q(
        npu_inst_pe_1_0_5_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_0_5_n99), .CK(
        npu_inst_pe_1_0_5_net4178), .RN(npu_inst_pe_1_0_5_n9), .Q(
        npu_inst_pe_1_0_5_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_0_5_n100), 
        .CK(npu_inst_pe_1_0_5_net4178), .RN(npu_inst_pe_1_0_5_n9), .Q(
        npu_inst_pe_1_0_5_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_0_5_n33), .CK(
        npu_inst_pe_1_0_5_net4178), .RN(npu_inst_pe_1_0_5_n9), .Q(
        npu_inst_pe_1_0_5_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_0_5_n101), 
        .CK(npu_inst_pe_1_0_5_net4178), .RN(npu_inst_pe_1_0_5_n9), .Q(
        npu_inst_pe_1_0_5_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_weight_reg_0_ ( .D(npu_inst_n112), .CK(
        npu_inst_pe_1_0_5_net4184), .RN(npu_inst_pe_1_0_5_n9), .Q(
        npu_inst_pe_1_0_5_int_q_weight_0_), .QN(npu_inst_pe_1_0_5_n27) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_weight_reg_1_ ( .D(npu_inst_n118), .CK(
        npu_inst_pe_1_0_5_net4184), .RN(npu_inst_pe_1_0_5_n9), .Q(
        npu_inst_pe_1_0_5_int_q_weight_1_), .QN(npu_inst_pe_1_0_5_n26) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_0_5_n113), 
        .CK(npu_inst_pe_1_0_5_net4184), .RN(npu_inst_pe_1_0_5_n9), .Q(
        npu_inst_pe_1_0_5_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_0_5_n107), 
        .CK(npu_inst_pe_1_0_5_net4184), .RN(npu_inst_pe_1_0_5_n9), .Q(
        npu_inst_pe_1_0_5_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_0_5_n112), 
        .CK(npu_inst_pe_1_0_5_net4184), .RN(npu_inst_pe_1_0_5_n10), .Q(
        npu_inst_pe_1_0_5_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_0_5_n106), 
        .CK(npu_inst_pe_1_0_5_net4184), .RN(npu_inst_pe_1_0_5_n10), .Q(
        npu_inst_pe_1_0_5_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_0_5_n111), 
        .CK(npu_inst_pe_1_0_5_net4184), .RN(npu_inst_pe_1_0_5_n10), .Q(
        npu_inst_pe_1_0_5_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_0_5_n105), 
        .CK(npu_inst_pe_1_0_5_net4184), .RN(npu_inst_pe_1_0_5_n10), .Q(
        npu_inst_pe_1_0_5_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_0_5_n110), 
        .CK(npu_inst_pe_1_0_5_net4184), .RN(npu_inst_pe_1_0_5_n10), .Q(
        npu_inst_pe_1_0_5_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_0_5_n104), 
        .CK(npu_inst_pe_1_0_5_net4184), .RN(npu_inst_pe_1_0_5_n10), .Q(
        npu_inst_pe_1_0_5_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_0_5_n109), 
        .CK(npu_inst_pe_1_0_5_net4184), .RN(npu_inst_pe_1_0_5_n10), .Q(
        npu_inst_pe_1_0_5_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_0_5_n103), 
        .CK(npu_inst_pe_1_0_5_net4184), .RN(npu_inst_pe_1_0_5_n10), .Q(
        npu_inst_pe_1_0_5_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_0_5_n108), 
        .CK(npu_inst_pe_1_0_5_net4184), .RN(npu_inst_pe_1_0_5_n10), .Q(
        npu_inst_pe_1_0_5_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_0_5_n102), 
        .CK(npu_inst_pe_1_0_5_net4184), .RN(npu_inst_pe_1_0_5_n10), .Q(
        npu_inst_pe_1_0_5_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_0_5_n86), 
        .CK(npu_inst_pe_1_0_5_net4184), .RN(npu_inst_pe_1_0_5_n10), .Q(
        npu_inst_pe_1_0_5_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_0_5_n87), 
        .CK(npu_inst_pe_1_0_5_net4184), .RN(npu_inst_pe_1_0_5_n10), .Q(
        npu_inst_pe_1_0_5_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_0_5_n88), 
        .CK(npu_inst_pe_1_0_5_net4184), .RN(npu_inst_pe_1_0_5_n11), .Q(
        npu_inst_pe_1_0_5_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_0_5_n89), 
        .CK(npu_inst_pe_1_0_5_net4184), .RN(npu_inst_pe_1_0_5_n11), .Q(
        npu_inst_pe_1_0_5_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_0_5_n90), 
        .CK(npu_inst_pe_1_0_5_net4184), .RN(npu_inst_pe_1_0_5_n11), .Q(
        npu_inst_pe_1_0_5_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_0_5_n91), 
        .CK(npu_inst_pe_1_0_5_net4184), .RN(npu_inst_pe_1_0_5_n11), .Q(
        npu_inst_pe_1_0_5_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_0_5_n92), 
        .CK(npu_inst_pe_1_0_5_net4184), .RN(npu_inst_pe_1_0_5_n11), .Q(
        npu_inst_pe_1_0_5_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_0_5_n93), 
        .CK(npu_inst_pe_1_0_5_net4184), .RN(npu_inst_pe_1_0_5_n11), .Q(
        npu_inst_pe_1_0_5_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_0_5_n94), 
        .CK(npu_inst_pe_1_0_5_net4184), .RN(npu_inst_pe_1_0_5_n11), .Q(
        npu_inst_pe_1_0_5_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_0_5_n95), 
        .CK(npu_inst_pe_1_0_5_net4184), .RN(npu_inst_pe_1_0_5_n11), .Q(
        npu_inst_pe_1_0_5_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_0_5_n96), 
        .CK(npu_inst_pe_1_0_5_net4184), .RN(npu_inst_pe_1_0_5_n11), .Q(
        npu_inst_pe_1_0_5_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_0_5_n97), 
        .CK(npu_inst_pe_1_0_5_net4184), .RN(npu_inst_pe_1_0_5_n11), .Q(
        npu_inst_pe_1_0_5_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_0_5_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_0_5_N84), .SE(1'b0), .GCK(npu_inst_pe_1_0_5_net4178) );
  CLKGATETST_X1 npu_inst_pe_1_0_5_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n66), .SE(1'b0), .GCK(npu_inst_pe_1_0_5_net4184) );
  MUX2_X1 npu_inst_pe_1_0_6_U162 ( .A(npu_inst_pe_1_0_6_n32), .B(
        npu_inst_pe_1_0_6_n29), .S(npu_inst_pe_1_0_6_n8), .Z(
        npu_inst_pe_1_0_6_N93) );
  MUX2_X1 npu_inst_pe_1_0_6_U161 ( .A(npu_inst_pe_1_0_6_n31), .B(
        npu_inst_pe_1_0_6_n30), .S(npu_inst_pe_1_0_6_n6), .Z(
        npu_inst_pe_1_0_6_n32) );
  MUX2_X1 npu_inst_pe_1_0_6_U160 ( .A(npu_inst_pe_1_0_6_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_0_6_int_q_reg_v_1__0_), .S(npu_inst_pe_1_0_6_n4), .Z(
        npu_inst_pe_1_0_6_n31) );
  MUX2_X1 npu_inst_pe_1_0_6_U159 ( .A(npu_inst_pe_1_0_6_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_0_6_int_q_reg_v_3__0_), .S(npu_inst_pe_1_0_6_n4), .Z(
        npu_inst_pe_1_0_6_n30) );
  MUX2_X1 npu_inst_pe_1_0_6_U158 ( .A(npu_inst_pe_1_0_6_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_0_6_int_q_reg_v_5__0_), .S(npu_inst_pe_1_0_6_n4), .Z(
        npu_inst_pe_1_0_6_n29) );
  MUX2_X1 npu_inst_pe_1_0_6_U157 ( .A(npu_inst_pe_1_0_6_n28), .B(
        npu_inst_pe_1_0_6_n23), .S(npu_inst_pe_1_0_6_n8), .Z(
        npu_inst_pe_1_0_6_N94) );
  MUX2_X1 npu_inst_pe_1_0_6_U156 ( .A(npu_inst_pe_1_0_6_n25), .B(
        npu_inst_pe_1_0_6_n24), .S(npu_inst_pe_1_0_6_n6), .Z(
        npu_inst_pe_1_0_6_n28) );
  MUX2_X1 npu_inst_pe_1_0_6_U155 ( .A(npu_inst_pe_1_0_6_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_0_6_int_q_reg_v_1__1_), .S(npu_inst_pe_1_0_6_n4), .Z(
        npu_inst_pe_1_0_6_n25) );
  MUX2_X1 npu_inst_pe_1_0_6_U154 ( .A(npu_inst_pe_1_0_6_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_0_6_int_q_reg_v_3__1_), .S(npu_inst_pe_1_0_6_n4), .Z(
        npu_inst_pe_1_0_6_n24) );
  MUX2_X1 npu_inst_pe_1_0_6_U153 ( .A(npu_inst_pe_1_0_6_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_0_6_int_q_reg_v_5__1_), .S(npu_inst_pe_1_0_6_n4), .Z(
        npu_inst_pe_1_0_6_n23) );
  MUX2_X1 npu_inst_pe_1_0_6_U152 ( .A(npu_inst_pe_1_0_6_n22), .B(
        npu_inst_pe_1_0_6_n19), .S(npu_inst_pe_1_0_6_n8), .Z(
        npu_inst_int_data_x_0__6__1_) );
  MUX2_X1 npu_inst_pe_1_0_6_U151 ( .A(npu_inst_pe_1_0_6_n21), .B(
        npu_inst_pe_1_0_6_n20), .S(npu_inst_pe_1_0_6_n6), .Z(
        npu_inst_pe_1_0_6_n22) );
  MUX2_X1 npu_inst_pe_1_0_6_U150 ( .A(npu_inst_pe_1_0_6_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_0_6_int_q_reg_h_1__1_), .S(npu_inst_pe_1_0_6_n4), .Z(
        npu_inst_pe_1_0_6_n21) );
  MUX2_X1 npu_inst_pe_1_0_6_U149 ( .A(npu_inst_pe_1_0_6_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_0_6_int_q_reg_h_3__1_), .S(npu_inst_pe_1_0_6_n4), .Z(
        npu_inst_pe_1_0_6_n20) );
  MUX2_X1 npu_inst_pe_1_0_6_U148 ( .A(npu_inst_pe_1_0_6_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_0_6_int_q_reg_h_5__1_), .S(npu_inst_pe_1_0_6_n4), .Z(
        npu_inst_pe_1_0_6_n19) );
  MUX2_X1 npu_inst_pe_1_0_6_U147 ( .A(npu_inst_pe_1_0_6_n18), .B(
        npu_inst_pe_1_0_6_n15), .S(npu_inst_pe_1_0_6_n8), .Z(
        npu_inst_int_data_x_0__6__0_) );
  MUX2_X1 npu_inst_pe_1_0_6_U146 ( .A(npu_inst_pe_1_0_6_n17), .B(
        npu_inst_pe_1_0_6_n16), .S(npu_inst_pe_1_0_6_n6), .Z(
        npu_inst_pe_1_0_6_n18) );
  MUX2_X1 npu_inst_pe_1_0_6_U145 ( .A(npu_inst_pe_1_0_6_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_0_6_int_q_reg_h_1__0_), .S(npu_inst_pe_1_0_6_n4), .Z(
        npu_inst_pe_1_0_6_n17) );
  MUX2_X1 npu_inst_pe_1_0_6_U144 ( .A(npu_inst_pe_1_0_6_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_0_6_int_q_reg_h_3__0_), .S(npu_inst_pe_1_0_6_n4), .Z(
        npu_inst_pe_1_0_6_n16) );
  MUX2_X1 npu_inst_pe_1_0_6_U143 ( .A(npu_inst_pe_1_0_6_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_0_6_int_q_reg_h_5__0_), .S(npu_inst_pe_1_0_6_n4), .Z(
        npu_inst_pe_1_0_6_n15) );
  XOR2_X1 npu_inst_pe_1_0_6_U142 ( .A(npu_inst_pe_1_0_6_int_data_0_), .B(
        npu_inst_pe_1_0_6_int_q_acc_0_), .Z(npu_inst_pe_1_0_6_N73) );
  AND2_X1 npu_inst_pe_1_0_6_U141 ( .A1(npu_inst_pe_1_0_6_int_q_acc_0_), .A2(
        npu_inst_pe_1_0_6_int_data_0_), .ZN(npu_inst_pe_1_0_6_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_0_6_U140 ( .A(npu_inst_pe_1_0_6_int_q_acc_0_), .B(
        npu_inst_pe_1_0_6_n13), .ZN(npu_inst_pe_1_0_6_N65) );
  OR2_X1 npu_inst_pe_1_0_6_U139 ( .A1(npu_inst_pe_1_0_6_n13), .A2(
        npu_inst_pe_1_0_6_int_q_acc_0_), .ZN(npu_inst_pe_1_0_6_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_0_6_U138 ( .A(npu_inst_pe_1_0_6_int_q_acc_2_), .B(
        npu_inst_pe_1_0_6_add_79_carry_2_), .Z(npu_inst_pe_1_0_6_N75) );
  AND2_X1 npu_inst_pe_1_0_6_U137 ( .A1(npu_inst_pe_1_0_6_add_79_carry_2_), 
        .A2(npu_inst_pe_1_0_6_int_q_acc_2_), .ZN(
        npu_inst_pe_1_0_6_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_0_6_U136 ( .A(npu_inst_pe_1_0_6_int_q_acc_3_), .B(
        npu_inst_pe_1_0_6_add_79_carry_3_), .Z(npu_inst_pe_1_0_6_N76) );
  AND2_X1 npu_inst_pe_1_0_6_U135 ( .A1(npu_inst_pe_1_0_6_add_79_carry_3_), 
        .A2(npu_inst_pe_1_0_6_int_q_acc_3_), .ZN(
        npu_inst_pe_1_0_6_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_0_6_U134 ( .A(npu_inst_pe_1_0_6_int_q_acc_4_), .B(
        npu_inst_pe_1_0_6_add_79_carry_4_), .Z(npu_inst_pe_1_0_6_N77) );
  AND2_X1 npu_inst_pe_1_0_6_U133 ( .A1(npu_inst_pe_1_0_6_add_79_carry_4_), 
        .A2(npu_inst_pe_1_0_6_int_q_acc_4_), .ZN(
        npu_inst_pe_1_0_6_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_0_6_U132 ( .A(npu_inst_pe_1_0_6_int_q_acc_5_), .B(
        npu_inst_pe_1_0_6_add_79_carry_5_), .Z(npu_inst_pe_1_0_6_N78) );
  AND2_X1 npu_inst_pe_1_0_6_U131 ( .A1(npu_inst_pe_1_0_6_add_79_carry_5_), 
        .A2(npu_inst_pe_1_0_6_int_q_acc_5_), .ZN(
        npu_inst_pe_1_0_6_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_0_6_U130 ( .A(npu_inst_pe_1_0_6_int_q_acc_6_), .B(
        npu_inst_pe_1_0_6_add_79_carry_6_), .Z(npu_inst_pe_1_0_6_N79) );
  AND2_X1 npu_inst_pe_1_0_6_U129 ( .A1(npu_inst_pe_1_0_6_add_79_carry_6_), 
        .A2(npu_inst_pe_1_0_6_int_q_acc_6_), .ZN(
        npu_inst_pe_1_0_6_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_0_6_U128 ( .A(npu_inst_pe_1_0_6_int_q_acc_7_), .B(
        npu_inst_pe_1_0_6_add_79_carry_7_), .Z(npu_inst_pe_1_0_6_N80) );
  XNOR2_X1 npu_inst_pe_1_0_6_U127 ( .A(npu_inst_pe_1_0_6_sub_77_carry_2_), .B(
        npu_inst_pe_1_0_6_int_q_acc_2_), .ZN(npu_inst_pe_1_0_6_N67) );
  OR2_X1 npu_inst_pe_1_0_6_U126 ( .A1(npu_inst_pe_1_0_6_int_q_acc_2_), .A2(
        npu_inst_pe_1_0_6_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_0_6_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_0_6_U125 ( .A(npu_inst_pe_1_0_6_sub_77_carry_3_), .B(
        npu_inst_pe_1_0_6_int_q_acc_3_), .ZN(npu_inst_pe_1_0_6_N68) );
  OR2_X1 npu_inst_pe_1_0_6_U124 ( .A1(npu_inst_pe_1_0_6_int_q_acc_3_), .A2(
        npu_inst_pe_1_0_6_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_0_6_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_0_6_U123 ( .A(npu_inst_pe_1_0_6_sub_77_carry_4_), .B(
        npu_inst_pe_1_0_6_int_q_acc_4_), .ZN(npu_inst_pe_1_0_6_N69) );
  OR2_X1 npu_inst_pe_1_0_6_U122 ( .A1(npu_inst_pe_1_0_6_int_q_acc_4_), .A2(
        npu_inst_pe_1_0_6_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_0_6_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_0_6_U121 ( .A(npu_inst_pe_1_0_6_sub_77_carry_5_), .B(
        npu_inst_pe_1_0_6_int_q_acc_5_), .ZN(npu_inst_pe_1_0_6_N70) );
  OR2_X1 npu_inst_pe_1_0_6_U120 ( .A1(npu_inst_pe_1_0_6_int_q_acc_5_), .A2(
        npu_inst_pe_1_0_6_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_0_6_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_0_6_U119 ( .A(npu_inst_pe_1_0_6_sub_77_carry_6_), .B(
        npu_inst_pe_1_0_6_int_q_acc_6_), .ZN(npu_inst_pe_1_0_6_N71) );
  OR2_X1 npu_inst_pe_1_0_6_U118 ( .A1(npu_inst_pe_1_0_6_int_q_acc_6_), .A2(
        npu_inst_pe_1_0_6_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_0_6_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_0_6_U117 ( .A(npu_inst_pe_1_0_6_int_q_acc_7_), .B(
        npu_inst_pe_1_0_6_sub_77_carry_7_), .ZN(npu_inst_pe_1_0_6_N72) );
  INV_X1 npu_inst_pe_1_0_6_U116 ( .A(npu_inst_n79), .ZN(npu_inst_pe_1_0_6_n7)
         );
  INV_X1 npu_inst_pe_1_0_6_U115 ( .A(npu_inst_pe_1_0_6_n7), .ZN(
        npu_inst_pe_1_0_6_n6) );
  INV_X1 npu_inst_pe_1_0_6_U114 ( .A(npu_inst_n60), .ZN(npu_inst_pe_1_0_6_n3)
         );
  AOI22_X1 npu_inst_pe_1_0_6_U113 ( .A1(npu_inst_int_data_y_1__6__0_), .A2(
        npu_inst_pe_1_0_6_n58), .B1(npu_inst_pe_1_0_6_n114), .B2(
        npu_inst_pe_1_0_6_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_0_6_n57) );
  INV_X1 npu_inst_pe_1_0_6_U112 ( .A(npu_inst_pe_1_0_6_n57), .ZN(
        npu_inst_pe_1_0_6_n108) );
  AOI22_X1 npu_inst_pe_1_0_6_U111 ( .A1(npu_inst_int_data_y_1__6__0_), .A2(
        npu_inst_pe_1_0_6_n54), .B1(npu_inst_pe_1_0_6_n115), .B2(
        npu_inst_pe_1_0_6_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_0_6_n53) );
  INV_X1 npu_inst_pe_1_0_6_U110 ( .A(npu_inst_pe_1_0_6_n53), .ZN(
        npu_inst_pe_1_0_6_n109) );
  AOI22_X1 npu_inst_pe_1_0_6_U107 ( .A1(npu_inst_int_data_y_1__6__0_), .A2(
        npu_inst_pe_1_0_6_n50), .B1(npu_inst_pe_1_0_6_n116), .B2(
        npu_inst_pe_1_0_6_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_0_6_n49) );
  INV_X1 npu_inst_pe_1_0_6_U106 ( .A(npu_inst_pe_1_0_6_n49), .ZN(
        npu_inst_pe_1_0_6_n110) );
  AOI22_X1 npu_inst_pe_1_0_6_U105 ( .A1(npu_inst_int_data_y_1__6__0_), .A2(
        npu_inst_pe_1_0_6_n46), .B1(npu_inst_pe_1_0_6_n117), .B2(
        npu_inst_pe_1_0_6_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_0_6_n45) );
  INV_X1 npu_inst_pe_1_0_6_U104 ( .A(npu_inst_pe_1_0_6_n45), .ZN(
        npu_inst_pe_1_0_6_n111) );
  AOI22_X1 npu_inst_pe_1_0_6_U103 ( .A1(npu_inst_int_data_y_1__6__0_), .A2(
        npu_inst_pe_1_0_6_n42), .B1(npu_inst_pe_1_0_6_n119), .B2(
        npu_inst_pe_1_0_6_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_0_6_n41) );
  INV_X1 npu_inst_pe_1_0_6_U102 ( .A(npu_inst_pe_1_0_6_n41), .ZN(
        npu_inst_pe_1_0_6_n112) );
  AOI22_X1 npu_inst_pe_1_0_6_U101 ( .A1(npu_inst_int_data_y_1__6__1_), .A2(
        npu_inst_pe_1_0_6_n58), .B1(npu_inst_pe_1_0_6_n114), .B2(
        npu_inst_pe_1_0_6_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_0_6_n59) );
  INV_X1 npu_inst_pe_1_0_6_U100 ( .A(npu_inst_pe_1_0_6_n59), .ZN(
        npu_inst_pe_1_0_6_n102) );
  AOI22_X1 npu_inst_pe_1_0_6_U99 ( .A1(npu_inst_int_data_y_1__6__1_), .A2(
        npu_inst_pe_1_0_6_n54), .B1(npu_inst_pe_1_0_6_n115), .B2(
        npu_inst_pe_1_0_6_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_0_6_n55) );
  INV_X1 npu_inst_pe_1_0_6_U98 ( .A(npu_inst_pe_1_0_6_n55), .ZN(
        npu_inst_pe_1_0_6_n103) );
  AOI22_X1 npu_inst_pe_1_0_6_U97 ( .A1(npu_inst_int_data_y_1__6__1_), .A2(
        npu_inst_pe_1_0_6_n50), .B1(npu_inst_pe_1_0_6_n116), .B2(
        npu_inst_pe_1_0_6_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_0_6_n51) );
  INV_X1 npu_inst_pe_1_0_6_U96 ( .A(npu_inst_pe_1_0_6_n51), .ZN(
        npu_inst_pe_1_0_6_n104) );
  AOI22_X1 npu_inst_pe_1_0_6_U95 ( .A1(npu_inst_int_data_y_1__6__1_), .A2(
        npu_inst_pe_1_0_6_n46), .B1(npu_inst_pe_1_0_6_n117), .B2(
        npu_inst_pe_1_0_6_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_0_6_n47) );
  INV_X1 npu_inst_pe_1_0_6_U94 ( .A(npu_inst_pe_1_0_6_n47), .ZN(
        npu_inst_pe_1_0_6_n105) );
  AOI22_X1 npu_inst_pe_1_0_6_U93 ( .A1(npu_inst_int_data_y_1__6__1_), .A2(
        npu_inst_pe_1_0_6_n42), .B1(npu_inst_pe_1_0_6_n119), .B2(
        npu_inst_pe_1_0_6_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_0_6_n43) );
  INV_X1 npu_inst_pe_1_0_6_U92 ( .A(npu_inst_pe_1_0_6_n43), .ZN(
        npu_inst_pe_1_0_6_n106) );
  AOI22_X1 npu_inst_pe_1_0_6_U91 ( .A1(npu_inst_pe_1_0_6_n38), .A2(
        npu_inst_int_data_y_1__6__1_), .B1(npu_inst_pe_1_0_6_n118), .B2(
        npu_inst_pe_1_0_6_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_0_6_n39) );
  INV_X1 npu_inst_pe_1_0_6_U90 ( .A(npu_inst_pe_1_0_6_n39), .ZN(
        npu_inst_pe_1_0_6_n107) );
  AOI22_X1 npu_inst_pe_1_0_6_U89 ( .A1(npu_inst_pe_1_0_6_n38), .A2(
        npu_inst_int_data_y_1__6__0_), .B1(npu_inst_pe_1_0_6_n118), .B2(
        npu_inst_pe_1_0_6_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_0_6_n37) );
  INV_X1 npu_inst_pe_1_0_6_U88 ( .A(npu_inst_pe_1_0_6_n37), .ZN(
        npu_inst_pe_1_0_6_n113) );
  AND2_X1 npu_inst_pe_1_0_6_U87 ( .A1(npu_inst_pe_1_0_6_n2), .A2(
        npu_inst_pe_1_0_6_int_q_acc_7_), .ZN(o_data[15]) );
  AND2_X1 npu_inst_pe_1_0_6_U86 ( .A1(npu_inst_pe_1_0_6_int_q_acc_6_), .A2(
        npu_inst_pe_1_0_6_n2), .ZN(o_data[14]) );
  AND2_X1 npu_inst_pe_1_0_6_U85 ( .A1(npu_inst_pe_1_0_6_int_q_acc_5_), .A2(
        npu_inst_pe_1_0_6_n2), .ZN(o_data[13]) );
  AND2_X1 npu_inst_pe_1_0_6_U84 ( .A1(npu_inst_pe_1_0_6_int_q_acc_4_), .A2(
        npu_inst_pe_1_0_6_n2), .ZN(o_data[12]) );
  AND2_X1 npu_inst_pe_1_0_6_U83 ( .A1(npu_inst_pe_1_0_6_int_q_acc_3_), .A2(
        npu_inst_pe_1_0_6_n2), .ZN(o_data[11]) );
  NAND2_X1 npu_inst_pe_1_0_6_U82 ( .A1(npu_inst_pe_1_0_6_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_0_6_n60), .ZN(npu_inst_pe_1_0_6_n74) );
  OAI21_X1 npu_inst_pe_1_0_6_U81 ( .B1(npu_inst_pe_1_0_6_n63), .B2(
        npu_inst_pe_1_0_6_n60), .A(npu_inst_pe_1_0_6_n74), .ZN(
        npu_inst_pe_1_0_6_n97) );
  NAND2_X1 npu_inst_pe_1_0_6_U80 ( .A1(npu_inst_pe_1_0_6_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_0_6_n60), .ZN(npu_inst_pe_1_0_6_n73) );
  OAI21_X1 npu_inst_pe_1_0_6_U79 ( .B1(npu_inst_pe_1_0_6_n61), .B2(
        npu_inst_pe_1_0_6_n60), .A(npu_inst_pe_1_0_6_n73), .ZN(
        npu_inst_pe_1_0_6_n96) );
  NAND2_X1 npu_inst_pe_1_0_6_U78 ( .A1(npu_inst_pe_1_0_6_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_0_6_n56), .ZN(npu_inst_pe_1_0_6_n72) );
  OAI21_X1 npu_inst_pe_1_0_6_U77 ( .B1(npu_inst_pe_1_0_6_n63), .B2(
        npu_inst_pe_1_0_6_n56), .A(npu_inst_pe_1_0_6_n72), .ZN(
        npu_inst_pe_1_0_6_n95) );
  NAND2_X1 npu_inst_pe_1_0_6_U76 ( .A1(npu_inst_pe_1_0_6_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_0_6_n56), .ZN(npu_inst_pe_1_0_6_n71) );
  OAI21_X1 npu_inst_pe_1_0_6_U75 ( .B1(npu_inst_pe_1_0_6_n61), .B2(
        npu_inst_pe_1_0_6_n56), .A(npu_inst_pe_1_0_6_n71), .ZN(
        npu_inst_pe_1_0_6_n94) );
  NAND2_X1 npu_inst_pe_1_0_6_U74 ( .A1(npu_inst_pe_1_0_6_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_0_6_n52), .ZN(npu_inst_pe_1_0_6_n70) );
  OAI21_X1 npu_inst_pe_1_0_6_U73 ( .B1(npu_inst_pe_1_0_6_n63), .B2(
        npu_inst_pe_1_0_6_n52), .A(npu_inst_pe_1_0_6_n70), .ZN(
        npu_inst_pe_1_0_6_n93) );
  NAND2_X1 npu_inst_pe_1_0_6_U72 ( .A1(npu_inst_pe_1_0_6_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_0_6_n52), .ZN(npu_inst_pe_1_0_6_n69) );
  OAI21_X1 npu_inst_pe_1_0_6_U71 ( .B1(npu_inst_pe_1_0_6_n61), .B2(
        npu_inst_pe_1_0_6_n52), .A(npu_inst_pe_1_0_6_n69), .ZN(
        npu_inst_pe_1_0_6_n92) );
  NAND2_X1 npu_inst_pe_1_0_6_U70 ( .A1(npu_inst_pe_1_0_6_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_0_6_n48), .ZN(npu_inst_pe_1_0_6_n68) );
  OAI21_X1 npu_inst_pe_1_0_6_U69 ( .B1(npu_inst_pe_1_0_6_n63), .B2(
        npu_inst_pe_1_0_6_n48), .A(npu_inst_pe_1_0_6_n68), .ZN(
        npu_inst_pe_1_0_6_n91) );
  NAND2_X1 npu_inst_pe_1_0_6_U68 ( .A1(npu_inst_pe_1_0_6_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_0_6_n48), .ZN(npu_inst_pe_1_0_6_n67) );
  OAI21_X1 npu_inst_pe_1_0_6_U67 ( .B1(npu_inst_pe_1_0_6_n61), .B2(
        npu_inst_pe_1_0_6_n48), .A(npu_inst_pe_1_0_6_n67), .ZN(
        npu_inst_pe_1_0_6_n90) );
  NAND2_X1 npu_inst_pe_1_0_6_U66 ( .A1(npu_inst_pe_1_0_6_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_0_6_n44), .ZN(npu_inst_pe_1_0_6_n66) );
  OAI21_X1 npu_inst_pe_1_0_6_U65 ( .B1(npu_inst_pe_1_0_6_n63), .B2(
        npu_inst_pe_1_0_6_n44), .A(npu_inst_pe_1_0_6_n66), .ZN(
        npu_inst_pe_1_0_6_n89) );
  NAND2_X1 npu_inst_pe_1_0_6_U64 ( .A1(npu_inst_pe_1_0_6_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_0_6_n44), .ZN(npu_inst_pe_1_0_6_n65) );
  OAI21_X1 npu_inst_pe_1_0_6_U63 ( .B1(npu_inst_pe_1_0_6_n61), .B2(
        npu_inst_pe_1_0_6_n44), .A(npu_inst_pe_1_0_6_n65), .ZN(
        npu_inst_pe_1_0_6_n88) );
  NAND2_X1 npu_inst_pe_1_0_6_U62 ( .A1(npu_inst_pe_1_0_6_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_0_6_n40), .ZN(npu_inst_pe_1_0_6_n64) );
  OAI21_X1 npu_inst_pe_1_0_6_U61 ( .B1(npu_inst_pe_1_0_6_n63), .B2(
        npu_inst_pe_1_0_6_n40), .A(npu_inst_pe_1_0_6_n64), .ZN(
        npu_inst_pe_1_0_6_n87) );
  NAND2_X1 npu_inst_pe_1_0_6_U60 ( .A1(npu_inst_pe_1_0_6_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_0_6_n40), .ZN(npu_inst_pe_1_0_6_n62) );
  OAI21_X1 npu_inst_pe_1_0_6_U59 ( .B1(npu_inst_pe_1_0_6_n61), .B2(
        npu_inst_pe_1_0_6_n40), .A(npu_inst_pe_1_0_6_n62), .ZN(
        npu_inst_pe_1_0_6_n86) );
  NOR3_X1 npu_inst_pe_1_0_6_U58 ( .A1(npu_inst_pe_1_0_6_n26), .A2(npu_inst_n60), .A3(npu_inst_int_ckg[57]), .ZN(npu_inst_pe_1_0_6_n85) );
  OR2_X1 npu_inst_pe_1_0_6_U57 ( .A1(npu_inst_pe_1_0_6_n85), .A2(
        npu_inst_pe_1_0_6_n2), .ZN(npu_inst_pe_1_0_6_N84) );
  AND2_X1 npu_inst_pe_1_0_6_U56 ( .A1(npu_inst_pe_1_0_6_int_q_acc_0_), .A2(
        npu_inst_pe_1_0_6_n1), .ZN(o_data[8]) );
  AND2_X1 npu_inst_pe_1_0_6_U55 ( .A1(npu_inst_pe_1_0_6_int_q_acc_1_), .A2(
        npu_inst_pe_1_0_6_n1), .ZN(o_data[9]) );
  AND2_X1 npu_inst_pe_1_0_6_U54 ( .A1(npu_inst_pe_1_0_6_int_q_acc_2_), .A2(
        npu_inst_pe_1_0_6_n1), .ZN(o_data[10]) );
  AOI222_X1 npu_inst_pe_1_0_6_U53 ( .A1(npu_inst_int_data_res_1__6__0_), .A2(
        npu_inst_pe_1_0_6_n1), .B1(npu_inst_pe_1_0_6_N73), .B2(
        npu_inst_pe_1_0_6_n76), .C1(npu_inst_pe_1_0_6_N65), .C2(
        npu_inst_pe_1_0_6_n77), .ZN(npu_inst_pe_1_0_6_n84) );
  INV_X1 npu_inst_pe_1_0_6_U52 ( .A(npu_inst_pe_1_0_6_n84), .ZN(
        npu_inst_pe_1_0_6_n101) );
  AOI222_X1 npu_inst_pe_1_0_6_U51 ( .A1(npu_inst_int_data_res_1__6__7_), .A2(
        npu_inst_pe_1_0_6_n1), .B1(npu_inst_pe_1_0_6_N80), .B2(
        npu_inst_pe_1_0_6_n76), .C1(npu_inst_pe_1_0_6_N72), .C2(
        npu_inst_pe_1_0_6_n77), .ZN(npu_inst_pe_1_0_6_n75) );
  INV_X1 npu_inst_pe_1_0_6_U50 ( .A(npu_inst_pe_1_0_6_n75), .ZN(
        npu_inst_pe_1_0_6_n33) );
  AOI222_X1 npu_inst_pe_1_0_6_U49 ( .A1(npu_inst_int_data_res_1__6__1_), .A2(
        npu_inst_pe_1_0_6_n1), .B1(npu_inst_pe_1_0_6_N74), .B2(
        npu_inst_pe_1_0_6_n76), .C1(npu_inst_pe_1_0_6_N66), .C2(
        npu_inst_pe_1_0_6_n77), .ZN(npu_inst_pe_1_0_6_n83) );
  INV_X1 npu_inst_pe_1_0_6_U48 ( .A(npu_inst_pe_1_0_6_n83), .ZN(
        npu_inst_pe_1_0_6_n100) );
  AOI222_X1 npu_inst_pe_1_0_6_U47 ( .A1(npu_inst_int_data_res_1__6__2_), .A2(
        npu_inst_pe_1_0_6_n1), .B1(npu_inst_pe_1_0_6_N75), .B2(
        npu_inst_pe_1_0_6_n76), .C1(npu_inst_pe_1_0_6_N67), .C2(
        npu_inst_pe_1_0_6_n77), .ZN(npu_inst_pe_1_0_6_n82) );
  INV_X1 npu_inst_pe_1_0_6_U46 ( .A(npu_inst_pe_1_0_6_n82), .ZN(
        npu_inst_pe_1_0_6_n99) );
  AOI222_X1 npu_inst_pe_1_0_6_U45 ( .A1(npu_inst_int_data_res_1__6__3_), .A2(
        npu_inst_pe_1_0_6_n1), .B1(npu_inst_pe_1_0_6_N76), .B2(
        npu_inst_pe_1_0_6_n76), .C1(npu_inst_pe_1_0_6_N68), .C2(
        npu_inst_pe_1_0_6_n77), .ZN(npu_inst_pe_1_0_6_n81) );
  INV_X1 npu_inst_pe_1_0_6_U44 ( .A(npu_inst_pe_1_0_6_n81), .ZN(
        npu_inst_pe_1_0_6_n98) );
  AOI222_X1 npu_inst_pe_1_0_6_U43 ( .A1(npu_inst_int_data_res_1__6__4_), .A2(
        npu_inst_pe_1_0_6_n1), .B1(npu_inst_pe_1_0_6_N77), .B2(
        npu_inst_pe_1_0_6_n76), .C1(npu_inst_pe_1_0_6_N69), .C2(
        npu_inst_pe_1_0_6_n77), .ZN(npu_inst_pe_1_0_6_n80) );
  INV_X1 npu_inst_pe_1_0_6_U42 ( .A(npu_inst_pe_1_0_6_n80), .ZN(
        npu_inst_pe_1_0_6_n36) );
  AOI222_X1 npu_inst_pe_1_0_6_U41 ( .A1(npu_inst_int_data_res_1__6__5_), .A2(
        npu_inst_pe_1_0_6_n1), .B1(npu_inst_pe_1_0_6_N78), .B2(
        npu_inst_pe_1_0_6_n76), .C1(npu_inst_pe_1_0_6_N70), .C2(
        npu_inst_pe_1_0_6_n77), .ZN(npu_inst_pe_1_0_6_n79) );
  INV_X1 npu_inst_pe_1_0_6_U40 ( .A(npu_inst_pe_1_0_6_n79), .ZN(
        npu_inst_pe_1_0_6_n35) );
  AOI222_X1 npu_inst_pe_1_0_6_U39 ( .A1(npu_inst_int_data_res_1__6__6_), .A2(
        npu_inst_pe_1_0_6_n1), .B1(npu_inst_pe_1_0_6_N79), .B2(
        npu_inst_pe_1_0_6_n76), .C1(npu_inst_pe_1_0_6_N71), .C2(
        npu_inst_pe_1_0_6_n77), .ZN(npu_inst_pe_1_0_6_n78) );
  INV_X1 npu_inst_pe_1_0_6_U38 ( .A(npu_inst_pe_1_0_6_n78), .ZN(
        npu_inst_pe_1_0_6_n34) );
  INV_X1 npu_inst_pe_1_0_6_U37 ( .A(npu_inst_pe_1_0_6_int_data_1_), .ZN(
        npu_inst_pe_1_0_6_n14) );
  AND2_X1 npu_inst_pe_1_0_6_U36 ( .A1(npu_inst_int_data_x_0__6__1_), .A2(
        npu_inst_pe_1_0_6_int_q_weight_1_), .ZN(npu_inst_pe_1_0_6_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_0_6_U35 ( .A1(npu_inst_int_data_x_0__6__0_), .A2(
        npu_inst_pe_1_0_6_int_q_weight_1_), .ZN(npu_inst_pe_1_0_6_int_data_0_)
         );
  AND2_X1 npu_inst_pe_1_0_6_U34 ( .A1(npu_inst_pe_1_0_6_N93), .A2(npu_inst_n60), .ZN(npu_inst_pe_1_0_6_o_data_v_0_) );
  AND2_X1 npu_inst_pe_1_0_6_U33 ( .A1(npu_inst_n60), .A2(npu_inst_pe_1_0_6_N94), .ZN(npu_inst_pe_1_0_6_o_data_v_1_) );
  AOI22_X1 npu_inst_pe_1_0_6_U32 ( .A1(npu_inst_n60), .A2(
        npu_inst_int_data_y_1__6__1_), .B1(npu_inst_pe_1_0_6_n3), .B2(
        npu_inst_int_data_x_0__7__1_), .ZN(npu_inst_pe_1_0_6_n63) );
  AOI22_X1 npu_inst_pe_1_0_6_U31 ( .A1(npu_inst_n60), .A2(
        npu_inst_int_data_y_1__6__0_), .B1(npu_inst_pe_1_0_6_n3), .B2(
        npu_inst_int_data_x_0__7__0_), .ZN(npu_inst_pe_1_0_6_n61) );
  INV_X1 npu_inst_pe_1_0_6_U30 ( .A(npu_inst_pe_1_0_6_int_data_0_), .ZN(
        npu_inst_pe_1_0_6_n13) );
  INV_X1 npu_inst_pe_1_0_6_U29 ( .A(npu_inst_n71), .ZN(npu_inst_pe_1_0_6_n5)
         );
  OR3_X1 npu_inst_pe_1_0_6_U28 ( .A1(npu_inst_pe_1_0_6_n6), .A2(
        npu_inst_pe_1_0_6_n8), .A3(npu_inst_pe_1_0_6_n5), .ZN(
        npu_inst_pe_1_0_6_n56) );
  OR3_X1 npu_inst_pe_1_0_6_U27 ( .A1(npu_inst_pe_1_0_6_n5), .A2(
        npu_inst_pe_1_0_6_n8), .A3(npu_inst_pe_1_0_6_n7), .ZN(
        npu_inst_pe_1_0_6_n48) );
  INV_X1 npu_inst_pe_1_0_6_U26 ( .A(npu_inst_pe_1_0_6_n5), .ZN(
        npu_inst_pe_1_0_6_n4) );
  INV_X1 npu_inst_pe_1_0_6_U25 ( .A(npu_inst_n126), .ZN(npu_inst_pe_1_0_6_n12)
         );
  OR3_X1 npu_inst_pe_1_0_6_U24 ( .A1(npu_inst_pe_1_0_6_n4), .A2(
        npu_inst_pe_1_0_6_n8), .A3(npu_inst_pe_1_0_6_n7), .ZN(
        npu_inst_pe_1_0_6_n52) );
  OR3_X1 npu_inst_pe_1_0_6_U23 ( .A1(npu_inst_pe_1_0_6_n6), .A2(
        npu_inst_pe_1_0_6_n8), .A3(npu_inst_pe_1_0_6_n4), .ZN(
        npu_inst_pe_1_0_6_n60) );
  NOR2_X1 npu_inst_pe_1_0_6_U22 ( .A1(npu_inst_pe_1_0_6_n60), .A2(
        npu_inst_pe_1_0_6_n3), .ZN(npu_inst_pe_1_0_6_n58) );
  NOR2_X1 npu_inst_pe_1_0_6_U21 ( .A1(npu_inst_pe_1_0_6_n56), .A2(
        npu_inst_pe_1_0_6_n3), .ZN(npu_inst_pe_1_0_6_n54) );
  NOR2_X1 npu_inst_pe_1_0_6_U20 ( .A1(npu_inst_pe_1_0_6_n52), .A2(
        npu_inst_pe_1_0_6_n3), .ZN(npu_inst_pe_1_0_6_n50) );
  NOR2_X1 npu_inst_pe_1_0_6_U19 ( .A1(npu_inst_pe_1_0_6_n48), .A2(
        npu_inst_pe_1_0_6_n3), .ZN(npu_inst_pe_1_0_6_n46) );
  NOR2_X1 npu_inst_pe_1_0_6_U18 ( .A1(npu_inst_pe_1_0_6_n40), .A2(
        npu_inst_pe_1_0_6_n3), .ZN(npu_inst_pe_1_0_6_n38) );
  NOR2_X1 npu_inst_pe_1_0_6_U17 ( .A1(npu_inst_pe_1_0_6_n44), .A2(
        npu_inst_pe_1_0_6_n3), .ZN(npu_inst_pe_1_0_6_n42) );
  BUF_X1 npu_inst_pe_1_0_6_U16 ( .A(npu_inst_n106), .Z(npu_inst_pe_1_0_6_n8)
         );
  BUF_X1 npu_inst_pe_1_0_6_U15 ( .A(npu_inst_pe_1_0_6_n12), .Z(
        npu_inst_pe_1_0_6_n11) );
  BUF_X1 npu_inst_pe_1_0_6_U14 ( .A(npu_inst_pe_1_0_6_n12), .Z(
        npu_inst_pe_1_0_6_n10) );
  BUF_X1 npu_inst_pe_1_0_6_U13 ( .A(npu_inst_pe_1_0_6_n12), .Z(
        npu_inst_pe_1_0_6_n9) );
  INV_X1 npu_inst_pe_1_0_6_U12 ( .A(npu_inst_pe_1_0_6_n38), .ZN(
        npu_inst_pe_1_0_6_n118) );
  INV_X1 npu_inst_pe_1_0_6_U11 ( .A(npu_inst_pe_1_0_6_n58), .ZN(
        npu_inst_pe_1_0_6_n114) );
  INV_X1 npu_inst_pe_1_0_6_U10 ( .A(npu_inst_pe_1_0_6_n54), .ZN(
        npu_inst_pe_1_0_6_n115) );
  INV_X1 npu_inst_pe_1_0_6_U9 ( .A(npu_inst_pe_1_0_6_n50), .ZN(
        npu_inst_pe_1_0_6_n116) );
  INV_X1 npu_inst_pe_1_0_6_U8 ( .A(npu_inst_pe_1_0_6_n46), .ZN(
        npu_inst_pe_1_0_6_n117) );
  INV_X1 npu_inst_pe_1_0_6_U7 ( .A(npu_inst_pe_1_0_6_n42), .ZN(
        npu_inst_pe_1_0_6_n119) );
  BUF_X1 npu_inst_pe_1_0_6_U6 ( .A(npu_inst_n35), .Z(npu_inst_pe_1_0_6_n2) );
  BUF_X1 npu_inst_pe_1_0_6_U5 ( .A(npu_inst_n35), .Z(npu_inst_pe_1_0_6_n1) );
  NOR2_X1 npu_inst_pe_1_0_6_U4 ( .A1(npu_inst_pe_1_0_6_int_q_weight_0_), .A2(
        npu_inst_pe_1_0_6_n1), .ZN(npu_inst_pe_1_0_6_n76) );
  NOR2_X1 npu_inst_pe_1_0_6_U3 ( .A1(npu_inst_pe_1_0_6_n27), .A2(
        npu_inst_pe_1_0_6_n1), .ZN(npu_inst_pe_1_0_6_n77) );
  FA_X1 npu_inst_pe_1_0_6_sub_77_U2_1 ( .A(npu_inst_pe_1_0_6_int_q_acc_1_), 
        .B(npu_inst_pe_1_0_6_n14), .CI(npu_inst_pe_1_0_6_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_0_6_sub_77_carry_2_), .S(npu_inst_pe_1_0_6_N66) );
  FA_X1 npu_inst_pe_1_0_6_add_79_U1_1 ( .A(npu_inst_pe_1_0_6_int_q_acc_1_), 
        .B(npu_inst_pe_1_0_6_int_data_1_), .CI(
        npu_inst_pe_1_0_6_add_79_carry_1_), .CO(
        npu_inst_pe_1_0_6_add_79_carry_2_), .S(npu_inst_pe_1_0_6_N74) );
  NAND3_X1 npu_inst_pe_1_0_6_U109 ( .A1(npu_inst_pe_1_0_6_n5), .A2(
        npu_inst_pe_1_0_6_n7), .A3(npu_inst_pe_1_0_6_n8), .ZN(
        npu_inst_pe_1_0_6_n44) );
  NAND3_X1 npu_inst_pe_1_0_6_U108 ( .A1(npu_inst_pe_1_0_6_n4), .A2(
        npu_inst_pe_1_0_6_n7), .A3(npu_inst_pe_1_0_6_n8), .ZN(
        npu_inst_pe_1_0_6_n40) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_0_6_n34), .CK(
        npu_inst_pe_1_0_6_net4155), .RN(npu_inst_pe_1_0_6_n9), .Q(
        npu_inst_pe_1_0_6_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_0_6_n35), .CK(
        npu_inst_pe_1_0_6_net4155), .RN(npu_inst_pe_1_0_6_n9), .Q(
        npu_inst_pe_1_0_6_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_0_6_n36), .CK(
        npu_inst_pe_1_0_6_net4155), .RN(npu_inst_pe_1_0_6_n9), .Q(
        npu_inst_pe_1_0_6_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_0_6_n98), .CK(
        npu_inst_pe_1_0_6_net4155), .RN(npu_inst_pe_1_0_6_n9), .Q(
        npu_inst_pe_1_0_6_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_0_6_n99), .CK(
        npu_inst_pe_1_0_6_net4155), .RN(npu_inst_pe_1_0_6_n9), .Q(
        npu_inst_pe_1_0_6_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_0_6_n100), 
        .CK(npu_inst_pe_1_0_6_net4155), .RN(npu_inst_pe_1_0_6_n9), .Q(
        npu_inst_pe_1_0_6_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_0_6_n33), .CK(
        npu_inst_pe_1_0_6_net4155), .RN(npu_inst_pe_1_0_6_n9), .Q(
        npu_inst_pe_1_0_6_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_0_6_n101), 
        .CK(npu_inst_pe_1_0_6_net4155), .RN(npu_inst_pe_1_0_6_n9), .Q(
        npu_inst_pe_1_0_6_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_weight_reg_0_ ( .D(npu_inst_n112), .CK(
        npu_inst_pe_1_0_6_net4161), .RN(npu_inst_pe_1_0_6_n9), .Q(
        npu_inst_pe_1_0_6_int_q_weight_0_), .QN(npu_inst_pe_1_0_6_n27) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_weight_reg_1_ ( .D(npu_inst_n118), .CK(
        npu_inst_pe_1_0_6_net4161), .RN(npu_inst_pe_1_0_6_n9), .Q(
        npu_inst_pe_1_0_6_int_q_weight_1_), .QN(npu_inst_pe_1_0_6_n26) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_0_6_n113), 
        .CK(npu_inst_pe_1_0_6_net4161), .RN(npu_inst_pe_1_0_6_n9), .Q(
        npu_inst_pe_1_0_6_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_0_6_n107), 
        .CK(npu_inst_pe_1_0_6_net4161), .RN(npu_inst_pe_1_0_6_n9), .Q(
        npu_inst_pe_1_0_6_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_0_6_n112), 
        .CK(npu_inst_pe_1_0_6_net4161), .RN(npu_inst_pe_1_0_6_n10), .Q(
        npu_inst_pe_1_0_6_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_0_6_n106), 
        .CK(npu_inst_pe_1_0_6_net4161), .RN(npu_inst_pe_1_0_6_n10), .Q(
        npu_inst_pe_1_0_6_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_0_6_n111), 
        .CK(npu_inst_pe_1_0_6_net4161), .RN(npu_inst_pe_1_0_6_n10), .Q(
        npu_inst_pe_1_0_6_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_0_6_n105), 
        .CK(npu_inst_pe_1_0_6_net4161), .RN(npu_inst_pe_1_0_6_n10), .Q(
        npu_inst_pe_1_0_6_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_0_6_n110), 
        .CK(npu_inst_pe_1_0_6_net4161), .RN(npu_inst_pe_1_0_6_n10), .Q(
        npu_inst_pe_1_0_6_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_0_6_n104), 
        .CK(npu_inst_pe_1_0_6_net4161), .RN(npu_inst_pe_1_0_6_n10), .Q(
        npu_inst_pe_1_0_6_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_0_6_n109), 
        .CK(npu_inst_pe_1_0_6_net4161), .RN(npu_inst_pe_1_0_6_n10), .Q(
        npu_inst_pe_1_0_6_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_0_6_n103), 
        .CK(npu_inst_pe_1_0_6_net4161), .RN(npu_inst_pe_1_0_6_n10), .Q(
        npu_inst_pe_1_0_6_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_0_6_n108), 
        .CK(npu_inst_pe_1_0_6_net4161), .RN(npu_inst_pe_1_0_6_n10), .Q(
        npu_inst_pe_1_0_6_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_0_6_n102), 
        .CK(npu_inst_pe_1_0_6_net4161), .RN(npu_inst_pe_1_0_6_n10), .Q(
        npu_inst_pe_1_0_6_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_0_6_n86), 
        .CK(npu_inst_pe_1_0_6_net4161), .RN(npu_inst_pe_1_0_6_n10), .Q(
        npu_inst_pe_1_0_6_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_0_6_n87), 
        .CK(npu_inst_pe_1_0_6_net4161), .RN(npu_inst_pe_1_0_6_n10), .Q(
        npu_inst_pe_1_0_6_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_0_6_n88), 
        .CK(npu_inst_pe_1_0_6_net4161), .RN(npu_inst_pe_1_0_6_n11), .Q(
        npu_inst_pe_1_0_6_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_0_6_n89), 
        .CK(npu_inst_pe_1_0_6_net4161), .RN(npu_inst_pe_1_0_6_n11), .Q(
        npu_inst_pe_1_0_6_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_0_6_n90), 
        .CK(npu_inst_pe_1_0_6_net4161), .RN(npu_inst_pe_1_0_6_n11), .Q(
        npu_inst_pe_1_0_6_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_0_6_n91), 
        .CK(npu_inst_pe_1_0_6_net4161), .RN(npu_inst_pe_1_0_6_n11), .Q(
        npu_inst_pe_1_0_6_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_0_6_n92), 
        .CK(npu_inst_pe_1_0_6_net4161), .RN(npu_inst_pe_1_0_6_n11), .Q(
        npu_inst_pe_1_0_6_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_0_6_n93), 
        .CK(npu_inst_pe_1_0_6_net4161), .RN(npu_inst_pe_1_0_6_n11), .Q(
        npu_inst_pe_1_0_6_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_0_6_n94), 
        .CK(npu_inst_pe_1_0_6_net4161), .RN(npu_inst_pe_1_0_6_n11), .Q(
        npu_inst_pe_1_0_6_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_0_6_n95), 
        .CK(npu_inst_pe_1_0_6_net4161), .RN(npu_inst_pe_1_0_6_n11), .Q(
        npu_inst_pe_1_0_6_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_0_6_n96), 
        .CK(npu_inst_pe_1_0_6_net4161), .RN(npu_inst_pe_1_0_6_n11), .Q(
        npu_inst_pe_1_0_6_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_0_6_n97), 
        .CK(npu_inst_pe_1_0_6_net4161), .RN(npu_inst_pe_1_0_6_n11), .Q(
        npu_inst_pe_1_0_6_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_0_6_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_0_6_N84), .SE(1'b0), .GCK(npu_inst_pe_1_0_6_net4155) );
  CLKGATETST_X1 npu_inst_pe_1_0_6_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n66), .SE(1'b0), .GCK(npu_inst_pe_1_0_6_net4161) );
  MUX2_X1 npu_inst_pe_1_0_7_U162 ( .A(npu_inst_pe_1_0_7_n32), .B(
        npu_inst_pe_1_0_7_n29), .S(npu_inst_pe_1_0_7_n8), .Z(
        npu_inst_pe_1_0_7_N93) );
  MUX2_X1 npu_inst_pe_1_0_7_U161 ( .A(npu_inst_pe_1_0_7_n31), .B(
        npu_inst_pe_1_0_7_n30), .S(npu_inst_pe_1_0_7_n6), .Z(
        npu_inst_pe_1_0_7_n32) );
  MUX2_X1 npu_inst_pe_1_0_7_U160 ( .A(npu_inst_pe_1_0_7_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_0_7_int_q_reg_v_1__0_), .S(npu_inst_pe_1_0_7_n4), .Z(
        npu_inst_pe_1_0_7_n31) );
  MUX2_X1 npu_inst_pe_1_0_7_U159 ( .A(npu_inst_pe_1_0_7_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_0_7_int_q_reg_v_3__0_), .S(npu_inst_pe_1_0_7_n4), .Z(
        npu_inst_pe_1_0_7_n30) );
  MUX2_X1 npu_inst_pe_1_0_7_U158 ( .A(npu_inst_pe_1_0_7_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_0_7_int_q_reg_v_5__0_), .S(npu_inst_pe_1_0_7_n4), .Z(
        npu_inst_pe_1_0_7_n29) );
  MUX2_X1 npu_inst_pe_1_0_7_U157 ( .A(npu_inst_pe_1_0_7_n28), .B(
        npu_inst_pe_1_0_7_n23), .S(npu_inst_pe_1_0_7_n8), .Z(
        npu_inst_pe_1_0_7_N94) );
  MUX2_X1 npu_inst_pe_1_0_7_U156 ( .A(npu_inst_pe_1_0_7_n25), .B(
        npu_inst_pe_1_0_7_n24), .S(npu_inst_pe_1_0_7_n6), .Z(
        npu_inst_pe_1_0_7_n28) );
  MUX2_X1 npu_inst_pe_1_0_7_U155 ( .A(npu_inst_pe_1_0_7_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_0_7_int_q_reg_v_1__1_), .S(npu_inst_pe_1_0_7_n4), .Z(
        npu_inst_pe_1_0_7_n25) );
  MUX2_X1 npu_inst_pe_1_0_7_U154 ( .A(npu_inst_pe_1_0_7_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_0_7_int_q_reg_v_3__1_), .S(npu_inst_pe_1_0_7_n4), .Z(
        npu_inst_pe_1_0_7_n24) );
  MUX2_X1 npu_inst_pe_1_0_7_U153 ( .A(npu_inst_pe_1_0_7_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_0_7_int_q_reg_v_5__1_), .S(npu_inst_pe_1_0_7_n4), .Z(
        npu_inst_pe_1_0_7_n23) );
  MUX2_X1 npu_inst_pe_1_0_7_U152 ( .A(npu_inst_pe_1_0_7_n22), .B(
        npu_inst_pe_1_0_7_n19), .S(npu_inst_pe_1_0_7_n8), .Z(
        npu_inst_int_data_x_0__7__1_) );
  MUX2_X1 npu_inst_pe_1_0_7_U151 ( .A(npu_inst_pe_1_0_7_n21), .B(
        npu_inst_pe_1_0_7_n20), .S(npu_inst_pe_1_0_7_n6), .Z(
        npu_inst_pe_1_0_7_n22) );
  MUX2_X1 npu_inst_pe_1_0_7_U150 ( .A(npu_inst_pe_1_0_7_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_0_7_int_q_reg_h_1__1_), .S(npu_inst_pe_1_0_7_n4), .Z(
        npu_inst_pe_1_0_7_n21) );
  MUX2_X1 npu_inst_pe_1_0_7_U149 ( .A(npu_inst_pe_1_0_7_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_0_7_int_q_reg_h_3__1_), .S(npu_inst_pe_1_0_7_n4), .Z(
        npu_inst_pe_1_0_7_n20) );
  MUX2_X1 npu_inst_pe_1_0_7_U148 ( .A(npu_inst_pe_1_0_7_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_0_7_int_q_reg_h_5__1_), .S(npu_inst_pe_1_0_7_n4), .Z(
        npu_inst_pe_1_0_7_n19) );
  MUX2_X1 npu_inst_pe_1_0_7_U147 ( .A(npu_inst_pe_1_0_7_n18), .B(
        npu_inst_pe_1_0_7_n15), .S(npu_inst_pe_1_0_7_n8), .Z(
        npu_inst_int_data_x_0__7__0_) );
  MUX2_X1 npu_inst_pe_1_0_7_U146 ( .A(npu_inst_pe_1_0_7_n17), .B(
        npu_inst_pe_1_0_7_n16), .S(npu_inst_pe_1_0_7_n6), .Z(
        npu_inst_pe_1_0_7_n18) );
  MUX2_X1 npu_inst_pe_1_0_7_U145 ( .A(npu_inst_pe_1_0_7_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_0_7_int_q_reg_h_1__0_), .S(npu_inst_pe_1_0_7_n4), .Z(
        npu_inst_pe_1_0_7_n17) );
  MUX2_X1 npu_inst_pe_1_0_7_U144 ( .A(npu_inst_pe_1_0_7_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_0_7_int_q_reg_h_3__0_), .S(npu_inst_pe_1_0_7_n4), .Z(
        npu_inst_pe_1_0_7_n16) );
  MUX2_X1 npu_inst_pe_1_0_7_U143 ( .A(npu_inst_pe_1_0_7_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_0_7_int_q_reg_h_5__0_), .S(npu_inst_pe_1_0_7_n4), .Z(
        npu_inst_pe_1_0_7_n15) );
  XOR2_X1 npu_inst_pe_1_0_7_U142 ( .A(npu_inst_pe_1_0_7_int_data_0_), .B(
        npu_inst_pe_1_0_7_int_q_acc_0_), .Z(npu_inst_pe_1_0_7_N73) );
  AND2_X1 npu_inst_pe_1_0_7_U141 ( .A1(npu_inst_pe_1_0_7_int_q_acc_0_), .A2(
        npu_inst_pe_1_0_7_int_data_0_), .ZN(npu_inst_pe_1_0_7_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_0_7_U140 ( .A(npu_inst_pe_1_0_7_int_q_acc_0_), .B(
        npu_inst_pe_1_0_7_n13), .ZN(npu_inst_pe_1_0_7_N65) );
  OR2_X1 npu_inst_pe_1_0_7_U139 ( .A1(npu_inst_pe_1_0_7_n13), .A2(
        npu_inst_pe_1_0_7_int_q_acc_0_), .ZN(npu_inst_pe_1_0_7_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_0_7_U138 ( .A(npu_inst_pe_1_0_7_int_q_acc_2_), .B(
        npu_inst_pe_1_0_7_add_79_carry_2_), .Z(npu_inst_pe_1_0_7_N75) );
  AND2_X1 npu_inst_pe_1_0_7_U137 ( .A1(npu_inst_pe_1_0_7_add_79_carry_2_), 
        .A2(npu_inst_pe_1_0_7_int_q_acc_2_), .ZN(
        npu_inst_pe_1_0_7_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_0_7_U136 ( .A(npu_inst_pe_1_0_7_int_q_acc_3_), .B(
        npu_inst_pe_1_0_7_add_79_carry_3_), .Z(npu_inst_pe_1_0_7_N76) );
  AND2_X1 npu_inst_pe_1_0_7_U135 ( .A1(npu_inst_pe_1_0_7_add_79_carry_3_), 
        .A2(npu_inst_pe_1_0_7_int_q_acc_3_), .ZN(
        npu_inst_pe_1_0_7_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_0_7_U134 ( .A(npu_inst_pe_1_0_7_int_q_acc_4_), .B(
        npu_inst_pe_1_0_7_add_79_carry_4_), .Z(npu_inst_pe_1_0_7_N77) );
  AND2_X1 npu_inst_pe_1_0_7_U133 ( .A1(npu_inst_pe_1_0_7_add_79_carry_4_), 
        .A2(npu_inst_pe_1_0_7_int_q_acc_4_), .ZN(
        npu_inst_pe_1_0_7_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_0_7_U132 ( .A(npu_inst_pe_1_0_7_int_q_acc_5_), .B(
        npu_inst_pe_1_0_7_add_79_carry_5_), .Z(npu_inst_pe_1_0_7_N78) );
  AND2_X1 npu_inst_pe_1_0_7_U131 ( .A1(npu_inst_pe_1_0_7_add_79_carry_5_), 
        .A2(npu_inst_pe_1_0_7_int_q_acc_5_), .ZN(
        npu_inst_pe_1_0_7_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_0_7_U130 ( .A(npu_inst_pe_1_0_7_int_q_acc_6_), .B(
        npu_inst_pe_1_0_7_add_79_carry_6_), .Z(npu_inst_pe_1_0_7_N79) );
  AND2_X1 npu_inst_pe_1_0_7_U129 ( .A1(npu_inst_pe_1_0_7_add_79_carry_6_), 
        .A2(npu_inst_pe_1_0_7_int_q_acc_6_), .ZN(
        npu_inst_pe_1_0_7_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_0_7_U128 ( .A(npu_inst_pe_1_0_7_int_q_acc_7_), .B(
        npu_inst_pe_1_0_7_add_79_carry_7_), .Z(npu_inst_pe_1_0_7_N80) );
  XNOR2_X1 npu_inst_pe_1_0_7_U127 ( .A(npu_inst_pe_1_0_7_sub_77_carry_2_), .B(
        npu_inst_pe_1_0_7_int_q_acc_2_), .ZN(npu_inst_pe_1_0_7_N67) );
  OR2_X1 npu_inst_pe_1_0_7_U126 ( .A1(npu_inst_pe_1_0_7_int_q_acc_2_), .A2(
        npu_inst_pe_1_0_7_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_0_7_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_0_7_U125 ( .A(npu_inst_pe_1_0_7_sub_77_carry_3_), .B(
        npu_inst_pe_1_0_7_int_q_acc_3_), .ZN(npu_inst_pe_1_0_7_N68) );
  OR2_X1 npu_inst_pe_1_0_7_U124 ( .A1(npu_inst_pe_1_0_7_int_q_acc_3_), .A2(
        npu_inst_pe_1_0_7_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_0_7_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_0_7_U123 ( .A(npu_inst_pe_1_0_7_sub_77_carry_4_), .B(
        npu_inst_pe_1_0_7_int_q_acc_4_), .ZN(npu_inst_pe_1_0_7_N69) );
  OR2_X1 npu_inst_pe_1_0_7_U122 ( .A1(npu_inst_pe_1_0_7_int_q_acc_4_), .A2(
        npu_inst_pe_1_0_7_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_0_7_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_0_7_U121 ( .A(npu_inst_pe_1_0_7_sub_77_carry_5_), .B(
        npu_inst_pe_1_0_7_int_q_acc_5_), .ZN(npu_inst_pe_1_0_7_N70) );
  OR2_X1 npu_inst_pe_1_0_7_U120 ( .A1(npu_inst_pe_1_0_7_int_q_acc_5_), .A2(
        npu_inst_pe_1_0_7_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_0_7_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_0_7_U119 ( .A(npu_inst_pe_1_0_7_sub_77_carry_6_), .B(
        npu_inst_pe_1_0_7_int_q_acc_6_), .ZN(npu_inst_pe_1_0_7_N71) );
  OR2_X1 npu_inst_pe_1_0_7_U118 ( .A1(npu_inst_pe_1_0_7_int_q_acc_6_), .A2(
        npu_inst_pe_1_0_7_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_0_7_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_0_7_U117 ( .A(npu_inst_pe_1_0_7_int_q_acc_7_), .B(
        npu_inst_pe_1_0_7_sub_77_carry_7_), .ZN(npu_inst_pe_1_0_7_N72) );
  INV_X1 npu_inst_pe_1_0_7_U116 ( .A(npu_inst_n79), .ZN(npu_inst_pe_1_0_7_n7)
         );
  INV_X1 npu_inst_pe_1_0_7_U115 ( .A(npu_inst_pe_1_0_7_n7), .ZN(
        npu_inst_pe_1_0_7_n6) );
  INV_X1 npu_inst_pe_1_0_7_U114 ( .A(npu_inst_n60), .ZN(npu_inst_pe_1_0_7_n3)
         );
  AOI22_X1 npu_inst_pe_1_0_7_U113 ( .A1(npu_inst_int_data_y_1__7__0_), .A2(
        npu_inst_pe_1_0_7_n58), .B1(npu_inst_pe_1_0_7_n114), .B2(
        npu_inst_pe_1_0_7_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_0_7_n57) );
  INV_X1 npu_inst_pe_1_0_7_U112 ( .A(npu_inst_pe_1_0_7_n57), .ZN(
        npu_inst_pe_1_0_7_n108) );
  AOI22_X1 npu_inst_pe_1_0_7_U111 ( .A1(npu_inst_int_data_y_1__7__0_), .A2(
        npu_inst_pe_1_0_7_n54), .B1(npu_inst_pe_1_0_7_n115), .B2(
        npu_inst_pe_1_0_7_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_0_7_n53) );
  INV_X1 npu_inst_pe_1_0_7_U110 ( .A(npu_inst_pe_1_0_7_n53), .ZN(
        npu_inst_pe_1_0_7_n109) );
  AOI22_X1 npu_inst_pe_1_0_7_U107 ( .A1(npu_inst_int_data_y_1__7__0_), .A2(
        npu_inst_pe_1_0_7_n50), .B1(npu_inst_pe_1_0_7_n116), .B2(
        npu_inst_pe_1_0_7_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_0_7_n49) );
  INV_X1 npu_inst_pe_1_0_7_U106 ( .A(npu_inst_pe_1_0_7_n49), .ZN(
        npu_inst_pe_1_0_7_n110) );
  AOI22_X1 npu_inst_pe_1_0_7_U105 ( .A1(npu_inst_int_data_y_1__7__0_), .A2(
        npu_inst_pe_1_0_7_n46), .B1(npu_inst_pe_1_0_7_n117), .B2(
        npu_inst_pe_1_0_7_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_0_7_n45) );
  INV_X1 npu_inst_pe_1_0_7_U104 ( .A(npu_inst_pe_1_0_7_n45), .ZN(
        npu_inst_pe_1_0_7_n111) );
  AOI22_X1 npu_inst_pe_1_0_7_U103 ( .A1(npu_inst_int_data_y_1__7__0_), .A2(
        npu_inst_pe_1_0_7_n42), .B1(npu_inst_pe_1_0_7_n119), .B2(
        npu_inst_pe_1_0_7_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_0_7_n41) );
  INV_X1 npu_inst_pe_1_0_7_U102 ( .A(npu_inst_pe_1_0_7_n41), .ZN(
        npu_inst_pe_1_0_7_n112) );
  AOI22_X1 npu_inst_pe_1_0_7_U101 ( .A1(npu_inst_int_data_y_1__7__1_), .A2(
        npu_inst_pe_1_0_7_n58), .B1(npu_inst_pe_1_0_7_n114), .B2(
        npu_inst_pe_1_0_7_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_0_7_n59) );
  INV_X1 npu_inst_pe_1_0_7_U100 ( .A(npu_inst_pe_1_0_7_n59), .ZN(
        npu_inst_pe_1_0_7_n102) );
  AOI22_X1 npu_inst_pe_1_0_7_U99 ( .A1(npu_inst_int_data_y_1__7__1_), .A2(
        npu_inst_pe_1_0_7_n54), .B1(npu_inst_pe_1_0_7_n115), .B2(
        npu_inst_pe_1_0_7_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_0_7_n55) );
  INV_X1 npu_inst_pe_1_0_7_U98 ( .A(npu_inst_pe_1_0_7_n55), .ZN(
        npu_inst_pe_1_0_7_n103) );
  AOI22_X1 npu_inst_pe_1_0_7_U97 ( .A1(npu_inst_int_data_y_1__7__1_), .A2(
        npu_inst_pe_1_0_7_n50), .B1(npu_inst_pe_1_0_7_n116), .B2(
        npu_inst_pe_1_0_7_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_0_7_n51) );
  INV_X1 npu_inst_pe_1_0_7_U96 ( .A(npu_inst_pe_1_0_7_n51), .ZN(
        npu_inst_pe_1_0_7_n104) );
  AOI22_X1 npu_inst_pe_1_0_7_U95 ( .A1(npu_inst_int_data_y_1__7__1_), .A2(
        npu_inst_pe_1_0_7_n46), .B1(npu_inst_pe_1_0_7_n117), .B2(
        npu_inst_pe_1_0_7_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_0_7_n47) );
  INV_X1 npu_inst_pe_1_0_7_U94 ( .A(npu_inst_pe_1_0_7_n47), .ZN(
        npu_inst_pe_1_0_7_n105) );
  AOI22_X1 npu_inst_pe_1_0_7_U93 ( .A1(npu_inst_int_data_y_1__7__1_), .A2(
        npu_inst_pe_1_0_7_n42), .B1(npu_inst_pe_1_0_7_n119), .B2(
        npu_inst_pe_1_0_7_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_0_7_n43) );
  INV_X1 npu_inst_pe_1_0_7_U92 ( .A(npu_inst_pe_1_0_7_n43), .ZN(
        npu_inst_pe_1_0_7_n106) );
  AOI22_X1 npu_inst_pe_1_0_7_U91 ( .A1(npu_inst_pe_1_0_7_n38), .A2(
        npu_inst_int_data_y_1__7__1_), .B1(npu_inst_pe_1_0_7_n118), .B2(
        npu_inst_pe_1_0_7_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_0_7_n39) );
  INV_X1 npu_inst_pe_1_0_7_U90 ( .A(npu_inst_pe_1_0_7_n39), .ZN(
        npu_inst_pe_1_0_7_n107) );
  AOI22_X1 npu_inst_pe_1_0_7_U89 ( .A1(npu_inst_pe_1_0_7_n38), .A2(
        npu_inst_int_data_y_1__7__0_), .B1(npu_inst_pe_1_0_7_n118), .B2(
        npu_inst_pe_1_0_7_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_0_7_n37) );
  INV_X1 npu_inst_pe_1_0_7_U88 ( .A(npu_inst_pe_1_0_7_n37), .ZN(
        npu_inst_pe_1_0_7_n113) );
  AND2_X1 npu_inst_pe_1_0_7_U87 ( .A1(npu_inst_pe_1_0_7_n2), .A2(
        npu_inst_pe_1_0_7_int_q_acc_7_), .ZN(o_data[7]) );
  AND2_X1 npu_inst_pe_1_0_7_U86 ( .A1(npu_inst_pe_1_0_7_int_q_acc_6_), .A2(
        npu_inst_pe_1_0_7_n2), .ZN(o_data[6]) );
  AND2_X1 npu_inst_pe_1_0_7_U85 ( .A1(npu_inst_pe_1_0_7_int_q_acc_5_), .A2(
        npu_inst_pe_1_0_7_n2), .ZN(o_data[5]) );
  AND2_X1 npu_inst_pe_1_0_7_U84 ( .A1(npu_inst_pe_1_0_7_int_q_acc_4_), .A2(
        npu_inst_pe_1_0_7_n2), .ZN(o_data[4]) );
  AND2_X1 npu_inst_pe_1_0_7_U83 ( .A1(npu_inst_pe_1_0_7_int_q_acc_3_), .A2(
        npu_inst_pe_1_0_7_n2), .ZN(o_data[3]) );
  NOR3_X1 npu_inst_pe_1_0_7_U82 ( .A1(npu_inst_pe_1_0_7_n26), .A2(npu_inst_n60), .A3(npu_inst_int_ckg[56]), .ZN(npu_inst_pe_1_0_7_n85) );
  OR2_X1 npu_inst_pe_1_0_7_U81 ( .A1(npu_inst_pe_1_0_7_n85), .A2(
        npu_inst_pe_1_0_7_n2), .ZN(npu_inst_pe_1_0_7_N84) );
  AND2_X1 npu_inst_pe_1_0_7_U80 ( .A1(npu_inst_pe_1_0_7_int_q_acc_0_), .A2(
        npu_inst_pe_1_0_7_n1), .ZN(o_data[0]) );
  AND2_X1 npu_inst_pe_1_0_7_U79 ( .A1(npu_inst_pe_1_0_7_int_q_acc_1_), .A2(
        npu_inst_pe_1_0_7_n1), .ZN(o_data[1]) );
  AND2_X1 npu_inst_pe_1_0_7_U78 ( .A1(npu_inst_pe_1_0_7_int_q_acc_2_), .A2(
        npu_inst_pe_1_0_7_n1), .ZN(o_data[2]) );
  AOI222_X1 npu_inst_pe_1_0_7_U77 ( .A1(npu_inst_int_data_res_1__7__0_), .A2(
        npu_inst_pe_1_0_7_n1), .B1(npu_inst_pe_1_0_7_N73), .B2(
        npu_inst_pe_1_0_7_n76), .C1(npu_inst_pe_1_0_7_N65), .C2(
        npu_inst_pe_1_0_7_n77), .ZN(npu_inst_pe_1_0_7_n84) );
  INV_X1 npu_inst_pe_1_0_7_U76 ( .A(npu_inst_pe_1_0_7_n84), .ZN(
        npu_inst_pe_1_0_7_n101) );
  AOI222_X1 npu_inst_pe_1_0_7_U75 ( .A1(npu_inst_int_data_res_1__7__7_), .A2(
        npu_inst_pe_1_0_7_n1), .B1(npu_inst_pe_1_0_7_N80), .B2(
        npu_inst_pe_1_0_7_n76), .C1(npu_inst_pe_1_0_7_N72), .C2(
        npu_inst_pe_1_0_7_n77), .ZN(npu_inst_pe_1_0_7_n75) );
  INV_X1 npu_inst_pe_1_0_7_U74 ( .A(npu_inst_pe_1_0_7_n75), .ZN(
        npu_inst_pe_1_0_7_n33) );
  AOI222_X1 npu_inst_pe_1_0_7_U73 ( .A1(npu_inst_int_data_res_1__7__1_), .A2(
        npu_inst_pe_1_0_7_n1), .B1(npu_inst_pe_1_0_7_N74), .B2(
        npu_inst_pe_1_0_7_n76), .C1(npu_inst_pe_1_0_7_N66), .C2(
        npu_inst_pe_1_0_7_n77), .ZN(npu_inst_pe_1_0_7_n83) );
  INV_X1 npu_inst_pe_1_0_7_U72 ( .A(npu_inst_pe_1_0_7_n83), .ZN(
        npu_inst_pe_1_0_7_n100) );
  AOI222_X1 npu_inst_pe_1_0_7_U71 ( .A1(npu_inst_int_data_res_1__7__2_), .A2(
        npu_inst_pe_1_0_7_n1), .B1(npu_inst_pe_1_0_7_N75), .B2(
        npu_inst_pe_1_0_7_n76), .C1(npu_inst_pe_1_0_7_N67), .C2(
        npu_inst_pe_1_0_7_n77), .ZN(npu_inst_pe_1_0_7_n82) );
  INV_X1 npu_inst_pe_1_0_7_U70 ( .A(npu_inst_pe_1_0_7_n82), .ZN(
        npu_inst_pe_1_0_7_n99) );
  AOI222_X1 npu_inst_pe_1_0_7_U69 ( .A1(npu_inst_int_data_res_1__7__3_), .A2(
        npu_inst_pe_1_0_7_n1), .B1(npu_inst_pe_1_0_7_N76), .B2(
        npu_inst_pe_1_0_7_n76), .C1(npu_inst_pe_1_0_7_N68), .C2(
        npu_inst_pe_1_0_7_n77), .ZN(npu_inst_pe_1_0_7_n81) );
  INV_X1 npu_inst_pe_1_0_7_U68 ( .A(npu_inst_pe_1_0_7_n81), .ZN(
        npu_inst_pe_1_0_7_n98) );
  AOI222_X1 npu_inst_pe_1_0_7_U67 ( .A1(npu_inst_int_data_res_1__7__4_), .A2(
        npu_inst_pe_1_0_7_n1), .B1(npu_inst_pe_1_0_7_N77), .B2(
        npu_inst_pe_1_0_7_n76), .C1(npu_inst_pe_1_0_7_N69), .C2(
        npu_inst_pe_1_0_7_n77), .ZN(npu_inst_pe_1_0_7_n80) );
  INV_X1 npu_inst_pe_1_0_7_U66 ( .A(npu_inst_pe_1_0_7_n80), .ZN(
        npu_inst_pe_1_0_7_n36) );
  AOI222_X1 npu_inst_pe_1_0_7_U65 ( .A1(npu_inst_int_data_res_1__7__5_), .A2(
        npu_inst_pe_1_0_7_n1), .B1(npu_inst_pe_1_0_7_N78), .B2(
        npu_inst_pe_1_0_7_n76), .C1(npu_inst_pe_1_0_7_N70), .C2(
        npu_inst_pe_1_0_7_n77), .ZN(npu_inst_pe_1_0_7_n79) );
  INV_X1 npu_inst_pe_1_0_7_U64 ( .A(npu_inst_pe_1_0_7_n79), .ZN(
        npu_inst_pe_1_0_7_n35) );
  AOI222_X1 npu_inst_pe_1_0_7_U63 ( .A1(npu_inst_int_data_res_1__7__6_), .A2(
        npu_inst_pe_1_0_7_n1), .B1(npu_inst_pe_1_0_7_N79), .B2(
        npu_inst_pe_1_0_7_n76), .C1(npu_inst_pe_1_0_7_N71), .C2(
        npu_inst_pe_1_0_7_n77), .ZN(npu_inst_pe_1_0_7_n78) );
  INV_X1 npu_inst_pe_1_0_7_U62 ( .A(npu_inst_pe_1_0_7_n78), .ZN(
        npu_inst_pe_1_0_7_n34) );
  INV_X1 npu_inst_pe_1_0_7_U61 ( .A(npu_inst_pe_1_0_7_int_data_1_), .ZN(
        npu_inst_pe_1_0_7_n14) );
  AND2_X1 npu_inst_pe_1_0_7_U60 ( .A1(npu_inst_int_data_x_0__7__1_), .A2(
        npu_inst_pe_1_0_7_int_q_weight_1_), .ZN(npu_inst_pe_1_0_7_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_0_7_U59 ( .A1(npu_inst_int_data_x_0__7__0_), .A2(
        npu_inst_pe_1_0_7_int_q_weight_1_), .ZN(npu_inst_pe_1_0_7_int_data_0_)
         );
  NAND2_X1 npu_inst_pe_1_0_7_U58 ( .A1(npu_inst_pe_1_0_7_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_0_7_n60), .ZN(npu_inst_pe_1_0_7_n74) );
  OAI21_X1 npu_inst_pe_1_0_7_U57 ( .B1(npu_inst_pe_1_0_7_n63), .B2(
        npu_inst_pe_1_0_7_n60), .A(npu_inst_pe_1_0_7_n74), .ZN(
        npu_inst_pe_1_0_7_n97) );
  NAND2_X1 npu_inst_pe_1_0_7_U56 ( .A1(npu_inst_pe_1_0_7_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_0_7_n60), .ZN(npu_inst_pe_1_0_7_n73) );
  OAI21_X1 npu_inst_pe_1_0_7_U55 ( .B1(npu_inst_pe_1_0_7_n61), .B2(
        npu_inst_pe_1_0_7_n60), .A(npu_inst_pe_1_0_7_n73), .ZN(
        npu_inst_pe_1_0_7_n96) );
  NAND2_X1 npu_inst_pe_1_0_7_U54 ( .A1(npu_inst_pe_1_0_7_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_0_7_n56), .ZN(npu_inst_pe_1_0_7_n72) );
  OAI21_X1 npu_inst_pe_1_0_7_U53 ( .B1(npu_inst_pe_1_0_7_n63), .B2(
        npu_inst_pe_1_0_7_n56), .A(npu_inst_pe_1_0_7_n72), .ZN(
        npu_inst_pe_1_0_7_n95) );
  NAND2_X1 npu_inst_pe_1_0_7_U52 ( .A1(npu_inst_pe_1_0_7_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_0_7_n56), .ZN(npu_inst_pe_1_0_7_n71) );
  OAI21_X1 npu_inst_pe_1_0_7_U51 ( .B1(npu_inst_pe_1_0_7_n61), .B2(
        npu_inst_pe_1_0_7_n56), .A(npu_inst_pe_1_0_7_n71), .ZN(
        npu_inst_pe_1_0_7_n94) );
  NAND2_X1 npu_inst_pe_1_0_7_U50 ( .A1(npu_inst_pe_1_0_7_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_0_7_n52), .ZN(npu_inst_pe_1_0_7_n70) );
  OAI21_X1 npu_inst_pe_1_0_7_U49 ( .B1(npu_inst_pe_1_0_7_n63), .B2(
        npu_inst_pe_1_0_7_n52), .A(npu_inst_pe_1_0_7_n70), .ZN(
        npu_inst_pe_1_0_7_n93) );
  NAND2_X1 npu_inst_pe_1_0_7_U48 ( .A1(npu_inst_pe_1_0_7_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_0_7_n52), .ZN(npu_inst_pe_1_0_7_n69) );
  OAI21_X1 npu_inst_pe_1_0_7_U47 ( .B1(npu_inst_pe_1_0_7_n61), .B2(
        npu_inst_pe_1_0_7_n52), .A(npu_inst_pe_1_0_7_n69), .ZN(
        npu_inst_pe_1_0_7_n92) );
  NAND2_X1 npu_inst_pe_1_0_7_U46 ( .A1(npu_inst_pe_1_0_7_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_0_7_n48), .ZN(npu_inst_pe_1_0_7_n68) );
  OAI21_X1 npu_inst_pe_1_0_7_U45 ( .B1(npu_inst_pe_1_0_7_n63), .B2(
        npu_inst_pe_1_0_7_n48), .A(npu_inst_pe_1_0_7_n68), .ZN(
        npu_inst_pe_1_0_7_n91) );
  NAND2_X1 npu_inst_pe_1_0_7_U44 ( .A1(npu_inst_pe_1_0_7_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_0_7_n48), .ZN(npu_inst_pe_1_0_7_n67) );
  OAI21_X1 npu_inst_pe_1_0_7_U43 ( .B1(npu_inst_pe_1_0_7_n61), .B2(
        npu_inst_pe_1_0_7_n48), .A(npu_inst_pe_1_0_7_n67), .ZN(
        npu_inst_pe_1_0_7_n90) );
  NAND2_X1 npu_inst_pe_1_0_7_U42 ( .A1(npu_inst_pe_1_0_7_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_0_7_n44), .ZN(npu_inst_pe_1_0_7_n66) );
  OAI21_X1 npu_inst_pe_1_0_7_U41 ( .B1(npu_inst_pe_1_0_7_n63), .B2(
        npu_inst_pe_1_0_7_n44), .A(npu_inst_pe_1_0_7_n66), .ZN(
        npu_inst_pe_1_0_7_n89) );
  NAND2_X1 npu_inst_pe_1_0_7_U40 ( .A1(npu_inst_pe_1_0_7_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_0_7_n44), .ZN(npu_inst_pe_1_0_7_n65) );
  OAI21_X1 npu_inst_pe_1_0_7_U39 ( .B1(npu_inst_pe_1_0_7_n61), .B2(
        npu_inst_pe_1_0_7_n44), .A(npu_inst_pe_1_0_7_n65), .ZN(
        npu_inst_pe_1_0_7_n88) );
  NAND2_X1 npu_inst_pe_1_0_7_U38 ( .A1(npu_inst_pe_1_0_7_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_0_7_n40), .ZN(npu_inst_pe_1_0_7_n64) );
  OAI21_X1 npu_inst_pe_1_0_7_U37 ( .B1(npu_inst_pe_1_0_7_n63), .B2(
        npu_inst_pe_1_0_7_n40), .A(npu_inst_pe_1_0_7_n64), .ZN(
        npu_inst_pe_1_0_7_n87) );
  NAND2_X1 npu_inst_pe_1_0_7_U36 ( .A1(npu_inst_pe_1_0_7_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_0_7_n40), .ZN(npu_inst_pe_1_0_7_n62) );
  OAI21_X1 npu_inst_pe_1_0_7_U35 ( .B1(npu_inst_pe_1_0_7_n61), .B2(
        npu_inst_pe_1_0_7_n40), .A(npu_inst_pe_1_0_7_n62), .ZN(
        npu_inst_pe_1_0_7_n86) );
  AND2_X1 npu_inst_pe_1_0_7_U34 ( .A1(npu_inst_pe_1_0_7_N93), .A2(npu_inst_n60), .ZN(npu_inst_pe_1_0_7_o_data_v_0_) );
  AND2_X1 npu_inst_pe_1_0_7_U33 ( .A1(npu_inst_n60), .A2(npu_inst_pe_1_0_7_N94), .ZN(npu_inst_pe_1_0_7_o_data_v_1_) );
  INV_X1 npu_inst_pe_1_0_7_U32 ( .A(npu_inst_pe_1_0_7_int_data_0_), .ZN(
        npu_inst_pe_1_0_7_n13) );
  AOI22_X1 npu_inst_pe_1_0_7_U31 ( .A1(npu_inst_n60), .A2(
        npu_inst_int_data_y_1__7__1_), .B1(npu_inst_pe_1_0_7_n3), .B2(
        int_i_data_h_npu1[1]), .ZN(npu_inst_pe_1_0_7_n63) );
  AOI22_X1 npu_inst_pe_1_0_7_U30 ( .A1(npu_inst_n60), .A2(
        npu_inst_int_data_y_1__7__0_), .B1(npu_inst_pe_1_0_7_n3), .B2(
        int_i_data_h_npu1[0]), .ZN(npu_inst_pe_1_0_7_n61) );
  INV_X1 npu_inst_pe_1_0_7_U29 ( .A(npu_inst_n71), .ZN(npu_inst_pe_1_0_7_n5)
         );
  OR3_X1 npu_inst_pe_1_0_7_U28 ( .A1(npu_inst_pe_1_0_7_n6), .A2(
        npu_inst_pe_1_0_7_n8), .A3(npu_inst_pe_1_0_7_n5), .ZN(
        npu_inst_pe_1_0_7_n56) );
  OR3_X1 npu_inst_pe_1_0_7_U27 ( .A1(npu_inst_pe_1_0_7_n5), .A2(
        npu_inst_pe_1_0_7_n8), .A3(npu_inst_pe_1_0_7_n7), .ZN(
        npu_inst_pe_1_0_7_n48) );
  INV_X1 npu_inst_pe_1_0_7_U26 ( .A(npu_inst_pe_1_0_7_n5), .ZN(
        npu_inst_pe_1_0_7_n4) );
  INV_X1 npu_inst_pe_1_0_7_U25 ( .A(npu_inst_n126), .ZN(npu_inst_pe_1_0_7_n12)
         );
  OR3_X1 npu_inst_pe_1_0_7_U24 ( .A1(npu_inst_pe_1_0_7_n4), .A2(
        npu_inst_pe_1_0_7_n8), .A3(npu_inst_pe_1_0_7_n7), .ZN(
        npu_inst_pe_1_0_7_n52) );
  OR3_X1 npu_inst_pe_1_0_7_U23 ( .A1(npu_inst_pe_1_0_7_n6), .A2(
        npu_inst_pe_1_0_7_n8), .A3(npu_inst_pe_1_0_7_n4), .ZN(
        npu_inst_pe_1_0_7_n60) );
  NOR2_X1 npu_inst_pe_1_0_7_U22 ( .A1(npu_inst_pe_1_0_7_n60), .A2(
        npu_inst_pe_1_0_7_n3), .ZN(npu_inst_pe_1_0_7_n58) );
  NOR2_X1 npu_inst_pe_1_0_7_U21 ( .A1(npu_inst_pe_1_0_7_n56), .A2(
        npu_inst_pe_1_0_7_n3), .ZN(npu_inst_pe_1_0_7_n54) );
  NOR2_X1 npu_inst_pe_1_0_7_U20 ( .A1(npu_inst_pe_1_0_7_n52), .A2(
        npu_inst_pe_1_0_7_n3), .ZN(npu_inst_pe_1_0_7_n50) );
  NOR2_X1 npu_inst_pe_1_0_7_U19 ( .A1(npu_inst_pe_1_0_7_n48), .A2(
        npu_inst_pe_1_0_7_n3), .ZN(npu_inst_pe_1_0_7_n46) );
  NOR2_X1 npu_inst_pe_1_0_7_U18 ( .A1(npu_inst_pe_1_0_7_n40), .A2(
        npu_inst_pe_1_0_7_n3), .ZN(npu_inst_pe_1_0_7_n38) );
  NOR2_X1 npu_inst_pe_1_0_7_U17 ( .A1(npu_inst_pe_1_0_7_n44), .A2(
        npu_inst_pe_1_0_7_n3), .ZN(npu_inst_pe_1_0_7_n42) );
  BUF_X1 npu_inst_pe_1_0_7_U16 ( .A(npu_inst_n106), .Z(npu_inst_pe_1_0_7_n8)
         );
  BUF_X1 npu_inst_pe_1_0_7_U15 ( .A(npu_inst_pe_1_0_7_n12), .Z(
        npu_inst_pe_1_0_7_n11) );
  BUF_X1 npu_inst_pe_1_0_7_U14 ( .A(npu_inst_pe_1_0_7_n12), .Z(
        npu_inst_pe_1_0_7_n10) );
  BUF_X1 npu_inst_pe_1_0_7_U13 ( .A(npu_inst_pe_1_0_7_n12), .Z(
        npu_inst_pe_1_0_7_n9) );
  INV_X1 npu_inst_pe_1_0_7_U12 ( .A(npu_inst_pe_1_0_7_n38), .ZN(
        npu_inst_pe_1_0_7_n118) );
  INV_X1 npu_inst_pe_1_0_7_U11 ( .A(npu_inst_pe_1_0_7_n58), .ZN(
        npu_inst_pe_1_0_7_n114) );
  INV_X1 npu_inst_pe_1_0_7_U10 ( .A(npu_inst_pe_1_0_7_n54), .ZN(
        npu_inst_pe_1_0_7_n115) );
  INV_X1 npu_inst_pe_1_0_7_U9 ( .A(npu_inst_pe_1_0_7_n50), .ZN(
        npu_inst_pe_1_0_7_n116) );
  INV_X1 npu_inst_pe_1_0_7_U8 ( .A(npu_inst_pe_1_0_7_n46), .ZN(
        npu_inst_pe_1_0_7_n117) );
  INV_X1 npu_inst_pe_1_0_7_U7 ( .A(npu_inst_pe_1_0_7_n42), .ZN(
        npu_inst_pe_1_0_7_n119) );
  BUF_X1 npu_inst_pe_1_0_7_U6 ( .A(npu_inst_n35), .Z(npu_inst_pe_1_0_7_n2) );
  BUF_X1 npu_inst_pe_1_0_7_U5 ( .A(npu_inst_n35), .Z(npu_inst_pe_1_0_7_n1) );
  NOR2_X1 npu_inst_pe_1_0_7_U4 ( .A1(npu_inst_pe_1_0_7_int_q_weight_0_), .A2(
        npu_inst_pe_1_0_7_n1), .ZN(npu_inst_pe_1_0_7_n76) );
  NOR2_X1 npu_inst_pe_1_0_7_U3 ( .A1(npu_inst_pe_1_0_7_n27), .A2(
        npu_inst_pe_1_0_7_n1), .ZN(npu_inst_pe_1_0_7_n77) );
  FA_X1 npu_inst_pe_1_0_7_sub_77_U2_1 ( .A(npu_inst_pe_1_0_7_int_q_acc_1_), 
        .B(npu_inst_pe_1_0_7_n14), .CI(npu_inst_pe_1_0_7_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_0_7_sub_77_carry_2_), .S(npu_inst_pe_1_0_7_N66) );
  FA_X1 npu_inst_pe_1_0_7_add_79_U1_1 ( .A(npu_inst_pe_1_0_7_int_q_acc_1_), 
        .B(npu_inst_pe_1_0_7_int_data_1_), .CI(
        npu_inst_pe_1_0_7_add_79_carry_1_), .CO(
        npu_inst_pe_1_0_7_add_79_carry_2_), .S(npu_inst_pe_1_0_7_N74) );
  NAND3_X1 npu_inst_pe_1_0_7_U109 ( .A1(npu_inst_pe_1_0_7_n5), .A2(
        npu_inst_pe_1_0_7_n7), .A3(npu_inst_pe_1_0_7_n8), .ZN(
        npu_inst_pe_1_0_7_n44) );
  NAND3_X1 npu_inst_pe_1_0_7_U108 ( .A1(npu_inst_pe_1_0_7_n4), .A2(
        npu_inst_pe_1_0_7_n7), .A3(npu_inst_pe_1_0_7_n8), .ZN(
        npu_inst_pe_1_0_7_n40) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_0_7_n34), .CK(
        npu_inst_pe_1_0_7_net4132), .RN(npu_inst_pe_1_0_7_n9), .Q(
        npu_inst_pe_1_0_7_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_0_7_n35), .CK(
        npu_inst_pe_1_0_7_net4132), .RN(npu_inst_pe_1_0_7_n9), .Q(
        npu_inst_pe_1_0_7_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_0_7_n36), .CK(
        npu_inst_pe_1_0_7_net4132), .RN(npu_inst_pe_1_0_7_n9), .Q(
        npu_inst_pe_1_0_7_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_0_7_n98), .CK(
        npu_inst_pe_1_0_7_net4132), .RN(npu_inst_pe_1_0_7_n9), .Q(
        npu_inst_pe_1_0_7_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_0_7_n99), .CK(
        npu_inst_pe_1_0_7_net4132), .RN(npu_inst_pe_1_0_7_n9), .Q(
        npu_inst_pe_1_0_7_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_0_7_n100), 
        .CK(npu_inst_pe_1_0_7_net4132), .RN(npu_inst_pe_1_0_7_n9), .Q(
        npu_inst_pe_1_0_7_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_0_7_n33), .CK(
        npu_inst_pe_1_0_7_net4132), .RN(npu_inst_pe_1_0_7_n9), .Q(
        npu_inst_pe_1_0_7_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_0_7_n101), 
        .CK(npu_inst_pe_1_0_7_net4132), .RN(npu_inst_pe_1_0_7_n9), .Q(
        npu_inst_pe_1_0_7_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_weight_reg_0_ ( .D(npu_inst_n112), .CK(
        npu_inst_pe_1_0_7_net4138), .RN(npu_inst_pe_1_0_7_n9), .Q(
        npu_inst_pe_1_0_7_int_q_weight_0_), .QN(npu_inst_pe_1_0_7_n27) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_weight_reg_1_ ( .D(npu_inst_n118), .CK(
        npu_inst_pe_1_0_7_net4138), .RN(npu_inst_pe_1_0_7_n9), .Q(
        npu_inst_pe_1_0_7_int_q_weight_1_), .QN(npu_inst_pe_1_0_7_n26) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_0_7_n113), 
        .CK(npu_inst_pe_1_0_7_net4138), .RN(npu_inst_pe_1_0_7_n9), .Q(
        npu_inst_pe_1_0_7_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_0_7_n107), 
        .CK(npu_inst_pe_1_0_7_net4138), .RN(npu_inst_pe_1_0_7_n9), .Q(
        npu_inst_pe_1_0_7_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_0_7_n112), 
        .CK(npu_inst_pe_1_0_7_net4138), .RN(npu_inst_pe_1_0_7_n10), .Q(
        npu_inst_pe_1_0_7_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_0_7_n106), 
        .CK(npu_inst_pe_1_0_7_net4138), .RN(npu_inst_pe_1_0_7_n10), .Q(
        npu_inst_pe_1_0_7_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_0_7_n111), 
        .CK(npu_inst_pe_1_0_7_net4138), .RN(npu_inst_pe_1_0_7_n10), .Q(
        npu_inst_pe_1_0_7_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_0_7_n105), 
        .CK(npu_inst_pe_1_0_7_net4138), .RN(npu_inst_pe_1_0_7_n10), .Q(
        npu_inst_pe_1_0_7_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_0_7_n110), 
        .CK(npu_inst_pe_1_0_7_net4138), .RN(npu_inst_pe_1_0_7_n10), .Q(
        npu_inst_pe_1_0_7_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_0_7_n104), 
        .CK(npu_inst_pe_1_0_7_net4138), .RN(npu_inst_pe_1_0_7_n10), .Q(
        npu_inst_pe_1_0_7_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_0_7_n109), 
        .CK(npu_inst_pe_1_0_7_net4138), .RN(npu_inst_pe_1_0_7_n10), .Q(
        npu_inst_pe_1_0_7_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_0_7_n103), 
        .CK(npu_inst_pe_1_0_7_net4138), .RN(npu_inst_pe_1_0_7_n10), .Q(
        npu_inst_pe_1_0_7_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_0_7_n108), 
        .CK(npu_inst_pe_1_0_7_net4138), .RN(npu_inst_pe_1_0_7_n10), .Q(
        npu_inst_pe_1_0_7_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_0_7_n102), 
        .CK(npu_inst_pe_1_0_7_net4138), .RN(npu_inst_pe_1_0_7_n10), .Q(
        npu_inst_pe_1_0_7_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_0_7_n86), 
        .CK(npu_inst_pe_1_0_7_net4138), .RN(npu_inst_pe_1_0_7_n10), .Q(
        npu_inst_pe_1_0_7_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_0_7_n87), 
        .CK(npu_inst_pe_1_0_7_net4138), .RN(npu_inst_pe_1_0_7_n10), .Q(
        npu_inst_pe_1_0_7_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_0_7_n88), 
        .CK(npu_inst_pe_1_0_7_net4138), .RN(npu_inst_pe_1_0_7_n11), .Q(
        npu_inst_pe_1_0_7_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_0_7_n89), 
        .CK(npu_inst_pe_1_0_7_net4138), .RN(npu_inst_pe_1_0_7_n11), .Q(
        npu_inst_pe_1_0_7_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_0_7_n90), 
        .CK(npu_inst_pe_1_0_7_net4138), .RN(npu_inst_pe_1_0_7_n11), .Q(
        npu_inst_pe_1_0_7_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_0_7_n91), 
        .CK(npu_inst_pe_1_0_7_net4138), .RN(npu_inst_pe_1_0_7_n11), .Q(
        npu_inst_pe_1_0_7_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_0_7_n92), 
        .CK(npu_inst_pe_1_0_7_net4138), .RN(npu_inst_pe_1_0_7_n11), .Q(
        npu_inst_pe_1_0_7_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_0_7_n93), 
        .CK(npu_inst_pe_1_0_7_net4138), .RN(npu_inst_pe_1_0_7_n11), .Q(
        npu_inst_pe_1_0_7_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_0_7_n94), 
        .CK(npu_inst_pe_1_0_7_net4138), .RN(npu_inst_pe_1_0_7_n11), .Q(
        npu_inst_pe_1_0_7_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_0_7_n95), 
        .CK(npu_inst_pe_1_0_7_net4138), .RN(npu_inst_pe_1_0_7_n11), .Q(
        npu_inst_pe_1_0_7_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_0_7_n96), 
        .CK(npu_inst_pe_1_0_7_net4138), .RN(npu_inst_pe_1_0_7_n11), .Q(
        npu_inst_pe_1_0_7_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_0_7_n97), 
        .CK(npu_inst_pe_1_0_7_net4138), .RN(npu_inst_pe_1_0_7_n11), .Q(
        npu_inst_pe_1_0_7_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_0_7_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_0_7_N84), .SE(1'b0), .GCK(npu_inst_pe_1_0_7_net4132) );
  CLKGATETST_X1 npu_inst_pe_1_0_7_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n66), .SE(1'b0), .GCK(npu_inst_pe_1_0_7_net4138) );
  MUX2_X1 npu_inst_pe_1_1_0_U162 ( .A(npu_inst_pe_1_1_0_n32), .B(
        npu_inst_pe_1_1_0_n29), .S(npu_inst_pe_1_1_0_n8), .Z(
        npu_inst_pe_1_1_0_N93) );
  MUX2_X1 npu_inst_pe_1_1_0_U161 ( .A(npu_inst_pe_1_1_0_n31), .B(
        npu_inst_pe_1_1_0_n30), .S(npu_inst_pe_1_1_0_n6), .Z(
        npu_inst_pe_1_1_0_n32) );
  MUX2_X1 npu_inst_pe_1_1_0_U160 ( .A(npu_inst_pe_1_1_0_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_1_0_int_q_reg_v_1__0_), .S(npu_inst_pe_1_1_0_n4), .Z(
        npu_inst_pe_1_1_0_n31) );
  MUX2_X1 npu_inst_pe_1_1_0_U159 ( .A(npu_inst_pe_1_1_0_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_1_0_int_q_reg_v_3__0_), .S(npu_inst_pe_1_1_0_n4), .Z(
        npu_inst_pe_1_1_0_n30) );
  MUX2_X1 npu_inst_pe_1_1_0_U158 ( .A(npu_inst_pe_1_1_0_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_1_0_int_q_reg_v_5__0_), .S(npu_inst_pe_1_1_0_n4), .Z(
        npu_inst_pe_1_1_0_n29) );
  MUX2_X1 npu_inst_pe_1_1_0_U157 ( .A(npu_inst_pe_1_1_0_n28), .B(
        npu_inst_pe_1_1_0_n23), .S(npu_inst_pe_1_1_0_n8), .Z(
        npu_inst_pe_1_1_0_N94) );
  MUX2_X1 npu_inst_pe_1_1_0_U156 ( .A(npu_inst_pe_1_1_0_n25), .B(
        npu_inst_pe_1_1_0_n24), .S(npu_inst_pe_1_1_0_n6), .Z(
        npu_inst_pe_1_1_0_n28) );
  MUX2_X1 npu_inst_pe_1_1_0_U155 ( .A(npu_inst_pe_1_1_0_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_1_0_int_q_reg_v_1__1_), .S(npu_inst_pe_1_1_0_n4), .Z(
        npu_inst_pe_1_1_0_n25) );
  MUX2_X1 npu_inst_pe_1_1_0_U154 ( .A(npu_inst_pe_1_1_0_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_1_0_int_q_reg_v_3__1_), .S(npu_inst_pe_1_1_0_n4), .Z(
        npu_inst_pe_1_1_0_n24) );
  MUX2_X1 npu_inst_pe_1_1_0_U153 ( .A(npu_inst_pe_1_1_0_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_1_0_int_q_reg_v_5__1_), .S(npu_inst_pe_1_1_0_n4), .Z(
        npu_inst_pe_1_1_0_n23) );
  MUX2_X1 npu_inst_pe_1_1_0_U152 ( .A(npu_inst_pe_1_1_0_n22), .B(
        npu_inst_pe_1_1_0_n19), .S(npu_inst_pe_1_1_0_n8), .Z(
        npu_inst_pe_1_1_0_o_data_h_1_) );
  MUX2_X1 npu_inst_pe_1_1_0_U151 ( .A(npu_inst_pe_1_1_0_n21), .B(
        npu_inst_pe_1_1_0_n20), .S(npu_inst_pe_1_1_0_n6), .Z(
        npu_inst_pe_1_1_0_n22) );
  MUX2_X1 npu_inst_pe_1_1_0_U150 ( .A(npu_inst_pe_1_1_0_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_1_0_int_q_reg_h_1__1_), .S(npu_inst_pe_1_1_0_n4), .Z(
        npu_inst_pe_1_1_0_n21) );
  MUX2_X1 npu_inst_pe_1_1_0_U149 ( .A(npu_inst_pe_1_1_0_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_1_0_int_q_reg_h_3__1_), .S(npu_inst_pe_1_1_0_n4), .Z(
        npu_inst_pe_1_1_0_n20) );
  MUX2_X1 npu_inst_pe_1_1_0_U148 ( .A(npu_inst_pe_1_1_0_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_1_0_int_q_reg_h_5__1_), .S(npu_inst_pe_1_1_0_n4), .Z(
        npu_inst_pe_1_1_0_n19) );
  MUX2_X1 npu_inst_pe_1_1_0_U147 ( .A(npu_inst_pe_1_1_0_n18), .B(
        npu_inst_pe_1_1_0_n15), .S(npu_inst_pe_1_1_0_n8), .Z(
        npu_inst_pe_1_1_0_o_data_h_0_) );
  MUX2_X1 npu_inst_pe_1_1_0_U146 ( .A(npu_inst_pe_1_1_0_n17), .B(
        npu_inst_pe_1_1_0_n16), .S(npu_inst_pe_1_1_0_n6), .Z(
        npu_inst_pe_1_1_0_n18) );
  MUX2_X1 npu_inst_pe_1_1_0_U145 ( .A(npu_inst_pe_1_1_0_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_1_0_int_q_reg_h_1__0_), .S(npu_inst_pe_1_1_0_n4), .Z(
        npu_inst_pe_1_1_0_n17) );
  MUX2_X1 npu_inst_pe_1_1_0_U144 ( .A(npu_inst_pe_1_1_0_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_1_0_int_q_reg_h_3__0_), .S(npu_inst_pe_1_1_0_n4), .Z(
        npu_inst_pe_1_1_0_n16) );
  MUX2_X1 npu_inst_pe_1_1_0_U143 ( .A(npu_inst_pe_1_1_0_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_1_0_int_q_reg_h_5__0_), .S(npu_inst_pe_1_1_0_n4), .Z(
        npu_inst_pe_1_1_0_n15) );
  XOR2_X1 npu_inst_pe_1_1_0_U142 ( .A(npu_inst_pe_1_1_0_int_data_0_), .B(
        npu_inst_pe_1_1_0_int_q_acc_0_), .Z(npu_inst_pe_1_1_0_N73) );
  AND2_X1 npu_inst_pe_1_1_0_U141 ( .A1(npu_inst_pe_1_1_0_int_q_acc_0_), .A2(
        npu_inst_pe_1_1_0_int_data_0_), .ZN(npu_inst_pe_1_1_0_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_1_0_U140 ( .A(npu_inst_pe_1_1_0_int_q_acc_0_), .B(
        npu_inst_pe_1_1_0_n13), .ZN(npu_inst_pe_1_1_0_N65) );
  OR2_X1 npu_inst_pe_1_1_0_U139 ( .A1(npu_inst_pe_1_1_0_n13), .A2(
        npu_inst_pe_1_1_0_int_q_acc_0_), .ZN(npu_inst_pe_1_1_0_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_1_0_U138 ( .A(npu_inst_pe_1_1_0_int_q_acc_2_), .B(
        npu_inst_pe_1_1_0_add_79_carry_2_), .Z(npu_inst_pe_1_1_0_N75) );
  AND2_X1 npu_inst_pe_1_1_0_U137 ( .A1(npu_inst_pe_1_1_0_add_79_carry_2_), 
        .A2(npu_inst_pe_1_1_0_int_q_acc_2_), .ZN(
        npu_inst_pe_1_1_0_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_1_0_U136 ( .A(npu_inst_pe_1_1_0_int_q_acc_3_), .B(
        npu_inst_pe_1_1_0_add_79_carry_3_), .Z(npu_inst_pe_1_1_0_N76) );
  AND2_X1 npu_inst_pe_1_1_0_U135 ( .A1(npu_inst_pe_1_1_0_add_79_carry_3_), 
        .A2(npu_inst_pe_1_1_0_int_q_acc_3_), .ZN(
        npu_inst_pe_1_1_0_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_1_0_U134 ( .A(npu_inst_pe_1_1_0_int_q_acc_4_), .B(
        npu_inst_pe_1_1_0_add_79_carry_4_), .Z(npu_inst_pe_1_1_0_N77) );
  AND2_X1 npu_inst_pe_1_1_0_U133 ( .A1(npu_inst_pe_1_1_0_add_79_carry_4_), 
        .A2(npu_inst_pe_1_1_0_int_q_acc_4_), .ZN(
        npu_inst_pe_1_1_0_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_1_0_U132 ( .A(npu_inst_pe_1_1_0_int_q_acc_5_), .B(
        npu_inst_pe_1_1_0_add_79_carry_5_), .Z(npu_inst_pe_1_1_0_N78) );
  AND2_X1 npu_inst_pe_1_1_0_U131 ( .A1(npu_inst_pe_1_1_0_add_79_carry_5_), 
        .A2(npu_inst_pe_1_1_0_int_q_acc_5_), .ZN(
        npu_inst_pe_1_1_0_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_1_0_U130 ( .A(npu_inst_pe_1_1_0_int_q_acc_6_), .B(
        npu_inst_pe_1_1_0_add_79_carry_6_), .Z(npu_inst_pe_1_1_0_N79) );
  AND2_X1 npu_inst_pe_1_1_0_U129 ( .A1(npu_inst_pe_1_1_0_add_79_carry_6_), 
        .A2(npu_inst_pe_1_1_0_int_q_acc_6_), .ZN(
        npu_inst_pe_1_1_0_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_1_0_U128 ( .A(npu_inst_pe_1_1_0_int_q_acc_7_), .B(
        npu_inst_pe_1_1_0_add_79_carry_7_), .Z(npu_inst_pe_1_1_0_N80) );
  XNOR2_X1 npu_inst_pe_1_1_0_U127 ( .A(npu_inst_pe_1_1_0_sub_77_carry_2_), .B(
        npu_inst_pe_1_1_0_int_q_acc_2_), .ZN(npu_inst_pe_1_1_0_N67) );
  OR2_X1 npu_inst_pe_1_1_0_U126 ( .A1(npu_inst_pe_1_1_0_int_q_acc_2_), .A2(
        npu_inst_pe_1_1_0_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_1_0_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_1_0_U125 ( .A(npu_inst_pe_1_1_0_sub_77_carry_3_), .B(
        npu_inst_pe_1_1_0_int_q_acc_3_), .ZN(npu_inst_pe_1_1_0_N68) );
  OR2_X1 npu_inst_pe_1_1_0_U124 ( .A1(npu_inst_pe_1_1_0_int_q_acc_3_), .A2(
        npu_inst_pe_1_1_0_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_1_0_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_1_0_U123 ( .A(npu_inst_pe_1_1_0_sub_77_carry_4_), .B(
        npu_inst_pe_1_1_0_int_q_acc_4_), .ZN(npu_inst_pe_1_1_0_N69) );
  OR2_X1 npu_inst_pe_1_1_0_U122 ( .A1(npu_inst_pe_1_1_0_int_q_acc_4_), .A2(
        npu_inst_pe_1_1_0_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_1_0_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_1_0_U121 ( .A(npu_inst_pe_1_1_0_sub_77_carry_5_), .B(
        npu_inst_pe_1_1_0_int_q_acc_5_), .ZN(npu_inst_pe_1_1_0_N70) );
  OR2_X1 npu_inst_pe_1_1_0_U120 ( .A1(npu_inst_pe_1_1_0_int_q_acc_5_), .A2(
        npu_inst_pe_1_1_0_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_1_0_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_1_0_U119 ( .A(npu_inst_pe_1_1_0_sub_77_carry_6_), .B(
        npu_inst_pe_1_1_0_int_q_acc_6_), .ZN(npu_inst_pe_1_1_0_N71) );
  OR2_X1 npu_inst_pe_1_1_0_U118 ( .A1(npu_inst_pe_1_1_0_int_q_acc_6_), .A2(
        npu_inst_pe_1_1_0_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_1_0_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_1_0_U117 ( .A(npu_inst_pe_1_1_0_int_q_acc_7_), .B(
        npu_inst_pe_1_1_0_sub_77_carry_7_), .ZN(npu_inst_pe_1_1_0_N72) );
  INV_X1 npu_inst_pe_1_1_0_U116 ( .A(npu_inst_n79), .ZN(npu_inst_pe_1_1_0_n7)
         );
  INV_X1 npu_inst_pe_1_1_0_U115 ( .A(npu_inst_pe_1_1_0_n7), .ZN(
        npu_inst_pe_1_1_0_n6) );
  INV_X1 npu_inst_pe_1_1_0_U114 ( .A(npu_inst_n59), .ZN(npu_inst_pe_1_1_0_n3)
         );
  AOI22_X1 npu_inst_pe_1_1_0_U113 ( .A1(npu_inst_int_data_y_2__0__0_), .A2(
        npu_inst_pe_1_1_0_n58), .B1(npu_inst_pe_1_1_0_n114), .B2(
        npu_inst_pe_1_1_0_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_1_0_n57) );
  INV_X1 npu_inst_pe_1_1_0_U112 ( .A(npu_inst_pe_1_1_0_n57), .ZN(
        npu_inst_pe_1_1_0_n108) );
  AOI22_X1 npu_inst_pe_1_1_0_U111 ( .A1(npu_inst_int_data_y_2__0__0_), .A2(
        npu_inst_pe_1_1_0_n54), .B1(npu_inst_pe_1_1_0_n115), .B2(
        npu_inst_pe_1_1_0_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_1_0_n53) );
  INV_X1 npu_inst_pe_1_1_0_U110 ( .A(npu_inst_pe_1_1_0_n53), .ZN(
        npu_inst_pe_1_1_0_n109) );
  AOI22_X1 npu_inst_pe_1_1_0_U107 ( .A1(npu_inst_int_data_y_2__0__0_), .A2(
        npu_inst_pe_1_1_0_n50), .B1(npu_inst_pe_1_1_0_n116), .B2(
        npu_inst_pe_1_1_0_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_1_0_n49) );
  INV_X1 npu_inst_pe_1_1_0_U106 ( .A(npu_inst_pe_1_1_0_n49), .ZN(
        npu_inst_pe_1_1_0_n110) );
  AOI22_X1 npu_inst_pe_1_1_0_U105 ( .A1(npu_inst_int_data_y_2__0__0_), .A2(
        npu_inst_pe_1_1_0_n46), .B1(npu_inst_pe_1_1_0_n117), .B2(
        npu_inst_pe_1_1_0_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_1_0_n45) );
  INV_X1 npu_inst_pe_1_1_0_U104 ( .A(npu_inst_pe_1_1_0_n45), .ZN(
        npu_inst_pe_1_1_0_n111) );
  AOI22_X1 npu_inst_pe_1_1_0_U103 ( .A1(npu_inst_int_data_y_2__0__0_), .A2(
        npu_inst_pe_1_1_0_n42), .B1(npu_inst_pe_1_1_0_n119), .B2(
        npu_inst_pe_1_1_0_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_1_0_n41) );
  INV_X1 npu_inst_pe_1_1_0_U102 ( .A(npu_inst_pe_1_1_0_n41), .ZN(
        npu_inst_pe_1_1_0_n112) );
  AOI22_X1 npu_inst_pe_1_1_0_U101 ( .A1(npu_inst_int_data_y_2__0__1_), .A2(
        npu_inst_pe_1_1_0_n58), .B1(npu_inst_pe_1_1_0_n114), .B2(
        npu_inst_pe_1_1_0_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_1_0_n59) );
  INV_X1 npu_inst_pe_1_1_0_U100 ( .A(npu_inst_pe_1_1_0_n59), .ZN(
        npu_inst_pe_1_1_0_n102) );
  AOI22_X1 npu_inst_pe_1_1_0_U99 ( .A1(npu_inst_int_data_y_2__0__1_), .A2(
        npu_inst_pe_1_1_0_n54), .B1(npu_inst_pe_1_1_0_n115), .B2(
        npu_inst_pe_1_1_0_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_1_0_n55) );
  INV_X1 npu_inst_pe_1_1_0_U98 ( .A(npu_inst_pe_1_1_0_n55), .ZN(
        npu_inst_pe_1_1_0_n103) );
  AOI22_X1 npu_inst_pe_1_1_0_U97 ( .A1(npu_inst_int_data_y_2__0__1_), .A2(
        npu_inst_pe_1_1_0_n50), .B1(npu_inst_pe_1_1_0_n116), .B2(
        npu_inst_pe_1_1_0_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_1_0_n51) );
  INV_X1 npu_inst_pe_1_1_0_U96 ( .A(npu_inst_pe_1_1_0_n51), .ZN(
        npu_inst_pe_1_1_0_n104) );
  AOI22_X1 npu_inst_pe_1_1_0_U95 ( .A1(npu_inst_int_data_y_2__0__1_), .A2(
        npu_inst_pe_1_1_0_n46), .B1(npu_inst_pe_1_1_0_n117), .B2(
        npu_inst_pe_1_1_0_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_1_0_n47) );
  INV_X1 npu_inst_pe_1_1_0_U94 ( .A(npu_inst_pe_1_1_0_n47), .ZN(
        npu_inst_pe_1_1_0_n105) );
  AOI22_X1 npu_inst_pe_1_1_0_U93 ( .A1(npu_inst_int_data_y_2__0__1_), .A2(
        npu_inst_pe_1_1_0_n42), .B1(npu_inst_pe_1_1_0_n119), .B2(
        npu_inst_pe_1_1_0_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_1_0_n43) );
  INV_X1 npu_inst_pe_1_1_0_U92 ( .A(npu_inst_pe_1_1_0_n43), .ZN(
        npu_inst_pe_1_1_0_n106) );
  AOI22_X1 npu_inst_pe_1_1_0_U91 ( .A1(npu_inst_pe_1_1_0_n38), .A2(
        npu_inst_int_data_y_2__0__1_), .B1(npu_inst_pe_1_1_0_n118), .B2(
        npu_inst_pe_1_1_0_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_1_0_n39) );
  INV_X1 npu_inst_pe_1_1_0_U90 ( .A(npu_inst_pe_1_1_0_n39), .ZN(
        npu_inst_pe_1_1_0_n107) );
  AOI22_X1 npu_inst_pe_1_1_0_U89 ( .A1(npu_inst_pe_1_1_0_n38), .A2(
        npu_inst_int_data_y_2__0__0_), .B1(npu_inst_pe_1_1_0_n118), .B2(
        npu_inst_pe_1_1_0_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_1_0_n37) );
  INV_X1 npu_inst_pe_1_1_0_U88 ( .A(npu_inst_pe_1_1_0_n37), .ZN(
        npu_inst_pe_1_1_0_n113) );
  NAND2_X1 npu_inst_pe_1_1_0_U87 ( .A1(npu_inst_pe_1_1_0_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_1_0_n60), .ZN(npu_inst_pe_1_1_0_n74) );
  OAI21_X1 npu_inst_pe_1_1_0_U86 ( .B1(npu_inst_pe_1_1_0_n63), .B2(
        npu_inst_pe_1_1_0_n60), .A(npu_inst_pe_1_1_0_n74), .ZN(
        npu_inst_pe_1_1_0_n97) );
  NAND2_X1 npu_inst_pe_1_1_0_U85 ( .A1(npu_inst_pe_1_1_0_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_1_0_n60), .ZN(npu_inst_pe_1_1_0_n73) );
  OAI21_X1 npu_inst_pe_1_1_0_U84 ( .B1(npu_inst_pe_1_1_0_n61), .B2(
        npu_inst_pe_1_1_0_n60), .A(npu_inst_pe_1_1_0_n73), .ZN(
        npu_inst_pe_1_1_0_n96) );
  NAND2_X1 npu_inst_pe_1_1_0_U83 ( .A1(npu_inst_pe_1_1_0_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_1_0_n56), .ZN(npu_inst_pe_1_1_0_n72) );
  OAI21_X1 npu_inst_pe_1_1_0_U82 ( .B1(npu_inst_pe_1_1_0_n63), .B2(
        npu_inst_pe_1_1_0_n56), .A(npu_inst_pe_1_1_0_n72), .ZN(
        npu_inst_pe_1_1_0_n95) );
  NAND2_X1 npu_inst_pe_1_1_0_U81 ( .A1(npu_inst_pe_1_1_0_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_1_0_n56), .ZN(npu_inst_pe_1_1_0_n71) );
  OAI21_X1 npu_inst_pe_1_1_0_U80 ( .B1(npu_inst_pe_1_1_0_n61), .B2(
        npu_inst_pe_1_1_0_n56), .A(npu_inst_pe_1_1_0_n71), .ZN(
        npu_inst_pe_1_1_0_n94) );
  NAND2_X1 npu_inst_pe_1_1_0_U79 ( .A1(npu_inst_pe_1_1_0_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_1_0_n52), .ZN(npu_inst_pe_1_1_0_n70) );
  OAI21_X1 npu_inst_pe_1_1_0_U78 ( .B1(npu_inst_pe_1_1_0_n63), .B2(
        npu_inst_pe_1_1_0_n52), .A(npu_inst_pe_1_1_0_n70), .ZN(
        npu_inst_pe_1_1_0_n93) );
  NAND2_X1 npu_inst_pe_1_1_0_U77 ( .A1(npu_inst_pe_1_1_0_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_1_0_n52), .ZN(npu_inst_pe_1_1_0_n69) );
  OAI21_X1 npu_inst_pe_1_1_0_U76 ( .B1(npu_inst_pe_1_1_0_n61), .B2(
        npu_inst_pe_1_1_0_n52), .A(npu_inst_pe_1_1_0_n69), .ZN(
        npu_inst_pe_1_1_0_n92) );
  NAND2_X1 npu_inst_pe_1_1_0_U75 ( .A1(npu_inst_pe_1_1_0_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_1_0_n48), .ZN(npu_inst_pe_1_1_0_n68) );
  OAI21_X1 npu_inst_pe_1_1_0_U74 ( .B1(npu_inst_pe_1_1_0_n63), .B2(
        npu_inst_pe_1_1_0_n48), .A(npu_inst_pe_1_1_0_n68), .ZN(
        npu_inst_pe_1_1_0_n91) );
  NAND2_X1 npu_inst_pe_1_1_0_U73 ( .A1(npu_inst_pe_1_1_0_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_1_0_n48), .ZN(npu_inst_pe_1_1_0_n67) );
  OAI21_X1 npu_inst_pe_1_1_0_U72 ( .B1(npu_inst_pe_1_1_0_n61), .B2(
        npu_inst_pe_1_1_0_n48), .A(npu_inst_pe_1_1_0_n67), .ZN(
        npu_inst_pe_1_1_0_n90) );
  NAND2_X1 npu_inst_pe_1_1_0_U71 ( .A1(npu_inst_pe_1_1_0_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_1_0_n44), .ZN(npu_inst_pe_1_1_0_n66) );
  OAI21_X1 npu_inst_pe_1_1_0_U70 ( .B1(npu_inst_pe_1_1_0_n63), .B2(
        npu_inst_pe_1_1_0_n44), .A(npu_inst_pe_1_1_0_n66), .ZN(
        npu_inst_pe_1_1_0_n89) );
  NAND2_X1 npu_inst_pe_1_1_0_U69 ( .A1(npu_inst_pe_1_1_0_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_1_0_n44), .ZN(npu_inst_pe_1_1_0_n65) );
  OAI21_X1 npu_inst_pe_1_1_0_U68 ( .B1(npu_inst_pe_1_1_0_n61), .B2(
        npu_inst_pe_1_1_0_n44), .A(npu_inst_pe_1_1_0_n65), .ZN(
        npu_inst_pe_1_1_0_n88) );
  NAND2_X1 npu_inst_pe_1_1_0_U67 ( .A1(npu_inst_pe_1_1_0_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_1_0_n40), .ZN(npu_inst_pe_1_1_0_n64) );
  OAI21_X1 npu_inst_pe_1_1_0_U66 ( .B1(npu_inst_pe_1_1_0_n63), .B2(
        npu_inst_pe_1_1_0_n40), .A(npu_inst_pe_1_1_0_n64), .ZN(
        npu_inst_pe_1_1_0_n87) );
  NAND2_X1 npu_inst_pe_1_1_0_U65 ( .A1(npu_inst_pe_1_1_0_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_1_0_n40), .ZN(npu_inst_pe_1_1_0_n62) );
  OAI21_X1 npu_inst_pe_1_1_0_U64 ( .B1(npu_inst_pe_1_1_0_n61), .B2(
        npu_inst_pe_1_1_0_n40), .A(npu_inst_pe_1_1_0_n62), .ZN(
        npu_inst_pe_1_1_0_n86) );
  AND2_X1 npu_inst_pe_1_1_0_U63 ( .A1(npu_inst_pe_1_1_0_N93), .A2(npu_inst_n59), .ZN(npu_inst_int_data_y_1__0__0_) );
  AND2_X1 npu_inst_pe_1_1_0_U62 ( .A1(npu_inst_n59), .A2(npu_inst_pe_1_1_0_N94), .ZN(npu_inst_int_data_y_1__0__1_) );
  NOR3_X1 npu_inst_pe_1_1_0_U61 ( .A1(npu_inst_pe_1_1_0_n26), .A2(npu_inst_n59), .A3(npu_inst_int_ckg[55]), .ZN(npu_inst_pe_1_1_0_n85) );
  OR2_X1 npu_inst_pe_1_1_0_U60 ( .A1(npu_inst_pe_1_1_0_n85), .A2(
        npu_inst_pe_1_1_0_n2), .ZN(npu_inst_pe_1_1_0_N84) );
  AND2_X1 npu_inst_pe_1_1_0_U59 ( .A1(npu_inst_pe_1_1_0_int_q_acc_0_), .A2(
        npu_inst_pe_1_1_0_n1), .ZN(npu_inst_int_data_res_1__0__0_) );
  AND2_X1 npu_inst_pe_1_1_0_U58 ( .A1(npu_inst_pe_1_1_0_n2), .A2(
        npu_inst_pe_1_1_0_int_q_acc_7_), .ZN(npu_inst_int_data_res_1__0__7_)
         );
  AND2_X1 npu_inst_pe_1_1_0_U57 ( .A1(npu_inst_pe_1_1_0_int_q_acc_1_), .A2(
        npu_inst_pe_1_1_0_n1), .ZN(npu_inst_int_data_res_1__0__1_) );
  AND2_X1 npu_inst_pe_1_1_0_U56 ( .A1(npu_inst_pe_1_1_0_int_q_acc_2_), .A2(
        npu_inst_pe_1_1_0_n1), .ZN(npu_inst_int_data_res_1__0__2_) );
  AND2_X1 npu_inst_pe_1_1_0_U55 ( .A1(npu_inst_pe_1_1_0_int_q_acc_3_), .A2(
        npu_inst_pe_1_1_0_n2), .ZN(npu_inst_int_data_res_1__0__3_) );
  AND2_X1 npu_inst_pe_1_1_0_U54 ( .A1(npu_inst_pe_1_1_0_int_q_acc_4_), .A2(
        npu_inst_pe_1_1_0_n2), .ZN(npu_inst_int_data_res_1__0__4_) );
  AND2_X1 npu_inst_pe_1_1_0_U53 ( .A1(npu_inst_pe_1_1_0_int_q_acc_5_), .A2(
        npu_inst_pe_1_1_0_n2), .ZN(npu_inst_int_data_res_1__0__5_) );
  AND2_X1 npu_inst_pe_1_1_0_U52 ( .A1(npu_inst_pe_1_1_0_int_q_acc_6_), .A2(
        npu_inst_pe_1_1_0_n2), .ZN(npu_inst_int_data_res_1__0__6_) );
  AOI222_X1 npu_inst_pe_1_1_0_U51 ( .A1(npu_inst_int_data_res_2__0__0_), .A2(
        npu_inst_pe_1_1_0_n1), .B1(npu_inst_pe_1_1_0_N73), .B2(
        npu_inst_pe_1_1_0_n76), .C1(npu_inst_pe_1_1_0_N65), .C2(
        npu_inst_pe_1_1_0_n77), .ZN(npu_inst_pe_1_1_0_n84) );
  INV_X1 npu_inst_pe_1_1_0_U50 ( .A(npu_inst_pe_1_1_0_n84), .ZN(
        npu_inst_pe_1_1_0_n101) );
  AOI222_X1 npu_inst_pe_1_1_0_U49 ( .A1(npu_inst_int_data_res_2__0__7_), .A2(
        npu_inst_pe_1_1_0_n1), .B1(npu_inst_pe_1_1_0_N80), .B2(
        npu_inst_pe_1_1_0_n76), .C1(npu_inst_pe_1_1_0_N72), .C2(
        npu_inst_pe_1_1_0_n77), .ZN(npu_inst_pe_1_1_0_n75) );
  INV_X1 npu_inst_pe_1_1_0_U48 ( .A(npu_inst_pe_1_1_0_n75), .ZN(
        npu_inst_pe_1_1_0_n33) );
  AOI222_X1 npu_inst_pe_1_1_0_U47 ( .A1(npu_inst_int_data_res_2__0__1_), .A2(
        npu_inst_pe_1_1_0_n1), .B1(npu_inst_pe_1_1_0_N74), .B2(
        npu_inst_pe_1_1_0_n76), .C1(npu_inst_pe_1_1_0_N66), .C2(
        npu_inst_pe_1_1_0_n77), .ZN(npu_inst_pe_1_1_0_n83) );
  INV_X1 npu_inst_pe_1_1_0_U46 ( .A(npu_inst_pe_1_1_0_n83), .ZN(
        npu_inst_pe_1_1_0_n100) );
  AOI222_X1 npu_inst_pe_1_1_0_U45 ( .A1(npu_inst_int_data_res_2__0__2_), .A2(
        npu_inst_pe_1_1_0_n1), .B1(npu_inst_pe_1_1_0_N75), .B2(
        npu_inst_pe_1_1_0_n76), .C1(npu_inst_pe_1_1_0_N67), .C2(
        npu_inst_pe_1_1_0_n77), .ZN(npu_inst_pe_1_1_0_n82) );
  INV_X1 npu_inst_pe_1_1_0_U44 ( .A(npu_inst_pe_1_1_0_n82), .ZN(
        npu_inst_pe_1_1_0_n99) );
  AOI222_X1 npu_inst_pe_1_1_0_U43 ( .A1(npu_inst_int_data_res_2__0__3_), .A2(
        npu_inst_pe_1_1_0_n1), .B1(npu_inst_pe_1_1_0_N76), .B2(
        npu_inst_pe_1_1_0_n76), .C1(npu_inst_pe_1_1_0_N68), .C2(
        npu_inst_pe_1_1_0_n77), .ZN(npu_inst_pe_1_1_0_n81) );
  INV_X1 npu_inst_pe_1_1_0_U42 ( .A(npu_inst_pe_1_1_0_n81), .ZN(
        npu_inst_pe_1_1_0_n98) );
  AOI222_X1 npu_inst_pe_1_1_0_U41 ( .A1(npu_inst_int_data_res_2__0__4_), .A2(
        npu_inst_pe_1_1_0_n1), .B1(npu_inst_pe_1_1_0_N77), .B2(
        npu_inst_pe_1_1_0_n76), .C1(npu_inst_pe_1_1_0_N69), .C2(
        npu_inst_pe_1_1_0_n77), .ZN(npu_inst_pe_1_1_0_n80) );
  INV_X1 npu_inst_pe_1_1_0_U40 ( .A(npu_inst_pe_1_1_0_n80), .ZN(
        npu_inst_pe_1_1_0_n36) );
  AOI222_X1 npu_inst_pe_1_1_0_U39 ( .A1(npu_inst_int_data_res_2__0__5_), .A2(
        npu_inst_pe_1_1_0_n1), .B1(npu_inst_pe_1_1_0_N78), .B2(
        npu_inst_pe_1_1_0_n76), .C1(npu_inst_pe_1_1_0_N70), .C2(
        npu_inst_pe_1_1_0_n77), .ZN(npu_inst_pe_1_1_0_n79) );
  INV_X1 npu_inst_pe_1_1_0_U38 ( .A(npu_inst_pe_1_1_0_n79), .ZN(
        npu_inst_pe_1_1_0_n35) );
  AOI222_X1 npu_inst_pe_1_1_0_U37 ( .A1(npu_inst_int_data_res_2__0__6_), .A2(
        npu_inst_pe_1_1_0_n1), .B1(npu_inst_pe_1_1_0_N79), .B2(
        npu_inst_pe_1_1_0_n76), .C1(npu_inst_pe_1_1_0_N71), .C2(
        npu_inst_pe_1_1_0_n77), .ZN(npu_inst_pe_1_1_0_n78) );
  INV_X1 npu_inst_pe_1_1_0_U36 ( .A(npu_inst_pe_1_1_0_n78), .ZN(
        npu_inst_pe_1_1_0_n34) );
  AND2_X1 npu_inst_pe_1_1_0_U35 ( .A1(npu_inst_pe_1_1_0_o_data_h_1_), .A2(
        npu_inst_pe_1_1_0_int_q_weight_1_), .ZN(npu_inst_pe_1_1_0_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_1_0_U34 ( .A1(npu_inst_pe_1_1_0_o_data_h_0_), .A2(
        npu_inst_pe_1_1_0_int_q_weight_1_), .ZN(npu_inst_pe_1_1_0_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_1_0_U33 ( .A(npu_inst_pe_1_1_0_int_data_1_), .ZN(
        npu_inst_pe_1_1_0_n14) );
  AOI22_X1 npu_inst_pe_1_1_0_U32 ( .A1(npu_inst_n59), .A2(
        npu_inst_int_data_y_2__0__1_), .B1(npu_inst_pe_1_1_0_n3), .B2(
        npu_inst_int_data_x_1__1__1_), .ZN(npu_inst_pe_1_1_0_n63) );
  AOI22_X1 npu_inst_pe_1_1_0_U31 ( .A1(npu_inst_n59), .A2(
        npu_inst_int_data_y_2__0__0_), .B1(npu_inst_pe_1_1_0_n3), .B2(
        npu_inst_int_data_x_1__1__0_), .ZN(npu_inst_pe_1_1_0_n61) );
  INV_X1 npu_inst_pe_1_1_0_U30 ( .A(npu_inst_pe_1_1_0_int_data_0_), .ZN(
        npu_inst_pe_1_1_0_n13) );
  INV_X1 npu_inst_pe_1_1_0_U29 ( .A(npu_inst_n71), .ZN(npu_inst_pe_1_1_0_n5)
         );
  OR3_X1 npu_inst_pe_1_1_0_U28 ( .A1(npu_inst_pe_1_1_0_n6), .A2(
        npu_inst_pe_1_1_0_n8), .A3(npu_inst_pe_1_1_0_n5), .ZN(
        npu_inst_pe_1_1_0_n56) );
  OR3_X1 npu_inst_pe_1_1_0_U27 ( .A1(npu_inst_pe_1_1_0_n5), .A2(
        npu_inst_pe_1_1_0_n8), .A3(npu_inst_pe_1_1_0_n7), .ZN(
        npu_inst_pe_1_1_0_n48) );
  INV_X1 npu_inst_pe_1_1_0_U26 ( .A(npu_inst_pe_1_1_0_n5), .ZN(
        npu_inst_pe_1_1_0_n4) );
  INV_X1 npu_inst_pe_1_1_0_U25 ( .A(npu_inst_n126), .ZN(npu_inst_pe_1_1_0_n12)
         );
  OR3_X1 npu_inst_pe_1_1_0_U24 ( .A1(npu_inst_pe_1_1_0_n4), .A2(
        npu_inst_pe_1_1_0_n8), .A3(npu_inst_pe_1_1_0_n7), .ZN(
        npu_inst_pe_1_1_0_n52) );
  OR3_X1 npu_inst_pe_1_1_0_U23 ( .A1(npu_inst_pe_1_1_0_n6), .A2(
        npu_inst_pe_1_1_0_n8), .A3(npu_inst_pe_1_1_0_n4), .ZN(
        npu_inst_pe_1_1_0_n60) );
  NOR2_X1 npu_inst_pe_1_1_0_U22 ( .A1(npu_inst_pe_1_1_0_n60), .A2(
        npu_inst_pe_1_1_0_n3), .ZN(npu_inst_pe_1_1_0_n58) );
  NOR2_X1 npu_inst_pe_1_1_0_U21 ( .A1(npu_inst_pe_1_1_0_n56), .A2(
        npu_inst_pe_1_1_0_n3), .ZN(npu_inst_pe_1_1_0_n54) );
  NOR2_X1 npu_inst_pe_1_1_0_U20 ( .A1(npu_inst_pe_1_1_0_n52), .A2(
        npu_inst_pe_1_1_0_n3), .ZN(npu_inst_pe_1_1_0_n50) );
  NOR2_X1 npu_inst_pe_1_1_0_U19 ( .A1(npu_inst_pe_1_1_0_n48), .A2(
        npu_inst_pe_1_1_0_n3), .ZN(npu_inst_pe_1_1_0_n46) );
  NOR2_X1 npu_inst_pe_1_1_0_U18 ( .A1(npu_inst_pe_1_1_0_n40), .A2(
        npu_inst_pe_1_1_0_n3), .ZN(npu_inst_pe_1_1_0_n38) );
  NOR2_X1 npu_inst_pe_1_1_0_U17 ( .A1(npu_inst_pe_1_1_0_n44), .A2(
        npu_inst_pe_1_1_0_n3), .ZN(npu_inst_pe_1_1_0_n42) );
  BUF_X1 npu_inst_pe_1_1_0_U16 ( .A(npu_inst_n105), .Z(npu_inst_pe_1_1_0_n8)
         );
  BUF_X1 npu_inst_pe_1_1_0_U15 ( .A(npu_inst_pe_1_1_0_n12), .Z(
        npu_inst_pe_1_1_0_n11) );
  BUF_X1 npu_inst_pe_1_1_0_U14 ( .A(npu_inst_pe_1_1_0_n12), .Z(
        npu_inst_pe_1_1_0_n10) );
  BUF_X1 npu_inst_pe_1_1_0_U13 ( .A(npu_inst_pe_1_1_0_n12), .Z(
        npu_inst_pe_1_1_0_n9) );
  INV_X1 npu_inst_pe_1_1_0_U12 ( .A(npu_inst_pe_1_1_0_n38), .ZN(
        npu_inst_pe_1_1_0_n118) );
  INV_X1 npu_inst_pe_1_1_0_U11 ( .A(npu_inst_pe_1_1_0_n58), .ZN(
        npu_inst_pe_1_1_0_n114) );
  INV_X1 npu_inst_pe_1_1_0_U10 ( .A(npu_inst_pe_1_1_0_n54), .ZN(
        npu_inst_pe_1_1_0_n115) );
  INV_X1 npu_inst_pe_1_1_0_U9 ( .A(npu_inst_pe_1_1_0_n50), .ZN(
        npu_inst_pe_1_1_0_n116) );
  INV_X1 npu_inst_pe_1_1_0_U8 ( .A(npu_inst_pe_1_1_0_n46), .ZN(
        npu_inst_pe_1_1_0_n117) );
  INV_X1 npu_inst_pe_1_1_0_U7 ( .A(npu_inst_pe_1_1_0_n42), .ZN(
        npu_inst_pe_1_1_0_n119) );
  BUF_X1 npu_inst_pe_1_1_0_U6 ( .A(npu_inst_n34), .Z(npu_inst_pe_1_1_0_n2) );
  BUF_X1 npu_inst_pe_1_1_0_U5 ( .A(npu_inst_n34), .Z(npu_inst_pe_1_1_0_n1) );
  NOR2_X1 npu_inst_pe_1_1_0_U4 ( .A1(npu_inst_pe_1_1_0_int_q_weight_0_), .A2(
        npu_inst_pe_1_1_0_n1), .ZN(npu_inst_pe_1_1_0_n76) );
  NOR2_X1 npu_inst_pe_1_1_0_U3 ( .A1(npu_inst_pe_1_1_0_n27), .A2(
        npu_inst_pe_1_1_0_n1), .ZN(npu_inst_pe_1_1_0_n77) );
  FA_X1 npu_inst_pe_1_1_0_sub_77_U2_1 ( .A(npu_inst_pe_1_1_0_int_q_acc_1_), 
        .B(npu_inst_pe_1_1_0_n14), .CI(npu_inst_pe_1_1_0_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_1_0_sub_77_carry_2_), .S(npu_inst_pe_1_1_0_N66) );
  FA_X1 npu_inst_pe_1_1_0_add_79_U1_1 ( .A(npu_inst_pe_1_1_0_int_q_acc_1_), 
        .B(npu_inst_pe_1_1_0_int_data_1_), .CI(
        npu_inst_pe_1_1_0_add_79_carry_1_), .CO(
        npu_inst_pe_1_1_0_add_79_carry_2_), .S(npu_inst_pe_1_1_0_N74) );
  NAND3_X1 npu_inst_pe_1_1_0_U109 ( .A1(npu_inst_pe_1_1_0_n5), .A2(
        npu_inst_pe_1_1_0_n7), .A3(npu_inst_pe_1_1_0_n8), .ZN(
        npu_inst_pe_1_1_0_n44) );
  NAND3_X1 npu_inst_pe_1_1_0_U108 ( .A1(npu_inst_pe_1_1_0_n4), .A2(
        npu_inst_pe_1_1_0_n7), .A3(npu_inst_pe_1_1_0_n8), .ZN(
        npu_inst_pe_1_1_0_n40) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_1_0_n34), .CK(
        npu_inst_pe_1_1_0_net4109), .RN(npu_inst_pe_1_1_0_n9), .Q(
        npu_inst_pe_1_1_0_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_1_0_n35), .CK(
        npu_inst_pe_1_1_0_net4109), .RN(npu_inst_pe_1_1_0_n9), .Q(
        npu_inst_pe_1_1_0_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_1_0_n36), .CK(
        npu_inst_pe_1_1_0_net4109), .RN(npu_inst_pe_1_1_0_n9), .Q(
        npu_inst_pe_1_1_0_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_1_0_n98), .CK(
        npu_inst_pe_1_1_0_net4109), .RN(npu_inst_pe_1_1_0_n9), .Q(
        npu_inst_pe_1_1_0_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_1_0_n99), .CK(
        npu_inst_pe_1_1_0_net4109), .RN(npu_inst_pe_1_1_0_n9), .Q(
        npu_inst_pe_1_1_0_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_1_0_n100), 
        .CK(npu_inst_pe_1_1_0_net4109), .RN(npu_inst_pe_1_1_0_n9), .Q(
        npu_inst_pe_1_1_0_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_1_0_n33), .CK(
        npu_inst_pe_1_1_0_net4109), .RN(npu_inst_pe_1_1_0_n9), .Q(
        npu_inst_pe_1_1_0_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_1_0_n101), 
        .CK(npu_inst_pe_1_1_0_net4109), .RN(npu_inst_pe_1_1_0_n9), .Q(
        npu_inst_pe_1_1_0_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_weight_reg_0_ ( .D(npu_inst_n112), .CK(
        npu_inst_pe_1_1_0_net4115), .RN(npu_inst_pe_1_1_0_n9), .Q(
        npu_inst_pe_1_1_0_int_q_weight_0_), .QN(npu_inst_pe_1_1_0_n27) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_weight_reg_1_ ( .D(npu_inst_n118), .CK(
        npu_inst_pe_1_1_0_net4115), .RN(npu_inst_pe_1_1_0_n9), .Q(
        npu_inst_pe_1_1_0_int_q_weight_1_), .QN(npu_inst_pe_1_1_0_n26) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_1_0_n113), 
        .CK(npu_inst_pe_1_1_0_net4115), .RN(npu_inst_pe_1_1_0_n9), .Q(
        npu_inst_pe_1_1_0_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_1_0_n107), 
        .CK(npu_inst_pe_1_1_0_net4115), .RN(npu_inst_pe_1_1_0_n9), .Q(
        npu_inst_pe_1_1_0_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_1_0_n112), 
        .CK(npu_inst_pe_1_1_0_net4115), .RN(npu_inst_pe_1_1_0_n10), .Q(
        npu_inst_pe_1_1_0_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_1_0_n106), 
        .CK(npu_inst_pe_1_1_0_net4115), .RN(npu_inst_pe_1_1_0_n10), .Q(
        npu_inst_pe_1_1_0_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_1_0_n111), 
        .CK(npu_inst_pe_1_1_0_net4115), .RN(npu_inst_pe_1_1_0_n10), .Q(
        npu_inst_pe_1_1_0_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_1_0_n105), 
        .CK(npu_inst_pe_1_1_0_net4115), .RN(npu_inst_pe_1_1_0_n10), .Q(
        npu_inst_pe_1_1_0_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_1_0_n110), 
        .CK(npu_inst_pe_1_1_0_net4115), .RN(npu_inst_pe_1_1_0_n10), .Q(
        npu_inst_pe_1_1_0_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_1_0_n104), 
        .CK(npu_inst_pe_1_1_0_net4115), .RN(npu_inst_pe_1_1_0_n10), .Q(
        npu_inst_pe_1_1_0_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_1_0_n109), 
        .CK(npu_inst_pe_1_1_0_net4115), .RN(npu_inst_pe_1_1_0_n10), .Q(
        npu_inst_pe_1_1_0_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_1_0_n103), 
        .CK(npu_inst_pe_1_1_0_net4115), .RN(npu_inst_pe_1_1_0_n10), .Q(
        npu_inst_pe_1_1_0_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_1_0_n108), 
        .CK(npu_inst_pe_1_1_0_net4115), .RN(npu_inst_pe_1_1_0_n10), .Q(
        npu_inst_pe_1_1_0_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_1_0_n102), 
        .CK(npu_inst_pe_1_1_0_net4115), .RN(npu_inst_pe_1_1_0_n10), .Q(
        npu_inst_pe_1_1_0_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_1_0_n86), 
        .CK(npu_inst_pe_1_1_0_net4115), .RN(npu_inst_pe_1_1_0_n10), .Q(
        npu_inst_pe_1_1_0_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_1_0_n87), 
        .CK(npu_inst_pe_1_1_0_net4115), .RN(npu_inst_pe_1_1_0_n10), .Q(
        npu_inst_pe_1_1_0_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_1_0_n88), 
        .CK(npu_inst_pe_1_1_0_net4115), .RN(npu_inst_pe_1_1_0_n11), .Q(
        npu_inst_pe_1_1_0_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_1_0_n89), 
        .CK(npu_inst_pe_1_1_0_net4115), .RN(npu_inst_pe_1_1_0_n11), .Q(
        npu_inst_pe_1_1_0_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_1_0_n90), 
        .CK(npu_inst_pe_1_1_0_net4115), .RN(npu_inst_pe_1_1_0_n11), .Q(
        npu_inst_pe_1_1_0_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_1_0_n91), 
        .CK(npu_inst_pe_1_1_0_net4115), .RN(npu_inst_pe_1_1_0_n11), .Q(
        npu_inst_pe_1_1_0_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_1_0_n92), 
        .CK(npu_inst_pe_1_1_0_net4115), .RN(npu_inst_pe_1_1_0_n11), .Q(
        npu_inst_pe_1_1_0_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_1_0_n93), 
        .CK(npu_inst_pe_1_1_0_net4115), .RN(npu_inst_pe_1_1_0_n11), .Q(
        npu_inst_pe_1_1_0_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_1_0_n94), 
        .CK(npu_inst_pe_1_1_0_net4115), .RN(npu_inst_pe_1_1_0_n11), .Q(
        npu_inst_pe_1_1_0_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_1_0_n95), 
        .CK(npu_inst_pe_1_1_0_net4115), .RN(npu_inst_pe_1_1_0_n11), .Q(
        npu_inst_pe_1_1_0_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_1_0_n96), 
        .CK(npu_inst_pe_1_1_0_net4115), .RN(npu_inst_pe_1_1_0_n11), .Q(
        npu_inst_pe_1_1_0_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_1_0_n97), 
        .CK(npu_inst_pe_1_1_0_net4115), .RN(npu_inst_pe_1_1_0_n11), .Q(
        npu_inst_pe_1_1_0_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_1_0_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_1_0_N84), .SE(1'b0), .GCK(npu_inst_pe_1_1_0_net4109) );
  CLKGATETST_X1 npu_inst_pe_1_1_0_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n66), .SE(1'b0), .GCK(npu_inst_pe_1_1_0_net4115) );
  MUX2_X1 npu_inst_pe_1_1_1_U162 ( .A(npu_inst_pe_1_1_1_n32), .B(
        npu_inst_pe_1_1_1_n29), .S(npu_inst_pe_1_1_1_n8), .Z(
        npu_inst_pe_1_1_1_N93) );
  MUX2_X1 npu_inst_pe_1_1_1_U161 ( .A(npu_inst_pe_1_1_1_n31), .B(
        npu_inst_pe_1_1_1_n30), .S(npu_inst_pe_1_1_1_n6), .Z(
        npu_inst_pe_1_1_1_n32) );
  MUX2_X1 npu_inst_pe_1_1_1_U160 ( .A(npu_inst_pe_1_1_1_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_1_1_int_q_reg_v_1__0_), .S(npu_inst_pe_1_1_1_n4), .Z(
        npu_inst_pe_1_1_1_n31) );
  MUX2_X1 npu_inst_pe_1_1_1_U159 ( .A(npu_inst_pe_1_1_1_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_1_1_int_q_reg_v_3__0_), .S(npu_inst_pe_1_1_1_n4), .Z(
        npu_inst_pe_1_1_1_n30) );
  MUX2_X1 npu_inst_pe_1_1_1_U158 ( .A(npu_inst_pe_1_1_1_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_1_1_int_q_reg_v_5__0_), .S(npu_inst_pe_1_1_1_n4), .Z(
        npu_inst_pe_1_1_1_n29) );
  MUX2_X1 npu_inst_pe_1_1_1_U157 ( .A(npu_inst_pe_1_1_1_n28), .B(
        npu_inst_pe_1_1_1_n23), .S(npu_inst_pe_1_1_1_n8), .Z(
        npu_inst_pe_1_1_1_N94) );
  MUX2_X1 npu_inst_pe_1_1_1_U156 ( .A(npu_inst_pe_1_1_1_n25), .B(
        npu_inst_pe_1_1_1_n24), .S(npu_inst_pe_1_1_1_n6), .Z(
        npu_inst_pe_1_1_1_n28) );
  MUX2_X1 npu_inst_pe_1_1_1_U155 ( .A(npu_inst_pe_1_1_1_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_1_1_int_q_reg_v_1__1_), .S(npu_inst_pe_1_1_1_n4), .Z(
        npu_inst_pe_1_1_1_n25) );
  MUX2_X1 npu_inst_pe_1_1_1_U154 ( .A(npu_inst_pe_1_1_1_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_1_1_int_q_reg_v_3__1_), .S(npu_inst_pe_1_1_1_n4), .Z(
        npu_inst_pe_1_1_1_n24) );
  MUX2_X1 npu_inst_pe_1_1_1_U153 ( .A(npu_inst_pe_1_1_1_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_1_1_int_q_reg_v_5__1_), .S(npu_inst_pe_1_1_1_n4), .Z(
        npu_inst_pe_1_1_1_n23) );
  MUX2_X1 npu_inst_pe_1_1_1_U152 ( .A(npu_inst_pe_1_1_1_n22), .B(
        npu_inst_pe_1_1_1_n19), .S(npu_inst_pe_1_1_1_n8), .Z(
        npu_inst_int_data_x_1__1__1_) );
  MUX2_X1 npu_inst_pe_1_1_1_U151 ( .A(npu_inst_pe_1_1_1_n21), .B(
        npu_inst_pe_1_1_1_n20), .S(npu_inst_pe_1_1_1_n6), .Z(
        npu_inst_pe_1_1_1_n22) );
  MUX2_X1 npu_inst_pe_1_1_1_U150 ( .A(npu_inst_pe_1_1_1_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_1_1_int_q_reg_h_1__1_), .S(npu_inst_pe_1_1_1_n4), .Z(
        npu_inst_pe_1_1_1_n21) );
  MUX2_X1 npu_inst_pe_1_1_1_U149 ( .A(npu_inst_pe_1_1_1_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_1_1_int_q_reg_h_3__1_), .S(npu_inst_pe_1_1_1_n4), .Z(
        npu_inst_pe_1_1_1_n20) );
  MUX2_X1 npu_inst_pe_1_1_1_U148 ( .A(npu_inst_pe_1_1_1_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_1_1_int_q_reg_h_5__1_), .S(npu_inst_pe_1_1_1_n4), .Z(
        npu_inst_pe_1_1_1_n19) );
  MUX2_X1 npu_inst_pe_1_1_1_U147 ( .A(npu_inst_pe_1_1_1_n18), .B(
        npu_inst_pe_1_1_1_n15), .S(npu_inst_pe_1_1_1_n8), .Z(
        npu_inst_int_data_x_1__1__0_) );
  MUX2_X1 npu_inst_pe_1_1_1_U146 ( .A(npu_inst_pe_1_1_1_n17), .B(
        npu_inst_pe_1_1_1_n16), .S(npu_inst_pe_1_1_1_n6), .Z(
        npu_inst_pe_1_1_1_n18) );
  MUX2_X1 npu_inst_pe_1_1_1_U145 ( .A(npu_inst_pe_1_1_1_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_1_1_int_q_reg_h_1__0_), .S(npu_inst_pe_1_1_1_n4), .Z(
        npu_inst_pe_1_1_1_n17) );
  MUX2_X1 npu_inst_pe_1_1_1_U144 ( .A(npu_inst_pe_1_1_1_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_1_1_int_q_reg_h_3__0_), .S(npu_inst_pe_1_1_1_n4), .Z(
        npu_inst_pe_1_1_1_n16) );
  MUX2_X1 npu_inst_pe_1_1_1_U143 ( .A(npu_inst_pe_1_1_1_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_1_1_int_q_reg_h_5__0_), .S(npu_inst_pe_1_1_1_n4), .Z(
        npu_inst_pe_1_1_1_n15) );
  XOR2_X1 npu_inst_pe_1_1_1_U142 ( .A(npu_inst_pe_1_1_1_int_data_0_), .B(
        npu_inst_pe_1_1_1_int_q_acc_0_), .Z(npu_inst_pe_1_1_1_N73) );
  AND2_X1 npu_inst_pe_1_1_1_U141 ( .A1(npu_inst_pe_1_1_1_int_q_acc_0_), .A2(
        npu_inst_pe_1_1_1_int_data_0_), .ZN(npu_inst_pe_1_1_1_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_1_1_U140 ( .A(npu_inst_pe_1_1_1_int_q_acc_0_), .B(
        npu_inst_pe_1_1_1_n13), .ZN(npu_inst_pe_1_1_1_N65) );
  OR2_X1 npu_inst_pe_1_1_1_U139 ( .A1(npu_inst_pe_1_1_1_n13), .A2(
        npu_inst_pe_1_1_1_int_q_acc_0_), .ZN(npu_inst_pe_1_1_1_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_1_1_U138 ( .A(npu_inst_pe_1_1_1_int_q_acc_2_), .B(
        npu_inst_pe_1_1_1_add_79_carry_2_), .Z(npu_inst_pe_1_1_1_N75) );
  AND2_X1 npu_inst_pe_1_1_1_U137 ( .A1(npu_inst_pe_1_1_1_add_79_carry_2_), 
        .A2(npu_inst_pe_1_1_1_int_q_acc_2_), .ZN(
        npu_inst_pe_1_1_1_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_1_1_U136 ( .A(npu_inst_pe_1_1_1_int_q_acc_3_), .B(
        npu_inst_pe_1_1_1_add_79_carry_3_), .Z(npu_inst_pe_1_1_1_N76) );
  AND2_X1 npu_inst_pe_1_1_1_U135 ( .A1(npu_inst_pe_1_1_1_add_79_carry_3_), 
        .A2(npu_inst_pe_1_1_1_int_q_acc_3_), .ZN(
        npu_inst_pe_1_1_1_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_1_1_U134 ( .A(npu_inst_pe_1_1_1_int_q_acc_4_), .B(
        npu_inst_pe_1_1_1_add_79_carry_4_), .Z(npu_inst_pe_1_1_1_N77) );
  AND2_X1 npu_inst_pe_1_1_1_U133 ( .A1(npu_inst_pe_1_1_1_add_79_carry_4_), 
        .A2(npu_inst_pe_1_1_1_int_q_acc_4_), .ZN(
        npu_inst_pe_1_1_1_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_1_1_U132 ( .A(npu_inst_pe_1_1_1_int_q_acc_5_), .B(
        npu_inst_pe_1_1_1_add_79_carry_5_), .Z(npu_inst_pe_1_1_1_N78) );
  AND2_X1 npu_inst_pe_1_1_1_U131 ( .A1(npu_inst_pe_1_1_1_add_79_carry_5_), 
        .A2(npu_inst_pe_1_1_1_int_q_acc_5_), .ZN(
        npu_inst_pe_1_1_1_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_1_1_U130 ( .A(npu_inst_pe_1_1_1_int_q_acc_6_), .B(
        npu_inst_pe_1_1_1_add_79_carry_6_), .Z(npu_inst_pe_1_1_1_N79) );
  AND2_X1 npu_inst_pe_1_1_1_U129 ( .A1(npu_inst_pe_1_1_1_add_79_carry_6_), 
        .A2(npu_inst_pe_1_1_1_int_q_acc_6_), .ZN(
        npu_inst_pe_1_1_1_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_1_1_U128 ( .A(npu_inst_pe_1_1_1_int_q_acc_7_), .B(
        npu_inst_pe_1_1_1_add_79_carry_7_), .Z(npu_inst_pe_1_1_1_N80) );
  XNOR2_X1 npu_inst_pe_1_1_1_U127 ( .A(npu_inst_pe_1_1_1_sub_77_carry_2_), .B(
        npu_inst_pe_1_1_1_int_q_acc_2_), .ZN(npu_inst_pe_1_1_1_N67) );
  OR2_X1 npu_inst_pe_1_1_1_U126 ( .A1(npu_inst_pe_1_1_1_int_q_acc_2_), .A2(
        npu_inst_pe_1_1_1_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_1_1_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_1_1_U125 ( .A(npu_inst_pe_1_1_1_sub_77_carry_3_), .B(
        npu_inst_pe_1_1_1_int_q_acc_3_), .ZN(npu_inst_pe_1_1_1_N68) );
  OR2_X1 npu_inst_pe_1_1_1_U124 ( .A1(npu_inst_pe_1_1_1_int_q_acc_3_), .A2(
        npu_inst_pe_1_1_1_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_1_1_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_1_1_U123 ( .A(npu_inst_pe_1_1_1_sub_77_carry_4_), .B(
        npu_inst_pe_1_1_1_int_q_acc_4_), .ZN(npu_inst_pe_1_1_1_N69) );
  OR2_X1 npu_inst_pe_1_1_1_U122 ( .A1(npu_inst_pe_1_1_1_int_q_acc_4_), .A2(
        npu_inst_pe_1_1_1_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_1_1_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_1_1_U121 ( .A(npu_inst_pe_1_1_1_sub_77_carry_5_), .B(
        npu_inst_pe_1_1_1_int_q_acc_5_), .ZN(npu_inst_pe_1_1_1_N70) );
  OR2_X1 npu_inst_pe_1_1_1_U120 ( .A1(npu_inst_pe_1_1_1_int_q_acc_5_), .A2(
        npu_inst_pe_1_1_1_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_1_1_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_1_1_U119 ( .A(npu_inst_pe_1_1_1_sub_77_carry_6_), .B(
        npu_inst_pe_1_1_1_int_q_acc_6_), .ZN(npu_inst_pe_1_1_1_N71) );
  OR2_X1 npu_inst_pe_1_1_1_U118 ( .A1(npu_inst_pe_1_1_1_int_q_acc_6_), .A2(
        npu_inst_pe_1_1_1_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_1_1_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_1_1_U117 ( .A(npu_inst_pe_1_1_1_int_q_acc_7_), .B(
        npu_inst_pe_1_1_1_sub_77_carry_7_), .ZN(npu_inst_pe_1_1_1_N72) );
  INV_X1 npu_inst_pe_1_1_1_U116 ( .A(npu_inst_n79), .ZN(npu_inst_pe_1_1_1_n7)
         );
  INV_X1 npu_inst_pe_1_1_1_U115 ( .A(npu_inst_pe_1_1_1_n7), .ZN(
        npu_inst_pe_1_1_1_n6) );
  INV_X1 npu_inst_pe_1_1_1_U114 ( .A(npu_inst_n59), .ZN(npu_inst_pe_1_1_1_n3)
         );
  AOI22_X1 npu_inst_pe_1_1_1_U113 ( .A1(npu_inst_int_data_y_2__1__0_), .A2(
        npu_inst_pe_1_1_1_n58), .B1(npu_inst_pe_1_1_1_n114), .B2(
        npu_inst_pe_1_1_1_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_1_1_n57) );
  INV_X1 npu_inst_pe_1_1_1_U112 ( .A(npu_inst_pe_1_1_1_n57), .ZN(
        npu_inst_pe_1_1_1_n108) );
  AOI22_X1 npu_inst_pe_1_1_1_U111 ( .A1(npu_inst_int_data_y_2__1__0_), .A2(
        npu_inst_pe_1_1_1_n54), .B1(npu_inst_pe_1_1_1_n115), .B2(
        npu_inst_pe_1_1_1_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_1_1_n53) );
  INV_X1 npu_inst_pe_1_1_1_U110 ( .A(npu_inst_pe_1_1_1_n53), .ZN(
        npu_inst_pe_1_1_1_n109) );
  AOI22_X1 npu_inst_pe_1_1_1_U107 ( .A1(npu_inst_int_data_y_2__1__0_), .A2(
        npu_inst_pe_1_1_1_n50), .B1(npu_inst_pe_1_1_1_n116), .B2(
        npu_inst_pe_1_1_1_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_1_1_n49) );
  INV_X1 npu_inst_pe_1_1_1_U106 ( .A(npu_inst_pe_1_1_1_n49), .ZN(
        npu_inst_pe_1_1_1_n110) );
  AOI22_X1 npu_inst_pe_1_1_1_U105 ( .A1(npu_inst_int_data_y_2__1__0_), .A2(
        npu_inst_pe_1_1_1_n46), .B1(npu_inst_pe_1_1_1_n117), .B2(
        npu_inst_pe_1_1_1_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_1_1_n45) );
  INV_X1 npu_inst_pe_1_1_1_U104 ( .A(npu_inst_pe_1_1_1_n45), .ZN(
        npu_inst_pe_1_1_1_n111) );
  AOI22_X1 npu_inst_pe_1_1_1_U103 ( .A1(npu_inst_int_data_y_2__1__0_), .A2(
        npu_inst_pe_1_1_1_n42), .B1(npu_inst_pe_1_1_1_n119), .B2(
        npu_inst_pe_1_1_1_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_1_1_n41) );
  INV_X1 npu_inst_pe_1_1_1_U102 ( .A(npu_inst_pe_1_1_1_n41), .ZN(
        npu_inst_pe_1_1_1_n112) );
  AOI22_X1 npu_inst_pe_1_1_1_U101 ( .A1(npu_inst_int_data_y_2__1__1_), .A2(
        npu_inst_pe_1_1_1_n58), .B1(npu_inst_pe_1_1_1_n114), .B2(
        npu_inst_pe_1_1_1_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_1_1_n59) );
  INV_X1 npu_inst_pe_1_1_1_U100 ( .A(npu_inst_pe_1_1_1_n59), .ZN(
        npu_inst_pe_1_1_1_n102) );
  AOI22_X1 npu_inst_pe_1_1_1_U99 ( .A1(npu_inst_int_data_y_2__1__1_), .A2(
        npu_inst_pe_1_1_1_n54), .B1(npu_inst_pe_1_1_1_n115), .B2(
        npu_inst_pe_1_1_1_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_1_1_n55) );
  INV_X1 npu_inst_pe_1_1_1_U98 ( .A(npu_inst_pe_1_1_1_n55), .ZN(
        npu_inst_pe_1_1_1_n103) );
  AOI22_X1 npu_inst_pe_1_1_1_U97 ( .A1(npu_inst_int_data_y_2__1__1_), .A2(
        npu_inst_pe_1_1_1_n50), .B1(npu_inst_pe_1_1_1_n116), .B2(
        npu_inst_pe_1_1_1_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_1_1_n51) );
  INV_X1 npu_inst_pe_1_1_1_U96 ( .A(npu_inst_pe_1_1_1_n51), .ZN(
        npu_inst_pe_1_1_1_n104) );
  AOI22_X1 npu_inst_pe_1_1_1_U95 ( .A1(npu_inst_int_data_y_2__1__1_), .A2(
        npu_inst_pe_1_1_1_n46), .B1(npu_inst_pe_1_1_1_n117), .B2(
        npu_inst_pe_1_1_1_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_1_1_n47) );
  INV_X1 npu_inst_pe_1_1_1_U94 ( .A(npu_inst_pe_1_1_1_n47), .ZN(
        npu_inst_pe_1_1_1_n105) );
  AOI22_X1 npu_inst_pe_1_1_1_U93 ( .A1(npu_inst_int_data_y_2__1__1_), .A2(
        npu_inst_pe_1_1_1_n42), .B1(npu_inst_pe_1_1_1_n119), .B2(
        npu_inst_pe_1_1_1_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_1_1_n43) );
  INV_X1 npu_inst_pe_1_1_1_U92 ( .A(npu_inst_pe_1_1_1_n43), .ZN(
        npu_inst_pe_1_1_1_n106) );
  AOI22_X1 npu_inst_pe_1_1_1_U91 ( .A1(npu_inst_pe_1_1_1_n38), .A2(
        npu_inst_int_data_y_2__1__1_), .B1(npu_inst_pe_1_1_1_n118), .B2(
        npu_inst_pe_1_1_1_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_1_1_n39) );
  INV_X1 npu_inst_pe_1_1_1_U90 ( .A(npu_inst_pe_1_1_1_n39), .ZN(
        npu_inst_pe_1_1_1_n107) );
  AOI22_X1 npu_inst_pe_1_1_1_U89 ( .A1(npu_inst_pe_1_1_1_n38), .A2(
        npu_inst_int_data_y_2__1__0_), .B1(npu_inst_pe_1_1_1_n118), .B2(
        npu_inst_pe_1_1_1_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_1_1_n37) );
  INV_X1 npu_inst_pe_1_1_1_U88 ( .A(npu_inst_pe_1_1_1_n37), .ZN(
        npu_inst_pe_1_1_1_n113) );
  NAND2_X1 npu_inst_pe_1_1_1_U87 ( .A1(npu_inst_pe_1_1_1_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_1_1_n60), .ZN(npu_inst_pe_1_1_1_n74) );
  OAI21_X1 npu_inst_pe_1_1_1_U86 ( .B1(npu_inst_pe_1_1_1_n63), .B2(
        npu_inst_pe_1_1_1_n60), .A(npu_inst_pe_1_1_1_n74), .ZN(
        npu_inst_pe_1_1_1_n97) );
  NAND2_X1 npu_inst_pe_1_1_1_U85 ( .A1(npu_inst_pe_1_1_1_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_1_1_n60), .ZN(npu_inst_pe_1_1_1_n73) );
  OAI21_X1 npu_inst_pe_1_1_1_U84 ( .B1(npu_inst_pe_1_1_1_n61), .B2(
        npu_inst_pe_1_1_1_n60), .A(npu_inst_pe_1_1_1_n73), .ZN(
        npu_inst_pe_1_1_1_n96) );
  NAND2_X1 npu_inst_pe_1_1_1_U83 ( .A1(npu_inst_pe_1_1_1_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_1_1_n56), .ZN(npu_inst_pe_1_1_1_n72) );
  OAI21_X1 npu_inst_pe_1_1_1_U82 ( .B1(npu_inst_pe_1_1_1_n63), .B2(
        npu_inst_pe_1_1_1_n56), .A(npu_inst_pe_1_1_1_n72), .ZN(
        npu_inst_pe_1_1_1_n95) );
  NAND2_X1 npu_inst_pe_1_1_1_U81 ( .A1(npu_inst_pe_1_1_1_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_1_1_n56), .ZN(npu_inst_pe_1_1_1_n71) );
  OAI21_X1 npu_inst_pe_1_1_1_U80 ( .B1(npu_inst_pe_1_1_1_n61), .B2(
        npu_inst_pe_1_1_1_n56), .A(npu_inst_pe_1_1_1_n71), .ZN(
        npu_inst_pe_1_1_1_n94) );
  NAND2_X1 npu_inst_pe_1_1_1_U79 ( .A1(npu_inst_pe_1_1_1_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_1_1_n52), .ZN(npu_inst_pe_1_1_1_n70) );
  OAI21_X1 npu_inst_pe_1_1_1_U78 ( .B1(npu_inst_pe_1_1_1_n63), .B2(
        npu_inst_pe_1_1_1_n52), .A(npu_inst_pe_1_1_1_n70), .ZN(
        npu_inst_pe_1_1_1_n93) );
  NAND2_X1 npu_inst_pe_1_1_1_U77 ( .A1(npu_inst_pe_1_1_1_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_1_1_n52), .ZN(npu_inst_pe_1_1_1_n69) );
  OAI21_X1 npu_inst_pe_1_1_1_U76 ( .B1(npu_inst_pe_1_1_1_n61), .B2(
        npu_inst_pe_1_1_1_n52), .A(npu_inst_pe_1_1_1_n69), .ZN(
        npu_inst_pe_1_1_1_n92) );
  NAND2_X1 npu_inst_pe_1_1_1_U75 ( .A1(npu_inst_pe_1_1_1_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_1_1_n48), .ZN(npu_inst_pe_1_1_1_n68) );
  OAI21_X1 npu_inst_pe_1_1_1_U74 ( .B1(npu_inst_pe_1_1_1_n63), .B2(
        npu_inst_pe_1_1_1_n48), .A(npu_inst_pe_1_1_1_n68), .ZN(
        npu_inst_pe_1_1_1_n91) );
  NAND2_X1 npu_inst_pe_1_1_1_U73 ( .A1(npu_inst_pe_1_1_1_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_1_1_n48), .ZN(npu_inst_pe_1_1_1_n67) );
  OAI21_X1 npu_inst_pe_1_1_1_U72 ( .B1(npu_inst_pe_1_1_1_n61), .B2(
        npu_inst_pe_1_1_1_n48), .A(npu_inst_pe_1_1_1_n67), .ZN(
        npu_inst_pe_1_1_1_n90) );
  NAND2_X1 npu_inst_pe_1_1_1_U71 ( .A1(npu_inst_pe_1_1_1_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_1_1_n44), .ZN(npu_inst_pe_1_1_1_n66) );
  OAI21_X1 npu_inst_pe_1_1_1_U70 ( .B1(npu_inst_pe_1_1_1_n63), .B2(
        npu_inst_pe_1_1_1_n44), .A(npu_inst_pe_1_1_1_n66), .ZN(
        npu_inst_pe_1_1_1_n89) );
  NAND2_X1 npu_inst_pe_1_1_1_U69 ( .A1(npu_inst_pe_1_1_1_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_1_1_n44), .ZN(npu_inst_pe_1_1_1_n65) );
  OAI21_X1 npu_inst_pe_1_1_1_U68 ( .B1(npu_inst_pe_1_1_1_n61), .B2(
        npu_inst_pe_1_1_1_n44), .A(npu_inst_pe_1_1_1_n65), .ZN(
        npu_inst_pe_1_1_1_n88) );
  NAND2_X1 npu_inst_pe_1_1_1_U67 ( .A1(npu_inst_pe_1_1_1_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_1_1_n40), .ZN(npu_inst_pe_1_1_1_n64) );
  OAI21_X1 npu_inst_pe_1_1_1_U66 ( .B1(npu_inst_pe_1_1_1_n63), .B2(
        npu_inst_pe_1_1_1_n40), .A(npu_inst_pe_1_1_1_n64), .ZN(
        npu_inst_pe_1_1_1_n87) );
  NAND2_X1 npu_inst_pe_1_1_1_U65 ( .A1(npu_inst_pe_1_1_1_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_1_1_n40), .ZN(npu_inst_pe_1_1_1_n62) );
  OAI21_X1 npu_inst_pe_1_1_1_U64 ( .B1(npu_inst_pe_1_1_1_n61), .B2(
        npu_inst_pe_1_1_1_n40), .A(npu_inst_pe_1_1_1_n62), .ZN(
        npu_inst_pe_1_1_1_n86) );
  AND2_X1 npu_inst_pe_1_1_1_U63 ( .A1(npu_inst_pe_1_1_1_N93), .A2(npu_inst_n59), .ZN(npu_inst_int_data_y_1__1__0_) );
  AND2_X1 npu_inst_pe_1_1_1_U62 ( .A1(npu_inst_n59), .A2(npu_inst_pe_1_1_1_N94), .ZN(npu_inst_int_data_y_1__1__1_) );
  NOR3_X1 npu_inst_pe_1_1_1_U61 ( .A1(npu_inst_pe_1_1_1_n26), .A2(npu_inst_n59), .A3(npu_inst_int_ckg[54]), .ZN(npu_inst_pe_1_1_1_n85) );
  OR2_X1 npu_inst_pe_1_1_1_U60 ( .A1(npu_inst_pe_1_1_1_n85), .A2(
        npu_inst_pe_1_1_1_n2), .ZN(npu_inst_pe_1_1_1_N84) );
  AND2_X1 npu_inst_pe_1_1_1_U59 ( .A1(npu_inst_pe_1_1_1_int_q_acc_0_), .A2(
        npu_inst_pe_1_1_1_n1), .ZN(npu_inst_int_data_res_1__1__0_) );
  AND2_X1 npu_inst_pe_1_1_1_U58 ( .A1(npu_inst_pe_1_1_1_n2), .A2(
        npu_inst_pe_1_1_1_int_q_acc_7_), .ZN(npu_inst_int_data_res_1__1__7_)
         );
  AND2_X1 npu_inst_pe_1_1_1_U57 ( .A1(npu_inst_pe_1_1_1_int_q_acc_1_), .A2(
        npu_inst_pe_1_1_1_n1), .ZN(npu_inst_int_data_res_1__1__1_) );
  AND2_X1 npu_inst_pe_1_1_1_U56 ( .A1(npu_inst_pe_1_1_1_int_q_acc_2_), .A2(
        npu_inst_pe_1_1_1_n1), .ZN(npu_inst_int_data_res_1__1__2_) );
  AND2_X1 npu_inst_pe_1_1_1_U55 ( .A1(npu_inst_pe_1_1_1_int_q_acc_3_), .A2(
        npu_inst_pe_1_1_1_n2), .ZN(npu_inst_int_data_res_1__1__3_) );
  AND2_X1 npu_inst_pe_1_1_1_U54 ( .A1(npu_inst_pe_1_1_1_int_q_acc_4_), .A2(
        npu_inst_pe_1_1_1_n2), .ZN(npu_inst_int_data_res_1__1__4_) );
  AND2_X1 npu_inst_pe_1_1_1_U53 ( .A1(npu_inst_pe_1_1_1_int_q_acc_5_), .A2(
        npu_inst_pe_1_1_1_n2), .ZN(npu_inst_int_data_res_1__1__5_) );
  AND2_X1 npu_inst_pe_1_1_1_U52 ( .A1(npu_inst_pe_1_1_1_int_q_acc_6_), .A2(
        npu_inst_pe_1_1_1_n2), .ZN(npu_inst_int_data_res_1__1__6_) );
  AOI222_X1 npu_inst_pe_1_1_1_U51 ( .A1(npu_inst_int_data_res_2__1__0_), .A2(
        npu_inst_pe_1_1_1_n1), .B1(npu_inst_pe_1_1_1_N73), .B2(
        npu_inst_pe_1_1_1_n76), .C1(npu_inst_pe_1_1_1_N65), .C2(
        npu_inst_pe_1_1_1_n77), .ZN(npu_inst_pe_1_1_1_n84) );
  INV_X1 npu_inst_pe_1_1_1_U50 ( .A(npu_inst_pe_1_1_1_n84), .ZN(
        npu_inst_pe_1_1_1_n101) );
  AOI222_X1 npu_inst_pe_1_1_1_U49 ( .A1(npu_inst_int_data_res_2__1__7_), .A2(
        npu_inst_pe_1_1_1_n1), .B1(npu_inst_pe_1_1_1_N80), .B2(
        npu_inst_pe_1_1_1_n76), .C1(npu_inst_pe_1_1_1_N72), .C2(
        npu_inst_pe_1_1_1_n77), .ZN(npu_inst_pe_1_1_1_n75) );
  INV_X1 npu_inst_pe_1_1_1_U48 ( .A(npu_inst_pe_1_1_1_n75), .ZN(
        npu_inst_pe_1_1_1_n33) );
  AOI222_X1 npu_inst_pe_1_1_1_U47 ( .A1(npu_inst_int_data_res_2__1__1_), .A2(
        npu_inst_pe_1_1_1_n1), .B1(npu_inst_pe_1_1_1_N74), .B2(
        npu_inst_pe_1_1_1_n76), .C1(npu_inst_pe_1_1_1_N66), .C2(
        npu_inst_pe_1_1_1_n77), .ZN(npu_inst_pe_1_1_1_n83) );
  INV_X1 npu_inst_pe_1_1_1_U46 ( .A(npu_inst_pe_1_1_1_n83), .ZN(
        npu_inst_pe_1_1_1_n100) );
  AOI222_X1 npu_inst_pe_1_1_1_U45 ( .A1(npu_inst_int_data_res_2__1__2_), .A2(
        npu_inst_pe_1_1_1_n1), .B1(npu_inst_pe_1_1_1_N75), .B2(
        npu_inst_pe_1_1_1_n76), .C1(npu_inst_pe_1_1_1_N67), .C2(
        npu_inst_pe_1_1_1_n77), .ZN(npu_inst_pe_1_1_1_n82) );
  INV_X1 npu_inst_pe_1_1_1_U44 ( .A(npu_inst_pe_1_1_1_n82), .ZN(
        npu_inst_pe_1_1_1_n99) );
  AOI222_X1 npu_inst_pe_1_1_1_U43 ( .A1(npu_inst_int_data_res_2__1__3_), .A2(
        npu_inst_pe_1_1_1_n1), .B1(npu_inst_pe_1_1_1_N76), .B2(
        npu_inst_pe_1_1_1_n76), .C1(npu_inst_pe_1_1_1_N68), .C2(
        npu_inst_pe_1_1_1_n77), .ZN(npu_inst_pe_1_1_1_n81) );
  INV_X1 npu_inst_pe_1_1_1_U42 ( .A(npu_inst_pe_1_1_1_n81), .ZN(
        npu_inst_pe_1_1_1_n98) );
  AOI222_X1 npu_inst_pe_1_1_1_U41 ( .A1(npu_inst_int_data_res_2__1__4_), .A2(
        npu_inst_pe_1_1_1_n1), .B1(npu_inst_pe_1_1_1_N77), .B2(
        npu_inst_pe_1_1_1_n76), .C1(npu_inst_pe_1_1_1_N69), .C2(
        npu_inst_pe_1_1_1_n77), .ZN(npu_inst_pe_1_1_1_n80) );
  INV_X1 npu_inst_pe_1_1_1_U40 ( .A(npu_inst_pe_1_1_1_n80), .ZN(
        npu_inst_pe_1_1_1_n36) );
  AOI222_X1 npu_inst_pe_1_1_1_U39 ( .A1(npu_inst_int_data_res_2__1__5_), .A2(
        npu_inst_pe_1_1_1_n1), .B1(npu_inst_pe_1_1_1_N78), .B2(
        npu_inst_pe_1_1_1_n76), .C1(npu_inst_pe_1_1_1_N70), .C2(
        npu_inst_pe_1_1_1_n77), .ZN(npu_inst_pe_1_1_1_n79) );
  INV_X1 npu_inst_pe_1_1_1_U38 ( .A(npu_inst_pe_1_1_1_n79), .ZN(
        npu_inst_pe_1_1_1_n35) );
  AOI222_X1 npu_inst_pe_1_1_1_U37 ( .A1(npu_inst_int_data_res_2__1__6_), .A2(
        npu_inst_pe_1_1_1_n1), .B1(npu_inst_pe_1_1_1_N79), .B2(
        npu_inst_pe_1_1_1_n76), .C1(npu_inst_pe_1_1_1_N71), .C2(
        npu_inst_pe_1_1_1_n77), .ZN(npu_inst_pe_1_1_1_n78) );
  INV_X1 npu_inst_pe_1_1_1_U36 ( .A(npu_inst_pe_1_1_1_n78), .ZN(
        npu_inst_pe_1_1_1_n34) );
  INV_X1 npu_inst_pe_1_1_1_U35 ( .A(npu_inst_pe_1_1_1_int_data_1_), .ZN(
        npu_inst_pe_1_1_1_n14) );
  AND2_X1 npu_inst_pe_1_1_1_U34 ( .A1(npu_inst_int_data_x_1__1__1_), .A2(
        npu_inst_pe_1_1_1_int_q_weight_1_), .ZN(npu_inst_pe_1_1_1_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_1_1_U33 ( .A1(npu_inst_int_data_x_1__1__0_), .A2(
        npu_inst_pe_1_1_1_int_q_weight_1_), .ZN(npu_inst_pe_1_1_1_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_1_1_U32 ( .A1(npu_inst_n59), .A2(
        npu_inst_int_data_y_2__1__1_), .B1(npu_inst_pe_1_1_1_n3), .B2(
        npu_inst_int_data_x_1__2__1_), .ZN(npu_inst_pe_1_1_1_n63) );
  AOI22_X1 npu_inst_pe_1_1_1_U31 ( .A1(npu_inst_n59), .A2(
        npu_inst_int_data_y_2__1__0_), .B1(npu_inst_pe_1_1_1_n3), .B2(
        npu_inst_int_data_x_1__2__0_), .ZN(npu_inst_pe_1_1_1_n61) );
  INV_X1 npu_inst_pe_1_1_1_U30 ( .A(npu_inst_pe_1_1_1_int_data_0_), .ZN(
        npu_inst_pe_1_1_1_n13) );
  INV_X1 npu_inst_pe_1_1_1_U29 ( .A(npu_inst_n71), .ZN(npu_inst_pe_1_1_1_n5)
         );
  OR3_X1 npu_inst_pe_1_1_1_U28 ( .A1(npu_inst_pe_1_1_1_n6), .A2(
        npu_inst_pe_1_1_1_n8), .A3(npu_inst_pe_1_1_1_n5), .ZN(
        npu_inst_pe_1_1_1_n56) );
  OR3_X1 npu_inst_pe_1_1_1_U27 ( .A1(npu_inst_pe_1_1_1_n5), .A2(
        npu_inst_pe_1_1_1_n8), .A3(npu_inst_pe_1_1_1_n7), .ZN(
        npu_inst_pe_1_1_1_n48) );
  INV_X1 npu_inst_pe_1_1_1_U26 ( .A(npu_inst_pe_1_1_1_n5), .ZN(
        npu_inst_pe_1_1_1_n4) );
  INV_X1 npu_inst_pe_1_1_1_U25 ( .A(npu_inst_n126), .ZN(npu_inst_pe_1_1_1_n12)
         );
  OR3_X1 npu_inst_pe_1_1_1_U24 ( .A1(npu_inst_pe_1_1_1_n4), .A2(
        npu_inst_pe_1_1_1_n8), .A3(npu_inst_pe_1_1_1_n7), .ZN(
        npu_inst_pe_1_1_1_n52) );
  OR3_X1 npu_inst_pe_1_1_1_U23 ( .A1(npu_inst_pe_1_1_1_n6), .A2(
        npu_inst_pe_1_1_1_n8), .A3(npu_inst_pe_1_1_1_n4), .ZN(
        npu_inst_pe_1_1_1_n60) );
  NOR2_X1 npu_inst_pe_1_1_1_U22 ( .A1(npu_inst_pe_1_1_1_n60), .A2(
        npu_inst_pe_1_1_1_n3), .ZN(npu_inst_pe_1_1_1_n58) );
  NOR2_X1 npu_inst_pe_1_1_1_U21 ( .A1(npu_inst_pe_1_1_1_n56), .A2(
        npu_inst_pe_1_1_1_n3), .ZN(npu_inst_pe_1_1_1_n54) );
  NOR2_X1 npu_inst_pe_1_1_1_U20 ( .A1(npu_inst_pe_1_1_1_n52), .A2(
        npu_inst_pe_1_1_1_n3), .ZN(npu_inst_pe_1_1_1_n50) );
  NOR2_X1 npu_inst_pe_1_1_1_U19 ( .A1(npu_inst_pe_1_1_1_n48), .A2(
        npu_inst_pe_1_1_1_n3), .ZN(npu_inst_pe_1_1_1_n46) );
  NOR2_X1 npu_inst_pe_1_1_1_U18 ( .A1(npu_inst_pe_1_1_1_n40), .A2(
        npu_inst_pe_1_1_1_n3), .ZN(npu_inst_pe_1_1_1_n38) );
  NOR2_X1 npu_inst_pe_1_1_1_U17 ( .A1(npu_inst_pe_1_1_1_n44), .A2(
        npu_inst_pe_1_1_1_n3), .ZN(npu_inst_pe_1_1_1_n42) );
  BUF_X1 npu_inst_pe_1_1_1_U16 ( .A(npu_inst_n105), .Z(npu_inst_pe_1_1_1_n8)
         );
  BUF_X1 npu_inst_pe_1_1_1_U15 ( .A(npu_inst_pe_1_1_1_n12), .Z(
        npu_inst_pe_1_1_1_n11) );
  BUF_X1 npu_inst_pe_1_1_1_U14 ( .A(npu_inst_pe_1_1_1_n12), .Z(
        npu_inst_pe_1_1_1_n10) );
  BUF_X1 npu_inst_pe_1_1_1_U13 ( .A(npu_inst_pe_1_1_1_n12), .Z(
        npu_inst_pe_1_1_1_n9) );
  INV_X1 npu_inst_pe_1_1_1_U12 ( .A(npu_inst_pe_1_1_1_n38), .ZN(
        npu_inst_pe_1_1_1_n118) );
  INV_X1 npu_inst_pe_1_1_1_U11 ( .A(npu_inst_pe_1_1_1_n58), .ZN(
        npu_inst_pe_1_1_1_n114) );
  INV_X1 npu_inst_pe_1_1_1_U10 ( .A(npu_inst_pe_1_1_1_n54), .ZN(
        npu_inst_pe_1_1_1_n115) );
  INV_X1 npu_inst_pe_1_1_1_U9 ( .A(npu_inst_pe_1_1_1_n50), .ZN(
        npu_inst_pe_1_1_1_n116) );
  INV_X1 npu_inst_pe_1_1_1_U8 ( .A(npu_inst_pe_1_1_1_n46), .ZN(
        npu_inst_pe_1_1_1_n117) );
  INV_X1 npu_inst_pe_1_1_1_U7 ( .A(npu_inst_pe_1_1_1_n42), .ZN(
        npu_inst_pe_1_1_1_n119) );
  BUF_X1 npu_inst_pe_1_1_1_U6 ( .A(npu_inst_n34), .Z(npu_inst_pe_1_1_1_n2) );
  BUF_X1 npu_inst_pe_1_1_1_U5 ( .A(npu_inst_n34), .Z(npu_inst_pe_1_1_1_n1) );
  NOR2_X1 npu_inst_pe_1_1_1_U4 ( .A1(npu_inst_pe_1_1_1_int_q_weight_0_), .A2(
        npu_inst_pe_1_1_1_n1), .ZN(npu_inst_pe_1_1_1_n76) );
  NOR2_X1 npu_inst_pe_1_1_1_U3 ( .A1(npu_inst_pe_1_1_1_n27), .A2(
        npu_inst_pe_1_1_1_n1), .ZN(npu_inst_pe_1_1_1_n77) );
  FA_X1 npu_inst_pe_1_1_1_sub_77_U2_1 ( .A(npu_inst_pe_1_1_1_int_q_acc_1_), 
        .B(npu_inst_pe_1_1_1_n14), .CI(npu_inst_pe_1_1_1_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_1_1_sub_77_carry_2_), .S(npu_inst_pe_1_1_1_N66) );
  FA_X1 npu_inst_pe_1_1_1_add_79_U1_1 ( .A(npu_inst_pe_1_1_1_int_q_acc_1_), 
        .B(npu_inst_pe_1_1_1_int_data_1_), .CI(
        npu_inst_pe_1_1_1_add_79_carry_1_), .CO(
        npu_inst_pe_1_1_1_add_79_carry_2_), .S(npu_inst_pe_1_1_1_N74) );
  NAND3_X1 npu_inst_pe_1_1_1_U109 ( .A1(npu_inst_pe_1_1_1_n5), .A2(
        npu_inst_pe_1_1_1_n7), .A3(npu_inst_pe_1_1_1_n8), .ZN(
        npu_inst_pe_1_1_1_n44) );
  NAND3_X1 npu_inst_pe_1_1_1_U108 ( .A1(npu_inst_pe_1_1_1_n4), .A2(
        npu_inst_pe_1_1_1_n7), .A3(npu_inst_pe_1_1_1_n8), .ZN(
        npu_inst_pe_1_1_1_n40) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_1_1_n34), .CK(
        npu_inst_pe_1_1_1_net4086), .RN(npu_inst_pe_1_1_1_n9), .Q(
        npu_inst_pe_1_1_1_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_1_1_n35), .CK(
        npu_inst_pe_1_1_1_net4086), .RN(npu_inst_pe_1_1_1_n9), .Q(
        npu_inst_pe_1_1_1_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_1_1_n36), .CK(
        npu_inst_pe_1_1_1_net4086), .RN(npu_inst_pe_1_1_1_n9), .Q(
        npu_inst_pe_1_1_1_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_1_1_n98), .CK(
        npu_inst_pe_1_1_1_net4086), .RN(npu_inst_pe_1_1_1_n9), .Q(
        npu_inst_pe_1_1_1_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_1_1_n99), .CK(
        npu_inst_pe_1_1_1_net4086), .RN(npu_inst_pe_1_1_1_n9), .Q(
        npu_inst_pe_1_1_1_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_1_1_n100), 
        .CK(npu_inst_pe_1_1_1_net4086), .RN(npu_inst_pe_1_1_1_n9), .Q(
        npu_inst_pe_1_1_1_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_1_1_n33), .CK(
        npu_inst_pe_1_1_1_net4086), .RN(npu_inst_pe_1_1_1_n9), .Q(
        npu_inst_pe_1_1_1_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_1_1_n101), 
        .CK(npu_inst_pe_1_1_1_net4086), .RN(npu_inst_pe_1_1_1_n9), .Q(
        npu_inst_pe_1_1_1_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_weight_reg_0_ ( .D(npu_inst_n112), .CK(
        npu_inst_pe_1_1_1_net4092), .RN(npu_inst_pe_1_1_1_n9), .Q(
        npu_inst_pe_1_1_1_int_q_weight_0_), .QN(npu_inst_pe_1_1_1_n27) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_weight_reg_1_ ( .D(npu_inst_n118), .CK(
        npu_inst_pe_1_1_1_net4092), .RN(npu_inst_pe_1_1_1_n9), .Q(
        npu_inst_pe_1_1_1_int_q_weight_1_), .QN(npu_inst_pe_1_1_1_n26) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_1_1_n113), 
        .CK(npu_inst_pe_1_1_1_net4092), .RN(npu_inst_pe_1_1_1_n9), .Q(
        npu_inst_pe_1_1_1_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_1_1_n107), 
        .CK(npu_inst_pe_1_1_1_net4092), .RN(npu_inst_pe_1_1_1_n9), .Q(
        npu_inst_pe_1_1_1_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_1_1_n112), 
        .CK(npu_inst_pe_1_1_1_net4092), .RN(npu_inst_pe_1_1_1_n10), .Q(
        npu_inst_pe_1_1_1_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_1_1_n106), 
        .CK(npu_inst_pe_1_1_1_net4092), .RN(npu_inst_pe_1_1_1_n10), .Q(
        npu_inst_pe_1_1_1_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_1_1_n111), 
        .CK(npu_inst_pe_1_1_1_net4092), .RN(npu_inst_pe_1_1_1_n10), .Q(
        npu_inst_pe_1_1_1_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_1_1_n105), 
        .CK(npu_inst_pe_1_1_1_net4092), .RN(npu_inst_pe_1_1_1_n10), .Q(
        npu_inst_pe_1_1_1_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_1_1_n110), 
        .CK(npu_inst_pe_1_1_1_net4092), .RN(npu_inst_pe_1_1_1_n10), .Q(
        npu_inst_pe_1_1_1_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_1_1_n104), 
        .CK(npu_inst_pe_1_1_1_net4092), .RN(npu_inst_pe_1_1_1_n10), .Q(
        npu_inst_pe_1_1_1_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_1_1_n109), 
        .CK(npu_inst_pe_1_1_1_net4092), .RN(npu_inst_pe_1_1_1_n10), .Q(
        npu_inst_pe_1_1_1_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_1_1_n103), 
        .CK(npu_inst_pe_1_1_1_net4092), .RN(npu_inst_pe_1_1_1_n10), .Q(
        npu_inst_pe_1_1_1_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_1_1_n108), 
        .CK(npu_inst_pe_1_1_1_net4092), .RN(npu_inst_pe_1_1_1_n10), .Q(
        npu_inst_pe_1_1_1_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_1_1_n102), 
        .CK(npu_inst_pe_1_1_1_net4092), .RN(npu_inst_pe_1_1_1_n10), .Q(
        npu_inst_pe_1_1_1_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_1_1_n86), 
        .CK(npu_inst_pe_1_1_1_net4092), .RN(npu_inst_pe_1_1_1_n10), .Q(
        npu_inst_pe_1_1_1_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_1_1_n87), 
        .CK(npu_inst_pe_1_1_1_net4092), .RN(npu_inst_pe_1_1_1_n10), .Q(
        npu_inst_pe_1_1_1_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_1_1_n88), 
        .CK(npu_inst_pe_1_1_1_net4092), .RN(npu_inst_pe_1_1_1_n11), .Q(
        npu_inst_pe_1_1_1_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_1_1_n89), 
        .CK(npu_inst_pe_1_1_1_net4092), .RN(npu_inst_pe_1_1_1_n11), .Q(
        npu_inst_pe_1_1_1_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_1_1_n90), 
        .CK(npu_inst_pe_1_1_1_net4092), .RN(npu_inst_pe_1_1_1_n11), .Q(
        npu_inst_pe_1_1_1_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_1_1_n91), 
        .CK(npu_inst_pe_1_1_1_net4092), .RN(npu_inst_pe_1_1_1_n11), .Q(
        npu_inst_pe_1_1_1_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_1_1_n92), 
        .CK(npu_inst_pe_1_1_1_net4092), .RN(npu_inst_pe_1_1_1_n11), .Q(
        npu_inst_pe_1_1_1_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_1_1_n93), 
        .CK(npu_inst_pe_1_1_1_net4092), .RN(npu_inst_pe_1_1_1_n11), .Q(
        npu_inst_pe_1_1_1_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_1_1_n94), 
        .CK(npu_inst_pe_1_1_1_net4092), .RN(npu_inst_pe_1_1_1_n11), .Q(
        npu_inst_pe_1_1_1_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_1_1_n95), 
        .CK(npu_inst_pe_1_1_1_net4092), .RN(npu_inst_pe_1_1_1_n11), .Q(
        npu_inst_pe_1_1_1_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_1_1_n96), 
        .CK(npu_inst_pe_1_1_1_net4092), .RN(npu_inst_pe_1_1_1_n11), .Q(
        npu_inst_pe_1_1_1_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_1_1_n97), 
        .CK(npu_inst_pe_1_1_1_net4092), .RN(npu_inst_pe_1_1_1_n11), .Q(
        npu_inst_pe_1_1_1_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_1_1_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_1_1_N84), .SE(1'b0), .GCK(npu_inst_pe_1_1_1_net4086) );
  CLKGATETST_X1 npu_inst_pe_1_1_1_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n65), .SE(1'b0), .GCK(npu_inst_pe_1_1_1_net4092) );
  MUX2_X1 npu_inst_pe_1_1_2_U162 ( .A(npu_inst_pe_1_1_2_n32), .B(
        npu_inst_pe_1_1_2_n29), .S(npu_inst_pe_1_1_2_n8), .Z(
        npu_inst_pe_1_1_2_N93) );
  MUX2_X1 npu_inst_pe_1_1_2_U161 ( .A(npu_inst_pe_1_1_2_n31), .B(
        npu_inst_pe_1_1_2_n30), .S(npu_inst_pe_1_1_2_n6), .Z(
        npu_inst_pe_1_1_2_n32) );
  MUX2_X1 npu_inst_pe_1_1_2_U160 ( .A(npu_inst_pe_1_1_2_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_1_2_int_q_reg_v_1__0_), .S(npu_inst_pe_1_1_2_n4), .Z(
        npu_inst_pe_1_1_2_n31) );
  MUX2_X1 npu_inst_pe_1_1_2_U159 ( .A(npu_inst_pe_1_1_2_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_1_2_int_q_reg_v_3__0_), .S(npu_inst_pe_1_1_2_n4), .Z(
        npu_inst_pe_1_1_2_n30) );
  MUX2_X1 npu_inst_pe_1_1_2_U158 ( .A(npu_inst_pe_1_1_2_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_1_2_int_q_reg_v_5__0_), .S(npu_inst_pe_1_1_2_n4), .Z(
        npu_inst_pe_1_1_2_n29) );
  MUX2_X1 npu_inst_pe_1_1_2_U157 ( .A(npu_inst_pe_1_1_2_n28), .B(
        npu_inst_pe_1_1_2_n23), .S(npu_inst_pe_1_1_2_n8), .Z(
        npu_inst_pe_1_1_2_N94) );
  MUX2_X1 npu_inst_pe_1_1_2_U156 ( .A(npu_inst_pe_1_1_2_n25), .B(
        npu_inst_pe_1_1_2_n24), .S(npu_inst_pe_1_1_2_n6), .Z(
        npu_inst_pe_1_1_2_n28) );
  MUX2_X1 npu_inst_pe_1_1_2_U155 ( .A(npu_inst_pe_1_1_2_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_1_2_int_q_reg_v_1__1_), .S(npu_inst_pe_1_1_2_n4), .Z(
        npu_inst_pe_1_1_2_n25) );
  MUX2_X1 npu_inst_pe_1_1_2_U154 ( .A(npu_inst_pe_1_1_2_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_1_2_int_q_reg_v_3__1_), .S(npu_inst_pe_1_1_2_n4), .Z(
        npu_inst_pe_1_1_2_n24) );
  MUX2_X1 npu_inst_pe_1_1_2_U153 ( .A(npu_inst_pe_1_1_2_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_1_2_int_q_reg_v_5__1_), .S(npu_inst_pe_1_1_2_n4), .Z(
        npu_inst_pe_1_1_2_n23) );
  MUX2_X1 npu_inst_pe_1_1_2_U152 ( .A(npu_inst_pe_1_1_2_n22), .B(
        npu_inst_pe_1_1_2_n19), .S(npu_inst_pe_1_1_2_n8), .Z(
        npu_inst_int_data_x_1__2__1_) );
  MUX2_X1 npu_inst_pe_1_1_2_U151 ( .A(npu_inst_pe_1_1_2_n21), .B(
        npu_inst_pe_1_1_2_n20), .S(npu_inst_pe_1_1_2_n6), .Z(
        npu_inst_pe_1_1_2_n22) );
  MUX2_X1 npu_inst_pe_1_1_2_U150 ( .A(npu_inst_pe_1_1_2_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_1_2_int_q_reg_h_1__1_), .S(npu_inst_pe_1_1_2_n4), .Z(
        npu_inst_pe_1_1_2_n21) );
  MUX2_X1 npu_inst_pe_1_1_2_U149 ( .A(npu_inst_pe_1_1_2_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_1_2_int_q_reg_h_3__1_), .S(npu_inst_pe_1_1_2_n4), .Z(
        npu_inst_pe_1_1_2_n20) );
  MUX2_X1 npu_inst_pe_1_1_2_U148 ( .A(npu_inst_pe_1_1_2_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_1_2_int_q_reg_h_5__1_), .S(npu_inst_pe_1_1_2_n4), .Z(
        npu_inst_pe_1_1_2_n19) );
  MUX2_X1 npu_inst_pe_1_1_2_U147 ( .A(npu_inst_pe_1_1_2_n18), .B(
        npu_inst_pe_1_1_2_n15), .S(npu_inst_pe_1_1_2_n8), .Z(
        npu_inst_int_data_x_1__2__0_) );
  MUX2_X1 npu_inst_pe_1_1_2_U146 ( .A(npu_inst_pe_1_1_2_n17), .B(
        npu_inst_pe_1_1_2_n16), .S(npu_inst_pe_1_1_2_n6), .Z(
        npu_inst_pe_1_1_2_n18) );
  MUX2_X1 npu_inst_pe_1_1_2_U145 ( .A(npu_inst_pe_1_1_2_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_1_2_int_q_reg_h_1__0_), .S(npu_inst_pe_1_1_2_n4), .Z(
        npu_inst_pe_1_1_2_n17) );
  MUX2_X1 npu_inst_pe_1_1_2_U144 ( .A(npu_inst_pe_1_1_2_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_1_2_int_q_reg_h_3__0_), .S(npu_inst_pe_1_1_2_n4), .Z(
        npu_inst_pe_1_1_2_n16) );
  MUX2_X1 npu_inst_pe_1_1_2_U143 ( .A(npu_inst_pe_1_1_2_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_1_2_int_q_reg_h_5__0_), .S(npu_inst_pe_1_1_2_n4), .Z(
        npu_inst_pe_1_1_2_n15) );
  XOR2_X1 npu_inst_pe_1_1_2_U142 ( .A(npu_inst_pe_1_1_2_int_data_0_), .B(
        npu_inst_pe_1_1_2_int_q_acc_0_), .Z(npu_inst_pe_1_1_2_N73) );
  AND2_X1 npu_inst_pe_1_1_2_U141 ( .A1(npu_inst_pe_1_1_2_int_q_acc_0_), .A2(
        npu_inst_pe_1_1_2_int_data_0_), .ZN(npu_inst_pe_1_1_2_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_1_2_U140 ( .A(npu_inst_pe_1_1_2_int_q_acc_0_), .B(
        npu_inst_pe_1_1_2_n13), .ZN(npu_inst_pe_1_1_2_N65) );
  OR2_X1 npu_inst_pe_1_1_2_U139 ( .A1(npu_inst_pe_1_1_2_n13), .A2(
        npu_inst_pe_1_1_2_int_q_acc_0_), .ZN(npu_inst_pe_1_1_2_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_1_2_U138 ( .A(npu_inst_pe_1_1_2_int_q_acc_2_), .B(
        npu_inst_pe_1_1_2_add_79_carry_2_), .Z(npu_inst_pe_1_1_2_N75) );
  AND2_X1 npu_inst_pe_1_1_2_U137 ( .A1(npu_inst_pe_1_1_2_add_79_carry_2_), 
        .A2(npu_inst_pe_1_1_2_int_q_acc_2_), .ZN(
        npu_inst_pe_1_1_2_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_1_2_U136 ( .A(npu_inst_pe_1_1_2_int_q_acc_3_), .B(
        npu_inst_pe_1_1_2_add_79_carry_3_), .Z(npu_inst_pe_1_1_2_N76) );
  AND2_X1 npu_inst_pe_1_1_2_U135 ( .A1(npu_inst_pe_1_1_2_add_79_carry_3_), 
        .A2(npu_inst_pe_1_1_2_int_q_acc_3_), .ZN(
        npu_inst_pe_1_1_2_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_1_2_U134 ( .A(npu_inst_pe_1_1_2_int_q_acc_4_), .B(
        npu_inst_pe_1_1_2_add_79_carry_4_), .Z(npu_inst_pe_1_1_2_N77) );
  AND2_X1 npu_inst_pe_1_1_2_U133 ( .A1(npu_inst_pe_1_1_2_add_79_carry_4_), 
        .A2(npu_inst_pe_1_1_2_int_q_acc_4_), .ZN(
        npu_inst_pe_1_1_2_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_1_2_U132 ( .A(npu_inst_pe_1_1_2_int_q_acc_5_), .B(
        npu_inst_pe_1_1_2_add_79_carry_5_), .Z(npu_inst_pe_1_1_2_N78) );
  AND2_X1 npu_inst_pe_1_1_2_U131 ( .A1(npu_inst_pe_1_1_2_add_79_carry_5_), 
        .A2(npu_inst_pe_1_1_2_int_q_acc_5_), .ZN(
        npu_inst_pe_1_1_2_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_1_2_U130 ( .A(npu_inst_pe_1_1_2_int_q_acc_6_), .B(
        npu_inst_pe_1_1_2_add_79_carry_6_), .Z(npu_inst_pe_1_1_2_N79) );
  AND2_X1 npu_inst_pe_1_1_2_U129 ( .A1(npu_inst_pe_1_1_2_add_79_carry_6_), 
        .A2(npu_inst_pe_1_1_2_int_q_acc_6_), .ZN(
        npu_inst_pe_1_1_2_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_1_2_U128 ( .A(npu_inst_pe_1_1_2_int_q_acc_7_), .B(
        npu_inst_pe_1_1_2_add_79_carry_7_), .Z(npu_inst_pe_1_1_2_N80) );
  XNOR2_X1 npu_inst_pe_1_1_2_U127 ( .A(npu_inst_pe_1_1_2_sub_77_carry_2_), .B(
        npu_inst_pe_1_1_2_int_q_acc_2_), .ZN(npu_inst_pe_1_1_2_N67) );
  OR2_X1 npu_inst_pe_1_1_2_U126 ( .A1(npu_inst_pe_1_1_2_int_q_acc_2_), .A2(
        npu_inst_pe_1_1_2_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_1_2_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_1_2_U125 ( .A(npu_inst_pe_1_1_2_sub_77_carry_3_), .B(
        npu_inst_pe_1_1_2_int_q_acc_3_), .ZN(npu_inst_pe_1_1_2_N68) );
  OR2_X1 npu_inst_pe_1_1_2_U124 ( .A1(npu_inst_pe_1_1_2_int_q_acc_3_), .A2(
        npu_inst_pe_1_1_2_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_1_2_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_1_2_U123 ( .A(npu_inst_pe_1_1_2_sub_77_carry_4_), .B(
        npu_inst_pe_1_1_2_int_q_acc_4_), .ZN(npu_inst_pe_1_1_2_N69) );
  OR2_X1 npu_inst_pe_1_1_2_U122 ( .A1(npu_inst_pe_1_1_2_int_q_acc_4_), .A2(
        npu_inst_pe_1_1_2_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_1_2_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_1_2_U121 ( .A(npu_inst_pe_1_1_2_sub_77_carry_5_), .B(
        npu_inst_pe_1_1_2_int_q_acc_5_), .ZN(npu_inst_pe_1_1_2_N70) );
  OR2_X1 npu_inst_pe_1_1_2_U120 ( .A1(npu_inst_pe_1_1_2_int_q_acc_5_), .A2(
        npu_inst_pe_1_1_2_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_1_2_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_1_2_U119 ( .A(npu_inst_pe_1_1_2_sub_77_carry_6_), .B(
        npu_inst_pe_1_1_2_int_q_acc_6_), .ZN(npu_inst_pe_1_1_2_N71) );
  OR2_X1 npu_inst_pe_1_1_2_U118 ( .A1(npu_inst_pe_1_1_2_int_q_acc_6_), .A2(
        npu_inst_pe_1_1_2_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_1_2_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_1_2_U117 ( .A(npu_inst_pe_1_1_2_int_q_acc_7_), .B(
        npu_inst_pe_1_1_2_sub_77_carry_7_), .ZN(npu_inst_pe_1_1_2_N72) );
  INV_X1 npu_inst_pe_1_1_2_U116 ( .A(npu_inst_n79), .ZN(npu_inst_pe_1_1_2_n7)
         );
  INV_X1 npu_inst_pe_1_1_2_U115 ( .A(npu_inst_pe_1_1_2_n7), .ZN(
        npu_inst_pe_1_1_2_n6) );
  INV_X1 npu_inst_pe_1_1_2_U114 ( .A(npu_inst_n59), .ZN(npu_inst_pe_1_1_2_n3)
         );
  AOI22_X1 npu_inst_pe_1_1_2_U113 ( .A1(npu_inst_int_data_y_2__2__0_), .A2(
        npu_inst_pe_1_1_2_n58), .B1(npu_inst_pe_1_1_2_n114), .B2(
        npu_inst_pe_1_1_2_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_1_2_n57) );
  INV_X1 npu_inst_pe_1_1_2_U112 ( .A(npu_inst_pe_1_1_2_n57), .ZN(
        npu_inst_pe_1_1_2_n108) );
  AOI22_X1 npu_inst_pe_1_1_2_U111 ( .A1(npu_inst_int_data_y_2__2__0_), .A2(
        npu_inst_pe_1_1_2_n54), .B1(npu_inst_pe_1_1_2_n115), .B2(
        npu_inst_pe_1_1_2_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_1_2_n53) );
  INV_X1 npu_inst_pe_1_1_2_U110 ( .A(npu_inst_pe_1_1_2_n53), .ZN(
        npu_inst_pe_1_1_2_n109) );
  AOI22_X1 npu_inst_pe_1_1_2_U107 ( .A1(npu_inst_int_data_y_2__2__0_), .A2(
        npu_inst_pe_1_1_2_n50), .B1(npu_inst_pe_1_1_2_n116), .B2(
        npu_inst_pe_1_1_2_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_1_2_n49) );
  INV_X1 npu_inst_pe_1_1_2_U106 ( .A(npu_inst_pe_1_1_2_n49), .ZN(
        npu_inst_pe_1_1_2_n110) );
  AOI22_X1 npu_inst_pe_1_1_2_U105 ( .A1(npu_inst_int_data_y_2__2__0_), .A2(
        npu_inst_pe_1_1_2_n46), .B1(npu_inst_pe_1_1_2_n117), .B2(
        npu_inst_pe_1_1_2_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_1_2_n45) );
  INV_X1 npu_inst_pe_1_1_2_U104 ( .A(npu_inst_pe_1_1_2_n45), .ZN(
        npu_inst_pe_1_1_2_n111) );
  AOI22_X1 npu_inst_pe_1_1_2_U103 ( .A1(npu_inst_int_data_y_2__2__0_), .A2(
        npu_inst_pe_1_1_2_n42), .B1(npu_inst_pe_1_1_2_n119), .B2(
        npu_inst_pe_1_1_2_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_1_2_n41) );
  INV_X1 npu_inst_pe_1_1_2_U102 ( .A(npu_inst_pe_1_1_2_n41), .ZN(
        npu_inst_pe_1_1_2_n112) );
  AOI22_X1 npu_inst_pe_1_1_2_U101 ( .A1(npu_inst_int_data_y_2__2__1_), .A2(
        npu_inst_pe_1_1_2_n58), .B1(npu_inst_pe_1_1_2_n114), .B2(
        npu_inst_pe_1_1_2_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_1_2_n59) );
  INV_X1 npu_inst_pe_1_1_2_U100 ( .A(npu_inst_pe_1_1_2_n59), .ZN(
        npu_inst_pe_1_1_2_n102) );
  AOI22_X1 npu_inst_pe_1_1_2_U99 ( .A1(npu_inst_int_data_y_2__2__1_), .A2(
        npu_inst_pe_1_1_2_n54), .B1(npu_inst_pe_1_1_2_n115), .B2(
        npu_inst_pe_1_1_2_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_1_2_n55) );
  INV_X1 npu_inst_pe_1_1_2_U98 ( .A(npu_inst_pe_1_1_2_n55), .ZN(
        npu_inst_pe_1_1_2_n103) );
  AOI22_X1 npu_inst_pe_1_1_2_U97 ( .A1(npu_inst_int_data_y_2__2__1_), .A2(
        npu_inst_pe_1_1_2_n50), .B1(npu_inst_pe_1_1_2_n116), .B2(
        npu_inst_pe_1_1_2_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_1_2_n51) );
  INV_X1 npu_inst_pe_1_1_2_U96 ( .A(npu_inst_pe_1_1_2_n51), .ZN(
        npu_inst_pe_1_1_2_n104) );
  AOI22_X1 npu_inst_pe_1_1_2_U95 ( .A1(npu_inst_int_data_y_2__2__1_), .A2(
        npu_inst_pe_1_1_2_n46), .B1(npu_inst_pe_1_1_2_n117), .B2(
        npu_inst_pe_1_1_2_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_1_2_n47) );
  INV_X1 npu_inst_pe_1_1_2_U94 ( .A(npu_inst_pe_1_1_2_n47), .ZN(
        npu_inst_pe_1_1_2_n105) );
  AOI22_X1 npu_inst_pe_1_1_2_U93 ( .A1(npu_inst_int_data_y_2__2__1_), .A2(
        npu_inst_pe_1_1_2_n42), .B1(npu_inst_pe_1_1_2_n119), .B2(
        npu_inst_pe_1_1_2_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_1_2_n43) );
  INV_X1 npu_inst_pe_1_1_2_U92 ( .A(npu_inst_pe_1_1_2_n43), .ZN(
        npu_inst_pe_1_1_2_n106) );
  AOI22_X1 npu_inst_pe_1_1_2_U91 ( .A1(npu_inst_pe_1_1_2_n38), .A2(
        npu_inst_int_data_y_2__2__1_), .B1(npu_inst_pe_1_1_2_n118), .B2(
        npu_inst_pe_1_1_2_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_1_2_n39) );
  INV_X1 npu_inst_pe_1_1_2_U90 ( .A(npu_inst_pe_1_1_2_n39), .ZN(
        npu_inst_pe_1_1_2_n107) );
  AOI22_X1 npu_inst_pe_1_1_2_U89 ( .A1(npu_inst_pe_1_1_2_n38), .A2(
        npu_inst_int_data_y_2__2__0_), .B1(npu_inst_pe_1_1_2_n118), .B2(
        npu_inst_pe_1_1_2_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_1_2_n37) );
  INV_X1 npu_inst_pe_1_1_2_U88 ( .A(npu_inst_pe_1_1_2_n37), .ZN(
        npu_inst_pe_1_1_2_n113) );
  NAND2_X1 npu_inst_pe_1_1_2_U87 ( .A1(npu_inst_pe_1_1_2_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_1_2_n60), .ZN(npu_inst_pe_1_1_2_n74) );
  OAI21_X1 npu_inst_pe_1_1_2_U86 ( .B1(npu_inst_pe_1_1_2_n63), .B2(
        npu_inst_pe_1_1_2_n60), .A(npu_inst_pe_1_1_2_n74), .ZN(
        npu_inst_pe_1_1_2_n97) );
  NAND2_X1 npu_inst_pe_1_1_2_U85 ( .A1(npu_inst_pe_1_1_2_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_1_2_n60), .ZN(npu_inst_pe_1_1_2_n73) );
  OAI21_X1 npu_inst_pe_1_1_2_U84 ( .B1(npu_inst_pe_1_1_2_n61), .B2(
        npu_inst_pe_1_1_2_n60), .A(npu_inst_pe_1_1_2_n73), .ZN(
        npu_inst_pe_1_1_2_n96) );
  NAND2_X1 npu_inst_pe_1_1_2_U83 ( .A1(npu_inst_pe_1_1_2_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_1_2_n56), .ZN(npu_inst_pe_1_1_2_n72) );
  OAI21_X1 npu_inst_pe_1_1_2_U82 ( .B1(npu_inst_pe_1_1_2_n63), .B2(
        npu_inst_pe_1_1_2_n56), .A(npu_inst_pe_1_1_2_n72), .ZN(
        npu_inst_pe_1_1_2_n95) );
  NAND2_X1 npu_inst_pe_1_1_2_U81 ( .A1(npu_inst_pe_1_1_2_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_1_2_n56), .ZN(npu_inst_pe_1_1_2_n71) );
  OAI21_X1 npu_inst_pe_1_1_2_U80 ( .B1(npu_inst_pe_1_1_2_n61), .B2(
        npu_inst_pe_1_1_2_n56), .A(npu_inst_pe_1_1_2_n71), .ZN(
        npu_inst_pe_1_1_2_n94) );
  NAND2_X1 npu_inst_pe_1_1_2_U79 ( .A1(npu_inst_pe_1_1_2_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_1_2_n52), .ZN(npu_inst_pe_1_1_2_n70) );
  OAI21_X1 npu_inst_pe_1_1_2_U78 ( .B1(npu_inst_pe_1_1_2_n63), .B2(
        npu_inst_pe_1_1_2_n52), .A(npu_inst_pe_1_1_2_n70), .ZN(
        npu_inst_pe_1_1_2_n93) );
  NAND2_X1 npu_inst_pe_1_1_2_U77 ( .A1(npu_inst_pe_1_1_2_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_1_2_n52), .ZN(npu_inst_pe_1_1_2_n69) );
  OAI21_X1 npu_inst_pe_1_1_2_U76 ( .B1(npu_inst_pe_1_1_2_n61), .B2(
        npu_inst_pe_1_1_2_n52), .A(npu_inst_pe_1_1_2_n69), .ZN(
        npu_inst_pe_1_1_2_n92) );
  NAND2_X1 npu_inst_pe_1_1_2_U75 ( .A1(npu_inst_pe_1_1_2_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_1_2_n48), .ZN(npu_inst_pe_1_1_2_n68) );
  OAI21_X1 npu_inst_pe_1_1_2_U74 ( .B1(npu_inst_pe_1_1_2_n63), .B2(
        npu_inst_pe_1_1_2_n48), .A(npu_inst_pe_1_1_2_n68), .ZN(
        npu_inst_pe_1_1_2_n91) );
  NAND2_X1 npu_inst_pe_1_1_2_U73 ( .A1(npu_inst_pe_1_1_2_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_1_2_n48), .ZN(npu_inst_pe_1_1_2_n67) );
  OAI21_X1 npu_inst_pe_1_1_2_U72 ( .B1(npu_inst_pe_1_1_2_n61), .B2(
        npu_inst_pe_1_1_2_n48), .A(npu_inst_pe_1_1_2_n67), .ZN(
        npu_inst_pe_1_1_2_n90) );
  NAND2_X1 npu_inst_pe_1_1_2_U71 ( .A1(npu_inst_pe_1_1_2_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_1_2_n44), .ZN(npu_inst_pe_1_1_2_n66) );
  OAI21_X1 npu_inst_pe_1_1_2_U70 ( .B1(npu_inst_pe_1_1_2_n63), .B2(
        npu_inst_pe_1_1_2_n44), .A(npu_inst_pe_1_1_2_n66), .ZN(
        npu_inst_pe_1_1_2_n89) );
  NAND2_X1 npu_inst_pe_1_1_2_U69 ( .A1(npu_inst_pe_1_1_2_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_1_2_n44), .ZN(npu_inst_pe_1_1_2_n65) );
  OAI21_X1 npu_inst_pe_1_1_2_U68 ( .B1(npu_inst_pe_1_1_2_n61), .B2(
        npu_inst_pe_1_1_2_n44), .A(npu_inst_pe_1_1_2_n65), .ZN(
        npu_inst_pe_1_1_2_n88) );
  NAND2_X1 npu_inst_pe_1_1_2_U67 ( .A1(npu_inst_pe_1_1_2_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_1_2_n40), .ZN(npu_inst_pe_1_1_2_n64) );
  OAI21_X1 npu_inst_pe_1_1_2_U66 ( .B1(npu_inst_pe_1_1_2_n63), .B2(
        npu_inst_pe_1_1_2_n40), .A(npu_inst_pe_1_1_2_n64), .ZN(
        npu_inst_pe_1_1_2_n87) );
  NAND2_X1 npu_inst_pe_1_1_2_U65 ( .A1(npu_inst_pe_1_1_2_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_1_2_n40), .ZN(npu_inst_pe_1_1_2_n62) );
  OAI21_X1 npu_inst_pe_1_1_2_U64 ( .B1(npu_inst_pe_1_1_2_n61), .B2(
        npu_inst_pe_1_1_2_n40), .A(npu_inst_pe_1_1_2_n62), .ZN(
        npu_inst_pe_1_1_2_n86) );
  AND2_X1 npu_inst_pe_1_1_2_U63 ( .A1(npu_inst_pe_1_1_2_N93), .A2(npu_inst_n59), .ZN(npu_inst_int_data_y_1__2__0_) );
  AND2_X1 npu_inst_pe_1_1_2_U62 ( .A1(npu_inst_n59), .A2(npu_inst_pe_1_1_2_N94), .ZN(npu_inst_int_data_y_1__2__1_) );
  NOR3_X1 npu_inst_pe_1_1_2_U61 ( .A1(npu_inst_pe_1_1_2_n26), .A2(npu_inst_n59), .A3(npu_inst_int_ckg[53]), .ZN(npu_inst_pe_1_1_2_n85) );
  OR2_X1 npu_inst_pe_1_1_2_U60 ( .A1(npu_inst_pe_1_1_2_n85), .A2(
        npu_inst_pe_1_1_2_n2), .ZN(npu_inst_pe_1_1_2_N84) );
  AND2_X1 npu_inst_pe_1_1_2_U59 ( .A1(npu_inst_pe_1_1_2_int_q_acc_0_), .A2(
        npu_inst_pe_1_1_2_n1), .ZN(npu_inst_int_data_res_1__2__0_) );
  AND2_X1 npu_inst_pe_1_1_2_U58 ( .A1(npu_inst_pe_1_1_2_n2), .A2(
        npu_inst_pe_1_1_2_int_q_acc_7_), .ZN(npu_inst_int_data_res_1__2__7_)
         );
  AND2_X1 npu_inst_pe_1_1_2_U57 ( .A1(npu_inst_pe_1_1_2_int_q_acc_1_), .A2(
        npu_inst_pe_1_1_2_n1), .ZN(npu_inst_int_data_res_1__2__1_) );
  AND2_X1 npu_inst_pe_1_1_2_U56 ( .A1(npu_inst_pe_1_1_2_int_q_acc_2_), .A2(
        npu_inst_pe_1_1_2_n1), .ZN(npu_inst_int_data_res_1__2__2_) );
  AND2_X1 npu_inst_pe_1_1_2_U55 ( .A1(npu_inst_pe_1_1_2_int_q_acc_3_), .A2(
        npu_inst_pe_1_1_2_n2), .ZN(npu_inst_int_data_res_1__2__3_) );
  AND2_X1 npu_inst_pe_1_1_2_U54 ( .A1(npu_inst_pe_1_1_2_int_q_acc_4_), .A2(
        npu_inst_pe_1_1_2_n2), .ZN(npu_inst_int_data_res_1__2__4_) );
  AND2_X1 npu_inst_pe_1_1_2_U53 ( .A1(npu_inst_pe_1_1_2_int_q_acc_5_), .A2(
        npu_inst_pe_1_1_2_n2), .ZN(npu_inst_int_data_res_1__2__5_) );
  AND2_X1 npu_inst_pe_1_1_2_U52 ( .A1(npu_inst_pe_1_1_2_int_q_acc_6_), .A2(
        npu_inst_pe_1_1_2_n2), .ZN(npu_inst_int_data_res_1__2__6_) );
  AOI222_X1 npu_inst_pe_1_1_2_U51 ( .A1(npu_inst_int_data_res_2__2__0_), .A2(
        npu_inst_pe_1_1_2_n1), .B1(npu_inst_pe_1_1_2_N73), .B2(
        npu_inst_pe_1_1_2_n76), .C1(npu_inst_pe_1_1_2_N65), .C2(
        npu_inst_pe_1_1_2_n77), .ZN(npu_inst_pe_1_1_2_n84) );
  INV_X1 npu_inst_pe_1_1_2_U50 ( .A(npu_inst_pe_1_1_2_n84), .ZN(
        npu_inst_pe_1_1_2_n101) );
  AOI222_X1 npu_inst_pe_1_1_2_U49 ( .A1(npu_inst_int_data_res_2__2__7_), .A2(
        npu_inst_pe_1_1_2_n1), .B1(npu_inst_pe_1_1_2_N80), .B2(
        npu_inst_pe_1_1_2_n76), .C1(npu_inst_pe_1_1_2_N72), .C2(
        npu_inst_pe_1_1_2_n77), .ZN(npu_inst_pe_1_1_2_n75) );
  INV_X1 npu_inst_pe_1_1_2_U48 ( .A(npu_inst_pe_1_1_2_n75), .ZN(
        npu_inst_pe_1_1_2_n33) );
  AOI222_X1 npu_inst_pe_1_1_2_U47 ( .A1(npu_inst_int_data_res_2__2__1_), .A2(
        npu_inst_pe_1_1_2_n1), .B1(npu_inst_pe_1_1_2_N74), .B2(
        npu_inst_pe_1_1_2_n76), .C1(npu_inst_pe_1_1_2_N66), .C2(
        npu_inst_pe_1_1_2_n77), .ZN(npu_inst_pe_1_1_2_n83) );
  INV_X1 npu_inst_pe_1_1_2_U46 ( .A(npu_inst_pe_1_1_2_n83), .ZN(
        npu_inst_pe_1_1_2_n100) );
  AOI222_X1 npu_inst_pe_1_1_2_U45 ( .A1(npu_inst_int_data_res_2__2__2_), .A2(
        npu_inst_pe_1_1_2_n1), .B1(npu_inst_pe_1_1_2_N75), .B2(
        npu_inst_pe_1_1_2_n76), .C1(npu_inst_pe_1_1_2_N67), .C2(
        npu_inst_pe_1_1_2_n77), .ZN(npu_inst_pe_1_1_2_n82) );
  INV_X1 npu_inst_pe_1_1_2_U44 ( .A(npu_inst_pe_1_1_2_n82), .ZN(
        npu_inst_pe_1_1_2_n99) );
  AOI222_X1 npu_inst_pe_1_1_2_U43 ( .A1(npu_inst_int_data_res_2__2__3_), .A2(
        npu_inst_pe_1_1_2_n1), .B1(npu_inst_pe_1_1_2_N76), .B2(
        npu_inst_pe_1_1_2_n76), .C1(npu_inst_pe_1_1_2_N68), .C2(
        npu_inst_pe_1_1_2_n77), .ZN(npu_inst_pe_1_1_2_n81) );
  INV_X1 npu_inst_pe_1_1_2_U42 ( .A(npu_inst_pe_1_1_2_n81), .ZN(
        npu_inst_pe_1_1_2_n98) );
  AOI222_X1 npu_inst_pe_1_1_2_U41 ( .A1(npu_inst_int_data_res_2__2__4_), .A2(
        npu_inst_pe_1_1_2_n1), .B1(npu_inst_pe_1_1_2_N77), .B2(
        npu_inst_pe_1_1_2_n76), .C1(npu_inst_pe_1_1_2_N69), .C2(
        npu_inst_pe_1_1_2_n77), .ZN(npu_inst_pe_1_1_2_n80) );
  INV_X1 npu_inst_pe_1_1_2_U40 ( .A(npu_inst_pe_1_1_2_n80), .ZN(
        npu_inst_pe_1_1_2_n36) );
  AOI222_X1 npu_inst_pe_1_1_2_U39 ( .A1(npu_inst_int_data_res_2__2__5_), .A2(
        npu_inst_pe_1_1_2_n1), .B1(npu_inst_pe_1_1_2_N78), .B2(
        npu_inst_pe_1_1_2_n76), .C1(npu_inst_pe_1_1_2_N70), .C2(
        npu_inst_pe_1_1_2_n77), .ZN(npu_inst_pe_1_1_2_n79) );
  INV_X1 npu_inst_pe_1_1_2_U38 ( .A(npu_inst_pe_1_1_2_n79), .ZN(
        npu_inst_pe_1_1_2_n35) );
  AOI222_X1 npu_inst_pe_1_1_2_U37 ( .A1(npu_inst_int_data_res_2__2__6_), .A2(
        npu_inst_pe_1_1_2_n1), .B1(npu_inst_pe_1_1_2_N79), .B2(
        npu_inst_pe_1_1_2_n76), .C1(npu_inst_pe_1_1_2_N71), .C2(
        npu_inst_pe_1_1_2_n77), .ZN(npu_inst_pe_1_1_2_n78) );
  INV_X1 npu_inst_pe_1_1_2_U36 ( .A(npu_inst_pe_1_1_2_n78), .ZN(
        npu_inst_pe_1_1_2_n34) );
  INV_X1 npu_inst_pe_1_1_2_U35 ( .A(npu_inst_pe_1_1_2_int_data_1_), .ZN(
        npu_inst_pe_1_1_2_n14) );
  AND2_X1 npu_inst_pe_1_1_2_U34 ( .A1(npu_inst_int_data_x_1__2__1_), .A2(
        npu_inst_pe_1_1_2_int_q_weight_1_), .ZN(npu_inst_pe_1_1_2_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_1_2_U33 ( .A1(npu_inst_int_data_x_1__2__0_), .A2(
        npu_inst_pe_1_1_2_int_q_weight_1_), .ZN(npu_inst_pe_1_1_2_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_1_2_U32 ( .A1(npu_inst_n59), .A2(
        npu_inst_int_data_y_2__2__1_), .B1(npu_inst_pe_1_1_2_n3), .B2(
        npu_inst_int_data_x_1__3__1_), .ZN(npu_inst_pe_1_1_2_n63) );
  AOI22_X1 npu_inst_pe_1_1_2_U31 ( .A1(npu_inst_n59), .A2(
        npu_inst_int_data_y_2__2__0_), .B1(npu_inst_pe_1_1_2_n3), .B2(
        npu_inst_int_data_x_1__3__0_), .ZN(npu_inst_pe_1_1_2_n61) );
  INV_X1 npu_inst_pe_1_1_2_U30 ( .A(npu_inst_pe_1_1_2_int_data_0_), .ZN(
        npu_inst_pe_1_1_2_n13) );
  INV_X1 npu_inst_pe_1_1_2_U29 ( .A(npu_inst_n71), .ZN(npu_inst_pe_1_1_2_n5)
         );
  OR3_X1 npu_inst_pe_1_1_2_U28 ( .A1(npu_inst_pe_1_1_2_n6), .A2(
        npu_inst_pe_1_1_2_n8), .A3(npu_inst_pe_1_1_2_n5), .ZN(
        npu_inst_pe_1_1_2_n56) );
  OR3_X1 npu_inst_pe_1_1_2_U27 ( .A1(npu_inst_pe_1_1_2_n5), .A2(
        npu_inst_pe_1_1_2_n8), .A3(npu_inst_pe_1_1_2_n7), .ZN(
        npu_inst_pe_1_1_2_n48) );
  INV_X1 npu_inst_pe_1_1_2_U26 ( .A(npu_inst_pe_1_1_2_n5), .ZN(
        npu_inst_pe_1_1_2_n4) );
  INV_X1 npu_inst_pe_1_1_2_U25 ( .A(npu_inst_n126), .ZN(npu_inst_pe_1_1_2_n12)
         );
  OR3_X1 npu_inst_pe_1_1_2_U24 ( .A1(npu_inst_pe_1_1_2_n4), .A2(
        npu_inst_pe_1_1_2_n8), .A3(npu_inst_pe_1_1_2_n7), .ZN(
        npu_inst_pe_1_1_2_n52) );
  OR3_X1 npu_inst_pe_1_1_2_U23 ( .A1(npu_inst_pe_1_1_2_n6), .A2(
        npu_inst_pe_1_1_2_n8), .A3(npu_inst_pe_1_1_2_n4), .ZN(
        npu_inst_pe_1_1_2_n60) );
  NOR2_X1 npu_inst_pe_1_1_2_U22 ( .A1(npu_inst_pe_1_1_2_n60), .A2(
        npu_inst_pe_1_1_2_n3), .ZN(npu_inst_pe_1_1_2_n58) );
  NOR2_X1 npu_inst_pe_1_1_2_U21 ( .A1(npu_inst_pe_1_1_2_n56), .A2(
        npu_inst_pe_1_1_2_n3), .ZN(npu_inst_pe_1_1_2_n54) );
  NOR2_X1 npu_inst_pe_1_1_2_U20 ( .A1(npu_inst_pe_1_1_2_n52), .A2(
        npu_inst_pe_1_1_2_n3), .ZN(npu_inst_pe_1_1_2_n50) );
  NOR2_X1 npu_inst_pe_1_1_2_U19 ( .A1(npu_inst_pe_1_1_2_n48), .A2(
        npu_inst_pe_1_1_2_n3), .ZN(npu_inst_pe_1_1_2_n46) );
  NOR2_X1 npu_inst_pe_1_1_2_U18 ( .A1(npu_inst_pe_1_1_2_n40), .A2(
        npu_inst_pe_1_1_2_n3), .ZN(npu_inst_pe_1_1_2_n38) );
  NOR2_X1 npu_inst_pe_1_1_2_U17 ( .A1(npu_inst_pe_1_1_2_n44), .A2(
        npu_inst_pe_1_1_2_n3), .ZN(npu_inst_pe_1_1_2_n42) );
  BUF_X1 npu_inst_pe_1_1_2_U16 ( .A(npu_inst_n105), .Z(npu_inst_pe_1_1_2_n8)
         );
  BUF_X1 npu_inst_pe_1_1_2_U15 ( .A(npu_inst_pe_1_1_2_n12), .Z(
        npu_inst_pe_1_1_2_n11) );
  BUF_X1 npu_inst_pe_1_1_2_U14 ( .A(npu_inst_pe_1_1_2_n12), .Z(
        npu_inst_pe_1_1_2_n10) );
  BUF_X1 npu_inst_pe_1_1_2_U13 ( .A(npu_inst_pe_1_1_2_n12), .Z(
        npu_inst_pe_1_1_2_n9) );
  INV_X1 npu_inst_pe_1_1_2_U12 ( .A(npu_inst_pe_1_1_2_n38), .ZN(
        npu_inst_pe_1_1_2_n118) );
  INV_X1 npu_inst_pe_1_1_2_U11 ( .A(npu_inst_pe_1_1_2_n58), .ZN(
        npu_inst_pe_1_1_2_n114) );
  INV_X1 npu_inst_pe_1_1_2_U10 ( .A(npu_inst_pe_1_1_2_n54), .ZN(
        npu_inst_pe_1_1_2_n115) );
  INV_X1 npu_inst_pe_1_1_2_U9 ( .A(npu_inst_pe_1_1_2_n50), .ZN(
        npu_inst_pe_1_1_2_n116) );
  INV_X1 npu_inst_pe_1_1_2_U8 ( .A(npu_inst_pe_1_1_2_n46), .ZN(
        npu_inst_pe_1_1_2_n117) );
  INV_X1 npu_inst_pe_1_1_2_U7 ( .A(npu_inst_pe_1_1_2_n42), .ZN(
        npu_inst_pe_1_1_2_n119) );
  BUF_X1 npu_inst_pe_1_1_2_U6 ( .A(npu_inst_n33), .Z(npu_inst_pe_1_1_2_n2) );
  BUF_X1 npu_inst_pe_1_1_2_U5 ( .A(npu_inst_n33), .Z(npu_inst_pe_1_1_2_n1) );
  NOR2_X1 npu_inst_pe_1_1_2_U4 ( .A1(npu_inst_pe_1_1_2_int_q_weight_0_), .A2(
        npu_inst_pe_1_1_2_n1), .ZN(npu_inst_pe_1_1_2_n76) );
  NOR2_X1 npu_inst_pe_1_1_2_U3 ( .A1(npu_inst_pe_1_1_2_n27), .A2(
        npu_inst_pe_1_1_2_n1), .ZN(npu_inst_pe_1_1_2_n77) );
  FA_X1 npu_inst_pe_1_1_2_sub_77_U2_1 ( .A(npu_inst_pe_1_1_2_int_q_acc_1_), 
        .B(npu_inst_pe_1_1_2_n14), .CI(npu_inst_pe_1_1_2_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_1_2_sub_77_carry_2_), .S(npu_inst_pe_1_1_2_N66) );
  FA_X1 npu_inst_pe_1_1_2_add_79_U1_1 ( .A(npu_inst_pe_1_1_2_int_q_acc_1_), 
        .B(npu_inst_pe_1_1_2_int_data_1_), .CI(
        npu_inst_pe_1_1_2_add_79_carry_1_), .CO(
        npu_inst_pe_1_1_2_add_79_carry_2_), .S(npu_inst_pe_1_1_2_N74) );
  NAND3_X1 npu_inst_pe_1_1_2_U109 ( .A1(npu_inst_pe_1_1_2_n5), .A2(
        npu_inst_pe_1_1_2_n7), .A3(npu_inst_pe_1_1_2_n8), .ZN(
        npu_inst_pe_1_1_2_n44) );
  NAND3_X1 npu_inst_pe_1_1_2_U108 ( .A1(npu_inst_pe_1_1_2_n4), .A2(
        npu_inst_pe_1_1_2_n7), .A3(npu_inst_pe_1_1_2_n8), .ZN(
        npu_inst_pe_1_1_2_n40) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_1_2_n34), .CK(
        npu_inst_pe_1_1_2_net4063), .RN(npu_inst_pe_1_1_2_n9), .Q(
        npu_inst_pe_1_1_2_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_1_2_n35), .CK(
        npu_inst_pe_1_1_2_net4063), .RN(npu_inst_pe_1_1_2_n9), .Q(
        npu_inst_pe_1_1_2_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_1_2_n36), .CK(
        npu_inst_pe_1_1_2_net4063), .RN(npu_inst_pe_1_1_2_n9), .Q(
        npu_inst_pe_1_1_2_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_1_2_n98), .CK(
        npu_inst_pe_1_1_2_net4063), .RN(npu_inst_pe_1_1_2_n9), .Q(
        npu_inst_pe_1_1_2_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_1_2_n99), .CK(
        npu_inst_pe_1_1_2_net4063), .RN(npu_inst_pe_1_1_2_n9), .Q(
        npu_inst_pe_1_1_2_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_1_2_n100), 
        .CK(npu_inst_pe_1_1_2_net4063), .RN(npu_inst_pe_1_1_2_n9), .Q(
        npu_inst_pe_1_1_2_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_1_2_n33), .CK(
        npu_inst_pe_1_1_2_net4063), .RN(npu_inst_pe_1_1_2_n9), .Q(
        npu_inst_pe_1_1_2_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_1_2_n101), 
        .CK(npu_inst_pe_1_1_2_net4063), .RN(npu_inst_pe_1_1_2_n9), .Q(
        npu_inst_pe_1_1_2_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_weight_reg_0_ ( .D(npu_inst_n112), .CK(
        npu_inst_pe_1_1_2_net4069), .RN(npu_inst_pe_1_1_2_n9), .Q(
        npu_inst_pe_1_1_2_int_q_weight_0_), .QN(npu_inst_pe_1_1_2_n27) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_weight_reg_1_ ( .D(npu_inst_n118), .CK(
        npu_inst_pe_1_1_2_net4069), .RN(npu_inst_pe_1_1_2_n9), .Q(
        npu_inst_pe_1_1_2_int_q_weight_1_), .QN(npu_inst_pe_1_1_2_n26) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_1_2_n113), 
        .CK(npu_inst_pe_1_1_2_net4069), .RN(npu_inst_pe_1_1_2_n9), .Q(
        npu_inst_pe_1_1_2_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_1_2_n107), 
        .CK(npu_inst_pe_1_1_2_net4069), .RN(npu_inst_pe_1_1_2_n9), .Q(
        npu_inst_pe_1_1_2_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_1_2_n112), 
        .CK(npu_inst_pe_1_1_2_net4069), .RN(npu_inst_pe_1_1_2_n10), .Q(
        npu_inst_pe_1_1_2_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_1_2_n106), 
        .CK(npu_inst_pe_1_1_2_net4069), .RN(npu_inst_pe_1_1_2_n10), .Q(
        npu_inst_pe_1_1_2_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_1_2_n111), 
        .CK(npu_inst_pe_1_1_2_net4069), .RN(npu_inst_pe_1_1_2_n10), .Q(
        npu_inst_pe_1_1_2_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_1_2_n105), 
        .CK(npu_inst_pe_1_1_2_net4069), .RN(npu_inst_pe_1_1_2_n10), .Q(
        npu_inst_pe_1_1_2_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_1_2_n110), 
        .CK(npu_inst_pe_1_1_2_net4069), .RN(npu_inst_pe_1_1_2_n10), .Q(
        npu_inst_pe_1_1_2_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_1_2_n104), 
        .CK(npu_inst_pe_1_1_2_net4069), .RN(npu_inst_pe_1_1_2_n10), .Q(
        npu_inst_pe_1_1_2_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_1_2_n109), 
        .CK(npu_inst_pe_1_1_2_net4069), .RN(npu_inst_pe_1_1_2_n10), .Q(
        npu_inst_pe_1_1_2_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_1_2_n103), 
        .CK(npu_inst_pe_1_1_2_net4069), .RN(npu_inst_pe_1_1_2_n10), .Q(
        npu_inst_pe_1_1_2_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_1_2_n108), 
        .CK(npu_inst_pe_1_1_2_net4069), .RN(npu_inst_pe_1_1_2_n10), .Q(
        npu_inst_pe_1_1_2_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_1_2_n102), 
        .CK(npu_inst_pe_1_1_2_net4069), .RN(npu_inst_pe_1_1_2_n10), .Q(
        npu_inst_pe_1_1_2_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_1_2_n86), 
        .CK(npu_inst_pe_1_1_2_net4069), .RN(npu_inst_pe_1_1_2_n10), .Q(
        npu_inst_pe_1_1_2_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_1_2_n87), 
        .CK(npu_inst_pe_1_1_2_net4069), .RN(npu_inst_pe_1_1_2_n10), .Q(
        npu_inst_pe_1_1_2_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_1_2_n88), 
        .CK(npu_inst_pe_1_1_2_net4069), .RN(npu_inst_pe_1_1_2_n11), .Q(
        npu_inst_pe_1_1_2_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_1_2_n89), 
        .CK(npu_inst_pe_1_1_2_net4069), .RN(npu_inst_pe_1_1_2_n11), .Q(
        npu_inst_pe_1_1_2_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_1_2_n90), 
        .CK(npu_inst_pe_1_1_2_net4069), .RN(npu_inst_pe_1_1_2_n11), .Q(
        npu_inst_pe_1_1_2_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_1_2_n91), 
        .CK(npu_inst_pe_1_1_2_net4069), .RN(npu_inst_pe_1_1_2_n11), .Q(
        npu_inst_pe_1_1_2_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_1_2_n92), 
        .CK(npu_inst_pe_1_1_2_net4069), .RN(npu_inst_pe_1_1_2_n11), .Q(
        npu_inst_pe_1_1_2_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_1_2_n93), 
        .CK(npu_inst_pe_1_1_2_net4069), .RN(npu_inst_pe_1_1_2_n11), .Q(
        npu_inst_pe_1_1_2_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_1_2_n94), 
        .CK(npu_inst_pe_1_1_2_net4069), .RN(npu_inst_pe_1_1_2_n11), .Q(
        npu_inst_pe_1_1_2_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_1_2_n95), 
        .CK(npu_inst_pe_1_1_2_net4069), .RN(npu_inst_pe_1_1_2_n11), .Q(
        npu_inst_pe_1_1_2_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_1_2_n96), 
        .CK(npu_inst_pe_1_1_2_net4069), .RN(npu_inst_pe_1_1_2_n11), .Q(
        npu_inst_pe_1_1_2_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_1_2_n97), 
        .CK(npu_inst_pe_1_1_2_net4069), .RN(npu_inst_pe_1_1_2_n11), .Q(
        npu_inst_pe_1_1_2_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_1_2_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_1_2_N84), .SE(1'b0), .GCK(npu_inst_pe_1_1_2_net4063) );
  CLKGATETST_X1 npu_inst_pe_1_1_2_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n65), .SE(1'b0), .GCK(npu_inst_pe_1_1_2_net4069) );
  MUX2_X1 npu_inst_pe_1_1_3_U162 ( .A(npu_inst_pe_1_1_3_n32), .B(
        npu_inst_pe_1_1_3_n29), .S(npu_inst_pe_1_1_3_n8), .Z(
        npu_inst_pe_1_1_3_N93) );
  MUX2_X1 npu_inst_pe_1_1_3_U161 ( .A(npu_inst_pe_1_1_3_n31), .B(
        npu_inst_pe_1_1_3_n30), .S(npu_inst_pe_1_1_3_n6), .Z(
        npu_inst_pe_1_1_3_n32) );
  MUX2_X1 npu_inst_pe_1_1_3_U160 ( .A(npu_inst_pe_1_1_3_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_1_3_int_q_reg_v_1__0_), .S(npu_inst_pe_1_1_3_n4), .Z(
        npu_inst_pe_1_1_3_n31) );
  MUX2_X1 npu_inst_pe_1_1_3_U159 ( .A(npu_inst_pe_1_1_3_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_1_3_int_q_reg_v_3__0_), .S(npu_inst_pe_1_1_3_n4), .Z(
        npu_inst_pe_1_1_3_n30) );
  MUX2_X1 npu_inst_pe_1_1_3_U158 ( .A(npu_inst_pe_1_1_3_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_1_3_int_q_reg_v_5__0_), .S(npu_inst_pe_1_1_3_n4), .Z(
        npu_inst_pe_1_1_3_n29) );
  MUX2_X1 npu_inst_pe_1_1_3_U157 ( .A(npu_inst_pe_1_1_3_n28), .B(
        npu_inst_pe_1_1_3_n23), .S(npu_inst_pe_1_1_3_n8), .Z(
        npu_inst_pe_1_1_3_N94) );
  MUX2_X1 npu_inst_pe_1_1_3_U156 ( .A(npu_inst_pe_1_1_3_n25), .B(
        npu_inst_pe_1_1_3_n24), .S(npu_inst_pe_1_1_3_n6), .Z(
        npu_inst_pe_1_1_3_n28) );
  MUX2_X1 npu_inst_pe_1_1_3_U155 ( .A(npu_inst_pe_1_1_3_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_1_3_int_q_reg_v_1__1_), .S(npu_inst_pe_1_1_3_n4), .Z(
        npu_inst_pe_1_1_3_n25) );
  MUX2_X1 npu_inst_pe_1_1_3_U154 ( .A(npu_inst_pe_1_1_3_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_1_3_int_q_reg_v_3__1_), .S(npu_inst_pe_1_1_3_n4), .Z(
        npu_inst_pe_1_1_3_n24) );
  MUX2_X1 npu_inst_pe_1_1_3_U153 ( .A(npu_inst_pe_1_1_3_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_1_3_int_q_reg_v_5__1_), .S(npu_inst_pe_1_1_3_n4), .Z(
        npu_inst_pe_1_1_3_n23) );
  MUX2_X1 npu_inst_pe_1_1_3_U152 ( .A(npu_inst_pe_1_1_3_n22), .B(
        npu_inst_pe_1_1_3_n19), .S(npu_inst_pe_1_1_3_n8), .Z(
        npu_inst_int_data_x_1__3__1_) );
  MUX2_X1 npu_inst_pe_1_1_3_U151 ( .A(npu_inst_pe_1_1_3_n21), .B(
        npu_inst_pe_1_1_3_n20), .S(npu_inst_pe_1_1_3_n6), .Z(
        npu_inst_pe_1_1_3_n22) );
  MUX2_X1 npu_inst_pe_1_1_3_U150 ( .A(npu_inst_pe_1_1_3_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_1_3_int_q_reg_h_1__1_), .S(npu_inst_pe_1_1_3_n4), .Z(
        npu_inst_pe_1_1_3_n21) );
  MUX2_X1 npu_inst_pe_1_1_3_U149 ( .A(npu_inst_pe_1_1_3_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_1_3_int_q_reg_h_3__1_), .S(npu_inst_pe_1_1_3_n4), .Z(
        npu_inst_pe_1_1_3_n20) );
  MUX2_X1 npu_inst_pe_1_1_3_U148 ( .A(npu_inst_pe_1_1_3_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_1_3_int_q_reg_h_5__1_), .S(npu_inst_pe_1_1_3_n4), .Z(
        npu_inst_pe_1_1_3_n19) );
  MUX2_X1 npu_inst_pe_1_1_3_U147 ( .A(npu_inst_pe_1_1_3_n18), .B(
        npu_inst_pe_1_1_3_n15), .S(npu_inst_pe_1_1_3_n8), .Z(
        npu_inst_int_data_x_1__3__0_) );
  MUX2_X1 npu_inst_pe_1_1_3_U146 ( .A(npu_inst_pe_1_1_3_n17), .B(
        npu_inst_pe_1_1_3_n16), .S(npu_inst_pe_1_1_3_n6), .Z(
        npu_inst_pe_1_1_3_n18) );
  MUX2_X1 npu_inst_pe_1_1_3_U145 ( .A(npu_inst_pe_1_1_3_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_1_3_int_q_reg_h_1__0_), .S(npu_inst_pe_1_1_3_n4), .Z(
        npu_inst_pe_1_1_3_n17) );
  MUX2_X1 npu_inst_pe_1_1_3_U144 ( .A(npu_inst_pe_1_1_3_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_1_3_int_q_reg_h_3__0_), .S(npu_inst_pe_1_1_3_n4), .Z(
        npu_inst_pe_1_1_3_n16) );
  MUX2_X1 npu_inst_pe_1_1_3_U143 ( .A(npu_inst_pe_1_1_3_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_1_3_int_q_reg_h_5__0_), .S(npu_inst_pe_1_1_3_n4), .Z(
        npu_inst_pe_1_1_3_n15) );
  XOR2_X1 npu_inst_pe_1_1_3_U142 ( .A(npu_inst_pe_1_1_3_int_data_0_), .B(
        npu_inst_pe_1_1_3_int_q_acc_0_), .Z(npu_inst_pe_1_1_3_N73) );
  AND2_X1 npu_inst_pe_1_1_3_U141 ( .A1(npu_inst_pe_1_1_3_int_q_acc_0_), .A2(
        npu_inst_pe_1_1_3_int_data_0_), .ZN(npu_inst_pe_1_1_3_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_1_3_U140 ( .A(npu_inst_pe_1_1_3_int_q_acc_0_), .B(
        npu_inst_pe_1_1_3_n13), .ZN(npu_inst_pe_1_1_3_N65) );
  OR2_X1 npu_inst_pe_1_1_3_U139 ( .A1(npu_inst_pe_1_1_3_n13), .A2(
        npu_inst_pe_1_1_3_int_q_acc_0_), .ZN(npu_inst_pe_1_1_3_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_1_3_U138 ( .A(npu_inst_pe_1_1_3_int_q_acc_2_), .B(
        npu_inst_pe_1_1_3_add_79_carry_2_), .Z(npu_inst_pe_1_1_3_N75) );
  AND2_X1 npu_inst_pe_1_1_3_U137 ( .A1(npu_inst_pe_1_1_3_add_79_carry_2_), 
        .A2(npu_inst_pe_1_1_3_int_q_acc_2_), .ZN(
        npu_inst_pe_1_1_3_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_1_3_U136 ( .A(npu_inst_pe_1_1_3_int_q_acc_3_), .B(
        npu_inst_pe_1_1_3_add_79_carry_3_), .Z(npu_inst_pe_1_1_3_N76) );
  AND2_X1 npu_inst_pe_1_1_3_U135 ( .A1(npu_inst_pe_1_1_3_add_79_carry_3_), 
        .A2(npu_inst_pe_1_1_3_int_q_acc_3_), .ZN(
        npu_inst_pe_1_1_3_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_1_3_U134 ( .A(npu_inst_pe_1_1_3_int_q_acc_4_), .B(
        npu_inst_pe_1_1_3_add_79_carry_4_), .Z(npu_inst_pe_1_1_3_N77) );
  AND2_X1 npu_inst_pe_1_1_3_U133 ( .A1(npu_inst_pe_1_1_3_add_79_carry_4_), 
        .A2(npu_inst_pe_1_1_3_int_q_acc_4_), .ZN(
        npu_inst_pe_1_1_3_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_1_3_U132 ( .A(npu_inst_pe_1_1_3_int_q_acc_5_), .B(
        npu_inst_pe_1_1_3_add_79_carry_5_), .Z(npu_inst_pe_1_1_3_N78) );
  AND2_X1 npu_inst_pe_1_1_3_U131 ( .A1(npu_inst_pe_1_1_3_add_79_carry_5_), 
        .A2(npu_inst_pe_1_1_3_int_q_acc_5_), .ZN(
        npu_inst_pe_1_1_3_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_1_3_U130 ( .A(npu_inst_pe_1_1_3_int_q_acc_6_), .B(
        npu_inst_pe_1_1_3_add_79_carry_6_), .Z(npu_inst_pe_1_1_3_N79) );
  AND2_X1 npu_inst_pe_1_1_3_U129 ( .A1(npu_inst_pe_1_1_3_add_79_carry_6_), 
        .A2(npu_inst_pe_1_1_3_int_q_acc_6_), .ZN(
        npu_inst_pe_1_1_3_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_1_3_U128 ( .A(npu_inst_pe_1_1_3_int_q_acc_7_), .B(
        npu_inst_pe_1_1_3_add_79_carry_7_), .Z(npu_inst_pe_1_1_3_N80) );
  XNOR2_X1 npu_inst_pe_1_1_3_U127 ( .A(npu_inst_pe_1_1_3_sub_77_carry_2_), .B(
        npu_inst_pe_1_1_3_int_q_acc_2_), .ZN(npu_inst_pe_1_1_3_N67) );
  OR2_X1 npu_inst_pe_1_1_3_U126 ( .A1(npu_inst_pe_1_1_3_int_q_acc_2_), .A2(
        npu_inst_pe_1_1_3_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_1_3_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_1_3_U125 ( .A(npu_inst_pe_1_1_3_sub_77_carry_3_), .B(
        npu_inst_pe_1_1_3_int_q_acc_3_), .ZN(npu_inst_pe_1_1_3_N68) );
  OR2_X1 npu_inst_pe_1_1_3_U124 ( .A1(npu_inst_pe_1_1_3_int_q_acc_3_), .A2(
        npu_inst_pe_1_1_3_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_1_3_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_1_3_U123 ( .A(npu_inst_pe_1_1_3_sub_77_carry_4_), .B(
        npu_inst_pe_1_1_3_int_q_acc_4_), .ZN(npu_inst_pe_1_1_3_N69) );
  OR2_X1 npu_inst_pe_1_1_3_U122 ( .A1(npu_inst_pe_1_1_3_int_q_acc_4_), .A2(
        npu_inst_pe_1_1_3_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_1_3_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_1_3_U121 ( .A(npu_inst_pe_1_1_3_sub_77_carry_5_), .B(
        npu_inst_pe_1_1_3_int_q_acc_5_), .ZN(npu_inst_pe_1_1_3_N70) );
  OR2_X1 npu_inst_pe_1_1_3_U120 ( .A1(npu_inst_pe_1_1_3_int_q_acc_5_), .A2(
        npu_inst_pe_1_1_3_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_1_3_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_1_3_U119 ( .A(npu_inst_pe_1_1_3_sub_77_carry_6_), .B(
        npu_inst_pe_1_1_3_int_q_acc_6_), .ZN(npu_inst_pe_1_1_3_N71) );
  OR2_X1 npu_inst_pe_1_1_3_U118 ( .A1(npu_inst_pe_1_1_3_int_q_acc_6_), .A2(
        npu_inst_pe_1_1_3_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_1_3_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_1_3_U117 ( .A(npu_inst_pe_1_1_3_int_q_acc_7_), .B(
        npu_inst_pe_1_1_3_sub_77_carry_7_), .ZN(npu_inst_pe_1_1_3_N72) );
  INV_X1 npu_inst_pe_1_1_3_U116 ( .A(npu_inst_n79), .ZN(npu_inst_pe_1_1_3_n7)
         );
  INV_X1 npu_inst_pe_1_1_3_U115 ( .A(npu_inst_pe_1_1_3_n7), .ZN(
        npu_inst_pe_1_1_3_n6) );
  INV_X1 npu_inst_pe_1_1_3_U114 ( .A(npu_inst_n59), .ZN(npu_inst_pe_1_1_3_n3)
         );
  AOI22_X1 npu_inst_pe_1_1_3_U113 ( .A1(npu_inst_int_data_y_2__3__0_), .A2(
        npu_inst_pe_1_1_3_n58), .B1(npu_inst_pe_1_1_3_n114), .B2(
        npu_inst_pe_1_1_3_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_1_3_n57) );
  INV_X1 npu_inst_pe_1_1_3_U112 ( .A(npu_inst_pe_1_1_3_n57), .ZN(
        npu_inst_pe_1_1_3_n108) );
  AOI22_X1 npu_inst_pe_1_1_3_U111 ( .A1(npu_inst_int_data_y_2__3__0_), .A2(
        npu_inst_pe_1_1_3_n54), .B1(npu_inst_pe_1_1_3_n115), .B2(
        npu_inst_pe_1_1_3_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_1_3_n53) );
  INV_X1 npu_inst_pe_1_1_3_U110 ( .A(npu_inst_pe_1_1_3_n53), .ZN(
        npu_inst_pe_1_1_3_n109) );
  AOI22_X1 npu_inst_pe_1_1_3_U107 ( .A1(npu_inst_int_data_y_2__3__0_), .A2(
        npu_inst_pe_1_1_3_n50), .B1(npu_inst_pe_1_1_3_n116), .B2(
        npu_inst_pe_1_1_3_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_1_3_n49) );
  INV_X1 npu_inst_pe_1_1_3_U106 ( .A(npu_inst_pe_1_1_3_n49), .ZN(
        npu_inst_pe_1_1_3_n110) );
  AOI22_X1 npu_inst_pe_1_1_3_U105 ( .A1(npu_inst_int_data_y_2__3__0_), .A2(
        npu_inst_pe_1_1_3_n46), .B1(npu_inst_pe_1_1_3_n117), .B2(
        npu_inst_pe_1_1_3_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_1_3_n45) );
  INV_X1 npu_inst_pe_1_1_3_U104 ( .A(npu_inst_pe_1_1_3_n45), .ZN(
        npu_inst_pe_1_1_3_n111) );
  AOI22_X1 npu_inst_pe_1_1_3_U103 ( .A1(npu_inst_int_data_y_2__3__0_), .A2(
        npu_inst_pe_1_1_3_n42), .B1(npu_inst_pe_1_1_3_n119), .B2(
        npu_inst_pe_1_1_3_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_1_3_n41) );
  INV_X1 npu_inst_pe_1_1_3_U102 ( .A(npu_inst_pe_1_1_3_n41), .ZN(
        npu_inst_pe_1_1_3_n112) );
  AOI22_X1 npu_inst_pe_1_1_3_U101 ( .A1(npu_inst_int_data_y_2__3__1_), .A2(
        npu_inst_pe_1_1_3_n58), .B1(npu_inst_pe_1_1_3_n114), .B2(
        npu_inst_pe_1_1_3_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_1_3_n59) );
  INV_X1 npu_inst_pe_1_1_3_U100 ( .A(npu_inst_pe_1_1_3_n59), .ZN(
        npu_inst_pe_1_1_3_n102) );
  AOI22_X1 npu_inst_pe_1_1_3_U99 ( .A1(npu_inst_int_data_y_2__3__1_), .A2(
        npu_inst_pe_1_1_3_n54), .B1(npu_inst_pe_1_1_3_n115), .B2(
        npu_inst_pe_1_1_3_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_1_3_n55) );
  INV_X1 npu_inst_pe_1_1_3_U98 ( .A(npu_inst_pe_1_1_3_n55), .ZN(
        npu_inst_pe_1_1_3_n103) );
  AOI22_X1 npu_inst_pe_1_1_3_U97 ( .A1(npu_inst_int_data_y_2__3__1_), .A2(
        npu_inst_pe_1_1_3_n50), .B1(npu_inst_pe_1_1_3_n116), .B2(
        npu_inst_pe_1_1_3_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_1_3_n51) );
  INV_X1 npu_inst_pe_1_1_3_U96 ( .A(npu_inst_pe_1_1_3_n51), .ZN(
        npu_inst_pe_1_1_3_n104) );
  AOI22_X1 npu_inst_pe_1_1_3_U95 ( .A1(npu_inst_int_data_y_2__3__1_), .A2(
        npu_inst_pe_1_1_3_n46), .B1(npu_inst_pe_1_1_3_n117), .B2(
        npu_inst_pe_1_1_3_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_1_3_n47) );
  INV_X1 npu_inst_pe_1_1_3_U94 ( .A(npu_inst_pe_1_1_3_n47), .ZN(
        npu_inst_pe_1_1_3_n105) );
  AOI22_X1 npu_inst_pe_1_1_3_U93 ( .A1(npu_inst_int_data_y_2__3__1_), .A2(
        npu_inst_pe_1_1_3_n42), .B1(npu_inst_pe_1_1_3_n119), .B2(
        npu_inst_pe_1_1_3_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_1_3_n43) );
  INV_X1 npu_inst_pe_1_1_3_U92 ( .A(npu_inst_pe_1_1_3_n43), .ZN(
        npu_inst_pe_1_1_3_n106) );
  AOI22_X1 npu_inst_pe_1_1_3_U91 ( .A1(npu_inst_pe_1_1_3_n38), .A2(
        npu_inst_int_data_y_2__3__1_), .B1(npu_inst_pe_1_1_3_n118), .B2(
        npu_inst_pe_1_1_3_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_1_3_n39) );
  INV_X1 npu_inst_pe_1_1_3_U90 ( .A(npu_inst_pe_1_1_3_n39), .ZN(
        npu_inst_pe_1_1_3_n107) );
  AOI22_X1 npu_inst_pe_1_1_3_U89 ( .A1(npu_inst_pe_1_1_3_n38), .A2(
        npu_inst_int_data_y_2__3__0_), .B1(npu_inst_pe_1_1_3_n118), .B2(
        npu_inst_pe_1_1_3_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_1_3_n37) );
  INV_X1 npu_inst_pe_1_1_3_U88 ( .A(npu_inst_pe_1_1_3_n37), .ZN(
        npu_inst_pe_1_1_3_n113) );
  NAND2_X1 npu_inst_pe_1_1_3_U87 ( .A1(npu_inst_pe_1_1_3_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_1_3_n60), .ZN(npu_inst_pe_1_1_3_n74) );
  OAI21_X1 npu_inst_pe_1_1_3_U86 ( .B1(npu_inst_pe_1_1_3_n63), .B2(
        npu_inst_pe_1_1_3_n60), .A(npu_inst_pe_1_1_3_n74), .ZN(
        npu_inst_pe_1_1_3_n97) );
  NAND2_X1 npu_inst_pe_1_1_3_U85 ( .A1(npu_inst_pe_1_1_3_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_1_3_n60), .ZN(npu_inst_pe_1_1_3_n73) );
  OAI21_X1 npu_inst_pe_1_1_3_U84 ( .B1(npu_inst_pe_1_1_3_n61), .B2(
        npu_inst_pe_1_1_3_n60), .A(npu_inst_pe_1_1_3_n73), .ZN(
        npu_inst_pe_1_1_3_n96) );
  NAND2_X1 npu_inst_pe_1_1_3_U83 ( .A1(npu_inst_pe_1_1_3_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_1_3_n56), .ZN(npu_inst_pe_1_1_3_n72) );
  OAI21_X1 npu_inst_pe_1_1_3_U82 ( .B1(npu_inst_pe_1_1_3_n63), .B2(
        npu_inst_pe_1_1_3_n56), .A(npu_inst_pe_1_1_3_n72), .ZN(
        npu_inst_pe_1_1_3_n95) );
  NAND2_X1 npu_inst_pe_1_1_3_U81 ( .A1(npu_inst_pe_1_1_3_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_1_3_n56), .ZN(npu_inst_pe_1_1_3_n71) );
  OAI21_X1 npu_inst_pe_1_1_3_U80 ( .B1(npu_inst_pe_1_1_3_n61), .B2(
        npu_inst_pe_1_1_3_n56), .A(npu_inst_pe_1_1_3_n71), .ZN(
        npu_inst_pe_1_1_3_n94) );
  NAND2_X1 npu_inst_pe_1_1_3_U79 ( .A1(npu_inst_pe_1_1_3_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_1_3_n52), .ZN(npu_inst_pe_1_1_3_n70) );
  OAI21_X1 npu_inst_pe_1_1_3_U78 ( .B1(npu_inst_pe_1_1_3_n63), .B2(
        npu_inst_pe_1_1_3_n52), .A(npu_inst_pe_1_1_3_n70), .ZN(
        npu_inst_pe_1_1_3_n93) );
  NAND2_X1 npu_inst_pe_1_1_3_U77 ( .A1(npu_inst_pe_1_1_3_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_1_3_n52), .ZN(npu_inst_pe_1_1_3_n69) );
  OAI21_X1 npu_inst_pe_1_1_3_U76 ( .B1(npu_inst_pe_1_1_3_n61), .B2(
        npu_inst_pe_1_1_3_n52), .A(npu_inst_pe_1_1_3_n69), .ZN(
        npu_inst_pe_1_1_3_n92) );
  NAND2_X1 npu_inst_pe_1_1_3_U75 ( .A1(npu_inst_pe_1_1_3_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_1_3_n48), .ZN(npu_inst_pe_1_1_3_n68) );
  OAI21_X1 npu_inst_pe_1_1_3_U74 ( .B1(npu_inst_pe_1_1_3_n63), .B2(
        npu_inst_pe_1_1_3_n48), .A(npu_inst_pe_1_1_3_n68), .ZN(
        npu_inst_pe_1_1_3_n91) );
  NAND2_X1 npu_inst_pe_1_1_3_U73 ( .A1(npu_inst_pe_1_1_3_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_1_3_n48), .ZN(npu_inst_pe_1_1_3_n67) );
  OAI21_X1 npu_inst_pe_1_1_3_U72 ( .B1(npu_inst_pe_1_1_3_n61), .B2(
        npu_inst_pe_1_1_3_n48), .A(npu_inst_pe_1_1_3_n67), .ZN(
        npu_inst_pe_1_1_3_n90) );
  NAND2_X1 npu_inst_pe_1_1_3_U71 ( .A1(npu_inst_pe_1_1_3_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_1_3_n44), .ZN(npu_inst_pe_1_1_3_n66) );
  OAI21_X1 npu_inst_pe_1_1_3_U70 ( .B1(npu_inst_pe_1_1_3_n63), .B2(
        npu_inst_pe_1_1_3_n44), .A(npu_inst_pe_1_1_3_n66), .ZN(
        npu_inst_pe_1_1_3_n89) );
  NAND2_X1 npu_inst_pe_1_1_3_U69 ( .A1(npu_inst_pe_1_1_3_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_1_3_n44), .ZN(npu_inst_pe_1_1_3_n65) );
  OAI21_X1 npu_inst_pe_1_1_3_U68 ( .B1(npu_inst_pe_1_1_3_n61), .B2(
        npu_inst_pe_1_1_3_n44), .A(npu_inst_pe_1_1_3_n65), .ZN(
        npu_inst_pe_1_1_3_n88) );
  NAND2_X1 npu_inst_pe_1_1_3_U67 ( .A1(npu_inst_pe_1_1_3_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_1_3_n40), .ZN(npu_inst_pe_1_1_3_n64) );
  OAI21_X1 npu_inst_pe_1_1_3_U66 ( .B1(npu_inst_pe_1_1_3_n63), .B2(
        npu_inst_pe_1_1_3_n40), .A(npu_inst_pe_1_1_3_n64), .ZN(
        npu_inst_pe_1_1_3_n87) );
  NAND2_X1 npu_inst_pe_1_1_3_U65 ( .A1(npu_inst_pe_1_1_3_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_1_3_n40), .ZN(npu_inst_pe_1_1_3_n62) );
  OAI21_X1 npu_inst_pe_1_1_3_U64 ( .B1(npu_inst_pe_1_1_3_n61), .B2(
        npu_inst_pe_1_1_3_n40), .A(npu_inst_pe_1_1_3_n62), .ZN(
        npu_inst_pe_1_1_3_n86) );
  AND2_X1 npu_inst_pe_1_1_3_U63 ( .A1(npu_inst_pe_1_1_3_N93), .A2(npu_inst_n59), .ZN(npu_inst_int_data_y_1__3__0_) );
  AND2_X1 npu_inst_pe_1_1_3_U62 ( .A1(npu_inst_n59), .A2(npu_inst_pe_1_1_3_N94), .ZN(npu_inst_int_data_y_1__3__1_) );
  NOR3_X1 npu_inst_pe_1_1_3_U61 ( .A1(npu_inst_pe_1_1_3_n26), .A2(npu_inst_n59), .A3(npu_inst_int_ckg[52]), .ZN(npu_inst_pe_1_1_3_n85) );
  OR2_X1 npu_inst_pe_1_1_3_U60 ( .A1(npu_inst_pe_1_1_3_n85), .A2(
        npu_inst_pe_1_1_3_n2), .ZN(npu_inst_pe_1_1_3_N84) );
  AND2_X1 npu_inst_pe_1_1_3_U59 ( .A1(npu_inst_pe_1_1_3_int_q_acc_0_), .A2(
        npu_inst_pe_1_1_3_n1), .ZN(npu_inst_int_data_res_1__3__0_) );
  AND2_X1 npu_inst_pe_1_1_3_U58 ( .A1(npu_inst_pe_1_1_3_n2), .A2(
        npu_inst_pe_1_1_3_int_q_acc_7_), .ZN(npu_inst_int_data_res_1__3__7_)
         );
  AND2_X1 npu_inst_pe_1_1_3_U57 ( .A1(npu_inst_pe_1_1_3_int_q_acc_1_), .A2(
        npu_inst_pe_1_1_3_n1), .ZN(npu_inst_int_data_res_1__3__1_) );
  AND2_X1 npu_inst_pe_1_1_3_U56 ( .A1(npu_inst_pe_1_1_3_int_q_acc_2_), .A2(
        npu_inst_pe_1_1_3_n1), .ZN(npu_inst_int_data_res_1__3__2_) );
  AND2_X1 npu_inst_pe_1_1_3_U55 ( .A1(npu_inst_pe_1_1_3_int_q_acc_3_), .A2(
        npu_inst_pe_1_1_3_n2), .ZN(npu_inst_int_data_res_1__3__3_) );
  AND2_X1 npu_inst_pe_1_1_3_U54 ( .A1(npu_inst_pe_1_1_3_int_q_acc_4_), .A2(
        npu_inst_pe_1_1_3_n2), .ZN(npu_inst_int_data_res_1__3__4_) );
  AND2_X1 npu_inst_pe_1_1_3_U53 ( .A1(npu_inst_pe_1_1_3_int_q_acc_5_), .A2(
        npu_inst_pe_1_1_3_n2), .ZN(npu_inst_int_data_res_1__3__5_) );
  AND2_X1 npu_inst_pe_1_1_3_U52 ( .A1(npu_inst_pe_1_1_3_int_q_acc_6_), .A2(
        npu_inst_pe_1_1_3_n2), .ZN(npu_inst_int_data_res_1__3__6_) );
  AOI222_X1 npu_inst_pe_1_1_3_U51 ( .A1(npu_inst_int_data_res_2__3__0_), .A2(
        npu_inst_pe_1_1_3_n1), .B1(npu_inst_pe_1_1_3_N73), .B2(
        npu_inst_pe_1_1_3_n76), .C1(npu_inst_pe_1_1_3_N65), .C2(
        npu_inst_pe_1_1_3_n77), .ZN(npu_inst_pe_1_1_3_n84) );
  INV_X1 npu_inst_pe_1_1_3_U50 ( .A(npu_inst_pe_1_1_3_n84), .ZN(
        npu_inst_pe_1_1_3_n101) );
  AOI222_X1 npu_inst_pe_1_1_3_U49 ( .A1(npu_inst_int_data_res_2__3__7_), .A2(
        npu_inst_pe_1_1_3_n1), .B1(npu_inst_pe_1_1_3_N80), .B2(
        npu_inst_pe_1_1_3_n76), .C1(npu_inst_pe_1_1_3_N72), .C2(
        npu_inst_pe_1_1_3_n77), .ZN(npu_inst_pe_1_1_3_n75) );
  INV_X1 npu_inst_pe_1_1_3_U48 ( .A(npu_inst_pe_1_1_3_n75), .ZN(
        npu_inst_pe_1_1_3_n33) );
  AOI222_X1 npu_inst_pe_1_1_3_U47 ( .A1(npu_inst_int_data_res_2__3__1_), .A2(
        npu_inst_pe_1_1_3_n1), .B1(npu_inst_pe_1_1_3_N74), .B2(
        npu_inst_pe_1_1_3_n76), .C1(npu_inst_pe_1_1_3_N66), .C2(
        npu_inst_pe_1_1_3_n77), .ZN(npu_inst_pe_1_1_3_n83) );
  INV_X1 npu_inst_pe_1_1_3_U46 ( .A(npu_inst_pe_1_1_3_n83), .ZN(
        npu_inst_pe_1_1_3_n100) );
  AOI222_X1 npu_inst_pe_1_1_3_U45 ( .A1(npu_inst_int_data_res_2__3__2_), .A2(
        npu_inst_pe_1_1_3_n1), .B1(npu_inst_pe_1_1_3_N75), .B2(
        npu_inst_pe_1_1_3_n76), .C1(npu_inst_pe_1_1_3_N67), .C2(
        npu_inst_pe_1_1_3_n77), .ZN(npu_inst_pe_1_1_3_n82) );
  INV_X1 npu_inst_pe_1_1_3_U44 ( .A(npu_inst_pe_1_1_3_n82), .ZN(
        npu_inst_pe_1_1_3_n99) );
  AOI222_X1 npu_inst_pe_1_1_3_U43 ( .A1(npu_inst_int_data_res_2__3__3_), .A2(
        npu_inst_pe_1_1_3_n1), .B1(npu_inst_pe_1_1_3_N76), .B2(
        npu_inst_pe_1_1_3_n76), .C1(npu_inst_pe_1_1_3_N68), .C2(
        npu_inst_pe_1_1_3_n77), .ZN(npu_inst_pe_1_1_3_n81) );
  INV_X1 npu_inst_pe_1_1_3_U42 ( .A(npu_inst_pe_1_1_3_n81), .ZN(
        npu_inst_pe_1_1_3_n98) );
  AOI222_X1 npu_inst_pe_1_1_3_U41 ( .A1(npu_inst_int_data_res_2__3__4_), .A2(
        npu_inst_pe_1_1_3_n1), .B1(npu_inst_pe_1_1_3_N77), .B2(
        npu_inst_pe_1_1_3_n76), .C1(npu_inst_pe_1_1_3_N69), .C2(
        npu_inst_pe_1_1_3_n77), .ZN(npu_inst_pe_1_1_3_n80) );
  INV_X1 npu_inst_pe_1_1_3_U40 ( .A(npu_inst_pe_1_1_3_n80), .ZN(
        npu_inst_pe_1_1_3_n36) );
  AOI222_X1 npu_inst_pe_1_1_3_U39 ( .A1(npu_inst_int_data_res_2__3__5_), .A2(
        npu_inst_pe_1_1_3_n1), .B1(npu_inst_pe_1_1_3_N78), .B2(
        npu_inst_pe_1_1_3_n76), .C1(npu_inst_pe_1_1_3_N70), .C2(
        npu_inst_pe_1_1_3_n77), .ZN(npu_inst_pe_1_1_3_n79) );
  INV_X1 npu_inst_pe_1_1_3_U38 ( .A(npu_inst_pe_1_1_3_n79), .ZN(
        npu_inst_pe_1_1_3_n35) );
  AOI222_X1 npu_inst_pe_1_1_3_U37 ( .A1(npu_inst_int_data_res_2__3__6_), .A2(
        npu_inst_pe_1_1_3_n1), .B1(npu_inst_pe_1_1_3_N79), .B2(
        npu_inst_pe_1_1_3_n76), .C1(npu_inst_pe_1_1_3_N71), .C2(
        npu_inst_pe_1_1_3_n77), .ZN(npu_inst_pe_1_1_3_n78) );
  INV_X1 npu_inst_pe_1_1_3_U36 ( .A(npu_inst_pe_1_1_3_n78), .ZN(
        npu_inst_pe_1_1_3_n34) );
  INV_X1 npu_inst_pe_1_1_3_U35 ( .A(npu_inst_pe_1_1_3_int_data_1_), .ZN(
        npu_inst_pe_1_1_3_n14) );
  AND2_X1 npu_inst_pe_1_1_3_U34 ( .A1(npu_inst_int_data_x_1__3__1_), .A2(
        npu_inst_pe_1_1_3_int_q_weight_1_), .ZN(npu_inst_pe_1_1_3_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_1_3_U33 ( .A1(npu_inst_int_data_x_1__3__0_), .A2(
        npu_inst_pe_1_1_3_int_q_weight_1_), .ZN(npu_inst_pe_1_1_3_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_1_3_U32 ( .A1(npu_inst_n59), .A2(
        npu_inst_int_data_y_2__3__1_), .B1(npu_inst_pe_1_1_3_n3), .B2(
        npu_inst_int_data_x_1__4__1_), .ZN(npu_inst_pe_1_1_3_n63) );
  AOI22_X1 npu_inst_pe_1_1_3_U31 ( .A1(npu_inst_n59), .A2(
        npu_inst_int_data_y_2__3__0_), .B1(npu_inst_pe_1_1_3_n3), .B2(
        npu_inst_int_data_x_1__4__0_), .ZN(npu_inst_pe_1_1_3_n61) );
  INV_X1 npu_inst_pe_1_1_3_U30 ( .A(npu_inst_pe_1_1_3_int_data_0_), .ZN(
        npu_inst_pe_1_1_3_n13) );
  INV_X1 npu_inst_pe_1_1_3_U29 ( .A(npu_inst_n71), .ZN(npu_inst_pe_1_1_3_n5)
         );
  OR3_X1 npu_inst_pe_1_1_3_U28 ( .A1(npu_inst_pe_1_1_3_n6), .A2(
        npu_inst_pe_1_1_3_n8), .A3(npu_inst_pe_1_1_3_n5), .ZN(
        npu_inst_pe_1_1_3_n56) );
  OR3_X1 npu_inst_pe_1_1_3_U27 ( .A1(npu_inst_pe_1_1_3_n5), .A2(
        npu_inst_pe_1_1_3_n8), .A3(npu_inst_pe_1_1_3_n7), .ZN(
        npu_inst_pe_1_1_3_n48) );
  INV_X1 npu_inst_pe_1_1_3_U26 ( .A(npu_inst_pe_1_1_3_n5), .ZN(
        npu_inst_pe_1_1_3_n4) );
  INV_X1 npu_inst_pe_1_1_3_U25 ( .A(npu_inst_n126), .ZN(npu_inst_pe_1_1_3_n12)
         );
  OR3_X1 npu_inst_pe_1_1_3_U24 ( .A1(npu_inst_pe_1_1_3_n4), .A2(
        npu_inst_pe_1_1_3_n8), .A3(npu_inst_pe_1_1_3_n7), .ZN(
        npu_inst_pe_1_1_3_n52) );
  OR3_X1 npu_inst_pe_1_1_3_U23 ( .A1(npu_inst_pe_1_1_3_n6), .A2(
        npu_inst_pe_1_1_3_n8), .A3(npu_inst_pe_1_1_3_n4), .ZN(
        npu_inst_pe_1_1_3_n60) );
  NOR2_X1 npu_inst_pe_1_1_3_U22 ( .A1(npu_inst_pe_1_1_3_n60), .A2(
        npu_inst_pe_1_1_3_n3), .ZN(npu_inst_pe_1_1_3_n58) );
  NOR2_X1 npu_inst_pe_1_1_3_U21 ( .A1(npu_inst_pe_1_1_3_n56), .A2(
        npu_inst_pe_1_1_3_n3), .ZN(npu_inst_pe_1_1_3_n54) );
  NOR2_X1 npu_inst_pe_1_1_3_U20 ( .A1(npu_inst_pe_1_1_3_n52), .A2(
        npu_inst_pe_1_1_3_n3), .ZN(npu_inst_pe_1_1_3_n50) );
  NOR2_X1 npu_inst_pe_1_1_3_U19 ( .A1(npu_inst_pe_1_1_3_n48), .A2(
        npu_inst_pe_1_1_3_n3), .ZN(npu_inst_pe_1_1_3_n46) );
  NOR2_X1 npu_inst_pe_1_1_3_U18 ( .A1(npu_inst_pe_1_1_3_n40), .A2(
        npu_inst_pe_1_1_3_n3), .ZN(npu_inst_pe_1_1_3_n38) );
  NOR2_X1 npu_inst_pe_1_1_3_U17 ( .A1(npu_inst_pe_1_1_3_n44), .A2(
        npu_inst_pe_1_1_3_n3), .ZN(npu_inst_pe_1_1_3_n42) );
  BUF_X1 npu_inst_pe_1_1_3_U16 ( .A(npu_inst_n105), .Z(npu_inst_pe_1_1_3_n8)
         );
  BUF_X1 npu_inst_pe_1_1_3_U15 ( .A(npu_inst_pe_1_1_3_n12), .Z(
        npu_inst_pe_1_1_3_n11) );
  BUF_X1 npu_inst_pe_1_1_3_U14 ( .A(npu_inst_pe_1_1_3_n12), .Z(
        npu_inst_pe_1_1_3_n10) );
  BUF_X1 npu_inst_pe_1_1_3_U13 ( .A(npu_inst_pe_1_1_3_n12), .Z(
        npu_inst_pe_1_1_3_n9) );
  INV_X1 npu_inst_pe_1_1_3_U12 ( .A(npu_inst_pe_1_1_3_n38), .ZN(
        npu_inst_pe_1_1_3_n118) );
  INV_X1 npu_inst_pe_1_1_3_U11 ( .A(npu_inst_pe_1_1_3_n58), .ZN(
        npu_inst_pe_1_1_3_n114) );
  INV_X1 npu_inst_pe_1_1_3_U10 ( .A(npu_inst_pe_1_1_3_n54), .ZN(
        npu_inst_pe_1_1_3_n115) );
  INV_X1 npu_inst_pe_1_1_3_U9 ( .A(npu_inst_pe_1_1_3_n50), .ZN(
        npu_inst_pe_1_1_3_n116) );
  INV_X1 npu_inst_pe_1_1_3_U8 ( .A(npu_inst_pe_1_1_3_n46), .ZN(
        npu_inst_pe_1_1_3_n117) );
  INV_X1 npu_inst_pe_1_1_3_U7 ( .A(npu_inst_pe_1_1_3_n42), .ZN(
        npu_inst_pe_1_1_3_n119) );
  BUF_X1 npu_inst_pe_1_1_3_U6 ( .A(npu_inst_n33), .Z(npu_inst_pe_1_1_3_n2) );
  BUF_X1 npu_inst_pe_1_1_3_U5 ( .A(npu_inst_n33), .Z(npu_inst_pe_1_1_3_n1) );
  NOR2_X1 npu_inst_pe_1_1_3_U4 ( .A1(npu_inst_pe_1_1_3_int_q_weight_0_), .A2(
        npu_inst_pe_1_1_3_n1), .ZN(npu_inst_pe_1_1_3_n76) );
  NOR2_X1 npu_inst_pe_1_1_3_U3 ( .A1(npu_inst_pe_1_1_3_n27), .A2(
        npu_inst_pe_1_1_3_n1), .ZN(npu_inst_pe_1_1_3_n77) );
  FA_X1 npu_inst_pe_1_1_3_sub_77_U2_1 ( .A(npu_inst_pe_1_1_3_int_q_acc_1_), 
        .B(npu_inst_pe_1_1_3_n14), .CI(npu_inst_pe_1_1_3_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_1_3_sub_77_carry_2_), .S(npu_inst_pe_1_1_3_N66) );
  FA_X1 npu_inst_pe_1_1_3_add_79_U1_1 ( .A(npu_inst_pe_1_1_3_int_q_acc_1_), 
        .B(npu_inst_pe_1_1_3_int_data_1_), .CI(
        npu_inst_pe_1_1_3_add_79_carry_1_), .CO(
        npu_inst_pe_1_1_3_add_79_carry_2_), .S(npu_inst_pe_1_1_3_N74) );
  NAND3_X1 npu_inst_pe_1_1_3_U109 ( .A1(npu_inst_pe_1_1_3_n5), .A2(
        npu_inst_pe_1_1_3_n7), .A3(npu_inst_pe_1_1_3_n8), .ZN(
        npu_inst_pe_1_1_3_n44) );
  NAND3_X1 npu_inst_pe_1_1_3_U108 ( .A1(npu_inst_pe_1_1_3_n4), .A2(
        npu_inst_pe_1_1_3_n7), .A3(npu_inst_pe_1_1_3_n8), .ZN(
        npu_inst_pe_1_1_3_n40) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_1_3_n34), .CK(
        npu_inst_pe_1_1_3_net4040), .RN(npu_inst_pe_1_1_3_n9), .Q(
        npu_inst_pe_1_1_3_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_1_3_n35), .CK(
        npu_inst_pe_1_1_3_net4040), .RN(npu_inst_pe_1_1_3_n9), .Q(
        npu_inst_pe_1_1_3_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_1_3_n36), .CK(
        npu_inst_pe_1_1_3_net4040), .RN(npu_inst_pe_1_1_3_n9), .Q(
        npu_inst_pe_1_1_3_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_1_3_n98), .CK(
        npu_inst_pe_1_1_3_net4040), .RN(npu_inst_pe_1_1_3_n9), .Q(
        npu_inst_pe_1_1_3_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_1_3_n99), .CK(
        npu_inst_pe_1_1_3_net4040), .RN(npu_inst_pe_1_1_3_n9), .Q(
        npu_inst_pe_1_1_3_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_1_3_n100), 
        .CK(npu_inst_pe_1_1_3_net4040), .RN(npu_inst_pe_1_1_3_n9), .Q(
        npu_inst_pe_1_1_3_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_1_3_n33), .CK(
        npu_inst_pe_1_1_3_net4040), .RN(npu_inst_pe_1_1_3_n9), .Q(
        npu_inst_pe_1_1_3_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_1_3_n101), 
        .CK(npu_inst_pe_1_1_3_net4040), .RN(npu_inst_pe_1_1_3_n9), .Q(
        npu_inst_pe_1_1_3_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_weight_reg_0_ ( .D(npu_inst_n112), .CK(
        npu_inst_pe_1_1_3_net4046), .RN(npu_inst_pe_1_1_3_n9), .Q(
        npu_inst_pe_1_1_3_int_q_weight_0_), .QN(npu_inst_pe_1_1_3_n27) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_weight_reg_1_ ( .D(npu_inst_n118), .CK(
        npu_inst_pe_1_1_3_net4046), .RN(npu_inst_pe_1_1_3_n9), .Q(
        npu_inst_pe_1_1_3_int_q_weight_1_), .QN(npu_inst_pe_1_1_3_n26) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_1_3_n113), 
        .CK(npu_inst_pe_1_1_3_net4046), .RN(npu_inst_pe_1_1_3_n9), .Q(
        npu_inst_pe_1_1_3_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_1_3_n107), 
        .CK(npu_inst_pe_1_1_3_net4046), .RN(npu_inst_pe_1_1_3_n9), .Q(
        npu_inst_pe_1_1_3_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_1_3_n112), 
        .CK(npu_inst_pe_1_1_3_net4046), .RN(npu_inst_pe_1_1_3_n10), .Q(
        npu_inst_pe_1_1_3_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_1_3_n106), 
        .CK(npu_inst_pe_1_1_3_net4046), .RN(npu_inst_pe_1_1_3_n10), .Q(
        npu_inst_pe_1_1_3_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_1_3_n111), 
        .CK(npu_inst_pe_1_1_3_net4046), .RN(npu_inst_pe_1_1_3_n10), .Q(
        npu_inst_pe_1_1_3_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_1_3_n105), 
        .CK(npu_inst_pe_1_1_3_net4046), .RN(npu_inst_pe_1_1_3_n10), .Q(
        npu_inst_pe_1_1_3_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_1_3_n110), 
        .CK(npu_inst_pe_1_1_3_net4046), .RN(npu_inst_pe_1_1_3_n10), .Q(
        npu_inst_pe_1_1_3_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_1_3_n104), 
        .CK(npu_inst_pe_1_1_3_net4046), .RN(npu_inst_pe_1_1_3_n10), .Q(
        npu_inst_pe_1_1_3_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_1_3_n109), 
        .CK(npu_inst_pe_1_1_3_net4046), .RN(npu_inst_pe_1_1_3_n10), .Q(
        npu_inst_pe_1_1_3_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_1_3_n103), 
        .CK(npu_inst_pe_1_1_3_net4046), .RN(npu_inst_pe_1_1_3_n10), .Q(
        npu_inst_pe_1_1_3_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_1_3_n108), 
        .CK(npu_inst_pe_1_1_3_net4046), .RN(npu_inst_pe_1_1_3_n10), .Q(
        npu_inst_pe_1_1_3_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_1_3_n102), 
        .CK(npu_inst_pe_1_1_3_net4046), .RN(npu_inst_pe_1_1_3_n10), .Q(
        npu_inst_pe_1_1_3_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_1_3_n86), 
        .CK(npu_inst_pe_1_1_3_net4046), .RN(npu_inst_pe_1_1_3_n10), .Q(
        npu_inst_pe_1_1_3_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_1_3_n87), 
        .CK(npu_inst_pe_1_1_3_net4046), .RN(npu_inst_pe_1_1_3_n10), .Q(
        npu_inst_pe_1_1_3_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_1_3_n88), 
        .CK(npu_inst_pe_1_1_3_net4046), .RN(npu_inst_pe_1_1_3_n11), .Q(
        npu_inst_pe_1_1_3_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_1_3_n89), 
        .CK(npu_inst_pe_1_1_3_net4046), .RN(npu_inst_pe_1_1_3_n11), .Q(
        npu_inst_pe_1_1_3_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_1_3_n90), 
        .CK(npu_inst_pe_1_1_3_net4046), .RN(npu_inst_pe_1_1_3_n11), .Q(
        npu_inst_pe_1_1_3_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_1_3_n91), 
        .CK(npu_inst_pe_1_1_3_net4046), .RN(npu_inst_pe_1_1_3_n11), .Q(
        npu_inst_pe_1_1_3_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_1_3_n92), 
        .CK(npu_inst_pe_1_1_3_net4046), .RN(npu_inst_pe_1_1_3_n11), .Q(
        npu_inst_pe_1_1_3_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_1_3_n93), 
        .CK(npu_inst_pe_1_1_3_net4046), .RN(npu_inst_pe_1_1_3_n11), .Q(
        npu_inst_pe_1_1_3_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_1_3_n94), 
        .CK(npu_inst_pe_1_1_3_net4046), .RN(npu_inst_pe_1_1_3_n11), .Q(
        npu_inst_pe_1_1_3_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_1_3_n95), 
        .CK(npu_inst_pe_1_1_3_net4046), .RN(npu_inst_pe_1_1_3_n11), .Q(
        npu_inst_pe_1_1_3_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_1_3_n96), 
        .CK(npu_inst_pe_1_1_3_net4046), .RN(npu_inst_pe_1_1_3_n11), .Q(
        npu_inst_pe_1_1_3_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_1_3_n97), 
        .CK(npu_inst_pe_1_1_3_net4046), .RN(npu_inst_pe_1_1_3_n11), .Q(
        npu_inst_pe_1_1_3_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_1_3_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_1_3_N84), .SE(1'b0), .GCK(npu_inst_pe_1_1_3_net4040) );
  CLKGATETST_X1 npu_inst_pe_1_1_3_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n65), .SE(1'b0), .GCK(npu_inst_pe_1_1_3_net4046) );
  MUX2_X1 npu_inst_pe_1_1_4_U162 ( .A(npu_inst_pe_1_1_4_n32), .B(
        npu_inst_pe_1_1_4_n29), .S(npu_inst_pe_1_1_4_n8), .Z(
        npu_inst_pe_1_1_4_N93) );
  MUX2_X1 npu_inst_pe_1_1_4_U161 ( .A(npu_inst_pe_1_1_4_n31), .B(
        npu_inst_pe_1_1_4_n30), .S(npu_inst_pe_1_1_4_n6), .Z(
        npu_inst_pe_1_1_4_n32) );
  MUX2_X1 npu_inst_pe_1_1_4_U160 ( .A(npu_inst_pe_1_1_4_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_1_4_int_q_reg_v_1__0_), .S(npu_inst_pe_1_1_4_n4), .Z(
        npu_inst_pe_1_1_4_n31) );
  MUX2_X1 npu_inst_pe_1_1_4_U159 ( .A(npu_inst_pe_1_1_4_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_1_4_int_q_reg_v_3__0_), .S(npu_inst_pe_1_1_4_n4), .Z(
        npu_inst_pe_1_1_4_n30) );
  MUX2_X1 npu_inst_pe_1_1_4_U158 ( .A(npu_inst_pe_1_1_4_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_1_4_int_q_reg_v_5__0_), .S(npu_inst_pe_1_1_4_n4), .Z(
        npu_inst_pe_1_1_4_n29) );
  MUX2_X1 npu_inst_pe_1_1_4_U157 ( .A(npu_inst_pe_1_1_4_n28), .B(
        npu_inst_pe_1_1_4_n23), .S(npu_inst_pe_1_1_4_n8), .Z(
        npu_inst_pe_1_1_4_N94) );
  MUX2_X1 npu_inst_pe_1_1_4_U156 ( .A(npu_inst_pe_1_1_4_n25), .B(
        npu_inst_pe_1_1_4_n24), .S(npu_inst_pe_1_1_4_n6), .Z(
        npu_inst_pe_1_1_4_n28) );
  MUX2_X1 npu_inst_pe_1_1_4_U155 ( .A(npu_inst_pe_1_1_4_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_1_4_int_q_reg_v_1__1_), .S(npu_inst_pe_1_1_4_n4), .Z(
        npu_inst_pe_1_1_4_n25) );
  MUX2_X1 npu_inst_pe_1_1_4_U154 ( .A(npu_inst_pe_1_1_4_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_1_4_int_q_reg_v_3__1_), .S(npu_inst_pe_1_1_4_n4), .Z(
        npu_inst_pe_1_1_4_n24) );
  MUX2_X1 npu_inst_pe_1_1_4_U153 ( .A(npu_inst_pe_1_1_4_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_1_4_int_q_reg_v_5__1_), .S(npu_inst_pe_1_1_4_n4), .Z(
        npu_inst_pe_1_1_4_n23) );
  MUX2_X1 npu_inst_pe_1_1_4_U152 ( .A(npu_inst_pe_1_1_4_n22), .B(
        npu_inst_pe_1_1_4_n19), .S(npu_inst_pe_1_1_4_n8), .Z(
        npu_inst_int_data_x_1__4__1_) );
  MUX2_X1 npu_inst_pe_1_1_4_U151 ( .A(npu_inst_pe_1_1_4_n21), .B(
        npu_inst_pe_1_1_4_n20), .S(npu_inst_pe_1_1_4_n6), .Z(
        npu_inst_pe_1_1_4_n22) );
  MUX2_X1 npu_inst_pe_1_1_4_U150 ( .A(npu_inst_pe_1_1_4_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_1_4_int_q_reg_h_1__1_), .S(npu_inst_pe_1_1_4_n4), .Z(
        npu_inst_pe_1_1_4_n21) );
  MUX2_X1 npu_inst_pe_1_1_4_U149 ( .A(npu_inst_pe_1_1_4_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_1_4_int_q_reg_h_3__1_), .S(npu_inst_pe_1_1_4_n4), .Z(
        npu_inst_pe_1_1_4_n20) );
  MUX2_X1 npu_inst_pe_1_1_4_U148 ( .A(npu_inst_pe_1_1_4_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_1_4_int_q_reg_h_5__1_), .S(npu_inst_pe_1_1_4_n4), .Z(
        npu_inst_pe_1_1_4_n19) );
  MUX2_X1 npu_inst_pe_1_1_4_U147 ( .A(npu_inst_pe_1_1_4_n18), .B(
        npu_inst_pe_1_1_4_n15), .S(npu_inst_pe_1_1_4_n8), .Z(
        npu_inst_int_data_x_1__4__0_) );
  MUX2_X1 npu_inst_pe_1_1_4_U146 ( .A(npu_inst_pe_1_1_4_n17), .B(
        npu_inst_pe_1_1_4_n16), .S(npu_inst_pe_1_1_4_n6), .Z(
        npu_inst_pe_1_1_4_n18) );
  MUX2_X1 npu_inst_pe_1_1_4_U145 ( .A(npu_inst_pe_1_1_4_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_1_4_int_q_reg_h_1__0_), .S(npu_inst_pe_1_1_4_n4), .Z(
        npu_inst_pe_1_1_4_n17) );
  MUX2_X1 npu_inst_pe_1_1_4_U144 ( .A(npu_inst_pe_1_1_4_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_1_4_int_q_reg_h_3__0_), .S(npu_inst_pe_1_1_4_n4), .Z(
        npu_inst_pe_1_1_4_n16) );
  MUX2_X1 npu_inst_pe_1_1_4_U143 ( .A(npu_inst_pe_1_1_4_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_1_4_int_q_reg_h_5__0_), .S(npu_inst_pe_1_1_4_n4), .Z(
        npu_inst_pe_1_1_4_n15) );
  XOR2_X1 npu_inst_pe_1_1_4_U142 ( .A(npu_inst_pe_1_1_4_int_data_0_), .B(
        npu_inst_pe_1_1_4_int_q_acc_0_), .Z(npu_inst_pe_1_1_4_N73) );
  AND2_X1 npu_inst_pe_1_1_4_U141 ( .A1(npu_inst_pe_1_1_4_int_q_acc_0_), .A2(
        npu_inst_pe_1_1_4_int_data_0_), .ZN(npu_inst_pe_1_1_4_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_1_4_U140 ( .A(npu_inst_pe_1_1_4_int_q_acc_0_), .B(
        npu_inst_pe_1_1_4_n13), .ZN(npu_inst_pe_1_1_4_N65) );
  OR2_X1 npu_inst_pe_1_1_4_U139 ( .A1(npu_inst_pe_1_1_4_n13), .A2(
        npu_inst_pe_1_1_4_int_q_acc_0_), .ZN(npu_inst_pe_1_1_4_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_1_4_U138 ( .A(npu_inst_pe_1_1_4_int_q_acc_2_), .B(
        npu_inst_pe_1_1_4_add_79_carry_2_), .Z(npu_inst_pe_1_1_4_N75) );
  AND2_X1 npu_inst_pe_1_1_4_U137 ( .A1(npu_inst_pe_1_1_4_add_79_carry_2_), 
        .A2(npu_inst_pe_1_1_4_int_q_acc_2_), .ZN(
        npu_inst_pe_1_1_4_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_1_4_U136 ( .A(npu_inst_pe_1_1_4_int_q_acc_3_), .B(
        npu_inst_pe_1_1_4_add_79_carry_3_), .Z(npu_inst_pe_1_1_4_N76) );
  AND2_X1 npu_inst_pe_1_1_4_U135 ( .A1(npu_inst_pe_1_1_4_add_79_carry_3_), 
        .A2(npu_inst_pe_1_1_4_int_q_acc_3_), .ZN(
        npu_inst_pe_1_1_4_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_1_4_U134 ( .A(npu_inst_pe_1_1_4_int_q_acc_4_), .B(
        npu_inst_pe_1_1_4_add_79_carry_4_), .Z(npu_inst_pe_1_1_4_N77) );
  AND2_X1 npu_inst_pe_1_1_4_U133 ( .A1(npu_inst_pe_1_1_4_add_79_carry_4_), 
        .A2(npu_inst_pe_1_1_4_int_q_acc_4_), .ZN(
        npu_inst_pe_1_1_4_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_1_4_U132 ( .A(npu_inst_pe_1_1_4_int_q_acc_5_), .B(
        npu_inst_pe_1_1_4_add_79_carry_5_), .Z(npu_inst_pe_1_1_4_N78) );
  AND2_X1 npu_inst_pe_1_1_4_U131 ( .A1(npu_inst_pe_1_1_4_add_79_carry_5_), 
        .A2(npu_inst_pe_1_1_4_int_q_acc_5_), .ZN(
        npu_inst_pe_1_1_4_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_1_4_U130 ( .A(npu_inst_pe_1_1_4_int_q_acc_6_), .B(
        npu_inst_pe_1_1_4_add_79_carry_6_), .Z(npu_inst_pe_1_1_4_N79) );
  AND2_X1 npu_inst_pe_1_1_4_U129 ( .A1(npu_inst_pe_1_1_4_add_79_carry_6_), 
        .A2(npu_inst_pe_1_1_4_int_q_acc_6_), .ZN(
        npu_inst_pe_1_1_4_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_1_4_U128 ( .A(npu_inst_pe_1_1_4_int_q_acc_7_), .B(
        npu_inst_pe_1_1_4_add_79_carry_7_), .Z(npu_inst_pe_1_1_4_N80) );
  XNOR2_X1 npu_inst_pe_1_1_4_U127 ( .A(npu_inst_pe_1_1_4_sub_77_carry_2_), .B(
        npu_inst_pe_1_1_4_int_q_acc_2_), .ZN(npu_inst_pe_1_1_4_N67) );
  OR2_X1 npu_inst_pe_1_1_4_U126 ( .A1(npu_inst_pe_1_1_4_int_q_acc_2_), .A2(
        npu_inst_pe_1_1_4_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_1_4_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_1_4_U125 ( .A(npu_inst_pe_1_1_4_sub_77_carry_3_), .B(
        npu_inst_pe_1_1_4_int_q_acc_3_), .ZN(npu_inst_pe_1_1_4_N68) );
  OR2_X1 npu_inst_pe_1_1_4_U124 ( .A1(npu_inst_pe_1_1_4_int_q_acc_3_), .A2(
        npu_inst_pe_1_1_4_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_1_4_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_1_4_U123 ( .A(npu_inst_pe_1_1_4_sub_77_carry_4_), .B(
        npu_inst_pe_1_1_4_int_q_acc_4_), .ZN(npu_inst_pe_1_1_4_N69) );
  OR2_X1 npu_inst_pe_1_1_4_U122 ( .A1(npu_inst_pe_1_1_4_int_q_acc_4_), .A2(
        npu_inst_pe_1_1_4_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_1_4_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_1_4_U121 ( .A(npu_inst_pe_1_1_4_sub_77_carry_5_), .B(
        npu_inst_pe_1_1_4_int_q_acc_5_), .ZN(npu_inst_pe_1_1_4_N70) );
  OR2_X1 npu_inst_pe_1_1_4_U120 ( .A1(npu_inst_pe_1_1_4_int_q_acc_5_), .A2(
        npu_inst_pe_1_1_4_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_1_4_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_1_4_U119 ( .A(npu_inst_pe_1_1_4_sub_77_carry_6_), .B(
        npu_inst_pe_1_1_4_int_q_acc_6_), .ZN(npu_inst_pe_1_1_4_N71) );
  OR2_X1 npu_inst_pe_1_1_4_U118 ( .A1(npu_inst_pe_1_1_4_int_q_acc_6_), .A2(
        npu_inst_pe_1_1_4_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_1_4_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_1_4_U117 ( .A(npu_inst_pe_1_1_4_int_q_acc_7_), .B(
        npu_inst_pe_1_1_4_sub_77_carry_7_), .ZN(npu_inst_pe_1_1_4_N72) );
  INV_X1 npu_inst_pe_1_1_4_U116 ( .A(npu_inst_n79), .ZN(npu_inst_pe_1_1_4_n7)
         );
  INV_X1 npu_inst_pe_1_1_4_U115 ( .A(npu_inst_pe_1_1_4_n7), .ZN(
        npu_inst_pe_1_1_4_n6) );
  INV_X1 npu_inst_pe_1_1_4_U114 ( .A(npu_inst_n59), .ZN(npu_inst_pe_1_1_4_n3)
         );
  AOI22_X1 npu_inst_pe_1_1_4_U113 ( .A1(npu_inst_int_data_y_2__4__0_), .A2(
        npu_inst_pe_1_1_4_n58), .B1(npu_inst_pe_1_1_4_n114), .B2(
        npu_inst_pe_1_1_4_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_1_4_n57) );
  INV_X1 npu_inst_pe_1_1_4_U112 ( .A(npu_inst_pe_1_1_4_n57), .ZN(
        npu_inst_pe_1_1_4_n108) );
  AOI22_X1 npu_inst_pe_1_1_4_U111 ( .A1(npu_inst_int_data_y_2__4__0_), .A2(
        npu_inst_pe_1_1_4_n54), .B1(npu_inst_pe_1_1_4_n115), .B2(
        npu_inst_pe_1_1_4_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_1_4_n53) );
  INV_X1 npu_inst_pe_1_1_4_U110 ( .A(npu_inst_pe_1_1_4_n53), .ZN(
        npu_inst_pe_1_1_4_n109) );
  AOI22_X1 npu_inst_pe_1_1_4_U107 ( .A1(npu_inst_int_data_y_2__4__0_), .A2(
        npu_inst_pe_1_1_4_n50), .B1(npu_inst_pe_1_1_4_n116), .B2(
        npu_inst_pe_1_1_4_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_1_4_n49) );
  INV_X1 npu_inst_pe_1_1_4_U106 ( .A(npu_inst_pe_1_1_4_n49), .ZN(
        npu_inst_pe_1_1_4_n110) );
  AOI22_X1 npu_inst_pe_1_1_4_U105 ( .A1(npu_inst_int_data_y_2__4__0_), .A2(
        npu_inst_pe_1_1_4_n46), .B1(npu_inst_pe_1_1_4_n117), .B2(
        npu_inst_pe_1_1_4_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_1_4_n45) );
  INV_X1 npu_inst_pe_1_1_4_U104 ( .A(npu_inst_pe_1_1_4_n45), .ZN(
        npu_inst_pe_1_1_4_n111) );
  AOI22_X1 npu_inst_pe_1_1_4_U103 ( .A1(npu_inst_int_data_y_2__4__0_), .A2(
        npu_inst_pe_1_1_4_n42), .B1(npu_inst_pe_1_1_4_n119), .B2(
        npu_inst_pe_1_1_4_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_1_4_n41) );
  INV_X1 npu_inst_pe_1_1_4_U102 ( .A(npu_inst_pe_1_1_4_n41), .ZN(
        npu_inst_pe_1_1_4_n112) );
  AOI22_X1 npu_inst_pe_1_1_4_U101 ( .A1(npu_inst_int_data_y_2__4__1_), .A2(
        npu_inst_pe_1_1_4_n58), .B1(npu_inst_pe_1_1_4_n114), .B2(
        npu_inst_pe_1_1_4_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_1_4_n59) );
  INV_X1 npu_inst_pe_1_1_4_U100 ( .A(npu_inst_pe_1_1_4_n59), .ZN(
        npu_inst_pe_1_1_4_n102) );
  AOI22_X1 npu_inst_pe_1_1_4_U99 ( .A1(npu_inst_int_data_y_2__4__1_), .A2(
        npu_inst_pe_1_1_4_n54), .B1(npu_inst_pe_1_1_4_n115), .B2(
        npu_inst_pe_1_1_4_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_1_4_n55) );
  INV_X1 npu_inst_pe_1_1_4_U98 ( .A(npu_inst_pe_1_1_4_n55), .ZN(
        npu_inst_pe_1_1_4_n103) );
  AOI22_X1 npu_inst_pe_1_1_4_U97 ( .A1(npu_inst_int_data_y_2__4__1_), .A2(
        npu_inst_pe_1_1_4_n50), .B1(npu_inst_pe_1_1_4_n116), .B2(
        npu_inst_pe_1_1_4_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_1_4_n51) );
  INV_X1 npu_inst_pe_1_1_4_U96 ( .A(npu_inst_pe_1_1_4_n51), .ZN(
        npu_inst_pe_1_1_4_n104) );
  AOI22_X1 npu_inst_pe_1_1_4_U95 ( .A1(npu_inst_int_data_y_2__4__1_), .A2(
        npu_inst_pe_1_1_4_n46), .B1(npu_inst_pe_1_1_4_n117), .B2(
        npu_inst_pe_1_1_4_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_1_4_n47) );
  INV_X1 npu_inst_pe_1_1_4_U94 ( .A(npu_inst_pe_1_1_4_n47), .ZN(
        npu_inst_pe_1_1_4_n105) );
  AOI22_X1 npu_inst_pe_1_1_4_U93 ( .A1(npu_inst_int_data_y_2__4__1_), .A2(
        npu_inst_pe_1_1_4_n42), .B1(npu_inst_pe_1_1_4_n119), .B2(
        npu_inst_pe_1_1_4_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_1_4_n43) );
  INV_X1 npu_inst_pe_1_1_4_U92 ( .A(npu_inst_pe_1_1_4_n43), .ZN(
        npu_inst_pe_1_1_4_n106) );
  AOI22_X1 npu_inst_pe_1_1_4_U91 ( .A1(npu_inst_pe_1_1_4_n38), .A2(
        npu_inst_int_data_y_2__4__1_), .B1(npu_inst_pe_1_1_4_n118), .B2(
        npu_inst_pe_1_1_4_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_1_4_n39) );
  INV_X1 npu_inst_pe_1_1_4_U90 ( .A(npu_inst_pe_1_1_4_n39), .ZN(
        npu_inst_pe_1_1_4_n107) );
  AOI22_X1 npu_inst_pe_1_1_4_U89 ( .A1(npu_inst_pe_1_1_4_n38), .A2(
        npu_inst_int_data_y_2__4__0_), .B1(npu_inst_pe_1_1_4_n118), .B2(
        npu_inst_pe_1_1_4_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_1_4_n37) );
  INV_X1 npu_inst_pe_1_1_4_U88 ( .A(npu_inst_pe_1_1_4_n37), .ZN(
        npu_inst_pe_1_1_4_n113) );
  NAND2_X1 npu_inst_pe_1_1_4_U87 ( .A1(npu_inst_pe_1_1_4_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_1_4_n60), .ZN(npu_inst_pe_1_1_4_n74) );
  OAI21_X1 npu_inst_pe_1_1_4_U86 ( .B1(npu_inst_pe_1_1_4_n63), .B2(
        npu_inst_pe_1_1_4_n60), .A(npu_inst_pe_1_1_4_n74), .ZN(
        npu_inst_pe_1_1_4_n97) );
  NAND2_X1 npu_inst_pe_1_1_4_U85 ( .A1(npu_inst_pe_1_1_4_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_1_4_n60), .ZN(npu_inst_pe_1_1_4_n73) );
  OAI21_X1 npu_inst_pe_1_1_4_U84 ( .B1(npu_inst_pe_1_1_4_n61), .B2(
        npu_inst_pe_1_1_4_n60), .A(npu_inst_pe_1_1_4_n73), .ZN(
        npu_inst_pe_1_1_4_n96) );
  NAND2_X1 npu_inst_pe_1_1_4_U83 ( .A1(npu_inst_pe_1_1_4_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_1_4_n56), .ZN(npu_inst_pe_1_1_4_n72) );
  OAI21_X1 npu_inst_pe_1_1_4_U82 ( .B1(npu_inst_pe_1_1_4_n63), .B2(
        npu_inst_pe_1_1_4_n56), .A(npu_inst_pe_1_1_4_n72), .ZN(
        npu_inst_pe_1_1_4_n95) );
  NAND2_X1 npu_inst_pe_1_1_4_U81 ( .A1(npu_inst_pe_1_1_4_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_1_4_n56), .ZN(npu_inst_pe_1_1_4_n71) );
  OAI21_X1 npu_inst_pe_1_1_4_U80 ( .B1(npu_inst_pe_1_1_4_n61), .B2(
        npu_inst_pe_1_1_4_n56), .A(npu_inst_pe_1_1_4_n71), .ZN(
        npu_inst_pe_1_1_4_n94) );
  NAND2_X1 npu_inst_pe_1_1_4_U79 ( .A1(npu_inst_pe_1_1_4_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_1_4_n52), .ZN(npu_inst_pe_1_1_4_n70) );
  OAI21_X1 npu_inst_pe_1_1_4_U78 ( .B1(npu_inst_pe_1_1_4_n63), .B2(
        npu_inst_pe_1_1_4_n52), .A(npu_inst_pe_1_1_4_n70), .ZN(
        npu_inst_pe_1_1_4_n93) );
  NAND2_X1 npu_inst_pe_1_1_4_U77 ( .A1(npu_inst_pe_1_1_4_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_1_4_n52), .ZN(npu_inst_pe_1_1_4_n69) );
  OAI21_X1 npu_inst_pe_1_1_4_U76 ( .B1(npu_inst_pe_1_1_4_n61), .B2(
        npu_inst_pe_1_1_4_n52), .A(npu_inst_pe_1_1_4_n69), .ZN(
        npu_inst_pe_1_1_4_n92) );
  NAND2_X1 npu_inst_pe_1_1_4_U75 ( .A1(npu_inst_pe_1_1_4_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_1_4_n48), .ZN(npu_inst_pe_1_1_4_n68) );
  OAI21_X1 npu_inst_pe_1_1_4_U74 ( .B1(npu_inst_pe_1_1_4_n63), .B2(
        npu_inst_pe_1_1_4_n48), .A(npu_inst_pe_1_1_4_n68), .ZN(
        npu_inst_pe_1_1_4_n91) );
  NAND2_X1 npu_inst_pe_1_1_4_U73 ( .A1(npu_inst_pe_1_1_4_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_1_4_n48), .ZN(npu_inst_pe_1_1_4_n67) );
  OAI21_X1 npu_inst_pe_1_1_4_U72 ( .B1(npu_inst_pe_1_1_4_n61), .B2(
        npu_inst_pe_1_1_4_n48), .A(npu_inst_pe_1_1_4_n67), .ZN(
        npu_inst_pe_1_1_4_n90) );
  NAND2_X1 npu_inst_pe_1_1_4_U71 ( .A1(npu_inst_pe_1_1_4_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_1_4_n44), .ZN(npu_inst_pe_1_1_4_n66) );
  OAI21_X1 npu_inst_pe_1_1_4_U70 ( .B1(npu_inst_pe_1_1_4_n63), .B2(
        npu_inst_pe_1_1_4_n44), .A(npu_inst_pe_1_1_4_n66), .ZN(
        npu_inst_pe_1_1_4_n89) );
  NAND2_X1 npu_inst_pe_1_1_4_U69 ( .A1(npu_inst_pe_1_1_4_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_1_4_n44), .ZN(npu_inst_pe_1_1_4_n65) );
  OAI21_X1 npu_inst_pe_1_1_4_U68 ( .B1(npu_inst_pe_1_1_4_n61), .B2(
        npu_inst_pe_1_1_4_n44), .A(npu_inst_pe_1_1_4_n65), .ZN(
        npu_inst_pe_1_1_4_n88) );
  NAND2_X1 npu_inst_pe_1_1_4_U67 ( .A1(npu_inst_pe_1_1_4_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_1_4_n40), .ZN(npu_inst_pe_1_1_4_n64) );
  OAI21_X1 npu_inst_pe_1_1_4_U66 ( .B1(npu_inst_pe_1_1_4_n63), .B2(
        npu_inst_pe_1_1_4_n40), .A(npu_inst_pe_1_1_4_n64), .ZN(
        npu_inst_pe_1_1_4_n87) );
  NAND2_X1 npu_inst_pe_1_1_4_U65 ( .A1(npu_inst_pe_1_1_4_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_1_4_n40), .ZN(npu_inst_pe_1_1_4_n62) );
  OAI21_X1 npu_inst_pe_1_1_4_U64 ( .B1(npu_inst_pe_1_1_4_n61), .B2(
        npu_inst_pe_1_1_4_n40), .A(npu_inst_pe_1_1_4_n62), .ZN(
        npu_inst_pe_1_1_4_n86) );
  AND2_X1 npu_inst_pe_1_1_4_U63 ( .A1(npu_inst_pe_1_1_4_N93), .A2(npu_inst_n59), .ZN(npu_inst_int_data_y_1__4__0_) );
  AND2_X1 npu_inst_pe_1_1_4_U62 ( .A1(npu_inst_n59), .A2(npu_inst_pe_1_1_4_N94), .ZN(npu_inst_int_data_y_1__4__1_) );
  NOR3_X1 npu_inst_pe_1_1_4_U61 ( .A1(npu_inst_pe_1_1_4_n26), .A2(npu_inst_n59), .A3(npu_inst_int_ckg[51]), .ZN(npu_inst_pe_1_1_4_n85) );
  OR2_X1 npu_inst_pe_1_1_4_U60 ( .A1(npu_inst_pe_1_1_4_n85), .A2(
        npu_inst_pe_1_1_4_n2), .ZN(npu_inst_pe_1_1_4_N84) );
  AND2_X1 npu_inst_pe_1_1_4_U59 ( .A1(npu_inst_pe_1_1_4_int_q_acc_0_), .A2(
        npu_inst_pe_1_1_4_n1), .ZN(npu_inst_int_data_res_1__4__0_) );
  AND2_X1 npu_inst_pe_1_1_4_U58 ( .A1(npu_inst_pe_1_1_4_n2), .A2(
        npu_inst_pe_1_1_4_int_q_acc_7_), .ZN(npu_inst_int_data_res_1__4__7_)
         );
  AND2_X1 npu_inst_pe_1_1_4_U57 ( .A1(npu_inst_pe_1_1_4_int_q_acc_1_), .A2(
        npu_inst_pe_1_1_4_n1), .ZN(npu_inst_int_data_res_1__4__1_) );
  AND2_X1 npu_inst_pe_1_1_4_U56 ( .A1(npu_inst_pe_1_1_4_int_q_acc_2_), .A2(
        npu_inst_pe_1_1_4_n1), .ZN(npu_inst_int_data_res_1__4__2_) );
  AND2_X1 npu_inst_pe_1_1_4_U55 ( .A1(npu_inst_pe_1_1_4_int_q_acc_3_), .A2(
        npu_inst_pe_1_1_4_n2), .ZN(npu_inst_int_data_res_1__4__3_) );
  AND2_X1 npu_inst_pe_1_1_4_U54 ( .A1(npu_inst_pe_1_1_4_int_q_acc_4_), .A2(
        npu_inst_pe_1_1_4_n2), .ZN(npu_inst_int_data_res_1__4__4_) );
  AND2_X1 npu_inst_pe_1_1_4_U53 ( .A1(npu_inst_pe_1_1_4_int_q_acc_5_), .A2(
        npu_inst_pe_1_1_4_n2), .ZN(npu_inst_int_data_res_1__4__5_) );
  AND2_X1 npu_inst_pe_1_1_4_U52 ( .A1(npu_inst_pe_1_1_4_int_q_acc_6_), .A2(
        npu_inst_pe_1_1_4_n2), .ZN(npu_inst_int_data_res_1__4__6_) );
  AOI222_X1 npu_inst_pe_1_1_4_U51 ( .A1(npu_inst_int_data_res_2__4__0_), .A2(
        npu_inst_pe_1_1_4_n1), .B1(npu_inst_pe_1_1_4_N73), .B2(
        npu_inst_pe_1_1_4_n76), .C1(npu_inst_pe_1_1_4_N65), .C2(
        npu_inst_pe_1_1_4_n77), .ZN(npu_inst_pe_1_1_4_n84) );
  INV_X1 npu_inst_pe_1_1_4_U50 ( .A(npu_inst_pe_1_1_4_n84), .ZN(
        npu_inst_pe_1_1_4_n101) );
  AOI222_X1 npu_inst_pe_1_1_4_U49 ( .A1(npu_inst_int_data_res_2__4__7_), .A2(
        npu_inst_pe_1_1_4_n1), .B1(npu_inst_pe_1_1_4_N80), .B2(
        npu_inst_pe_1_1_4_n76), .C1(npu_inst_pe_1_1_4_N72), .C2(
        npu_inst_pe_1_1_4_n77), .ZN(npu_inst_pe_1_1_4_n75) );
  INV_X1 npu_inst_pe_1_1_4_U48 ( .A(npu_inst_pe_1_1_4_n75), .ZN(
        npu_inst_pe_1_1_4_n33) );
  AOI222_X1 npu_inst_pe_1_1_4_U47 ( .A1(npu_inst_int_data_res_2__4__1_), .A2(
        npu_inst_pe_1_1_4_n1), .B1(npu_inst_pe_1_1_4_N74), .B2(
        npu_inst_pe_1_1_4_n76), .C1(npu_inst_pe_1_1_4_N66), .C2(
        npu_inst_pe_1_1_4_n77), .ZN(npu_inst_pe_1_1_4_n83) );
  INV_X1 npu_inst_pe_1_1_4_U46 ( .A(npu_inst_pe_1_1_4_n83), .ZN(
        npu_inst_pe_1_1_4_n100) );
  AOI222_X1 npu_inst_pe_1_1_4_U45 ( .A1(npu_inst_int_data_res_2__4__2_), .A2(
        npu_inst_pe_1_1_4_n1), .B1(npu_inst_pe_1_1_4_N75), .B2(
        npu_inst_pe_1_1_4_n76), .C1(npu_inst_pe_1_1_4_N67), .C2(
        npu_inst_pe_1_1_4_n77), .ZN(npu_inst_pe_1_1_4_n82) );
  INV_X1 npu_inst_pe_1_1_4_U44 ( .A(npu_inst_pe_1_1_4_n82), .ZN(
        npu_inst_pe_1_1_4_n99) );
  AOI222_X1 npu_inst_pe_1_1_4_U43 ( .A1(npu_inst_int_data_res_2__4__3_), .A2(
        npu_inst_pe_1_1_4_n1), .B1(npu_inst_pe_1_1_4_N76), .B2(
        npu_inst_pe_1_1_4_n76), .C1(npu_inst_pe_1_1_4_N68), .C2(
        npu_inst_pe_1_1_4_n77), .ZN(npu_inst_pe_1_1_4_n81) );
  INV_X1 npu_inst_pe_1_1_4_U42 ( .A(npu_inst_pe_1_1_4_n81), .ZN(
        npu_inst_pe_1_1_4_n98) );
  AOI222_X1 npu_inst_pe_1_1_4_U41 ( .A1(npu_inst_int_data_res_2__4__4_), .A2(
        npu_inst_pe_1_1_4_n1), .B1(npu_inst_pe_1_1_4_N77), .B2(
        npu_inst_pe_1_1_4_n76), .C1(npu_inst_pe_1_1_4_N69), .C2(
        npu_inst_pe_1_1_4_n77), .ZN(npu_inst_pe_1_1_4_n80) );
  INV_X1 npu_inst_pe_1_1_4_U40 ( .A(npu_inst_pe_1_1_4_n80), .ZN(
        npu_inst_pe_1_1_4_n36) );
  AOI222_X1 npu_inst_pe_1_1_4_U39 ( .A1(npu_inst_int_data_res_2__4__5_), .A2(
        npu_inst_pe_1_1_4_n1), .B1(npu_inst_pe_1_1_4_N78), .B2(
        npu_inst_pe_1_1_4_n76), .C1(npu_inst_pe_1_1_4_N70), .C2(
        npu_inst_pe_1_1_4_n77), .ZN(npu_inst_pe_1_1_4_n79) );
  INV_X1 npu_inst_pe_1_1_4_U38 ( .A(npu_inst_pe_1_1_4_n79), .ZN(
        npu_inst_pe_1_1_4_n35) );
  AOI222_X1 npu_inst_pe_1_1_4_U37 ( .A1(npu_inst_int_data_res_2__4__6_), .A2(
        npu_inst_pe_1_1_4_n1), .B1(npu_inst_pe_1_1_4_N79), .B2(
        npu_inst_pe_1_1_4_n76), .C1(npu_inst_pe_1_1_4_N71), .C2(
        npu_inst_pe_1_1_4_n77), .ZN(npu_inst_pe_1_1_4_n78) );
  INV_X1 npu_inst_pe_1_1_4_U36 ( .A(npu_inst_pe_1_1_4_n78), .ZN(
        npu_inst_pe_1_1_4_n34) );
  INV_X1 npu_inst_pe_1_1_4_U35 ( .A(npu_inst_pe_1_1_4_int_data_1_), .ZN(
        npu_inst_pe_1_1_4_n14) );
  AND2_X1 npu_inst_pe_1_1_4_U34 ( .A1(npu_inst_int_data_x_1__4__1_), .A2(
        npu_inst_pe_1_1_4_int_q_weight_1_), .ZN(npu_inst_pe_1_1_4_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_1_4_U33 ( .A1(npu_inst_int_data_x_1__4__0_), .A2(
        npu_inst_pe_1_1_4_int_q_weight_1_), .ZN(npu_inst_pe_1_1_4_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_1_4_U32 ( .A1(npu_inst_n59), .A2(
        npu_inst_int_data_y_2__4__1_), .B1(npu_inst_pe_1_1_4_n3), .B2(
        npu_inst_int_data_x_1__5__1_), .ZN(npu_inst_pe_1_1_4_n63) );
  AOI22_X1 npu_inst_pe_1_1_4_U31 ( .A1(npu_inst_n59), .A2(
        npu_inst_int_data_y_2__4__0_), .B1(npu_inst_pe_1_1_4_n3), .B2(
        npu_inst_int_data_x_1__5__0_), .ZN(npu_inst_pe_1_1_4_n61) );
  INV_X1 npu_inst_pe_1_1_4_U30 ( .A(npu_inst_pe_1_1_4_int_data_0_), .ZN(
        npu_inst_pe_1_1_4_n13) );
  INV_X1 npu_inst_pe_1_1_4_U29 ( .A(npu_inst_n71), .ZN(npu_inst_pe_1_1_4_n5)
         );
  OR3_X1 npu_inst_pe_1_1_4_U28 ( .A1(npu_inst_pe_1_1_4_n6), .A2(
        npu_inst_pe_1_1_4_n8), .A3(npu_inst_pe_1_1_4_n5), .ZN(
        npu_inst_pe_1_1_4_n56) );
  OR3_X1 npu_inst_pe_1_1_4_U27 ( .A1(npu_inst_pe_1_1_4_n5), .A2(
        npu_inst_pe_1_1_4_n8), .A3(npu_inst_pe_1_1_4_n7), .ZN(
        npu_inst_pe_1_1_4_n48) );
  INV_X1 npu_inst_pe_1_1_4_U26 ( .A(npu_inst_pe_1_1_4_n5), .ZN(
        npu_inst_pe_1_1_4_n4) );
  INV_X1 npu_inst_pe_1_1_4_U25 ( .A(npu_inst_n126), .ZN(npu_inst_pe_1_1_4_n12)
         );
  OR3_X1 npu_inst_pe_1_1_4_U24 ( .A1(npu_inst_pe_1_1_4_n4), .A2(
        npu_inst_pe_1_1_4_n8), .A3(npu_inst_pe_1_1_4_n7), .ZN(
        npu_inst_pe_1_1_4_n52) );
  OR3_X1 npu_inst_pe_1_1_4_U23 ( .A1(npu_inst_pe_1_1_4_n6), .A2(
        npu_inst_pe_1_1_4_n8), .A3(npu_inst_pe_1_1_4_n4), .ZN(
        npu_inst_pe_1_1_4_n60) );
  NOR2_X1 npu_inst_pe_1_1_4_U22 ( .A1(npu_inst_pe_1_1_4_n60), .A2(
        npu_inst_pe_1_1_4_n3), .ZN(npu_inst_pe_1_1_4_n58) );
  NOR2_X1 npu_inst_pe_1_1_4_U21 ( .A1(npu_inst_pe_1_1_4_n56), .A2(
        npu_inst_pe_1_1_4_n3), .ZN(npu_inst_pe_1_1_4_n54) );
  NOR2_X1 npu_inst_pe_1_1_4_U20 ( .A1(npu_inst_pe_1_1_4_n52), .A2(
        npu_inst_pe_1_1_4_n3), .ZN(npu_inst_pe_1_1_4_n50) );
  NOR2_X1 npu_inst_pe_1_1_4_U19 ( .A1(npu_inst_pe_1_1_4_n48), .A2(
        npu_inst_pe_1_1_4_n3), .ZN(npu_inst_pe_1_1_4_n46) );
  NOR2_X1 npu_inst_pe_1_1_4_U18 ( .A1(npu_inst_pe_1_1_4_n40), .A2(
        npu_inst_pe_1_1_4_n3), .ZN(npu_inst_pe_1_1_4_n38) );
  NOR2_X1 npu_inst_pe_1_1_4_U17 ( .A1(npu_inst_pe_1_1_4_n44), .A2(
        npu_inst_pe_1_1_4_n3), .ZN(npu_inst_pe_1_1_4_n42) );
  BUF_X1 npu_inst_pe_1_1_4_U16 ( .A(npu_inst_n104), .Z(npu_inst_pe_1_1_4_n8)
         );
  BUF_X1 npu_inst_pe_1_1_4_U15 ( .A(npu_inst_pe_1_1_4_n12), .Z(
        npu_inst_pe_1_1_4_n11) );
  BUF_X1 npu_inst_pe_1_1_4_U14 ( .A(npu_inst_pe_1_1_4_n12), .Z(
        npu_inst_pe_1_1_4_n10) );
  BUF_X1 npu_inst_pe_1_1_4_U13 ( .A(npu_inst_pe_1_1_4_n12), .Z(
        npu_inst_pe_1_1_4_n9) );
  INV_X1 npu_inst_pe_1_1_4_U12 ( .A(npu_inst_pe_1_1_4_n38), .ZN(
        npu_inst_pe_1_1_4_n118) );
  INV_X1 npu_inst_pe_1_1_4_U11 ( .A(npu_inst_pe_1_1_4_n58), .ZN(
        npu_inst_pe_1_1_4_n114) );
  INV_X1 npu_inst_pe_1_1_4_U10 ( .A(npu_inst_pe_1_1_4_n54), .ZN(
        npu_inst_pe_1_1_4_n115) );
  INV_X1 npu_inst_pe_1_1_4_U9 ( .A(npu_inst_pe_1_1_4_n50), .ZN(
        npu_inst_pe_1_1_4_n116) );
  INV_X1 npu_inst_pe_1_1_4_U8 ( .A(npu_inst_pe_1_1_4_n46), .ZN(
        npu_inst_pe_1_1_4_n117) );
  INV_X1 npu_inst_pe_1_1_4_U7 ( .A(npu_inst_pe_1_1_4_n42), .ZN(
        npu_inst_pe_1_1_4_n119) );
  BUF_X1 npu_inst_pe_1_1_4_U6 ( .A(npu_inst_n32), .Z(npu_inst_pe_1_1_4_n2) );
  BUF_X1 npu_inst_pe_1_1_4_U5 ( .A(npu_inst_n32), .Z(npu_inst_pe_1_1_4_n1) );
  NOR2_X1 npu_inst_pe_1_1_4_U4 ( .A1(npu_inst_pe_1_1_4_int_q_weight_0_), .A2(
        npu_inst_pe_1_1_4_n1), .ZN(npu_inst_pe_1_1_4_n76) );
  NOR2_X1 npu_inst_pe_1_1_4_U3 ( .A1(npu_inst_pe_1_1_4_n27), .A2(
        npu_inst_pe_1_1_4_n1), .ZN(npu_inst_pe_1_1_4_n77) );
  FA_X1 npu_inst_pe_1_1_4_sub_77_U2_1 ( .A(npu_inst_pe_1_1_4_int_q_acc_1_), 
        .B(npu_inst_pe_1_1_4_n14), .CI(npu_inst_pe_1_1_4_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_1_4_sub_77_carry_2_), .S(npu_inst_pe_1_1_4_N66) );
  FA_X1 npu_inst_pe_1_1_4_add_79_U1_1 ( .A(npu_inst_pe_1_1_4_int_q_acc_1_), 
        .B(npu_inst_pe_1_1_4_int_data_1_), .CI(
        npu_inst_pe_1_1_4_add_79_carry_1_), .CO(
        npu_inst_pe_1_1_4_add_79_carry_2_), .S(npu_inst_pe_1_1_4_N74) );
  NAND3_X1 npu_inst_pe_1_1_4_U109 ( .A1(npu_inst_pe_1_1_4_n5), .A2(
        npu_inst_pe_1_1_4_n7), .A3(npu_inst_pe_1_1_4_n8), .ZN(
        npu_inst_pe_1_1_4_n44) );
  NAND3_X1 npu_inst_pe_1_1_4_U108 ( .A1(npu_inst_pe_1_1_4_n4), .A2(
        npu_inst_pe_1_1_4_n7), .A3(npu_inst_pe_1_1_4_n8), .ZN(
        npu_inst_pe_1_1_4_n40) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_1_4_n34), .CK(
        npu_inst_pe_1_1_4_net4017), .RN(npu_inst_pe_1_1_4_n9), .Q(
        npu_inst_pe_1_1_4_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_1_4_n35), .CK(
        npu_inst_pe_1_1_4_net4017), .RN(npu_inst_pe_1_1_4_n9), .Q(
        npu_inst_pe_1_1_4_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_1_4_n36), .CK(
        npu_inst_pe_1_1_4_net4017), .RN(npu_inst_pe_1_1_4_n9), .Q(
        npu_inst_pe_1_1_4_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_1_4_n98), .CK(
        npu_inst_pe_1_1_4_net4017), .RN(npu_inst_pe_1_1_4_n9), .Q(
        npu_inst_pe_1_1_4_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_1_4_n99), .CK(
        npu_inst_pe_1_1_4_net4017), .RN(npu_inst_pe_1_1_4_n9), .Q(
        npu_inst_pe_1_1_4_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_1_4_n100), 
        .CK(npu_inst_pe_1_1_4_net4017), .RN(npu_inst_pe_1_1_4_n9), .Q(
        npu_inst_pe_1_1_4_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_1_4_n33), .CK(
        npu_inst_pe_1_1_4_net4017), .RN(npu_inst_pe_1_1_4_n9), .Q(
        npu_inst_pe_1_1_4_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_1_4_n101), 
        .CK(npu_inst_pe_1_1_4_net4017), .RN(npu_inst_pe_1_1_4_n9), .Q(
        npu_inst_pe_1_1_4_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_weight_reg_0_ ( .D(npu_inst_n112), .CK(
        npu_inst_pe_1_1_4_net4023), .RN(npu_inst_pe_1_1_4_n9), .Q(
        npu_inst_pe_1_1_4_int_q_weight_0_), .QN(npu_inst_pe_1_1_4_n27) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_weight_reg_1_ ( .D(npu_inst_n118), .CK(
        npu_inst_pe_1_1_4_net4023), .RN(npu_inst_pe_1_1_4_n9), .Q(
        npu_inst_pe_1_1_4_int_q_weight_1_), .QN(npu_inst_pe_1_1_4_n26) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_1_4_n113), 
        .CK(npu_inst_pe_1_1_4_net4023), .RN(npu_inst_pe_1_1_4_n9), .Q(
        npu_inst_pe_1_1_4_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_1_4_n107), 
        .CK(npu_inst_pe_1_1_4_net4023), .RN(npu_inst_pe_1_1_4_n9), .Q(
        npu_inst_pe_1_1_4_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_1_4_n112), 
        .CK(npu_inst_pe_1_1_4_net4023), .RN(npu_inst_pe_1_1_4_n10), .Q(
        npu_inst_pe_1_1_4_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_1_4_n106), 
        .CK(npu_inst_pe_1_1_4_net4023), .RN(npu_inst_pe_1_1_4_n10), .Q(
        npu_inst_pe_1_1_4_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_1_4_n111), 
        .CK(npu_inst_pe_1_1_4_net4023), .RN(npu_inst_pe_1_1_4_n10), .Q(
        npu_inst_pe_1_1_4_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_1_4_n105), 
        .CK(npu_inst_pe_1_1_4_net4023), .RN(npu_inst_pe_1_1_4_n10), .Q(
        npu_inst_pe_1_1_4_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_1_4_n110), 
        .CK(npu_inst_pe_1_1_4_net4023), .RN(npu_inst_pe_1_1_4_n10), .Q(
        npu_inst_pe_1_1_4_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_1_4_n104), 
        .CK(npu_inst_pe_1_1_4_net4023), .RN(npu_inst_pe_1_1_4_n10), .Q(
        npu_inst_pe_1_1_4_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_1_4_n109), 
        .CK(npu_inst_pe_1_1_4_net4023), .RN(npu_inst_pe_1_1_4_n10), .Q(
        npu_inst_pe_1_1_4_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_1_4_n103), 
        .CK(npu_inst_pe_1_1_4_net4023), .RN(npu_inst_pe_1_1_4_n10), .Q(
        npu_inst_pe_1_1_4_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_1_4_n108), 
        .CK(npu_inst_pe_1_1_4_net4023), .RN(npu_inst_pe_1_1_4_n10), .Q(
        npu_inst_pe_1_1_4_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_1_4_n102), 
        .CK(npu_inst_pe_1_1_4_net4023), .RN(npu_inst_pe_1_1_4_n10), .Q(
        npu_inst_pe_1_1_4_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_1_4_n86), 
        .CK(npu_inst_pe_1_1_4_net4023), .RN(npu_inst_pe_1_1_4_n10), .Q(
        npu_inst_pe_1_1_4_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_1_4_n87), 
        .CK(npu_inst_pe_1_1_4_net4023), .RN(npu_inst_pe_1_1_4_n10), .Q(
        npu_inst_pe_1_1_4_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_1_4_n88), 
        .CK(npu_inst_pe_1_1_4_net4023), .RN(npu_inst_pe_1_1_4_n11), .Q(
        npu_inst_pe_1_1_4_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_1_4_n89), 
        .CK(npu_inst_pe_1_1_4_net4023), .RN(npu_inst_pe_1_1_4_n11), .Q(
        npu_inst_pe_1_1_4_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_1_4_n90), 
        .CK(npu_inst_pe_1_1_4_net4023), .RN(npu_inst_pe_1_1_4_n11), .Q(
        npu_inst_pe_1_1_4_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_1_4_n91), 
        .CK(npu_inst_pe_1_1_4_net4023), .RN(npu_inst_pe_1_1_4_n11), .Q(
        npu_inst_pe_1_1_4_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_1_4_n92), 
        .CK(npu_inst_pe_1_1_4_net4023), .RN(npu_inst_pe_1_1_4_n11), .Q(
        npu_inst_pe_1_1_4_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_1_4_n93), 
        .CK(npu_inst_pe_1_1_4_net4023), .RN(npu_inst_pe_1_1_4_n11), .Q(
        npu_inst_pe_1_1_4_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_1_4_n94), 
        .CK(npu_inst_pe_1_1_4_net4023), .RN(npu_inst_pe_1_1_4_n11), .Q(
        npu_inst_pe_1_1_4_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_1_4_n95), 
        .CK(npu_inst_pe_1_1_4_net4023), .RN(npu_inst_pe_1_1_4_n11), .Q(
        npu_inst_pe_1_1_4_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_1_4_n96), 
        .CK(npu_inst_pe_1_1_4_net4023), .RN(npu_inst_pe_1_1_4_n11), .Q(
        npu_inst_pe_1_1_4_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_1_4_n97), 
        .CK(npu_inst_pe_1_1_4_net4023), .RN(npu_inst_pe_1_1_4_n11), .Q(
        npu_inst_pe_1_1_4_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_1_4_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_1_4_N84), .SE(1'b0), .GCK(npu_inst_pe_1_1_4_net4017) );
  CLKGATETST_X1 npu_inst_pe_1_1_4_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n65), .SE(1'b0), .GCK(npu_inst_pe_1_1_4_net4023) );
  MUX2_X1 npu_inst_pe_1_1_5_U162 ( .A(npu_inst_pe_1_1_5_n32), .B(
        npu_inst_pe_1_1_5_n29), .S(npu_inst_pe_1_1_5_n8), .Z(
        npu_inst_pe_1_1_5_N93) );
  MUX2_X1 npu_inst_pe_1_1_5_U161 ( .A(npu_inst_pe_1_1_5_n31), .B(
        npu_inst_pe_1_1_5_n30), .S(npu_inst_pe_1_1_5_n6), .Z(
        npu_inst_pe_1_1_5_n32) );
  MUX2_X1 npu_inst_pe_1_1_5_U160 ( .A(npu_inst_pe_1_1_5_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_1_5_int_q_reg_v_1__0_), .S(npu_inst_pe_1_1_5_n4), .Z(
        npu_inst_pe_1_1_5_n31) );
  MUX2_X1 npu_inst_pe_1_1_5_U159 ( .A(npu_inst_pe_1_1_5_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_1_5_int_q_reg_v_3__0_), .S(npu_inst_pe_1_1_5_n4), .Z(
        npu_inst_pe_1_1_5_n30) );
  MUX2_X1 npu_inst_pe_1_1_5_U158 ( .A(npu_inst_pe_1_1_5_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_1_5_int_q_reg_v_5__0_), .S(npu_inst_pe_1_1_5_n4), .Z(
        npu_inst_pe_1_1_5_n29) );
  MUX2_X1 npu_inst_pe_1_1_5_U157 ( .A(npu_inst_pe_1_1_5_n28), .B(
        npu_inst_pe_1_1_5_n23), .S(npu_inst_pe_1_1_5_n8), .Z(
        npu_inst_pe_1_1_5_N94) );
  MUX2_X1 npu_inst_pe_1_1_5_U156 ( .A(npu_inst_pe_1_1_5_n25), .B(
        npu_inst_pe_1_1_5_n24), .S(npu_inst_pe_1_1_5_n6), .Z(
        npu_inst_pe_1_1_5_n28) );
  MUX2_X1 npu_inst_pe_1_1_5_U155 ( .A(npu_inst_pe_1_1_5_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_1_5_int_q_reg_v_1__1_), .S(npu_inst_pe_1_1_5_n4), .Z(
        npu_inst_pe_1_1_5_n25) );
  MUX2_X1 npu_inst_pe_1_1_5_U154 ( .A(npu_inst_pe_1_1_5_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_1_5_int_q_reg_v_3__1_), .S(npu_inst_pe_1_1_5_n4), .Z(
        npu_inst_pe_1_1_5_n24) );
  MUX2_X1 npu_inst_pe_1_1_5_U153 ( .A(npu_inst_pe_1_1_5_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_1_5_int_q_reg_v_5__1_), .S(npu_inst_pe_1_1_5_n4), .Z(
        npu_inst_pe_1_1_5_n23) );
  MUX2_X1 npu_inst_pe_1_1_5_U152 ( .A(npu_inst_pe_1_1_5_n22), .B(
        npu_inst_pe_1_1_5_n19), .S(npu_inst_pe_1_1_5_n8), .Z(
        npu_inst_int_data_x_1__5__1_) );
  MUX2_X1 npu_inst_pe_1_1_5_U151 ( .A(npu_inst_pe_1_1_5_n21), .B(
        npu_inst_pe_1_1_5_n20), .S(npu_inst_pe_1_1_5_n6), .Z(
        npu_inst_pe_1_1_5_n22) );
  MUX2_X1 npu_inst_pe_1_1_5_U150 ( .A(npu_inst_pe_1_1_5_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_1_5_int_q_reg_h_1__1_), .S(npu_inst_pe_1_1_5_n4), .Z(
        npu_inst_pe_1_1_5_n21) );
  MUX2_X1 npu_inst_pe_1_1_5_U149 ( .A(npu_inst_pe_1_1_5_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_1_5_int_q_reg_h_3__1_), .S(npu_inst_pe_1_1_5_n4), .Z(
        npu_inst_pe_1_1_5_n20) );
  MUX2_X1 npu_inst_pe_1_1_5_U148 ( .A(npu_inst_pe_1_1_5_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_1_5_int_q_reg_h_5__1_), .S(npu_inst_pe_1_1_5_n4), .Z(
        npu_inst_pe_1_1_5_n19) );
  MUX2_X1 npu_inst_pe_1_1_5_U147 ( .A(npu_inst_pe_1_1_5_n18), .B(
        npu_inst_pe_1_1_5_n15), .S(npu_inst_pe_1_1_5_n8), .Z(
        npu_inst_int_data_x_1__5__0_) );
  MUX2_X1 npu_inst_pe_1_1_5_U146 ( .A(npu_inst_pe_1_1_5_n17), .B(
        npu_inst_pe_1_1_5_n16), .S(npu_inst_pe_1_1_5_n6), .Z(
        npu_inst_pe_1_1_5_n18) );
  MUX2_X1 npu_inst_pe_1_1_5_U145 ( .A(npu_inst_pe_1_1_5_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_1_5_int_q_reg_h_1__0_), .S(npu_inst_pe_1_1_5_n4), .Z(
        npu_inst_pe_1_1_5_n17) );
  MUX2_X1 npu_inst_pe_1_1_5_U144 ( .A(npu_inst_pe_1_1_5_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_1_5_int_q_reg_h_3__0_), .S(npu_inst_pe_1_1_5_n4), .Z(
        npu_inst_pe_1_1_5_n16) );
  MUX2_X1 npu_inst_pe_1_1_5_U143 ( .A(npu_inst_pe_1_1_5_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_1_5_int_q_reg_h_5__0_), .S(npu_inst_pe_1_1_5_n4), .Z(
        npu_inst_pe_1_1_5_n15) );
  XOR2_X1 npu_inst_pe_1_1_5_U142 ( .A(npu_inst_pe_1_1_5_int_data_0_), .B(
        npu_inst_pe_1_1_5_int_q_acc_0_), .Z(npu_inst_pe_1_1_5_N73) );
  AND2_X1 npu_inst_pe_1_1_5_U141 ( .A1(npu_inst_pe_1_1_5_int_q_acc_0_), .A2(
        npu_inst_pe_1_1_5_int_data_0_), .ZN(npu_inst_pe_1_1_5_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_1_5_U140 ( .A(npu_inst_pe_1_1_5_int_q_acc_0_), .B(
        npu_inst_pe_1_1_5_n13), .ZN(npu_inst_pe_1_1_5_N65) );
  OR2_X1 npu_inst_pe_1_1_5_U139 ( .A1(npu_inst_pe_1_1_5_n13), .A2(
        npu_inst_pe_1_1_5_int_q_acc_0_), .ZN(npu_inst_pe_1_1_5_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_1_5_U138 ( .A(npu_inst_pe_1_1_5_int_q_acc_2_), .B(
        npu_inst_pe_1_1_5_add_79_carry_2_), .Z(npu_inst_pe_1_1_5_N75) );
  AND2_X1 npu_inst_pe_1_1_5_U137 ( .A1(npu_inst_pe_1_1_5_add_79_carry_2_), 
        .A2(npu_inst_pe_1_1_5_int_q_acc_2_), .ZN(
        npu_inst_pe_1_1_5_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_1_5_U136 ( .A(npu_inst_pe_1_1_5_int_q_acc_3_), .B(
        npu_inst_pe_1_1_5_add_79_carry_3_), .Z(npu_inst_pe_1_1_5_N76) );
  AND2_X1 npu_inst_pe_1_1_5_U135 ( .A1(npu_inst_pe_1_1_5_add_79_carry_3_), 
        .A2(npu_inst_pe_1_1_5_int_q_acc_3_), .ZN(
        npu_inst_pe_1_1_5_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_1_5_U134 ( .A(npu_inst_pe_1_1_5_int_q_acc_4_), .B(
        npu_inst_pe_1_1_5_add_79_carry_4_), .Z(npu_inst_pe_1_1_5_N77) );
  AND2_X1 npu_inst_pe_1_1_5_U133 ( .A1(npu_inst_pe_1_1_5_add_79_carry_4_), 
        .A2(npu_inst_pe_1_1_5_int_q_acc_4_), .ZN(
        npu_inst_pe_1_1_5_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_1_5_U132 ( .A(npu_inst_pe_1_1_5_int_q_acc_5_), .B(
        npu_inst_pe_1_1_5_add_79_carry_5_), .Z(npu_inst_pe_1_1_5_N78) );
  AND2_X1 npu_inst_pe_1_1_5_U131 ( .A1(npu_inst_pe_1_1_5_add_79_carry_5_), 
        .A2(npu_inst_pe_1_1_5_int_q_acc_5_), .ZN(
        npu_inst_pe_1_1_5_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_1_5_U130 ( .A(npu_inst_pe_1_1_5_int_q_acc_6_), .B(
        npu_inst_pe_1_1_5_add_79_carry_6_), .Z(npu_inst_pe_1_1_5_N79) );
  AND2_X1 npu_inst_pe_1_1_5_U129 ( .A1(npu_inst_pe_1_1_5_add_79_carry_6_), 
        .A2(npu_inst_pe_1_1_5_int_q_acc_6_), .ZN(
        npu_inst_pe_1_1_5_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_1_5_U128 ( .A(npu_inst_pe_1_1_5_int_q_acc_7_), .B(
        npu_inst_pe_1_1_5_add_79_carry_7_), .Z(npu_inst_pe_1_1_5_N80) );
  XNOR2_X1 npu_inst_pe_1_1_5_U127 ( .A(npu_inst_pe_1_1_5_sub_77_carry_2_), .B(
        npu_inst_pe_1_1_5_int_q_acc_2_), .ZN(npu_inst_pe_1_1_5_N67) );
  OR2_X1 npu_inst_pe_1_1_5_U126 ( .A1(npu_inst_pe_1_1_5_int_q_acc_2_), .A2(
        npu_inst_pe_1_1_5_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_1_5_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_1_5_U125 ( .A(npu_inst_pe_1_1_5_sub_77_carry_3_), .B(
        npu_inst_pe_1_1_5_int_q_acc_3_), .ZN(npu_inst_pe_1_1_5_N68) );
  OR2_X1 npu_inst_pe_1_1_5_U124 ( .A1(npu_inst_pe_1_1_5_int_q_acc_3_), .A2(
        npu_inst_pe_1_1_5_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_1_5_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_1_5_U123 ( .A(npu_inst_pe_1_1_5_sub_77_carry_4_), .B(
        npu_inst_pe_1_1_5_int_q_acc_4_), .ZN(npu_inst_pe_1_1_5_N69) );
  OR2_X1 npu_inst_pe_1_1_5_U122 ( .A1(npu_inst_pe_1_1_5_int_q_acc_4_), .A2(
        npu_inst_pe_1_1_5_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_1_5_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_1_5_U121 ( .A(npu_inst_pe_1_1_5_sub_77_carry_5_), .B(
        npu_inst_pe_1_1_5_int_q_acc_5_), .ZN(npu_inst_pe_1_1_5_N70) );
  OR2_X1 npu_inst_pe_1_1_5_U120 ( .A1(npu_inst_pe_1_1_5_int_q_acc_5_), .A2(
        npu_inst_pe_1_1_5_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_1_5_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_1_5_U119 ( .A(npu_inst_pe_1_1_5_sub_77_carry_6_), .B(
        npu_inst_pe_1_1_5_int_q_acc_6_), .ZN(npu_inst_pe_1_1_5_N71) );
  OR2_X1 npu_inst_pe_1_1_5_U118 ( .A1(npu_inst_pe_1_1_5_int_q_acc_6_), .A2(
        npu_inst_pe_1_1_5_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_1_5_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_1_5_U117 ( .A(npu_inst_pe_1_1_5_int_q_acc_7_), .B(
        npu_inst_pe_1_1_5_sub_77_carry_7_), .ZN(npu_inst_pe_1_1_5_N72) );
  INV_X1 npu_inst_pe_1_1_5_U116 ( .A(npu_inst_n79), .ZN(npu_inst_pe_1_1_5_n7)
         );
  INV_X1 npu_inst_pe_1_1_5_U115 ( .A(npu_inst_pe_1_1_5_n7), .ZN(
        npu_inst_pe_1_1_5_n6) );
  INV_X1 npu_inst_pe_1_1_5_U114 ( .A(npu_inst_n59), .ZN(npu_inst_pe_1_1_5_n3)
         );
  AOI22_X1 npu_inst_pe_1_1_5_U113 ( .A1(npu_inst_int_data_y_2__5__0_), .A2(
        npu_inst_pe_1_1_5_n58), .B1(npu_inst_pe_1_1_5_n114), .B2(
        npu_inst_pe_1_1_5_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_1_5_n57) );
  INV_X1 npu_inst_pe_1_1_5_U112 ( .A(npu_inst_pe_1_1_5_n57), .ZN(
        npu_inst_pe_1_1_5_n108) );
  AOI22_X1 npu_inst_pe_1_1_5_U111 ( .A1(npu_inst_int_data_y_2__5__0_), .A2(
        npu_inst_pe_1_1_5_n54), .B1(npu_inst_pe_1_1_5_n115), .B2(
        npu_inst_pe_1_1_5_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_1_5_n53) );
  INV_X1 npu_inst_pe_1_1_5_U110 ( .A(npu_inst_pe_1_1_5_n53), .ZN(
        npu_inst_pe_1_1_5_n109) );
  AOI22_X1 npu_inst_pe_1_1_5_U107 ( .A1(npu_inst_int_data_y_2__5__0_), .A2(
        npu_inst_pe_1_1_5_n50), .B1(npu_inst_pe_1_1_5_n116), .B2(
        npu_inst_pe_1_1_5_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_1_5_n49) );
  INV_X1 npu_inst_pe_1_1_5_U106 ( .A(npu_inst_pe_1_1_5_n49), .ZN(
        npu_inst_pe_1_1_5_n110) );
  AOI22_X1 npu_inst_pe_1_1_5_U105 ( .A1(npu_inst_int_data_y_2__5__0_), .A2(
        npu_inst_pe_1_1_5_n46), .B1(npu_inst_pe_1_1_5_n117), .B2(
        npu_inst_pe_1_1_5_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_1_5_n45) );
  INV_X1 npu_inst_pe_1_1_5_U104 ( .A(npu_inst_pe_1_1_5_n45), .ZN(
        npu_inst_pe_1_1_5_n111) );
  AOI22_X1 npu_inst_pe_1_1_5_U103 ( .A1(npu_inst_int_data_y_2__5__0_), .A2(
        npu_inst_pe_1_1_5_n42), .B1(npu_inst_pe_1_1_5_n119), .B2(
        npu_inst_pe_1_1_5_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_1_5_n41) );
  INV_X1 npu_inst_pe_1_1_5_U102 ( .A(npu_inst_pe_1_1_5_n41), .ZN(
        npu_inst_pe_1_1_5_n112) );
  AOI22_X1 npu_inst_pe_1_1_5_U101 ( .A1(npu_inst_int_data_y_2__5__1_), .A2(
        npu_inst_pe_1_1_5_n58), .B1(npu_inst_pe_1_1_5_n114), .B2(
        npu_inst_pe_1_1_5_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_1_5_n59) );
  INV_X1 npu_inst_pe_1_1_5_U100 ( .A(npu_inst_pe_1_1_5_n59), .ZN(
        npu_inst_pe_1_1_5_n102) );
  AOI22_X1 npu_inst_pe_1_1_5_U99 ( .A1(npu_inst_int_data_y_2__5__1_), .A2(
        npu_inst_pe_1_1_5_n54), .B1(npu_inst_pe_1_1_5_n115), .B2(
        npu_inst_pe_1_1_5_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_1_5_n55) );
  INV_X1 npu_inst_pe_1_1_5_U98 ( .A(npu_inst_pe_1_1_5_n55), .ZN(
        npu_inst_pe_1_1_5_n103) );
  AOI22_X1 npu_inst_pe_1_1_5_U97 ( .A1(npu_inst_int_data_y_2__5__1_), .A2(
        npu_inst_pe_1_1_5_n50), .B1(npu_inst_pe_1_1_5_n116), .B2(
        npu_inst_pe_1_1_5_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_1_5_n51) );
  INV_X1 npu_inst_pe_1_1_5_U96 ( .A(npu_inst_pe_1_1_5_n51), .ZN(
        npu_inst_pe_1_1_5_n104) );
  AOI22_X1 npu_inst_pe_1_1_5_U95 ( .A1(npu_inst_int_data_y_2__5__1_), .A2(
        npu_inst_pe_1_1_5_n46), .B1(npu_inst_pe_1_1_5_n117), .B2(
        npu_inst_pe_1_1_5_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_1_5_n47) );
  INV_X1 npu_inst_pe_1_1_5_U94 ( .A(npu_inst_pe_1_1_5_n47), .ZN(
        npu_inst_pe_1_1_5_n105) );
  AOI22_X1 npu_inst_pe_1_1_5_U93 ( .A1(npu_inst_int_data_y_2__5__1_), .A2(
        npu_inst_pe_1_1_5_n42), .B1(npu_inst_pe_1_1_5_n119), .B2(
        npu_inst_pe_1_1_5_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_1_5_n43) );
  INV_X1 npu_inst_pe_1_1_5_U92 ( .A(npu_inst_pe_1_1_5_n43), .ZN(
        npu_inst_pe_1_1_5_n106) );
  AOI22_X1 npu_inst_pe_1_1_5_U91 ( .A1(npu_inst_pe_1_1_5_n38), .A2(
        npu_inst_int_data_y_2__5__1_), .B1(npu_inst_pe_1_1_5_n118), .B2(
        npu_inst_pe_1_1_5_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_1_5_n39) );
  INV_X1 npu_inst_pe_1_1_5_U90 ( .A(npu_inst_pe_1_1_5_n39), .ZN(
        npu_inst_pe_1_1_5_n107) );
  AOI22_X1 npu_inst_pe_1_1_5_U89 ( .A1(npu_inst_pe_1_1_5_n38), .A2(
        npu_inst_int_data_y_2__5__0_), .B1(npu_inst_pe_1_1_5_n118), .B2(
        npu_inst_pe_1_1_5_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_1_5_n37) );
  INV_X1 npu_inst_pe_1_1_5_U88 ( .A(npu_inst_pe_1_1_5_n37), .ZN(
        npu_inst_pe_1_1_5_n113) );
  NAND2_X1 npu_inst_pe_1_1_5_U87 ( .A1(npu_inst_pe_1_1_5_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_1_5_n60), .ZN(npu_inst_pe_1_1_5_n74) );
  OAI21_X1 npu_inst_pe_1_1_5_U86 ( .B1(npu_inst_pe_1_1_5_n63), .B2(
        npu_inst_pe_1_1_5_n60), .A(npu_inst_pe_1_1_5_n74), .ZN(
        npu_inst_pe_1_1_5_n97) );
  NAND2_X1 npu_inst_pe_1_1_5_U85 ( .A1(npu_inst_pe_1_1_5_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_1_5_n60), .ZN(npu_inst_pe_1_1_5_n73) );
  OAI21_X1 npu_inst_pe_1_1_5_U84 ( .B1(npu_inst_pe_1_1_5_n61), .B2(
        npu_inst_pe_1_1_5_n60), .A(npu_inst_pe_1_1_5_n73), .ZN(
        npu_inst_pe_1_1_5_n96) );
  NAND2_X1 npu_inst_pe_1_1_5_U83 ( .A1(npu_inst_pe_1_1_5_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_1_5_n56), .ZN(npu_inst_pe_1_1_5_n72) );
  OAI21_X1 npu_inst_pe_1_1_5_U82 ( .B1(npu_inst_pe_1_1_5_n63), .B2(
        npu_inst_pe_1_1_5_n56), .A(npu_inst_pe_1_1_5_n72), .ZN(
        npu_inst_pe_1_1_5_n95) );
  NAND2_X1 npu_inst_pe_1_1_5_U81 ( .A1(npu_inst_pe_1_1_5_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_1_5_n56), .ZN(npu_inst_pe_1_1_5_n71) );
  OAI21_X1 npu_inst_pe_1_1_5_U80 ( .B1(npu_inst_pe_1_1_5_n61), .B2(
        npu_inst_pe_1_1_5_n56), .A(npu_inst_pe_1_1_5_n71), .ZN(
        npu_inst_pe_1_1_5_n94) );
  NAND2_X1 npu_inst_pe_1_1_5_U79 ( .A1(npu_inst_pe_1_1_5_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_1_5_n52), .ZN(npu_inst_pe_1_1_5_n70) );
  OAI21_X1 npu_inst_pe_1_1_5_U78 ( .B1(npu_inst_pe_1_1_5_n63), .B2(
        npu_inst_pe_1_1_5_n52), .A(npu_inst_pe_1_1_5_n70), .ZN(
        npu_inst_pe_1_1_5_n93) );
  NAND2_X1 npu_inst_pe_1_1_5_U77 ( .A1(npu_inst_pe_1_1_5_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_1_5_n52), .ZN(npu_inst_pe_1_1_5_n69) );
  OAI21_X1 npu_inst_pe_1_1_5_U76 ( .B1(npu_inst_pe_1_1_5_n61), .B2(
        npu_inst_pe_1_1_5_n52), .A(npu_inst_pe_1_1_5_n69), .ZN(
        npu_inst_pe_1_1_5_n92) );
  NAND2_X1 npu_inst_pe_1_1_5_U75 ( .A1(npu_inst_pe_1_1_5_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_1_5_n48), .ZN(npu_inst_pe_1_1_5_n68) );
  OAI21_X1 npu_inst_pe_1_1_5_U74 ( .B1(npu_inst_pe_1_1_5_n63), .B2(
        npu_inst_pe_1_1_5_n48), .A(npu_inst_pe_1_1_5_n68), .ZN(
        npu_inst_pe_1_1_5_n91) );
  NAND2_X1 npu_inst_pe_1_1_5_U73 ( .A1(npu_inst_pe_1_1_5_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_1_5_n48), .ZN(npu_inst_pe_1_1_5_n67) );
  OAI21_X1 npu_inst_pe_1_1_5_U72 ( .B1(npu_inst_pe_1_1_5_n61), .B2(
        npu_inst_pe_1_1_5_n48), .A(npu_inst_pe_1_1_5_n67), .ZN(
        npu_inst_pe_1_1_5_n90) );
  NAND2_X1 npu_inst_pe_1_1_5_U71 ( .A1(npu_inst_pe_1_1_5_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_1_5_n44), .ZN(npu_inst_pe_1_1_5_n66) );
  OAI21_X1 npu_inst_pe_1_1_5_U70 ( .B1(npu_inst_pe_1_1_5_n63), .B2(
        npu_inst_pe_1_1_5_n44), .A(npu_inst_pe_1_1_5_n66), .ZN(
        npu_inst_pe_1_1_5_n89) );
  NAND2_X1 npu_inst_pe_1_1_5_U69 ( .A1(npu_inst_pe_1_1_5_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_1_5_n44), .ZN(npu_inst_pe_1_1_5_n65) );
  OAI21_X1 npu_inst_pe_1_1_5_U68 ( .B1(npu_inst_pe_1_1_5_n61), .B2(
        npu_inst_pe_1_1_5_n44), .A(npu_inst_pe_1_1_5_n65), .ZN(
        npu_inst_pe_1_1_5_n88) );
  NAND2_X1 npu_inst_pe_1_1_5_U67 ( .A1(npu_inst_pe_1_1_5_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_1_5_n40), .ZN(npu_inst_pe_1_1_5_n64) );
  OAI21_X1 npu_inst_pe_1_1_5_U66 ( .B1(npu_inst_pe_1_1_5_n63), .B2(
        npu_inst_pe_1_1_5_n40), .A(npu_inst_pe_1_1_5_n64), .ZN(
        npu_inst_pe_1_1_5_n87) );
  NAND2_X1 npu_inst_pe_1_1_5_U65 ( .A1(npu_inst_pe_1_1_5_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_1_5_n40), .ZN(npu_inst_pe_1_1_5_n62) );
  OAI21_X1 npu_inst_pe_1_1_5_U64 ( .B1(npu_inst_pe_1_1_5_n61), .B2(
        npu_inst_pe_1_1_5_n40), .A(npu_inst_pe_1_1_5_n62), .ZN(
        npu_inst_pe_1_1_5_n86) );
  AND2_X1 npu_inst_pe_1_1_5_U63 ( .A1(npu_inst_pe_1_1_5_N93), .A2(npu_inst_n59), .ZN(npu_inst_int_data_y_1__5__0_) );
  AND2_X1 npu_inst_pe_1_1_5_U62 ( .A1(npu_inst_n59), .A2(npu_inst_pe_1_1_5_N94), .ZN(npu_inst_int_data_y_1__5__1_) );
  NOR3_X1 npu_inst_pe_1_1_5_U61 ( .A1(npu_inst_pe_1_1_5_n26), .A2(npu_inst_n59), .A3(npu_inst_int_ckg[50]), .ZN(npu_inst_pe_1_1_5_n85) );
  OR2_X1 npu_inst_pe_1_1_5_U60 ( .A1(npu_inst_pe_1_1_5_n85), .A2(
        npu_inst_pe_1_1_5_n2), .ZN(npu_inst_pe_1_1_5_N84) );
  AND2_X1 npu_inst_pe_1_1_5_U59 ( .A1(npu_inst_pe_1_1_5_int_q_acc_0_), .A2(
        npu_inst_pe_1_1_5_n1), .ZN(npu_inst_int_data_res_1__5__0_) );
  AND2_X1 npu_inst_pe_1_1_5_U58 ( .A1(npu_inst_pe_1_1_5_n2), .A2(
        npu_inst_pe_1_1_5_int_q_acc_7_), .ZN(npu_inst_int_data_res_1__5__7_)
         );
  AND2_X1 npu_inst_pe_1_1_5_U57 ( .A1(npu_inst_pe_1_1_5_int_q_acc_1_), .A2(
        npu_inst_pe_1_1_5_n1), .ZN(npu_inst_int_data_res_1__5__1_) );
  AND2_X1 npu_inst_pe_1_1_5_U56 ( .A1(npu_inst_pe_1_1_5_int_q_acc_2_), .A2(
        npu_inst_pe_1_1_5_n1), .ZN(npu_inst_int_data_res_1__5__2_) );
  AND2_X1 npu_inst_pe_1_1_5_U55 ( .A1(npu_inst_pe_1_1_5_int_q_acc_3_), .A2(
        npu_inst_pe_1_1_5_n2), .ZN(npu_inst_int_data_res_1__5__3_) );
  AND2_X1 npu_inst_pe_1_1_5_U54 ( .A1(npu_inst_pe_1_1_5_int_q_acc_4_), .A2(
        npu_inst_pe_1_1_5_n2), .ZN(npu_inst_int_data_res_1__5__4_) );
  AND2_X1 npu_inst_pe_1_1_5_U53 ( .A1(npu_inst_pe_1_1_5_int_q_acc_5_), .A2(
        npu_inst_pe_1_1_5_n2), .ZN(npu_inst_int_data_res_1__5__5_) );
  AND2_X1 npu_inst_pe_1_1_5_U52 ( .A1(npu_inst_pe_1_1_5_int_q_acc_6_), .A2(
        npu_inst_pe_1_1_5_n2), .ZN(npu_inst_int_data_res_1__5__6_) );
  AOI222_X1 npu_inst_pe_1_1_5_U51 ( .A1(npu_inst_int_data_res_2__5__0_), .A2(
        npu_inst_pe_1_1_5_n1), .B1(npu_inst_pe_1_1_5_N73), .B2(
        npu_inst_pe_1_1_5_n76), .C1(npu_inst_pe_1_1_5_N65), .C2(
        npu_inst_pe_1_1_5_n77), .ZN(npu_inst_pe_1_1_5_n84) );
  INV_X1 npu_inst_pe_1_1_5_U50 ( .A(npu_inst_pe_1_1_5_n84), .ZN(
        npu_inst_pe_1_1_5_n101) );
  AOI222_X1 npu_inst_pe_1_1_5_U49 ( .A1(npu_inst_int_data_res_2__5__7_), .A2(
        npu_inst_pe_1_1_5_n1), .B1(npu_inst_pe_1_1_5_N80), .B2(
        npu_inst_pe_1_1_5_n76), .C1(npu_inst_pe_1_1_5_N72), .C2(
        npu_inst_pe_1_1_5_n77), .ZN(npu_inst_pe_1_1_5_n75) );
  INV_X1 npu_inst_pe_1_1_5_U48 ( .A(npu_inst_pe_1_1_5_n75), .ZN(
        npu_inst_pe_1_1_5_n33) );
  AOI222_X1 npu_inst_pe_1_1_5_U47 ( .A1(npu_inst_int_data_res_2__5__1_), .A2(
        npu_inst_pe_1_1_5_n1), .B1(npu_inst_pe_1_1_5_N74), .B2(
        npu_inst_pe_1_1_5_n76), .C1(npu_inst_pe_1_1_5_N66), .C2(
        npu_inst_pe_1_1_5_n77), .ZN(npu_inst_pe_1_1_5_n83) );
  INV_X1 npu_inst_pe_1_1_5_U46 ( .A(npu_inst_pe_1_1_5_n83), .ZN(
        npu_inst_pe_1_1_5_n100) );
  AOI222_X1 npu_inst_pe_1_1_5_U45 ( .A1(npu_inst_int_data_res_2__5__2_), .A2(
        npu_inst_pe_1_1_5_n1), .B1(npu_inst_pe_1_1_5_N75), .B2(
        npu_inst_pe_1_1_5_n76), .C1(npu_inst_pe_1_1_5_N67), .C2(
        npu_inst_pe_1_1_5_n77), .ZN(npu_inst_pe_1_1_5_n82) );
  INV_X1 npu_inst_pe_1_1_5_U44 ( .A(npu_inst_pe_1_1_5_n82), .ZN(
        npu_inst_pe_1_1_5_n99) );
  AOI222_X1 npu_inst_pe_1_1_5_U43 ( .A1(npu_inst_int_data_res_2__5__3_), .A2(
        npu_inst_pe_1_1_5_n1), .B1(npu_inst_pe_1_1_5_N76), .B2(
        npu_inst_pe_1_1_5_n76), .C1(npu_inst_pe_1_1_5_N68), .C2(
        npu_inst_pe_1_1_5_n77), .ZN(npu_inst_pe_1_1_5_n81) );
  INV_X1 npu_inst_pe_1_1_5_U42 ( .A(npu_inst_pe_1_1_5_n81), .ZN(
        npu_inst_pe_1_1_5_n98) );
  AOI222_X1 npu_inst_pe_1_1_5_U41 ( .A1(npu_inst_int_data_res_2__5__4_), .A2(
        npu_inst_pe_1_1_5_n1), .B1(npu_inst_pe_1_1_5_N77), .B2(
        npu_inst_pe_1_1_5_n76), .C1(npu_inst_pe_1_1_5_N69), .C2(
        npu_inst_pe_1_1_5_n77), .ZN(npu_inst_pe_1_1_5_n80) );
  INV_X1 npu_inst_pe_1_1_5_U40 ( .A(npu_inst_pe_1_1_5_n80), .ZN(
        npu_inst_pe_1_1_5_n36) );
  AOI222_X1 npu_inst_pe_1_1_5_U39 ( .A1(npu_inst_int_data_res_2__5__5_), .A2(
        npu_inst_pe_1_1_5_n1), .B1(npu_inst_pe_1_1_5_N78), .B2(
        npu_inst_pe_1_1_5_n76), .C1(npu_inst_pe_1_1_5_N70), .C2(
        npu_inst_pe_1_1_5_n77), .ZN(npu_inst_pe_1_1_5_n79) );
  INV_X1 npu_inst_pe_1_1_5_U38 ( .A(npu_inst_pe_1_1_5_n79), .ZN(
        npu_inst_pe_1_1_5_n35) );
  AOI222_X1 npu_inst_pe_1_1_5_U37 ( .A1(npu_inst_int_data_res_2__5__6_), .A2(
        npu_inst_pe_1_1_5_n1), .B1(npu_inst_pe_1_1_5_N79), .B2(
        npu_inst_pe_1_1_5_n76), .C1(npu_inst_pe_1_1_5_N71), .C2(
        npu_inst_pe_1_1_5_n77), .ZN(npu_inst_pe_1_1_5_n78) );
  INV_X1 npu_inst_pe_1_1_5_U36 ( .A(npu_inst_pe_1_1_5_n78), .ZN(
        npu_inst_pe_1_1_5_n34) );
  INV_X1 npu_inst_pe_1_1_5_U35 ( .A(npu_inst_pe_1_1_5_int_data_1_), .ZN(
        npu_inst_pe_1_1_5_n14) );
  AND2_X1 npu_inst_pe_1_1_5_U34 ( .A1(npu_inst_int_data_x_1__5__1_), .A2(
        npu_inst_pe_1_1_5_int_q_weight_1_), .ZN(npu_inst_pe_1_1_5_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_1_5_U33 ( .A1(npu_inst_int_data_x_1__5__0_), .A2(
        npu_inst_pe_1_1_5_int_q_weight_1_), .ZN(npu_inst_pe_1_1_5_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_1_5_U32 ( .A1(npu_inst_n59), .A2(
        npu_inst_int_data_y_2__5__1_), .B1(npu_inst_pe_1_1_5_n3), .B2(
        npu_inst_int_data_x_1__6__1_), .ZN(npu_inst_pe_1_1_5_n63) );
  AOI22_X1 npu_inst_pe_1_1_5_U31 ( .A1(npu_inst_n59), .A2(
        npu_inst_int_data_y_2__5__0_), .B1(npu_inst_pe_1_1_5_n3), .B2(
        npu_inst_int_data_x_1__6__0_), .ZN(npu_inst_pe_1_1_5_n61) );
  INV_X1 npu_inst_pe_1_1_5_U30 ( .A(npu_inst_pe_1_1_5_int_data_0_), .ZN(
        npu_inst_pe_1_1_5_n13) );
  INV_X1 npu_inst_pe_1_1_5_U29 ( .A(npu_inst_n71), .ZN(npu_inst_pe_1_1_5_n5)
         );
  OR3_X1 npu_inst_pe_1_1_5_U28 ( .A1(npu_inst_pe_1_1_5_n6), .A2(
        npu_inst_pe_1_1_5_n8), .A3(npu_inst_pe_1_1_5_n5), .ZN(
        npu_inst_pe_1_1_5_n56) );
  OR3_X1 npu_inst_pe_1_1_5_U27 ( .A1(npu_inst_pe_1_1_5_n5), .A2(
        npu_inst_pe_1_1_5_n8), .A3(npu_inst_pe_1_1_5_n7), .ZN(
        npu_inst_pe_1_1_5_n48) );
  INV_X1 npu_inst_pe_1_1_5_U26 ( .A(npu_inst_pe_1_1_5_n5), .ZN(
        npu_inst_pe_1_1_5_n4) );
  INV_X1 npu_inst_pe_1_1_5_U25 ( .A(npu_inst_n126), .ZN(npu_inst_pe_1_1_5_n12)
         );
  OR3_X1 npu_inst_pe_1_1_5_U24 ( .A1(npu_inst_pe_1_1_5_n4), .A2(
        npu_inst_pe_1_1_5_n8), .A3(npu_inst_pe_1_1_5_n7), .ZN(
        npu_inst_pe_1_1_5_n52) );
  OR3_X1 npu_inst_pe_1_1_5_U23 ( .A1(npu_inst_pe_1_1_5_n6), .A2(
        npu_inst_pe_1_1_5_n8), .A3(npu_inst_pe_1_1_5_n4), .ZN(
        npu_inst_pe_1_1_5_n60) );
  NOR2_X1 npu_inst_pe_1_1_5_U22 ( .A1(npu_inst_pe_1_1_5_n60), .A2(
        npu_inst_pe_1_1_5_n3), .ZN(npu_inst_pe_1_1_5_n58) );
  NOR2_X1 npu_inst_pe_1_1_5_U21 ( .A1(npu_inst_pe_1_1_5_n56), .A2(
        npu_inst_pe_1_1_5_n3), .ZN(npu_inst_pe_1_1_5_n54) );
  NOR2_X1 npu_inst_pe_1_1_5_U20 ( .A1(npu_inst_pe_1_1_5_n52), .A2(
        npu_inst_pe_1_1_5_n3), .ZN(npu_inst_pe_1_1_5_n50) );
  NOR2_X1 npu_inst_pe_1_1_5_U19 ( .A1(npu_inst_pe_1_1_5_n48), .A2(
        npu_inst_pe_1_1_5_n3), .ZN(npu_inst_pe_1_1_5_n46) );
  NOR2_X1 npu_inst_pe_1_1_5_U18 ( .A1(npu_inst_pe_1_1_5_n40), .A2(
        npu_inst_pe_1_1_5_n3), .ZN(npu_inst_pe_1_1_5_n38) );
  NOR2_X1 npu_inst_pe_1_1_5_U17 ( .A1(npu_inst_pe_1_1_5_n44), .A2(
        npu_inst_pe_1_1_5_n3), .ZN(npu_inst_pe_1_1_5_n42) );
  BUF_X1 npu_inst_pe_1_1_5_U16 ( .A(npu_inst_n104), .Z(npu_inst_pe_1_1_5_n8)
         );
  BUF_X1 npu_inst_pe_1_1_5_U15 ( .A(npu_inst_pe_1_1_5_n12), .Z(
        npu_inst_pe_1_1_5_n11) );
  BUF_X1 npu_inst_pe_1_1_5_U14 ( .A(npu_inst_pe_1_1_5_n12), .Z(
        npu_inst_pe_1_1_5_n10) );
  BUF_X1 npu_inst_pe_1_1_5_U13 ( .A(npu_inst_pe_1_1_5_n12), .Z(
        npu_inst_pe_1_1_5_n9) );
  INV_X1 npu_inst_pe_1_1_5_U12 ( .A(npu_inst_pe_1_1_5_n38), .ZN(
        npu_inst_pe_1_1_5_n118) );
  INV_X1 npu_inst_pe_1_1_5_U11 ( .A(npu_inst_pe_1_1_5_n58), .ZN(
        npu_inst_pe_1_1_5_n114) );
  INV_X1 npu_inst_pe_1_1_5_U10 ( .A(npu_inst_pe_1_1_5_n54), .ZN(
        npu_inst_pe_1_1_5_n115) );
  INV_X1 npu_inst_pe_1_1_5_U9 ( .A(npu_inst_pe_1_1_5_n50), .ZN(
        npu_inst_pe_1_1_5_n116) );
  INV_X1 npu_inst_pe_1_1_5_U8 ( .A(npu_inst_pe_1_1_5_n46), .ZN(
        npu_inst_pe_1_1_5_n117) );
  INV_X1 npu_inst_pe_1_1_5_U7 ( .A(npu_inst_pe_1_1_5_n42), .ZN(
        npu_inst_pe_1_1_5_n119) );
  BUF_X1 npu_inst_pe_1_1_5_U6 ( .A(npu_inst_n32), .Z(npu_inst_pe_1_1_5_n2) );
  BUF_X1 npu_inst_pe_1_1_5_U5 ( .A(npu_inst_n32), .Z(npu_inst_pe_1_1_5_n1) );
  NOR2_X1 npu_inst_pe_1_1_5_U4 ( .A1(npu_inst_pe_1_1_5_int_q_weight_0_), .A2(
        npu_inst_pe_1_1_5_n1), .ZN(npu_inst_pe_1_1_5_n76) );
  NOR2_X1 npu_inst_pe_1_1_5_U3 ( .A1(npu_inst_pe_1_1_5_n27), .A2(
        npu_inst_pe_1_1_5_n1), .ZN(npu_inst_pe_1_1_5_n77) );
  FA_X1 npu_inst_pe_1_1_5_sub_77_U2_1 ( .A(npu_inst_pe_1_1_5_int_q_acc_1_), 
        .B(npu_inst_pe_1_1_5_n14), .CI(npu_inst_pe_1_1_5_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_1_5_sub_77_carry_2_), .S(npu_inst_pe_1_1_5_N66) );
  FA_X1 npu_inst_pe_1_1_5_add_79_U1_1 ( .A(npu_inst_pe_1_1_5_int_q_acc_1_), 
        .B(npu_inst_pe_1_1_5_int_data_1_), .CI(
        npu_inst_pe_1_1_5_add_79_carry_1_), .CO(
        npu_inst_pe_1_1_5_add_79_carry_2_), .S(npu_inst_pe_1_1_5_N74) );
  NAND3_X1 npu_inst_pe_1_1_5_U109 ( .A1(npu_inst_pe_1_1_5_n5), .A2(
        npu_inst_pe_1_1_5_n7), .A3(npu_inst_pe_1_1_5_n8), .ZN(
        npu_inst_pe_1_1_5_n44) );
  NAND3_X1 npu_inst_pe_1_1_5_U108 ( .A1(npu_inst_pe_1_1_5_n4), .A2(
        npu_inst_pe_1_1_5_n7), .A3(npu_inst_pe_1_1_5_n8), .ZN(
        npu_inst_pe_1_1_5_n40) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_1_5_n34), .CK(
        npu_inst_pe_1_1_5_net3994), .RN(npu_inst_pe_1_1_5_n9), .Q(
        npu_inst_pe_1_1_5_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_1_5_n35), .CK(
        npu_inst_pe_1_1_5_net3994), .RN(npu_inst_pe_1_1_5_n9), .Q(
        npu_inst_pe_1_1_5_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_1_5_n36), .CK(
        npu_inst_pe_1_1_5_net3994), .RN(npu_inst_pe_1_1_5_n9), .Q(
        npu_inst_pe_1_1_5_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_1_5_n98), .CK(
        npu_inst_pe_1_1_5_net3994), .RN(npu_inst_pe_1_1_5_n9), .Q(
        npu_inst_pe_1_1_5_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_1_5_n99), .CK(
        npu_inst_pe_1_1_5_net3994), .RN(npu_inst_pe_1_1_5_n9), .Q(
        npu_inst_pe_1_1_5_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_1_5_n100), 
        .CK(npu_inst_pe_1_1_5_net3994), .RN(npu_inst_pe_1_1_5_n9), .Q(
        npu_inst_pe_1_1_5_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_1_5_n33), .CK(
        npu_inst_pe_1_1_5_net3994), .RN(npu_inst_pe_1_1_5_n9), .Q(
        npu_inst_pe_1_1_5_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_1_5_n101), 
        .CK(npu_inst_pe_1_1_5_net3994), .RN(npu_inst_pe_1_1_5_n9), .Q(
        npu_inst_pe_1_1_5_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_weight_reg_0_ ( .D(npu_inst_n112), .CK(
        npu_inst_pe_1_1_5_net4000), .RN(npu_inst_pe_1_1_5_n9), .Q(
        npu_inst_pe_1_1_5_int_q_weight_0_), .QN(npu_inst_pe_1_1_5_n27) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_weight_reg_1_ ( .D(npu_inst_n118), .CK(
        npu_inst_pe_1_1_5_net4000), .RN(npu_inst_pe_1_1_5_n9), .Q(
        npu_inst_pe_1_1_5_int_q_weight_1_), .QN(npu_inst_pe_1_1_5_n26) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_1_5_n113), 
        .CK(npu_inst_pe_1_1_5_net4000), .RN(npu_inst_pe_1_1_5_n9), .Q(
        npu_inst_pe_1_1_5_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_1_5_n107), 
        .CK(npu_inst_pe_1_1_5_net4000), .RN(npu_inst_pe_1_1_5_n9), .Q(
        npu_inst_pe_1_1_5_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_1_5_n112), 
        .CK(npu_inst_pe_1_1_5_net4000), .RN(npu_inst_pe_1_1_5_n10), .Q(
        npu_inst_pe_1_1_5_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_1_5_n106), 
        .CK(npu_inst_pe_1_1_5_net4000), .RN(npu_inst_pe_1_1_5_n10), .Q(
        npu_inst_pe_1_1_5_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_1_5_n111), 
        .CK(npu_inst_pe_1_1_5_net4000), .RN(npu_inst_pe_1_1_5_n10), .Q(
        npu_inst_pe_1_1_5_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_1_5_n105), 
        .CK(npu_inst_pe_1_1_5_net4000), .RN(npu_inst_pe_1_1_5_n10), .Q(
        npu_inst_pe_1_1_5_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_1_5_n110), 
        .CK(npu_inst_pe_1_1_5_net4000), .RN(npu_inst_pe_1_1_5_n10), .Q(
        npu_inst_pe_1_1_5_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_1_5_n104), 
        .CK(npu_inst_pe_1_1_5_net4000), .RN(npu_inst_pe_1_1_5_n10), .Q(
        npu_inst_pe_1_1_5_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_1_5_n109), 
        .CK(npu_inst_pe_1_1_5_net4000), .RN(npu_inst_pe_1_1_5_n10), .Q(
        npu_inst_pe_1_1_5_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_1_5_n103), 
        .CK(npu_inst_pe_1_1_5_net4000), .RN(npu_inst_pe_1_1_5_n10), .Q(
        npu_inst_pe_1_1_5_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_1_5_n108), 
        .CK(npu_inst_pe_1_1_5_net4000), .RN(npu_inst_pe_1_1_5_n10), .Q(
        npu_inst_pe_1_1_5_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_1_5_n102), 
        .CK(npu_inst_pe_1_1_5_net4000), .RN(npu_inst_pe_1_1_5_n10), .Q(
        npu_inst_pe_1_1_5_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_1_5_n86), 
        .CK(npu_inst_pe_1_1_5_net4000), .RN(npu_inst_pe_1_1_5_n10), .Q(
        npu_inst_pe_1_1_5_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_1_5_n87), 
        .CK(npu_inst_pe_1_1_5_net4000), .RN(npu_inst_pe_1_1_5_n10), .Q(
        npu_inst_pe_1_1_5_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_1_5_n88), 
        .CK(npu_inst_pe_1_1_5_net4000), .RN(npu_inst_pe_1_1_5_n11), .Q(
        npu_inst_pe_1_1_5_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_1_5_n89), 
        .CK(npu_inst_pe_1_1_5_net4000), .RN(npu_inst_pe_1_1_5_n11), .Q(
        npu_inst_pe_1_1_5_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_1_5_n90), 
        .CK(npu_inst_pe_1_1_5_net4000), .RN(npu_inst_pe_1_1_5_n11), .Q(
        npu_inst_pe_1_1_5_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_1_5_n91), 
        .CK(npu_inst_pe_1_1_5_net4000), .RN(npu_inst_pe_1_1_5_n11), .Q(
        npu_inst_pe_1_1_5_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_1_5_n92), 
        .CK(npu_inst_pe_1_1_5_net4000), .RN(npu_inst_pe_1_1_5_n11), .Q(
        npu_inst_pe_1_1_5_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_1_5_n93), 
        .CK(npu_inst_pe_1_1_5_net4000), .RN(npu_inst_pe_1_1_5_n11), .Q(
        npu_inst_pe_1_1_5_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_1_5_n94), 
        .CK(npu_inst_pe_1_1_5_net4000), .RN(npu_inst_pe_1_1_5_n11), .Q(
        npu_inst_pe_1_1_5_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_1_5_n95), 
        .CK(npu_inst_pe_1_1_5_net4000), .RN(npu_inst_pe_1_1_5_n11), .Q(
        npu_inst_pe_1_1_5_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_1_5_n96), 
        .CK(npu_inst_pe_1_1_5_net4000), .RN(npu_inst_pe_1_1_5_n11), .Q(
        npu_inst_pe_1_1_5_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_1_5_n97), 
        .CK(npu_inst_pe_1_1_5_net4000), .RN(npu_inst_pe_1_1_5_n11), .Q(
        npu_inst_pe_1_1_5_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_1_5_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_1_5_N84), .SE(1'b0), .GCK(npu_inst_pe_1_1_5_net3994) );
  CLKGATETST_X1 npu_inst_pe_1_1_5_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n65), .SE(1'b0), .GCK(npu_inst_pe_1_1_5_net4000) );
  MUX2_X1 npu_inst_pe_1_1_6_U162 ( .A(npu_inst_pe_1_1_6_n32), .B(
        npu_inst_pe_1_1_6_n29), .S(npu_inst_pe_1_1_6_n8), .Z(
        npu_inst_pe_1_1_6_N93) );
  MUX2_X1 npu_inst_pe_1_1_6_U161 ( .A(npu_inst_pe_1_1_6_n31), .B(
        npu_inst_pe_1_1_6_n30), .S(npu_inst_pe_1_1_6_n6), .Z(
        npu_inst_pe_1_1_6_n32) );
  MUX2_X1 npu_inst_pe_1_1_6_U160 ( .A(npu_inst_pe_1_1_6_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_1_6_int_q_reg_v_1__0_), .S(npu_inst_pe_1_1_6_n4), .Z(
        npu_inst_pe_1_1_6_n31) );
  MUX2_X1 npu_inst_pe_1_1_6_U159 ( .A(npu_inst_pe_1_1_6_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_1_6_int_q_reg_v_3__0_), .S(npu_inst_pe_1_1_6_n4), .Z(
        npu_inst_pe_1_1_6_n30) );
  MUX2_X1 npu_inst_pe_1_1_6_U158 ( .A(npu_inst_pe_1_1_6_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_1_6_int_q_reg_v_5__0_), .S(npu_inst_pe_1_1_6_n4), .Z(
        npu_inst_pe_1_1_6_n29) );
  MUX2_X1 npu_inst_pe_1_1_6_U157 ( .A(npu_inst_pe_1_1_6_n28), .B(
        npu_inst_pe_1_1_6_n23), .S(npu_inst_pe_1_1_6_n8), .Z(
        npu_inst_pe_1_1_6_N94) );
  MUX2_X1 npu_inst_pe_1_1_6_U156 ( .A(npu_inst_pe_1_1_6_n25), .B(
        npu_inst_pe_1_1_6_n24), .S(npu_inst_pe_1_1_6_n6), .Z(
        npu_inst_pe_1_1_6_n28) );
  MUX2_X1 npu_inst_pe_1_1_6_U155 ( .A(npu_inst_pe_1_1_6_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_1_6_int_q_reg_v_1__1_), .S(npu_inst_pe_1_1_6_n4), .Z(
        npu_inst_pe_1_1_6_n25) );
  MUX2_X1 npu_inst_pe_1_1_6_U154 ( .A(npu_inst_pe_1_1_6_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_1_6_int_q_reg_v_3__1_), .S(npu_inst_pe_1_1_6_n4), .Z(
        npu_inst_pe_1_1_6_n24) );
  MUX2_X1 npu_inst_pe_1_1_6_U153 ( .A(npu_inst_pe_1_1_6_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_1_6_int_q_reg_v_5__1_), .S(npu_inst_pe_1_1_6_n4), .Z(
        npu_inst_pe_1_1_6_n23) );
  MUX2_X1 npu_inst_pe_1_1_6_U152 ( .A(npu_inst_pe_1_1_6_n22), .B(
        npu_inst_pe_1_1_6_n19), .S(npu_inst_pe_1_1_6_n8), .Z(
        npu_inst_int_data_x_1__6__1_) );
  MUX2_X1 npu_inst_pe_1_1_6_U151 ( .A(npu_inst_pe_1_1_6_n21), .B(
        npu_inst_pe_1_1_6_n20), .S(npu_inst_pe_1_1_6_n6), .Z(
        npu_inst_pe_1_1_6_n22) );
  MUX2_X1 npu_inst_pe_1_1_6_U150 ( .A(npu_inst_pe_1_1_6_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_1_6_int_q_reg_h_1__1_), .S(npu_inst_pe_1_1_6_n4), .Z(
        npu_inst_pe_1_1_6_n21) );
  MUX2_X1 npu_inst_pe_1_1_6_U149 ( .A(npu_inst_pe_1_1_6_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_1_6_int_q_reg_h_3__1_), .S(npu_inst_pe_1_1_6_n4), .Z(
        npu_inst_pe_1_1_6_n20) );
  MUX2_X1 npu_inst_pe_1_1_6_U148 ( .A(npu_inst_pe_1_1_6_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_1_6_int_q_reg_h_5__1_), .S(npu_inst_pe_1_1_6_n4), .Z(
        npu_inst_pe_1_1_6_n19) );
  MUX2_X1 npu_inst_pe_1_1_6_U147 ( .A(npu_inst_pe_1_1_6_n18), .B(
        npu_inst_pe_1_1_6_n15), .S(npu_inst_pe_1_1_6_n8), .Z(
        npu_inst_int_data_x_1__6__0_) );
  MUX2_X1 npu_inst_pe_1_1_6_U146 ( .A(npu_inst_pe_1_1_6_n17), .B(
        npu_inst_pe_1_1_6_n16), .S(npu_inst_pe_1_1_6_n6), .Z(
        npu_inst_pe_1_1_6_n18) );
  MUX2_X1 npu_inst_pe_1_1_6_U145 ( .A(npu_inst_pe_1_1_6_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_1_6_int_q_reg_h_1__0_), .S(npu_inst_pe_1_1_6_n4), .Z(
        npu_inst_pe_1_1_6_n17) );
  MUX2_X1 npu_inst_pe_1_1_6_U144 ( .A(npu_inst_pe_1_1_6_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_1_6_int_q_reg_h_3__0_), .S(npu_inst_pe_1_1_6_n4), .Z(
        npu_inst_pe_1_1_6_n16) );
  MUX2_X1 npu_inst_pe_1_1_6_U143 ( .A(npu_inst_pe_1_1_6_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_1_6_int_q_reg_h_5__0_), .S(npu_inst_pe_1_1_6_n4), .Z(
        npu_inst_pe_1_1_6_n15) );
  XOR2_X1 npu_inst_pe_1_1_6_U142 ( .A(npu_inst_pe_1_1_6_int_data_0_), .B(
        npu_inst_pe_1_1_6_int_q_acc_0_), .Z(npu_inst_pe_1_1_6_N73) );
  AND2_X1 npu_inst_pe_1_1_6_U141 ( .A1(npu_inst_pe_1_1_6_int_q_acc_0_), .A2(
        npu_inst_pe_1_1_6_int_data_0_), .ZN(npu_inst_pe_1_1_6_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_1_6_U140 ( .A(npu_inst_pe_1_1_6_int_q_acc_0_), .B(
        npu_inst_pe_1_1_6_n13), .ZN(npu_inst_pe_1_1_6_N65) );
  OR2_X1 npu_inst_pe_1_1_6_U139 ( .A1(npu_inst_pe_1_1_6_n13), .A2(
        npu_inst_pe_1_1_6_int_q_acc_0_), .ZN(npu_inst_pe_1_1_6_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_1_6_U138 ( .A(npu_inst_pe_1_1_6_int_q_acc_2_), .B(
        npu_inst_pe_1_1_6_add_79_carry_2_), .Z(npu_inst_pe_1_1_6_N75) );
  AND2_X1 npu_inst_pe_1_1_6_U137 ( .A1(npu_inst_pe_1_1_6_add_79_carry_2_), 
        .A2(npu_inst_pe_1_1_6_int_q_acc_2_), .ZN(
        npu_inst_pe_1_1_6_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_1_6_U136 ( .A(npu_inst_pe_1_1_6_int_q_acc_3_), .B(
        npu_inst_pe_1_1_6_add_79_carry_3_), .Z(npu_inst_pe_1_1_6_N76) );
  AND2_X1 npu_inst_pe_1_1_6_U135 ( .A1(npu_inst_pe_1_1_6_add_79_carry_3_), 
        .A2(npu_inst_pe_1_1_6_int_q_acc_3_), .ZN(
        npu_inst_pe_1_1_6_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_1_6_U134 ( .A(npu_inst_pe_1_1_6_int_q_acc_4_), .B(
        npu_inst_pe_1_1_6_add_79_carry_4_), .Z(npu_inst_pe_1_1_6_N77) );
  AND2_X1 npu_inst_pe_1_1_6_U133 ( .A1(npu_inst_pe_1_1_6_add_79_carry_4_), 
        .A2(npu_inst_pe_1_1_6_int_q_acc_4_), .ZN(
        npu_inst_pe_1_1_6_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_1_6_U132 ( .A(npu_inst_pe_1_1_6_int_q_acc_5_), .B(
        npu_inst_pe_1_1_6_add_79_carry_5_), .Z(npu_inst_pe_1_1_6_N78) );
  AND2_X1 npu_inst_pe_1_1_6_U131 ( .A1(npu_inst_pe_1_1_6_add_79_carry_5_), 
        .A2(npu_inst_pe_1_1_6_int_q_acc_5_), .ZN(
        npu_inst_pe_1_1_6_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_1_6_U130 ( .A(npu_inst_pe_1_1_6_int_q_acc_6_), .B(
        npu_inst_pe_1_1_6_add_79_carry_6_), .Z(npu_inst_pe_1_1_6_N79) );
  AND2_X1 npu_inst_pe_1_1_6_U129 ( .A1(npu_inst_pe_1_1_6_add_79_carry_6_), 
        .A2(npu_inst_pe_1_1_6_int_q_acc_6_), .ZN(
        npu_inst_pe_1_1_6_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_1_6_U128 ( .A(npu_inst_pe_1_1_6_int_q_acc_7_), .B(
        npu_inst_pe_1_1_6_add_79_carry_7_), .Z(npu_inst_pe_1_1_6_N80) );
  XNOR2_X1 npu_inst_pe_1_1_6_U127 ( .A(npu_inst_pe_1_1_6_sub_77_carry_2_), .B(
        npu_inst_pe_1_1_6_int_q_acc_2_), .ZN(npu_inst_pe_1_1_6_N67) );
  OR2_X1 npu_inst_pe_1_1_6_U126 ( .A1(npu_inst_pe_1_1_6_int_q_acc_2_), .A2(
        npu_inst_pe_1_1_6_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_1_6_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_1_6_U125 ( .A(npu_inst_pe_1_1_6_sub_77_carry_3_), .B(
        npu_inst_pe_1_1_6_int_q_acc_3_), .ZN(npu_inst_pe_1_1_6_N68) );
  OR2_X1 npu_inst_pe_1_1_6_U124 ( .A1(npu_inst_pe_1_1_6_int_q_acc_3_), .A2(
        npu_inst_pe_1_1_6_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_1_6_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_1_6_U123 ( .A(npu_inst_pe_1_1_6_sub_77_carry_4_), .B(
        npu_inst_pe_1_1_6_int_q_acc_4_), .ZN(npu_inst_pe_1_1_6_N69) );
  OR2_X1 npu_inst_pe_1_1_6_U122 ( .A1(npu_inst_pe_1_1_6_int_q_acc_4_), .A2(
        npu_inst_pe_1_1_6_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_1_6_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_1_6_U121 ( .A(npu_inst_pe_1_1_6_sub_77_carry_5_), .B(
        npu_inst_pe_1_1_6_int_q_acc_5_), .ZN(npu_inst_pe_1_1_6_N70) );
  OR2_X1 npu_inst_pe_1_1_6_U120 ( .A1(npu_inst_pe_1_1_6_int_q_acc_5_), .A2(
        npu_inst_pe_1_1_6_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_1_6_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_1_6_U119 ( .A(npu_inst_pe_1_1_6_sub_77_carry_6_), .B(
        npu_inst_pe_1_1_6_int_q_acc_6_), .ZN(npu_inst_pe_1_1_6_N71) );
  OR2_X1 npu_inst_pe_1_1_6_U118 ( .A1(npu_inst_pe_1_1_6_int_q_acc_6_), .A2(
        npu_inst_pe_1_1_6_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_1_6_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_1_6_U117 ( .A(npu_inst_pe_1_1_6_int_q_acc_7_), .B(
        npu_inst_pe_1_1_6_sub_77_carry_7_), .ZN(npu_inst_pe_1_1_6_N72) );
  INV_X1 npu_inst_pe_1_1_6_U116 ( .A(npu_inst_n79), .ZN(npu_inst_pe_1_1_6_n7)
         );
  INV_X1 npu_inst_pe_1_1_6_U115 ( .A(npu_inst_pe_1_1_6_n7), .ZN(
        npu_inst_pe_1_1_6_n6) );
  INV_X1 npu_inst_pe_1_1_6_U114 ( .A(npu_inst_n59), .ZN(npu_inst_pe_1_1_6_n3)
         );
  AOI22_X1 npu_inst_pe_1_1_6_U113 ( .A1(npu_inst_int_data_y_2__6__0_), .A2(
        npu_inst_pe_1_1_6_n58), .B1(npu_inst_pe_1_1_6_n114), .B2(
        npu_inst_pe_1_1_6_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_1_6_n57) );
  INV_X1 npu_inst_pe_1_1_6_U112 ( .A(npu_inst_pe_1_1_6_n57), .ZN(
        npu_inst_pe_1_1_6_n108) );
  AOI22_X1 npu_inst_pe_1_1_6_U111 ( .A1(npu_inst_int_data_y_2__6__0_), .A2(
        npu_inst_pe_1_1_6_n54), .B1(npu_inst_pe_1_1_6_n115), .B2(
        npu_inst_pe_1_1_6_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_1_6_n53) );
  INV_X1 npu_inst_pe_1_1_6_U110 ( .A(npu_inst_pe_1_1_6_n53), .ZN(
        npu_inst_pe_1_1_6_n109) );
  AOI22_X1 npu_inst_pe_1_1_6_U107 ( .A1(npu_inst_int_data_y_2__6__0_), .A2(
        npu_inst_pe_1_1_6_n50), .B1(npu_inst_pe_1_1_6_n116), .B2(
        npu_inst_pe_1_1_6_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_1_6_n49) );
  INV_X1 npu_inst_pe_1_1_6_U106 ( .A(npu_inst_pe_1_1_6_n49), .ZN(
        npu_inst_pe_1_1_6_n110) );
  AOI22_X1 npu_inst_pe_1_1_6_U105 ( .A1(npu_inst_int_data_y_2__6__0_), .A2(
        npu_inst_pe_1_1_6_n46), .B1(npu_inst_pe_1_1_6_n117), .B2(
        npu_inst_pe_1_1_6_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_1_6_n45) );
  INV_X1 npu_inst_pe_1_1_6_U104 ( .A(npu_inst_pe_1_1_6_n45), .ZN(
        npu_inst_pe_1_1_6_n111) );
  AOI22_X1 npu_inst_pe_1_1_6_U103 ( .A1(npu_inst_int_data_y_2__6__0_), .A2(
        npu_inst_pe_1_1_6_n42), .B1(npu_inst_pe_1_1_6_n119), .B2(
        npu_inst_pe_1_1_6_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_1_6_n41) );
  INV_X1 npu_inst_pe_1_1_6_U102 ( .A(npu_inst_pe_1_1_6_n41), .ZN(
        npu_inst_pe_1_1_6_n112) );
  AOI22_X1 npu_inst_pe_1_1_6_U101 ( .A1(npu_inst_int_data_y_2__6__1_), .A2(
        npu_inst_pe_1_1_6_n58), .B1(npu_inst_pe_1_1_6_n114), .B2(
        npu_inst_pe_1_1_6_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_1_6_n59) );
  INV_X1 npu_inst_pe_1_1_6_U100 ( .A(npu_inst_pe_1_1_6_n59), .ZN(
        npu_inst_pe_1_1_6_n102) );
  AOI22_X1 npu_inst_pe_1_1_6_U99 ( .A1(npu_inst_int_data_y_2__6__1_), .A2(
        npu_inst_pe_1_1_6_n54), .B1(npu_inst_pe_1_1_6_n115), .B2(
        npu_inst_pe_1_1_6_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_1_6_n55) );
  INV_X1 npu_inst_pe_1_1_6_U98 ( .A(npu_inst_pe_1_1_6_n55), .ZN(
        npu_inst_pe_1_1_6_n103) );
  AOI22_X1 npu_inst_pe_1_1_6_U97 ( .A1(npu_inst_int_data_y_2__6__1_), .A2(
        npu_inst_pe_1_1_6_n50), .B1(npu_inst_pe_1_1_6_n116), .B2(
        npu_inst_pe_1_1_6_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_1_6_n51) );
  INV_X1 npu_inst_pe_1_1_6_U96 ( .A(npu_inst_pe_1_1_6_n51), .ZN(
        npu_inst_pe_1_1_6_n104) );
  AOI22_X1 npu_inst_pe_1_1_6_U95 ( .A1(npu_inst_int_data_y_2__6__1_), .A2(
        npu_inst_pe_1_1_6_n46), .B1(npu_inst_pe_1_1_6_n117), .B2(
        npu_inst_pe_1_1_6_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_1_6_n47) );
  INV_X1 npu_inst_pe_1_1_6_U94 ( .A(npu_inst_pe_1_1_6_n47), .ZN(
        npu_inst_pe_1_1_6_n105) );
  AOI22_X1 npu_inst_pe_1_1_6_U93 ( .A1(npu_inst_int_data_y_2__6__1_), .A2(
        npu_inst_pe_1_1_6_n42), .B1(npu_inst_pe_1_1_6_n119), .B2(
        npu_inst_pe_1_1_6_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_1_6_n43) );
  INV_X1 npu_inst_pe_1_1_6_U92 ( .A(npu_inst_pe_1_1_6_n43), .ZN(
        npu_inst_pe_1_1_6_n106) );
  AOI22_X1 npu_inst_pe_1_1_6_U91 ( .A1(npu_inst_pe_1_1_6_n38), .A2(
        npu_inst_int_data_y_2__6__1_), .B1(npu_inst_pe_1_1_6_n118), .B2(
        npu_inst_pe_1_1_6_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_1_6_n39) );
  INV_X1 npu_inst_pe_1_1_6_U90 ( .A(npu_inst_pe_1_1_6_n39), .ZN(
        npu_inst_pe_1_1_6_n107) );
  AOI22_X1 npu_inst_pe_1_1_6_U89 ( .A1(npu_inst_pe_1_1_6_n38), .A2(
        npu_inst_int_data_y_2__6__0_), .B1(npu_inst_pe_1_1_6_n118), .B2(
        npu_inst_pe_1_1_6_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_1_6_n37) );
  INV_X1 npu_inst_pe_1_1_6_U88 ( .A(npu_inst_pe_1_1_6_n37), .ZN(
        npu_inst_pe_1_1_6_n113) );
  NAND2_X1 npu_inst_pe_1_1_6_U87 ( .A1(npu_inst_pe_1_1_6_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_1_6_n60), .ZN(npu_inst_pe_1_1_6_n74) );
  OAI21_X1 npu_inst_pe_1_1_6_U86 ( .B1(npu_inst_pe_1_1_6_n63), .B2(
        npu_inst_pe_1_1_6_n60), .A(npu_inst_pe_1_1_6_n74), .ZN(
        npu_inst_pe_1_1_6_n97) );
  NAND2_X1 npu_inst_pe_1_1_6_U85 ( .A1(npu_inst_pe_1_1_6_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_1_6_n60), .ZN(npu_inst_pe_1_1_6_n73) );
  OAI21_X1 npu_inst_pe_1_1_6_U84 ( .B1(npu_inst_pe_1_1_6_n61), .B2(
        npu_inst_pe_1_1_6_n60), .A(npu_inst_pe_1_1_6_n73), .ZN(
        npu_inst_pe_1_1_6_n96) );
  NAND2_X1 npu_inst_pe_1_1_6_U83 ( .A1(npu_inst_pe_1_1_6_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_1_6_n56), .ZN(npu_inst_pe_1_1_6_n72) );
  OAI21_X1 npu_inst_pe_1_1_6_U82 ( .B1(npu_inst_pe_1_1_6_n63), .B2(
        npu_inst_pe_1_1_6_n56), .A(npu_inst_pe_1_1_6_n72), .ZN(
        npu_inst_pe_1_1_6_n95) );
  NAND2_X1 npu_inst_pe_1_1_6_U81 ( .A1(npu_inst_pe_1_1_6_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_1_6_n56), .ZN(npu_inst_pe_1_1_6_n71) );
  OAI21_X1 npu_inst_pe_1_1_6_U80 ( .B1(npu_inst_pe_1_1_6_n61), .B2(
        npu_inst_pe_1_1_6_n56), .A(npu_inst_pe_1_1_6_n71), .ZN(
        npu_inst_pe_1_1_6_n94) );
  NAND2_X1 npu_inst_pe_1_1_6_U79 ( .A1(npu_inst_pe_1_1_6_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_1_6_n52), .ZN(npu_inst_pe_1_1_6_n70) );
  OAI21_X1 npu_inst_pe_1_1_6_U78 ( .B1(npu_inst_pe_1_1_6_n63), .B2(
        npu_inst_pe_1_1_6_n52), .A(npu_inst_pe_1_1_6_n70), .ZN(
        npu_inst_pe_1_1_6_n93) );
  NAND2_X1 npu_inst_pe_1_1_6_U77 ( .A1(npu_inst_pe_1_1_6_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_1_6_n52), .ZN(npu_inst_pe_1_1_6_n69) );
  OAI21_X1 npu_inst_pe_1_1_6_U76 ( .B1(npu_inst_pe_1_1_6_n61), .B2(
        npu_inst_pe_1_1_6_n52), .A(npu_inst_pe_1_1_6_n69), .ZN(
        npu_inst_pe_1_1_6_n92) );
  NAND2_X1 npu_inst_pe_1_1_6_U75 ( .A1(npu_inst_pe_1_1_6_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_1_6_n48), .ZN(npu_inst_pe_1_1_6_n68) );
  OAI21_X1 npu_inst_pe_1_1_6_U74 ( .B1(npu_inst_pe_1_1_6_n63), .B2(
        npu_inst_pe_1_1_6_n48), .A(npu_inst_pe_1_1_6_n68), .ZN(
        npu_inst_pe_1_1_6_n91) );
  NAND2_X1 npu_inst_pe_1_1_6_U73 ( .A1(npu_inst_pe_1_1_6_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_1_6_n48), .ZN(npu_inst_pe_1_1_6_n67) );
  OAI21_X1 npu_inst_pe_1_1_6_U72 ( .B1(npu_inst_pe_1_1_6_n61), .B2(
        npu_inst_pe_1_1_6_n48), .A(npu_inst_pe_1_1_6_n67), .ZN(
        npu_inst_pe_1_1_6_n90) );
  NAND2_X1 npu_inst_pe_1_1_6_U71 ( .A1(npu_inst_pe_1_1_6_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_1_6_n44), .ZN(npu_inst_pe_1_1_6_n66) );
  OAI21_X1 npu_inst_pe_1_1_6_U70 ( .B1(npu_inst_pe_1_1_6_n63), .B2(
        npu_inst_pe_1_1_6_n44), .A(npu_inst_pe_1_1_6_n66), .ZN(
        npu_inst_pe_1_1_6_n89) );
  NAND2_X1 npu_inst_pe_1_1_6_U69 ( .A1(npu_inst_pe_1_1_6_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_1_6_n44), .ZN(npu_inst_pe_1_1_6_n65) );
  OAI21_X1 npu_inst_pe_1_1_6_U68 ( .B1(npu_inst_pe_1_1_6_n61), .B2(
        npu_inst_pe_1_1_6_n44), .A(npu_inst_pe_1_1_6_n65), .ZN(
        npu_inst_pe_1_1_6_n88) );
  NAND2_X1 npu_inst_pe_1_1_6_U67 ( .A1(npu_inst_pe_1_1_6_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_1_6_n40), .ZN(npu_inst_pe_1_1_6_n64) );
  OAI21_X1 npu_inst_pe_1_1_6_U66 ( .B1(npu_inst_pe_1_1_6_n63), .B2(
        npu_inst_pe_1_1_6_n40), .A(npu_inst_pe_1_1_6_n64), .ZN(
        npu_inst_pe_1_1_6_n87) );
  NAND2_X1 npu_inst_pe_1_1_6_U65 ( .A1(npu_inst_pe_1_1_6_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_1_6_n40), .ZN(npu_inst_pe_1_1_6_n62) );
  OAI21_X1 npu_inst_pe_1_1_6_U64 ( .B1(npu_inst_pe_1_1_6_n61), .B2(
        npu_inst_pe_1_1_6_n40), .A(npu_inst_pe_1_1_6_n62), .ZN(
        npu_inst_pe_1_1_6_n86) );
  AND2_X1 npu_inst_pe_1_1_6_U63 ( .A1(npu_inst_pe_1_1_6_N93), .A2(npu_inst_n59), .ZN(npu_inst_int_data_y_1__6__0_) );
  AND2_X1 npu_inst_pe_1_1_6_U62 ( .A1(npu_inst_n59), .A2(npu_inst_pe_1_1_6_N94), .ZN(npu_inst_int_data_y_1__6__1_) );
  NOR3_X1 npu_inst_pe_1_1_6_U61 ( .A1(npu_inst_pe_1_1_6_n26), .A2(npu_inst_n59), .A3(npu_inst_int_ckg[49]), .ZN(npu_inst_pe_1_1_6_n85) );
  OR2_X1 npu_inst_pe_1_1_6_U60 ( .A1(npu_inst_pe_1_1_6_n85), .A2(
        npu_inst_pe_1_1_6_n2), .ZN(npu_inst_pe_1_1_6_N84) );
  AND2_X1 npu_inst_pe_1_1_6_U59 ( .A1(npu_inst_pe_1_1_6_int_q_acc_0_), .A2(
        npu_inst_pe_1_1_6_n1), .ZN(npu_inst_int_data_res_1__6__0_) );
  AND2_X1 npu_inst_pe_1_1_6_U58 ( .A1(npu_inst_pe_1_1_6_n2), .A2(
        npu_inst_pe_1_1_6_int_q_acc_7_), .ZN(npu_inst_int_data_res_1__6__7_)
         );
  AND2_X1 npu_inst_pe_1_1_6_U57 ( .A1(npu_inst_pe_1_1_6_int_q_acc_1_), .A2(
        npu_inst_pe_1_1_6_n1), .ZN(npu_inst_int_data_res_1__6__1_) );
  AND2_X1 npu_inst_pe_1_1_6_U56 ( .A1(npu_inst_pe_1_1_6_int_q_acc_2_), .A2(
        npu_inst_pe_1_1_6_n1), .ZN(npu_inst_int_data_res_1__6__2_) );
  AND2_X1 npu_inst_pe_1_1_6_U55 ( .A1(npu_inst_pe_1_1_6_int_q_acc_3_), .A2(
        npu_inst_pe_1_1_6_n2), .ZN(npu_inst_int_data_res_1__6__3_) );
  AND2_X1 npu_inst_pe_1_1_6_U54 ( .A1(npu_inst_pe_1_1_6_int_q_acc_4_), .A2(
        npu_inst_pe_1_1_6_n2), .ZN(npu_inst_int_data_res_1__6__4_) );
  AND2_X1 npu_inst_pe_1_1_6_U53 ( .A1(npu_inst_pe_1_1_6_int_q_acc_5_), .A2(
        npu_inst_pe_1_1_6_n2), .ZN(npu_inst_int_data_res_1__6__5_) );
  AND2_X1 npu_inst_pe_1_1_6_U52 ( .A1(npu_inst_pe_1_1_6_int_q_acc_6_), .A2(
        npu_inst_pe_1_1_6_n2), .ZN(npu_inst_int_data_res_1__6__6_) );
  AOI222_X1 npu_inst_pe_1_1_6_U51 ( .A1(npu_inst_int_data_res_2__6__0_), .A2(
        npu_inst_pe_1_1_6_n1), .B1(npu_inst_pe_1_1_6_N73), .B2(
        npu_inst_pe_1_1_6_n76), .C1(npu_inst_pe_1_1_6_N65), .C2(
        npu_inst_pe_1_1_6_n77), .ZN(npu_inst_pe_1_1_6_n84) );
  INV_X1 npu_inst_pe_1_1_6_U50 ( .A(npu_inst_pe_1_1_6_n84), .ZN(
        npu_inst_pe_1_1_6_n101) );
  AOI222_X1 npu_inst_pe_1_1_6_U49 ( .A1(npu_inst_int_data_res_2__6__7_), .A2(
        npu_inst_pe_1_1_6_n1), .B1(npu_inst_pe_1_1_6_N80), .B2(
        npu_inst_pe_1_1_6_n76), .C1(npu_inst_pe_1_1_6_N72), .C2(
        npu_inst_pe_1_1_6_n77), .ZN(npu_inst_pe_1_1_6_n75) );
  INV_X1 npu_inst_pe_1_1_6_U48 ( .A(npu_inst_pe_1_1_6_n75), .ZN(
        npu_inst_pe_1_1_6_n33) );
  AOI222_X1 npu_inst_pe_1_1_6_U47 ( .A1(npu_inst_int_data_res_2__6__1_), .A2(
        npu_inst_pe_1_1_6_n1), .B1(npu_inst_pe_1_1_6_N74), .B2(
        npu_inst_pe_1_1_6_n76), .C1(npu_inst_pe_1_1_6_N66), .C2(
        npu_inst_pe_1_1_6_n77), .ZN(npu_inst_pe_1_1_6_n83) );
  INV_X1 npu_inst_pe_1_1_6_U46 ( .A(npu_inst_pe_1_1_6_n83), .ZN(
        npu_inst_pe_1_1_6_n100) );
  AOI222_X1 npu_inst_pe_1_1_6_U45 ( .A1(npu_inst_int_data_res_2__6__2_), .A2(
        npu_inst_pe_1_1_6_n1), .B1(npu_inst_pe_1_1_6_N75), .B2(
        npu_inst_pe_1_1_6_n76), .C1(npu_inst_pe_1_1_6_N67), .C2(
        npu_inst_pe_1_1_6_n77), .ZN(npu_inst_pe_1_1_6_n82) );
  INV_X1 npu_inst_pe_1_1_6_U44 ( .A(npu_inst_pe_1_1_6_n82), .ZN(
        npu_inst_pe_1_1_6_n99) );
  AOI222_X1 npu_inst_pe_1_1_6_U43 ( .A1(npu_inst_int_data_res_2__6__3_), .A2(
        npu_inst_pe_1_1_6_n1), .B1(npu_inst_pe_1_1_6_N76), .B2(
        npu_inst_pe_1_1_6_n76), .C1(npu_inst_pe_1_1_6_N68), .C2(
        npu_inst_pe_1_1_6_n77), .ZN(npu_inst_pe_1_1_6_n81) );
  INV_X1 npu_inst_pe_1_1_6_U42 ( .A(npu_inst_pe_1_1_6_n81), .ZN(
        npu_inst_pe_1_1_6_n98) );
  AOI222_X1 npu_inst_pe_1_1_6_U41 ( .A1(npu_inst_int_data_res_2__6__4_), .A2(
        npu_inst_pe_1_1_6_n1), .B1(npu_inst_pe_1_1_6_N77), .B2(
        npu_inst_pe_1_1_6_n76), .C1(npu_inst_pe_1_1_6_N69), .C2(
        npu_inst_pe_1_1_6_n77), .ZN(npu_inst_pe_1_1_6_n80) );
  INV_X1 npu_inst_pe_1_1_6_U40 ( .A(npu_inst_pe_1_1_6_n80), .ZN(
        npu_inst_pe_1_1_6_n36) );
  AOI222_X1 npu_inst_pe_1_1_6_U39 ( .A1(npu_inst_int_data_res_2__6__5_), .A2(
        npu_inst_pe_1_1_6_n1), .B1(npu_inst_pe_1_1_6_N78), .B2(
        npu_inst_pe_1_1_6_n76), .C1(npu_inst_pe_1_1_6_N70), .C2(
        npu_inst_pe_1_1_6_n77), .ZN(npu_inst_pe_1_1_6_n79) );
  INV_X1 npu_inst_pe_1_1_6_U38 ( .A(npu_inst_pe_1_1_6_n79), .ZN(
        npu_inst_pe_1_1_6_n35) );
  AOI222_X1 npu_inst_pe_1_1_6_U37 ( .A1(npu_inst_int_data_res_2__6__6_), .A2(
        npu_inst_pe_1_1_6_n1), .B1(npu_inst_pe_1_1_6_N79), .B2(
        npu_inst_pe_1_1_6_n76), .C1(npu_inst_pe_1_1_6_N71), .C2(
        npu_inst_pe_1_1_6_n77), .ZN(npu_inst_pe_1_1_6_n78) );
  INV_X1 npu_inst_pe_1_1_6_U36 ( .A(npu_inst_pe_1_1_6_n78), .ZN(
        npu_inst_pe_1_1_6_n34) );
  INV_X1 npu_inst_pe_1_1_6_U35 ( .A(npu_inst_pe_1_1_6_int_data_1_), .ZN(
        npu_inst_pe_1_1_6_n14) );
  AND2_X1 npu_inst_pe_1_1_6_U34 ( .A1(npu_inst_int_data_x_1__6__1_), .A2(
        npu_inst_pe_1_1_6_int_q_weight_1_), .ZN(npu_inst_pe_1_1_6_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_1_6_U33 ( .A1(npu_inst_int_data_x_1__6__0_), .A2(
        npu_inst_pe_1_1_6_int_q_weight_1_), .ZN(npu_inst_pe_1_1_6_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_1_6_U32 ( .A1(npu_inst_n59), .A2(
        npu_inst_int_data_y_2__6__1_), .B1(npu_inst_pe_1_1_6_n3), .B2(
        npu_inst_int_data_x_1__7__1_), .ZN(npu_inst_pe_1_1_6_n63) );
  AOI22_X1 npu_inst_pe_1_1_6_U31 ( .A1(npu_inst_n59), .A2(
        npu_inst_int_data_y_2__6__0_), .B1(npu_inst_pe_1_1_6_n3), .B2(
        npu_inst_int_data_x_1__7__0_), .ZN(npu_inst_pe_1_1_6_n61) );
  INV_X1 npu_inst_pe_1_1_6_U30 ( .A(npu_inst_pe_1_1_6_int_data_0_), .ZN(
        npu_inst_pe_1_1_6_n13) );
  INV_X1 npu_inst_pe_1_1_6_U29 ( .A(npu_inst_n71), .ZN(npu_inst_pe_1_1_6_n5)
         );
  OR3_X1 npu_inst_pe_1_1_6_U28 ( .A1(npu_inst_pe_1_1_6_n6), .A2(
        npu_inst_pe_1_1_6_n8), .A3(npu_inst_pe_1_1_6_n5), .ZN(
        npu_inst_pe_1_1_6_n56) );
  OR3_X1 npu_inst_pe_1_1_6_U27 ( .A1(npu_inst_pe_1_1_6_n5), .A2(
        npu_inst_pe_1_1_6_n8), .A3(npu_inst_pe_1_1_6_n7), .ZN(
        npu_inst_pe_1_1_6_n48) );
  INV_X1 npu_inst_pe_1_1_6_U26 ( .A(npu_inst_pe_1_1_6_n5), .ZN(
        npu_inst_pe_1_1_6_n4) );
  INV_X1 npu_inst_pe_1_1_6_U25 ( .A(npu_inst_n126), .ZN(npu_inst_pe_1_1_6_n12)
         );
  OR3_X1 npu_inst_pe_1_1_6_U24 ( .A1(npu_inst_pe_1_1_6_n4), .A2(
        npu_inst_pe_1_1_6_n8), .A3(npu_inst_pe_1_1_6_n7), .ZN(
        npu_inst_pe_1_1_6_n52) );
  OR3_X1 npu_inst_pe_1_1_6_U23 ( .A1(npu_inst_pe_1_1_6_n6), .A2(
        npu_inst_pe_1_1_6_n8), .A3(npu_inst_pe_1_1_6_n4), .ZN(
        npu_inst_pe_1_1_6_n60) );
  NOR2_X1 npu_inst_pe_1_1_6_U22 ( .A1(npu_inst_pe_1_1_6_n60), .A2(
        npu_inst_pe_1_1_6_n3), .ZN(npu_inst_pe_1_1_6_n58) );
  NOR2_X1 npu_inst_pe_1_1_6_U21 ( .A1(npu_inst_pe_1_1_6_n56), .A2(
        npu_inst_pe_1_1_6_n3), .ZN(npu_inst_pe_1_1_6_n54) );
  NOR2_X1 npu_inst_pe_1_1_6_U20 ( .A1(npu_inst_pe_1_1_6_n52), .A2(
        npu_inst_pe_1_1_6_n3), .ZN(npu_inst_pe_1_1_6_n50) );
  NOR2_X1 npu_inst_pe_1_1_6_U19 ( .A1(npu_inst_pe_1_1_6_n48), .A2(
        npu_inst_pe_1_1_6_n3), .ZN(npu_inst_pe_1_1_6_n46) );
  NOR2_X1 npu_inst_pe_1_1_6_U18 ( .A1(npu_inst_pe_1_1_6_n40), .A2(
        npu_inst_pe_1_1_6_n3), .ZN(npu_inst_pe_1_1_6_n38) );
  NOR2_X1 npu_inst_pe_1_1_6_U17 ( .A1(npu_inst_pe_1_1_6_n44), .A2(
        npu_inst_pe_1_1_6_n3), .ZN(npu_inst_pe_1_1_6_n42) );
  BUF_X1 npu_inst_pe_1_1_6_U16 ( .A(npu_inst_n104), .Z(npu_inst_pe_1_1_6_n8)
         );
  BUF_X1 npu_inst_pe_1_1_6_U15 ( .A(npu_inst_pe_1_1_6_n12), .Z(
        npu_inst_pe_1_1_6_n11) );
  BUF_X1 npu_inst_pe_1_1_6_U14 ( .A(npu_inst_pe_1_1_6_n12), .Z(
        npu_inst_pe_1_1_6_n10) );
  BUF_X1 npu_inst_pe_1_1_6_U13 ( .A(npu_inst_pe_1_1_6_n12), .Z(
        npu_inst_pe_1_1_6_n9) );
  INV_X1 npu_inst_pe_1_1_6_U12 ( .A(npu_inst_pe_1_1_6_n38), .ZN(
        npu_inst_pe_1_1_6_n118) );
  INV_X1 npu_inst_pe_1_1_6_U11 ( .A(npu_inst_pe_1_1_6_n58), .ZN(
        npu_inst_pe_1_1_6_n114) );
  INV_X1 npu_inst_pe_1_1_6_U10 ( .A(npu_inst_pe_1_1_6_n54), .ZN(
        npu_inst_pe_1_1_6_n115) );
  INV_X1 npu_inst_pe_1_1_6_U9 ( .A(npu_inst_pe_1_1_6_n50), .ZN(
        npu_inst_pe_1_1_6_n116) );
  INV_X1 npu_inst_pe_1_1_6_U8 ( .A(npu_inst_pe_1_1_6_n46), .ZN(
        npu_inst_pe_1_1_6_n117) );
  INV_X1 npu_inst_pe_1_1_6_U7 ( .A(npu_inst_pe_1_1_6_n42), .ZN(
        npu_inst_pe_1_1_6_n119) );
  BUF_X1 npu_inst_pe_1_1_6_U6 ( .A(npu_inst_n31), .Z(npu_inst_pe_1_1_6_n2) );
  BUF_X1 npu_inst_pe_1_1_6_U5 ( .A(npu_inst_n31), .Z(npu_inst_pe_1_1_6_n1) );
  NOR2_X1 npu_inst_pe_1_1_6_U4 ( .A1(npu_inst_pe_1_1_6_int_q_weight_0_), .A2(
        npu_inst_pe_1_1_6_n1), .ZN(npu_inst_pe_1_1_6_n76) );
  NOR2_X1 npu_inst_pe_1_1_6_U3 ( .A1(npu_inst_pe_1_1_6_n27), .A2(
        npu_inst_pe_1_1_6_n1), .ZN(npu_inst_pe_1_1_6_n77) );
  FA_X1 npu_inst_pe_1_1_6_sub_77_U2_1 ( .A(npu_inst_pe_1_1_6_int_q_acc_1_), 
        .B(npu_inst_pe_1_1_6_n14), .CI(npu_inst_pe_1_1_6_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_1_6_sub_77_carry_2_), .S(npu_inst_pe_1_1_6_N66) );
  FA_X1 npu_inst_pe_1_1_6_add_79_U1_1 ( .A(npu_inst_pe_1_1_6_int_q_acc_1_), 
        .B(npu_inst_pe_1_1_6_int_data_1_), .CI(
        npu_inst_pe_1_1_6_add_79_carry_1_), .CO(
        npu_inst_pe_1_1_6_add_79_carry_2_), .S(npu_inst_pe_1_1_6_N74) );
  NAND3_X1 npu_inst_pe_1_1_6_U109 ( .A1(npu_inst_pe_1_1_6_n5), .A2(
        npu_inst_pe_1_1_6_n7), .A3(npu_inst_pe_1_1_6_n8), .ZN(
        npu_inst_pe_1_1_6_n44) );
  NAND3_X1 npu_inst_pe_1_1_6_U108 ( .A1(npu_inst_pe_1_1_6_n4), .A2(
        npu_inst_pe_1_1_6_n7), .A3(npu_inst_pe_1_1_6_n8), .ZN(
        npu_inst_pe_1_1_6_n40) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_1_6_n34), .CK(
        npu_inst_pe_1_1_6_net3971), .RN(npu_inst_pe_1_1_6_n9), .Q(
        npu_inst_pe_1_1_6_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_1_6_n35), .CK(
        npu_inst_pe_1_1_6_net3971), .RN(npu_inst_pe_1_1_6_n9), .Q(
        npu_inst_pe_1_1_6_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_1_6_n36), .CK(
        npu_inst_pe_1_1_6_net3971), .RN(npu_inst_pe_1_1_6_n9), .Q(
        npu_inst_pe_1_1_6_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_1_6_n98), .CK(
        npu_inst_pe_1_1_6_net3971), .RN(npu_inst_pe_1_1_6_n9), .Q(
        npu_inst_pe_1_1_6_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_1_6_n99), .CK(
        npu_inst_pe_1_1_6_net3971), .RN(npu_inst_pe_1_1_6_n9), .Q(
        npu_inst_pe_1_1_6_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_1_6_n100), 
        .CK(npu_inst_pe_1_1_6_net3971), .RN(npu_inst_pe_1_1_6_n9), .Q(
        npu_inst_pe_1_1_6_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_1_6_n33), .CK(
        npu_inst_pe_1_1_6_net3971), .RN(npu_inst_pe_1_1_6_n9), .Q(
        npu_inst_pe_1_1_6_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_1_6_n101), 
        .CK(npu_inst_pe_1_1_6_net3971), .RN(npu_inst_pe_1_1_6_n9), .Q(
        npu_inst_pe_1_1_6_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_weight_reg_0_ ( .D(npu_inst_n112), .CK(
        npu_inst_pe_1_1_6_net3977), .RN(npu_inst_pe_1_1_6_n9), .Q(
        npu_inst_pe_1_1_6_int_q_weight_0_), .QN(npu_inst_pe_1_1_6_n27) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_weight_reg_1_ ( .D(npu_inst_n118), .CK(
        npu_inst_pe_1_1_6_net3977), .RN(npu_inst_pe_1_1_6_n9), .Q(
        npu_inst_pe_1_1_6_int_q_weight_1_), .QN(npu_inst_pe_1_1_6_n26) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_1_6_n113), 
        .CK(npu_inst_pe_1_1_6_net3977), .RN(npu_inst_pe_1_1_6_n9), .Q(
        npu_inst_pe_1_1_6_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_1_6_n107), 
        .CK(npu_inst_pe_1_1_6_net3977), .RN(npu_inst_pe_1_1_6_n9), .Q(
        npu_inst_pe_1_1_6_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_1_6_n112), 
        .CK(npu_inst_pe_1_1_6_net3977), .RN(npu_inst_pe_1_1_6_n10), .Q(
        npu_inst_pe_1_1_6_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_1_6_n106), 
        .CK(npu_inst_pe_1_1_6_net3977), .RN(npu_inst_pe_1_1_6_n10), .Q(
        npu_inst_pe_1_1_6_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_1_6_n111), 
        .CK(npu_inst_pe_1_1_6_net3977), .RN(npu_inst_pe_1_1_6_n10), .Q(
        npu_inst_pe_1_1_6_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_1_6_n105), 
        .CK(npu_inst_pe_1_1_6_net3977), .RN(npu_inst_pe_1_1_6_n10), .Q(
        npu_inst_pe_1_1_6_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_1_6_n110), 
        .CK(npu_inst_pe_1_1_6_net3977), .RN(npu_inst_pe_1_1_6_n10), .Q(
        npu_inst_pe_1_1_6_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_1_6_n104), 
        .CK(npu_inst_pe_1_1_6_net3977), .RN(npu_inst_pe_1_1_6_n10), .Q(
        npu_inst_pe_1_1_6_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_1_6_n109), 
        .CK(npu_inst_pe_1_1_6_net3977), .RN(npu_inst_pe_1_1_6_n10), .Q(
        npu_inst_pe_1_1_6_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_1_6_n103), 
        .CK(npu_inst_pe_1_1_6_net3977), .RN(npu_inst_pe_1_1_6_n10), .Q(
        npu_inst_pe_1_1_6_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_1_6_n108), 
        .CK(npu_inst_pe_1_1_6_net3977), .RN(npu_inst_pe_1_1_6_n10), .Q(
        npu_inst_pe_1_1_6_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_1_6_n102), 
        .CK(npu_inst_pe_1_1_6_net3977), .RN(npu_inst_pe_1_1_6_n10), .Q(
        npu_inst_pe_1_1_6_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_1_6_n86), 
        .CK(npu_inst_pe_1_1_6_net3977), .RN(npu_inst_pe_1_1_6_n10), .Q(
        npu_inst_pe_1_1_6_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_1_6_n87), 
        .CK(npu_inst_pe_1_1_6_net3977), .RN(npu_inst_pe_1_1_6_n10), .Q(
        npu_inst_pe_1_1_6_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_1_6_n88), 
        .CK(npu_inst_pe_1_1_6_net3977), .RN(npu_inst_pe_1_1_6_n11), .Q(
        npu_inst_pe_1_1_6_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_1_6_n89), 
        .CK(npu_inst_pe_1_1_6_net3977), .RN(npu_inst_pe_1_1_6_n11), .Q(
        npu_inst_pe_1_1_6_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_1_6_n90), 
        .CK(npu_inst_pe_1_1_6_net3977), .RN(npu_inst_pe_1_1_6_n11), .Q(
        npu_inst_pe_1_1_6_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_1_6_n91), 
        .CK(npu_inst_pe_1_1_6_net3977), .RN(npu_inst_pe_1_1_6_n11), .Q(
        npu_inst_pe_1_1_6_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_1_6_n92), 
        .CK(npu_inst_pe_1_1_6_net3977), .RN(npu_inst_pe_1_1_6_n11), .Q(
        npu_inst_pe_1_1_6_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_1_6_n93), 
        .CK(npu_inst_pe_1_1_6_net3977), .RN(npu_inst_pe_1_1_6_n11), .Q(
        npu_inst_pe_1_1_6_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_1_6_n94), 
        .CK(npu_inst_pe_1_1_6_net3977), .RN(npu_inst_pe_1_1_6_n11), .Q(
        npu_inst_pe_1_1_6_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_1_6_n95), 
        .CK(npu_inst_pe_1_1_6_net3977), .RN(npu_inst_pe_1_1_6_n11), .Q(
        npu_inst_pe_1_1_6_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_1_6_n96), 
        .CK(npu_inst_pe_1_1_6_net3977), .RN(npu_inst_pe_1_1_6_n11), .Q(
        npu_inst_pe_1_1_6_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_1_6_n97), 
        .CK(npu_inst_pe_1_1_6_net3977), .RN(npu_inst_pe_1_1_6_n11), .Q(
        npu_inst_pe_1_1_6_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_1_6_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_1_6_N84), .SE(1'b0), .GCK(npu_inst_pe_1_1_6_net3971) );
  CLKGATETST_X1 npu_inst_pe_1_1_6_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n65), .SE(1'b0), .GCK(npu_inst_pe_1_1_6_net3977) );
  MUX2_X1 npu_inst_pe_1_1_7_U162 ( .A(npu_inst_pe_1_1_7_n32), .B(
        npu_inst_pe_1_1_7_n29), .S(npu_inst_pe_1_1_7_n8), .Z(
        npu_inst_pe_1_1_7_N93) );
  MUX2_X1 npu_inst_pe_1_1_7_U161 ( .A(npu_inst_pe_1_1_7_n31), .B(
        npu_inst_pe_1_1_7_n30), .S(npu_inst_pe_1_1_7_n6), .Z(
        npu_inst_pe_1_1_7_n32) );
  MUX2_X1 npu_inst_pe_1_1_7_U160 ( .A(npu_inst_pe_1_1_7_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_1_7_int_q_reg_v_1__0_), .S(npu_inst_pe_1_1_7_n4), .Z(
        npu_inst_pe_1_1_7_n31) );
  MUX2_X1 npu_inst_pe_1_1_7_U159 ( .A(npu_inst_pe_1_1_7_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_1_7_int_q_reg_v_3__0_), .S(npu_inst_pe_1_1_7_n4), .Z(
        npu_inst_pe_1_1_7_n30) );
  MUX2_X1 npu_inst_pe_1_1_7_U158 ( .A(npu_inst_pe_1_1_7_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_1_7_int_q_reg_v_5__0_), .S(npu_inst_pe_1_1_7_n4), .Z(
        npu_inst_pe_1_1_7_n29) );
  MUX2_X1 npu_inst_pe_1_1_7_U157 ( .A(npu_inst_pe_1_1_7_n28), .B(
        npu_inst_pe_1_1_7_n23), .S(npu_inst_pe_1_1_7_n8), .Z(
        npu_inst_pe_1_1_7_N94) );
  MUX2_X1 npu_inst_pe_1_1_7_U156 ( .A(npu_inst_pe_1_1_7_n25), .B(
        npu_inst_pe_1_1_7_n24), .S(npu_inst_pe_1_1_7_n6), .Z(
        npu_inst_pe_1_1_7_n28) );
  MUX2_X1 npu_inst_pe_1_1_7_U155 ( .A(npu_inst_pe_1_1_7_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_1_7_int_q_reg_v_1__1_), .S(npu_inst_pe_1_1_7_n4), .Z(
        npu_inst_pe_1_1_7_n25) );
  MUX2_X1 npu_inst_pe_1_1_7_U154 ( .A(npu_inst_pe_1_1_7_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_1_7_int_q_reg_v_3__1_), .S(npu_inst_pe_1_1_7_n4), .Z(
        npu_inst_pe_1_1_7_n24) );
  MUX2_X1 npu_inst_pe_1_1_7_U153 ( .A(npu_inst_pe_1_1_7_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_1_7_int_q_reg_v_5__1_), .S(npu_inst_pe_1_1_7_n4), .Z(
        npu_inst_pe_1_1_7_n23) );
  MUX2_X1 npu_inst_pe_1_1_7_U152 ( .A(npu_inst_pe_1_1_7_n22), .B(
        npu_inst_pe_1_1_7_n19), .S(npu_inst_pe_1_1_7_n8), .Z(
        npu_inst_int_data_x_1__7__1_) );
  MUX2_X1 npu_inst_pe_1_1_7_U151 ( .A(npu_inst_pe_1_1_7_n21), .B(
        npu_inst_pe_1_1_7_n20), .S(npu_inst_pe_1_1_7_n6), .Z(
        npu_inst_pe_1_1_7_n22) );
  MUX2_X1 npu_inst_pe_1_1_7_U150 ( .A(npu_inst_pe_1_1_7_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_1_7_int_q_reg_h_1__1_), .S(npu_inst_pe_1_1_7_n4), .Z(
        npu_inst_pe_1_1_7_n21) );
  MUX2_X1 npu_inst_pe_1_1_7_U149 ( .A(npu_inst_pe_1_1_7_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_1_7_int_q_reg_h_3__1_), .S(npu_inst_pe_1_1_7_n4), .Z(
        npu_inst_pe_1_1_7_n20) );
  MUX2_X1 npu_inst_pe_1_1_7_U148 ( .A(npu_inst_pe_1_1_7_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_1_7_int_q_reg_h_5__1_), .S(npu_inst_pe_1_1_7_n4), .Z(
        npu_inst_pe_1_1_7_n19) );
  MUX2_X1 npu_inst_pe_1_1_7_U147 ( .A(npu_inst_pe_1_1_7_n18), .B(
        npu_inst_pe_1_1_7_n15), .S(npu_inst_pe_1_1_7_n8), .Z(
        npu_inst_int_data_x_1__7__0_) );
  MUX2_X1 npu_inst_pe_1_1_7_U146 ( .A(npu_inst_pe_1_1_7_n17), .B(
        npu_inst_pe_1_1_7_n16), .S(npu_inst_pe_1_1_7_n6), .Z(
        npu_inst_pe_1_1_7_n18) );
  MUX2_X1 npu_inst_pe_1_1_7_U145 ( .A(npu_inst_pe_1_1_7_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_1_7_int_q_reg_h_1__0_), .S(npu_inst_pe_1_1_7_n4), .Z(
        npu_inst_pe_1_1_7_n17) );
  MUX2_X1 npu_inst_pe_1_1_7_U144 ( .A(npu_inst_pe_1_1_7_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_1_7_int_q_reg_h_3__0_), .S(npu_inst_pe_1_1_7_n4), .Z(
        npu_inst_pe_1_1_7_n16) );
  MUX2_X1 npu_inst_pe_1_1_7_U143 ( .A(npu_inst_pe_1_1_7_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_1_7_int_q_reg_h_5__0_), .S(npu_inst_pe_1_1_7_n4), .Z(
        npu_inst_pe_1_1_7_n15) );
  XOR2_X1 npu_inst_pe_1_1_7_U142 ( .A(npu_inst_pe_1_1_7_int_data_0_), .B(
        npu_inst_pe_1_1_7_int_q_acc_0_), .Z(npu_inst_pe_1_1_7_N73) );
  AND2_X1 npu_inst_pe_1_1_7_U141 ( .A1(npu_inst_pe_1_1_7_int_q_acc_0_), .A2(
        npu_inst_pe_1_1_7_int_data_0_), .ZN(npu_inst_pe_1_1_7_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_1_7_U140 ( .A(npu_inst_pe_1_1_7_int_q_acc_0_), .B(
        npu_inst_pe_1_1_7_n13), .ZN(npu_inst_pe_1_1_7_N65) );
  OR2_X1 npu_inst_pe_1_1_7_U139 ( .A1(npu_inst_pe_1_1_7_n13), .A2(
        npu_inst_pe_1_1_7_int_q_acc_0_), .ZN(npu_inst_pe_1_1_7_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_1_7_U138 ( .A(npu_inst_pe_1_1_7_int_q_acc_2_), .B(
        npu_inst_pe_1_1_7_add_79_carry_2_), .Z(npu_inst_pe_1_1_7_N75) );
  AND2_X1 npu_inst_pe_1_1_7_U137 ( .A1(npu_inst_pe_1_1_7_add_79_carry_2_), 
        .A2(npu_inst_pe_1_1_7_int_q_acc_2_), .ZN(
        npu_inst_pe_1_1_7_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_1_7_U136 ( .A(npu_inst_pe_1_1_7_int_q_acc_3_), .B(
        npu_inst_pe_1_1_7_add_79_carry_3_), .Z(npu_inst_pe_1_1_7_N76) );
  AND2_X1 npu_inst_pe_1_1_7_U135 ( .A1(npu_inst_pe_1_1_7_add_79_carry_3_), 
        .A2(npu_inst_pe_1_1_7_int_q_acc_3_), .ZN(
        npu_inst_pe_1_1_7_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_1_7_U134 ( .A(npu_inst_pe_1_1_7_int_q_acc_4_), .B(
        npu_inst_pe_1_1_7_add_79_carry_4_), .Z(npu_inst_pe_1_1_7_N77) );
  AND2_X1 npu_inst_pe_1_1_7_U133 ( .A1(npu_inst_pe_1_1_7_add_79_carry_4_), 
        .A2(npu_inst_pe_1_1_7_int_q_acc_4_), .ZN(
        npu_inst_pe_1_1_7_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_1_7_U132 ( .A(npu_inst_pe_1_1_7_int_q_acc_5_), .B(
        npu_inst_pe_1_1_7_add_79_carry_5_), .Z(npu_inst_pe_1_1_7_N78) );
  AND2_X1 npu_inst_pe_1_1_7_U131 ( .A1(npu_inst_pe_1_1_7_add_79_carry_5_), 
        .A2(npu_inst_pe_1_1_7_int_q_acc_5_), .ZN(
        npu_inst_pe_1_1_7_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_1_7_U130 ( .A(npu_inst_pe_1_1_7_int_q_acc_6_), .B(
        npu_inst_pe_1_1_7_add_79_carry_6_), .Z(npu_inst_pe_1_1_7_N79) );
  AND2_X1 npu_inst_pe_1_1_7_U129 ( .A1(npu_inst_pe_1_1_7_add_79_carry_6_), 
        .A2(npu_inst_pe_1_1_7_int_q_acc_6_), .ZN(
        npu_inst_pe_1_1_7_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_1_7_U128 ( .A(npu_inst_pe_1_1_7_int_q_acc_7_), .B(
        npu_inst_pe_1_1_7_add_79_carry_7_), .Z(npu_inst_pe_1_1_7_N80) );
  XNOR2_X1 npu_inst_pe_1_1_7_U127 ( .A(npu_inst_pe_1_1_7_sub_77_carry_2_), .B(
        npu_inst_pe_1_1_7_int_q_acc_2_), .ZN(npu_inst_pe_1_1_7_N67) );
  OR2_X1 npu_inst_pe_1_1_7_U126 ( .A1(npu_inst_pe_1_1_7_int_q_acc_2_), .A2(
        npu_inst_pe_1_1_7_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_1_7_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_1_7_U125 ( .A(npu_inst_pe_1_1_7_sub_77_carry_3_), .B(
        npu_inst_pe_1_1_7_int_q_acc_3_), .ZN(npu_inst_pe_1_1_7_N68) );
  OR2_X1 npu_inst_pe_1_1_7_U124 ( .A1(npu_inst_pe_1_1_7_int_q_acc_3_), .A2(
        npu_inst_pe_1_1_7_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_1_7_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_1_7_U123 ( .A(npu_inst_pe_1_1_7_sub_77_carry_4_), .B(
        npu_inst_pe_1_1_7_int_q_acc_4_), .ZN(npu_inst_pe_1_1_7_N69) );
  OR2_X1 npu_inst_pe_1_1_7_U122 ( .A1(npu_inst_pe_1_1_7_int_q_acc_4_), .A2(
        npu_inst_pe_1_1_7_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_1_7_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_1_7_U121 ( .A(npu_inst_pe_1_1_7_sub_77_carry_5_), .B(
        npu_inst_pe_1_1_7_int_q_acc_5_), .ZN(npu_inst_pe_1_1_7_N70) );
  OR2_X1 npu_inst_pe_1_1_7_U120 ( .A1(npu_inst_pe_1_1_7_int_q_acc_5_), .A2(
        npu_inst_pe_1_1_7_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_1_7_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_1_7_U119 ( .A(npu_inst_pe_1_1_7_sub_77_carry_6_), .B(
        npu_inst_pe_1_1_7_int_q_acc_6_), .ZN(npu_inst_pe_1_1_7_N71) );
  OR2_X1 npu_inst_pe_1_1_7_U118 ( .A1(npu_inst_pe_1_1_7_int_q_acc_6_), .A2(
        npu_inst_pe_1_1_7_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_1_7_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_1_7_U117 ( .A(npu_inst_pe_1_1_7_int_q_acc_7_), .B(
        npu_inst_pe_1_1_7_sub_77_carry_7_), .ZN(npu_inst_pe_1_1_7_N72) );
  INV_X1 npu_inst_pe_1_1_7_U116 ( .A(npu_inst_n79), .ZN(npu_inst_pe_1_1_7_n7)
         );
  INV_X1 npu_inst_pe_1_1_7_U115 ( .A(npu_inst_pe_1_1_7_n7), .ZN(
        npu_inst_pe_1_1_7_n6) );
  INV_X1 npu_inst_pe_1_1_7_U114 ( .A(npu_inst_n58), .ZN(npu_inst_pe_1_1_7_n3)
         );
  AOI22_X1 npu_inst_pe_1_1_7_U113 ( .A1(npu_inst_int_data_y_2__7__0_), .A2(
        npu_inst_pe_1_1_7_n58), .B1(npu_inst_pe_1_1_7_n114), .B2(
        npu_inst_pe_1_1_7_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_1_7_n57) );
  INV_X1 npu_inst_pe_1_1_7_U112 ( .A(npu_inst_pe_1_1_7_n57), .ZN(
        npu_inst_pe_1_1_7_n108) );
  AOI22_X1 npu_inst_pe_1_1_7_U111 ( .A1(npu_inst_int_data_y_2__7__0_), .A2(
        npu_inst_pe_1_1_7_n54), .B1(npu_inst_pe_1_1_7_n115), .B2(
        npu_inst_pe_1_1_7_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_1_7_n53) );
  INV_X1 npu_inst_pe_1_1_7_U110 ( .A(npu_inst_pe_1_1_7_n53), .ZN(
        npu_inst_pe_1_1_7_n109) );
  AOI22_X1 npu_inst_pe_1_1_7_U107 ( .A1(npu_inst_int_data_y_2__7__0_), .A2(
        npu_inst_pe_1_1_7_n50), .B1(npu_inst_pe_1_1_7_n116), .B2(
        npu_inst_pe_1_1_7_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_1_7_n49) );
  INV_X1 npu_inst_pe_1_1_7_U106 ( .A(npu_inst_pe_1_1_7_n49), .ZN(
        npu_inst_pe_1_1_7_n110) );
  AOI22_X1 npu_inst_pe_1_1_7_U105 ( .A1(npu_inst_int_data_y_2__7__0_), .A2(
        npu_inst_pe_1_1_7_n46), .B1(npu_inst_pe_1_1_7_n117), .B2(
        npu_inst_pe_1_1_7_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_1_7_n45) );
  INV_X1 npu_inst_pe_1_1_7_U104 ( .A(npu_inst_pe_1_1_7_n45), .ZN(
        npu_inst_pe_1_1_7_n111) );
  AOI22_X1 npu_inst_pe_1_1_7_U103 ( .A1(npu_inst_int_data_y_2__7__0_), .A2(
        npu_inst_pe_1_1_7_n42), .B1(npu_inst_pe_1_1_7_n119), .B2(
        npu_inst_pe_1_1_7_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_1_7_n41) );
  INV_X1 npu_inst_pe_1_1_7_U102 ( .A(npu_inst_pe_1_1_7_n41), .ZN(
        npu_inst_pe_1_1_7_n112) );
  AOI22_X1 npu_inst_pe_1_1_7_U101 ( .A1(npu_inst_int_data_y_2__7__1_), .A2(
        npu_inst_pe_1_1_7_n58), .B1(npu_inst_pe_1_1_7_n114), .B2(
        npu_inst_pe_1_1_7_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_1_7_n59) );
  INV_X1 npu_inst_pe_1_1_7_U100 ( .A(npu_inst_pe_1_1_7_n59), .ZN(
        npu_inst_pe_1_1_7_n102) );
  AOI22_X1 npu_inst_pe_1_1_7_U99 ( .A1(npu_inst_int_data_y_2__7__1_), .A2(
        npu_inst_pe_1_1_7_n54), .B1(npu_inst_pe_1_1_7_n115), .B2(
        npu_inst_pe_1_1_7_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_1_7_n55) );
  INV_X1 npu_inst_pe_1_1_7_U98 ( .A(npu_inst_pe_1_1_7_n55), .ZN(
        npu_inst_pe_1_1_7_n103) );
  AOI22_X1 npu_inst_pe_1_1_7_U97 ( .A1(npu_inst_int_data_y_2__7__1_), .A2(
        npu_inst_pe_1_1_7_n50), .B1(npu_inst_pe_1_1_7_n116), .B2(
        npu_inst_pe_1_1_7_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_1_7_n51) );
  INV_X1 npu_inst_pe_1_1_7_U96 ( .A(npu_inst_pe_1_1_7_n51), .ZN(
        npu_inst_pe_1_1_7_n104) );
  AOI22_X1 npu_inst_pe_1_1_7_U95 ( .A1(npu_inst_int_data_y_2__7__1_), .A2(
        npu_inst_pe_1_1_7_n46), .B1(npu_inst_pe_1_1_7_n117), .B2(
        npu_inst_pe_1_1_7_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_1_7_n47) );
  INV_X1 npu_inst_pe_1_1_7_U94 ( .A(npu_inst_pe_1_1_7_n47), .ZN(
        npu_inst_pe_1_1_7_n105) );
  AOI22_X1 npu_inst_pe_1_1_7_U93 ( .A1(npu_inst_int_data_y_2__7__1_), .A2(
        npu_inst_pe_1_1_7_n42), .B1(npu_inst_pe_1_1_7_n119), .B2(
        npu_inst_pe_1_1_7_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_1_7_n43) );
  INV_X1 npu_inst_pe_1_1_7_U92 ( .A(npu_inst_pe_1_1_7_n43), .ZN(
        npu_inst_pe_1_1_7_n106) );
  AOI22_X1 npu_inst_pe_1_1_7_U91 ( .A1(npu_inst_pe_1_1_7_n38), .A2(
        npu_inst_int_data_y_2__7__1_), .B1(npu_inst_pe_1_1_7_n118), .B2(
        npu_inst_pe_1_1_7_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_1_7_n39) );
  INV_X1 npu_inst_pe_1_1_7_U90 ( .A(npu_inst_pe_1_1_7_n39), .ZN(
        npu_inst_pe_1_1_7_n107) );
  AOI22_X1 npu_inst_pe_1_1_7_U89 ( .A1(npu_inst_pe_1_1_7_n38), .A2(
        npu_inst_int_data_y_2__7__0_), .B1(npu_inst_pe_1_1_7_n118), .B2(
        npu_inst_pe_1_1_7_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_1_7_n37) );
  INV_X1 npu_inst_pe_1_1_7_U88 ( .A(npu_inst_pe_1_1_7_n37), .ZN(
        npu_inst_pe_1_1_7_n113) );
  AND2_X1 npu_inst_pe_1_1_7_U87 ( .A1(npu_inst_pe_1_1_7_N93), .A2(npu_inst_n58), .ZN(npu_inst_int_data_y_1__7__0_) );
  AND2_X1 npu_inst_pe_1_1_7_U86 ( .A1(npu_inst_n58), .A2(npu_inst_pe_1_1_7_N94), .ZN(npu_inst_int_data_y_1__7__1_) );
  NOR3_X1 npu_inst_pe_1_1_7_U85 ( .A1(npu_inst_pe_1_1_7_n26), .A2(npu_inst_n58), .A3(npu_inst_int_ckg[48]), .ZN(npu_inst_pe_1_1_7_n85) );
  OR2_X1 npu_inst_pe_1_1_7_U84 ( .A1(npu_inst_pe_1_1_7_n85), .A2(
        npu_inst_pe_1_1_7_n2), .ZN(npu_inst_pe_1_1_7_N84) );
  AND2_X1 npu_inst_pe_1_1_7_U83 ( .A1(npu_inst_pe_1_1_7_int_q_acc_0_), .A2(
        npu_inst_pe_1_1_7_n1), .ZN(npu_inst_int_data_res_1__7__0_) );
  AND2_X1 npu_inst_pe_1_1_7_U82 ( .A1(npu_inst_pe_1_1_7_n2), .A2(
        npu_inst_pe_1_1_7_int_q_acc_7_), .ZN(npu_inst_int_data_res_1__7__7_)
         );
  AND2_X1 npu_inst_pe_1_1_7_U81 ( .A1(npu_inst_pe_1_1_7_int_q_acc_1_), .A2(
        npu_inst_pe_1_1_7_n1), .ZN(npu_inst_int_data_res_1__7__1_) );
  AND2_X1 npu_inst_pe_1_1_7_U80 ( .A1(npu_inst_pe_1_1_7_int_q_acc_2_), .A2(
        npu_inst_pe_1_1_7_n1), .ZN(npu_inst_int_data_res_1__7__2_) );
  AND2_X1 npu_inst_pe_1_1_7_U79 ( .A1(npu_inst_pe_1_1_7_int_q_acc_3_), .A2(
        npu_inst_pe_1_1_7_n2), .ZN(npu_inst_int_data_res_1__7__3_) );
  AND2_X1 npu_inst_pe_1_1_7_U78 ( .A1(npu_inst_pe_1_1_7_int_q_acc_4_), .A2(
        npu_inst_pe_1_1_7_n2), .ZN(npu_inst_int_data_res_1__7__4_) );
  AND2_X1 npu_inst_pe_1_1_7_U77 ( .A1(npu_inst_pe_1_1_7_int_q_acc_5_), .A2(
        npu_inst_pe_1_1_7_n2), .ZN(npu_inst_int_data_res_1__7__5_) );
  AND2_X1 npu_inst_pe_1_1_7_U76 ( .A1(npu_inst_pe_1_1_7_int_q_acc_6_), .A2(
        npu_inst_pe_1_1_7_n2), .ZN(npu_inst_int_data_res_1__7__6_) );
  AOI222_X1 npu_inst_pe_1_1_7_U75 ( .A1(npu_inst_int_data_res_2__7__0_), .A2(
        npu_inst_pe_1_1_7_n1), .B1(npu_inst_pe_1_1_7_N73), .B2(
        npu_inst_pe_1_1_7_n76), .C1(npu_inst_pe_1_1_7_N65), .C2(
        npu_inst_pe_1_1_7_n77), .ZN(npu_inst_pe_1_1_7_n84) );
  INV_X1 npu_inst_pe_1_1_7_U74 ( .A(npu_inst_pe_1_1_7_n84), .ZN(
        npu_inst_pe_1_1_7_n101) );
  AOI222_X1 npu_inst_pe_1_1_7_U73 ( .A1(npu_inst_int_data_res_2__7__7_), .A2(
        npu_inst_pe_1_1_7_n1), .B1(npu_inst_pe_1_1_7_N80), .B2(
        npu_inst_pe_1_1_7_n76), .C1(npu_inst_pe_1_1_7_N72), .C2(
        npu_inst_pe_1_1_7_n77), .ZN(npu_inst_pe_1_1_7_n75) );
  INV_X1 npu_inst_pe_1_1_7_U72 ( .A(npu_inst_pe_1_1_7_n75), .ZN(
        npu_inst_pe_1_1_7_n33) );
  AOI222_X1 npu_inst_pe_1_1_7_U71 ( .A1(npu_inst_int_data_res_2__7__1_), .A2(
        npu_inst_pe_1_1_7_n1), .B1(npu_inst_pe_1_1_7_N74), .B2(
        npu_inst_pe_1_1_7_n76), .C1(npu_inst_pe_1_1_7_N66), .C2(
        npu_inst_pe_1_1_7_n77), .ZN(npu_inst_pe_1_1_7_n83) );
  INV_X1 npu_inst_pe_1_1_7_U70 ( .A(npu_inst_pe_1_1_7_n83), .ZN(
        npu_inst_pe_1_1_7_n100) );
  AOI222_X1 npu_inst_pe_1_1_7_U69 ( .A1(npu_inst_int_data_res_2__7__2_), .A2(
        npu_inst_pe_1_1_7_n1), .B1(npu_inst_pe_1_1_7_N75), .B2(
        npu_inst_pe_1_1_7_n76), .C1(npu_inst_pe_1_1_7_N67), .C2(
        npu_inst_pe_1_1_7_n77), .ZN(npu_inst_pe_1_1_7_n82) );
  INV_X1 npu_inst_pe_1_1_7_U68 ( .A(npu_inst_pe_1_1_7_n82), .ZN(
        npu_inst_pe_1_1_7_n99) );
  AOI222_X1 npu_inst_pe_1_1_7_U67 ( .A1(npu_inst_int_data_res_2__7__3_), .A2(
        npu_inst_pe_1_1_7_n1), .B1(npu_inst_pe_1_1_7_N76), .B2(
        npu_inst_pe_1_1_7_n76), .C1(npu_inst_pe_1_1_7_N68), .C2(
        npu_inst_pe_1_1_7_n77), .ZN(npu_inst_pe_1_1_7_n81) );
  INV_X1 npu_inst_pe_1_1_7_U66 ( .A(npu_inst_pe_1_1_7_n81), .ZN(
        npu_inst_pe_1_1_7_n98) );
  AOI222_X1 npu_inst_pe_1_1_7_U65 ( .A1(npu_inst_int_data_res_2__7__4_), .A2(
        npu_inst_pe_1_1_7_n1), .B1(npu_inst_pe_1_1_7_N77), .B2(
        npu_inst_pe_1_1_7_n76), .C1(npu_inst_pe_1_1_7_N69), .C2(
        npu_inst_pe_1_1_7_n77), .ZN(npu_inst_pe_1_1_7_n80) );
  INV_X1 npu_inst_pe_1_1_7_U64 ( .A(npu_inst_pe_1_1_7_n80), .ZN(
        npu_inst_pe_1_1_7_n36) );
  AOI222_X1 npu_inst_pe_1_1_7_U63 ( .A1(npu_inst_int_data_res_2__7__5_), .A2(
        npu_inst_pe_1_1_7_n1), .B1(npu_inst_pe_1_1_7_N78), .B2(
        npu_inst_pe_1_1_7_n76), .C1(npu_inst_pe_1_1_7_N70), .C2(
        npu_inst_pe_1_1_7_n77), .ZN(npu_inst_pe_1_1_7_n79) );
  INV_X1 npu_inst_pe_1_1_7_U62 ( .A(npu_inst_pe_1_1_7_n79), .ZN(
        npu_inst_pe_1_1_7_n35) );
  AOI222_X1 npu_inst_pe_1_1_7_U61 ( .A1(npu_inst_int_data_res_2__7__6_), .A2(
        npu_inst_pe_1_1_7_n1), .B1(npu_inst_pe_1_1_7_N79), .B2(
        npu_inst_pe_1_1_7_n76), .C1(npu_inst_pe_1_1_7_N71), .C2(
        npu_inst_pe_1_1_7_n77), .ZN(npu_inst_pe_1_1_7_n78) );
  INV_X1 npu_inst_pe_1_1_7_U60 ( .A(npu_inst_pe_1_1_7_n78), .ZN(
        npu_inst_pe_1_1_7_n34) );
  INV_X1 npu_inst_pe_1_1_7_U59 ( .A(npu_inst_pe_1_1_7_int_data_1_), .ZN(
        npu_inst_pe_1_1_7_n14) );
  AND2_X1 npu_inst_pe_1_1_7_U58 ( .A1(npu_inst_int_data_x_1__7__1_), .A2(
        npu_inst_pe_1_1_7_int_q_weight_1_), .ZN(npu_inst_pe_1_1_7_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_1_7_U57 ( .A1(npu_inst_int_data_x_1__7__0_), .A2(
        npu_inst_pe_1_1_7_int_q_weight_1_), .ZN(npu_inst_pe_1_1_7_int_data_0_)
         );
  NAND2_X1 npu_inst_pe_1_1_7_U56 ( .A1(npu_inst_pe_1_1_7_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_1_7_n60), .ZN(npu_inst_pe_1_1_7_n74) );
  OAI21_X1 npu_inst_pe_1_1_7_U55 ( .B1(npu_inst_pe_1_1_7_n63), .B2(
        npu_inst_pe_1_1_7_n60), .A(npu_inst_pe_1_1_7_n74), .ZN(
        npu_inst_pe_1_1_7_n97) );
  NAND2_X1 npu_inst_pe_1_1_7_U54 ( .A1(npu_inst_pe_1_1_7_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_1_7_n60), .ZN(npu_inst_pe_1_1_7_n73) );
  OAI21_X1 npu_inst_pe_1_1_7_U53 ( .B1(npu_inst_pe_1_1_7_n61), .B2(
        npu_inst_pe_1_1_7_n60), .A(npu_inst_pe_1_1_7_n73), .ZN(
        npu_inst_pe_1_1_7_n96) );
  NAND2_X1 npu_inst_pe_1_1_7_U52 ( .A1(npu_inst_pe_1_1_7_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_1_7_n56), .ZN(npu_inst_pe_1_1_7_n72) );
  OAI21_X1 npu_inst_pe_1_1_7_U51 ( .B1(npu_inst_pe_1_1_7_n63), .B2(
        npu_inst_pe_1_1_7_n56), .A(npu_inst_pe_1_1_7_n72), .ZN(
        npu_inst_pe_1_1_7_n95) );
  NAND2_X1 npu_inst_pe_1_1_7_U50 ( .A1(npu_inst_pe_1_1_7_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_1_7_n56), .ZN(npu_inst_pe_1_1_7_n71) );
  OAI21_X1 npu_inst_pe_1_1_7_U49 ( .B1(npu_inst_pe_1_1_7_n61), .B2(
        npu_inst_pe_1_1_7_n56), .A(npu_inst_pe_1_1_7_n71), .ZN(
        npu_inst_pe_1_1_7_n94) );
  NAND2_X1 npu_inst_pe_1_1_7_U48 ( .A1(npu_inst_pe_1_1_7_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_1_7_n52), .ZN(npu_inst_pe_1_1_7_n70) );
  OAI21_X1 npu_inst_pe_1_1_7_U47 ( .B1(npu_inst_pe_1_1_7_n63), .B2(
        npu_inst_pe_1_1_7_n52), .A(npu_inst_pe_1_1_7_n70), .ZN(
        npu_inst_pe_1_1_7_n93) );
  NAND2_X1 npu_inst_pe_1_1_7_U46 ( .A1(npu_inst_pe_1_1_7_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_1_7_n52), .ZN(npu_inst_pe_1_1_7_n69) );
  OAI21_X1 npu_inst_pe_1_1_7_U45 ( .B1(npu_inst_pe_1_1_7_n61), .B2(
        npu_inst_pe_1_1_7_n52), .A(npu_inst_pe_1_1_7_n69), .ZN(
        npu_inst_pe_1_1_7_n92) );
  NAND2_X1 npu_inst_pe_1_1_7_U44 ( .A1(npu_inst_pe_1_1_7_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_1_7_n48), .ZN(npu_inst_pe_1_1_7_n68) );
  OAI21_X1 npu_inst_pe_1_1_7_U43 ( .B1(npu_inst_pe_1_1_7_n63), .B2(
        npu_inst_pe_1_1_7_n48), .A(npu_inst_pe_1_1_7_n68), .ZN(
        npu_inst_pe_1_1_7_n91) );
  NAND2_X1 npu_inst_pe_1_1_7_U42 ( .A1(npu_inst_pe_1_1_7_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_1_7_n48), .ZN(npu_inst_pe_1_1_7_n67) );
  OAI21_X1 npu_inst_pe_1_1_7_U41 ( .B1(npu_inst_pe_1_1_7_n61), .B2(
        npu_inst_pe_1_1_7_n48), .A(npu_inst_pe_1_1_7_n67), .ZN(
        npu_inst_pe_1_1_7_n90) );
  NAND2_X1 npu_inst_pe_1_1_7_U40 ( .A1(npu_inst_pe_1_1_7_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_1_7_n44), .ZN(npu_inst_pe_1_1_7_n66) );
  OAI21_X1 npu_inst_pe_1_1_7_U39 ( .B1(npu_inst_pe_1_1_7_n63), .B2(
        npu_inst_pe_1_1_7_n44), .A(npu_inst_pe_1_1_7_n66), .ZN(
        npu_inst_pe_1_1_7_n89) );
  NAND2_X1 npu_inst_pe_1_1_7_U38 ( .A1(npu_inst_pe_1_1_7_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_1_7_n44), .ZN(npu_inst_pe_1_1_7_n65) );
  OAI21_X1 npu_inst_pe_1_1_7_U37 ( .B1(npu_inst_pe_1_1_7_n61), .B2(
        npu_inst_pe_1_1_7_n44), .A(npu_inst_pe_1_1_7_n65), .ZN(
        npu_inst_pe_1_1_7_n88) );
  NAND2_X1 npu_inst_pe_1_1_7_U36 ( .A1(npu_inst_pe_1_1_7_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_1_7_n40), .ZN(npu_inst_pe_1_1_7_n64) );
  OAI21_X1 npu_inst_pe_1_1_7_U35 ( .B1(npu_inst_pe_1_1_7_n63), .B2(
        npu_inst_pe_1_1_7_n40), .A(npu_inst_pe_1_1_7_n64), .ZN(
        npu_inst_pe_1_1_7_n87) );
  NAND2_X1 npu_inst_pe_1_1_7_U34 ( .A1(npu_inst_pe_1_1_7_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_1_7_n40), .ZN(npu_inst_pe_1_1_7_n62) );
  OAI21_X1 npu_inst_pe_1_1_7_U33 ( .B1(npu_inst_pe_1_1_7_n61), .B2(
        npu_inst_pe_1_1_7_n40), .A(npu_inst_pe_1_1_7_n62), .ZN(
        npu_inst_pe_1_1_7_n86) );
  INV_X1 npu_inst_pe_1_1_7_U32 ( .A(npu_inst_pe_1_1_7_int_data_0_), .ZN(
        npu_inst_pe_1_1_7_n13) );
  AOI22_X1 npu_inst_pe_1_1_7_U31 ( .A1(npu_inst_n58), .A2(
        npu_inst_int_data_y_2__7__1_), .B1(npu_inst_pe_1_1_7_n3), .B2(
        int_i_data_h_npu2[1]), .ZN(npu_inst_pe_1_1_7_n63) );
  INV_X1 npu_inst_pe_1_1_7_U30 ( .A(npu_inst_n71), .ZN(npu_inst_pe_1_1_7_n5)
         );
  AOI22_X1 npu_inst_pe_1_1_7_U29 ( .A1(npu_inst_n58), .A2(
        npu_inst_int_data_y_2__7__0_), .B1(npu_inst_pe_1_1_7_n3), .B2(
        int_i_data_h_npu2[0]), .ZN(npu_inst_pe_1_1_7_n61) );
  OR3_X1 npu_inst_pe_1_1_7_U28 ( .A1(npu_inst_pe_1_1_7_n6), .A2(
        npu_inst_pe_1_1_7_n8), .A3(npu_inst_pe_1_1_7_n5), .ZN(
        npu_inst_pe_1_1_7_n56) );
  OR3_X1 npu_inst_pe_1_1_7_U27 ( .A1(npu_inst_pe_1_1_7_n5), .A2(
        npu_inst_pe_1_1_7_n8), .A3(npu_inst_pe_1_1_7_n7), .ZN(
        npu_inst_pe_1_1_7_n48) );
  INV_X1 npu_inst_pe_1_1_7_U26 ( .A(npu_inst_pe_1_1_7_n5), .ZN(
        npu_inst_pe_1_1_7_n4) );
  INV_X1 npu_inst_pe_1_1_7_U25 ( .A(npu_inst_n126), .ZN(npu_inst_pe_1_1_7_n12)
         );
  OR3_X1 npu_inst_pe_1_1_7_U24 ( .A1(npu_inst_pe_1_1_7_n4), .A2(
        npu_inst_pe_1_1_7_n8), .A3(npu_inst_pe_1_1_7_n7), .ZN(
        npu_inst_pe_1_1_7_n52) );
  OR3_X1 npu_inst_pe_1_1_7_U23 ( .A1(npu_inst_pe_1_1_7_n6), .A2(
        npu_inst_pe_1_1_7_n8), .A3(npu_inst_pe_1_1_7_n4), .ZN(
        npu_inst_pe_1_1_7_n60) );
  NOR2_X1 npu_inst_pe_1_1_7_U22 ( .A1(npu_inst_pe_1_1_7_n60), .A2(
        npu_inst_pe_1_1_7_n3), .ZN(npu_inst_pe_1_1_7_n58) );
  NOR2_X1 npu_inst_pe_1_1_7_U21 ( .A1(npu_inst_pe_1_1_7_n56), .A2(
        npu_inst_pe_1_1_7_n3), .ZN(npu_inst_pe_1_1_7_n54) );
  NOR2_X1 npu_inst_pe_1_1_7_U20 ( .A1(npu_inst_pe_1_1_7_n52), .A2(
        npu_inst_pe_1_1_7_n3), .ZN(npu_inst_pe_1_1_7_n50) );
  NOR2_X1 npu_inst_pe_1_1_7_U19 ( .A1(npu_inst_pe_1_1_7_n48), .A2(
        npu_inst_pe_1_1_7_n3), .ZN(npu_inst_pe_1_1_7_n46) );
  NOR2_X1 npu_inst_pe_1_1_7_U18 ( .A1(npu_inst_pe_1_1_7_n40), .A2(
        npu_inst_pe_1_1_7_n3), .ZN(npu_inst_pe_1_1_7_n38) );
  NOR2_X1 npu_inst_pe_1_1_7_U17 ( .A1(npu_inst_pe_1_1_7_n44), .A2(
        npu_inst_pe_1_1_7_n3), .ZN(npu_inst_pe_1_1_7_n42) );
  BUF_X1 npu_inst_pe_1_1_7_U16 ( .A(npu_inst_n104), .Z(npu_inst_pe_1_1_7_n8)
         );
  BUF_X1 npu_inst_pe_1_1_7_U15 ( .A(npu_inst_pe_1_1_7_n12), .Z(
        npu_inst_pe_1_1_7_n11) );
  BUF_X1 npu_inst_pe_1_1_7_U14 ( .A(npu_inst_pe_1_1_7_n12), .Z(
        npu_inst_pe_1_1_7_n10) );
  BUF_X1 npu_inst_pe_1_1_7_U13 ( .A(npu_inst_pe_1_1_7_n12), .Z(
        npu_inst_pe_1_1_7_n9) );
  INV_X1 npu_inst_pe_1_1_7_U12 ( .A(npu_inst_pe_1_1_7_n38), .ZN(
        npu_inst_pe_1_1_7_n118) );
  INV_X1 npu_inst_pe_1_1_7_U11 ( .A(npu_inst_pe_1_1_7_n58), .ZN(
        npu_inst_pe_1_1_7_n114) );
  INV_X1 npu_inst_pe_1_1_7_U10 ( .A(npu_inst_pe_1_1_7_n54), .ZN(
        npu_inst_pe_1_1_7_n115) );
  INV_X1 npu_inst_pe_1_1_7_U9 ( .A(npu_inst_pe_1_1_7_n50), .ZN(
        npu_inst_pe_1_1_7_n116) );
  INV_X1 npu_inst_pe_1_1_7_U8 ( .A(npu_inst_pe_1_1_7_n46), .ZN(
        npu_inst_pe_1_1_7_n117) );
  INV_X1 npu_inst_pe_1_1_7_U7 ( .A(npu_inst_pe_1_1_7_n42), .ZN(
        npu_inst_pe_1_1_7_n119) );
  BUF_X1 npu_inst_pe_1_1_7_U6 ( .A(npu_inst_n31), .Z(npu_inst_pe_1_1_7_n2) );
  BUF_X1 npu_inst_pe_1_1_7_U5 ( .A(npu_inst_n31), .Z(npu_inst_pe_1_1_7_n1) );
  NOR2_X1 npu_inst_pe_1_1_7_U4 ( .A1(npu_inst_pe_1_1_7_int_q_weight_0_), .A2(
        npu_inst_pe_1_1_7_n1), .ZN(npu_inst_pe_1_1_7_n76) );
  NOR2_X1 npu_inst_pe_1_1_7_U3 ( .A1(npu_inst_pe_1_1_7_n27), .A2(
        npu_inst_pe_1_1_7_n1), .ZN(npu_inst_pe_1_1_7_n77) );
  FA_X1 npu_inst_pe_1_1_7_sub_77_U2_1 ( .A(npu_inst_pe_1_1_7_int_q_acc_1_), 
        .B(npu_inst_pe_1_1_7_n14), .CI(npu_inst_pe_1_1_7_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_1_7_sub_77_carry_2_), .S(npu_inst_pe_1_1_7_N66) );
  FA_X1 npu_inst_pe_1_1_7_add_79_U1_1 ( .A(npu_inst_pe_1_1_7_int_q_acc_1_), 
        .B(npu_inst_pe_1_1_7_int_data_1_), .CI(
        npu_inst_pe_1_1_7_add_79_carry_1_), .CO(
        npu_inst_pe_1_1_7_add_79_carry_2_), .S(npu_inst_pe_1_1_7_N74) );
  NAND3_X1 npu_inst_pe_1_1_7_U109 ( .A1(npu_inst_pe_1_1_7_n5), .A2(
        npu_inst_pe_1_1_7_n7), .A3(npu_inst_pe_1_1_7_n8), .ZN(
        npu_inst_pe_1_1_7_n44) );
  NAND3_X1 npu_inst_pe_1_1_7_U108 ( .A1(npu_inst_pe_1_1_7_n4), .A2(
        npu_inst_pe_1_1_7_n7), .A3(npu_inst_pe_1_1_7_n8), .ZN(
        npu_inst_pe_1_1_7_n40) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_1_7_n34), .CK(
        npu_inst_pe_1_1_7_net3948), .RN(npu_inst_pe_1_1_7_n9), .Q(
        npu_inst_pe_1_1_7_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_1_7_n35), .CK(
        npu_inst_pe_1_1_7_net3948), .RN(npu_inst_pe_1_1_7_n9), .Q(
        npu_inst_pe_1_1_7_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_1_7_n36), .CK(
        npu_inst_pe_1_1_7_net3948), .RN(npu_inst_pe_1_1_7_n9), .Q(
        npu_inst_pe_1_1_7_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_1_7_n98), .CK(
        npu_inst_pe_1_1_7_net3948), .RN(npu_inst_pe_1_1_7_n9), .Q(
        npu_inst_pe_1_1_7_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_1_7_n99), .CK(
        npu_inst_pe_1_1_7_net3948), .RN(npu_inst_pe_1_1_7_n9), .Q(
        npu_inst_pe_1_1_7_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_1_7_n100), 
        .CK(npu_inst_pe_1_1_7_net3948), .RN(npu_inst_pe_1_1_7_n9), .Q(
        npu_inst_pe_1_1_7_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_1_7_n33), .CK(
        npu_inst_pe_1_1_7_net3948), .RN(npu_inst_pe_1_1_7_n9), .Q(
        npu_inst_pe_1_1_7_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_1_7_n101), 
        .CK(npu_inst_pe_1_1_7_net3948), .RN(npu_inst_pe_1_1_7_n9), .Q(
        npu_inst_pe_1_1_7_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_weight_reg_0_ ( .D(npu_inst_n112), .CK(
        npu_inst_pe_1_1_7_net3954), .RN(npu_inst_pe_1_1_7_n9), .Q(
        npu_inst_pe_1_1_7_int_q_weight_0_), .QN(npu_inst_pe_1_1_7_n27) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_weight_reg_1_ ( .D(npu_inst_n118), .CK(
        npu_inst_pe_1_1_7_net3954), .RN(npu_inst_pe_1_1_7_n9), .Q(
        npu_inst_pe_1_1_7_int_q_weight_1_), .QN(npu_inst_pe_1_1_7_n26) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_1_7_n113), 
        .CK(npu_inst_pe_1_1_7_net3954), .RN(npu_inst_pe_1_1_7_n9), .Q(
        npu_inst_pe_1_1_7_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_1_7_n107), 
        .CK(npu_inst_pe_1_1_7_net3954), .RN(npu_inst_pe_1_1_7_n9), .Q(
        npu_inst_pe_1_1_7_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_1_7_n112), 
        .CK(npu_inst_pe_1_1_7_net3954), .RN(npu_inst_pe_1_1_7_n10), .Q(
        npu_inst_pe_1_1_7_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_1_7_n106), 
        .CK(npu_inst_pe_1_1_7_net3954), .RN(npu_inst_pe_1_1_7_n10), .Q(
        npu_inst_pe_1_1_7_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_1_7_n111), 
        .CK(npu_inst_pe_1_1_7_net3954), .RN(npu_inst_pe_1_1_7_n10), .Q(
        npu_inst_pe_1_1_7_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_1_7_n105), 
        .CK(npu_inst_pe_1_1_7_net3954), .RN(npu_inst_pe_1_1_7_n10), .Q(
        npu_inst_pe_1_1_7_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_1_7_n110), 
        .CK(npu_inst_pe_1_1_7_net3954), .RN(npu_inst_pe_1_1_7_n10), .Q(
        npu_inst_pe_1_1_7_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_1_7_n104), 
        .CK(npu_inst_pe_1_1_7_net3954), .RN(npu_inst_pe_1_1_7_n10), .Q(
        npu_inst_pe_1_1_7_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_1_7_n109), 
        .CK(npu_inst_pe_1_1_7_net3954), .RN(npu_inst_pe_1_1_7_n10), .Q(
        npu_inst_pe_1_1_7_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_1_7_n103), 
        .CK(npu_inst_pe_1_1_7_net3954), .RN(npu_inst_pe_1_1_7_n10), .Q(
        npu_inst_pe_1_1_7_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_1_7_n108), 
        .CK(npu_inst_pe_1_1_7_net3954), .RN(npu_inst_pe_1_1_7_n10), .Q(
        npu_inst_pe_1_1_7_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_1_7_n102), 
        .CK(npu_inst_pe_1_1_7_net3954), .RN(npu_inst_pe_1_1_7_n10), .Q(
        npu_inst_pe_1_1_7_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_1_7_n86), 
        .CK(npu_inst_pe_1_1_7_net3954), .RN(npu_inst_pe_1_1_7_n10), .Q(
        npu_inst_pe_1_1_7_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_1_7_n87), 
        .CK(npu_inst_pe_1_1_7_net3954), .RN(npu_inst_pe_1_1_7_n10), .Q(
        npu_inst_pe_1_1_7_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_1_7_n88), 
        .CK(npu_inst_pe_1_1_7_net3954), .RN(npu_inst_pe_1_1_7_n11), .Q(
        npu_inst_pe_1_1_7_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_1_7_n89), 
        .CK(npu_inst_pe_1_1_7_net3954), .RN(npu_inst_pe_1_1_7_n11), .Q(
        npu_inst_pe_1_1_7_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_1_7_n90), 
        .CK(npu_inst_pe_1_1_7_net3954), .RN(npu_inst_pe_1_1_7_n11), .Q(
        npu_inst_pe_1_1_7_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_1_7_n91), 
        .CK(npu_inst_pe_1_1_7_net3954), .RN(npu_inst_pe_1_1_7_n11), .Q(
        npu_inst_pe_1_1_7_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_1_7_n92), 
        .CK(npu_inst_pe_1_1_7_net3954), .RN(npu_inst_pe_1_1_7_n11), .Q(
        npu_inst_pe_1_1_7_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_1_7_n93), 
        .CK(npu_inst_pe_1_1_7_net3954), .RN(npu_inst_pe_1_1_7_n11), .Q(
        npu_inst_pe_1_1_7_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_1_7_n94), 
        .CK(npu_inst_pe_1_1_7_net3954), .RN(npu_inst_pe_1_1_7_n11), .Q(
        npu_inst_pe_1_1_7_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_1_7_n95), 
        .CK(npu_inst_pe_1_1_7_net3954), .RN(npu_inst_pe_1_1_7_n11), .Q(
        npu_inst_pe_1_1_7_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_1_7_n96), 
        .CK(npu_inst_pe_1_1_7_net3954), .RN(npu_inst_pe_1_1_7_n11), .Q(
        npu_inst_pe_1_1_7_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_1_7_n97), 
        .CK(npu_inst_pe_1_1_7_net3954), .RN(npu_inst_pe_1_1_7_n11), .Q(
        npu_inst_pe_1_1_7_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_1_7_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_1_7_N84), .SE(1'b0), .GCK(npu_inst_pe_1_1_7_net3948) );
  CLKGATETST_X1 npu_inst_pe_1_1_7_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n65), .SE(1'b0), .GCK(npu_inst_pe_1_1_7_net3954) );
  MUX2_X1 npu_inst_pe_1_2_0_U161 ( .A(npu_inst_pe_1_2_0_n31), .B(
        npu_inst_pe_1_2_0_n28), .S(npu_inst_pe_1_2_0_n7), .Z(
        npu_inst_pe_1_2_0_N93) );
  MUX2_X1 npu_inst_pe_1_2_0_U160 ( .A(npu_inst_pe_1_2_0_n30), .B(
        npu_inst_pe_1_2_0_n29), .S(npu_inst_n78), .Z(npu_inst_pe_1_2_0_n31) );
  MUX2_X1 npu_inst_pe_1_2_0_U159 ( .A(npu_inst_pe_1_2_0_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_2_0_int_q_reg_v_1__0_), .S(npu_inst_pe_1_2_0_n4), .Z(
        npu_inst_pe_1_2_0_n30) );
  MUX2_X1 npu_inst_pe_1_2_0_U158 ( .A(npu_inst_pe_1_2_0_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_2_0_int_q_reg_v_3__0_), .S(npu_inst_pe_1_2_0_n4), .Z(
        npu_inst_pe_1_2_0_n29) );
  MUX2_X1 npu_inst_pe_1_2_0_U157 ( .A(npu_inst_pe_1_2_0_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_2_0_int_q_reg_v_5__0_), .S(npu_inst_pe_1_2_0_n4), .Z(
        npu_inst_pe_1_2_0_n28) );
  MUX2_X1 npu_inst_pe_1_2_0_U156 ( .A(npu_inst_pe_1_2_0_n25), .B(
        npu_inst_pe_1_2_0_n22), .S(npu_inst_pe_1_2_0_n7), .Z(
        npu_inst_pe_1_2_0_N94) );
  MUX2_X1 npu_inst_pe_1_2_0_U155 ( .A(npu_inst_pe_1_2_0_n24), .B(
        npu_inst_pe_1_2_0_n23), .S(npu_inst_n78), .Z(npu_inst_pe_1_2_0_n25) );
  MUX2_X1 npu_inst_pe_1_2_0_U154 ( .A(npu_inst_pe_1_2_0_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_2_0_int_q_reg_v_1__1_), .S(npu_inst_pe_1_2_0_n4), .Z(
        npu_inst_pe_1_2_0_n24) );
  MUX2_X1 npu_inst_pe_1_2_0_U153 ( .A(npu_inst_pe_1_2_0_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_2_0_int_q_reg_v_3__1_), .S(npu_inst_pe_1_2_0_n4), .Z(
        npu_inst_pe_1_2_0_n23) );
  MUX2_X1 npu_inst_pe_1_2_0_U152 ( .A(npu_inst_pe_1_2_0_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_2_0_int_q_reg_v_5__1_), .S(npu_inst_pe_1_2_0_n4), .Z(
        npu_inst_pe_1_2_0_n22) );
  MUX2_X1 npu_inst_pe_1_2_0_U151 ( .A(npu_inst_pe_1_2_0_n21), .B(
        npu_inst_pe_1_2_0_n18), .S(npu_inst_pe_1_2_0_n7), .Z(
        npu_inst_pe_1_2_0_o_data_h_1_) );
  MUX2_X1 npu_inst_pe_1_2_0_U150 ( .A(npu_inst_pe_1_2_0_n20), .B(
        npu_inst_pe_1_2_0_n19), .S(npu_inst_n78), .Z(npu_inst_pe_1_2_0_n21) );
  MUX2_X1 npu_inst_pe_1_2_0_U149 ( .A(npu_inst_pe_1_2_0_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_2_0_int_q_reg_h_1__1_), .S(npu_inst_pe_1_2_0_n4), .Z(
        npu_inst_pe_1_2_0_n20) );
  MUX2_X1 npu_inst_pe_1_2_0_U148 ( .A(npu_inst_pe_1_2_0_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_2_0_int_q_reg_h_3__1_), .S(npu_inst_pe_1_2_0_n4), .Z(
        npu_inst_pe_1_2_0_n19) );
  MUX2_X1 npu_inst_pe_1_2_0_U147 ( .A(npu_inst_pe_1_2_0_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_2_0_int_q_reg_h_5__1_), .S(npu_inst_pe_1_2_0_n4), .Z(
        npu_inst_pe_1_2_0_n18) );
  MUX2_X1 npu_inst_pe_1_2_0_U146 ( .A(npu_inst_pe_1_2_0_n17), .B(
        npu_inst_pe_1_2_0_n14), .S(npu_inst_pe_1_2_0_n7), .Z(
        npu_inst_pe_1_2_0_o_data_h_0_) );
  MUX2_X1 npu_inst_pe_1_2_0_U145 ( .A(npu_inst_pe_1_2_0_n16), .B(
        npu_inst_pe_1_2_0_n15), .S(npu_inst_n78), .Z(npu_inst_pe_1_2_0_n17) );
  MUX2_X1 npu_inst_pe_1_2_0_U144 ( .A(npu_inst_pe_1_2_0_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_2_0_int_q_reg_h_1__0_), .S(npu_inst_pe_1_2_0_n4), .Z(
        npu_inst_pe_1_2_0_n16) );
  MUX2_X1 npu_inst_pe_1_2_0_U143 ( .A(npu_inst_pe_1_2_0_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_2_0_int_q_reg_h_3__0_), .S(npu_inst_pe_1_2_0_n4), .Z(
        npu_inst_pe_1_2_0_n15) );
  MUX2_X1 npu_inst_pe_1_2_0_U142 ( .A(npu_inst_pe_1_2_0_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_2_0_int_q_reg_h_5__0_), .S(npu_inst_pe_1_2_0_n4), .Z(
        npu_inst_pe_1_2_0_n14) );
  XOR2_X1 npu_inst_pe_1_2_0_U141 ( .A(npu_inst_pe_1_2_0_int_data_0_), .B(
        npu_inst_pe_1_2_0_int_q_acc_0_), .Z(npu_inst_pe_1_2_0_N73) );
  AND2_X1 npu_inst_pe_1_2_0_U140 ( .A1(npu_inst_pe_1_2_0_int_q_acc_0_), .A2(
        npu_inst_pe_1_2_0_int_data_0_), .ZN(npu_inst_pe_1_2_0_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_2_0_U139 ( .A(npu_inst_pe_1_2_0_int_q_acc_0_), .B(
        npu_inst_pe_1_2_0_n12), .ZN(npu_inst_pe_1_2_0_N65) );
  OR2_X1 npu_inst_pe_1_2_0_U138 ( .A1(npu_inst_pe_1_2_0_n12), .A2(
        npu_inst_pe_1_2_0_int_q_acc_0_), .ZN(npu_inst_pe_1_2_0_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_2_0_U137 ( .A(npu_inst_pe_1_2_0_int_q_acc_2_), .B(
        npu_inst_pe_1_2_0_add_79_carry_2_), .Z(npu_inst_pe_1_2_0_N75) );
  AND2_X1 npu_inst_pe_1_2_0_U136 ( .A1(npu_inst_pe_1_2_0_add_79_carry_2_), 
        .A2(npu_inst_pe_1_2_0_int_q_acc_2_), .ZN(
        npu_inst_pe_1_2_0_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_2_0_U135 ( .A(npu_inst_pe_1_2_0_int_q_acc_3_), .B(
        npu_inst_pe_1_2_0_add_79_carry_3_), .Z(npu_inst_pe_1_2_0_N76) );
  AND2_X1 npu_inst_pe_1_2_0_U134 ( .A1(npu_inst_pe_1_2_0_add_79_carry_3_), 
        .A2(npu_inst_pe_1_2_0_int_q_acc_3_), .ZN(
        npu_inst_pe_1_2_0_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_2_0_U133 ( .A(npu_inst_pe_1_2_0_int_q_acc_4_), .B(
        npu_inst_pe_1_2_0_add_79_carry_4_), .Z(npu_inst_pe_1_2_0_N77) );
  AND2_X1 npu_inst_pe_1_2_0_U132 ( .A1(npu_inst_pe_1_2_0_add_79_carry_4_), 
        .A2(npu_inst_pe_1_2_0_int_q_acc_4_), .ZN(
        npu_inst_pe_1_2_0_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_2_0_U131 ( .A(npu_inst_pe_1_2_0_int_q_acc_5_), .B(
        npu_inst_pe_1_2_0_add_79_carry_5_), .Z(npu_inst_pe_1_2_0_N78) );
  AND2_X1 npu_inst_pe_1_2_0_U130 ( .A1(npu_inst_pe_1_2_0_add_79_carry_5_), 
        .A2(npu_inst_pe_1_2_0_int_q_acc_5_), .ZN(
        npu_inst_pe_1_2_0_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_2_0_U129 ( .A(npu_inst_pe_1_2_0_int_q_acc_6_), .B(
        npu_inst_pe_1_2_0_add_79_carry_6_), .Z(npu_inst_pe_1_2_0_N79) );
  AND2_X1 npu_inst_pe_1_2_0_U128 ( .A1(npu_inst_pe_1_2_0_add_79_carry_6_), 
        .A2(npu_inst_pe_1_2_0_int_q_acc_6_), .ZN(
        npu_inst_pe_1_2_0_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_2_0_U127 ( .A(npu_inst_pe_1_2_0_int_q_acc_7_), .B(
        npu_inst_pe_1_2_0_add_79_carry_7_), .Z(npu_inst_pe_1_2_0_N80) );
  XNOR2_X1 npu_inst_pe_1_2_0_U126 ( .A(npu_inst_pe_1_2_0_sub_77_carry_2_), .B(
        npu_inst_pe_1_2_0_int_q_acc_2_), .ZN(npu_inst_pe_1_2_0_N67) );
  OR2_X1 npu_inst_pe_1_2_0_U125 ( .A1(npu_inst_pe_1_2_0_int_q_acc_2_), .A2(
        npu_inst_pe_1_2_0_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_2_0_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_2_0_U124 ( .A(npu_inst_pe_1_2_0_sub_77_carry_3_), .B(
        npu_inst_pe_1_2_0_int_q_acc_3_), .ZN(npu_inst_pe_1_2_0_N68) );
  OR2_X1 npu_inst_pe_1_2_0_U123 ( .A1(npu_inst_pe_1_2_0_int_q_acc_3_), .A2(
        npu_inst_pe_1_2_0_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_2_0_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_2_0_U122 ( .A(npu_inst_pe_1_2_0_sub_77_carry_4_), .B(
        npu_inst_pe_1_2_0_int_q_acc_4_), .ZN(npu_inst_pe_1_2_0_N69) );
  OR2_X1 npu_inst_pe_1_2_0_U121 ( .A1(npu_inst_pe_1_2_0_int_q_acc_4_), .A2(
        npu_inst_pe_1_2_0_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_2_0_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_2_0_U120 ( .A(npu_inst_pe_1_2_0_sub_77_carry_5_), .B(
        npu_inst_pe_1_2_0_int_q_acc_5_), .ZN(npu_inst_pe_1_2_0_N70) );
  OR2_X1 npu_inst_pe_1_2_0_U119 ( .A1(npu_inst_pe_1_2_0_int_q_acc_5_), .A2(
        npu_inst_pe_1_2_0_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_2_0_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_2_0_U118 ( .A(npu_inst_pe_1_2_0_sub_77_carry_6_), .B(
        npu_inst_pe_1_2_0_int_q_acc_6_), .ZN(npu_inst_pe_1_2_0_N71) );
  OR2_X1 npu_inst_pe_1_2_0_U117 ( .A1(npu_inst_pe_1_2_0_int_q_acc_6_), .A2(
        npu_inst_pe_1_2_0_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_2_0_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_2_0_U116 ( .A(npu_inst_pe_1_2_0_int_q_acc_7_), .B(
        npu_inst_pe_1_2_0_sub_77_carry_7_), .ZN(npu_inst_pe_1_2_0_N72) );
  INV_X1 npu_inst_pe_1_2_0_U115 ( .A(npu_inst_n78), .ZN(npu_inst_pe_1_2_0_n6)
         );
  INV_X1 npu_inst_pe_1_2_0_U114 ( .A(npu_inst_n58), .ZN(npu_inst_pe_1_2_0_n3)
         );
  AOI22_X1 npu_inst_pe_1_2_0_U113 ( .A1(npu_inst_int_data_y_3__0__0_), .A2(
        npu_inst_pe_1_2_0_n58), .B1(npu_inst_pe_1_2_0_n113), .B2(
        npu_inst_pe_1_2_0_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_2_0_n57) );
  INV_X1 npu_inst_pe_1_2_0_U112 ( .A(npu_inst_pe_1_2_0_n57), .ZN(
        npu_inst_pe_1_2_0_n107) );
  AOI22_X1 npu_inst_pe_1_2_0_U111 ( .A1(npu_inst_int_data_y_3__0__0_), .A2(
        npu_inst_pe_1_2_0_n54), .B1(npu_inst_pe_1_2_0_n114), .B2(
        npu_inst_pe_1_2_0_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_2_0_n53) );
  INV_X1 npu_inst_pe_1_2_0_U110 ( .A(npu_inst_pe_1_2_0_n53), .ZN(
        npu_inst_pe_1_2_0_n108) );
  AOI22_X1 npu_inst_pe_1_2_0_U107 ( .A1(npu_inst_int_data_y_3__0__0_), .A2(
        npu_inst_pe_1_2_0_n50), .B1(npu_inst_pe_1_2_0_n115), .B2(
        npu_inst_pe_1_2_0_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_2_0_n49) );
  INV_X1 npu_inst_pe_1_2_0_U106 ( .A(npu_inst_pe_1_2_0_n49), .ZN(
        npu_inst_pe_1_2_0_n109) );
  AOI22_X1 npu_inst_pe_1_2_0_U105 ( .A1(npu_inst_int_data_y_3__0__0_), .A2(
        npu_inst_pe_1_2_0_n46), .B1(npu_inst_pe_1_2_0_n116), .B2(
        npu_inst_pe_1_2_0_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_2_0_n45) );
  INV_X1 npu_inst_pe_1_2_0_U104 ( .A(npu_inst_pe_1_2_0_n45), .ZN(
        npu_inst_pe_1_2_0_n110) );
  AOI22_X1 npu_inst_pe_1_2_0_U103 ( .A1(npu_inst_int_data_y_3__0__0_), .A2(
        npu_inst_pe_1_2_0_n42), .B1(npu_inst_pe_1_2_0_n118), .B2(
        npu_inst_pe_1_2_0_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_2_0_n41) );
  INV_X1 npu_inst_pe_1_2_0_U102 ( .A(npu_inst_pe_1_2_0_n41), .ZN(
        npu_inst_pe_1_2_0_n111) );
  AOI22_X1 npu_inst_pe_1_2_0_U101 ( .A1(npu_inst_int_data_y_3__0__1_), .A2(
        npu_inst_pe_1_2_0_n58), .B1(npu_inst_pe_1_2_0_n113), .B2(
        npu_inst_pe_1_2_0_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_2_0_n59) );
  INV_X1 npu_inst_pe_1_2_0_U100 ( .A(npu_inst_pe_1_2_0_n59), .ZN(
        npu_inst_pe_1_2_0_n101) );
  AOI22_X1 npu_inst_pe_1_2_0_U99 ( .A1(npu_inst_int_data_y_3__0__1_), .A2(
        npu_inst_pe_1_2_0_n54), .B1(npu_inst_pe_1_2_0_n114), .B2(
        npu_inst_pe_1_2_0_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_2_0_n55) );
  INV_X1 npu_inst_pe_1_2_0_U98 ( .A(npu_inst_pe_1_2_0_n55), .ZN(
        npu_inst_pe_1_2_0_n102) );
  AOI22_X1 npu_inst_pe_1_2_0_U97 ( .A1(npu_inst_int_data_y_3__0__1_), .A2(
        npu_inst_pe_1_2_0_n50), .B1(npu_inst_pe_1_2_0_n115), .B2(
        npu_inst_pe_1_2_0_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_2_0_n51) );
  INV_X1 npu_inst_pe_1_2_0_U96 ( .A(npu_inst_pe_1_2_0_n51), .ZN(
        npu_inst_pe_1_2_0_n103) );
  AOI22_X1 npu_inst_pe_1_2_0_U95 ( .A1(npu_inst_int_data_y_3__0__1_), .A2(
        npu_inst_pe_1_2_0_n46), .B1(npu_inst_pe_1_2_0_n116), .B2(
        npu_inst_pe_1_2_0_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_2_0_n47) );
  INV_X1 npu_inst_pe_1_2_0_U94 ( .A(npu_inst_pe_1_2_0_n47), .ZN(
        npu_inst_pe_1_2_0_n104) );
  AOI22_X1 npu_inst_pe_1_2_0_U93 ( .A1(npu_inst_int_data_y_3__0__1_), .A2(
        npu_inst_pe_1_2_0_n42), .B1(npu_inst_pe_1_2_0_n118), .B2(
        npu_inst_pe_1_2_0_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_2_0_n43) );
  INV_X1 npu_inst_pe_1_2_0_U92 ( .A(npu_inst_pe_1_2_0_n43), .ZN(
        npu_inst_pe_1_2_0_n105) );
  AOI22_X1 npu_inst_pe_1_2_0_U91 ( .A1(npu_inst_pe_1_2_0_n38), .A2(
        npu_inst_int_data_y_3__0__1_), .B1(npu_inst_pe_1_2_0_n117), .B2(
        npu_inst_pe_1_2_0_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_2_0_n39) );
  INV_X1 npu_inst_pe_1_2_0_U90 ( .A(npu_inst_pe_1_2_0_n39), .ZN(
        npu_inst_pe_1_2_0_n106) );
  AOI22_X1 npu_inst_pe_1_2_0_U89 ( .A1(npu_inst_pe_1_2_0_n38), .A2(
        npu_inst_int_data_y_3__0__0_), .B1(npu_inst_pe_1_2_0_n117), .B2(
        npu_inst_pe_1_2_0_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_2_0_n37) );
  INV_X1 npu_inst_pe_1_2_0_U88 ( .A(npu_inst_pe_1_2_0_n37), .ZN(
        npu_inst_pe_1_2_0_n112) );
  NAND2_X1 npu_inst_pe_1_2_0_U87 ( .A1(npu_inst_pe_1_2_0_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_2_0_n60), .ZN(npu_inst_pe_1_2_0_n74) );
  OAI21_X1 npu_inst_pe_1_2_0_U86 ( .B1(npu_inst_pe_1_2_0_n63), .B2(
        npu_inst_pe_1_2_0_n60), .A(npu_inst_pe_1_2_0_n74), .ZN(
        npu_inst_pe_1_2_0_n97) );
  NAND2_X1 npu_inst_pe_1_2_0_U85 ( .A1(npu_inst_pe_1_2_0_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_2_0_n60), .ZN(npu_inst_pe_1_2_0_n73) );
  OAI21_X1 npu_inst_pe_1_2_0_U84 ( .B1(npu_inst_pe_1_2_0_n61), .B2(
        npu_inst_pe_1_2_0_n60), .A(npu_inst_pe_1_2_0_n73), .ZN(
        npu_inst_pe_1_2_0_n96) );
  NAND2_X1 npu_inst_pe_1_2_0_U83 ( .A1(npu_inst_pe_1_2_0_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_2_0_n56), .ZN(npu_inst_pe_1_2_0_n72) );
  OAI21_X1 npu_inst_pe_1_2_0_U82 ( .B1(npu_inst_pe_1_2_0_n63), .B2(
        npu_inst_pe_1_2_0_n56), .A(npu_inst_pe_1_2_0_n72), .ZN(
        npu_inst_pe_1_2_0_n95) );
  NAND2_X1 npu_inst_pe_1_2_0_U81 ( .A1(npu_inst_pe_1_2_0_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_2_0_n56), .ZN(npu_inst_pe_1_2_0_n71) );
  OAI21_X1 npu_inst_pe_1_2_0_U80 ( .B1(npu_inst_pe_1_2_0_n61), .B2(
        npu_inst_pe_1_2_0_n56), .A(npu_inst_pe_1_2_0_n71), .ZN(
        npu_inst_pe_1_2_0_n94) );
  NAND2_X1 npu_inst_pe_1_2_0_U79 ( .A1(npu_inst_pe_1_2_0_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_2_0_n52), .ZN(npu_inst_pe_1_2_0_n70) );
  OAI21_X1 npu_inst_pe_1_2_0_U78 ( .B1(npu_inst_pe_1_2_0_n63), .B2(
        npu_inst_pe_1_2_0_n52), .A(npu_inst_pe_1_2_0_n70), .ZN(
        npu_inst_pe_1_2_0_n93) );
  NAND2_X1 npu_inst_pe_1_2_0_U77 ( .A1(npu_inst_pe_1_2_0_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_2_0_n52), .ZN(npu_inst_pe_1_2_0_n69) );
  OAI21_X1 npu_inst_pe_1_2_0_U76 ( .B1(npu_inst_pe_1_2_0_n61), .B2(
        npu_inst_pe_1_2_0_n52), .A(npu_inst_pe_1_2_0_n69), .ZN(
        npu_inst_pe_1_2_0_n92) );
  NAND2_X1 npu_inst_pe_1_2_0_U75 ( .A1(npu_inst_pe_1_2_0_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_2_0_n48), .ZN(npu_inst_pe_1_2_0_n68) );
  OAI21_X1 npu_inst_pe_1_2_0_U74 ( .B1(npu_inst_pe_1_2_0_n63), .B2(
        npu_inst_pe_1_2_0_n48), .A(npu_inst_pe_1_2_0_n68), .ZN(
        npu_inst_pe_1_2_0_n91) );
  NAND2_X1 npu_inst_pe_1_2_0_U73 ( .A1(npu_inst_pe_1_2_0_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_2_0_n48), .ZN(npu_inst_pe_1_2_0_n67) );
  OAI21_X1 npu_inst_pe_1_2_0_U72 ( .B1(npu_inst_pe_1_2_0_n61), .B2(
        npu_inst_pe_1_2_0_n48), .A(npu_inst_pe_1_2_0_n67), .ZN(
        npu_inst_pe_1_2_0_n90) );
  NAND2_X1 npu_inst_pe_1_2_0_U71 ( .A1(npu_inst_pe_1_2_0_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_2_0_n44), .ZN(npu_inst_pe_1_2_0_n66) );
  OAI21_X1 npu_inst_pe_1_2_0_U70 ( .B1(npu_inst_pe_1_2_0_n63), .B2(
        npu_inst_pe_1_2_0_n44), .A(npu_inst_pe_1_2_0_n66), .ZN(
        npu_inst_pe_1_2_0_n89) );
  NAND2_X1 npu_inst_pe_1_2_0_U69 ( .A1(npu_inst_pe_1_2_0_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_2_0_n44), .ZN(npu_inst_pe_1_2_0_n65) );
  OAI21_X1 npu_inst_pe_1_2_0_U68 ( .B1(npu_inst_pe_1_2_0_n61), .B2(
        npu_inst_pe_1_2_0_n44), .A(npu_inst_pe_1_2_0_n65), .ZN(
        npu_inst_pe_1_2_0_n88) );
  NAND2_X1 npu_inst_pe_1_2_0_U67 ( .A1(npu_inst_pe_1_2_0_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_2_0_n40), .ZN(npu_inst_pe_1_2_0_n64) );
  OAI21_X1 npu_inst_pe_1_2_0_U66 ( .B1(npu_inst_pe_1_2_0_n63), .B2(
        npu_inst_pe_1_2_0_n40), .A(npu_inst_pe_1_2_0_n64), .ZN(
        npu_inst_pe_1_2_0_n87) );
  NAND2_X1 npu_inst_pe_1_2_0_U65 ( .A1(npu_inst_pe_1_2_0_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_2_0_n40), .ZN(npu_inst_pe_1_2_0_n62) );
  OAI21_X1 npu_inst_pe_1_2_0_U64 ( .B1(npu_inst_pe_1_2_0_n61), .B2(
        npu_inst_pe_1_2_0_n40), .A(npu_inst_pe_1_2_0_n62), .ZN(
        npu_inst_pe_1_2_0_n86) );
  AND2_X1 npu_inst_pe_1_2_0_U63 ( .A1(npu_inst_pe_1_2_0_N93), .A2(npu_inst_n58), .ZN(npu_inst_int_data_y_2__0__0_) );
  AND2_X1 npu_inst_pe_1_2_0_U62 ( .A1(npu_inst_n58), .A2(npu_inst_pe_1_2_0_N94), .ZN(npu_inst_int_data_y_2__0__1_) );
  NOR3_X1 npu_inst_pe_1_2_0_U61 ( .A1(npu_inst_pe_1_2_0_n26), .A2(npu_inst_n58), .A3(npu_inst_int_ckg[47]), .ZN(npu_inst_pe_1_2_0_n85) );
  OR2_X1 npu_inst_pe_1_2_0_U60 ( .A1(npu_inst_pe_1_2_0_n85), .A2(
        npu_inst_pe_1_2_0_n2), .ZN(npu_inst_pe_1_2_0_N84) );
  AND2_X1 npu_inst_pe_1_2_0_U59 ( .A1(npu_inst_pe_1_2_0_int_q_acc_0_), .A2(
        npu_inst_pe_1_2_0_n1), .ZN(npu_inst_int_data_res_2__0__0_) );
  AND2_X1 npu_inst_pe_1_2_0_U58 ( .A1(npu_inst_pe_1_2_0_n2), .A2(
        npu_inst_pe_1_2_0_int_q_acc_7_), .ZN(npu_inst_int_data_res_2__0__7_)
         );
  AND2_X1 npu_inst_pe_1_2_0_U57 ( .A1(npu_inst_pe_1_2_0_int_q_acc_1_), .A2(
        npu_inst_pe_1_2_0_n1), .ZN(npu_inst_int_data_res_2__0__1_) );
  AND2_X1 npu_inst_pe_1_2_0_U56 ( .A1(npu_inst_pe_1_2_0_int_q_acc_2_), .A2(
        npu_inst_pe_1_2_0_n1), .ZN(npu_inst_int_data_res_2__0__2_) );
  AND2_X1 npu_inst_pe_1_2_0_U55 ( .A1(npu_inst_pe_1_2_0_int_q_acc_3_), .A2(
        npu_inst_pe_1_2_0_n2), .ZN(npu_inst_int_data_res_2__0__3_) );
  AND2_X1 npu_inst_pe_1_2_0_U54 ( .A1(npu_inst_pe_1_2_0_int_q_acc_4_), .A2(
        npu_inst_pe_1_2_0_n2), .ZN(npu_inst_int_data_res_2__0__4_) );
  AND2_X1 npu_inst_pe_1_2_0_U53 ( .A1(npu_inst_pe_1_2_0_int_q_acc_5_), .A2(
        npu_inst_pe_1_2_0_n2), .ZN(npu_inst_int_data_res_2__0__5_) );
  AND2_X1 npu_inst_pe_1_2_0_U52 ( .A1(npu_inst_pe_1_2_0_int_q_acc_6_), .A2(
        npu_inst_pe_1_2_0_n2), .ZN(npu_inst_int_data_res_2__0__6_) );
  AOI222_X1 npu_inst_pe_1_2_0_U51 ( .A1(npu_inst_int_data_res_3__0__0_), .A2(
        npu_inst_pe_1_2_0_n1), .B1(npu_inst_pe_1_2_0_N73), .B2(
        npu_inst_pe_1_2_0_n76), .C1(npu_inst_pe_1_2_0_N65), .C2(
        npu_inst_pe_1_2_0_n77), .ZN(npu_inst_pe_1_2_0_n84) );
  INV_X1 npu_inst_pe_1_2_0_U50 ( .A(npu_inst_pe_1_2_0_n84), .ZN(
        npu_inst_pe_1_2_0_n100) );
  AOI222_X1 npu_inst_pe_1_2_0_U49 ( .A1(npu_inst_int_data_res_3__0__7_), .A2(
        npu_inst_pe_1_2_0_n1), .B1(npu_inst_pe_1_2_0_N80), .B2(
        npu_inst_pe_1_2_0_n76), .C1(npu_inst_pe_1_2_0_N72), .C2(
        npu_inst_pe_1_2_0_n77), .ZN(npu_inst_pe_1_2_0_n75) );
  INV_X1 npu_inst_pe_1_2_0_U48 ( .A(npu_inst_pe_1_2_0_n75), .ZN(
        npu_inst_pe_1_2_0_n32) );
  AOI222_X1 npu_inst_pe_1_2_0_U47 ( .A1(npu_inst_int_data_res_3__0__1_), .A2(
        npu_inst_pe_1_2_0_n1), .B1(npu_inst_pe_1_2_0_N74), .B2(
        npu_inst_pe_1_2_0_n76), .C1(npu_inst_pe_1_2_0_N66), .C2(
        npu_inst_pe_1_2_0_n77), .ZN(npu_inst_pe_1_2_0_n83) );
  INV_X1 npu_inst_pe_1_2_0_U46 ( .A(npu_inst_pe_1_2_0_n83), .ZN(
        npu_inst_pe_1_2_0_n99) );
  AOI222_X1 npu_inst_pe_1_2_0_U45 ( .A1(npu_inst_int_data_res_3__0__2_), .A2(
        npu_inst_pe_1_2_0_n1), .B1(npu_inst_pe_1_2_0_N75), .B2(
        npu_inst_pe_1_2_0_n76), .C1(npu_inst_pe_1_2_0_N67), .C2(
        npu_inst_pe_1_2_0_n77), .ZN(npu_inst_pe_1_2_0_n82) );
  INV_X1 npu_inst_pe_1_2_0_U44 ( .A(npu_inst_pe_1_2_0_n82), .ZN(
        npu_inst_pe_1_2_0_n98) );
  AOI222_X1 npu_inst_pe_1_2_0_U43 ( .A1(npu_inst_int_data_res_3__0__3_), .A2(
        npu_inst_pe_1_2_0_n1), .B1(npu_inst_pe_1_2_0_N76), .B2(
        npu_inst_pe_1_2_0_n76), .C1(npu_inst_pe_1_2_0_N68), .C2(
        npu_inst_pe_1_2_0_n77), .ZN(npu_inst_pe_1_2_0_n81) );
  INV_X1 npu_inst_pe_1_2_0_U42 ( .A(npu_inst_pe_1_2_0_n81), .ZN(
        npu_inst_pe_1_2_0_n36) );
  AOI222_X1 npu_inst_pe_1_2_0_U41 ( .A1(npu_inst_int_data_res_3__0__4_), .A2(
        npu_inst_pe_1_2_0_n1), .B1(npu_inst_pe_1_2_0_N77), .B2(
        npu_inst_pe_1_2_0_n76), .C1(npu_inst_pe_1_2_0_N69), .C2(
        npu_inst_pe_1_2_0_n77), .ZN(npu_inst_pe_1_2_0_n80) );
  INV_X1 npu_inst_pe_1_2_0_U40 ( .A(npu_inst_pe_1_2_0_n80), .ZN(
        npu_inst_pe_1_2_0_n35) );
  AOI222_X1 npu_inst_pe_1_2_0_U39 ( .A1(npu_inst_int_data_res_3__0__5_), .A2(
        npu_inst_pe_1_2_0_n1), .B1(npu_inst_pe_1_2_0_N78), .B2(
        npu_inst_pe_1_2_0_n76), .C1(npu_inst_pe_1_2_0_N70), .C2(
        npu_inst_pe_1_2_0_n77), .ZN(npu_inst_pe_1_2_0_n79) );
  INV_X1 npu_inst_pe_1_2_0_U38 ( .A(npu_inst_pe_1_2_0_n79), .ZN(
        npu_inst_pe_1_2_0_n34) );
  AOI222_X1 npu_inst_pe_1_2_0_U37 ( .A1(npu_inst_int_data_res_3__0__6_), .A2(
        npu_inst_pe_1_2_0_n1), .B1(npu_inst_pe_1_2_0_N79), .B2(
        npu_inst_pe_1_2_0_n76), .C1(npu_inst_pe_1_2_0_N71), .C2(
        npu_inst_pe_1_2_0_n77), .ZN(npu_inst_pe_1_2_0_n78) );
  INV_X1 npu_inst_pe_1_2_0_U36 ( .A(npu_inst_pe_1_2_0_n78), .ZN(
        npu_inst_pe_1_2_0_n33) );
  AND2_X1 npu_inst_pe_1_2_0_U35 ( .A1(npu_inst_pe_1_2_0_o_data_h_1_), .A2(
        npu_inst_pe_1_2_0_int_q_weight_1_), .ZN(npu_inst_pe_1_2_0_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_2_0_U34 ( .A1(npu_inst_pe_1_2_0_o_data_h_0_), .A2(
        npu_inst_pe_1_2_0_int_q_weight_1_), .ZN(npu_inst_pe_1_2_0_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_2_0_U33 ( .A(npu_inst_pe_1_2_0_int_data_1_), .ZN(
        npu_inst_pe_1_2_0_n13) );
  AOI22_X1 npu_inst_pe_1_2_0_U32 ( .A1(npu_inst_n58), .A2(
        npu_inst_int_data_y_3__0__1_), .B1(npu_inst_pe_1_2_0_n3), .B2(
        npu_inst_int_data_x_2__1__1_), .ZN(npu_inst_pe_1_2_0_n63) );
  AOI22_X1 npu_inst_pe_1_2_0_U31 ( .A1(npu_inst_n58), .A2(
        npu_inst_int_data_y_3__0__0_), .B1(npu_inst_pe_1_2_0_n3), .B2(
        npu_inst_int_data_x_2__1__0_), .ZN(npu_inst_pe_1_2_0_n61) );
  INV_X1 npu_inst_pe_1_2_0_U30 ( .A(npu_inst_pe_1_2_0_int_data_0_), .ZN(
        npu_inst_pe_1_2_0_n12) );
  INV_X1 npu_inst_pe_1_2_0_U29 ( .A(npu_inst_n70), .ZN(npu_inst_pe_1_2_0_n5)
         );
  OR3_X1 npu_inst_pe_1_2_0_U28 ( .A1(npu_inst_n78), .A2(npu_inst_pe_1_2_0_n7), 
        .A3(npu_inst_pe_1_2_0_n5), .ZN(npu_inst_pe_1_2_0_n56) );
  OR3_X1 npu_inst_pe_1_2_0_U27 ( .A1(npu_inst_pe_1_2_0_n5), .A2(
        npu_inst_pe_1_2_0_n7), .A3(npu_inst_pe_1_2_0_n6), .ZN(
        npu_inst_pe_1_2_0_n48) );
  INV_X1 npu_inst_pe_1_2_0_U26 ( .A(npu_inst_pe_1_2_0_n5), .ZN(
        npu_inst_pe_1_2_0_n4) );
  INV_X1 npu_inst_pe_1_2_0_U25 ( .A(npu_inst_n125), .ZN(npu_inst_pe_1_2_0_n11)
         );
  OR3_X1 npu_inst_pe_1_2_0_U24 ( .A1(npu_inst_pe_1_2_0_n4), .A2(
        npu_inst_pe_1_2_0_n7), .A3(npu_inst_pe_1_2_0_n6), .ZN(
        npu_inst_pe_1_2_0_n52) );
  OR3_X1 npu_inst_pe_1_2_0_U23 ( .A1(npu_inst_n78), .A2(npu_inst_pe_1_2_0_n7), 
        .A3(npu_inst_pe_1_2_0_n4), .ZN(npu_inst_pe_1_2_0_n60) );
  NOR2_X1 npu_inst_pe_1_2_0_U22 ( .A1(npu_inst_pe_1_2_0_n60), .A2(
        npu_inst_pe_1_2_0_n3), .ZN(npu_inst_pe_1_2_0_n58) );
  NOR2_X1 npu_inst_pe_1_2_0_U21 ( .A1(npu_inst_pe_1_2_0_n56), .A2(
        npu_inst_pe_1_2_0_n3), .ZN(npu_inst_pe_1_2_0_n54) );
  NOR2_X1 npu_inst_pe_1_2_0_U20 ( .A1(npu_inst_pe_1_2_0_n52), .A2(
        npu_inst_pe_1_2_0_n3), .ZN(npu_inst_pe_1_2_0_n50) );
  NOR2_X1 npu_inst_pe_1_2_0_U19 ( .A1(npu_inst_pe_1_2_0_n48), .A2(
        npu_inst_pe_1_2_0_n3), .ZN(npu_inst_pe_1_2_0_n46) );
  NOR2_X1 npu_inst_pe_1_2_0_U18 ( .A1(npu_inst_pe_1_2_0_n40), .A2(
        npu_inst_pe_1_2_0_n3), .ZN(npu_inst_pe_1_2_0_n38) );
  NOR2_X1 npu_inst_pe_1_2_0_U17 ( .A1(npu_inst_pe_1_2_0_n44), .A2(
        npu_inst_pe_1_2_0_n3), .ZN(npu_inst_pe_1_2_0_n42) );
  BUF_X1 npu_inst_pe_1_2_0_U16 ( .A(npu_inst_n103), .Z(npu_inst_pe_1_2_0_n7)
         );
  BUF_X1 npu_inst_pe_1_2_0_U15 ( .A(npu_inst_pe_1_2_0_n11), .Z(
        npu_inst_pe_1_2_0_n10) );
  BUF_X1 npu_inst_pe_1_2_0_U14 ( .A(npu_inst_pe_1_2_0_n11), .Z(
        npu_inst_pe_1_2_0_n9) );
  BUF_X1 npu_inst_pe_1_2_0_U13 ( .A(npu_inst_pe_1_2_0_n11), .Z(
        npu_inst_pe_1_2_0_n8) );
  INV_X1 npu_inst_pe_1_2_0_U12 ( .A(npu_inst_pe_1_2_0_n38), .ZN(
        npu_inst_pe_1_2_0_n117) );
  INV_X1 npu_inst_pe_1_2_0_U11 ( .A(npu_inst_pe_1_2_0_n58), .ZN(
        npu_inst_pe_1_2_0_n113) );
  INV_X1 npu_inst_pe_1_2_0_U10 ( .A(npu_inst_pe_1_2_0_n54), .ZN(
        npu_inst_pe_1_2_0_n114) );
  INV_X1 npu_inst_pe_1_2_0_U9 ( .A(npu_inst_pe_1_2_0_n50), .ZN(
        npu_inst_pe_1_2_0_n115) );
  INV_X1 npu_inst_pe_1_2_0_U8 ( .A(npu_inst_pe_1_2_0_n46), .ZN(
        npu_inst_pe_1_2_0_n116) );
  INV_X1 npu_inst_pe_1_2_0_U7 ( .A(npu_inst_pe_1_2_0_n42), .ZN(
        npu_inst_pe_1_2_0_n118) );
  BUF_X1 npu_inst_pe_1_2_0_U6 ( .A(npu_inst_n30), .Z(npu_inst_pe_1_2_0_n2) );
  BUF_X1 npu_inst_pe_1_2_0_U5 ( .A(npu_inst_n30), .Z(npu_inst_pe_1_2_0_n1) );
  NOR2_X1 npu_inst_pe_1_2_0_U4 ( .A1(npu_inst_pe_1_2_0_int_q_weight_0_), .A2(
        npu_inst_pe_1_2_0_n1), .ZN(npu_inst_pe_1_2_0_n76) );
  NOR2_X1 npu_inst_pe_1_2_0_U3 ( .A1(npu_inst_pe_1_2_0_n27), .A2(
        npu_inst_pe_1_2_0_n1), .ZN(npu_inst_pe_1_2_0_n77) );
  FA_X1 npu_inst_pe_1_2_0_sub_77_U2_1 ( .A(npu_inst_pe_1_2_0_int_q_acc_1_), 
        .B(npu_inst_pe_1_2_0_n13), .CI(npu_inst_pe_1_2_0_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_2_0_sub_77_carry_2_), .S(npu_inst_pe_1_2_0_N66) );
  FA_X1 npu_inst_pe_1_2_0_add_79_U1_1 ( .A(npu_inst_pe_1_2_0_int_q_acc_1_), 
        .B(npu_inst_pe_1_2_0_int_data_1_), .CI(
        npu_inst_pe_1_2_0_add_79_carry_1_), .CO(
        npu_inst_pe_1_2_0_add_79_carry_2_), .S(npu_inst_pe_1_2_0_N74) );
  NAND3_X1 npu_inst_pe_1_2_0_U109 ( .A1(npu_inst_pe_1_2_0_n5), .A2(
        npu_inst_pe_1_2_0_n6), .A3(npu_inst_pe_1_2_0_n7), .ZN(
        npu_inst_pe_1_2_0_n44) );
  NAND3_X1 npu_inst_pe_1_2_0_U108 ( .A1(npu_inst_pe_1_2_0_n4), .A2(
        npu_inst_pe_1_2_0_n6), .A3(npu_inst_pe_1_2_0_n7), .ZN(
        npu_inst_pe_1_2_0_n40) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_2_0_n33), .CK(
        npu_inst_pe_1_2_0_net3925), .RN(npu_inst_pe_1_2_0_n8), .Q(
        npu_inst_pe_1_2_0_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_2_0_n34), .CK(
        npu_inst_pe_1_2_0_net3925), .RN(npu_inst_pe_1_2_0_n8), .Q(
        npu_inst_pe_1_2_0_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_2_0_n35), .CK(
        npu_inst_pe_1_2_0_net3925), .RN(npu_inst_pe_1_2_0_n8), .Q(
        npu_inst_pe_1_2_0_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_2_0_n36), .CK(
        npu_inst_pe_1_2_0_net3925), .RN(npu_inst_pe_1_2_0_n8), .Q(
        npu_inst_pe_1_2_0_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_2_0_n98), .CK(
        npu_inst_pe_1_2_0_net3925), .RN(npu_inst_pe_1_2_0_n8), .Q(
        npu_inst_pe_1_2_0_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_2_0_n99), .CK(
        npu_inst_pe_1_2_0_net3925), .RN(npu_inst_pe_1_2_0_n8), .Q(
        npu_inst_pe_1_2_0_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_2_0_n32), .CK(
        npu_inst_pe_1_2_0_net3925), .RN(npu_inst_pe_1_2_0_n8), .Q(
        npu_inst_pe_1_2_0_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_2_0_n100), 
        .CK(npu_inst_pe_1_2_0_net3925), .RN(npu_inst_pe_1_2_0_n8), .Q(
        npu_inst_pe_1_2_0_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_weight_reg_0_ ( .D(npu_inst_n111), .CK(
        npu_inst_pe_1_2_0_net3931), .RN(npu_inst_pe_1_2_0_n8), .Q(
        npu_inst_pe_1_2_0_int_q_weight_0_), .QN(npu_inst_pe_1_2_0_n27) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_weight_reg_1_ ( .D(npu_inst_n117), .CK(
        npu_inst_pe_1_2_0_net3931), .RN(npu_inst_pe_1_2_0_n8), .Q(
        npu_inst_pe_1_2_0_int_q_weight_1_), .QN(npu_inst_pe_1_2_0_n26) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_2_0_n112), 
        .CK(npu_inst_pe_1_2_0_net3931), .RN(npu_inst_pe_1_2_0_n8), .Q(
        npu_inst_pe_1_2_0_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_2_0_n106), 
        .CK(npu_inst_pe_1_2_0_net3931), .RN(npu_inst_pe_1_2_0_n8), .Q(
        npu_inst_pe_1_2_0_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_2_0_n111), 
        .CK(npu_inst_pe_1_2_0_net3931), .RN(npu_inst_pe_1_2_0_n9), .Q(
        npu_inst_pe_1_2_0_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_2_0_n105), 
        .CK(npu_inst_pe_1_2_0_net3931), .RN(npu_inst_pe_1_2_0_n9), .Q(
        npu_inst_pe_1_2_0_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_2_0_n110), 
        .CK(npu_inst_pe_1_2_0_net3931), .RN(npu_inst_pe_1_2_0_n9), .Q(
        npu_inst_pe_1_2_0_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_2_0_n104), 
        .CK(npu_inst_pe_1_2_0_net3931), .RN(npu_inst_pe_1_2_0_n9), .Q(
        npu_inst_pe_1_2_0_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_2_0_n109), 
        .CK(npu_inst_pe_1_2_0_net3931), .RN(npu_inst_pe_1_2_0_n9), .Q(
        npu_inst_pe_1_2_0_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_2_0_n103), 
        .CK(npu_inst_pe_1_2_0_net3931), .RN(npu_inst_pe_1_2_0_n9), .Q(
        npu_inst_pe_1_2_0_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_2_0_n108), 
        .CK(npu_inst_pe_1_2_0_net3931), .RN(npu_inst_pe_1_2_0_n9), .Q(
        npu_inst_pe_1_2_0_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_2_0_n102), 
        .CK(npu_inst_pe_1_2_0_net3931), .RN(npu_inst_pe_1_2_0_n9), .Q(
        npu_inst_pe_1_2_0_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_2_0_n107), 
        .CK(npu_inst_pe_1_2_0_net3931), .RN(npu_inst_pe_1_2_0_n9), .Q(
        npu_inst_pe_1_2_0_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_2_0_n101), 
        .CK(npu_inst_pe_1_2_0_net3931), .RN(npu_inst_pe_1_2_0_n9), .Q(
        npu_inst_pe_1_2_0_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_2_0_n86), 
        .CK(npu_inst_pe_1_2_0_net3931), .RN(npu_inst_pe_1_2_0_n9), .Q(
        npu_inst_pe_1_2_0_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_2_0_n87), 
        .CK(npu_inst_pe_1_2_0_net3931), .RN(npu_inst_pe_1_2_0_n9), .Q(
        npu_inst_pe_1_2_0_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_2_0_n88), 
        .CK(npu_inst_pe_1_2_0_net3931), .RN(npu_inst_pe_1_2_0_n10), .Q(
        npu_inst_pe_1_2_0_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_2_0_n89), 
        .CK(npu_inst_pe_1_2_0_net3931), .RN(npu_inst_pe_1_2_0_n10), .Q(
        npu_inst_pe_1_2_0_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_2_0_n90), 
        .CK(npu_inst_pe_1_2_0_net3931), .RN(npu_inst_pe_1_2_0_n10), .Q(
        npu_inst_pe_1_2_0_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_2_0_n91), 
        .CK(npu_inst_pe_1_2_0_net3931), .RN(npu_inst_pe_1_2_0_n10), .Q(
        npu_inst_pe_1_2_0_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_2_0_n92), 
        .CK(npu_inst_pe_1_2_0_net3931), .RN(npu_inst_pe_1_2_0_n10), .Q(
        npu_inst_pe_1_2_0_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_2_0_n93), 
        .CK(npu_inst_pe_1_2_0_net3931), .RN(npu_inst_pe_1_2_0_n10), .Q(
        npu_inst_pe_1_2_0_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_2_0_n94), 
        .CK(npu_inst_pe_1_2_0_net3931), .RN(npu_inst_pe_1_2_0_n10), .Q(
        npu_inst_pe_1_2_0_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_2_0_n95), 
        .CK(npu_inst_pe_1_2_0_net3931), .RN(npu_inst_pe_1_2_0_n10), .Q(
        npu_inst_pe_1_2_0_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_2_0_n96), 
        .CK(npu_inst_pe_1_2_0_net3931), .RN(npu_inst_pe_1_2_0_n10), .Q(
        npu_inst_pe_1_2_0_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_2_0_n97), 
        .CK(npu_inst_pe_1_2_0_net3931), .RN(npu_inst_pe_1_2_0_n10), .Q(
        npu_inst_pe_1_2_0_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_2_0_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_2_0_N84), .SE(1'b0), .GCK(npu_inst_pe_1_2_0_net3925) );
  CLKGATETST_X1 npu_inst_pe_1_2_0_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n65), .SE(1'b0), .GCK(npu_inst_pe_1_2_0_net3931) );
  MUX2_X1 npu_inst_pe_1_2_1_U162 ( .A(npu_inst_pe_1_2_1_n32), .B(
        npu_inst_pe_1_2_1_n29), .S(npu_inst_pe_1_2_1_n8), .Z(
        npu_inst_pe_1_2_1_N93) );
  MUX2_X1 npu_inst_pe_1_2_1_U161 ( .A(npu_inst_pe_1_2_1_n31), .B(
        npu_inst_pe_1_2_1_n30), .S(npu_inst_pe_1_2_1_n6), .Z(
        npu_inst_pe_1_2_1_n32) );
  MUX2_X1 npu_inst_pe_1_2_1_U160 ( .A(npu_inst_pe_1_2_1_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_2_1_int_q_reg_v_1__0_), .S(npu_inst_pe_1_2_1_n4), .Z(
        npu_inst_pe_1_2_1_n31) );
  MUX2_X1 npu_inst_pe_1_2_1_U159 ( .A(npu_inst_pe_1_2_1_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_2_1_int_q_reg_v_3__0_), .S(npu_inst_pe_1_2_1_n4), .Z(
        npu_inst_pe_1_2_1_n30) );
  MUX2_X1 npu_inst_pe_1_2_1_U158 ( .A(npu_inst_pe_1_2_1_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_2_1_int_q_reg_v_5__0_), .S(npu_inst_pe_1_2_1_n4), .Z(
        npu_inst_pe_1_2_1_n29) );
  MUX2_X1 npu_inst_pe_1_2_1_U157 ( .A(npu_inst_pe_1_2_1_n28), .B(
        npu_inst_pe_1_2_1_n23), .S(npu_inst_pe_1_2_1_n8), .Z(
        npu_inst_pe_1_2_1_N94) );
  MUX2_X1 npu_inst_pe_1_2_1_U156 ( .A(npu_inst_pe_1_2_1_n25), .B(
        npu_inst_pe_1_2_1_n24), .S(npu_inst_pe_1_2_1_n6), .Z(
        npu_inst_pe_1_2_1_n28) );
  MUX2_X1 npu_inst_pe_1_2_1_U155 ( .A(npu_inst_pe_1_2_1_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_2_1_int_q_reg_v_1__1_), .S(npu_inst_pe_1_2_1_n4), .Z(
        npu_inst_pe_1_2_1_n25) );
  MUX2_X1 npu_inst_pe_1_2_1_U154 ( .A(npu_inst_pe_1_2_1_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_2_1_int_q_reg_v_3__1_), .S(npu_inst_pe_1_2_1_n4), .Z(
        npu_inst_pe_1_2_1_n24) );
  MUX2_X1 npu_inst_pe_1_2_1_U153 ( .A(npu_inst_pe_1_2_1_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_2_1_int_q_reg_v_5__1_), .S(npu_inst_pe_1_2_1_n4), .Z(
        npu_inst_pe_1_2_1_n23) );
  MUX2_X1 npu_inst_pe_1_2_1_U152 ( .A(npu_inst_pe_1_2_1_n22), .B(
        npu_inst_pe_1_2_1_n19), .S(npu_inst_pe_1_2_1_n8), .Z(
        npu_inst_int_data_x_2__1__1_) );
  MUX2_X1 npu_inst_pe_1_2_1_U151 ( .A(npu_inst_pe_1_2_1_n21), .B(
        npu_inst_pe_1_2_1_n20), .S(npu_inst_pe_1_2_1_n6), .Z(
        npu_inst_pe_1_2_1_n22) );
  MUX2_X1 npu_inst_pe_1_2_1_U150 ( .A(npu_inst_pe_1_2_1_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_2_1_int_q_reg_h_1__1_), .S(npu_inst_pe_1_2_1_n4), .Z(
        npu_inst_pe_1_2_1_n21) );
  MUX2_X1 npu_inst_pe_1_2_1_U149 ( .A(npu_inst_pe_1_2_1_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_2_1_int_q_reg_h_3__1_), .S(npu_inst_pe_1_2_1_n4), .Z(
        npu_inst_pe_1_2_1_n20) );
  MUX2_X1 npu_inst_pe_1_2_1_U148 ( .A(npu_inst_pe_1_2_1_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_2_1_int_q_reg_h_5__1_), .S(npu_inst_pe_1_2_1_n4), .Z(
        npu_inst_pe_1_2_1_n19) );
  MUX2_X1 npu_inst_pe_1_2_1_U147 ( .A(npu_inst_pe_1_2_1_n18), .B(
        npu_inst_pe_1_2_1_n15), .S(npu_inst_pe_1_2_1_n8), .Z(
        npu_inst_int_data_x_2__1__0_) );
  MUX2_X1 npu_inst_pe_1_2_1_U146 ( .A(npu_inst_pe_1_2_1_n17), .B(
        npu_inst_pe_1_2_1_n16), .S(npu_inst_pe_1_2_1_n6), .Z(
        npu_inst_pe_1_2_1_n18) );
  MUX2_X1 npu_inst_pe_1_2_1_U145 ( .A(npu_inst_pe_1_2_1_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_2_1_int_q_reg_h_1__0_), .S(npu_inst_pe_1_2_1_n4), .Z(
        npu_inst_pe_1_2_1_n17) );
  MUX2_X1 npu_inst_pe_1_2_1_U144 ( .A(npu_inst_pe_1_2_1_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_2_1_int_q_reg_h_3__0_), .S(npu_inst_pe_1_2_1_n4), .Z(
        npu_inst_pe_1_2_1_n16) );
  MUX2_X1 npu_inst_pe_1_2_1_U143 ( .A(npu_inst_pe_1_2_1_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_2_1_int_q_reg_h_5__0_), .S(npu_inst_pe_1_2_1_n4), .Z(
        npu_inst_pe_1_2_1_n15) );
  XOR2_X1 npu_inst_pe_1_2_1_U142 ( .A(npu_inst_pe_1_2_1_int_data_0_), .B(
        npu_inst_pe_1_2_1_int_q_acc_0_), .Z(npu_inst_pe_1_2_1_N73) );
  AND2_X1 npu_inst_pe_1_2_1_U141 ( .A1(npu_inst_pe_1_2_1_int_q_acc_0_), .A2(
        npu_inst_pe_1_2_1_int_data_0_), .ZN(npu_inst_pe_1_2_1_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_2_1_U140 ( .A(npu_inst_pe_1_2_1_int_q_acc_0_), .B(
        npu_inst_pe_1_2_1_n13), .ZN(npu_inst_pe_1_2_1_N65) );
  OR2_X1 npu_inst_pe_1_2_1_U139 ( .A1(npu_inst_pe_1_2_1_n13), .A2(
        npu_inst_pe_1_2_1_int_q_acc_0_), .ZN(npu_inst_pe_1_2_1_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_2_1_U138 ( .A(npu_inst_pe_1_2_1_int_q_acc_2_), .B(
        npu_inst_pe_1_2_1_add_79_carry_2_), .Z(npu_inst_pe_1_2_1_N75) );
  AND2_X1 npu_inst_pe_1_2_1_U137 ( .A1(npu_inst_pe_1_2_1_add_79_carry_2_), 
        .A2(npu_inst_pe_1_2_1_int_q_acc_2_), .ZN(
        npu_inst_pe_1_2_1_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_2_1_U136 ( .A(npu_inst_pe_1_2_1_int_q_acc_3_), .B(
        npu_inst_pe_1_2_1_add_79_carry_3_), .Z(npu_inst_pe_1_2_1_N76) );
  AND2_X1 npu_inst_pe_1_2_1_U135 ( .A1(npu_inst_pe_1_2_1_add_79_carry_3_), 
        .A2(npu_inst_pe_1_2_1_int_q_acc_3_), .ZN(
        npu_inst_pe_1_2_1_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_2_1_U134 ( .A(npu_inst_pe_1_2_1_int_q_acc_4_), .B(
        npu_inst_pe_1_2_1_add_79_carry_4_), .Z(npu_inst_pe_1_2_1_N77) );
  AND2_X1 npu_inst_pe_1_2_1_U133 ( .A1(npu_inst_pe_1_2_1_add_79_carry_4_), 
        .A2(npu_inst_pe_1_2_1_int_q_acc_4_), .ZN(
        npu_inst_pe_1_2_1_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_2_1_U132 ( .A(npu_inst_pe_1_2_1_int_q_acc_5_), .B(
        npu_inst_pe_1_2_1_add_79_carry_5_), .Z(npu_inst_pe_1_2_1_N78) );
  AND2_X1 npu_inst_pe_1_2_1_U131 ( .A1(npu_inst_pe_1_2_1_add_79_carry_5_), 
        .A2(npu_inst_pe_1_2_1_int_q_acc_5_), .ZN(
        npu_inst_pe_1_2_1_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_2_1_U130 ( .A(npu_inst_pe_1_2_1_int_q_acc_6_), .B(
        npu_inst_pe_1_2_1_add_79_carry_6_), .Z(npu_inst_pe_1_2_1_N79) );
  AND2_X1 npu_inst_pe_1_2_1_U129 ( .A1(npu_inst_pe_1_2_1_add_79_carry_6_), 
        .A2(npu_inst_pe_1_2_1_int_q_acc_6_), .ZN(
        npu_inst_pe_1_2_1_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_2_1_U128 ( .A(npu_inst_pe_1_2_1_int_q_acc_7_), .B(
        npu_inst_pe_1_2_1_add_79_carry_7_), .Z(npu_inst_pe_1_2_1_N80) );
  XNOR2_X1 npu_inst_pe_1_2_1_U127 ( .A(npu_inst_pe_1_2_1_sub_77_carry_2_), .B(
        npu_inst_pe_1_2_1_int_q_acc_2_), .ZN(npu_inst_pe_1_2_1_N67) );
  OR2_X1 npu_inst_pe_1_2_1_U126 ( .A1(npu_inst_pe_1_2_1_int_q_acc_2_), .A2(
        npu_inst_pe_1_2_1_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_2_1_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_2_1_U125 ( .A(npu_inst_pe_1_2_1_sub_77_carry_3_), .B(
        npu_inst_pe_1_2_1_int_q_acc_3_), .ZN(npu_inst_pe_1_2_1_N68) );
  OR2_X1 npu_inst_pe_1_2_1_U124 ( .A1(npu_inst_pe_1_2_1_int_q_acc_3_), .A2(
        npu_inst_pe_1_2_1_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_2_1_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_2_1_U123 ( .A(npu_inst_pe_1_2_1_sub_77_carry_4_), .B(
        npu_inst_pe_1_2_1_int_q_acc_4_), .ZN(npu_inst_pe_1_2_1_N69) );
  OR2_X1 npu_inst_pe_1_2_1_U122 ( .A1(npu_inst_pe_1_2_1_int_q_acc_4_), .A2(
        npu_inst_pe_1_2_1_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_2_1_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_2_1_U121 ( .A(npu_inst_pe_1_2_1_sub_77_carry_5_), .B(
        npu_inst_pe_1_2_1_int_q_acc_5_), .ZN(npu_inst_pe_1_2_1_N70) );
  OR2_X1 npu_inst_pe_1_2_1_U120 ( .A1(npu_inst_pe_1_2_1_int_q_acc_5_), .A2(
        npu_inst_pe_1_2_1_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_2_1_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_2_1_U119 ( .A(npu_inst_pe_1_2_1_sub_77_carry_6_), .B(
        npu_inst_pe_1_2_1_int_q_acc_6_), .ZN(npu_inst_pe_1_2_1_N71) );
  OR2_X1 npu_inst_pe_1_2_1_U118 ( .A1(npu_inst_pe_1_2_1_int_q_acc_6_), .A2(
        npu_inst_pe_1_2_1_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_2_1_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_2_1_U117 ( .A(npu_inst_pe_1_2_1_int_q_acc_7_), .B(
        npu_inst_pe_1_2_1_sub_77_carry_7_), .ZN(npu_inst_pe_1_2_1_N72) );
  INV_X1 npu_inst_pe_1_2_1_U116 ( .A(npu_inst_n78), .ZN(npu_inst_pe_1_2_1_n7)
         );
  INV_X1 npu_inst_pe_1_2_1_U115 ( .A(npu_inst_pe_1_2_1_n7), .ZN(
        npu_inst_pe_1_2_1_n6) );
  INV_X1 npu_inst_pe_1_2_1_U114 ( .A(npu_inst_n58), .ZN(npu_inst_pe_1_2_1_n3)
         );
  AOI22_X1 npu_inst_pe_1_2_1_U113 ( .A1(npu_inst_int_data_y_3__1__0_), .A2(
        npu_inst_pe_1_2_1_n58), .B1(npu_inst_pe_1_2_1_n114), .B2(
        npu_inst_pe_1_2_1_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_2_1_n57) );
  INV_X1 npu_inst_pe_1_2_1_U112 ( .A(npu_inst_pe_1_2_1_n57), .ZN(
        npu_inst_pe_1_2_1_n108) );
  AOI22_X1 npu_inst_pe_1_2_1_U111 ( .A1(npu_inst_int_data_y_3__1__0_), .A2(
        npu_inst_pe_1_2_1_n54), .B1(npu_inst_pe_1_2_1_n115), .B2(
        npu_inst_pe_1_2_1_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_2_1_n53) );
  INV_X1 npu_inst_pe_1_2_1_U110 ( .A(npu_inst_pe_1_2_1_n53), .ZN(
        npu_inst_pe_1_2_1_n109) );
  AOI22_X1 npu_inst_pe_1_2_1_U107 ( .A1(npu_inst_int_data_y_3__1__0_), .A2(
        npu_inst_pe_1_2_1_n50), .B1(npu_inst_pe_1_2_1_n116), .B2(
        npu_inst_pe_1_2_1_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_2_1_n49) );
  INV_X1 npu_inst_pe_1_2_1_U106 ( .A(npu_inst_pe_1_2_1_n49), .ZN(
        npu_inst_pe_1_2_1_n110) );
  AOI22_X1 npu_inst_pe_1_2_1_U105 ( .A1(npu_inst_int_data_y_3__1__0_), .A2(
        npu_inst_pe_1_2_1_n46), .B1(npu_inst_pe_1_2_1_n117), .B2(
        npu_inst_pe_1_2_1_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_2_1_n45) );
  INV_X1 npu_inst_pe_1_2_1_U104 ( .A(npu_inst_pe_1_2_1_n45), .ZN(
        npu_inst_pe_1_2_1_n111) );
  AOI22_X1 npu_inst_pe_1_2_1_U103 ( .A1(npu_inst_int_data_y_3__1__0_), .A2(
        npu_inst_pe_1_2_1_n42), .B1(npu_inst_pe_1_2_1_n119), .B2(
        npu_inst_pe_1_2_1_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_2_1_n41) );
  INV_X1 npu_inst_pe_1_2_1_U102 ( .A(npu_inst_pe_1_2_1_n41), .ZN(
        npu_inst_pe_1_2_1_n112) );
  AOI22_X1 npu_inst_pe_1_2_1_U101 ( .A1(npu_inst_int_data_y_3__1__1_), .A2(
        npu_inst_pe_1_2_1_n58), .B1(npu_inst_pe_1_2_1_n114), .B2(
        npu_inst_pe_1_2_1_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_2_1_n59) );
  INV_X1 npu_inst_pe_1_2_1_U100 ( .A(npu_inst_pe_1_2_1_n59), .ZN(
        npu_inst_pe_1_2_1_n102) );
  AOI22_X1 npu_inst_pe_1_2_1_U99 ( .A1(npu_inst_int_data_y_3__1__1_), .A2(
        npu_inst_pe_1_2_1_n54), .B1(npu_inst_pe_1_2_1_n115), .B2(
        npu_inst_pe_1_2_1_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_2_1_n55) );
  INV_X1 npu_inst_pe_1_2_1_U98 ( .A(npu_inst_pe_1_2_1_n55), .ZN(
        npu_inst_pe_1_2_1_n103) );
  AOI22_X1 npu_inst_pe_1_2_1_U97 ( .A1(npu_inst_int_data_y_3__1__1_), .A2(
        npu_inst_pe_1_2_1_n50), .B1(npu_inst_pe_1_2_1_n116), .B2(
        npu_inst_pe_1_2_1_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_2_1_n51) );
  INV_X1 npu_inst_pe_1_2_1_U96 ( .A(npu_inst_pe_1_2_1_n51), .ZN(
        npu_inst_pe_1_2_1_n104) );
  AOI22_X1 npu_inst_pe_1_2_1_U95 ( .A1(npu_inst_int_data_y_3__1__1_), .A2(
        npu_inst_pe_1_2_1_n46), .B1(npu_inst_pe_1_2_1_n117), .B2(
        npu_inst_pe_1_2_1_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_2_1_n47) );
  INV_X1 npu_inst_pe_1_2_1_U94 ( .A(npu_inst_pe_1_2_1_n47), .ZN(
        npu_inst_pe_1_2_1_n105) );
  AOI22_X1 npu_inst_pe_1_2_1_U93 ( .A1(npu_inst_int_data_y_3__1__1_), .A2(
        npu_inst_pe_1_2_1_n42), .B1(npu_inst_pe_1_2_1_n119), .B2(
        npu_inst_pe_1_2_1_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_2_1_n43) );
  INV_X1 npu_inst_pe_1_2_1_U92 ( .A(npu_inst_pe_1_2_1_n43), .ZN(
        npu_inst_pe_1_2_1_n106) );
  AOI22_X1 npu_inst_pe_1_2_1_U91 ( .A1(npu_inst_pe_1_2_1_n38), .A2(
        npu_inst_int_data_y_3__1__1_), .B1(npu_inst_pe_1_2_1_n118), .B2(
        npu_inst_pe_1_2_1_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_2_1_n39) );
  INV_X1 npu_inst_pe_1_2_1_U90 ( .A(npu_inst_pe_1_2_1_n39), .ZN(
        npu_inst_pe_1_2_1_n107) );
  AOI22_X1 npu_inst_pe_1_2_1_U89 ( .A1(npu_inst_pe_1_2_1_n38), .A2(
        npu_inst_int_data_y_3__1__0_), .B1(npu_inst_pe_1_2_1_n118), .B2(
        npu_inst_pe_1_2_1_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_2_1_n37) );
  INV_X1 npu_inst_pe_1_2_1_U88 ( .A(npu_inst_pe_1_2_1_n37), .ZN(
        npu_inst_pe_1_2_1_n113) );
  NAND2_X1 npu_inst_pe_1_2_1_U87 ( .A1(npu_inst_pe_1_2_1_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_2_1_n60), .ZN(npu_inst_pe_1_2_1_n74) );
  OAI21_X1 npu_inst_pe_1_2_1_U86 ( .B1(npu_inst_pe_1_2_1_n63), .B2(
        npu_inst_pe_1_2_1_n60), .A(npu_inst_pe_1_2_1_n74), .ZN(
        npu_inst_pe_1_2_1_n97) );
  NAND2_X1 npu_inst_pe_1_2_1_U85 ( .A1(npu_inst_pe_1_2_1_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_2_1_n60), .ZN(npu_inst_pe_1_2_1_n73) );
  OAI21_X1 npu_inst_pe_1_2_1_U84 ( .B1(npu_inst_pe_1_2_1_n61), .B2(
        npu_inst_pe_1_2_1_n60), .A(npu_inst_pe_1_2_1_n73), .ZN(
        npu_inst_pe_1_2_1_n96) );
  NAND2_X1 npu_inst_pe_1_2_1_U83 ( .A1(npu_inst_pe_1_2_1_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_2_1_n56), .ZN(npu_inst_pe_1_2_1_n72) );
  OAI21_X1 npu_inst_pe_1_2_1_U82 ( .B1(npu_inst_pe_1_2_1_n63), .B2(
        npu_inst_pe_1_2_1_n56), .A(npu_inst_pe_1_2_1_n72), .ZN(
        npu_inst_pe_1_2_1_n95) );
  NAND2_X1 npu_inst_pe_1_2_1_U81 ( .A1(npu_inst_pe_1_2_1_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_2_1_n56), .ZN(npu_inst_pe_1_2_1_n71) );
  OAI21_X1 npu_inst_pe_1_2_1_U80 ( .B1(npu_inst_pe_1_2_1_n61), .B2(
        npu_inst_pe_1_2_1_n56), .A(npu_inst_pe_1_2_1_n71), .ZN(
        npu_inst_pe_1_2_1_n94) );
  NAND2_X1 npu_inst_pe_1_2_1_U79 ( .A1(npu_inst_pe_1_2_1_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_2_1_n52), .ZN(npu_inst_pe_1_2_1_n70) );
  OAI21_X1 npu_inst_pe_1_2_1_U78 ( .B1(npu_inst_pe_1_2_1_n63), .B2(
        npu_inst_pe_1_2_1_n52), .A(npu_inst_pe_1_2_1_n70), .ZN(
        npu_inst_pe_1_2_1_n93) );
  NAND2_X1 npu_inst_pe_1_2_1_U77 ( .A1(npu_inst_pe_1_2_1_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_2_1_n52), .ZN(npu_inst_pe_1_2_1_n69) );
  OAI21_X1 npu_inst_pe_1_2_1_U76 ( .B1(npu_inst_pe_1_2_1_n61), .B2(
        npu_inst_pe_1_2_1_n52), .A(npu_inst_pe_1_2_1_n69), .ZN(
        npu_inst_pe_1_2_1_n92) );
  NAND2_X1 npu_inst_pe_1_2_1_U75 ( .A1(npu_inst_pe_1_2_1_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_2_1_n48), .ZN(npu_inst_pe_1_2_1_n68) );
  OAI21_X1 npu_inst_pe_1_2_1_U74 ( .B1(npu_inst_pe_1_2_1_n63), .B2(
        npu_inst_pe_1_2_1_n48), .A(npu_inst_pe_1_2_1_n68), .ZN(
        npu_inst_pe_1_2_1_n91) );
  NAND2_X1 npu_inst_pe_1_2_1_U73 ( .A1(npu_inst_pe_1_2_1_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_2_1_n48), .ZN(npu_inst_pe_1_2_1_n67) );
  OAI21_X1 npu_inst_pe_1_2_1_U72 ( .B1(npu_inst_pe_1_2_1_n61), .B2(
        npu_inst_pe_1_2_1_n48), .A(npu_inst_pe_1_2_1_n67), .ZN(
        npu_inst_pe_1_2_1_n90) );
  NAND2_X1 npu_inst_pe_1_2_1_U71 ( .A1(npu_inst_pe_1_2_1_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_2_1_n44), .ZN(npu_inst_pe_1_2_1_n66) );
  OAI21_X1 npu_inst_pe_1_2_1_U70 ( .B1(npu_inst_pe_1_2_1_n63), .B2(
        npu_inst_pe_1_2_1_n44), .A(npu_inst_pe_1_2_1_n66), .ZN(
        npu_inst_pe_1_2_1_n89) );
  NAND2_X1 npu_inst_pe_1_2_1_U69 ( .A1(npu_inst_pe_1_2_1_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_2_1_n44), .ZN(npu_inst_pe_1_2_1_n65) );
  OAI21_X1 npu_inst_pe_1_2_1_U68 ( .B1(npu_inst_pe_1_2_1_n61), .B2(
        npu_inst_pe_1_2_1_n44), .A(npu_inst_pe_1_2_1_n65), .ZN(
        npu_inst_pe_1_2_1_n88) );
  NAND2_X1 npu_inst_pe_1_2_1_U67 ( .A1(npu_inst_pe_1_2_1_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_2_1_n40), .ZN(npu_inst_pe_1_2_1_n64) );
  OAI21_X1 npu_inst_pe_1_2_1_U66 ( .B1(npu_inst_pe_1_2_1_n63), .B2(
        npu_inst_pe_1_2_1_n40), .A(npu_inst_pe_1_2_1_n64), .ZN(
        npu_inst_pe_1_2_1_n87) );
  NAND2_X1 npu_inst_pe_1_2_1_U65 ( .A1(npu_inst_pe_1_2_1_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_2_1_n40), .ZN(npu_inst_pe_1_2_1_n62) );
  OAI21_X1 npu_inst_pe_1_2_1_U64 ( .B1(npu_inst_pe_1_2_1_n61), .B2(
        npu_inst_pe_1_2_1_n40), .A(npu_inst_pe_1_2_1_n62), .ZN(
        npu_inst_pe_1_2_1_n86) );
  AND2_X1 npu_inst_pe_1_2_1_U63 ( .A1(npu_inst_pe_1_2_1_N93), .A2(npu_inst_n58), .ZN(npu_inst_int_data_y_2__1__0_) );
  AND2_X1 npu_inst_pe_1_2_1_U62 ( .A1(npu_inst_n58), .A2(npu_inst_pe_1_2_1_N94), .ZN(npu_inst_int_data_y_2__1__1_) );
  NOR3_X1 npu_inst_pe_1_2_1_U61 ( .A1(npu_inst_pe_1_2_1_n26), .A2(npu_inst_n58), .A3(npu_inst_int_ckg[46]), .ZN(npu_inst_pe_1_2_1_n85) );
  OR2_X1 npu_inst_pe_1_2_1_U60 ( .A1(npu_inst_pe_1_2_1_n85), .A2(
        npu_inst_pe_1_2_1_n2), .ZN(npu_inst_pe_1_2_1_N84) );
  AND2_X1 npu_inst_pe_1_2_1_U59 ( .A1(npu_inst_pe_1_2_1_int_q_acc_0_), .A2(
        npu_inst_pe_1_2_1_n1), .ZN(npu_inst_int_data_res_2__1__0_) );
  AND2_X1 npu_inst_pe_1_2_1_U58 ( .A1(npu_inst_pe_1_2_1_n2), .A2(
        npu_inst_pe_1_2_1_int_q_acc_7_), .ZN(npu_inst_int_data_res_2__1__7_)
         );
  AND2_X1 npu_inst_pe_1_2_1_U57 ( .A1(npu_inst_pe_1_2_1_int_q_acc_1_), .A2(
        npu_inst_pe_1_2_1_n1), .ZN(npu_inst_int_data_res_2__1__1_) );
  AND2_X1 npu_inst_pe_1_2_1_U56 ( .A1(npu_inst_pe_1_2_1_int_q_acc_2_), .A2(
        npu_inst_pe_1_2_1_n1), .ZN(npu_inst_int_data_res_2__1__2_) );
  AND2_X1 npu_inst_pe_1_2_1_U55 ( .A1(npu_inst_pe_1_2_1_int_q_acc_3_), .A2(
        npu_inst_pe_1_2_1_n2), .ZN(npu_inst_int_data_res_2__1__3_) );
  AND2_X1 npu_inst_pe_1_2_1_U54 ( .A1(npu_inst_pe_1_2_1_int_q_acc_4_), .A2(
        npu_inst_pe_1_2_1_n2), .ZN(npu_inst_int_data_res_2__1__4_) );
  AND2_X1 npu_inst_pe_1_2_1_U53 ( .A1(npu_inst_pe_1_2_1_int_q_acc_5_), .A2(
        npu_inst_pe_1_2_1_n2), .ZN(npu_inst_int_data_res_2__1__5_) );
  AND2_X1 npu_inst_pe_1_2_1_U52 ( .A1(npu_inst_pe_1_2_1_int_q_acc_6_), .A2(
        npu_inst_pe_1_2_1_n2), .ZN(npu_inst_int_data_res_2__1__6_) );
  AOI222_X1 npu_inst_pe_1_2_1_U51 ( .A1(npu_inst_int_data_res_3__1__0_), .A2(
        npu_inst_pe_1_2_1_n1), .B1(npu_inst_pe_1_2_1_N73), .B2(
        npu_inst_pe_1_2_1_n76), .C1(npu_inst_pe_1_2_1_N65), .C2(
        npu_inst_pe_1_2_1_n77), .ZN(npu_inst_pe_1_2_1_n84) );
  INV_X1 npu_inst_pe_1_2_1_U50 ( .A(npu_inst_pe_1_2_1_n84), .ZN(
        npu_inst_pe_1_2_1_n101) );
  AOI222_X1 npu_inst_pe_1_2_1_U49 ( .A1(npu_inst_int_data_res_3__1__7_), .A2(
        npu_inst_pe_1_2_1_n1), .B1(npu_inst_pe_1_2_1_N80), .B2(
        npu_inst_pe_1_2_1_n76), .C1(npu_inst_pe_1_2_1_N72), .C2(
        npu_inst_pe_1_2_1_n77), .ZN(npu_inst_pe_1_2_1_n75) );
  INV_X1 npu_inst_pe_1_2_1_U48 ( .A(npu_inst_pe_1_2_1_n75), .ZN(
        npu_inst_pe_1_2_1_n33) );
  AOI222_X1 npu_inst_pe_1_2_1_U47 ( .A1(npu_inst_int_data_res_3__1__1_), .A2(
        npu_inst_pe_1_2_1_n1), .B1(npu_inst_pe_1_2_1_N74), .B2(
        npu_inst_pe_1_2_1_n76), .C1(npu_inst_pe_1_2_1_N66), .C2(
        npu_inst_pe_1_2_1_n77), .ZN(npu_inst_pe_1_2_1_n83) );
  INV_X1 npu_inst_pe_1_2_1_U46 ( .A(npu_inst_pe_1_2_1_n83), .ZN(
        npu_inst_pe_1_2_1_n100) );
  AOI222_X1 npu_inst_pe_1_2_1_U45 ( .A1(npu_inst_int_data_res_3__1__2_), .A2(
        npu_inst_pe_1_2_1_n1), .B1(npu_inst_pe_1_2_1_N75), .B2(
        npu_inst_pe_1_2_1_n76), .C1(npu_inst_pe_1_2_1_N67), .C2(
        npu_inst_pe_1_2_1_n77), .ZN(npu_inst_pe_1_2_1_n82) );
  INV_X1 npu_inst_pe_1_2_1_U44 ( .A(npu_inst_pe_1_2_1_n82), .ZN(
        npu_inst_pe_1_2_1_n99) );
  AOI222_X1 npu_inst_pe_1_2_1_U43 ( .A1(npu_inst_int_data_res_3__1__3_), .A2(
        npu_inst_pe_1_2_1_n1), .B1(npu_inst_pe_1_2_1_N76), .B2(
        npu_inst_pe_1_2_1_n76), .C1(npu_inst_pe_1_2_1_N68), .C2(
        npu_inst_pe_1_2_1_n77), .ZN(npu_inst_pe_1_2_1_n81) );
  INV_X1 npu_inst_pe_1_2_1_U42 ( .A(npu_inst_pe_1_2_1_n81), .ZN(
        npu_inst_pe_1_2_1_n98) );
  AOI222_X1 npu_inst_pe_1_2_1_U41 ( .A1(npu_inst_int_data_res_3__1__4_), .A2(
        npu_inst_pe_1_2_1_n1), .B1(npu_inst_pe_1_2_1_N77), .B2(
        npu_inst_pe_1_2_1_n76), .C1(npu_inst_pe_1_2_1_N69), .C2(
        npu_inst_pe_1_2_1_n77), .ZN(npu_inst_pe_1_2_1_n80) );
  INV_X1 npu_inst_pe_1_2_1_U40 ( .A(npu_inst_pe_1_2_1_n80), .ZN(
        npu_inst_pe_1_2_1_n36) );
  AOI222_X1 npu_inst_pe_1_2_1_U39 ( .A1(npu_inst_int_data_res_3__1__5_), .A2(
        npu_inst_pe_1_2_1_n1), .B1(npu_inst_pe_1_2_1_N78), .B2(
        npu_inst_pe_1_2_1_n76), .C1(npu_inst_pe_1_2_1_N70), .C2(
        npu_inst_pe_1_2_1_n77), .ZN(npu_inst_pe_1_2_1_n79) );
  INV_X1 npu_inst_pe_1_2_1_U38 ( .A(npu_inst_pe_1_2_1_n79), .ZN(
        npu_inst_pe_1_2_1_n35) );
  AOI222_X1 npu_inst_pe_1_2_1_U37 ( .A1(npu_inst_int_data_res_3__1__6_), .A2(
        npu_inst_pe_1_2_1_n1), .B1(npu_inst_pe_1_2_1_N79), .B2(
        npu_inst_pe_1_2_1_n76), .C1(npu_inst_pe_1_2_1_N71), .C2(
        npu_inst_pe_1_2_1_n77), .ZN(npu_inst_pe_1_2_1_n78) );
  INV_X1 npu_inst_pe_1_2_1_U36 ( .A(npu_inst_pe_1_2_1_n78), .ZN(
        npu_inst_pe_1_2_1_n34) );
  INV_X1 npu_inst_pe_1_2_1_U35 ( .A(npu_inst_pe_1_2_1_int_data_1_), .ZN(
        npu_inst_pe_1_2_1_n14) );
  AND2_X1 npu_inst_pe_1_2_1_U34 ( .A1(npu_inst_int_data_x_2__1__1_), .A2(
        npu_inst_pe_1_2_1_int_q_weight_1_), .ZN(npu_inst_pe_1_2_1_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_2_1_U33 ( .A1(npu_inst_int_data_x_2__1__0_), .A2(
        npu_inst_pe_1_2_1_int_q_weight_1_), .ZN(npu_inst_pe_1_2_1_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_2_1_U32 ( .A1(npu_inst_n58), .A2(
        npu_inst_int_data_y_3__1__1_), .B1(npu_inst_pe_1_2_1_n3), .B2(
        npu_inst_int_data_x_2__2__1_), .ZN(npu_inst_pe_1_2_1_n63) );
  AOI22_X1 npu_inst_pe_1_2_1_U31 ( .A1(npu_inst_n58), .A2(
        npu_inst_int_data_y_3__1__0_), .B1(npu_inst_pe_1_2_1_n3), .B2(
        npu_inst_int_data_x_2__2__0_), .ZN(npu_inst_pe_1_2_1_n61) );
  INV_X1 npu_inst_pe_1_2_1_U30 ( .A(npu_inst_pe_1_2_1_int_data_0_), .ZN(
        npu_inst_pe_1_2_1_n13) );
  INV_X1 npu_inst_pe_1_2_1_U29 ( .A(npu_inst_n70), .ZN(npu_inst_pe_1_2_1_n5)
         );
  OR3_X1 npu_inst_pe_1_2_1_U28 ( .A1(npu_inst_pe_1_2_1_n6), .A2(
        npu_inst_pe_1_2_1_n8), .A3(npu_inst_pe_1_2_1_n5), .ZN(
        npu_inst_pe_1_2_1_n56) );
  OR3_X1 npu_inst_pe_1_2_1_U27 ( .A1(npu_inst_pe_1_2_1_n5), .A2(
        npu_inst_pe_1_2_1_n8), .A3(npu_inst_pe_1_2_1_n7), .ZN(
        npu_inst_pe_1_2_1_n48) );
  INV_X1 npu_inst_pe_1_2_1_U26 ( .A(npu_inst_pe_1_2_1_n5), .ZN(
        npu_inst_pe_1_2_1_n4) );
  INV_X1 npu_inst_pe_1_2_1_U25 ( .A(npu_inst_n125), .ZN(npu_inst_pe_1_2_1_n12)
         );
  OR3_X1 npu_inst_pe_1_2_1_U24 ( .A1(npu_inst_pe_1_2_1_n4), .A2(
        npu_inst_pe_1_2_1_n8), .A3(npu_inst_pe_1_2_1_n7), .ZN(
        npu_inst_pe_1_2_1_n52) );
  OR3_X1 npu_inst_pe_1_2_1_U23 ( .A1(npu_inst_pe_1_2_1_n6), .A2(
        npu_inst_pe_1_2_1_n8), .A3(npu_inst_pe_1_2_1_n4), .ZN(
        npu_inst_pe_1_2_1_n60) );
  NOR2_X1 npu_inst_pe_1_2_1_U22 ( .A1(npu_inst_pe_1_2_1_n60), .A2(
        npu_inst_pe_1_2_1_n3), .ZN(npu_inst_pe_1_2_1_n58) );
  NOR2_X1 npu_inst_pe_1_2_1_U21 ( .A1(npu_inst_pe_1_2_1_n56), .A2(
        npu_inst_pe_1_2_1_n3), .ZN(npu_inst_pe_1_2_1_n54) );
  NOR2_X1 npu_inst_pe_1_2_1_U20 ( .A1(npu_inst_pe_1_2_1_n52), .A2(
        npu_inst_pe_1_2_1_n3), .ZN(npu_inst_pe_1_2_1_n50) );
  NOR2_X1 npu_inst_pe_1_2_1_U19 ( .A1(npu_inst_pe_1_2_1_n48), .A2(
        npu_inst_pe_1_2_1_n3), .ZN(npu_inst_pe_1_2_1_n46) );
  NOR2_X1 npu_inst_pe_1_2_1_U18 ( .A1(npu_inst_pe_1_2_1_n40), .A2(
        npu_inst_pe_1_2_1_n3), .ZN(npu_inst_pe_1_2_1_n38) );
  NOR2_X1 npu_inst_pe_1_2_1_U17 ( .A1(npu_inst_pe_1_2_1_n44), .A2(
        npu_inst_pe_1_2_1_n3), .ZN(npu_inst_pe_1_2_1_n42) );
  BUF_X1 npu_inst_pe_1_2_1_U16 ( .A(npu_inst_n103), .Z(npu_inst_pe_1_2_1_n8)
         );
  BUF_X1 npu_inst_pe_1_2_1_U15 ( .A(npu_inst_pe_1_2_1_n12), .Z(
        npu_inst_pe_1_2_1_n11) );
  BUF_X1 npu_inst_pe_1_2_1_U14 ( .A(npu_inst_pe_1_2_1_n12), .Z(
        npu_inst_pe_1_2_1_n10) );
  BUF_X1 npu_inst_pe_1_2_1_U13 ( .A(npu_inst_pe_1_2_1_n12), .Z(
        npu_inst_pe_1_2_1_n9) );
  INV_X1 npu_inst_pe_1_2_1_U12 ( .A(npu_inst_pe_1_2_1_n38), .ZN(
        npu_inst_pe_1_2_1_n118) );
  INV_X1 npu_inst_pe_1_2_1_U11 ( .A(npu_inst_pe_1_2_1_n58), .ZN(
        npu_inst_pe_1_2_1_n114) );
  INV_X1 npu_inst_pe_1_2_1_U10 ( .A(npu_inst_pe_1_2_1_n54), .ZN(
        npu_inst_pe_1_2_1_n115) );
  INV_X1 npu_inst_pe_1_2_1_U9 ( .A(npu_inst_pe_1_2_1_n50), .ZN(
        npu_inst_pe_1_2_1_n116) );
  INV_X1 npu_inst_pe_1_2_1_U8 ( .A(npu_inst_pe_1_2_1_n46), .ZN(
        npu_inst_pe_1_2_1_n117) );
  INV_X1 npu_inst_pe_1_2_1_U7 ( .A(npu_inst_pe_1_2_1_n42), .ZN(
        npu_inst_pe_1_2_1_n119) );
  BUF_X1 npu_inst_pe_1_2_1_U6 ( .A(npu_inst_n30), .Z(npu_inst_pe_1_2_1_n2) );
  BUF_X1 npu_inst_pe_1_2_1_U5 ( .A(npu_inst_n30), .Z(npu_inst_pe_1_2_1_n1) );
  NOR2_X1 npu_inst_pe_1_2_1_U4 ( .A1(npu_inst_pe_1_2_1_int_q_weight_0_), .A2(
        npu_inst_pe_1_2_1_n1), .ZN(npu_inst_pe_1_2_1_n76) );
  NOR2_X1 npu_inst_pe_1_2_1_U3 ( .A1(npu_inst_pe_1_2_1_n27), .A2(
        npu_inst_pe_1_2_1_n1), .ZN(npu_inst_pe_1_2_1_n77) );
  FA_X1 npu_inst_pe_1_2_1_sub_77_U2_1 ( .A(npu_inst_pe_1_2_1_int_q_acc_1_), 
        .B(npu_inst_pe_1_2_1_n14), .CI(npu_inst_pe_1_2_1_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_2_1_sub_77_carry_2_), .S(npu_inst_pe_1_2_1_N66) );
  FA_X1 npu_inst_pe_1_2_1_add_79_U1_1 ( .A(npu_inst_pe_1_2_1_int_q_acc_1_), 
        .B(npu_inst_pe_1_2_1_int_data_1_), .CI(
        npu_inst_pe_1_2_1_add_79_carry_1_), .CO(
        npu_inst_pe_1_2_1_add_79_carry_2_), .S(npu_inst_pe_1_2_1_N74) );
  NAND3_X1 npu_inst_pe_1_2_1_U109 ( .A1(npu_inst_pe_1_2_1_n5), .A2(
        npu_inst_pe_1_2_1_n7), .A3(npu_inst_pe_1_2_1_n8), .ZN(
        npu_inst_pe_1_2_1_n44) );
  NAND3_X1 npu_inst_pe_1_2_1_U108 ( .A1(npu_inst_pe_1_2_1_n4), .A2(
        npu_inst_pe_1_2_1_n7), .A3(npu_inst_pe_1_2_1_n8), .ZN(
        npu_inst_pe_1_2_1_n40) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_2_1_n34), .CK(
        npu_inst_pe_1_2_1_net3902), .RN(npu_inst_pe_1_2_1_n9), .Q(
        npu_inst_pe_1_2_1_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_2_1_n35), .CK(
        npu_inst_pe_1_2_1_net3902), .RN(npu_inst_pe_1_2_1_n9), .Q(
        npu_inst_pe_1_2_1_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_2_1_n36), .CK(
        npu_inst_pe_1_2_1_net3902), .RN(npu_inst_pe_1_2_1_n9), .Q(
        npu_inst_pe_1_2_1_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_2_1_n98), .CK(
        npu_inst_pe_1_2_1_net3902), .RN(npu_inst_pe_1_2_1_n9), .Q(
        npu_inst_pe_1_2_1_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_2_1_n99), .CK(
        npu_inst_pe_1_2_1_net3902), .RN(npu_inst_pe_1_2_1_n9), .Q(
        npu_inst_pe_1_2_1_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_2_1_n100), 
        .CK(npu_inst_pe_1_2_1_net3902), .RN(npu_inst_pe_1_2_1_n9), .Q(
        npu_inst_pe_1_2_1_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_2_1_n33), .CK(
        npu_inst_pe_1_2_1_net3902), .RN(npu_inst_pe_1_2_1_n9), .Q(
        npu_inst_pe_1_2_1_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_2_1_n101), 
        .CK(npu_inst_pe_1_2_1_net3902), .RN(npu_inst_pe_1_2_1_n9), .Q(
        npu_inst_pe_1_2_1_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_weight_reg_0_ ( .D(npu_inst_n111), .CK(
        npu_inst_pe_1_2_1_net3908), .RN(npu_inst_pe_1_2_1_n9), .Q(
        npu_inst_pe_1_2_1_int_q_weight_0_), .QN(npu_inst_pe_1_2_1_n27) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_weight_reg_1_ ( .D(npu_inst_n117), .CK(
        npu_inst_pe_1_2_1_net3908), .RN(npu_inst_pe_1_2_1_n9), .Q(
        npu_inst_pe_1_2_1_int_q_weight_1_), .QN(npu_inst_pe_1_2_1_n26) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_2_1_n113), 
        .CK(npu_inst_pe_1_2_1_net3908), .RN(npu_inst_pe_1_2_1_n9), .Q(
        npu_inst_pe_1_2_1_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_2_1_n107), 
        .CK(npu_inst_pe_1_2_1_net3908), .RN(npu_inst_pe_1_2_1_n9), .Q(
        npu_inst_pe_1_2_1_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_2_1_n112), 
        .CK(npu_inst_pe_1_2_1_net3908), .RN(npu_inst_pe_1_2_1_n10), .Q(
        npu_inst_pe_1_2_1_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_2_1_n106), 
        .CK(npu_inst_pe_1_2_1_net3908), .RN(npu_inst_pe_1_2_1_n10), .Q(
        npu_inst_pe_1_2_1_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_2_1_n111), 
        .CK(npu_inst_pe_1_2_1_net3908), .RN(npu_inst_pe_1_2_1_n10), .Q(
        npu_inst_pe_1_2_1_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_2_1_n105), 
        .CK(npu_inst_pe_1_2_1_net3908), .RN(npu_inst_pe_1_2_1_n10), .Q(
        npu_inst_pe_1_2_1_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_2_1_n110), 
        .CK(npu_inst_pe_1_2_1_net3908), .RN(npu_inst_pe_1_2_1_n10), .Q(
        npu_inst_pe_1_2_1_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_2_1_n104), 
        .CK(npu_inst_pe_1_2_1_net3908), .RN(npu_inst_pe_1_2_1_n10), .Q(
        npu_inst_pe_1_2_1_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_2_1_n109), 
        .CK(npu_inst_pe_1_2_1_net3908), .RN(npu_inst_pe_1_2_1_n10), .Q(
        npu_inst_pe_1_2_1_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_2_1_n103), 
        .CK(npu_inst_pe_1_2_1_net3908), .RN(npu_inst_pe_1_2_1_n10), .Q(
        npu_inst_pe_1_2_1_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_2_1_n108), 
        .CK(npu_inst_pe_1_2_1_net3908), .RN(npu_inst_pe_1_2_1_n10), .Q(
        npu_inst_pe_1_2_1_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_2_1_n102), 
        .CK(npu_inst_pe_1_2_1_net3908), .RN(npu_inst_pe_1_2_1_n10), .Q(
        npu_inst_pe_1_2_1_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_2_1_n86), 
        .CK(npu_inst_pe_1_2_1_net3908), .RN(npu_inst_pe_1_2_1_n10), .Q(
        npu_inst_pe_1_2_1_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_2_1_n87), 
        .CK(npu_inst_pe_1_2_1_net3908), .RN(npu_inst_pe_1_2_1_n10), .Q(
        npu_inst_pe_1_2_1_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_2_1_n88), 
        .CK(npu_inst_pe_1_2_1_net3908), .RN(npu_inst_pe_1_2_1_n11), .Q(
        npu_inst_pe_1_2_1_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_2_1_n89), 
        .CK(npu_inst_pe_1_2_1_net3908), .RN(npu_inst_pe_1_2_1_n11), .Q(
        npu_inst_pe_1_2_1_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_2_1_n90), 
        .CK(npu_inst_pe_1_2_1_net3908), .RN(npu_inst_pe_1_2_1_n11), .Q(
        npu_inst_pe_1_2_1_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_2_1_n91), 
        .CK(npu_inst_pe_1_2_1_net3908), .RN(npu_inst_pe_1_2_1_n11), .Q(
        npu_inst_pe_1_2_1_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_2_1_n92), 
        .CK(npu_inst_pe_1_2_1_net3908), .RN(npu_inst_pe_1_2_1_n11), .Q(
        npu_inst_pe_1_2_1_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_2_1_n93), 
        .CK(npu_inst_pe_1_2_1_net3908), .RN(npu_inst_pe_1_2_1_n11), .Q(
        npu_inst_pe_1_2_1_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_2_1_n94), 
        .CK(npu_inst_pe_1_2_1_net3908), .RN(npu_inst_pe_1_2_1_n11), .Q(
        npu_inst_pe_1_2_1_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_2_1_n95), 
        .CK(npu_inst_pe_1_2_1_net3908), .RN(npu_inst_pe_1_2_1_n11), .Q(
        npu_inst_pe_1_2_1_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_2_1_n96), 
        .CK(npu_inst_pe_1_2_1_net3908), .RN(npu_inst_pe_1_2_1_n11), .Q(
        npu_inst_pe_1_2_1_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_2_1_n97), 
        .CK(npu_inst_pe_1_2_1_net3908), .RN(npu_inst_pe_1_2_1_n11), .Q(
        npu_inst_pe_1_2_1_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_2_1_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_2_1_N84), .SE(1'b0), .GCK(npu_inst_pe_1_2_1_net3902) );
  CLKGATETST_X1 npu_inst_pe_1_2_1_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n65), .SE(1'b0), .GCK(npu_inst_pe_1_2_1_net3908) );
  MUX2_X1 npu_inst_pe_1_2_2_U162 ( .A(npu_inst_pe_1_2_2_n32), .B(
        npu_inst_pe_1_2_2_n29), .S(npu_inst_pe_1_2_2_n8), .Z(
        npu_inst_pe_1_2_2_N93) );
  MUX2_X1 npu_inst_pe_1_2_2_U161 ( .A(npu_inst_pe_1_2_2_n31), .B(
        npu_inst_pe_1_2_2_n30), .S(npu_inst_pe_1_2_2_n6), .Z(
        npu_inst_pe_1_2_2_n32) );
  MUX2_X1 npu_inst_pe_1_2_2_U160 ( .A(npu_inst_pe_1_2_2_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_2_2_int_q_reg_v_1__0_), .S(npu_inst_pe_1_2_2_n4), .Z(
        npu_inst_pe_1_2_2_n31) );
  MUX2_X1 npu_inst_pe_1_2_2_U159 ( .A(npu_inst_pe_1_2_2_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_2_2_int_q_reg_v_3__0_), .S(npu_inst_pe_1_2_2_n4), .Z(
        npu_inst_pe_1_2_2_n30) );
  MUX2_X1 npu_inst_pe_1_2_2_U158 ( .A(npu_inst_pe_1_2_2_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_2_2_int_q_reg_v_5__0_), .S(npu_inst_pe_1_2_2_n4), .Z(
        npu_inst_pe_1_2_2_n29) );
  MUX2_X1 npu_inst_pe_1_2_2_U157 ( .A(npu_inst_pe_1_2_2_n28), .B(
        npu_inst_pe_1_2_2_n23), .S(npu_inst_pe_1_2_2_n8), .Z(
        npu_inst_pe_1_2_2_N94) );
  MUX2_X1 npu_inst_pe_1_2_2_U156 ( .A(npu_inst_pe_1_2_2_n25), .B(
        npu_inst_pe_1_2_2_n24), .S(npu_inst_pe_1_2_2_n6), .Z(
        npu_inst_pe_1_2_2_n28) );
  MUX2_X1 npu_inst_pe_1_2_2_U155 ( .A(npu_inst_pe_1_2_2_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_2_2_int_q_reg_v_1__1_), .S(npu_inst_pe_1_2_2_n4), .Z(
        npu_inst_pe_1_2_2_n25) );
  MUX2_X1 npu_inst_pe_1_2_2_U154 ( .A(npu_inst_pe_1_2_2_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_2_2_int_q_reg_v_3__1_), .S(npu_inst_pe_1_2_2_n4), .Z(
        npu_inst_pe_1_2_2_n24) );
  MUX2_X1 npu_inst_pe_1_2_2_U153 ( .A(npu_inst_pe_1_2_2_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_2_2_int_q_reg_v_5__1_), .S(npu_inst_pe_1_2_2_n4), .Z(
        npu_inst_pe_1_2_2_n23) );
  MUX2_X1 npu_inst_pe_1_2_2_U152 ( .A(npu_inst_pe_1_2_2_n22), .B(
        npu_inst_pe_1_2_2_n19), .S(npu_inst_pe_1_2_2_n8), .Z(
        npu_inst_int_data_x_2__2__1_) );
  MUX2_X1 npu_inst_pe_1_2_2_U151 ( .A(npu_inst_pe_1_2_2_n21), .B(
        npu_inst_pe_1_2_2_n20), .S(npu_inst_pe_1_2_2_n6), .Z(
        npu_inst_pe_1_2_2_n22) );
  MUX2_X1 npu_inst_pe_1_2_2_U150 ( .A(npu_inst_pe_1_2_2_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_2_2_int_q_reg_h_1__1_), .S(npu_inst_pe_1_2_2_n4), .Z(
        npu_inst_pe_1_2_2_n21) );
  MUX2_X1 npu_inst_pe_1_2_2_U149 ( .A(npu_inst_pe_1_2_2_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_2_2_int_q_reg_h_3__1_), .S(npu_inst_pe_1_2_2_n4), .Z(
        npu_inst_pe_1_2_2_n20) );
  MUX2_X1 npu_inst_pe_1_2_2_U148 ( .A(npu_inst_pe_1_2_2_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_2_2_int_q_reg_h_5__1_), .S(npu_inst_pe_1_2_2_n4), .Z(
        npu_inst_pe_1_2_2_n19) );
  MUX2_X1 npu_inst_pe_1_2_2_U147 ( .A(npu_inst_pe_1_2_2_n18), .B(
        npu_inst_pe_1_2_2_n15), .S(npu_inst_pe_1_2_2_n8), .Z(
        npu_inst_int_data_x_2__2__0_) );
  MUX2_X1 npu_inst_pe_1_2_2_U146 ( .A(npu_inst_pe_1_2_2_n17), .B(
        npu_inst_pe_1_2_2_n16), .S(npu_inst_pe_1_2_2_n6), .Z(
        npu_inst_pe_1_2_2_n18) );
  MUX2_X1 npu_inst_pe_1_2_2_U145 ( .A(npu_inst_pe_1_2_2_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_2_2_int_q_reg_h_1__0_), .S(npu_inst_pe_1_2_2_n4), .Z(
        npu_inst_pe_1_2_2_n17) );
  MUX2_X1 npu_inst_pe_1_2_2_U144 ( .A(npu_inst_pe_1_2_2_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_2_2_int_q_reg_h_3__0_), .S(npu_inst_pe_1_2_2_n4), .Z(
        npu_inst_pe_1_2_2_n16) );
  MUX2_X1 npu_inst_pe_1_2_2_U143 ( .A(npu_inst_pe_1_2_2_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_2_2_int_q_reg_h_5__0_), .S(npu_inst_pe_1_2_2_n4), .Z(
        npu_inst_pe_1_2_2_n15) );
  XOR2_X1 npu_inst_pe_1_2_2_U142 ( .A(npu_inst_pe_1_2_2_int_data_0_), .B(
        npu_inst_pe_1_2_2_int_q_acc_0_), .Z(npu_inst_pe_1_2_2_N73) );
  AND2_X1 npu_inst_pe_1_2_2_U141 ( .A1(npu_inst_pe_1_2_2_int_q_acc_0_), .A2(
        npu_inst_pe_1_2_2_int_data_0_), .ZN(npu_inst_pe_1_2_2_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_2_2_U140 ( .A(npu_inst_pe_1_2_2_int_q_acc_0_), .B(
        npu_inst_pe_1_2_2_n13), .ZN(npu_inst_pe_1_2_2_N65) );
  OR2_X1 npu_inst_pe_1_2_2_U139 ( .A1(npu_inst_pe_1_2_2_n13), .A2(
        npu_inst_pe_1_2_2_int_q_acc_0_), .ZN(npu_inst_pe_1_2_2_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_2_2_U138 ( .A(npu_inst_pe_1_2_2_int_q_acc_2_), .B(
        npu_inst_pe_1_2_2_add_79_carry_2_), .Z(npu_inst_pe_1_2_2_N75) );
  AND2_X1 npu_inst_pe_1_2_2_U137 ( .A1(npu_inst_pe_1_2_2_add_79_carry_2_), 
        .A2(npu_inst_pe_1_2_2_int_q_acc_2_), .ZN(
        npu_inst_pe_1_2_2_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_2_2_U136 ( .A(npu_inst_pe_1_2_2_int_q_acc_3_), .B(
        npu_inst_pe_1_2_2_add_79_carry_3_), .Z(npu_inst_pe_1_2_2_N76) );
  AND2_X1 npu_inst_pe_1_2_2_U135 ( .A1(npu_inst_pe_1_2_2_add_79_carry_3_), 
        .A2(npu_inst_pe_1_2_2_int_q_acc_3_), .ZN(
        npu_inst_pe_1_2_2_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_2_2_U134 ( .A(npu_inst_pe_1_2_2_int_q_acc_4_), .B(
        npu_inst_pe_1_2_2_add_79_carry_4_), .Z(npu_inst_pe_1_2_2_N77) );
  AND2_X1 npu_inst_pe_1_2_2_U133 ( .A1(npu_inst_pe_1_2_2_add_79_carry_4_), 
        .A2(npu_inst_pe_1_2_2_int_q_acc_4_), .ZN(
        npu_inst_pe_1_2_2_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_2_2_U132 ( .A(npu_inst_pe_1_2_2_int_q_acc_5_), .B(
        npu_inst_pe_1_2_2_add_79_carry_5_), .Z(npu_inst_pe_1_2_2_N78) );
  AND2_X1 npu_inst_pe_1_2_2_U131 ( .A1(npu_inst_pe_1_2_2_add_79_carry_5_), 
        .A2(npu_inst_pe_1_2_2_int_q_acc_5_), .ZN(
        npu_inst_pe_1_2_2_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_2_2_U130 ( .A(npu_inst_pe_1_2_2_int_q_acc_6_), .B(
        npu_inst_pe_1_2_2_add_79_carry_6_), .Z(npu_inst_pe_1_2_2_N79) );
  AND2_X1 npu_inst_pe_1_2_2_U129 ( .A1(npu_inst_pe_1_2_2_add_79_carry_6_), 
        .A2(npu_inst_pe_1_2_2_int_q_acc_6_), .ZN(
        npu_inst_pe_1_2_2_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_2_2_U128 ( .A(npu_inst_pe_1_2_2_int_q_acc_7_), .B(
        npu_inst_pe_1_2_2_add_79_carry_7_), .Z(npu_inst_pe_1_2_2_N80) );
  XNOR2_X1 npu_inst_pe_1_2_2_U127 ( .A(npu_inst_pe_1_2_2_sub_77_carry_2_), .B(
        npu_inst_pe_1_2_2_int_q_acc_2_), .ZN(npu_inst_pe_1_2_2_N67) );
  OR2_X1 npu_inst_pe_1_2_2_U126 ( .A1(npu_inst_pe_1_2_2_int_q_acc_2_), .A2(
        npu_inst_pe_1_2_2_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_2_2_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_2_2_U125 ( .A(npu_inst_pe_1_2_2_sub_77_carry_3_), .B(
        npu_inst_pe_1_2_2_int_q_acc_3_), .ZN(npu_inst_pe_1_2_2_N68) );
  OR2_X1 npu_inst_pe_1_2_2_U124 ( .A1(npu_inst_pe_1_2_2_int_q_acc_3_), .A2(
        npu_inst_pe_1_2_2_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_2_2_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_2_2_U123 ( .A(npu_inst_pe_1_2_2_sub_77_carry_4_), .B(
        npu_inst_pe_1_2_2_int_q_acc_4_), .ZN(npu_inst_pe_1_2_2_N69) );
  OR2_X1 npu_inst_pe_1_2_2_U122 ( .A1(npu_inst_pe_1_2_2_int_q_acc_4_), .A2(
        npu_inst_pe_1_2_2_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_2_2_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_2_2_U121 ( .A(npu_inst_pe_1_2_2_sub_77_carry_5_), .B(
        npu_inst_pe_1_2_2_int_q_acc_5_), .ZN(npu_inst_pe_1_2_2_N70) );
  OR2_X1 npu_inst_pe_1_2_2_U120 ( .A1(npu_inst_pe_1_2_2_int_q_acc_5_), .A2(
        npu_inst_pe_1_2_2_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_2_2_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_2_2_U119 ( .A(npu_inst_pe_1_2_2_sub_77_carry_6_), .B(
        npu_inst_pe_1_2_2_int_q_acc_6_), .ZN(npu_inst_pe_1_2_2_N71) );
  OR2_X1 npu_inst_pe_1_2_2_U118 ( .A1(npu_inst_pe_1_2_2_int_q_acc_6_), .A2(
        npu_inst_pe_1_2_2_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_2_2_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_2_2_U117 ( .A(npu_inst_pe_1_2_2_int_q_acc_7_), .B(
        npu_inst_pe_1_2_2_sub_77_carry_7_), .ZN(npu_inst_pe_1_2_2_N72) );
  INV_X1 npu_inst_pe_1_2_2_U116 ( .A(npu_inst_n78), .ZN(npu_inst_pe_1_2_2_n7)
         );
  INV_X1 npu_inst_pe_1_2_2_U115 ( .A(npu_inst_pe_1_2_2_n7), .ZN(
        npu_inst_pe_1_2_2_n6) );
  INV_X1 npu_inst_pe_1_2_2_U114 ( .A(npu_inst_n58), .ZN(npu_inst_pe_1_2_2_n3)
         );
  AOI22_X1 npu_inst_pe_1_2_2_U113 ( .A1(npu_inst_int_data_y_3__2__0_), .A2(
        npu_inst_pe_1_2_2_n58), .B1(npu_inst_pe_1_2_2_n114), .B2(
        npu_inst_pe_1_2_2_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_2_2_n57) );
  INV_X1 npu_inst_pe_1_2_2_U112 ( .A(npu_inst_pe_1_2_2_n57), .ZN(
        npu_inst_pe_1_2_2_n108) );
  AOI22_X1 npu_inst_pe_1_2_2_U111 ( .A1(npu_inst_int_data_y_3__2__0_), .A2(
        npu_inst_pe_1_2_2_n54), .B1(npu_inst_pe_1_2_2_n115), .B2(
        npu_inst_pe_1_2_2_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_2_2_n53) );
  INV_X1 npu_inst_pe_1_2_2_U110 ( .A(npu_inst_pe_1_2_2_n53), .ZN(
        npu_inst_pe_1_2_2_n109) );
  AOI22_X1 npu_inst_pe_1_2_2_U107 ( .A1(npu_inst_int_data_y_3__2__0_), .A2(
        npu_inst_pe_1_2_2_n50), .B1(npu_inst_pe_1_2_2_n116), .B2(
        npu_inst_pe_1_2_2_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_2_2_n49) );
  INV_X1 npu_inst_pe_1_2_2_U106 ( .A(npu_inst_pe_1_2_2_n49), .ZN(
        npu_inst_pe_1_2_2_n110) );
  AOI22_X1 npu_inst_pe_1_2_2_U105 ( .A1(npu_inst_int_data_y_3__2__0_), .A2(
        npu_inst_pe_1_2_2_n46), .B1(npu_inst_pe_1_2_2_n117), .B2(
        npu_inst_pe_1_2_2_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_2_2_n45) );
  INV_X1 npu_inst_pe_1_2_2_U104 ( .A(npu_inst_pe_1_2_2_n45), .ZN(
        npu_inst_pe_1_2_2_n111) );
  AOI22_X1 npu_inst_pe_1_2_2_U103 ( .A1(npu_inst_int_data_y_3__2__0_), .A2(
        npu_inst_pe_1_2_2_n42), .B1(npu_inst_pe_1_2_2_n119), .B2(
        npu_inst_pe_1_2_2_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_2_2_n41) );
  INV_X1 npu_inst_pe_1_2_2_U102 ( .A(npu_inst_pe_1_2_2_n41), .ZN(
        npu_inst_pe_1_2_2_n112) );
  AOI22_X1 npu_inst_pe_1_2_2_U101 ( .A1(npu_inst_int_data_y_3__2__1_), .A2(
        npu_inst_pe_1_2_2_n58), .B1(npu_inst_pe_1_2_2_n114), .B2(
        npu_inst_pe_1_2_2_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_2_2_n59) );
  INV_X1 npu_inst_pe_1_2_2_U100 ( .A(npu_inst_pe_1_2_2_n59), .ZN(
        npu_inst_pe_1_2_2_n102) );
  AOI22_X1 npu_inst_pe_1_2_2_U99 ( .A1(npu_inst_int_data_y_3__2__1_), .A2(
        npu_inst_pe_1_2_2_n54), .B1(npu_inst_pe_1_2_2_n115), .B2(
        npu_inst_pe_1_2_2_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_2_2_n55) );
  INV_X1 npu_inst_pe_1_2_2_U98 ( .A(npu_inst_pe_1_2_2_n55), .ZN(
        npu_inst_pe_1_2_2_n103) );
  AOI22_X1 npu_inst_pe_1_2_2_U97 ( .A1(npu_inst_int_data_y_3__2__1_), .A2(
        npu_inst_pe_1_2_2_n50), .B1(npu_inst_pe_1_2_2_n116), .B2(
        npu_inst_pe_1_2_2_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_2_2_n51) );
  INV_X1 npu_inst_pe_1_2_2_U96 ( .A(npu_inst_pe_1_2_2_n51), .ZN(
        npu_inst_pe_1_2_2_n104) );
  AOI22_X1 npu_inst_pe_1_2_2_U95 ( .A1(npu_inst_int_data_y_3__2__1_), .A2(
        npu_inst_pe_1_2_2_n46), .B1(npu_inst_pe_1_2_2_n117), .B2(
        npu_inst_pe_1_2_2_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_2_2_n47) );
  INV_X1 npu_inst_pe_1_2_2_U94 ( .A(npu_inst_pe_1_2_2_n47), .ZN(
        npu_inst_pe_1_2_2_n105) );
  AOI22_X1 npu_inst_pe_1_2_2_U93 ( .A1(npu_inst_int_data_y_3__2__1_), .A2(
        npu_inst_pe_1_2_2_n42), .B1(npu_inst_pe_1_2_2_n119), .B2(
        npu_inst_pe_1_2_2_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_2_2_n43) );
  INV_X1 npu_inst_pe_1_2_2_U92 ( .A(npu_inst_pe_1_2_2_n43), .ZN(
        npu_inst_pe_1_2_2_n106) );
  AOI22_X1 npu_inst_pe_1_2_2_U91 ( .A1(npu_inst_pe_1_2_2_n38), .A2(
        npu_inst_int_data_y_3__2__1_), .B1(npu_inst_pe_1_2_2_n118), .B2(
        npu_inst_pe_1_2_2_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_2_2_n39) );
  INV_X1 npu_inst_pe_1_2_2_U90 ( .A(npu_inst_pe_1_2_2_n39), .ZN(
        npu_inst_pe_1_2_2_n107) );
  AOI22_X1 npu_inst_pe_1_2_2_U89 ( .A1(npu_inst_pe_1_2_2_n38), .A2(
        npu_inst_int_data_y_3__2__0_), .B1(npu_inst_pe_1_2_2_n118), .B2(
        npu_inst_pe_1_2_2_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_2_2_n37) );
  INV_X1 npu_inst_pe_1_2_2_U88 ( .A(npu_inst_pe_1_2_2_n37), .ZN(
        npu_inst_pe_1_2_2_n113) );
  NAND2_X1 npu_inst_pe_1_2_2_U87 ( .A1(npu_inst_pe_1_2_2_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_2_2_n60), .ZN(npu_inst_pe_1_2_2_n74) );
  OAI21_X1 npu_inst_pe_1_2_2_U86 ( .B1(npu_inst_pe_1_2_2_n63), .B2(
        npu_inst_pe_1_2_2_n60), .A(npu_inst_pe_1_2_2_n74), .ZN(
        npu_inst_pe_1_2_2_n97) );
  NAND2_X1 npu_inst_pe_1_2_2_U85 ( .A1(npu_inst_pe_1_2_2_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_2_2_n60), .ZN(npu_inst_pe_1_2_2_n73) );
  OAI21_X1 npu_inst_pe_1_2_2_U84 ( .B1(npu_inst_pe_1_2_2_n61), .B2(
        npu_inst_pe_1_2_2_n60), .A(npu_inst_pe_1_2_2_n73), .ZN(
        npu_inst_pe_1_2_2_n96) );
  NAND2_X1 npu_inst_pe_1_2_2_U83 ( .A1(npu_inst_pe_1_2_2_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_2_2_n56), .ZN(npu_inst_pe_1_2_2_n72) );
  OAI21_X1 npu_inst_pe_1_2_2_U82 ( .B1(npu_inst_pe_1_2_2_n63), .B2(
        npu_inst_pe_1_2_2_n56), .A(npu_inst_pe_1_2_2_n72), .ZN(
        npu_inst_pe_1_2_2_n95) );
  NAND2_X1 npu_inst_pe_1_2_2_U81 ( .A1(npu_inst_pe_1_2_2_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_2_2_n56), .ZN(npu_inst_pe_1_2_2_n71) );
  OAI21_X1 npu_inst_pe_1_2_2_U80 ( .B1(npu_inst_pe_1_2_2_n61), .B2(
        npu_inst_pe_1_2_2_n56), .A(npu_inst_pe_1_2_2_n71), .ZN(
        npu_inst_pe_1_2_2_n94) );
  NAND2_X1 npu_inst_pe_1_2_2_U79 ( .A1(npu_inst_pe_1_2_2_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_2_2_n52), .ZN(npu_inst_pe_1_2_2_n70) );
  OAI21_X1 npu_inst_pe_1_2_2_U78 ( .B1(npu_inst_pe_1_2_2_n63), .B2(
        npu_inst_pe_1_2_2_n52), .A(npu_inst_pe_1_2_2_n70), .ZN(
        npu_inst_pe_1_2_2_n93) );
  NAND2_X1 npu_inst_pe_1_2_2_U77 ( .A1(npu_inst_pe_1_2_2_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_2_2_n52), .ZN(npu_inst_pe_1_2_2_n69) );
  OAI21_X1 npu_inst_pe_1_2_2_U76 ( .B1(npu_inst_pe_1_2_2_n61), .B2(
        npu_inst_pe_1_2_2_n52), .A(npu_inst_pe_1_2_2_n69), .ZN(
        npu_inst_pe_1_2_2_n92) );
  NAND2_X1 npu_inst_pe_1_2_2_U75 ( .A1(npu_inst_pe_1_2_2_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_2_2_n48), .ZN(npu_inst_pe_1_2_2_n68) );
  OAI21_X1 npu_inst_pe_1_2_2_U74 ( .B1(npu_inst_pe_1_2_2_n63), .B2(
        npu_inst_pe_1_2_2_n48), .A(npu_inst_pe_1_2_2_n68), .ZN(
        npu_inst_pe_1_2_2_n91) );
  NAND2_X1 npu_inst_pe_1_2_2_U73 ( .A1(npu_inst_pe_1_2_2_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_2_2_n48), .ZN(npu_inst_pe_1_2_2_n67) );
  OAI21_X1 npu_inst_pe_1_2_2_U72 ( .B1(npu_inst_pe_1_2_2_n61), .B2(
        npu_inst_pe_1_2_2_n48), .A(npu_inst_pe_1_2_2_n67), .ZN(
        npu_inst_pe_1_2_2_n90) );
  NAND2_X1 npu_inst_pe_1_2_2_U71 ( .A1(npu_inst_pe_1_2_2_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_2_2_n44), .ZN(npu_inst_pe_1_2_2_n66) );
  OAI21_X1 npu_inst_pe_1_2_2_U70 ( .B1(npu_inst_pe_1_2_2_n63), .B2(
        npu_inst_pe_1_2_2_n44), .A(npu_inst_pe_1_2_2_n66), .ZN(
        npu_inst_pe_1_2_2_n89) );
  NAND2_X1 npu_inst_pe_1_2_2_U69 ( .A1(npu_inst_pe_1_2_2_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_2_2_n44), .ZN(npu_inst_pe_1_2_2_n65) );
  OAI21_X1 npu_inst_pe_1_2_2_U68 ( .B1(npu_inst_pe_1_2_2_n61), .B2(
        npu_inst_pe_1_2_2_n44), .A(npu_inst_pe_1_2_2_n65), .ZN(
        npu_inst_pe_1_2_2_n88) );
  NAND2_X1 npu_inst_pe_1_2_2_U67 ( .A1(npu_inst_pe_1_2_2_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_2_2_n40), .ZN(npu_inst_pe_1_2_2_n64) );
  OAI21_X1 npu_inst_pe_1_2_2_U66 ( .B1(npu_inst_pe_1_2_2_n63), .B2(
        npu_inst_pe_1_2_2_n40), .A(npu_inst_pe_1_2_2_n64), .ZN(
        npu_inst_pe_1_2_2_n87) );
  NAND2_X1 npu_inst_pe_1_2_2_U65 ( .A1(npu_inst_pe_1_2_2_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_2_2_n40), .ZN(npu_inst_pe_1_2_2_n62) );
  OAI21_X1 npu_inst_pe_1_2_2_U64 ( .B1(npu_inst_pe_1_2_2_n61), .B2(
        npu_inst_pe_1_2_2_n40), .A(npu_inst_pe_1_2_2_n62), .ZN(
        npu_inst_pe_1_2_2_n86) );
  AND2_X1 npu_inst_pe_1_2_2_U63 ( .A1(npu_inst_pe_1_2_2_N93), .A2(npu_inst_n58), .ZN(npu_inst_int_data_y_2__2__0_) );
  AND2_X1 npu_inst_pe_1_2_2_U62 ( .A1(npu_inst_n58), .A2(npu_inst_pe_1_2_2_N94), .ZN(npu_inst_int_data_y_2__2__1_) );
  NOR3_X1 npu_inst_pe_1_2_2_U61 ( .A1(npu_inst_pe_1_2_2_n26), .A2(npu_inst_n58), .A3(npu_inst_int_ckg[45]), .ZN(npu_inst_pe_1_2_2_n85) );
  OR2_X1 npu_inst_pe_1_2_2_U60 ( .A1(npu_inst_pe_1_2_2_n85), .A2(
        npu_inst_pe_1_2_2_n2), .ZN(npu_inst_pe_1_2_2_N84) );
  AND2_X1 npu_inst_pe_1_2_2_U59 ( .A1(npu_inst_pe_1_2_2_int_q_acc_0_), .A2(
        npu_inst_pe_1_2_2_n1), .ZN(npu_inst_int_data_res_2__2__0_) );
  AND2_X1 npu_inst_pe_1_2_2_U58 ( .A1(npu_inst_pe_1_2_2_n2), .A2(
        npu_inst_pe_1_2_2_int_q_acc_7_), .ZN(npu_inst_int_data_res_2__2__7_)
         );
  AND2_X1 npu_inst_pe_1_2_2_U57 ( .A1(npu_inst_pe_1_2_2_int_q_acc_1_), .A2(
        npu_inst_pe_1_2_2_n1), .ZN(npu_inst_int_data_res_2__2__1_) );
  AND2_X1 npu_inst_pe_1_2_2_U56 ( .A1(npu_inst_pe_1_2_2_int_q_acc_2_), .A2(
        npu_inst_pe_1_2_2_n1), .ZN(npu_inst_int_data_res_2__2__2_) );
  AND2_X1 npu_inst_pe_1_2_2_U55 ( .A1(npu_inst_pe_1_2_2_int_q_acc_3_), .A2(
        npu_inst_pe_1_2_2_n2), .ZN(npu_inst_int_data_res_2__2__3_) );
  AND2_X1 npu_inst_pe_1_2_2_U54 ( .A1(npu_inst_pe_1_2_2_int_q_acc_4_), .A2(
        npu_inst_pe_1_2_2_n2), .ZN(npu_inst_int_data_res_2__2__4_) );
  AND2_X1 npu_inst_pe_1_2_2_U53 ( .A1(npu_inst_pe_1_2_2_int_q_acc_5_), .A2(
        npu_inst_pe_1_2_2_n2), .ZN(npu_inst_int_data_res_2__2__5_) );
  AND2_X1 npu_inst_pe_1_2_2_U52 ( .A1(npu_inst_pe_1_2_2_int_q_acc_6_), .A2(
        npu_inst_pe_1_2_2_n2), .ZN(npu_inst_int_data_res_2__2__6_) );
  AOI222_X1 npu_inst_pe_1_2_2_U51 ( .A1(npu_inst_int_data_res_3__2__0_), .A2(
        npu_inst_pe_1_2_2_n1), .B1(npu_inst_pe_1_2_2_N73), .B2(
        npu_inst_pe_1_2_2_n76), .C1(npu_inst_pe_1_2_2_N65), .C2(
        npu_inst_pe_1_2_2_n77), .ZN(npu_inst_pe_1_2_2_n84) );
  INV_X1 npu_inst_pe_1_2_2_U50 ( .A(npu_inst_pe_1_2_2_n84), .ZN(
        npu_inst_pe_1_2_2_n101) );
  AOI222_X1 npu_inst_pe_1_2_2_U49 ( .A1(npu_inst_int_data_res_3__2__7_), .A2(
        npu_inst_pe_1_2_2_n1), .B1(npu_inst_pe_1_2_2_N80), .B2(
        npu_inst_pe_1_2_2_n76), .C1(npu_inst_pe_1_2_2_N72), .C2(
        npu_inst_pe_1_2_2_n77), .ZN(npu_inst_pe_1_2_2_n75) );
  INV_X1 npu_inst_pe_1_2_2_U48 ( .A(npu_inst_pe_1_2_2_n75), .ZN(
        npu_inst_pe_1_2_2_n33) );
  AOI222_X1 npu_inst_pe_1_2_2_U47 ( .A1(npu_inst_int_data_res_3__2__1_), .A2(
        npu_inst_pe_1_2_2_n1), .B1(npu_inst_pe_1_2_2_N74), .B2(
        npu_inst_pe_1_2_2_n76), .C1(npu_inst_pe_1_2_2_N66), .C2(
        npu_inst_pe_1_2_2_n77), .ZN(npu_inst_pe_1_2_2_n83) );
  INV_X1 npu_inst_pe_1_2_2_U46 ( .A(npu_inst_pe_1_2_2_n83), .ZN(
        npu_inst_pe_1_2_2_n100) );
  AOI222_X1 npu_inst_pe_1_2_2_U45 ( .A1(npu_inst_int_data_res_3__2__2_), .A2(
        npu_inst_pe_1_2_2_n1), .B1(npu_inst_pe_1_2_2_N75), .B2(
        npu_inst_pe_1_2_2_n76), .C1(npu_inst_pe_1_2_2_N67), .C2(
        npu_inst_pe_1_2_2_n77), .ZN(npu_inst_pe_1_2_2_n82) );
  INV_X1 npu_inst_pe_1_2_2_U44 ( .A(npu_inst_pe_1_2_2_n82), .ZN(
        npu_inst_pe_1_2_2_n99) );
  AOI222_X1 npu_inst_pe_1_2_2_U43 ( .A1(npu_inst_int_data_res_3__2__3_), .A2(
        npu_inst_pe_1_2_2_n1), .B1(npu_inst_pe_1_2_2_N76), .B2(
        npu_inst_pe_1_2_2_n76), .C1(npu_inst_pe_1_2_2_N68), .C2(
        npu_inst_pe_1_2_2_n77), .ZN(npu_inst_pe_1_2_2_n81) );
  INV_X1 npu_inst_pe_1_2_2_U42 ( .A(npu_inst_pe_1_2_2_n81), .ZN(
        npu_inst_pe_1_2_2_n98) );
  AOI222_X1 npu_inst_pe_1_2_2_U41 ( .A1(npu_inst_int_data_res_3__2__4_), .A2(
        npu_inst_pe_1_2_2_n1), .B1(npu_inst_pe_1_2_2_N77), .B2(
        npu_inst_pe_1_2_2_n76), .C1(npu_inst_pe_1_2_2_N69), .C2(
        npu_inst_pe_1_2_2_n77), .ZN(npu_inst_pe_1_2_2_n80) );
  INV_X1 npu_inst_pe_1_2_2_U40 ( .A(npu_inst_pe_1_2_2_n80), .ZN(
        npu_inst_pe_1_2_2_n36) );
  AOI222_X1 npu_inst_pe_1_2_2_U39 ( .A1(npu_inst_int_data_res_3__2__5_), .A2(
        npu_inst_pe_1_2_2_n1), .B1(npu_inst_pe_1_2_2_N78), .B2(
        npu_inst_pe_1_2_2_n76), .C1(npu_inst_pe_1_2_2_N70), .C2(
        npu_inst_pe_1_2_2_n77), .ZN(npu_inst_pe_1_2_2_n79) );
  INV_X1 npu_inst_pe_1_2_2_U38 ( .A(npu_inst_pe_1_2_2_n79), .ZN(
        npu_inst_pe_1_2_2_n35) );
  AOI222_X1 npu_inst_pe_1_2_2_U37 ( .A1(npu_inst_int_data_res_3__2__6_), .A2(
        npu_inst_pe_1_2_2_n1), .B1(npu_inst_pe_1_2_2_N79), .B2(
        npu_inst_pe_1_2_2_n76), .C1(npu_inst_pe_1_2_2_N71), .C2(
        npu_inst_pe_1_2_2_n77), .ZN(npu_inst_pe_1_2_2_n78) );
  INV_X1 npu_inst_pe_1_2_2_U36 ( .A(npu_inst_pe_1_2_2_n78), .ZN(
        npu_inst_pe_1_2_2_n34) );
  INV_X1 npu_inst_pe_1_2_2_U35 ( .A(npu_inst_pe_1_2_2_int_data_1_), .ZN(
        npu_inst_pe_1_2_2_n14) );
  AND2_X1 npu_inst_pe_1_2_2_U34 ( .A1(npu_inst_int_data_x_2__2__1_), .A2(
        npu_inst_pe_1_2_2_int_q_weight_1_), .ZN(npu_inst_pe_1_2_2_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_2_2_U33 ( .A1(npu_inst_int_data_x_2__2__0_), .A2(
        npu_inst_pe_1_2_2_int_q_weight_1_), .ZN(npu_inst_pe_1_2_2_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_2_2_U32 ( .A1(npu_inst_n58), .A2(
        npu_inst_int_data_y_3__2__1_), .B1(npu_inst_pe_1_2_2_n3), .B2(
        npu_inst_int_data_x_2__3__1_), .ZN(npu_inst_pe_1_2_2_n63) );
  AOI22_X1 npu_inst_pe_1_2_2_U31 ( .A1(npu_inst_n58), .A2(
        npu_inst_int_data_y_3__2__0_), .B1(npu_inst_pe_1_2_2_n3), .B2(
        npu_inst_int_data_x_2__3__0_), .ZN(npu_inst_pe_1_2_2_n61) );
  INV_X1 npu_inst_pe_1_2_2_U30 ( .A(npu_inst_pe_1_2_2_int_data_0_), .ZN(
        npu_inst_pe_1_2_2_n13) );
  INV_X1 npu_inst_pe_1_2_2_U29 ( .A(npu_inst_n70), .ZN(npu_inst_pe_1_2_2_n5)
         );
  OR3_X1 npu_inst_pe_1_2_2_U28 ( .A1(npu_inst_pe_1_2_2_n6), .A2(
        npu_inst_pe_1_2_2_n8), .A3(npu_inst_pe_1_2_2_n5), .ZN(
        npu_inst_pe_1_2_2_n56) );
  OR3_X1 npu_inst_pe_1_2_2_U27 ( .A1(npu_inst_pe_1_2_2_n5), .A2(
        npu_inst_pe_1_2_2_n8), .A3(npu_inst_pe_1_2_2_n7), .ZN(
        npu_inst_pe_1_2_2_n48) );
  INV_X1 npu_inst_pe_1_2_2_U26 ( .A(npu_inst_pe_1_2_2_n5), .ZN(
        npu_inst_pe_1_2_2_n4) );
  INV_X1 npu_inst_pe_1_2_2_U25 ( .A(npu_inst_n125), .ZN(npu_inst_pe_1_2_2_n12)
         );
  OR3_X1 npu_inst_pe_1_2_2_U24 ( .A1(npu_inst_pe_1_2_2_n4), .A2(
        npu_inst_pe_1_2_2_n8), .A3(npu_inst_pe_1_2_2_n7), .ZN(
        npu_inst_pe_1_2_2_n52) );
  OR3_X1 npu_inst_pe_1_2_2_U23 ( .A1(npu_inst_pe_1_2_2_n6), .A2(
        npu_inst_pe_1_2_2_n8), .A3(npu_inst_pe_1_2_2_n4), .ZN(
        npu_inst_pe_1_2_2_n60) );
  NOR2_X1 npu_inst_pe_1_2_2_U22 ( .A1(npu_inst_pe_1_2_2_n60), .A2(
        npu_inst_pe_1_2_2_n3), .ZN(npu_inst_pe_1_2_2_n58) );
  NOR2_X1 npu_inst_pe_1_2_2_U21 ( .A1(npu_inst_pe_1_2_2_n56), .A2(
        npu_inst_pe_1_2_2_n3), .ZN(npu_inst_pe_1_2_2_n54) );
  NOR2_X1 npu_inst_pe_1_2_2_U20 ( .A1(npu_inst_pe_1_2_2_n52), .A2(
        npu_inst_pe_1_2_2_n3), .ZN(npu_inst_pe_1_2_2_n50) );
  NOR2_X1 npu_inst_pe_1_2_2_U19 ( .A1(npu_inst_pe_1_2_2_n48), .A2(
        npu_inst_pe_1_2_2_n3), .ZN(npu_inst_pe_1_2_2_n46) );
  NOR2_X1 npu_inst_pe_1_2_2_U18 ( .A1(npu_inst_pe_1_2_2_n40), .A2(
        npu_inst_pe_1_2_2_n3), .ZN(npu_inst_pe_1_2_2_n38) );
  NOR2_X1 npu_inst_pe_1_2_2_U17 ( .A1(npu_inst_pe_1_2_2_n44), .A2(
        npu_inst_pe_1_2_2_n3), .ZN(npu_inst_pe_1_2_2_n42) );
  BUF_X1 npu_inst_pe_1_2_2_U16 ( .A(npu_inst_n103), .Z(npu_inst_pe_1_2_2_n8)
         );
  BUF_X1 npu_inst_pe_1_2_2_U15 ( .A(npu_inst_pe_1_2_2_n12), .Z(
        npu_inst_pe_1_2_2_n11) );
  BUF_X1 npu_inst_pe_1_2_2_U14 ( .A(npu_inst_pe_1_2_2_n12), .Z(
        npu_inst_pe_1_2_2_n10) );
  BUF_X1 npu_inst_pe_1_2_2_U13 ( .A(npu_inst_pe_1_2_2_n12), .Z(
        npu_inst_pe_1_2_2_n9) );
  INV_X1 npu_inst_pe_1_2_2_U12 ( .A(npu_inst_pe_1_2_2_n38), .ZN(
        npu_inst_pe_1_2_2_n118) );
  INV_X1 npu_inst_pe_1_2_2_U11 ( .A(npu_inst_pe_1_2_2_n58), .ZN(
        npu_inst_pe_1_2_2_n114) );
  INV_X1 npu_inst_pe_1_2_2_U10 ( .A(npu_inst_pe_1_2_2_n54), .ZN(
        npu_inst_pe_1_2_2_n115) );
  INV_X1 npu_inst_pe_1_2_2_U9 ( .A(npu_inst_pe_1_2_2_n50), .ZN(
        npu_inst_pe_1_2_2_n116) );
  INV_X1 npu_inst_pe_1_2_2_U8 ( .A(npu_inst_pe_1_2_2_n46), .ZN(
        npu_inst_pe_1_2_2_n117) );
  INV_X1 npu_inst_pe_1_2_2_U7 ( .A(npu_inst_pe_1_2_2_n42), .ZN(
        npu_inst_pe_1_2_2_n119) );
  BUF_X1 npu_inst_pe_1_2_2_U6 ( .A(npu_inst_n29), .Z(npu_inst_pe_1_2_2_n2) );
  BUF_X1 npu_inst_pe_1_2_2_U5 ( .A(npu_inst_n29), .Z(npu_inst_pe_1_2_2_n1) );
  NOR2_X1 npu_inst_pe_1_2_2_U4 ( .A1(npu_inst_pe_1_2_2_int_q_weight_0_), .A2(
        npu_inst_pe_1_2_2_n1), .ZN(npu_inst_pe_1_2_2_n76) );
  NOR2_X1 npu_inst_pe_1_2_2_U3 ( .A1(npu_inst_pe_1_2_2_n27), .A2(
        npu_inst_pe_1_2_2_n1), .ZN(npu_inst_pe_1_2_2_n77) );
  FA_X1 npu_inst_pe_1_2_2_sub_77_U2_1 ( .A(npu_inst_pe_1_2_2_int_q_acc_1_), 
        .B(npu_inst_pe_1_2_2_n14), .CI(npu_inst_pe_1_2_2_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_2_2_sub_77_carry_2_), .S(npu_inst_pe_1_2_2_N66) );
  FA_X1 npu_inst_pe_1_2_2_add_79_U1_1 ( .A(npu_inst_pe_1_2_2_int_q_acc_1_), 
        .B(npu_inst_pe_1_2_2_int_data_1_), .CI(
        npu_inst_pe_1_2_2_add_79_carry_1_), .CO(
        npu_inst_pe_1_2_2_add_79_carry_2_), .S(npu_inst_pe_1_2_2_N74) );
  NAND3_X1 npu_inst_pe_1_2_2_U109 ( .A1(npu_inst_pe_1_2_2_n5), .A2(
        npu_inst_pe_1_2_2_n7), .A3(npu_inst_pe_1_2_2_n8), .ZN(
        npu_inst_pe_1_2_2_n44) );
  NAND3_X1 npu_inst_pe_1_2_2_U108 ( .A1(npu_inst_pe_1_2_2_n4), .A2(
        npu_inst_pe_1_2_2_n7), .A3(npu_inst_pe_1_2_2_n8), .ZN(
        npu_inst_pe_1_2_2_n40) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_2_2_n34), .CK(
        npu_inst_pe_1_2_2_net3879), .RN(npu_inst_pe_1_2_2_n9), .Q(
        npu_inst_pe_1_2_2_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_2_2_n35), .CK(
        npu_inst_pe_1_2_2_net3879), .RN(npu_inst_pe_1_2_2_n9), .Q(
        npu_inst_pe_1_2_2_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_2_2_n36), .CK(
        npu_inst_pe_1_2_2_net3879), .RN(npu_inst_pe_1_2_2_n9), .Q(
        npu_inst_pe_1_2_2_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_2_2_n98), .CK(
        npu_inst_pe_1_2_2_net3879), .RN(npu_inst_pe_1_2_2_n9), .Q(
        npu_inst_pe_1_2_2_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_2_2_n99), .CK(
        npu_inst_pe_1_2_2_net3879), .RN(npu_inst_pe_1_2_2_n9), .Q(
        npu_inst_pe_1_2_2_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_2_2_n100), 
        .CK(npu_inst_pe_1_2_2_net3879), .RN(npu_inst_pe_1_2_2_n9), .Q(
        npu_inst_pe_1_2_2_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_2_2_n33), .CK(
        npu_inst_pe_1_2_2_net3879), .RN(npu_inst_pe_1_2_2_n9), .Q(
        npu_inst_pe_1_2_2_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_2_2_n101), 
        .CK(npu_inst_pe_1_2_2_net3879), .RN(npu_inst_pe_1_2_2_n9), .Q(
        npu_inst_pe_1_2_2_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_weight_reg_0_ ( .D(npu_inst_n111), .CK(
        npu_inst_pe_1_2_2_net3885), .RN(npu_inst_pe_1_2_2_n9), .Q(
        npu_inst_pe_1_2_2_int_q_weight_0_), .QN(npu_inst_pe_1_2_2_n27) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_weight_reg_1_ ( .D(npu_inst_n117), .CK(
        npu_inst_pe_1_2_2_net3885), .RN(npu_inst_pe_1_2_2_n9), .Q(
        npu_inst_pe_1_2_2_int_q_weight_1_), .QN(npu_inst_pe_1_2_2_n26) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_2_2_n113), 
        .CK(npu_inst_pe_1_2_2_net3885), .RN(npu_inst_pe_1_2_2_n9), .Q(
        npu_inst_pe_1_2_2_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_2_2_n107), 
        .CK(npu_inst_pe_1_2_2_net3885), .RN(npu_inst_pe_1_2_2_n9), .Q(
        npu_inst_pe_1_2_2_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_2_2_n112), 
        .CK(npu_inst_pe_1_2_2_net3885), .RN(npu_inst_pe_1_2_2_n10), .Q(
        npu_inst_pe_1_2_2_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_2_2_n106), 
        .CK(npu_inst_pe_1_2_2_net3885), .RN(npu_inst_pe_1_2_2_n10), .Q(
        npu_inst_pe_1_2_2_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_2_2_n111), 
        .CK(npu_inst_pe_1_2_2_net3885), .RN(npu_inst_pe_1_2_2_n10), .Q(
        npu_inst_pe_1_2_2_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_2_2_n105), 
        .CK(npu_inst_pe_1_2_2_net3885), .RN(npu_inst_pe_1_2_2_n10), .Q(
        npu_inst_pe_1_2_2_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_2_2_n110), 
        .CK(npu_inst_pe_1_2_2_net3885), .RN(npu_inst_pe_1_2_2_n10), .Q(
        npu_inst_pe_1_2_2_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_2_2_n104), 
        .CK(npu_inst_pe_1_2_2_net3885), .RN(npu_inst_pe_1_2_2_n10), .Q(
        npu_inst_pe_1_2_2_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_2_2_n109), 
        .CK(npu_inst_pe_1_2_2_net3885), .RN(npu_inst_pe_1_2_2_n10), .Q(
        npu_inst_pe_1_2_2_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_2_2_n103), 
        .CK(npu_inst_pe_1_2_2_net3885), .RN(npu_inst_pe_1_2_2_n10), .Q(
        npu_inst_pe_1_2_2_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_2_2_n108), 
        .CK(npu_inst_pe_1_2_2_net3885), .RN(npu_inst_pe_1_2_2_n10), .Q(
        npu_inst_pe_1_2_2_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_2_2_n102), 
        .CK(npu_inst_pe_1_2_2_net3885), .RN(npu_inst_pe_1_2_2_n10), .Q(
        npu_inst_pe_1_2_2_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_2_2_n86), 
        .CK(npu_inst_pe_1_2_2_net3885), .RN(npu_inst_pe_1_2_2_n10), .Q(
        npu_inst_pe_1_2_2_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_2_2_n87), 
        .CK(npu_inst_pe_1_2_2_net3885), .RN(npu_inst_pe_1_2_2_n10), .Q(
        npu_inst_pe_1_2_2_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_2_2_n88), 
        .CK(npu_inst_pe_1_2_2_net3885), .RN(npu_inst_pe_1_2_2_n11), .Q(
        npu_inst_pe_1_2_2_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_2_2_n89), 
        .CK(npu_inst_pe_1_2_2_net3885), .RN(npu_inst_pe_1_2_2_n11), .Q(
        npu_inst_pe_1_2_2_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_2_2_n90), 
        .CK(npu_inst_pe_1_2_2_net3885), .RN(npu_inst_pe_1_2_2_n11), .Q(
        npu_inst_pe_1_2_2_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_2_2_n91), 
        .CK(npu_inst_pe_1_2_2_net3885), .RN(npu_inst_pe_1_2_2_n11), .Q(
        npu_inst_pe_1_2_2_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_2_2_n92), 
        .CK(npu_inst_pe_1_2_2_net3885), .RN(npu_inst_pe_1_2_2_n11), .Q(
        npu_inst_pe_1_2_2_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_2_2_n93), 
        .CK(npu_inst_pe_1_2_2_net3885), .RN(npu_inst_pe_1_2_2_n11), .Q(
        npu_inst_pe_1_2_2_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_2_2_n94), 
        .CK(npu_inst_pe_1_2_2_net3885), .RN(npu_inst_pe_1_2_2_n11), .Q(
        npu_inst_pe_1_2_2_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_2_2_n95), 
        .CK(npu_inst_pe_1_2_2_net3885), .RN(npu_inst_pe_1_2_2_n11), .Q(
        npu_inst_pe_1_2_2_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_2_2_n96), 
        .CK(npu_inst_pe_1_2_2_net3885), .RN(npu_inst_pe_1_2_2_n11), .Q(
        npu_inst_pe_1_2_2_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_2_2_n97), 
        .CK(npu_inst_pe_1_2_2_net3885), .RN(npu_inst_pe_1_2_2_n11), .Q(
        npu_inst_pe_1_2_2_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_2_2_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_2_2_N84), .SE(1'b0), .GCK(npu_inst_pe_1_2_2_net3879) );
  CLKGATETST_X1 npu_inst_pe_1_2_2_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n65), .SE(1'b0), .GCK(npu_inst_pe_1_2_2_net3885) );
  MUX2_X1 npu_inst_pe_1_2_3_U162 ( .A(npu_inst_pe_1_2_3_n32), .B(
        npu_inst_pe_1_2_3_n29), .S(npu_inst_pe_1_2_3_n8), .Z(
        npu_inst_pe_1_2_3_N93) );
  MUX2_X1 npu_inst_pe_1_2_3_U161 ( .A(npu_inst_pe_1_2_3_n31), .B(
        npu_inst_pe_1_2_3_n30), .S(npu_inst_pe_1_2_3_n6), .Z(
        npu_inst_pe_1_2_3_n32) );
  MUX2_X1 npu_inst_pe_1_2_3_U160 ( .A(npu_inst_pe_1_2_3_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_2_3_int_q_reg_v_1__0_), .S(npu_inst_pe_1_2_3_n4), .Z(
        npu_inst_pe_1_2_3_n31) );
  MUX2_X1 npu_inst_pe_1_2_3_U159 ( .A(npu_inst_pe_1_2_3_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_2_3_int_q_reg_v_3__0_), .S(npu_inst_pe_1_2_3_n4), .Z(
        npu_inst_pe_1_2_3_n30) );
  MUX2_X1 npu_inst_pe_1_2_3_U158 ( .A(npu_inst_pe_1_2_3_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_2_3_int_q_reg_v_5__0_), .S(npu_inst_pe_1_2_3_n4), .Z(
        npu_inst_pe_1_2_3_n29) );
  MUX2_X1 npu_inst_pe_1_2_3_U157 ( .A(npu_inst_pe_1_2_3_n28), .B(
        npu_inst_pe_1_2_3_n23), .S(npu_inst_pe_1_2_3_n8), .Z(
        npu_inst_pe_1_2_3_N94) );
  MUX2_X1 npu_inst_pe_1_2_3_U156 ( .A(npu_inst_pe_1_2_3_n25), .B(
        npu_inst_pe_1_2_3_n24), .S(npu_inst_pe_1_2_3_n6), .Z(
        npu_inst_pe_1_2_3_n28) );
  MUX2_X1 npu_inst_pe_1_2_3_U155 ( .A(npu_inst_pe_1_2_3_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_2_3_int_q_reg_v_1__1_), .S(npu_inst_pe_1_2_3_n4), .Z(
        npu_inst_pe_1_2_3_n25) );
  MUX2_X1 npu_inst_pe_1_2_3_U154 ( .A(npu_inst_pe_1_2_3_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_2_3_int_q_reg_v_3__1_), .S(npu_inst_pe_1_2_3_n4), .Z(
        npu_inst_pe_1_2_3_n24) );
  MUX2_X1 npu_inst_pe_1_2_3_U153 ( .A(npu_inst_pe_1_2_3_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_2_3_int_q_reg_v_5__1_), .S(npu_inst_pe_1_2_3_n4), .Z(
        npu_inst_pe_1_2_3_n23) );
  MUX2_X1 npu_inst_pe_1_2_3_U152 ( .A(npu_inst_pe_1_2_3_n22), .B(
        npu_inst_pe_1_2_3_n19), .S(npu_inst_pe_1_2_3_n8), .Z(
        npu_inst_int_data_x_2__3__1_) );
  MUX2_X1 npu_inst_pe_1_2_3_U151 ( .A(npu_inst_pe_1_2_3_n21), .B(
        npu_inst_pe_1_2_3_n20), .S(npu_inst_pe_1_2_3_n6), .Z(
        npu_inst_pe_1_2_3_n22) );
  MUX2_X1 npu_inst_pe_1_2_3_U150 ( .A(npu_inst_pe_1_2_3_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_2_3_int_q_reg_h_1__1_), .S(npu_inst_pe_1_2_3_n4), .Z(
        npu_inst_pe_1_2_3_n21) );
  MUX2_X1 npu_inst_pe_1_2_3_U149 ( .A(npu_inst_pe_1_2_3_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_2_3_int_q_reg_h_3__1_), .S(npu_inst_pe_1_2_3_n4), .Z(
        npu_inst_pe_1_2_3_n20) );
  MUX2_X1 npu_inst_pe_1_2_3_U148 ( .A(npu_inst_pe_1_2_3_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_2_3_int_q_reg_h_5__1_), .S(npu_inst_pe_1_2_3_n4), .Z(
        npu_inst_pe_1_2_3_n19) );
  MUX2_X1 npu_inst_pe_1_2_3_U147 ( .A(npu_inst_pe_1_2_3_n18), .B(
        npu_inst_pe_1_2_3_n15), .S(npu_inst_pe_1_2_3_n8), .Z(
        npu_inst_int_data_x_2__3__0_) );
  MUX2_X1 npu_inst_pe_1_2_3_U146 ( .A(npu_inst_pe_1_2_3_n17), .B(
        npu_inst_pe_1_2_3_n16), .S(npu_inst_pe_1_2_3_n6), .Z(
        npu_inst_pe_1_2_3_n18) );
  MUX2_X1 npu_inst_pe_1_2_3_U145 ( .A(npu_inst_pe_1_2_3_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_2_3_int_q_reg_h_1__0_), .S(npu_inst_pe_1_2_3_n4), .Z(
        npu_inst_pe_1_2_3_n17) );
  MUX2_X1 npu_inst_pe_1_2_3_U144 ( .A(npu_inst_pe_1_2_3_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_2_3_int_q_reg_h_3__0_), .S(npu_inst_pe_1_2_3_n4), .Z(
        npu_inst_pe_1_2_3_n16) );
  MUX2_X1 npu_inst_pe_1_2_3_U143 ( .A(npu_inst_pe_1_2_3_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_2_3_int_q_reg_h_5__0_), .S(npu_inst_pe_1_2_3_n4), .Z(
        npu_inst_pe_1_2_3_n15) );
  XOR2_X1 npu_inst_pe_1_2_3_U142 ( .A(npu_inst_pe_1_2_3_int_data_0_), .B(
        npu_inst_pe_1_2_3_int_q_acc_0_), .Z(npu_inst_pe_1_2_3_N73) );
  AND2_X1 npu_inst_pe_1_2_3_U141 ( .A1(npu_inst_pe_1_2_3_int_q_acc_0_), .A2(
        npu_inst_pe_1_2_3_int_data_0_), .ZN(npu_inst_pe_1_2_3_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_2_3_U140 ( .A(npu_inst_pe_1_2_3_int_q_acc_0_), .B(
        npu_inst_pe_1_2_3_n13), .ZN(npu_inst_pe_1_2_3_N65) );
  OR2_X1 npu_inst_pe_1_2_3_U139 ( .A1(npu_inst_pe_1_2_3_n13), .A2(
        npu_inst_pe_1_2_3_int_q_acc_0_), .ZN(npu_inst_pe_1_2_3_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_2_3_U138 ( .A(npu_inst_pe_1_2_3_int_q_acc_2_), .B(
        npu_inst_pe_1_2_3_add_79_carry_2_), .Z(npu_inst_pe_1_2_3_N75) );
  AND2_X1 npu_inst_pe_1_2_3_U137 ( .A1(npu_inst_pe_1_2_3_add_79_carry_2_), 
        .A2(npu_inst_pe_1_2_3_int_q_acc_2_), .ZN(
        npu_inst_pe_1_2_3_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_2_3_U136 ( .A(npu_inst_pe_1_2_3_int_q_acc_3_), .B(
        npu_inst_pe_1_2_3_add_79_carry_3_), .Z(npu_inst_pe_1_2_3_N76) );
  AND2_X1 npu_inst_pe_1_2_3_U135 ( .A1(npu_inst_pe_1_2_3_add_79_carry_3_), 
        .A2(npu_inst_pe_1_2_3_int_q_acc_3_), .ZN(
        npu_inst_pe_1_2_3_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_2_3_U134 ( .A(npu_inst_pe_1_2_3_int_q_acc_4_), .B(
        npu_inst_pe_1_2_3_add_79_carry_4_), .Z(npu_inst_pe_1_2_3_N77) );
  AND2_X1 npu_inst_pe_1_2_3_U133 ( .A1(npu_inst_pe_1_2_3_add_79_carry_4_), 
        .A2(npu_inst_pe_1_2_3_int_q_acc_4_), .ZN(
        npu_inst_pe_1_2_3_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_2_3_U132 ( .A(npu_inst_pe_1_2_3_int_q_acc_5_), .B(
        npu_inst_pe_1_2_3_add_79_carry_5_), .Z(npu_inst_pe_1_2_3_N78) );
  AND2_X1 npu_inst_pe_1_2_3_U131 ( .A1(npu_inst_pe_1_2_3_add_79_carry_5_), 
        .A2(npu_inst_pe_1_2_3_int_q_acc_5_), .ZN(
        npu_inst_pe_1_2_3_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_2_3_U130 ( .A(npu_inst_pe_1_2_3_int_q_acc_6_), .B(
        npu_inst_pe_1_2_3_add_79_carry_6_), .Z(npu_inst_pe_1_2_3_N79) );
  AND2_X1 npu_inst_pe_1_2_3_U129 ( .A1(npu_inst_pe_1_2_3_add_79_carry_6_), 
        .A2(npu_inst_pe_1_2_3_int_q_acc_6_), .ZN(
        npu_inst_pe_1_2_3_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_2_3_U128 ( .A(npu_inst_pe_1_2_3_int_q_acc_7_), .B(
        npu_inst_pe_1_2_3_add_79_carry_7_), .Z(npu_inst_pe_1_2_3_N80) );
  XNOR2_X1 npu_inst_pe_1_2_3_U127 ( .A(npu_inst_pe_1_2_3_sub_77_carry_2_), .B(
        npu_inst_pe_1_2_3_int_q_acc_2_), .ZN(npu_inst_pe_1_2_3_N67) );
  OR2_X1 npu_inst_pe_1_2_3_U126 ( .A1(npu_inst_pe_1_2_3_int_q_acc_2_), .A2(
        npu_inst_pe_1_2_3_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_2_3_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_2_3_U125 ( .A(npu_inst_pe_1_2_3_sub_77_carry_3_), .B(
        npu_inst_pe_1_2_3_int_q_acc_3_), .ZN(npu_inst_pe_1_2_3_N68) );
  OR2_X1 npu_inst_pe_1_2_3_U124 ( .A1(npu_inst_pe_1_2_3_int_q_acc_3_), .A2(
        npu_inst_pe_1_2_3_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_2_3_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_2_3_U123 ( .A(npu_inst_pe_1_2_3_sub_77_carry_4_), .B(
        npu_inst_pe_1_2_3_int_q_acc_4_), .ZN(npu_inst_pe_1_2_3_N69) );
  OR2_X1 npu_inst_pe_1_2_3_U122 ( .A1(npu_inst_pe_1_2_3_int_q_acc_4_), .A2(
        npu_inst_pe_1_2_3_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_2_3_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_2_3_U121 ( .A(npu_inst_pe_1_2_3_sub_77_carry_5_), .B(
        npu_inst_pe_1_2_3_int_q_acc_5_), .ZN(npu_inst_pe_1_2_3_N70) );
  OR2_X1 npu_inst_pe_1_2_3_U120 ( .A1(npu_inst_pe_1_2_3_int_q_acc_5_), .A2(
        npu_inst_pe_1_2_3_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_2_3_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_2_3_U119 ( .A(npu_inst_pe_1_2_3_sub_77_carry_6_), .B(
        npu_inst_pe_1_2_3_int_q_acc_6_), .ZN(npu_inst_pe_1_2_3_N71) );
  OR2_X1 npu_inst_pe_1_2_3_U118 ( .A1(npu_inst_pe_1_2_3_int_q_acc_6_), .A2(
        npu_inst_pe_1_2_3_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_2_3_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_2_3_U117 ( .A(npu_inst_pe_1_2_3_int_q_acc_7_), .B(
        npu_inst_pe_1_2_3_sub_77_carry_7_), .ZN(npu_inst_pe_1_2_3_N72) );
  INV_X1 npu_inst_pe_1_2_3_U116 ( .A(npu_inst_n78), .ZN(npu_inst_pe_1_2_3_n7)
         );
  INV_X1 npu_inst_pe_1_2_3_U115 ( .A(npu_inst_pe_1_2_3_n7), .ZN(
        npu_inst_pe_1_2_3_n6) );
  INV_X1 npu_inst_pe_1_2_3_U114 ( .A(npu_inst_n58), .ZN(npu_inst_pe_1_2_3_n3)
         );
  AOI22_X1 npu_inst_pe_1_2_3_U113 ( .A1(npu_inst_int_data_y_3__3__0_), .A2(
        npu_inst_pe_1_2_3_n58), .B1(npu_inst_pe_1_2_3_n114), .B2(
        npu_inst_pe_1_2_3_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_2_3_n57) );
  INV_X1 npu_inst_pe_1_2_3_U112 ( .A(npu_inst_pe_1_2_3_n57), .ZN(
        npu_inst_pe_1_2_3_n108) );
  AOI22_X1 npu_inst_pe_1_2_3_U111 ( .A1(npu_inst_int_data_y_3__3__0_), .A2(
        npu_inst_pe_1_2_3_n54), .B1(npu_inst_pe_1_2_3_n115), .B2(
        npu_inst_pe_1_2_3_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_2_3_n53) );
  INV_X1 npu_inst_pe_1_2_3_U110 ( .A(npu_inst_pe_1_2_3_n53), .ZN(
        npu_inst_pe_1_2_3_n109) );
  AOI22_X1 npu_inst_pe_1_2_3_U107 ( .A1(npu_inst_int_data_y_3__3__0_), .A2(
        npu_inst_pe_1_2_3_n50), .B1(npu_inst_pe_1_2_3_n116), .B2(
        npu_inst_pe_1_2_3_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_2_3_n49) );
  INV_X1 npu_inst_pe_1_2_3_U106 ( .A(npu_inst_pe_1_2_3_n49), .ZN(
        npu_inst_pe_1_2_3_n110) );
  AOI22_X1 npu_inst_pe_1_2_3_U105 ( .A1(npu_inst_int_data_y_3__3__0_), .A2(
        npu_inst_pe_1_2_3_n46), .B1(npu_inst_pe_1_2_3_n117), .B2(
        npu_inst_pe_1_2_3_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_2_3_n45) );
  INV_X1 npu_inst_pe_1_2_3_U104 ( .A(npu_inst_pe_1_2_3_n45), .ZN(
        npu_inst_pe_1_2_3_n111) );
  AOI22_X1 npu_inst_pe_1_2_3_U103 ( .A1(npu_inst_int_data_y_3__3__0_), .A2(
        npu_inst_pe_1_2_3_n42), .B1(npu_inst_pe_1_2_3_n119), .B2(
        npu_inst_pe_1_2_3_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_2_3_n41) );
  INV_X1 npu_inst_pe_1_2_3_U102 ( .A(npu_inst_pe_1_2_3_n41), .ZN(
        npu_inst_pe_1_2_3_n112) );
  AOI22_X1 npu_inst_pe_1_2_3_U101 ( .A1(npu_inst_int_data_y_3__3__1_), .A2(
        npu_inst_pe_1_2_3_n58), .B1(npu_inst_pe_1_2_3_n114), .B2(
        npu_inst_pe_1_2_3_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_2_3_n59) );
  INV_X1 npu_inst_pe_1_2_3_U100 ( .A(npu_inst_pe_1_2_3_n59), .ZN(
        npu_inst_pe_1_2_3_n102) );
  AOI22_X1 npu_inst_pe_1_2_3_U99 ( .A1(npu_inst_int_data_y_3__3__1_), .A2(
        npu_inst_pe_1_2_3_n54), .B1(npu_inst_pe_1_2_3_n115), .B2(
        npu_inst_pe_1_2_3_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_2_3_n55) );
  INV_X1 npu_inst_pe_1_2_3_U98 ( .A(npu_inst_pe_1_2_3_n55), .ZN(
        npu_inst_pe_1_2_3_n103) );
  AOI22_X1 npu_inst_pe_1_2_3_U97 ( .A1(npu_inst_int_data_y_3__3__1_), .A2(
        npu_inst_pe_1_2_3_n50), .B1(npu_inst_pe_1_2_3_n116), .B2(
        npu_inst_pe_1_2_3_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_2_3_n51) );
  INV_X1 npu_inst_pe_1_2_3_U96 ( .A(npu_inst_pe_1_2_3_n51), .ZN(
        npu_inst_pe_1_2_3_n104) );
  AOI22_X1 npu_inst_pe_1_2_3_U95 ( .A1(npu_inst_int_data_y_3__3__1_), .A2(
        npu_inst_pe_1_2_3_n46), .B1(npu_inst_pe_1_2_3_n117), .B2(
        npu_inst_pe_1_2_3_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_2_3_n47) );
  INV_X1 npu_inst_pe_1_2_3_U94 ( .A(npu_inst_pe_1_2_3_n47), .ZN(
        npu_inst_pe_1_2_3_n105) );
  AOI22_X1 npu_inst_pe_1_2_3_U93 ( .A1(npu_inst_int_data_y_3__3__1_), .A2(
        npu_inst_pe_1_2_3_n42), .B1(npu_inst_pe_1_2_3_n119), .B2(
        npu_inst_pe_1_2_3_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_2_3_n43) );
  INV_X1 npu_inst_pe_1_2_3_U92 ( .A(npu_inst_pe_1_2_3_n43), .ZN(
        npu_inst_pe_1_2_3_n106) );
  AOI22_X1 npu_inst_pe_1_2_3_U91 ( .A1(npu_inst_pe_1_2_3_n38), .A2(
        npu_inst_int_data_y_3__3__1_), .B1(npu_inst_pe_1_2_3_n118), .B2(
        npu_inst_pe_1_2_3_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_2_3_n39) );
  INV_X1 npu_inst_pe_1_2_3_U90 ( .A(npu_inst_pe_1_2_3_n39), .ZN(
        npu_inst_pe_1_2_3_n107) );
  AOI22_X1 npu_inst_pe_1_2_3_U89 ( .A1(npu_inst_pe_1_2_3_n38), .A2(
        npu_inst_int_data_y_3__3__0_), .B1(npu_inst_pe_1_2_3_n118), .B2(
        npu_inst_pe_1_2_3_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_2_3_n37) );
  INV_X1 npu_inst_pe_1_2_3_U88 ( .A(npu_inst_pe_1_2_3_n37), .ZN(
        npu_inst_pe_1_2_3_n113) );
  NAND2_X1 npu_inst_pe_1_2_3_U87 ( .A1(npu_inst_pe_1_2_3_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_2_3_n60), .ZN(npu_inst_pe_1_2_3_n74) );
  OAI21_X1 npu_inst_pe_1_2_3_U86 ( .B1(npu_inst_pe_1_2_3_n63), .B2(
        npu_inst_pe_1_2_3_n60), .A(npu_inst_pe_1_2_3_n74), .ZN(
        npu_inst_pe_1_2_3_n97) );
  NAND2_X1 npu_inst_pe_1_2_3_U85 ( .A1(npu_inst_pe_1_2_3_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_2_3_n60), .ZN(npu_inst_pe_1_2_3_n73) );
  OAI21_X1 npu_inst_pe_1_2_3_U84 ( .B1(npu_inst_pe_1_2_3_n61), .B2(
        npu_inst_pe_1_2_3_n60), .A(npu_inst_pe_1_2_3_n73), .ZN(
        npu_inst_pe_1_2_3_n96) );
  NAND2_X1 npu_inst_pe_1_2_3_U83 ( .A1(npu_inst_pe_1_2_3_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_2_3_n56), .ZN(npu_inst_pe_1_2_3_n72) );
  OAI21_X1 npu_inst_pe_1_2_3_U82 ( .B1(npu_inst_pe_1_2_3_n63), .B2(
        npu_inst_pe_1_2_3_n56), .A(npu_inst_pe_1_2_3_n72), .ZN(
        npu_inst_pe_1_2_3_n95) );
  NAND2_X1 npu_inst_pe_1_2_3_U81 ( .A1(npu_inst_pe_1_2_3_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_2_3_n56), .ZN(npu_inst_pe_1_2_3_n71) );
  OAI21_X1 npu_inst_pe_1_2_3_U80 ( .B1(npu_inst_pe_1_2_3_n61), .B2(
        npu_inst_pe_1_2_3_n56), .A(npu_inst_pe_1_2_3_n71), .ZN(
        npu_inst_pe_1_2_3_n94) );
  NAND2_X1 npu_inst_pe_1_2_3_U79 ( .A1(npu_inst_pe_1_2_3_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_2_3_n52), .ZN(npu_inst_pe_1_2_3_n70) );
  OAI21_X1 npu_inst_pe_1_2_3_U78 ( .B1(npu_inst_pe_1_2_3_n63), .B2(
        npu_inst_pe_1_2_3_n52), .A(npu_inst_pe_1_2_3_n70), .ZN(
        npu_inst_pe_1_2_3_n93) );
  NAND2_X1 npu_inst_pe_1_2_3_U77 ( .A1(npu_inst_pe_1_2_3_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_2_3_n52), .ZN(npu_inst_pe_1_2_3_n69) );
  OAI21_X1 npu_inst_pe_1_2_3_U76 ( .B1(npu_inst_pe_1_2_3_n61), .B2(
        npu_inst_pe_1_2_3_n52), .A(npu_inst_pe_1_2_3_n69), .ZN(
        npu_inst_pe_1_2_3_n92) );
  NAND2_X1 npu_inst_pe_1_2_3_U75 ( .A1(npu_inst_pe_1_2_3_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_2_3_n48), .ZN(npu_inst_pe_1_2_3_n68) );
  OAI21_X1 npu_inst_pe_1_2_3_U74 ( .B1(npu_inst_pe_1_2_3_n63), .B2(
        npu_inst_pe_1_2_3_n48), .A(npu_inst_pe_1_2_3_n68), .ZN(
        npu_inst_pe_1_2_3_n91) );
  NAND2_X1 npu_inst_pe_1_2_3_U73 ( .A1(npu_inst_pe_1_2_3_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_2_3_n48), .ZN(npu_inst_pe_1_2_3_n67) );
  OAI21_X1 npu_inst_pe_1_2_3_U72 ( .B1(npu_inst_pe_1_2_3_n61), .B2(
        npu_inst_pe_1_2_3_n48), .A(npu_inst_pe_1_2_3_n67), .ZN(
        npu_inst_pe_1_2_3_n90) );
  NAND2_X1 npu_inst_pe_1_2_3_U71 ( .A1(npu_inst_pe_1_2_3_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_2_3_n44), .ZN(npu_inst_pe_1_2_3_n66) );
  OAI21_X1 npu_inst_pe_1_2_3_U70 ( .B1(npu_inst_pe_1_2_3_n63), .B2(
        npu_inst_pe_1_2_3_n44), .A(npu_inst_pe_1_2_3_n66), .ZN(
        npu_inst_pe_1_2_3_n89) );
  NAND2_X1 npu_inst_pe_1_2_3_U69 ( .A1(npu_inst_pe_1_2_3_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_2_3_n44), .ZN(npu_inst_pe_1_2_3_n65) );
  OAI21_X1 npu_inst_pe_1_2_3_U68 ( .B1(npu_inst_pe_1_2_3_n61), .B2(
        npu_inst_pe_1_2_3_n44), .A(npu_inst_pe_1_2_3_n65), .ZN(
        npu_inst_pe_1_2_3_n88) );
  NAND2_X1 npu_inst_pe_1_2_3_U67 ( .A1(npu_inst_pe_1_2_3_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_2_3_n40), .ZN(npu_inst_pe_1_2_3_n64) );
  OAI21_X1 npu_inst_pe_1_2_3_U66 ( .B1(npu_inst_pe_1_2_3_n63), .B2(
        npu_inst_pe_1_2_3_n40), .A(npu_inst_pe_1_2_3_n64), .ZN(
        npu_inst_pe_1_2_3_n87) );
  NAND2_X1 npu_inst_pe_1_2_3_U65 ( .A1(npu_inst_pe_1_2_3_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_2_3_n40), .ZN(npu_inst_pe_1_2_3_n62) );
  OAI21_X1 npu_inst_pe_1_2_3_U64 ( .B1(npu_inst_pe_1_2_3_n61), .B2(
        npu_inst_pe_1_2_3_n40), .A(npu_inst_pe_1_2_3_n62), .ZN(
        npu_inst_pe_1_2_3_n86) );
  AND2_X1 npu_inst_pe_1_2_3_U63 ( .A1(npu_inst_pe_1_2_3_N93), .A2(npu_inst_n58), .ZN(npu_inst_int_data_y_2__3__0_) );
  AND2_X1 npu_inst_pe_1_2_3_U62 ( .A1(npu_inst_n58), .A2(npu_inst_pe_1_2_3_N94), .ZN(npu_inst_int_data_y_2__3__1_) );
  NOR3_X1 npu_inst_pe_1_2_3_U61 ( .A1(npu_inst_pe_1_2_3_n26), .A2(npu_inst_n58), .A3(npu_inst_int_ckg[44]), .ZN(npu_inst_pe_1_2_3_n85) );
  OR2_X1 npu_inst_pe_1_2_3_U60 ( .A1(npu_inst_pe_1_2_3_n85), .A2(
        npu_inst_pe_1_2_3_n2), .ZN(npu_inst_pe_1_2_3_N84) );
  AND2_X1 npu_inst_pe_1_2_3_U59 ( .A1(npu_inst_pe_1_2_3_int_q_acc_0_), .A2(
        npu_inst_pe_1_2_3_n1), .ZN(npu_inst_int_data_res_2__3__0_) );
  AND2_X1 npu_inst_pe_1_2_3_U58 ( .A1(npu_inst_pe_1_2_3_n2), .A2(
        npu_inst_pe_1_2_3_int_q_acc_7_), .ZN(npu_inst_int_data_res_2__3__7_)
         );
  AND2_X1 npu_inst_pe_1_2_3_U57 ( .A1(npu_inst_pe_1_2_3_int_q_acc_1_), .A2(
        npu_inst_pe_1_2_3_n1), .ZN(npu_inst_int_data_res_2__3__1_) );
  AND2_X1 npu_inst_pe_1_2_3_U56 ( .A1(npu_inst_pe_1_2_3_int_q_acc_2_), .A2(
        npu_inst_pe_1_2_3_n1), .ZN(npu_inst_int_data_res_2__3__2_) );
  AND2_X1 npu_inst_pe_1_2_3_U55 ( .A1(npu_inst_pe_1_2_3_int_q_acc_3_), .A2(
        npu_inst_pe_1_2_3_n2), .ZN(npu_inst_int_data_res_2__3__3_) );
  AND2_X1 npu_inst_pe_1_2_3_U54 ( .A1(npu_inst_pe_1_2_3_int_q_acc_4_), .A2(
        npu_inst_pe_1_2_3_n2), .ZN(npu_inst_int_data_res_2__3__4_) );
  AND2_X1 npu_inst_pe_1_2_3_U53 ( .A1(npu_inst_pe_1_2_3_int_q_acc_5_), .A2(
        npu_inst_pe_1_2_3_n2), .ZN(npu_inst_int_data_res_2__3__5_) );
  AND2_X1 npu_inst_pe_1_2_3_U52 ( .A1(npu_inst_pe_1_2_3_int_q_acc_6_), .A2(
        npu_inst_pe_1_2_3_n2), .ZN(npu_inst_int_data_res_2__3__6_) );
  AOI222_X1 npu_inst_pe_1_2_3_U51 ( .A1(npu_inst_int_data_res_3__3__0_), .A2(
        npu_inst_pe_1_2_3_n1), .B1(npu_inst_pe_1_2_3_N73), .B2(
        npu_inst_pe_1_2_3_n76), .C1(npu_inst_pe_1_2_3_N65), .C2(
        npu_inst_pe_1_2_3_n77), .ZN(npu_inst_pe_1_2_3_n84) );
  INV_X1 npu_inst_pe_1_2_3_U50 ( .A(npu_inst_pe_1_2_3_n84), .ZN(
        npu_inst_pe_1_2_3_n101) );
  AOI222_X1 npu_inst_pe_1_2_3_U49 ( .A1(npu_inst_int_data_res_3__3__7_), .A2(
        npu_inst_pe_1_2_3_n1), .B1(npu_inst_pe_1_2_3_N80), .B2(
        npu_inst_pe_1_2_3_n76), .C1(npu_inst_pe_1_2_3_N72), .C2(
        npu_inst_pe_1_2_3_n77), .ZN(npu_inst_pe_1_2_3_n75) );
  INV_X1 npu_inst_pe_1_2_3_U48 ( .A(npu_inst_pe_1_2_3_n75), .ZN(
        npu_inst_pe_1_2_3_n33) );
  AOI222_X1 npu_inst_pe_1_2_3_U47 ( .A1(npu_inst_int_data_res_3__3__1_), .A2(
        npu_inst_pe_1_2_3_n1), .B1(npu_inst_pe_1_2_3_N74), .B2(
        npu_inst_pe_1_2_3_n76), .C1(npu_inst_pe_1_2_3_N66), .C2(
        npu_inst_pe_1_2_3_n77), .ZN(npu_inst_pe_1_2_3_n83) );
  INV_X1 npu_inst_pe_1_2_3_U46 ( .A(npu_inst_pe_1_2_3_n83), .ZN(
        npu_inst_pe_1_2_3_n100) );
  AOI222_X1 npu_inst_pe_1_2_3_U45 ( .A1(npu_inst_int_data_res_3__3__2_), .A2(
        npu_inst_pe_1_2_3_n1), .B1(npu_inst_pe_1_2_3_N75), .B2(
        npu_inst_pe_1_2_3_n76), .C1(npu_inst_pe_1_2_3_N67), .C2(
        npu_inst_pe_1_2_3_n77), .ZN(npu_inst_pe_1_2_3_n82) );
  INV_X1 npu_inst_pe_1_2_3_U44 ( .A(npu_inst_pe_1_2_3_n82), .ZN(
        npu_inst_pe_1_2_3_n99) );
  AOI222_X1 npu_inst_pe_1_2_3_U43 ( .A1(npu_inst_int_data_res_3__3__3_), .A2(
        npu_inst_pe_1_2_3_n1), .B1(npu_inst_pe_1_2_3_N76), .B2(
        npu_inst_pe_1_2_3_n76), .C1(npu_inst_pe_1_2_3_N68), .C2(
        npu_inst_pe_1_2_3_n77), .ZN(npu_inst_pe_1_2_3_n81) );
  INV_X1 npu_inst_pe_1_2_3_U42 ( .A(npu_inst_pe_1_2_3_n81), .ZN(
        npu_inst_pe_1_2_3_n98) );
  AOI222_X1 npu_inst_pe_1_2_3_U41 ( .A1(npu_inst_int_data_res_3__3__4_), .A2(
        npu_inst_pe_1_2_3_n1), .B1(npu_inst_pe_1_2_3_N77), .B2(
        npu_inst_pe_1_2_3_n76), .C1(npu_inst_pe_1_2_3_N69), .C2(
        npu_inst_pe_1_2_3_n77), .ZN(npu_inst_pe_1_2_3_n80) );
  INV_X1 npu_inst_pe_1_2_3_U40 ( .A(npu_inst_pe_1_2_3_n80), .ZN(
        npu_inst_pe_1_2_3_n36) );
  AOI222_X1 npu_inst_pe_1_2_3_U39 ( .A1(npu_inst_int_data_res_3__3__5_), .A2(
        npu_inst_pe_1_2_3_n1), .B1(npu_inst_pe_1_2_3_N78), .B2(
        npu_inst_pe_1_2_3_n76), .C1(npu_inst_pe_1_2_3_N70), .C2(
        npu_inst_pe_1_2_3_n77), .ZN(npu_inst_pe_1_2_3_n79) );
  INV_X1 npu_inst_pe_1_2_3_U38 ( .A(npu_inst_pe_1_2_3_n79), .ZN(
        npu_inst_pe_1_2_3_n35) );
  AOI222_X1 npu_inst_pe_1_2_3_U37 ( .A1(npu_inst_int_data_res_3__3__6_), .A2(
        npu_inst_pe_1_2_3_n1), .B1(npu_inst_pe_1_2_3_N79), .B2(
        npu_inst_pe_1_2_3_n76), .C1(npu_inst_pe_1_2_3_N71), .C2(
        npu_inst_pe_1_2_3_n77), .ZN(npu_inst_pe_1_2_3_n78) );
  INV_X1 npu_inst_pe_1_2_3_U36 ( .A(npu_inst_pe_1_2_3_n78), .ZN(
        npu_inst_pe_1_2_3_n34) );
  INV_X1 npu_inst_pe_1_2_3_U35 ( .A(npu_inst_pe_1_2_3_int_data_1_), .ZN(
        npu_inst_pe_1_2_3_n14) );
  AND2_X1 npu_inst_pe_1_2_3_U34 ( .A1(npu_inst_int_data_x_2__3__1_), .A2(
        npu_inst_pe_1_2_3_int_q_weight_1_), .ZN(npu_inst_pe_1_2_3_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_2_3_U33 ( .A1(npu_inst_int_data_x_2__3__0_), .A2(
        npu_inst_pe_1_2_3_int_q_weight_1_), .ZN(npu_inst_pe_1_2_3_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_2_3_U32 ( .A1(npu_inst_n58), .A2(
        npu_inst_int_data_y_3__3__1_), .B1(npu_inst_pe_1_2_3_n3), .B2(
        npu_inst_int_data_x_2__4__1_), .ZN(npu_inst_pe_1_2_3_n63) );
  AOI22_X1 npu_inst_pe_1_2_3_U31 ( .A1(npu_inst_n58), .A2(
        npu_inst_int_data_y_3__3__0_), .B1(npu_inst_pe_1_2_3_n3), .B2(
        npu_inst_int_data_x_2__4__0_), .ZN(npu_inst_pe_1_2_3_n61) );
  INV_X1 npu_inst_pe_1_2_3_U30 ( .A(npu_inst_pe_1_2_3_int_data_0_), .ZN(
        npu_inst_pe_1_2_3_n13) );
  INV_X1 npu_inst_pe_1_2_3_U29 ( .A(npu_inst_n70), .ZN(npu_inst_pe_1_2_3_n5)
         );
  OR3_X1 npu_inst_pe_1_2_3_U28 ( .A1(npu_inst_pe_1_2_3_n6), .A2(
        npu_inst_pe_1_2_3_n8), .A3(npu_inst_pe_1_2_3_n5), .ZN(
        npu_inst_pe_1_2_3_n56) );
  OR3_X1 npu_inst_pe_1_2_3_U27 ( .A1(npu_inst_pe_1_2_3_n5), .A2(
        npu_inst_pe_1_2_3_n8), .A3(npu_inst_pe_1_2_3_n7), .ZN(
        npu_inst_pe_1_2_3_n48) );
  INV_X1 npu_inst_pe_1_2_3_U26 ( .A(npu_inst_pe_1_2_3_n5), .ZN(
        npu_inst_pe_1_2_3_n4) );
  INV_X1 npu_inst_pe_1_2_3_U25 ( .A(npu_inst_n125), .ZN(npu_inst_pe_1_2_3_n12)
         );
  OR3_X1 npu_inst_pe_1_2_3_U24 ( .A1(npu_inst_pe_1_2_3_n4), .A2(
        npu_inst_pe_1_2_3_n8), .A3(npu_inst_pe_1_2_3_n7), .ZN(
        npu_inst_pe_1_2_3_n52) );
  OR3_X1 npu_inst_pe_1_2_3_U23 ( .A1(npu_inst_pe_1_2_3_n6), .A2(
        npu_inst_pe_1_2_3_n8), .A3(npu_inst_pe_1_2_3_n4), .ZN(
        npu_inst_pe_1_2_3_n60) );
  NOR2_X1 npu_inst_pe_1_2_3_U22 ( .A1(npu_inst_pe_1_2_3_n60), .A2(
        npu_inst_pe_1_2_3_n3), .ZN(npu_inst_pe_1_2_3_n58) );
  NOR2_X1 npu_inst_pe_1_2_3_U21 ( .A1(npu_inst_pe_1_2_3_n56), .A2(
        npu_inst_pe_1_2_3_n3), .ZN(npu_inst_pe_1_2_3_n54) );
  NOR2_X1 npu_inst_pe_1_2_3_U20 ( .A1(npu_inst_pe_1_2_3_n52), .A2(
        npu_inst_pe_1_2_3_n3), .ZN(npu_inst_pe_1_2_3_n50) );
  NOR2_X1 npu_inst_pe_1_2_3_U19 ( .A1(npu_inst_pe_1_2_3_n48), .A2(
        npu_inst_pe_1_2_3_n3), .ZN(npu_inst_pe_1_2_3_n46) );
  NOR2_X1 npu_inst_pe_1_2_3_U18 ( .A1(npu_inst_pe_1_2_3_n40), .A2(
        npu_inst_pe_1_2_3_n3), .ZN(npu_inst_pe_1_2_3_n38) );
  NOR2_X1 npu_inst_pe_1_2_3_U17 ( .A1(npu_inst_pe_1_2_3_n44), .A2(
        npu_inst_pe_1_2_3_n3), .ZN(npu_inst_pe_1_2_3_n42) );
  BUF_X1 npu_inst_pe_1_2_3_U16 ( .A(npu_inst_n103), .Z(npu_inst_pe_1_2_3_n8)
         );
  BUF_X1 npu_inst_pe_1_2_3_U15 ( .A(npu_inst_pe_1_2_3_n12), .Z(
        npu_inst_pe_1_2_3_n11) );
  BUF_X1 npu_inst_pe_1_2_3_U14 ( .A(npu_inst_pe_1_2_3_n12), .Z(
        npu_inst_pe_1_2_3_n10) );
  BUF_X1 npu_inst_pe_1_2_3_U13 ( .A(npu_inst_pe_1_2_3_n12), .Z(
        npu_inst_pe_1_2_3_n9) );
  INV_X1 npu_inst_pe_1_2_3_U12 ( .A(npu_inst_pe_1_2_3_n38), .ZN(
        npu_inst_pe_1_2_3_n118) );
  INV_X1 npu_inst_pe_1_2_3_U11 ( .A(npu_inst_pe_1_2_3_n58), .ZN(
        npu_inst_pe_1_2_3_n114) );
  INV_X1 npu_inst_pe_1_2_3_U10 ( .A(npu_inst_pe_1_2_3_n54), .ZN(
        npu_inst_pe_1_2_3_n115) );
  INV_X1 npu_inst_pe_1_2_3_U9 ( .A(npu_inst_pe_1_2_3_n50), .ZN(
        npu_inst_pe_1_2_3_n116) );
  INV_X1 npu_inst_pe_1_2_3_U8 ( .A(npu_inst_pe_1_2_3_n46), .ZN(
        npu_inst_pe_1_2_3_n117) );
  INV_X1 npu_inst_pe_1_2_3_U7 ( .A(npu_inst_pe_1_2_3_n42), .ZN(
        npu_inst_pe_1_2_3_n119) );
  BUF_X1 npu_inst_pe_1_2_3_U6 ( .A(npu_inst_n29), .Z(npu_inst_pe_1_2_3_n2) );
  BUF_X1 npu_inst_pe_1_2_3_U5 ( .A(npu_inst_n29), .Z(npu_inst_pe_1_2_3_n1) );
  NOR2_X1 npu_inst_pe_1_2_3_U4 ( .A1(npu_inst_pe_1_2_3_int_q_weight_0_), .A2(
        npu_inst_pe_1_2_3_n1), .ZN(npu_inst_pe_1_2_3_n76) );
  NOR2_X1 npu_inst_pe_1_2_3_U3 ( .A1(npu_inst_pe_1_2_3_n27), .A2(
        npu_inst_pe_1_2_3_n1), .ZN(npu_inst_pe_1_2_3_n77) );
  FA_X1 npu_inst_pe_1_2_3_sub_77_U2_1 ( .A(npu_inst_pe_1_2_3_int_q_acc_1_), 
        .B(npu_inst_pe_1_2_3_n14), .CI(npu_inst_pe_1_2_3_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_2_3_sub_77_carry_2_), .S(npu_inst_pe_1_2_3_N66) );
  FA_X1 npu_inst_pe_1_2_3_add_79_U1_1 ( .A(npu_inst_pe_1_2_3_int_q_acc_1_), 
        .B(npu_inst_pe_1_2_3_int_data_1_), .CI(
        npu_inst_pe_1_2_3_add_79_carry_1_), .CO(
        npu_inst_pe_1_2_3_add_79_carry_2_), .S(npu_inst_pe_1_2_3_N74) );
  NAND3_X1 npu_inst_pe_1_2_3_U109 ( .A1(npu_inst_pe_1_2_3_n5), .A2(
        npu_inst_pe_1_2_3_n7), .A3(npu_inst_pe_1_2_3_n8), .ZN(
        npu_inst_pe_1_2_3_n44) );
  NAND3_X1 npu_inst_pe_1_2_3_U108 ( .A1(npu_inst_pe_1_2_3_n4), .A2(
        npu_inst_pe_1_2_3_n7), .A3(npu_inst_pe_1_2_3_n8), .ZN(
        npu_inst_pe_1_2_3_n40) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_2_3_n34), .CK(
        npu_inst_pe_1_2_3_net3856), .RN(npu_inst_pe_1_2_3_n9), .Q(
        npu_inst_pe_1_2_3_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_2_3_n35), .CK(
        npu_inst_pe_1_2_3_net3856), .RN(npu_inst_pe_1_2_3_n9), .Q(
        npu_inst_pe_1_2_3_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_2_3_n36), .CK(
        npu_inst_pe_1_2_3_net3856), .RN(npu_inst_pe_1_2_3_n9), .Q(
        npu_inst_pe_1_2_3_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_2_3_n98), .CK(
        npu_inst_pe_1_2_3_net3856), .RN(npu_inst_pe_1_2_3_n9), .Q(
        npu_inst_pe_1_2_3_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_2_3_n99), .CK(
        npu_inst_pe_1_2_3_net3856), .RN(npu_inst_pe_1_2_3_n9), .Q(
        npu_inst_pe_1_2_3_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_2_3_n100), 
        .CK(npu_inst_pe_1_2_3_net3856), .RN(npu_inst_pe_1_2_3_n9), .Q(
        npu_inst_pe_1_2_3_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_2_3_n33), .CK(
        npu_inst_pe_1_2_3_net3856), .RN(npu_inst_pe_1_2_3_n9), .Q(
        npu_inst_pe_1_2_3_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_2_3_n101), 
        .CK(npu_inst_pe_1_2_3_net3856), .RN(npu_inst_pe_1_2_3_n9), .Q(
        npu_inst_pe_1_2_3_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_weight_reg_0_ ( .D(npu_inst_n111), .CK(
        npu_inst_pe_1_2_3_net3862), .RN(npu_inst_pe_1_2_3_n9), .Q(
        npu_inst_pe_1_2_3_int_q_weight_0_), .QN(npu_inst_pe_1_2_3_n27) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_weight_reg_1_ ( .D(npu_inst_n117), .CK(
        npu_inst_pe_1_2_3_net3862), .RN(npu_inst_pe_1_2_3_n9), .Q(
        npu_inst_pe_1_2_3_int_q_weight_1_), .QN(npu_inst_pe_1_2_3_n26) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_2_3_n113), 
        .CK(npu_inst_pe_1_2_3_net3862), .RN(npu_inst_pe_1_2_3_n9), .Q(
        npu_inst_pe_1_2_3_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_2_3_n107), 
        .CK(npu_inst_pe_1_2_3_net3862), .RN(npu_inst_pe_1_2_3_n9), .Q(
        npu_inst_pe_1_2_3_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_2_3_n112), 
        .CK(npu_inst_pe_1_2_3_net3862), .RN(npu_inst_pe_1_2_3_n10), .Q(
        npu_inst_pe_1_2_3_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_2_3_n106), 
        .CK(npu_inst_pe_1_2_3_net3862), .RN(npu_inst_pe_1_2_3_n10), .Q(
        npu_inst_pe_1_2_3_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_2_3_n111), 
        .CK(npu_inst_pe_1_2_3_net3862), .RN(npu_inst_pe_1_2_3_n10), .Q(
        npu_inst_pe_1_2_3_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_2_3_n105), 
        .CK(npu_inst_pe_1_2_3_net3862), .RN(npu_inst_pe_1_2_3_n10), .Q(
        npu_inst_pe_1_2_3_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_2_3_n110), 
        .CK(npu_inst_pe_1_2_3_net3862), .RN(npu_inst_pe_1_2_3_n10), .Q(
        npu_inst_pe_1_2_3_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_2_3_n104), 
        .CK(npu_inst_pe_1_2_3_net3862), .RN(npu_inst_pe_1_2_3_n10), .Q(
        npu_inst_pe_1_2_3_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_2_3_n109), 
        .CK(npu_inst_pe_1_2_3_net3862), .RN(npu_inst_pe_1_2_3_n10), .Q(
        npu_inst_pe_1_2_3_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_2_3_n103), 
        .CK(npu_inst_pe_1_2_3_net3862), .RN(npu_inst_pe_1_2_3_n10), .Q(
        npu_inst_pe_1_2_3_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_2_3_n108), 
        .CK(npu_inst_pe_1_2_3_net3862), .RN(npu_inst_pe_1_2_3_n10), .Q(
        npu_inst_pe_1_2_3_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_2_3_n102), 
        .CK(npu_inst_pe_1_2_3_net3862), .RN(npu_inst_pe_1_2_3_n10), .Q(
        npu_inst_pe_1_2_3_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_2_3_n86), 
        .CK(npu_inst_pe_1_2_3_net3862), .RN(npu_inst_pe_1_2_3_n10), .Q(
        npu_inst_pe_1_2_3_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_2_3_n87), 
        .CK(npu_inst_pe_1_2_3_net3862), .RN(npu_inst_pe_1_2_3_n10), .Q(
        npu_inst_pe_1_2_3_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_2_3_n88), 
        .CK(npu_inst_pe_1_2_3_net3862), .RN(npu_inst_pe_1_2_3_n11), .Q(
        npu_inst_pe_1_2_3_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_2_3_n89), 
        .CK(npu_inst_pe_1_2_3_net3862), .RN(npu_inst_pe_1_2_3_n11), .Q(
        npu_inst_pe_1_2_3_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_2_3_n90), 
        .CK(npu_inst_pe_1_2_3_net3862), .RN(npu_inst_pe_1_2_3_n11), .Q(
        npu_inst_pe_1_2_3_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_2_3_n91), 
        .CK(npu_inst_pe_1_2_3_net3862), .RN(npu_inst_pe_1_2_3_n11), .Q(
        npu_inst_pe_1_2_3_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_2_3_n92), 
        .CK(npu_inst_pe_1_2_3_net3862), .RN(npu_inst_pe_1_2_3_n11), .Q(
        npu_inst_pe_1_2_3_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_2_3_n93), 
        .CK(npu_inst_pe_1_2_3_net3862), .RN(npu_inst_pe_1_2_3_n11), .Q(
        npu_inst_pe_1_2_3_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_2_3_n94), 
        .CK(npu_inst_pe_1_2_3_net3862), .RN(npu_inst_pe_1_2_3_n11), .Q(
        npu_inst_pe_1_2_3_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_2_3_n95), 
        .CK(npu_inst_pe_1_2_3_net3862), .RN(npu_inst_pe_1_2_3_n11), .Q(
        npu_inst_pe_1_2_3_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_2_3_n96), 
        .CK(npu_inst_pe_1_2_3_net3862), .RN(npu_inst_pe_1_2_3_n11), .Q(
        npu_inst_pe_1_2_3_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_2_3_n97), 
        .CK(npu_inst_pe_1_2_3_net3862), .RN(npu_inst_pe_1_2_3_n11), .Q(
        npu_inst_pe_1_2_3_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_2_3_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_2_3_N84), .SE(1'b0), .GCK(npu_inst_pe_1_2_3_net3856) );
  CLKGATETST_X1 npu_inst_pe_1_2_3_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n65), .SE(1'b0), .GCK(npu_inst_pe_1_2_3_net3862) );
  MUX2_X1 npu_inst_pe_1_2_4_U162 ( .A(npu_inst_pe_1_2_4_n32), .B(
        npu_inst_pe_1_2_4_n29), .S(npu_inst_pe_1_2_4_n8), .Z(
        npu_inst_pe_1_2_4_N93) );
  MUX2_X1 npu_inst_pe_1_2_4_U161 ( .A(npu_inst_pe_1_2_4_n31), .B(
        npu_inst_pe_1_2_4_n30), .S(npu_inst_pe_1_2_4_n6), .Z(
        npu_inst_pe_1_2_4_n32) );
  MUX2_X1 npu_inst_pe_1_2_4_U160 ( .A(npu_inst_pe_1_2_4_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_2_4_int_q_reg_v_1__0_), .S(npu_inst_pe_1_2_4_n4), .Z(
        npu_inst_pe_1_2_4_n31) );
  MUX2_X1 npu_inst_pe_1_2_4_U159 ( .A(npu_inst_pe_1_2_4_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_2_4_int_q_reg_v_3__0_), .S(npu_inst_pe_1_2_4_n4), .Z(
        npu_inst_pe_1_2_4_n30) );
  MUX2_X1 npu_inst_pe_1_2_4_U158 ( .A(npu_inst_pe_1_2_4_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_2_4_int_q_reg_v_5__0_), .S(npu_inst_pe_1_2_4_n4), .Z(
        npu_inst_pe_1_2_4_n29) );
  MUX2_X1 npu_inst_pe_1_2_4_U157 ( .A(npu_inst_pe_1_2_4_n28), .B(
        npu_inst_pe_1_2_4_n23), .S(npu_inst_pe_1_2_4_n8), .Z(
        npu_inst_pe_1_2_4_N94) );
  MUX2_X1 npu_inst_pe_1_2_4_U156 ( .A(npu_inst_pe_1_2_4_n25), .B(
        npu_inst_pe_1_2_4_n24), .S(npu_inst_pe_1_2_4_n6), .Z(
        npu_inst_pe_1_2_4_n28) );
  MUX2_X1 npu_inst_pe_1_2_4_U155 ( .A(npu_inst_pe_1_2_4_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_2_4_int_q_reg_v_1__1_), .S(npu_inst_pe_1_2_4_n4), .Z(
        npu_inst_pe_1_2_4_n25) );
  MUX2_X1 npu_inst_pe_1_2_4_U154 ( .A(npu_inst_pe_1_2_4_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_2_4_int_q_reg_v_3__1_), .S(npu_inst_pe_1_2_4_n4), .Z(
        npu_inst_pe_1_2_4_n24) );
  MUX2_X1 npu_inst_pe_1_2_4_U153 ( .A(npu_inst_pe_1_2_4_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_2_4_int_q_reg_v_5__1_), .S(npu_inst_pe_1_2_4_n4), .Z(
        npu_inst_pe_1_2_4_n23) );
  MUX2_X1 npu_inst_pe_1_2_4_U152 ( .A(npu_inst_pe_1_2_4_n22), .B(
        npu_inst_pe_1_2_4_n19), .S(npu_inst_pe_1_2_4_n8), .Z(
        npu_inst_int_data_x_2__4__1_) );
  MUX2_X1 npu_inst_pe_1_2_4_U151 ( .A(npu_inst_pe_1_2_4_n21), .B(
        npu_inst_pe_1_2_4_n20), .S(npu_inst_pe_1_2_4_n6), .Z(
        npu_inst_pe_1_2_4_n22) );
  MUX2_X1 npu_inst_pe_1_2_4_U150 ( .A(npu_inst_pe_1_2_4_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_2_4_int_q_reg_h_1__1_), .S(npu_inst_pe_1_2_4_n4), .Z(
        npu_inst_pe_1_2_4_n21) );
  MUX2_X1 npu_inst_pe_1_2_4_U149 ( .A(npu_inst_pe_1_2_4_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_2_4_int_q_reg_h_3__1_), .S(npu_inst_pe_1_2_4_n4), .Z(
        npu_inst_pe_1_2_4_n20) );
  MUX2_X1 npu_inst_pe_1_2_4_U148 ( .A(npu_inst_pe_1_2_4_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_2_4_int_q_reg_h_5__1_), .S(npu_inst_pe_1_2_4_n4), .Z(
        npu_inst_pe_1_2_4_n19) );
  MUX2_X1 npu_inst_pe_1_2_4_U147 ( .A(npu_inst_pe_1_2_4_n18), .B(
        npu_inst_pe_1_2_4_n15), .S(npu_inst_pe_1_2_4_n8), .Z(
        npu_inst_int_data_x_2__4__0_) );
  MUX2_X1 npu_inst_pe_1_2_4_U146 ( .A(npu_inst_pe_1_2_4_n17), .B(
        npu_inst_pe_1_2_4_n16), .S(npu_inst_pe_1_2_4_n6), .Z(
        npu_inst_pe_1_2_4_n18) );
  MUX2_X1 npu_inst_pe_1_2_4_U145 ( .A(npu_inst_pe_1_2_4_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_2_4_int_q_reg_h_1__0_), .S(npu_inst_pe_1_2_4_n4), .Z(
        npu_inst_pe_1_2_4_n17) );
  MUX2_X1 npu_inst_pe_1_2_4_U144 ( .A(npu_inst_pe_1_2_4_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_2_4_int_q_reg_h_3__0_), .S(npu_inst_pe_1_2_4_n4), .Z(
        npu_inst_pe_1_2_4_n16) );
  MUX2_X1 npu_inst_pe_1_2_4_U143 ( .A(npu_inst_pe_1_2_4_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_2_4_int_q_reg_h_5__0_), .S(npu_inst_pe_1_2_4_n4), .Z(
        npu_inst_pe_1_2_4_n15) );
  XOR2_X1 npu_inst_pe_1_2_4_U142 ( .A(npu_inst_pe_1_2_4_int_data_0_), .B(
        npu_inst_pe_1_2_4_int_q_acc_0_), .Z(npu_inst_pe_1_2_4_N73) );
  AND2_X1 npu_inst_pe_1_2_4_U141 ( .A1(npu_inst_pe_1_2_4_int_q_acc_0_), .A2(
        npu_inst_pe_1_2_4_int_data_0_), .ZN(npu_inst_pe_1_2_4_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_2_4_U140 ( .A(npu_inst_pe_1_2_4_int_q_acc_0_), .B(
        npu_inst_pe_1_2_4_n13), .ZN(npu_inst_pe_1_2_4_N65) );
  OR2_X1 npu_inst_pe_1_2_4_U139 ( .A1(npu_inst_pe_1_2_4_n13), .A2(
        npu_inst_pe_1_2_4_int_q_acc_0_), .ZN(npu_inst_pe_1_2_4_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_2_4_U138 ( .A(npu_inst_pe_1_2_4_int_q_acc_2_), .B(
        npu_inst_pe_1_2_4_add_79_carry_2_), .Z(npu_inst_pe_1_2_4_N75) );
  AND2_X1 npu_inst_pe_1_2_4_U137 ( .A1(npu_inst_pe_1_2_4_add_79_carry_2_), 
        .A2(npu_inst_pe_1_2_4_int_q_acc_2_), .ZN(
        npu_inst_pe_1_2_4_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_2_4_U136 ( .A(npu_inst_pe_1_2_4_int_q_acc_3_), .B(
        npu_inst_pe_1_2_4_add_79_carry_3_), .Z(npu_inst_pe_1_2_4_N76) );
  AND2_X1 npu_inst_pe_1_2_4_U135 ( .A1(npu_inst_pe_1_2_4_add_79_carry_3_), 
        .A2(npu_inst_pe_1_2_4_int_q_acc_3_), .ZN(
        npu_inst_pe_1_2_4_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_2_4_U134 ( .A(npu_inst_pe_1_2_4_int_q_acc_4_), .B(
        npu_inst_pe_1_2_4_add_79_carry_4_), .Z(npu_inst_pe_1_2_4_N77) );
  AND2_X1 npu_inst_pe_1_2_4_U133 ( .A1(npu_inst_pe_1_2_4_add_79_carry_4_), 
        .A2(npu_inst_pe_1_2_4_int_q_acc_4_), .ZN(
        npu_inst_pe_1_2_4_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_2_4_U132 ( .A(npu_inst_pe_1_2_4_int_q_acc_5_), .B(
        npu_inst_pe_1_2_4_add_79_carry_5_), .Z(npu_inst_pe_1_2_4_N78) );
  AND2_X1 npu_inst_pe_1_2_4_U131 ( .A1(npu_inst_pe_1_2_4_add_79_carry_5_), 
        .A2(npu_inst_pe_1_2_4_int_q_acc_5_), .ZN(
        npu_inst_pe_1_2_4_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_2_4_U130 ( .A(npu_inst_pe_1_2_4_int_q_acc_6_), .B(
        npu_inst_pe_1_2_4_add_79_carry_6_), .Z(npu_inst_pe_1_2_4_N79) );
  AND2_X1 npu_inst_pe_1_2_4_U129 ( .A1(npu_inst_pe_1_2_4_add_79_carry_6_), 
        .A2(npu_inst_pe_1_2_4_int_q_acc_6_), .ZN(
        npu_inst_pe_1_2_4_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_2_4_U128 ( .A(npu_inst_pe_1_2_4_int_q_acc_7_), .B(
        npu_inst_pe_1_2_4_add_79_carry_7_), .Z(npu_inst_pe_1_2_4_N80) );
  XNOR2_X1 npu_inst_pe_1_2_4_U127 ( .A(npu_inst_pe_1_2_4_sub_77_carry_2_), .B(
        npu_inst_pe_1_2_4_int_q_acc_2_), .ZN(npu_inst_pe_1_2_4_N67) );
  OR2_X1 npu_inst_pe_1_2_4_U126 ( .A1(npu_inst_pe_1_2_4_int_q_acc_2_), .A2(
        npu_inst_pe_1_2_4_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_2_4_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_2_4_U125 ( .A(npu_inst_pe_1_2_4_sub_77_carry_3_), .B(
        npu_inst_pe_1_2_4_int_q_acc_3_), .ZN(npu_inst_pe_1_2_4_N68) );
  OR2_X1 npu_inst_pe_1_2_4_U124 ( .A1(npu_inst_pe_1_2_4_int_q_acc_3_), .A2(
        npu_inst_pe_1_2_4_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_2_4_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_2_4_U123 ( .A(npu_inst_pe_1_2_4_sub_77_carry_4_), .B(
        npu_inst_pe_1_2_4_int_q_acc_4_), .ZN(npu_inst_pe_1_2_4_N69) );
  OR2_X1 npu_inst_pe_1_2_4_U122 ( .A1(npu_inst_pe_1_2_4_int_q_acc_4_), .A2(
        npu_inst_pe_1_2_4_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_2_4_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_2_4_U121 ( .A(npu_inst_pe_1_2_4_sub_77_carry_5_), .B(
        npu_inst_pe_1_2_4_int_q_acc_5_), .ZN(npu_inst_pe_1_2_4_N70) );
  OR2_X1 npu_inst_pe_1_2_4_U120 ( .A1(npu_inst_pe_1_2_4_int_q_acc_5_), .A2(
        npu_inst_pe_1_2_4_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_2_4_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_2_4_U119 ( .A(npu_inst_pe_1_2_4_sub_77_carry_6_), .B(
        npu_inst_pe_1_2_4_int_q_acc_6_), .ZN(npu_inst_pe_1_2_4_N71) );
  OR2_X1 npu_inst_pe_1_2_4_U118 ( .A1(npu_inst_pe_1_2_4_int_q_acc_6_), .A2(
        npu_inst_pe_1_2_4_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_2_4_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_2_4_U117 ( .A(npu_inst_pe_1_2_4_int_q_acc_7_), .B(
        npu_inst_pe_1_2_4_sub_77_carry_7_), .ZN(npu_inst_pe_1_2_4_N72) );
  INV_X1 npu_inst_pe_1_2_4_U116 ( .A(npu_inst_n78), .ZN(npu_inst_pe_1_2_4_n7)
         );
  INV_X1 npu_inst_pe_1_2_4_U115 ( .A(npu_inst_pe_1_2_4_n7), .ZN(
        npu_inst_pe_1_2_4_n6) );
  INV_X1 npu_inst_pe_1_2_4_U114 ( .A(npu_inst_n58), .ZN(npu_inst_pe_1_2_4_n3)
         );
  AOI22_X1 npu_inst_pe_1_2_4_U113 ( .A1(npu_inst_int_data_y_3__4__0_), .A2(
        npu_inst_pe_1_2_4_n58), .B1(npu_inst_pe_1_2_4_n114), .B2(
        npu_inst_pe_1_2_4_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_2_4_n57) );
  INV_X1 npu_inst_pe_1_2_4_U112 ( .A(npu_inst_pe_1_2_4_n57), .ZN(
        npu_inst_pe_1_2_4_n108) );
  AOI22_X1 npu_inst_pe_1_2_4_U111 ( .A1(npu_inst_int_data_y_3__4__0_), .A2(
        npu_inst_pe_1_2_4_n54), .B1(npu_inst_pe_1_2_4_n115), .B2(
        npu_inst_pe_1_2_4_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_2_4_n53) );
  INV_X1 npu_inst_pe_1_2_4_U110 ( .A(npu_inst_pe_1_2_4_n53), .ZN(
        npu_inst_pe_1_2_4_n109) );
  AOI22_X1 npu_inst_pe_1_2_4_U107 ( .A1(npu_inst_int_data_y_3__4__0_), .A2(
        npu_inst_pe_1_2_4_n50), .B1(npu_inst_pe_1_2_4_n116), .B2(
        npu_inst_pe_1_2_4_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_2_4_n49) );
  INV_X1 npu_inst_pe_1_2_4_U106 ( .A(npu_inst_pe_1_2_4_n49), .ZN(
        npu_inst_pe_1_2_4_n110) );
  AOI22_X1 npu_inst_pe_1_2_4_U105 ( .A1(npu_inst_int_data_y_3__4__0_), .A2(
        npu_inst_pe_1_2_4_n46), .B1(npu_inst_pe_1_2_4_n117), .B2(
        npu_inst_pe_1_2_4_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_2_4_n45) );
  INV_X1 npu_inst_pe_1_2_4_U104 ( .A(npu_inst_pe_1_2_4_n45), .ZN(
        npu_inst_pe_1_2_4_n111) );
  AOI22_X1 npu_inst_pe_1_2_4_U103 ( .A1(npu_inst_int_data_y_3__4__0_), .A2(
        npu_inst_pe_1_2_4_n42), .B1(npu_inst_pe_1_2_4_n119), .B2(
        npu_inst_pe_1_2_4_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_2_4_n41) );
  INV_X1 npu_inst_pe_1_2_4_U102 ( .A(npu_inst_pe_1_2_4_n41), .ZN(
        npu_inst_pe_1_2_4_n112) );
  AOI22_X1 npu_inst_pe_1_2_4_U101 ( .A1(npu_inst_int_data_y_3__4__1_), .A2(
        npu_inst_pe_1_2_4_n58), .B1(npu_inst_pe_1_2_4_n114), .B2(
        npu_inst_pe_1_2_4_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_2_4_n59) );
  INV_X1 npu_inst_pe_1_2_4_U100 ( .A(npu_inst_pe_1_2_4_n59), .ZN(
        npu_inst_pe_1_2_4_n102) );
  AOI22_X1 npu_inst_pe_1_2_4_U99 ( .A1(npu_inst_int_data_y_3__4__1_), .A2(
        npu_inst_pe_1_2_4_n54), .B1(npu_inst_pe_1_2_4_n115), .B2(
        npu_inst_pe_1_2_4_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_2_4_n55) );
  INV_X1 npu_inst_pe_1_2_4_U98 ( .A(npu_inst_pe_1_2_4_n55), .ZN(
        npu_inst_pe_1_2_4_n103) );
  AOI22_X1 npu_inst_pe_1_2_4_U97 ( .A1(npu_inst_int_data_y_3__4__1_), .A2(
        npu_inst_pe_1_2_4_n50), .B1(npu_inst_pe_1_2_4_n116), .B2(
        npu_inst_pe_1_2_4_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_2_4_n51) );
  INV_X1 npu_inst_pe_1_2_4_U96 ( .A(npu_inst_pe_1_2_4_n51), .ZN(
        npu_inst_pe_1_2_4_n104) );
  AOI22_X1 npu_inst_pe_1_2_4_U95 ( .A1(npu_inst_int_data_y_3__4__1_), .A2(
        npu_inst_pe_1_2_4_n46), .B1(npu_inst_pe_1_2_4_n117), .B2(
        npu_inst_pe_1_2_4_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_2_4_n47) );
  INV_X1 npu_inst_pe_1_2_4_U94 ( .A(npu_inst_pe_1_2_4_n47), .ZN(
        npu_inst_pe_1_2_4_n105) );
  AOI22_X1 npu_inst_pe_1_2_4_U93 ( .A1(npu_inst_int_data_y_3__4__1_), .A2(
        npu_inst_pe_1_2_4_n42), .B1(npu_inst_pe_1_2_4_n119), .B2(
        npu_inst_pe_1_2_4_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_2_4_n43) );
  INV_X1 npu_inst_pe_1_2_4_U92 ( .A(npu_inst_pe_1_2_4_n43), .ZN(
        npu_inst_pe_1_2_4_n106) );
  AOI22_X1 npu_inst_pe_1_2_4_U91 ( .A1(npu_inst_pe_1_2_4_n38), .A2(
        npu_inst_int_data_y_3__4__1_), .B1(npu_inst_pe_1_2_4_n118), .B2(
        npu_inst_pe_1_2_4_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_2_4_n39) );
  INV_X1 npu_inst_pe_1_2_4_U90 ( .A(npu_inst_pe_1_2_4_n39), .ZN(
        npu_inst_pe_1_2_4_n107) );
  AOI22_X1 npu_inst_pe_1_2_4_U89 ( .A1(npu_inst_pe_1_2_4_n38), .A2(
        npu_inst_int_data_y_3__4__0_), .B1(npu_inst_pe_1_2_4_n118), .B2(
        npu_inst_pe_1_2_4_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_2_4_n37) );
  INV_X1 npu_inst_pe_1_2_4_U88 ( .A(npu_inst_pe_1_2_4_n37), .ZN(
        npu_inst_pe_1_2_4_n113) );
  NAND2_X1 npu_inst_pe_1_2_4_U87 ( .A1(npu_inst_pe_1_2_4_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_2_4_n60), .ZN(npu_inst_pe_1_2_4_n74) );
  OAI21_X1 npu_inst_pe_1_2_4_U86 ( .B1(npu_inst_pe_1_2_4_n63), .B2(
        npu_inst_pe_1_2_4_n60), .A(npu_inst_pe_1_2_4_n74), .ZN(
        npu_inst_pe_1_2_4_n97) );
  NAND2_X1 npu_inst_pe_1_2_4_U85 ( .A1(npu_inst_pe_1_2_4_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_2_4_n60), .ZN(npu_inst_pe_1_2_4_n73) );
  OAI21_X1 npu_inst_pe_1_2_4_U84 ( .B1(npu_inst_pe_1_2_4_n61), .B2(
        npu_inst_pe_1_2_4_n60), .A(npu_inst_pe_1_2_4_n73), .ZN(
        npu_inst_pe_1_2_4_n96) );
  NAND2_X1 npu_inst_pe_1_2_4_U83 ( .A1(npu_inst_pe_1_2_4_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_2_4_n56), .ZN(npu_inst_pe_1_2_4_n72) );
  OAI21_X1 npu_inst_pe_1_2_4_U82 ( .B1(npu_inst_pe_1_2_4_n63), .B2(
        npu_inst_pe_1_2_4_n56), .A(npu_inst_pe_1_2_4_n72), .ZN(
        npu_inst_pe_1_2_4_n95) );
  NAND2_X1 npu_inst_pe_1_2_4_U81 ( .A1(npu_inst_pe_1_2_4_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_2_4_n56), .ZN(npu_inst_pe_1_2_4_n71) );
  OAI21_X1 npu_inst_pe_1_2_4_U80 ( .B1(npu_inst_pe_1_2_4_n61), .B2(
        npu_inst_pe_1_2_4_n56), .A(npu_inst_pe_1_2_4_n71), .ZN(
        npu_inst_pe_1_2_4_n94) );
  NAND2_X1 npu_inst_pe_1_2_4_U79 ( .A1(npu_inst_pe_1_2_4_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_2_4_n52), .ZN(npu_inst_pe_1_2_4_n70) );
  OAI21_X1 npu_inst_pe_1_2_4_U78 ( .B1(npu_inst_pe_1_2_4_n63), .B2(
        npu_inst_pe_1_2_4_n52), .A(npu_inst_pe_1_2_4_n70), .ZN(
        npu_inst_pe_1_2_4_n93) );
  NAND2_X1 npu_inst_pe_1_2_4_U77 ( .A1(npu_inst_pe_1_2_4_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_2_4_n52), .ZN(npu_inst_pe_1_2_4_n69) );
  OAI21_X1 npu_inst_pe_1_2_4_U76 ( .B1(npu_inst_pe_1_2_4_n61), .B2(
        npu_inst_pe_1_2_4_n52), .A(npu_inst_pe_1_2_4_n69), .ZN(
        npu_inst_pe_1_2_4_n92) );
  NAND2_X1 npu_inst_pe_1_2_4_U75 ( .A1(npu_inst_pe_1_2_4_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_2_4_n48), .ZN(npu_inst_pe_1_2_4_n68) );
  OAI21_X1 npu_inst_pe_1_2_4_U74 ( .B1(npu_inst_pe_1_2_4_n63), .B2(
        npu_inst_pe_1_2_4_n48), .A(npu_inst_pe_1_2_4_n68), .ZN(
        npu_inst_pe_1_2_4_n91) );
  NAND2_X1 npu_inst_pe_1_2_4_U73 ( .A1(npu_inst_pe_1_2_4_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_2_4_n48), .ZN(npu_inst_pe_1_2_4_n67) );
  OAI21_X1 npu_inst_pe_1_2_4_U72 ( .B1(npu_inst_pe_1_2_4_n61), .B2(
        npu_inst_pe_1_2_4_n48), .A(npu_inst_pe_1_2_4_n67), .ZN(
        npu_inst_pe_1_2_4_n90) );
  NAND2_X1 npu_inst_pe_1_2_4_U71 ( .A1(npu_inst_pe_1_2_4_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_2_4_n44), .ZN(npu_inst_pe_1_2_4_n66) );
  OAI21_X1 npu_inst_pe_1_2_4_U70 ( .B1(npu_inst_pe_1_2_4_n63), .B2(
        npu_inst_pe_1_2_4_n44), .A(npu_inst_pe_1_2_4_n66), .ZN(
        npu_inst_pe_1_2_4_n89) );
  NAND2_X1 npu_inst_pe_1_2_4_U69 ( .A1(npu_inst_pe_1_2_4_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_2_4_n44), .ZN(npu_inst_pe_1_2_4_n65) );
  OAI21_X1 npu_inst_pe_1_2_4_U68 ( .B1(npu_inst_pe_1_2_4_n61), .B2(
        npu_inst_pe_1_2_4_n44), .A(npu_inst_pe_1_2_4_n65), .ZN(
        npu_inst_pe_1_2_4_n88) );
  NAND2_X1 npu_inst_pe_1_2_4_U67 ( .A1(npu_inst_pe_1_2_4_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_2_4_n40), .ZN(npu_inst_pe_1_2_4_n64) );
  OAI21_X1 npu_inst_pe_1_2_4_U66 ( .B1(npu_inst_pe_1_2_4_n63), .B2(
        npu_inst_pe_1_2_4_n40), .A(npu_inst_pe_1_2_4_n64), .ZN(
        npu_inst_pe_1_2_4_n87) );
  NAND2_X1 npu_inst_pe_1_2_4_U65 ( .A1(npu_inst_pe_1_2_4_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_2_4_n40), .ZN(npu_inst_pe_1_2_4_n62) );
  OAI21_X1 npu_inst_pe_1_2_4_U64 ( .B1(npu_inst_pe_1_2_4_n61), .B2(
        npu_inst_pe_1_2_4_n40), .A(npu_inst_pe_1_2_4_n62), .ZN(
        npu_inst_pe_1_2_4_n86) );
  AND2_X1 npu_inst_pe_1_2_4_U63 ( .A1(npu_inst_pe_1_2_4_N93), .A2(npu_inst_n58), .ZN(npu_inst_int_data_y_2__4__0_) );
  AND2_X1 npu_inst_pe_1_2_4_U62 ( .A1(npu_inst_n58), .A2(npu_inst_pe_1_2_4_N94), .ZN(npu_inst_int_data_y_2__4__1_) );
  NOR3_X1 npu_inst_pe_1_2_4_U61 ( .A1(npu_inst_pe_1_2_4_n26), .A2(npu_inst_n58), .A3(npu_inst_int_ckg[43]), .ZN(npu_inst_pe_1_2_4_n85) );
  OR2_X1 npu_inst_pe_1_2_4_U60 ( .A1(npu_inst_pe_1_2_4_n85), .A2(
        npu_inst_pe_1_2_4_n2), .ZN(npu_inst_pe_1_2_4_N84) );
  AND2_X1 npu_inst_pe_1_2_4_U59 ( .A1(npu_inst_pe_1_2_4_int_q_acc_0_), .A2(
        npu_inst_pe_1_2_4_n1), .ZN(npu_inst_int_data_res_2__4__0_) );
  AND2_X1 npu_inst_pe_1_2_4_U58 ( .A1(npu_inst_pe_1_2_4_n2), .A2(
        npu_inst_pe_1_2_4_int_q_acc_7_), .ZN(npu_inst_int_data_res_2__4__7_)
         );
  AND2_X1 npu_inst_pe_1_2_4_U57 ( .A1(npu_inst_pe_1_2_4_int_q_acc_1_), .A2(
        npu_inst_pe_1_2_4_n1), .ZN(npu_inst_int_data_res_2__4__1_) );
  AND2_X1 npu_inst_pe_1_2_4_U56 ( .A1(npu_inst_pe_1_2_4_int_q_acc_2_), .A2(
        npu_inst_pe_1_2_4_n1), .ZN(npu_inst_int_data_res_2__4__2_) );
  AND2_X1 npu_inst_pe_1_2_4_U55 ( .A1(npu_inst_pe_1_2_4_int_q_acc_3_), .A2(
        npu_inst_pe_1_2_4_n2), .ZN(npu_inst_int_data_res_2__4__3_) );
  AND2_X1 npu_inst_pe_1_2_4_U54 ( .A1(npu_inst_pe_1_2_4_int_q_acc_4_), .A2(
        npu_inst_pe_1_2_4_n2), .ZN(npu_inst_int_data_res_2__4__4_) );
  AND2_X1 npu_inst_pe_1_2_4_U53 ( .A1(npu_inst_pe_1_2_4_int_q_acc_5_), .A2(
        npu_inst_pe_1_2_4_n2), .ZN(npu_inst_int_data_res_2__4__5_) );
  AND2_X1 npu_inst_pe_1_2_4_U52 ( .A1(npu_inst_pe_1_2_4_int_q_acc_6_), .A2(
        npu_inst_pe_1_2_4_n2), .ZN(npu_inst_int_data_res_2__4__6_) );
  AOI222_X1 npu_inst_pe_1_2_4_U51 ( .A1(npu_inst_int_data_res_3__4__0_), .A2(
        npu_inst_pe_1_2_4_n1), .B1(npu_inst_pe_1_2_4_N73), .B2(
        npu_inst_pe_1_2_4_n76), .C1(npu_inst_pe_1_2_4_N65), .C2(
        npu_inst_pe_1_2_4_n77), .ZN(npu_inst_pe_1_2_4_n84) );
  INV_X1 npu_inst_pe_1_2_4_U50 ( .A(npu_inst_pe_1_2_4_n84), .ZN(
        npu_inst_pe_1_2_4_n101) );
  AOI222_X1 npu_inst_pe_1_2_4_U49 ( .A1(npu_inst_int_data_res_3__4__7_), .A2(
        npu_inst_pe_1_2_4_n1), .B1(npu_inst_pe_1_2_4_N80), .B2(
        npu_inst_pe_1_2_4_n76), .C1(npu_inst_pe_1_2_4_N72), .C2(
        npu_inst_pe_1_2_4_n77), .ZN(npu_inst_pe_1_2_4_n75) );
  INV_X1 npu_inst_pe_1_2_4_U48 ( .A(npu_inst_pe_1_2_4_n75), .ZN(
        npu_inst_pe_1_2_4_n33) );
  AOI222_X1 npu_inst_pe_1_2_4_U47 ( .A1(npu_inst_int_data_res_3__4__1_), .A2(
        npu_inst_pe_1_2_4_n1), .B1(npu_inst_pe_1_2_4_N74), .B2(
        npu_inst_pe_1_2_4_n76), .C1(npu_inst_pe_1_2_4_N66), .C2(
        npu_inst_pe_1_2_4_n77), .ZN(npu_inst_pe_1_2_4_n83) );
  INV_X1 npu_inst_pe_1_2_4_U46 ( .A(npu_inst_pe_1_2_4_n83), .ZN(
        npu_inst_pe_1_2_4_n100) );
  AOI222_X1 npu_inst_pe_1_2_4_U45 ( .A1(npu_inst_int_data_res_3__4__2_), .A2(
        npu_inst_pe_1_2_4_n1), .B1(npu_inst_pe_1_2_4_N75), .B2(
        npu_inst_pe_1_2_4_n76), .C1(npu_inst_pe_1_2_4_N67), .C2(
        npu_inst_pe_1_2_4_n77), .ZN(npu_inst_pe_1_2_4_n82) );
  INV_X1 npu_inst_pe_1_2_4_U44 ( .A(npu_inst_pe_1_2_4_n82), .ZN(
        npu_inst_pe_1_2_4_n99) );
  AOI222_X1 npu_inst_pe_1_2_4_U43 ( .A1(npu_inst_int_data_res_3__4__3_), .A2(
        npu_inst_pe_1_2_4_n1), .B1(npu_inst_pe_1_2_4_N76), .B2(
        npu_inst_pe_1_2_4_n76), .C1(npu_inst_pe_1_2_4_N68), .C2(
        npu_inst_pe_1_2_4_n77), .ZN(npu_inst_pe_1_2_4_n81) );
  INV_X1 npu_inst_pe_1_2_4_U42 ( .A(npu_inst_pe_1_2_4_n81), .ZN(
        npu_inst_pe_1_2_4_n98) );
  AOI222_X1 npu_inst_pe_1_2_4_U41 ( .A1(npu_inst_int_data_res_3__4__4_), .A2(
        npu_inst_pe_1_2_4_n1), .B1(npu_inst_pe_1_2_4_N77), .B2(
        npu_inst_pe_1_2_4_n76), .C1(npu_inst_pe_1_2_4_N69), .C2(
        npu_inst_pe_1_2_4_n77), .ZN(npu_inst_pe_1_2_4_n80) );
  INV_X1 npu_inst_pe_1_2_4_U40 ( .A(npu_inst_pe_1_2_4_n80), .ZN(
        npu_inst_pe_1_2_4_n36) );
  AOI222_X1 npu_inst_pe_1_2_4_U39 ( .A1(npu_inst_int_data_res_3__4__5_), .A2(
        npu_inst_pe_1_2_4_n1), .B1(npu_inst_pe_1_2_4_N78), .B2(
        npu_inst_pe_1_2_4_n76), .C1(npu_inst_pe_1_2_4_N70), .C2(
        npu_inst_pe_1_2_4_n77), .ZN(npu_inst_pe_1_2_4_n79) );
  INV_X1 npu_inst_pe_1_2_4_U38 ( .A(npu_inst_pe_1_2_4_n79), .ZN(
        npu_inst_pe_1_2_4_n35) );
  AOI222_X1 npu_inst_pe_1_2_4_U37 ( .A1(npu_inst_int_data_res_3__4__6_), .A2(
        npu_inst_pe_1_2_4_n1), .B1(npu_inst_pe_1_2_4_N79), .B2(
        npu_inst_pe_1_2_4_n76), .C1(npu_inst_pe_1_2_4_N71), .C2(
        npu_inst_pe_1_2_4_n77), .ZN(npu_inst_pe_1_2_4_n78) );
  INV_X1 npu_inst_pe_1_2_4_U36 ( .A(npu_inst_pe_1_2_4_n78), .ZN(
        npu_inst_pe_1_2_4_n34) );
  INV_X1 npu_inst_pe_1_2_4_U35 ( .A(npu_inst_pe_1_2_4_int_data_1_), .ZN(
        npu_inst_pe_1_2_4_n14) );
  AND2_X1 npu_inst_pe_1_2_4_U34 ( .A1(npu_inst_int_data_x_2__4__1_), .A2(
        npu_inst_pe_1_2_4_int_q_weight_1_), .ZN(npu_inst_pe_1_2_4_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_2_4_U33 ( .A1(npu_inst_int_data_x_2__4__0_), .A2(
        npu_inst_pe_1_2_4_int_q_weight_1_), .ZN(npu_inst_pe_1_2_4_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_2_4_U32 ( .A1(npu_inst_n58), .A2(
        npu_inst_int_data_y_3__4__1_), .B1(npu_inst_pe_1_2_4_n3), .B2(
        npu_inst_int_data_x_2__5__1_), .ZN(npu_inst_pe_1_2_4_n63) );
  AOI22_X1 npu_inst_pe_1_2_4_U31 ( .A1(npu_inst_n58), .A2(
        npu_inst_int_data_y_3__4__0_), .B1(npu_inst_pe_1_2_4_n3), .B2(
        npu_inst_int_data_x_2__5__0_), .ZN(npu_inst_pe_1_2_4_n61) );
  INV_X1 npu_inst_pe_1_2_4_U30 ( .A(npu_inst_pe_1_2_4_int_data_0_), .ZN(
        npu_inst_pe_1_2_4_n13) );
  INV_X1 npu_inst_pe_1_2_4_U29 ( .A(npu_inst_n70), .ZN(npu_inst_pe_1_2_4_n5)
         );
  OR3_X1 npu_inst_pe_1_2_4_U28 ( .A1(npu_inst_pe_1_2_4_n6), .A2(
        npu_inst_pe_1_2_4_n8), .A3(npu_inst_pe_1_2_4_n5), .ZN(
        npu_inst_pe_1_2_4_n56) );
  OR3_X1 npu_inst_pe_1_2_4_U27 ( .A1(npu_inst_pe_1_2_4_n5), .A2(
        npu_inst_pe_1_2_4_n8), .A3(npu_inst_pe_1_2_4_n7), .ZN(
        npu_inst_pe_1_2_4_n48) );
  INV_X1 npu_inst_pe_1_2_4_U26 ( .A(npu_inst_pe_1_2_4_n5), .ZN(
        npu_inst_pe_1_2_4_n4) );
  INV_X1 npu_inst_pe_1_2_4_U25 ( .A(npu_inst_n125), .ZN(npu_inst_pe_1_2_4_n12)
         );
  OR3_X1 npu_inst_pe_1_2_4_U24 ( .A1(npu_inst_pe_1_2_4_n4), .A2(
        npu_inst_pe_1_2_4_n8), .A3(npu_inst_pe_1_2_4_n7), .ZN(
        npu_inst_pe_1_2_4_n52) );
  OR3_X1 npu_inst_pe_1_2_4_U23 ( .A1(npu_inst_pe_1_2_4_n6), .A2(
        npu_inst_pe_1_2_4_n8), .A3(npu_inst_pe_1_2_4_n4), .ZN(
        npu_inst_pe_1_2_4_n60) );
  NOR2_X1 npu_inst_pe_1_2_4_U22 ( .A1(npu_inst_pe_1_2_4_n60), .A2(
        npu_inst_pe_1_2_4_n3), .ZN(npu_inst_pe_1_2_4_n58) );
  NOR2_X1 npu_inst_pe_1_2_4_U21 ( .A1(npu_inst_pe_1_2_4_n56), .A2(
        npu_inst_pe_1_2_4_n3), .ZN(npu_inst_pe_1_2_4_n54) );
  NOR2_X1 npu_inst_pe_1_2_4_U20 ( .A1(npu_inst_pe_1_2_4_n52), .A2(
        npu_inst_pe_1_2_4_n3), .ZN(npu_inst_pe_1_2_4_n50) );
  NOR2_X1 npu_inst_pe_1_2_4_U19 ( .A1(npu_inst_pe_1_2_4_n48), .A2(
        npu_inst_pe_1_2_4_n3), .ZN(npu_inst_pe_1_2_4_n46) );
  NOR2_X1 npu_inst_pe_1_2_4_U18 ( .A1(npu_inst_pe_1_2_4_n40), .A2(
        npu_inst_pe_1_2_4_n3), .ZN(npu_inst_pe_1_2_4_n38) );
  NOR2_X1 npu_inst_pe_1_2_4_U17 ( .A1(npu_inst_pe_1_2_4_n44), .A2(
        npu_inst_pe_1_2_4_n3), .ZN(npu_inst_pe_1_2_4_n42) );
  BUF_X1 npu_inst_pe_1_2_4_U16 ( .A(npu_inst_n102), .Z(npu_inst_pe_1_2_4_n8)
         );
  BUF_X1 npu_inst_pe_1_2_4_U15 ( .A(npu_inst_pe_1_2_4_n12), .Z(
        npu_inst_pe_1_2_4_n11) );
  BUF_X1 npu_inst_pe_1_2_4_U14 ( .A(npu_inst_pe_1_2_4_n12), .Z(
        npu_inst_pe_1_2_4_n10) );
  BUF_X1 npu_inst_pe_1_2_4_U13 ( .A(npu_inst_pe_1_2_4_n12), .Z(
        npu_inst_pe_1_2_4_n9) );
  INV_X1 npu_inst_pe_1_2_4_U12 ( .A(npu_inst_pe_1_2_4_n38), .ZN(
        npu_inst_pe_1_2_4_n118) );
  INV_X1 npu_inst_pe_1_2_4_U11 ( .A(npu_inst_pe_1_2_4_n58), .ZN(
        npu_inst_pe_1_2_4_n114) );
  INV_X1 npu_inst_pe_1_2_4_U10 ( .A(npu_inst_pe_1_2_4_n54), .ZN(
        npu_inst_pe_1_2_4_n115) );
  INV_X1 npu_inst_pe_1_2_4_U9 ( .A(npu_inst_pe_1_2_4_n50), .ZN(
        npu_inst_pe_1_2_4_n116) );
  INV_X1 npu_inst_pe_1_2_4_U8 ( .A(npu_inst_pe_1_2_4_n46), .ZN(
        npu_inst_pe_1_2_4_n117) );
  INV_X1 npu_inst_pe_1_2_4_U7 ( .A(npu_inst_pe_1_2_4_n42), .ZN(
        npu_inst_pe_1_2_4_n119) );
  BUF_X1 npu_inst_pe_1_2_4_U6 ( .A(npu_inst_n28), .Z(npu_inst_pe_1_2_4_n2) );
  BUF_X1 npu_inst_pe_1_2_4_U5 ( .A(npu_inst_n28), .Z(npu_inst_pe_1_2_4_n1) );
  NOR2_X1 npu_inst_pe_1_2_4_U4 ( .A1(npu_inst_pe_1_2_4_int_q_weight_0_), .A2(
        npu_inst_pe_1_2_4_n1), .ZN(npu_inst_pe_1_2_4_n76) );
  NOR2_X1 npu_inst_pe_1_2_4_U3 ( .A1(npu_inst_pe_1_2_4_n27), .A2(
        npu_inst_pe_1_2_4_n1), .ZN(npu_inst_pe_1_2_4_n77) );
  FA_X1 npu_inst_pe_1_2_4_sub_77_U2_1 ( .A(npu_inst_pe_1_2_4_int_q_acc_1_), 
        .B(npu_inst_pe_1_2_4_n14), .CI(npu_inst_pe_1_2_4_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_2_4_sub_77_carry_2_), .S(npu_inst_pe_1_2_4_N66) );
  FA_X1 npu_inst_pe_1_2_4_add_79_U1_1 ( .A(npu_inst_pe_1_2_4_int_q_acc_1_), 
        .B(npu_inst_pe_1_2_4_int_data_1_), .CI(
        npu_inst_pe_1_2_4_add_79_carry_1_), .CO(
        npu_inst_pe_1_2_4_add_79_carry_2_), .S(npu_inst_pe_1_2_4_N74) );
  NAND3_X1 npu_inst_pe_1_2_4_U109 ( .A1(npu_inst_pe_1_2_4_n5), .A2(
        npu_inst_pe_1_2_4_n7), .A3(npu_inst_pe_1_2_4_n8), .ZN(
        npu_inst_pe_1_2_4_n44) );
  NAND3_X1 npu_inst_pe_1_2_4_U108 ( .A1(npu_inst_pe_1_2_4_n4), .A2(
        npu_inst_pe_1_2_4_n7), .A3(npu_inst_pe_1_2_4_n8), .ZN(
        npu_inst_pe_1_2_4_n40) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_2_4_n34), .CK(
        npu_inst_pe_1_2_4_net3833), .RN(npu_inst_pe_1_2_4_n9), .Q(
        npu_inst_pe_1_2_4_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_2_4_n35), .CK(
        npu_inst_pe_1_2_4_net3833), .RN(npu_inst_pe_1_2_4_n9), .Q(
        npu_inst_pe_1_2_4_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_2_4_n36), .CK(
        npu_inst_pe_1_2_4_net3833), .RN(npu_inst_pe_1_2_4_n9), .Q(
        npu_inst_pe_1_2_4_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_2_4_n98), .CK(
        npu_inst_pe_1_2_4_net3833), .RN(npu_inst_pe_1_2_4_n9), .Q(
        npu_inst_pe_1_2_4_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_2_4_n99), .CK(
        npu_inst_pe_1_2_4_net3833), .RN(npu_inst_pe_1_2_4_n9), .Q(
        npu_inst_pe_1_2_4_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_2_4_n100), 
        .CK(npu_inst_pe_1_2_4_net3833), .RN(npu_inst_pe_1_2_4_n9), .Q(
        npu_inst_pe_1_2_4_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_2_4_n33), .CK(
        npu_inst_pe_1_2_4_net3833), .RN(npu_inst_pe_1_2_4_n9), .Q(
        npu_inst_pe_1_2_4_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_2_4_n101), 
        .CK(npu_inst_pe_1_2_4_net3833), .RN(npu_inst_pe_1_2_4_n9), .Q(
        npu_inst_pe_1_2_4_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_weight_reg_0_ ( .D(npu_inst_n111), .CK(
        npu_inst_pe_1_2_4_net3839), .RN(npu_inst_pe_1_2_4_n9), .Q(
        npu_inst_pe_1_2_4_int_q_weight_0_), .QN(npu_inst_pe_1_2_4_n27) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_weight_reg_1_ ( .D(npu_inst_n117), .CK(
        npu_inst_pe_1_2_4_net3839), .RN(npu_inst_pe_1_2_4_n9), .Q(
        npu_inst_pe_1_2_4_int_q_weight_1_), .QN(npu_inst_pe_1_2_4_n26) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_2_4_n113), 
        .CK(npu_inst_pe_1_2_4_net3839), .RN(npu_inst_pe_1_2_4_n9), .Q(
        npu_inst_pe_1_2_4_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_2_4_n107), 
        .CK(npu_inst_pe_1_2_4_net3839), .RN(npu_inst_pe_1_2_4_n9), .Q(
        npu_inst_pe_1_2_4_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_2_4_n112), 
        .CK(npu_inst_pe_1_2_4_net3839), .RN(npu_inst_pe_1_2_4_n10), .Q(
        npu_inst_pe_1_2_4_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_2_4_n106), 
        .CK(npu_inst_pe_1_2_4_net3839), .RN(npu_inst_pe_1_2_4_n10), .Q(
        npu_inst_pe_1_2_4_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_2_4_n111), 
        .CK(npu_inst_pe_1_2_4_net3839), .RN(npu_inst_pe_1_2_4_n10), .Q(
        npu_inst_pe_1_2_4_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_2_4_n105), 
        .CK(npu_inst_pe_1_2_4_net3839), .RN(npu_inst_pe_1_2_4_n10), .Q(
        npu_inst_pe_1_2_4_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_2_4_n110), 
        .CK(npu_inst_pe_1_2_4_net3839), .RN(npu_inst_pe_1_2_4_n10), .Q(
        npu_inst_pe_1_2_4_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_2_4_n104), 
        .CK(npu_inst_pe_1_2_4_net3839), .RN(npu_inst_pe_1_2_4_n10), .Q(
        npu_inst_pe_1_2_4_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_2_4_n109), 
        .CK(npu_inst_pe_1_2_4_net3839), .RN(npu_inst_pe_1_2_4_n10), .Q(
        npu_inst_pe_1_2_4_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_2_4_n103), 
        .CK(npu_inst_pe_1_2_4_net3839), .RN(npu_inst_pe_1_2_4_n10), .Q(
        npu_inst_pe_1_2_4_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_2_4_n108), 
        .CK(npu_inst_pe_1_2_4_net3839), .RN(npu_inst_pe_1_2_4_n10), .Q(
        npu_inst_pe_1_2_4_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_2_4_n102), 
        .CK(npu_inst_pe_1_2_4_net3839), .RN(npu_inst_pe_1_2_4_n10), .Q(
        npu_inst_pe_1_2_4_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_2_4_n86), 
        .CK(npu_inst_pe_1_2_4_net3839), .RN(npu_inst_pe_1_2_4_n10), .Q(
        npu_inst_pe_1_2_4_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_2_4_n87), 
        .CK(npu_inst_pe_1_2_4_net3839), .RN(npu_inst_pe_1_2_4_n10), .Q(
        npu_inst_pe_1_2_4_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_2_4_n88), 
        .CK(npu_inst_pe_1_2_4_net3839), .RN(npu_inst_pe_1_2_4_n11), .Q(
        npu_inst_pe_1_2_4_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_2_4_n89), 
        .CK(npu_inst_pe_1_2_4_net3839), .RN(npu_inst_pe_1_2_4_n11), .Q(
        npu_inst_pe_1_2_4_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_2_4_n90), 
        .CK(npu_inst_pe_1_2_4_net3839), .RN(npu_inst_pe_1_2_4_n11), .Q(
        npu_inst_pe_1_2_4_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_2_4_n91), 
        .CK(npu_inst_pe_1_2_4_net3839), .RN(npu_inst_pe_1_2_4_n11), .Q(
        npu_inst_pe_1_2_4_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_2_4_n92), 
        .CK(npu_inst_pe_1_2_4_net3839), .RN(npu_inst_pe_1_2_4_n11), .Q(
        npu_inst_pe_1_2_4_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_2_4_n93), 
        .CK(npu_inst_pe_1_2_4_net3839), .RN(npu_inst_pe_1_2_4_n11), .Q(
        npu_inst_pe_1_2_4_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_2_4_n94), 
        .CK(npu_inst_pe_1_2_4_net3839), .RN(npu_inst_pe_1_2_4_n11), .Q(
        npu_inst_pe_1_2_4_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_2_4_n95), 
        .CK(npu_inst_pe_1_2_4_net3839), .RN(npu_inst_pe_1_2_4_n11), .Q(
        npu_inst_pe_1_2_4_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_2_4_n96), 
        .CK(npu_inst_pe_1_2_4_net3839), .RN(npu_inst_pe_1_2_4_n11), .Q(
        npu_inst_pe_1_2_4_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_2_4_n97), 
        .CK(npu_inst_pe_1_2_4_net3839), .RN(npu_inst_pe_1_2_4_n11), .Q(
        npu_inst_pe_1_2_4_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_2_4_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_2_4_N84), .SE(1'b0), .GCK(npu_inst_pe_1_2_4_net3833) );
  CLKGATETST_X1 npu_inst_pe_1_2_4_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n64), .SE(1'b0), .GCK(npu_inst_pe_1_2_4_net3839) );
  MUX2_X1 npu_inst_pe_1_2_5_U162 ( .A(npu_inst_pe_1_2_5_n32), .B(
        npu_inst_pe_1_2_5_n29), .S(npu_inst_pe_1_2_5_n8), .Z(
        npu_inst_pe_1_2_5_N93) );
  MUX2_X1 npu_inst_pe_1_2_5_U161 ( .A(npu_inst_pe_1_2_5_n31), .B(
        npu_inst_pe_1_2_5_n30), .S(npu_inst_pe_1_2_5_n6), .Z(
        npu_inst_pe_1_2_5_n32) );
  MUX2_X1 npu_inst_pe_1_2_5_U160 ( .A(npu_inst_pe_1_2_5_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_2_5_int_q_reg_v_1__0_), .S(npu_inst_pe_1_2_5_n4), .Z(
        npu_inst_pe_1_2_5_n31) );
  MUX2_X1 npu_inst_pe_1_2_5_U159 ( .A(npu_inst_pe_1_2_5_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_2_5_int_q_reg_v_3__0_), .S(npu_inst_pe_1_2_5_n4), .Z(
        npu_inst_pe_1_2_5_n30) );
  MUX2_X1 npu_inst_pe_1_2_5_U158 ( .A(npu_inst_pe_1_2_5_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_2_5_int_q_reg_v_5__0_), .S(npu_inst_pe_1_2_5_n4), .Z(
        npu_inst_pe_1_2_5_n29) );
  MUX2_X1 npu_inst_pe_1_2_5_U157 ( .A(npu_inst_pe_1_2_5_n28), .B(
        npu_inst_pe_1_2_5_n23), .S(npu_inst_pe_1_2_5_n8), .Z(
        npu_inst_pe_1_2_5_N94) );
  MUX2_X1 npu_inst_pe_1_2_5_U156 ( .A(npu_inst_pe_1_2_5_n25), .B(
        npu_inst_pe_1_2_5_n24), .S(npu_inst_pe_1_2_5_n6), .Z(
        npu_inst_pe_1_2_5_n28) );
  MUX2_X1 npu_inst_pe_1_2_5_U155 ( .A(npu_inst_pe_1_2_5_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_2_5_int_q_reg_v_1__1_), .S(npu_inst_pe_1_2_5_n4), .Z(
        npu_inst_pe_1_2_5_n25) );
  MUX2_X1 npu_inst_pe_1_2_5_U154 ( .A(npu_inst_pe_1_2_5_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_2_5_int_q_reg_v_3__1_), .S(npu_inst_pe_1_2_5_n4), .Z(
        npu_inst_pe_1_2_5_n24) );
  MUX2_X1 npu_inst_pe_1_2_5_U153 ( .A(npu_inst_pe_1_2_5_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_2_5_int_q_reg_v_5__1_), .S(npu_inst_pe_1_2_5_n4), .Z(
        npu_inst_pe_1_2_5_n23) );
  MUX2_X1 npu_inst_pe_1_2_5_U152 ( .A(npu_inst_pe_1_2_5_n22), .B(
        npu_inst_pe_1_2_5_n19), .S(npu_inst_pe_1_2_5_n8), .Z(
        npu_inst_int_data_x_2__5__1_) );
  MUX2_X1 npu_inst_pe_1_2_5_U151 ( .A(npu_inst_pe_1_2_5_n21), .B(
        npu_inst_pe_1_2_5_n20), .S(npu_inst_pe_1_2_5_n6), .Z(
        npu_inst_pe_1_2_5_n22) );
  MUX2_X1 npu_inst_pe_1_2_5_U150 ( .A(npu_inst_pe_1_2_5_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_2_5_int_q_reg_h_1__1_), .S(npu_inst_pe_1_2_5_n4), .Z(
        npu_inst_pe_1_2_5_n21) );
  MUX2_X1 npu_inst_pe_1_2_5_U149 ( .A(npu_inst_pe_1_2_5_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_2_5_int_q_reg_h_3__1_), .S(npu_inst_pe_1_2_5_n4), .Z(
        npu_inst_pe_1_2_5_n20) );
  MUX2_X1 npu_inst_pe_1_2_5_U148 ( .A(npu_inst_pe_1_2_5_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_2_5_int_q_reg_h_5__1_), .S(npu_inst_pe_1_2_5_n4), .Z(
        npu_inst_pe_1_2_5_n19) );
  MUX2_X1 npu_inst_pe_1_2_5_U147 ( .A(npu_inst_pe_1_2_5_n18), .B(
        npu_inst_pe_1_2_5_n15), .S(npu_inst_pe_1_2_5_n8), .Z(
        npu_inst_int_data_x_2__5__0_) );
  MUX2_X1 npu_inst_pe_1_2_5_U146 ( .A(npu_inst_pe_1_2_5_n17), .B(
        npu_inst_pe_1_2_5_n16), .S(npu_inst_pe_1_2_5_n6), .Z(
        npu_inst_pe_1_2_5_n18) );
  MUX2_X1 npu_inst_pe_1_2_5_U145 ( .A(npu_inst_pe_1_2_5_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_2_5_int_q_reg_h_1__0_), .S(npu_inst_pe_1_2_5_n4), .Z(
        npu_inst_pe_1_2_5_n17) );
  MUX2_X1 npu_inst_pe_1_2_5_U144 ( .A(npu_inst_pe_1_2_5_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_2_5_int_q_reg_h_3__0_), .S(npu_inst_pe_1_2_5_n4), .Z(
        npu_inst_pe_1_2_5_n16) );
  MUX2_X1 npu_inst_pe_1_2_5_U143 ( .A(npu_inst_pe_1_2_5_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_2_5_int_q_reg_h_5__0_), .S(npu_inst_pe_1_2_5_n4), .Z(
        npu_inst_pe_1_2_5_n15) );
  XOR2_X1 npu_inst_pe_1_2_5_U142 ( .A(npu_inst_pe_1_2_5_int_data_0_), .B(
        npu_inst_pe_1_2_5_int_q_acc_0_), .Z(npu_inst_pe_1_2_5_N73) );
  AND2_X1 npu_inst_pe_1_2_5_U141 ( .A1(npu_inst_pe_1_2_5_int_q_acc_0_), .A2(
        npu_inst_pe_1_2_5_int_data_0_), .ZN(npu_inst_pe_1_2_5_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_2_5_U140 ( .A(npu_inst_pe_1_2_5_int_q_acc_0_), .B(
        npu_inst_pe_1_2_5_n13), .ZN(npu_inst_pe_1_2_5_N65) );
  OR2_X1 npu_inst_pe_1_2_5_U139 ( .A1(npu_inst_pe_1_2_5_n13), .A2(
        npu_inst_pe_1_2_5_int_q_acc_0_), .ZN(npu_inst_pe_1_2_5_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_2_5_U138 ( .A(npu_inst_pe_1_2_5_int_q_acc_2_), .B(
        npu_inst_pe_1_2_5_add_79_carry_2_), .Z(npu_inst_pe_1_2_5_N75) );
  AND2_X1 npu_inst_pe_1_2_5_U137 ( .A1(npu_inst_pe_1_2_5_add_79_carry_2_), 
        .A2(npu_inst_pe_1_2_5_int_q_acc_2_), .ZN(
        npu_inst_pe_1_2_5_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_2_5_U136 ( .A(npu_inst_pe_1_2_5_int_q_acc_3_), .B(
        npu_inst_pe_1_2_5_add_79_carry_3_), .Z(npu_inst_pe_1_2_5_N76) );
  AND2_X1 npu_inst_pe_1_2_5_U135 ( .A1(npu_inst_pe_1_2_5_add_79_carry_3_), 
        .A2(npu_inst_pe_1_2_5_int_q_acc_3_), .ZN(
        npu_inst_pe_1_2_5_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_2_5_U134 ( .A(npu_inst_pe_1_2_5_int_q_acc_4_), .B(
        npu_inst_pe_1_2_5_add_79_carry_4_), .Z(npu_inst_pe_1_2_5_N77) );
  AND2_X1 npu_inst_pe_1_2_5_U133 ( .A1(npu_inst_pe_1_2_5_add_79_carry_4_), 
        .A2(npu_inst_pe_1_2_5_int_q_acc_4_), .ZN(
        npu_inst_pe_1_2_5_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_2_5_U132 ( .A(npu_inst_pe_1_2_5_int_q_acc_5_), .B(
        npu_inst_pe_1_2_5_add_79_carry_5_), .Z(npu_inst_pe_1_2_5_N78) );
  AND2_X1 npu_inst_pe_1_2_5_U131 ( .A1(npu_inst_pe_1_2_5_add_79_carry_5_), 
        .A2(npu_inst_pe_1_2_5_int_q_acc_5_), .ZN(
        npu_inst_pe_1_2_5_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_2_5_U130 ( .A(npu_inst_pe_1_2_5_int_q_acc_6_), .B(
        npu_inst_pe_1_2_5_add_79_carry_6_), .Z(npu_inst_pe_1_2_5_N79) );
  AND2_X1 npu_inst_pe_1_2_5_U129 ( .A1(npu_inst_pe_1_2_5_add_79_carry_6_), 
        .A2(npu_inst_pe_1_2_5_int_q_acc_6_), .ZN(
        npu_inst_pe_1_2_5_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_2_5_U128 ( .A(npu_inst_pe_1_2_5_int_q_acc_7_), .B(
        npu_inst_pe_1_2_5_add_79_carry_7_), .Z(npu_inst_pe_1_2_5_N80) );
  XNOR2_X1 npu_inst_pe_1_2_5_U127 ( .A(npu_inst_pe_1_2_5_sub_77_carry_2_), .B(
        npu_inst_pe_1_2_5_int_q_acc_2_), .ZN(npu_inst_pe_1_2_5_N67) );
  OR2_X1 npu_inst_pe_1_2_5_U126 ( .A1(npu_inst_pe_1_2_5_int_q_acc_2_), .A2(
        npu_inst_pe_1_2_5_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_2_5_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_2_5_U125 ( .A(npu_inst_pe_1_2_5_sub_77_carry_3_), .B(
        npu_inst_pe_1_2_5_int_q_acc_3_), .ZN(npu_inst_pe_1_2_5_N68) );
  OR2_X1 npu_inst_pe_1_2_5_U124 ( .A1(npu_inst_pe_1_2_5_int_q_acc_3_), .A2(
        npu_inst_pe_1_2_5_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_2_5_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_2_5_U123 ( .A(npu_inst_pe_1_2_5_sub_77_carry_4_), .B(
        npu_inst_pe_1_2_5_int_q_acc_4_), .ZN(npu_inst_pe_1_2_5_N69) );
  OR2_X1 npu_inst_pe_1_2_5_U122 ( .A1(npu_inst_pe_1_2_5_int_q_acc_4_), .A2(
        npu_inst_pe_1_2_5_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_2_5_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_2_5_U121 ( .A(npu_inst_pe_1_2_5_sub_77_carry_5_), .B(
        npu_inst_pe_1_2_5_int_q_acc_5_), .ZN(npu_inst_pe_1_2_5_N70) );
  OR2_X1 npu_inst_pe_1_2_5_U120 ( .A1(npu_inst_pe_1_2_5_int_q_acc_5_), .A2(
        npu_inst_pe_1_2_5_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_2_5_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_2_5_U119 ( .A(npu_inst_pe_1_2_5_sub_77_carry_6_), .B(
        npu_inst_pe_1_2_5_int_q_acc_6_), .ZN(npu_inst_pe_1_2_5_N71) );
  OR2_X1 npu_inst_pe_1_2_5_U118 ( .A1(npu_inst_pe_1_2_5_int_q_acc_6_), .A2(
        npu_inst_pe_1_2_5_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_2_5_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_2_5_U117 ( .A(npu_inst_pe_1_2_5_int_q_acc_7_), .B(
        npu_inst_pe_1_2_5_sub_77_carry_7_), .ZN(npu_inst_pe_1_2_5_N72) );
  INV_X1 npu_inst_pe_1_2_5_U116 ( .A(npu_inst_n78), .ZN(npu_inst_pe_1_2_5_n7)
         );
  INV_X1 npu_inst_pe_1_2_5_U115 ( .A(npu_inst_pe_1_2_5_n7), .ZN(
        npu_inst_pe_1_2_5_n6) );
  INV_X1 npu_inst_pe_1_2_5_U114 ( .A(npu_inst_n58), .ZN(npu_inst_pe_1_2_5_n3)
         );
  AOI22_X1 npu_inst_pe_1_2_5_U113 ( .A1(npu_inst_int_data_y_3__5__0_), .A2(
        npu_inst_pe_1_2_5_n58), .B1(npu_inst_pe_1_2_5_n114), .B2(
        npu_inst_pe_1_2_5_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_2_5_n57) );
  INV_X1 npu_inst_pe_1_2_5_U112 ( .A(npu_inst_pe_1_2_5_n57), .ZN(
        npu_inst_pe_1_2_5_n108) );
  AOI22_X1 npu_inst_pe_1_2_5_U111 ( .A1(npu_inst_int_data_y_3__5__0_), .A2(
        npu_inst_pe_1_2_5_n54), .B1(npu_inst_pe_1_2_5_n115), .B2(
        npu_inst_pe_1_2_5_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_2_5_n53) );
  INV_X1 npu_inst_pe_1_2_5_U110 ( .A(npu_inst_pe_1_2_5_n53), .ZN(
        npu_inst_pe_1_2_5_n109) );
  AOI22_X1 npu_inst_pe_1_2_5_U107 ( .A1(npu_inst_int_data_y_3__5__0_), .A2(
        npu_inst_pe_1_2_5_n50), .B1(npu_inst_pe_1_2_5_n116), .B2(
        npu_inst_pe_1_2_5_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_2_5_n49) );
  INV_X1 npu_inst_pe_1_2_5_U106 ( .A(npu_inst_pe_1_2_5_n49), .ZN(
        npu_inst_pe_1_2_5_n110) );
  AOI22_X1 npu_inst_pe_1_2_5_U105 ( .A1(npu_inst_int_data_y_3__5__0_), .A2(
        npu_inst_pe_1_2_5_n46), .B1(npu_inst_pe_1_2_5_n117), .B2(
        npu_inst_pe_1_2_5_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_2_5_n45) );
  INV_X1 npu_inst_pe_1_2_5_U104 ( .A(npu_inst_pe_1_2_5_n45), .ZN(
        npu_inst_pe_1_2_5_n111) );
  AOI22_X1 npu_inst_pe_1_2_5_U103 ( .A1(npu_inst_int_data_y_3__5__0_), .A2(
        npu_inst_pe_1_2_5_n42), .B1(npu_inst_pe_1_2_5_n119), .B2(
        npu_inst_pe_1_2_5_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_2_5_n41) );
  INV_X1 npu_inst_pe_1_2_5_U102 ( .A(npu_inst_pe_1_2_5_n41), .ZN(
        npu_inst_pe_1_2_5_n112) );
  AOI22_X1 npu_inst_pe_1_2_5_U101 ( .A1(npu_inst_int_data_y_3__5__1_), .A2(
        npu_inst_pe_1_2_5_n58), .B1(npu_inst_pe_1_2_5_n114), .B2(
        npu_inst_pe_1_2_5_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_2_5_n59) );
  INV_X1 npu_inst_pe_1_2_5_U100 ( .A(npu_inst_pe_1_2_5_n59), .ZN(
        npu_inst_pe_1_2_5_n102) );
  AOI22_X1 npu_inst_pe_1_2_5_U99 ( .A1(npu_inst_int_data_y_3__5__1_), .A2(
        npu_inst_pe_1_2_5_n54), .B1(npu_inst_pe_1_2_5_n115), .B2(
        npu_inst_pe_1_2_5_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_2_5_n55) );
  INV_X1 npu_inst_pe_1_2_5_U98 ( .A(npu_inst_pe_1_2_5_n55), .ZN(
        npu_inst_pe_1_2_5_n103) );
  AOI22_X1 npu_inst_pe_1_2_5_U97 ( .A1(npu_inst_int_data_y_3__5__1_), .A2(
        npu_inst_pe_1_2_5_n50), .B1(npu_inst_pe_1_2_5_n116), .B2(
        npu_inst_pe_1_2_5_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_2_5_n51) );
  INV_X1 npu_inst_pe_1_2_5_U96 ( .A(npu_inst_pe_1_2_5_n51), .ZN(
        npu_inst_pe_1_2_5_n104) );
  AOI22_X1 npu_inst_pe_1_2_5_U95 ( .A1(npu_inst_int_data_y_3__5__1_), .A2(
        npu_inst_pe_1_2_5_n46), .B1(npu_inst_pe_1_2_5_n117), .B2(
        npu_inst_pe_1_2_5_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_2_5_n47) );
  INV_X1 npu_inst_pe_1_2_5_U94 ( .A(npu_inst_pe_1_2_5_n47), .ZN(
        npu_inst_pe_1_2_5_n105) );
  AOI22_X1 npu_inst_pe_1_2_5_U93 ( .A1(npu_inst_int_data_y_3__5__1_), .A2(
        npu_inst_pe_1_2_5_n42), .B1(npu_inst_pe_1_2_5_n119), .B2(
        npu_inst_pe_1_2_5_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_2_5_n43) );
  INV_X1 npu_inst_pe_1_2_5_U92 ( .A(npu_inst_pe_1_2_5_n43), .ZN(
        npu_inst_pe_1_2_5_n106) );
  AOI22_X1 npu_inst_pe_1_2_5_U91 ( .A1(npu_inst_pe_1_2_5_n38), .A2(
        npu_inst_int_data_y_3__5__1_), .B1(npu_inst_pe_1_2_5_n118), .B2(
        npu_inst_pe_1_2_5_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_2_5_n39) );
  INV_X1 npu_inst_pe_1_2_5_U90 ( .A(npu_inst_pe_1_2_5_n39), .ZN(
        npu_inst_pe_1_2_5_n107) );
  AOI22_X1 npu_inst_pe_1_2_5_U89 ( .A1(npu_inst_pe_1_2_5_n38), .A2(
        npu_inst_int_data_y_3__5__0_), .B1(npu_inst_pe_1_2_5_n118), .B2(
        npu_inst_pe_1_2_5_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_2_5_n37) );
  INV_X1 npu_inst_pe_1_2_5_U88 ( .A(npu_inst_pe_1_2_5_n37), .ZN(
        npu_inst_pe_1_2_5_n113) );
  NAND2_X1 npu_inst_pe_1_2_5_U87 ( .A1(npu_inst_pe_1_2_5_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_2_5_n60), .ZN(npu_inst_pe_1_2_5_n74) );
  OAI21_X1 npu_inst_pe_1_2_5_U86 ( .B1(npu_inst_pe_1_2_5_n63), .B2(
        npu_inst_pe_1_2_5_n60), .A(npu_inst_pe_1_2_5_n74), .ZN(
        npu_inst_pe_1_2_5_n97) );
  NAND2_X1 npu_inst_pe_1_2_5_U85 ( .A1(npu_inst_pe_1_2_5_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_2_5_n60), .ZN(npu_inst_pe_1_2_5_n73) );
  OAI21_X1 npu_inst_pe_1_2_5_U84 ( .B1(npu_inst_pe_1_2_5_n61), .B2(
        npu_inst_pe_1_2_5_n60), .A(npu_inst_pe_1_2_5_n73), .ZN(
        npu_inst_pe_1_2_5_n96) );
  NAND2_X1 npu_inst_pe_1_2_5_U83 ( .A1(npu_inst_pe_1_2_5_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_2_5_n56), .ZN(npu_inst_pe_1_2_5_n72) );
  OAI21_X1 npu_inst_pe_1_2_5_U82 ( .B1(npu_inst_pe_1_2_5_n63), .B2(
        npu_inst_pe_1_2_5_n56), .A(npu_inst_pe_1_2_5_n72), .ZN(
        npu_inst_pe_1_2_5_n95) );
  NAND2_X1 npu_inst_pe_1_2_5_U81 ( .A1(npu_inst_pe_1_2_5_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_2_5_n56), .ZN(npu_inst_pe_1_2_5_n71) );
  OAI21_X1 npu_inst_pe_1_2_5_U80 ( .B1(npu_inst_pe_1_2_5_n61), .B2(
        npu_inst_pe_1_2_5_n56), .A(npu_inst_pe_1_2_5_n71), .ZN(
        npu_inst_pe_1_2_5_n94) );
  NAND2_X1 npu_inst_pe_1_2_5_U79 ( .A1(npu_inst_pe_1_2_5_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_2_5_n52), .ZN(npu_inst_pe_1_2_5_n70) );
  OAI21_X1 npu_inst_pe_1_2_5_U78 ( .B1(npu_inst_pe_1_2_5_n63), .B2(
        npu_inst_pe_1_2_5_n52), .A(npu_inst_pe_1_2_5_n70), .ZN(
        npu_inst_pe_1_2_5_n93) );
  NAND2_X1 npu_inst_pe_1_2_5_U77 ( .A1(npu_inst_pe_1_2_5_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_2_5_n52), .ZN(npu_inst_pe_1_2_5_n69) );
  OAI21_X1 npu_inst_pe_1_2_5_U76 ( .B1(npu_inst_pe_1_2_5_n61), .B2(
        npu_inst_pe_1_2_5_n52), .A(npu_inst_pe_1_2_5_n69), .ZN(
        npu_inst_pe_1_2_5_n92) );
  NAND2_X1 npu_inst_pe_1_2_5_U75 ( .A1(npu_inst_pe_1_2_5_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_2_5_n48), .ZN(npu_inst_pe_1_2_5_n68) );
  OAI21_X1 npu_inst_pe_1_2_5_U74 ( .B1(npu_inst_pe_1_2_5_n63), .B2(
        npu_inst_pe_1_2_5_n48), .A(npu_inst_pe_1_2_5_n68), .ZN(
        npu_inst_pe_1_2_5_n91) );
  NAND2_X1 npu_inst_pe_1_2_5_U73 ( .A1(npu_inst_pe_1_2_5_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_2_5_n48), .ZN(npu_inst_pe_1_2_5_n67) );
  OAI21_X1 npu_inst_pe_1_2_5_U72 ( .B1(npu_inst_pe_1_2_5_n61), .B2(
        npu_inst_pe_1_2_5_n48), .A(npu_inst_pe_1_2_5_n67), .ZN(
        npu_inst_pe_1_2_5_n90) );
  NAND2_X1 npu_inst_pe_1_2_5_U71 ( .A1(npu_inst_pe_1_2_5_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_2_5_n44), .ZN(npu_inst_pe_1_2_5_n66) );
  OAI21_X1 npu_inst_pe_1_2_5_U70 ( .B1(npu_inst_pe_1_2_5_n63), .B2(
        npu_inst_pe_1_2_5_n44), .A(npu_inst_pe_1_2_5_n66), .ZN(
        npu_inst_pe_1_2_5_n89) );
  NAND2_X1 npu_inst_pe_1_2_5_U69 ( .A1(npu_inst_pe_1_2_5_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_2_5_n44), .ZN(npu_inst_pe_1_2_5_n65) );
  OAI21_X1 npu_inst_pe_1_2_5_U68 ( .B1(npu_inst_pe_1_2_5_n61), .B2(
        npu_inst_pe_1_2_5_n44), .A(npu_inst_pe_1_2_5_n65), .ZN(
        npu_inst_pe_1_2_5_n88) );
  NAND2_X1 npu_inst_pe_1_2_5_U67 ( .A1(npu_inst_pe_1_2_5_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_2_5_n40), .ZN(npu_inst_pe_1_2_5_n64) );
  OAI21_X1 npu_inst_pe_1_2_5_U66 ( .B1(npu_inst_pe_1_2_5_n63), .B2(
        npu_inst_pe_1_2_5_n40), .A(npu_inst_pe_1_2_5_n64), .ZN(
        npu_inst_pe_1_2_5_n87) );
  NAND2_X1 npu_inst_pe_1_2_5_U65 ( .A1(npu_inst_pe_1_2_5_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_2_5_n40), .ZN(npu_inst_pe_1_2_5_n62) );
  OAI21_X1 npu_inst_pe_1_2_5_U64 ( .B1(npu_inst_pe_1_2_5_n61), .B2(
        npu_inst_pe_1_2_5_n40), .A(npu_inst_pe_1_2_5_n62), .ZN(
        npu_inst_pe_1_2_5_n86) );
  AND2_X1 npu_inst_pe_1_2_5_U63 ( .A1(npu_inst_pe_1_2_5_N93), .A2(npu_inst_n58), .ZN(npu_inst_int_data_y_2__5__0_) );
  AND2_X1 npu_inst_pe_1_2_5_U62 ( .A1(npu_inst_n58), .A2(npu_inst_pe_1_2_5_N94), .ZN(npu_inst_int_data_y_2__5__1_) );
  NOR3_X1 npu_inst_pe_1_2_5_U61 ( .A1(npu_inst_pe_1_2_5_n26), .A2(npu_inst_n58), .A3(npu_inst_int_ckg[42]), .ZN(npu_inst_pe_1_2_5_n85) );
  OR2_X1 npu_inst_pe_1_2_5_U60 ( .A1(npu_inst_pe_1_2_5_n85), .A2(
        npu_inst_pe_1_2_5_n2), .ZN(npu_inst_pe_1_2_5_N84) );
  AND2_X1 npu_inst_pe_1_2_5_U59 ( .A1(npu_inst_pe_1_2_5_int_q_acc_0_), .A2(
        npu_inst_pe_1_2_5_n1), .ZN(npu_inst_int_data_res_2__5__0_) );
  AND2_X1 npu_inst_pe_1_2_5_U58 ( .A1(npu_inst_pe_1_2_5_n2), .A2(
        npu_inst_pe_1_2_5_int_q_acc_7_), .ZN(npu_inst_int_data_res_2__5__7_)
         );
  AND2_X1 npu_inst_pe_1_2_5_U57 ( .A1(npu_inst_pe_1_2_5_int_q_acc_1_), .A2(
        npu_inst_pe_1_2_5_n1), .ZN(npu_inst_int_data_res_2__5__1_) );
  AND2_X1 npu_inst_pe_1_2_5_U56 ( .A1(npu_inst_pe_1_2_5_int_q_acc_2_), .A2(
        npu_inst_pe_1_2_5_n1), .ZN(npu_inst_int_data_res_2__5__2_) );
  AND2_X1 npu_inst_pe_1_2_5_U55 ( .A1(npu_inst_pe_1_2_5_int_q_acc_3_), .A2(
        npu_inst_pe_1_2_5_n2), .ZN(npu_inst_int_data_res_2__5__3_) );
  AND2_X1 npu_inst_pe_1_2_5_U54 ( .A1(npu_inst_pe_1_2_5_int_q_acc_4_), .A2(
        npu_inst_pe_1_2_5_n2), .ZN(npu_inst_int_data_res_2__5__4_) );
  AND2_X1 npu_inst_pe_1_2_5_U53 ( .A1(npu_inst_pe_1_2_5_int_q_acc_5_), .A2(
        npu_inst_pe_1_2_5_n2), .ZN(npu_inst_int_data_res_2__5__5_) );
  AND2_X1 npu_inst_pe_1_2_5_U52 ( .A1(npu_inst_pe_1_2_5_int_q_acc_6_), .A2(
        npu_inst_pe_1_2_5_n2), .ZN(npu_inst_int_data_res_2__5__6_) );
  AOI222_X1 npu_inst_pe_1_2_5_U51 ( .A1(npu_inst_int_data_res_3__5__0_), .A2(
        npu_inst_pe_1_2_5_n1), .B1(npu_inst_pe_1_2_5_N73), .B2(
        npu_inst_pe_1_2_5_n76), .C1(npu_inst_pe_1_2_5_N65), .C2(
        npu_inst_pe_1_2_5_n77), .ZN(npu_inst_pe_1_2_5_n84) );
  INV_X1 npu_inst_pe_1_2_5_U50 ( .A(npu_inst_pe_1_2_5_n84), .ZN(
        npu_inst_pe_1_2_5_n101) );
  AOI222_X1 npu_inst_pe_1_2_5_U49 ( .A1(npu_inst_int_data_res_3__5__7_), .A2(
        npu_inst_pe_1_2_5_n1), .B1(npu_inst_pe_1_2_5_N80), .B2(
        npu_inst_pe_1_2_5_n76), .C1(npu_inst_pe_1_2_5_N72), .C2(
        npu_inst_pe_1_2_5_n77), .ZN(npu_inst_pe_1_2_5_n75) );
  INV_X1 npu_inst_pe_1_2_5_U48 ( .A(npu_inst_pe_1_2_5_n75), .ZN(
        npu_inst_pe_1_2_5_n33) );
  AOI222_X1 npu_inst_pe_1_2_5_U47 ( .A1(npu_inst_int_data_res_3__5__1_), .A2(
        npu_inst_pe_1_2_5_n1), .B1(npu_inst_pe_1_2_5_N74), .B2(
        npu_inst_pe_1_2_5_n76), .C1(npu_inst_pe_1_2_5_N66), .C2(
        npu_inst_pe_1_2_5_n77), .ZN(npu_inst_pe_1_2_5_n83) );
  INV_X1 npu_inst_pe_1_2_5_U46 ( .A(npu_inst_pe_1_2_5_n83), .ZN(
        npu_inst_pe_1_2_5_n100) );
  AOI222_X1 npu_inst_pe_1_2_5_U45 ( .A1(npu_inst_int_data_res_3__5__2_), .A2(
        npu_inst_pe_1_2_5_n1), .B1(npu_inst_pe_1_2_5_N75), .B2(
        npu_inst_pe_1_2_5_n76), .C1(npu_inst_pe_1_2_5_N67), .C2(
        npu_inst_pe_1_2_5_n77), .ZN(npu_inst_pe_1_2_5_n82) );
  INV_X1 npu_inst_pe_1_2_5_U44 ( .A(npu_inst_pe_1_2_5_n82), .ZN(
        npu_inst_pe_1_2_5_n99) );
  AOI222_X1 npu_inst_pe_1_2_5_U43 ( .A1(npu_inst_int_data_res_3__5__3_), .A2(
        npu_inst_pe_1_2_5_n1), .B1(npu_inst_pe_1_2_5_N76), .B2(
        npu_inst_pe_1_2_5_n76), .C1(npu_inst_pe_1_2_5_N68), .C2(
        npu_inst_pe_1_2_5_n77), .ZN(npu_inst_pe_1_2_5_n81) );
  INV_X1 npu_inst_pe_1_2_5_U42 ( .A(npu_inst_pe_1_2_5_n81), .ZN(
        npu_inst_pe_1_2_5_n98) );
  AOI222_X1 npu_inst_pe_1_2_5_U41 ( .A1(npu_inst_int_data_res_3__5__4_), .A2(
        npu_inst_pe_1_2_5_n1), .B1(npu_inst_pe_1_2_5_N77), .B2(
        npu_inst_pe_1_2_5_n76), .C1(npu_inst_pe_1_2_5_N69), .C2(
        npu_inst_pe_1_2_5_n77), .ZN(npu_inst_pe_1_2_5_n80) );
  INV_X1 npu_inst_pe_1_2_5_U40 ( .A(npu_inst_pe_1_2_5_n80), .ZN(
        npu_inst_pe_1_2_5_n36) );
  AOI222_X1 npu_inst_pe_1_2_5_U39 ( .A1(npu_inst_int_data_res_3__5__5_), .A2(
        npu_inst_pe_1_2_5_n1), .B1(npu_inst_pe_1_2_5_N78), .B2(
        npu_inst_pe_1_2_5_n76), .C1(npu_inst_pe_1_2_5_N70), .C2(
        npu_inst_pe_1_2_5_n77), .ZN(npu_inst_pe_1_2_5_n79) );
  INV_X1 npu_inst_pe_1_2_5_U38 ( .A(npu_inst_pe_1_2_5_n79), .ZN(
        npu_inst_pe_1_2_5_n35) );
  AOI222_X1 npu_inst_pe_1_2_5_U37 ( .A1(npu_inst_int_data_res_3__5__6_), .A2(
        npu_inst_pe_1_2_5_n1), .B1(npu_inst_pe_1_2_5_N79), .B2(
        npu_inst_pe_1_2_5_n76), .C1(npu_inst_pe_1_2_5_N71), .C2(
        npu_inst_pe_1_2_5_n77), .ZN(npu_inst_pe_1_2_5_n78) );
  INV_X1 npu_inst_pe_1_2_5_U36 ( .A(npu_inst_pe_1_2_5_n78), .ZN(
        npu_inst_pe_1_2_5_n34) );
  INV_X1 npu_inst_pe_1_2_5_U35 ( .A(npu_inst_pe_1_2_5_int_data_1_), .ZN(
        npu_inst_pe_1_2_5_n14) );
  AND2_X1 npu_inst_pe_1_2_5_U34 ( .A1(npu_inst_int_data_x_2__5__1_), .A2(
        npu_inst_pe_1_2_5_int_q_weight_1_), .ZN(npu_inst_pe_1_2_5_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_2_5_U33 ( .A1(npu_inst_int_data_x_2__5__0_), .A2(
        npu_inst_pe_1_2_5_int_q_weight_1_), .ZN(npu_inst_pe_1_2_5_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_2_5_U32 ( .A1(npu_inst_n58), .A2(
        npu_inst_int_data_y_3__5__1_), .B1(npu_inst_pe_1_2_5_n3), .B2(
        npu_inst_int_data_x_2__6__1_), .ZN(npu_inst_pe_1_2_5_n63) );
  AOI22_X1 npu_inst_pe_1_2_5_U31 ( .A1(npu_inst_n58), .A2(
        npu_inst_int_data_y_3__5__0_), .B1(npu_inst_pe_1_2_5_n3), .B2(
        npu_inst_int_data_x_2__6__0_), .ZN(npu_inst_pe_1_2_5_n61) );
  INV_X1 npu_inst_pe_1_2_5_U30 ( .A(npu_inst_pe_1_2_5_int_data_0_), .ZN(
        npu_inst_pe_1_2_5_n13) );
  INV_X1 npu_inst_pe_1_2_5_U29 ( .A(npu_inst_n70), .ZN(npu_inst_pe_1_2_5_n5)
         );
  OR3_X1 npu_inst_pe_1_2_5_U28 ( .A1(npu_inst_pe_1_2_5_n6), .A2(
        npu_inst_pe_1_2_5_n8), .A3(npu_inst_pe_1_2_5_n5), .ZN(
        npu_inst_pe_1_2_5_n56) );
  OR3_X1 npu_inst_pe_1_2_5_U27 ( .A1(npu_inst_pe_1_2_5_n5), .A2(
        npu_inst_pe_1_2_5_n8), .A3(npu_inst_pe_1_2_5_n7), .ZN(
        npu_inst_pe_1_2_5_n48) );
  INV_X1 npu_inst_pe_1_2_5_U26 ( .A(npu_inst_pe_1_2_5_n5), .ZN(
        npu_inst_pe_1_2_5_n4) );
  INV_X1 npu_inst_pe_1_2_5_U25 ( .A(npu_inst_n125), .ZN(npu_inst_pe_1_2_5_n12)
         );
  OR3_X1 npu_inst_pe_1_2_5_U24 ( .A1(npu_inst_pe_1_2_5_n4), .A2(
        npu_inst_pe_1_2_5_n8), .A3(npu_inst_pe_1_2_5_n7), .ZN(
        npu_inst_pe_1_2_5_n52) );
  OR3_X1 npu_inst_pe_1_2_5_U23 ( .A1(npu_inst_pe_1_2_5_n6), .A2(
        npu_inst_pe_1_2_5_n8), .A3(npu_inst_pe_1_2_5_n4), .ZN(
        npu_inst_pe_1_2_5_n60) );
  NOR2_X1 npu_inst_pe_1_2_5_U22 ( .A1(npu_inst_pe_1_2_5_n60), .A2(
        npu_inst_pe_1_2_5_n3), .ZN(npu_inst_pe_1_2_5_n58) );
  NOR2_X1 npu_inst_pe_1_2_5_U21 ( .A1(npu_inst_pe_1_2_5_n56), .A2(
        npu_inst_pe_1_2_5_n3), .ZN(npu_inst_pe_1_2_5_n54) );
  NOR2_X1 npu_inst_pe_1_2_5_U20 ( .A1(npu_inst_pe_1_2_5_n52), .A2(
        npu_inst_pe_1_2_5_n3), .ZN(npu_inst_pe_1_2_5_n50) );
  NOR2_X1 npu_inst_pe_1_2_5_U19 ( .A1(npu_inst_pe_1_2_5_n48), .A2(
        npu_inst_pe_1_2_5_n3), .ZN(npu_inst_pe_1_2_5_n46) );
  NOR2_X1 npu_inst_pe_1_2_5_U18 ( .A1(npu_inst_pe_1_2_5_n40), .A2(
        npu_inst_pe_1_2_5_n3), .ZN(npu_inst_pe_1_2_5_n38) );
  NOR2_X1 npu_inst_pe_1_2_5_U17 ( .A1(npu_inst_pe_1_2_5_n44), .A2(
        npu_inst_pe_1_2_5_n3), .ZN(npu_inst_pe_1_2_5_n42) );
  BUF_X1 npu_inst_pe_1_2_5_U16 ( .A(npu_inst_n102), .Z(npu_inst_pe_1_2_5_n8)
         );
  BUF_X1 npu_inst_pe_1_2_5_U15 ( .A(npu_inst_pe_1_2_5_n12), .Z(
        npu_inst_pe_1_2_5_n11) );
  BUF_X1 npu_inst_pe_1_2_5_U14 ( .A(npu_inst_pe_1_2_5_n12), .Z(
        npu_inst_pe_1_2_5_n10) );
  BUF_X1 npu_inst_pe_1_2_5_U13 ( .A(npu_inst_pe_1_2_5_n12), .Z(
        npu_inst_pe_1_2_5_n9) );
  INV_X1 npu_inst_pe_1_2_5_U12 ( .A(npu_inst_pe_1_2_5_n38), .ZN(
        npu_inst_pe_1_2_5_n118) );
  INV_X1 npu_inst_pe_1_2_5_U11 ( .A(npu_inst_pe_1_2_5_n58), .ZN(
        npu_inst_pe_1_2_5_n114) );
  INV_X1 npu_inst_pe_1_2_5_U10 ( .A(npu_inst_pe_1_2_5_n54), .ZN(
        npu_inst_pe_1_2_5_n115) );
  INV_X1 npu_inst_pe_1_2_5_U9 ( .A(npu_inst_pe_1_2_5_n50), .ZN(
        npu_inst_pe_1_2_5_n116) );
  INV_X1 npu_inst_pe_1_2_5_U8 ( .A(npu_inst_pe_1_2_5_n46), .ZN(
        npu_inst_pe_1_2_5_n117) );
  INV_X1 npu_inst_pe_1_2_5_U7 ( .A(npu_inst_pe_1_2_5_n42), .ZN(
        npu_inst_pe_1_2_5_n119) );
  BUF_X1 npu_inst_pe_1_2_5_U6 ( .A(npu_inst_n28), .Z(npu_inst_pe_1_2_5_n2) );
  BUF_X1 npu_inst_pe_1_2_5_U5 ( .A(npu_inst_n28), .Z(npu_inst_pe_1_2_5_n1) );
  NOR2_X1 npu_inst_pe_1_2_5_U4 ( .A1(npu_inst_pe_1_2_5_int_q_weight_0_), .A2(
        npu_inst_pe_1_2_5_n1), .ZN(npu_inst_pe_1_2_5_n76) );
  NOR2_X1 npu_inst_pe_1_2_5_U3 ( .A1(npu_inst_pe_1_2_5_n27), .A2(
        npu_inst_pe_1_2_5_n1), .ZN(npu_inst_pe_1_2_5_n77) );
  FA_X1 npu_inst_pe_1_2_5_sub_77_U2_1 ( .A(npu_inst_pe_1_2_5_int_q_acc_1_), 
        .B(npu_inst_pe_1_2_5_n14), .CI(npu_inst_pe_1_2_5_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_2_5_sub_77_carry_2_), .S(npu_inst_pe_1_2_5_N66) );
  FA_X1 npu_inst_pe_1_2_5_add_79_U1_1 ( .A(npu_inst_pe_1_2_5_int_q_acc_1_), 
        .B(npu_inst_pe_1_2_5_int_data_1_), .CI(
        npu_inst_pe_1_2_5_add_79_carry_1_), .CO(
        npu_inst_pe_1_2_5_add_79_carry_2_), .S(npu_inst_pe_1_2_5_N74) );
  NAND3_X1 npu_inst_pe_1_2_5_U109 ( .A1(npu_inst_pe_1_2_5_n5), .A2(
        npu_inst_pe_1_2_5_n7), .A3(npu_inst_pe_1_2_5_n8), .ZN(
        npu_inst_pe_1_2_5_n44) );
  NAND3_X1 npu_inst_pe_1_2_5_U108 ( .A1(npu_inst_pe_1_2_5_n4), .A2(
        npu_inst_pe_1_2_5_n7), .A3(npu_inst_pe_1_2_5_n8), .ZN(
        npu_inst_pe_1_2_5_n40) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_2_5_n34), .CK(
        npu_inst_pe_1_2_5_net3810), .RN(npu_inst_pe_1_2_5_n9), .Q(
        npu_inst_pe_1_2_5_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_2_5_n35), .CK(
        npu_inst_pe_1_2_5_net3810), .RN(npu_inst_pe_1_2_5_n9), .Q(
        npu_inst_pe_1_2_5_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_2_5_n36), .CK(
        npu_inst_pe_1_2_5_net3810), .RN(npu_inst_pe_1_2_5_n9), .Q(
        npu_inst_pe_1_2_5_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_2_5_n98), .CK(
        npu_inst_pe_1_2_5_net3810), .RN(npu_inst_pe_1_2_5_n9), .Q(
        npu_inst_pe_1_2_5_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_2_5_n99), .CK(
        npu_inst_pe_1_2_5_net3810), .RN(npu_inst_pe_1_2_5_n9), .Q(
        npu_inst_pe_1_2_5_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_2_5_n100), 
        .CK(npu_inst_pe_1_2_5_net3810), .RN(npu_inst_pe_1_2_5_n9), .Q(
        npu_inst_pe_1_2_5_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_2_5_n33), .CK(
        npu_inst_pe_1_2_5_net3810), .RN(npu_inst_pe_1_2_5_n9), .Q(
        npu_inst_pe_1_2_5_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_2_5_n101), 
        .CK(npu_inst_pe_1_2_5_net3810), .RN(npu_inst_pe_1_2_5_n9), .Q(
        npu_inst_pe_1_2_5_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_weight_reg_0_ ( .D(npu_inst_n111), .CK(
        npu_inst_pe_1_2_5_net3816), .RN(npu_inst_pe_1_2_5_n9), .Q(
        npu_inst_pe_1_2_5_int_q_weight_0_), .QN(npu_inst_pe_1_2_5_n27) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_weight_reg_1_ ( .D(npu_inst_n117), .CK(
        npu_inst_pe_1_2_5_net3816), .RN(npu_inst_pe_1_2_5_n9), .Q(
        npu_inst_pe_1_2_5_int_q_weight_1_), .QN(npu_inst_pe_1_2_5_n26) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_2_5_n113), 
        .CK(npu_inst_pe_1_2_5_net3816), .RN(npu_inst_pe_1_2_5_n9), .Q(
        npu_inst_pe_1_2_5_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_2_5_n107), 
        .CK(npu_inst_pe_1_2_5_net3816), .RN(npu_inst_pe_1_2_5_n9), .Q(
        npu_inst_pe_1_2_5_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_2_5_n112), 
        .CK(npu_inst_pe_1_2_5_net3816), .RN(npu_inst_pe_1_2_5_n10), .Q(
        npu_inst_pe_1_2_5_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_2_5_n106), 
        .CK(npu_inst_pe_1_2_5_net3816), .RN(npu_inst_pe_1_2_5_n10), .Q(
        npu_inst_pe_1_2_5_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_2_5_n111), 
        .CK(npu_inst_pe_1_2_5_net3816), .RN(npu_inst_pe_1_2_5_n10), .Q(
        npu_inst_pe_1_2_5_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_2_5_n105), 
        .CK(npu_inst_pe_1_2_5_net3816), .RN(npu_inst_pe_1_2_5_n10), .Q(
        npu_inst_pe_1_2_5_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_2_5_n110), 
        .CK(npu_inst_pe_1_2_5_net3816), .RN(npu_inst_pe_1_2_5_n10), .Q(
        npu_inst_pe_1_2_5_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_2_5_n104), 
        .CK(npu_inst_pe_1_2_5_net3816), .RN(npu_inst_pe_1_2_5_n10), .Q(
        npu_inst_pe_1_2_5_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_2_5_n109), 
        .CK(npu_inst_pe_1_2_5_net3816), .RN(npu_inst_pe_1_2_5_n10), .Q(
        npu_inst_pe_1_2_5_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_2_5_n103), 
        .CK(npu_inst_pe_1_2_5_net3816), .RN(npu_inst_pe_1_2_5_n10), .Q(
        npu_inst_pe_1_2_5_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_2_5_n108), 
        .CK(npu_inst_pe_1_2_5_net3816), .RN(npu_inst_pe_1_2_5_n10), .Q(
        npu_inst_pe_1_2_5_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_2_5_n102), 
        .CK(npu_inst_pe_1_2_5_net3816), .RN(npu_inst_pe_1_2_5_n10), .Q(
        npu_inst_pe_1_2_5_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_2_5_n86), 
        .CK(npu_inst_pe_1_2_5_net3816), .RN(npu_inst_pe_1_2_5_n10), .Q(
        npu_inst_pe_1_2_5_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_2_5_n87), 
        .CK(npu_inst_pe_1_2_5_net3816), .RN(npu_inst_pe_1_2_5_n10), .Q(
        npu_inst_pe_1_2_5_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_2_5_n88), 
        .CK(npu_inst_pe_1_2_5_net3816), .RN(npu_inst_pe_1_2_5_n11), .Q(
        npu_inst_pe_1_2_5_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_2_5_n89), 
        .CK(npu_inst_pe_1_2_5_net3816), .RN(npu_inst_pe_1_2_5_n11), .Q(
        npu_inst_pe_1_2_5_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_2_5_n90), 
        .CK(npu_inst_pe_1_2_5_net3816), .RN(npu_inst_pe_1_2_5_n11), .Q(
        npu_inst_pe_1_2_5_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_2_5_n91), 
        .CK(npu_inst_pe_1_2_5_net3816), .RN(npu_inst_pe_1_2_5_n11), .Q(
        npu_inst_pe_1_2_5_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_2_5_n92), 
        .CK(npu_inst_pe_1_2_5_net3816), .RN(npu_inst_pe_1_2_5_n11), .Q(
        npu_inst_pe_1_2_5_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_2_5_n93), 
        .CK(npu_inst_pe_1_2_5_net3816), .RN(npu_inst_pe_1_2_5_n11), .Q(
        npu_inst_pe_1_2_5_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_2_5_n94), 
        .CK(npu_inst_pe_1_2_5_net3816), .RN(npu_inst_pe_1_2_5_n11), .Q(
        npu_inst_pe_1_2_5_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_2_5_n95), 
        .CK(npu_inst_pe_1_2_5_net3816), .RN(npu_inst_pe_1_2_5_n11), .Q(
        npu_inst_pe_1_2_5_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_2_5_n96), 
        .CK(npu_inst_pe_1_2_5_net3816), .RN(npu_inst_pe_1_2_5_n11), .Q(
        npu_inst_pe_1_2_5_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_2_5_n97), 
        .CK(npu_inst_pe_1_2_5_net3816), .RN(npu_inst_pe_1_2_5_n11), .Q(
        npu_inst_pe_1_2_5_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_2_5_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_2_5_N84), .SE(1'b0), .GCK(npu_inst_pe_1_2_5_net3810) );
  CLKGATETST_X1 npu_inst_pe_1_2_5_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n64), .SE(1'b0), .GCK(npu_inst_pe_1_2_5_net3816) );
  MUX2_X1 npu_inst_pe_1_2_6_U162 ( .A(npu_inst_pe_1_2_6_n32), .B(
        npu_inst_pe_1_2_6_n29), .S(npu_inst_pe_1_2_6_n8), .Z(
        npu_inst_pe_1_2_6_N93) );
  MUX2_X1 npu_inst_pe_1_2_6_U161 ( .A(npu_inst_pe_1_2_6_n31), .B(
        npu_inst_pe_1_2_6_n30), .S(npu_inst_pe_1_2_6_n6), .Z(
        npu_inst_pe_1_2_6_n32) );
  MUX2_X1 npu_inst_pe_1_2_6_U160 ( .A(npu_inst_pe_1_2_6_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_2_6_int_q_reg_v_1__0_), .S(npu_inst_pe_1_2_6_n4), .Z(
        npu_inst_pe_1_2_6_n31) );
  MUX2_X1 npu_inst_pe_1_2_6_U159 ( .A(npu_inst_pe_1_2_6_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_2_6_int_q_reg_v_3__0_), .S(npu_inst_pe_1_2_6_n4), .Z(
        npu_inst_pe_1_2_6_n30) );
  MUX2_X1 npu_inst_pe_1_2_6_U158 ( .A(npu_inst_pe_1_2_6_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_2_6_int_q_reg_v_5__0_), .S(npu_inst_pe_1_2_6_n4), .Z(
        npu_inst_pe_1_2_6_n29) );
  MUX2_X1 npu_inst_pe_1_2_6_U157 ( .A(npu_inst_pe_1_2_6_n28), .B(
        npu_inst_pe_1_2_6_n23), .S(npu_inst_pe_1_2_6_n8), .Z(
        npu_inst_pe_1_2_6_N94) );
  MUX2_X1 npu_inst_pe_1_2_6_U156 ( .A(npu_inst_pe_1_2_6_n25), .B(
        npu_inst_pe_1_2_6_n24), .S(npu_inst_pe_1_2_6_n6), .Z(
        npu_inst_pe_1_2_6_n28) );
  MUX2_X1 npu_inst_pe_1_2_6_U155 ( .A(npu_inst_pe_1_2_6_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_2_6_int_q_reg_v_1__1_), .S(npu_inst_pe_1_2_6_n4), .Z(
        npu_inst_pe_1_2_6_n25) );
  MUX2_X1 npu_inst_pe_1_2_6_U154 ( .A(npu_inst_pe_1_2_6_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_2_6_int_q_reg_v_3__1_), .S(npu_inst_pe_1_2_6_n4), .Z(
        npu_inst_pe_1_2_6_n24) );
  MUX2_X1 npu_inst_pe_1_2_6_U153 ( .A(npu_inst_pe_1_2_6_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_2_6_int_q_reg_v_5__1_), .S(npu_inst_pe_1_2_6_n4), .Z(
        npu_inst_pe_1_2_6_n23) );
  MUX2_X1 npu_inst_pe_1_2_6_U152 ( .A(npu_inst_pe_1_2_6_n22), .B(
        npu_inst_pe_1_2_6_n19), .S(npu_inst_pe_1_2_6_n8), .Z(
        npu_inst_int_data_x_2__6__1_) );
  MUX2_X1 npu_inst_pe_1_2_6_U151 ( .A(npu_inst_pe_1_2_6_n21), .B(
        npu_inst_pe_1_2_6_n20), .S(npu_inst_pe_1_2_6_n6), .Z(
        npu_inst_pe_1_2_6_n22) );
  MUX2_X1 npu_inst_pe_1_2_6_U150 ( .A(npu_inst_pe_1_2_6_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_2_6_int_q_reg_h_1__1_), .S(npu_inst_pe_1_2_6_n4), .Z(
        npu_inst_pe_1_2_6_n21) );
  MUX2_X1 npu_inst_pe_1_2_6_U149 ( .A(npu_inst_pe_1_2_6_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_2_6_int_q_reg_h_3__1_), .S(npu_inst_pe_1_2_6_n4), .Z(
        npu_inst_pe_1_2_6_n20) );
  MUX2_X1 npu_inst_pe_1_2_6_U148 ( .A(npu_inst_pe_1_2_6_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_2_6_int_q_reg_h_5__1_), .S(npu_inst_pe_1_2_6_n4), .Z(
        npu_inst_pe_1_2_6_n19) );
  MUX2_X1 npu_inst_pe_1_2_6_U147 ( .A(npu_inst_pe_1_2_6_n18), .B(
        npu_inst_pe_1_2_6_n15), .S(npu_inst_pe_1_2_6_n8), .Z(
        npu_inst_int_data_x_2__6__0_) );
  MUX2_X1 npu_inst_pe_1_2_6_U146 ( .A(npu_inst_pe_1_2_6_n17), .B(
        npu_inst_pe_1_2_6_n16), .S(npu_inst_pe_1_2_6_n6), .Z(
        npu_inst_pe_1_2_6_n18) );
  MUX2_X1 npu_inst_pe_1_2_6_U145 ( .A(npu_inst_pe_1_2_6_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_2_6_int_q_reg_h_1__0_), .S(npu_inst_pe_1_2_6_n4), .Z(
        npu_inst_pe_1_2_6_n17) );
  MUX2_X1 npu_inst_pe_1_2_6_U144 ( .A(npu_inst_pe_1_2_6_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_2_6_int_q_reg_h_3__0_), .S(npu_inst_pe_1_2_6_n4), .Z(
        npu_inst_pe_1_2_6_n16) );
  MUX2_X1 npu_inst_pe_1_2_6_U143 ( .A(npu_inst_pe_1_2_6_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_2_6_int_q_reg_h_5__0_), .S(npu_inst_pe_1_2_6_n4), .Z(
        npu_inst_pe_1_2_6_n15) );
  XOR2_X1 npu_inst_pe_1_2_6_U142 ( .A(npu_inst_pe_1_2_6_int_data_0_), .B(
        npu_inst_pe_1_2_6_int_q_acc_0_), .Z(npu_inst_pe_1_2_6_N73) );
  AND2_X1 npu_inst_pe_1_2_6_U141 ( .A1(npu_inst_pe_1_2_6_int_q_acc_0_), .A2(
        npu_inst_pe_1_2_6_int_data_0_), .ZN(npu_inst_pe_1_2_6_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_2_6_U140 ( .A(npu_inst_pe_1_2_6_int_q_acc_0_), .B(
        npu_inst_pe_1_2_6_n13), .ZN(npu_inst_pe_1_2_6_N65) );
  OR2_X1 npu_inst_pe_1_2_6_U139 ( .A1(npu_inst_pe_1_2_6_n13), .A2(
        npu_inst_pe_1_2_6_int_q_acc_0_), .ZN(npu_inst_pe_1_2_6_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_2_6_U138 ( .A(npu_inst_pe_1_2_6_int_q_acc_2_), .B(
        npu_inst_pe_1_2_6_add_79_carry_2_), .Z(npu_inst_pe_1_2_6_N75) );
  AND2_X1 npu_inst_pe_1_2_6_U137 ( .A1(npu_inst_pe_1_2_6_add_79_carry_2_), 
        .A2(npu_inst_pe_1_2_6_int_q_acc_2_), .ZN(
        npu_inst_pe_1_2_6_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_2_6_U136 ( .A(npu_inst_pe_1_2_6_int_q_acc_3_), .B(
        npu_inst_pe_1_2_6_add_79_carry_3_), .Z(npu_inst_pe_1_2_6_N76) );
  AND2_X1 npu_inst_pe_1_2_6_U135 ( .A1(npu_inst_pe_1_2_6_add_79_carry_3_), 
        .A2(npu_inst_pe_1_2_6_int_q_acc_3_), .ZN(
        npu_inst_pe_1_2_6_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_2_6_U134 ( .A(npu_inst_pe_1_2_6_int_q_acc_4_), .B(
        npu_inst_pe_1_2_6_add_79_carry_4_), .Z(npu_inst_pe_1_2_6_N77) );
  AND2_X1 npu_inst_pe_1_2_6_U133 ( .A1(npu_inst_pe_1_2_6_add_79_carry_4_), 
        .A2(npu_inst_pe_1_2_6_int_q_acc_4_), .ZN(
        npu_inst_pe_1_2_6_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_2_6_U132 ( .A(npu_inst_pe_1_2_6_int_q_acc_5_), .B(
        npu_inst_pe_1_2_6_add_79_carry_5_), .Z(npu_inst_pe_1_2_6_N78) );
  AND2_X1 npu_inst_pe_1_2_6_U131 ( .A1(npu_inst_pe_1_2_6_add_79_carry_5_), 
        .A2(npu_inst_pe_1_2_6_int_q_acc_5_), .ZN(
        npu_inst_pe_1_2_6_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_2_6_U130 ( .A(npu_inst_pe_1_2_6_int_q_acc_6_), .B(
        npu_inst_pe_1_2_6_add_79_carry_6_), .Z(npu_inst_pe_1_2_6_N79) );
  AND2_X1 npu_inst_pe_1_2_6_U129 ( .A1(npu_inst_pe_1_2_6_add_79_carry_6_), 
        .A2(npu_inst_pe_1_2_6_int_q_acc_6_), .ZN(
        npu_inst_pe_1_2_6_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_2_6_U128 ( .A(npu_inst_pe_1_2_6_int_q_acc_7_), .B(
        npu_inst_pe_1_2_6_add_79_carry_7_), .Z(npu_inst_pe_1_2_6_N80) );
  XNOR2_X1 npu_inst_pe_1_2_6_U127 ( .A(npu_inst_pe_1_2_6_sub_77_carry_2_), .B(
        npu_inst_pe_1_2_6_int_q_acc_2_), .ZN(npu_inst_pe_1_2_6_N67) );
  OR2_X1 npu_inst_pe_1_2_6_U126 ( .A1(npu_inst_pe_1_2_6_int_q_acc_2_), .A2(
        npu_inst_pe_1_2_6_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_2_6_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_2_6_U125 ( .A(npu_inst_pe_1_2_6_sub_77_carry_3_), .B(
        npu_inst_pe_1_2_6_int_q_acc_3_), .ZN(npu_inst_pe_1_2_6_N68) );
  OR2_X1 npu_inst_pe_1_2_6_U124 ( .A1(npu_inst_pe_1_2_6_int_q_acc_3_), .A2(
        npu_inst_pe_1_2_6_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_2_6_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_2_6_U123 ( .A(npu_inst_pe_1_2_6_sub_77_carry_4_), .B(
        npu_inst_pe_1_2_6_int_q_acc_4_), .ZN(npu_inst_pe_1_2_6_N69) );
  OR2_X1 npu_inst_pe_1_2_6_U122 ( .A1(npu_inst_pe_1_2_6_int_q_acc_4_), .A2(
        npu_inst_pe_1_2_6_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_2_6_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_2_6_U121 ( .A(npu_inst_pe_1_2_6_sub_77_carry_5_), .B(
        npu_inst_pe_1_2_6_int_q_acc_5_), .ZN(npu_inst_pe_1_2_6_N70) );
  OR2_X1 npu_inst_pe_1_2_6_U120 ( .A1(npu_inst_pe_1_2_6_int_q_acc_5_), .A2(
        npu_inst_pe_1_2_6_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_2_6_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_2_6_U119 ( .A(npu_inst_pe_1_2_6_sub_77_carry_6_), .B(
        npu_inst_pe_1_2_6_int_q_acc_6_), .ZN(npu_inst_pe_1_2_6_N71) );
  OR2_X1 npu_inst_pe_1_2_6_U118 ( .A1(npu_inst_pe_1_2_6_int_q_acc_6_), .A2(
        npu_inst_pe_1_2_6_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_2_6_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_2_6_U117 ( .A(npu_inst_pe_1_2_6_int_q_acc_7_), .B(
        npu_inst_pe_1_2_6_sub_77_carry_7_), .ZN(npu_inst_pe_1_2_6_N72) );
  INV_X1 npu_inst_pe_1_2_6_U116 ( .A(npu_inst_n78), .ZN(npu_inst_pe_1_2_6_n7)
         );
  INV_X1 npu_inst_pe_1_2_6_U115 ( .A(npu_inst_pe_1_2_6_n7), .ZN(
        npu_inst_pe_1_2_6_n6) );
  INV_X1 npu_inst_pe_1_2_6_U114 ( .A(npu_inst_n57), .ZN(npu_inst_pe_1_2_6_n3)
         );
  AOI22_X1 npu_inst_pe_1_2_6_U113 ( .A1(npu_inst_int_data_y_3__6__0_), .A2(
        npu_inst_pe_1_2_6_n58), .B1(npu_inst_pe_1_2_6_n114), .B2(
        npu_inst_pe_1_2_6_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_2_6_n57) );
  INV_X1 npu_inst_pe_1_2_6_U112 ( .A(npu_inst_pe_1_2_6_n57), .ZN(
        npu_inst_pe_1_2_6_n108) );
  AOI22_X1 npu_inst_pe_1_2_6_U111 ( .A1(npu_inst_int_data_y_3__6__0_), .A2(
        npu_inst_pe_1_2_6_n54), .B1(npu_inst_pe_1_2_6_n115), .B2(
        npu_inst_pe_1_2_6_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_2_6_n53) );
  INV_X1 npu_inst_pe_1_2_6_U110 ( .A(npu_inst_pe_1_2_6_n53), .ZN(
        npu_inst_pe_1_2_6_n109) );
  AOI22_X1 npu_inst_pe_1_2_6_U107 ( .A1(npu_inst_int_data_y_3__6__0_), .A2(
        npu_inst_pe_1_2_6_n50), .B1(npu_inst_pe_1_2_6_n116), .B2(
        npu_inst_pe_1_2_6_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_2_6_n49) );
  INV_X1 npu_inst_pe_1_2_6_U106 ( .A(npu_inst_pe_1_2_6_n49), .ZN(
        npu_inst_pe_1_2_6_n110) );
  AOI22_X1 npu_inst_pe_1_2_6_U105 ( .A1(npu_inst_int_data_y_3__6__0_), .A2(
        npu_inst_pe_1_2_6_n46), .B1(npu_inst_pe_1_2_6_n117), .B2(
        npu_inst_pe_1_2_6_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_2_6_n45) );
  INV_X1 npu_inst_pe_1_2_6_U104 ( .A(npu_inst_pe_1_2_6_n45), .ZN(
        npu_inst_pe_1_2_6_n111) );
  AOI22_X1 npu_inst_pe_1_2_6_U103 ( .A1(npu_inst_int_data_y_3__6__0_), .A2(
        npu_inst_pe_1_2_6_n42), .B1(npu_inst_pe_1_2_6_n119), .B2(
        npu_inst_pe_1_2_6_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_2_6_n41) );
  INV_X1 npu_inst_pe_1_2_6_U102 ( .A(npu_inst_pe_1_2_6_n41), .ZN(
        npu_inst_pe_1_2_6_n112) );
  AOI22_X1 npu_inst_pe_1_2_6_U101 ( .A1(npu_inst_int_data_y_3__6__1_), .A2(
        npu_inst_pe_1_2_6_n58), .B1(npu_inst_pe_1_2_6_n114), .B2(
        npu_inst_pe_1_2_6_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_2_6_n59) );
  INV_X1 npu_inst_pe_1_2_6_U100 ( .A(npu_inst_pe_1_2_6_n59), .ZN(
        npu_inst_pe_1_2_6_n102) );
  AOI22_X1 npu_inst_pe_1_2_6_U99 ( .A1(npu_inst_int_data_y_3__6__1_), .A2(
        npu_inst_pe_1_2_6_n54), .B1(npu_inst_pe_1_2_6_n115), .B2(
        npu_inst_pe_1_2_6_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_2_6_n55) );
  INV_X1 npu_inst_pe_1_2_6_U98 ( .A(npu_inst_pe_1_2_6_n55), .ZN(
        npu_inst_pe_1_2_6_n103) );
  AOI22_X1 npu_inst_pe_1_2_6_U97 ( .A1(npu_inst_int_data_y_3__6__1_), .A2(
        npu_inst_pe_1_2_6_n50), .B1(npu_inst_pe_1_2_6_n116), .B2(
        npu_inst_pe_1_2_6_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_2_6_n51) );
  INV_X1 npu_inst_pe_1_2_6_U96 ( .A(npu_inst_pe_1_2_6_n51), .ZN(
        npu_inst_pe_1_2_6_n104) );
  AOI22_X1 npu_inst_pe_1_2_6_U95 ( .A1(npu_inst_int_data_y_3__6__1_), .A2(
        npu_inst_pe_1_2_6_n46), .B1(npu_inst_pe_1_2_6_n117), .B2(
        npu_inst_pe_1_2_6_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_2_6_n47) );
  INV_X1 npu_inst_pe_1_2_6_U94 ( .A(npu_inst_pe_1_2_6_n47), .ZN(
        npu_inst_pe_1_2_6_n105) );
  AOI22_X1 npu_inst_pe_1_2_6_U93 ( .A1(npu_inst_int_data_y_3__6__1_), .A2(
        npu_inst_pe_1_2_6_n42), .B1(npu_inst_pe_1_2_6_n119), .B2(
        npu_inst_pe_1_2_6_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_2_6_n43) );
  INV_X1 npu_inst_pe_1_2_6_U92 ( .A(npu_inst_pe_1_2_6_n43), .ZN(
        npu_inst_pe_1_2_6_n106) );
  AOI22_X1 npu_inst_pe_1_2_6_U91 ( .A1(npu_inst_pe_1_2_6_n38), .A2(
        npu_inst_int_data_y_3__6__1_), .B1(npu_inst_pe_1_2_6_n118), .B2(
        npu_inst_pe_1_2_6_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_2_6_n39) );
  INV_X1 npu_inst_pe_1_2_6_U90 ( .A(npu_inst_pe_1_2_6_n39), .ZN(
        npu_inst_pe_1_2_6_n107) );
  AOI22_X1 npu_inst_pe_1_2_6_U89 ( .A1(npu_inst_pe_1_2_6_n38), .A2(
        npu_inst_int_data_y_3__6__0_), .B1(npu_inst_pe_1_2_6_n118), .B2(
        npu_inst_pe_1_2_6_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_2_6_n37) );
  INV_X1 npu_inst_pe_1_2_6_U88 ( .A(npu_inst_pe_1_2_6_n37), .ZN(
        npu_inst_pe_1_2_6_n113) );
  NAND2_X1 npu_inst_pe_1_2_6_U87 ( .A1(npu_inst_pe_1_2_6_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_2_6_n60), .ZN(npu_inst_pe_1_2_6_n74) );
  OAI21_X1 npu_inst_pe_1_2_6_U86 ( .B1(npu_inst_pe_1_2_6_n63), .B2(
        npu_inst_pe_1_2_6_n60), .A(npu_inst_pe_1_2_6_n74), .ZN(
        npu_inst_pe_1_2_6_n97) );
  NAND2_X1 npu_inst_pe_1_2_6_U85 ( .A1(npu_inst_pe_1_2_6_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_2_6_n60), .ZN(npu_inst_pe_1_2_6_n73) );
  OAI21_X1 npu_inst_pe_1_2_6_U84 ( .B1(npu_inst_pe_1_2_6_n61), .B2(
        npu_inst_pe_1_2_6_n60), .A(npu_inst_pe_1_2_6_n73), .ZN(
        npu_inst_pe_1_2_6_n96) );
  NAND2_X1 npu_inst_pe_1_2_6_U83 ( .A1(npu_inst_pe_1_2_6_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_2_6_n56), .ZN(npu_inst_pe_1_2_6_n72) );
  OAI21_X1 npu_inst_pe_1_2_6_U82 ( .B1(npu_inst_pe_1_2_6_n63), .B2(
        npu_inst_pe_1_2_6_n56), .A(npu_inst_pe_1_2_6_n72), .ZN(
        npu_inst_pe_1_2_6_n95) );
  NAND2_X1 npu_inst_pe_1_2_6_U81 ( .A1(npu_inst_pe_1_2_6_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_2_6_n56), .ZN(npu_inst_pe_1_2_6_n71) );
  OAI21_X1 npu_inst_pe_1_2_6_U80 ( .B1(npu_inst_pe_1_2_6_n61), .B2(
        npu_inst_pe_1_2_6_n56), .A(npu_inst_pe_1_2_6_n71), .ZN(
        npu_inst_pe_1_2_6_n94) );
  NAND2_X1 npu_inst_pe_1_2_6_U79 ( .A1(npu_inst_pe_1_2_6_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_2_6_n52), .ZN(npu_inst_pe_1_2_6_n70) );
  OAI21_X1 npu_inst_pe_1_2_6_U78 ( .B1(npu_inst_pe_1_2_6_n63), .B2(
        npu_inst_pe_1_2_6_n52), .A(npu_inst_pe_1_2_6_n70), .ZN(
        npu_inst_pe_1_2_6_n93) );
  NAND2_X1 npu_inst_pe_1_2_6_U77 ( .A1(npu_inst_pe_1_2_6_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_2_6_n52), .ZN(npu_inst_pe_1_2_6_n69) );
  OAI21_X1 npu_inst_pe_1_2_6_U76 ( .B1(npu_inst_pe_1_2_6_n61), .B2(
        npu_inst_pe_1_2_6_n52), .A(npu_inst_pe_1_2_6_n69), .ZN(
        npu_inst_pe_1_2_6_n92) );
  NAND2_X1 npu_inst_pe_1_2_6_U75 ( .A1(npu_inst_pe_1_2_6_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_2_6_n48), .ZN(npu_inst_pe_1_2_6_n68) );
  OAI21_X1 npu_inst_pe_1_2_6_U74 ( .B1(npu_inst_pe_1_2_6_n63), .B2(
        npu_inst_pe_1_2_6_n48), .A(npu_inst_pe_1_2_6_n68), .ZN(
        npu_inst_pe_1_2_6_n91) );
  NAND2_X1 npu_inst_pe_1_2_6_U73 ( .A1(npu_inst_pe_1_2_6_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_2_6_n48), .ZN(npu_inst_pe_1_2_6_n67) );
  OAI21_X1 npu_inst_pe_1_2_6_U72 ( .B1(npu_inst_pe_1_2_6_n61), .B2(
        npu_inst_pe_1_2_6_n48), .A(npu_inst_pe_1_2_6_n67), .ZN(
        npu_inst_pe_1_2_6_n90) );
  NAND2_X1 npu_inst_pe_1_2_6_U71 ( .A1(npu_inst_pe_1_2_6_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_2_6_n44), .ZN(npu_inst_pe_1_2_6_n66) );
  OAI21_X1 npu_inst_pe_1_2_6_U70 ( .B1(npu_inst_pe_1_2_6_n63), .B2(
        npu_inst_pe_1_2_6_n44), .A(npu_inst_pe_1_2_6_n66), .ZN(
        npu_inst_pe_1_2_6_n89) );
  NAND2_X1 npu_inst_pe_1_2_6_U69 ( .A1(npu_inst_pe_1_2_6_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_2_6_n44), .ZN(npu_inst_pe_1_2_6_n65) );
  OAI21_X1 npu_inst_pe_1_2_6_U68 ( .B1(npu_inst_pe_1_2_6_n61), .B2(
        npu_inst_pe_1_2_6_n44), .A(npu_inst_pe_1_2_6_n65), .ZN(
        npu_inst_pe_1_2_6_n88) );
  NAND2_X1 npu_inst_pe_1_2_6_U67 ( .A1(npu_inst_pe_1_2_6_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_2_6_n40), .ZN(npu_inst_pe_1_2_6_n64) );
  OAI21_X1 npu_inst_pe_1_2_6_U66 ( .B1(npu_inst_pe_1_2_6_n63), .B2(
        npu_inst_pe_1_2_6_n40), .A(npu_inst_pe_1_2_6_n64), .ZN(
        npu_inst_pe_1_2_6_n87) );
  NAND2_X1 npu_inst_pe_1_2_6_U65 ( .A1(npu_inst_pe_1_2_6_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_2_6_n40), .ZN(npu_inst_pe_1_2_6_n62) );
  OAI21_X1 npu_inst_pe_1_2_6_U64 ( .B1(npu_inst_pe_1_2_6_n61), .B2(
        npu_inst_pe_1_2_6_n40), .A(npu_inst_pe_1_2_6_n62), .ZN(
        npu_inst_pe_1_2_6_n86) );
  AND2_X1 npu_inst_pe_1_2_6_U63 ( .A1(npu_inst_pe_1_2_6_N93), .A2(npu_inst_n57), .ZN(npu_inst_int_data_y_2__6__0_) );
  AND2_X1 npu_inst_pe_1_2_6_U62 ( .A1(npu_inst_n57), .A2(npu_inst_pe_1_2_6_N94), .ZN(npu_inst_int_data_y_2__6__1_) );
  NOR3_X1 npu_inst_pe_1_2_6_U61 ( .A1(npu_inst_pe_1_2_6_n26), .A2(npu_inst_n57), .A3(npu_inst_int_ckg[41]), .ZN(npu_inst_pe_1_2_6_n85) );
  OR2_X1 npu_inst_pe_1_2_6_U60 ( .A1(npu_inst_pe_1_2_6_n85), .A2(
        npu_inst_pe_1_2_6_n2), .ZN(npu_inst_pe_1_2_6_N84) );
  AND2_X1 npu_inst_pe_1_2_6_U59 ( .A1(npu_inst_pe_1_2_6_int_q_acc_0_), .A2(
        npu_inst_pe_1_2_6_n1), .ZN(npu_inst_int_data_res_2__6__0_) );
  AND2_X1 npu_inst_pe_1_2_6_U58 ( .A1(npu_inst_pe_1_2_6_n2), .A2(
        npu_inst_pe_1_2_6_int_q_acc_7_), .ZN(npu_inst_int_data_res_2__6__7_)
         );
  AND2_X1 npu_inst_pe_1_2_6_U57 ( .A1(npu_inst_pe_1_2_6_int_q_acc_1_), .A2(
        npu_inst_pe_1_2_6_n1), .ZN(npu_inst_int_data_res_2__6__1_) );
  AND2_X1 npu_inst_pe_1_2_6_U56 ( .A1(npu_inst_pe_1_2_6_int_q_acc_2_), .A2(
        npu_inst_pe_1_2_6_n1), .ZN(npu_inst_int_data_res_2__6__2_) );
  AND2_X1 npu_inst_pe_1_2_6_U55 ( .A1(npu_inst_pe_1_2_6_int_q_acc_3_), .A2(
        npu_inst_pe_1_2_6_n2), .ZN(npu_inst_int_data_res_2__6__3_) );
  AND2_X1 npu_inst_pe_1_2_6_U54 ( .A1(npu_inst_pe_1_2_6_int_q_acc_4_), .A2(
        npu_inst_pe_1_2_6_n2), .ZN(npu_inst_int_data_res_2__6__4_) );
  AND2_X1 npu_inst_pe_1_2_6_U53 ( .A1(npu_inst_pe_1_2_6_int_q_acc_5_), .A2(
        npu_inst_pe_1_2_6_n2), .ZN(npu_inst_int_data_res_2__6__5_) );
  AND2_X1 npu_inst_pe_1_2_6_U52 ( .A1(npu_inst_pe_1_2_6_int_q_acc_6_), .A2(
        npu_inst_pe_1_2_6_n2), .ZN(npu_inst_int_data_res_2__6__6_) );
  AOI222_X1 npu_inst_pe_1_2_6_U51 ( .A1(npu_inst_int_data_res_3__6__0_), .A2(
        npu_inst_pe_1_2_6_n1), .B1(npu_inst_pe_1_2_6_N73), .B2(
        npu_inst_pe_1_2_6_n76), .C1(npu_inst_pe_1_2_6_N65), .C2(
        npu_inst_pe_1_2_6_n77), .ZN(npu_inst_pe_1_2_6_n84) );
  INV_X1 npu_inst_pe_1_2_6_U50 ( .A(npu_inst_pe_1_2_6_n84), .ZN(
        npu_inst_pe_1_2_6_n101) );
  AOI222_X1 npu_inst_pe_1_2_6_U49 ( .A1(npu_inst_int_data_res_3__6__7_), .A2(
        npu_inst_pe_1_2_6_n1), .B1(npu_inst_pe_1_2_6_N80), .B2(
        npu_inst_pe_1_2_6_n76), .C1(npu_inst_pe_1_2_6_N72), .C2(
        npu_inst_pe_1_2_6_n77), .ZN(npu_inst_pe_1_2_6_n75) );
  INV_X1 npu_inst_pe_1_2_6_U48 ( .A(npu_inst_pe_1_2_6_n75), .ZN(
        npu_inst_pe_1_2_6_n33) );
  AOI222_X1 npu_inst_pe_1_2_6_U47 ( .A1(npu_inst_int_data_res_3__6__1_), .A2(
        npu_inst_pe_1_2_6_n1), .B1(npu_inst_pe_1_2_6_N74), .B2(
        npu_inst_pe_1_2_6_n76), .C1(npu_inst_pe_1_2_6_N66), .C2(
        npu_inst_pe_1_2_6_n77), .ZN(npu_inst_pe_1_2_6_n83) );
  INV_X1 npu_inst_pe_1_2_6_U46 ( .A(npu_inst_pe_1_2_6_n83), .ZN(
        npu_inst_pe_1_2_6_n100) );
  AOI222_X1 npu_inst_pe_1_2_6_U45 ( .A1(npu_inst_int_data_res_3__6__2_), .A2(
        npu_inst_pe_1_2_6_n1), .B1(npu_inst_pe_1_2_6_N75), .B2(
        npu_inst_pe_1_2_6_n76), .C1(npu_inst_pe_1_2_6_N67), .C2(
        npu_inst_pe_1_2_6_n77), .ZN(npu_inst_pe_1_2_6_n82) );
  INV_X1 npu_inst_pe_1_2_6_U44 ( .A(npu_inst_pe_1_2_6_n82), .ZN(
        npu_inst_pe_1_2_6_n99) );
  AOI222_X1 npu_inst_pe_1_2_6_U43 ( .A1(npu_inst_int_data_res_3__6__3_), .A2(
        npu_inst_pe_1_2_6_n1), .B1(npu_inst_pe_1_2_6_N76), .B2(
        npu_inst_pe_1_2_6_n76), .C1(npu_inst_pe_1_2_6_N68), .C2(
        npu_inst_pe_1_2_6_n77), .ZN(npu_inst_pe_1_2_6_n81) );
  INV_X1 npu_inst_pe_1_2_6_U42 ( .A(npu_inst_pe_1_2_6_n81), .ZN(
        npu_inst_pe_1_2_6_n98) );
  AOI222_X1 npu_inst_pe_1_2_6_U41 ( .A1(npu_inst_int_data_res_3__6__4_), .A2(
        npu_inst_pe_1_2_6_n1), .B1(npu_inst_pe_1_2_6_N77), .B2(
        npu_inst_pe_1_2_6_n76), .C1(npu_inst_pe_1_2_6_N69), .C2(
        npu_inst_pe_1_2_6_n77), .ZN(npu_inst_pe_1_2_6_n80) );
  INV_X1 npu_inst_pe_1_2_6_U40 ( .A(npu_inst_pe_1_2_6_n80), .ZN(
        npu_inst_pe_1_2_6_n36) );
  AOI222_X1 npu_inst_pe_1_2_6_U39 ( .A1(npu_inst_int_data_res_3__6__5_), .A2(
        npu_inst_pe_1_2_6_n1), .B1(npu_inst_pe_1_2_6_N78), .B2(
        npu_inst_pe_1_2_6_n76), .C1(npu_inst_pe_1_2_6_N70), .C2(
        npu_inst_pe_1_2_6_n77), .ZN(npu_inst_pe_1_2_6_n79) );
  INV_X1 npu_inst_pe_1_2_6_U38 ( .A(npu_inst_pe_1_2_6_n79), .ZN(
        npu_inst_pe_1_2_6_n35) );
  AOI222_X1 npu_inst_pe_1_2_6_U37 ( .A1(npu_inst_int_data_res_3__6__6_), .A2(
        npu_inst_pe_1_2_6_n1), .B1(npu_inst_pe_1_2_6_N79), .B2(
        npu_inst_pe_1_2_6_n76), .C1(npu_inst_pe_1_2_6_N71), .C2(
        npu_inst_pe_1_2_6_n77), .ZN(npu_inst_pe_1_2_6_n78) );
  INV_X1 npu_inst_pe_1_2_6_U36 ( .A(npu_inst_pe_1_2_6_n78), .ZN(
        npu_inst_pe_1_2_6_n34) );
  INV_X1 npu_inst_pe_1_2_6_U35 ( .A(npu_inst_pe_1_2_6_int_data_1_), .ZN(
        npu_inst_pe_1_2_6_n14) );
  AND2_X1 npu_inst_pe_1_2_6_U34 ( .A1(npu_inst_int_data_x_2__6__1_), .A2(
        npu_inst_pe_1_2_6_int_q_weight_1_), .ZN(npu_inst_pe_1_2_6_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_2_6_U33 ( .A1(npu_inst_int_data_x_2__6__0_), .A2(
        npu_inst_pe_1_2_6_int_q_weight_1_), .ZN(npu_inst_pe_1_2_6_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_2_6_U32 ( .A1(npu_inst_n57), .A2(
        npu_inst_int_data_y_3__6__1_), .B1(npu_inst_pe_1_2_6_n3), .B2(
        npu_inst_int_data_x_2__7__1_), .ZN(npu_inst_pe_1_2_6_n63) );
  AOI22_X1 npu_inst_pe_1_2_6_U31 ( .A1(npu_inst_n57), .A2(
        npu_inst_int_data_y_3__6__0_), .B1(npu_inst_pe_1_2_6_n3), .B2(
        npu_inst_int_data_x_2__7__0_), .ZN(npu_inst_pe_1_2_6_n61) );
  INV_X1 npu_inst_pe_1_2_6_U30 ( .A(npu_inst_pe_1_2_6_int_data_0_), .ZN(
        npu_inst_pe_1_2_6_n13) );
  INV_X1 npu_inst_pe_1_2_6_U29 ( .A(npu_inst_n70), .ZN(npu_inst_pe_1_2_6_n5)
         );
  OR3_X1 npu_inst_pe_1_2_6_U28 ( .A1(npu_inst_pe_1_2_6_n6), .A2(
        npu_inst_pe_1_2_6_n8), .A3(npu_inst_pe_1_2_6_n5), .ZN(
        npu_inst_pe_1_2_6_n56) );
  OR3_X1 npu_inst_pe_1_2_6_U27 ( .A1(npu_inst_pe_1_2_6_n5), .A2(
        npu_inst_pe_1_2_6_n8), .A3(npu_inst_pe_1_2_6_n7), .ZN(
        npu_inst_pe_1_2_6_n48) );
  INV_X1 npu_inst_pe_1_2_6_U26 ( .A(npu_inst_pe_1_2_6_n5), .ZN(
        npu_inst_pe_1_2_6_n4) );
  INV_X1 npu_inst_pe_1_2_6_U25 ( .A(npu_inst_n125), .ZN(npu_inst_pe_1_2_6_n12)
         );
  OR3_X1 npu_inst_pe_1_2_6_U24 ( .A1(npu_inst_pe_1_2_6_n4), .A2(
        npu_inst_pe_1_2_6_n8), .A3(npu_inst_pe_1_2_6_n7), .ZN(
        npu_inst_pe_1_2_6_n52) );
  OR3_X1 npu_inst_pe_1_2_6_U23 ( .A1(npu_inst_pe_1_2_6_n6), .A2(
        npu_inst_pe_1_2_6_n8), .A3(npu_inst_pe_1_2_6_n4), .ZN(
        npu_inst_pe_1_2_6_n60) );
  NOR2_X1 npu_inst_pe_1_2_6_U22 ( .A1(npu_inst_pe_1_2_6_n60), .A2(
        npu_inst_pe_1_2_6_n3), .ZN(npu_inst_pe_1_2_6_n58) );
  NOR2_X1 npu_inst_pe_1_2_6_U21 ( .A1(npu_inst_pe_1_2_6_n56), .A2(
        npu_inst_pe_1_2_6_n3), .ZN(npu_inst_pe_1_2_6_n54) );
  NOR2_X1 npu_inst_pe_1_2_6_U20 ( .A1(npu_inst_pe_1_2_6_n52), .A2(
        npu_inst_pe_1_2_6_n3), .ZN(npu_inst_pe_1_2_6_n50) );
  NOR2_X1 npu_inst_pe_1_2_6_U19 ( .A1(npu_inst_pe_1_2_6_n48), .A2(
        npu_inst_pe_1_2_6_n3), .ZN(npu_inst_pe_1_2_6_n46) );
  NOR2_X1 npu_inst_pe_1_2_6_U18 ( .A1(npu_inst_pe_1_2_6_n40), .A2(
        npu_inst_pe_1_2_6_n3), .ZN(npu_inst_pe_1_2_6_n38) );
  NOR2_X1 npu_inst_pe_1_2_6_U17 ( .A1(npu_inst_pe_1_2_6_n44), .A2(
        npu_inst_pe_1_2_6_n3), .ZN(npu_inst_pe_1_2_6_n42) );
  BUF_X1 npu_inst_pe_1_2_6_U16 ( .A(npu_inst_n102), .Z(npu_inst_pe_1_2_6_n8)
         );
  BUF_X1 npu_inst_pe_1_2_6_U15 ( .A(npu_inst_pe_1_2_6_n12), .Z(
        npu_inst_pe_1_2_6_n11) );
  BUF_X1 npu_inst_pe_1_2_6_U14 ( .A(npu_inst_pe_1_2_6_n12), .Z(
        npu_inst_pe_1_2_6_n10) );
  BUF_X1 npu_inst_pe_1_2_6_U13 ( .A(npu_inst_pe_1_2_6_n12), .Z(
        npu_inst_pe_1_2_6_n9) );
  INV_X1 npu_inst_pe_1_2_6_U12 ( .A(npu_inst_pe_1_2_6_n38), .ZN(
        npu_inst_pe_1_2_6_n118) );
  INV_X1 npu_inst_pe_1_2_6_U11 ( .A(npu_inst_pe_1_2_6_n58), .ZN(
        npu_inst_pe_1_2_6_n114) );
  INV_X1 npu_inst_pe_1_2_6_U10 ( .A(npu_inst_pe_1_2_6_n54), .ZN(
        npu_inst_pe_1_2_6_n115) );
  INV_X1 npu_inst_pe_1_2_6_U9 ( .A(npu_inst_pe_1_2_6_n50), .ZN(
        npu_inst_pe_1_2_6_n116) );
  INV_X1 npu_inst_pe_1_2_6_U8 ( .A(npu_inst_pe_1_2_6_n46), .ZN(
        npu_inst_pe_1_2_6_n117) );
  INV_X1 npu_inst_pe_1_2_6_U7 ( .A(npu_inst_pe_1_2_6_n42), .ZN(
        npu_inst_pe_1_2_6_n119) );
  BUF_X1 npu_inst_pe_1_2_6_U6 ( .A(npu_inst_n27), .Z(npu_inst_pe_1_2_6_n2) );
  BUF_X1 npu_inst_pe_1_2_6_U5 ( .A(npu_inst_n27), .Z(npu_inst_pe_1_2_6_n1) );
  NOR2_X1 npu_inst_pe_1_2_6_U4 ( .A1(npu_inst_pe_1_2_6_int_q_weight_0_), .A2(
        npu_inst_pe_1_2_6_n1), .ZN(npu_inst_pe_1_2_6_n76) );
  NOR2_X1 npu_inst_pe_1_2_6_U3 ( .A1(npu_inst_pe_1_2_6_n27), .A2(
        npu_inst_pe_1_2_6_n1), .ZN(npu_inst_pe_1_2_6_n77) );
  FA_X1 npu_inst_pe_1_2_6_sub_77_U2_1 ( .A(npu_inst_pe_1_2_6_int_q_acc_1_), 
        .B(npu_inst_pe_1_2_6_n14), .CI(npu_inst_pe_1_2_6_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_2_6_sub_77_carry_2_), .S(npu_inst_pe_1_2_6_N66) );
  FA_X1 npu_inst_pe_1_2_6_add_79_U1_1 ( .A(npu_inst_pe_1_2_6_int_q_acc_1_), 
        .B(npu_inst_pe_1_2_6_int_data_1_), .CI(
        npu_inst_pe_1_2_6_add_79_carry_1_), .CO(
        npu_inst_pe_1_2_6_add_79_carry_2_), .S(npu_inst_pe_1_2_6_N74) );
  NAND3_X1 npu_inst_pe_1_2_6_U109 ( .A1(npu_inst_pe_1_2_6_n5), .A2(
        npu_inst_pe_1_2_6_n7), .A3(npu_inst_pe_1_2_6_n8), .ZN(
        npu_inst_pe_1_2_6_n44) );
  NAND3_X1 npu_inst_pe_1_2_6_U108 ( .A1(npu_inst_pe_1_2_6_n4), .A2(
        npu_inst_pe_1_2_6_n7), .A3(npu_inst_pe_1_2_6_n8), .ZN(
        npu_inst_pe_1_2_6_n40) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_2_6_n34), .CK(
        npu_inst_pe_1_2_6_net3787), .RN(npu_inst_pe_1_2_6_n9), .Q(
        npu_inst_pe_1_2_6_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_2_6_n35), .CK(
        npu_inst_pe_1_2_6_net3787), .RN(npu_inst_pe_1_2_6_n9), .Q(
        npu_inst_pe_1_2_6_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_2_6_n36), .CK(
        npu_inst_pe_1_2_6_net3787), .RN(npu_inst_pe_1_2_6_n9), .Q(
        npu_inst_pe_1_2_6_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_2_6_n98), .CK(
        npu_inst_pe_1_2_6_net3787), .RN(npu_inst_pe_1_2_6_n9), .Q(
        npu_inst_pe_1_2_6_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_2_6_n99), .CK(
        npu_inst_pe_1_2_6_net3787), .RN(npu_inst_pe_1_2_6_n9), .Q(
        npu_inst_pe_1_2_6_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_2_6_n100), 
        .CK(npu_inst_pe_1_2_6_net3787), .RN(npu_inst_pe_1_2_6_n9), .Q(
        npu_inst_pe_1_2_6_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_2_6_n33), .CK(
        npu_inst_pe_1_2_6_net3787), .RN(npu_inst_pe_1_2_6_n9), .Q(
        npu_inst_pe_1_2_6_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_2_6_n101), 
        .CK(npu_inst_pe_1_2_6_net3787), .RN(npu_inst_pe_1_2_6_n9), .Q(
        npu_inst_pe_1_2_6_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_weight_reg_0_ ( .D(npu_inst_n111), .CK(
        npu_inst_pe_1_2_6_net3793), .RN(npu_inst_pe_1_2_6_n9), .Q(
        npu_inst_pe_1_2_6_int_q_weight_0_), .QN(npu_inst_pe_1_2_6_n27) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_weight_reg_1_ ( .D(npu_inst_n117), .CK(
        npu_inst_pe_1_2_6_net3793), .RN(npu_inst_pe_1_2_6_n9), .Q(
        npu_inst_pe_1_2_6_int_q_weight_1_), .QN(npu_inst_pe_1_2_6_n26) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_2_6_n113), 
        .CK(npu_inst_pe_1_2_6_net3793), .RN(npu_inst_pe_1_2_6_n9), .Q(
        npu_inst_pe_1_2_6_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_2_6_n107), 
        .CK(npu_inst_pe_1_2_6_net3793), .RN(npu_inst_pe_1_2_6_n9), .Q(
        npu_inst_pe_1_2_6_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_2_6_n112), 
        .CK(npu_inst_pe_1_2_6_net3793), .RN(npu_inst_pe_1_2_6_n10), .Q(
        npu_inst_pe_1_2_6_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_2_6_n106), 
        .CK(npu_inst_pe_1_2_6_net3793), .RN(npu_inst_pe_1_2_6_n10), .Q(
        npu_inst_pe_1_2_6_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_2_6_n111), 
        .CK(npu_inst_pe_1_2_6_net3793), .RN(npu_inst_pe_1_2_6_n10), .Q(
        npu_inst_pe_1_2_6_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_2_6_n105), 
        .CK(npu_inst_pe_1_2_6_net3793), .RN(npu_inst_pe_1_2_6_n10), .Q(
        npu_inst_pe_1_2_6_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_2_6_n110), 
        .CK(npu_inst_pe_1_2_6_net3793), .RN(npu_inst_pe_1_2_6_n10), .Q(
        npu_inst_pe_1_2_6_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_2_6_n104), 
        .CK(npu_inst_pe_1_2_6_net3793), .RN(npu_inst_pe_1_2_6_n10), .Q(
        npu_inst_pe_1_2_6_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_2_6_n109), 
        .CK(npu_inst_pe_1_2_6_net3793), .RN(npu_inst_pe_1_2_6_n10), .Q(
        npu_inst_pe_1_2_6_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_2_6_n103), 
        .CK(npu_inst_pe_1_2_6_net3793), .RN(npu_inst_pe_1_2_6_n10), .Q(
        npu_inst_pe_1_2_6_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_2_6_n108), 
        .CK(npu_inst_pe_1_2_6_net3793), .RN(npu_inst_pe_1_2_6_n10), .Q(
        npu_inst_pe_1_2_6_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_2_6_n102), 
        .CK(npu_inst_pe_1_2_6_net3793), .RN(npu_inst_pe_1_2_6_n10), .Q(
        npu_inst_pe_1_2_6_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_2_6_n86), 
        .CK(npu_inst_pe_1_2_6_net3793), .RN(npu_inst_pe_1_2_6_n10), .Q(
        npu_inst_pe_1_2_6_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_2_6_n87), 
        .CK(npu_inst_pe_1_2_6_net3793), .RN(npu_inst_pe_1_2_6_n10), .Q(
        npu_inst_pe_1_2_6_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_2_6_n88), 
        .CK(npu_inst_pe_1_2_6_net3793), .RN(npu_inst_pe_1_2_6_n11), .Q(
        npu_inst_pe_1_2_6_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_2_6_n89), 
        .CK(npu_inst_pe_1_2_6_net3793), .RN(npu_inst_pe_1_2_6_n11), .Q(
        npu_inst_pe_1_2_6_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_2_6_n90), 
        .CK(npu_inst_pe_1_2_6_net3793), .RN(npu_inst_pe_1_2_6_n11), .Q(
        npu_inst_pe_1_2_6_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_2_6_n91), 
        .CK(npu_inst_pe_1_2_6_net3793), .RN(npu_inst_pe_1_2_6_n11), .Q(
        npu_inst_pe_1_2_6_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_2_6_n92), 
        .CK(npu_inst_pe_1_2_6_net3793), .RN(npu_inst_pe_1_2_6_n11), .Q(
        npu_inst_pe_1_2_6_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_2_6_n93), 
        .CK(npu_inst_pe_1_2_6_net3793), .RN(npu_inst_pe_1_2_6_n11), .Q(
        npu_inst_pe_1_2_6_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_2_6_n94), 
        .CK(npu_inst_pe_1_2_6_net3793), .RN(npu_inst_pe_1_2_6_n11), .Q(
        npu_inst_pe_1_2_6_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_2_6_n95), 
        .CK(npu_inst_pe_1_2_6_net3793), .RN(npu_inst_pe_1_2_6_n11), .Q(
        npu_inst_pe_1_2_6_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_2_6_n96), 
        .CK(npu_inst_pe_1_2_6_net3793), .RN(npu_inst_pe_1_2_6_n11), .Q(
        npu_inst_pe_1_2_6_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_2_6_n97), 
        .CK(npu_inst_pe_1_2_6_net3793), .RN(npu_inst_pe_1_2_6_n11), .Q(
        npu_inst_pe_1_2_6_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_2_6_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_2_6_N84), .SE(1'b0), .GCK(npu_inst_pe_1_2_6_net3787) );
  CLKGATETST_X1 npu_inst_pe_1_2_6_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n64), .SE(1'b0), .GCK(npu_inst_pe_1_2_6_net3793) );
  MUX2_X1 npu_inst_pe_1_2_7_U162 ( .A(npu_inst_pe_1_2_7_n32), .B(
        npu_inst_pe_1_2_7_n29), .S(npu_inst_pe_1_2_7_n8), .Z(
        npu_inst_pe_1_2_7_N93) );
  MUX2_X1 npu_inst_pe_1_2_7_U161 ( .A(npu_inst_pe_1_2_7_n31), .B(
        npu_inst_pe_1_2_7_n30), .S(npu_inst_pe_1_2_7_n6), .Z(
        npu_inst_pe_1_2_7_n32) );
  MUX2_X1 npu_inst_pe_1_2_7_U160 ( .A(npu_inst_pe_1_2_7_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_2_7_int_q_reg_v_1__0_), .S(npu_inst_pe_1_2_7_n4), .Z(
        npu_inst_pe_1_2_7_n31) );
  MUX2_X1 npu_inst_pe_1_2_7_U159 ( .A(npu_inst_pe_1_2_7_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_2_7_int_q_reg_v_3__0_), .S(npu_inst_pe_1_2_7_n4), .Z(
        npu_inst_pe_1_2_7_n30) );
  MUX2_X1 npu_inst_pe_1_2_7_U158 ( .A(npu_inst_pe_1_2_7_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_2_7_int_q_reg_v_5__0_), .S(npu_inst_pe_1_2_7_n4), .Z(
        npu_inst_pe_1_2_7_n29) );
  MUX2_X1 npu_inst_pe_1_2_7_U157 ( .A(npu_inst_pe_1_2_7_n28), .B(
        npu_inst_pe_1_2_7_n23), .S(npu_inst_pe_1_2_7_n8), .Z(
        npu_inst_pe_1_2_7_N94) );
  MUX2_X1 npu_inst_pe_1_2_7_U156 ( .A(npu_inst_pe_1_2_7_n25), .B(
        npu_inst_pe_1_2_7_n24), .S(npu_inst_pe_1_2_7_n6), .Z(
        npu_inst_pe_1_2_7_n28) );
  MUX2_X1 npu_inst_pe_1_2_7_U155 ( .A(npu_inst_pe_1_2_7_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_2_7_int_q_reg_v_1__1_), .S(npu_inst_pe_1_2_7_n4), .Z(
        npu_inst_pe_1_2_7_n25) );
  MUX2_X1 npu_inst_pe_1_2_7_U154 ( .A(npu_inst_pe_1_2_7_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_2_7_int_q_reg_v_3__1_), .S(npu_inst_pe_1_2_7_n4), .Z(
        npu_inst_pe_1_2_7_n24) );
  MUX2_X1 npu_inst_pe_1_2_7_U153 ( .A(npu_inst_pe_1_2_7_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_2_7_int_q_reg_v_5__1_), .S(npu_inst_pe_1_2_7_n4), .Z(
        npu_inst_pe_1_2_7_n23) );
  MUX2_X1 npu_inst_pe_1_2_7_U152 ( .A(npu_inst_pe_1_2_7_n22), .B(
        npu_inst_pe_1_2_7_n19), .S(npu_inst_pe_1_2_7_n8), .Z(
        npu_inst_int_data_x_2__7__1_) );
  MUX2_X1 npu_inst_pe_1_2_7_U151 ( .A(npu_inst_pe_1_2_7_n21), .B(
        npu_inst_pe_1_2_7_n20), .S(npu_inst_pe_1_2_7_n6), .Z(
        npu_inst_pe_1_2_7_n22) );
  MUX2_X1 npu_inst_pe_1_2_7_U150 ( .A(npu_inst_pe_1_2_7_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_2_7_int_q_reg_h_1__1_), .S(npu_inst_pe_1_2_7_n4), .Z(
        npu_inst_pe_1_2_7_n21) );
  MUX2_X1 npu_inst_pe_1_2_7_U149 ( .A(npu_inst_pe_1_2_7_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_2_7_int_q_reg_h_3__1_), .S(npu_inst_pe_1_2_7_n4), .Z(
        npu_inst_pe_1_2_7_n20) );
  MUX2_X1 npu_inst_pe_1_2_7_U148 ( .A(npu_inst_pe_1_2_7_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_2_7_int_q_reg_h_5__1_), .S(npu_inst_pe_1_2_7_n4), .Z(
        npu_inst_pe_1_2_7_n19) );
  MUX2_X1 npu_inst_pe_1_2_7_U147 ( .A(npu_inst_pe_1_2_7_n18), .B(
        npu_inst_pe_1_2_7_n15), .S(npu_inst_pe_1_2_7_n8), .Z(
        npu_inst_int_data_x_2__7__0_) );
  MUX2_X1 npu_inst_pe_1_2_7_U146 ( .A(npu_inst_pe_1_2_7_n17), .B(
        npu_inst_pe_1_2_7_n16), .S(npu_inst_pe_1_2_7_n6), .Z(
        npu_inst_pe_1_2_7_n18) );
  MUX2_X1 npu_inst_pe_1_2_7_U145 ( .A(npu_inst_pe_1_2_7_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_2_7_int_q_reg_h_1__0_), .S(npu_inst_pe_1_2_7_n4), .Z(
        npu_inst_pe_1_2_7_n17) );
  MUX2_X1 npu_inst_pe_1_2_7_U144 ( .A(npu_inst_pe_1_2_7_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_2_7_int_q_reg_h_3__0_), .S(npu_inst_pe_1_2_7_n4), .Z(
        npu_inst_pe_1_2_7_n16) );
  MUX2_X1 npu_inst_pe_1_2_7_U143 ( .A(npu_inst_pe_1_2_7_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_2_7_int_q_reg_h_5__0_), .S(npu_inst_pe_1_2_7_n4), .Z(
        npu_inst_pe_1_2_7_n15) );
  XOR2_X1 npu_inst_pe_1_2_7_U142 ( .A(npu_inst_pe_1_2_7_int_data_0_), .B(
        npu_inst_pe_1_2_7_int_q_acc_0_), .Z(npu_inst_pe_1_2_7_N73) );
  AND2_X1 npu_inst_pe_1_2_7_U141 ( .A1(npu_inst_pe_1_2_7_int_q_acc_0_), .A2(
        npu_inst_pe_1_2_7_int_data_0_), .ZN(npu_inst_pe_1_2_7_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_2_7_U140 ( .A(npu_inst_pe_1_2_7_int_q_acc_0_), .B(
        npu_inst_pe_1_2_7_n13), .ZN(npu_inst_pe_1_2_7_N65) );
  OR2_X1 npu_inst_pe_1_2_7_U139 ( .A1(npu_inst_pe_1_2_7_n13), .A2(
        npu_inst_pe_1_2_7_int_q_acc_0_), .ZN(npu_inst_pe_1_2_7_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_2_7_U138 ( .A(npu_inst_pe_1_2_7_int_q_acc_2_), .B(
        npu_inst_pe_1_2_7_add_79_carry_2_), .Z(npu_inst_pe_1_2_7_N75) );
  AND2_X1 npu_inst_pe_1_2_7_U137 ( .A1(npu_inst_pe_1_2_7_add_79_carry_2_), 
        .A2(npu_inst_pe_1_2_7_int_q_acc_2_), .ZN(
        npu_inst_pe_1_2_7_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_2_7_U136 ( .A(npu_inst_pe_1_2_7_int_q_acc_3_), .B(
        npu_inst_pe_1_2_7_add_79_carry_3_), .Z(npu_inst_pe_1_2_7_N76) );
  AND2_X1 npu_inst_pe_1_2_7_U135 ( .A1(npu_inst_pe_1_2_7_add_79_carry_3_), 
        .A2(npu_inst_pe_1_2_7_int_q_acc_3_), .ZN(
        npu_inst_pe_1_2_7_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_2_7_U134 ( .A(npu_inst_pe_1_2_7_int_q_acc_4_), .B(
        npu_inst_pe_1_2_7_add_79_carry_4_), .Z(npu_inst_pe_1_2_7_N77) );
  AND2_X1 npu_inst_pe_1_2_7_U133 ( .A1(npu_inst_pe_1_2_7_add_79_carry_4_), 
        .A2(npu_inst_pe_1_2_7_int_q_acc_4_), .ZN(
        npu_inst_pe_1_2_7_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_2_7_U132 ( .A(npu_inst_pe_1_2_7_int_q_acc_5_), .B(
        npu_inst_pe_1_2_7_add_79_carry_5_), .Z(npu_inst_pe_1_2_7_N78) );
  AND2_X1 npu_inst_pe_1_2_7_U131 ( .A1(npu_inst_pe_1_2_7_add_79_carry_5_), 
        .A2(npu_inst_pe_1_2_7_int_q_acc_5_), .ZN(
        npu_inst_pe_1_2_7_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_2_7_U130 ( .A(npu_inst_pe_1_2_7_int_q_acc_6_), .B(
        npu_inst_pe_1_2_7_add_79_carry_6_), .Z(npu_inst_pe_1_2_7_N79) );
  AND2_X1 npu_inst_pe_1_2_7_U129 ( .A1(npu_inst_pe_1_2_7_add_79_carry_6_), 
        .A2(npu_inst_pe_1_2_7_int_q_acc_6_), .ZN(
        npu_inst_pe_1_2_7_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_2_7_U128 ( .A(npu_inst_pe_1_2_7_int_q_acc_7_), .B(
        npu_inst_pe_1_2_7_add_79_carry_7_), .Z(npu_inst_pe_1_2_7_N80) );
  XNOR2_X1 npu_inst_pe_1_2_7_U127 ( .A(npu_inst_pe_1_2_7_sub_77_carry_2_), .B(
        npu_inst_pe_1_2_7_int_q_acc_2_), .ZN(npu_inst_pe_1_2_7_N67) );
  OR2_X1 npu_inst_pe_1_2_7_U126 ( .A1(npu_inst_pe_1_2_7_int_q_acc_2_), .A2(
        npu_inst_pe_1_2_7_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_2_7_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_2_7_U125 ( .A(npu_inst_pe_1_2_7_sub_77_carry_3_), .B(
        npu_inst_pe_1_2_7_int_q_acc_3_), .ZN(npu_inst_pe_1_2_7_N68) );
  OR2_X1 npu_inst_pe_1_2_7_U124 ( .A1(npu_inst_pe_1_2_7_int_q_acc_3_), .A2(
        npu_inst_pe_1_2_7_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_2_7_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_2_7_U123 ( .A(npu_inst_pe_1_2_7_sub_77_carry_4_), .B(
        npu_inst_pe_1_2_7_int_q_acc_4_), .ZN(npu_inst_pe_1_2_7_N69) );
  OR2_X1 npu_inst_pe_1_2_7_U122 ( .A1(npu_inst_pe_1_2_7_int_q_acc_4_), .A2(
        npu_inst_pe_1_2_7_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_2_7_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_2_7_U121 ( .A(npu_inst_pe_1_2_7_sub_77_carry_5_), .B(
        npu_inst_pe_1_2_7_int_q_acc_5_), .ZN(npu_inst_pe_1_2_7_N70) );
  OR2_X1 npu_inst_pe_1_2_7_U120 ( .A1(npu_inst_pe_1_2_7_int_q_acc_5_), .A2(
        npu_inst_pe_1_2_7_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_2_7_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_2_7_U119 ( .A(npu_inst_pe_1_2_7_sub_77_carry_6_), .B(
        npu_inst_pe_1_2_7_int_q_acc_6_), .ZN(npu_inst_pe_1_2_7_N71) );
  OR2_X1 npu_inst_pe_1_2_7_U118 ( .A1(npu_inst_pe_1_2_7_int_q_acc_6_), .A2(
        npu_inst_pe_1_2_7_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_2_7_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_2_7_U117 ( .A(npu_inst_pe_1_2_7_int_q_acc_7_), .B(
        npu_inst_pe_1_2_7_sub_77_carry_7_), .ZN(npu_inst_pe_1_2_7_N72) );
  INV_X1 npu_inst_pe_1_2_7_U116 ( .A(npu_inst_n78), .ZN(npu_inst_pe_1_2_7_n7)
         );
  INV_X1 npu_inst_pe_1_2_7_U115 ( .A(npu_inst_pe_1_2_7_n7), .ZN(
        npu_inst_pe_1_2_7_n6) );
  INV_X1 npu_inst_pe_1_2_7_U114 ( .A(npu_inst_n57), .ZN(npu_inst_pe_1_2_7_n3)
         );
  AOI22_X1 npu_inst_pe_1_2_7_U113 ( .A1(npu_inst_int_data_y_3__7__0_), .A2(
        npu_inst_pe_1_2_7_n58), .B1(npu_inst_pe_1_2_7_n114), .B2(
        npu_inst_pe_1_2_7_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_2_7_n57) );
  INV_X1 npu_inst_pe_1_2_7_U112 ( .A(npu_inst_pe_1_2_7_n57), .ZN(
        npu_inst_pe_1_2_7_n108) );
  AOI22_X1 npu_inst_pe_1_2_7_U111 ( .A1(npu_inst_int_data_y_3__7__0_), .A2(
        npu_inst_pe_1_2_7_n54), .B1(npu_inst_pe_1_2_7_n115), .B2(
        npu_inst_pe_1_2_7_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_2_7_n53) );
  INV_X1 npu_inst_pe_1_2_7_U110 ( .A(npu_inst_pe_1_2_7_n53), .ZN(
        npu_inst_pe_1_2_7_n109) );
  AOI22_X1 npu_inst_pe_1_2_7_U107 ( .A1(npu_inst_int_data_y_3__7__0_), .A2(
        npu_inst_pe_1_2_7_n50), .B1(npu_inst_pe_1_2_7_n116), .B2(
        npu_inst_pe_1_2_7_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_2_7_n49) );
  INV_X1 npu_inst_pe_1_2_7_U106 ( .A(npu_inst_pe_1_2_7_n49), .ZN(
        npu_inst_pe_1_2_7_n110) );
  AOI22_X1 npu_inst_pe_1_2_7_U105 ( .A1(npu_inst_int_data_y_3__7__0_), .A2(
        npu_inst_pe_1_2_7_n46), .B1(npu_inst_pe_1_2_7_n117), .B2(
        npu_inst_pe_1_2_7_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_2_7_n45) );
  INV_X1 npu_inst_pe_1_2_7_U104 ( .A(npu_inst_pe_1_2_7_n45), .ZN(
        npu_inst_pe_1_2_7_n111) );
  AOI22_X1 npu_inst_pe_1_2_7_U103 ( .A1(npu_inst_int_data_y_3__7__0_), .A2(
        npu_inst_pe_1_2_7_n42), .B1(npu_inst_pe_1_2_7_n119), .B2(
        npu_inst_pe_1_2_7_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_2_7_n41) );
  INV_X1 npu_inst_pe_1_2_7_U102 ( .A(npu_inst_pe_1_2_7_n41), .ZN(
        npu_inst_pe_1_2_7_n112) );
  AOI22_X1 npu_inst_pe_1_2_7_U101 ( .A1(npu_inst_int_data_y_3__7__1_), .A2(
        npu_inst_pe_1_2_7_n58), .B1(npu_inst_pe_1_2_7_n114), .B2(
        npu_inst_pe_1_2_7_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_2_7_n59) );
  INV_X1 npu_inst_pe_1_2_7_U100 ( .A(npu_inst_pe_1_2_7_n59), .ZN(
        npu_inst_pe_1_2_7_n102) );
  AOI22_X1 npu_inst_pe_1_2_7_U99 ( .A1(npu_inst_int_data_y_3__7__1_), .A2(
        npu_inst_pe_1_2_7_n54), .B1(npu_inst_pe_1_2_7_n115), .B2(
        npu_inst_pe_1_2_7_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_2_7_n55) );
  INV_X1 npu_inst_pe_1_2_7_U98 ( .A(npu_inst_pe_1_2_7_n55), .ZN(
        npu_inst_pe_1_2_7_n103) );
  AOI22_X1 npu_inst_pe_1_2_7_U97 ( .A1(npu_inst_int_data_y_3__7__1_), .A2(
        npu_inst_pe_1_2_7_n50), .B1(npu_inst_pe_1_2_7_n116), .B2(
        npu_inst_pe_1_2_7_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_2_7_n51) );
  INV_X1 npu_inst_pe_1_2_7_U96 ( .A(npu_inst_pe_1_2_7_n51), .ZN(
        npu_inst_pe_1_2_7_n104) );
  AOI22_X1 npu_inst_pe_1_2_7_U95 ( .A1(npu_inst_int_data_y_3__7__1_), .A2(
        npu_inst_pe_1_2_7_n46), .B1(npu_inst_pe_1_2_7_n117), .B2(
        npu_inst_pe_1_2_7_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_2_7_n47) );
  INV_X1 npu_inst_pe_1_2_7_U94 ( .A(npu_inst_pe_1_2_7_n47), .ZN(
        npu_inst_pe_1_2_7_n105) );
  AOI22_X1 npu_inst_pe_1_2_7_U93 ( .A1(npu_inst_int_data_y_3__7__1_), .A2(
        npu_inst_pe_1_2_7_n42), .B1(npu_inst_pe_1_2_7_n119), .B2(
        npu_inst_pe_1_2_7_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_2_7_n43) );
  INV_X1 npu_inst_pe_1_2_7_U92 ( .A(npu_inst_pe_1_2_7_n43), .ZN(
        npu_inst_pe_1_2_7_n106) );
  AOI22_X1 npu_inst_pe_1_2_7_U91 ( .A1(npu_inst_pe_1_2_7_n38), .A2(
        npu_inst_int_data_y_3__7__1_), .B1(npu_inst_pe_1_2_7_n118), .B2(
        npu_inst_pe_1_2_7_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_2_7_n39) );
  INV_X1 npu_inst_pe_1_2_7_U90 ( .A(npu_inst_pe_1_2_7_n39), .ZN(
        npu_inst_pe_1_2_7_n107) );
  AOI22_X1 npu_inst_pe_1_2_7_U89 ( .A1(npu_inst_pe_1_2_7_n38), .A2(
        npu_inst_int_data_y_3__7__0_), .B1(npu_inst_pe_1_2_7_n118), .B2(
        npu_inst_pe_1_2_7_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_2_7_n37) );
  INV_X1 npu_inst_pe_1_2_7_U88 ( .A(npu_inst_pe_1_2_7_n37), .ZN(
        npu_inst_pe_1_2_7_n113) );
  AND2_X1 npu_inst_pe_1_2_7_U87 ( .A1(npu_inst_pe_1_2_7_N93), .A2(npu_inst_n57), .ZN(npu_inst_int_data_y_2__7__0_) );
  AND2_X1 npu_inst_pe_1_2_7_U86 ( .A1(npu_inst_n57), .A2(npu_inst_pe_1_2_7_N94), .ZN(npu_inst_int_data_y_2__7__1_) );
  NOR3_X1 npu_inst_pe_1_2_7_U85 ( .A1(npu_inst_pe_1_2_7_n26), .A2(npu_inst_n57), .A3(npu_inst_int_ckg[40]), .ZN(npu_inst_pe_1_2_7_n85) );
  OR2_X1 npu_inst_pe_1_2_7_U84 ( .A1(npu_inst_pe_1_2_7_n85), .A2(
        npu_inst_pe_1_2_7_n2), .ZN(npu_inst_pe_1_2_7_N84) );
  AND2_X1 npu_inst_pe_1_2_7_U83 ( .A1(npu_inst_pe_1_2_7_int_q_acc_0_), .A2(
        npu_inst_pe_1_2_7_n1), .ZN(npu_inst_int_data_res_2__7__0_) );
  AND2_X1 npu_inst_pe_1_2_7_U82 ( .A1(npu_inst_pe_1_2_7_n2), .A2(
        npu_inst_pe_1_2_7_int_q_acc_7_), .ZN(npu_inst_int_data_res_2__7__7_)
         );
  AND2_X1 npu_inst_pe_1_2_7_U81 ( .A1(npu_inst_pe_1_2_7_int_q_acc_1_), .A2(
        npu_inst_pe_1_2_7_n1), .ZN(npu_inst_int_data_res_2__7__1_) );
  AND2_X1 npu_inst_pe_1_2_7_U80 ( .A1(npu_inst_pe_1_2_7_int_q_acc_2_), .A2(
        npu_inst_pe_1_2_7_n1), .ZN(npu_inst_int_data_res_2__7__2_) );
  AND2_X1 npu_inst_pe_1_2_7_U79 ( .A1(npu_inst_pe_1_2_7_int_q_acc_3_), .A2(
        npu_inst_pe_1_2_7_n2), .ZN(npu_inst_int_data_res_2__7__3_) );
  AND2_X1 npu_inst_pe_1_2_7_U78 ( .A1(npu_inst_pe_1_2_7_int_q_acc_4_), .A2(
        npu_inst_pe_1_2_7_n2), .ZN(npu_inst_int_data_res_2__7__4_) );
  AND2_X1 npu_inst_pe_1_2_7_U77 ( .A1(npu_inst_pe_1_2_7_int_q_acc_5_), .A2(
        npu_inst_pe_1_2_7_n2), .ZN(npu_inst_int_data_res_2__7__5_) );
  AND2_X1 npu_inst_pe_1_2_7_U76 ( .A1(npu_inst_pe_1_2_7_int_q_acc_6_), .A2(
        npu_inst_pe_1_2_7_n2), .ZN(npu_inst_int_data_res_2__7__6_) );
  AOI222_X1 npu_inst_pe_1_2_7_U75 ( .A1(npu_inst_int_data_res_3__7__0_), .A2(
        npu_inst_pe_1_2_7_n1), .B1(npu_inst_pe_1_2_7_N73), .B2(
        npu_inst_pe_1_2_7_n76), .C1(npu_inst_pe_1_2_7_N65), .C2(
        npu_inst_pe_1_2_7_n77), .ZN(npu_inst_pe_1_2_7_n84) );
  INV_X1 npu_inst_pe_1_2_7_U74 ( .A(npu_inst_pe_1_2_7_n84), .ZN(
        npu_inst_pe_1_2_7_n101) );
  AOI222_X1 npu_inst_pe_1_2_7_U73 ( .A1(npu_inst_int_data_res_3__7__7_), .A2(
        npu_inst_pe_1_2_7_n1), .B1(npu_inst_pe_1_2_7_N80), .B2(
        npu_inst_pe_1_2_7_n76), .C1(npu_inst_pe_1_2_7_N72), .C2(
        npu_inst_pe_1_2_7_n77), .ZN(npu_inst_pe_1_2_7_n75) );
  INV_X1 npu_inst_pe_1_2_7_U72 ( .A(npu_inst_pe_1_2_7_n75), .ZN(
        npu_inst_pe_1_2_7_n33) );
  AOI222_X1 npu_inst_pe_1_2_7_U71 ( .A1(npu_inst_int_data_res_3__7__1_), .A2(
        npu_inst_pe_1_2_7_n1), .B1(npu_inst_pe_1_2_7_N74), .B2(
        npu_inst_pe_1_2_7_n76), .C1(npu_inst_pe_1_2_7_N66), .C2(
        npu_inst_pe_1_2_7_n77), .ZN(npu_inst_pe_1_2_7_n83) );
  INV_X1 npu_inst_pe_1_2_7_U70 ( .A(npu_inst_pe_1_2_7_n83), .ZN(
        npu_inst_pe_1_2_7_n100) );
  AOI222_X1 npu_inst_pe_1_2_7_U69 ( .A1(npu_inst_int_data_res_3__7__2_), .A2(
        npu_inst_pe_1_2_7_n1), .B1(npu_inst_pe_1_2_7_N75), .B2(
        npu_inst_pe_1_2_7_n76), .C1(npu_inst_pe_1_2_7_N67), .C2(
        npu_inst_pe_1_2_7_n77), .ZN(npu_inst_pe_1_2_7_n82) );
  INV_X1 npu_inst_pe_1_2_7_U68 ( .A(npu_inst_pe_1_2_7_n82), .ZN(
        npu_inst_pe_1_2_7_n99) );
  AOI222_X1 npu_inst_pe_1_2_7_U67 ( .A1(npu_inst_int_data_res_3__7__3_), .A2(
        npu_inst_pe_1_2_7_n1), .B1(npu_inst_pe_1_2_7_N76), .B2(
        npu_inst_pe_1_2_7_n76), .C1(npu_inst_pe_1_2_7_N68), .C2(
        npu_inst_pe_1_2_7_n77), .ZN(npu_inst_pe_1_2_7_n81) );
  INV_X1 npu_inst_pe_1_2_7_U66 ( .A(npu_inst_pe_1_2_7_n81), .ZN(
        npu_inst_pe_1_2_7_n98) );
  AOI222_X1 npu_inst_pe_1_2_7_U65 ( .A1(npu_inst_int_data_res_3__7__4_), .A2(
        npu_inst_pe_1_2_7_n1), .B1(npu_inst_pe_1_2_7_N77), .B2(
        npu_inst_pe_1_2_7_n76), .C1(npu_inst_pe_1_2_7_N69), .C2(
        npu_inst_pe_1_2_7_n77), .ZN(npu_inst_pe_1_2_7_n80) );
  INV_X1 npu_inst_pe_1_2_7_U64 ( .A(npu_inst_pe_1_2_7_n80), .ZN(
        npu_inst_pe_1_2_7_n36) );
  AOI222_X1 npu_inst_pe_1_2_7_U63 ( .A1(npu_inst_int_data_res_3__7__5_), .A2(
        npu_inst_pe_1_2_7_n1), .B1(npu_inst_pe_1_2_7_N78), .B2(
        npu_inst_pe_1_2_7_n76), .C1(npu_inst_pe_1_2_7_N70), .C2(
        npu_inst_pe_1_2_7_n77), .ZN(npu_inst_pe_1_2_7_n79) );
  INV_X1 npu_inst_pe_1_2_7_U62 ( .A(npu_inst_pe_1_2_7_n79), .ZN(
        npu_inst_pe_1_2_7_n35) );
  AOI222_X1 npu_inst_pe_1_2_7_U61 ( .A1(npu_inst_int_data_res_3__7__6_), .A2(
        npu_inst_pe_1_2_7_n1), .B1(npu_inst_pe_1_2_7_N79), .B2(
        npu_inst_pe_1_2_7_n76), .C1(npu_inst_pe_1_2_7_N71), .C2(
        npu_inst_pe_1_2_7_n77), .ZN(npu_inst_pe_1_2_7_n78) );
  INV_X1 npu_inst_pe_1_2_7_U60 ( .A(npu_inst_pe_1_2_7_n78), .ZN(
        npu_inst_pe_1_2_7_n34) );
  INV_X1 npu_inst_pe_1_2_7_U59 ( .A(npu_inst_pe_1_2_7_int_data_1_), .ZN(
        npu_inst_pe_1_2_7_n14) );
  AND2_X1 npu_inst_pe_1_2_7_U58 ( .A1(npu_inst_int_data_x_2__7__1_), .A2(
        npu_inst_pe_1_2_7_int_q_weight_1_), .ZN(npu_inst_pe_1_2_7_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_2_7_U57 ( .A1(npu_inst_int_data_x_2__7__0_), .A2(
        npu_inst_pe_1_2_7_int_q_weight_1_), .ZN(npu_inst_pe_1_2_7_int_data_0_)
         );
  NAND2_X1 npu_inst_pe_1_2_7_U56 ( .A1(npu_inst_pe_1_2_7_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_2_7_n60), .ZN(npu_inst_pe_1_2_7_n74) );
  OAI21_X1 npu_inst_pe_1_2_7_U55 ( .B1(npu_inst_pe_1_2_7_n63), .B2(
        npu_inst_pe_1_2_7_n60), .A(npu_inst_pe_1_2_7_n74), .ZN(
        npu_inst_pe_1_2_7_n97) );
  NAND2_X1 npu_inst_pe_1_2_7_U54 ( .A1(npu_inst_pe_1_2_7_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_2_7_n60), .ZN(npu_inst_pe_1_2_7_n73) );
  OAI21_X1 npu_inst_pe_1_2_7_U53 ( .B1(npu_inst_pe_1_2_7_n61), .B2(
        npu_inst_pe_1_2_7_n60), .A(npu_inst_pe_1_2_7_n73), .ZN(
        npu_inst_pe_1_2_7_n96) );
  NAND2_X1 npu_inst_pe_1_2_7_U52 ( .A1(npu_inst_pe_1_2_7_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_2_7_n56), .ZN(npu_inst_pe_1_2_7_n72) );
  OAI21_X1 npu_inst_pe_1_2_7_U51 ( .B1(npu_inst_pe_1_2_7_n63), .B2(
        npu_inst_pe_1_2_7_n56), .A(npu_inst_pe_1_2_7_n72), .ZN(
        npu_inst_pe_1_2_7_n95) );
  NAND2_X1 npu_inst_pe_1_2_7_U50 ( .A1(npu_inst_pe_1_2_7_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_2_7_n56), .ZN(npu_inst_pe_1_2_7_n71) );
  OAI21_X1 npu_inst_pe_1_2_7_U49 ( .B1(npu_inst_pe_1_2_7_n61), .B2(
        npu_inst_pe_1_2_7_n56), .A(npu_inst_pe_1_2_7_n71), .ZN(
        npu_inst_pe_1_2_7_n94) );
  NAND2_X1 npu_inst_pe_1_2_7_U48 ( .A1(npu_inst_pe_1_2_7_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_2_7_n52), .ZN(npu_inst_pe_1_2_7_n70) );
  OAI21_X1 npu_inst_pe_1_2_7_U47 ( .B1(npu_inst_pe_1_2_7_n63), .B2(
        npu_inst_pe_1_2_7_n52), .A(npu_inst_pe_1_2_7_n70), .ZN(
        npu_inst_pe_1_2_7_n93) );
  NAND2_X1 npu_inst_pe_1_2_7_U46 ( .A1(npu_inst_pe_1_2_7_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_2_7_n52), .ZN(npu_inst_pe_1_2_7_n69) );
  OAI21_X1 npu_inst_pe_1_2_7_U45 ( .B1(npu_inst_pe_1_2_7_n61), .B2(
        npu_inst_pe_1_2_7_n52), .A(npu_inst_pe_1_2_7_n69), .ZN(
        npu_inst_pe_1_2_7_n92) );
  NAND2_X1 npu_inst_pe_1_2_7_U44 ( .A1(npu_inst_pe_1_2_7_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_2_7_n48), .ZN(npu_inst_pe_1_2_7_n68) );
  OAI21_X1 npu_inst_pe_1_2_7_U43 ( .B1(npu_inst_pe_1_2_7_n63), .B2(
        npu_inst_pe_1_2_7_n48), .A(npu_inst_pe_1_2_7_n68), .ZN(
        npu_inst_pe_1_2_7_n91) );
  NAND2_X1 npu_inst_pe_1_2_7_U42 ( .A1(npu_inst_pe_1_2_7_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_2_7_n48), .ZN(npu_inst_pe_1_2_7_n67) );
  OAI21_X1 npu_inst_pe_1_2_7_U41 ( .B1(npu_inst_pe_1_2_7_n61), .B2(
        npu_inst_pe_1_2_7_n48), .A(npu_inst_pe_1_2_7_n67), .ZN(
        npu_inst_pe_1_2_7_n90) );
  NAND2_X1 npu_inst_pe_1_2_7_U40 ( .A1(npu_inst_pe_1_2_7_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_2_7_n44), .ZN(npu_inst_pe_1_2_7_n66) );
  OAI21_X1 npu_inst_pe_1_2_7_U39 ( .B1(npu_inst_pe_1_2_7_n63), .B2(
        npu_inst_pe_1_2_7_n44), .A(npu_inst_pe_1_2_7_n66), .ZN(
        npu_inst_pe_1_2_7_n89) );
  NAND2_X1 npu_inst_pe_1_2_7_U38 ( .A1(npu_inst_pe_1_2_7_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_2_7_n44), .ZN(npu_inst_pe_1_2_7_n65) );
  OAI21_X1 npu_inst_pe_1_2_7_U37 ( .B1(npu_inst_pe_1_2_7_n61), .B2(
        npu_inst_pe_1_2_7_n44), .A(npu_inst_pe_1_2_7_n65), .ZN(
        npu_inst_pe_1_2_7_n88) );
  NAND2_X1 npu_inst_pe_1_2_7_U36 ( .A1(npu_inst_pe_1_2_7_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_2_7_n40), .ZN(npu_inst_pe_1_2_7_n64) );
  OAI21_X1 npu_inst_pe_1_2_7_U35 ( .B1(npu_inst_pe_1_2_7_n63), .B2(
        npu_inst_pe_1_2_7_n40), .A(npu_inst_pe_1_2_7_n64), .ZN(
        npu_inst_pe_1_2_7_n87) );
  NAND2_X1 npu_inst_pe_1_2_7_U34 ( .A1(npu_inst_pe_1_2_7_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_2_7_n40), .ZN(npu_inst_pe_1_2_7_n62) );
  OAI21_X1 npu_inst_pe_1_2_7_U33 ( .B1(npu_inst_pe_1_2_7_n61), .B2(
        npu_inst_pe_1_2_7_n40), .A(npu_inst_pe_1_2_7_n62), .ZN(
        npu_inst_pe_1_2_7_n86) );
  INV_X1 npu_inst_pe_1_2_7_U32 ( .A(npu_inst_pe_1_2_7_int_data_0_), .ZN(
        npu_inst_pe_1_2_7_n13) );
  AOI22_X1 npu_inst_pe_1_2_7_U31 ( .A1(npu_inst_n57), .A2(
        npu_inst_int_data_y_3__7__1_), .B1(npu_inst_pe_1_2_7_n3), .B2(
        int_i_data_h_npu3[1]), .ZN(npu_inst_pe_1_2_7_n63) );
  AOI22_X1 npu_inst_pe_1_2_7_U30 ( .A1(npu_inst_n57), .A2(
        npu_inst_int_data_y_3__7__0_), .B1(npu_inst_pe_1_2_7_n3), .B2(
        int_i_data_h_npu3[0]), .ZN(npu_inst_pe_1_2_7_n61) );
  INV_X1 npu_inst_pe_1_2_7_U29 ( .A(npu_inst_n70), .ZN(npu_inst_pe_1_2_7_n5)
         );
  OR3_X1 npu_inst_pe_1_2_7_U28 ( .A1(npu_inst_pe_1_2_7_n6), .A2(
        npu_inst_pe_1_2_7_n8), .A3(npu_inst_pe_1_2_7_n5), .ZN(
        npu_inst_pe_1_2_7_n56) );
  OR3_X1 npu_inst_pe_1_2_7_U27 ( .A1(npu_inst_pe_1_2_7_n5), .A2(
        npu_inst_pe_1_2_7_n8), .A3(npu_inst_pe_1_2_7_n7), .ZN(
        npu_inst_pe_1_2_7_n48) );
  INV_X1 npu_inst_pe_1_2_7_U26 ( .A(npu_inst_pe_1_2_7_n5), .ZN(
        npu_inst_pe_1_2_7_n4) );
  INV_X1 npu_inst_pe_1_2_7_U25 ( .A(npu_inst_n125), .ZN(npu_inst_pe_1_2_7_n12)
         );
  OR3_X1 npu_inst_pe_1_2_7_U24 ( .A1(npu_inst_pe_1_2_7_n4), .A2(
        npu_inst_pe_1_2_7_n8), .A3(npu_inst_pe_1_2_7_n7), .ZN(
        npu_inst_pe_1_2_7_n52) );
  OR3_X1 npu_inst_pe_1_2_7_U23 ( .A1(npu_inst_pe_1_2_7_n6), .A2(
        npu_inst_pe_1_2_7_n8), .A3(npu_inst_pe_1_2_7_n4), .ZN(
        npu_inst_pe_1_2_7_n60) );
  NOR2_X1 npu_inst_pe_1_2_7_U22 ( .A1(npu_inst_pe_1_2_7_n60), .A2(
        npu_inst_pe_1_2_7_n3), .ZN(npu_inst_pe_1_2_7_n58) );
  NOR2_X1 npu_inst_pe_1_2_7_U21 ( .A1(npu_inst_pe_1_2_7_n56), .A2(
        npu_inst_pe_1_2_7_n3), .ZN(npu_inst_pe_1_2_7_n54) );
  NOR2_X1 npu_inst_pe_1_2_7_U20 ( .A1(npu_inst_pe_1_2_7_n52), .A2(
        npu_inst_pe_1_2_7_n3), .ZN(npu_inst_pe_1_2_7_n50) );
  NOR2_X1 npu_inst_pe_1_2_7_U19 ( .A1(npu_inst_pe_1_2_7_n48), .A2(
        npu_inst_pe_1_2_7_n3), .ZN(npu_inst_pe_1_2_7_n46) );
  NOR2_X1 npu_inst_pe_1_2_7_U18 ( .A1(npu_inst_pe_1_2_7_n40), .A2(
        npu_inst_pe_1_2_7_n3), .ZN(npu_inst_pe_1_2_7_n38) );
  NOR2_X1 npu_inst_pe_1_2_7_U17 ( .A1(npu_inst_pe_1_2_7_n44), .A2(
        npu_inst_pe_1_2_7_n3), .ZN(npu_inst_pe_1_2_7_n42) );
  BUF_X1 npu_inst_pe_1_2_7_U16 ( .A(npu_inst_n102), .Z(npu_inst_pe_1_2_7_n8)
         );
  BUF_X1 npu_inst_pe_1_2_7_U15 ( .A(npu_inst_pe_1_2_7_n12), .Z(
        npu_inst_pe_1_2_7_n11) );
  BUF_X1 npu_inst_pe_1_2_7_U14 ( .A(npu_inst_pe_1_2_7_n12), .Z(
        npu_inst_pe_1_2_7_n10) );
  BUF_X1 npu_inst_pe_1_2_7_U13 ( .A(npu_inst_pe_1_2_7_n12), .Z(
        npu_inst_pe_1_2_7_n9) );
  INV_X1 npu_inst_pe_1_2_7_U12 ( .A(npu_inst_pe_1_2_7_n38), .ZN(
        npu_inst_pe_1_2_7_n118) );
  INV_X1 npu_inst_pe_1_2_7_U11 ( .A(npu_inst_pe_1_2_7_n58), .ZN(
        npu_inst_pe_1_2_7_n114) );
  INV_X1 npu_inst_pe_1_2_7_U10 ( .A(npu_inst_pe_1_2_7_n54), .ZN(
        npu_inst_pe_1_2_7_n115) );
  INV_X1 npu_inst_pe_1_2_7_U9 ( .A(npu_inst_pe_1_2_7_n50), .ZN(
        npu_inst_pe_1_2_7_n116) );
  INV_X1 npu_inst_pe_1_2_7_U8 ( .A(npu_inst_pe_1_2_7_n46), .ZN(
        npu_inst_pe_1_2_7_n117) );
  INV_X1 npu_inst_pe_1_2_7_U7 ( .A(npu_inst_pe_1_2_7_n42), .ZN(
        npu_inst_pe_1_2_7_n119) );
  BUF_X1 npu_inst_pe_1_2_7_U6 ( .A(npu_inst_n27), .Z(npu_inst_pe_1_2_7_n2) );
  BUF_X1 npu_inst_pe_1_2_7_U5 ( .A(npu_inst_n27), .Z(npu_inst_pe_1_2_7_n1) );
  NOR2_X1 npu_inst_pe_1_2_7_U4 ( .A1(npu_inst_pe_1_2_7_int_q_weight_0_), .A2(
        npu_inst_pe_1_2_7_n1), .ZN(npu_inst_pe_1_2_7_n76) );
  NOR2_X1 npu_inst_pe_1_2_7_U3 ( .A1(npu_inst_pe_1_2_7_n27), .A2(
        npu_inst_pe_1_2_7_n1), .ZN(npu_inst_pe_1_2_7_n77) );
  FA_X1 npu_inst_pe_1_2_7_sub_77_U2_1 ( .A(npu_inst_pe_1_2_7_int_q_acc_1_), 
        .B(npu_inst_pe_1_2_7_n14), .CI(npu_inst_pe_1_2_7_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_2_7_sub_77_carry_2_), .S(npu_inst_pe_1_2_7_N66) );
  FA_X1 npu_inst_pe_1_2_7_add_79_U1_1 ( .A(npu_inst_pe_1_2_7_int_q_acc_1_), 
        .B(npu_inst_pe_1_2_7_int_data_1_), .CI(
        npu_inst_pe_1_2_7_add_79_carry_1_), .CO(
        npu_inst_pe_1_2_7_add_79_carry_2_), .S(npu_inst_pe_1_2_7_N74) );
  NAND3_X1 npu_inst_pe_1_2_7_U109 ( .A1(npu_inst_pe_1_2_7_n5), .A2(
        npu_inst_pe_1_2_7_n7), .A3(npu_inst_pe_1_2_7_n8), .ZN(
        npu_inst_pe_1_2_7_n44) );
  NAND3_X1 npu_inst_pe_1_2_7_U108 ( .A1(npu_inst_pe_1_2_7_n4), .A2(
        npu_inst_pe_1_2_7_n7), .A3(npu_inst_pe_1_2_7_n8), .ZN(
        npu_inst_pe_1_2_7_n40) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_2_7_n34), .CK(
        npu_inst_pe_1_2_7_net3764), .RN(npu_inst_pe_1_2_7_n9), .Q(
        npu_inst_pe_1_2_7_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_2_7_n35), .CK(
        npu_inst_pe_1_2_7_net3764), .RN(npu_inst_pe_1_2_7_n9), .Q(
        npu_inst_pe_1_2_7_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_2_7_n36), .CK(
        npu_inst_pe_1_2_7_net3764), .RN(npu_inst_pe_1_2_7_n9), .Q(
        npu_inst_pe_1_2_7_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_2_7_n98), .CK(
        npu_inst_pe_1_2_7_net3764), .RN(npu_inst_pe_1_2_7_n9), .Q(
        npu_inst_pe_1_2_7_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_2_7_n99), .CK(
        npu_inst_pe_1_2_7_net3764), .RN(npu_inst_pe_1_2_7_n9), .Q(
        npu_inst_pe_1_2_7_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_2_7_n100), 
        .CK(npu_inst_pe_1_2_7_net3764), .RN(npu_inst_pe_1_2_7_n9), .Q(
        npu_inst_pe_1_2_7_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_2_7_n33), .CK(
        npu_inst_pe_1_2_7_net3764), .RN(npu_inst_pe_1_2_7_n9), .Q(
        npu_inst_pe_1_2_7_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_2_7_n101), 
        .CK(npu_inst_pe_1_2_7_net3764), .RN(npu_inst_pe_1_2_7_n9), .Q(
        npu_inst_pe_1_2_7_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_weight_reg_0_ ( .D(npu_inst_n111), .CK(
        npu_inst_pe_1_2_7_net3770), .RN(npu_inst_pe_1_2_7_n9), .Q(
        npu_inst_pe_1_2_7_int_q_weight_0_), .QN(npu_inst_pe_1_2_7_n27) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_weight_reg_1_ ( .D(npu_inst_n117), .CK(
        npu_inst_pe_1_2_7_net3770), .RN(npu_inst_pe_1_2_7_n9), .Q(
        npu_inst_pe_1_2_7_int_q_weight_1_), .QN(npu_inst_pe_1_2_7_n26) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_2_7_n113), 
        .CK(npu_inst_pe_1_2_7_net3770), .RN(npu_inst_pe_1_2_7_n9), .Q(
        npu_inst_pe_1_2_7_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_2_7_n107), 
        .CK(npu_inst_pe_1_2_7_net3770), .RN(npu_inst_pe_1_2_7_n9), .Q(
        npu_inst_pe_1_2_7_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_2_7_n112), 
        .CK(npu_inst_pe_1_2_7_net3770), .RN(npu_inst_pe_1_2_7_n10), .Q(
        npu_inst_pe_1_2_7_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_2_7_n106), 
        .CK(npu_inst_pe_1_2_7_net3770), .RN(npu_inst_pe_1_2_7_n10), .Q(
        npu_inst_pe_1_2_7_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_2_7_n111), 
        .CK(npu_inst_pe_1_2_7_net3770), .RN(npu_inst_pe_1_2_7_n10), .Q(
        npu_inst_pe_1_2_7_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_2_7_n105), 
        .CK(npu_inst_pe_1_2_7_net3770), .RN(npu_inst_pe_1_2_7_n10), .Q(
        npu_inst_pe_1_2_7_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_2_7_n110), 
        .CK(npu_inst_pe_1_2_7_net3770), .RN(npu_inst_pe_1_2_7_n10), .Q(
        npu_inst_pe_1_2_7_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_2_7_n104), 
        .CK(npu_inst_pe_1_2_7_net3770), .RN(npu_inst_pe_1_2_7_n10), .Q(
        npu_inst_pe_1_2_7_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_2_7_n109), 
        .CK(npu_inst_pe_1_2_7_net3770), .RN(npu_inst_pe_1_2_7_n10), .Q(
        npu_inst_pe_1_2_7_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_2_7_n103), 
        .CK(npu_inst_pe_1_2_7_net3770), .RN(npu_inst_pe_1_2_7_n10), .Q(
        npu_inst_pe_1_2_7_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_2_7_n108), 
        .CK(npu_inst_pe_1_2_7_net3770), .RN(npu_inst_pe_1_2_7_n10), .Q(
        npu_inst_pe_1_2_7_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_2_7_n102), 
        .CK(npu_inst_pe_1_2_7_net3770), .RN(npu_inst_pe_1_2_7_n10), .Q(
        npu_inst_pe_1_2_7_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_2_7_n86), 
        .CK(npu_inst_pe_1_2_7_net3770), .RN(npu_inst_pe_1_2_7_n10), .Q(
        npu_inst_pe_1_2_7_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_2_7_n87), 
        .CK(npu_inst_pe_1_2_7_net3770), .RN(npu_inst_pe_1_2_7_n10), .Q(
        npu_inst_pe_1_2_7_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_2_7_n88), 
        .CK(npu_inst_pe_1_2_7_net3770), .RN(npu_inst_pe_1_2_7_n11), .Q(
        npu_inst_pe_1_2_7_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_2_7_n89), 
        .CK(npu_inst_pe_1_2_7_net3770), .RN(npu_inst_pe_1_2_7_n11), .Q(
        npu_inst_pe_1_2_7_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_2_7_n90), 
        .CK(npu_inst_pe_1_2_7_net3770), .RN(npu_inst_pe_1_2_7_n11), .Q(
        npu_inst_pe_1_2_7_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_2_7_n91), 
        .CK(npu_inst_pe_1_2_7_net3770), .RN(npu_inst_pe_1_2_7_n11), .Q(
        npu_inst_pe_1_2_7_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_2_7_n92), 
        .CK(npu_inst_pe_1_2_7_net3770), .RN(npu_inst_pe_1_2_7_n11), .Q(
        npu_inst_pe_1_2_7_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_2_7_n93), 
        .CK(npu_inst_pe_1_2_7_net3770), .RN(npu_inst_pe_1_2_7_n11), .Q(
        npu_inst_pe_1_2_7_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_2_7_n94), 
        .CK(npu_inst_pe_1_2_7_net3770), .RN(npu_inst_pe_1_2_7_n11), .Q(
        npu_inst_pe_1_2_7_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_2_7_n95), 
        .CK(npu_inst_pe_1_2_7_net3770), .RN(npu_inst_pe_1_2_7_n11), .Q(
        npu_inst_pe_1_2_7_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_2_7_n96), 
        .CK(npu_inst_pe_1_2_7_net3770), .RN(npu_inst_pe_1_2_7_n11), .Q(
        npu_inst_pe_1_2_7_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_2_7_n97), 
        .CK(npu_inst_pe_1_2_7_net3770), .RN(npu_inst_pe_1_2_7_n11), .Q(
        npu_inst_pe_1_2_7_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_2_7_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_2_7_N84), .SE(1'b0), .GCK(npu_inst_pe_1_2_7_net3764) );
  CLKGATETST_X1 npu_inst_pe_1_2_7_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n64), .SE(1'b0), .GCK(npu_inst_pe_1_2_7_net3770) );
  MUX2_X1 npu_inst_pe_1_3_0_U162 ( .A(npu_inst_pe_1_3_0_n32), .B(
        npu_inst_pe_1_3_0_n29), .S(npu_inst_pe_1_3_0_n8), .Z(
        npu_inst_pe_1_3_0_N93) );
  MUX2_X1 npu_inst_pe_1_3_0_U161 ( .A(npu_inst_pe_1_3_0_n31), .B(
        npu_inst_pe_1_3_0_n30), .S(npu_inst_pe_1_3_0_n6), .Z(
        npu_inst_pe_1_3_0_n32) );
  MUX2_X1 npu_inst_pe_1_3_0_U160 ( .A(npu_inst_pe_1_3_0_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_3_0_int_q_reg_v_1__0_), .S(npu_inst_pe_1_3_0_n4), .Z(
        npu_inst_pe_1_3_0_n31) );
  MUX2_X1 npu_inst_pe_1_3_0_U159 ( .A(npu_inst_pe_1_3_0_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_3_0_int_q_reg_v_3__0_), .S(npu_inst_pe_1_3_0_n4), .Z(
        npu_inst_pe_1_3_0_n30) );
  MUX2_X1 npu_inst_pe_1_3_0_U158 ( .A(npu_inst_pe_1_3_0_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_3_0_int_q_reg_v_5__0_), .S(npu_inst_pe_1_3_0_n4), .Z(
        npu_inst_pe_1_3_0_n29) );
  MUX2_X1 npu_inst_pe_1_3_0_U157 ( .A(npu_inst_pe_1_3_0_n28), .B(
        npu_inst_pe_1_3_0_n23), .S(npu_inst_pe_1_3_0_n8), .Z(
        npu_inst_pe_1_3_0_N94) );
  MUX2_X1 npu_inst_pe_1_3_0_U156 ( .A(npu_inst_pe_1_3_0_n25), .B(
        npu_inst_pe_1_3_0_n24), .S(npu_inst_pe_1_3_0_n6), .Z(
        npu_inst_pe_1_3_0_n28) );
  MUX2_X1 npu_inst_pe_1_3_0_U155 ( .A(npu_inst_pe_1_3_0_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_3_0_int_q_reg_v_1__1_), .S(npu_inst_pe_1_3_0_n4), .Z(
        npu_inst_pe_1_3_0_n25) );
  MUX2_X1 npu_inst_pe_1_3_0_U154 ( .A(npu_inst_pe_1_3_0_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_3_0_int_q_reg_v_3__1_), .S(npu_inst_pe_1_3_0_n4), .Z(
        npu_inst_pe_1_3_0_n24) );
  MUX2_X1 npu_inst_pe_1_3_0_U153 ( .A(npu_inst_pe_1_3_0_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_3_0_int_q_reg_v_5__1_), .S(npu_inst_pe_1_3_0_n4), .Z(
        npu_inst_pe_1_3_0_n23) );
  MUX2_X1 npu_inst_pe_1_3_0_U152 ( .A(npu_inst_pe_1_3_0_n22), .B(
        npu_inst_pe_1_3_0_n19), .S(npu_inst_pe_1_3_0_n8), .Z(
        npu_inst_pe_1_3_0_o_data_h_1_) );
  MUX2_X1 npu_inst_pe_1_3_0_U151 ( .A(npu_inst_pe_1_3_0_n21), .B(
        npu_inst_pe_1_3_0_n20), .S(npu_inst_pe_1_3_0_n6), .Z(
        npu_inst_pe_1_3_0_n22) );
  MUX2_X1 npu_inst_pe_1_3_0_U150 ( .A(npu_inst_pe_1_3_0_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_3_0_int_q_reg_h_1__1_), .S(npu_inst_pe_1_3_0_n4), .Z(
        npu_inst_pe_1_3_0_n21) );
  MUX2_X1 npu_inst_pe_1_3_0_U149 ( .A(npu_inst_pe_1_3_0_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_3_0_int_q_reg_h_3__1_), .S(npu_inst_pe_1_3_0_n4), .Z(
        npu_inst_pe_1_3_0_n20) );
  MUX2_X1 npu_inst_pe_1_3_0_U148 ( .A(npu_inst_pe_1_3_0_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_3_0_int_q_reg_h_5__1_), .S(npu_inst_pe_1_3_0_n4), .Z(
        npu_inst_pe_1_3_0_n19) );
  MUX2_X1 npu_inst_pe_1_3_0_U147 ( .A(npu_inst_pe_1_3_0_n18), .B(
        npu_inst_pe_1_3_0_n15), .S(npu_inst_pe_1_3_0_n8), .Z(
        npu_inst_pe_1_3_0_o_data_h_0_) );
  MUX2_X1 npu_inst_pe_1_3_0_U146 ( .A(npu_inst_pe_1_3_0_n17), .B(
        npu_inst_pe_1_3_0_n16), .S(npu_inst_pe_1_3_0_n6), .Z(
        npu_inst_pe_1_3_0_n18) );
  MUX2_X1 npu_inst_pe_1_3_0_U145 ( .A(npu_inst_pe_1_3_0_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_3_0_int_q_reg_h_1__0_), .S(npu_inst_pe_1_3_0_n4), .Z(
        npu_inst_pe_1_3_0_n17) );
  MUX2_X1 npu_inst_pe_1_3_0_U144 ( .A(npu_inst_pe_1_3_0_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_3_0_int_q_reg_h_3__0_), .S(npu_inst_pe_1_3_0_n4), .Z(
        npu_inst_pe_1_3_0_n16) );
  MUX2_X1 npu_inst_pe_1_3_0_U143 ( .A(npu_inst_pe_1_3_0_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_3_0_int_q_reg_h_5__0_), .S(npu_inst_pe_1_3_0_n4), .Z(
        npu_inst_pe_1_3_0_n15) );
  XOR2_X1 npu_inst_pe_1_3_0_U142 ( .A(npu_inst_pe_1_3_0_int_data_0_), .B(
        npu_inst_pe_1_3_0_int_q_acc_0_), .Z(npu_inst_pe_1_3_0_N73) );
  AND2_X1 npu_inst_pe_1_3_0_U141 ( .A1(npu_inst_pe_1_3_0_int_q_acc_0_), .A2(
        npu_inst_pe_1_3_0_int_data_0_), .ZN(npu_inst_pe_1_3_0_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_3_0_U140 ( .A(npu_inst_pe_1_3_0_int_q_acc_0_), .B(
        npu_inst_pe_1_3_0_n13), .ZN(npu_inst_pe_1_3_0_N65) );
  OR2_X1 npu_inst_pe_1_3_0_U139 ( .A1(npu_inst_pe_1_3_0_n13), .A2(
        npu_inst_pe_1_3_0_int_q_acc_0_), .ZN(npu_inst_pe_1_3_0_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_3_0_U138 ( .A(npu_inst_pe_1_3_0_int_q_acc_2_), .B(
        npu_inst_pe_1_3_0_add_79_carry_2_), .Z(npu_inst_pe_1_3_0_N75) );
  AND2_X1 npu_inst_pe_1_3_0_U137 ( .A1(npu_inst_pe_1_3_0_add_79_carry_2_), 
        .A2(npu_inst_pe_1_3_0_int_q_acc_2_), .ZN(
        npu_inst_pe_1_3_0_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_3_0_U136 ( .A(npu_inst_pe_1_3_0_int_q_acc_3_), .B(
        npu_inst_pe_1_3_0_add_79_carry_3_), .Z(npu_inst_pe_1_3_0_N76) );
  AND2_X1 npu_inst_pe_1_3_0_U135 ( .A1(npu_inst_pe_1_3_0_add_79_carry_3_), 
        .A2(npu_inst_pe_1_3_0_int_q_acc_3_), .ZN(
        npu_inst_pe_1_3_0_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_3_0_U134 ( .A(npu_inst_pe_1_3_0_int_q_acc_4_), .B(
        npu_inst_pe_1_3_0_add_79_carry_4_), .Z(npu_inst_pe_1_3_0_N77) );
  AND2_X1 npu_inst_pe_1_3_0_U133 ( .A1(npu_inst_pe_1_3_0_add_79_carry_4_), 
        .A2(npu_inst_pe_1_3_0_int_q_acc_4_), .ZN(
        npu_inst_pe_1_3_0_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_3_0_U132 ( .A(npu_inst_pe_1_3_0_int_q_acc_5_), .B(
        npu_inst_pe_1_3_0_add_79_carry_5_), .Z(npu_inst_pe_1_3_0_N78) );
  AND2_X1 npu_inst_pe_1_3_0_U131 ( .A1(npu_inst_pe_1_3_0_add_79_carry_5_), 
        .A2(npu_inst_pe_1_3_0_int_q_acc_5_), .ZN(
        npu_inst_pe_1_3_0_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_3_0_U130 ( .A(npu_inst_pe_1_3_0_int_q_acc_6_), .B(
        npu_inst_pe_1_3_0_add_79_carry_6_), .Z(npu_inst_pe_1_3_0_N79) );
  AND2_X1 npu_inst_pe_1_3_0_U129 ( .A1(npu_inst_pe_1_3_0_add_79_carry_6_), 
        .A2(npu_inst_pe_1_3_0_int_q_acc_6_), .ZN(
        npu_inst_pe_1_3_0_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_3_0_U128 ( .A(npu_inst_pe_1_3_0_int_q_acc_7_), .B(
        npu_inst_pe_1_3_0_add_79_carry_7_), .Z(npu_inst_pe_1_3_0_N80) );
  XNOR2_X1 npu_inst_pe_1_3_0_U127 ( .A(npu_inst_pe_1_3_0_sub_77_carry_2_), .B(
        npu_inst_pe_1_3_0_int_q_acc_2_), .ZN(npu_inst_pe_1_3_0_N67) );
  OR2_X1 npu_inst_pe_1_3_0_U126 ( .A1(npu_inst_pe_1_3_0_int_q_acc_2_), .A2(
        npu_inst_pe_1_3_0_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_3_0_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_3_0_U125 ( .A(npu_inst_pe_1_3_0_sub_77_carry_3_), .B(
        npu_inst_pe_1_3_0_int_q_acc_3_), .ZN(npu_inst_pe_1_3_0_N68) );
  OR2_X1 npu_inst_pe_1_3_0_U124 ( .A1(npu_inst_pe_1_3_0_int_q_acc_3_), .A2(
        npu_inst_pe_1_3_0_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_3_0_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_3_0_U123 ( .A(npu_inst_pe_1_3_0_sub_77_carry_4_), .B(
        npu_inst_pe_1_3_0_int_q_acc_4_), .ZN(npu_inst_pe_1_3_0_N69) );
  OR2_X1 npu_inst_pe_1_3_0_U122 ( .A1(npu_inst_pe_1_3_0_int_q_acc_4_), .A2(
        npu_inst_pe_1_3_0_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_3_0_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_3_0_U121 ( .A(npu_inst_pe_1_3_0_sub_77_carry_5_), .B(
        npu_inst_pe_1_3_0_int_q_acc_5_), .ZN(npu_inst_pe_1_3_0_N70) );
  OR2_X1 npu_inst_pe_1_3_0_U120 ( .A1(npu_inst_pe_1_3_0_int_q_acc_5_), .A2(
        npu_inst_pe_1_3_0_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_3_0_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_3_0_U119 ( .A(npu_inst_pe_1_3_0_sub_77_carry_6_), .B(
        npu_inst_pe_1_3_0_int_q_acc_6_), .ZN(npu_inst_pe_1_3_0_N71) );
  OR2_X1 npu_inst_pe_1_3_0_U118 ( .A1(npu_inst_pe_1_3_0_int_q_acc_6_), .A2(
        npu_inst_pe_1_3_0_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_3_0_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_3_0_U117 ( .A(npu_inst_pe_1_3_0_int_q_acc_7_), .B(
        npu_inst_pe_1_3_0_sub_77_carry_7_), .ZN(npu_inst_pe_1_3_0_N72) );
  INV_X1 npu_inst_pe_1_3_0_U116 ( .A(npu_inst_n78), .ZN(npu_inst_pe_1_3_0_n7)
         );
  INV_X1 npu_inst_pe_1_3_0_U115 ( .A(npu_inst_pe_1_3_0_n7), .ZN(
        npu_inst_pe_1_3_0_n6) );
  INV_X1 npu_inst_pe_1_3_0_U114 ( .A(npu_inst_n57), .ZN(npu_inst_pe_1_3_0_n3)
         );
  AOI22_X1 npu_inst_pe_1_3_0_U113 ( .A1(npu_inst_int_data_y_4__0__0_), .A2(
        npu_inst_pe_1_3_0_n58), .B1(npu_inst_pe_1_3_0_n114), .B2(
        npu_inst_pe_1_3_0_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_3_0_n57) );
  INV_X1 npu_inst_pe_1_3_0_U112 ( .A(npu_inst_pe_1_3_0_n57), .ZN(
        npu_inst_pe_1_3_0_n108) );
  AOI22_X1 npu_inst_pe_1_3_0_U111 ( .A1(npu_inst_int_data_y_4__0__0_), .A2(
        npu_inst_pe_1_3_0_n54), .B1(npu_inst_pe_1_3_0_n115), .B2(
        npu_inst_pe_1_3_0_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_3_0_n53) );
  INV_X1 npu_inst_pe_1_3_0_U110 ( .A(npu_inst_pe_1_3_0_n53), .ZN(
        npu_inst_pe_1_3_0_n109) );
  AOI22_X1 npu_inst_pe_1_3_0_U107 ( .A1(npu_inst_int_data_y_4__0__0_), .A2(
        npu_inst_pe_1_3_0_n50), .B1(npu_inst_pe_1_3_0_n116), .B2(
        npu_inst_pe_1_3_0_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_3_0_n49) );
  INV_X1 npu_inst_pe_1_3_0_U106 ( .A(npu_inst_pe_1_3_0_n49), .ZN(
        npu_inst_pe_1_3_0_n110) );
  AOI22_X1 npu_inst_pe_1_3_0_U105 ( .A1(npu_inst_int_data_y_4__0__0_), .A2(
        npu_inst_pe_1_3_0_n46), .B1(npu_inst_pe_1_3_0_n117), .B2(
        npu_inst_pe_1_3_0_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_3_0_n45) );
  INV_X1 npu_inst_pe_1_3_0_U104 ( .A(npu_inst_pe_1_3_0_n45), .ZN(
        npu_inst_pe_1_3_0_n111) );
  AOI22_X1 npu_inst_pe_1_3_0_U103 ( .A1(npu_inst_int_data_y_4__0__0_), .A2(
        npu_inst_pe_1_3_0_n42), .B1(npu_inst_pe_1_3_0_n119), .B2(
        npu_inst_pe_1_3_0_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_3_0_n41) );
  INV_X1 npu_inst_pe_1_3_0_U102 ( .A(npu_inst_pe_1_3_0_n41), .ZN(
        npu_inst_pe_1_3_0_n112) );
  AOI22_X1 npu_inst_pe_1_3_0_U101 ( .A1(npu_inst_int_data_y_4__0__1_), .A2(
        npu_inst_pe_1_3_0_n58), .B1(npu_inst_pe_1_3_0_n114), .B2(
        npu_inst_pe_1_3_0_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_3_0_n59) );
  INV_X1 npu_inst_pe_1_3_0_U100 ( .A(npu_inst_pe_1_3_0_n59), .ZN(
        npu_inst_pe_1_3_0_n102) );
  AOI22_X1 npu_inst_pe_1_3_0_U99 ( .A1(npu_inst_int_data_y_4__0__1_), .A2(
        npu_inst_pe_1_3_0_n54), .B1(npu_inst_pe_1_3_0_n115), .B2(
        npu_inst_pe_1_3_0_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_3_0_n55) );
  INV_X1 npu_inst_pe_1_3_0_U98 ( .A(npu_inst_pe_1_3_0_n55), .ZN(
        npu_inst_pe_1_3_0_n103) );
  AOI22_X1 npu_inst_pe_1_3_0_U97 ( .A1(npu_inst_int_data_y_4__0__1_), .A2(
        npu_inst_pe_1_3_0_n50), .B1(npu_inst_pe_1_3_0_n116), .B2(
        npu_inst_pe_1_3_0_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_3_0_n51) );
  INV_X1 npu_inst_pe_1_3_0_U96 ( .A(npu_inst_pe_1_3_0_n51), .ZN(
        npu_inst_pe_1_3_0_n104) );
  AOI22_X1 npu_inst_pe_1_3_0_U95 ( .A1(npu_inst_int_data_y_4__0__1_), .A2(
        npu_inst_pe_1_3_0_n46), .B1(npu_inst_pe_1_3_0_n117), .B2(
        npu_inst_pe_1_3_0_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_3_0_n47) );
  INV_X1 npu_inst_pe_1_3_0_U94 ( .A(npu_inst_pe_1_3_0_n47), .ZN(
        npu_inst_pe_1_3_0_n105) );
  AOI22_X1 npu_inst_pe_1_3_0_U93 ( .A1(npu_inst_int_data_y_4__0__1_), .A2(
        npu_inst_pe_1_3_0_n42), .B1(npu_inst_pe_1_3_0_n119), .B2(
        npu_inst_pe_1_3_0_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_3_0_n43) );
  INV_X1 npu_inst_pe_1_3_0_U92 ( .A(npu_inst_pe_1_3_0_n43), .ZN(
        npu_inst_pe_1_3_0_n106) );
  AOI22_X1 npu_inst_pe_1_3_0_U91 ( .A1(npu_inst_pe_1_3_0_n38), .A2(
        npu_inst_int_data_y_4__0__1_), .B1(npu_inst_pe_1_3_0_n118), .B2(
        npu_inst_pe_1_3_0_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_3_0_n39) );
  INV_X1 npu_inst_pe_1_3_0_U90 ( .A(npu_inst_pe_1_3_0_n39), .ZN(
        npu_inst_pe_1_3_0_n107) );
  AOI22_X1 npu_inst_pe_1_3_0_U89 ( .A1(npu_inst_pe_1_3_0_n38), .A2(
        npu_inst_int_data_y_4__0__0_), .B1(npu_inst_pe_1_3_0_n118), .B2(
        npu_inst_pe_1_3_0_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_3_0_n37) );
  INV_X1 npu_inst_pe_1_3_0_U88 ( .A(npu_inst_pe_1_3_0_n37), .ZN(
        npu_inst_pe_1_3_0_n113) );
  NAND2_X1 npu_inst_pe_1_3_0_U87 ( .A1(npu_inst_pe_1_3_0_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_3_0_n60), .ZN(npu_inst_pe_1_3_0_n74) );
  OAI21_X1 npu_inst_pe_1_3_0_U86 ( .B1(npu_inst_pe_1_3_0_n63), .B2(
        npu_inst_pe_1_3_0_n60), .A(npu_inst_pe_1_3_0_n74), .ZN(
        npu_inst_pe_1_3_0_n97) );
  NAND2_X1 npu_inst_pe_1_3_0_U85 ( .A1(npu_inst_pe_1_3_0_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_3_0_n60), .ZN(npu_inst_pe_1_3_0_n73) );
  OAI21_X1 npu_inst_pe_1_3_0_U84 ( .B1(npu_inst_pe_1_3_0_n61), .B2(
        npu_inst_pe_1_3_0_n60), .A(npu_inst_pe_1_3_0_n73), .ZN(
        npu_inst_pe_1_3_0_n96) );
  NAND2_X1 npu_inst_pe_1_3_0_U83 ( .A1(npu_inst_pe_1_3_0_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_3_0_n56), .ZN(npu_inst_pe_1_3_0_n72) );
  OAI21_X1 npu_inst_pe_1_3_0_U82 ( .B1(npu_inst_pe_1_3_0_n63), .B2(
        npu_inst_pe_1_3_0_n56), .A(npu_inst_pe_1_3_0_n72), .ZN(
        npu_inst_pe_1_3_0_n95) );
  NAND2_X1 npu_inst_pe_1_3_0_U81 ( .A1(npu_inst_pe_1_3_0_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_3_0_n56), .ZN(npu_inst_pe_1_3_0_n71) );
  OAI21_X1 npu_inst_pe_1_3_0_U80 ( .B1(npu_inst_pe_1_3_0_n61), .B2(
        npu_inst_pe_1_3_0_n56), .A(npu_inst_pe_1_3_0_n71), .ZN(
        npu_inst_pe_1_3_0_n94) );
  NAND2_X1 npu_inst_pe_1_3_0_U79 ( .A1(npu_inst_pe_1_3_0_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_3_0_n52), .ZN(npu_inst_pe_1_3_0_n70) );
  OAI21_X1 npu_inst_pe_1_3_0_U78 ( .B1(npu_inst_pe_1_3_0_n63), .B2(
        npu_inst_pe_1_3_0_n52), .A(npu_inst_pe_1_3_0_n70), .ZN(
        npu_inst_pe_1_3_0_n93) );
  NAND2_X1 npu_inst_pe_1_3_0_U77 ( .A1(npu_inst_pe_1_3_0_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_3_0_n52), .ZN(npu_inst_pe_1_3_0_n69) );
  OAI21_X1 npu_inst_pe_1_3_0_U76 ( .B1(npu_inst_pe_1_3_0_n61), .B2(
        npu_inst_pe_1_3_0_n52), .A(npu_inst_pe_1_3_0_n69), .ZN(
        npu_inst_pe_1_3_0_n92) );
  NAND2_X1 npu_inst_pe_1_3_0_U75 ( .A1(npu_inst_pe_1_3_0_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_3_0_n48), .ZN(npu_inst_pe_1_3_0_n68) );
  OAI21_X1 npu_inst_pe_1_3_0_U74 ( .B1(npu_inst_pe_1_3_0_n63), .B2(
        npu_inst_pe_1_3_0_n48), .A(npu_inst_pe_1_3_0_n68), .ZN(
        npu_inst_pe_1_3_0_n91) );
  NAND2_X1 npu_inst_pe_1_3_0_U73 ( .A1(npu_inst_pe_1_3_0_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_3_0_n48), .ZN(npu_inst_pe_1_3_0_n67) );
  OAI21_X1 npu_inst_pe_1_3_0_U72 ( .B1(npu_inst_pe_1_3_0_n61), .B2(
        npu_inst_pe_1_3_0_n48), .A(npu_inst_pe_1_3_0_n67), .ZN(
        npu_inst_pe_1_3_0_n90) );
  NAND2_X1 npu_inst_pe_1_3_0_U71 ( .A1(npu_inst_pe_1_3_0_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_3_0_n44), .ZN(npu_inst_pe_1_3_0_n66) );
  OAI21_X1 npu_inst_pe_1_3_0_U70 ( .B1(npu_inst_pe_1_3_0_n63), .B2(
        npu_inst_pe_1_3_0_n44), .A(npu_inst_pe_1_3_0_n66), .ZN(
        npu_inst_pe_1_3_0_n89) );
  NAND2_X1 npu_inst_pe_1_3_0_U69 ( .A1(npu_inst_pe_1_3_0_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_3_0_n44), .ZN(npu_inst_pe_1_3_0_n65) );
  OAI21_X1 npu_inst_pe_1_3_0_U68 ( .B1(npu_inst_pe_1_3_0_n61), .B2(
        npu_inst_pe_1_3_0_n44), .A(npu_inst_pe_1_3_0_n65), .ZN(
        npu_inst_pe_1_3_0_n88) );
  NAND2_X1 npu_inst_pe_1_3_0_U67 ( .A1(npu_inst_pe_1_3_0_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_3_0_n40), .ZN(npu_inst_pe_1_3_0_n64) );
  OAI21_X1 npu_inst_pe_1_3_0_U66 ( .B1(npu_inst_pe_1_3_0_n63), .B2(
        npu_inst_pe_1_3_0_n40), .A(npu_inst_pe_1_3_0_n64), .ZN(
        npu_inst_pe_1_3_0_n87) );
  NAND2_X1 npu_inst_pe_1_3_0_U65 ( .A1(npu_inst_pe_1_3_0_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_3_0_n40), .ZN(npu_inst_pe_1_3_0_n62) );
  OAI21_X1 npu_inst_pe_1_3_0_U64 ( .B1(npu_inst_pe_1_3_0_n61), .B2(
        npu_inst_pe_1_3_0_n40), .A(npu_inst_pe_1_3_0_n62), .ZN(
        npu_inst_pe_1_3_0_n86) );
  AND2_X1 npu_inst_pe_1_3_0_U63 ( .A1(npu_inst_pe_1_3_0_N93), .A2(npu_inst_n57), .ZN(npu_inst_int_data_y_3__0__0_) );
  AND2_X1 npu_inst_pe_1_3_0_U62 ( .A1(npu_inst_n57), .A2(npu_inst_pe_1_3_0_N94), .ZN(npu_inst_int_data_y_3__0__1_) );
  NOR3_X1 npu_inst_pe_1_3_0_U61 ( .A1(npu_inst_pe_1_3_0_n26), .A2(npu_inst_n57), .A3(npu_inst_int_ckg[39]), .ZN(npu_inst_pe_1_3_0_n85) );
  OR2_X1 npu_inst_pe_1_3_0_U60 ( .A1(npu_inst_pe_1_3_0_n85), .A2(
        npu_inst_pe_1_3_0_n2), .ZN(npu_inst_pe_1_3_0_N84) );
  AND2_X1 npu_inst_pe_1_3_0_U59 ( .A1(npu_inst_pe_1_3_0_int_q_acc_0_), .A2(
        npu_inst_pe_1_3_0_n1), .ZN(npu_inst_int_data_res_3__0__0_) );
  AND2_X1 npu_inst_pe_1_3_0_U58 ( .A1(npu_inst_pe_1_3_0_n2), .A2(
        npu_inst_pe_1_3_0_int_q_acc_7_), .ZN(npu_inst_int_data_res_3__0__7_)
         );
  AND2_X1 npu_inst_pe_1_3_0_U57 ( .A1(npu_inst_pe_1_3_0_int_q_acc_1_), .A2(
        npu_inst_pe_1_3_0_n1), .ZN(npu_inst_int_data_res_3__0__1_) );
  AND2_X1 npu_inst_pe_1_3_0_U56 ( .A1(npu_inst_pe_1_3_0_int_q_acc_2_), .A2(
        npu_inst_pe_1_3_0_n1), .ZN(npu_inst_int_data_res_3__0__2_) );
  AND2_X1 npu_inst_pe_1_3_0_U55 ( .A1(npu_inst_pe_1_3_0_int_q_acc_3_), .A2(
        npu_inst_pe_1_3_0_n2), .ZN(npu_inst_int_data_res_3__0__3_) );
  AND2_X1 npu_inst_pe_1_3_0_U54 ( .A1(npu_inst_pe_1_3_0_int_q_acc_4_), .A2(
        npu_inst_pe_1_3_0_n2), .ZN(npu_inst_int_data_res_3__0__4_) );
  AND2_X1 npu_inst_pe_1_3_0_U53 ( .A1(npu_inst_pe_1_3_0_int_q_acc_5_), .A2(
        npu_inst_pe_1_3_0_n2), .ZN(npu_inst_int_data_res_3__0__5_) );
  AND2_X1 npu_inst_pe_1_3_0_U52 ( .A1(npu_inst_pe_1_3_0_int_q_acc_6_), .A2(
        npu_inst_pe_1_3_0_n2), .ZN(npu_inst_int_data_res_3__0__6_) );
  AOI222_X1 npu_inst_pe_1_3_0_U51 ( .A1(npu_inst_int_data_res_4__0__0_), .A2(
        npu_inst_pe_1_3_0_n1), .B1(npu_inst_pe_1_3_0_N73), .B2(
        npu_inst_pe_1_3_0_n76), .C1(npu_inst_pe_1_3_0_N65), .C2(
        npu_inst_pe_1_3_0_n77), .ZN(npu_inst_pe_1_3_0_n84) );
  INV_X1 npu_inst_pe_1_3_0_U50 ( .A(npu_inst_pe_1_3_0_n84), .ZN(
        npu_inst_pe_1_3_0_n101) );
  AOI222_X1 npu_inst_pe_1_3_0_U49 ( .A1(npu_inst_int_data_res_4__0__7_), .A2(
        npu_inst_pe_1_3_0_n1), .B1(npu_inst_pe_1_3_0_N80), .B2(
        npu_inst_pe_1_3_0_n76), .C1(npu_inst_pe_1_3_0_N72), .C2(
        npu_inst_pe_1_3_0_n77), .ZN(npu_inst_pe_1_3_0_n75) );
  INV_X1 npu_inst_pe_1_3_0_U48 ( .A(npu_inst_pe_1_3_0_n75), .ZN(
        npu_inst_pe_1_3_0_n33) );
  AOI222_X1 npu_inst_pe_1_3_0_U47 ( .A1(npu_inst_int_data_res_4__0__1_), .A2(
        npu_inst_pe_1_3_0_n1), .B1(npu_inst_pe_1_3_0_N74), .B2(
        npu_inst_pe_1_3_0_n76), .C1(npu_inst_pe_1_3_0_N66), .C2(
        npu_inst_pe_1_3_0_n77), .ZN(npu_inst_pe_1_3_0_n83) );
  INV_X1 npu_inst_pe_1_3_0_U46 ( .A(npu_inst_pe_1_3_0_n83), .ZN(
        npu_inst_pe_1_3_0_n100) );
  AOI222_X1 npu_inst_pe_1_3_0_U45 ( .A1(npu_inst_int_data_res_4__0__2_), .A2(
        npu_inst_pe_1_3_0_n1), .B1(npu_inst_pe_1_3_0_N75), .B2(
        npu_inst_pe_1_3_0_n76), .C1(npu_inst_pe_1_3_0_N67), .C2(
        npu_inst_pe_1_3_0_n77), .ZN(npu_inst_pe_1_3_0_n82) );
  INV_X1 npu_inst_pe_1_3_0_U44 ( .A(npu_inst_pe_1_3_0_n82), .ZN(
        npu_inst_pe_1_3_0_n99) );
  AOI222_X1 npu_inst_pe_1_3_0_U43 ( .A1(npu_inst_int_data_res_4__0__3_), .A2(
        npu_inst_pe_1_3_0_n1), .B1(npu_inst_pe_1_3_0_N76), .B2(
        npu_inst_pe_1_3_0_n76), .C1(npu_inst_pe_1_3_0_N68), .C2(
        npu_inst_pe_1_3_0_n77), .ZN(npu_inst_pe_1_3_0_n81) );
  INV_X1 npu_inst_pe_1_3_0_U42 ( .A(npu_inst_pe_1_3_0_n81), .ZN(
        npu_inst_pe_1_3_0_n98) );
  AOI222_X1 npu_inst_pe_1_3_0_U41 ( .A1(npu_inst_int_data_res_4__0__4_), .A2(
        npu_inst_pe_1_3_0_n1), .B1(npu_inst_pe_1_3_0_N77), .B2(
        npu_inst_pe_1_3_0_n76), .C1(npu_inst_pe_1_3_0_N69), .C2(
        npu_inst_pe_1_3_0_n77), .ZN(npu_inst_pe_1_3_0_n80) );
  INV_X1 npu_inst_pe_1_3_0_U40 ( .A(npu_inst_pe_1_3_0_n80), .ZN(
        npu_inst_pe_1_3_0_n36) );
  AOI222_X1 npu_inst_pe_1_3_0_U39 ( .A1(npu_inst_int_data_res_4__0__5_), .A2(
        npu_inst_pe_1_3_0_n1), .B1(npu_inst_pe_1_3_0_N78), .B2(
        npu_inst_pe_1_3_0_n76), .C1(npu_inst_pe_1_3_0_N70), .C2(
        npu_inst_pe_1_3_0_n77), .ZN(npu_inst_pe_1_3_0_n79) );
  INV_X1 npu_inst_pe_1_3_0_U38 ( .A(npu_inst_pe_1_3_0_n79), .ZN(
        npu_inst_pe_1_3_0_n35) );
  AOI222_X1 npu_inst_pe_1_3_0_U37 ( .A1(npu_inst_int_data_res_4__0__6_), .A2(
        npu_inst_pe_1_3_0_n1), .B1(npu_inst_pe_1_3_0_N79), .B2(
        npu_inst_pe_1_3_0_n76), .C1(npu_inst_pe_1_3_0_N71), .C2(
        npu_inst_pe_1_3_0_n77), .ZN(npu_inst_pe_1_3_0_n78) );
  INV_X1 npu_inst_pe_1_3_0_U36 ( .A(npu_inst_pe_1_3_0_n78), .ZN(
        npu_inst_pe_1_3_0_n34) );
  AND2_X1 npu_inst_pe_1_3_0_U35 ( .A1(npu_inst_pe_1_3_0_o_data_h_1_), .A2(
        npu_inst_pe_1_3_0_int_q_weight_1_), .ZN(npu_inst_pe_1_3_0_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_3_0_U34 ( .A1(npu_inst_pe_1_3_0_o_data_h_0_), .A2(
        npu_inst_pe_1_3_0_int_q_weight_1_), .ZN(npu_inst_pe_1_3_0_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_3_0_U33 ( .A(npu_inst_pe_1_3_0_int_data_1_), .ZN(
        npu_inst_pe_1_3_0_n14) );
  AOI22_X1 npu_inst_pe_1_3_0_U32 ( .A1(npu_inst_n57), .A2(
        npu_inst_int_data_y_4__0__1_), .B1(npu_inst_pe_1_3_0_n3), .B2(
        npu_inst_int_data_x_3__1__1_), .ZN(npu_inst_pe_1_3_0_n63) );
  AOI22_X1 npu_inst_pe_1_3_0_U31 ( .A1(npu_inst_n57), .A2(
        npu_inst_int_data_y_4__0__0_), .B1(npu_inst_pe_1_3_0_n3), .B2(
        npu_inst_int_data_x_3__1__0_), .ZN(npu_inst_pe_1_3_0_n61) );
  INV_X1 npu_inst_pe_1_3_0_U30 ( .A(npu_inst_pe_1_3_0_int_data_0_), .ZN(
        npu_inst_pe_1_3_0_n13) );
  INV_X1 npu_inst_pe_1_3_0_U29 ( .A(npu_inst_n70), .ZN(npu_inst_pe_1_3_0_n5)
         );
  OR3_X1 npu_inst_pe_1_3_0_U28 ( .A1(npu_inst_pe_1_3_0_n6), .A2(
        npu_inst_pe_1_3_0_n8), .A3(npu_inst_pe_1_3_0_n5), .ZN(
        npu_inst_pe_1_3_0_n56) );
  OR3_X1 npu_inst_pe_1_3_0_U27 ( .A1(npu_inst_pe_1_3_0_n5), .A2(
        npu_inst_pe_1_3_0_n8), .A3(npu_inst_pe_1_3_0_n7), .ZN(
        npu_inst_pe_1_3_0_n48) );
  INV_X1 npu_inst_pe_1_3_0_U26 ( .A(npu_inst_pe_1_3_0_n5), .ZN(
        npu_inst_pe_1_3_0_n4) );
  INV_X1 npu_inst_pe_1_3_0_U25 ( .A(npu_inst_n125), .ZN(npu_inst_pe_1_3_0_n12)
         );
  OR3_X1 npu_inst_pe_1_3_0_U24 ( .A1(npu_inst_pe_1_3_0_n4), .A2(
        npu_inst_pe_1_3_0_n8), .A3(npu_inst_pe_1_3_0_n7), .ZN(
        npu_inst_pe_1_3_0_n52) );
  OR3_X1 npu_inst_pe_1_3_0_U23 ( .A1(npu_inst_pe_1_3_0_n6), .A2(
        npu_inst_pe_1_3_0_n8), .A3(npu_inst_pe_1_3_0_n4), .ZN(
        npu_inst_pe_1_3_0_n60) );
  NOR2_X1 npu_inst_pe_1_3_0_U22 ( .A1(npu_inst_pe_1_3_0_n60), .A2(
        npu_inst_pe_1_3_0_n3), .ZN(npu_inst_pe_1_3_0_n58) );
  NOR2_X1 npu_inst_pe_1_3_0_U21 ( .A1(npu_inst_pe_1_3_0_n56), .A2(
        npu_inst_pe_1_3_0_n3), .ZN(npu_inst_pe_1_3_0_n54) );
  NOR2_X1 npu_inst_pe_1_3_0_U20 ( .A1(npu_inst_pe_1_3_0_n52), .A2(
        npu_inst_pe_1_3_0_n3), .ZN(npu_inst_pe_1_3_0_n50) );
  NOR2_X1 npu_inst_pe_1_3_0_U19 ( .A1(npu_inst_pe_1_3_0_n48), .A2(
        npu_inst_pe_1_3_0_n3), .ZN(npu_inst_pe_1_3_0_n46) );
  NOR2_X1 npu_inst_pe_1_3_0_U18 ( .A1(npu_inst_pe_1_3_0_n40), .A2(
        npu_inst_pe_1_3_0_n3), .ZN(npu_inst_pe_1_3_0_n38) );
  NOR2_X1 npu_inst_pe_1_3_0_U17 ( .A1(npu_inst_pe_1_3_0_n44), .A2(
        npu_inst_pe_1_3_0_n3), .ZN(npu_inst_pe_1_3_0_n42) );
  BUF_X1 npu_inst_pe_1_3_0_U16 ( .A(npu_inst_n101), .Z(npu_inst_pe_1_3_0_n8)
         );
  BUF_X1 npu_inst_pe_1_3_0_U15 ( .A(npu_inst_pe_1_3_0_n12), .Z(
        npu_inst_pe_1_3_0_n11) );
  BUF_X1 npu_inst_pe_1_3_0_U14 ( .A(npu_inst_pe_1_3_0_n12), .Z(
        npu_inst_pe_1_3_0_n10) );
  BUF_X1 npu_inst_pe_1_3_0_U13 ( .A(npu_inst_pe_1_3_0_n12), .Z(
        npu_inst_pe_1_3_0_n9) );
  INV_X1 npu_inst_pe_1_3_0_U12 ( .A(npu_inst_pe_1_3_0_n38), .ZN(
        npu_inst_pe_1_3_0_n118) );
  INV_X1 npu_inst_pe_1_3_0_U11 ( .A(npu_inst_pe_1_3_0_n58), .ZN(
        npu_inst_pe_1_3_0_n114) );
  INV_X1 npu_inst_pe_1_3_0_U10 ( .A(npu_inst_pe_1_3_0_n54), .ZN(
        npu_inst_pe_1_3_0_n115) );
  INV_X1 npu_inst_pe_1_3_0_U9 ( .A(npu_inst_pe_1_3_0_n50), .ZN(
        npu_inst_pe_1_3_0_n116) );
  INV_X1 npu_inst_pe_1_3_0_U8 ( .A(npu_inst_pe_1_3_0_n46), .ZN(
        npu_inst_pe_1_3_0_n117) );
  INV_X1 npu_inst_pe_1_3_0_U7 ( .A(npu_inst_pe_1_3_0_n42), .ZN(
        npu_inst_pe_1_3_0_n119) );
  BUF_X1 npu_inst_pe_1_3_0_U6 ( .A(npu_inst_n26), .Z(npu_inst_pe_1_3_0_n2) );
  BUF_X1 npu_inst_pe_1_3_0_U5 ( .A(npu_inst_n26), .Z(npu_inst_pe_1_3_0_n1) );
  NOR2_X1 npu_inst_pe_1_3_0_U4 ( .A1(npu_inst_pe_1_3_0_int_q_weight_0_), .A2(
        npu_inst_pe_1_3_0_n1), .ZN(npu_inst_pe_1_3_0_n76) );
  NOR2_X1 npu_inst_pe_1_3_0_U3 ( .A1(npu_inst_pe_1_3_0_n27), .A2(
        npu_inst_pe_1_3_0_n1), .ZN(npu_inst_pe_1_3_0_n77) );
  FA_X1 npu_inst_pe_1_3_0_sub_77_U2_1 ( .A(npu_inst_pe_1_3_0_int_q_acc_1_), 
        .B(npu_inst_pe_1_3_0_n14), .CI(npu_inst_pe_1_3_0_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_3_0_sub_77_carry_2_), .S(npu_inst_pe_1_3_0_N66) );
  FA_X1 npu_inst_pe_1_3_0_add_79_U1_1 ( .A(npu_inst_pe_1_3_0_int_q_acc_1_), 
        .B(npu_inst_pe_1_3_0_int_data_1_), .CI(
        npu_inst_pe_1_3_0_add_79_carry_1_), .CO(
        npu_inst_pe_1_3_0_add_79_carry_2_), .S(npu_inst_pe_1_3_0_N74) );
  NAND3_X1 npu_inst_pe_1_3_0_U109 ( .A1(npu_inst_pe_1_3_0_n5), .A2(
        npu_inst_pe_1_3_0_n7), .A3(npu_inst_pe_1_3_0_n8), .ZN(
        npu_inst_pe_1_3_0_n44) );
  NAND3_X1 npu_inst_pe_1_3_0_U108 ( .A1(npu_inst_pe_1_3_0_n4), .A2(
        npu_inst_pe_1_3_0_n7), .A3(npu_inst_pe_1_3_0_n8), .ZN(
        npu_inst_pe_1_3_0_n40) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_3_0_n34), .CK(
        npu_inst_pe_1_3_0_net3741), .RN(npu_inst_pe_1_3_0_n9), .Q(
        npu_inst_pe_1_3_0_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_3_0_n35), .CK(
        npu_inst_pe_1_3_0_net3741), .RN(npu_inst_pe_1_3_0_n9), .Q(
        npu_inst_pe_1_3_0_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_3_0_n36), .CK(
        npu_inst_pe_1_3_0_net3741), .RN(npu_inst_pe_1_3_0_n9), .Q(
        npu_inst_pe_1_3_0_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_3_0_n98), .CK(
        npu_inst_pe_1_3_0_net3741), .RN(npu_inst_pe_1_3_0_n9), .Q(
        npu_inst_pe_1_3_0_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_3_0_n99), .CK(
        npu_inst_pe_1_3_0_net3741), .RN(npu_inst_pe_1_3_0_n9), .Q(
        npu_inst_pe_1_3_0_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_3_0_n100), 
        .CK(npu_inst_pe_1_3_0_net3741), .RN(npu_inst_pe_1_3_0_n9), .Q(
        npu_inst_pe_1_3_0_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_3_0_n33), .CK(
        npu_inst_pe_1_3_0_net3741), .RN(npu_inst_pe_1_3_0_n9), .Q(
        npu_inst_pe_1_3_0_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_3_0_n101), 
        .CK(npu_inst_pe_1_3_0_net3741), .RN(npu_inst_pe_1_3_0_n9), .Q(
        npu_inst_pe_1_3_0_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_weight_reg_0_ ( .D(npu_inst_n111), .CK(
        npu_inst_pe_1_3_0_net3747), .RN(npu_inst_pe_1_3_0_n9), .Q(
        npu_inst_pe_1_3_0_int_q_weight_0_), .QN(npu_inst_pe_1_3_0_n27) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_weight_reg_1_ ( .D(npu_inst_n117), .CK(
        npu_inst_pe_1_3_0_net3747), .RN(npu_inst_pe_1_3_0_n9), .Q(
        npu_inst_pe_1_3_0_int_q_weight_1_), .QN(npu_inst_pe_1_3_0_n26) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_3_0_n113), 
        .CK(npu_inst_pe_1_3_0_net3747), .RN(npu_inst_pe_1_3_0_n9), .Q(
        npu_inst_pe_1_3_0_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_3_0_n107), 
        .CK(npu_inst_pe_1_3_0_net3747), .RN(npu_inst_pe_1_3_0_n9), .Q(
        npu_inst_pe_1_3_0_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_3_0_n112), 
        .CK(npu_inst_pe_1_3_0_net3747), .RN(npu_inst_pe_1_3_0_n10), .Q(
        npu_inst_pe_1_3_0_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_3_0_n106), 
        .CK(npu_inst_pe_1_3_0_net3747), .RN(npu_inst_pe_1_3_0_n10), .Q(
        npu_inst_pe_1_3_0_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_3_0_n111), 
        .CK(npu_inst_pe_1_3_0_net3747), .RN(npu_inst_pe_1_3_0_n10), .Q(
        npu_inst_pe_1_3_0_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_3_0_n105), 
        .CK(npu_inst_pe_1_3_0_net3747), .RN(npu_inst_pe_1_3_0_n10), .Q(
        npu_inst_pe_1_3_0_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_3_0_n110), 
        .CK(npu_inst_pe_1_3_0_net3747), .RN(npu_inst_pe_1_3_0_n10), .Q(
        npu_inst_pe_1_3_0_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_3_0_n104), 
        .CK(npu_inst_pe_1_3_0_net3747), .RN(npu_inst_pe_1_3_0_n10), .Q(
        npu_inst_pe_1_3_0_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_3_0_n109), 
        .CK(npu_inst_pe_1_3_0_net3747), .RN(npu_inst_pe_1_3_0_n10), .Q(
        npu_inst_pe_1_3_0_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_3_0_n103), 
        .CK(npu_inst_pe_1_3_0_net3747), .RN(npu_inst_pe_1_3_0_n10), .Q(
        npu_inst_pe_1_3_0_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_3_0_n108), 
        .CK(npu_inst_pe_1_3_0_net3747), .RN(npu_inst_pe_1_3_0_n10), .Q(
        npu_inst_pe_1_3_0_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_3_0_n102), 
        .CK(npu_inst_pe_1_3_0_net3747), .RN(npu_inst_pe_1_3_0_n10), .Q(
        npu_inst_pe_1_3_0_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_3_0_n86), 
        .CK(npu_inst_pe_1_3_0_net3747), .RN(npu_inst_pe_1_3_0_n10), .Q(
        npu_inst_pe_1_3_0_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_3_0_n87), 
        .CK(npu_inst_pe_1_3_0_net3747), .RN(npu_inst_pe_1_3_0_n10), .Q(
        npu_inst_pe_1_3_0_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_3_0_n88), 
        .CK(npu_inst_pe_1_3_0_net3747), .RN(npu_inst_pe_1_3_0_n11), .Q(
        npu_inst_pe_1_3_0_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_3_0_n89), 
        .CK(npu_inst_pe_1_3_0_net3747), .RN(npu_inst_pe_1_3_0_n11), .Q(
        npu_inst_pe_1_3_0_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_3_0_n90), 
        .CK(npu_inst_pe_1_3_0_net3747), .RN(npu_inst_pe_1_3_0_n11), .Q(
        npu_inst_pe_1_3_0_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_3_0_n91), 
        .CK(npu_inst_pe_1_3_0_net3747), .RN(npu_inst_pe_1_3_0_n11), .Q(
        npu_inst_pe_1_3_0_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_3_0_n92), 
        .CK(npu_inst_pe_1_3_0_net3747), .RN(npu_inst_pe_1_3_0_n11), .Q(
        npu_inst_pe_1_3_0_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_3_0_n93), 
        .CK(npu_inst_pe_1_3_0_net3747), .RN(npu_inst_pe_1_3_0_n11), .Q(
        npu_inst_pe_1_3_0_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_3_0_n94), 
        .CK(npu_inst_pe_1_3_0_net3747), .RN(npu_inst_pe_1_3_0_n11), .Q(
        npu_inst_pe_1_3_0_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_3_0_n95), 
        .CK(npu_inst_pe_1_3_0_net3747), .RN(npu_inst_pe_1_3_0_n11), .Q(
        npu_inst_pe_1_3_0_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_3_0_n96), 
        .CK(npu_inst_pe_1_3_0_net3747), .RN(npu_inst_pe_1_3_0_n11), .Q(
        npu_inst_pe_1_3_0_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_3_0_n97), 
        .CK(npu_inst_pe_1_3_0_net3747), .RN(npu_inst_pe_1_3_0_n11), .Q(
        npu_inst_pe_1_3_0_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_3_0_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_3_0_N84), .SE(1'b0), .GCK(npu_inst_pe_1_3_0_net3741) );
  CLKGATETST_X1 npu_inst_pe_1_3_0_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n64), .SE(1'b0), .GCK(npu_inst_pe_1_3_0_net3747) );
  MUX2_X1 npu_inst_pe_1_3_1_U162 ( .A(npu_inst_pe_1_3_1_n32), .B(
        npu_inst_pe_1_3_1_n29), .S(npu_inst_pe_1_3_1_n8), .Z(
        npu_inst_pe_1_3_1_N93) );
  MUX2_X1 npu_inst_pe_1_3_1_U161 ( .A(npu_inst_pe_1_3_1_n31), .B(
        npu_inst_pe_1_3_1_n30), .S(npu_inst_pe_1_3_1_n6), .Z(
        npu_inst_pe_1_3_1_n32) );
  MUX2_X1 npu_inst_pe_1_3_1_U160 ( .A(npu_inst_pe_1_3_1_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_3_1_int_q_reg_v_1__0_), .S(npu_inst_pe_1_3_1_n4), .Z(
        npu_inst_pe_1_3_1_n31) );
  MUX2_X1 npu_inst_pe_1_3_1_U159 ( .A(npu_inst_pe_1_3_1_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_3_1_int_q_reg_v_3__0_), .S(npu_inst_pe_1_3_1_n4), .Z(
        npu_inst_pe_1_3_1_n30) );
  MUX2_X1 npu_inst_pe_1_3_1_U158 ( .A(npu_inst_pe_1_3_1_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_3_1_int_q_reg_v_5__0_), .S(npu_inst_pe_1_3_1_n4), .Z(
        npu_inst_pe_1_3_1_n29) );
  MUX2_X1 npu_inst_pe_1_3_1_U157 ( .A(npu_inst_pe_1_3_1_n28), .B(
        npu_inst_pe_1_3_1_n23), .S(npu_inst_pe_1_3_1_n8), .Z(
        npu_inst_pe_1_3_1_N94) );
  MUX2_X1 npu_inst_pe_1_3_1_U156 ( .A(npu_inst_pe_1_3_1_n25), .B(
        npu_inst_pe_1_3_1_n24), .S(npu_inst_pe_1_3_1_n6), .Z(
        npu_inst_pe_1_3_1_n28) );
  MUX2_X1 npu_inst_pe_1_3_1_U155 ( .A(npu_inst_pe_1_3_1_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_3_1_int_q_reg_v_1__1_), .S(npu_inst_pe_1_3_1_n4), .Z(
        npu_inst_pe_1_3_1_n25) );
  MUX2_X1 npu_inst_pe_1_3_1_U154 ( .A(npu_inst_pe_1_3_1_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_3_1_int_q_reg_v_3__1_), .S(npu_inst_pe_1_3_1_n4), .Z(
        npu_inst_pe_1_3_1_n24) );
  MUX2_X1 npu_inst_pe_1_3_1_U153 ( .A(npu_inst_pe_1_3_1_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_3_1_int_q_reg_v_5__1_), .S(npu_inst_pe_1_3_1_n4), .Z(
        npu_inst_pe_1_3_1_n23) );
  MUX2_X1 npu_inst_pe_1_3_1_U152 ( .A(npu_inst_pe_1_3_1_n22), .B(
        npu_inst_pe_1_3_1_n19), .S(npu_inst_pe_1_3_1_n8), .Z(
        npu_inst_int_data_x_3__1__1_) );
  MUX2_X1 npu_inst_pe_1_3_1_U151 ( .A(npu_inst_pe_1_3_1_n21), .B(
        npu_inst_pe_1_3_1_n20), .S(npu_inst_pe_1_3_1_n6), .Z(
        npu_inst_pe_1_3_1_n22) );
  MUX2_X1 npu_inst_pe_1_3_1_U150 ( .A(npu_inst_pe_1_3_1_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_3_1_int_q_reg_h_1__1_), .S(npu_inst_pe_1_3_1_n4), .Z(
        npu_inst_pe_1_3_1_n21) );
  MUX2_X1 npu_inst_pe_1_3_1_U149 ( .A(npu_inst_pe_1_3_1_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_3_1_int_q_reg_h_3__1_), .S(npu_inst_pe_1_3_1_n4), .Z(
        npu_inst_pe_1_3_1_n20) );
  MUX2_X1 npu_inst_pe_1_3_1_U148 ( .A(npu_inst_pe_1_3_1_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_3_1_int_q_reg_h_5__1_), .S(npu_inst_pe_1_3_1_n4), .Z(
        npu_inst_pe_1_3_1_n19) );
  MUX2_X1 npu_inst_pe_1_3_1_U147 ( .A(npu_inst_pe_1_3_1_n18), .B(
        npu_inst_pe_1_3_1_n15), .S(npu_inst_pe_1_3_1_n8), .Z(
        npu_inst_int_data_x_3__1__0_) );
  MUX2_X1 npu_inst_pe_1_3_1_U146 ( .A(npu_inst_pe_1_3_1_n17), .B(
        npu_inst_pe_1_3_1_n16), .S(npu_inst_pe_1_3_1_n6), .Z(
        npu_inst_pe_1_3_1_n18) );
  MUX2_X1 npu_inst_pe_1_3_1_U145 ( .A(npu_inst_pe_1_3_1_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_3_1_int_q_reg_h_1__0_), .S(npu_inst_pe_1_3_1_n4), .Z(
        npu_inst_pe_1_3_1_n17) );
  MUX2_X1 npu_inst_pe_1_3_1_U144 ( .A(npu_inst_pe_1_3_1_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_3_1_int_q_reg_h_3__0_), .S(npu_inst_pe_1_3_1_n4), .Z(
        npu_inst_pe_1_3_1_n16) );
  MUX2_X1 npu_inst_pe_1_3_1_U143 ( .A(npu_inst_pe_1_3_1_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_3_1_int_q_reg_h_5__0_), .S(npu_inst_pe_1_3_1_n4), .Z(
        npu_inst_pe_1_3_1_n15) );
  XOR2_X1 npu_inst_pe_1_3_1_U142 ( .A(npu_inst_pe_1_3_1_int_data_0_), .B(
        npu_inst_pe_1_3_1_int_q_acc_0_), .Z(npu_inst_pe_1_3_1_N73) );
  AND2_X1 npu_inst_pe_1_3_1_U141 ( .A1(npu_inst_pe_1_3_1_int_q_acc_0_), .A2(
        npu_inst_pe_1_3_1_int_data_0_), .ZN(npu_inst_pe_1_3_1_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_3_1_U140 ( .A(npu_inst_pe_1_3_1_int_q_acc_0_), .B(
        npu_inst_pe_1_3_1_n13), .ZN(npu_inst_pe_1_3_1_N65) );
  OR2_X1 npu_inst_pe_1_3_1_U139 ( .A1(npu_inst_pe_1_3_1_n13), .A2(
        npu_inst_pe_1_3_1_int_q_acc_0_), .ZN(npu_inst_pe_1_3_1_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_3_1_U138 ( .A(npu_inst_pe_1_3_1_int_q_acc_2_), .B(
        npu_inst_pe_1_3_1_add_79_carry_2_), .Z(npu_inst_pe_1_3_1_N75) );
  AND2_X1 npu_inst_pe_1_3_1_U137 ( .A1(npu_inst_pe_1_3_1_add_79_carry_2_), 
        .A2(npu_inst_pe_1_3_1_int_q_acc_2_), .ZN(
        npu_inst_pe_1_3_1_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_3_1_U136 ( .A(npu_inst_pe_1_3_1_int_q_acc_3_), .B(
        npu_inst_pe_1_3_1_add_79_carry_3_), .Z(npu_inst_pe_1_3_1_N76) );
  AND2_X1 npu_inst_pe_1_3_1_U135 ( .A1(npu_inst_pe_1_3_1_add_79_carry_3_), 
        .A2(npu_inst_pe_1_3_1_int_q_acc_3_), .ZN(
        npu_inst_pe_1_3_1_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_3_1_U134 ( .A(npu_inst_pe_1_3_1_int_q_acc_4_), .B(
        npu_inst_pe_1_3_1_add_79_carry_4_), .Z(npu_inst_pe_1_3_1_N77) );
  AND2_X1 npu_inst_pe_1_3_1_U133 ( .A1(npu_inst_pe_1_3_1_add_79_carry_4_), 
        .A2(npu_inst_pe_1_3_1_int_q_acc_4_), .ZN(
        npu_inst_pe_1_3_1_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_3_1_U132 ( .A(npu_inst_pe_1_3_1_int_q_acc_5_), .B(
        npu_inst_pe_1_3_1_add_79_carry_5_), .Z(npu_inst_pe_1_3_1_N78) );
  AND2_X1 npu_inst_pe_1_3_1_U131 ( .A1(npu_inst_pe_1_3_1_add_79_carry_5_), 
        .A2(npu_inst_pe_1_3_1_int_q_acc_5_), .ZN(
        npu_inst_pe_1_3_1_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_3_1_U130 ( .A(npu_inst_pe_1_3_1_int_q_acc_6_), .B(
        npu_inst_pe_1_3_1_add_79_carry_6_), .Z(npu_inst_pe_1_3_1_N79) );
  AND2_X1 npu_inst_pe_1_3_1_U129 ( .A1(npu_inst_pe_1_3_1_add_79_carry_6_), 
        .A2(npu_inst_pe_1_3_1_int_q_acc_6_), .ZN(
        npu_inst_pe_1_3_1_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_3_1_U128 ( .A(npu_inst_pe_1_3_1_int_q_acc_7_), .B(
        npu_inst_pe_1_3_1_add_79_carry_7_), .Z(npu_inst_pe_1_3_1_N80) );
  XNOR2_X1 npu_inst_pe_1_3_1_U127 ( .A(npu_inst_pe_1_3_1_sub_77_carry_2_), .B(
        npu_inst_pe_1_3_1_int_q_acc_2_), .ZN(npu_inst_pe_1_3_1_N67) );
  OR2_X1 npu_inst_pe_1_3_1_U126 ( .A1(npu_inst_pe_1_3_1_int_q_acc_2_), .A2(
        npu_inst_pe_1_3_1_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_3_1_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_3_1_U125 ( .A(npu_inst_pe_1_3_1_sub_77_carry_3_), .B(
        npu_inst_pe_1_3_1_int_q_acc_3_), .ZN(npu_inst_pe_1_3_1_N68) );
  OR2_X1 npu_inst_pe_1_3_1_U124 ( .A1(npu_inst_pe_1_3_1_int_q_acc_3_), .A2(
        npu_inst_pe_1_3_1_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_3_1_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_3_1_U123 ( .A(npu_inst_pe_1_3_1_sub_77_carry_4_), .B(
        npu_inst_pe_1_3_1_int_q_acc_4_), .ZN(npu_inst_pe_1_3_1_N69) );
  OR2_X1 npu_inst_pe_1_3_1_U122 ( .A1(npu_inst_pe_1_3_1_int_q_acc_4_), .A2(
        npu_inst_pe_1_3_1_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_3_1_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_3_1_U121 ( .A(npu_inst_pe_1_3_1_sub_77_carry_5_), .B(
        npu_inst_pe_1_3_1_int_q_acc_5_), .ZN(npu_inst_pe_1_3_1_N70) );
  OR2_X1 npu_inst_pe_1_3_1_U120 ( .A1(npu_inst_pe_1_3_1_int_q_acc_5_), .A2(
        npu_inst_pe_1_3_1_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_3_1_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_3_1_U119 ( .A(npu_inst_pe_1_3_1_sub_77_carry_6_), .B(
        npu_inst_pe_1_3_1_int_q_acc_6_), .ZN(npu_inst_pe_1_3_1_N71) );
  OR2_X1 npu_inst_pe_1_3_1_U118 ( .A1(npu_inst_pe_1_3_1_int_q_acc_6_), .A2(
        npu_inst_pe_1_3_1_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_3_1_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_3_1_U117 ( .A(npu_inst_pe_1_3_1_int_q_acc_7_), .B(
        npu_inst_pe_1_3_1_sub_77_carry_7_), .ZN(npu_inst_pe_1_3_1_N72) );
  INV_X1 npu_inst_pe_1_3_1_U116 ( .A(npu_inst_n78), .ZN(npu_inst_pe_1_3_1_n7)
         );
  INV_X1 npu_inst_pe_1_3_1_U115 ( .A(npu_inst_pe_1_3_1_n7), .ZN(
        npu_inst_pe_1_3_1_n6) );
  INV_X1 npu_inst_pe_1_3_1_U114 ( .A(npu_inst_n57), .ZN(npu_inst_pe_1_3_1_n3)
         );
  AOI22_X1 npu_inst_pe_1_3_1_U113 ( .A1(npu_inst_int_data_y_4__1__0_), .A2(
        npu_inst_pe_1_3_1_n58), .B1(npu_inst_pe_1_3_1_n114), .B2(
        npu_inst_pe_1_3_1_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_3_1_n57) );
  INV_X1 npu_inst_pe_1_3_1_U112 ( .A(npu_inst_pe_1_3_1_n57), .ZN(
        npu_inst_pe_1_3_1_n108) );
  AOI22_X1 npu_inst_pe_1_3_1_U111 ( .A1(npu_inst_int_data_y_4__1__0_), .A2(
        npu_inst_pe_1_3_1_n54), .B1(npu_inst_pe_1_3_1_n115), .B2(
        npu_inst_pe_1_3_1_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_3_1_n53) );
  INV_X1 npu_inst_pe_1_3_1_U110 ( .A(npu_inst_pe_1_3_1_n53), .ZN(
        npu_inst_pe_1_3_1_n109) );
  AOI22_X1 npu_inst_pe_1_3_1_U107 ( .A1(npu_inst_int_data_y_4__1__0_), .A2(
        npu_inst_pe_1_3_1_n50), .B1(npu_inst_pe_1_3_1_n116), .B2(
        npu_inst_pe_1_3_1_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_3_1_n49) );
  INV_X1 npu_inst_pe_1_3_1_U106 ( .A(npu_inst_pe_1_3_1_n49), .ZN(
        npu_inst_pe_1_3_1_n110) );
  AOI22_X1 npu_inst_pe_1_3_1_U105 ( .A1(npu_inst_int_data_y_4__1__0_), .A2(
        npu_inst_pe_1_3_1_n46), .B1(npu_inst_pe_1_3_1_n117), .B2(
        npu_inst_pe_1_3_1_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_3_1_n45) );
  INV_X1 npu_inst_pe_1_3_1_U104 ( .A(npu_inst_pe_1_3_1_n45), .ZN(
        npu_inst_pe_1_3_1_n111) );
  AOI22_X1 npu_inst_pe_1_3_1_U103 ( .A1(npu_inst_int_data_y_4__1__0_), .A2(
        npu_inst_pe_1_3_1_n42), .B1(npu_inst_pe_1_3_1_n119), .B2(
        npu_inst_pe_1_3_1_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_3_1_n41) );
  INV_X1 npu_inst_pe_1_3_1_U102 ( .A(npu_inst_pe_1_3_1_n41), .ZN(
        npu_inst_pe_1_3_1_n112) );
  AOI22_X1 npu_inst_pe_1_3_1_U101 ( .A1(npu_inst_int_data_y_4__1__1_), .A2(
        npu_inst_pe_1_3_1_n58), .B1(npu_inst_pe_1_3_1_n114), .B2(
        npu_inst_pe_1_3_1_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_3_1_n59) );
  INV_X1 npu_inst_pe_1_3_1_U100 ( .A(npu_inst_pe_1_3_1_n59), .ZN(
        npu_inst_pe_1_3_1_n102) );
  AOI22_X1 npu_inst_pe_1_3_1_U99 ( .A1(npu_inst_int_data_y_4__1__1_), .A2(
        npu_inst_pe_1_3_1_n54), .B1(npu_inst_pe_1_3_1_n115), .B2(
        npu_inst_pe_1_3_1_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_3_1_n55) );
  INV_X1 npu_inst_pe_1_3_1_U98 ( .A(npu_inst_pe_1_3_1_n55), .ZN(
        npu_inst_pe_1_3_1_n103) );
  AOI22_X1 npu_inst_pe_1_3_1_U97 ( .A1(npu_inst_int_data_y_4__1__1_), .A2(
        npu_inst_pe_1_3_1_n50), .B1(npu_inst_pe_1_3_1_n116), .B2(
        npu_inst_pe_1_3_1_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_3_1_n51) );
  INV_X1 npu_inst_pe_1_3_1_U96 ( .A(npu_inst_pe_1_3_1_n51), .ZN(
        npu_inst_pe_1_3_1_n104) );
  AOI22_X1 npu_inst_pe_1_3_1_U95 ( .A1(npu_inst_int_data_y_4__1__1_), .A2(
        npu_inst_pe_1_3_1_n46), .B1(npu_inst_pe_1_3_1_n117), .B2(
        npu_inst_pe_1_3_1_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_3_1_n47) );
  INV_X1 npu_inst_pe_1_3_1_U94 ( .A(npu_inst_pe_1_3_1_n47), .ZN(
        npu_inst_pe_1_3_1_n105) );
  AOI22_X1 npu_inst_pe_1_3_1_U93 ( .A1(npu_inst_int_data_y_4__1__1_), .A2(
        npu_inst_pe_1_3_1_n42), .B1(npu_inst_pe_1_3_1_n119), .B2(
        npu_inst_pe_1_3_1_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_3_1_n43) );
  INV_X1 npu_inst_pe_1_3_1_U92 ( .A(npu_inst_pe_1_3_1_n43), .ZN(
        npu_inst_pe_1_3_1_n106) );
  AOI22_X1 npu_inst_pe_1_3_1_U91 ( .A1(npu_inst_pe_1_3_1_n38), .A2(
        npu_inst_int_data_y_4__1__1_), .B1(npu_inst_pe_1_3_1_n118), .B2(
        npu_inst_pe_1_3_1_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_3_1_n39) );
  INV_X1 npu_inst_pe_1_3_1_U90 ( .A(npu_inst_pe_1_3_1_n39), .ZN(
        npu_inst_pe_1_3_1_n107) );
  AOI22_X1 npu_inst_pe_1_3_1_U89 ( .A1(npu_inst_pe_1_3_1_n38), .A2(
        npu_inst_int_data_y_4__1__0_), .B1(npu_inst_pe_1_3_1_n118), .B2(
        npu_inst_pe_1_3_1_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_3_1_n37) );
  INV_X1 npu_inst_pe_1_3_1_U88 ( .A(npu_inst_pe_1_3_1_n37), .ZN(
        npu_inst_pe_1_3_1_n113) );
  NAND2_X1 npu_inst_pe_1_3_1_U87 ( .A1(npu_inst_pe_1_3_1_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_3_1_n60), .ZN(npu_inst_pe_1_3_1_n74) );
  OAI21_X1 npu_inst_pe_1_3_1_U86 ( .B1(npu_inst_pe_1_3_1_n63), .B2(
        npu_inst_pe_1_3_1_n60), .A(npu_inst_pe_1_3_1_n74), .ZN(
        npu_inst_pe_1_3_1_n97) );
  NAND2_X1 npu_inst_pe_1_3_1_U85 ( .A1(npu_inst_pe_1_3_1_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_3_1_n60), .ZN(npu_inst_pe_1_3_1_n73) );
  OAI21_X1 npu_inst_pe_1_3_1_U84 ( .B1(npu_inst_pe_1_3_1_n61), .B2(
        npu_inst_pe_1_3_1_n60), .A(npu_inst_pe_1_3_1_n73), .ZN(
        npu_inst_pe_1_3_1_n96) );
  NAND2_X1 npu_inst_pe_1_3_1_U83 ( .A1(npu_inst_pe_1_3_1_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_3_1_n56), .ZN(npu_inst_pe_1_3_1_n72) );
  OAI21_X1 npu_inst_pe_1_3_1_U82 ( .B1(npu_inst_pe_1_3_1_n63), .B2(
        npu_inst_pe_1_3_1_n56), .A(npu_inst_pe_1_3_1_n72), .ZN(
        npu_inst_pe_1_3_1_n95) );
  NAND2_X1 npu_inst_pe_1_3_1_U81 ( .A1(npu_inst_pe_1_3_1_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_3_1_n56), .ZN(npu_inst_pe_1_3_1_n71) );
  OAI21_X1 npu_inst_pe_1_3_1_U80 ( .B1(npu_inst_pe_1_3_1_n61), .B2(
        npu_inst_pe_1_3_1_n56), .A(npu_inst_pe_1_3_1_n71), .ZN(
        npu_inst_pe_1_3_1_n94) );
  NAND2_X1 npu_inst_pe_1_3_1_U79 ( .A1(npu_inst_pe_1_3_1_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_3_1_n52), .ZN(npu_inst_pe_1_3_1_n70) );
  OAI21_X1 npu_inst_pe_1_3_1_U78 ( .B1(npu_inst_pe_1_3_1_n63), .B2(
        npu_inst_pe_1_3_1_n52), .A(npu_inst_pe_1_3_1_n70), .ZN(
        npu_inst_pe_1_3_1_n93) );
  NAND2_X1 npu_inst_pe_1_3_1_U77 ( .A1(npu_inst_pe_1_3_1_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_3_1_n52), .ZN(npu_inst_pe_1_3_1_n69) );
  OAI21_X1 npu_inst_pe_1_3_1_U76 ( .B1(npu_inst_pe_1_3_1_n61), .B2(
        npu_inst_pe_1_3_1_n52), .A(npu_inst_pe_1_3_1_n69), .ZN(
        npu_inst_pe_1_3_1_n92) );
  NAND2_X1 npu_inst_pe_1_3_1_U75 ( .A1(npu_inst_pe_1_3_1_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_3_1_n48), .ZN(npu_inst_pe_1_3_1_n68) );
  OAI21_X1 npu_inst_pe_1_3_1_U74 ( .B1(npu_inst_pe_1_3_1_n63), .B2(
        npu_inst_pe_1_3_1_n48), .A(npu_inst_pe_1_3_1_n68), .ZN(
        npu_inst_pe_1_3_1_n91) );
  NAND2_X1 npu_inst_pe_1_3_1_U73 ( .A1(npu_inst_pe_1_3_1_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_3_1_n48), .ZN(npu_inst_pe_1_3_1_n67) );
  OAI21_X1 npu_inst_pe_1_3_1_U72 ( .B1(npu_inst_pe_1_3_1_n61), .B2(
        npu_inst_pe_1_3_1_n48), .A(npu_inst_pe_1_3_1_n67), .ZN(
        npu_inst_pe_1_3_1_n90) );
  NAND2_X1 npu_inst_pe_1_3_1_U71 ( .A1(npu_inst_pe_1_3_1_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_3_1_n44), .ZN(npu_inst_pe_1_3_1_n66) );
  OAI21_X1 npu_inst_pe_1_3_1_U70 ( .B1(npu_inst_pe_1_3_1_n63), .B2(
        npu_inst_pe_1_3_1_n44), .A(npu_inst_pe_1_3_1_n66), .ZN(
        npu_inst_pe_1_3_1_n89) );
  NAND2_X1 npu_inst_pe_1_3_1_U69 ( .A1(npu_inst_pe_1_3_1_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_3_1_n44), .ZN(npu_inst_pe_1_3_1_n65) );
  OAI21_X1 npu_inst_pe_1_3_1_U68 ( .B1(npu_inst_pe_1_3_1_n61), .B2(
        npu_inst_pe_1_3_1_n44), .A(npu_inst_pe_1_3_1_n65), .ZN(
        npu_inst_pe_1_3_1_n88) );
  NAND2_X1 npu_inst_pe_1_3_1_U67 ( .A1(npu_inst_pe_1_3_1_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_3_1_n40), .ZN(npu_inst_pe_1_3_1_n64) );
  OAI21_X1 npu_inst_pe_1_3_1_U66 ( .B1(npu_inst_pe_1_3_1_n63), .B2(
        npu_inst_pe_1_3_1_n40), .A(npu_inst_pe_1_3_1_n64), .ZN(
        npu_inst_pe_1_3_1_n87) );
  NAND2_X1 npu_inst_pe_1_3_1_U65 ( .A1(npu_inst_pe_1_3_1_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_3_1_n40), .ZN(npu_inst_pe_1_3_1_n62) );
  OAI21_X1 npu_inst_pe_1_3_1_U64 ( .B1(npu_inst_pe_1_3_1_n61), .B2(
        npu_inst_pe_1_3_1_n40), .A(npu_inst_pe_1_3_1_n62), .ZN(
        npu_inst_pe_1_3_1_n86) );
  AND2_X1 npu_inst_pe_1_3_1_U63 ( .A1(npu_inst_pe_1_3_1_N93), .A2(npu_inst_n57), .ZN(npu_inst_int_data_y_3__1__0_) );
  AND2_X1 npu_inst_pe_1_3_1_U62 ( .A1(npu_inst_n57), .A2(npu_inst_pe_1_3_1_N94), .ZN(npu_inst_int_data_y_3__1__1_) );
  NOR3_X1 npu_inst_pe_1_3_1_U61 ( .A1(npu_inst_pe_1_3_1_n26), .A2(npu_inst_n57), .A3(npu_inst_int_ckg[38]), .ZN(npu_inst_pe_1_3_1_n85) );
  OR2_X1 npu_inst_pe_1_3_1_U60 ( .A1(npu_inst_pe_1_3_1_n85), .A2(
        npu_inst_pe_1_3_1_n2), .ZN(npu_inst_pe_1_3_1_N84) );
  AND2_X1 npu_inst_pe_1_3_1_U59 ( .A1(npu_inst_pe_1_3_1_int_q_acc_0_), .A2(
        npu_inst_pe_1_3_1_n1), .ZN(npu_inst_int_data_res_3__1__0_) );
  AND2_X1 npu_inst_pe_1_3_1_U58 ( .A1(npu_inst_pe_1_3_1_n2), .A2(
        npu_inst_pe_1_3_1_int_q_acc_7_), .ZN(npu_inst_int_data_res_3__1__7_)
         );
  AND2_X1 npu_inst_pe_1_3_1_U57 ( .A1(npu_inst_pe_1_3_1_int_q_acc_1_), .A2(
        npu_inst_pe_1_3_1_n1), .ZN(npu_inst_int_data_res_3__1__1_) );
  AND2_X1 npu_inst_pe_1_3_1_U56 ( .A1(npu_inst_pe_1_3_1_int_q_acc_2_), .A2(
        npu_inst_pe_1_3_1_n1), .ZN(npu_inst_int_data_res_3__1__2_) );
  AND2_X1 npu_inst_pe_1_3_1_U55 ( .A1(npu_inst_pe_1_3_1_int_q_acc_3_), .A2(
        npu_inst_pe_1_3_1_n2), .ZN(npu_inst_int_data_res_3__1__3_) );
  AND2_X1 npu_inst_pe_1_3_1_U54 ( .A1(npu_inst_pe_1_3_1_int_q_acc_4_), .A2(
        npu_inst_pe_1_3_1_n2), .ZN(npu_inst_int_data_res_3__1__4_) );
  AND2_X1 npu_inst_pe_1_3_1_U53 ( .A1(npu_inst_pe_1_3_1_int_q_acc_5_), .A2(
        npu_inst_pe_1_3_1_n2), .ZN(npu_inst_int_data_res_3__1__5_) );
  AND2_X1 npu_inst_pe_1_3_1_U52 ( .A1(npu_inst_pe_1_3_1_int_q_acc_6_), .A2(
        npu_inst_pe_1_3_1_n2), .ZN(npu_inst_int_data_res_3__1__6_) );
  AOI222_X1 npu_inst_pe_1_3_1_U51 ( .A1(npu_inst_int_data_res_4__1__0_), .A2(
        npu_inst_pe_1_3_1_n1), .B1(npu_inst_pe_1_3_1_N73), .B2(
        npu_inst_pe_1_3_1_n76), .C1(npu_inst_pe_1_3_1_N65), .C2(
        npu_inst_pe_1_3_1_n77), .ZN(npu_inst_pe_1_3_1_n84) );
  INV_X1 npu_inst_pe_1_3_1_U50 ( .A(npu_inst_pe_1_3_1_n84), .ZN(
        npu_inst_pe_1_3_1_n101) );
  AOI222_X1 npu_inst_pe_1_3_1_U49 ( .A1(npu_inst_int_data_res_4__1__7_), .A2(
        npu_inst_pe_1_3_1_n1), .B1(npu_inst_pe_1_3_1_N80), .B2(
        npu_inst_pe_1_3_1_n76), .C1(npu_inst_pe_1_3_1_N72), .C2(
        npu_inst_pe_1_3_1_n77), .ZN(npu_inst_pe_1_3_1_n75) );
  INV_X1 npu_inst_pe_1_3_1_U48 ( .A(npu_inst_pe_1_3_1_n75), .ZN(
        npu_inst_pe_1_3_1_n33) );
  AOI222_X1 npu_inst_pe_1_3_1_U47 ( .A1(npu_inst_int_data_res_4__1__1_), .A2(
        npu_inst_pe_1_3_1_n1), .B1(npu_inst_pe_1_3_1_N74), .B2(
        npu_inst_pe_1_3_1_n76), .C1(npu_inst_pe_1_3_1_N66), .C2(
        npu_inst_pe_1_3_1_n77), .ZN(npu_inst_pe_1_3_1_n83) );
  INV_X1 npu_inst_pe_1_3_1_U46 ( .A(npu_inst_pe_1_3_1_n83), .ZN(
        npu_inst_pe_1_3_1_n100) );
  AOI222_X1 npu_inst_pe_1_3_1_U45 ( .A1(npu_inst_int_data_res_4__1__2_), .A2(
        npu_inst_pe_1_3_1_n1), .B1(npu_inst_pe_1_3_1_N75), .B2(
        npu_inst_pe_1_3_1_n76), .C1(npu_inst_pe_1_3_1_N67), .C2(
        npu_inst_pe_1_3_1_n77), .ZN(npu_inst_pe_1_3_1_n82) );
  INV_X1 npu_inst_pe_1_3_1_U44 ( .A(npu_inst_pe_1_3_1_n82), .ZN(
        npu_inst_pe_1_3_1_n99) );
  AOI222_X1 npu_inst_pe_1_3_1_U43 ( .A1(npu_inst_int_data_res_4__1__3_), .A2(
        npu_inst_pe_1_3_1_n1), .B1(npu_inst_pe_1_3_1_N76), .B2(
        npu_inst_pe_1_3_1_n76), .C1(npu_inst_pe_1_3_1_N68), .C2(
        npu_inst_pe_1_3_1_n77), .ZN(npu_inst_pe_1_3_1_n81) );
  INV_X1 npu_inst_pe_1_3_1_U42 ( .A(npu_inst_pe_1_3_1_n81), .ZN(
        npu_inst_pe_1_3_1_n98) );
  AOI222_X1 npu_inst_pe_1_3_1_U41 ( .A1(npu_inst_int_data_res_4__1__4_), .A2(
        npu_inst_pe_1_3_1_n1), .B1(npu_inst_pe_1_3_1_N77), .B2(
        npu_inst_pe_1_3_1_n76), .C1(npu_inst_pe_1_3_1_N69), .C2(
        npu_inst_pe_1_3_1_n77), .ZN(npu_inst_pe_1_3_1_n80) );
  INV_X1 npu_inst_pe_1_3_1_U40 ( .A(npu_inst_pe_1_3_1_n80), .ZN(
        npu_inst_pe_1_3_1_n36) );
  AOI222_X1 npu_inst_pe_1_3_1_U39 ( .A1(npu_inst_int_data_res_4__1__5_), .A2(
        npu_inst_pe_1_3_1_n1), .B1(npu_inst_pe_1_3_1_N78), .B2(
        npu_inst_pe_1_3_1_n76), .C1(npu_inst_pe_1_3_1_N70), .C2(
        npu_inst_pe_1_3_1_n77), .ZN(npu_inst_pe_1_3_1_n79) );
  INV_X1 npu_inst_pe_1_3_1_U38 ( .A(npu_inst_pe_1_3_1_n79), .ZN(
        npu_inst_pe_1_3_1_n35) );
  AOI222_X1 npu_inst_pe_1_3_1_U37 ( .A1(npu_inst_int_data_res_4__1__6_), .A2(
        npu_inst_pe_1_3_1_n1), .B1(npu_inst_pe_1_3_1_N79), .B2(
        npu_inst_pe_1_3_1_n76), .C1(npu_inst_pe_1_3_1_N71), .C2(
        npu_inst_pe_1_3_1_n77), .ZN(npu_inst_pe_1_3_1_n78) );
  INV_X1 npu_inst_pe_1_3_1_U36 ( .A(npu_inst_pe_1_3_1_n78), .ZN(
        npu_inst_pe_1_3_1_n34) );
  INV_X1 npu_inst_pe_1_3_1_U35 ( .A(npu_inst_pe_1_3_1_int_data_1_), .ZN(
        npu_inst_pe_1_3_1_n14) );
  AND2_X1 npu_inst_pe_1_3_1_U34 ( .A1(npu_inst_int_data_x_3__1__1_), .A2(
        npu_inst_pe_1_3_1_int_q_weight_1_), .ZN(npu_inst_pe_1_3_1_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_3_1_U33 ( .A1(npu_inst_int_data_x_3__1__0_), .A2(
        npu_inst_pe_1_3_1_int_q_weight_1_), .ZN(npu_inst_pe_1_3_1_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_3_1_U32 ( .A1(npu_inst_n57), .A2(
        npu_inst_int_data_y_4__1__1_), .B1(npu_inst_pe_1_3_1_n3), .B2(
        npu_inst_int_data_x_3__2__1_), .ZN(npu_inst_pe_1_3_1_n63) );
  AOI22_X1 npu_inst_pe_1_3_1_U31 ( .A1(npu_inst_n57), .A2(
        npu_inst_int_data_y_4__1__0_), .B1(npu_inst_pe_1_3_1_n3), .B2(
        npu_inst_int_data_x_3__2__0_), .ZN(npu_inst_pe_1_3_1_n61) );
  INV_X1 npu_inst_pe_1_3_1_U30 ( .A(npu_inst_pe_1_3_1_int_data_0_), .ZN(
        npu_inst_pe_1_3_1_n13) );
  INV_X1 npu_inst_pe_1_3_1_U29 ( .A(npu_inst_n70), .ZN(npu_inst_pe_1_3_1_n5)
         );
  OR3_X1 npu_inst_pe_1_3_1_U28 ( .A1(npu_inst_pe_1_3_1_n6), .A2(
        npu_inst_pe_1_3_1_n8), .A3(npu_inst_pe_1_3_1_n5), .ZN(
        npu_inst_pe_1_3_1_n56) );
  OR3_X1 npu_inst_pe_1_3_1_U27 ( .A1(npu_inst_pe_1_3_1_n5), .A2(
        npu_inst_pe_1_3_1_n8), .A3(npu_inst_pe_1_3_1_n7), .ZN(
        npu_inst_pe_1_3_1_n48) );
  INV_X1 npu_inst_pe_1_3_1_U26 ( .A(npu_inst_pe_1_3_1_n5), .ZN(
        npu_inst_pe_1_3_1_n4) );
  INV_X1 npu_inst_pe_1_3_1_U25 ( .A(npu_inst_n125), .ZN(npu_inst_pe_1_3_1_n12)
         );
  OR3_X1 npu_inst_pe_1_3_1_U24 ( .A1(npu_inst_pe_1_3_1_n4), .A2(
        npu_inst_pe_1_3_1_n8), .A3(npu_inst_pe_1_3_1_n7), .ZN(
        npu_inst_pe_1_3_1_n52) );
  OR3_X1 npu_inst_pe_1_3_1_U23 ( .A1(npu_inst_pe_1_3_1_n6), .A2(
        npu_inst_pe_1_3_1_n8), .A3(npu_inst_pe_1_3_1_n4), .ZN(
        npu_inst_pe_1_3_1_n60) );
  NOR2_X1 npu_inst_pe_1_3_1_U22 ( .A1(npu_inst_pe_1_3_1_n60), .A2(
        npu_inst_pe_1_3_1_n3), .ZN(npu_inst_pe_1_3_1_n58) );
  NOR2_X1 npu_inst_pe_1_3_1_U21 ( .A1(npu_inst_pe_1_3_1_n56), .A2(
        npu_inst_pe_1_3_1_n3), .ZN(npu_inst_pe_1_3_1_n54) );
  NOR2_X1 npu_inst_pe_1_3_1_U20 ( .A1(npu_inst_pe_1_3_1_n52), .A2(
        npu_inst_pe_1_3_1_n3), .ZN(npu_inst_pe_1_3_1_n50) );
  NOR2_X1 npu_inst_pe_1_3_1_U19 ( .A1(npu_inst_pe_1_3_1_n48), .A2(
        npu_inst_pe_1_3_1_n3), .ZN(npu_inst_pe_1_3_1_n46) );
  NOR2_X1 npu_inst_pe_1_3_1_U18 ( .A1(npu_inst_pe_1_3_1_n40), .A2(
        npu_inst_pe_1_3_1_n3), .ZN(npu_inst_pe_1_3_1_n38) );
  NOR2_X1 npu_inst_pe_1_3_1_U17 ( .A1(npu_inst_pe_1_3_1_n44), .A2(
        npu_inst_pe_1_3_1_n3), .ZN(npu_inst_pe_1_3_1_n42) );
  BUF_X1 npu_inst_pe_1_3_1_U16 ( .A(npu_inst_n101), .Z(npu_inst_pe_1_3_1_n8)
         );
  BUF_X1 npu_inst_pe_1_3_1_U15 ( .A(npu_inst_pe_1_3_1_n12), .Z(
        npu_inst_pe_1_3_1_n11) );
  BUF_X1 npu_inst_pe_1_3_1_U14 ( .A(npu_inst_pe_1_3_1_n12), .Z(
        npu_inst_pe_1_3_1_n10) );
  BUF_X1 npu_inst_pe_1_3_1_U13 ( .A(npu_inst_pe_1_3_1_n12), .Z(
        npu_inst_pe_1_3_1_n9) );
  INV_X1 npu_inst_pe_1_3_1_U12 ( .A(npu_inst_pe_1_3_1_n38), .ZN(
        npu_inst_pe_1_3_1_n118) );
  INV_X1 npu_inst_pe_1_3_1_U11 ( .A(npu_inst_pe_1_3_1_n58), .ZN(
        npu_inst_pe_1_3_1_n114) );
  INV_X1 npu_inst_pe_1_3_1_U10 ( .A(npu_inst_pe_1_3_1_n54), .ZN(
        npu_inst_pe_1_3_1_n115) );
  INV_X1 npu_inst_pe_1_3_1_U9 ( .A(npu_inst_pe_1_3_1_n50), .ZN(
        npu_inst_pe_1_3_1_n116) );
  INV_X1 npu_inst_pe_1_3_1_U8 ( .A(npu_inst_pe_1_3_1_n46), .ZN(
        npu_inst_pe_1_3_1_n117) );
  INV_X1 npu_inst_pe_1_3_1_U7 ( .A(npu_inst_pe_1_3_1_n42), .ZN(
        npu_inst_pe_1_3_1_n119) );
  BUF_X1 npu_inst_pe_1_3_1_U6 ( .A(npu_inst_n26), .Z(npu_inst_pe_1_3_1_n2) );
  BUF_X1 npu_inst_pe_1_3_1_U5 ( .A(npu_inst_n26), .Z(npu_inst_pe_1_3_1_n1) );
  NOR2_X1 npu_inst_pe_1_3_1_U4 ( .A1(npu_inst_pe_1_3_1_int_q_weight_0_), .A2(
        npu_inst_pe_1_3_1_n1), .ZN(npu_inst_pe_1_3_1_n76) );
  NOR2_X1 npu_inst_pe_1_3_1_U3 ( .A1(npu_inst_pe_1_3_1_n27), .A2(
        npu_inst_pe_1_3_1_n1), .ZN(npu_inst_pe_1_3_1_n77) );
  FA_X1 npu_inst_pe_1_3_1_sub_77_U2_1 ( .A(npu_inst_pe_1_3_1_int_q_acc_1_), 
        .B(npu_inst_pe_1_3_1_n14), .CI(npu_inst_pe_1_3_1_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_3_1_sub_77_carry_2_), .S(npu_inst_pe_1_3_1_N66) );
  FA_X1 npu_inst_pe_1_3_1_add_79_U1_1 ( .A(npu_inst_pe_1_3_1_int_q_acc_1_), 
        .B(npu_inst_pe_1_3_1_int_data_1_), .CI(
        npu_inst_pe_1_3_1_add_79_carry_1_), .CO(
        npu_inst_pe_1_3_1_add_79_carry_2_), .S(npu_inst_pe_1_3_1_N74) );
  NAND3_X1 npu_inst_pe_1_3_1_U109 ( .A1(npu_inst_pe_1_3_1_n5), .A2(
        npu_inst_pe_1_3_1_n7), .A3(npu_inst_pe_1_3_1_n8), .ZN(
        npu_inst_pe_1_3_1_n44) );
  NAND3_X1 npu_inst_pe_1_3_1_U108 ( .A1(npu_inst_pe_1_3_1_n4), .A2(
        npu_inst_pe_1_3_1_n7), .A3(npu_inst_pe_1_3_1_n8), .ZN(
        npu_inst_pe_1_3_1_n40) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_3_1_n34), .CK(
        npu_inst_pe_1_3_1_net3718), .RN(npu_inst_pe_1_3_1_n9), .Q(
        npu_inst_pe_1_3_1_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_3_1_n35), .CK(
        npu_inst_pe_1_3_1_net3718), .RN(npu_inst_pe_1_3_1_n9), .Q(
        npu_inst_pe_1_3_1_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_3_1_n36), .CK(
        npu_inst_pe_1_3_1_net3718), .RN(npu_inst_pe_1_3_1_n9), .Q(
        npu_inst_pe_1_3_1_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_3_1_n98), .CK(
        npu_inst_pe_1_3_1_net3718), .RN(npu_inst_pe_1_3_1_n9), .Q(
        npu_inst_pe_1_3_1_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_3_1_n99), .CK(
        npu_inst_pe_1_3_1_net3718), .RN(npu_inst_pe_1_3_1_n9), .Q(
        npu_inst_pe_1_3_1_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_3_1_n100), 
        .CK(npu_inst_pe_1_3_1_net3718), .RN(npu_inst_pe_1_3_1_n9), .Q(
        npu_inst_pe_1_3_1_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_3_1_n33), .CK(
        npu_inst_pe_1_3_1_net3718), .RN(npu_inst_pe_1_3_1_n9), .Q(
        npu_inst_pe_1_3_1_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_3_1_n101), 
        .CK(npu_inst_pe_1_3_1_net3718), .RN(npu_inst_pe_1_3_1_n9), .Q(
        npu_inst_pe_1_3_1_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_weight_reg_0_ ( .D(npu_inst_n111), .CK(
        npu_inst_pe_1_3_1_net3724), .RN(npu_inst_pe_1_3_1_n9), .Q(
        npu_inst_pe_1_3_1_int_q_weight_0_), .QN(npu_inst_pe_1_3_1_n27) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_weight_reg_1_ ( .D(npu_inst_n117), .CK(
        npu_inst_pe_1_3_1_net3724), .RN(npu_inst_pe_1_3_1_n9), .Q(
        npu_inst_pe_1_3_1_int_q_weight_1_), .QN(npu_inst_pe_1_3_1_n26) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_3_1_n113), 
        .CK(npu_inst_pe_1_3_1_net3724), .RN(npu_inst_pe_1_3_1_n9), .Q(
        npu_inst_pe_1_3_1_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_3_1_n107), 
        .CK(npu_inst_pe_1_3_1_net3724), .RN(npu_inst_pe_1_3_1_n9), .Q(
        npu_inst_pe_1_3_1_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_3_1_n112), 
        .CK(npu_inst_pe_1_3_1_net3724), .RN(npu_inst_pe_1_3_1_n10), .Q(
        npu_inst_pe_1_3_1_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_3_1_n106), 
        .CK(npu_inst_pe_1_3_1_net3724), .RN(npu_inst_pe_1_3_1_n10), .Q(
        npu_inst_pe_1_3_1_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_3_1_n111), 
        .CK(npu_inst_pe_1_3_1_net3724), .RN(npu_inst_pe_1_3_1_n10), .Q(
        npu_inst_pe_1_3_1_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_3_1_n105), 
        .CK(npu_inst_pe_1_3_1_net3724), .RN(npu_inst_pe_1_3_1_n10), .Q(
        npu_inst_pe_1_3_1_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_3_1_n110), 
        .CK(npu_inst_pe_1_3_1_net3724), .RN(npu_inst_pe_1_3_1_n10), .Q(
        npu_inst_pe_1_3_1_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_3_1_n104), 
        .CK(npu_inst_pe_1_3_1_net3724), .RN(npu_inst_pe_1_3_1_n10), .Q(
        npu_inst_pe_1_3_1_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_3_1_n109), 
        .CK(npu_inst_pe_1_3_1_net3724), .RN(npu_inst_pe_1_3_1_n10), .Q(
        npu_inst_pe_1_3_1_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_3_1_n103), 
        .CK(npu_inst_pe_1_3_1_net3724), .RN(npu_inst_pe_1_3_1_n10), .Q(
        npu_inst_pe_1_3_1_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_3_1_n108), 
        .CK(npu_inst_pe_1_3_1_net3724), .RN(npu_inst_pe_1_3_1_n10), .Q(
        npu_inst_pe_1_3_1_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_3_1_n102), 
        .CK(npu_inst_pe_1_3_1_net3724), .RN(npu_inst_pe_1_3_1_n10), .Q(
        npu_inst_pe_1_3_1_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_3_1_n86), 
        .CK(npu_inst_pe_1_3_1_net3724), .RN(npu_inst_pe_1_3_1_n10), .Q(
        npu_inst_pe_1_3_1_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_3_1_n87), 
        .CK(npu_inst_pe_1_3_1_net3724), .RN(npu_inst_pe_1_3_1_n10), .Q(
        npu_inst_pe_1_3_1_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_3_1_n88), 
        .CK(npu_inst_pe_1_3_1_net3724), .RN(npu_inst_pe_1_3_1_n11), .Q(
        npu_inst_pe_1_3_1_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_3_1_n89), 
        .CK(npu_inst_pe_1_3_1_net3724), .RN(npu_inst_pe_1_3_1_n11), .Q(
        npu_inst_pe_1_3_1_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_3_1_n90), 
        .CK(npu_inst_pe_1_3_1_net3724), .RN(npu_inst_pe_1_3_1_n11), .Q(
        npu_inst_pe_1_3_1_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_3_1_n91), 
        .CK(npu_inst_pe_1_3_1_net3724), .RN(npu_inst_pe_1_3_1_n11), .Q(
        npu_inst_pe_1_3_1_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_3_1_n92), 
        .CK(npu_inst_pe_1_3_1_net3724), .RN(npu_inst_pe_1_3_1_n11), .Q(
        npu_inst_pe_1_3_1_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_3_1_n93), 
        .CK(npu_inst_pe_1_3_1_net3724), .RN(npu_inst_pe_1_3_1_n11), .Q(
        npu_inst_pe_1_3_1_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_3_1_n94), 
        .CK(npu_inst_pe_1_3_1_net3724), .RN(npu_inst_pe_1_3_1_n11), .Q(
        npu_inst_pe_1_3_1_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_3_1_n95), 
        .CK(npu_inst_pe_1_3_1_net3724), .RN(npu_inst_pe_1_3_1_n11), .Q(
        npu_inst_pe_1_3_1_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_3_1_n96), 
        .CK(npu_inst_pe_1_3_1_net3724), .RN(npu_inst_pe_1_3_1_n11), .Q(
        npu_inst_pe_1_3_1_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_3_1_n97), 
        .CK(npu_inst_pe_1_3_1_net3724), .RN(npu_inst_pe_1_3_1_n11), .Q(
        npu_inst_pe_1_3_1_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_3_1_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_3_1_N84), .SE(1'b0), .GCK(npu_inst_pe_1_3_1_net3718) );
  CLKGATETST_X1 npu_inst_pe_1_3_1_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n64), .SE(1'b0), .GCK(npu_inst_pe_1_3_1_net3724) );
  MUX2_X1 npu_inst_pe_1_3_2_U162 ( .A(npu_inst_pe_1_3_2_n32), .B(
        npu_inst_pe_1_3_2_n29), .S(npu_inst_pe_1_3_2_n8), .Z(
        npu_inst_pe_1_3_2_N93) );
  MUX2_X1 npu_inst_pe_1_3_2_U161 ( .A(npu_inst_pe_1_3_2_n31), .B(
        npu_inst_pe_1_3_2_n30), .S(npu_inst_pe_1_3_2_n6), .Z(
        npu_inst_pe_1_3_2_n32) );
  MUX2_X1 npu_inst_pe_1_3_2_U160 ( .A(npu_inst_pe_1_3_2_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_3_2_int_q_reg_v_1__0_), .S(npu_inst_pe_1_3_2_n4), .Z(
        npu_inst_pe_1_3_2_n31) );
  MUX2_X1 npu_inst_pe_1_3_2_U159 ( .A(npu_inst_pe_1_3_2_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_3_2_int_q_reg_v_3__0_), .S(npu_inst_pe_1_3_2_n4), .Z(
        npu_inst_pe_1_3_2_n30) );
  MUX2_X1 npu_inst_pe_1_3_2_U158 ( .A(npu_inst_pe_1_3_2_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_3_2_int_q_reg_v_5__0_), .S(npu_inst_pe_1_3_2_n4), .Z(
        npu_inst_pe_1_3_2_n29) );
  MUX2_X1 npu_inst_pe_1_3_2_U157 ( .A(npu_inst_pe_1_3_2_n28), .B(
        npu_inst_pe_1_3_2_n23), .S(npu_inst_pe_1_3_2_n8), .Z(
        npu_inst_pe_1_3_2_N94) );
  MUX2_X1 npu_inst_pe_1_3_2_U156 ( .A(npu_inst_pe_1_3_2_n25), .B(
        npu_inst_pe_1_3_2_n24), .S(npu_inst_pe_1_3_2_n6), .Z(
        npu_inst_pe_1_3_2_n28) );
  MUX2_X1 npu_inst_pe_1_3_2_U155 ( .A(npu_inst_pe_1_3_2_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_3_2_int_q_reg_v_1__1_), .S(npu_inst_pe_1_3_2_n4), .Z(
        npu_inst_pe_1_3_2_n25) );
  MUX2_X1 npu_inst_pe_1_3_2_U154 ( .A(npu_inst_pe_1_3_2_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_3_2_int_q_reg_v_3__1_), .S(npu_inst_pe_1_3_2_n4), .Z(
        npu_inst_pe_1_3_2_n24) );
  MUX2_X1 npu_inst_pe_1_3_2_U153 ( .A(npu_inst_pe_1_3_2_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_3_2_int_q_reg_v_5__1_), .S(npu_inst_pe_1_3_2_n4), .Z(
        npu_inst_pe_1_3_2_n23) );
  MUX2_X1 npu_inst_pe_1_3_2_U152 ( .A(npu_inst_pe_1_3_2_n22), .B(
        npu_inst_pe_1_3_2_n19), .S(npu_inst_pe_1_3_2_n8), .Z(
        npu_inst_int_data_x_3__2__1_) );
  MUX2_X1 npu_inst_pe_1_3_2_U151 ( .A(npu_inst_pe_1_3_2_n21), .B(
        npu_inst_pe_1_3_2_n20), .S(npu_inst_pe_1_3_2_n6), .Z(
        npu_inst_pe_1_3_2_n22) );
  MUX2_X1 npu_inst_pe_1_3_2_U150 ( .A(npu_inst_pe_1_3_2_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_3_2_int_q_reg_h_1__1_), .S(npu_inst_pe_1_3_2_n4), .Z(
        npu_inst_pe_1_3_2_n21) );
  MUX2_X1 npu_inst_pe_1_3_2_U149 ( .A(npu_inst_pe_1_3_2_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_3_2_int_q_reg_h_3__1_), .S(npu_inst_pe_1_3_2_n4), .Z(
        npu_inst_pe_1_3_2_n20) );
  MUX2_X1 npu_inst_pe_1_3_2_U148 ( .A(npu_inst_pe_1_3_2_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_3_2_int_q_reg_h_5__1_), .S(npu_inst_pe_1_3_2_n4), .Z(
        npu_inst_pe_1_3_2_n19) );
  MUX2_X1 npu_inst_pe_1_3_2_U147 ( .A(npu_inst_pe_1_3_2_n18), .B(
        npu_inst_pe_1_3_2_n15), .S(npu_inst_pe_1_3_2_n8), .Z(
        npu_inst_int_data_x_3__2__0_) );
  MUX2_X1 npu_inst_pe_1_3_2_U146 ( .A(npu_inst_pe_1_3_2_n17), .B(
        npu_inst_pe_1_3_2_n16), .S(npu_inst_pe_1_3_2_n6), .Z(
        npu_inst_pe_1_3_2_n18) );
  MUX2_X1 npu_inst_pe_1_3_2_U145 ( .A(npu_inst_pe_1_3_2_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_3_2_int_q_reg_h_1__0_), .S(npu_inst_pe_1_3_2_n4), .Z(
        npu_inst_pe_1_3_2_n17) );
  MUX2_X1 npu_inst_pe_1_3_2_U144 ( .A(npu_inst_pe_1_3_2_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_3_2_int_q_reg_h_3__0_), .S(npu_inst_pe_1_3_2_n4), .Z(
        npu_inst_pe_1_3_2_n16) );
  MUX2_X1 npu_inst_pe_1_3_2_U143 ( .A(npu_inst_pe_1_3_2_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_3_2_int_q_reg_h_5__0_), .S(npu_inst_pe_1_3_2_n4), .Z(
        npu_inst_pe_1_3_2_n15) );
  XOR2_X1 npu_inst_pe_1_3_2_U142 ( .A(npu_inst_pe_1_3_2_int_data_0_), .B(
        npu_inst_pe_1_3_2_int_q_acc_0_), .Z(npu_inst_pe_1_3_2_N73) );
  AND2_X1 npu_inst_pe_1_3_2_U141 ( .A1(npu_inst_pe_1_3_2_int_q_acc_0_), .A2(
        npu_inst_pe_1_3_2_int_data_0_), .ZN(npu_inst_pe_1_3_2_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_3_2_U140 ( .A(npu_inst_pe_1_3_2_int_q_acc_0_), .B(
        npu_inst_pe_1_3_2_n13), .ZN(npu_inst_pe_1_3_2_N65) );
  OR2_X1 npu_inst_pe_1_3_2_U139 ( .A1(npu_inst_pe_1_3_2_n13), .A2(
        npu_inst_pe_1_3_2_int_q_acc_0_), .ZN(npu_inst_pe_1_3_2_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_3_2_U138 ( .A(npu_inst_pe_1_3_2_int_q_acc_2_), .B(
        npu_inst_pe_1_3_2_add_79_carry_2_), .Z(npu_inst_pe_1_3_2_N75) );
  AND2_X1 npu_inst_pe_1_3_2_U137 ( .A1(npu_inst_pe_1_3_2_add_79_carry_2_), 
        .A2(npu_inst_pe_1_3_2_int_q_acc_2_), .ZN(
        npu_inst_pe_1_3_2_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_3_2_U136 ( .A(npu_inst_pe_1_3_2_int_q_acc_3_), .B(
        npu_inst_pe_1_3_2_add_79_carry_3_), .Z(npu_inst_pe_1_3_2_N76) );
  AND2_X1 npu_inst_pe_1_3_2_U135 ( .A1(npu_inst_pe_1_3_2_add_79_carry_3_), 
        .A2(npu_inst_pe_1_3_2_int_q_acc_3_), .ZN(
        npu_inst_pe_1_3_2_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_3_2_U134 ( .A(npu_inst_pe_1_3_2_int_q_acc_4_), .B(
        npu_inst_pe_1_3_2_add_79_carry_4_), .Z(npu_inst_pe_1_3_2_N77) );
  AND2_X1 npu_inst_pe_1_3_2_U133 ( .A1(npu_inst_pe_1_3_2_add_79_carry_4_), 
        .A2(npu_inst_pe_1_3_2_int_q_acc_4_), .ZN(
        npu_inst_pe_1_3_2_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_3_2_U132 ( .A(npu_inst_pe_1_3_2_int_q_acc_5_), .B(
        npu_inst_pe_1_3_2_add_79_carry_5_), .Z(npu_inst_pe_1_3_2_N78) );
  AND2_X1 npu_inst_pe_1_3_2_U131 ( .A1(npu_inst_pe_1_3_2_add_79_carry_5_), 
        .A2(npu_inst_pe_1_3_2_int_q_acc_5_), .ZN(
        npu_inst_pe_1_3_2_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_3_2_U130 ( .A(npu_inst_pe_1_3_2_int_q_acc_6_), .B(
        npu_inst_pe_1_3_2_add_79_carry_6_), .Z(npu_inst_pe_1_3_2_N79) );
  AND2_X1 npu_inst_pe_1_3_2_U129 ( .A1(npu_inst_pe_1_3_2_add_79_carry_6_), 
        .A2(npu_inst_pe_1_3_2_int_q_acc_6_), .ZN(
        npu_inst_pe_1_3_2_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_3_2_U128 ( .A(npu_inst_pe_1_3_2_int_q_acc_7_), .B(
        npu_inst_pe_1_3_2_add_79_carry_7_), .Z(npu_inst_pe_1_3_2_N80) );
  XNOR2_X1 npu_inst_pe_1_3_2_U127 ( .A(npu_inst_pe_1_3_2_sub_77_carry_2_), .B(
        npu_inst_pe_1_3_2_int_q_acc_2_), .ZN(npu_inst_pe_1_3_2_N67) );
  OR2_X1 npu_inst_pe_1_3_2_U126 ( .A1(npu_inst_pe_1_3_2_int_q_acc_2_), .A2(
        npu_inst_pe_1_3_2_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_3_2_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_3_2_U125 ( .A(npu_inst_pe_1_3_2_sub_77_carry_3_), .B(
        npu_inst_pe_1_3_2_int_q_acc_3_), .ZN(npu_inst_pe_1_3_2_N68) );
  OR2_X1 npu_inst_pe_1_3_2_U124 ( .A1(npu_inst_pe_1_3_2_int_q_acc_3_), .A2(
        npu_inst_pe_1_3_2_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_3_2_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_3_2_U123 ( .A(npu_inst_pe_1_3_2_sub_77_carry_4_), .B(
        npu_inst_pe_1_3_2_int_q_acc_4_), .ZN(npu_inst_pe_1_3_2_N69) );
  OR2_X1 npu_inst_pe_1_3_2_U122 ( .A1(npu_inst_pe_1_3_2_int_q_acc_4_), .A2(
        npu_inst_pe_1_3_2_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_3_2_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_3_2_U121 ( .A(npu_inst_pe_1_3_2_sub_77_carry_5_), .B(
        npu_inst_pe_1_3_2_int_q_acc_5_), .ZN(npu_inst_pe_1_3_2_N70) );
  OR2_X1 npu_inst_pe_1_3_2_U120 ( .A1(npu_inst_pe_1_3_2_int_q_acc_5_), .A2(
        npu_inst_pe_1_3_2_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_3_2_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_3_2_U119 ( .A(npu_inst_pe_1_3_2_sub_77_carry_6_), .B(
        npu_inst_pe_1_3_2_int_q_acc_6_), .ZN(npu_inst_pe_1_3_2_N71) );
  OR2_X1 npu_inst_pe_1_3_2_U118 ( .A1(npu_inst_pe_1_3_2_int_q_acc_6_), .A2(
        npu_inst_pe_1_3_2_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_3_2_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_3_2_U117 ( .A(npu_inst_pe_1_3_2_int_q_acc_7_), .B(
        npu_inst_pe_1_3_2_sub_77_carry_7_), .ZN(npu_inst_pe_1_3_2_N72) );
  INV_X1 npu_inst_pe_1_3_2_U116 ( .A(npu_inst_n78), .ZN(npu_inst_pe_1_3_2_n7)
         );
  INV_X1 npu_inst_pe_1_3_2_U115 ( .A(npu_inst_pe_1_3_2_n7), .ZN(
        npu_inst_pe_1_3_2_n6) );
  INV_X1 npu_inst_pe_1_3_2_U114 ( .A(npu_inst_n57), .ZN(npu_inst_pe_1_3_2_n3)
         );
  AOI22_X1 npu_inst_pe_1_3_2_U113 ( .A1(npu_inst_int_data_y_4__2__0_), .A2(
        npu_inst_pe_1_3_2_n58), .B1(npu_inst_pe_1_3_2_n114), .B2(
        npu_inst_pe_1_3_2_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_3_2_n57) );
  INV_X1 npu_inst_pe_1_3_2_U112 ( .A(npu_inst_pe_1_3_2_n57), .ZN(
        npu_inst_pe_1_3_2_n108) );
  AOI22_X1 npu_inst_pe_1_3_2_U111 ( .A1(npu_inst_int_data_y_4__2__0_), .A2(
        npu_inst_pe_1_3_2_n54), .B1(npu_inst_pe_1_3_2_n115), .B2(
        npu_inst_pe_1_3_2_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_3_2_n53) );
  INV_X1 npu_inst_pe_1_3_2_U110 ( .A(npu_inst_pe_1_3_2_n53), .ZN(
        npu_inst_pe_1_3_2_n109) );
  AOI22_X1 npu_inst_pe_1_3_2_U107 ( .A1(npu_inst_int_data_y_4__2__0_), .A2(
        npu_inst_pe_1_3_2_n50), .B1(npu_inst_pe_1_3_2_n116), .B2(
        npu_inst_pe_1_3_2_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_3_2_n49) );
  INV_X1 npu_inst_pe_1_3_2_U106 ( .A(npu_inst_pe_1_3_2_n49), .ZN(
        npu_inst_pe_1_3_2_n110) );
  AOI22_X1 npu_inst_pe_1_3_2_U105 ( .A1(npu_inst_int_data_y_4__2__0_), .A2(
        npu_inst_pe_1_3_2_n46), .B1(npu_inst_pe_1_3_2_n117), .B2(
        npu_inst_pe_1_3_2_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_3_2_n45) );
  INV_X1 npu_inst_pe_1_3_2_U104 ( .A(npu_inst_pe_1_3_2_n45), .ZN(
        npu_inst_pe_1_3_2_n111) );
  AOI22_X1 npu_inst_pe_1_3_2_U103 ( .A1(npu_inst_int_data_y_4__2__0_), .A2(
        npu_inst_pe_1_3_2_n42), .B1(npu_inst_pe_1_3_2_n119), .B2(
        npu_inst_pe_1_3_2_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_3_2_n41) );
  INV_X1 npu_inst_pe_1_3_2_U102 ( .A(npu_inst_pe_1_3_2_n41), .ZN(
        npu_inst_pe_1_3_2_n112) );
  AOI22_X1 npu_inst_pe_1_3_2_U101 ( .A1(npu_inst_int_data_y_4__2__1_), .A2(
        npu_inst_pe_1_3_2_n58), .B1(npu_inst_pe_1_3_2_n114), .B2(
        npu_inst_pe_1_3_2_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_3_2_n59) );
  INV_X1 npu_inst_pe_1_3_2_U100 ( .A(npu_inst_pe_1_3_2_n59), .ZN(
        npu_inst_pe_1_3_2_n102) );
  AOI22_X1 npu_inst_pe_1_3_2_U99 ( .A1(npu_inst_int_data_y_4__2__1_), .A2(
        npu_inst_pe_1_3_2_n54), .B1(npu_inst_pe_1_3_2_n115), .B2(
        npu_inst_pe_1_3_2_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_3_2_n55) );
  INV_X1 npu_inst_pe_1_3_2_U98 ( .A(npu_inst_pe_1_3_2_n55), .ZN(
        npu_inst_pe_1_3_2_n103) );
  AOI22_X1 npu_inst_pe_1_3_2_U97 ( .A1(npu_inst_int_data_y_4__2__1_), .A2(
        npu_inst_pe_1_3_2_n50), .B1(npu_inst_pe_1_3_2_n116), .B2(
        npu_inst_pe_1_3_2_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_3_2_n51) );
  INV_X1 npu_inst_pe_1_3_2_U96 ( .A(npu_inst_pe_1_3_2_n51), .ZN(
        npu_inst_pe_1_3_2_n104) );
  AOI22_X1 npu_inst_pe_1_3_2_U95 ( .A1(npu_inst_int_data_y_4__2__1_), .A2(
        npu_inst_pe_1_3_2_n46), .B1(npu_inst_pe_1_3_2_n117), .B2(
        npu_inst_pe_1_3_2_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_3_2_n47) );
  INV_X1 npu_inst_pe_1_3_2_U94 ( .A(npu_inst_pe_1_3_2_n47), .ZN(
        npu_inst_pe_1_3_2_n105) );
  AOI22_X1 npu_inst_pe_1_3_2_U93 ( .A1(npu_inst_int_data_y_4__2__1_), .A2(
        npu_inst_pe_1_3_2_n42), .B1(npu_inst_pe_1_3_2_n119), .B2(
        npu_inst_pe_1_3_2_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_3_2_n43) );
  INV_X1 npu_inst_pe_1_3_2_U92 ( .A(npu_inst_pe_1_3_2_n43), .ZN(
        npu_inst_pe_1_3_2_n106) );
  AOI22_X1 npu_inst_pe_1_3_2_U91 ( .A1(npu_inst_pe_1_3_2_n38), .A2(
        npu_inst_int_data_y_4__2__1_), .B1(npu_inst_pe_1_3_2_n118), .B2(
        npu_inst_pe_1_3_2_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_3_2_n39) );
  INV_X1 npu_inst_pe_1_3_2_U90 ( .A(npu_inst_pe_1_3_2_n39), .ZN(
        npu_inst_pe_1_3_2_n107) );
  AOI22_X1 npu_inst_pe_1_3_2_U89 ( .A1(npu_inst_pe_1_3_2_n38), .A2(
        npu_inst_int_data_y_4__2__0_), .B1(npu_inst_pe_1_3_2_n118), .B2(
        npu_inst_pe_1_3_2_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_3_2_n37) );
  INV_X1 npu_inst_pe_1_3_2_U88 ( .A(npu_inst_pe_1_3_2_n37), .ZN(
        npu_inst_pe_1_3_2_n113) );
  NAND2_X1 npu_inst_pe_1_3_2_U87 ( .A1(npu_inst_pe_1_3_2_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_3_2_n60), .ZN(npu_inst_pe_1_3_2_n74) );
  OAI21_X1 npu_inst_pe_1_3_2_U86 ( .B1(npu_inst_pe_1_3_2_n63), .B2(
        npu_inst_pe_1_3_2_n60), .A(npu_inst_pe_1_3_2_n74), .ZN(
        npu_inst_pe_1_3_2_n97) );
  NAND2_X1 npu_inst_pe_1_3_2_U85 ( .A1(npu_inst_pe_1_3_2_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_3_2_n60), .ZN(npu_inst_pe_1_3_2_n73) );
  OAI21_X1 npu_inst_pe_1_3_2_U84 ( .B1(npu_inst_pe_1_3_2_n61), .B2(
        npu_inst_pe_1_3_2_n60), .A(npu_inst_pe_1_3_2_n73), .ZN(
        npu_inst_pe_1_3_2_n96) );
  NAND2_X1 npu_inst_pe_1_3_2_U83 ( .A1(npu_inst_pe_1_3_2_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_3_2_n56), .ZN(npu_inst_pe_1_3_2_n72) );
  OAI21_X1 npu_inst_pe_1_3_2_U82 ( .B1(npu_inst_pe_1_3_2_n63), .B2(
        npu_inst_pe_1_3_2_n56), .A(npu_inst_pe_1_3_2_n72), .ZN(
        npu_inst_pe_1_3_2_n95) );
  NAND2_X1 npu_inst_pe_1_3_2_U81 ( .A1(npu_inst_pe_1_3_2_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_3_2_n56), .ZN(npu_inst_pe_1_3_2_n71) );
  OAI21_X1 npu_inst_pe_1_3_2_U80 ( .B1(npu_inst_pe_1_3_2_n61), .B2(
        npu_inst_pe_1_3_2_n56), .A(npu_inst_pe_1_3_2_n71), .ZN(
        npu_inst_pe_1_3_2_n94) );
  NAND2_X1 npu_inst_pe_1_3_2_U79 ( .A1(npu_inst_pe_1_3_2_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_3_2_n52), .ZN(npu_inst_pe_1_3_2_n70) );
  OAI21_X1 npu_inst_pe_1_3_2_U78 ( .B1(npu_inst_pe_1_3_2_n63), .B2(
        npu_inst_pe_1_3_2_n52), .A(npu_inst_pe_1_3_2_n70), .ZN(
        npu_inst_pe_1_3_2_n93) );
  NAND2_X1 npu_inst_pe_1_3_2_U77 ( .A1(npu_inst_pe_1_3_2_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_3_2_n52), .ZN(npu_inst_pe_1_3_2_n69) );
  OAI21_X1 npu_inst_pe_1_3_2_U76 ( .B1(npu_inst_pe_1_3_2_n61), .B2(
        npu_inst_pe_1_3_2_n52), .A(npu_inst_pe_1_3_2_n69), .ZN(
        npu_inst_pe_1_3_2_n92) );
  NAND2_X1 npu_inst_pe_1_3_2_U75 ( .A1(npu_inst_pe_1_3_2_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_3_2_n48), .ZN(npu_inst_pe_1_3_2_n68) );
  OAI21_X1 npu_inst_pe_1_3_2_U74 ( .B1(npu_inst_pe_1_3_2_n63), .B2(
        npu_inst_pe_1_3_2_n48), .A(npu_inst_pe_1_3_2_n68), .ZN(
        npu_inst_pe_1_3_2_n91) );
  NAND2_X1 npu_inst_pe_1_3_2_U73 ( .A1(npu_inst_pe_1_3_2_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_3_2_n48), .ZN(npu_inst_pe_1_3_2_n67) );
  OAI21_X1 npu_inst_pe_1_3_2_U72 ( .B1(npu_inst_pe_1_3_2_n61), .B2(
        npu_inst_pe_1_3_2_n48), .A(npu_inst_pe_1_3_2_n67), .ZN(
        npu_inst_pe_1_3_2_n90) );
  NAND2_X1 npu_inst_pe_1_3_2_U71 ( .A1(npu_inst_pe_1_3_2_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_3_2_n44), .ZN(npu_inst_pe_1_3_2_n66) );
  OAI21_X1 npu_inst_pe_1_3_2_U70 ( .B1(npu_inst_pe_1_3_2_n63), .B2(
        npu_inst_pe_1_3_2_n44), .A(npu_inst_pe_1_3_2_n66), .ZN(
        npu_inst_pe_1_3_2_n89) );
  NAND2_X1 npu_inst_pe_1_3_2_U69 ( .A1(npu_inst_pe_1_3_2_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_3_2_n44), .ZN(npu_inst_pe_1_3_2_n65) );
  OAI21_X1 npu_inst_pe_1_3_2_U68 ( .B1(npu_inst_pe_1_3_2_n61), .B2(
        npu_inst_pe_1_3_2_n44), .A(npu_inst_pe_1_3_2_n65), .ZN(
        npu_inst_pe_1_3_2_n88) );
  NAND2_X1 npu_inst_pe_1_3_2_U67 ( .A1(npu_inst_pe_1_3_2_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_3_2_n40), .ZN(npu_inst_pe_1_3_2_n64) );
  OAI21_X1 npu_inst_pe_1_3_2_U66 ( .B1(npu_inst_pe_1_3_2_n63), .B2(
        npu_inst_pe_1_3_2_n40), .A(npu_inst_pe_1_3_2_n64), .ZN(
        npu_inst_pe_1_3_2_n87) );
  NAND2_X1 npu_inst_pe_1_3_2_U65 ( .A1(npu_inst_pe_1_3_2_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_3_2_n40), .ZN(npu_inst_pe_1_3_2_n62) );
  OAI21_X1 npu_inst_pe_1_3_2_U64 ( .B1(npu_inst_pe_1_3_2_n61), .B2(
        npu_inst_pe_1_3_2_n40), .A(npu_inst_pe_1_3_2_n62), .ZN(
        npu_inst_pe_1_3_2_n86) );
  AND2_X1 npu_inst_pe_1_3_2_U63 ( .A1(npu_inst_pe_1_3_2_N93), .A2(npu_inst_n57), .ZN(npu_inst_int_data_y_3__2__0_) );
  AND2_X1 npu_inst_pe_1_3_2_U62 ( .A1(npu_inst_n57), .A2(npu_inst_pe_1_3_2_N94), .ZN(npu_inst_int_data_y_3__2__1_) );
  NOR3_X1 npu_inst_pe_1_3_2_U61 ( .A1(npu_inst_pe_1_3_2_n26), .A2(npu_inst_n57), .A3(npu_inst_int_ckg[37]), .ZN(npu_inst_pe_1_3_2_n85) );
  OR2_X1 npu_inst_pe_1_3_2_U60 ( .A1(npu_inst_pe_1_3_2_n85), .A2(
        npu_inst_pe_1_3_2_n2), .ZN(npu_inst_pe_1_3_2_N84) );
  AND2_X1 npu_inst_pe_1_3_2_U59 ( .A1(npu_inst_pe_1_3_2_int_q_acc_0_), .A2(
        npu_inst_pe_1_3_2_n1), .ZN(npu_inst_int_data_res_3__2__0_) );
  AND2_X1 npu_inst_pe_1_3_2_U58 ( .A1(npu_inst_pe_1_3_2_n2), .A2(
        npu_inst_pe_1_3_2_int_q_acc_7_), .ZN(npu_inst_int_data_res_3__2__7_)
         );
  AND2_X1 npu_inst_pe_1_3_2_U57 ( .A1(npu_inst_pe_1_3_2_int_q_acc_1_), .A2(
        npu_inst_pe_1_3_2_n1), .ZN(npu_inst_int_data_res_3__2__1_) );
  AND2_X1 npu_inst_pe_1_3_2_U56 ( .A1(npu_inst_pe_1_3_2_int_q_acc_2_), .A2(
        npu_inst_pe_1_3_2_n1), .ZN(npu_inst_int_data_res_3__2__2_) );
  AND2_X1 npu_inst_pe_1_3_2_U55 ( .A1(npu_inst_pe_1_3_2_int_q_acc_3_), .A2(
        npu_inst_pe_1_3_2_n2), .ZN(npu_inst_int_data_res_3__2__3_) );
  AND2_X1 npu_inst_pe_1_3_2_U54 ( .A1(npu_inst_pe_1_3_2_int_q_acc_4_), .A2(
        npu_inst_pe_1_3_2_n2), .ZN(npu_inst_int_data_res_3__2__4_) );
  AND2_X1 npu_inst_pe_1_3_2_U53 ( .A1(npu_inst_pe_1_3_2_int_q_acc_5_), .A2(
        npu_inst_pe_1_3_2_n2), .ZN(npu_inst_int_data_res_3__2__5_) );
  AND2_X1 npu_inst_pe_1_3_2_U52 ( .A1(npu_inst_pe_1_3_2_int_q_acc_6_), .A2(
        npu_inst_pe_1_3_2_n2), .ZN(npu_inst_int_data_res_3__2__6_) );
  AOI222_X1 npu_inst_pe_1_3_2_U51 ( .A1(npu_inst_int_data_res_4__2__0_), .A2(
        npu_inst_pe_1_3_2_n1), .B1(npu_inst_pe_1_3_2_N73), .B2(
        npu_inst_pe_1_3_2_n76), .C1(npu_inst_pe_1_3_2_N65), .C2(
        npu_inst_pe_1_3_2_n77), .ZN(npu_inst_pe_1_3_2_n84) );
  INV_X1 npu_inst_pe_1_3_2_U50 ( .A(npu_inst_pe_1_3_2_n84), .ZN(
        npu_inst_pe_1_3_2_n101) );
  AOI222_X1 npu_inst_pe_1_3_2_U49 ( .A1(npu_inst_int_data_res_4__2__7_), .A2(
        npu_inst_pe_1_3_2_n1), .B1(npu_inst_pe_1_3_2_N80), .B2(
        npu_inst_pe_1_3_2_n76), .C1(npu_inst_pe_1_3_2_N72), .C2(
        npu_inst_pe_1_3_2_n77), .ZN(npu_inst_pe_1_3_2_n75) );
  INV_X1 npu_inst_pe_1_3_2_U48 ( .A(npu_inst_pe_1_3_2_n75), .ZN(
        npu_inst_pe_1_3_2_n33) );
  AOI222_X1 npu_inst_pe_1_3_2_U47 ( .A1(npu_inst_int_data_res_4__2__1_), .A2(
        npu_inst_pe_1_3_2_n1), .B1(npu_inst_pe_1_3_2_N74), .B2(
        npu_inst_pe_1_3_2_n76), .C1(npu_inst_pe_1_3_2_N66), .C2(
        npu_inst_pe_1_3_2_n77), .ZN(npu_inst_pe_1_3_2_n83) );
  INV_X1 npu_inst_pe_1_3_2_U46 ( .A(npu_inst_pe_1_3_2_n83), .ZN(
        npu_inst_pe_1_3_2_n100) );
  AOI222_X1 npu_inst_pe_1_3_2_U45 ( .A1(npu_inst_int_data_res_4__2__2_), .A2(
        npu_inst_pe_1_3_2_n1), .B1(npu_inst_pe_1_3_2_N75), .B2(
        npu_inst_pe_1_3_2_n76), .C1(npu_inst_pe_1_3_2_N67), .C2(
        npu_inst_pe_1_3_2_n77), .ZN(npu_inst_pe_1_3_2_n82) );
  INV_X1 npu_inst_pe_1_3_2_U44 ( .A(npu_inst_pe_1_3_2_n82), .ZN(
        npu_inst_pe_1_3_2_n99) );
  AOI222_X1 npu_inst_pe_1_3_2_U43 ( .A1(npu_inst_int_data_res_4__2__3_), .A2(
        npu_inst_pe_1_3_2_n1), .B1(npu_inst_pe_1_3_2_N76), .B2(
        npu_inst_pe_1_3_2_n76), .C1(npu_inst_pe_1_3_2_N68), .C2(
        npu_inst_pe_1_3_2_n77), .ZN(npu_inst_pe_1_3_2_n81) );
  INV_X1 npu_inst_pe_1_3_2_U42 ( .A(npu_inst_pe_1_3_2_n81), .ZN(
        npu_inst_pe_1_3_2_n98) );
  AOI222_X1 npu_inst_pe_1_3_2_U41 ( .A1(npu_inst_int_data_res_4__2__4_), .A2(
        npu_inst_pe_1_3_2_n1), .B1(npu_inst_pe_1_3_2_N77), .B2(
        npu_inst_pe_1_3_2_n76), .C1(npu_inst_pe_1_3_2_N69), .C2(
        npu_inst_pe_1_3_2_n77), .ZN(npu_inst_pe_1_3_2_n80) );
  INV_X1 npu_inst_pe_1_3_2_U40 ( .A(npu_inst_pe_1_3_2_n80), .ZN(
        npu_inst_pe_1_3_2_n36) );
  AOI222_X1 npu_inst_pe_1_3_2_U39 ( .A1(npu_inst_int_data_res_4__2__5_), .A2(
        npu_inst_pe_1_3_2_n1), .B1(npu_inst_pe_1_3_2_N78), .B2(
        npu_inst_pe_1_3_2_n76), .C1(npu_inst_pe_1_3_2_N70), .C2(
        npu_inst_pe_1_3_2_n77), .ZN(npu_inst_pe_1_3_2_n79) );
  INV_X1 npu_inst_pe_1_3_2_U38 ( .A(npu_inst_pe_1_3_2_n79), .ZN(
        npu_inst_pe_1_3_2_n35) );
  AOI222_X1 npu_inst_pe_1_3_2_U37 ( .A1(npu_inst_int_data_res_4__2__6_), .A2(
        npu_inst_pe_1_3_2_n1), .B1(npu_inst_pe_1_3_2_N79), .B2(
        npu_inst_pe_1_3_2_n76), .C1(npu_inst_pe_1_3_2_N71), .C2(
        npu_inst_pe_1_3_2_n77), .ZN(npu_inst_pe_1_3_2_n78) );
  INV_X1 npu_inst_pe_1_3_2_U36 ( .A(npu_inst_pe_1_3_2_n78), .ZN(
        npu_inst_pe_1_3_2_n34) );
  INV_X1 npu_inst_pe_1_3_2_U35 ( .A(npu_inst_pe_1_3_2_int_data_1_), .ZN(
        npu_inst_pe_1_3_2_n14) );
  AND2_X1 npu_inst_pe_1_3_2_U34 ( .A1(npu_inst_int_data_x_3__2__1_), .A2(
        npu_inst_pe_1_3_2_int_q_weight_1_), .ZN(npu_inst_pe_1_3_2_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_3_2_U33 ( .A1(npu_inst_int_data_x_3__2__0_), .A2(
        npu_inst_pe_1_3_2_int_q_weight_1_), .ZN(npu_inst_pe_1_3_2_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_3_2_U32 ( .A1(npu_inst_n57), .A2(
        npu_inst_int_data_y_4__2__1_), .B1(npu_inst_pe_1_3_2_n3), .B2(
        npu_inst_int_data_x_3__3__1_), .ZN(npu_inst_pe_1_3_2_n63) );
  AOI22_X1 npu_inst_pe_1_3_2_U31 ( .A1(npu_inst_n57), .A2(
        npu_inst_int_data_y_4__2__0_), .B1(npu_inst_pe_1_3_2_n3), .B2(
        npu_inst_int_data_x_3__3__0_), .ZN(npu_inst_pe_1_3_2_n61) );
  INV_X1 npu_inst_pe_1_3_2_U30 ( .A(npu_inst_pe_1_3_2_int_data_0_), .ZN(
        npu_inst_pe_1_3_2_n13) );
  INV_X1 npu_inst_pe_1_3_2_U29 ( .A(npu_inst_n70), .ZN(npu_inst_pe_1_3_2_n5)
         );
  OR3_X1 npu_inst_pe_1_3_2_U28 ( .A1(npu_inst_pe_1_3_2_n6), .A2(
        npu_inst_pe_1_3_2_n8), .A3(npu_inst_pe_1_3_2_n5), .ZN(
        npu_inst_pe_1_3_2_n56) );
  OR3_X1 npu_inst_pe_1_3_2_U27 ( .A1(npu_inst_pe_1_3_2_n5), .A2(
        npu_inst_pe_1_3_2_n8), .A3(npu_inst_pe_1_3_2_n7), .ZN(
        npu_inst_pe_1_3_2_n48) );
  INV_X1 npu_inst_pe_1_3_2_U26 ( .A(npu_inst_pe_1_3_2_n5), .ZN(
        npu_inst_pe_1_3_2_n4) );
  INV_X1 npu_inst_pe_1_3_2_U25 ( .A(npu_inst_n125), .ZN(npu_inst_pe_1_3_2_n12)
         );
  OR3_X1 npu_inst_pe_1_3_2_U24 ( .A1(npu_inst_pe_1_3_2_n4), .A2(
        npu_inst_pe_1_3_2_n8), .A3(npu_inst_pe_1_3_2_n7), .ZN(
        npu_inst_pe_1_3_2_n52) );
  OR3_X1 npu_inst_pe_1_3_2_U23 ( .A1(npu_inst_pe_1_3_2_n6), .A2(
        npu_inst_pe_1_3_2_n8), .A3(npu_inst_pe_1_3_2_n4), .ZN(
        npu_inst_pe_1_3_2_n60) );
  NOR2_X1 npu_inst_pe_1_3_2_U22 ( .A1(npu_inst_pe_1_3_2_n60), .A2(
        npu_inst_pe_1_3_2_n3), .ZN(npu_inst_pe_1_3_2_n58) );
  NOR2_X1 npu_inst_pe_1_3_2_U21 ( .A1(npu_inst_pe_1_3_2_n56), .A2(
        npu_inst_pe_1_3_2_n3), .ZN(npu_inst_pe_1_3_2_n54) );
  NOR2_X1 npu_inst_pe_1_3_2_U20 ( .A1(npu_inst_pe_1_3_2_n52), .A2(
        npu_inst_pe_1_3_2_n3), .ZN(npu_inst_pe_1_3_2_n50) );
  NOR2_X1 npu_inst_pe_1_3_2_U19 ( .A1(npu_inst_pe_1_3_2_n48), .A2(
        npu_inst_pe_1_3_2_n3), .ZN(npu_inst_pe_1_3_2_n46) );
  NOR2_X1 npu_inst_pe_1_3_2_U18 ( .A1(npu_inst_pe_1_3_2_n40), .A2(
        npu_inst_pe_1_3_2_n3), .ZN(npu_inst_pe_1_3_2_n38) );
  NOR2_X1 npu_inst_pe_1_3_2_U17 ( .A1(npu_inst_pe_1_3_2_n44), .A2(
        npu_inst_pe_1_3_2_n3), .ZN(npu_inst_pe_1_3_2_n42) );
  BUF_X1 npu_inst_pe_1_3_2_U16 ( .A(npu_inst_n101), .Z(npu_inst_pe_1_3_2_n8)
         );
  BUF_X1 npu_inst_pe_1_3_2_U15 ( .A(npu_inst_pe_1_3_2_n12), .Z(
        npu_inst_pe_1_3_2_n11) );
  BUF_X1 npu_inst_pe_1_3_2_U14 ( .A(npu_inst_pe_1_3_2_n12), .Z(
        npu_inst_pe_1_3_2_n10) );
  BUF_X1 npu_inst_pe_1_3_2_U13 ( .A(npu_inst_pe_1_3_2_n12), .Z(
        npu_inst_pe_1_3_2_n9) );
  INV_X1 npu_inst_pe_1_3_2_U12 ( .A(npu_inst_pe_1_3_2_n38), .ZN(
        npu_inst_pe_1_3_2_n118) );
  INV_X1 npu_inst_pe_1_3_2_U11 ( .A(npu_inst_pe_1_3_2_n58), .ZN(
        npu_inst_pe_1_3_2_n114) );
  INV_X1 npu_inst_pe_1_3_2_U10 ( .A(npu_inst_pe_1_3_2_n54), .ZN(
        npu_inst_pe_1_3_2_n115) );
  INV_X1 npu_inst_pe_1_3_2_U9 ( .A(npu_inst_pe_1_3_2_n50), .ZN(
        npu_inst_pe_1_3_2_n116) );
  INV_X1 npu_inst_pe_1_3_2_U8 ( .A(npu_inst_pe_1_3_2_n46), .ZN(
        npu_inst_pe_1_3_2_n117) );
  INV_X1 npu_inst_pe_1_3_2_U7 ( .A(npu_inst_pe_1_3_2_n42), .ZN(
        npu_inst_pe_1_3_2_n119) );
  BUF_X1 npu_inst_pe_1_3_2_U6 ( .A(npu_inst_n25), .Z(npu_inst_pe_1_3_2_n2) );
  BUF_X1 npu_inst_pe_1_3_2_U5 ( .A(npu_inst_n25), .Z(npu_inst_pe_1_3_2_n1) );
  NOR2_X1 npu_inst_pe_1_3_2_U4 ( .A1(npu_inst_pe_1_3_2_int_q_weight_0_), .A2(
        npu_inst_pe_1_3_2_n1), .ZN(npu_inst_pe_1_3_2_n76) );
  NOR2_X1 npu_inst_pe_1_3_2_U3 ( .A1(npu_inst_pe_1_3_2_n27), .A2(
        npu_inst_pe_1_3_2_n1), .ZN(npu_inst_pe_1_3_2_n77) );
  FA_X1 npu_inst_pe_1_3_2_sub_77_U2_1 ( .A(npu_inst_pe_1_3_2_int_q_acc_1_), 
        .B(npu_inst_pe_1_3_2_n14), .CI(npu_inst_pe_1_3_2_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_3_2_sub_77_carry_2_), .S(npu_inst_pe_1_3_2_N66) );
  FA_X1 npu_inst_pe_1_3_2_add_79_U1_1 ( .A(npu_inst_pe_1_3_2_int_q_acc_1_), 
        .B(npu_inst_pe_1_3_2_int_data_1_), .CI(
        npu_inst_pe_1_3_2_add_79_carry_1_), .CO(
        npu_inst_pe_1_3_2_add_79_carry_2_), .S(npu_inst_pe_1_3_2_N74) );
  NAND3_X1 npu_inst_pe_1_3_2_U109 ( .A1(npu_inst_pe_1_3_2_n5), .A2(
        npu_inst_pe_1_3_2_n7), .A3(npu_inst_pe_1_3_2_n8), .ZN(
        npu_inst_pe_1_3_2_n44) );
  NAND3_X1 npu_inst_pe_1_3_2_U108 ( .A1(npu_inst_pe_1_3_2_n4), .A2(
        npu_inst_pe_1_3_2_n7), .A3(npu_inst_pe_1_3_2_n8), .ZN(
        npu_inst_pe_1_3_2_n40) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_3_2_n34), .CK(
        npu_inst_pe_1_3_2_net3695), .RN(npu_inst_pe_1_3_2_n9), .Q(
        npu_inst_pe_1_3_2_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_3_2_n35), .CK(
        npu_inst_pe_1_3_2_net3695), .RN(npu_inst_pe_1_3_2_n9), .Q(
        npu_inst_pe_1_3_2_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_3_2_n36), .CK(
        npu_inst_pe_1_3_2_net3695), .RN(npu_inst_pe_1_3_2_n9), .Q(
        npu_inst_pe_1_3_2_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_3_2_n98), .CK(
        npu_inst_pe_1_3_2_net3695), .RN(npu_inst_pe_1_3_2_n9), .Q(
        npu_inst_pe_1_3_2_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_3_2_n99), .CK(
        npu_inst_pe_1_3_2_net3695), .RN(npu_inst_pe_1_3_2_n9), .Q(
        npu_inst_pe_1_3_2_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_3_2_n100), 
        .CK(npu_inst_pe_1_3_2_net3695), .RN(npu_inst_pe_1_3_2_n9), .Q(
        npu_inst_pe_1_3_2_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_3_2_n33), .CK(
        npu_inst_pe_1_3_2_net3695), .RN(npu_inst_pe_1_3_2_n9), .Q(
        npu_inst_pe_1_3_2_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_3_2_n101), 
        .CK(npu_inst_pe_1_3_2_net3695), .RN(npu_inst_pe_1_3_2_n9), .Q(
        npu_inst_pe_1_3_2_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_weight_reg_0_ ( .D(npu_inst_n111), .CK(
        npu_inst_pe_1_3_2_net3701), .RN(npu_inst_pe_1_3_2_n9), .Q(
        npu_inst_pe_1_3_2_int_q_weight_0_), .QN(npu_inst_pe_1_3_2_n27) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_weight_reg_1_ ( .D(npu_inst_n117), .CK(
        npu_inst_pe_1_3_2_net3701), .RN(npu_inst_pe_1_3_2_n9), .Q(
        npu_inst_pe_1_3_2_int_q_weight_1_), .QN(npu_inst_pe_1_3_2_n26) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_3_2_n113), 
        .CK(npu_inst_pe_1_3_2_net3701), .RN(npu_inst_pe_1_3_2_n9), .Q(
        npu_inst_pe_1_3_2_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_3_2_n107), 
        .CK(npu_inst_pe_1_3_2_net3701), .RN(npu_inst_pe_1_3_2_n9), .Q(
        npu_inst_pe_1_3_2_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_3_2_n112), 
        .CK(npu_inst_pe_1_3_2_net3701), .RN(npu_inst_pe_1_3_2_n10), .Q(
        npu_inst_pe_1_3_2_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_3_2_n106), 
        .CK(npu_inst_pe_1_3_2_net3701), .RN(npu_inst_pe_1_3_2_n10), .Q(
        npu_inst_pe_1_3_2_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_3_2_n111), 
        .CK(npu_inst_pe_1_3_2_net3701), .RN(npu_inst_pe_1_3_2_n10), .Q(
        npu_inst_pe_1_3_2_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_3_2_n105), 
        .CK(npu_inst_pe_1_3_2_net3701), .RN(npu_inst_pe_1_3_2_n10), .Q(
        npu_inst_pe_1_3_2_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_3_2_n110), 
        .CK(npu_inst_pe_1_3_2_net3701), .RN(npu_inst_pe_1_3_2_n10), .Q(
        npu_inst_pe_1_3_2_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_3_2_n104), 
        .CK(npu_inst_pe_1_3_2_net3701), .RN(npu_inst_pe_1_3_2_n10), .Q(
        npu_inst_pe_1_3_2_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_3_2_n109), 
        .CK(npu_inst_pe_1_3_2_net3701), .RN(npu_inst_pe_1_3_2_n10), .Q(
        npu_inst_pe_1_3_2_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_3_2_n103), 
        .CK(npu_inst_pe_1_3_2_net3701), .RN(npu_inst_pe_1_3_2_n10), .Q(
        npu_inst_pe_1_3_2_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_3_2_n108), 
        .CK(npu_inst_pe_1_3_2_net3701), .RN(npu_inst_pe_1_3_2_n10), .Q(
        npu_inst_pe_1_3_2_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_3_2_n102), 
        .CK(npu_inst_pe_1_3_2_net3701), .RN(npu_inst_pe_1_3_2_n10), .Q(
        npu_inst_pe_1_3_2_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_3_2_n86), 
        .CK(npu_inst_pe_1_3_2_net3701), .RN(npu_inst_pe_1_3_2_n10), .Q(
        npu_inst_pe_1_3_2_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_3_2_n87), 
        .CK(npu_inst_pe_1_3_2_net3701), .RN(npu_inst_pe_1_3_2_n10), .Q(
        npu_inst_pe_1_3_2_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_3_2_n88), 
        .CK(npu_inst_pe_1_3_2_net3701), .RN(npu_inst_pe_1_3_2_n11), .Q(
        npu_inst_pe_1_3_2_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_3_2_n89), 
        .CK(npu_inst_pe_1_3_2_net3701), .RN(npu_inst_pe_1_3_2_n11), .Q(
        npu_inst_pe_1_3_2_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_3_2_n90), 
        .CK(npu_inst_pe_1_3_2_net3701), .RN(npu_inst_pe_1_3_2_n11), .Q(
        npu_inst_pe_1_3_2_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_3_2_n91), 
        .CK(npu_inst_pe_1_3_2_net3701), .RN(npu_inst_pe_1_3_2_n11), .Q(
        npu_inst_pe_1_3_2_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_3_2_n92), 
        .CK(npu_inst_pe_1_3_2_net3701), .RN(npu_inst_pe_1_3_2_n11), .Q(
        npu_inst_pe_1_3_2_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_3_2_n93), 
        .CK(npu_inst_pe_1_3_2_net3701), .RN(npu_inst_pe_1_3_2_n11), .Q(
        npu_inst_pe_1_3_2_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_3_2_n94), 
        .CK(npu_inst_pe_1_3_2_net3701), .RN(npu_inst_pe_1_3_2_n11), .Q(
        npu_inst_pe_1_3_2_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_3_2_n95), 
        .CK(npu_inst_pe_1_3_2_net3701), .RN(npu_inst_pe_1_3_2_n11), .Q(
        npu_inst_pe_1_3_2_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_3_2_n96), 
        .CK(npu_inst_pe_1_3_2_net3701), .RN(npu_inst_pe_1_3_2_n11), .Q(
        npu_inst_pe_1_3_2_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_3_2_n97), 
        .CK(npu_inst_pe_1_3_2_net3701), .RN(npu_inst_pe_1_3_2_n11), .Q(
        npu_inst_pe_1_3_2_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_3_2_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_3_2_N84), .SE(1'b0), .GCK(npu_inst_pe_1_3_2_net3695) );
  CLKGATETST_X1 npu_inst_pe_1_3_2_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n64), .SE(1'b0), .GCK(npu_inst_pe_1_3_2_net3701) );
  MUX2_X1 npu_inst_pe_1_3_3_U162 ( .A(npu_inst_pe_1_3_3_n32), .B(
        npu_inst_pe_1_3_3_n29), .S(npu_inst_pe_1_3_3_n8), .Z(
        npu_inst_pe_1_3_3_N93) );
  MUX2_X1 npu_inst_pe_1_3_3_U161 ( .A(npu_inst_pe_1_3_3_n31), .B(
        npu_inst_pe_1_3_3_n30), .S(npu_inst_pe_1_3_3_n6), .Z(
        npu_inst_pe_1_3_3_n32) );
  MUX2_X1 npu_inst_pe_1_3_3_U160 ( .A(npu_inst_pe_1_3_3_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_3_3_int_q_reg_v_1__0_), .S(npu_inst_pe_1_3_3_n4), .Z(
        npu_inst_pe_1_3_3_n31) );
  MUX2_X1 npu_inst_pe_1_3_3_U159 ( .A(npu_inst_pe_1_3_3_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_3_3_int_q_reg_v_3__0_), .S(npu_inst_pe_1_3_3_n4), .Z(
        npu_inst_pe_1_3_3_n30) );
  MUX2_X1 npu_inst_pe_1_3_3_U158 ( .A(npu_inst_pe_1_3_3_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_3_3_int_q_reg_v_5__0_), .S(npu_inst_pe_1_3_3_n4), .Z(
        npu_inst_pe_1_3_3_n29) );
  MUX2_X1 npu_inst_pe_1_3_3_U157 ( .A(npu_inst_pe_1_3_3_n28), .B(
        npu_inst_pe_1_3_3_n23), .S(npu_inst_pe_1_3_3_n8), .Z(
        npu_inst_pe_1_3_3_N94) );
  MUX2_X1 npu_inst_pe_1_3_3_U156 ( .A(npu_inst_pe_1_3_3_n25), .B(
        npu_inst_pe_1_3_3_n24), .S(npu_inst_pe_1_3_3_n6), .Z(
        npu_inst_pe_1_3_3_n28) );
  MUX2_X1 npu_inst_pe_1_3_3_U155 ( .A(npu_inst_pe_1_3_3_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_3_3_int_q_reg_v_1__1_), .S(npu_inst_pe_1_3_3_n4), .Z(
        npu_inst_pe_1_3_3_n25) );
  MUX2_X1 npu_inst_pe_1_3_3_U154 ( .A(npu_inst_pe_1_3_3_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_3_3_int_q_reg_v_3__1_), .S(npu_inst_pe_1_3_3_n4), .Z(
        npu_inst_pe_1_3_3_n24) );
  MUX2_X1 npu_inst_pe_1_3_3_U153 ( .A(npu_inst_pe_1_3_3_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_3_3_int_q_reg_v_5__1_), .S(npu_inst_pe_1_3_3_n4), .Z(
        npu_inst_pe_1_3_3_n23) );
  MUX2_X1 npu_inst_pe_1_3_3_U152 ( .A(npu_inst_pe_1_3_3_n22), .B(
        npu_inst_pe_1_3_3_n19), .S(npu_inst_pe_1_3_3_n8), .Z(
        npu_inst_int_data_x_3__3__1_) );
  MUX2_X1 npu_inst_pe_1_3_3_U151 ( .A(npu_inst_pe_1_3_3_n21), .B(
        npu_inst_pe_1_3_3_n20), .S(npu_inst_pe_1_3_3_n6), .Z(
        npu_inst_pe_1_3_3_n22) );
  MUX2_X1 npu_inst_pe_1_3_3_U150 ( .A(npu_inst_pe_1_3_3_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_3_3_int_q_reg_h_1__1_), .S(npu_inst_pe_1_3_3_n4), .Z(
        npu_inst_pe_1_3_3_n21) );
  MUX2_X1 npu_inst_pe_1_3_3_U149 ( .A(npu_inst_pe_1_3_3_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_3_3_int_q_reg_h_3__1_), .S(npu_inst_pe_1_3_3_n4), .Z(
        npu_inst_pe_1_3_3_n20) );
  MUX2_X1 npu_inst_pe_1_3_3_U148 ( .A(npu_inst_pe_1_3_3_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_3_3_int_q_reg_h_5__1_), .S(npu_inst_pe_1_3_3_n4), .Z(
        npu_inst_pe_1_3_3_n19) );
  MUX2_X1 npu_inst_pe_1_3_3_U147 ( .A(npu_inst_pe_1_3_3_n18), .B(
        npu_inst_pe_1_3_3_n15), .S(npu_inst_pe_1_3_3_n8), .Z(
        npu_inst_int_data_x_3__3__0_) );
  MUX2_X1 npu_inst_pe_1_3_3_U146 ( .A(npu_inst_pe_1_3_3_n17), .B(
        npu_inst_pe_1_3_3_n16), .S(npu_inst_pe_1_3_3_n6), .Z(
        npu_inst_pe_1_3_3_n18) );
  MUX2_X1 npu_inst_pe_1_3_3_U145 ( .A(npu_inst_pe_1_3_3_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_3_3_int_q_reg_h_1__0_), .S(npu_inst_pe_1_3_3_n4), .Z(
        npu_inst_pe_1_3_3_n17) );
  MUX2_X1 npu_inst_pe_1_3_3_U144 ( .A(npu_inst_pe_1_3_3_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_3_3_int_q_reg_h_3__0_), .S(npu_inst_pe_1_3_3_n4), .Z(
        npu_inst_pe_1_3_3_n16) );
  MUX2_X1 npu_inst_pe_1_3_3_U143 ( .A(npu_inst_pe_1_3_3_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_3_3_int_q_reg_h_5__0_), .S(npu_inst_pe_1_3_3_n4), .Z(
        npu_inst_pe_1_3_3_n15) );
  XOR2_X1 npu_inst_pe_1_3_3_U142 ( .A(npu_inst_pe_1_3_3_int_data_0_), .B(
        npu_inst_pe_1_3_3_int_q_acc_0_), .Z(npu_inst_pe_1_3_3_N73) );
  AND2_X1 npu_inst_pe_1_3_3_U141 ( .A1(npu_inst_pe_1_3_3_int_q_acc_0_), .A2(
        npu_inst_pe_1_3_3_int_data_0_), .ZN(npu_inst_pe_1_3_3_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_3_3_U140 ( .A(npu_inst_pe_1_3_3_int_q_acc_0_), .B(
        npu_inst_pe_1_3_3_n13), .ZN(npu_inst_pe_1_3_3_N65) );
  OR2_X1 npu_inst_pe_1_3_3_U139 ( .A1(npu_inst_pe_1_3_3_n13), .A2(
        npu_inst_pe_1_3_3_int_q_acc_0_), .ZN(npu_inst_pe_1_3_3_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_3_3_U138 ( .A(npu_inst_pe_1_3_3_int_q_acc_2_), .B(
        npu_inst_pe_1_3_3_add_79_carry_2_), .Z(npu_inst_pe_1_3_3_N75) );
  AND2_X1 npu_inst_pe_1_3_3_U137 ( .A1(npu_inst_pe_1_3_3_add_79_carry_2_), 
        .A2(npu_inst_pe_1_3_3_int_q_acc_2_), .ZN(
        npu_inst_pe_1_3_3_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_3_3_U136 ( .A(npu_inst_pe_1_3_3_int_q_acc_3_), .B(
        npu_inst_pe_1_3_3_add_79_carry_3_), .Z(npu_inst_pe_1_3_3_N76) );
  AND2_X1 npu_inst_pe_1_3_3_U135 ( .A1(npu_inst_pe_1_3_3_add_79_carry_3_), 
        .A2(npu_inst_pe_1_3_3_int_q_acc_3_), .ZN(
        npu_inst_pe_1_3_3_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_3_3_U134 ( .A(npu_inst_pe_1_3_3_int_q_acc_4_), .B(
        npu_inst_pe_1_3_3_add_79_carry_4_), .Z(npu_inst_pe_1_3_3_N77) );
  AND2_X1 npu_inst_pe_1_3_3_U133 ( .A1(npu_inst_pe_1_3_3_add_79_carry_4_), 
        .A2(npu_inst_pe_1_3_3_int_q_acc_4_), .ZN(
        npu_inst_pe_1_3_3_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_3_3_U132 ( .A(npu_inst_pe_1_3_3_int_q_acc_5_), .B(
        npu_inst_pe_1_3_3_add_79_carry_5_), .Z(npu_inst_pe_1_3_3_N78) );
  AND2_X1 npu_inst_pe_1_3_3_U131 ( .A1(npu_inst_pe_1_3_3_add_79_carry_5_), 
        .A2(npu_inst_pe_1_3_3_int_q_acc_5_), .ZN(
        npu_inst_pe_1_3_3_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_3_3_U130 ( .A(npu_inst_pe_1_3_3_int_q_acc_6_), .B(
        npu_inst_pe_1_3_3_add_79_carry_6_), .Z(npu_inst_pe_1_3_3_N79) );
  AND2_X1 npu_inst_pe_1_3_3_U129 ( .A1(npu_inst_pe_1_3_3_add_79_carry_6_), 
        .A2(npu_inst_pe_1_3_3_int_q_acc_6_), .ZN(
        npu_inst_pe_1_3_3_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_3_3_U128 ( .A(npu_inst_pe_1_3_3_int_q_acc_7_), .B(
        npu_inst_pe_1_3_3_add_79_carry_7_), .Z(npu_inst_pe_1_3_3_N80) );
  XNOR2_X1 npu_inst_pe_1_3_3_U127 ( .A(npu_inst_pe_1_3_3_sub_77_carry_2_), .B(
        npu_inst_pe_1_3_3_int_q_acc_2_), .ZN(npu_inst_pe_1_3_3_N67) );
  OR2_X1 npu_inst_pe_1_3_3_U126 ( .A1(npu_inst_pe_1_3_3_int_q_acc_2_), .A2(
        npu_inst_pe_1_3_3_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_3_3_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_3_3_U125 ( .A(npu_inst_pe_1_3_3_sub_77_carry_3_), .B(
        npu_inst_pe_1_3_3_int_q_acc_3_), .ZN(npu_inst_pe_1_3_3_N68) );
  OR2_X1 npu_inst_pe_1_3_3_U124 ( .A1(npu_inst_pe_1_3_3_int_q_acc_3_), .A2(
        npu_inst_pe_1_3_3_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_3_3_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_3_3_U123 ( .A(npu_inst_pe_1_3_3_sub_77_carry_4_), .B(
        npu_inst_pe_1_3_3_int_q_acc_4_), .ZN(npu_inst_pe_1_3_3_N69) );
  OR2_X1 npu_inst_pe_1_3_3_U122 ( .A1(npu_inst_pe_1_3_3_int_q_acc_4_), .A2(
        npu_inst_pe_1_3_3_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_3_3_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_3_3_U121 ( .A(npu_inst_pe_1_3_3_sub_77_carry_5_), .B(
        npu_inst_pe_1_3_3_int_q_acc_5_), .ZN(npu_inst_pe_1_3_3_N70) );
  OR2_X1 npu_inst_pe_1_3_3_U120 ( .A1(npu_inst_pe_1_3_3_int_q_acc_5_), .A2(
        npu_inst_pe_1_3_3_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_3_3_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_3_3_U119 ( .A(npu_inst_pe_1_3_3_sub_77_carry_6_), .B(
        npu_inst_pe_1_3_3_int_q_acc_6_), .ZN(npu_inst_pe_1_3_3_N71) );
  OR2_X1 npu_inst_pe_1_3_3_U118 ( .A1(npu_inst_pe_1_3_3_int_q_acc_6_), .A2(
        npu_inst_pe_1_3_3_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_3_3_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_3_3_U117 ( .A(npu_inst_pe_1_3_3_int_q_acc_7_), .B(
        npu_inst_pe_1_3_3_sub_77_carry_7_), .ZN(npu_inst_pe_1_3_3_N72) );
  INV_X1 npu_inst_pe_1_3_3_U116 ( .A(npu_inst_n78), .ZN(npu_inst_pe_1_3_3_n7)
         );
  INV_X1 npu_inst_pe_1_3_3_U115 ( .A(npu_inst_pe_1_3_3_n7), .ZN(
        npu_inst_pe_1_3_3_n6) );
  INV_X1 npu_inst_pe_1_3_3_U114 ( .A(npu_inst_n57), .ZN(npu_inst_pe_1_3_3_n3)
         );
  AOI22_X1 npu_inst_pe_1_3_3_U113 ( .A1(npu_inst_int_data_y_4__3__0_), .A2(
        npu_inst_pe_1_3_3_n58), .B1(npu_inst_pe_1_3_3_n114), .B2(
        npu_inst_pe_1_3_3_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_3_3_n57) );
  INV_X1 npu_inst_pe_1_3_3_U112 ( .A(npu_inst_pe_1_3_3_n57), .ZN(
        npu_inst_pe_1_3_3_n108) );
  AOI22_X1 npu_inst_pe_1_3_3_U111 ( .A1(npu_inst_int_data_y_4__3__0_), .A2(
        npu_inst_pe_1_3_3_n54), .B1(npu_inst_pe_1_3_3_n115), .B2(
        npu_inst_pe_1_3_3_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_3_3_n53) );
  INV_X1 npu_inst_pe_1_3_3_U110 ( .A(npu_inst_pe_1_3_3_n53), .ZN(
        npu_inst_pe_1_3_3_n109) );
  AOI22_X1 npu_inst_pe_1_3_3_U107 ( .A1(npu_inst_int_data_y_4__3__0_), .A2(
        npu_inst_pe_1_3_3_n50), .B1(npu_inst_pe_1_3_3_n116), .B2(
        npu_inst_pe_1_3_3_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_3_3_n49) );
  INV_X1 npu_inst_pe_1_3_3_U106 ( .A(npu_inst_pe_1_3_3_n49), .ZN(
        npu_inst_pe_1_3_3_n110) );
  AOI22_X1 npu_inst_pe_1_3_3_U105 ( .A1(npu_inst_int_data_y_4__3__0_), .A2(
        npu_inst_pe_1_3_3_n46), .B1(npu_inst_pe_1_3_3_n117), .B2(
        npu_inst_pe_1_3_3_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_3_3_n45) );
  INV_X1 npu_inst_pe_1_3_3_U104 ( .A(npu_inst_pe_1_3_3_n45), .ZN(
        npu_inst_pe_1_3_3_n111) );
  AOI22_X1 npu_inst_pe_1_3_3_U103 ( .A1(npu_inst_int_data_y_4__3__0_), .A2(
        npu_inst_pe_1_3_3_n42), .B1(npu_inst_pe_1_3_3_n119), .B2(
        npu_inst_pe_1_3_3_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_3_3_n41) );
  INV_X1 npu_inst_pe_1_3_3_U102 ( .A(npu_inst_pe_1_3_3_n41), .ZN(
        npu_inst_pe_1_3_3_n112) );
  AOI22_X1 npu_inst_pe_1_3_3_U101 ( .A1(npu_inst_int_data_y_4__3__1_), .A2(
        npu_inst_pe_1_3_3_n58), .B1(npu_inst_pe_1_3_3_n114), .B2(
        npu_inst_pe_1_3_3_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_3_3_n59) );
  INV_X1 npu_inst_pe_1_3_3_U100 ( .A(npu_inst_pe_1_3_3_n59), .ZN(
        npu_inst_pe_1_3_3_n102) );
  AOI22_X1 npu_inst_pe_1_3_3_U99 ( .A1(npu_inst_int_data_y_4__3__1_), .A2(
        npu_inst_pe_1_3_3_n54), .B1(npu_inst_pe_1_3_3_n115), .B2(
        npu_inst_pe_1_3_3_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_3_3_n55) );
  INV_X1 npu_inst_pe_1_3_3_U98 ( .A(npu_inst_pe_1_3_3_n55), .ZN(
        npu_inst_pe_1_3_3_n103) );
  AOI22_X1 npu_inst_pe_1_3_3_U97 ( .A1(npu_inst_int_data_y_4__3__1_), .A2(
        npu_inst_pe_1_3_3_n50), .B1(npu_inst_pe_1_3_3_n116), .B2(
        npu_inst_pe_1_3_3_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_3_3_n51) );
  INV_X1 npu_inst_pe_1_3_3_U96 ( .A(npu_inst_pe_1_3_3_n51), .ZN(
        npu_inst_pe_1_3_3_n104) );
  AOI22_X1 npu_inst_pe_1_3_3_U95 ( .A1(npu_inst_int_data_y_4__3__1_), .A2(
        npu_inst_pe_1_3_3_n46), .B1(npu_inst_pe_1_3_3_n117), .B2(
        npu_inst_pe_1_3_3_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_3_3_n47) );
  INV_X1 npu_inst_pe_1_3_3_U94 ( .A(npu_inst_pe_1_3_3_n47), .ZN(
        npu_inst_pe_1_3_3_n105) );
  AOI22_X1 npu_inst_pe_1_3_3_U93 ( .A1(npu_inst_int_data_y_4__3__1_), .A2(
        npu_inst_pe_1_3_3_n42), .B1(npu_inst_pe_1_3_3_n119), .B2(
        npu_inst_pe_1_3_3_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_3_3_n43) );
  INV_X1 npu_inst_pe_1_3_3_U92 ( .A(npu_inst_pe_1_3_3_n43), .ZN(
        npu_inst_pe_1_3_3_n106) );
  AOI22_X1 npu_inst_pe_1_3_3_U91 ( .A1(npu_inst_pe_1_3_3_n38), .A2(
        npu_inst_int_data_y_4__3__1_), .B1(npu_inst_pe_1_3_3_n118), .B2(
        npu_inst_pe_1_3_3_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_3_3_n39) );
  INV_X1 npu_inst_pe_1_3_3_U90 ( .A(npu_inst_pe_1_3_3_n39), .ZN(
        npu_inst_pe_1_3_3_n107) );
  AOI22_X1 npu_inst_pe_1_3_3_U89 ( .A1(npu_inst_pe_1_3_3_n38), .A2(
        npu_inst_int_data_y_4__3__0_), .B1(npu_inst_pe_1_3_3_n118), .B2(
        npu_inst_pe_1_3_3_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_3_3_n37) );
  INV_X1 npu_inst_pe_1_3_3_U88 ( .A(npu_inst_pe_1_3_3_n37), .ZN(
        npu_inst_pe_1_3_3_n113) );
  NAND2_X1 npu_inst_pe_1_3_3_U87 ( .A1(npu_inst_pe_1_3_3_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_3_3_n60), .ZN(npu_inst_pe_1_3_3_n74) );
  OAI21_X1 npu_inst_pe_1_3_3_U86 ( .B1(npu_inst_pe_1_3_3_n63), .B2(
        npu_inst_pe_1_3_3_n60), .A(npu_inst_pe_1_3_3_n74), .ZN(
        npu_inst_pe_1_3_3_n97) );
  NAND2_X1 npu_inst_pe_1_3_3_U85 ( .A1(npu_inst_pe_1_3_3_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_3_3_n60), .ZN(npu_inst_pe_1_3_3_n73) );
  OAI21_X1 npu_inst_pe_1_3_3_U84 ( .B1(npu_inst_pe_1_3_3_n61), .B2(
        npu_inst_pe_1_3_3_n60), .A(npu_inst_pe_1_3_3_n73), .ZN(
        npu_inst_pe_1_3_3_n96) );
  NAND2_X1 npu_inst_pe_1_3_3_U83 ( .A1(npu_inst_pe_1_3_3_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_3_3_n56), .ZN(npu_inst_pe_1_3_3_n72) );
  OAI21_X1 npu_inst_pe_1_3_3_U82 ( .B1(npu_inst_pe_1_3_3_n63), .B2(
        npu_inst_pe_1_3_3_n56), .A(npu_inst_pe_1_3_3_n72), .ZN(
        npu_inst_pe_1_3_3_n95) );
  NAND2_X1 npu_inst_pe_1_3_3_U81 ( .A1(npu_inst_pe_1_3_3_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_3_3_n56), .ZN(npu_inst_pe_1_3_3_n71) );
  OAI21_X1 npu_inst_pe_1_3_3_U80 ( .B1(npu_inst_pe_1_3_3_n61), .B2(
        npu_inst_pe_1_3_3_n56), .A(npu_inst_pe_1_3_3_n71), .ZN(
        npu_inst_pe_1_3_3_n94) );
  NAND2_X1 npu_inst_pe_1_3_3_U79 ( .A1(npu_inst_pe_1_3_3_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_3_3_n52), .ZN(npu_inst_pe_1_3_3_n70) );
  OAI21_X1 npu_inst_pe_1_3_3_U78 ( .B1(npu_inst_pe_1_3_3_n63), .B2(
        npu_inst_pe_1_3_3_n52), .A(npu_inst_pe_1_3_3_n70), .ZN(
        npu_inst_pe_1_3_3_n93) );
  NAND2_X1 npu_inst_pe_1_3_3_U77 ( .A1(npu_inst_pe_1_3_3_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_3_3_n52), .ZN(npu_inst_pe_1_3_3_n69) );
  OAI21_X1 npu_inst_pe_1_3_3_U76 ( .B1(npu_inst_pe_1_3_3_n61), .B2(
        npu_inst_pe_1_3_3_n52), .A(npu_inst_pe_1_3_3_n69), .ZN(
        npu_inst_pe_1_3_3_n92) );
  NAND2_X1 npu_inst_pe_1_3_3_U75 ( .A1(npu_inst_pe_1_3_3_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_3_3_n48), .ZN(npu_inst_pe_1_3_3_n68) );
  OAI21_X1 npu_inst_pe_1_3_3_U74 ( .B1(npu_inst_pe_1_3_3_n63), .B2(
        npu_inst_pe_1_3_3_n48), .A(npu_inst_pe_1_3_3_n68), .ZN(
        npu_inst_pe_1_3_3_n91) );
  NAND2_X1 npu_inst_pe_1_3_3_U73 ( .A1(npu_inst_pe_1_3_3_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_3_3_n48), .ZN(npu_inst_pe_1_3_3_n67) );
  OAI21_X1 npu_inst_pe_1_3_3_U72 ( .B1(npu_inst_pe_1_3_3_n61), .B2(
        npu_inst_pe_1_3_3_n48), .A(npu_inst_pe_1_3_3_n67), .ZN(
        npu_inst_pe_1_3_3_n90) );
  NAND2_X1 npu_inst_pe_1_3_3_U71 ( .A1(npu_inst_pe_1_3_3_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_3_3_n44), .ZN(npu_inst_pe_1_3_3_n66) );
  OAI21_X1 npu_inst_pe_1_3_3_U70 ( .B1(npu_inst_pe_1_3_3_n63), .B2(
        npu_inst_pe_1_3_3_n44), .A(npu_inst_pe_1_3_3_n66), .ZN(
        npu_inst_pe_1_3_3_n89) );
  NAND2_X1 npu_inst_pe_1_3_3_U69 ( .A1(npu_inst_pe_1_3_3_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_3_3_n44), .ZN(npu_inst_pe_1_3_3_n65) );
  OAI21_X1 npu_inst_pe_1_3_3_U68 ( .B1(npu_inst_pe_1_3_3_n61), .B2(
        npu_inst_pe_1_3_3_n44), .A(npu_inst_pe_1_3_3_n65), .ZN(
        npu_inst_pe_1_3_3_n88) );
  NAND2_X1 npu_inst_pe_1_3_3_U67 ( .A1(npu_inst_pe_1_3_3_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_3_3_n40), .ZN(npu_inst_pe_1_3_3_n64) );
  OAI21_X1 npu_inst_pe_1_3_3_U66 ( .B1(npu_inst_pe_1_3_3_n63), .B2(
        npu_inst_pe_1_3_3_n40), .A(npu_inst_pe_1_3_3_n64), .ZN(
        npu_inst_pe_1_3_3_n87) );
  NAND2_X1 npu_inst_pe_1_3_3_U65 ( .A1(npu_inst_pe_1_3_3_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_3_3_n40), .ZN(npu_inst_pe_1_3_3_n62) );
  OAI21_X1 npu_inst_pe_1_3_3_U64 ( .B1(npu_inst_pe_1_3_3_n61), .B2(
        npu_inst_pe_1_3_3_n40), .A(npu_inst_pe_1_3_3_n62), .ZN(
        npu_inst_pe_1_3_3_n86) );
  AND2_X1 npu_inst_pe_1_3_3_U63 ( .A1(npu_inst_pe_1_3_3_N93), .A2(npu_inst_n57), .ZN(npu_inst_int_data_y_3__3__0_) );
  AND2_X1 npu_inst_pe_1_3_3_U62 ( .A1(npu_inst_n57), .A2(npu_inst_pe_1_3_3_N94), .ZN(npu_inst_int_data_y_3__3__1_) );
  NOR3_X1 npu_inst_pe_1_3_3_U61 ( .A1(npu_inst_pe_1_3_3_n26), .A2(npu_inst_n57), .A3(npu_inst_int_ckg[36]), .ZN(npu_inst_pe_1_3_3_n85) );
  OR2_X1 npu_inst_pe_1_3_3_U60 ( .A1(npu_inst_pe_1_3_3_n85), .A2(
        npu_inst_pe_1_3_3_n2), .ZN(npu_inst_pe_1_3_3_N84) );
  AND2_X1 npu_inst_pe_1_3_3_U59 ( .A1(npu_inst_pe_1_3_3_int_q_acc_0_), .A2(
        npu_inst_pe_1_3_3_n1), .ZN(npu_inst_int_data_res_3__3__0_) );
  AND2_X1 npu_inst_pe_1_3_3_U58 ( .A1(npu_inst_pe_1_3_3_n2), .A2(
        npu_inst_pe_1_3_3_int_q_acc_7_), .ZN(npu_inst_int_data_res_3__3__7_)
         );
  AND2_X1 npu_inst_pe_1_3_3_U57 ( .A1(npu_inst_pe_1_3_3_int_q_acc_1_), .A2(
        npu_inst_pe_1_3_3_n1), .ZN(npu_inst_int_data_res_3__3__1_) );
  AND2_X1 npu_inst_pe_1_3_3_U56 ( .A1(npu_inst_pe_1_3_3_int_q_acc_2_), .A2(
        npu_inst_pe_1_3_3_n1), .ZN(npu_inst_int_data_res_3__3__2_) );
  AND2_X1 npu_inst_pe_1_3_3_U55 ( .A1(npu_inst_pe_1_3_3_int_q_acc_3_), .A2(
        npu_inst_pe_1_3_3_n2), .ZN(npu_inst_int_data_res_3__3__3_) );
  AND2_X1 npu_inst_pe_1_3_3_U54 ( .A1(npu_inst_pe_1_3_3_int_q_acc_4_), .A2(
        npu_inst_pe_1_3_3_n2), .ZN(npu_inst_int_data_res_3__3__4_) );
  AND2_X1 npu_inst_pe_1_3_3_U53 ( .A1(npu_inst_pe_1_3_3_int_q_acc_5_), .A2(
        npu_inst_pe_1_3_3_n2), .ZN(npu_inst_int_data_res_3__3__5_) );
  AND2_X1 npu_inst_pe_1_3_3_U52 ( .A1(npu_inst_pe_1_3_3_int_q_acc_6_), .A2(
        npu_inst_pe_1_3_3_n2), .ZN(npu_inst_int_data_res_3__3__6_) );
  AOI222_X1 npu_inst_pe_1_3_3_U51 ( .A1(npu_inst_int_data_res_4__3__0_), .A2(
        npu_inst_pe_1_3_3_n1), .B1(npu_inst_pe_1_3_3_N73), .B2(
        npu_inst_pe_1_3_3_n76), .C1(npu_inst_pe_1_3_3_N65), .C2(
        npu_inst_pe_1_3_3_n77), .ZN(npu_inst_pe_1_3_3_n84) );
  INV_X1 npu_inst_pe_1_3_3_U50 ( .A(npu_inst_pe_1_3_3_n84), .ZN(
        npu_inst_pe_1_3_3_n101) );
  AOI222_X1 npu_inst_pe_1_3_3_U49 ( .A1(npu_inst_int_data_res_4__3__7_), .A2(
        npu_inst_pe_1_3_3_n1), .B1(npu_inst_pe_1_3_3_N80), .B2(
        npu_inst_pe_1_3_3_n76), .C1(npu_inst_pe_1_3_3_N72), .C2(
        npu_inst_pe_1_3_3_n77), .ZN(npu_inst_pe_1_3_3_n75) );
  INV_X1 npu_inst_pe_1_3_3_U48 ( .A(npu_inst_pe_1_3_3_n75), .ZN(
        npu_inst_pe_1_3_3_n33) );
  AOI222_X1 npu_inst_pe_1_3_3_U47 ( .A1(npu_inst_int_data_res_4__3__1_), .A2(
        npu_inst_pe_1_3_3_n1), .B1(npu_inst_pe_1_3_3_N74), .B2(
        npu_inst_pe_1_3_3_n76), .C1(npu_inst_pe_1_3_3_N66), .C2(
        npu_inst_pe_1_3_3_n77), .ZN(npu_inst_pe_1_3_3_n83) );
  INV_X1 npu_inst_pe_1_3_3_U46 ( .A(npu_inst_pe_1_3_3_n83), .ZN(
        npu_inst_pe_1_3_3_n100) );
  AOI222_X1 npu_inst_pe_1_3_3_U45 ( .A1(npu_inst_int_data_res_4__3__2_), .A2(
        npu_inst_pe_1_3_3_n1), .B1(npu_inst_pe_1_3_3_N75), .B2(
        npu_inst_pe_1_3_3_n76), .C1(npu_inst_pe_1_3_3_N67), .C2(
        npu_inst_pe_1_3_3_n77), .ZN(npu_inst_pe_1_3_3_n82) );
  INV_X1 npu_inst_pe_1_3_3_U44 ( .A(npu_inst_pe_1_3_3_n82), .ZN(
        npu_inst_pe_1_3_3_n99) );
  AOI222_X1 npu_inst_pe_1_3_3_U43 ( .A1(npu_inst_int_data_res_4__3__3_), .A2(
        npu_inst_pe_1_3_3_n1), .B1(npu_inst_pe_1_3_3_N76), .B2(
        npu_inst_pe_1_3_3_n76), .C1(npu_inst_pe_1_3_3_N68), .C2(
        npu_inst_pe_1_3_3_n77), .ZN(npu_inst_pe_1_3_3_n81) );
  INV_X1 npu_inst_pe_1_3_3_U42 ( .A(npu_inst_pe_1_3_3_n81), .ZN(
        npu_inst_pe_1_3_3_n98) );
  AOI222_X1 npu_inst_pe_1_3_3_U41 ( .A1(npu_inst_int_data_res_4__3__4_), .A2(
        npu_inst_pe_1_3_3_n1), .B1(npu_inst_pe_1_3_3_N77), .B2(
        npu_inst_pe_1_3_3_n76), .C1(npu_inst_pe_1_3_3_N69), .C2(
        npu_inst_pe_1_3_3_n77), .ZN(npu_inst_pe_1_3_3_n80) );
  INV_X1 npu_inst_pe_1_3_3_U40 ( .A(npu_inst_pe_1_3_3_n80), .ZN(
        npu_inst_pe_1_3_3_n36) );
  AOI222_X1 npu_inst_pe_1_3_3_U39 ( .A1(npu_inst_int_data_res_4__3__5_), .A2(
        npu_inst_pe_1_3_3_n1), .B1(npu_inst_pe_1_3_3_N78), .B2(
        npu_inst_pe_1_3_3_n76), .C1(npu_inst_pe_1_3_3_N70), .C2(
        npu_inst_pe_1_3_3_n77), .ZN(npu_inst_pe_1_3_3_n79) );
  INV_X1 npu_inst_pe_1_3_3_U38 ( .A(npu_inst_pe_1_3_3_n79), .ZN(
        npu_inst_pe_1_3_3_n35) );
  AOI222_X1 npu_inst_pe_1_3_3_U37 ( .A1(npu_inst_int_data_res_4__3__6_), .A2(
        npu_inst_pe_1_3_3_n1), .B1(npu_inst_pe_1_3_3_N79), .B2(
        npu_inst_pe_1_3_3_n76), .C1(npu_inst_pe_1_3_3_N71), .C2(
        npu_inst_pe_1_3_3_n77), .ZN(npu_inst_pe_1_3_3_n78) );
  INV_X1 npu_inst_pe_1_3_3_U36 ( .A(npu_inst_pe_1_3_3_n78), .ZN(
        npu_inst_pe_1_3_3_n34) );
  INV_X1 npu_inst_pe_1_3_3_U35 ( .A(npu_inst_pe_1_3_3_int_data_1_), .ZN(
        npu_inst_pe_1_3_3_n14) );
  AND2_X1 npu_inst_pe_1_3_3_U34 ( .A1(npu_inst_int_data_x_3__3__1_), .A2(
        npu_inst_pe_1_3_3_int_q_weight_1_), .ZN(npu_inst_pe_1_3_3_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_3_3_U33 ( .A1(npu_inst_int_data_x_3__3__0_), .A2(
        npu_inst_pe_1_3_3_int_q_weight_1_), .ZN(npu_inst_pe_1_3_3_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_3_3_U32 ( .A1(npu_inst_n57), .A2(
        npu_inst_int_data_y_4__3__1_), .B1(npu_inst_pe_1_3_3_n3), .B2(
        npu_inst_int_data_x_3__4__1_), .ZN(npu_inst_pe_1_3_3_n63) );
  AOI22_X1 npu_inst_pe_1_3_3_U31 ( .A1(npu_inst_n57), .A2(
        npu_inst_int_data_y_4__3__0_), .B1(npu_inst_pe_1_3_3_n3), .B2(
        npu_inst_int_data_x_3__4__0_), .ZN(npu_inst_pe_1_3_3_n61) );
  INV_X1 npu_inst_pe_1_3_3_U30 ( .A(npu_inst_pe_1_3_3_int_data_0_), .ZN(
        npu_inst_pe_1_3_3_n13) );
  INV_X1 npu_inst_pe_1_3_3_U29 ( .A(npu_inst_n70), .ZN(npu_inst_pe_1_3_3_n5)
         );
  OR3_X1 npu_inst_pe_1_3_3_U28 ( .A1(npu_inst_pe_1_3_3_n6), .A2(
        npu_inst_pe_1_3_3_n8), .A3(npu_inst_pe_1_3_3_n5), .ZN(
        npu_inst_pe_1_3_3_n56) );
  OR3_X1 npu_inst_pe_1_3_3_U27 ( .A1(npu_inst_pe_1_3_3_n5), .A2(
        npu_inst_pe_1_3_3_n8), .A3(npu_inst_pe_1_3_3_n7), .ZN(
        npu_inst_pe_1_3_3_n48) );
  INV_X1 npu_inst_pe_1_3_3_U26 ( .A(npu_inst_pe_1_3_3_n5), .ZN(
        npu_inst_pe_1_3_3_n4) );
  INV_X1 npu_inst_pe_1_3_3_U25 ( .A(npu_inst_n125), .ZN(npu_inst_pe_1_3_3_n12)
         );
  OR3_X1 npu_inst_pe_1_3_3_U24 ( .A1(npu_inst_pe_1_3_3_n4), .A2(
        npu_inst_pe_1_3_3_n8), .A3(npu_inst_pe_1_3_3_n7), .ZN(
        npu_inst_pe_1_3_3_n52) );
  OR3_X1 npu_inst_pe_1_3_3_U23 ( .A1(npu_inst_pe_1_3_3_n6), .A2(
        npu_inst_pe_1_3_3_n8), .A3(npu_inst_pe_1_3_3_n4), .ZN(
        npu_inst_pe_1_3_3_n60) );
  NOR2_X1 npu_inst_pe_1_3_3_U22 ( .A1(npu_inst_pe_1_3_3_n60), .A2(
        npu_inst_pe_1_3_3_n3), .ZN(npu_inst_pe_1_3_3_n58) );
  NOR2_X1 npu_inst_pe_1_3_3_U21 ( .A1(npu_inst_pe_1_3_3_n56), .A2(
        npu_inst_pe_1_3_3_n3), .ZN(npu_inst_pe_1_3_3_n54) );
  NOR2_X1 npu_inst_pe_1_3_3_U20 ( .A1(npu_inst_pe_1_3_3_n52), .A2(
        npu_inst_pe_1_3_3_n3), .ZN(npu_inst_pe_1_3_3_n50) );
  NOR2_X1 npu_inst_pe_1_3_3_U19 ( .A1(npu_inst_pe_1_3_3_n48), .A2(
        npu_inst_pe_1_3_3_n3), .ZN(npu_inst_pe_1_3_3_n46) );
  NOR2_X1 npu_inst_pe_1_3_3_U18 ( .A1(npu_inst_pe_1_3_3_n40), .A2(
        npu_inst_pe_1_3_3_n3), .ZN(npu_inst_pe_1_3_3_n38) );
  NOR2_X1 npu_inst_pe_1_3_3_U17 ( .A1(npu_inst_pe_1_3_3_n44), .A2(
        npu_inst_pe_1_3_3_n3), .ZN(npu_inst_pe_1_3_3_n42) );
  BUF_X1 npu_inst_pe_1_3_3_U16 ( .A(npu_inst_n101), .Z(npu_inst_pe_1_3_3_n8)
         );
  BUF_X1 npu_inst_pe_1_3_3_U15 ( .A(npu_inst_pe_1_3_3_n12), .Z(
        npu_inst_pe_1_3_3_n11) );
  BUF_X1 npu_inst_pe_1_3_3_U14 ( .A(npu_inst_pe_1_3_3_n12), .Z(
        npu_inst_pe_1_3_3_n10) );
  BUF_X1 npu_inst_pe_1_3_3_U13 ( .A(npu_inst_pe_1_3_3_n12), .Z(
        npu_inst_pe_1_3_3_n9) );
  INV_X1 npu_inst_pe_1_3_3_U12 ( .A(npu_inst_pe_1_3_3_n38), .ZN(
        npu_inst_pe_1_3_3_n118) );
  INV_X1 npu_inst_pe_1_3_3_U11 ( .A(npu_inst_pe_1_3_3_n58), .ZN(
        npu_inst_pe_1_3_3_n114) );
  INV_X1 npu_inst_pe_1_3_3_U10 ( .A(npu_inst_pe_1_3_3_n54), .ZN(
        npu_inst_pe_1_3_3_n115) );
  INV_X1 npu_inst_pe_1_3_3_U9 ( .A(npu_inst_pe_1_3_3_n50), .ZN(
        npu_inst_pe_1_3_3_n116) );
  INV_X1 npu_inst_pe_1_3_3_U8 ( .A(npu_inst_pe_1_3_3_n46), .ZN(
        npu_inst_pe_1_3_3_n117) );
  INV_X1 npu_inst_pe_1_3_3_U7 ( .A(npu_inst_pe_1_3_3_n42), .ZN(
        npu_inst_pe_1_3_3_n119) );
  BUF_X1 npu_inst_pe_1_3_3_U6 ( .A(npu_inst_n25), .Z(npu_inst_pe_1_3_3_n2) );
  BUF_X1 npu_inst_pe_1_3_3_U5 ( .A(npu_inst_n25), .Z(npu_inst_pe_1_3_3_n1) );
  NOR2_X1 npu_inst_pe_1_3_3_U4 ( .A1(npu_inst_pe_1_3_3_int_q_weight_0_), .A2(
        npu_inst_pe_1_3_3_n1), .ZN(npu_inst_pe_1_3_3_n76) );
  NOR2_X1 npu_inst_pe_1_3_3_U3 ( .A1(npu_inst_pe_1_3_3_n27), .A2(
        npu_inst_pe_1_3_3_n1), .ZN(npu_inst_pe_1_3_3_n77) );
  FA_X1 npu_inst_pe_1_3_3_sub_77_U2_1 ( .A(npu_inst_pe_1_3_3_int_q_acc_1_), 
        .B(npu_inst_pe_1_3_3_n14), .CI(npu_inst_pe_1_3_3_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_3_3_sub_77_carry_2_), .S(npu_inst_pe_1_3_3_N66) );
  FA_X1 npu_inst_pe_1_3_3_add_79_U1_1 ( .A(npu_inst_pe_1_3_3_int_q_acc_1_), 
        .B(npu_inst_pe_1_3_3_int_data_1_), .CI(
        npu_inst_pe_1_3_3_add_79_carry_1_), .CO(
        npu_inst_pe_1_3_3_add_79_carry_2_), .S(npu_inst_pe_1_3_3_N74) );
  NAND3_X1 npu_inst_pe_1_3_3_U109 ( .A1(npu_inst_pe_1_3_3_n5), .A2(
        npu_inst_pe_1_3_3_n7), .A3(npu_inst_pe_1_3_3_n8), .ZN(
        npu_inst_pe_1_3_3_n44) );
  NAND3_X1 npu_inst_pe_1_3_3_U108 ( .A1(npu_inst_pe_1_3_3_n4), .A2(
        npu_inst_pe_1_3_3_n7), .A3(npu_inst_pe_1_3_3_n8), .ZN(
        npu_inst_pe_1_3_3_n40) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_3_3_n34), .CK(
        npu_inst_pe_1_3_3_net3672), .RN(npu_inst_pe_1_3_3_n9), .Q(
        npu_inst_pe_1_3_3_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_3_3_n35), .CK(
        npu_inst_pe_1_3_3_net3672), .RN(npu_inst_pe_1_3_3_n9), .Q(
        npu_inst_pe_1_3_3_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_3_3_n36), .CK(
        npu_inst_pe_1_3_3_net3672), .RN(npu_inst_pe_1_3_3_n9), .Q(
        npu_inst_pe_1_3_3_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_3_3_n98), .CK(
        npu_inst_pe_1_3_3_net3672), .RN(npu_inst_pe_1_3_3_n9), .Q(
        npu_inst_pe_1_3_3_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_3_3_n99), .CK(
        npu_inst_pe_1_3_3_net3672), .RN(npu_inst_pe_1_3_3_n9), .Q(
        npu_inst_pe_1_3_3_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_3_3_n100), 
        .CK(npu_inst_pe_1_3_3_net3672), .RN(npu_inst_pe_1_3_3_n9), .Q(
        npu_inst_pe_1_3_3_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_3_3_n33), .CK(
        npu_inst_pe_1_3_3_net3672), .RN(npu_inst_pe_1_3_3_n9), .Q(
        npu_inst_pe_1_3_3_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_3_3_n101), 
        .CK(npu_inst_pe_1_3_3_net3672), .RN(npu_inst_pe_1_3_3_n9), .Q(
        npu_inst_pe_1_3_3_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_weight_reg_0_ ( .D(npu_inst_n111), .CK(
        npu_inst_pe_1_3_3_net3678), .RN(npu_inst_pe_1_3_3_n9), .Q(
        npu_inst_pe_1_3_3_int_q_weight_0_), .QN(npu_inst_pe_1_3_3_n27) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_weight_reg_1_ ( .D(npu_inst_n117), .CK(
        npu_inst_pe_1_3_3_net3678), .RN(npu_inst_pe_1_3_3_n9), .Q(
        npu_inst_pe_1_3_3_int_q_weight_1_), .QN(npu_inst_pe_1_3_3_n26) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_3_3_n113), 
        .CK(npu_inst_pe_1_3_3_net3678), .RN(npu_inst_pe_1_3_3_n9), .Q(
        npu_inst_pe_1_3_3_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_3_3_n107), 
        .CK(npu_inst_pe_1_3_3_net3678), .RN(npu_inst_pe_1_3_3_n9), .Q(
        npu_inst_pe_1_3_3_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_3_3_n112), 
        .CK(npu_inst_pe_1_3_3_net3678), .RN(npu_inst_pe_1_3_3_n10), .Q(
        npu_inst_pe_1_3_3_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_3_3_n106), 
        .CK(npu_inst_pe_1_3_3_net3678), .RN(npu_inst_pe_1_3_3_n10), .Q(
        npu_inst_pe_1_3_3_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_3_3_n111), 
        .CK(npu_inst_pe_1_3_3_net3678), .RN(npu_inst_pe_1_3_3_n10), .Q(
        npu_inst_pe_1_3_3_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_3_3_n105), 
        .CK(npu_inst_pe_1_3_3_net3678), .RN(npu_inst_pe_1_3_3_n10), .Q(
        npu_inst_pe_1_3_3_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_3_3_n110), 
        .CK(npu_inst_pe_1_3_3_net3678), .RN(npu_inst_pe_1_3_3_n10), .Q(
        npu_inst_pe_1_3_3_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_3_3_n104), 
        .CK(npu_inst_pe_1_3_3_net3678), .RN(npu_inst_pe_1_3_3_n10), .Q(
        npu_inst_pe_1_3_3_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_3_3_n109), 
        .CK(npu_inst_pe_1_3_3_net3678), .RN(npu_inst_pe_1_3_3_n10), .Q(
        npu_inst_pe_1_3_3_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_3_3_n103), 
        .CK(npu_inst_pe_1_3_3_net3678), .RN(npu_inst_pe_1_3_3_n10), .Q(
        npu_inst_pe_1_3_3_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_3_3_n108), 
        .CK(npu_inst_pe_1_3_3_net3678), .RN(npu_inst_pe_1_3_3_n10), .Q(
        npu_inst_pe_1_3_3_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_3_3_n102), 
        .CK(npu_inst_pe_1_3_3_net3678), .RN(npu_inst_pe_1_3_3_n10), .Q(
        npu_inst_pe_1_3_3_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_3_3_n86), 
        .CK(npu_inst_pe_1_3_3_net3678), .RN(npu_inst_pe_1_3_3_n10), .Q(
        npu_inst_pe_1_3_3_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_3_3_n87), 
        .CK(npu_inst_pe_1_3_3_net3678), .RN(npu_inst_pe_1_3_3_n10), .Q(
        npu_inst_pe_1_3_3_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_3_3_n88), 
        .CK(npu_inst_pe_1_3_3_net3678), .RN(npu_inst_pe_1_3_3_n11), .Q(
        npu_inst_pe_1_3_3_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_3_3_n89), 
        .CK(npu_inst_pe_1_3_3_net3678), .RN(npu_inst_pe_1_3_3_n11), .Q(
        npu_inst_pe_1_3_3_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_3_3_n90), 
        .CK(npu_inst_pe_1_3_3_net3678), .RN(npu_inst_pe_1_3_3_n11), .Q(
        npu_inst_pe_1_3_3_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_3_3_n91), 
        .CK(npu_inst_pe_1_3_3_net3678), .RN(npu_inst_pe_1_3_3_n11), .Q(
        npu_inst_pe_1_3_3_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_3_3_n92), 
        .CK(npu_inst_pe_1_3_3_net3678), .RN(npu_inst_pe_1_3_3_n11), .Q(
        npu_inst_pe_1_3_3_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_3_3_n93), 
        .CK(npu_inst_pe_1_3_3_net3678), .RN(npu_inst_pe_1_3_3_n11), .Q(
        npu_inst_pe_1_3_3_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_3_3_n94), 
        .CK(npu_inst_pe_1_3_3_net3678), .RN(npu_inst_pe_1_3_3_n11), .Q(
        npu_inst_pe_1_3_3_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_3_3_n95), 
        .CK(npu_inst_pe_1_3_3_net3678), .RN(npu_inst_pe_1_3_3_n11), .Q(
        npu_inst_pe_1_3_3_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_3_3_n96), 
        .CK(npu_inst_pe_1_3_3_net3678), .RN(npu_inst_pe_1_3_3_n11), .Q(
        npu_inst_pe_1_3_3_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_3_3_n97), 
        .CK(npu_inst_pe_1_3_3_net3678), .RN(npu_inst_pe_1_3_3_n11), .Q(
        npu_inst_pe_1_3_3_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_3_3_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_3_3_N84), .SE(1'b0), .GCK(npu_inst_pe_1_3_3_net3672) );
  CLKGATETST_X1 npu_inst_pe_1_3_3_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n64), .SE(1'b0), .GCK(npu_inst_pe_1_3_3_net3678) );
  MUX2_X1 npu_inst_pe_1_3_4_U161 ( .A(npu_inst_pe_1_3_4_n31), .B(
        npu_inst_pe_1_3_4_n28), .S(npu_inst_pe_1_3_4_n7), .Z(
        npu_inst_pe_1_3_4_N93) );
  MUX2_X1 npu_inst_pe_1_3_4_U160 ( .A(npu_inst_pe_1_3_4_n30), .B(
        npu_inst_pe_1_3_4_n29), .S(npu_inst_n77), .Z(npu_inst_pe_1_3_4_n31) );
  MUX2_X1 npu_inst_pe_1_3_4_U159 ( .A(npu_inst_pe_1_3_4_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_3_4_int_q_reg_v_1__0_), .S(npu_inst_pe_1_3_4_n4), .Z(
        npu_inst_pe_1_3_4_n30) );
  MUX2_X1 npu_inst_pe_1_3_4_U158 ( .A(npu_inst_pe_1_3_4_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_3_4_int_q_reg_v_3__0_), .S(npu_inst_pe_1_3_4_n4), .Z(
        npu_inst_pe_1_3_4_n29) );
  MUX2_X1 npu_inst_pe_1_3_4_U157 ( .A(npu_inst_pe_1_3_4_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_3_4_int_q_reg_v_5__0_), .S(npu_inst_pe_1_3_4_n4), .Z(
        npu_inst_pe_1_3_4_n28) );
  MUX2_X1 npu_inst_pe_1_3_4_U156 ( .A(npu_inst_pe_1_3_4_n25), .B(
        npu_inst_pe_1_3_4_n22), .S(npu_inst_pe_1_3_4_n7), .Z(
        npu_inst_pe_1_3_4_N94) );
  MUX2_X1 npu_inst_pe_1_3_4_U155 ( .A(npu_inst_pe_1_3_4_n24), .B(
        npu_inst_pe_1_3_4_n23), .S(npu_inst_n77), .Z(npu_inst_pe_1_3_4_n25) );
  MUX2_X1 npu_inst_pe_1_3_4_U154 ( .A(npu_inst_pe_1_3_4_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_3_4_int_q_reg_v_1__1_), .S(npu_inst_pe_1_3_4_n4), .Z(
        npu_inst_pe_1_3_4_n24) );
  MUX2_X1 npu_inst_pe_1_3_4_U153 ( .A(npu_inst_pe_1_3_4_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_3_4_int_q_reg_v_3__1_), .S(npu_inst_pe_1_3_4_n4), .Z(
        npu_inst_pe_1_3_4_n23) );
  MUX2_X1 npu_inst_pe_1_3_4_U152 ( .A(npu_inst_pe_1_3_4_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_3_4_int_q_reg_v_5__1_), .S(npu_inst_pe_1_3_4_n4), .Z(
        npu_inst_pe_1_3_4_n22) );
  MUX2_X1 npu_inst_pe_1_3_4_U151 ( .A(npu_inst_pe_1_3_4_n21), .B(
        npu_inst_pe_1_3_4_n18), .S(npu_inst_pe_1_3_4_n7), .Z(
        npu_inst_int_data_x_3__4__1_) );
  MUX2_X1 npu_inst_pe_1_3_4_U150 ( .A(npu_inst_pe_1_3_4_n20), .B(
        npu_inst_pe_1_3_4_n19), .S(npu_inst_n77), .Z(npu_inst_pe_1_3_4_n21) );
  MUX2_X1 npu_inst_pe_1_3_4_U149 ( .A(npu_inst_pe_1_3_4_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_3_4_int_q_reg_h_1__1_), .S(npu_inst_pe_1_3_4_n4), .Z(
        npu_inst_pe_1_3_4_n20) );
  MUX2_X1 npu_inst_pe_1_3_4_U148 ( .A(npu_inst_pe_1_3_4_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_3_4_int_q_reg_h_3__1_), .S(npu_inst_pe_1_3_4_n4), .Z(
        npu_inst_pe_1_3_4_n19) );
  MUX2_X1 npu_inst_pe_1_3_4_U147 ( .A(npu_inst_pe_1_3_4_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_3_4_int_q_reg_h_5__1_), .S(npu_inst_pe_1_3_4_n4), .Z(
        npu_inst_pe_1_3_4_n18) );
  MUX2_X1 npu_inst_pe_1_3_4_U146 ( .A(npu_inst_pe_1_3_4_n17), .B(
        npu_inst_pe_1_3_4_n14), .S(npu_inst_pe_1_3_4_n7), .Z(
        npu_inst_int_data_x_3__4__0_) );
  MUX2_X1 npu_inst_pe_1_3_4_U145 ( .A(npu_inst_pe_1_3_4_n16), .B(
        npu_inst_pe_1_3_4_n15), .S(npu_inst_n77), .Z(npu_inst_pe_1_3_4_n17) );
  MUX2_X1 npu_inst_pe_1_3_4_U144 ( .A(npu_inst_pe_1_3_4_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_3_4_int_q_reg_h_1__0_), .S(npu_inst_pe_1_3_4_n4), .Z(
        npu_inst_pe_1_3_4_n16) );
  MUX2_X1 npu_inst_pe_1_3_4_U143 ( .A(npu_inst_pe_1_3_4_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_3_4_int_q_reg_h_3__0_), .S(npu_inst_pe_1_3_4_n4), .Z(
        npu_inst_pe_1_3_4_n15) );
  MUX2_X1 npu_inst_pe_1_3_4_U142 ( .A(npu_inst_pe_1_3_4_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_3_4_int_q_reg_h_5__0_), .S(npu_inst_pe_1_3_4_n4), .Z(
        npu_inst_pe_1_3_4_n14) );
  XOR2_X1 npu_inst_pe_1_3_4_U141 ( .A(npu_inst_pe_1_3_4_int_data_0_), .B(
        npu_inst_pe_1_3_4_int_q_acc_0_), .Z(npu_inst_pe_1_3_4_N73) );
  AND2_X1 npu_inst_pe_1_3_4_U140 ( .A1(npu_inst_pe_1_3_4_int_q_acc_0_), .A2(
        npu_inst_pe_1_3_4_int_data_0_), .ZN(npu_inst_pe_1_3_4_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_3_4_U139 ( .A(npu_inst_pe_1_3_4_int_q_acc_0_), .B(
        npu_inst_pe_1_3_4_n12), .ZN(npu_inst_pe_1_3_4_N65) );
  OR2_X1 npu_inst_pe_1_3_4_U138 ( .A1(npu_inst_pe_1_3_4_n12), .A2(
        npu_inst_pe_1_3_4_int_q_acc_0_), .ZN(npu_inst_pe_1_3_4_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_3_4_U137 ( .A(npu_inst_pe_1_3_4_int_q_acc_2_), .B(
        npu_inst_pe_1_3_4_add_79_carry_2_), .Z(npu_inst_pe_1_3_4_N75) );
  AND2_X1 npu_inst_pe_1_3_4_U136 ( .A1(npu_inst_pe_1_3_4_add_79_carry_2_), 
        .A2(npu_inst_pe_1_3_4_int_q_acc_2_), .ZN(
        npu_inst_pe_1_3_4_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_3_4_U135 ( .A(npu_inst_pe_1_3_4_int_q_acc_3_), .B(
        npu_inst_pe_1_3_4_add_79_carry_3_), .Z(npu_inst_pe_1_3_4_N76) );
  AND2_X1 npu_inst_pe_1_3_4_U134 ( .A1(npu_inst_pe_1_3_4_add_79_carry_3_), 
        .A2(npu_inst_pe_1_3_4_int_q_acc_3_), .ZN(
        npu_inst_pe_1_3_4_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_3_4_U133 ( .A(npu_inst_pe_1_3_4_int_q_acc_4_), .B(
        npu_inst_pe_1_3_4_add_79_carry_4_), .Z(npu_inst_pe_1_3_4_N77) );
  AND2_X1 npu_inst_pe_1_3_4_U132 ( .A1(npu_inst_pe_1_3_4_add_79_carry_4_), 
        .A2(npu_inst_pe_1_3_4_int_q_acc_4_), .ZN(
        npu_inst_pe_1_3_4_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_3_4_U131 ( .A(npu_inst_pe_1_3_4_int_q_acc_5_), .B(
        npu_inst_pe_1_3_4_add_79_carry_5_), .Z(npu_inst_pe_1_3_4_N78) );
  AND2_X1 npu_inst_pe_1_3_4_U130 ( .A1(npu_inst_pe_1_3_4_add_79_carry_5_), 
        .A2(npu_inst_pe_1_3_4_int_q_acc_5_), .ZN(
        npu_inst_pe_1_3_4_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_3_4_U129 ( .A(npu_inst_pe_1_3_4_int_q_acc_6_), .B(
        npu_inst_pe_1_3_4_add_79_carry_6_), .Z(npu_inst_pe_1_3_4_N79) );
  AND2_X1 npu_inst_pe_1_3_4_U128 ( .A1(npu_inst_pe_1_3_4_add_79_carry_6_), 
        .A2(npu_inst_pe_1_3_4_int_q_acc_6_), .ZN(
        npu_inst_pe_1_3_4_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_3_4_U127 ( .A(npu_inst_pe_1_3_4_int_q_acc_7_), .B(
        npu_inst_pe_1_3_4_add_79_carry_7_), .Z(npu_inst_pe_1_3_4_N80) );
  XNOR2_X1 npu_inst_pe_1_3_4_U126 ( .A(npu_inst_pe_1_3_4_sub_77_carry_2_), .B(
        npu_inst_pe_1_3_4_int_q_acc_2_), .ZN(npu_inst_pe_1_3_4_N67) );
  OR2_X1 npu_inst_pe_1_3_4_U125 ( .A1(npu_inst_pe_1_3_4_int_q_acc_2_), .A2(
        npu_inst_pe_1_3_4_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_3_4_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_3_4_U124 ( .A(npu_inst_pe_1_3_4_sub_77_carry_3_), .B(
        npu_inst_pe_1_3_4_int_q_acc_3_), .ZN(npu_inst_pe_1_3_4_N68) );
  OR2_X1 npu_inst_pe_1_3_4_U123 ( .A1(npu_inst_pe_1_3_4_int_q_acc_3_), .A2(
        npu_inst_pe_1_3_4_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_3_4_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_3_4_U122 ( .A(npu_inst_pe_1_3_4_sub_77_carry_4_), .B(
        npu_inst_pe_1_3_4_int_q_acc_4_), .ZN(npu_inst_pe_1_3_4_N69) );
  OR2_X1 npu_inst_pe_1_3_4_U121 ( .A1(npu_inst_pe_1_3_4_int_q_acc_4_), .A2(
        npu_inst_pe_1_3_4_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_3_4_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_3_4_U120 ( .A(npu_inst_pe_1_3_4_sub_77_carry_5_), .B(
        npu_inst_pe_1_3_4_int_q_acc_5_), .ZN(npu_inst_pe_1_3_4_N70) );
  OR2_X1 npu_inst_pe_1_3_4_U119 ( .A1(npu_inst_pe_1_3_4_int_q_acc_5_), .A2(
        npu_inst_pe_1_3_4_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_3_4_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_3_4_U118 ( .A(npu_inst_pe_1_3_4_sub_77_carry_6_), .B(
        npu_inst_pe_1_3_4_int_q_acc_6_), .ZN(npu_inst_pe_1_3_4_N71) );
  OR2_X1 npu_inst_pe_1_3_4_U117 ( .A1(npu_inst_pe_1_3_4_int_q_acc_6_), .A2(
        npu_inst_pe_1_3_4_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_3_4_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_3_4_U116 ( .A(npu_inst_pe_1_3_4_int_q_acc_7_), .B(
        npu_inst_pe_1_3_4_sub_77_carry_7_), .ZN(npu_inst_pe_1_3_4_N72) );
  INV_X1 npu_inst_pe_1_3_4_U115 ( .A(npu_inst_n77), .ZN(npu_inst_pe_1_3_4_n6)
         );
  INV_X1 npu_inst_pe_1_3_4_U114 ( .A(npu_inst_n57), .ZN(npu_inst_pe_1_3_4_n3)
         );
  AOI22_X1 npu_inst_pe_1_3_4_U113 ( .A1(npu_inst_int_data_y_4__4__0_), .A2(
        npu_inst_pe_1_3_4_n58), .B1(npu_inst_pe_1_3_4_n113), .B2(
        npu_inst_pe_1_3_4_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_3_4_n57) );
  INV_X1 npu_inst_pe_1_3_4_U112 ( .A(npu_inst_pe_1_3_4_n57), .ZN(
        npu_inst_pe_1_3_4_n107) );
  AOI22_X1 npu_inst_pe_1_3_4_U111 ( .A1(npu_inst_int_data_y_4__4__0_), .A2(
        npu_inst_pe_1_3_4_n54), .B1(npu_inst_pe_1_3_4_n114), .B2(
        npu_inst_pe_1_3_4_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_3_4_n53) );
  INV_X1 npu_inst_pe_1_3_4_U110 ( .A(npu_inst_pe_1_3_4_n53), .ZN(
        npu_inst_pe_1_3_4_n108) );
  AOI22_X1 npu_inst_pe_1_3_4_U107 ( .A1(npu_inst_int_data_y_4__4__0_), .A2(
        npu_inst_pe_1_3_4_n50), .B1(npu_inst_pe_1_3_4_n115), .B2(
        npu_inst_pe_1_3_4_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_3_4_n49) );
  INV_X1 npu_inst_pe_1_3_4_U106 ( .A(npu_inst_pe_1_3_4_n49), .ZN(
        npu_inst_pe_1_3_4_n109) );
  AOI22_X1 npu_inst_pe_1_3_4_U105 ( .A1(npu_inst_int_data_y_4__4__0_), .A2(
        npu_inst_pe_1_3_4_n46), .B1(npu_inst_pe_1_3_4_n116), .B2(
        npu_inst_pe_1_3_4_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_3_4_n45) );
  INV_X1 npu_inst_pe_1_3_4_U104 ( .A(npu_inst_pe_1_3_4_n45), .ZN(
        npu_inst_pe_1_3_4_n110) );
  AOI22_X1 npu_inst_pe_1_3_4_U103 ( .A1(npu_inst_int_data_y_4__4__0_), .A2(
        npu_inst_pe_1_3_4_n42), .B1(npu_inst_pe_1_3_4_n118), .B2(
        npu_inst_pe_1_3_4_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_3_4_n41) );
  INV_X1 npu_inst_pe_1_3_4_U102 ( .A(npu_inst_pe_1_3_4_n41), .ZN(
        npu_inst_pe_1_3_4_n111) );
  AOI22_X1 npu_inst_pe_1_3_4_U101 ( .A1(npu_inst_int_data_y_4__4__1_), .A2(
        npu_inst_pe_1_3_4_n58), .B1(npu_inst_pe_1_3_4_n113), .B2(
        npu_inst_pe_1_3_4_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_3_4_n59) );
  INV_X1 npu_inst_pe_1_3_4_U100 ( .A(npu_inst_pe_1_3_4_n59), .ZN(
        npu_inst_pe_1_3_4_n101) );
  AOI22_X1 npu_inst_pe_1_3_4_U99 ( .A1(npu_inst_int_data_y_4__4__1_), .A2(
        npu_inst_pe_1_3_4_n54), .B1(npu_inst_pe_1_3_4_n114), .B2(
        npu_inst_pe_1_3_4_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_3_4_n55) );
  INV_X1 npu_inst_pe_1_3_4_U98 ( .A(npu_inst_pe_1_3_4_n55), .ZN(
        npu_inst_pe_1_3_4_n102) );
  AOI22_X1 npu_inst_pe_1_3_4_U97 ( .A1(npu_inst_int_data_y_4__4__1_), .A2(
        npu_inst_pe_1_3_4_n50), .B1(npu_inst_pe_1_3_4_n115), .B2(
        npu_inst_pe_1_3_4_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_3_4_n51) );
  INV_X1 npu_inst_pe_1_3_4_U96 ( .A(npu_inst_pe_1_3_4_n51), .ZN(
        npu_inst_pe_1_3_4_n103) );
  AOI22_X1 npu_inst_pe_1_3_4_U95 ( .A1(npu_inst_int_data_y_4__4__1_), .A2(
        npu_inst_pe_1_3_4_n46), .B1(npu_inst_pe_1_3_4_n116), .B2(
        npu_inst_pe_1_3_4_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_3_4_n47) );
  INV_X1 npu_inst_pe_1_3_4_U94 ( .A(npu_inst_pe_1_3_4_n47), .ZN(
        npu_inst_pe_1_3_4_n104) );
  AOI22_X1 npu_inst_pe_1_3_4_U93 ( .A1(npu_inst_int_data_y_4__4__1_), .A2(
        npu_inst_pe_1_3_4_n42), .B1(npu_inst_pe_1_3_4_n118), .B2(
        npu_inst_pe_1_3_4_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_3_4_n43) );
  INV_X1 npu_inst_pe_1_3_4_U92 ( .A(npu_inst_pe_1_3_4_n43), .ZN(
        npu_inst_pe_1_3_4_n105) );
  AOI22_X1 npu_inst_pe_1_3_4_U91 ( .A1(npu_inst_pe_1_3_4_n38), .A2(
        npu_inst_int_data_y_4__4__1_), .B1(npu_inst_pe_1_3_4_n117), .B2(
        npu_inst_pe_1_3_4_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_3_4_n39) );
  INV_X1 npu_inst_pe_1_3_4_U90 ( .A(npu_inst_pe_1_3_4_n39), .ZN(
        npu_inst_pe_1_3_4_n106) );
  AOI22_X1 npu_inst_pe_1_3_4_U89 ( .A1(npu_inst_pe_1_3_4_n38), .A2(
        npu_inst_int_data_y_4__4__0_), .B1(npu_inst_pe_1_3_4_n117), .B2(
        npu_inst_pe_1_3_4_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_3_4_n37) );
  INV_X1 npu_inst_pe_1_3_4_U88 ( .A(npu_inst_pe_1_3_4_n37), .ZN(
        npu_inst_pe_1_3_4_n112) );
  NAND2_X1 npu_inst_pe_1_3_4_U87 ( .A1(npu_inst_pe_1_3_4_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_3_4_n60), .ZN(npu_inst_pe_1_3_4_n74) );
  OAI21_X1 npu_inst_pe_1_3_4_U86 ( .B1(npu_inst_pe_1_3_4_n63), .B2(
        npu_inst_pe_1_3_4_n60), .A(npu_inst_pe_1_3_4_n74), .ZN(
        npu_inst_pe_1_3_4_n97) );
  NAND2_X1 npu_inst_pe_1_3_4_U85 ( .A1(npu_inst_pe_1_3_4_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_3_4_n60), .ZN(npu_inst_pe_1_3_4_n73) );
  OAI21_X1 npu_inst_pe_1_3_4_U84 ( .B1(npu_inst_pe_1_3_4_n61), .B2(
        npu_inst_pe_1_3_4_n60), .A(npu_inst_pe_1_3_4_n73), .ZN(
        npu_inst_pe_1_3_4_n96) );
  NAND2_X1 npu_inst_pe_1_3_4_U83 ( .A1(npu_inst_pe_1_3_4_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_3_4_n56), .ZN(npu_inst_pe_1_3_4_n72) );
  OAI21_X1 npu_inst_pe_1_3_4_U82 ( .B1(npu_inst_pe_1_3_4_n63), .B2(
        npu_inst_pe_1_3_4_n56), .A(npu_inst_pe_1_3_4_n72), .ZN(
        npu_inst_pe_1_3_4_n95) );
  NAND2_X1 npu_inst_pe_1_3_4_U81 ( .A1(npu_inst_pe_1_3_4_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_3_4_n56), .ZN(npu_inst_pe_1_3_4_n71) );
  OAI21_X1 npu_inst_pe_1_3_4_U80 ( .B1(npu_inst_pe_1_3_4_n61), .B2(
        npu_inst_pe_1_3_4_n56), .A(npu_inst_pe_1_3_4_n71), .ZN(
        npu_inst_pe_1_3_4_n94) );
  NAND2_X1 npu_inst_pe_1_3_4_U79 ( .A1(npu_inst_pe_1_3_4_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_3_4_n52), .ZN(npu_inst_pe_1_3_4_n70) );
  OAI21_X1 npu_inst_pe_1_3_4_U78 ( .B1(npu_inst_pe_1_3_4_n63), .B2(
        npu_inst_pe_1_3_4_n52), .A(npu_inst_pe_1_3_4_n70), .ZN(
        npu_inst_pe_1_3_4_n93) );
  NAND2_X1 npu_inst_pe_1_3_4_U77 ( .A1(npu_inst_pe_1_3_4_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_3_4_n52), .ZN(npu_inst_pe_1_3_4_n69) );
  OAI21_X1 npu_inst_pe_1_3_4_U76 ( .B1(npu_inst_pe_1_3_4_n61), .B2(
        npu_inst_pe_1_3_4_n52), .A(npu_inst_pe_1_3_4_n69), .ZN(
        npu_inst_pe_1_3_4_n92) );
  NAND2_X1 npu_inst_pe_1_3_4_U75 ( .A1(npu_inst_pe_1_3_4_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_3_4_n48), .ZN(npu_inst_pe_1_3_4_n68) );
  OAI21_X1 npu_inst_pe_1_3_4_U74 ( .B1(npu_inst_pe_1_3_4_n63), .B2(
        npu_inst_pe_1_3_4_n48), .A(npu_inst_pe_1_3_4_n68), .ZN(
        npu_inst_pe_1_3_4_n91) );
  NAND2_X1 npu_inst_pe_1_3_4_U73 ( .A1(npu_inst_pe_1_3_4_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_3_4_n48), .ZN(npu_inst_pe_1_3_4_n67) );
  OAI21_X1 npu_inst_pe_1_3_4_U72 ( .B1(npu_inst_pe_1_3_4_n61), .B2(
        npu_inst_pe_1_3_4_n48), .A(npu_inst_pe_1_3_4_n67), .ZN(
        npu_inst_pe_1_3_4_n90) );
  NAND2_X1 npu_inst_pe_1_3_4_U71 ( .A1(npu_inst_pe_1_3_4_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_3_4_n44), .ZN(npu_inst_pe_1_3_4_n66) );
  OAI21_X1 npu_inst_pe_1_3_4_U70 ( .B1(npu_inst_pe_1_3_4_n63), .B2(
        npu_inst_pe_1_3_4_n44), .A(npu_inst_pe_1_3_4_n66), .ZN(
        npu_inst_pe_1_3_4_n89) );
  NAND2_X1 npu_inst_pe_1_3_4_U69 ( .A1(npu_inst_pe_1_3_4_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_3_4_n44), .ZN(npu_inst_pe_1_3_4_n65) );
  OAI21_X1 npu_inst_pe_1_3_4_U68 ( .B1(npu_inst_pe_1_3_4_n61), .B2(
        npu_inst_pe_1_3_4_n44), .A(npu_inst_pe_1_3_4_n65), .ZN(
        npu_inst_pe_1_3_4_n88) );
  NAND2_X1 npu_inst_pe_1_3_4_U67 ( .A1(npu_inst_pe_1_3_4_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_3_4_n40), .ZN(npu_inst_pe_1_3_4_n64) );
  OAI21_X1 npu_inst_pe_1_3_4_U66 ( .B1(npu_inst_pe_1_3_4_n63), .B2(
        npu_inst_pe_1_3_4_n40), .A(npu_inst_pe_1_3_4_n64), .ZN(
        npu_inst_pe_1_3_4_n87) );
  NAND2_X1 npu_inst_pe_1_3_4_U65 ( .A1(npu_inst_pe_1_3_4_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_3_4_n40), .ZN(npu_inst_pe_1_3_4_n62) );
  OAI21_X1 npu_inst_pe_1_3_4_U64 ( .B1(npu_inst_pe_1_3_4_n61), .B2(
        npu_inst_pe_1_3_4_n40), .A(npu_inst_pe_1_3_4_n62), .ZN(
        npu_inst_pe_1_3_4_n86) );
  AND2_X1 npu_inst_pe_1_3_4_U63 ( .A1(npu_inst_pe_1_3_4_N93), .A2(npu_inst_n57), .ZN(npu_inst_int_data_y_3__4__0_) );
  AND2_X1 npu_inst_pe_1_3_4_U62 ( .A1(npu_inst_n57), .A2(npu_inst_pe_1_3_4_N94), .ZN(npu_inst_int_data_y_3__4__1_) );
  NOR3_X1 npu_inst_pe_1_3_4_U61 ( .A1(npu_inst_pe_1_3_4_n26), .A2(npu_inst_n57), .A3(npu_inst_int_ckg[35]), .ZN(npu_inst_pe_1_3_4_n85) );
  OR2_X1 npu_inst_pe_1_3_4_U60 ( .A1(npu_inst_pe_1_3_4_n85), .A2(
        npu_inst_pe_1_3_4_n2), .ZN(npu_inst_pe_1_3_4_N84) );
  AND2_X1 npu_inst_pe_1_3_4_U59 ( .A1(npu_inst_pe_1_3_4_int_q_acc_0_), .A2(
        npu_inst_pe_1_3_4_n1), .ZN(npu_inst_int_data_res_3__4__0_) );
  AND2_X1 npu_inst_pe_1_3_4_U58 ( .A1(npu_inst_pe_1_3_4_n2), .A2(
        npu_inst_pe_1_3_4_int_q_acc_7_), .ZN(npu_inst_int_data_res_3__4__7_)
         );
  AND2_X1 npu_inst_pe_1_3_4_U57 ( .A1(npu_inst_pe_1_3_4_int_q_acc_1_), .A2(
        npu_inst_pe_1_3_4_n1), .ZN(npu_inst_int_data_res_3__4__1_) );
  AND2_X1 npu_inst_pe_1_3_4_U56 ( .A1(npu_inst_pe_1_3_4_int_q_acc_2_), .A2(
        npu_inst_pe_1_3_4_n1), .ZN(npu_inst_int_data_res_3__4__2_) );
  AND2_X1 npu_inst_pe_1_3_4_U55 ( .A1(npu_inst_pe_1_3_4_int_q_acc_3_), .A2(
        npu_inst_pe_1_3_4_n2), .ZN(npu_inst_int_data_res_3__4__3_) );
  AND2_X1 npu_inst_pe_1_3_4_U54 ( .A1(npu_inst_pe_1_3_4_int_q_acc_4_), .A2(
        npu_inst_pe_1_3_4_n2), .ZN(npu_inst_int_data_res_3__4__4_) );
  AND2_X1 npu_inst_pe_1_3_4_U53 ( .A1(npu_inst_pe_1_3_4_int_q_acc_5_), .A2(
        npu_inst_pe_1_3_4_n2), .ZN(npu_inst_int_data_res_3__4__5_) );
  AND2_X1 npu_inst_pe_1_3_4_U52 ( .A1(npu_inst_pe_1_3_4_int_q_acc_6_), .A2(
        npu_inst_pe_1_3_4_n2), .ZN(npu_inst_int_data_res_3__4__6_) );
  AOI222_X1 npu_inst_pe_1_3_4_U51 ( .A1(npu_inst_int_data_res_4__4__0_), .A2(
        npu_inst_pe_1_3_4_n1), .B1(npu_inst_pe_1_3_4_N73), .B2(
        npu_inst_pe_1_3_4_n76), .C1(npu_inst_pe_1_3_4_N65), .C2(
        npu_inst_pe_1_3_4_n77), .ZN(npu_inst_pe_1_3_4_n84) );
  INV_X1 npu_inst_pe_1_3_4_U50 ( .A(npu_inst_pe_1_3_4_n84), .ZN(
        npu_inst_pe_1_3_4_n100) );
  AOI222_X1 npu_inst_pe_1_3_4_U49 ( .A1(npu_inst_int_data_res_4__4__7_), .A2(
        npu_inst_pe_1_3_4_n1), .B1(npu_inst_pe_1_3_4_N80), .B2(
        npu_inst_pe_1_3_4_n76), .C1(npu_inst_pe_1_3_4_N72), .C2(
        npu_inst_pe_1_3_4_n77), .ZN(npu_inst_pe_1_3_4_n75) );
  INV_X1 npu_inst_pe_1_3_4_U48 ( .A(npu_inst_pe_1_3_4_n75), .ZN(
        npu_inst_pe_1_3_4_n32) );
  AOI222_X1 npu_inst_pe_1_3_4_U47 ( .A1(npu_inst_int_data_res_4__4__1_), .A2(
        npu_inst_pe_1_3_4_n1), .B1(npu_inst_pe_1_3_4_N74), .B2(
        npu_inst_pe_1_3_4_n76), .C1(npu_inst_pe_1_3_4_N66), .C2(
        npu_inst_pe_1_3_4_n77), .ZN(npu_inst_pe_1_3_4_n83) );
  INV_X1 npu_inst_pe_1_3_4_U46 ( .A(npu_inst_pe_1_3_4_n83), .ZN(
        npu_inst_pe_1_3_4_n99) );
  AOI222_X1 npu_inst_pe_1_3_4_U45 ( .A1(npu_inst_int_data_res_4__4__2_), .A2(
        npu_inst_pe_1_3_4_n1), .B1(npu_inst_pe_1_3_4_N75), .B2(
        npu_inst_pe_1_3_4_n76), .C1(npu_inst_pe_1_3_4_N67), .C2(
        npu_inst_pe_1_3_4_n77), .ZN(npu_inst_pe_1_3_4_n82) );
  INV_X1 npu_inst_pe_1_3_4_U44 ( .A(npu_inst_pe_1_3_4_n82), .ZN(
        npu_inst_pe_1_3_4_n98) );
  AOI222_X1 npu_inst_pe_1_3_4_U43 ( .A1(npu_inst_int_data_res_4__4__3_), .A2(
        npu_inst_pe_1_3_4_n1), .B1(npu_inst_pe_1_3_4_N76), .B2(
        npu_inst_pe_1_3_4_n76), .C1(npu_inst_pe_1_3_4_N68), .C2(
        npu_inst_pe_1_3_4_n77), .ZN(npu_inst_pe_1_3_4_n81) );
  INV_X1 npu_inst_pe_1_3_4_U42 ( .A(npu_inst_pe_1_3_4_n81), .ZN(
        npu_inst_pe_1_3_4_n36) );
  AOI222_X1 npu_inst_pe_1_3_4_U41 ( .A1(npu_inst_int_data_res_4__4__4_), .A2(
        npu_inst_pe_1_3_4_n1), .B1(npu_inst_pe_1_3_4_N77), .B2(
        npu_inst_pe_1_3_4_n76), .C1(npu_inst_pe_1_3_4_N69), .C2(
        npu_inst_pe_1_3_4_n77), .ZN(npu_inst_pe_1_3_4_n80) );
  INV_X1 npu_inst_pe_1_3_4_U40 ( .A(npu_inst_pe_1_3_4_n80), .ZN(
        npu_inst_pe_1_3_4_n35) );
  AOI222_X1 npu_inst_pe_1_3_4_U39 ( .A1(npu_inst_int_data_res_4__4__5_), .A2(
        npu_inst_pe_1_3_4_n1), .B1(npu_inst_pe_1_3_4_N78), .B2(
        npu_inst_pe_1_3_4_n76), .C1(npu_inst_pe_1_3_4_N70), .C2(
        npu_inst_pe_1_3_4_n77), .ZN(npu_inst_pe_1_3_4_n79) );
  INV_X1 npu_inst_pe_1_3_4_U38 ( .A(npu_inst_pe_1_3_4_n79), .ZN(
        npu_inst_pe_1_3_4_n34) );
  AOI222_X1 npu_inst_pe_1_3_4_U37 ( .A1(npu_inst_int_data_res_4__4__6_), .A2(
        npu_inst_pe_1_3_4_n1), .B1(npu_inst_pe_1_3_4_N79), .B2(
        npu_inst_pe_1_3_4_n76), .C1(npu_inst_pe_1_3_4_N71), .C2(
        npu_inst_pe_1_3_4_n77), .ZN(npu_inst_pe_1_3_4_n78) );
  INV_X1 npu_inst_pe_1_3_4_U36 ( .A(npu_inst_pe_1_3_4_n78), .ZN(
        npu_inst_pe_1_3_4_n33) );
  INV_X1 npu_inst_pe_1_3_4_U35 ( .A(npu_inst_pe_1_3_4_int_data_1_), .ZN(
        npu_inst_pe_1_3_4_n13) );
  AND2_X1 npu_inst_pe_1_3_4_U34 ( .A1(npu_inst_int_data_x_3__4__1_), .A2(
        npu_inst_pe_1_3_4_int_q_weight_1_), .ZN(npu_inst_pe_1_3_4_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_3_4_U33 ( .A1(npu_inst_int_data_x_3__4__0_), .A2(
        npu_inst_pe_1_3_4_int_q_weight_1_), .ZN(npu_inst_pe_1_3_4_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_3_4_U32 ( .A1(npu_inst_n57), .A2(
        npu_inst_int_data_y_4__4__1_), .B1(npu_inst_pe_1_3_4_n3), .B2(
        npu_inst_int_data_x_3__5__1_), .ZN(npu_inst_pe_1_3_4_n63) );
  AOI22_X1 npu_inst_pe_1_3_4_U31 ( .A1(npu_inst_n57), .A2(
        npu_inst_int_data_y_4__4__0_), .B1(npu_inst_pe_1_3_4_n3), .B2(
        npu_inst_int_data_x_3__5__0_), .ZN(npu_inst_pe_1_3_4_n61) );
  INV_X1 npu_inst_pe_1_3_4_U30 ( .A(npu_inst_pe_1_3_4_int_data_0_), .ZN(
        npu_inst_pe_1_3_4_n12) );
  INV_X1 npu_inst_pe_1_3_4_U29 ( .A(npu_inst_n69), .ZN(npu_inst_pe_1_3_4_n5)
         );
  OR3_X1 npu_inst_pe_1_3_4_U28 ( .A1(npu_inst_n77), .A2(npu_inst_pe_1_3_4_n7), 
        .A3(npu_inst_pe_1_3_4_n5), .ZN(npu_inst_pe_1_3_4_n56) );
  OR3_X1 npu_inst_pe_1_3_4_U27 ( .A1(npu_inst_pe_1_3_4_n5), .A2(
        npu_inst_pe_1_3_4_n7), .A3(npu_inst_pe_1_3_4_n6), .ZN(
        npu_inst_pe_1_3_4_n48) );
  INV_X1 npu_inst_pe_1_3_4_U26 ( .A(npu_inst_pe_1_3_4_n5), .ZN(
        npu_inst_pe_1_3_4_n4) );
  INV_X1 npu_inst_pe_1_3_4_U25 ( .A(npu_inst_n124), .ZN(npu_inst_pe_1_3_4_n11)
         );
  OR3_X1 npu_inst_pe_1_3_4_U24 ( .A1(npu_inst_pe_1_3_4_n4), .A2(
        npu_inst_pe_1_3_4_n7), .A3(npu_inst_pe_1_3_4_n6), .ZN(
        npu_inst_pe_1_3_4_n52) );
  OR3_X1 npu_inst_pe_1_3_4_U23 ( .A1(npu_inst_n77), .A2(npu_inst_pe_1_3_4_n7), 
        .A3(npu_inst_pe_1_3_4_n4), .ZN(npu_inst_pe_1_3_4_n60) );
  NOR2_X1 npu_inst_pe_1_3_4_U22 ( .A1(npu_inst_pe_1_3_4_n60), .A2(
        npu_inst_pe_1_3_4_n3), .ZN(npu_inst_pe_1_3_4_n58) );
  NOR2_X1 npu_inst_pe_1_3_4_U21 ( .A1(npu_inst_pe_1_3_4_n56), .A2(
        npu_inst_pe_1_3_4_n3), .ZN(npu_inst_pe_1_3_4_n54) );
  NOR2_X1 npu_inst_pe_1_3_4_U20 ( .A1(npu_inst_pe_1_3_4_n52), .A2(
        npu_inst_pe_1_3_4_n3), .ZN(npu_inst_pe_1_3_4_n50) );
  NOR2_X1 npu_inst_pe_1_3_4_U19 ( .A1(npu_inst_pe_1_3_4_n48), .A2(
        npu_inst_pe_1_3_4_n3), .ZN(npu_inst_pe_1_3_4_n46) );
  NOR2_X1 npu_inst_pe_1_3_4_U18 ( .A1(npu_inst_pe_1_3_4_n40), .A2(
        npu_inst_pe_1_3_4_n3), .ZN(npu_inst_pe_1_3_4_n38) );
  NOR2_X1 npu_inst_pe_1_3_4_U17 ( .A1(npu_inst_pe_1_3_4_n44), .A2(
        npu_inst_pe_1_3_4_n3), .ZN(npu_inst_pe_1_3_4_n42) );
  BUF_X1 npu_inst_pe_1_3_4_U16 ( .A(npu_inst_n100), .Z(npu_inst_pe_1_3_4_n7)
         );
  BUF_X1 npu_inst_pe_1_3_4_U15 ( .A(npu_inst_pe_1_3_4_n11), .Z(
        npu_inst_pe_1_3_4_n10) );
  BUF_X1 npu_inst_pe_1_3_4_U14 ( .A(npu_inst_pe_1_3_4_n11), .Z(
        npu_inst_pe_1_3_4_n9) );
  BUF_X1 npu_inst_pe_1_3_4_U13 ( .A(npu_inst_pe_1_3_4_n11), .Z(
        npu_inst_pe_1_3_4_n8) );
  INV_X1 npu_inst_pe_1_3_4_U12 ( .A(npu_inst_pe_1_3_4_n38), .ZN(
        npu_inst_pe_1_3_4_n117) );
  INV_X1 npu_inst_pe_1_3_4_U11 ( .A(npu_inst_pe_1_3_4_n58), .ZN(
        npu_inst_pe_1_3_4_n113) );
  INV_X1 npu_inst_pe_1_3_4_U10 ( .A(npu_inst_pe_1_3_4_n54), .ZN(
        npu_inst_pe_1_3_4_n114) );
  INV_X1 npu_inst_pe_1_3_4_U9 ( .A(npu_inst_pe_1_3_4_n50), .ZN(
        npu_inst_pe_1_3_4_n115) );
  INV_X1 npu_inst_pe_1_3_4_U8 ( .A(npu_inst_pe_1_3_4_n46), .ZN(
        npu_inst_pe_1_3_4_n116) );
  INV_X1 npu_inst_pe_1_3_4_U7 ( .A(npu_inst_pe_1_3_4_n42), .ZN(
        npu_inst_pe_1_3_4_n118) );
  BUF_X1 npu_inst_pe_1_3_4_U6 ( .A(npu_inst_n24), .Z(npu_inst_pe_1_3_4_n2) );
  BUF_X1 npu_inst_pe_1_3_4_U5 ( .A(npu_inst_n24), .Z(npu_inst_pe_1_3_4_n1) );
  NOR2_X1 npu_inst_pe_1_3_4_U4 ( .A1(npu_inst_pe_1_3_4_int_q_weight_0_), .A2(
        npu_inst_pe_1_3_4_n1), .ZN(npu_inst_pe_1_3_4_n76) );
  NOR2_X1 npu_inst_pe_1_3_4_U3 ( .A1(npu_inst_pe_1_3_4_n27), .A2(
        npu_inst_pe_1_3_4_n1), .ZN(npu_inst_pe_1_3_4_n77) );
  FA_X1 npu_inst_pe_1_3_4_sub_77_U2_1 ( .A(npu_inst_pe_1_3_4_int_q_acc_1_), 
        .B(npu_inst_pe_1_3_4_n13), .CI(npu_inst_pe_1_3_4_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_3_4_sub_77_carry_2_), .S(npu_inst_pe_1_3_4_N66) );
  FA_X1 npu_inst_pe_1_3_4_add_79_U1_1 ( .A(npu_inst_pe_1_3_4_int_q_acc_1_), 
        .B(npu_inst_pe_1_3_4_int_data_1_), .CI(
        npu_inst_pe_1_3_4_add_79_carry_1_), .CO(
        npu_inst_pe_1_3_4_add_79_carry_2_), .S(npu_inst_pe_1_3_4_N74) );
  NAND3_X1 npu_inst_pe_1_3_4_U109 ( .A1(npu_inst_pe_1_3_4_n5), .A2(
        npu_inst_pe_1_3_4_n6), .A3(npu_inst_pe_1_3_4_n7), .ZN(
        npu_inst_pe_1_3_4_n44) );
  NAND3_X1 npu_inst_pe_1_3_4_U108 ( .A1(npu_inst_pe_1_3_4_n4), .A2(
        npu_inst_pe_1_3_4_n6), .A3(npu_inst_pe_1_3_4_n7), .ZN(
        npu_inst_pe_1_3_4_n40) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_3_4_n33), .CK(
        npu_inst_pe_1_3_4_net3649), .RN(npu_inst_pe_1_3_4_n8), .Q(
        npu_inst_pe_1_3_4_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_3_4_n34), .CK(
        npu_inst_pe_1_3_4_net3649), .RN(npu_inst_pe_1_3_4_n8), .Q(
        npu_inst_pe_1_3_4_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_3_4_n35), .CK(
        npu_inst_pe_1_3_4_net3649), .RN(npu_inst_pe_1_3_4_n8), .Q(
        npu_inst_pe_1_3_4_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_3_4_n36), .CK(
        npu_inst_pe_1_3_4_net3649), .RN(npu_inst_pe_1_3_4_n8), .Q(
        npu_inst_pe_1_3_4_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_3_4_n98), .CK(
        npu_inst_pe_1_3_4_net3649), .RN(npu_inst_pe_1_3_4_n8), .Q(
        npu_inst_pe_1_3_4_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_3_4_n99), .CK(
        npu_inst_pe_1_3_4_net3649), .RN(npu_inst_pe_1_3_4_n8), .Q(
        npu_inst_pe_1_3_4_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_3_4_n32), .CK(
        npu_inst_pe_1_3_4_net3649), .RN(npu_inst_pe_1_3_4_n8), .Q(
        npu_inst_pe_1_3_4_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_3_4_n100), 
        .CK(npu_inst_pe_1_3_4_net3649), .RN(npu_inst_pe_1_3_4_n8), .Q(
        npu_inst_pe_1_3_4_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_weight_reg_0_ ( .D(npu_inst_n110), .CK(
        npu_inst_pe_1_3_4_net3655), .RN(npu_inst_pe_1_3_4_n8), .Q(
        npu_inst_pe_1_3_4_int_q_weight_0_), .QN(npu_inst_pe_1_3_4_n27) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_weight_reg_1_ ( .D(npu_inst_n116), .CK(
        npu_inst_pe_1_3_4_net3655), .RN(npu_inst_pe_1_3_4_n8), .Q(
        npu_inst_pe_1_3_4_int_q_weight_1_), .QN(npu_inst_pe_1_3_4_n26) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_3_4_n112), 
        .CK(npu_inst_pe_1_3_4_net3655), .RN(npu_inst_pe_1_3_4_n8), .Q(
        npu_inst_pe_1_3_4_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_3_4_n106), 
        .CK(npu_inst_pe_1_3_4_net3655), .RN(npu_inst_pe_1_3_4_n8), .Q(
        npu_inst_pe_1_3_4_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_3_4_n111), 
        .CK(npu_inst_pe_1_3_4_net3655), .RN(npu_inst_pe_1_3_4_n9), .Q(
        npu_inst_pe_1_3_4_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_3_4_n105), 
        .CK(npu_inst_pe_1_3_4_net3655), .RN(npu_inst_pe_1_3_4_n9), .Q(
        npu_inst_pe_1_3_4_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_3_4_n110), 
        .CK(npu_inst_pe_1_3_4_net3655), .RN(npu_inst_pe_1_3_4_n9), .Q(
        npu_inst_pe_1_3_4_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_3_4_n104), 
        .CK(npu_inst_pe_1_3_4_net3655), .RN(npu_inst_pe_1_3_4_n9), .Q(
        npu_inst_pe_1_3_4_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_3_4_n109), 
        .CK(npu_inst_pe_1_3_4_net3655), .RN(npu_inst_pe_1_3_4_n9), .Q(
        npu_inst_pe_1_3_4_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_3_4_n103), 
        .CK(npu_inst_pe_1_3_4_net3655), .RN(npu_inst_pe_1_3_4_n9), .Q(
        npu_inst_pe_1_3_4_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_3_4_n108), 
        .CK(npu_inst_pe_1_3_4_net3655), .RN(npu_inst_pe_1_3_4_n9), .Q(
        npu_inst_pe_1_3_4_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_3_4_n102), 
        .CK(npu_inst_pe_1_3_4_net3655), .RN(npu_inst_pe_1_3_4_n9), .Q(
        npu_inst_pe_1_3_4_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_3_4_n107), 
        .CK(npu_inst_pe_1_3_4_net3655), .RN(npu_inst_pe_1_3_4_n9), .Q(
        npu_inst_pe_1_3_4_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_3_4_n101), 
        .CK(npu_inst_pe_1_3_4_net3655), .RN(npu_inst_pe_1_3_4_n9), .Q(
        npu_inst_pe_1_3_4_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_3_4_n86), 
        .CK(npu_inst_pe_1_3_4_net3655), .RN(npu_inst_pe_1_3_4_n9), .Q(
        npu_inst_pe_1_3_4_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_3_4_n87), 
        .CK(npu_inst_pe_1_3_4_net3655), .RN(npu_inst_pe_1_3_4_n9), .Q(
        npu_inst_pe_1_3_4_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_3_4_n88), 
        .CK(npu_inst_pe_1_3_4_net3655), .RN(npu_inst_pe_1_3_4_n10), .Q(
        npu_inst_pe_1_3_4_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_3_4_n89), 
        .CK(npu_inst_pe_1_3_4_net3655), .RN(npu_inst_pe_1_3_4_n10), .Q(
        npu_inst_pe_1_3_4_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_3_4_n90), 
        .CK(npu_inst_pe_1_3_4_net3655), .RN(npu_inst_pe_1_3_4_n10), .Q(
        npu_inst_pe_1_3_4_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_3_4_n91), 
        .CK(npu_inst_pe_1_3_4_net3655), .RN(npu_inst_pe_1_3_4_n10), .Q(
        npu_inst_pe_1_3_4_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_3_4_n92), 
        .CK(npu_inst_pe_1_3_4_net3655), .RN(npu_inst_pe_1_3_4_n10), .Q(
        npu_inst_pe_1_3_4_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_3_4_n93), 
        .CK(npu_inst_pe_1_3_4_net3655), .RN(npu_inst_pe_1_3_4_n10), .Q(
        npu_inst_pe_1_3_4_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_3_4_n94), 
        .CK(npu_inst_pe_1_3_4_net3655), .RN(npu_inst_pe_1_3_4_n10), .Q(
        npu_inst_pe_1_3_4_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_3_4_n95), 
        .CK(npu_inst_pe_1_3_4_net3655), .RN(npu_inst_pe_1_3_4_n10), .Q(
        npu_inst_pe_1_3_4_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_3_4_n96), 
        .CK(npu_inst_pe_1_3_4_net3655), .RN(npu_inst_pe_1_3_4_n10), .Q(
        npu_inst_pe_1_3_4_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_3_4_n97), 
        .CK(npu_inst_pe_1_3_4_net3655), .RN(npu_inst_pe_1_3_4_n10), .Q(
        npu_inst_pe_1_3_4_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_3_4_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_3_4_N84), .SE(1'b0), .GCK(npu_inst_pe_1_3_4_net3649) );
  CLKGATETST_X1 npu_inst_pe_1_3_4_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n64), .SE(1'b0), .GCK(npu_inst_pe_1_3_4_net3655) );
  MUX2_X1 npu_inst_pe_1_3_5_U162 ( .A(npu_inst_pe_1_3_5_n32), .B(
        npu_inst_pe_1_3_5_n29), .S(npu_inst_pe_1_3_5_n8), .Z(
        npu_inst_pe_1_3_5_N93) );
  MUX2_X1 npu_inst_pe_1_3_5_U161 ( .A(npu_inst_pe_1_3_5_n31), .B(
        npu_inst_pe_1_3_5_n30), .S(npu_inst_pe_1_3_5_n6), .Z(
        npu_inst_pe_1_3_5_n32) );
  MUX2_X1 npu_inst_pe_1_3_5_U160 ( .A(npu_inst_pe_1_3_5_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_3_5_int_q_reg_v_1__0_), .S(npu_inst_pe_1_3_5_n4), .Z(
        npu_inst_pe_1_3_5_n31) );
  MUX2_X1 npu_inst_pe_1_3_5_U159 ( .A(npu_inst_pe_1_3_5_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_3_5_int_q_reg_v_3__0_), .S(npu_inst_pe_1_3_5_n4), .Z(
        npu_inst_pe_1_3_5_n30) );
  MUX2_X1 npu_inst_pe_1_3_5_U158 ( .A(npu_inst_pe_1_3_5_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_3_5_int_q_reg_v_5__0_), .S(npu_inst_pe_1_3_5_n4), .Z(
        npu_inst_pe_1_3_5_n29) );
  MUX2_X1 npu_inst_pe_1_3_5_U157 ( .A(npu_inst_pe_1_3_5_n28), .B(
        npu_inst_pe_1_3_5_n23), .S(npu_inst_pe_1_3_5_n8), .Z(
        npu_inst_pe_1_3_5_N94) );
  MUX2_X1 npu_inst_pe_1_3_5_U156 ( .A(npu_inst_pe_1_3_5_n25), .B(
        npu_inst_pe_1_3_5_n24), .S(npu_inst_pe_1_3_5_n6), .Z(
        npu_inst_pe_1_3_5_n28) );
  MUX2_X1 npu_inst_pe_1_3_5_U155 ( .A(npu_inst_pe_1_3_5_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_3_5_int_q_reg_v_1__1_), .S(npu_inst_pe_1_3_5_n4), .Z(
        npu_inst_pe_1_3_5_n25) );
  MUX2_X1 npu_inst_pe_1_3_5_U154 ( .A(npu_inst_pe_1_3_5_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_3_5_int_q_reg_v_3__1_), .S(npu_inst_pe_1_3_5_n4), .Z(
        npu_inst_pe_1_3_5_n24) );
  MUX2_X1 npu_inst_pe_1_3_5_U153 ( .A(npu_inst_pe_1_3_5_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_3_5_int_q_reg_v_5__1_), .S(npu_inst_pe_1_3_5_n4), .Z(
        npu_inst_pe_1_3_5_n23) );
  MUX2_X1 npu_inst_pe_1_3_5_U152 ( .A(npu_inst_pe_1_3_5_n22), .B(
        npu_inst_pe_1_3_5_n19), .S(npu_inst_pe_1_3_5_n8), .Z(
        npu_inst_int_data_x_3__5__1_) );
  MUX2_X1 npu_inst_pe_1_3_5_U151 ( .A(npu_inst_pe_1_3_5_n21), .B(
        npu_inst_pe_1_3_5_n20), .S(npu_inst_pe_1_3_5_n6), .Z(
        npu_inst_pe_1_3_5_n22) );
  MUX2_X1 npu_inst_pe_1_3_5_U150 ( .A(npu_inst_pe_1_3_5_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_3_5_int_q_reg_h_1__1_), .S(npu_inst_pe_1_3_5_n4), .Z(
        npu_inst_pe_1_3_5_n21) );
  MUX2_X1 npu_inst_pe_1_3_5_U149 ( .A(npu_inst_pe_1_3_5_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_3_5_int_q_reg_h_3__1_), .S(npu_inst_pe_1_3_5_n4), .Z(
        npu_inst_pe_1_3_5_n20) );
  MUX2_X1 npu_inst_pe_1_3_5_U148 ( .A(npu_inst_pe_1_3_5_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_3_5_int_q_reg_h_5__1_), .S(npu_inst_pe_1_3_5_n4), .Z(
        npu_inst_pe_1_3_5_n19) );
  MUX2_X1 npu_inst_pe_1_3_5_U147 ( .A(npu_inst_pe_1_3_5_n18), .B(
        npu_inst_pe_1_3_5_n15), .S(npu_inst_pe_1_3_5_n8), .Z(
        npu_inst_int_data_x_3__5__0_) );
  MUX2_X1 npu_inst_pe_1_3_5_U146 ( .A(npu_inst_pe_1_3_5_n17), .B(
        npu_inst_pe_1_3_5_n16), .S(npu_inst_pe_1_3_5_n6), .Z(
        npu_inst_pe_1_3_5_n18) );
  MUX2_X1 npu_inst_pe_1_3_5_U145 ( .A(npu_inst_pe_1_3_5_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_3_5_int_q_reg_h_1__0_), .S(npu_inst_pe_1_3_5_n4), .Z(
        npu_inst_pe_1_3_5_n17) );
  MUX2_X1 npu_inst_pe_1_3_5_U144 ( .A(npu_inst_pe_1_3_5_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_3_5_int_q_reg_h_3__0_), .S(npu_inst_pe_1_3_5_n4), .Z(
        npu_inst_pe_1_3_5_n16) );
  MUX2_X1 npu_inst_pe_1_3_5_U143 ( .A(npu_inst_pe_1_3_5_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_3_5_int_q_reg_h_5__0_), .S(npu_inst_pe_1_3_5_n4), .Z(
        npu_inst_pe_1_3_5_n15) );
  XOR2_X1 npu_inst_pe_1_3_5_U142 ( .A(npu_inst_pe_1_3_5_int_data_0_), .B(
        npu_inst_pe_1_3_5_int_q_acc_0_), .Z(npu_inst_pe_1_3_5_N73) );
  AND2_X1 npu_inst_pe_1_3_5_U141 ( .A1(npu_inst_pe_1_3_5_int_q_acc_0_), .A2(
        npu_inst_pe_1_3_5_int_data_0_), .ZN(npu_inst_pe_1_3_5_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_3_5_U140 ( .A(npu_inst_pe_1_3_5_int_q_acc_0_), .B(
        npu_inst_pe_1_3_5_n13), .ZN(npu_inst_pe_1_3_5_N65) );
  OR2_X1 npu_inst_pe_1_3_5_U139 ( .A1(npu_inst_pe_1_3_5_n13), .A2(
        npu_inst_pe_1_3_5_int_q_acc_0_), .ZN(npu_inst_pe_1_3_5_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_3_5_U138 ( .A(npu_inst_pe_1_3_5_int_q_acc_2_), .B(
        npu_inst_pe_1_3_5_add_79_carry_2_), .Z(npu_inst_pe_1_3_5_N75) );
  AND2_X1 npu_inst_pe_1_3_5_U137 ( .A1(npu_inst_pe_1_3_5_add_79_carry_2_), 
        .A2(npu_inst_pe_1_3_5_int_q_acc_2_), .ZN(
        npu_inst_pe_1_3_5_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_3_5_U136 ( .A(npu_inst_pe_1_3_5_int_q_acc_3_), .B(
        npu_inst_pe_1_3_5_add_79_carry_3_), .Z(npu_inst_pe_1_3_5_N76) );
  AND2_X1 npu_inst_pe_1_3_5_U135 ( .A1(npu_inst_pe_1_3_5_add_79_carry_3_), 
        .A2(npu_inst_pe_1_3_5_int_q_acc_3_), .ZN(
        npu_inst_pe_1_3_5_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_3_5_U134 ( .A(npu_inst_pe_1_3_5_int_q_acc_4_), .B(
        npu_inst_pe_1_3_5_add_79_carry_4_), .Z(npu_inst_pe_1_3_5_N77) );
  AND2_X1 npu_inst_pe_1_3_5_U133 ( .A1(npu_inst_pe_1_3_5_add_79_carry_4_), 
        .A2(npu_inst_pe_1_3_5_int_q_acc_4_), .ZN(
        npu_inst_pe_1_3_5_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_3_5_U132 ( .A(npu_inst_pe_1_3_5_int_q_acc_5_), .B(
        npu_inst_pe_1_3_5_add_79_carry_5_), .Z(npu_inst_pe_1_3_5_N78) );
  AND2_X1 npu_inst_pe_1_3_5_U131 ( .A1(npu_inst_pe_1_3_5_add_79_carry_5_), 
        .A2(npu_inst_pe_1_3_5_int_q_acc_5_), .ZN(
        npu_inst_pe_1_3_5_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_3_5_U130 ( .A(npu_inst_pe_1_3_5_int_q_acc_6_), .B(
        npu_inst_pe_1_3_5_add_79_carry_6_), .Z(npu_inst_pe_1_3_5_N79) );
  AND2_X1 npu_inst_pe_1_3_5_U129 ( .A1(npu_inst_pe_1_3_5_add_79_carry_6_), 
        .A2(npu_inst_pe_1_3_5_int_q_acc_6_), .ZN(
        npu_inst_pe_1_3_5_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_3_5_U128 ( .A(npu_inst_pe_1_3_5_int_q_acc_7_), .B(
        npu_inst_pe_1_3_5_add_79_carry_7_), .Z(npu_inst_pe_1_3_5_N80) );
  XNOR2_X1 npu_inst_pe_1_3_5_U127 ( .A(npu_inst_pe_1_3_5_sub_77_carry_2_), .B(
        npu_inst_pe_1_3_5_int_q_acc_2_), .ZN(npu_inst_pe_1_3_5_N67) );
  OR2_X1 npu_inst_pe_1_3_5_U126 ( .A1(npu_inst_pe_1_3_5_int_q_acc_2_), .A2(
        npu_inst_pe_1_3_5_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_3_5_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_3_5_U125 ( .A(npu_inst_pe_1_3_5_sub_77_carry_3_), .B(
        npu_inst_pe_1_3_5_int_q_acc_3_), .ZN(npu_inst_pe_1_3_5_N68) );
  OR2_X1 npu_inst_pe_1_3_5_U124 ( .A1(npu_inst_pe_1_3_5_int_q_acc_3_), .A2(
        npu_inst_pe_1_3_5_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_3_5_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_3_5_U123 ( .A(npu_inst_pe_1_3_5_sub_77_carry_4_), .B(
        npu_inst_pe_1_3_5_int_q_acc_4_), .ZN(npu_inst_pe_1_3_5_N69) );
  OR2_X1 npu_inst_pe_1_3_5_U122 ( .A1(npu_inst_pe_1_3_5_int_q_acc_4_), .A2(
        npu_inst_pe_1_3_5_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_3_5_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_3_5_U121 ( .A(npu_inst_pe_1_3_5_sub_77_carry_5_), .B(
        npu_inst_pe_1_3_5_int_q_acc_5_), .ZN(npu_inst_pe_1_3_5_N70) );
  OR2_X1 npu_inst_pe_1_3_5_U120 ( .A1(npu_inst_pe_1_3_5_int_q_acc_5_), .A2(
        npu_inst_pe_1_3_5_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_3_5_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_3_5_U119 ( .A(npu_inst_pe_1_3_5_sub_77_carry_6_), .B(
        npu_inst_pe_1_3_5_int_q_acc_6_), .ZN(npu_inst_pe_1_3_5_N71) );
  OR2_X1 npu_inst_pe_1_3_5_U118 ( .A1(npu_inst_pe_1_3_5_int_q_acc_6_), .A2(
        npu_inst_pe_1_3_5_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_3_5_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_3_5_U117 ( .A(npu_inst_pe_1_3_5_int_q_acc_7_), .B(
        npu_inst_pe_1_3_5_sub_77_carry_7_), .ZN(npu_inst_pe_1_3_5_N72) );
  INV_X1 npu_inst_pe_1_3_5_U116 ( .A(npu_inst_n77), .ZN(npu_inst_pe_1_3_5_n7)
         );
  INV_X1 npu_inst_pe_1_3_5_U115 ( .A(npu_inst_pe_1_3_5_n7), .ZN(
        npu_inst_pe_1_3_5_n6) );
  INV_X1 npu_inst_pe_1_3_5_U114 ( .A(npu_inst_n56), .ZN(npu_inst_pe_1_3_5_n3)
         );
  AOI22_X1 npu_inst_pe_1_3_5_U113 ( .A1(npu_inst_int_data_y_4__5__0_), .A2(
        npu_inst_pe_1_3_5_n58), .B1(npu_inst_pe_1_3_5_n114), .B2(
        npu_inst_pe_1_3_5_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_3_5_n57) );
  INV_X1 npu_inst_pe_1_3_5_U112 ( .A(npu_inst_pe_1_3_5_n57), .ZN(
        npu_inst_pe_1_3_5_n108) );
  AOI22_X1 npu_inst_pe_1_3_5_U111 ( .A1(npu_inst_int_data_y_4__5__0_), .A2(
        npu_inst_pe_1_3_5_n54), .B1(npu_inst_pe_1_3_5_n115), .B2(
        npu_inst_pe_1_3_5_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_3_5_n53) );
  INV_X1 npu_inst_pe_1_3_5_U110 ( .A(npu_inst_pe_1_3_5_n53), .ZN(
        npu_inst_pe_1_3_5_n109) );
  AOI22_X1 npu_inst_pe_1_3_5_U107 ( .A1(npu_inst_int_data_y_4__5__0_), .A2(
        npu_inst_pe_1_3_5_n50), .B1(npu_inst_pe_1_3_5_n116), .B2(
        npu_inst_pe_1_3_5_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_3_5_n49) );
  INV_X1 npu_inst_pe_1_3_5_U106 ( .A(npu_inst_pe_1_3_5_n49), .ZN(
        npu_inst_pe_1_3_5_n110) );
  AOI22_X1 npu_inst_pe_1_3_5_U105 ( .A1(npu_inst_int_data_y_4__5__0_), .A2(
        npu_inst_pe_1_3_5_n46), .B1(npu_inst_pe_1_3_5_n117), .B2(
        npu_inst_pe_1_3_5_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_3_5_n45) );
  INV_X1 npu_inst_pe_1_3_5_U104 ( .A(npu_inst_pe_1_3_5_n45), .ZN(
        npu_inst_pe_1_3_5_n111) );
  AOI22_X1 npu_inst_pe_1_3_5_U103 ( .A1(npu_inst_int_data_y_4__5__0_), .A2(
        npu_inst_pe_1_3_5_n42), .B1(npu_inst_pe_1_3_5_n119), .B2(
        npu_inst_pe_1_3_5_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_3_5_n41) );
  INV_X1 npu_inst_pe_1_3_5_U102 ( .A(npu_inst_pe_1_3_5_n41), .ZN(
        npu_inst_pe_1_3_5_n112) );
  AOI22_X1 npu_inst_pe_1_3_5_U101 ( .A1(npu_inst_int_data_y_4__5__1_), .A2(
        npu_inst_pe_1_3_5_n58), .B1(npu_inst_pe_1_3_5_n114), .B2(
        npu_inst_pe_1_3_5_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_3_5_n59) );
  INV_X1 npu_inst_pe_1_3_5_U100 ( .A(npu_inst_pe_1_3_5_n59), .ZN(
        npu_inst_pe_1_3_5_n102) );
  AOI22_X1 npu_inst_pe_1_3_5_U99 ( .A1(npu_inst_int_data_y_4__5__1_), .A2(
        npu_inst_pe_1_3_5_n54), .B1(npu_inst_pe_1_3_5_n115), .B2(
        npu_inst_pe_1_3_5_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_3_5_n55) );
  INV_X1 npu_inst_pe_1_3_5_U98 ( .A(npu_inst_pe_1_3_5_n55), .ZN(
        npu_inst_pe_1_3_5_n103) );
  AOI22_X1 npu_inst_pe_1_3_5_U97 ( .A1(npu_inst_int_data_y_4__5__1_), .A2(
        npu_inst_pe_1_3_5_n50), .B1(npu_inst_pe_1_3_5_n116), .B2(
        npu_inst_pe_1_3_5_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_3_5_n51) );
  INV_X1 npu_inst_pe_1_3_5_U96 ( .A(npu_inst_pe_1_3_5_n51), .ZN(
        npu_inst_pe_1_3_5_n104) );
  AOI22_X1 npu_inst_pe_1_3_5_U95 ( .A1(npu_inst_int_data_y_4__5__1_), .A2(
        npu_inst_pe_1_3_5_n46), .B1(npu_inst_pe_1_3_5_n117), .B2(
        npu_inst_pe_1_3_5_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_3_5_n47) );
  INV_X1 npu_inst_pe_1_3_5_U94 ( .A(npu_inst_pe_1_3_5_n47), .ZN(
        npu_inst_pe_1_3_5_n105) );
  AOI22_X1 npu_inst_pe_1_3_5_U93 ( .A1(npu_inst_int_data_y_4__5__1_), .A2(
        npu_inst_pe_1_3_5_n42), .B1(npu_inst_pe_1_3_5_n119), .B2(
        npu_inst_pe_1_3_5_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_3_5_n43) );
  INV_X1 npu_inst_pe_1_3_5_U92 ( .A(npu_inst_pe_1_3_5_n43), .ZN(
        npu_inst_pe_1_3_5_n106) );
  AOI22_X1 npu_inst_pe_1_3_5_U91 ( .A1(npu_inst_pe_1_3_5_n38), .A2(
        npu_inst_int_data_y_4__5__1_), .B1(npu_inst_pe_1_3_5_n118), .B2(
        npu_inst_pe_1_3_5_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_3_5_n39) );
  INV_X1 npu_inst_pe_1_3_5_U90 ( .A(npu_inst_pe_1_3_5_n39), .ZN(
        npu_inst_pe_1_3_5_n107) );
  AOI22_X1 npu_inst_pe_1_3_5_U89 ( .A1(npu_inst_pe_1_3_5_n38), .A2(
        npu_inst_int_data_y_4__5__0_), .B1(npu_inst_pe_1_3_5_n118), .B2(
        npu_inst_pe_1_3_5_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_3_5_n37) );
  INV_X1 npu_inst_pe_1_3_5_U88 ( .A(npu_inst_pe_1_3_5_n37), .ZN(
        npu_inst_pe_1_3_5_n113) );
  NAND2_X1 npu_inst_pe_1_3_5_U87 ( .A1(npu_inst_pe_1_3_5_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_3_5_n60), .ZN(npu_inst_pe_1_3_5_n74) );
  OAI21_X1 npu_inst_pe_1_3_5_U86 ( .B1(npu_inst_pe_1_3_5_n63), .B2(
        npu_inst_pe_1_3_5_n60), .A(npu_inst_pe_1_3_5_n74), .ZN(
        npu_inst_pe_1_3_5_n97) );
  NAND2_X1 npu_inst_pe_1_3_5_U85 ( .A1(npu_inst_pe_1_3_5_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_3_5_n60), .ZN(npu_inst_pe_1_3_5_n73) );
  OAI21_X1 npu_inst_pe_1_3_5_U84 ( .B1(npu_inst_pe_1_3_5_n61), .B2(
        npu_inst_pe_1_3_5_n60), .A(npu_inst_pe_1_3_5_n73), .ZN(
        npu_inst_pe_1_3_5_n96) );
  NAND2_X1 npu_inst_pe_1_3_5_U83 ( .A1(npu_inst_pe_1_3_5_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_3_5_n56), .ZN(npu_inst_pe_1_3_5_n72) );
  OAI21_X1 npu_inst_pe_1_3_5_U82 ( .B1(npu_inst_pe_1_3_5_n63), .B2(
        npu_inst_pe_1_3_5_n56), .A(npu_inst_pe_1_3_5_n72), .ZN(
        npu_inst_pe_1_3_5_n95) );
  NAND2_X1 npu_inst_pe_1_3_5_U81 ( .A1(npu_inst_pe_1_3_5_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_3_5_n56), .ZN(npu_inst_pe_1_3_5_n71) );
  OAI21_X1 npu_inst_pe_1_3_5_U80 ( .B1(npu_inst_pe_1_3_5_n61), .B2(
        npu_inst_pe_1_3_5_n56), .A(npu_inst_pe_1_3_5_n71), .ZN(
        npu_inst_pe_1_3_5_n94) );
  NAND2_X1 npu_inst_pe_1_3_5_U79 ( .A1(npu_inst_pe_1_3_5_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_3_5_n52), .ZN(npu_inst_pe_1_3_5_n70) );
  OAI21_X1 npu_inst_pe_1_3_5_U78 ( .B1(npu_inst_pe_1_3_5_n63), .B2(
        npu_inst_pe_1_3_5_n52), .A(npu_inst_pe_1_3_5_n70), .ZN(
        npu_inst_pe_1_3_5_n93) );
  NAND2_X1 npu_inst_pe_1_3_5_U77 ( .A1(npu_inst_pe_1_3_5_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_3_5_n52), .ZN(npu_inst_pe_1_3_5_n69) );
  OAI21_X1 npu_inst_pe_1_3_5_U76 ( .B1(npu_inst_pe_1_3_5_n61), .B2(
        npu_inst_pe_1_3_5_n52), .A(npu_inst_pe_1_3_5_n69), .ZN(
        npu_inst_pe_1_3_5_n92) );
  NAND2_X1 npu_inst_pe_1_3_5_U75 ( .A1(npu_inst_pe_1_3_5_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_3_5_n48), .ZN(npu_inst_pe_1_3_5_n68) );
  OAI21_X1 npu_inst_pe_1_3_5_U74 ( .B1(npu_inst_pe_1_3_5_n63), .B2(
        npu_inst_pe_1_3_5_n48), .A(npu_inst_pe_1_3_5_n68), .ZN(
        npu_inst_pe_1_3_5_n91) );
  NAND2_X1 npu_inst_pe_1_3_5_U73 ( .A1(npu_inst_pe_1_3_5_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_3_5_n48), .ZN(npu_inst_pe_1_3_5_n67) );
  OAI21_X1 npu_inst_pe_1_3_5_U72 ( .B1(npu_inst_pe_1_3_5_n61), .B2(
        npu_inst_pe_1_3_5_n48), .A(npu_inst_pe_1_3_5_n67), .ZN(
        npu_inst_pe_1_3_5_n90) );
  NAND2_X1 npu_inst_pe_1_3_5_U71 ( .A1(npu_inst_pe_1_3_5_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_3_5_n44), .ZN(npu_inst_pe_1_3_5_n66) );
  OAI21_X1 npu_inst_pe_1_3_5_U70 ( .B1(npu_inst_pe_1_3_5_n63), .B2(
        npu_inst_pe_1_3_5_n44), .A(npu_inst_pe_1_3_5_n66), .ZN(
        npu_inst_pe_1_3_5_n89) );
  NAND2_X1 npu_inst_pe_1_3_5_U69 ( .A1(npu_inst_pe_1_3_5_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_3_5_n44), .ZN(npu_inst_pe_1_3_5_n65) );
  OAI21_X1 npu_inst_pe_1_3_5_U68 ( .B1(npu_inst_pe_1_3_5_n61), .B2(
        npu_inst_pe_1_3_5_n44), .A(npu_inst_pe_1_3_5_n65), .ZN(
        npu_inst_pe_1_3_5_n88) );
  NAND2_X1 npu_inst_pe_1_3_5_U67 ( .A1(npu_inst_pe_1_3_5_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_3_5_n40), .ZN(npu_inst_pe_1_3_5_n64) );
  OAI21_X1 npu_inst_pe_1_3_5_U66 ( .B1(npu_inst_pe_1_3_5_n63), .B2(
        npu_inst_pe_1_3_5_n40), .A(npu_inst_pe_1_3_5_n64), .ZN(
        npu_inst_pe_1_3_5_n87) );
  NAND2_X1 npu_inst_pe_1_3_5_U65 ( .A1(npu_inst_pe_1_3_5_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_3_5_n40), .ZN(npu_inst_pe_1_3_5_n62) );
  OAI21_X1 npu_inst_pe_1_3_5_U64 ( .B1(npu_inst_pe_1_3_5_n61), .B2(
        npu_inst_pe_1_3_5_n40), .A(npu_inst_pe_1_3_5_n62), .ZN(
        npu_inst_pe_1_3_5_n86) );
  AND2_X1 npu_inst_pe_1_3_5_U63 ( .A1(npu_inst_pe_1_3_5_N93), .A2(npu_inst_n56), .ZN(npu_inst_int_data_y_3__5__0_) );
  AND2_X1 npu_inst_pe_1_3_5_U62 ( .A1(npu_inst_n56), .A2(npu_inst_pe_1_3_5_N94), .ZN(npu_inst_int_data_y_3__5__1_) );
  NOR3_X1 npu_inst_pe_1_3_5_U61 ( .A1(npu_inst_pe_1_3_5_n26), .A2(npu_inst_n56), .A3(npu_inst_int_ckg[34]), .ZN(npu_inst_pe_1_3_5_n85) );
  OR2_X1 npu_inst_pe_1_3_5_U60 ( .A1(npu_inst_pe_1_3_5_n85), .A2(
        npu_inst_pe_1_3_5_n2), .ZN(npu_inst_pe_1_3_5_N84) );
  AND2_X1 npu_inst_pe_1_3_5_U59 ( .A1(npu_inst_pe_1_3_5_int_q_acc_0_), .A2(
        npu_inst_pe_1_3_5_n1), .ZN(npu_inst_int_data_res_3__5__0_) );
  AND2_X1 npu_inst_pe_1_3_5_U58 ( .A1(npu_inst_pe_1_3_5_n2), .A2(
        npu_inst_pe_1_3_5_int_q_acc_7_), .ZN(npu_inst_int_data_res_3__5__7_)
         );
  AND2_X1 npu_inst_pe_1_3_5_U57 ( .A1(npu_inst_pe_1_3_5_int_q_acc_1_), .A2(
        npu_inst_pe_1_3_5_n1), .ZN(npu_inst_int_data_res_3__5__1_) );
  AND2_X1 npu_inst_pe_1_3_5_U56 ( .A1(npu_inst_pe_1_3_5_int_q_acc_2_), .A2(
        npu_inst_pe_1_3_5_n1), .ZN(npu_inst_int_data_res_3__5__2_) );
  AND2_X1 npu_inst_pe_1_3_5_U55 ( .A1(npu_inst_pe_1_3_5_int_q_acc_3_), .A2(
        npu_inst_pe_1_3_5_n2), .ZN(npu_inst_int_data_res_3__5__3_) );
  AND2_X1 npu_inst_pe_1_3_5_U54 ( .A1(npu_inst_pe_1_3_5_int_q_acc_4_), .A2(
        npu_inst_pe_1_3_5_n2), .ZN(npu_inst_int_data_res_3__5__4_) );
  AND2_X1 npu_inst_pe_1_3_5_U53 ( .A1(npu_inst_pe_1_3_5_int_q_acc_5_), .A2(
        npu_inst_pe_1_3_5_n2), .ZN(npu_inst_int_data_res_3__5__5_) );
  AND2_X1 npu_inst_pe_1_3_5_U52 ( .A1(npu_inst_pe_1_3_5_int_q_acc_6_), .A2(
        npu_inst_pe_1_3_5_n2), .ZN(npu_inst_int_data_res_3__5__6_) );
  AOI222_X1 npu_inst_pe_1_3_5_U51 ( .A1(npu_inst_int_data_res_4__5__0_), .A2(
        npu_inst_pe_1_3_5_n1), .B1(npu_inst_pe_1_3_5_N73), .B2(
        npu_inst_pe_1_3_5_n76), .C1(npu_inst_pe_1_3_5_N65), .C2(
        npu_inst_pe_1_3_5_n77), .ZN(npu_inst_pe_1_3_5_n84) );
  INV_X1 npu_inst_pe_1_3_5_U50 ( .A(npu_inst_pe_1_3_5_n84), .ZN(
        npu_inst_pe_1_3_5_n101) );
  AOI222_X1 npu_inst_pe_1_3_5_U49 ( .A1(npu_inst_int_data_res_4__5__7_), .A2(
        npu_inst_pe_1_3_5_n1), .B1(npu_inst_pe_1_3_5_N80), .B2(
        npu_inst_pe_1_3_5_n76), .C1(npu_inst_pe_1_3_5_N72), .C2(
        npu_inst_pe_1_3_5_n77), .ZN(npu_inst_pe_1_3_5_n75) );
  INV_X1 npu_inst_pe_1_3_5_U48 ( .A(npu_inst_pe_1_3_5_n75), .ZN(
        npu_inst_pe_1_3_5_n33) );
  AOI222_X1 npu_inst_pe_1_3_5_U47 ( .A1(npu_inst_int_data_res_4__5__1_), .A2(
        npu_inst_pe_1_3_5_n1), .B1(npu_inst_pe_1_3_5_N74), .B2(
        npu_inst_pe_1_3_5_n76), .C1(npu_inst_pe_1_3_5_N66), .C2(
        npu_inst_pe_1_3_5_n77), .ZN(npu_inst_pe_1_3_5_n83) );
  INV_X1 npu_inst_pe_1_3_5_U46 ( .A(npu_inst_pe_1_3_5_n83), .ZN(
        npu_inst_pe_1_3_5_n100) );
  AOI222_X1 npu_inst_pe_1_3_5_U45 ( .A1(npu_inst_int_data_res_4__5__2_), .A2(
        npu_inst_pe_1_3_5_n1), .B1(npu_inst_pe_1_3_5_N75), .B2(
        npu_inst_pe_1_3_5_n76), .C1(npu_inst_pe_1_3_5_N67), .C2(
        npu_inst_pe_1_3_5_n77), .ZN(npu_inst_pe_1_3_5_n82) );
  INV_X1 npu_inst_pe_1_3_5_U44 ( .A(npu_inst_pe_1_3_5_n82), .ZN(
        npu_inst_pe_1_3_5_n99) );
  AOI222_X1 npu_inst_pe_1_3_5_U43 ( .A1(npu_inst_int_data_res_4__5__3_), .A2(
        npu_inst_pe_1_3_5_n1), .B1(npu_inst_pe_1_3_5_N76), .B2(
        npu_inst_pe_1_3_5_n76), .C1(npu_inst_pe_1_3_5_N68), .C2(
        npu_inst_pe_1_3_5_n77), .ZN(npu_inst_pe_1_3_5_n81) );
  INV_X1 npu_inst_pe_1_3_5_U42 ( .A(npu_inst_pe_1_3_5_n81), .ZN(
        npu_inst_pe_1_3_5_n98) );
  AOI222_X1 npu_inst_pe_1_3_5_U41 ( .A1(npu_inst_int_data_res_4__5__4_), .A2(
        npu_inst_pe_1_3_5_n1), .B1(npu_inst_pe_1_3_5_N77), .B2(
        npu_inst_pe_1_3_5_n76), .C1(npu_inst_pe_1_3_5_N69), .C2(
        npu_inst_pe_1_3_5_n77), .ZN(npu_inst_pe_1_3_5_n80) );
  INV_X1 npu_inst_pe_1_3_5_U40 ( .A(npu_inst_pe_1_3_5_n80), .ZN(
        npu_inst_pe_1_3_5_n36) );
  AOI222_X1 npu_inst_pe_1_3_5_U39 ( .A1(npu_inst_int_data_res_4__5__5_), .A2(
        npu_inst_pe_1_3_5_n1), .B1(npu_inst_pe_1_3_5_N78), .B2(
        npu_inst_pe_1_3_5_n76), .C1(npu_inst_pe_1_3_5_N70), .C2(
        npu_inst_pe_1_3_5_n77), .ZN(npu_inst_pe_1_3_5_n79) );
  INV_X1 npu_inst_pe_1_3_5_U38 ( .A(npu_inst_pe_1_3_5_n79), .ZN(
        npu_inst_pe_1_3_5_n35) );
  AOI222_X1 npu_inst_pe_1_3_5_U37 ( .A1(npu_inst_int_data_res_4__5__6_), .A2(
        npu_inst_pe_1_3_5_n1), .B1(npu_inst_pe_1_3_5_N79), .B2(
        npu_inst_pe_1_3_5_n76), .C1(npu_inst_pe_1_3_5_N71), .C2(
        npu_inst_pe_1_3_5_n77), .ZN(npu_inst_pe_1_3_5_n78) );
  INV_X1 npu_inst_pe_1_3_5_U36 ( .A(npu_inst_pe_1_3_5_n78), .ZN(
        npu_inst_pe_1_3_5_n34) );
  INV_X1 npu_inst_pe_1_3_5_U35 ( .A(npu_inst_pe_1_3_5_int_data_1_), .ZN(
        npu_inst_pe_1_3_5_n14) );
  AND2_X1 npu_inst_pe_1_3_5_U34 ( .A1(npu_inst_int_data_x_3__5__1_), .A2(
        npu_inst_pe_1_3_5_int_q_weight_1_), .ZN(npu_inst_pe_1_3_5_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_3_5_U33 ( .A1(npu_inst_int_data_x_3__5__0_), .A2(
        npu_inst_pe_1_3_5_int_q_weight_1_), .ZN(npu_inst_pe_1_3_5_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_3_5_U32 ( .A1(npu_inst_n56), .A2(
        npu_inst_int_data_y_4__5__1_), .B1(npu_inst_pe_1_3_5_n3), .B2(
        npu_inst_int_data_x_3__6__1_), .ZN(npu_inst_pe_1_3_5_n63) );
  AOI22_X1 npu_inst_pe_1_3_5_U31 ( .A1(npu_inst_n56), .A2(
        npu_inst_int_data_y_4__5__0_), .B1(npu_inst_pe_1_3_5_n3), .B2(
        npu_inst_int_data_x_3__6__0_), .ZN(npu_inst_pe_1_3_5_n61) );
  INV_X1 npu_inst_pe_1_3_5_U30 ( .A(npu_inst_pe_1_3_5_int_data_0_), .ZN(
        npu_inst_pe_1_3_5_n13) );
  INV_X1 npu_inst_pe_1_3_5_U29 ( .A(npu_inst_n69), .ZN(npu_inst_pe_1_3_5_n5)
         );
  OR3_X1 npu_inst_pe_1_3_5_U28 ( .A1(npu_inst_pe_1_3_5_n6), .A2(
        npu_inst_pe_1_3_5_n8), .A3(npu_inst_pe_1_3_5_n5), .ZN(
        npu_inst_pe_1_3_5_n56) );
  OR3_X1 npu_inst_pe_1_3_5_U27 ( .A1(npu_inst_pe_1_3_5_n5), .A2(
        npu_inst_pe_1_3_5_n8), .A3(npu_inst_pe_1_3_5_n7), .ZN(
        npu_inst_pe_1_3_5_n48) );
  INV_X1 npu_inst_pe_1_3_5_U26 ( .A(npu_inst_pe_1_3_5_n5), .ZN(
        npu_inst_pe_1_3_5_n4) );
  INV_X1 npu_inst_pe_1_3_5_U25 ( .A(npu_inst_n124), .ZN(npu_inst_pe_1_3_5_n12)
         );
  OR3_X1 npu_inst_pe_1_3_5_U24 ( .A1(npu_inst_pe_1_3_5_n4), .A2(
        npu_inst_pe_1_3_5_n8), .A3(npu_inst_pe_1_3_5_n7), .ZN(
        npu_inst_pe_1_3_5_n52) );
  OR3_X1 npu_inst_pe_1_3_5_U23 ( .A1(npu_inst_pe_1_3_5_n6), .A2(
        npu_inst_pe_1_3_5_n8), .A3(npu_inst_pe_1_3_5_n4), .ZN(
        npu_inst_pe_1_3_5_n60) );
  NOR2_X1 npu_inst_pe_1_3_5_U22 ( .A1(npu_inst_pe_1_3_5_n60), .A2(
        npu_inst_pe_1_3_5_n3), .ZN(npu_inst_pe_1_3_5_n58) );
  NOR2_X1 npu_inst_pe_1_3_5_U21 ( .A1(npu_inst_pe_1_3_5_n56), .A2(
        npu_inst_pe_1_3_5_n3), .ZN(npu_inst_pe_1_3_5_n54) );
  NOR2_X1 npu_inst_pe_1_3_5_U20 ( .A1(npu_inst_pe_1_3_5_n52), .A2(
        npu_inst_pe_1_3_5_n3), .ZN(npu_inst_pe_1_3_5_n50) );
  NOR2_X1 npu_inst_pe_1_3_5_U19 ( .A1(npu_inst_pe_1_3_5_n48), .A2(
        npu_inst_pe_1_3_5_n3), .ZN(npu_inst_pe_1_3_5_n46) );
  NOR2_X1 npu_inst_pe_1_3_5_U18 ( .A1(npu_inst_pe_1_3_5_n40), .A2(
        npu_inst_pe_1_3_5_n3), .ZN(npu_inst_pe_1_3_5_n38) );
  NOR2_X1 npu_inst_pe_1_3_5_U17 ( .A1(npu_inst_pe_1_3_5_n44), .A2(
        npu_inst_pe_1_3_5_n3), .ZN(npu_inst_pe_1_3_5_n42) );
  BUF_X1 npu_inst_pe_1_3_5_U16 ( .A(npu_inst_n100), .Z(npu_inst_pe_1_3_5_n8)
         );
  BUF_X1 npu_inst_pe_1_3_5_U15 ( .A(npu_inst_pe_1_3_5_n12), .Z(
        npu_inst_pe_1_3_5_n11) );
  BUF_X1 npu_inst_pe_1_3_5_U14 ( .A(npu_inst_pe_1_3_5_n12), .Z(
        npu_inst_pe_1_3_5_n10) );
  BUF_X1 npu_inst_pe_1_3_5_U13 ( .A(npu_inst_pe_1_3_5_n12), .Z(
        npu_inst_pe_1_3_5_n9) );
  INV_X1 npu_inst_pe_1_3_5_U12 ( .A(npu_inst_pe_1_3_5_n38), .ZN(
        npu_inst_pe_1_3_5_n118) );
  INV_X1 npu_inst_pe_1_3_5_U11 ( .A(npu_inst_pe_1_3_5_n58), .ZN(
        npu_inst_pe_1_3_5_n114) );
  INV_X1 npu_inst_pe_1_3_5_U10 ( .A(npu_inst_pe_1_3_5_n54), .ZN(
        npu_inst_pe_1_3_5_n115) );
  INV_X1 npu_inst_pe_1_3_5_U9 ( .A(npu_inst_pe_1_3_5_n50), .ZN(
        npu_inst_pe_1_3_5_n116) );
  INV_X1 npu_inst_pe_1_3_5_U8 ( .A(npu_inst_pe_1_3_5_n46), .ZN(
        npu_inst_pe_1_3_5_n117) );
  INV_X1 npu_inst_pe_1_3_5_U7 ( .A(npu_inst_pe_1_3_5_n42), .ZN(
        npu_inst_pe_1_3_5_n119) );
  BUF_X1 npu_inst_pe_1_3_5_U6 ( .A(npu_inst_n24), .Z(npu_inst_pe_1_3_5_n2) );
  BUF_X1 npu_inst_pe_1_3_5_U5 ( .A(npu_inst_n24), .Z(npu_inst_pe_1_3_5_n1) );
  NOR2_X1 npu_inst_pe_1_3_5_U4 ( .A1(npu_inst_pe_1_3_5_int_q_weight_0_), .A2(
        npu_inst_pe_1_3_5_n1), .ZN(npu_inst_pe_1_3_5_n76) );
  NOR2_X1 npu_inst_pe_1_3_5_U3 ( .A1(npu_inst_pe_1_3_5_n27), .A2(
        npu_inst_pe_1_3_5_n1), .ZN(npu_inst_pe_1_3_5_n77) );
  FA_X1 npu_inst_pe_1_3_5_sub_77_U2_1 ( .A(npu_inst_pe_1_3_5_int_q_acc_1_), 
        .B(npu_inst_pe_1_3_5_n14), .CI(npu_inst_pe_1_3_5_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_3_5_sub_77_carry_2_), .S(npu_inst_pe_1_3_5_N66) );
  FA_X1 npu_inst_pe_1_3_5_add_79_U1_1 ( .A(npu_inst_pe_1_3_5_int_q_acc_1_), 
        .B(npu_inst_pe_1_3_5_int_data_1_), .CI(
        npu_inst_pe_1_3_5_add_79_carry_1_), .CO(
        npu_inst_pe_1_3_5_add_79_carry_2_), .S(npu_inst_pe_1_3_5_N74) );
  NAND3_X1 npu_inst_pe_1_3_5_U109 ( .A1(npu_inst_pe_1_3_5_n5), .A2(
        npu_inst_pe_1_3_5_n7), .A3(npu_inst_pe_1_3_5_n8), .ZN(
        npu_inst_pe_1_3_5_n44) );
  NAND3_X1 npu_inst_pe_1_3_5_U108 ( .A1(npu_inst_pe_1_3_5_n4), .A2(
        npu_inst_pe_1_3_5_n7), .A3(npu_inst_pe_1_3_5_n8), .ZN(
        npu_inst_pe_1_3_5_n40) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_3_5_n34), .CK(
        npu_inst_pe_1_3_5_net3626), .RN(npu_inst_pe_1_3_5_n9), .Q(
        npu_inst_pe_1_3_5_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_3_5_n35), .CK(
        npu_inst_pe_1_3_5_net3626), .RN(npu_inst_pe_1_3_5_n9), .Q(
        npu_inst_pe_1_3_5_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_3_5_n36), .CK(
        npu_inst_pe_1_3_5_net3626), .RN(npu_inst_pe_1_3_5_n9), .Q(
        npu_inst_pe_1_3_5_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_3_5_n98), .CK(
        npu_inst_pe_1_3_5_net3626), .RN(npu_inst_pe_1_3_5_n9), .Q(
        npu_inst_pe_1_3_5_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_3_5_n99), .CK(
        npu_inst_pe_1_3_5_net3626), .RN(npu_inst_pe_1_3_5_n9), .Q(
        npu_inst_pe_1_3_5_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_3_5_n100), 
        .CK(npu_inst_pe_1_3_5_net3626), .RN(npu_inst_pe_1_3_5_n9), .Q(
        npu_inst_pe_1_3_5_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_3_5_n33), .CK(
        npu_inst_pe_1_3_5_net3626), .RN(npu_inst_pe_1_3_5_n9), .Q(
        npu_inst_pe_1_3_5_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_3_5_n101), 
        .CK(npu_inst_pe_1_3_5_net3626), .RN(npu_inst_pe_1_3_5_n9), .Q(
        npu_inst_pe_1_3_5_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_weight_reg_0_ ( .D(npu_inst_n110), .CK(
        npu_inst_pe_1_3_5_net3632), .RN(npu_inst_pe_1_3_5_n9), .Q(
        npu_inst_pe_1_3_5_int_q_weight_0_), .QN(npu_inst_pe_1_3_5_n27) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_weight_reg_1_ ( .D(npu_inst_n116), .CK(
        npu_inst_pe_1_3_5_net3632), .RN(npu_inst_pe_1_3_5_n9), .Q(
        npu_inst_pe_1_3_5_int_q_weight_1_), .QN(npu_inst_pe_1_3_5_n26) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_3_5_n113), 
        .CK(npu_inst_pe_1_3_5_net3632), .RN(npu_inst_pe_1_3_5_n9), .Q(
        npu_inst_pe_1_3_5_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_3_5_n107), 
        .CK(npu_inst_pe_1_3_5_net3632), .RN(npu_inst_pe_1_3_5_n9), .Q(
        npu_inst_pe_1_3_5_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_3_5_n112), 
        .CK(npu_inst_pe_1_3_5_net3632), .RN(npu_inst_pe_1_3_5_n10), .Q(
        npu_inst_pe_1_3_5_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_3_5_n106), 
        .CK(npu_inst_pe_1_3_5_net3632), .RN(npu_inst_pe_1_3_5_n10), .Q(
        npu_inst_pe_1_3_5_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_3_5_n111), 
        .CK(npu_inst_pe_1_3_5_net3632), .RN(npu_inst_pe_1_3_5_n10), .Q(
        npu_inst_pe_1_3_5_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_3_5_n105), 
        .CK(npu_inst_pe_1_3_5_net3632), .RN(npu_inst_pe_1_3_5_n10), .Q(
        npu_inst_pe_1_3_5_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_3_5_n110), 
        .CK(npu_inst_pe_1_3_5_net3632), .RN(npu_inst_pe_1_3_5_n10), .Q(
        npu_inst_pe_1_3_5_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_3_5_n104), 
        .CK(npu_inst_pe_1_3_5_net3632), .RN(npu_inst_pe_1_3_5_n10), .Q(
        npu_inst_pe_1_3_5_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_3_5_n109), 
        .CK(npu_inst_pe_1_3_5_net3632), .RN(npu_inst_pe_1_3_5_n10), .Q(
        npu_inst_pe_1_3_5_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_3_5_n103), 
        .CK(npu_inst_pe_1_3_5_net3632), .RN(npu_inst_pe_1_3_5_n10), .Q(
        npu_inst_pe_1_3_5_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_3_5_n108), 
        .CK(npu_inst_pe_1_3_5_net3632), .RN(npu_inst_pe_1_3_5_n10), .Q(
        npu_inst_pe_1_3_5_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_3_5_n102), 
        .CK(npu_inst_pe_1_3_5_net3632), .RN(npu_inst_pe_1_3_5_n10), .Q(
        npu_inst_pe_1_3_5_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_3_5_n86), 
        .CK(npu_inst_pe_1_3_5_net3632), .RN(npu_inst_pe_1_3_5_n10), .Q(
        npu_inst_pe_1_3_5_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_3_5_n87), 
        .CK(npu_inst_pe_1_3_5_net3632), .RN(npu_inst_pe_1_3_5_n10), .Q(
        npu_inst_pe_1_3_5_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_3_5_n88), 
        .CK(npu_inst_pe_1_3_5_net3632), .RN(npu_inst_pe_1_3_5_n11), .Q(
        npu_inst_pe_1_3_5_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_3_5_n89), 
        .CK(npu_inst_pe_1_3_5_net3632), .RN(npu_inst_pe_1_3_5_n11), .Q(
        npu_inst_pe_1_3_5_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_3_5_n90), 
        .CK(npu_inst_pe_1_3_5_net3632), .RN(npu_inst_pe_1_3_5_n11), .Q(
        npu_inst_pe_1_3_5_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_3_5_n91), 
        .CK(npu_inst_pe_1_3_5_net3632), .RN(npu_inst_pe_1_3_5_n11), .Q(
        npu_inst_pe_1_3_5_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_3_5_n92), 
        .CK(npu_inst_pe_1_3_5_net3632), .RN(npu_inst_pe_1_3_5_n11), .Q(
        npu_inst_pe_1_3_5_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_3_5_n93), 
        .CK(npu_inst_pe_1_3_5_net3632), .RN(npu_inst_pe_1_3_5_n11), .Q(
        npu_inst_pe_1_3_5_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_3_5_n94), 
        .CK(npu_inst_pe_1_3_5_net3632), .RN(npu_inst_pe_1_3_5_n11), .Q(
        npu_inst_pe_1_3_5_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_3_5_n95), 
        .CK(npu_inst_pe_1_3_5_net3632), .RN(npu_inst_pe_1_3_5_n11), .Q(
        npu_inst_pe_1_3_5_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_3_5_n96), 
        .CK(npu_inst_pe_1_3_5_net3632), .RN(npu_inst_pe_1_3_5_n11), .Q(
        npu_inst_pe_1_3_5_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_3_5_n97), 
        .CK(npu_inst_pe_1_3_5_net3632), .RN(npu_inst_pe_1_3_5_n11), .Q(
        npu_inst_pe_1_3_5_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_3_5_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_3_5_N84), .SE(1'b0), .GCK(npu_inst_pe_1_3_5_net3626) );
  CLKGATETST_X1 npu_inst_pe_1_3_5_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n64), .SE(1'b0), .GCK(npu_inst_pe_1_3_5_net3632) );
  MUX2_X1 npu_inst_pe_1_3_6_U162 ( .A(npu_inst_pe_1_3_6_n32), .B(
        npu_inst_pe_1_3_6_n29), .S(npu_inst_pe_1_3_6_n8), .Z(
        npu_inst_pe_1_3_6_N93) );
  MUX2_X1 npu_inst_pe_1_3_6_U161 ( .A(npu_inst_pe_1_3_6_n31), .B(
        npu_inst_pe_1_3_6_n30), .S(npu_inst_pe_1_3_6_n6), .Z(
        npu_inst_pe_1_3_6_n32) );
  MUX2_X1 npu_inst_pe_1_3_6_U160 ( .A(npu_inst_pe_1_3_6_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_3_6_int_q_reg_v_1__0_), .S(npu_inst_pe_1_3_6_n4), .Z(
        npu_inst_pe_1_3_6_n31) );
  MUX2_X1 npu_inst_pe_1_3_6_U159 ( .A(npu_inst_pe_1_3_6_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_3_6_int_q_reg_v_3__0_), .S(npu_inst_pe_1_3_6_n4), .Z(
        npu_inst_pe_1_3_6_n30) );
  MUX2_X1 npu_inst_pe_1_3_6_U158 ( .A(npu_inst_pe_1_3_6_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_3_6_int_q_reg_v_5__0_), .S(npu_inst_pe_1_3_6_n4), .Z(
        npu_inst_pe_1_3_6_n29) );
  MUX2_X1 npu_inst_pe_1_3_6_U157 ( .A(npu_inst_pe_1_3_6_n28), .B(
        npu_inst_pe_1_3_6_n23), .S(npu_inst_pe_1_3_6_n8), .Z(
        npu_inst_pe_1_3_6_N94) );
  MUX2_X1 npu_inst_pe_1_3_6_U156 ( .A(npu_inst_pe_1_3_6_n25), .B(
        npu_inst_pe_1_3_6_n24), .S(npu_inst_pe_1_3_6_n6), .Z(
        npu_inst_pe_1_3_6_n28) );
  MUX2_X1 npu_inst_pe_1_3_6_U155 ( .A(npu_inst_pe_1_3_6_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_3_6_int_q_reg_v_1__1_), .S(npu_inst_pe_1_3_6_n4), .Z(
        npu_inst_pe_1_3_6_n25) );
  MUX2_X1 npu_inst_pe_1_3_6_U154 ( .A(npu_inst_pe_1_3_6_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_3_6_int_q_reg_v_3__1_), .S(npu_inst_pe_1_3_6_n4), .Z(
        npu_inst_pe_1_3_6_n24) );
  MUX2_X1 npu_inst_pe_1_3_6_U153 ( .A(npu_inst_pe_1_3_6_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_3_6_int_q_reg_v_5__1_), .S(npu_inst_pe_1_3_6_n4), .Z(
        npu_inst_pe_1_3_6_n23) );
  MUX2_X1 npu_inst_pe_1_3_6_U152 ( .A(npu_inst_pe_1_3_6_n22), .B(
        npu_inst_pe_1_3_6_n19), .S(npu_inst_pe_1_3_6_n8), .Z(
        npu_inst_int_data_x_3__6__1_) );
  MUX2_X1 npu_inst_pe_1_3_6_U151 ( .A(npu_inst_pe_1_3_6_n21), .B(
        npu_inst_pe_1_3_6_n20), .S(npu_inst_pe_1_3_6_n6), .Z(
        npu_inst_pe_1_3_6_n22) );
  MUX2_X1 npu_inst_pe_1_3_6_U150 ( .A(npu_inst_pe_1_3_6_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_3_6_int_q_reg_h_1__1_), .S(npu_inst_pe_1_3_6_n4), .Z(
        npu_inst_pe_1_3_6_n21) );
  MUX2_X1 npu_inst_pe_1_3_6_U149 ( .A(npu_inst_pe_1_3_6_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_3_6_int_q_reg_h_3__1_), .S(npu_inst_pe_1_3_6_n4), .Z(
        npu_inst_pe_1_3_6_n20) );
  MUX2_X1 npu_inst_pe_1_3_6_U148 ( .A(npu_inst_pe_1_3_6_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_3_6_int_q_reg_h_5__1_), .S(npu_inst_pe_1_3_6_n4), .Z(
        npu_inst_pe_1_3_6_n19) );
  MUX2_X1 npu_inst_pe_1_3_6_U147 ( .A(npu_inst_pe_1_3_6_n18), .B(
        npu_inst_pe_1_3_6_n15), .S(npu_inst_pe_1_3_6_n8), .Z(
        npu_inst_int_data_x_3__6__0_) );
  MUX2_X1 npu_inst_pe_1_3_6_U146 ( .A(npu_inst_pe_1_3_6_n17), .B(
        npu_inst_pe_1_3_6_n16), .S(npu_inst_pe_1_3_6_n6), .Z(
        npu_inst_pe_1_3_6_n18) );
  MUX2_X1 npu_inst_pe_1_3_6_U145 ( .A(npu_inst_pe_1_3_6_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_3_6_int_q_reg_h_1__0_), .S(npu_inst_pe_1_3_6_n4), .Z(
        npu_inst_pe_1_3_6_n17) );
  MUX2_X1 npu_inst_pe_1_3_6_U144 ( .A(npu_inst_pe_1_3_6_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_3_6_int_q_reg_h_3__0_), .S(npu_inst_pe_1_3_6_n4), .Z(
        npu_inst_pe_1_3_6_n16) );
  MUX2_X1 npu_inst_pe_1_3_6_U143 ( .A(npu_inst_pe_1_3_6_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_3_6_int_q_reg_h_5__0_), .S(npu_inst_pe_1_3_6_n4), .Z(
        npu_inst_pe_1_3_6_n15) );
  XOR2_X1 npu_inst_pe_1_3_6_U142 ( .A(npu_inst_pe_1_3_6_int_data_0_), .B(
        npu_inst_pe_1_3_6_int_q_acc_0_), .Z(npu_inst_pe_1_3_6_N73) );
  AND2_X1 npu_inst_pe_1_3_6_U141 ( .A1(npu_inst_pe_1_3_6_int_q_acc_0_), .A2(
        npu_inst_pe_1_3_6_int_data_0_), .ZN(npu_inst_pe_1_3_6_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_3_6_U140 ( .A(npu_inst_pe_1_3_6_int_q_acc_0_), .B(
        npu_inst_pe_1_3_6_n13), .ZN(npu_inst_pe_1_3_6_N65) );
  OR2_X1 npu_inst_pe_1_3_6_U139 ( .A1(npu_inst_pe_1_3_6_n13), .A2(
        npu_inst_pe_1_3_6_int_q_acc_0_), .ZN(npu_inst_pe_1_3_6_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_3_6_U138 ( .A(npu_inst_pe_1_3_6_int_q_acc_2_), .B(
        npu_inst_pe_1_3_6_add_79_carry_2_), .Z(npu_inst_pe_1_3_6_N75) );
  AND2_X1 npu_inst_pe_1_3_6_U137 ( .A1(npu_inst_pe_1_3_6_add_79_carry_2_), 
        .A2(npu_inst_pe_1_3_6_int_q_acc_2_), .ZN(
        npu_inst_pe_1_3_6_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_3_6_U136 ( .A(npu_inst_pe_1_3_6_int_q_acc_3_), .B(
        npu_inst_pe_1_3_6_add_79_carry_3_), .Z(npu_inst_pe_1_3_6_N76) );
  AND2_X1 npu_inst_pe_1_3_6_U135 ( .A1(npu_inst_pe_1_3_6_add_79_carry_3_), 
        .A2(npu_inst_pe_1_3_6_int_q_acc_3_), .ZN(
        npu_inst_pe_1_3_6_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_3_6_U134 ( .A(npu_inst_pe_1_3_6_int_q_acc_4_), .B(
        npu_inst_pe_1_3_6_add_79_carry_4_), .Z(npu_inst_pe_1_3_6_N77) );
  AND2_X1 npu_inst_pe_1_3_6_U133 ( .A1(npu_inst_pe_1_3_6_add_79_carry_4_), 
        .A2(npu_inst_pe_1_3_6_int_q_acc_4_), .ZN(
        npu_inst_pe_1_3_6_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_3_6_U132 ( .A(npu_inst_pe_1_3_6_int_q_acc_5_), .B(
        npu_inst_pe_1_3_6_add_79_carry_5_), .Z(npu_inst_pe_1_3_6_N78) );
  AND2_X1 npu_inst_pe_1_3_6_U131 ( .A1(npu_inst_pe_1_3_6_add_79_carry_5_), 
        .A2(npu_inst_pe_1_3_6_int_q_acc_5_), .ZN(
        npu_inst_pe_1_3_6_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_3_6_U130 ( .A(npu_inst_pe_1_3_6_int_q_acc_6_), .B(
        npu_inst_pe_1_3_6_add_79_carry_6_), .Z(npu_inst_pe_1_3_6_N79) );
  AND2_X1 npu_inst_pe_1_3_6_U129 ( .A1(npu_inst_pe_1_3_6_add_79_carry_6_), 
        .A2(npu_inst_pe_1_3_6_int_q_acc_6_), .ZN(
        npu_inst_pe_1_3_6_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_3_6_U128 ( .A(npu_inst_pe_1_3_6_int_q_acc_7_), .B(
        npu_inst_pe_1_3_6_add_79_carry_7_), .Z(npu_inst_pe_1_3_6_N80) );
  XNOR2_X1 npu_inst_pe_1_3_6_U127 ( .A(npu_inst_pe_1_3_6_sub_77_carry_2_), .B(
        npu_inst_pe_1_3_6_int_q_acc_2_), .ZN(npu_inst_pe_1_3_6_N67) );
  OR2_X1 npu_inst_pe_1_3_6_U126 ( .A1(npu_inst_pe_1_3_6_int_q_acc_2_), .A2(
        npu_inst_pe_1_3_6_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_3_6_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_3_6_U125 ( .A(npu_inst_pe_1_3_6_sub_77_carry_3_), .B(
        npu_inst_pe_1_3_6_int_q_acc_3_), .ZN(npu_inst_pe_1_3_6_N68) );
  OR2_X1 npu_inst_pe_1_3_6_U124 ( .A1(npu_inst_pe_1_3_6_int_q_acc_3_), .A2(
        npu_inst_pe_1_3_6_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_3_6_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_3_6_U123 ( .A(npu_inst_pe_1_3_6_sub_77_carry_4_), .B(
        npu_inst_pe_1_3_6_int_q_acc_4_), .ZN(npu_inst_pe_1_3_6_N69) );
  OR2_X1 npu_inst_pe_1_3_6_U122 ( .A1(npu_inst_pe_1_3_6_int_q_acc_4_), .A2(
        npu_inst_pe_1_3_6_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_3_6_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_3_6_U121 ( .A(npu_inst_pe_1_3_6_sub_77_carry_5_), .B(
        npu_inst_pe_1_3_6_int_q_acc_5_), .ZN(npu_inst_pe_1_3_6_N70) );
  OR2_X1 npu_inst_pe_1_3_6_U120 ( .A1(npu_inst_pe_1_3_6_int_q_acc_5_), .A2(
        npu_inst_pe_1_3_6_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_3_6_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_3_6_U119 ( .A(npu_inst_pe_1_3_6_sub_77_carry_6_), .B(
        npu_inst_pe_1_3_6_int_q_acc_6_), .ZN(npu_inst_pe_1_3_6_N71) );
  OR2_X1 npu_inst_pe_1_3_6_U118 ( .A1(npu_inst_pe_1_3_6_int_q_acc_6_), .A2(
        npu_inst_pe_1_3_6_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_3_6_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_3_6_U117 ( .A(npu_inst_pe_1_3_6_int_q_acc_7_), .B(
        npu_inst_pe_1_3_6_sub_77_carry_7_), .ZN(npu_inst_pe_1_3_6_N72) );
  INV_X1 npu_inst_pe_1_3_6_U116 ( .A(npu_inst_n77), .ZN(npu_inst_pe_1_3_6_n7)
         );
  INV_X1 npu_inst_pe_1_3_6_U115 ( .A(npu_inst_pe_1_3_6_n7), .ZN(
        npu_inst_pe_1_3_6_n6) );
  INV_X1 npu_inst_pe_1_3_6_U114 ( .A(npu_inst_n56), .ZN(npu_inst_pe_1_3_6_n3)
         );
  AOI22_X1 npu_inst_pe_1_3_6_U113 ( .A1(npu_inst_int_data_y_4__6__0_), .A2(
        npu_inst_pe_1_3_6_n58), .B1(npu_inst_pe_1_3_6_n114), .B2(
        npu_inst_pe_1_3_6_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_3_6_n57) );
  INV_X1 npu_inst_pe_1_3_6_U112 ( .A(npu_inst_pe_1_3_6_n57), .ZN(
        npu_inst_pe_1_3_6_n108) );
  AOI22_X1 npu_inst_pe_1_3_6_U111 ( .A1(npu_inst_int_data_y_4__6__0_), .A2(
        npu_inst_pe_1_3_6_n54), .B1(npu_inst_pe_1_3_6_n115), .B2(
        npu_inst_pe_1_3_6_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_3_6_n53) );
  INV_X1 npu_inst_pe_1_3_6_U110 ( .A(npu_inst_pe_1_3_6_n53), .ZN(
        npu_inst_pe_1_3_6_n109) );
  AOI22_X1 npu_inst_pe_1_3_6_U107 ( .A1(npu_inst_int_data_y_4__6__0_), .A2(
        npu_inst_pe_1_3_6_n50), .B1(npu_inst_pe_1_3_6_n116), .B2(
        npu_inst_pe_1_3_6_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_3_6_n49) );
  INV_X1 npu_inst_pe_1_3_6_U106 ( .A(npu_inst_pe_1_3_6_n49), .ZN(
        npu_inst_pe_1_3_6_n110) );
  AOI22_X1 npu_inst_pe_1_3_6_U105 ( .A1(npu_inst_int_data_y_4__6__0_), .A2(
        npu_inst_pe_1_3_6_n46), .B1(npu_inst_pe_1_3_6_n117), .B2(
        npu_inst_pe_1_3_6_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_3_6_n45) );
  INV_X1 npu_inst_pe_1_3_6_U104 ( .A(npu_inst_pe_1_3_6_n45), .ZN(
        npu_inst_pe_1_3_6_n111) );
  AOI22_X1 npu_inst_pe_1_3_6_U103 ( .A1(npu_inst_int_data_y_4__6__0_), .A2(
        npu_inst_pe_1_3_6_n42), .B1(npu_inst_pe_1_3_6_n119), .B2(
        npu_inst_pe_1_3_6_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_3_6_n41) );
  INV_X1 npu_inst_pe_1_3_6_U102 ( .A(npu_inst_pe_1_3_6_n41), .ZN(
        npu_inst_pe_1_3_6_n112) );
  AOI22_X1 npu_inst_pe_1_3_6_U101 ( .A1(npu_inst_int_data_y_4__6__1_), .A2(
        npu_inst_pe_1_3_6_n58), .B1(npu_inst_pe_1_3_6_n114), .B2(
        npu_inst_pe_1_3_6_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_3_6_n59) );
  INV_X1 npu_inst_pe_1_3_6_U100 ( .A(npu_inst_pe_1_3_6_n59), .ZN(
        npu_inst_pe_1_3_6_n102) );
  AOI22_X1 npu_inst_pe_1_3_6_U99 ( .A1(npu_inst_int_data_y_4__6__1_), .A2(
        npu_inst_pe_1_3_6_n54), .B1(npu_inst_pe_1_3_6_n115), .B2(
        npu_inst_pe_1_3_6_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_3_6_n55) );
  INV_X1 npu_inst_pe_1_3_6_U98 ( .A(npu_inst_pe_1_3_6_n55), .ZN(
        npu_inst_pe_1_3_6_n103) );
  AOI22_X1 npu_inst_pe_1_3_6_U97 ( .A1(npu_inst_int_data_y_4__6__1_), .A2(
        npu_inst_pe_1_3_6_n50), .B1(npu_inst_pe_1_3_6_n116), .B2(
        npu_inst_pe_1_3_6_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_3_6_n51) );
  INV_X1 npu_inst_pe_1_3_6_U96 ( .A(npu_inst_pe_1_3_6_n51), .ZN(
        npu_inst_pe_1_3_6_n104) );
  AOI22_X1 npu_inst_pe_1_3_6_U95 ( .A1(npu_inst_int_data_y_4__6__1_), .A2(
        npu_inst_pe_1_3_6_n46), .B1(npu_inst_pe_1_3_6_n117), .B2(
        npu_inst_pe_1_3_6_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_3_6_n47) );
  INV_X1 npu_inst_pe_1_3_6_U94 ( .A(npu_inst_pe_1_3_6_n47), .ZN(
        npu_inst_pe_1_3_6_n105) );
  AOI22_X1 npu_inst_pe_1_3_6_U93 ( .A1(npu_inst_int_data_y_4__6__1_), .A2(
        npu_inst_pe_1_3_6_n42), .B1(npu_inst_pe_1_3_6_n119), .B2(
        npu_inst_pe_1_3_6_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_3_6_n43) );
  INV_X1 npu_inst_pe_1_3_6_U92 ( .A(npu_inst_pe_1_3_6_n43), .ZN(
        npu_inst_pe_1_3_6_n106) );
  AOI22_X1 npu_inst_pe_1_3_6_U91 ( .A1(npu_inst_pe_1_3_6_n38), .A2(
        npu_inst_int_data_y_4__6__1_), .B1(npu_inst_pe_1_3_6_n118), .B2(
        npu_inst_pe_1_3_6_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_3_6_n39) );
  INV_X1 npu_inst_pe_1_3_6_U90 ( .A(npu_inst_pe_1_3_6_n39), .ZN(
        npu_inst_pe_1_3_6_n107) );
  AOI22_X1 npu_inst_pe_1_3_6_U89 ( .A1(npu_inst_pe_1_3_6_n38), .A2(
        npu_inst_int_data_y_4__6__0_), .B1(npu_inst_pe_1_3_6_n118), .B2(
        npu_inst_pe_1_3_6_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_3_6_n37) );
  INV_X1 npu_inst_pe_1_3_6_U88 ( .A(npu_inst_pe_1_3_6_n37), .ZN(
        npu_inst_pe_1_3_6_n113) );
  NAND2_X1 npu_inst_pe_1_3_6_U87 ( .A1(npu_inst_pe_1_3_6_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_3_6_n60), .ZN(npu_inst_pe_1_3_6_n74) );
  OAI21_X1 npu_inst_pe_1_3_6_U86 ( .B1(npu_inst_pe_1_3_6_n63), .B2(
        npu_inst_pe_1_3_6_n60), .A(npu_inst_pe_1_3_6_n74), .ZN(
        npu_inst_pe_1_3_6_n97) );
  NAND2_X1 npu_inst_pe_1_3_6_U85 ( .A1(npu_inst_pe_1_3_6_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_3_6_n60), .ZN(npu_inst_pe_1_3_6_n73) );
  OAI21_X1 npu_inst_pe_1_3_6_U84 ( .B1(npu_inst_pe_1_3_6_n61), .B2(
        npu_inst_pe_1_3_6_n60), .A(npu_inst_pe_1_3_6_n73), .ZN(
        npu_inst_pe_1_3_6_n96) );
  NAND2_X1 npu_inst_pe_1_3_6_U83 ( .A1(npu_inst_pe_1_3_6_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_3_6_n56), .ZN(npu_inst_pe_1_3_6_n72) );
  OAI21_X1 npu_inst_pe_1_3_6_U82 ( .B1(npu_inst_pe_1_3_6_n63), .B2(
        npu_inst_pe_1_3_6_n56), .A(npu_inst_pe_1_3_6_n72), .ZN(
        npu_inst_pe_1_3_6_n95) );
  NAND2_X1 npu_inst_pe_1_3_6_U81 ( .A1(npu_inst_pe_1_3_6_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_3_6_n56), .ZN(npu_inst_pe_1_3_6_n71) );
  OAI21_X1 npu_inst_pe_1_3_6_U80 ( .B1(npu_inst_pe_1_3_6_n61), .B2(
        npu_inst_pe_1_3_6_n56), .A(npu_inst_pe_1_3_6_n71), .ZN(
        npu_inst_pe_1_3_6_n94) );
  NAND2_X1 npu_inst_pe_1_3_6_U79 ( .A1(npu_inst_pe_1_3_6_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_3_6_n52), .ZN(npu_inst_pe_1_3_6_n70) );
  OAI21_X1 npu_inst_pe_1_3_6_U78 ( .B1(npu_inst_pe_1_3_6_n63), .B2(
        npu_inst_pe_1_3_6_n52), .A(npu_inst_pe_1_3_6_n70), .ZN(
        npu_inst_pe_1_3_6_n93) );
  NAND2_X1 npu_inst_pe_1_3_6_U77 ( .A1(npu_inst_pe_1_3_6_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_3_6_n52), .ZN(npu_inst_pe_1_3_6_n69) );
  OAI21_X1 npu_inst_pe_1_3_6_U76 ( .B1(npu_inst_pe_1_3_6_n61), .B2(
        npu_inst_pe_1_3_6_n52), .A(npu_inst_pe_1_3_6_n69), .ZN(
        npu_inst_pe_1_3_6_n92) );
  NAND2_X1 npu_inst_pe_1_3_6_U75 ( .A1(npu_inst_pe_1_3_6_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_3_6_n48), .ZN(npu_inst_pe_1_3_6_n68) );
  OAI21_X1 npu_inst_pe_1_3_6_U74 ( .B1(npu_inst_pe_1_3_6_n63), .B2(
        npu_inst_pe_1_3_6_n48), .A(npu_inst_pe_1_3_6_n68), .ZN(
        npu_inst_pe_1_3_6_n91) );
  NAND2_X1 npu_inst_pe_1_3_6_U73 ( .A1(npu_inst_pe_1_3_6_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_3_6_n48), .ZN(npu_inst_pe_1_3_6_n67) );
  OAI21_X1 npu_inst_pe_1_3_6_U72 ( .B1(npu_inst_pe_1_3_6_n61), .B2(
        npu_inst_pe_1_3_6_n48), .A(npu_inst_pe_1_3_6_n67), .ZN(
        npu_inst_pe_1_3_6_n90) );
  NAND2_X1 npu_inst_pe_1_3_6_U71 ( .A1(npu_inst_pe_1_3_6_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_3_6_n44), .ZN(npu_inst_pe_1_3_6_n66) );
  OAI21_X1 npu_inst_pe_1_3_6_U70 ( .B1(npu_inst_pe_1_3_6_n63), .B2(
        npu_inst_pe_1_3_6_n44), .A(npu_inst_pe_1_3_6_n66), .ZN(
        npu_inst_pe_1_3_6_n89) );
  NAND2_X1 npu_inst_pe_1_3_6_U69 ( .A1(npu_inst_pe_1_3_6_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_3_6_n44), .ZN(npu_inst_pe_1_3_6_n65) );
  OAI21_X1 npu_inst_pe_1_3_6_U68 ( .B1(npu_inst_pe_1_3_6_n61), .B2(
        npu_inst_pe_1_3_6_n44), .A(npu_inst_pe_1_3_6_n65), .ZN(
        npu_inst_pe_1_3_6_n88) );
  NAND2_X1 npu_inst_pe_1_3_6_U67 ( .A1(npu_inst_pe_1_3_6_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_3_6_n40), .ZN(npu_inst_pe_1_3_6_n64) );
  OAI21_X1 npu_inst_pe_1_3_6_U66 ( .B1(npu_inst_pe_1_3_6_n63), .B2(
        npu_inst_pe_1_3_6_n40), .A(npu_inst_pe_1_3_6_n64), .ZN(
        npu_inst_pe_1_3_6_n87) );
  NAND2_X1 npu_inst_pe_1_3_6_U65 ( .A1(npu_inst_pe_1_3_6_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_3_6_n40), .ZN(npu_inst_pe_1_3_6_n62) );
  OAI21_X1 npu_inst_pe_1_3_6_U64 ( .B1(npu_inst_pe_1_3_6_n61), .B2(
        npu_inst_pe_1_3_6_n40), .A(npu_inst_pe_1_3_6_n62), .ZN(
        npu_inst_pe_1_3_6_n86) );
  AND2_X1 npu_inst_pe_1_3_6_U63 ( .A1(npu_inst_pe_1_3_6_N93), .A2(npu_inst_n56), .ZN(npu_inst_int_data_y_3__6__0_) );
  AND2_X1 npu_inst_pe_1_3_6_U62 ( .A1(npu_inst_n56), .A2(npu_inst_pe_1_3_6_N94), .ZN(npu_inst_int_data_y_3__6__1_) );
  NOR3_X1 npu_inst_pe_1_3_6_U61 ( .A1(npu_inst_pe_1_3_6_n26), .A2(npu_inst_n56), .A3(npu_inst_int_ckg[33]), .ZN(npu_inst_pe_1_3_6_n85) );
  OR2_X1 npu_inst_pe_1_3_6_U60 ( .A1(npu_inst_pe_1_3_6_n85), .A2(
        npu_inst_pe_1_3_6_n2), .ZN(npu_inst_pe_1_3_6_N84) );
  AND2_X1 npu_inst_pe_1_3_6_U59 ( .A1(npu_inst_pe_1_3_6_int_q_acc_0_), .A2(
        npu_inst_pe_1_3_6_n1), .ZN(npu_inst_int_data_res_3__6__0_) );
  AND2_X1 npu_inst_pe_1_3_6_U58 ( .A1(npu_inst_pe_1_3_6_n2), .A2(
        npu_inst_pe_1_3_6_int_q_acc_7_), .ZN(npu_inst_int_data_res_3__6__7_)
         );
  AND2_X1 npu_inst_pe_1_3_6_U57 ( .A1(npu_inst_pe_1_3_6_int_q_acc_1_), .A2(
        npu_inst_pe_1_3_6_n1), .ZN(npu_inst_int_data_res_3__6__1_) );
  AND2_X1 npu_inst_pe_1_3_6_U56 ( .A1(npu_inst_pe_1_3_6_int_q_acc_2_), .A2(
        npu_inst_pe_1_3_6_n1), .ZN(npu_inst_int_data_res_3__6__2_) );
  AND2_X1 npu_inst_pe_1_3_6_U55 ( .A1(npu_inst_pe_1_3_6_int_q_acc_3_), .A2(
        npu_inst_pe_1_3_6_n2), .ZN(npu_inst_int_data_res_3__6__3_) );
  AND2_X1 npu_inst_pe_1_3_6_U54 ( .A1(npu_inst_pe_1_3_6_int_q_acc_4_), .A2(
        npu_inst_pe_1_3_6_n2), .ZN(npu_inst_int_data_res_3__6__4_) );
  AND2_X1 npu_inst_pe_1_3_6_U53 ( .A1(npu_inst_pe_1_3_6_int_q_acc_5_), .A2(
        npu_inst_pe_1_3_6_n2), .ZN(npu_inst_int_data_res_3__6__5_) );
  AND2_X1 npu_inst_pe_1_3_6_U52 ( .A1(npu_inst_pe_1_3_6_int_q_acc_6_), .A2(
        npu_inst_pe_1_3_6_n2), .ZN(npu_inst_int_data_res_3__6__6_) );
  AOI222_X1 npu_inst_pe_1_3_6_U51 ( .A1(npu_inst_int_data_res_4__6__0_), .A2(
        npu_inst_pe_1_3_6_n1), .B1(npu_inst_pe_1_3_6_N73), .B2(
        npu_inst_pe_1_3_6_n76), .C1(npu_inst_pe_1_3_6_N65), .C2(
        npu_inst_pe_1_3_6_n77), .ZN(npu_inst_pe_1_3_6_n84) );
  INV_X1 npu_inst_pe_1_3_6_U50 ( .A(npu_inst_pe_1_3_6_n84), .ZN(
        npu_inst_pe_1_3_6_n101) );
  AOI222_X1 npu_inst_pe_1_3_6_U49 ( .A1(npu_inst_int_data_res_4__6__7_), .A2(
        npu_inst_pe_1_3_6_n1), .B1(npu_inst_pe_1_3_6_N80), .B2(
        npu_inst_pe_1_3_6_n76), .C1(npu_inst_pe_1_3_6_N72), .C2(
        npu_inst_pe_1_3_6_n77), .ZN(npu_inst_pe_1_3_6_n75) );
  INV_X1 npu_inst_pe_1_3_6_U48 ( .A(npu_inst_pe_1_3_6_n75), .ZN(
        npu_inst_pe_1_3_6_n33) );
  AOI222_X1 npu_inst_pe_1_3_6_U47 ( .A1(npu_inst_int_data_res_4__6__1_), .A2(
        npu_inst_pe_1_3_6_n1), .B1(npu_inst_pe_1_3_6_N74), .B2(
        npu_inst_pe_1_3_6_n76), .C1(npu_inst_pe_1_3_6_N66), .C2(
        npu_inst_pe_1_3_6_n77), .ZN(npu_inst_pe_1_3_6_n83) );
  INV_X1 npu_inst_pe_1_3_6_U46 ( .A(npu_inst_pe_1_3_6_n83), .ZN(
        npu_inst_pe_1_3_6_n100) );
  AOI222_X1 npu_inst_pe_1_3_6_U45 ( .A1(npu_inst_int_data_res_4__6__2_), .A2(
        npu_inst_pe_1_3_6_n1), .B1(npu_inst_pe_1_3_6_N75), .B2(
        npu_inst_pe_1_3_6_n76), .C1(npu_inst_pe_1_3_6_N67), .C2(
        npu_inst_pe_1_3_6_n77), .ZN(npu_inst_pe_1_3_6_n82) );
  INV_X1 npu_inst_pe_1_3_6_U44 ( .A(npu_inst_pe_1_3_6_n82), .ZN(
        npu_inst_pe_1_3_6_n99) );
  AOI222_X1 npu_inst_pe_1_3_6_U43 ( .A1(npu_inst_int_data_res_4__6__3_), .A2(
        npu_inst_pe_1_3_6_n1), .B1(npu_inst_pe_1_3_6_N76), .B2(
        npu_inst_pe_1_3_6_n76), .C1(npu_inst_pe_1_3_6_N68), .C2(
        npu_inst_pe_1_3_6_n77), .ZN(npu_inst_pe_1_3_6_n81) );
  INV_X1 npu_inst_pe_1_3_6_U42 ( .A(npu_inst_pe_1_3_6_n81), .ZN(
        npu_inst_pe_1_3_6_n98) );
  AOI222_X1 npu_inst_pe_1_3_6_U41 ( .A1(npu_inst_int_data_res_4__6__4_), .A2(
        npu_inst_pe_1_3_6_n1), .B1(npu_inst_pe_1_3_6_N77), .B2(
        npu_inst_pe_1_3_6_n76), .C1(npu_inst_pe_1_3_6_N69), .C2(
        npu_inst_pe_1_3_6_n77), .ZN(npu_inst_pe_1_3_6_n80) );
  INV_X1 npu_inst_pe_1_3_6_U40 ( .A(npu_inst_pe_1_3_6_n80), .ZN(
        npu_inst_pe_1_3_6_n36) );
  AOI222_X1 npu_inst_pe_1_3_6_U39 ( .A1(npu_inst_int_data_res_4__6__5_), .A2(
        npu_inst_pe_1_3_6_n1), .B1(npu_inst_pe_1_3_6_N78), .B2(
        npu_inst_pe_1_3_6_n76), .C1(npu_inst_pe_1_3_6_N70), .C2(
        npu_inst_pe_1_3_6_n77), .ZN(npu_inst_pe_1_3_6_n79) );
  INV_X1 npu_inst_pe_1_3_6_U38 ( .A(npu_inst_pe_1_3_6_n79), .ZN(
        npu_inst_pe_1_3_6_n35) );
  AOI222_X1 npu_inst_pe_1_3_6_U37 ( .A1(npu_inst_int_data_res_4__6__6_), .A2(
        npu_inst_pe_1_3_6_n1), .B1(npu_inst_pe_1_3_6_N79), .B2(
        npu_inst_pe_1_3_6_n76), .C1(npu_inst_pe_1_3_6_N71), .C2(
        npu_inst_pe_1_3_6_n77), .ZN(npu_inst_pe_1_3_6_n78) );
  INV_X1 npu_inst_pe_1_3_6_U36 ( .A(npu_inst_pe_1_3_6_n78), .ZN(
        npu_inst_pe_1_3_6_n34) );
  INV_X1 npu_inst_pe_1_3_6_U35 ( .A(npu_inst_pe_1_3_6_int_data_1_), .ZN(
        npu_inst_pe_1_3_6_n14) );
  AND2_X1 npu_inst_pe_1_3_6_U34 ( .A1(npu_inst_int_data_x_3__6__1_), .A2(
        npu_inst_pe_1_3_6_int_q_weight_1_), .ZN(npu_inst_pe_1_3_6_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_3_6_U33 ( .A1(npu_inst_int_data_x_3__6__0_), .A2(
        npu_inst_pe_1_3_6_int_q_weight_1_), .ZN(npu_inst_pe_1_3_6_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_3_6_U32 ( .A1(npu_inst_n56), .A2(
        npu_inst_int_data_y_4__6__1_), .B1(npu_inst_pe_1_3_6_n3), .B2(
        npu_inst_int_data_x_3__7__1_), .ZN(npu_inst_pe_1_3_6_n63) );
  AOI22_X1 npu_inst_pe_1_3_6_U31 ( .A1(npu_inst_n56), .A2(
        npu_inst_int_data_y_4__6__0_), .B1(npu_inst_pe_1_3_6_n3), .B2(
        npu_inst_int_data_x_3__7__0_), .ZN(npu_inst_pe_1_3_6_n61) );
  INV_X1 npu_inst_pe_1_3_6_U30 ( .A(npu_inst_pe_1_3_6_int_data_0_), .ZN(
        npu_inst_pe_1_3_6_n13) );
  INV_X1 npu_inst_pe_1_3_6_U29 ( .A(npu_inst_n69), .ZN(npu_inst_pe_1_3_6_n5)
         );
  OR3_X1 npu_inst_pe_1_3_6_U28 ( .A1(npu_inst_pe_1_3_6_n6), .A2(
        npu_inst_pe_1_3_6_n8), .A3(npu_inst_pe_1_3_6_n5), .ZN(
        npu_inst_pe_1_3_6_n56) );
  OR3_X1 npu_inst_pe_1_3_6_U27 ( .A1(npu_inst_pe_1_3_6_n5), .A2(
        npu_inst_pe_1_3_6_n8), .A3(npu_inst_pe_1_3_6_n7), .ZN(
        npu_inst_pe_1_3_6_n48) );
  INV_X1 npu_inst_pe_1_3_6_U26 ( .A(npu_inst_pe_1_3_6_n5), .ZN(
        npu_inst_pe_1_3_6_n4) );
  INV_X1 npu_inst_pe_1_3_6_U25 ( .A(npu_inst_n124), .ZN(npu_inst_pe_1_3_6_n12)
         );
  OR3_X1 npu_inst_pe_1_3_6_U24 ( .A1(npu_inst_pe_1_3_6_n4), .A2(
        npu_inst_pe_1_3_6_n8), .A3(npu_inst_pe_1_3_6_n7), .ZN(
        npu_inst_pe_1_3_6_n52) );
  OR3_X1 npu_inst_pe_1_3_6_U23 ( .A1(npu_inst_pe_1_3_6_n6), .A2(
        npu_inst_pe_1_3_6_n8), .A3(npu_inst_pe_1_3_6_n4), .ZN(
        npu_inst_pe_1_3_6_n60) );
  NOR2_X1 npu_inst_pe_1_3_6_U22 ( .A1(npu_inst_pe_1_3_6_n60), .A2(
        npu_inst_pe_1_3_6_n3), .ZN(npu_inst_pe_1_3_6_n58) );
  NOR2_X1 npu_inst_pe_1_3_6_U21 ( .A1(npu_inst_pe_1_3_6_n56), .A2(
        npu_inst_pe_1_3_6_n3), .ZN(npu_inst_pe_1_3_6_n54) );
  NOR2_X1 npu_inst_pe_1_3_6_U20 ( .A1(npu_inst_pe_1_3_6_n52), .A2(
        npu_inst_pe_1_3_6_n3), .ZN(npu_inst_pe_1_3_6_n50) );
  NOR2_X1 npu_inst_pe_1_3_6_U19 ( .A1(npu_inst_pe_1_3_6_n48), .A2(
        npu_inst_pe_1_3_6_n3), .ZN(npu_inst_pe_1_3_6_n46) );
  NOR2_X1 npu_inst_pe_1_3_6_U18 ( .A1(npu_inst_pe_1_3_6_n40), .A2(
        npu_inst_pe_1_3_6_n3), .ZN(npu_inst_pe_1_3_6_n38) );
  NOR2_X1 npu_inst_pe_1_3_6_U17 ( .A1(npu_inst_pe_1_3_6_n44), .A2(
        npu_inst_pe_1_3_6_n3), .ZN(npu_inst_pe_1_3_6_n42) );
  BUF_X1 npu_inst_pe_1_3_6_U16 ( .A(npu_inst_n100), .Z(npu_inst_pe_1_3_6_n8)
         );
  BUF_X1 npu_inst_pe_1_3_6_U15 ( .A(npu_inst_pe_1_3_6_n12), .Z(
        npu_inst_pe_1_3_6_n11) );
  BUF_X1 npu_inst_pe_1_3_6_U14 ( .A(npu_inst_pe_1_3_6_n12), .Z(
        npu_inst_pe_1_3_6_n10) );
  BUF_X1 npu_inst_pe_1_3_6_U13 ( .A(npu_inst_pe_1_3_6_n12), .Z(
        npu_inst_pe_1_3_6_n9) );
  INV_X1 npu_inst_pe_1_3_6_U12 ( .A(npu_inst_pe_1_3_6_n38), .ZN(
        npu_inst_pe_1_3_6_n118) );
  INV_X1 npu_inst_pe_1_3_6_U11 ( .A(npu_inst_pe_1_3_6_n58), .ZN(
        npu_inst_pe_1_3_6_n114) );
  INV_X1 npu_inst_pe_1_3_6_U10 ( .A(npu_inst_pe_1_3_6_n54), .ZN(
        npu_inst_pe_1_3_6_n115) );
  INV_X1 npu_inst_pe_1_3_6_U9 ( .A(npu_inst_pe_1_3_6_n50), .ZN(
        npu_inst_pe_1_3_6_n116) );
  INV_X1 npu_inst_pe_1_3_6_U8 ( .A(npu_inst_pe_1_3_6_n46), .ZN(
        npu_inst_pe_1_3_6_n117) );
  INV_X1 npu_inst_pe_1_3_6_U7 ( .A(npu_inst_pe_1_3_6_n42), .ZN(
        npu_inst_pe_1_3_6_n119) );
  BUF_X1 npu_inst_pe_1_3_6_U6 ( .A(npu_inst_n23), .Z(npu_inst_pe_1_3_6_n2) );
  BUF_X1 npu_inst_pe_1_3_6_U5 ( .A(npu_inst_n23), .Z(npu_inst_pe_1_3_6_n1) );
  NOR2_X1 npu_inst_pe_1_3_6_U4 ( .A1(npu_inst_pe_1_3_6_int_q_weight_0_), .A2(
        npu_inst_pe_1_3_6_n1), .ZN(npu_inst_pe_1_3_6_n76) );
  NOR2_X1 npu_inst_pe_1_3_6_U3 ( .A1(npu_inst_pe_1_3_6_n27), .A2(
        npu_inst_pe_1_3_6_n1), .ZN(npu_inst_pe_1_3_6_n77) );
  FA_X1 npu_inst_pe_1_3_6_sub_77_U2_1 ( .A(npu_inst_pe_1_3_6_int_q_acc_1_), 
        .B(npu_inst_pe_1_3_6_n14), .CI(npu_inst_pe_1_3_6_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_3_6_sub_77_carry_2_), .S(npu_inst_pe_1_3_6_N66) );
  FA_X1 npu_inst_pe_1_3_6_add_79_U1_1 ( .A(npu_inst_pe_1_3_6_int_q_acc_1_), 
        .B(npu_inst_pe_1_3_6_int_data_1_), .CI(
        npu_inst_pe_1_3_6_add_79_carry_1_), .CO(
        npu_inst_pe_1_3_6_add_79_carry_2_), .S(npu_inst_pe_1_3_6_N74) );
  NAND3_X1 npu_inst_pe_1_3_6_U109 ( .A1(npu_inst_pe_1_3_6_n5), .A2(
        npu_inst_pe_1_3_6_n7), .A3(npu_inst_pe_1_3_6_n8), .ZN(
        npu_inst_pe_1_3_6_n44) );
  NAND3_X1 npu_inst_pe_1_3_6_U108 ( .A1(npu_inst_pe_1_3_6_n4), .A2(
        npu_inst_pe_1_3_6_n7), .A3(npu_inst_pe_1_3_6_n8), .ZN(
        npu_inst_pe_1_3_6_n40) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_3_6_n34), .CK(
        npu_inst_pe_1_3_6_net3603), .RN(npu_inst_pe_1_3_6_n9), .Q(
        npu_inst_pe_1_3_6_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_3_6_n35), .CK(
        npu_inst_pe_1_3_6_net3603), .RN(npu_inst_pe_1_3_6_n9), .Q(
        npu_inst_pe_1_3_6_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_3_6_n36), .CK(
        npu_inst_pe_1_3_6_net3603), .RN(npu_inst_pe_1_3_6_n9), .Q(
        npu_inst_pe_1_3_6_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_3_6_n98), .CK(
        npu_inst_pe_1_3_6_net3603), .RN(npu_inst_pe_1_3_6_n9), .Q(
        npu_inst_pe_1_3_6_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_3_6_n99), .CK(
        npu_inst_pe_1_3_6_net3603), .RN(npu_inst_pe_1_3_6_n9), .Q(
        npu_inst_pe_1_3_6_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_3_6_n100), 
        .CK(npu_inst_pe_1_3_6_net3603), .RN(npu_inst_pe_1_3_6_n9), .Q(
        npu_inst_pe_1_3_6_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_3_6_n33), .CK(
        npu_inst_pe_1_3_6_net3603), .RN(npu_inst_pe_1_3_6_n9), .Q(
        npu_inst_pe_1_3_6_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_3_6_n101), 
        .CK(npu_inst_pe_1_3_6_net3603), .RN(npu_inst_pe_1_3_6_n9), .Q(
        npu_inst_pe_1_3_6_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_weight_reg_0_ ( .D(npu_inst_n110), .CK(
        npu_inst_pe_1_3_6_net3609), .RN(npu_inst_pe_1_3_6_n9), .Q(
        npu_inst_pe_1_3_6_int_q_weight_0_), .QN(npu_inst_pe_1_3_6_n27) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_weight_reg_1_ ( .D(npu_inst_n116), .CK(
        npu_inst_pe_1_3_6_net3609), .RN(npu_inst_pe_1_3_6_n9), .Q(
        npu_inst_pe_1_3_6_int_q_weight_1_), .QN(npu_inst_pe_1_3_6_n26) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_3_6_n113), 
        .CK(npu_inst_pe_1_3_6_net3609), .RN(npu_inst_pe_1_3_6_n9), .Q(
        npu_inst_pe_1_3_6_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_3_6_n107), 
        .CK(npu_inst_pe_1_3_6_net3609), .RN(npu_inst_pe_1_3_6_n9), .Q(
        npu_inst_pe_1_3_6_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_3_6_n112), 
        .CK(npu_inst_pe_1_3_6_net3609), .RN(npu_inst_pe_1_3_6_n10), .Q(
        npu_inst_pe_1_3_6_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_3_6_n106), 
        .CK(npu_inst_pe_1_3_6_net3609), .RN(npu_inst_pe_1_3_6_n10), .Q(
        npu_inst_pe_1_3_6_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_3_6_n111), 
        .CK(npu_inst_pe_1_3_6_net3609), .RN(npu_inst_pe_1_3_6_n10), .Q(
        npu_inst_pe_1_3_6_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_3_6_n105), 
        .CK(npu_inst_pe_1_3_6_net3609), .RN(npu_inst_pe_1_3_6_n10), .Q(
        npu_inst_pe_1_3_6_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_3_6_n110), 
        .CK(npu_inst_pe_1_3_6_net3609), .RN(npu_inst_pe_1_3_6_n10), .Q(
        npu_inst_pe_1_3_6_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_3_6_n104), 
        .CK(npu_inst_pe_1_3_6_net3609), .RN(npu_inst_pe_1_3_6_n10), .Q(
        npu_inst_pe_1_3_6_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_3_6_n109), 
        .CK(npu_inst_pe_1_3_6_net3609), .RN(npu_inst_pe_1_3_6_n10), .Q(
        npu_inst_pe_1_3_6_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_3_6_n103), 
        .CK(npu_inst_pe_1_3_6_net3609), .RN(npu_inst_pe_1_3_6_n10), .Q(
        npu_inst_pe_1_3_6_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_3_6_n108), 
        .CK(npu_inst_pe_1_3_6_net3609), .RN(npu_inst_pe_1_3_6_n10), .Q(
        npu_inst_pe_1_3_6_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_3_6_n102), 
        .CK(npu_inst_pe_1_3_6_net3609), .RN(npu_inst_pe_1_3_6_n10), .Q(
        npu_inst_pe_1_3_6_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_3_6_n86), 
        .CK(npu_inst_pe_1_3_6_net3609), .RN(npu_inst_pe_1_3_6_n10), .Q(
        npu_inst_pe_1_3_6_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_3_6_n87), 
        .CK(npu_inst_pe_1_3_6_net3609), .RN(npu_inst_pe_1_3_6_n10), .Q(
        npu_inst_pe_1_3_6_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_3_6_n88), 
        .CK(npu_inst_pe_1_3_6_net3609), .RN(npu_inst_pe_1_3_6_n11), .Q(
        npu_inst_pe_1_3_6_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_3_6_n89), 
        .CK(npu_inst_pe_1_3_6_net3609), .RN(npu_inst_pe_1_3_6_n11), .Q(
        npu_inst_pe_1_3_6_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_3_6_n90), 
        .CK(npu_inst_pe_1_3_6_net3609), .RN(npu_inst_pe_1_3_6_n11), .Q(
        npu_inst_pe_1_3_6_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_3_6_n91), 
        .CK(npu_inst_pe_1_3_6_net3609), .RN(npu_inst_pe_1_3_6_n11), .Q(
        npu_inst_pe_1_3_6_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_3_6_n92), 
        .CK(npu_inst_pe_1_3_6_net3609), .RN(npu_inst_pe_1_3_6_n11), .Q(
        npu_inst_pe_1_3_6_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_3_6_n93), 
        .CK(npu_inst_pe_1_3_6_net3609), .RN(npu_inst_pe_1_3_6_n11), .Q(
        npu_inst_pe_1_3_6_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_3_6_n94), 
        .CK(npu_inst_pe_1_3_6_net3609), .RN(npu_inst_pe_1_3_6_n11), .Q(
        npu_inst_pe_1_3_6_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_3_6_n95), 
        .CK(npu_inst_pe_1_3_6_net3609), .RN(npu_inst_pe_1_3_6_n11), .Q(
        npu_inst_pe_1_3_6_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_3_6_n96), 
        .CK(npu_inst_pe_1_3_6_net3609), .RN(npu_inst_pe_1_3_6_n11), .Q(
        npu_inst_pe_1_3_6_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_3_6_n97), 
        .CK(npu_inst_pe_1_3_6_net3609), .RN(npu_inst_pe_1_3_6_n11), .Q(
        npu_inst_pe_1_3_6_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_3_6_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_3_6_N84), .SE(1'b0), .GCK(npu_inst_pe_1_3_6_net3603) );
  CLKGATETST_X1 npu_inst_pe_1_3_6_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n64), .SE(1'b0), .GCK(npu_inst_pe_1_3_6_net3609) );
  MUX2_X1 npu_inst_pe_1_3_7_U162 ( .A(npu_inst_pe_1_3_7_n32), .B(
        npu_inst_pe_1_3_7_n29), .S(npu_inst_pe_1_3_7_n8), .Z(
        npu_inst_pe_1_3_7_N93) );
  MUX2_X1 npu_inst_pe_1_3_7_U161 ( .A(npu_inst_pe_1_3_7_n31), .B(
        npu_inst_pe_1_3_7_n30), .S(npu_inst_pe_1_3_7_n6), .Z(
        npu_inst_pe_1_3_7_n32) );
  MUX2_X1 npu_inst_pe_1_3_7_U160 ( .A(npu_inst_pe_1_3_7_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_3_7_int_q_reg_v_1__0_), .S(npu_inst_pe_1_3_7_n4), .Z(
        npu_inst_pe_1_3_7_n31) );
  MUX2_X1 npu_inst_pe_1_3_7_U159 ( .A(npu_inst_pe_1_3_7_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_3_7_int_q_reg_v_3__0_), .S(npu_inst_pe_1_3_7_n4), .Z(
        npu_inst_pe_1_3_7_n30) );
  MUX2_X1 npu_inst_pe_1_3_7_U158 ( .A(npu_inst_pe_1_3_7_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_3_7_int_q_reg_v_5__0_), .S(npu_inst_pe_1_3_7_n4), .Z(
        npu_inst_pe_1_3_7_n29) );
  MUX2_X1 npu_inst_pe_1_3_7_U157 ( .A(npu_inst_pe_1_3_7_n28), .B(
        npu_inst_pe_1_3_7_n23), .S(npu_inst_pe_1_3_7_n8), .Z(
        npu_inst_pe_1_3_7_N94) );
  MUX2_X1 npu_inst_pe_1_3_7_U156 ( .A(npu_inst_pe_1_3_7_n25), .B(
        npu_inst_pe_1_3_7_n24), .S(npu_inst_pe_1_3_7_n6), .Z(
        npu_inst_pe_1_3_7_n28) );
  MUX2_X1 npu_inst_pe_1_3_7_U155 ( .A(npu_inst_pe_1_3_7_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_3_7_int_q_reg_v_1__1_), .S(npu_inst_pe_1_3_7_n4), .Z(
        npu_inst_pe_1_3_7_n25) );
  MUX2_X1 npu_inst_pe_1_3_7_U154 ( .A(npu_inst_pe_1_3_7_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_3_7_int_q_reg_v_3__1_), .S(npu_inst_pe_1_3_7_n4), .Z(
        npu_inst_pe_1_3_7_n24) );
  MUX2_X1 npu_inst_pe_1_3_7_U153 ( .A(npu_inst_pe_1_3_7_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_3_7_int_q_reg_v_5__1_), .S(npu_inst_pe_1_3_7_n4), .Z(
        npu_inst_pe_1_3_7_n23) );
  MUX2_X1 npu_inst_pe_1_3_7_U152 ( .A(npu_inst_pe_1_3_7_n22), .B(
        npu_inst_pe_1_3_7_n19), .S(npu_inst_pe_1_3_7_n8), .Z(
        npu_inst_int_data_x_3__7__1_) );
  MUX2_X1 npu_inst_pe_1_3_7_U151 ( .A(npu_inst_pe_1_3_7_n21), .B(
        npu_inst_pe_1_3_7_n20), .S(npu_inst_pe_1_3_7_n6), .Z(
        npu_inst_pe_1_3_7_n22) );
  MUX2_X1 npu_inst_pe_1_3_7_U150 ( .A(npu_inst_pe_1_3_7_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_3_7_int_q_reg_h_1__1_), .S(npu_inst_pe_1_3_7_n4), .Z(
        npu_inst_pe_1_3_7_n21) );
  MUX2_X1 npu_inst_pe_1_3_7_U149 ( .A(npu_inst_pe_1_3_7_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_3_7_int_q_reg_h_3__1_), .S(npu_inst_pe_1_3_7_n4), .Z(
        npu_inst_pe_1_3_7_n20) );
  MUX2_X1 npu_inst_pe_1_3_7_U148 ( .A(npu_inst_pe_1_3_7_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_3_7_int_q_reg_h_5__1_), .S(npu_inst_pe_1_3_7_n4), .Z(
        npu_inst_pe_1_3_7_n19) );
  MUX2_X1 npu_inst_pe_1_3_7_U147 ( .A(npu_inst_pe_1_3_7_n18), .B(
        npu_inst_pe_1_3_7_n15), .S(npu_inst_pe_1_3_7_n8), .Z(
        npu_inst_int_data_x_3__7__0_) );
  MUX2_X1 npu_inst_pe_1_3_7_U146 ( .A(npu_inst_pe_1_3_7_n17), .B(
        npu_inst_pe_1_3_7_n16), .S(npu_inst_pe_1_3_7_n6), .Z(
        npu_inst_pe_1_3_7_n18) );
  MUX2_X1 npu_inst_pe_1_3_7_U145 ( .A(npu_inst_pe_1_3_7_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_3_7_int_q_reg_h_1__0_), .S(npu_inst_pe_1_3_7_n4), .Z(
        npu_inst_pe_1_3_7_n17) );
  MUX2_X1 npu_inst_pe_1_3_7_U144 ( .A(npu_inst_pe_1_3_7_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_3_7_int_q_reg_h_3__0_), .S(npu_inst_pe_1_3_7_n4), .Z(
        npu_inst_pe_1_3_7_n16) );
  MUX2_X1 npu_inst_pe_1_3_7_U143 ( .A(npu_inst_pe_1_3_7_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_3_7_int_q_reg_h_5__0_), .S(npu_inst_pe_1_3_7_n4), .Z(
        npu_inst_pe_1_3_7_n15) );
  XOR2_X1 npu_inst_pe_1_3_7_U142 ( .A(npu_inst_pe_1_3_7_int_data_0_), .B(
        npu_inst_pe_1_3_7_int_q_acc_0_), .Z(npu_inst_pe_1_3_7_N73) );
  AND2_X1 npu_inst_pe_1_3_7_U141 ( .A1(npu_inst_pe_1_3_7_int_q_acc_0_), .A2(
        npu_inst_pe_1_3_7_int_data_0_), .ZN(npu_inst_pe_1_3_7_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_3_7_U140 ( .A(npu_inst_pe_1_3_7_int_q_acc_0_), .B(
        npu_inst_pe_1_3_7_n13), .ZN(npu_inst_pe_1_3_7_N65) );
  OR2_X1 npu_inst_pe_1_3_7_U139 ( .A1(npu_inst_pe_1_3_7_n13), .A2(
        npu_inst_pe_1_3_7_int_q_acc_0_), .ZN(npu_inst_pe_1_3_7_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_3_7_U138 ( .A(npu_inst_pe_1_3_7_int_q_acc_2_), .B(
        npu_inst_pe_1_3_7_add_79_carry_2_), .Z(npu_inst_pe_1_3_7_N75) );
  AND2_X1 npu_inst_pe_1_3_7_U137 ( .A1(npu_inst_pe_1_3_7_add_79_carry_2_), 
        .A2(npu_inst_pe_1_3_7_int_q_acc_2_), .ZN(
        npu_inst_pe_1_3_7_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_3_7_U136 ( .A(npu_inst_pe_1_3_7_int_q_acc_3_), .B(
        npu_inst_pe_1_3_7_add_79_carry_3_), .Z(npu_inst_pe_1_3_7_N76) );
  AND2_X1 npu_inst_pe_1_3_7_U135 ( .A1(npu_inst_pe_1_3_7_add_79_carry_3_), 
        .A2(npu_inst_pe_1_3_7_int_q_acc_3_), .ZN(
        npu_inst_pe_1_3_7_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_3_7_U134 ( .A(npu_inst_pe_1_3_7_int_q_acc_4_), .B(
        npu_inst_pe_1_3_7_add_79_carry_4_), .Z(npu_inst_pe_1_3_7_N77) );
  AND2_X1 npu_inst_pe_1_3_7_U133 ( .A1(npu_inst_pe_1_3_7_add_79_carry_4_), 
        .A2(npu_inst_pe_1_3_7_int_q_acc_4_), .ZN(
        npu_inst_pe_1_3_7_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_3_7_U132 ( .A(npu_inst_pe_1_3_7_int_q_acc_5_), .B(
        npu_inst_pe_1_3_7_add_79_carry_5_), .Z(npu_inst_pe_1_3_7_N78) );
  AND2_X1 npu_inst_pe_1_3_7_U131 ( .A1(npu_inst_pe_1_3_7_add_79_carry_5_), 
        .A2(npu_inst_pe_1_3_7_int_q_acc_5_), .ZN(
        npu_inst_pe_1_3_7_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_3_7_U130 ( .A(npu_inst_pe_1_3_7_int_q_acc_6_), .B(
        npu_inst_pe_1_3_7_add_79_carry_6_), .Z(npu_inst_pe_1_3_7_N79) );
  AND2_X1 npu_inst_pe_1_3_7_U129 ( .A1(npu_inst_pe_1_3_7_add_79_carry_6_), 
        .A2(npu_inst_pe_1_3_7_int_q_acc_6_), .ZN(
        npu_inst_pe_1_3_7_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_3_7_U128 ( .A(npu_inst_pe_1_3_7_int_q_acc_7_), .B(
        npu_inst_pe_1_3_7_add_79_carry_7_), .Z(npu_inst_pe_1_3_7_N80) );
  XNOR2_X1 npu_inst_pe_1_3_7_U127 ( .A(npu_inst_pe_1_3_7_sub_77_carry_2_), .B(
        npu_inst_pe_1_3_7_int_q_acc_2_), .ZN(npu_inst_pe_1_3_7_N67) );
  OR2_X1 npu_inst_pe_1_3_7_U126 ( .A1(npu_inst_pe_1_3_7_int_q_acc_2_), .A2(
        npu_inst_pe_1_3_7_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_3_7_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_3_7_U125 ( .A(npu_inst_pe_1_3_7_sub_77_carry_3_), .B(
        npu_inst_pe_1_3_7_int_q_acc_3_), .ZN(npu_inst_pe_1_3_7_N68) );
  OR2_X1 npu_inst_pe_1_3_7_U124 ( .A1(npu_inst_pe_1_3_7_int_q_acc_3_), .A2(
        npu_inst_pe_1_3_7_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_3_7_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_3_7_U123 ( .A(npu_inst_pe_1_3_7_sub_77_carry_4_), .B(
        npu_inst_pe_1_3_7_int_q_acc_4_), .ZN(npu_inst_pe_1_3_7_N69) );
  OR2_X1 npu_inst_pe_1_3_7_U122 ( .A1(npu_inst_pe_1_3_7_int_q_acc_4_), .A2(
        npu_inst_pe_1_3_7_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_3_7_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_3_7_U121 ( .A(npu_inst_pe_1_3_7_sub_77_carry_5_), .B(
        npu_inst_pe_1_3_7_int_q_acc_5_), .ZN(npu_inst_pe_1_3_7_N70) );
  OR2_X1 npu_inst_pe_1_3_7_U120 ( .A1(npu_inst_pe_1_3_7_int_q_acc_5_), .A2(
        npu_inst_pe_1_3_7_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_3_7_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_3_7_U119 ( .A(npu_inst_pe_1_3_7_sub_77_carry_6_), .B(
        npu_inst_pe_1_3_7_int_q_acc_6_), .ZN(npu_inst_pe_1_3_7_N71) );
  OR2_X1 npu_inst_pe_1_3_7_U118 ( .A1(npu_inst_pe_1_3_7_int_q_acc_6_), .A2(
        npu_inst_pe_1_3_7_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_3_7_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_3_7_U117 ( .A(npu_inst_pe_1_3_7_int_q_acc_7_), .B(
        npu_inst_pe_1_3_7_sub_77_carry_7_), .ZN(npu_inst_pe_1_3_7_N72) );
  INV_X1 npu_inst_pe_1_3_7_U116 ( .A(npu_inst_n77), .ZN(npu_inst_pe_1_3_7_n7)
         );
  INV_X1 npu_inst_pe_1_3_7_U115 ( .A(npu_inst_pe_1_3_7_n7), .ZN(
        npu_inst_pe_1_3_7_n6) );
  INV_X1 npu_inst_pe_1_3_7_U114 ( .A(npu_inst_n56), .ZN(npu_inst_pe_1_3_7_n3)
         );
  AOI22_X1 npu_inst_pe_1_3_7_U113 ( .A1(npu_inst_int_data_y_4__7__0_), .A2(
        npu_inst_pe_1_3_7_n58), .B1(npu_inst_pe_1_3_7_n114), .B2(
        npu_inst_pe_1_3_7_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_3_7_n57) );
  INV_X1 npu_inst_pe_1_3_7_U112 ( .A(npu_inst_pe_1_3_7_n57), .ZN(
        npu_inst_pe_1_3_7_n108) );
  AOI22_X1 npu_inst_pe_1_3_7_U111 ( .A1(npu_inst_int_data_y_4__7__0_), .A2(
        npu_inst_pe_1_3_7_n54), .B1(npu_inst_pe_1_3_7_n115), .B2(
        npu_inst_pe_1_3_7_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_3_7_n53) );
  INV_X1 npu_inst_pe_1_3_7_U110 ( .A(npu_inst_pe_1_3_7_n53), .ZN(
        npu_inst_pe_1_3_7_n109) );
  AOI22_X1 npu_inst_pe_1_3_7_U107 ( .A1(npu_inst_int_data_y_4__7__0_), .A2(
        npu_inst_pe_1_3_7_n50), .B1(npu_inst_pe_1_3_7_n116), .B2(
        npu_inst_pe_1_3_7_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_3_7_n49) );
  INV_X1 npu_inst_pe_1_3_7_U106 ( .A(npu_inst_pe_1_3_7_n49), .ZN(
        npu_inst_pe_1_3_7_n110) );
  AOI22_X1 npu_inst_pe_1_3_7_U105 ( .A1(npu_inst_int_data_y_4__7__0_), .A2(
        npu_inst_pe_1_3_7_n46), .B1(npu_inst_pe_1_3_7_n117), .B2(
        npu_inst_pe_1_3_7_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_3_7_n45) );
  INV_X1 npu_inst_pe_1_3_7_U104 ( .A(npu_inst_pe_1_3_7_n45), .ZN(
        npu_inst_pe_1_3_7_n111) );
  AOI22_X1 npu_inst_pe_1_3_7_U103 ( .A1(npu_inst_int_data_y_4__7__0_), .A2(
        npu_inst_pe_1_3_7_n42), .B1(npu_inst_pe_1_3_7_n119), .B2(
        npu_inst_pe_1_3_7_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_3_7_n41) );
  INV_X1 npu_inst_pe_1_3_7_U102 ( .A(npu_inst_pe_1_3_7_n41), .ZN(
        npu_inst_pe_1_3_7_n112) );
  AOI22_X1 npu_inst_pe_1_3_7_U101 ( .A1(npu_inst_int_data_y_4__7__1_), .A2(
        npu_inst_pe_1_3_7_n58), .B1(npu_inst_pe_1_3_7_n114), .B2(
        npu_inst_pe_1_3_7_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_3_7_n59) );
  INV_X1 npu_inst_pe_1_3_7_U100 ( .A(npu_inst_pe_1_3_7_n59), .ZN(
        npu_inst_pe_1_3_7_n102) );
  AOI22_X1 npu_inst_pe_1_3_7_U99 ( .A1(npu_inst_int_data_y_4__7__1_), .A2(
        npu_inst_pe_1_3_7_n54), .B1(npu_inst_pe_1_3_7_n115), .B2(
        npu_inst_pe_1_3_7_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_3_7_n55) );
  INV_X1 npu_inst_pe_1_3_7_U98 ( .A(npu_inst_pe_1_3_7_n55), .ZN(
        npu_inst_pe_1_3_7_n103) );
  AOI22_X1 npu_inst_pe_1_3_7_U97 ( .A1(npu_inst_int_data_y_4__7__1_), .A2(
        npu_inst_pe_1_3_7_n50), .B1(npu_inst_pe_1_3_7_n116), .B2(
        npu_inst_pe_1_3_7_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_3_7_n51) );
  INV_X1 npu_inst_pe_1_3_7_U96 ( .A(npu_inst_pe_1_3_7_n51), .ZN(
        npu_inst_pe_1_3_7_n104) );
  AOI22_X1 npu_inst_pe_1_3_7_U95 ( .A1(npu_inst_int_data_y_4__7__1_), .A2(
        npu_inst_pe_1_3_7_n46), .B1(npu_inst_pe_1_3_7_n117), .B2(
        npu_inst_pe_1_3_7_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_3_7_n47) );
  INV_X1 npu_inst_pe_1_3_7_U94 ( .A(npu_inst_pe_1_3_7_n47), .ZN(
        npu_inst_pe_1_3_7_n105) );
  AOI22_X1 npu_inst_pe_1_3_7_U93 ( .A1(npu_inst_int_data_y_4__7__1_), .A2(
        npu_inst_pe_1_3_7_n42), .B1(npu_inst_pe_1_3_7_n119), .B2(
        npu_inst_pe_1_3_7_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_3_7_n43) );
  INV_X1 npu_inst_pe_1_3_7_U92 ( .A(npu_inst_pe_1_3_7_n43), .ZN(
        npu_inst_pe_1_3_7_n106) );
  AOI22_X1 npu_inst_pe_1_3_7_U91 ( .A1(npu_inst_pe_1_3_7_n38), .A2(
        npu_inst_int_data_y_4__7__1_), .B1(npu_inst_pe_1_3_7_n118), .B2(
        npu_inst_pe_1_3_7_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_3_7_n39) );
  INV_X1 npu_inst_pe_1_3_7_U90 ( .A(npu_inst_pe_1_3_7_n39), .ZN(
        npu_inst_pe_1_3_7_n107) );
  AOI22_X1 npu_inst_pe_1_3_7_U89 ( .A1(npu_inst_pe_1_3_7_n38), .A2(
        npu_inst_int_data_y_4__7__0_), .B1(npu_inst_pe_1_3_7_n118), .B2(
        npu_inst_pe_1_3_7_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_3_7_n37) );
  INV_X1 npu_inst_pe_1_3_7_U88 ( .A(npu_inst_pe_1_3_7_n37), .ZN(
        npu_inst_pe_1_3_7_n113) );
  AND2_X1 npu_inst_pe_1_3_7_U87 ( .A1(npu_inst_pe_1_3_7_N93), .A2(npu_inst_n56), .ZN(npu_inst_int_data_y_3__7__0_) );
  AND2_X1 npu_inst_pe_1_3_7_U86 ( .A1(npu_inst_n56), .A2(npu_inst_pe_1_3_7_N94), .ZN(npu_inst_int_data_y_3__7__1_) );
  NOR3_X1 npu_inst_pe_1_3_7_U85 ( .A1(npu_inst_pe_1_3_7_n26), .A2(npu_inst_n56), .A3(npu_inst_int_ckg[32]), .ZN(npu_inst_pe_1_3_7_n85) );
  OR2_X1 npu_inst_pe_1_3_7_U84 ( .A1(npu_inst_pe_1_3_7_n85), .A2(
        npu_inst_pe_1_3_7_n2), .ZN(npu_inst_pe_1_3_7_N84) );
  AND2_X1 npu_inst_pe_1_3_7_U83 ( .A1(npu_inst_pe_1_3_7_int_q_acc_0_), .A2(
        npu_inst_pe_1_3_7_n1), .ZN(npu_inst_int_data_res_3__7__0_) );
  AND2_X1 npu_inst_pe_1_3_7_U82 ( .A1(npu_inst_pe_1_3_7_n2), .A2(
        npu_inst_pe_1_3_7_int_q_acc_7_), .ZN(npu_inst_int_data_res_3__7__7_)
         );
  AND2_X1 npu_inst_pe_1_3_7_U81 ( .A1(npu_inst_pe_1_3_7_int_q_acc_1_), .A2(
        npu_inst_pe_1_3_7_n1), .ZN(npu_inst_int_data_res_3__7__1_) );
  AND2_X1 npu_inst_pe_1_3_7_U80 ( .A1(npu_inst_pe_1_3_7_int_q_acc_2_), .A2(
        npu_inst_pe_1_3_7_n1), .ZN(npu_inst_int_data_res_3__7__2_) );
  AND2_X1 npu_inst_pe_1_3_7_U79 ( .A1(npu_inst_pe_1_3_7_int_q_acc_3_), .A2(
        npu_inst_pe_1_3_7_n2), .ZN(npu_inst_int_data_res_3__7__3_) );
  AND2_X1 npu_inst_pe_1_3_7_U78 ( .A1(npu_inst_pe_1_3_7_int_q_acc_4_), .A2(
        npu_inst_pe_1_3_7_n2), .ZN(npu_inst_int_data_res_3__7__4_) );
  AND2_X1 npu_inst_pe_1_3_7_U77 ( .A1(npu_inst_pe_1_3_7_int_q_acc_5_), .A2(
        npu_inst_pe_1_3_7_n2), .ZN(npu_inst_int_data_res_3__7__5_) );
  AND2_X1 npu_inst_pe_1_3_7_U76 ( .A1(npu_inst_pe_1_3_7_int_q_acc_6_), .A2(
        npu_inst_pe_1_3_7_n2), .ZN(npu_inst_int_data_res_3__7__6_) );
  AOI222_X1 npu_inst_pe_1_3_7_U75 ( .A1(npu_inst_int_data_res_4__7__0_), .A2(
        npu_inst_pe_1_3_7_n1), .B1(npu_inst_pe_1_3_7_N73), .B2(
        npu_inst_pe_1_3_7_n76), .C1(npu_inst_pe_1_3_7_N65), .C2(
        npu_inst_pe_1_3_7_n77), .ZN(npu_inst_pe_1_3_7_n84) );
  INV_X1 npu_inst_pe_1_3_7_U74 ( .A(npu_inst_pe_1_3_7_n84), .ZN(
        npu_inst_pe_1_3_7_n101) );
  AOI222_X1 npu_inst_pe_1_3_7_U73 ( .A1(npu_inst_int_data_res_4__7__7_), .A2(
        npu_inst_pe_1_3_7_n1), .B1(npu_inst_pe_1_3_7_N80), .B2(
        npu_inst_pe_1_3_7_n76), .C1(npu_inst_pe_1_3_7_N72), .C2(
        npu_inst_pe_1_3_7_n77), .ZN(npu_inst_pe_1_3_7_n75) );
  INV_X1 npu_inst_pe_1_3_7_U72 ( .A(npu_inst_pe_1_3_7_n75), .ZN(
        npu_inst_pe_1_3_7_n33) );
  AOI222_X1 npu_inst_pe_1_3_7_U71 ( .A1(npu_inst_int_data_res_4__7__1_), .A2(
        npu_inst_pe_1_3_7_n1), .B1(npu_inst_pe_1_3_7_N74), .B2(
        npu_inst_pe_1_3_7_n76), .C1(npu_inst_pe_1_3_7_N66), .C2(
        npu_inst_pe_1_3_7_n77), .ZN(npu_inst_pe_1_3_7_n83) );
  INV_X1 npu_inst_pe_1_3_7_U70 ( .A(npu_inst_pe_1_3_7_n83), .ZN(
        npu_inst_pe_1_3_7_n100) );
  AOI222_X1 npu_inst_pe_1_3_7_U69 ( .A1(npu_inst_int_data_res_4__7__2_), .A2(
        npu_inst_pe_1_3_7_n1), .B1(npu_inst_pe_1_3_7_N75), .B2(
        npu_inst_pe_1_3_7_n76), .C1(npu_inst_pe_1_3_7_N67), .C2(
        npu_inst_pe_1_3_7_n77), .ZN(npu_inst_pe_1_3_7_n82) );
  INV_X1 npu_inst_pe_1_3_7_U68 ( .A(npu_inst_pe_1_3_7_n82), .ZN(
        npu_inst_pe_1_3_7_n99) );
  AOI222_X1 npu_inst_pe_1_3_7_U67 ( .A1(npu_inst_int_data_res_4__7__3_), .A2(
        npu_inst_pe_1_3_7_n1), .B1(npu_inst_pe_1_3_7_N76), .B2(
        npu_inst_pe_1_3_7_n76), .C1(npu_inst_pe_1_3_7_N68), .C2(
        npu_inst_pe_1_3_7_n77), .ZN(npu_inst_pe_1_3_7_n81) );
  INV_X1 npu_inst_pe_1_3_7_U66 ( .A(npu_inst_pe_1_3_7_n81), .ZN(
        npu_inst_pe_1_3_7_n98) );
  AOI222_X1 npu_inst_pe_1_3_7_U65 ( .A1(npu_inst_int_data_res_4__7__4_), .A2(
        npu_inst_pe_1_3_7_n1), .B1(npu_inst_pe_1_3_7_N77), .B2(
        npu_inst_pe_1_3_7_n76), .C1(npu_inst_pe_1_3_7_N69), .C2(
        npu_inst_pe_1_3_7_n77), .ZN(npu_inst_pe_1_3_7_n80) );
  INV_X1 npu_inst_pe_1_3_7_U64 ( .A(npu_inst_pe_1_3_7_n80), .ZN(
        npu_inst_pe_1_3_7_n36) );
  AOI222_X1 npu_inst_pe_1_3_7_U63 ( .A1(npu_inst_int_data_res_4__7__5_), .A2(
        npu_inst_pe_1_3_7_n1), .B1(npu_inst_pe_1_3_7_N78), .B2(
        npu_inst_pe_1_3_7_n76), .C1(npu_inst_pe_1_3_7_N70), .C2(
        npu_inst_pe_1_3_7_n77), .ZN(npu_inst_pe_1_3_7_n79) );
  INV_X1 npu_inst_pe_1_3_7_U62 ( .A(npu_inst_pe_1_3_7_n79), .ZN(
        npu_inst_pe_1_3_7_n35) );
  AOI222_X1 npu_inst_pe_1_3_7_U61 ( .A1(npu_inst_int_data_res_4__7__6_), .A2(
        npu_inst_pe_1_3_7_n1), .B1(npu_inst_pe_1_3_7_N79), .B2(
        npu_inst_pe_1_3_7_n76), .C1(npu_inst_pe_1_3_7_N71), .C2(
        npu_inst_pe_1_3_7_n77), .ZN(npu_inst_pe_1_3_7_n78) );
  INV_X1 npu_inst_pe_1_3_7_U60 ( .A(npu_inst_pe_1_3_7_n78), .ZN(
        npu_inst_pe_1_3_7_n34) );
  INV_X1 npu_inst_pe_1_3_7_U59 ( .A(npu_inst_pe_1_3_7_int_data_1_), .ZN(
        npu_inst_pe_1_3_7_n14) );
  AND2_X1 npu_inst_pe_1_3_7_U58 ( .A1(npu_inst_int_data_x_3__7__1_), .A2(
        npu_inst_pe_1_3_7_int_q_weight_1_), .ZN(npu_inst_pe_1_3_7_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_3_7_U57 ( .A1(npu_inst_int_data_x_3__7__0_), .A2(
        npu_inst_pe_1_3_7_int_q_weight_1_), .ZN(npu_inst_pe_1_3_7_int_data_0_)
         );
  NAND2_X1 npu_inst_pe_1_3_7_U56 ( .A1(npu_inst_pe_1_3_7_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_3_7_n60), .ZN(npu_inst_pe_1_3_7_n74) );
  OAI21_X1 npu_inst_pe_1_3_7_U55 ( .B1(npu_inst_pe_1_3_7_n63), .B2(
        npu_inst_pe_1_3_7_n60), .A(npu_inst_pe_1_3_7_n74), .ZN(
        npu_inst_pe_1_3_7_n97) );
  NAND2_X1 npu_inst_pe_1_3_7_U54 ( .A1(npu_inst_pe_1_3_7_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_3_7_n60), .ZN(npu_inst_pe_1_3_7_n73) );
  OAI21_X1 npu_inst_pe_1_3_7_U53 ( .B1(npu_inst_pe_1_3_7_n61), .B2(
        npu_inst_pe_1_3_7_n60), .A(npu_inst_pe_1_3_7_n73), .ZN(
        npu_inst_pe_1_3_7_n96) );
  NAND2_X1 npu_inst_pe_1_3_7_U52 ( .A1(npu_inst_pe_1_3_7_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_3_7_n56), .ZN(npu_inst_pe_1_3_7_n72) );
  OAI21_X1 npu_inst_pe_1_3_7_U51 ( .B1(npu_inst_pe_1_3_7_n63), .B2(
        npu_inst_pe_1_3_7_n56), .A(npu_inst_pe_1_3_7_n72), .ZN(
        npu_inst_pe_1_3_7_n95) );
  NAND2_X1 npu_inst_pe_1_3_7_U50 ( .A1(npu_inst_pe_1_3_7_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_3_7_n56), .ZN(npu_inst_pe_1_3_7_n71) );
  OAI21_X1 npu_inst_pe_1_3_7_U49 ( .B1(npu_inst_pe_1_3_7_n61), .B2(
        npu_inst_pe_1_3_7_n56), .A(npu_inst_pe_1_3_7_n71), .ZN(
        npu_inst_pe_1_3_7_n94) );
  NAND2_X1 npu_inst_pe_1_3_7_U48 ( .A1(npu_inst_pe_1_3_7_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_3_7_n52), .ZN(npu_inst_pe_1_3_7_n70) );
  OAI21_X1 npu_inst_pe_1_3_7_U47 ( .B1(npu_inst_pe_1_3_7_n63), .B2(
        npu_inst_pe_1_3_7_n52), .A(npu_inst_pe_1_3_7_n70), .ZN(
        npu_inst_pe_1_3_7_n93) );
  NAND2_X1 npu_inst_pe_1_3_7_U46 ( .A1(npu_inst_pe_1_3_7_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_3_7_n52), .ZN(npu_inst_pe_1_3_7_n69) );
  OAI21_X1 npu_inst_pe_1_3_7_U45 ( .B1(npu_inst_pe_1_3_7_n61), .B2(
        npu_inst_pe_1_3_7_n52), .A(npu_inst_pe_1_3_7_n69), .ZN(
        npu_inst_pe_1_3_7_n92) );
  NAND2_X1 npu_inst_pe_1_3_7_U44 ( .A1(npu_inst_pe_1_3_7_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_3_7_n48), .ZN(npu_inst_pe_1_3_7_n68) );
  OAI21_X1 npu_inst_pe_1_3_7_U43 ( .B1(npu_inst_pe_1_3_7_n63), .B2(
        npu_inst_pe_1_3_7_n48), .A(npu_inst_pe_1_3_7_n68), .ZN(
        npu_inst_pe_1_3_7_n91) );
  NAND2_X1 npu_inst_pe_1_3_7_U42 ( .A1(npu_inst_pe_1_3_7_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_3_7_n48), .ZN(npu_inst_pe_1_3_7_n67) );
  OAI21_X1 npu_inst_pe_1_3_7_U41 ( .B1(npu_inst_pe_1_3_7_n61), .B2(
        npu_inst_pe_1_3_7_n48), .A(npu_inst_pe_1_3_7_n67), .ZN(
        npu_inst_pe_1_3_7_n90) );
  NAND2_X1 npu_inst_pe_1_3_7_U40 ( .A1(npu_inst_pe_1_3_7_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_3_7_n44), .ZN(npu_inst_pe_1_3_7_n66) );
  OAI21_X1 npu_inst_pe_1_3_7_U39 ( .B1(npu_inst_pe_1_3_7_n63), .B2(
        npu_inst_pe_1_3_7_n44), .A(npu_inst_pe_1_3_7_n66), .ZN(
        npu_inst_pe_1_3_7_n89) );
  NAND2_X1 npu_inst_pe_1_3_7_U38 ( .A1(npu_inst_pe_1_3_7_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_3_7_n44), .ZN(npu_inst_pe_1_3_7_n65) );
  OAI21_X1 npu_inst_pe_1_3_7_U37 ( .B1(npu_inst_pe_1_3_7_n61), .B2(
        npu_inst_pe_1_3_7_n44), .A(npu_inst_pe_1_3_7_n65), .ZN(
        npu_inst_pe_1_3_7_n88) );
  NAND2_X1 npu_inst_pe_1_3_7_U36 ( .A1(npu_inst_pe_1_3_7_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_3_7_n40), .ZN(npu_inst_pe_1_3_7_n64) );
  OAI21_X1 npu_inst_pe_1_3_7_U35 ( .B1(npu_inst_pe_1_3_7_n63), .B2(
        npu_inst_pe_1_3_7_n40), .A(npu_inst_pe_1_3_7_n64), .ZN(
        npu_inst_pe_1_3_7_n87) );
  NAND2_X1 npu_inst_pe_1_3_7_U34 ( .A1(npu_inst_pe_1_3_7_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_3_7_n40), .ZN(npu_inst_pe_1_3_7_n62) );
  OAI21_X1 npu_inst_pe_1_3_7_U33 ( .B1(npu_inst_pe_1_3_7_n61), .B2(
        npu_inst_pe_1_3_7_n40), .A(npu_inst_pe_1_3_7_n62), .ZN(
        npu_inst_pe_1_3_7_n86) );
  INV_X1 npu_inst_pe_1_3_7_U32 ( .A(npu_inst_pe_1_3_7_int_data_0_), .ZN(
        npu_inst_pe_1_3_7_n13) );
  INV_X1 npu_inst_pe_1_3_7_U31 ( .A(npu_inst_n69), .ZN(npu_inst_pe_1_3_7_n5)
         );
  AOI22_X1 npu_inst_pe_1_3_7_U30 ( .A1(npu_inst_n56), .A2(
        npu_inst_int_data_y_4__7__1_), .B1(npu_inst_pe_1_3_7_n3), .B2(
        int_i_data_h_npu4[1]), .ZN(npu_inst_pe_1_3_7_n63) );
  AOI22_X1 npu_inst_pe_1_3_7_U29 ( .A1(npu_inst_n56), .A2(
        npu_inst_int_data_y_4__7__0_), .B1(npu_inst_pe_1_3_7_n3), .B2(
        int_i_data_h_npu4[0]), .ZN(npu_inst_pe_1_3_7_n61) );
  OR3_X1 npu_inst_pe_1_3_7_U28 ( .A1(npu_inst_pe_1_3_7_n6), .A2(
        npu_inst_pe_1_3_7_n8), .A3(npu_inst_pe_1_3_7_n5), .ZN(
        npu_inst_pe_1_3_7_n56) );
  OR3_X1 npu_inst_pe_1_3_7_U27 ( .A1(npu_inst_pe_1_3_7_n5), .A2(
        npu_inst_pe_1_3_7_n8), .A3(npu_inst_pe_1_3_7_n7), .ZN(
        npu_inst_pe_1_3_7_n48) );
  INV_X1 npu_inst_pe_1_3_7_U26 ( .A(npu_inst_pe_1_3_7_n5), .ZN(
        npu_inst_pe_1_3_7_n4) );
  INV_X1 npu_inst_pe_1_3_7_U25 ( .A(npu_inst_n124), .ZN(npu_inst_pe_1_3_7_n12)
         );
  OR3_X1 npu_inst_pe_1_3_7_U24 ( .A1(npu_inst_pe_1_3_7_n4), .A2(
        npu_inst_pe_1_3_7_n8), .A3(npu_inst_pe_1_3_7_n7), .ZN(
        npu_inst_pe_1_3_7_n52) );
  OR3_X1 npu_inst_pe_1_3_7_U23 ( .A1(npu_inst_pe_1_3_7_n6), .A2(
        npu_inst_pe_1_3_7_n8), .A3(npu_inst_pe_1_3_7_n4), .ZN(
        npu_inst_pe_1_3_7_n60) );
  NOR2_X1 npu_inst_pe_1_3_7_U22 ( .A1(npu_inst_pe_1_3_7_n60), .A2(
        npu_inst_pe_1_3_7_n3), .ZN(npu_inst_pe_1_3_7_n58) );
  NOR2_X1 npu_inst_pe_1_3_7_U21 ( .A1(npu_inst_pe_1_3_7_n56), .A2(
        npu_inst_pe_1_3_7_n3), .ZN(npu_inst_pe_1_3_7_n54) );
  NOR2_X1 npu_inst_pe_1_3_7_U20 ( .A1(npu_inst_pe_1_3_7_n52), .A2(
        npu_inst_pe_1_3_7_n3), .ZN(npu_inst_pe_1_3_7_n50) );
  NOR2_X1 npu_inst_pe_1_3_7_U19 ( .A1(npu_inst_pe_1_3_7_n48), .A2(
        npu_inst_pe_1_3_7_n3), .ZN(npu_inst_pe_1_3_7_n46) );
  NOR2_X1 npu_inst_pe_1_3_7_U18 ( .A1(npu_inst_pe_1_3_7_n40), .A2(
        npu_inst_pe_1_3_7_n3), .ZN(npu_inst_pe_1_3_7_n38) );
  NOR2_X1 npu_inst_pe_1_3_7_U17 ( .A1(npu_inst_pe_1_3_7_n44), .A2(
        npu_inst_pe_1_3_7_n3), .ZN(npu_inst_pe_1_3_7_n42) );
  BUF_X1 npu_inst_pe_1_3_7_U16 ( .A(npu_inst_n100), .Z(npu_inst_pe_1_3_7_n8)
         );
  BUF_X1 npu_inst_pe_1_3_7_U15 ( .A(npu_inst_pe_1_3_7_n12), .Z(
        npu_inst_pe_1_3_7_n11) );
  BUF_X1 npu_inst_pe_1_3_7_U14 ( .A(npu_inst_pe_1_3_7_n12), .Z(
        npu_inst_pe_1_3_7_n10) );
  BUF_X1 npu_inst_pe_1_3_7_U13 ( .A(npu_inst_pe_1_3_7_n12), .Z(
        npu_inst_pe_1_3_7_n9) );
  INV_X1 npu_inst_pe_1_3_7_U12 ( .A(npu_inst_pe_1_3_7_n38), .ZN(
        npu_inst_pe_1_3_7_n118) );
  INV_X1 npu_inst_pe_1_3_7_U11 ( .A(npu_inst_pe_1_3_7_n58), .ZN(
        npu_inst_pe_1_3_7_n114) );
  INV_X1 npu_inst_pe_1_3_7_U10 ( .A(npu_inst_pe_1_3_7_n54), .ZN(
        npu_inst_pe_1_3_7_n115) );
  INV_X1 npu_inst_pe_1_3_7_U9 ( .A(npu_inst_pe_1_3_7_n50), .ZN(
        npu_inst_pe_1_3_7_n116) );
  INV_X1 npu_inst_pe_1_3_7_U8 ( .A(npu_inst_pe_1_3_7_n46), .ZN(
        npu_inst_pe_1_3_7_n117) );
  INV_X1 npu_inst_pe_1_3_7_U7 ( .A(npu_inst_pe_1_3_7_n42), .ZN(
        npu_inst_pe_1_3_7_n119) );
  BUF_X1 npu_inst_pe_1_3_7_U6 ( .A(npu_inst_n23), .Z(npu_inst_pe_1_3_7_n2) );
  BUF_X1 npu_inst_pe_1_3_7_U5 ( .A(npu_inst_n23), .Z(npu_inst_pe_1_3_7_n1) );
  NOR2_X1 npu_inst_pe_1_3_7_U4 ( .A1(npu_inst_pe_1_3_7_int_q_weight_0_), .A2(
        npu_inst_pe_1_3_7_n1), .ZN(npu_inst_pe_1_3_7_n76) );
  NOR2_X1 npu_inst_pe_1_3_7_U3 ( .A1(npu_inst_pe_1_3_7_n27), .A2(
        npu_inst_pe_1_3_7_n1), .ZN(npu_inst_pe_1_3_7_n77) );
  FA_X1 npu_inst_pe_1_3_7_sub_77_U2_1 ( .A(npu_inst_pe_1_3_7_int_q_acc_1_), 
        .B(npu_inst_pe_1_3_7_n14), .CI(npu_inst_pe_1_3_7_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_3_7_sub_77_carry_2_), .S(npu_inst_pe_1_3_7_N66) );
  FA_X1 npu_inst_pe_1_3_7_add_79_U1_1 ( .A(npu_inst_pe_1_3_7_int_q_acc_1_), 
        .B(npu_inst_pe_1_3_7_int_data_1_), .CI(
        npu_inst_pe_1_3_7_add_79_carry_1_), .CO(
        npu_inst_pe_1_3_7_add_79_carry_2_), .S(npu_inst_pe_1_3_7_N74) );
  NAND3_X1 npu_inst_pe_1_3_7_U109 ( .A1(npu_inst_pe_1_3_7_n5), .A2(
        npu_inst_pe_1_3_7_n7), .A3(npu_inst_pe_1_3_7_n8), .ZN(
        npu_inst_pe_1_3_7_n44) );
  NAND3_X1 npu_inst_pe_1_3_7_U108 ( .A1(npu_inst_pe_1_3_7_n4), .A2(
        npu_inst_pe_1_3_7_n7), .A3(npu_inst_pe_1_3_7_n8), .ZN(
        npu_inst_pe_1_3_7_n40) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_3_7_n34), .CK(
        npu_inst_pe_1_3_7_net3580), .RN(npu_inst_pe_1_3_7_n9), .Q(
        npu_inst_pe_1_3_7_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_3_7_n35), .CK(
        npu_inst_pe_1_3_7_net3580), .RN(npu_inst_pe_1_3_7_n9), .Q(
        npu_inst_pe_1_3_7_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_3_7_n36), .CK(
        npu_inst_pe_1_3_7_net3580), .RN(npu_inst_pe_1_3_7_n9), .Q(
        npu_inst_pe_1_3_7_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_3_7_n98), .CK(
        npu_inst_pe_1_3_7_net3580), .RN(npu_inst_pe_1_3_7_n9), .Q(
        npu_inst_pe_1_3_7_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_3_7_n99), .CK(
        npu_inst_pe_1_3_7_net3580), .RN(npu_inst_pe_1_3_7_n9), .Q(
        npu_inst_pe_1_3_7_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_3_7_n100), 
        .CK(npu_inst_pe_1_3_7_net3580), .RN(npu_inst_pe_1_3_7_n9), .Q(
        npu_inst_pe_1_3_7_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_3_7_n33), .CK(
        npu_inst_pe_1_3_7_net3580), .RN(npu_inst_pe_1_3_7_n9), .Q(
        npu_inst_pe_1_3_7_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_3_7_n101), 
        .CK(npu_inst_pe_1_3_7_net3580), .RN(npu_inst_pe_1_3_7_n9), .Q(
        npu_inst_pe_1_3_7_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_weight_reg_0_ ( .D(npu_inst_n110), .CK(
        npu_inst_pe_1_3_7_net3586), .RN(npu_inst_pe_1_3_7_n9), .Q(
        npu_inst_pe_1_3_7_int_q_weight_0_), .QN(npu_inst_pe_1_3_7_n27) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_weight_reg_1_ ( .D(npu_inst_n116), .CK(
        npu_inst_pe_1_3_7_net3586), .RN(npu_inst_pe_1_3_7_n9), .Q(
        npu_inst_pe_1_3_7_int_q_weight_1_), .QN(npu_inst_pe_1_3_7_n26) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_3_7_n113), 
        .CK(npu_inst_pe_1_3_7_net3586), .RN(npu_inst_pe_1_3_7_n9), .Q(
        npu_inst_pe_1_3_7_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_3_7_n107), 
        .CK(npu_inst_pe_1_3_7_net3586), .RN(npu_inst_pe_1_3_7_n9), .Q(
        npu_inst_pe_1_3_7_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_3_7_n112), 
        .CK(npu_inst_pe_1_3_7_net3586), .RN(npu_inst_pe_1_3_7_n10), .Q(
        npu_inst_pe_1_3_7_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_3_7_n106), 
        .CK(npu_inst_pe_1_3_7_net3586), .RN(npu_inst_pe_1_3_7_n10), .Q(
        npu_inst_pe_1_3_7_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_3_7_n111), 
        .CK(npu_inst_pe_1_3_7_net3586), .RN(npu_inst_pe_1_3_7_n10), .Q(
        npu_inst_pe_1_3_7_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_3_7_n105), 
        .CK(npu_inst_pe_1_3_7_net3586), .RN(npu_inst_pe_1_3_7_n10), .Q(
        npu_inst_pe_1_3_7_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_3_7_n110), 
        .CK(npu_inst_pe_1_3_7_net3586), .RN(npu_inst_pe_1_3_7_n10), .Q(
        npu_inst_pe_1_3_7_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_3_7_n104), 
        .CK(npu_inst_pe_1_3_7_net3586), .RN(npu_inst_pe_1_3_7_n10), .Q(
        npu_inst_pe_1_3_7_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_3_7_n109), 
        .CK(npu_inst_pe_1_3_7_net3586), .RN(npu_inst_pe_1_3_7_n10), .Q(
        npu_inst_pe_1_3_7_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_3_7_n103), 
        .CK(npu_inst_pe_1_3_7_net3586), .RN(npu_inst_pe_1_3_7_n10), .Q(
        npu_inst_pe_1_3_7_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_3_7_n108), 
        .CK(npu_inst_pe_1_3_7_net3586), .RN(npu_inst_pe_1_3_7_n10), .Q(
        npu_inst_pe_1_3_7_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_3_7_n102), 
        .CK(npu_inst_pe_1_3_7_net3586), .RN(npu_inst_pe_1_3_7_n10), .Q(
        npu_inst_pe_1_3_7_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_3_7_n86), 
        .CK(npu_inst_pe_1_3_7_net3586), .RN(npu_inst_pe_1_3_7_n10), .Q(
        npu_inst_pe_1_3_7_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_3_7_n87), 
        .CK(npu_inst_pe_1_3_7_net3586), .RN(npu_inst_pe_1_3_7_n10), .Q(
        npu_inst_pe_1_3_7_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_3_7_n88), 
        .CK(npu_inst_pe_1_3_7_net3586), .RN(npu_inst_pe_1_3_7_n11), .Q(
        npu_inst_pe_1_3_7_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_3_7_n89), 
        .CK(npu_inst_pe_1_3_7_net3586), .RN(npu_inst_pe_1_3_7_n11), .Q(
        npu_inst_pe_1_3_7_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_3_7_n90), 
        .CK(npu_inst_pe_1_3_7_net3586), .RN(npu_inst_pe_1_3_7_n11), .Q(
        npu_inst_pe_1_3_7_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_3_7_n91), 
        .CK(npu_inst_pe_1_3_7_net3586), .RN(npu_inst_pe_1_3_7_n11), .Q(
        npu_inst_pe_1_3_7_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_3_7_n92), 
        .CK(npu_inst_pe_1_3_7_net3586), .RN(npu_inst_pe_1_3_7_n11), .Q(
        npu_inst_pe_1_3_7_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_3_7_n93), 
        .CK(npu_inst_pe_1_3_7_net3586), .RN(npu_inst_pe_1_3_7_n11), .Q(
        npu_inst_pe_1_3_7_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_3_7_n94), 
        .CK(npu_inst_pe_1_3_7_net3586), .RN(npu_inst_pe_1_3_7_n11), .Q(
        npu_inst_pe_1_3_7_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_3_7_n95), 
        .CK(npu_inst_pe_1_3_7_net3586), .RN(npu_inst_pe_1_3_7_n11), .Q(
        npu_inst_pe_1_3_7_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_3_7_n96), 
        .CK(npu_inst_pe_1_3_7_net3586), .RN(npu_inst_pe_1_3_7_n11), .Q(
        npu_inst_pe_1_3_7_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_3_7_n97), 
        .CK(npu_inst_pe_1_3_7_net3586), .RN(npu_inst_pe_1_3_7_n11), .Q(
        npu_inst_pe_1_3_7_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_3_7_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_3_7_N84), .SE(1'b0), .GCK(npu_inst_pe_1_3_7_net3580) );
  CLKGATETST_X1 npu_inst_pe_1_3_7_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n63), .SE(1'b0), .GCK(npu_inst_pe_1_3_7_net3586) );
  MUX2_X1 npu_inst_pe_1_4_0_U162 ( .A(npu_inst_pe_1_4_0_n32), .B(
        npu_inst_pe_1_4_0_n29), .S(npu_inst_pe_1_4_0_n8), .Z(
        npu_inst_pe_1_4_0_N93) );
  MUX2_X1 npu_inst_pe_1_4_0_U161 ( .A(npu_inst_pe_1_4_0_n31), .B(
        npu_inst_pe_1_4_0_n30), .S(npu_inst_pe_1_4_0_n6), .Z(
        npu_inst_pe_1_4_0_n32) );
  MUX2_X1 npu_inst_pe_1_4_0_U160 ( .A(npu_inst_pe_1_4_0_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_4_0_int_q_reg_v_1__0_), .S(npu_inst_pe_1_4_0_n4), .Z(
        npu_inst_pe_1_4_0_n31) );
  MUX2_X1 npu_inst_pe_1_4_0_U159 ( .A(npu_inst_pe_1_4_0_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_4_0_int_q_reg_v_3__0_), .S(npu_inst_pe_1_4_0_n4), .Z(
        npu_inst_pe_1_4_0_n30) );
  MUX2_X1 npu_inst_pe_1_4_0_U158 ( .A(npu_inst_pe_1_4_0_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_4_0_int_q_reg_v_5__0_), .S(npu_inst_pe_1_4_0_n4), .Z(
        npu_inst_pe_1_4_0_n29) );
  MUX2_X1 npu_inst_pe_1_4_0_U157 ( .A(npu_inst_pe_1_4_0_n28), .B(
        npu_inst_pe_1_4_0_n23), .S(npu_inst_pe_1_4_0_n8), .Z(
        npu_inst_pe_1_4_0_N94) );
  MUX2_X1 npu_inst_pe_1_4_0_U156 ( .A(npu_inst_pe_1_4_0_n25), .B(
        npu_inst_pe_1_4_0_n24), .S(npu_inst_pe_1_4_0_n6), .Z(
        npu_inst_pe_1_4_0_n28) );
  MUX2_X1 npu_inst_pe_1_4_0_U155 ( .A(npu_inst_pe_1_4_0_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_4_0_int_q_reg_v_1__1_), .S(npu_inst_pe_1_4_0_n4), .Z(
        npu_inst_pe_1_4_0_n25) );
  MUX2_X1 npu_inst_pe_1_4_0_U154 ( .A(npu_inst_pe_1_4_0_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_4_0_int_q_reg_v_3__1_), .S(npu_inst_pe_1_4_0_n4), .Z(
        npu_inst_pe_1_4_0_n24) );
  MUX2_X1 npu_inst_pe_1_4_0_U153 ( .A(npu_inst_pe_1_4_0_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_4_0_int_q_reg_v_5__1_), .S(npu_inst_pe_1_4_0_n4), .Z(
        npu_inst_pe_1_4_0_n23) );
  MUX2_X1 npu_inst_pe_1_4_0_U152 ( .A(npu_inst_pe_1_4_0_n22), .B(
        npu_inst_pe_1_4_0_n19), .S(npu_inst_pe_1_4_0_n8), .Z(
        npu_inst_pe_1_4_0_o_data_h_1_) );
  MUX2_X1 npu_inst_pe_1_4_0_U151 ( .A(npu_inst_pe_1_4_0_n21), .B(
        npu_inst_pe_1_4_0_n20), .S(npu_inst_pe_1_4_0_n6), .Z(
        npu_inst_pe_1_4_0_n22) );
  MUX2_X1 npu_inst_pe_1_4_0_U150 ( .A(npu_inst_pe_1_4_0_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_4_0_int_q_reg_h_1__1_), .S(npu_inst_pe_1_4_0_n4), .Z(
        npu_inst_pe_1_4_0_n21) );
  MUX2_X1 npu_inst_pe_1_4_0_U149 ( .A(npu_inst_pe_1_4_0_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_4_0_int_q_reg_h_3__1_), .S(npu_inst_pe_1_4_0_n4), .Z(
        npu_inst_pe_1_4_0_n20) );
  MUX2_X1 npu_inst_pe_1_4_0_U148 ( .A(npu_inst_pe_1_4_0_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_4_0_int_q_reg_h_5__1_), .S(npu_inst_pe_1_4_0_n4), .Z(
        npu_inst_pe_1_4_0_n19) );
  MUX2_X1 npu_inst_pe_1_4_0_U147 ( .A(npu_inst_pe_1_4_0_n18), .B(
        npu_inst_pe_1_4_0_n15), .S(npu_inst_pe_1_4_0_n8), .Z(
        npu_inst_pe_1_4_0_o_data_h_0_) );
  MUX2_X1 npu_inst_pe_1_4_0_U146 ( .A(npu_inst_pe_1_4_0_n17), .B(
        npu_inst_pe_1_4_0_n16), .S(npu_inst_pe_1_4_0_n6), .Z(
        npu_inst_pe_1_4_0_n18) );
  MUX2_X1 npu_inst_pe_1_4_0_U145 ( .A(npu_inst_pe_1_4_0_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_4_0_int_q_reg_h_1__0_), .S(npu_inst_pe_1_4_0_n4), .Z(
        npu_inst_pe_1_4_0_n17) );
  MUX2_X1 npu_inst_pe_1_4_0_U144 ( .A(npu_inst_pe_1_4_0_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_4_0_int_q_reg_h_3__0_), .S(npu_inst_pe_1_4_0_n4), .Z(
        npu_inst_pe_1_4_0_n16) );
  MUX2_X1 npu_inst_pe_1_4_0_U143 ( .A(npu_inst_pe_1_4_0_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_4_0_int_q_reg_h_5__0_), .S(npu_inst_pe_1_4_0_n4), .Z(
        npu_inst_pe_1_4_0_n15) );
  XOR2_X1 npu_inst_pe_1_4_0_U142 ( .A(npu_inst_pe_1_4_0_int_data_0_), .B(
        npu_inst_pe_1_4_0_int_q_acc_0_), .Z(npu_inst_pe_1_4_0_N73) );
  AND2_X1 npu_inst_pe_1_4_0_U141 ( .A1(npu_inst_pe_1_4_0_int_q_acc_0_), .A2(
        npu_inst_pe_1_4_0_int_data_0_), .ZN(npu_inst_pe_1_4_0_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_4_0_U140 ( .A(npu_inst_pe_1_4_0_int_q_acc_0_), .B(
        npu_inst_pe_1_4_0_n13), .ZN(npu_inst_pe_1_4_0_N65) );
  OR2_X1 npu_inst_pe_1_4_0_U139 ( .A1(npu_inst_pe_1_4_0_n13), .A2(
        npu_inst_pe_1_4_0_int_q_acc_0_), .ZN(npu_inst_pe_1_4_0_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_4_0_U138 ( .A(npu_inst_pe_1_4_0_int_q_acc_2_), .B(
        npu_inst_pe_1_4_0_add_79_carry_2_), .Z(npu_inst_pe_1_4_0_N75) );
  AND2_X1 npu_inst_pe_1_4_0_U137 ( .A1(npu_inst_pe_1_4_0_add_79_carry_2_), 
        .A2(npu_inst_pe_1_4_0_int_q_acc_2_), .ZN(
        npu_inst_pe_1_4_0_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_4_0_U136 ( .A(npu_inst_pe_1_4_0_int_q_acc_3_), .B(
        npu_inst_pe_1_4_0_add_79_carry_3_), .Z(npu_inst_pe_1_4_0_N76) );
  AND2_X1 npu_inst_pe_1_4_0_U135 ( .A1(npu_inst_pe_1_4_0_add_79_carry_3_), 
        .A2(npu_inst_pe_1_4_0_int_q_acc_3_), .ZN(
        npu_inst_pe_1_4_0_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_4_0_U134 ( .A(npu_inst_pe_1_4_0_int_q_acc_4_), .B(
        npu_inst_pe_1_4_0_add_79_carry_4_), .Z(npu_inst_pe_1_4_0_N77) );
  AND2_X1 npu_inst_pe_1_4_0_U133 ( .A1(npu_inst_pe_1_4_0_add_79_carry_4_), 
        .A2(npu_inst_pe_1_4_0_int_q_acc_4_), .ZN(
        npu_inst_pe_1_4_0_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_4_0_U132 ( .A(npu_inst_pe_1_4_0_int_q_acc_5_), .B(
        npu_inst_pe_1_4_0_add_79_carry_5_), .Z(npu_inst_pe_1_4_0_N78) );
  AND2_X1 npu_inst_pe_1_4_0_U131 ( .A1(npu_inst_pe_1_4_0_add_79_carry_5_), 
        .A2(npu_inst_pe_1_4_0_int_q_acc_5_), .ZN(
        npu_inst_pe_1_4_0_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_4_0_U130 ( .A(npu_inst_pe_1_4_0_int_q_acc_6_), .B(
        npu_inst_pe_1_4_0_add_79_carry_6_), .Z(npu_inst_pe_1_4_0_N79) );
  AND2_X1 npu_inst_pe_1_4_0_U129 ( .A1(npu_inst_pe_1_4_0_add_79_carry_6_), 
        .A2(npu_inst_pe_1_4_0_int_q_acc_6_), .ZN(
        npu_inst_pe_1_4_0_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_4_0_U128 ( .A(npu_inst_pe_1_4_0_int_q_acc_7_), .B(
        npu_inst_pe_1_4_0_add_79_carry_7_), .Z(npu_inst_pe_1_4_0_N80) );
  XNOR2_X1 npu_inst_pe_1_4_0_U127 ( .A(npu_inst_pe_1_4_0_sub_77_carry_2_), .B(
        npu_inst_pe_1_4_0_int_q_acc_2_), .ZN(npu_inst_pe_1_4_0_N67) );
  OR2_X1 npu_inst_pe_1_4_0_U126 ( .A1(npu_inst_pe_1_4_0_int_q_acc_2_), .A2(
        npu_inst_pe_1_4_0_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_4_0_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_4_0_U125 ( .A(npu_inst_pe_1_4_0_sub_77_carry_3_), .B(
        npu_inst_pe_1_4_0_int_q_acc_3_), .ZN(npu_inst_pe_1_4_0_N68) );
  OR2_X1 npu_inst_pe_1_4_0_U124 ( .A1(npu_inst_pe_1_4_0_int_q_acc_3_), .A2(
        npu_inst_pe_1_4_0_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_4_0_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_4_0_U123 ( .A(npu_inst_pe_1_4_0_sub_77_carry_4_), .B(
        npu_inst_pe_1_4_0_int_q_acc_4_), .ZN(npu_inst_pe_1_4_0_N69) );
  OR2_X1 npu_inst_pe_1_4_0_U122 ( .A1(npu_inst_pe_1_4_0_int_q_acc_4_), .A2(
        npu_inst_pe_1_4_0_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_4_0_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_4_0_U121 ( .A(npu_inst_pe_1_4_0_sub_77_carry_5_), .B(
        npu_inst_pe_1_4_0_int_q_acc_5_), .ZN(npu_inst_pe_1_4_0_N70) );
  OR2_X1 npu_inst_pe_1_4_0_U120 ( .A1(npu_inst_pe_1_4_0_int_q_acc_5_), .A2(
        npu_inst_pe_1_4_0_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_4_0_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_4_0_U119 ( .A(npu_inst_pe_1_4_0_sub_77_carry_6_), .B(
        npu_inst_pe_1_4_0_int_q_acc_6_), .ZN(npu_inst_pe_1_4_0_N71) );
  OR2_X1 npu_inst_pe_1_4_0_U118 ( .A1(npu_inst_pe_1_4_0_int_q_acc_6_), .A2(
        npu_inst_pe_1_4_0_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_4_0_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_4_0_U117 ( .A(npu_inst_pe_1_4_0_int_q_acc_7_), .B(
        npu_inst_pe_1_4_0_sub_77_carry_7_), .ZN(npu_inst_pe_1_4_0_N72) );
  INV_X1 npu_inst_pe_1_4_0_U116 ( .A(npu_inst_n77), .ZN(npu_inst_pe_1_4_0_n7)
         );
  INV_X1 npu_inst_pe_1_4_0_U115 ( .A(npu_inst_pe_1_4_0_n7), .ZN(
        npu_inst_pe_1_4_0_n6) );
  INV_X1 npu_inst_pe_1_4_0_U114 ( .A(npu_inst_n56), .ZN(npu_inst_pe_1_4_0_n3)
         );
  AOI22_X1 npu_inst_pe_1_4_0_U113 ( .A1(npu_inst_int_data_y_5__0__0_), .A2(
        npu_inst_pe_1_4_0_n58), .B1(npu_inst_pe_1_4_0_n114), .B2(
        npu_inst_pe_1_4_0_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_4_0_n57) );
  INV_X1 npu_inst_pe_1_4_0_U112 ( .A(npu_inst_pe_1_4_0_n57), .ZN(
        npu_inst_pe_1_4_0_n108) );
  AOI22_X1 npu_inst_pe_1_4_0_U111 ( .A1(npu_inst_int_data_y_5__0__0_), .A2(
        npu_inst_pe_1_4_0_n54), .B1(npu_inst_pe_1_4_0_n115), .B2(
        npu_inst_pe_1_4_0_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_4_0_n53) );
  INV_X1 npu_inst_pe_1_4_0_U110 ( .A(npu_inst_pe_1_4_0_n53), .ZN(
        npu_inst_pe_1_4_0_n109) );
  AOI22_X1 npu_inst_pe_1_4_0_U107 ( .A1(npu_inst_int_data_y_5__0__0_), .A2(
        npu_inst_pe_1_4_0_n50), .B1(npu_inst_pe_1_4_0_n116), .B2(
        npu_inst_pe_1_4_0_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_4_0_n49) );
  INV_X1 npu_inst_pe_1_4_0_U106 ( .A(npu_inst_pe_1_4_0_n49), .ZN(
        npu_inst_pe_1_4_0_n110) );
  AOI22_X1 npu_inst_pe_1_4_0_U105 ( .A1(npu_inst_int_data_y_5__0__0_), .A2(
        npu_inst_pe_1_4_0_n46), .B1(npu_inst_pe_1_4_0_n117), .B2(
        npu_inst_pe_1_4_0_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_4_0_n45) );
  INV_X1 npu_inst_pe_1_4_0_U104 ( .A(npu_inst_pe_1_4_0_n45), .ZN(
        npu_inst_pe_1_4_0_n111) );
  AOI22_X1 npu_inst_pe_1_4_0_U103 ( .A1(npu_inst_int_data_y_5__0__0_), .A2(
        npu_inst_pe_1_4_0_n42), .B1(npu_inst_pe_1_4_0_n119), .B2(
        npu_inst_pe_1_4_0_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_4_0_n41) );
  INV_X1 npu_inst_pe_1_4_0_U102 ( .A(npu_inst_pe_1_4_0_n41), .ZN(
        npu_inst_pe_1_4_0_n112) );
  AOI22_X1 npu_inst_pe_1_4_0_U101 ( .A1(npu_inst_int_data_y_5__0__1_), .A2(
        npu_inst_pe_1_4_0_n58), .B1(npu_inst_pe_1_4_0_n114), .B2(
        npu_inst_pe_1_4_0_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_4_0_n59) );
  INV_X1 npu_inst_pe_1_4_0_U100 ( .A(npu_inst_pe_1_4_0_n59), .ZN(
        npu_inst_pe_1_4_0_n102) );
  AOI22_X1 npu_inst_pe_1_4_0_U99 ( .A1(npu_inst_int_data_y_5__0__1_), .A2(
        npu_inst_pe_1_4_0_n54), .B1(npu_inst_pe_1_4_0_n115), .B2(
        npu_inst_pe_1_4_0_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_4_0_n55) );
  INV_X1 npu_inst_pe_1_4_0_U98 ( .A(npu_inst_pe_1_4_0_n55), .ZN(
        npu_inst_pe_1_4_0_n103) );
  AOI22_X1 npu_inst_pe_1_4_0_U97 ( .A1(npu_inst_int_data_y_5__0__1_), .A2(
        npu_inst_pe_1_4_0_n50), .B1(npu_inst_pe_1_4_0_n116), .B2(
        npu_inst_pe_1_4_0_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_4_0_n51) );
  INV_X1 npu_inst_pe_1_4_0_U96 ( .A(npu_inst_pe_1_4_0_n51), .ZN(
        npu_inst_pe_1_4_0_n104) );
  AOI22_X1 npu_inst_pe_1_4_0_U95 ( .A1(npu_inst_int_data_y_5__0__1_), .A2(
        npu_inst_pe_1_4_0_n46), .B1(npu_inst_pe_1_4_0_n117), .B2(
        npu_inst_pe_1_4_0_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_4_0_n47) );
  INV_X1 npu_inst_pe_1_4_0_U94 ( .A(npu_inst_pe_1_4_0_n47), .ZN(
        npu_inst_pe_1_4_0_n105) );
  AOI22_X1 npu_inst_pe_1_4_0_U93 ( .A1(npu_inst_int_data_y_5__0__1_), .A2(
        npu_inst_pe_1_4_0_n42), .B1(npu_inst_pe_1_4_0_n119), .B2(
        npu_inst_pe_1_4_0_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_4_0_n43) );
  INV_X1 npu_inst_pe_1_4_0_U92 ( .A(npu_inst_pe_1_4_0_n43), .ZN(
        npu_inst_pe_1_4_0_n106) );
  AOI22_X1 npu_inst_pe_1_4_0_U91 ( .A1(npu_inst_pe_1_4_0_n38), .A2(
        npu_inst_int_data_y_5__0__1_), .B1(npu_inst_pe_1_4_0_n118), .B2(
        npu_inst_pe_1_4_0_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_4_0_n39) );
  INV_X1 npu_inst_pe_1_4_0_U90 ( .A(npu_inst_pe_1_4_0_n39), .ZN(
        npu_inst_pe_1_4_0_n107) );
  AOI22_X1 npu_inst_pe_1_4_0_U89 ( .A1(npu_inst_pe_1_4_0_n38), .A2(
        npu_inst_int_data_y_5__0__0_), .B1(npu_inst_pe_1_4_0_n118), .B2(
        npu_inst_pe_1_4_0_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_4_0_n37) );
  INV_X1 npu_inst_pe_1_4_0_U88 ( .A(npu_inst_pe_1_4_0_n37), .ZN(
        npu_inst_pe_1_4_0_n113) );
  NOR3_X1 npu_inst_pe_1_4_0_U87 ( .A1(npu_inst_pe_1_4_0_n26), .A2(npu_inst_n56), .A3(npu_inst_int_ckg[31]), .ZN(npu_inst_pe_1_4_0_n85) );
  OR2_X1 npu_inst_pe_1_4_0_U86 ( .A1(npu_inst_pe_1_4_0_n85), .A2(
        npu_inst_pe_1_4_0_n2), .ZN(npu_inst_pe_1_4_0_N84) );
  NAND2_X1 npu_inst_pe_1_4_0_U85 ( .A1(npu_inst_pe_1_4_0_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_4_0_n60), .ZN(npu_inst_pe_1_4_0_n74) );
  OAI21_X1 npu_inst_pe_1_4_0_U84 ( .B1(npu_inst_pe_1_4_0_n63), .B2(
        npu_inst_pe_1_4_0_n60), .A(npu_inst_pe_1_4_0_n74), .ZN(
        npu_inst_pe_1_4_0_n97) );
  NAND2_X1 npu_inst_pe_1_4_0_U83 ( .A1(npu_inst_pe_1_4_0_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_4_0_n60), .ZN(npu_inst_pe_1_4_0_n73) );
  OAI21_X1 npu_inst_pe_1_4_0_U82 ( .B1(npu_inst_pe_1_4_0_n61), .B2(
        npu_inst_pe_1_4_0_n60), .A(npu_inst_pe_1_4_0_n73), .ZN(
        npu_inst_pe_1_4_0_n96) );
  NAND2_X1 npu_inst_pe_1_4_0_U81 ( .A1(npu_inst_pe_1_4_0_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_4_0_n56), .ZN(npu_inst_pe_1_4_0_n72) );
  OAI21_X1 npu_inst_pe_1_4_0_U80 ( .B1(npu_inst_pe_1_4_0_n63), .B2(
        npu_inst_pe_1_4_0_n56), .A(npu_inst_pe_1_4_0_n72), .ZN(
        npu_inst_pe_1_4_0_n95) );
  NAND2_X1 npu_inst_pe_1_4_0_U79 ( .A1(npu_inst_pe_1_4_0_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_4_0_n56), .ZN(npu_inst_pe_1_4_0_n71) );
  OAI21_X1 npu_inst_pe_1_4_0_U78 ( .B1(npu_inst_pe_1_4_0_n61), .B2(
        npu_inst_pe_1_4_0_n56), .A(npu_inst_pe_1_4_0_n71), .ZN(
        npu_inst_pe_1_4_0_n94) );
  NAND2_X1 npu_inst_pe_1_4_0_U77 ( .A1(npu_inst_pe_1_4_0_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_4_0_n52), .ZN(npu_inst_pe_1_4_0_n70) );
  OAI21_X1 npu_inst_pe_1_4_0_U76 ( .B1(npu_inst_pe_1_4_0_n63), .B2(
        npu_inst_pe_1_4_0_n52), .A(npu_inst_pe_1_4_0_n70), .ZN(
        npu_inst_pe_1_4_0_n93) );
  NAND2_X1 npu_inst_pe_1_4_0_U75 ( .A1(npu_inst_pe_1_4_0_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_4_0_n52), .ZN(npu_inst_pe_1_4_0_n69) );
  OAI21_X1 npu_inst_pe_1_4_0_U74 ( .B1(npu_inst_pe_1_4_0_n61), .B2(
        npu_inst_pe_1_4_0_n52), .A(npu_inst_pe_1_4_0_n69), .ZN(
        npu_inst_pe_1_4_0_n92) );
  NAND2_X1 npu_inst_pe_1_4_0_U73 ( .A1(npu_inst_pe_1_4_0_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_4_0_n48), .ZN(npu_inst_pe_1_4_0_n68) );
  OAI21_X1 npu_inst_pe_1_4_0_U72 ( .B1(npu_inst_pe_1_4_0_n63), .B2(
        npu_inst_pe_1_4_0_n48), .A(npu_inst_pe_1_4_0_n68), .ZN(
        npu_inst_pe_1_4_0_n91) );
  NAND2_X1 npu_inst_pe_1_4_0_U71 ( .A1(npu_inst_pe_1_4_0_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_4_0_n48), .ZN(npu_inst_pe_1_4_0_n67) );
  OAI21_X1 npu_inst_pe_1_4_0_U70 ( .B1(npu_inst_pe_1_4_0_n61), .B2(
        npu_inst_pe_1_4_0_n48), .A(npu_inst_pe_1_4_0_n67), .ZN(
        npu_inst_pe_1_4_0_n90) );
  NAND2_X1 npu_inst_pe_1_4_0_U69 ( .A1(npu_inst_pe_1_4_0_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_4_0_n44), .ZN(npu_inst_pe_1_4_0_n66) );
  OAI21_X1 npu_inst_pe_1_4_0_U68 ( .B1(npu_inst_pe_1_4_0_n63), .B2(
        npu_inst_pe_1_4_0_n44), .A(npu_inst_pe_1_4_0_n66), .ZN(
        npu_inst_pe_1_4_0_n89) );
  NAND2_X1 npu_inst_pe_1_4_0_U67 ( .A1(npu_inst_pe_1_4_0_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_4_0_n44), .ZN(npu_inst_pe_1_4_0_n65) );
  OAI21_X1 npu_inst_pe_1_4_0_U66 ( .B1(npu_inst_pe_1_4_0_n61), .B2(
        npu_inst_pe_1_4_0_n44), .A(npu_inst_pe_1_4_0_n65), .ZN(
        npu_inst_pe_1_4_0_n88) );
  NAND2_X1 npu_inst_pe_1_4_0_U65 ( .A1(npu_inst_pe_1_4_0_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_4_0_n40), .ZN(npu_inst_pe_1_4_0_n64) );
  OAI21_X1 npu_inst_pe_1_4_0_U64 ( .B1(npu_inst_pe_1_4_0_n63), .B2(
        npu_inst_pe_1_4_0_n40), .A(npu_inst_pe_1_4_0_n64), .ZN(
        npu_inst_pe_1_4_0_n87) );
  NAND2_X1 npu_inst_pe_1_4_0_U63 ( .A1(npu_inst_pe_1_4_0_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_4_0_n40), .ZN(npu_inst_pe_1_4_0_n62) );
  OAI21_X1 npu_inst_pe_1_4_0_U62 ( .B1(npu_inst_pe_1_4_0_n61), .B2(
        npu_inst_pe_1_4_0_n40), .A(npu_inst_pe_1_4_0_n62), .ZN(
        npu_inst_pe_1_4_0_n86) );
  AND2_X1 npu_inst_pe_1_4_0_U61 ( .A1(npu_inst_pe_1_4_0_N93), .A2(npu_inst_n56), .ZN(npu_inst_int_data_y_4__0__0_) );
  AND2_X1 npu_inst_pe_1_4_0_U60 ( .A1(npu_inst_n56), .A2(npu_inst_pe_1_4_0_N94), .ZN(npu_inst_int_data_y_4__0__1_) );
  AND2_X1 npu_inst_pe_1_4_0_U59 ( .A1(npu_inst_pe_1_4_0_int_q_acc_0_), .A2(
        npu_inst_pe_1_4_0_n1), .ZN(npu_inst_int_data_res_4__0__0_) );
  AND2_X1 npu_inst_pe_1_4_0_U58 ( .A1(npu_inst_pe_1_4_0_n2), .A2(
        npu_inst_pe_1_4_0_int_q_acc_7_), .ZN(npu_inst_int_data_res_4__0__7_)
         );
  AND2_X1 npu_inst_pe_1_4_0_U57 ( .A1(npu_inst_pe_1_4_0_int_q_acc_1_), .A2(
        npu_inst_pe_1_4_0_n1), .ZN(npu_inst_int_data_res_4__0__1_) );
  AND2_X1 npu_inst_pe_1_4_0_U56 ( .A1(npu_inst_pe_1_4_0_int_q_acc_2_), .A2(
        npu_inst_pe_1_4_0_n1), .ZN(npu_inst_int_data_res_4__0__2_) );
  AND2_X1 npu_inst_pe_1_4_0_U55 ( .A1(npu_inst_pe_1_4_0_int_q_acc_3_), .A2(
        npu_inst_pe_1_4_0_n2), .ZN(npu_inst_int_data_res_4__0__3_) );
  AND2_X1 npu_inst_pe_1_4_0_U54 ( .A1(npu_inst_pe_1_4_0_int_q_acc_4_), .A2(
        npu_inst_pe_1_4_0_n2), .ZN(npu_inst_int_data_res_4__0__4_) );
  AND2_X1 npu_inst_pe_1_4_0_U53 ( .A1(npu_inst_pe_1_4_0_int_q_acc_5_), .A2(
        npu_inst_pe_1_4_0_n2), .ZN(npu_inst_int_data_res_4__0__5_) );
  AND2_X1 npu_inst_pe_1_4_0_U52 ( .A1(npu_inst_pe_1_4_0_int_q_acc_6_), .A2(
        npu_inst_pe_1_4_0_n2), .ZN(npu_inst_int_data_res_4__0__6_) );
  AOI222_X1 npu_inst_pe_1_4_0_U51 ( .A1(npu_inst_int_data_res_5__0__0_), .A2(
        npu_inst_pe_1_4_0_n1), .B1(npu_inst_pe_1_4_0_N73), .B2(
        npu_inst_pe_1_4_0_n76), .C1(npu_inst_pe_1_4_0_N65), .C2(
        npu_inst_pe_1_4_0_n77), .ZN(npu_inst_pe_1_4_0_n84) );
  INV_X1 npu_inst_pe_1_4_0_U50 ( .A(npu_inst_pe_1_4_0_n84), .ZN(
        npu_inst_pe_1_4_0_n101) );
  AOI222_X1 npu_inst_pe_1_4_0_U49 ( .A1(npu_inst_int_data_res_5__0__7_), .A2(
        npu_inst_pe_1_4_0_n1), .B1(npu_inst_pe_1_4_0_N80), .B2(
        npu_inst_pe_1_4_0_n76), .C1(npu_inst_pe_1_4_0_N72), .C2(
        npu_inst_pe_1_4_0_n77), .ZN(npu_inst_pe_1_4_0_n75) );
  INV_X1 npu_inst_pe_1_4_0_U48 ( .A(npu_inst_pe_1_4_0_n75), .ZN(
        npu_inst_pe_1_4_0_n33) );
  AOI222_X1 npu_inst_pe_1_4_0_U47 ( .A1(npu_inst_int_data_res_5__0__1_), .A2(
        npu_inst_pe_1_4_0_n1), .B1(npu_inst_pe_1_4_0_N74), .B2(
        npu_inst_pe_1_4_0_n76), .C1(npu_inst_pe_1_4_0_N66), .C2(
        npu_inst_pe_1_4_0_n77), .ZN(npu_inst_pe_1_4_0_n83) );
  INV_X1 npu_inst_pe_1_4_0_U46 ( .A(npu_inst_pe_1_4_0_n83), .ZN(
        npu_inst_pe_1_4_0_n100) );
  AOI222_X1 npu_inst_pe_1_4_0_U45 ( .A1(npu_inst_int_data_res_5__0__2_), .A2(
        npu_inst_pe_1_4_0_n1), .B1(npu_inst_pe_1_4_0_N75), .B2(
        npu_inst_pe_1_4_0_n76), .C1(npu_inst_pe_1_4_0_N67), .C2(
        npu_inst_pe_1_4_0_n77), .ZN(npu_inst_pe_1_4_0_n82) );
  INV_X1 npu_inst_pe_1_4_0_U44 ( .A(npu_inst_pe_1_4_0_n82), .ZN(
        npu_inst_pe_1_4_0_n99) );
  AOI222_X1 npu_inst_pe_1_4_0_U43 ( .A1(npu_inst_int_data_res_5__0__3_), .A2(
        npu_inst_pe_1_4_0_n1), .B1(npu_inst_pe_1_4_0_N76), .B2(
        npu_inst_pe_1_4_0_n76), .C1(npu_inst_pe_1_4_0_N68), .C2(
        npu_inst_pe_1_4_0_n77), .ZN(npu_inst_pe_1_4_0_n81) );
  INV_X1 npu_inst_pe_1_4_0_U42 ( .A(npu_inst_pe_1_4_0_n81), .ZN(
        npu_inst_pe_1_4_0_n98) );
  AOI222_X1 npu_inst_pe_1_4_0_U41 ( .A1(npu_inst_int_data_res_5__0__4_), .A2(
        npu_inst_pe_1_4_0_n1), .B1(npu_inst_pe_1_4_0_N77), .B2(
        npu_inst_pe_1_4_0_n76), .C1(npu_inst_pe_1_4_0_N69), .C2(
        npu_inst_pe_1_4_0_n77), .ZN(npu_inst_pe_1_4_0_n80) );
  INV_X1 npu_inst_pe_1_4_0_U40 ( .A(npu_inst_pe_1_4_0_n80), .ZN(
        npu_inst_pe_1_4_0_n36) );
  AOI222_X1 npu_inst_pe_1_4_0_U39 ( .A1(npu_inst_int_data_res_5__0__5_), .A2(
        npu_inst_pe_1_4_0_n1), .B1(npu_inst_pe_1_4_0_N78), .B2(
        npu_inst_pe_1_4_0_n76), .C1(npu_inst_pe_1_4_0_N70), .C2(
        npu_inst_pe_1_4_0_n77), .ZN(npu_inst_pe_1_4_0_n79) );
  INV_X1 npu_inst_pe_1_4_0_U38 ( .A(npu_inst_pe_1_4_0_n79), .ZN(
        npu_inst_pe_1_4_0_n35) );
  AOI222_X1 npu_inst_pe_1_4_0_U37 ( .A1(npu_inst_int_data_res_5__0__6_), .A2(
        npu_inst_pe_1_4_0_n1), .B1(npu_inst_pe_1_4_0_N79), .B2(
        npu_inst_pe_1_4_0_n76), .C1(npu_inst_pe_1_4_0_N71), .C2(
        npu_inst_pe_1_4_0_n77), .ZN(npu_inst_pe_1_4_0_n78) );
  INV_X1 npu_inst_pe_1_4_0_U36 ( .A(npu_inst_pe_1_4_0_n78), .ZN(
        npu_inst_pe_1_4_0_n34) );
  AND2_X1 npu_inst_pe_1_4_0_U35 ( .A1(npu_inst_pe_1_4_0_o_data_h_1_), .A2(
        npu_inst_pe_1_4_0_int_q_weight_1_), .ZN(npu_inst_pe_1_4_0_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_4_0_U34 ( .A1(npu_inst_pe_1_4_0_o_data_h_0_), .A2(
        npu_inst_pe_1_4_0_int_q_weight_1_), .ZN(npu_inst_pe_1_4_0_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_4_0_U33 ( .A(npu_inst_pe_1_4_0_int_data_1_), .ZN(
        npu_inst_pe_1_4_0_n14) );
  AOI22_X1 npu_inst_pe_1_4_0_U32 ( .A1(npu_inst_n56), .A2(
        npu_inst_int_data_y_5__0__1_), .B1(npu_inst_pe_1_4_0_n3), .B2(
        npu_inst_int_data_x_4__1__1_), .ZN(npu_inst_pe_1_4_0_n63) );
  AOI22_X1 npu_inst_pe_1_4_0_U31 ( .A1(npu_inst_n56), .A2(
        npu_inst_int_data_y_5__0__0_), .B1(npu_inst_pe_1_4_0_n3), .B2(
        npu_inst_int_data_x_4__1__0_), .ZN(npu_inst_pe_1_4_0_n61) );
  INV_X1 npu_inst_pe_1_4_0_U30 ( .A(npu_inst_pe_1_4_0_int_data_0_), .ZN(
        npu_inst_pe_1_4_0_n13) );
  INV_X1 npu_inst_pe_1_4_0_U29 ( .A(npu_inst_n69), .ZN(npu_inst_pe_1_4_0_n5)
         );
  OR3_X1 npu_inst_pe_1_4_0_U28 ( .A1(npu_inst_pe_1_4_0_n6), .A2(
        npu_inst_pe_1_4_0_n8), .A3(npu_inst_pe_1_4_0_n5), .ZN(
        npu_inst_pe_1_4_0_n56) );
  OR3_X1 npu_inst_pe_1_4_0_U27 ( .A1(npu_inst_pe_1_4_0_n5), .A2(
        npu_inst_pe_1_4_0_n8), .A3(npu_inst_pe_1_4_0_n7), .ZN(
        npu_inst_pe_1_4_0_n48) );
  INV_X1 npu_inst_pe_1_4_0_U26 ( .A(npu_inst_pe_1_4_0_n5), .ZN(
        npu_inst_pe_1_4_0_n4) );
  INV_X1 npu_inst_pe_1_4_0_U25 ( .A(npu_inst_n124), .ZN(npu_inst_pe_1_4_0_n12)
         );
  OR3_X1 npu_inst_pe_1_4_0_U24 ( .A1(npu_inst_pe_1_4_0_n4), .A2(
        npu_inst_pe_1_4_0_n8), .A3(npu_inst_pe_1_4_0_n7), .ZN(
        npu_inst_pe_1_4_0_n52) );
  OR3_X1 npu_inst_pe_1_4_0_U23 ( .A1(npu_inst_pe_1_4_0_n6), .A2(
        npu_inst_pe_1_4_0_n8), .A3(npu_inst_pe_1_4_0_n4), .ZN(
        npu_inst_pe_1_4_0_n60) );
  NOR2_X1 npu_inst_pe_1_4_0_U22 ( .A1(npu_inst_pe_1_4_0_n60), .A2(
        npu_inst_pe_1_4_0_n3), .ZN(npu_inst_pe_1_4_0_n58) );
  NOR2_X1 npu_inst_pe_1_4_0_U21 ( .A1(npu_inst_pe_1_4_0_n56), .A2(
        npu_inst_pe_1_4_0_n3), .ZN(npu_inst_pe_1_4_0_n54) );
  NOR2_X1 npu_inst_pe_1_4_0_U20 ( .A1(npu_inst_pe_1_4_0_n52), .A2(
        npu_inst_pe_1_4_0_n3), .ZN(npu_inst_pe_1_4_0_n50) );
  NOR2_X1 npu_inst_pe_1_4_0_U19 ( .A1(npu_inst_pe_1_4_0_n48), .A2(
        npu_inst_pe_1_4_0_n3), .ZN(npu_inst_pe_1_4_0_n46) );
  NOR2_X1 npu_inst_pe_1_4_0_U18 ( .A1(npu_inst_pe_1_4_0_n40), .A2(
        npu_inst_pe_1_4_0_n3), .ZN(npu_inst_pe_1_4_0_n38) );
  NOR2_X1 npu_inst_pe_1_4_0_U17 ( .A1(npu_inst_pe_1_4_0_n44), .A2(
        npu_inst_pe_1_4_0_n3), .ZN(npu_inst_pe_1_4_0_n42) );
  BUF_X1 npu_inst_pe_1_4_0_U16 ( .A(npu_inst_n99), .Z(npu_inst_pe_1_4_0_n8) );
  BUF_X1 npu_inst_pe_1_4_0_U15 ( .A(npu_inst_pe_1_4_0_n12), .Z(
        npu_inst_pe_1_4_0_n11) );
  BUF_X1 npu_inst_pe_1_4_0_U14 ( .A(npu_inst_pe_1_4_0_n12), .Z(
        npu_inst_pe_1_4_0_n10) );
  BUF_X1 npu_inst_pe_1_4_0_U13 ( .A(npu_inst_pe_1_4_0_n12), .Z(
        npu_inst_pe_1_4_0_n9) );
  INV_X1 npu_inst_pe_1_4_0_U12 ( .A(npu_inst_pe_1_4_0_n38), .ZN(
        npu_inst_pe_1_4_0_n118) );
  INV_X1 npu_inst_pe_1_4_0_U11 ( .A(npu_inst_pe_1_4_0_n58), .ZN(
        npu_inst_pe_1_4_0_n114) );
  INV_X1 npu_inst_pe_1_4_0_U10 ( .A(npu_inst_pe_1_4_0_n54), .ZN(
        npu_inst_pe_1_4_0_n115) );
  INV_X1 npu_inst_pe_1_4_0_U9 ( .A(npu_inst_pe_1_4_0_n50), .ZN(
        npu_inst_pe_1_4_0_n116) );
  INV_X1 npu_inst_pe_1_4_0_U8 ( .A(npu_inst_pe_1_4_0_n46), .ZN(
        npu_inst_pe_1_4_0_n117) );
  INV_X1 npu_inst_pe_1_4_0_U7 ( .A(npu_inst_pe_1_4_0_n42), .ZN(
        npu_inst_pe_1_4_0_n119) );
  BUF_X1 npu_inst_pe_1_4_0_U6 ( .A(npu_inst_n22), .Z(npu_inst_pe_1_4_0_n2) );
  BUF_X1 npu_inst_pe_1_4_0_U5 ( .A(npu_inst_n22), .Z(npu_inst_pe_1_4_0_n1) );
  NOR2_X1 npu_inst_pe_1_4_0_U4 ( .A1(npu_inst_pe_1_4_0_int_q_weight_0_), .A2(
        npu_inst_pe_1_4_0_n1), .ZN(npu_inst_pe_1_4_0_n76) );
  NOR2_X1 npu_inst_pe_1_4_0_U3 ( .A1(npu_inst_pe_1_4_0_n27), .A2(
        npu_inst_pe_1_4_0_n1), .ZN(npu_inst_pe_1_4_0_n77) );
  FA_X1 npu_inst_pe_1_4_0_sub_77_U2_1 ( .A(npu_inst_pe_1_4_0_int_q_acc_1_), 
        .B(npu_inst_pe_1_4_0_n14), .CI(npu_inst_pe_1_4_0_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_4_0_sub_77_carry_2_), .S(npu_inst_pe_1_4_0_N66) );
  FA_X1 npu_inst_pe_1_4_0_add_79_U1_1 ( .A(npu_inst_pe_1_4_0_int_q_acc_1_), 
        .B(npu_inst_pe_1_4_0_int_data_1_), .CI(
        npu_inst_pe_1_4_0_add_79_carry_1_), .CO(
        npu_inst_pe_1_4_0_add_79_carry_2_), .S(npu_inst_pe_1_4_0_N74) );
  NAND3_X1 npu_inst_pe_1_4_0_U109 ( .A1(npu_inst_pe_1_4_0_n5), .A2(
        npu_inst_pe_1_4_0_n7), .A3(npu_inst_pe_1_4_0_n8), .ZN(
        npu_inst_pe_1_4_0_n44) );
  NAND3_X1 npu_inst_pe_1_4_0_U108 ( .A1(npu_inst_pe_1_4_0_n4), .A2(
        npu_inst_pe_1_4_0_n7), .A3(npu_inst_pe_1_4_0_n8), .ZN(
        npu_inst_pe_1_4_0_n40) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_4_0_n34), .CK(
        npu_inst_pe_1_4_0_net3557), .RN(npu_inst_pe_1_4_0_n9), .Q(
        npu_inst_pe_1_4_0_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_4_0_n35), .CK(
        npu_inst_pe_1_4_0_net3557), .RN(npu_inst_pe_1_4_0_n9), .Q(
        npu_inst_pe_1_4_0_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_4_0_n36), .CK(
        npu_inst_pe_1_4_0_net3557), .RN(npu_inst_pe_1_4_0_n9), .Q(
        npu_inst_pe_1_4_0_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_4_0_n98), .CK(
        npu_inst_pe_1_4_0_net3557), .RN(npu_inst_pe_1_4_0_n9), .Q(
        npu_inst_pe_1_4_0_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_4_0_n99), .CK(
        npu_inst_pe_1_4_0_net3557), .RN(npu_inst_pe_1_4_0_n9), .Q(
        npu_inst_pe_1_4_0_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_4_0_n100), 
        .CK(npu_inst_pe_1_4_0_net3557), .RN(npu_inst_pe_1_4_0_n9), .Q(
        npu_inst_pe_1_4_0_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_4_0_n33), .CK(
        npu_inst_pe_1_4_0_net3557), .RN(npu_inst_pe_1_4_0_n9), .Q(
        npu_inst_pe_1_4_0_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_4_0_n101), 
        .CK(npu_inst_pe_1_4_0_net3557), .RN(npu_inst_pe_1_4_0_n9), .Q(
        npu_inst_pe_1_4_0_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_weight_reg_0_ ( .D(npu_inst_n110), .CK(
        npu_inst_pe_1_4_0_net3563), .RN(npu_inst_pe_1_4_0_n9), .Q(
        npu_inst_pe_1_4_0_int_q_weight_0_), .QN(npu_inst_pe_1_4_0_n27) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_weight_reg_1_ ( .D(npu_inst_n116), .CK(
        npu_inst_pe_1_4_0_net3563), .RN(npu_inst_pe_1_4_0_n9), .Q(
        npu_inst_pe_1_4_0_int_q_weight_1_), .QN(npu_inst_pe_1_4_0_n26) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_4_0_n113), 
        .CK(npu_inst_pe_1_4_0_net3563), .RN(npu_inst_pe_1_4_0_n9), .Q(
        npu_inst_pe_1_4_0_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_4_0_n107), 
        .CK(npu_inst_pe_1_4_0_net3563), .RN(npu_inst_pe_1_4_0_n9), .Q(
        npu_inst_pe_1_4_0_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_4_0_n112), 
        .CK(npu_inst_pe_1_4_0_net3563), .RN(npu_inst_pe_1_4_0_n10), .Q(
        npu_inst_pe_1_4_0_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_4_0_n106), 
        .CK(npu_inst_pe_1_4_0_net3563), .RN(npu_inst_pe_1_4_0_n10), .Q(
        npu_inst_pe_1_4_0_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_4_0_n111), 
        .CK(npu_inst_pe_1_4_0_net3563), .RN(npu_inst_pe_1_4_0_n10), .Q(
        npu_inst_pe_1_4_0_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_4_0_n105), 
        .CK(npu_inst_pe_1_4_0_net3563), .RN(npu_inst_pe_1_4_0_n10), .Q(
        npu_inst_pe_1_4_0_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_4_0_n110), 
        .CK(npu_inst_pe_1_4_0_net3563), .RN(npu_inst_pe_1_4_0_n10), .Q(
        npu_inst_pe_1_4_0_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_4_0_n104), 
        .CK(npu_inst_pe_1_4_0_net3563), .RN(npu_inst_pe_1_4_0_n10), .Q(
        npu_inst_pe_1_4_0_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_4_0_n109), 
        .CK(npu_inst_pe_1_4_0_net3563), .RN(npu_inst_pe_1_4_0_n10), .Q(
        npu_inst_pe_1_4_0_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_4_0_n103), 
        .CK(npu_inst_pe_1_4_0_net3563), .RN(npu_inst_pe_1_4_0_n10), .Q(
        npu_inst_pe_1_4_0_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_4_0_n108), 
        .CK(npu_inst_pe_1_4_0_net3563), .RN(npu_inst_pe_1_4_0_n10), .Q(
        npu_inst_pe_1_4_0_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_4_0_n102), 
        .CK(npu_inst_pe_1_4_0_net3563), .RN(npu_inst_pe_1_4_0_n10), .Q(
        npu_inst_pe_1_4_0_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_4_0_n86), 
        .CK(npu_inst_pe_1_4_0_net3563), .RN(npu_inst_pe_1_4_0_n10), .Q(
        npu_inst_pe_1_4_0_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_4_0_n87), 
        .CK(npu_inst_pe_1_4_0_net3563), .RN(npu_inst_pe_1_4_0_n10), .Q(
        npu_inst_pe_1_4_0_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_4_0_n88), 
        .CK(npu_inst_pe_1_4_0_net3563), .RN(npu_inst_pe_1_4_0_n11), .Q(
        npu_inst_pe_1_4_0_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_4_0_n89), 
        .CK(npu_inst_pe_1_4_0_net3563), .RN(npu_inst_pe_1_4_0_n11), .Q(
        npu_inst_pe_1_4_0_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_4_0_n90), 
        .CK(npu_inst_pe_1_4_0_net3563), .RN(npu_inst_pe_1_4_0_n11), .Q(
        npu_inst_pe_1_4_0_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_4_0_n91), 
        .CK(npu_inst_pe_1_4_0_net3563), .RN(npu_inst_pe_1_4_0_n11), .Q(
        npu_inst_pe_1_4_0_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_4_0_n92), 
        .CK(npu_inst_pe_1_4_0_net3563), .RN(npu_inst_pe_1_4_0_n11), .Q(
        npu_inst_pe_1_4_0_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_4_0_n93), 
        .CK(npu_inst_pe_1_4_0_net3563), .RN(npu_inst_pe_1_4_0_n11), .Q(
        npu_inst_pe_1_4_0_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_4_0_n94), 
        .CK(npu_inst_pe_1_4_0_net3563), .RN(npu_inst_pe_1_4_0_n11), .Q(
        npu_inst_pe_1_4_0_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_4_0_n95), 
        .CK(npu_inst_pe_1_4_0_net3563), .RN(npu_inst_pe_1_4_0_n11), .Q(
        npu_inst_pe_1_4_0_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_4_0_n96), 
        .CK(npu_inst_pe_1_4_0_net3563), .RN(npu_inst_pe_1_4_0_n11), .Q(
        npu_inst_pe_1_4_0_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_4_0_n97), 
        .CK(npu_inst_pe_1_4_0_net3563), .RN(npu_inst_pe_1_4_0_n11), .Q(
        npu_inst_pe_1_4_0_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_4_0_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_4_0_N84), .SE(1'b0), .GCK(npu_inst_pe_1_4_0_net3557) );
  CLKGATETST_X1 npu_inst_pe_1_4_0_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n63), .SE(1'b0), .GCK(npu_inst_pe_1_4_0_net3563) );
  MUX2_X1 npu_inst_pe_1_4_1_U162 ( .A(npu_inst_pe_1_4_1_n32), .B(
        npu_inst_pe_1_4_1_n29), .S(npu_inst_pe_1_4_1_n8), .Z(
        npu_inst_pe_1_4_1_N93) );
  MUX2_X1 npu_inst_pe_1_4_1_U161 ( .A(npu_inst_pe_1_4_1_n31), .B(
        npu_inst_pe_1_4_1_n30), .S(npu_inst_pe_1_4_1_n6), .Z(
        npu_inst_pe_1_4_1_n32) );
  MUX2_X1 npu_inst_pe_1_4_1_U160 ( .A(npu_inst_pe_1_4_1_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_4_1_int_q_reg_v_1__0_), .S(npu_inst_pe_1_4_1_n4), .Z(
        npu_inst_pe_1_4_1_n31) );
  MUX2_X1 npu_inst_pe_1_4_1_U159 ( .A(npu_inst_pe_1_4_1_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_4_1_int_q_reg_v_3__0_), .S(npu_inst_pe_1_4_1_n4), .Z(
        npu_inst_pe_1_4_1_n30) );
  MUX2_X1 npu_inst_pe_1_4_1_U158 ( .A(npu_inst_pe_1_4_1_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_4_1_int_q_reg_v_5__0_), .S(npu_inst_pe_1_4_1_n4), .Z(
        npu_inst_pe_1_4_1_n29) );
  MUX2_X1 npu_inst_pe_1_4_1_U157 ( .A(npu_inst_pe_1_4_1_n28), .B(
        npu_inst_pe_1_4_1_n23), .S(npu_inst_pe_1_4_1_n8), .Z(
        npu_inst_pe_1_4_1_N94) );
  MUX2_X1 npu_inst_pe_1_4_1_U156 ( .A(npu_inst_pe_1_4_1_n25), .B(
        npu_inst_pe_1_4_1_n24), .S(npu_inst_pe_1_4_1_n6), .Z(
        npu_inst_pe_1_4_1_n28) );
  MUX2_X1 npu_inst_pe_1_4_1_U155 ( .A(npu_inst_pe_1_4_1_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_4_1_int_q_reg_v_1__1_), .S(npu_inst_pe_1_4_1_n4), .Z(
        npu_inst_pe_1_4_1_n25) );
  MUX2_X1 npu_inst_pe_1_4_1_U154 ( .A(npu_inst_pe_1_4_1_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_4_1_int_q_reg_v_3__1_), .S(npu_inst_pe_1_4_1_n4), .Z(
        npu_inst_pe_1_4_1_n24) );
  MUX2_X1 npu_inst_pe_1_4_1_U153 ( .A(npu_inst_pe_1_4_1_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_4_1_int_q_reg_v_5__1_), .S(npu_inst_pe_1_4_1_n4), .Z(
        npu_inst_pe_1_4_1_n23) );
  MUX2_X1 npu_inst_pe_1_4_1_U152 ( .A(npu_inst_pe_1_4_1_n22), .B(
        npu_inst_pe_1_4_1_n19), .S(npu_inst_pe_1_4_1_n8), .Z(
        npu_inst_int_data_x_4__1__1_) );
  MUX2_X1 npu_inst_pe_1_4_1_U151 ( .A(npu_inst_pe_1_4_1_n21), .B(
        npu_inst_pe_1_4_1_n20), .S(npu_inst_pe_1_4_1_n6), .Z(
        npu_inst_pe_1_4_1_n22) );
  MUX2_X1 npu_inst_pe_1_4_1_U150 ( .A(npu_inst_pe_1_4_1_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_4_1_int_q_reg_h_1__1_), .S(npu_inst_pe_1_4_1_n4), .Z(
        npu_inst_pe_1_4_1_n21) );
  MUX2_X1 npu_inst_pe_1_4_1_U149 ( .A(npu_inst_pe_1_4_1_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_4_1_int_q_reg_h_3__1_), .S(npu_inst_pe_1_4_1_n4), .Z(
        npu_inst_pe_1_4_1_n20) );
  MUX2_X1 npu_inst_pe_1_4_1_U148 ( .A(npu_inst_pe_1_4_1_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_4_1_int_q_reg_h_5__1_), .S(npu_inst_pe_1_4_1_n4), .Z(
        npu_inst_pe_1_4_1_n19) );
  MUX2_X1 npu_inst_pe_1_4_1_U147 ( .A(npu_inst_pe_1_4_1_n18), .B(
        npu_inst_pe_1_4_1_n15), .S(npu_inst_pe_1_4_1_n8), .Z(
        npu_inst_int_data_x_4__1__0_) );
  MUX2_X1 npu_inst_pe_1_4_1_U146 ( .A(npu_inst_pe_1_4_1_n17), .B(
        npu_inst_pe_1_4_1_n16), .S(npu_inst_pe_1_4_1_n6), .Z(
        npu_inst_pe_1_4_1_n18) );
  MUX2_X1 npu_inst_pe_1_4_1_U145 ( .A(npu_inst_pe_1_4_1_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_4_1_int_q_reg_h_1__0_), .S(npu_inst_pe_1_4_1_n4), .Z(
        npu_inst_pe_1_4_1_n17) );
  MUX2_X1 npu_inst_pe_1_4_1_U144 ( .A(npu_inst_pe_1_4_1_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_4_1_int_q_reg_h_3__0_), .S(npu_inst_pe_1_4_1_n4), .Z(
        npu_inst_pe_1_4_1_n16) );
  MUX2_X1 npu_inst_pe_1_4_1_U143 ( .A(npu_inst_pe_1_4_1_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_4_1_int_q_reg_h_5__0_), .S(npu_inst_pe_1_4_1_n4), .Z(
        npu_inst_pe_1_4_1_n15) );
  XOR2_X1 npu_inst_pe_1_4_1_U142 ( .A(npu_inst_pe_1_4_1_int_data_0_), .B(
        npu_inst_pe_1_4_1_int_q_acc_0_), .Z(npu_inst_pe_1_4_1_N73) );
  AND2_X1 npu_inst_pe_1_4_1_U141 ( .A1(npu_inst_pe_1_4_1_int_q_acc_0_), .A2(
        npu_inst_pe_1_4_1_int_data_0_), .ZN(npu_inst_pe_1_4_1_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_4_1_U140 ( .A(npu_inst_pe_1_4_1_int_q_acc_0_), .B(
        npu_inst_pe_1_4_1_n13), .ZN(npu_inst_pe_1_4_1_N65) );
  OR2_X1 npu_inst_pe_1_4_1_U139 ( .A1(npu_inst_pe_1_4_1_n13), .A2(
        npu_inst_pe_1_4_1_int_q_acc_0_), .ZN(npu_inst_pe_1_4_1_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_4_1_U138 ( .A(npu_inst_pe_1_4_1_int_q_acc_2_), .B(
        npu_inst_pe_1_4_1_add_79_carry_2_), .Z(npu_inst_pe_1_4_1_N75) );
  AND2_X1 npu_inst_pe_1_4_1_U137 ( .A1(npu_inst_pe_1_4_1_add_79_carry_2_), 
        .A2(npu_inst_pe_1_4_1_int_q_acc_2_), .ZN(
        npu_inst_pe_1_4_1_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_4_1_U136 ( .A(npu_inst_pe_1_4_1_int_q_acc_3_), .B(
        npu_inst_pe_1_4_1_add_79_carry_3_), .Z(npu_inst_pe_1_4_1_N76) );
  AND2_X1 npu_inst_pe_1_4_1_U135 ( .A1(npu_inst_pe_1_4_1_add_79_carry_3_), 
        .A2(npu_inst_pe_1_4_1_int_q_acc_3_), .ZN(
        npu_inst_pe_1_4_1_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_4_1_U134 ( .A(npu_inst_pe_1_4_1_int_q_acc_4_), .B(
        npu_inst_pe_1_4_1_add_79_carry_4_), .Z(npu_inst_pe_1_4_1_N77) );
  AND2_X1 npu_inst_pe_1_4_1_U133 ( .A1(npu_inst_pe_1_4_1_add_79_carry_4_), 
        .A2(npu_inst_pe_1_4_1_int_q_acc_4_), .ZN(
        npu_inst_pe_1_4_1_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_4_1_U132 ( .A(npu_inst_pe_1_4_1_int_q_acc_5_), .B(
        npu_inst_pe_1_4_1_add_79_carry_5_), .Z(npu_inst_pe_1_4_1_N78) );
  AND2_X1 npu_inst_pe_1_4_1_U131 ( .A1(npu_inst_pe_1_4_1_add_79_carry_5_), 
        .A2(npu_inst_pe_1_4_1_int_q_acc_5_), .ZN(
        npu_inst_pe_1_4_1_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_4_1_U130 ( .A(npu_inst_pe_1_4_1_int_q_acc_6_), .B(
        npu_inst_pe_1_4_1_add_79_carry_6_), .Z(npu_inst_pe_1_4_1_N79) );
  AND2_X1 npu_inst_pe_1_4_1_U129 ( .A1(npu_inst_pe_1_4_1_add_79_carry_6_), 
        .A2(npu_inst_pe_1_4_1_int_q_acc_6_), .ZN(
        npu_inst_pe_1_4_1_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_4_1_U128 ( .A(npu_inst_pe_1_4_1_int_q_acc_7_), .B(
        npu_inst_pe_1_4_1_add_79_carry_7_), .Z(npu_inst_pe_1_4_1_N80) );
  XNOR2_X1 npu_inst_pe_1_4_1_U127 ( .A(npu_inst_pe_1_4_1_sub_77_carry_2_), .B(
        npu_inst_pe_1_4_1_int_q_acc_2_), .ZN(npu_inst_pe_1_4_1_N67) );
  OR2_X1 npu_inst_pe_1_4_1_U126 ( .A1(npu_inst_pe_1_4_1_int_q_acc_2_), .A2(
        npu_inst_pe_1_4_1_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_4_1_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_4_1_U125 ( .A(npu_inst_pe_1_4_1_sub_77_carry_3_), .B(
        npu_inst_pe_1_4_1_int_q_acc_3_), .ZN(npu_inst_pe_1_4_1_N68) );
  OR2_X1 npu_inst_pe_1_4_1_U124 ( .A1(npu_inst_pe_1_4_1_int_q_acc_3_), .A2(
        npu_inst_pe_1_4_1_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_4_1_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_4_1_U123 ( .A(npu_inst_pe_1_4_1_sub_77_carry_4_), .B(
        npu_inst_pe_1_4_1_int_q_acc_4_), .ZN(npu_inst_pe_1_4_1_N69) );
  OR2_X1 npu_inst_pe_1_4_1_U122 ( .A1(npu_inst_pe_1_4_1_int_q_acc_4_), .A2(
        npu_inst_pe_1_4_1_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_4_1_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_4_1_U121 ( .A(npu_inst_pe_1_4_1_sub_77_carry_5_), .B(
        npu_inst_pe_1_4_1_int_q_acc_5_), .ZN(npu_inst_pe_1_4_1_N70) );
  OR2_X1 npu_inst_pe_1_4_1_U120 ( .A1(npu_inst_pe_1_4_1_int_q_acc_5_), .A2(
        npu_inst_pe_1_4_1_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_4_1_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_4_1_U119 ( .A(npu_inst_pe_1_4_1_sub_77_carry_6_), .B(
        npu_inst_pe_1_4_1_int_q_acc_6_), .ZN(npu_inst_pe_1_4_1_N71) );
  OR2_X1 npu_inst_pe_1_4_1_U118 ( .A1(npu_inst_pe_1_4_1_int_q_acc_6_), .A2(
        npu_inst_pe_1_4_1_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_4_1_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_4_1_U117 ( .A(npu_inst_pe_1_4_1_int_q_acc_7_), .B(
        npu_inst_pe_1_4_1_sub_77_carry_7_), .ZN(npu_inst_pe_1_4_1_N72) );
  INV_X1 npu_inst_pe_1_4_1_U116 ( .A(npu_inst_n77), .ZN(npu_inst_pe_1_4_1_n7)
         );
  INV_X1 npu_inst_pe_1_4_1_U115 ( .A(npu_inst_pe_1_4_1_n7), .ZN(
        npu_inst_pe_1_4_1_n6) );
  INV_X1 npu_inst_pe_1_4_1_U114 ( .A(npu_inst_n56), .ZN(npu_inst_pe_1_4_1_n3)
         );
  AOI22_X1 npu_inst_pe_1_4_1_U113 ( .A1(npu_inst_int_data_y_5__1__0_), .A2(
        npu_inst_pe_1_4_1_n58), .B1(npu_inst_pe_1_4_1_n114), .B2(
        npu_inst_pe_1_4_1_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_4_1_n57) );
  INV_X1 npu_inst_pe_1_4_1_U112 ( .A(npu_inst_pe_1_4_1_n57), .ZN(
        npu_inst_pe_1_4_1_n108) );
  AOI22_X1 npu_inst_pe_1_4_1_U111 ( .A1(npu_inst_int_data_y_5__1__0_), .A2(
        npu_inst_pe_1_4_1_n54), .B1(npu_inst_pe_1_4_1_n115), .B2(
        npu_inst_pe_1_4_1_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_4_1_n53) );
  INV_X1 npu_inst_pe_1_4_1_U110 ( .A(npu_inst_pe_1_4_1_n53), .ZN(
        npu_inst_pe_1_4_1_n109) );
  AOI22_X1 npu_inst_pe_1_4_1_U107 ( .A1(npu_inst_int_data_y_5__1__0_), .A2(
        npu_inst_pe_1_4_1_n50), .B1(npu_inst_pe_1_4_1_n116), .B2(
        npu_inst_pe_1_4_1_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_4_1_n49) );
  INV_X1 npu_inst_pe_1_4_1_U106 ( .A(npu_inst_pe_1_4_1_n49), .ZN(
        npu_inst_pe_1_4_1_n110) );
  AOI22_X1 npu_inst_pe_1_4_1_U105 ( .A1(npu_inst_int_data_y_5__1__0_), .A2(
        npu_inst_pe_1_4_1_n46), .B1(npu_inst_pe_1_4_1_n117), .B2(
        npu_inst_pe_1_4_1_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_4_1_n45) );
  INV_X1 npu_inst_pe_1_4_1_U104 ( .A(npu_inst_pe_1_4_1_n45), .ZN(
        npu_inst_pe_1_4_1_n111) );
  AOI22_X1 npu_inst_pe_1_4_1_U103 ( .A1(npu_inst_int_data_y_5__1__0_), .A2(
        npu_inst_pe_1_4_1_n42), .B1(npu_inst_pe_1_4_1_n119), .B2(
        npu_inst_pe_1_4_1_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_4_1_n41) );
  INV_X1 npu_inst_pe_1_4_1_U102 ( .A(npu_inst_pe_1_4_1_n41), .ZN(
        npu_inst_pe_1_4_1_n112) );
  AOI22_X1 npu_inst_pe_1_4_1_U101 ( .A1(npu_inst_int_data_y_5__1__1_), .A2(
        npu_inst_pe_1_4_1_n58), .B1(npu_inst_pe_1_4_1_n114), .B2(
        npu_inst_pe_1_4_1_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_4_1_n59) );
  INV_X1 npu_inst_pe_1_4_1_U100 ( .A(npu_inst_pe_1_4_1_n59), .ZN(
        npu_inst_pe_1_4_1_n102) );
  AOI22_X1 npu_inst_pe_1_4_1_U99 ( .A1(npu_inst_int_data_y_5__1__1_), .A2(
        npu_inst_pe_1_4_1_n54), .B1(npu_inst_pe_1_4_1_n115), .B2(
        npu_inst_pe_1_4_1_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_4_1_n55) );
  INV_X1 npu_inst_pe_1_4_1_U98 ( .A(npu_inst_pe_1_4_1_n55), .ZN(
        npu_inst_pe_1_4_1_n103) );
  AOI22_X1 npu_inst_pe_1_4_1_U97 ( .A1(npu_inst_int_data_y_5__1__1_), .A2(
        npu_inst_pe_1_4_1_n50), .B1(npu_inst_pe_1_4_1_n116), .B2(
        npu_inst_pe_1_4_1_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_4_1_n51) );
  INV_X1 npu_inst_pe_1_4_1_U96 ( .A(npu_inst_pe_1_4_1_n51), .ZN(
        npu_inst_pe_1_4_1_n104) );
  AOI22_X1 npu_inst_pe_1_4_1_U95 ( .A1(npu_inst_int_data_y_5__1__1_), .A2(
        npu_inst_pe_1_4_1_n46), .B1(npu_inst_pe_1_4_1_n117), .B2(
        npu_inst_pe_1_4_1_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_4_1_n47) );
  INV_X1 npu_inst_pe_1_4_1_U94 ( .A(npu_inst_pe_1_4_1_n47), .ZN(
        npu_inst_pe_1_4_1_n105) );
  AOI22_X1 npu_inst_pe_1_4_1_U93 ( .A1(npu_inst_int_data_y_5__1__1_), .A2(
        npu_inst_pe_1_4_1_n42), .B1(npu_inst_pe_1_4_1_n119), .B2(
        npu_inst_pe_1_4_1_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_4_1_n43) );
  INV_X1 npu_inst_pe_1_4_1_U92 ( .A(npu_inst_pe_1_4_1_n43), .ZN(
        npu_inst_pe_1_4_1_n106) );
  AOI22_X1 npu_inst_pe_1_4_1_U91 ( .A1(npu_inst_pe_1_4_1_n38), .A2(
        npu_inst_int_data_y_5__1__1_), .B1(npu_inst_pe_1_4_1_n118), .B2(
        npu_inst_pe_1_4_1_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_4_1_n39) );
  INV_X1 npu_inst_pe_1_4_1_U90 ( .A(npu_inst_pe_1_4_1_n39), .ZN(
        npu_inst_pe_1_4_1_n107) );
  AOI22_X1 npu_inst_pe_1_4_1_U89 ( .A1(npu_inst_pe_1_4_1_n38), .A2(
        npu_inst_int_data_y_5__1__0_), .B1(npu_inst_pe_1_4_1_n118), .B2(
        npu_inst_pe_1_4_1_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_4_1_n37) );
  INV_X1 npu_inst_pe_1_4_1_U88 ( .A(npu_inst_pe_1_4_1_n37), .ZN(
        npu_inst_pe_1_4_1_n113) );
  NAND2_X1 npu_inst_pe_1_4_1_U87 ( .A1(npu_inst_pe_1_4_1_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_4_1_n60), .ZN(npu_inst_pe_1_4_1_n74) );
  OAI21_X1 npu_inst_pe_1_4_1_U86 ( .B1(npu_inst_pe_1_4_1_n63), .B2(
        npu_inst_pe_1_4_1_n60), .A(npu_inst_pe_1_4_1_n74), .ZN(
        npu_inst_pe_1_4_1_n97) );
  NAND2_X1 npu_inst_pe_1_4_1_U85 ( .A1(npu_inst_pe_1_4_1_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_4_1_n60), .ZN(npu_inst_pe_1_4_1_n73) );
  OAI21_X1 npu_inst_pe_1_4_1_U84 ( .B1(npu_inst_pe_1_4_1_n61), .B2(
        npu_inst_pe_1_4_1_n60), .A(npu_inst_pe_1_4_1_n73), .ZN(
        npu_inst_pe_1_4_1_n96) );
  NAND2_X1 npu_inst_pe_1_4_1_U83 ( .A1(npu_inst_pe_1_4_1_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_4_1_n56), .ZN(npu_inst_pe_1_4_1_n72) );
  OAI21_X1 npu_inst_pe_1_4_1_U82 ( .B1(npu_inst_pe_1_4_1_n63), .B2(
        npu_inst_pe_1_4_1_n56), .A(npu_inst_pe_1_4_1_n72), .ZN(
        npu_inst_pe_1_4_1_n95) );
  NAND2_X1 npu_inst_pe_1_4_1_U81 ( .A1(npu_inst_pe_1_4_1_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_4_1_n56), .ZN(npu_inst_pe_1_4_1_n71) );
  OAI21_X1 npu_inst_pe_1_4_1_U80 ( .B1(npu_inst_pe_1_4_1_n61), .B2(
        npu_inst_pe_1_4_1_n56), .A(npu_inst_pe_1_4_1_n71), .ZN(
        npu_inst_pe_1_4_1_n94) );
  NAND2_X1 npu_inst_pe_1_4_1_U79 ( .A1(npu_inst_pe_1_4_1_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_4_1_n52), .ZN(npu_inst_pe_1_4_1_n70) );
  OAI21_X1 npu_inst_pe_1_4_1_U78 ( .B1(npu_inst_pe_1_4_1_n63), .B2(
        npu_inst_pe_1_4_1_n52), .A(npu_inst_pe_1_4_1_n70), .ZN(
        npu_inst_pe_1_4_1_n93) );
  NAND2_X1 npu_inst_pe_1_4_1_U77 ( .A1(npu_inst_pe_1_4_1_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_4_1_n52), .ZN(npu_inst_pe_1_4_1_n69) );
  OAI21_X1 npu_inst_pe_1_4_1_U76 ( .B1(npu_inst_pe_1_4_1_n61), .B2(
        npu_inst_pe_1_4_1_n52), .A(npu_inst_pe_1_4_1_n69), .ZN(
        npu_inst_pe_1_4_1_n92) );
  NAND2_X1 npu_inst_pe_1_4_1_U75 ( .A1(npu_inst_pe_1_4_1_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_4_1_n48), .ZN(npu_inst_pe_1_4_1_n68) );
  OAI21_X1 npu_inst_pe_1_4_1_U74 ( .B1(npu_inst_pe_1_4_1_n63), .B2(
        npu_inst_pe_1_4_1_n48), .A(npu_inst_pe_1_4_1_n68), .ZN(
        npu_inst_pe_1_4_1_n91) );
  NAND2_X1 npu_inst_pe_1_4_1_U73 ( .A1(npu_inst_pe_1_4_1_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_4_1_n48), .ZN(npu_inst_pe_1_4_1_n67) );
  OAI21_X1 npu_inst_pe_1_4_1_U72 ( .B1(npu_inst_pe_1_4_1_n61), .B2(
        npu_inst_pe_1_4_1_n48), .A(npu_inst_pe_1_4_1_n67), .ZN(
        npu_inst_pe_1_4_1_n90) );
  NAND2_X1 npu_inst_pe_1_4_1_U71 ( .A1(npu_inst_pe_1_4_1_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_4_1_n44), .ZN(npu_inst_pe_1_4_1_n66) );
  OAI21_X1 npu_inst_pe_1_4_1_U70 ( .B1(npu_inst_pe_1_4_1_n63), .B2(
        npu_inst_pe_1_4_1_n44), .A(npu_inst_pe_1_4_1_n66), .ZN(
        npu_inst_pe_1_4_1_n89) );
  NAND2_X1 npu_inst_pe_1_4_1_U69 ( .A1(npu_inst_pe_1_4_1_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_4_1_n44), .ZN(npu_inst_pe_1_4_1_n65) );
  OAI21_X1 npu_inst_pe_1_4_1_U68 ( .B1(npu_inst_pe_1_4_1_n61), .B2(
        npu_inst_pe_1_4_1_n44), .A(npu_inst_pe_1_4_1_n65), .ZN(
        npu_inst_pe_1_4_1_n88) );
  NAND2_X1 npu_inst_pe_1_4_1_U67 ( .A1(npu_inst_pe_1_4_1_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_4_1_n40), .ZN(npu_inst_pe_1_4_1_n64) );
  OAI21_X1 npu_inst_pe_1_4_1_U66 ( .B1(npu_inst_pe_1_4_1_n63), .B2(
        npu_inst_pe_1_4_1_n40), .A(npu_inst_pe_1_4_1_n64), .ZN(
        npu_inst_pe_1_4_1_n87) );
  NAND2_X1 npu_inst_pe_1_4_1_U65 ( .A1(npu_inst_pe_1_4_1_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_4_1_n40), .ZN(npu_inst_pe_1_4_1_n62) );
  OAI21_X1 npu_inst_pe_1_4_1_U64 ( .B1(npu_inst_pe_1_4_1_n61), .B2(
        npu_inst_pe_1_4_1_n40), .A(npu_inst_pe_1_4_1_n62), .ZN(
        npu_inst_pe_1_4_1_n86) );
  AND2_X1 npu_inst_pe_1_4_1_U63 ( .A1(npu_inst_pe_1_4_1_N93), .A2(npu_inst_n56), .ZN(npu_inst_int_data_y_4__1__0_) );
  AND2_X1 npu_inst_pe_1_4_1_U62 ( .A1(npu_inst_n56), .A2(npu_inst_pe_1_4_1_N94), .ZN(npu_inst_int_data_y_4__1__1_) );
  NOR3_X1 npu_inst_pe_1_4_1_U61 ( .A1(npu_inst_pe_1_4_1_n26), .A2(npu_inst_n56), .A3(npu_inst_int_ckg[30]), .ZN(npu_inst_pe_1_4_1_n85) );
  OR2_X1 npu_inst_pe_1_4_1_U60 ( .A1(npu_inst_pe_1_4_1_n85), .A2(
        npu_inst_pe_1_4_1_n2), .ZN(npu_inst_pe_1_4_1_N84) );
  AND2_X1 npu_inst_pe_1_4_1_U59 ( .A1(npu_inst_pe_1_4_1_int_q_acc_0_), .A2(
        npu_inst_pe_1_4_1_n1), .ZN(npu_inst_int_data_res_4__1__0_) );
  AND2_X1 npu_inst_pe_1_4_1_U58 ( .A1(npu_inst_pe_1_4_1_n2), .A2(
        npu_inst_pe_1_4_1_int_q_acc_7_), .ZN(npu_inst_int_data_res_4__1__7_)
         );
  AND2_X1 npu_inst_pe_1_4_1_U57 ( .A1(npu_inst_pe_1_4_1_int_q_acc_1_), .A2(
        npu_inst_pe_1_4_1_n1), .ZN(npu_inst_int_data_res_4__1__1_) );
  AND2_X1 npu_inst_pe_1_4_1_U56 ( .A1(npu_inst_pe_1_4_1_int_q_acc_2_), .A2(
        npu_inst_pe_1_4_1_n1), .ZN(npu_inst_int_data_res_4__1__2_) );
  AND2_X1 npu_inst_pe_1_4_1_U55 ( .A1(npu_inst_pe_1_4_1_int_q_acc_3_), .A2(
        npu_inst_pe_1_4_1_n2), .ZN(npu_inst_int_data_res_4__1__3_) );
  AND2_X1 npu_inst_pe_1_4_1_U54 ( .A1(npu_inst_pe_1_4_1_int_q_acc_4_), .A2(
        npu_inst_pe_1_4_1_n2), .ZN(npu_inst_int_data_res_4__1__4_) );
  AND2_X1 npu_inst_pe_1_4_1_U53 ( .A1(npu_inst_pe_1_4_1_int_q_acc_5_), .A2(
        npu_inst_pe_1_4_1_n2), .ZN(npu_inst_int_data_res_4__1__5_) );
  AND2_X1 npu_inst_pe_1_4_1_U52 ( .A1(npu_inst_pe_1_4_1_int_q_acc_6_), .A2(
        npu_inst_pe_1_4_1_n2), .ZN(npu_inst_int_data_res_4__1__6_) );
  AOI222_X1 npu_inst_pe_1_4_1_U51 ( .A1(npu_inst_int_data_res_5__1__0_), .A2(
        npu_inst_pe_1_4_1_n1), .B1(npu_inst_pe_1_4_1_N73), .B2(
        npu_inst_pe_1_4_1_n76), .C1(npu_inst_pe_1_4_1_N65), .C2(
        npu_inst_pe_1_4_1_n77), .ZN(npu_inst_pe_1_4_1_n84) );
  INV_X1 npu_inst_pe_1_4_1_U50 ( .A(npu_inst_pe_1_4_1_n84), .ZN(
        npu_inst_pe_1_4_1_n101) );
  AOI222_X1 npu_inst_pe_1_4_1_U49 ( .A1(npu_inst_int_data_res_5__1__7_), .A2(
        npu_inst_pe_1_4_1_n1), .B1(npu_inst_pe_1_4_1_N80), .B2(
        npu_inst_pe_1_4_1_n76), .C1(npu_inst_pe_1_4_1_N72), .C2(
        npu_inst_pe_1_4_1_n77), .ZN(npu_inst_pe_1_4_1_n75) );
  INV_X1 npu_inst_pe_1_4_1_U48 ( .A(npu_inst_pe_1_4_1_n75), .ZN(
        npu_inst_pe_1_4_1_n33) );
  AOI222_X1 npu_inst_pe_1_4_1_U47 ( .A1(npu_inst_int_data_res_5__1__1_), .A2(
        npu_inst_pe_1_4_1_n1), .B1(npu_inst_pe_1_4_1_N74), .B2(
        npu_inst_pe_1_4_1_n76), .C1(npu_inst_pe_1_4_1_N66), .C2(
        npu_inst_pe_1_4_1_n77), .ZN(npu_inst_pe_1_4_1_n83) );
  INV_X1 npu_inst_pe_1_4_1_U46 ( .A(npu_inst_pe_1_4_1_n83), .ZN(
        npu_inst_pe_1_4_1_n100) );
  AOI222_X1 npu_inst_pe_1_4_1_U45 ( .A1(npu_inst_int_data_res_5__1__2_), .A2(
        npu_inst_pe_1_4_1_n1), .B1(npu_inst_pe_1_4_1_N75), .B2(
        npu_inst_pe_1_4_1_n76), .C1(npu_inst_pe_1_4_1_N67), .C2(
        npu_inst_pe_1_4_1_n77), .ZN(npu_inst_pe_1_4_1_n82) );
  INV_X1 npu_inst_pe_1_4_1_U44 ( .A(npu_inst_pe_1_4_1_n82), .ZN(
        npu_inst_pe_1_4_1_n99) );
  AOI222_X1 npu_inst_pe_1_4_1_U43 ( .A1(npu_inst_int_data_res_5__1__3_), .A2(
        npu_inst_pe_1_4_1_n1), .B1(npu_inst_pe_1_4_1_N76), .B2(
        npu_inst_pe_1_4_1_n76), .C1(npu_inst_pe_1_4_1_N68), .C2(
        npu_inst_pe_1_4_1_n77), .ZN(npu_inst_pe_1_4_1_n81) );
  INV_X1 npu_inst_pe_1_4_1_U42 ( .A(npu_inst_pe_1_4_1_n81), .ZN(
        npu_inst_pe_1_4_1_n98) );
  AOI222_X1 npu_inst_pe_1_4_1_U41 ( .A1(npu_inst_int_data_res_5__1__4_), .A2(
        npu_inst_pe_1_4_1_n1), .B1(npu_inst_pe_1_4_1_N77), .B2(
        npu_inst_pe_1_4_1_n76), .C1(npu_inst_pe_1_4_1_N69), .C2(
        npu_inst_pe_1_4_1_n77), .ZN(npu_inst_pe_1_4_1_n80) );
  INV_X1 npu_inst_pe_1_4_1_U40 ( .A(npu_inst_pe_1_4_1_n80), .ZN(
        npu_inst_pe_1_4_1_n36) );
  AOI222_X1 npu_inst_pe_1_4_1_U39 ( .A1(npu_inst_int_data_res_5__1__5_), .A2(
        npu_inst_pe_1_4_1_n1), .B1(npu_inst_pe_1_4_1_N78), .B2(
        npu_inst_pe_1_4_1_n76), .C1(npu_inst_pe_1_4_1_N70), .C2(
        npu_inst_pe_1_4_1_n77), .ZN(npu_inst_pe_1_4_1_n79) );
  INV_X1 npu_inst_pe_1_4_1_U38 ( .A(npu_inst_pe_1_4_1_n79), .ZN(
        npu_inst_pe_1_4_1_n35) );
  AOI222_X1 npu_inst_pe_1_4_1_U37 ( .A1(npu_inst_int_data_res_5__1__6_), .A2(
        npu_inst_pe_1_4_1_n1), .B1(npu_inst_pe_1_4_1_N79), .B2(
        npu_inst_pe_1_4_1_n76), .C1(npu_inst_pe_1_4_1_N71), .C2(
        npu_inst_pe_1_4_1_n77), .ZN(npu_inst_pe_1_4_1_n78) );
  INV_X1 npu_inst_pe_1_4_1_U36 ( .A(npu_inst_pe_1_4_1_n78), .ZN(
        npu_inst_pe_1_4_1_n34) );
  INV_X1 npu_inst_pe_1_4_1_U35 ( .A(npu_inst_pe_1_4_1_int_data_1_), .ZN(
        npu_inst_pe_1_4_1_n14) );
  AND2_X1 npu_inst_pe_1_4_1_U34 ( .A1(npu_inst_int_data_x_4__1__1_), .A2(
        npu_inst_pe_1_4_1_int_q_weight_1_), .ZN(npu_inst_pe_1_4_1_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_4_1_U33 ( .A1(npu_inst_int_data_x_4__1__0_), .A2(
        npu_inst_pe_1_4_1_int_q_weight_1_), .ZN(npu_inst_pe_1_4_1_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_4_1_U32 ( .A1(npu_inst_n56), .A2(
        npu_inst_int_data_y_5__1__1_), .B1(npu_inst_pe_1_4_1_n3), .B2(
        npu_inst_int_data_x_4__2__1_), .ZN(npu_inst_pe_1_4_1_n63) );
  AOI22_X1 npu_inst_pe_1_4_1_U31 ( .A1(npu_inst_n56), .A2(
        npu_inst_int_data_y_5__1__0_), .B1(npu_inst_pe_1_4_1_n3), .B2(
        npu_inst_int_data_x_4__2__0_), .ZN(npu_inst_pe_1_4_1_n61) );
  INV_X1 npu_inst_pe_1_4_1_U30 ( .A(npu_inst_pe_1_4_1_int_data_0_), .ZN(
        npu_inst_pe_1_4_1_n13) );
  INV_X1 npu_inst_pe_1_4_1_U29 ( .A(npu_inst_n69), .ZN(npu_inst_pe_1_4_1_n5)
         );
  OR3_X1 npu_inst_pe_1_4_1_U28 ( .A1(npu_inst_pe_1_4_1_n6), .A2(
        npu_inst_pe_1_4_1_n8), .A3(npu_inst_pe_1_4_1_n5), .ZN(
        npu_inst_pe_1_4_1_n56) );
  OR3_X1 npu_inst_pe_1_4_1_U27 ( .A1(npu_inst_pe_1_4_1_n5), .A2(
        npu_inst_pe_1_4_1_n8), .A3(npu_inst_pe_1_4_1_n7), .ZN(
        npu_inst_pe_1_4_1_n48) );
  INV_X1 npu_inst_pe_1_4_1_U26 ( .A(npu_inst_pe_1_4_1_n5), .ZN(
        npu_inst_pe_1_4_1_n4) );
  INV_X1 npu_inst_pe_1_4_1_U25 ( .A(npu_inst_n124), .ZN(npu_inst_pe_1_4_1_n12)
         );
  OR3_X1 npu_inst_pe_1_4_1_U24 ( .A1(npu_inst_pe_1_4_1_n4), .A2(
        npu_inst_pe_1_4_1_n8), .A3(npu_inst_pe_1_4_1_n7), .ZN(
        npu_inst_pe_1_4_1_n52) );
  OR3_X1 npu_inst_pe_1_4_1_U23 ( .A1(npu_inst_pe_1_4_1_n6), .A2(
        npu_inst_pe_1_4_1_n8), .A3(npu_inst_pe_1_4_1_n4), .ZN(
        npu_inst_pe_1_4_1_n60) );
  NOR2_X1 npu_inst_pe_1_4_1_U22 ( .A1(npu_inst_pe_1_4_1_n60), .A2(
        npu_inst_pe_1_4_1_n3), .ZN(npu_inst_pe_1_4_1_n58) );
  NOR2_X1 npu_inst_pe_1_4_1_U21 ( .A1(npu_inst_pe_1_4_1_n56), .A2(
        npu_inst_pe_1_4_1_n3), .ZN(npu_inst_pe_1_4_1_n54) );
  NOR2_X1 npu_inst_pe_1_4_1_U20 ( .A1(npu_inst_pe_1_4_1_n52), .A2(
        npu_inst_pe_1_4_1_n3), .ZN(npu_inst_pe_1_4_1_n50) );
  NOR2_X1 npu_inst_pe_1_4_1_U19 ( .A1(npu_inst_pe_1_4_1_n48), .A2(
        npu_inst_pe_1_4_1_n3), .ZN(npu_inst_pe_1_4_1_n46) );
  NOR2_X1 npu_inst_pe_1_4_1_U18 ( .A1(npu_inst_pe_1_4_1_n40), .A2(
        npu_inst_pe_1_4_1_n3), .ZN(npu_inst_pe_1_4_1_n38) );
  NOR2_X1 npu_inst_pe_1_4_1_U17 ( .A1(npu_inst_pe_1_4_1_n44), .A2(
        npu_inst_pe_1_4_1_n3), .ZN(npu_inst_pe_1_4_1_n42) );
  BUF_X1 npu_inst_pe_1_4_1_U16 ( .A(npu_inst_n99), .Z(npu_inst_pe_1_4_1_n8) );
  BUF_X1 npu_inst_pe_1_4_1_U15 ( .A(npu_inst_pe_1_4_1_n12), .Z(
        npu_inst_pe_1_4_1_n11) );
  BUF_X1 npu_inst_pe_1_4_1_U14 ( .A(npu_inst_pe_1_4_1_n12), .Z(
        npu_inst_pe_1_4_1_n10) );
  BUF_X1 npu_inst_pe_1_4_1_U13 ( .A(npu_inst_pe_1_4_1_n12), .Z(
        npu_inst_pe_1_4_1_n9) );
  INV_X1 npu_inst_pe_1_4_1_U12 ( .A(npu_inst_pe_1_4_1_n38), .ZN(
        npu_inst_pe_1_4_1_n118) );
  INV_X1 npu_inst_pe_1_4_1_U11 ( .A(npu_inst_pe_1_4_1_n58), .ZN(
        npu_inst_pe_1_4_1_n114) );
  INV_X1 npu_inst_pe_1_4_1_U10 ( .A(npu_inst_pe_1_4_1_n54), .ZN(
        npu_inst_pe_1_4_1_n115) );
  INV_X1 npu_inst_pe_1_4_1_U9 ( .A(npu_inst_pe_1_4_1_n50), .ZN(
        npu_inst_pe_1_4_1_n116) );
  INV_X1 npu_inst_pe_1_4_1_U8 ( .A(npu_inst_pe_1_4_1_n46), .ZN(
        npu_inst_pe_1_4_1_n117) );
  INV_X1 npu_inst_pe_1_4_1_U7 ( .A(npu_inst_pe_1_4_1_n42), .ZN(
        npu_inst_pe_1_4_1_n119) );
  BUF_X1 npu_inst_pe_1_4_1_U6 ( .A(npu_inst_n22), .Z(npu_inst_pe_1_4_1_n2) );
  BUF_X1 npu_inst_pe_1_4_1_U5 ( .A(npu_inst_n22), .Z(npu_inst_pe_1_4_1_n1) );
  NOR2_X1 npu_inst_pe_1_4_1_U4 ( .A1(npu_inst_pe_1_4_1_int_q_weight_0_), .A2(
        npu_inst_pe_1_4_1_n1), .ZN(npu_inst_pe_1_4_1_n76) );
  NOR2_X1 npu_inst_pe_1_4_1_U3 ( .A1(npu_inst_pe_1_4_1_n27), .A2(
        npu_inst_pe_1_4_1_n1), .ZN(npu_inst_pe_1_4_1_n77) );
  FA_X1 npu_inst_pe_1_4_1_sub_77_U2_1 ( .A(npu_inst_pe_1_4_1_int_q_acc_1_), 
        .B(npu_inst_pe_1_4_1_n14), .CI(npu_inst_pe_1_4_1_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_4_1_sub_77_carry_2_), .S(npu_inst_pe_1_4_1_N66) );
  FA_X1 npu_inst_pe_1_4_1_add_79_U1_1 ( .A(npu_inst_pe_1_4_1_int_q_acc_1_), 
        .B(npu_inst_pe_1_4_1_int_data_1_), .CI(
        npu_inst_pe_1_4_1_add_79_carry_1_), .CO(
        npu_inst_pe_1_4_1_add_79_carry_2_), .S(npu_inst_pe_1_4_1_N74) );
  NAND3_X1 npu_inst_pe_1_4_1_U109 ( .A1(npu_inst_pe_1_4_1_n5), .A2(
        npu_inst_pe_1_4_1_n7), .A3(npu_inst_pe_1_4_1_n8), .ZN(
        npu_inst_pe_1_4_1_n44) );
  NAND3_X1 npu_inst_pe_1_4_1_U108 ( .A1(npu_inst_pe_1_4_1_n4), .A2(
        npu_inst_pe_1_4_1_n7), .A3(npu_inst_pe_1_4_1_n8), .ZN(
        npu_inst_pe_1_4_1_n40) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_4_1_n34), .CK(
        npu_inst_pe_1_4_1_net3534), .RN(npu_inst_pe_1_4_1_n9), .Q(
        npu_inst_pe_1_4_1_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_4_1_n35), .CK(
        npu_inst_pe_1_4_1_net3534), .RN(npu_inst_pe_1_4_1_n9), .Q(
        npu_inst_pe_1_4_1_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_4_1_n36), .CK(
        npu_inst_pe_1_4_1_net3534), .RN(npu_inst_pe_1_4_1_n9), .Q(
        npu_inst_pe_1_4_1_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_4_1_n98), .CK(
        npu_inst_pe_1_4_1_net3534), .RN(npu_inst_pe_1_4_1_n9), .Q(
        npu_inst_pe_1_4_1_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_4_1_n99), .CK(
        npu_inst_pe_1_4_1_net3534), .RN(npu_inst_pe_1_4_1_n9), .Q(
        npu_inst_pe_1_4_1_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_4_1_n100), 
        .CK(npu_inst_pe_1_4_1_net3534), .RN(npu_inst_pe_1_4_1_n9), .Q(
        npu_inst_pe_1_4_1_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_4_1_n33), .CK(
        npu_inst_pe_1_4_1_net3534), .RN(npu_inst_pe_1_4_1_n9), .Q(
        npu_inst_pe_1_4_1_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_4_1_n101), 
        .CK(npu_inst_pe_1_4_1_net3534), .RN(npu_inst_pe_1_4_1_n9), .Q(
        npu_inst_pe_1_4_1_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_weight_reg_0_ ( .D(npu_inst_n110), .CK(
        npu_inst_pe_1_4_1_net3540), .RN(npu_inst_pe_1_4_1_n9), .Q(
        npu_inst_pe_1_4_1_int_q_weight_0_), .QN(npu_inst_pe_1_4_1_n27) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_weight_reg_1_ ( .D(npu_inst_n116), .CK(
        npu_inst_pe_1_4_1_net3540), .RN(npu_inst_pe_1_4_1_n9), .Q(
        npu_inst_pe_1_4_1_int_q_weight_1_), .QN(npu_inst_pe_1_4_1_n26) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_4_1_n113), 
        .CK(npu_inst_pe_1_4_1_net3540), .RN(npu_inst_pe_1_4_1_n9), .Q(
        npu_inst_pe_1_4_1_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_4_1_n107), 
        .CK(npu_inst_pe_1_4_1_net3540), .RN(npu_inst_pe_1_4_1_n9), .Q(
        npu_inst_pe_1_4_1_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_4_1_n112), 
        .CK(npu_inst_pe_1_4_1_net3540), .RN(npu_inst_pe_1_4_1_n10), .Q(
        npu_inst_pe_1_4_1_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_4_1_n106), 
        .CK(npu_inst_pe_1_4_1_net3540), .RN(npu_inst_pe_1_4_1_n10), .Q(
        npu_inst_pe_1_4_1_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_4_1_n111), 
        .CK(npu_inst_pe_1_4_1_net3540), .RN(npu_inst_pe_1_4_1_n10), .Q(
        npu_inst_pe_1_4_1_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_4_1_n105), 
        .CK(npu_inst_pe_1_4_1_net3540), .RN(npu_inst_pe_1_4_1_n10), .Q(
        npu_inst_pe_1_4_1_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_4_1_n110), 
        .CK(npu_inst_pe_1_4_1_net3540), .RN(npu_inst_pe_1_4_1_n10), .Q(
        npu_inst_pe_1_4_1_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_4_1_n104), 
        .CK(npu_inst_pe_1_4_1_net3540), .RN(npu_inst_pe_1_4_1_n10), .Q(
        npu_inst_pe_1_4_1_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_4_1_n109), 
        .CK(npu_inst_pe_1_4_1_net3540), .RN(npu_inst_pe_1_4_1_n10), .Q(
        npu_inst_pe_1_4_1_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_4_1_n103), 
        .CK(npu_inst_pe_1_4_1_net3540), .RN(npu_inst_pe_1_4_1_n10), .Q(
        npu_inst_pe_1_4_1_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_4_1_n108), 
        .CK(npu_inst_pe_1_4_1_net3540), .RN(npu_inst_pe_1_4_1_n10), .Q(
        npu_inst_pe_1_4_1_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_4_1_n102), 
        .CK(npu_inst_pe_1_4_1_net3540), .RN(npu_inst_pe_1_4_1_n10), .Q(
        npu_inst_pe_1_4_1_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_4_1_n86), 
        .CK(npu_inst_pe_1_4_1_net3540), .RN(npu_inst_pe_1_4_1_n10), .Q(
        npu_inst_pe_1_4_1_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_4_1_n87), 
        .CK(npu_inst_pe_1_4_1_net3540), .RN(npu_inst_pe_1_4_1_n10), .Q(
        npu_inst_pe_1_4_1_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_4_1_n88), 
        .CK(npu_inst_pe_1_4_1_net3540), .RN(npu_inst_pe_1_4_1_n11), .Q(
        npu_inst_pe_1_4_1_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_4_1_n89), 
        .CK(npu_inst_pe_1_4_1_net3540), .RN(npu_inst_pe_1_4_1_n11), .Q(
        npu_inst_pe_1_4_1_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_4_1_n90), 
        .CK(npu_inst_pe_1_4_1_net3540), .RN(npu_inst_pe_1_4_1_n11), .Q(
        npu_inst_pe_1_4_1_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_4_1_n91), 
        .CK(npu_inst_pe_1_4_1_net3540), .RN(npu_inst_pe_1_4_1_n11), .Q(
        npu_inst_pe_1_4_1_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_4_1_n92), 
        .CK(npu_inst_pe_1_4_1_net3540), .RN(npu_inst_pe_1_4_1_n11), .Q(
        npu_inst_pe_1_4_1_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_4_1_n93), 
        .CK(npu_inst_pe_1_4_1_net3540), .RN(npu_inst_pe_1_4_1_n11), .Q(
        npu_inst_pe_1_4_1_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_4_1_n94), 
        .CK(npu_inst_pe_1_4_1_net3540), .RN(npu_inst_pe_1_4_1_n11), .Q(
        npu_inst_pe_1_4_1_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_4_1_n95), 
        .CK(npu_inst_pe_1_4_1_net3540), .RN(npu_inst_pe_1_4_1_n11), .Q(
        npu_inst_pe_1_4_1_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_4_1_n96), 
        .CK(npu_inst_pe_1_4_1_net3540), .RN(npu_inst_pe_1_4_1_n11), .Q(
        npu_inst_pe_1_4_1_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_4_1_n97), 
        .CK(npu_inst_pe_1_4_1_net3540), .RN(npu_inst_pe_1_4_1_n11), .Q(
        npu_inst_pe_1_4_1_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_4_1_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_4_1_N84), .SE(1'b0), .GCK(npu_inst_pe_1_4_1_net3534) );
  CLKGATETST_X1 npu_inst_pe_1_4_1_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n63), .SE(1'b0), .GCK(npu_inst_pe_1_4_1_net3540) );
  MUX2_X1 npu_inst_pe_1_4_2_U162 ( .A(npu_inst_pe_1_4_2_n32), .B(
        npu_inst_pe_1_4_2_n29), .S(npu_inst_pe_1_4_2_n8), .Z(
        npu_inst_pe_1_4_2_N93) );
  MUX2_X1 npu_inst_pe_1_4_2_U161 ( .A(npu_inst_pe_1_4_2_n31), .B(
        npu_inst_pe_1_4_2_n30), .S(npu_inst_pe_1_4_2_n6), .Z(
        npu_inst_pe_1_4_2_n32) );
  MUX2_X1 npu_inst_pe_1_4_2_U160 ( .A(npu_inst_pe_1_4_2_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_4_2_int_q_reg_v_1__0_), .S(npu_inst_pe_1_4_2_n4), .Z(
        npu_inst_pe_1_4_2_n31) );
  MUX2_X1 npu_inst_pe_1_4_2_U159 ( .A(npu_inst_pe_1_4_2_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_4_2_int_q_reg_v_3__0_), .S(npu_inst_pe_1_4_2_n4), .Z(
        npu_inst_pe_1_4_2_n30) );
  MUX2_X1 npu_inst_pe_1_4_2_U158 ( .A(npu_inst_pe_1_4_2_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_4_2_int_q_reg_v_5__0_), .S(npu_inst_pe_1_4_2_n4), .Z(
        npu_inst_pe_1_4_2_n29) );
  MUX2_X1 npu_inst_pe_1_4_2_U157 ( .A(npu_inst_pe_1_4_2_n28), .B(
        npu_inst_pe_1_4_2_n23), .S(npu_inst_pe_1_4_2_n8), .Z(
        npu_inst_pe_1_4_2_N94) );
  MUX2_X1 npu_inst_pe_1_4_2_U156 ( .A(npu_inst_pe_1_4_2_n25), .B(
        npu_inst_pe_1_4_2_n24), .S(npu_inst_pe_1_4_2_n6), .Z(
        npu_inst_pe_1_4_2_n28) );
  MUX2_X1 npu_inst_pe_1_4_2_U155 ( .A(npu_inst_pe_1_4_2_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_4_2_int_q_reg_v_1__1_), .S(npu_inst_pe_1_4_2_n4), .Z(
        npu_inst_pe_1_4_2_n25) );
  MUX2_X1 npu_inst_pe_1_4_2_U154 ( .A(npu_inst_pe_1_4_2_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_4_2_int_q_reg_v_3__1_), .S(npu_inst_pe_1_4_2_n4), .Z(
        npu_inst_pe_1_4_2_n24) );
  MUX2_X1 npu_inst_pe_1_4_2_U153 ( .A(npu_inst_pe_1_4_2_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_4_2_int_q_reg_v_5__1_), .S(npu_inst_pe_1_4_2_n4), .Z(
        npu_inst_pe_1_4_2_n23) );
  MUX2_X1 npu_inst_pe_1_4_2_U152 ( .A(npu_inst_pe_1_4_2_n22), .B(
        npu_inst_pe_1_4_2_n19), .S(npu_inst_pe_1_4_2_n8), .Z(
        npu_inst_int_data_x_4__2__1_) );
  MUX2_X1 npu_inst_pe_1_4_2_U151 ( .A(npu_inst_pe_1_4_2_n21), .B(
        npu_inst_pe_1_4_2_n20), .S(npu_inst_pe_1_4_2_n6), .Z(
        npu_inst_pe_1_4_2_n22) );
  MUX2_X1 npu_inst_pe_1_4_2_U150 ( .A(npu_inst_pe_1_4_2_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_4_2_int_q_reg_h_1__1_), .S(npu_inst_pe_1_4_2_n4), .Z(
        npu_inst_pe_1_4_2_n21) );
  MUX2_X1 npu_inst_pe_1_4_2_U149 ( .A(npu_inst_pe_1_4_2_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_4_2_int_q_reg_h_3__1_), .S(npu_inst_pe_1_4_2_n4), .Z(
        npu_inst_pe_1_4_2_n20) );
  MUX2_X1 npu_inst_pe_1_4_2_U148 ( .A(npu_inst_pe_1_4_2_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_4_2_int_q_reg_h_5__1_), .S(npu_inst_pe_1_4_2_n4), .Z(
        npu_inst_pe_1_4_2_n19) );
  MUX2_X1 npu_inst_pe_1_4_2_U147 ( .A(npu_inst_pe_1_4_2_n18), .B(
        npu_inst_pe_1_4_2_n15), .S(npu_inst_pe_1_4_2_n8), .Z(
        npu_inst_int_data_x_4__2__0_) );
  MUX2_X1 npu_inst_pe_1_4_2_U146 ( .A(npu_inst_pe_1_4_2_n17), .B(
        npu_inst_pe_1_4_2_n16), .S(npu_inst_pe_1_4_2_n6), .Z(
        npu_inst_pe_1_4_2_n18) );
  MUX2_X1 npu_inst_pe_1_4_2_U145 ( .A(npu_inst_pe_1_4_2_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_4_2_int_q_reg_h_1__0_), .S(npu_inst_pe_1_4_2_n4), .Z(
        npu_inst_pe_1_4_2_n17) );
  MUX2_X1 npu_inst_pe_1_4_2_U144 ( .A(npu_inst_pe_1_4_2_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_4_2_int_q_reg_h_3__0_), .S(npu_inst_pe_1_4_2_n4), .Z(
        npu_inst_pe_1_4_2_n16) );
  MUX2_X1 npu_inst_pe_1_4_2_U143 ( .A(npu_inst_pe_1_4_2_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_4_2_int_q_reg_h_5__0_), .S(npu_inst_pe_1_4_2_n4), .Z(
        npu_inst_pe_1_4_2_n15) );
  XOR2_X1 npu_inst_pe_1_4_2_U142 ( .A(npu_inst_pe_1_4_2_int_data_0_), .B(
        npu_inst_pe_1_4_2_int_q_acc_0_), .Z(npu_inst_pe_1_4_2_N73) );
  AND2_X1 npu_inst_pe_1_4_2_U141 ( .A1(npu_inst_pe_1_4_2_int_q_acc_0_), .A2(
        npu_inst_pe_1_4_2_int_data_0_), .ZN(npu_inst_pe_1_4_2_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_4_2_U140 ( .A(npu_inst_pe_1_4_2_int_q_acc_0_), .B(
        npu_inst_pe_1_4_2_n13), .ZN(npu_inst_pe_1_4_2_N65) );
  OR2_X1 npu_inst_pe_1_4_2_U139 ( .A1(npu_inst_pe_1_4_2_n13), .A2(
        npu_inst_pe_1_4_2_int_q_acc_0_), .ZN(npu_inst_pe_1_4_2_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_4_2_U138 ( .A(npu_inst_pe_1_4_2_int_q_acc_2_), .B(
        npu_inst_pe_1_4_2_add_79_carry_2_), .Z(npu_inst_pe_1_4_2_N75) );
  AND2_X1 npu_inst_pe_1_4_2_U137 ( .A1(npu_inst_pe_1_4_2_add_79_carry_2_), 
        .A2(npu_inst_pe_1_4_2_int_q_acc_2_), .ZN(
        npu_inst_pe_1_4_2_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_4_2_U136 ( .A(npu_inst_pe_1_4_2_int_q_acc_3_), .B(
        npu_inst_pe_1_4_2_add_79_carry_3_), .Z(npu_inst_pe_1_4_2_N76) );
  AND2_X1 npu_inst_pe_1_4_2_U135 ( .A1(npu_inst_pe_1_4_2_add_79_carry_3_), 
        .A2(npu_inst_pe_1_4_2_int_q_acc_3_), .ZN(
        npu_inst_pe_1_4_2_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_4_2_U134 ( .A(npu_inst_pe_1_4_2_int_q_acc_4_), .B(
        npu_inst_pe_1_4_2_add_79_carry_4_), .Z(npu_inst_pe_1_4_2_N77) );
  AND2_X1 npu_inst_pe_1_4_2_U133 ( .A1(npu_inst_pe_1_4_2_add_79_carry_4_), 
        .A2(npu_inst_pe_1_4_2_int_q_acc_4_), .ZN(
        npu_inst_pe_1_4_2_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_4_2_U132 ( .A(npu_inst_pe_1_4_2_int_q_acc_5_), .B(
        npu_inst_pe_1_4_2_add_79_carry_5_), .Z(npu_inst_pe_1_4_2_N78) );
  AND2_X1 npu_inst_pe_1_4_2_U131 ( .A1(npu_inst_pe_1_4_2_add_79_carry_5_), 
        .A2(npu_inst_pe_1_4_2_int_q_acc_5_), .ZN(
        npu_inst_pe_1_4_2_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_4_2_U130 ( .A(npu_inst_pe_1_4_2_int_q_acc_6_), .B(
        npu_inst_pe_1_4_2_add_79_carry_6_), .Z(npu_inst_pe_1_4_2_N79) );
  AND2_X1 npu_inst_pe_1_4_2_U129 ( .A1(npu_inst_pe_1_4_2_add_79_carry_6_), 
        .A2(npu_inst_pe_1_4_2_int_q_acc_6_), .ZN(
        npu_inst_pe_1_4_2_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_4_2_U128 ( .A(npu_inst_pe_1_4_2_int_q_acc_7_), .B(
        npu_inst_pe_1_4_2_add_79_carry_7_), .Z(npu_inst_pe_1_4_2_N80) );
  XNOR2_X1 npu_inst_pe_1_4_2_U127 ( .A(npu_inst_pe_1_4_2_sub_77_carry_2_), .B(
        npu_inst_pe_1_4_2_int_q_acc_2_), .ZN(npu_inst_pe_1_4_2_N67) );
  OR2_X1 npu_inst_pe_1_4_2_U126 ( .A1(npu_inst_pe_1_4_2_int_q_acc_2_), .A2(
        npu_inst_pe_1_4_2_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_4_2_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_4_2_U125 ( .A(npu_inst_pe_1_4_2_sub_77_carry_3_), .B(
        npu_inst_pe_1_4_2_int_q_acc_3_), .ZN(npu_inst_pe_1_4_2_N68) );
  OR2_X1 npu_inst_pe_1_4_2_U124 ( .A1(npu_inst_pe_1_4_2_int_q_acc_3_), .A2(
        npu_inst_pe_1_4_2_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_4_2_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_4_2_U123 ( .A(npu_inst_pe_1_4_2_sub_77_carry_4_), .B(
        npu_inst_pe_1_4_2_int_q_acc_4_), .ZN(npu_inst_pe_1_4_2_N69) );
  OR2_X1 npu_inst_pe_1_4_2_U122 ( .A1(npu_inst_pe_1_4_2_int_q_acc_4_), .A2(
        npu_inst_pe_1_4_2_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_4_2_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_4_2_U121 ( .A(npu_inst_pe_1_4_2_sub_77_carry_5_), .B(
        npu_inst_pe_1_4_2_int_q_acc_5_), .ZN(npu_inst_pe_1_4_2_N70) );
  OR2_X1 npu_inst_pe_1_4_2_U120 ( .A1(npu_inst_pe_1_4_2_int_q_acc_5_), .A2(
        npu_inst_pe_1_4_2_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_4_2_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_4_2_U119 ( .A(npu_inst_pe_1_4_2_sub_77_carry_6_), .B(
        npu_inst_pe_1_4_2_int_q_acc_6_), .ZN(npu_inst_pe_1_4_2_N71) );
  OR2_X1 npu_inst_pe_1_4_2_U118 ( .A1(npu_inst_pe_1_4_2_int_q_acc_6_), .A2(
        npu_inst_pe_1_4_2_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_4_2_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_4_2_U117 ( .A(npu_inst_pe_1_4_2_int_q_acc_7_), .B(
        npu_inst_pe_1_4_2_sub_77_carry_7_), .ZN(npu_inst_pe_1_4_2_N72) );
  INV_X1 npu_inst_pe_1_4_2_U116 ( .A(npu_inst_n77), .ZN(npu_inst_pe_1_4_2_n7)
         );
  INV_X1 npu_inst_pe_1_4_2_U115 ( .A(npu_inst_pe_1_4_2_n7), .ZN(
        npu_inst_pe_1_4_2_n6) );
  INV_X1 npu_inst_pe_1_4_2_U114 ( .A(npu_inst_n56), .ZN(npu_inst_pe_1_4_2_n3)
         );
  AOI22_X1 npu_inst_pe_1_4_2_U113 ( .A1(npu_inst_int_data_y_5__2__0_), .A2(
        npu_inst_pe_1_4_2_n58), .B1(npu_inst_pe_1_4_2_n114), .B2(
        npu_inst_pe_1_4_2_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_4_2_n57) );
  INV_X1 npu_inst_pe_1_4_2_U112 ( .A(npu_inst_pe_1_4_2_n57), .ZN(
        npu_inst_pe_1_4_2_n108) );
  AOI22_X1 npu_inst_pe_1_4_2_U111 ( .A1(npu_inst_int_data_y_5__2__0_), .A2(
        npu_inst_pe_1_4_2_n54), .B1(npu_inst_pe_1_4_2_n115), .B2(
        npu_inst_pe_1_4_2_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_4_2_n53) );
  INV_X1 npu_inst_pe_1_4_2_U110 ( .A(npu_inst_pe_1_4_2_n53), .ZN(
        npu_inst_pe_1_4_2_n109) );
  AOI22_X1 npu_inst_pe_1_4_2_U107 ( .A1(npu_inst_int_data_y_5__2__0_), .A2(
        npu_inst_pe_1_4_2_n50), .B1(npu_inst_pe_1_4_2_n116), .B2(
        npu_inst_pe_1_4_2_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_4_2_n49) );
  INV_X1 npu_inst_pe_1_4_2_U106 ( .A(npu_inst_pe_1_4_2_n49), .ZN(
        npu_inst_pe_1_4_2_n110) );
  AOI22_X1 npu_inst_pe_1_4_2_U105 ( .A1(npu_inst_int_data_y_5__2__0_), .A2(
        npu_inst_pe_1_4_2_n46), .B1(npu_inst_pe_1_4_2_n117), .B2(
        npu_inst_pe_1_4_2_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_4_2_n45) );
  INV_X1 npu_inst_pe_1_4_2_U104 ( .A(npu_inst_pe_1_4_2_n45), .ZN(
        npu_inst_pe_1_4_2_n111) );
  AOI22_X1 npu_inst_pe_1_4_2_U103 ( .A1(npu_inst_int_data_y_5__2__0_), .A2(
        npu_inst_pe_1_4_2_n42), .B1(npu_inst_pe_1_4_2_n119), .B2(
        npu_inst_pe_1_4_2_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_4_2_n41) );
  INV_X1 npu_inst_pe_1_4_2_U102 ( .A(npu_inst_pe_1_4_2_n41), .ZN(
        npu_inst_pe_1_4_2_n112) );
  AOI22_X1 npu_inst_pe_1_4_2_U101 ( .A1(npu_inst_int_data_y_5__2__1_), .A2(
        npu_inst_pe_1_4_2_n58), .B1(npu_inst_pe_1_4_2_n114), .B2(
        npu_inst_pe_1_4_2_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_4_2_n59) );
  INV_X1 npu_inst_pe_1_4_2_U100 ( .A(npu_inst_pe_1_4_2_n59), .ZN(
        npu_inst_pe_1_4_2_n102) );
  AOI22_X1 npu_inst_pe_1_4_2_U99 ( .A1(npu_inst_int_data_y_5__2__1_), .A2(
        npu_inst_pe_1_4_2_n54), .B1(npu_inst_pe_1_4_2_n115), .B2(
        npu_inst_pe_1_4_2_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_4_2_n55) );
  INV_X1 npu_inst_pe_1_4_2_U98 ( .A(npu_inst_pe_1_4_2_n55), .ZN(
        npu_inst_pe_1_4_2_n103) );
  AOI22_X1 npu_inst_pe_1_4_2_U97 ( .A1(npu_inst_int_data_y_5__2__1_), .A2(
        npu_inst_pe_1_4_2_n50), .B1(npu_inst_pe_1_4_2_n116), .B2(
        npu_inst_pe_1_4_2_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_4_2_n51) );
  INV_X1 npu_inst_pe_1_4_2_U96 ( .A(npu_inst_pe_1_4_2_n51), .ZN(
        npu_inst_pe_1_4_2_n104) );
  AOI22_X1 npu_inst_pe_1_4_2_U95 ( .A1(npu_inst_int_data_y_5__2__1_), .A2(
        npu_inst_pe_1_4_2_n46), .B1(npu_inst_pe_1_4_2_n117), .B2(
        npu_inst_pe_1_4_2_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_4_2_n47) );
  INV_X1 npu_inst_pe_1_4_2_U94 ( .A(npu_inst_pe_1_4_2_n47), .ZN(
        npu_inst_pe_1_4_2_n105) );
  AOI22_X1 npu_inst_pe_1_4_2_U93 ( .A1(npu_inst_int_data_y_5__2__1_), .A2(
        npu_inst_pe_1_4_2_n42), .B1(npu_inst_pe_1_4_2_n119), .B2(
        npu_inst_pe_1_4_2_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_4_2_n43) );
  INV_X1 npu_inst_pe_1_4_2_U92 ( .A(npu_inst_pe_1_4_2_n43), .ZN(
        npu_inst_pe_1_4_2_n106) );
  AOI22_X1 npu_inst_pe_1_4_2_U91 ( .A1(npu_inst_pe_1_4_2_n38), .A2(
        npu_inst_int_data_y_5__2__1_), .B1(npu_inst_pe_1_4_2_n118), .B2(
        npu_inst_pe_1_4_2_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_4_2_n39) );
  INV_X1 npu_inst_pe_1_4_2_U90 ( .A(npu_inst_pe_1_4_2_n39), .ZN(
        npu_inst_pe_1_4_2_n107) );
  AOI22_X1 npu_inst_pe_1_4_2_U89 ( .A1(npu_inst_pe_1_4_2_n38), .A2(
        npu_inst_int_data_y_5__2__0_), .B1(npu_inst_pe_1_4_2_n118), .B2(
        npu_inst_pe_1_4_2_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_4_2_n37) );
  INV_X1 npu_inst_pe_1_4_2_U88 ( .A(npu_inst_pe_1_4_2_n37), .ZN(
        npu_inst_pe_1_4_2_n113) );
  NAND2_X1 npu_inst_pe_1_4_2_U87 ( .A1(npu_inst_pe_1_4_2_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_4_2_n60), .ZN(npu_inst_pe_1_4_2_n74) );
  OAI21_X1 npu_inst_pe_1_4_2_U86 ( .B1(npu_inst_pe_1_4_2_n63), .B2(
        npu_inst_pe_1_4_2_n60), .A(npu_inst_pe_1_4_2_n74), .ZN(
        npu_inst_pe_1_4_2_n97) );
  NAND2_X1 npu_inst_pe_1_4_2_U85 ( .A1(npu_inst_pe_1_4_2_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_4_2_n60), .ZN(npu_inst_pe_1_4_2_n73) );
  OAI21_X1 npu_inst_pe_1_4_2_U84 ( .B1(npu_inst_pe_1_4_2_n61), .B2(
        npu_inst_pe_1_4_2_n60), .A(npu_inst_pe_1_4_2_n73), .ZN(
        npu_inst_pe_1_4_2_n96) );
  NAND2_X1 npu_inst_pe_1_4_2_U83 ( .A1(npu_inst_pe_1_4_2_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_4_2_n56), .ZN(npu_inst_pe_1_4_2_n72) );
  OAI21_X1 npu_inst_pe_1_4_2_U82 ( .B1(npu_inst_pe_1_4_2_n63), .B2(
        npu_inst_pe_1_4_2_n56), .A(npu_inst_pe_1_4_2_n72), .ZN(
        npu_inst_pe_1_4_2_n95) );
  NAND2_X1 npu_inst_pe_1_4_2_U81 ( .A1(npu_inst_pe_1_4_2_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_4_2_n56), .ZN(npu_inst_pe_1_4_2_n71) );
  OAI21_X1 npu_inst_pe_1_4_2_U80 ( .B1(npu_inst_pe_1_4_2_n61), .B2(
        npu_inst_pe_1_4_2_n56), .A(npu_inst_pe_1_4_2_n71), .ZN(
        npu_inst_pe_1_4_2_n94) );
  NAND2_X1 npu_inst_pe_1_4_2_U79 ( .A1(npu_inst_pe_1_4_2_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_4_2_n52), .ZN(npu_inst_pe_1_4_2_n70) );
  OAI21_X1 npu_inst_pe_1_4_2_U78 ( .B1(npu_inst_pe_1_4_2_n63), .B2(
        npu_inst_pe_1_4_2_n52), .A(npu_inst_pe_1_4_2_n70), .ZN(
        npu_inst_pe_1_4_2_n93) );
  NAND2_X1 npu_inst_pe_1_4_2_U77 ( .A1(npu_inst_pe_1_4_2_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_4_2_n52), .ZN(npu_inst_pe_1_4_2_n69) );
  OAI21_X1 npu_inst_pe_1_4_2_U76 ( .B1(npu_inst_pe_1_4_2_n61), .B2(
        npu_inst_pe_1_4_2_n52), .A(npu_inst_pe_1_4_2_n69), .ZN(
        npu_inst_pe_1_4_2_n92) );
  NAND2_X1 npu_inst_pe_1_4_2_U75 ( .A1(npu_inst_pe_1_4_2_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_4_2_n48), .ZN(npu_inst_pe_1_4_2_n68) );
  OAI21_X1 npu_inst_pe_1_4_2_U74 ( .B1(npu_inst_pe_1_4_2_n63), .B2(
        npu_inst_pe_1_4_2_n48), .A(npu_inst_pe_1_4_2_n68), .ZN(
        npu_inst_pe_1_4_2_n91) );
  NAND2_X1 npu_inst_pe_1_4_2_U73 ( .A1(npu_inst_pe_1_4_2_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_4_2_n48), .ZN(npu_inst_pe_1_4_2_n67) );
  OAI21_X1 npu_inst_pe_1_4_2_U72 ( .B1(npu_inst_pe_1_4_2_n61), .B2(
        npu_inst_pe_1_4_2_n48), .A(npu_inst_pe_1_4_2_n67), .ZN(
        npu_inst_pe_1_4_2_n90) );
  NAND2_X1 npu_inst_pe_1_4_2_U71 ( .A1(npu_inst_pe_1_4_2_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_4_2_n44), .ZN(npu_inst_pe_1_4_2_n66) );
  OAI21_X1 npu_inst_pe_1_4_2_U70 ( .B1(npu_inst_pe_1_4_2_n63), .B2(
        npu_inst_pe_1_4_2_n44), .A(npu_inst_pe_1_4_2_n66), .ZN(
        npu_inst_pe_1_4_2_n89) );
  NAND2_X1 npu_inst_pe_1_4_2_U69 ( .A1(npu_inst_pe_1_4_2_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_4_2_n44), .ZN(npu_inst_pe_1_4_2_n65) );
  OAI21_X1 npu_inst_pe_1_4_2_U68 ( .B1(npu_inst_pe_1_4_2_n61), .B2(
        npu_inst_pe_1_4_2_n44), .A(npu_inst_pe_1_4_2_n65), .ZN(
        npu_inst_pe_1_4_2_n88) );
  NAND2_X1 npu_inst_pe_1_4_2_U67 ( .A1(npu_inst_pe_1_4_2_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_4_2_n40), .ZN(npu_inst_pe_1_4_2_n64) );
  OAI21_X1 npu_inst_pe_1_4_2_U66 ( .B1(npu_inst_pe_1_4_2_n63), .B2(
        npu_inst_pe_1_4_2_n40), .A(npu_inst_pe_1_4_2_n64), .ZN(
        npu_inst_pe_1_4_2_n87) );
  NAND2_X1 npu_inst_pe_1_4_2_U65 ( .A1(npu_inst_pe_1_4_2_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_4_2_n40), .ZN(npu_inst_pe_1_4_2_n62) );
  OAI21_X1 npu_inst_pe_1_4_2_U64 ( .B1(npu_inst_pe_1_4_2_n61), .B2(
        npu_inst_pe_1_4_2_n40), .A(npu_inst_pe_1_4_2_n62), .ZN(
        npu_inst_pe_1_4_2_n86) );
  AND2_X1 npu_inst_pe_1_4_2_U63 ( .A1(npu_inst_pe_1_4_2_N93), .A2(npu_inst_n56), .ZN(npu_inst_int_data_y_4__2__0_) );
  AND2_X1 npu_inst_pe_1_4_2_U62 ( .A1(npu_inst_n56), .A2(npu_inst_pe_1_4_2_N94), .ZN(npu_inst_int_data_y_4__2__1_) );
  NOR3_X1 npu_inst_pe_1_4_2_U61 ( .A1(npu_inst_pe_1_4_2_n26), .A2(npu_inst_n56), .A3(npu_inst_int_ckg[29]), .ZN(npu_inst_pe_1_4_2_n85) );
  OR2_X1 npu_inst_pe_1_4_2_U60 ( .A1(npu_inst_pe_1_4_2_n85), .A2(
        npu_inst_pe_1_4_2_n2), .ZN(npu_inst_pe_1_4_2_N84) );
  AND2_X1 npu_inst_pe_1_4_2_U59 ( .A1(npu_inst_pe_1_4_2_int_q_acc_0_), .A2(
        npu_inst_pe_1_4_2_n1), .ZN(npu_inst_int_data_res_4__2__0_) );
  AND2_X1 npu_inst_pe_1_4_2_U58 ( .A1(npu_inst_pe_1_4_2_n2), .A2(
        npu_inst_pe_1_4_2_int_q_acc_7_), .ZN(npu_inst_int_data_res_4__2__7_)
         );
  AND2_X1 npu_inst_pe_1_4_2_U57 ( .A1(npu_inst_pe_1_4_2_int_q_acc_1_), .A2(
        npu_inst_pe_1_4_2_n1), .ZN(npu_inst_int_data_res_4__2__1_) );
  AND2_X1 npu_inst_pe_1_4_2_U56 ( .A1(npu_inst_pe_1_4_2_int_q_acc_2_), .A2(
        npu_inst_pe_1_4_2_n1), .ZN(npu_inst_int_data_res_4__2__2_) );
  AND2_X1 npu_inst_pe_1_4_2_U55 ( .A1(npu_inst_pe_1_4_2_int_q_acc_3_), .A2(
        npu_inst_pe_1_4_2_n2), .ZN(npu_inst_int_data_res_4__2__3_) );
  AND2_X1 npu_inst_pe_1_4_2_U54 ( .A1(npu_inst_pe_1_4_2_int_q_acc_4_), .A2(
        npu_inst_pe_1_4_2_n2), .ZN(npu_inst_int_data_res_4__2__4_) );
  AND2_X1 npu_inst_pe_1_4_2_U53 ( .A1(npu_inst_pe_1_4_2_int_q_acc_5_), .A2(
        npu_inst_pe_1_4_2_n2), .ZN(npu_inst_int_data_res_4__2__5_) );
  AND2_X1 npu_inst_pe_1_4_2_U52 ( .A1(npu_inst_pe_1_4_2_int_q_acc_6_), .A2(
        npu_inst_pe_1_4_2_n2), .ZN(npu_inst_int_data_res_4__2__6_) );
  AOI222_X1 npu_inst_pe_1_4_2_U51 ( .A1(npu_inst_int_data_res_5__2__0_), .A2(
        npu_inst_pe_1_4_2_n1), .B1(npu_inst_pe_1_4_2_N73), .B2(
        npu_inst_pe_1_4_2_n76), .C1(npu_inst_pe_1_4_2_N65), .C2(
        npu_inst_pe_1_4_2_n77), .ZN(npu_inst_pe_1_4_2_n84) );
  INV_X1 npu_inst_pe_1_4_2_U50 ( .A(npu_inst_pe_1_4_2_n84), .ZN(
        npu_inst_pe_1_4_2_n101) );
  AOI222_X1 npu_inst_pe_1_4_2_U49 ( .A1(npu_inst_int_data_res_5__2__7_), .A2(
        npu_inst_pe_1_4_2_n1), .B1(npu_inst_pe_1_4_2_N80), .B2(
        npu_inst_pe_1_4_2_n76), .C1(npu_inst_pe_1_4_2_N72), .C2(
        npu_inst_pe_1_4_2_n77), .ZN(npu_inst_pe_1_4_2_n75) );
  INV_X1 npu_inst_pe_1_4_2_U48 ( .A(npu_inst_pe_1_4_2_n75), .ZN(
        npu_inst_pe_1_4_2_n33) );
  AOI222_X1 npu_inst_pe_1_4_2_U47 ( .A1(npu_inst_int_data_res_5__2__1_), .A2(
        npu_inst_pe_1_4_2_n1), .B1(npu_inst_pe_1_4_2_N74), .B2(
        npu_inst_pe_1_4_2_n76), .C1(npu_inst_pe_1_4_2_N66), .C2(
        npu_inst_pe_1_4_2_n77), .ZN(npu_inst_pe_1_4_2_n83) );
  INV_X1 npu_inst_pe_1_4_2_U46 ( .A(npu_inst_pe_1_4_2_n83), .ZN(
        npu_inst_pe_1_4_2_n100) );
  AOI222_X1 npu_inst_pe_1_4_2_U45 ( .A1(npu_inst_int_data_res_5__2__2_), .A2(
        npu_inst_pe_1_4_2_n1), .B1(npu_inst_pe_1_4_2_N75), .B2(
        npu_inst_pe_1_4_2_n76), .C1(npu_inst_pe_1_4_2_N67), .C2(
        npu_inst_pe_1_4_2_n77), .ZN(npu_inst_pe_1_4_2_n82) );
  INV_X1 npu_inst_pe_1_4_2_U44 ( .A(npu_inst_pe_1_4_2_n82), .ZN(
        npu_inst_pe_1_4_2_n99) );
  AOI222_X1 npu_inst_pe_1_4_2_U43 ( .A1(npu_inst_int_data_res_5__2__3_), .A2(
        npu_inst_pe_1_4_2_n1), .B1(npu_inst_pe_1_4_2_N76), .B2(
        npu_inst_pe_1_4_2_n76), .C1(npu_inst_pe_1_4_2_N68), .C2(
        npu_inst_pe_1_4_2_n77), .ZN(npu_inst_pe_1_4_2_n81) );
  INV_X1 npu_inst_pe_1_4_2_U42 ( .A(npu_inst_pe_1_4_2_n81), .ZN(
        npu_inst_pe_1_4_2_n98) );
  AOI222_X1 npu_inst_pe_1_4_2_U41 ( .A1(npu_inst_int_data_res_5__2__4_), .A2(
        npu_inst_pe_1_4_2_n1), .B1(npu_inst_pe_1_4_2_N77), .B2(
        npu_inst_pe_1_4_2_n76), .C1(npu_inst_pe_1_4_2_N69), .C2(
        npu_inst_pe_1_4_2_n77), .ZN(npu_inst_pe_1_4_2_n80) );
  INV_X1 npu_inst_pe_1_4_2_U40 ( .A(npu_inst_pe_1_4_2_n80), .ZN(
        npu_inst_pe_1_4_2_n36) );
  AOI222_X1 npu_inst_pe_1_4_2_U39 ( .A1(npu_inst_int_data_res_5__2__5_), .A2(
        npu_inst_pe_1_4_2_n1), .B1(npu_inst_pe_1_4_2_N78), .B2(
        npu_inst_pe_1_4_2_n76), .C1(npu_inst_pe_1_4_2_N70), .C2(
        npu_inst_pe_1_4_2_n77), .ZN(npu_inst_pe_1_4_2_n79) );
  INV_X1 npu_inst_pe_1_4_2_U38 ( .A(npu_inst_pe_1_4_2_n79), .ZN(
        npu_inst_pe_1_4_2_n35) );
  AOI222_X1 npu_inst_pe_1_4_2_U37 ( .A1(npu_inst_int_data_res_5__2__6_), .A2(
        npu_inst_pe_1_4_2_n1), .B1(npu_inst_pe_1_4_2_N79), .B2(
        npu_inst_pe_1_4_2_n76), .C1(npu_inst_pe_1_4_2_N71), .C2(
        npu_inst_pe_1_4_2_n77), .ZN(npu_inst_pe_1_4_2_n78) );
  INV_X1 npu_inst_pe_1_4_2_U36 ( .A(npu_inst_pe_1_4_2_n78), .ZN(
        npu_inst_pe_1_4_2_n34) );
  INV_X1 npu_inst_pe_1_4_2_U35 ( .A(npu_inst_pe_1_4_2_int_data_1_), .ZN(
        npu_inst_pe_1_4_2_n14) );
  AND2_X1 npu_inst_pe_1_4_2_U34 ( .A1(npu_inst_int_data_x_4__2__1_), .A2(
        npu_inst_pe_1_4_2_int_q_weight_1_), .ZN(npu_inst_pe_1_4_2_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_4_2_U33 ( .A1(npu_inst_int_data_x_4__2__0_), .A2(
        npu_inst_pe_1_4_2_int_q_weight_1_), .ZN(npu_inst_pe_1_4_2_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_4_2_U32 ( .A1(npu_inst_n56), .A2(
        npu_inst_int_data_y_5__2__1_), .B1(npu_inst_pe_1_4_2_n3), .B2(
        npu_inst_int_data_x_4__3__1_), .ZN(npu_inst_pe_1_4_2_n63) );
  AOI22_X1 npu_inst_pe_1_4_2_U31 ( .A1(npu_inst_n56), .A2(
        npu_inst_int_data_y_5__2__0_), .B1(npu_inst_pe_1_4_2_n3), .B2(
        npu_inst_int_data_x_4__3__0_), .ZN(npu_inst_pe_1_4_2_n61) );
  INV_X1 npu_inst_pe_1_4_2_U30 ( .A(npu_inst_pe_1_4_2_int_data_0_), .ZN(
        npu_inst_pe_1_4_2_n13) );
  INV_X1 npu_inst_pe_1_4_2_U29 ( .A(npu_inst_n69), .ZN(npu_inst_pe_1_4_2_n5)
         );
  OR3_X1 npu_inst_pe_1_4_2_U28 ( .A1(npu_inst_pe_1_4_2_n6), .A2(
        npu_inst_pe_1_4_2_n8), .A3(npu_inst_pe_1_4_2_n5), .ZN(
        npu_inst_pe_1_4_2_n56) );
  OR3_X1 npu_inst_pe_1_4_2_U27 ( .A1(npu_inst_pe_1_4_2_n5), .A2(
        npu_inst_pe_1_4_2_n8), .A3(npu_inst_pe_1_4_2_n7), .ZN(
        npu_inst_pe_1_4_2_n48) );
  INV_X1 npu_inst_pe_1_4_2_U26 ( .A(npu_inst_pe_1_4_2_n5), .ZN(
        npu_inst_pe_1_4_2_n4) );
  INV_X1 npu_inst_pe_1_4_2_U25 ( .A(npu_inst_n124), .ZN(npu_inst_pe_1_4_2_n12)
         );
  OR3_X1 npu_inst_pe_1_4_2_U24 ( .A1(npu_inst_pe_1_4_2_n4), .A2(
        npu_inst_pe_1_4_2_n8), .A3(npu_inst_pe_1_4_2_n7), .ZN(
        npu_inst_pe_1_4_2_n52) );
  OR3_X1 npu_inst_pe_1_4_2_U23 ( .A1(npu_inst_pe_1_4_2_n6), .A2(
        npu_inst_pe_1_4_2_n8), .A3(npu_inst_pe_1_4_2_n4), .ZN(
        npu_inst_pe_1_4_2_n60) );
  NOR2_X1 npu_inst_pe_1_4_2_U22 ( .A1(npu_inst_pe_1_4_2_n60), .A2(
        npu_inst_pe_1_4_2_n3), .ZN(npu_inst_pe_1_4_2_n58) );
  NOR2_X1 npu_inst_pe_1_4_2_U21 ( .A1(npu_inst_pe_1_4_2_n56), .A2(
        npu_inst_pe_1_4_2_n3), .ZN(npu_inst_pe_1_4_2_n54) );
  NOR2_X1 npu_inst_pe_1_4_2_U20 ( .A1(npu_inst_pe_1_4_2_n52), .A2(
        npu_inst_pe_1_4_2_n3), .ZN(npu_inst_pe_1_4_2_n50) );
  NOR2_X1 npu_inst_pe_1_4_2_U19 ( .A1(npu_inst_pe_1_4_2_n48), .A2(
        npu_inst_pe_1_4_2_n3), .ZN(npu_inst_pe_1_4_2_n46) );
  NOR2_X1 npu_inst_pe_1_4_2_U18 ( .A1(npu_inst_pe_1_4_2_n40), .A2(
        npu_inst_pe_1_4_2_n3), .ZN(npu_inst_pe_1_4_2_n38) );
  NOR2_X1 npu_inst_pe_1_4_2_U17 ( .A1(npu_inst_pe_1_4_2_n44), .A2(
        npu_inst_pe_1_4_2_n3), .ZN(npu_inst_pe_1_4_2_n42) );
  BUF_X1 npu_inst_pe_1_4_2_U16 ( .A(npu_inst_n99), .Z(npu_inst_pe_1_4_2_n8) );
  BUF_X1 npu_inst_pe_1_4_2_U15 ( .A(npu_inst_pe_1_4_2_n12), .Z(
        npu_inst_pe_1_4_2_n11) );
  BUF_X1 npu_inst_pe_1_4_2_U14 ( .A(npu_inst_pe_1_4_2_n12), .Z(
        npu_inst_pe_1_4_2_n10) );
  BUF_X1 npu_inst_pe_1_4_2_U13 ( .A(npu_inst_pe_1_4_2_n12), .Z(
        npu_inst_pe_1_4_2_n9) );
  INV_X1 npu_inst_pe_1_4_2_U12 ( .A(npu_inst_pe_1_4_2_n38), .ZN(
        npu_inst_pe_1_4_2_n118) );
  INV_X1 npu_inst_pe_1_4_2_U11 ( .A(npu_inst_pe_1_4_2_n58), .ZN(
        npu_inst_pe_1_4_2_n114) );
  INV_X1 npu_inst_pe_1_4_2_U10 ( .A(npu_inst_pe_1_4_2_n54), .ZN(
        npu_inst_pe_1_4_2_n115) );
  INV_X1 npu_inst_pe_1_4_2_U9 ( .A(npu_inst_pe_1_4_2_n50), .ZN(
        npu_inst_pe_1_4_2_n116) );
  INV_X1 npu_inst_pe_1_4_2_U8 ( .A(npu_inst_pe_1_4_2_n46), .ZN(
        npu_inst_pe_1_4_2_n117) );
  INV_X1 npu_inst_pe_1_4_2_U7 ( .A(npu_inst_pe_1_4_2_n42), .ZN(
        npu_inst_pe_1_4_2_n119) );
  BUF_X1 npu_inst_pe_1_4_2_U6 ( .A(npu_inst_n21), .Z(npu_inst_pe_1_4_2_n2) );
  BUF_X1 npu_inst_pe_1_4_2_U5 ( .A(npu_inst_n21), .Z(npu_inst_pe_1_4_2_n1) );
  NOR2_X1 npu_inst_pe_1_4_2_U4 ( .A1(npu_inst_pe_1_4_2_int_q_weight_0_), .A2(
        npu_inst_pe_1_4_2_n1), .ZN(npu_inst_pe_1_4_2_n76) );
  NOR2_X1 npu_inst_pe_1_4_2_U3 ( .A1(npu_inst_pe_1_4_2_n27), .A2(
        npu_inst_pe_1_4_2_n1), .ZN(npu_inst_pe_1_4_2_n77) );
  FA_X1 npu_inst_pe_1_4_2_sub_77_U2_1 ( .A(npu_inst_pe_1_4_2_int_q_acc_1_), 
        .B(npu_inst_pe_1_4_2_n14), .CI(npu_inst_pe_1_4_2_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_4_2_sub_77_carry_2_), .S(npu_inst_pe_1_4_2_N66) );
  FA_X1 npu_inst_pe_1_4_2_add_79_U1_1 ( .A(npu_inst_pe_1_4_2_int_q_acc_1_), 
        .B(npu_inst_pe_1_4_2_int_data_1_), .CI(
        npu_inst_pe_1_4_2_add_79_carry_1_), .CO(
        npu_inst_pe_1_4_2_add_79_carry_2_), .S(npu_inst_pe_1_4_2_N74) );
  NAND3_X1 npu_inst_pe_1_4_2_U109 ( .A1(npu_inst_pe_1_4_2_n5), .A2(
        npu_inst_pe_1_4_2_n7), .A3(npu_inst_pe_1_4_2_n8), .ZN(
        npu_inst_pe_1_4_2_n44) );
  NAND3_X1 npu_inst_pe_1_4_2_U108 ( .A1(npu_inst_pe_1_4_2_n4), .A2(
        npu_inst_pe_1_4_2_n7), .A3(npu_inst_pe_1_4_2_n8), .ZN(
        npu_inst_pe_1_4_2_n40) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_4_2_n34), .CK(
        npu_inst_pe_1_4_2_net3511), .RN(npu_inst_pe_1_4_2_n9), .Q(
        npu_inst_pe_1_4_2_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_4_2_n35), .CK(
        npu_inst_pe_1_4_2_net3511), .RN(npu_inst_pe_1_4_2_n9), .Q(
        npu_inst_pe_1_4_2_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_4_2_n36), .CK(
        npu_inst_pe_1_4_2_net3511), .RN(npu_inst_pe_1_4_2_n9), .Q(
        npu_inst_pe_1_4_2_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_4_2_n98), .CK(
        npu_inst_pe_1_4_2_net3511), .RN(npu_inst_pe_1_4_2_n9), .Q(
        npu_inst_pe_1_4_2_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_4_2_n99), .CK(
        npu_inst_pe_1_4_2_net3511), .RN(npu_inst_pe_1_4_2_n9), .Q(
        npu_inst_pe_1_4_2_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_4_2_n100), 
        .CK(npu_inst_pe_1_4_2_net3511), .RN(npu_inst_pe_1_4_2_n9), .Q(
        npu_inst_pe_1_4_2_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_4_2_n33), .CK(
        npu_inst_pe_1_4_2_net3511), .RN(npu_inst_pe_1_4_2_n9), .Q(
        npu_inst_pe_1_4_2_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_4_2_n101), 
        .CK(npu_inst_pe_1_4_2_net3511), .RN(npu_inst_pe_1_4_2_n9), .Q(
        npu_inst_pe_1_4_2_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_weight_reg_0_ ( .D(npu_inst_n110), .CK(
        npu_inst_pe_1_4_2_net3517), .RN(npu_inst_pe_1_4_2_n9), .Q(
        npu_inst_pe_1_4_2_int_q_weight_0_), .QN(npu_inst_pe_1_4_2_n27) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_weight_reg_1_ ( .D(npu_inst_n116), .CK(
        npu_inst_pe_1_4_2_net3517), .RN(npu_inst_pe_1_4_2_n9), .Q(
        npu_inst_pe_1_4_2_int_q_weight_1_), .QN(npu_inst_pe_1_4_2_n26) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_4_2_n113), 
        .CK(npu_inst_pe_1_4_2_net3517), .RN(npu_inst_pe_1_4_2_n9), .Q(
        npu_inst_pe_1_4_2_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_4_2_n107), 
        .CK(npu_inst_pe_1_4_2_net3517), .RN(npu_inst_pe_1_4_2_n9), .Q(
        npu_inst_pe_1_4_2_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_4_2_n112), 
        .CK(npu_inst_pe_1_4_2_net3517), .RN(npu_inst_pe_1_4_2_n10), .Q(
        npu_inst_pe_1_4_2_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_4_2_n106), 
        .CK(npu_inst_pe_1_4_2_net3517), .RN(npu_inst_pe_1_4_2_n10), .Q(
        npu_inst_pe_1_4_2_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_4_2_n111), 
        .CK(npu_inst_pe_1_4_2_net3517), .RN(npu_inst_pe_1_4_2_n10), .Q(
        npu_inst_pe_1_4_2_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_4_2_n105), 
        .CK(npu_inst_pe_1_4_2_net3517), .RN(npu_inst_pe_1_4_2_n10), .Q(
        npu_inst_pe_1_4_2_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_4_2_n110), 
        .CK(npu_inst_pe_1_4_2_net3517), .RN(npu_inst_pe_1_4_2_n10), .Q(
        npu_inst_pe_1_4_2_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_4_2_n104), 
        .CK(npu_inst_pe_1_4_2_net3517), .RN(npu_inst_pe_1_4_2_n10), .Q(
        npu_inst_pe_1_4_2_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_4_2_n109), 
        .CK(npu_inst_pe_1_4_2_net3517), .RN(npu_inst_pe_1_4_2_n10), .Q(
        npu_inst_pe_1_4_2_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_4_2_n103), 
        .CK(npu_inst_pe_1_4_2_net3517), .RN(npu_inst_pe_1_4_2_n10), .Q(
        npu_inst_pe_1_4_2_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_4_2_n108), 
        .CK(npu_inst_pe_1_4_2_net3517), .RN(npu_inst_pe_1_4_2_n10), .Q(
        npu_inst_pe_1_4_2_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_4_2_n102), 
        .CK(npu_inst_pe_1_4_2_net3517), .RN(npu_inst_pe_1_4_2_n10), .Q(
        npu_inst_pe_1_4_2_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_4_2_n86), 
        .CK(npu_inst_pe_1_4_2_net3517), .RN(npu_inst_pe_1_4_2_n10), .Q(
        npu_inst_pe_1_4_2_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_4_2_n87), 
        .CK(npu_inst_pe_1_4_2_net3517), .RN(npu_inst_pe_1_4_2_n10), .Q(
        npu_inst_pe_1_4_2_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_4_2_n88), 
        .CK(npu_inst_pe_1_4_2_net3517), .RN(npu_inst_pe_1_4_2_n11), .Q(
        npu_inst_pe_1_4_2_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_4_2_n89), 
        .CK(npu_inst_pe_1_4_2_net3517), .RN(npu_inst_pe_1_4_2_n11), .Q(
        npu_inst_pe_1_4_2_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_4_2_n90), 
        .CK(npu_inst_pe_1_4_2_net3517), .RN(npu_inst_pe_1_4_2_n11), .Q(
        npu_inst_pe_1_4_2_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_4_2_n91), 
        .CK(npu_inst_pe_1_4_2_net3517), .RN(npu_inst_pe_1_4_2_n11), .Q(
        npu_inst_pe_1_4_2_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_4_2_n92), 
        .CK(npu_inst_pe_1_4_2_net3517), .RN(npu_inst_pe_1_4_2_n11), .Q(
        npu_inst_pe_1_4_2_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_4_2_n93), 
        .CK(npu_inst_pe_1_4_2_net3517), .RN(npu_inst_pe_1_4_2_n11), .Q(
        npu_inst_pe_1_4_2_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_4_2_n94), 
        .CK(npu_inst_pe_1_4_2_net3517), .RN(npu_inst_pe_1_4_2_n11), .Q(
        npu_inst_pe_1_4_2_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_4_2_n95), 
        .CK(npu_inst_pe_1_4_2_net3517), .RN(npu_inst_pe_1_4_2_n11), .Q(
        npu_inst_pe_1_4_2_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_4_2_n96), 
        .CK(npu_inst_pe_1_4_2_net3517), .RN(npu_inst_pe_1_4_2_n11), .Q(
        npu_inst_pe_1_4_2_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_4_2_n97), 
        .CK(npu_inst_pe_1_4_2_net3517), .RN(npu_inst_pe_1_4_2_n11), .Q(
        npu_inst_pe_1_4_2_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_4_2_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_4_2_N84), .SE(1'b0), .GCK(npu_inst_pe_1_4_2_net3511) );
  CLKGATETST_X1 npu_inst_pe_1_4_2_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n63), .SE(1'b0), .GCK(npu_inst_pe_1_4_2_net3517) );
  MUX2_X1 npu_inst_pe_1_4_3_U162 ( .A(npu_inst_pe_1_4_3_n32), .B(
        npu_inst_pe_1_4_3_n29), .S(npu_inst_pe_1_4_3_n8), .Z(
        npu_inst_pe_1_4_3_N93) );
  MUX2_X1 npu_inst_pe_1_4_3_U161 ( .A(npu_inst_pe_1_4_3_n31), .B(
        npu_inst_pe_1_4_3_n30), .S(npu_inst_pe_1_4_3_n6), .Z(
        npu_inst_pe_1_4_3_n32) );
  MUX2_X1 npu_inst_pe_1_4_3_U160 ( .A(npu_inst_pe_1_4_3_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_4_3_int_q_reg_v_1__0_), .S(npu_inst_pe_1_4_3_n4), .Z(
        npu_inst_pe_1_4_3_n31) );
  MUX2_X1 npu_inst_pe_1_4_3_U159 ( .A(npu_inst_pe_1_4_3_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_4_3_int_q_reg_v_3__0_), .S(npu_inst_pe_1_4_3_n4), .Z(
        npu_inst_pe_1_4_3_n30) );
  MUX2_X1 npu_inst_pe_1_4_3_U158 ( .A(npu_inst_pe_1_4_3_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_4_3_int_q_reg_v_5__0_), .S(npu_inst_pe_1_4_3_n4), .Z(
        npu_inst_pe_1_4_3_n29) );
  MUX2_X1 npu_inst_pe_1_4_3_U157 ( .A(npu_inst_pe_1_4_3_n28), .B(
        npu_inst_pe_1_4_3_n23), .S(npu_inst_pe_1_4_3_n8), .Z(
        npu_inst_pe_1_4_3_N94) );
  MUX2_X1 npu_inst_pe_1_4_3_U156 ( .A(npu_inst_pe_1_4_3_n25), .B(
        npu_inst_pe_1_4_3_n24), .S(npu_inst_pe_1_4_3_n6), .Z(
        npu_inst_pe_1_4_3_n28) );
  MUX2_X1 npu_inst_pe_1_4_3_U155 ( .A(npu_inst_pe_1_4_3_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_4_3_int_q_reg_v_1__1_), .S(npu_inst_pe_1_4_3_n4), .Z(
        npu_inst_pe_1_4_3_n25) );
  MUX2_X1 npu_inst_pe_1_4_3_U154 ( .A(npu_inst_pe_1_4_3_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_4_3_int_q_reg_v_3__1_), .S(npu_inst_pe_1_4_3_n4), .Z(
        npu_inst_pe_1_4_3_n24) );
  MUX2_X1 npu_inst_pe_1_4_3_U153 ( .A(npu_inst_pe_1_4_3_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_4_3_int_q_reg_v_5__1_), .S(npu_inst_pe_1_4_3_n4), .Z(
        npu_inst_pe_1_4_3_n23) );
  MUX2_X1 npu_inst_pe_1_4_3_U152 ( .A(npu_inst_pe_1_4_3_n22), .B(
        npu_inst_pe_1_4_3_n19), .S(npu_inst_pe_1_4_3_n8), .Z(
        npu_inst_int_data_x_4__3__1_) );
  MUX2_X1 npu_inst_pe_1_4_3_U151 ( .A(npu_inst_pe_1_4_3_n21), .B(
        npu_inst_pe_1_4_3_n20), .S(npu_inst_pe_1_4_3_n6), .Z(
        npu_inst_pe_1_4_3_n22) );
  MUX2_X1 npu_inst_pe_1_4_3_U150 ( .A(npu_inst_pe_1_4_3_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_4_3_int_q_reg_h_1__1_), .S(npu_inst_pe_1_4_3_n4), .Z(
        npu_inst_pe_1_4_3_n21) );
  MUX2_X1 npu_inst_pe_1_4_3_U149 ( .A(npu_inst_pe_1_4_3_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_4_3_int_q_reg_h_3__1_), .S(npu_inst_pe_1_4_3_n4), .Z(
        npu_inst_pe_1_4_3_n20) );
  MUX2_X1 npu_inst_pe_1_4_3_U148 ( .A(npu_inst_pe_1_4_3_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_4_3_int_q_reg_h_5__1_), .S(npu_inst_pe_1_4_3_n4), .Z(
        npu_inst_pe_1_4_3_n19) );
  MUX2_X1 npu_inst_pe_1_4_3_U147 ( .A(npu_inst_pe_1_4_3_n18), .B(
        npu_inst_pe_1_4_3_n15), .S(npu_inst_pe_1_4_3_n8), .Z(
        npu_inst_int_data_x_4__3__0_) );
  MUX2_X1 npu_inst_pe_1_4_3_U146 ( .A(npu_inst_pe_1_4_3_n17), .B(
        npu_inst_pe_1_4_3_n16), .S(npu_inst_pe_1_4_3_n6), .Z(
        npu_inst_pe_1_4_3_n18) );
  MUX2_X1 npu_inst_pe_1_4_3_U145 ( .A(npu_inst_pe_1_4_3_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_4_3_int_q_reg_h_1__0_), .S(npu_inst_pe_1_4_3_n4), .Z(
        npu_inst_pe_1_4_3_n17) );
  MUX2_X1 npu_inst_pe_1_4_3_U144 ( .A(npu_inst_pe_1_4_3_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_4_3_int_q_reg_h_3__0_), .S(npu_inst_pe_1_4_3_n4), .Z(
        npu_inst_pe_1_4_3_n16) );
  MUX2_X1 npu_inst_pe_1_4_3_U143 ( .A(npu_inst_pe_1_4_3_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_4_3_int_q_reg_h_5__0_), .S(npu_inst_pe_1_4_3_n4), .Z(
        npu_inst_pe_1_4_3_n15) );
  XOR2_X1 npu_inst_pe_1_4_3_U142 ( .A(npu_inst_pe_1_4_3_int_data_0_), .B(
        npu_inst_pe_1_4_3_int_q_acc_0_), .Z(npu_inst_pe_1_4_3_N73) );
  AND2_X1 npu_inst_pe_1_4_3_U141 ( .A1(npu_inst_pe_1_4_3_int_q_acc_0_), .A2(
        npu_inst_pe_1_4_3_int_data_0_), .ZN(npu_inst_pe_1_4_3_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_4_3_U140 ( .A(npu_inst_pe_1_4_3_int_q_acc_0_), .B(
        npu_inst_pe_1_4_3_n13), .ZN(npu_inst_pe_1_4_3_N65) );
  OR2_X1 npu_inst_pe_1_4_3_U139 ( .A1(npu_inst_pe_1_4_3_n13), .A2(
        npu_inst_pe_1_4_3_int_q_acc_0_), .ZN(npu_inst_pe_1_4_3_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_4_3_U138 ( .A(npu_inst_pe_1_4_3_int_q_acc_2_), .B(
        npu_inst_pe_1_4_3_add_79_carry_2_), .Z(npu_inst_pe_1_4_3_N75) );
  AND2_X1 npu_inst_pe_1_4_3_U137 ( .A1(npu_inst_pe_1_4_3_add_79_carry_2_), 
        .A2(npu_inst_pe_1_4_3_int_q_acc_2_), .ZN(
        npu_inst_pe_1_4_3_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_4_3_U136 ( .A(npu_inst_pe_1_4_3_int_q_acc_3_), .B(
        npu_inst_pe_1_4_3_add_79_carry_3_), .Z(npu_inst_pe_1_4_3_N76) );
  AND2_X1 npu_inst_pe_1_4_3_U135 ( .A1(npu_inst_pe_1_4_3_add_79_carry_3_), 
        .A2(npu_inst_pe_1_4_3_int_q_acc_3_), .ZN(
        npu_inst_pe_1_4_3_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_4_3_U134 ( .A(npu_inst_pe_1_4_3_int_q_acc_4_), .B(
        npu_inst_pe_1_4_3_add_79_carry_4_), .Z(npu_inst_pe_1_4_3_N77) );
  AND2_X1 npu_inst_pe_1_4_3_U133 ( .A1(npu_inst_pe_1_4_3_add_79_carry_4_), 
        .A2(npu_inst_pe_1_4_3_int_q_acc_4_), .ZN(
        npu_inst_pe_1_4_3_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_4_3_U132 ( .A(npu_inst_pe_1_4_3_int_q_acc_5_), .B(
        npu_inst_pe_1_4_3_add_79_carry_5_), .Z(npu_inst_pe_1_4_3_N78) );
  AND2_X1 npu_inst_pe_1_4_3_U131 ( .A1(npu_inst_pe_1_4_3_add_79_carry_5_), 
        .A2(npu_inst_pe_1_4_3_int_q_acc_5_), .ZN(
        npu_inst_pe_1_4_3_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_4_3_U130 ( .A(npu_inst_pe_1_4_3_int_q_acc_6_), .B(
        npu_inst_pe_1_4_3_add_79_carry_6_), .Z(npu_inst_pe_1_4_3_N79) );
  AND2_X1 npu_inst_pe_1_4_3_U129 ( .A1(npu_inst_pe_1_4_3_add_79_carry_6_), 
        .A2(npu_inst_pe_1_4_3_int_q_acc_6_), .ZN(
        npu_inst_pe_1_4_3_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_4_3_U128 ( .A(npu_inst_pe_1_4_3_int_q_acc_7_), .B(
        npu_inst_pe_1_4_3_add_79_carry_7_), .Z(npu_inst_pe_1_4_3_N80) );
  XNOR2_X1 npu_inst_pe_1_4_3_U127 ( .A(npu_inst_pe_1_4_3_sub_77_carry_2_), .B(
        npu_inst_pe_1_4_3_int_q_acc_2_), .ZN(npu_inst_pe_1_4_3_N67) );
  OR2_X1 npu_inst_pe_1_4_3_U126 ( .A1(npu_inst_pe_1_4_3_int_q_acc_2_), .A2(
        npu_inst_pe_1_4_3_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_4_3_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_4_3_U125 ( .A(npu_inst_pe_1_4_3_sub_77_carry_3_), .B(
        npu_inst_pe_1_4_3_int_q_acc_3_), .ZN(npu_inst_pe_1_4_3_N68) );
  OR2_X1 npu_inst_pe_1_4_3_U124 ( .A1(npu_inst_pe_1_4_3_int_q_acc_3_), .A2(
        npu_inst_pe_1_4_3_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_4_3_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_4_3_U123 ( .A(npu_inst_pe_1_4_3_sub_77_carry_4_), .B(
        npu_inst_pe_1_4_3_int_q_acc_4_), .ZN(npu_inst_pe_1_4_3_N69) );
  OR2_X1 npu_inst_pe_1_4_3_U122 ( .A1(npu_inst_pe_1_4_3_int_q_acc_4_), .A2(
        npu_inst_pe_1_4_3_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_4_3_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_4_3_U121 ( .A(npu_inst_pe_1_4_3_sub_77_carry_5_), .B(
        npu_inst_pe_1_4_3_int_q_acc_5_), .ZN(npu_inst_pe_1_4_3_N70) );
  OR2_X1 npu_inst_pe_1_4_3_U120 ( .A1(npu_inst_pe_1_4_3_int_q_acc_5_), .A2(
        npu_inst_pe_1_4_3_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_4_3_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_4_3_U119 ( .A(npu_inst_pe_1_4_3_sub_77_carry_6_), .B(
        npu_inst_pe_1_4_3_int_q_acc_6_), .ZN(npu_inst_pe_1_4_3_N71) );
  OR2_X1 npu_inst_pe_1_4_3_U118 ( .A1(npu_inst_pe_1_4_3_int_q_acc_6_), .A2(
        npu_inst_pe_1_4_3_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_4_3_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_4_3_U117 ( .A(npu_inst_pe_1_4_3_int_q_acc_7_), .B(
        npu_inst_pe_1_4_3_sub_77_carry_7_), .ZN(npu_inst_pe_1_4_3_N72) );
  INV_X1 npu_inst_pe_1_4_3_U116 ( .A(npu_inst_n77), .ZN(npu_inst_pe_1_4_3_n7)
         );
  INV_X1 npu_inst_pe_1_4_3_U115 ( .A(npu_inst_pe_1_4_3_n7), .ZN(
        npu_inst_pe_1_4_3_n6) );
  INV_X1 npu_inst_pe_1_4_3_U114 ( .A(npu_inst_n56), .ZN(npu_inst_pe_1_4_3_n3)
         );
  AOI22_X1 npu_inst_pe_1_4_3_U113 ( .A1(npu_inst_int_data_y_5__3__0_), .A2(
        npu_inst_pe_1_4_3_n58), .B1(npu_inst_pe_1_4_3_n114), .B2(
        npu_inst_pe_1_4_3_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_4_3_n57) );
  INV_X1 npu_inst_pe_1_4_3_U112 ( .A(npu_inst_pe_1_4_3_n57), .ZN(
        npu_inst_pe_1_4_3_n108) );
  AOI22_X1 npu_inst_pe_1_4_3_U111 ( .A1(npu_inst_int_data_y_5__3__0_), .A2(
        npu_inst_pe_1_4_3_n54), .B1(npu_inst_pe_1_4_3_n115), .B2(
        npu_inst_pe_1_4_3_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_4_3_n53) );
  INV_X1 npu_inst_pe_1_4_3_U110 ( .A(npu_inst_pe_1_4_3_n53), .ZN(
        npu_inst_pe_1_4_3_n109) );
  AOI22_X1 npu_inst_pe_1_4_3_U107 ( .A1(npu_inst_int_data_y_5__3__0_), .A2(
        npu_inst_pe_1_4_3_n50), .B1(npu_inst_pe_1_4_3_n116), .B2(
        npu_inst_pe_1_4_3_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_4_3_n49) );
  INV_X1 npu_inst_pe_1_4_3_U106 ( .A(npu_inst_pe_1_4_3_n49), .ZN(
        npu_inst_pe_1_4_3_n110) );
  AOI22_X1 npu_inst_pe_1_4_3_U105 ( .A1(npu_inst_int_data_y_5__3__0_), .A2(
        npu_inst_pe_1_4_3_n46), .B1(npu_inst_pe_1_4_3_n117), .B2(
        npu_inst_pe_1_4_3_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_4_3_n45) );
  INV_X1 npu_inst_pe_1_4_3_U104 ( .A(npu_inst_pe_1_4_3_n45), .ZN(
        npu_inst_pe_1_4_3_n111) );
  AOI22_X1 npu_inst_pe_1_4_3_U103 ( .A1(npu_inst_int_data_y_5__3__0_), .A2(
        npu_inst_pe_1_4_3_n42), .B1(npu_inst_pe_1_4_3_n119), .B2(
        npu_inst_pe_1_4_3_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_4_3_n41) );
  INV_X1 npu_inst_pe_1_4_3_U102 ( .A(npu_inst_pe_1_4_3_n41), .ZN(
        npu_inst_pe_1_4_3_n112) );
  AOI22_X1 npu_inst_pe_1_4_3_U101 ( .A1(npu_inst_int_data_y_5__3__1_), .A2(
        npu_inst_pe_1_4_3_n58), .B1(npu_inst_pe_1_4_3_n114), .B2(
        npu_inst_pe_1_4_3_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_4_3_n59) );
  INV_X1 npu_inst_pe_1_4_3_U100 ( .A(npu_inst_pe_1_4_3_n59), .ZN(
        npu_inst_pe_1_4_3_n102) );
  AOI22_X1 npu_inst_pe_1_4_3_U99 ( .A1(npu_inst_int_data_y_5__3__1_), .A2(
        npu_inst_pe_1_4_3_n54), .B1(npu_inst_pe_1_4_3_n115), .B2(
        npu_inst_pe_1_4_3_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_4_3_n55) );
  INV_X1 npu_inst_pe_1_4_3_U98 ( .A(npu_inst_pe_1_4_3_n55), .ZN(
        npu_inst_pe_1_4_3_n103) );
  AOI22_X1 npu_inst_pe_1_4_3_U97 ( .A1(npu_inst_int_data_y_5__3__1_), .A2(
        npu_inst_pe_1_4_3_n50), .B1(npu_inst_pe_1_4_3_n116), .B2(
        npu_inst_pe_1_4_3_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_4_3_n51) );
  INV_X1 npu_inst_pe_1_4_3_U96 ( .A(npu_inst_pe_1_4_3_n51), .ZN(
        npu_inst_pe_1_4_3_n104) );
  AOI22_X1 npu_inst_pe_1_4_3_U95 ( .A1(npu_inst_int_data_y_5__3__1_), .A2(
        npu_inst_pe_1_4_3_n46), .B1(npu_inst_pe_1_4_3_n117), .B2(
        npu_inst_pe_1_4_3_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_4_3_n47) );
  INV_X1 npu_inst_pe_1_4_3_U94 ( .A(npu_inst_pe_1_4_3_n47), .ZN(
        npu_inst_pe_1_4_3_n105) );
  AOI22_X1 npu_inst_pe_1_4_3_U93 ( .A1(npu_inst_int_data_y_5__3__1_), .A2(
        npu_inst_pe_1_4_3_n42), .B1(npu_inst_pe_1_4_3_n119), .B2(
        npu_inst_pe_1_4_3_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_4_3_n43) );
  INV_X1 npu_inst_pe_1_4_3_U92 ( .A(npu_inst_pe_1_4_3_n43), .ZN(
        npu_inst_pe_1_4_3_n106) );
  AOI22_X1 npu_inst_pe_1_4_3_U91 ( .A1(npu_inst_pe_1_4_3_n38), .A2(
        npu_inst_int_data_y_5__3__1_), .B1(npu_inst_pe_1_4_3_n118), .B2(
        npu_inst_pe_1_4_3_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_4_3_n39) );
  INV_X1 npu_inst_pe_1_4_3_U90 ( .A(npu_inst_pe_1_4_3_n39), .ZN(
        npu_inst_pe_1_4_3_n107) );
  AOI22_X1 npu_inst_pe_1_4_3_U89 ( .A1(npu_inst_pe_1_4_3_n38), .A2(
        npu_inst_int_data_y_5__3__0_), .B1(npu_inst_pe_1_4_3_n118), .B2(
        npu_inst_pe_1_4_3_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_4_3_n37) );
  INV_X1 npu_inst_pe_1_4_3_U88 ( .A(npu_inst_pe_1_4_3_n37), .ZN(
        npu_inst_pe_1_4_3_n113) );
  NAND2_X1 npu_inst_pe_1_4_3_U87 ( .A1(npu_inst_pe_1_4_3_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_4_3_n60), .ZN(npu_inst_pe_1_4_3_n74) );
  OAI21_X1 npu_inst_pe_1_4_3_U86 ( .B1(npu_inst_pe_1_4_3_n63), .B2(
        npu_inst_pe_1_4_3_n60), .A(npu_inst_pe_1_4_3_n74), .ZN(
        npu_inst_pe_1_4_3_n97) );
  NAND2_X1 npu_inst_pe_1_4_3_U85 ( .A1(npu_inst_pe_1_4_3_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_4_3_n60), .ZN(npu_inst_pe_1_4_3_n73) );
  OAI21_X1 npu_inst_pe_1_4_3_U84 ( .B1(npu_inst_pe_1_4_3_n61), .B2(
        npu_inst_pe_1_4_3_n60), .A(npu_inst_pe_1_4_3_n73), .ZN(
        npu_inst_pe_1_4_3_n96) );
  NAND2_X1 npu_inst_pe_1_4_3_U83 ( .A1(npu_inst_pe_1_4_3_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_4_3_n56), .ZN(npu_inst_pe_1_4_3_n72) );
  OAI21_X1 npu_inst_pe_1_4_3_U82 ( .B1(npu_inst_pe_1_4_3_n63), .B2(
        npu_inst_pe_1_4_3_n56), .A(npu_inst_pe_1_4_3_n72), .ZN(
        npu_inst_pe_1_4_3_n95) );
  NAND2_X1 npu_inst_pe_1_4_3_U81 ( .A1(npu_inst_pe_1_4_3_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_4_3_n56), .ZN(npu_inst_pe_1_4_3_n71) );
  OAI21_X1 npu_inst_pe_1_4_3_U80 ( .B1(npu_inst_pe_1_4_3_n61), .B2(
        npu_inst_pe_1_4_3_n56), .A(npu_inst_pe_1_4_3_n71), .ZN(
        npu_inst_pe_1_4_3_n94) );
  NAND2_X1 npu_inst_pe_1_4_3_U79 ( .A1(npu_inst_pe_1_4_3_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_4_3_n52), .ZN(npu_inst_pe_1_4_3_n70) );
  OAI21_X1 npu_inst_pe_1_4_3_U78 ( .B1(npu_inst_pe_1_4_3_n63), .B2(
        npu_inst_pe_1_4_3_n52), .A(npu_inst_pe_1_4_3_n70), .ZN(
        npu_inst_pe_1_4_3_n93) );
  NAND2_X1 npu_inst_pe_1_4_3_U77 ( .A1(npu_inst_pe_1_4_3_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_4_3_n52), .ZN(npu_inst_pe_1_4_3_n69) );
  OAI21_X1 npu_inst_pe_1_4_3_U76 ( .B1(npu_inst_pe_1_4_3_n61), .B2(
        npu_inst_pe_1_4_3_n52), .A(npu_inst_pe_1_4_3_n69), .ZN(
        npu_inst_pe_1_4_3_n92) );
  NAND2_X1 npu_inst_pe_1_4_3_U75 ( .A1(npu_inst_pe_1_4_3_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_4_3_n48), .ZN(npu_inst_pe_1_4_3_n68) );
  OAI21_X1 npu_inst_pe_1_4_3_U74 ( .B1(npu_inst_pe_1_4_3_n63), .B2(
        npu_inst_pe_1_4_3_n48), .A(npu_inst_pe_1_4_3_n68), .ZN(
        npu_inst_pe_1_4_3_n91) );
  NAND2_X1 npu_inst_pe_1_4_3_U73 ( .A1(npu_inst_pe_1_4_3_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_4_3_n48), .ZN(npu_inst_pe_1_4_3_n67) );
  OAI21_X1 npu_inst_pe_1_4_3_U72 ( .B1(npu_inst_pe_1_4_3_n61), .B2(
        npu_inst_pe_1_4_3_n48), .A(npu_inst_pe_1_4_3_n67), .ZN(
        npu_inst_pe_1_4_3_n90) );
  NAND2_X1 npu_inst_pe_1_4_3_U71 ( .A1(npu_inst_pe_1_4_3_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_4_3_n44), .ZN(npu_inst_pe_1_4_3_n66) );
  OAI21_X1 npu_inst_pe_1_4_3_U70 ( .B1(npu_inst_pe_1_4_3_n63), .B2(
        npu_inst_pe_1_4_3_n44), .A(npu_inst_pe_1_4_3_n66), .ZN(
        npu_inst_pe_1_4_3_n89) );
  NAND2_X1 npu_inst_pe_1_4_3_U69 ( .A1(npu_inst_pe_1_4_3_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_4_3_n44), .ZN(npu_inst_pe_1_4_3_n65) );
  OAI21_X1 npu_inst_pe_1_4_3_U68 ( .B1(npu_inst_pe_1_4_3_n61), .B2(
        npu_inst_pe_1_4_3_n44), .A(npu_inst_pe_1_4_3_n65), .ZN(
        npu_inst_pe_1_4_3_n88) );
  NAND2_X1 npu_inst_pe_1_4_3_U67 ( .A1(npu_inst_pe_1_4_3_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_4_3_n40), .ZN(npu_inst_pe_1_4_3_n64) );
  OAI21_X1 npu_inst_pe_1_4_3_U66 ( .B1(npu_inst_pe_1_4_3_n63), .B2(
        npu_inst_pe_1_4_3_n40), .A(npu_inst_pe_1_4_3_n64), .ZN(
        npu_inst_pe_1_4_3_n87) );
  NAND2_X1 npu_inst_pe_1_4_3_U65 ( .A1(npu_inst_pe_1_4_3_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_4_3_n40), .ZN(npu_inst_pe_1_4_3_n62) );
  OAI21_X1 npu_inst_pe_1_4_3_U64 ( .B1(npu_inst_pe_1_4_3_n61), .B2(
        npu_inst_pe_1_4_3_n40), .A(npu_inst_pe_1_4_3_n62), .ZN(
        npu_inst_pe_1_4_3_n86) );
  AND2_X1 npu_inst_pe_1_4_3_U63 ( .A1(npu_inst_pe_1_4_3_N93), .A2(npu_inst_n56), .ZN(npu_inst_int_data_y_4__3__0_) );
  AND2_X1 npu_inst_pe_1_4_3_U62 ( .A1(npu_inst_n56), .A2(npu_inst_pe_1_4_3_N94), .ZN(npu_inst_int_data_y_4__3__1_) );
  NOR3_X1 npu_inst_pe_1_4_3_U61 ( .A1(npu_inst_pe_1_4_3_n26), .A2(npu_inst_n56), .A3(npu_inst_int_ckg[28]), .ZN(npu_inst_pe_1_4_3_n85) );
  OR2_X1 npu_inst_pe_1_4_3_U60 ( .A1(npu_inst_pe_1_4_3_n85), .A2(
        npu_inst_pe_1_4_3_n2), .ZN(npu_inst_pe_1_4_3_N84) );
  AND2_X1 npu_inst_pe_1_4_3_U59 ( .A1(npu_inst_pe_1_4_3_int_q_acc_0_), .A2(
        npu_inst_pe_1_4_3_n1), .ZN(npu_inst_int_data_res_4__3__0_) );
  AND2_X1 npu_inst_pe_1_4_3_U58 ( .A1(npu_inst_pe_1_4_3_n2), .A2(
        npu_inst_pe_1_4_3_int_q_acc_7_), .ZN(npu_inst_int_data_res_4__3__7_)
         );
  AND2_X1 npu_inst_pe_1_4_3_U57 ( .A1(npu_inst_pe_1_4_3_int_q_acc_1_), .A2(
        npu_inst_pe_1_4_3_n1), .ZN(npu_inst_int_data_res_4__3__1_) );
  AND2_X1 npu_inst_pe_1_4_3_U56 ( .A1(npu_inst_pe_1_4_3_int_q_acc_2_), .A2(
        npu_inst_pe_1_4_3_n1), .ZN(npu_inst_int_data_res_4__3__2_) );
  AND2_X1 npu_inst_pe_1_4_3_U55 ( .A1(npu_inst_pe_1_4_3_int_q_acc_3_), .A2(
        npu_inst_pe_1_4_3_n2), .ZN(npu_inst_int_data_res_4__3__3_) );
  AND2_X1 npu_inst_pe_1_4_3_U54 ( .A1(npu_inst_pe_1_4_3_int_q_acc_4_), .A2(
        npu_inst_pe_1_4_3_n2), .ZN(npu_inst_int_data_res_4__3__4_) );
  AND2_X1 npu_inst_pe_1_4_3_U53 ( .A1(npu_inst_pe_1_4_3_int_q_acc_5_), .A2(
        npu_inst_pe_1_4_3_n2), .ZN(npu_inst_int_data_res_4__3__5_) );
  AND2_X1 npu_inst_pe_1_4_3_U52 ( .A1(npu_inst_pe_1_4_3_int_q_acc_6_), .A2(
        npu_inst_pe_1_4_3_n2), .ZN(npu_inst_int_data_res_4__3__6_) );
  AOI222_X1 npu_inst_pe_1_4_3_U51 ( .A1(npu_inst_int_data_res_5__3__0_), .A2(
        npu_inst_pe_1_4_3_n1), .B1(npu_inst_pe_1_4_3_N73), .B2(
        npu_inst_pe_1_4_3_n76), .C1(npu_inst_pe_1_4_3_N65), .C2(
        npu_inst_pe_1_4_3_n77), .ZN(npu_inst_pe_1_4_3_n84) );
  INV_X1 npu_inst_pe_1_4_3_U50 ( .A(npu_inst_pe_1_4_3_n84), .ZN(
        npu_inst_pe_1_4_3_n101) );
  AOI222_X1 npu_inst_pe_1_4_3_U49 ( .A1(npu_inst_int_data_res_5__3__7_), .A2(
        npu_inst_pe_1_4_3_n1), .B1(npu_inst_pe_1_4_3_N80), .B2(
        npu_inst_pe_1_4_3_n76), .C1(npu_inst_pe_1_4_3_N72), .C2(
        npu_inst_pe_1_4_3_n77), .ZN(npu_inst_pe_1_4_3_n75) );
  INV_X1 npu_inst_pe_1_4_3_U48 ( .A(npu_inst_pe_1_4_3_n75), .ZN(
        npu_inst_pe_1_4_3_n33) );
  AOI222_X1 npu_inst_pe_1_4_3_U47 ( .A1(npu_inst_int_data_res_5__3__1_), .A2(
        npu_inst_pe_1_4_3_n1), .B1(npu_inst_pe_1_4_3_N74), .B2(
        npu_inst_pe_1_4_3_n76), .C1(npu_inst_pe_1_4_3_N66), .C2(
        npu_inst_pe_1_4_3_n77), .ZN(npu_inst_pe_1_4_3_n83) );
  INV_X1 npu_inst_pe_1_4_3_U46 ( .A(npu_inst_pe_1_4_3_n83), .ZN(
        npu_inst_pe_1_4_3_n100) );
  AOI222_X1 npu_inst_pe_1_4_3_U45 ( .A1(npu_inst_int_data_res_5__3__2_), .A2(
        npu_inst_pe_1_4_3_n1), .B1(npu_inst_pe_1_4_3_N75), .B2(
        npu_inst_pe_1_4_3_n76), .C1(npu_inst_pe_1_4_3_N67), .C2(
        npu_inst_pe_1_4_3_n77), .ZN(npu_inst_pe_1_4_3_n82) );
  INV_X1 npu_inst_pe_1_4_3_U44 ( .A(npu_inst_pe_1_4_3_n82), .ZN(
        npu_inst_pe_1_4_3_n99) );
  AOI222_X1 npu_inst_pe_1_4_3_U43 ( .A1(npu_inst_int_data_res_5__3__3_), .A2(
        npu_inst_pe_1_4_3_n1), .B1(npu_inst_pe_1_4_3_N76), .B2(
        npu_inst_pe_1_4_3_n76), .C1(npu_inst_pe_1_4_3_N68), .C2(
        npu_inst_pe_1_4_3_n77), .ZN(npu_inst_pe_1_4_3_n81) );
  INV_X1 npu_inst_pe_1_4_3_U42 ( .A(npu_inst_pe_1_4_3_n81), .ZN(
        npu_inst_pe_1_4_3_n98) );
  AOI222_X1 npu_inst_pe_1_4_3_U41 ( .A1(npu_inst_int_data_res_5__3__4_), .A2(
        npu_inst_pe_1_4_3_n1), .B1(npu_inst_pe_1_4_3_N77), .B2(
        npu_inst_pe_1_4_3_n76), .C1(npu_inst_pe_1_4_3_N69), .C2(
        npu_inst_pe_1_4_3_n77), .ZN(npu_inst_pe_1_4_3_n80) );
  INV_X1 npu_inst_pe_1_4_3_U40 ( .A(npu_inst_pe_1_4_3_n80), .ZN(
        npu_inst_pe_1_4_3_n36) );
  AOI222_X1 npu_inst_pe_1_4_3_U39 ( .A1(npu_inst_int_data_res_5__3__5_), .A2(
        npu_inst_pe_1_4_3_n1), .B1(npu_inst_pe_1_4_3_N78), .B2(
        npu_inst_pe_1_4_3_n76), .C1(npu_inst_pe_1_4_3_N70), .C2(
        npu_inst_pe_1_4_3_n77), .ZN(npu_inst_pe_1_4_3_n79) );
  INV_X1 npu_inst_pe_1_4_3_U38 ( .A(npu_inst_pe_1_4_3_n79), .ZN(
        npu_inst_pe_1_4_3_n35) );
  AOI222_X1 npu_inst_pe_1_4_3_U37 ( .A1(npu_inst_int_data_res_5__3__6_), .A2(
        npu_inst_pe_1_4_3_n1), .B1(npu_inst_pe_1_4_3_N79), .B2(
        npu_inst_pe_1_4_3_n76), .C1(npu_inst_pe_1_4_3_N71), .C2(
        npu_inst_pe_1_4_3_n77), .ZN(npu_inst_pe_1_4_3_n78) );
  INV_X1 npu_inst_pe_1_4_3_U36 ( .A(npu_inst_pe_1_4_3_n78), .ZN(
        npu_inst_pe_1_4_3_n34) );
  INV_X1 npu_inst_pe_1_4_3_U35 ( .A(npu_inst_pe_1_4_3_int_data_1_), .ZN(
        npu_inst_pe_1_4_3_n14) );
  AND2_X1 npu_inst_pe_1_4_3_U34 ( .A1(npu_inst_int_data_x_4__3__1_), .A2(
        npu_inst_pe_1_4_3_int_q_weight_1_), .ZN(npu_inst_pe_1_4_3_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_4_3_U33 ( .A1(npu_inst_int_data_x_4__3__0_), .A2(
        npu_inst_pe_1_4_3_int_q_weight_1_), .ZN(npu_inst_pe_1_4_3_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_4_3_U32 ( .A1(npu_inst_n56), .A2(
        npu_inst_int_data_y_5__3__1_), .B1(npu_inst_pe_1_4_3_n3), .B2(
        npu_inst_int_data_x_4__4__1_), .ZN(npu_inst_pe_1_4_3_n63) );
  AOI22_X1 npu_inst_pe_1_4_3_U31 ( .A1(npu_inst_n56), .A2(
        npu_inst_int_data_y_5__3__0_), .B1(npu_inst_pe_1_4_3_n3), .B2(
        npu_inst_int_data_x_4__4__0_), .ZN(npu_inst_pe_1_4_3_n61) );
  INV_X1 npu_inst_pe_1_4_3_U30 ( .A(npu_inst_pe_1_4_3_int_data_0_), .ZN(
        npu_inst_pe_1_4_3_n13) );
  INV_X1 npu_inst_pe_1_4_3_U29 ( .A(npu_inst_n69), .ZN(npu_inst_pe_1_4_3_n5)
         );
  OR3_X1 npu_inst_pe_1_4_3_U28 ( .A1(npu_inst_pe_1_4_3_n6), .A2(
        npu_inst_pe_1_4_3_n8), .A3(npu_inst_pe_1_4_3_n5), .ZN(
        npu_inst_pe_1_4_3_n56) );
  OR3_X1 npu_inst_pe_1_4_3_U27 ( .A1(npu_inst_pe_1_4_3_n5), .A2(
        npu_inst_pe_1_4_3_n8), .A3(npu_inst_pe_1_4_3_n7), .ZN(
        npu_inst_pe_1_4_3_n48) );
  INV_X1 npu_inst_pe_1_4_3_U26 ( .A(npu_inst_pe_1_4_3_n5), .ZN(
        npu_inst_pe_1_4_3_n4) );
  INV_X1 npu_inst_pe_1_4_3_U25 ( .A(npu_inst_n124), .ZN(npu_inst_pe_1_4_3_n12)
         );
  OR3_X1 npu_inst_pe_1_4_3_U24 ( .A1(npu_inst_pe_1_4_3_n4), .A2(
        npu_inst_pe_1_4_3_n8), .A3(npu_inst_pe_1_4_3_n7), .ZN(
        npu_inst_pe_1_4_3_n52) );
  OR3_X1 npu_inst_pe_1_4_3_U23 ( .A1(npu_inst_pe_1_4_3_n6), .A2(
        npu_inst_pe_1_4_3_n8), .A3(npu_inst_pe_1_4_3_n4), .ZN(
        npu_inst_pe_1_4_3_n60) );
  NOR2_X1 npu_inst_pe_1_4_3_U22 ( .A1(npu_inst_pe_1_4_3_n60), .A2(
        npu_inst_pe_1_4_3_n3), .ZN(npu_inst_pe_1_4_3_n58) );
  NOR2_X1 npu_inst_pe_1_4_3_U21 ( .A1(npu_inst_pe_1_4_3_n56), .A2(
        npu_inst_pe_1_4_3_n3), .ZN(npu_inst_pe_1_4_3_n54) );
  NOR2_X1 npu_inst_pe_1_4_3_U20 ( .A1(npu_inst_pe_1_4_3_n52), .A2(
        npu_inst_pe_1_4_3_n3), .ZN(npu_inst_pe_1_4_3_n50) );
  NOR2_X1 npu_inst_pe_1_4_3_U19 ( .A1(npu_inst_pe_1_4_3_n48), .A2(
        npu_inst_pe_1_4_3_n3), .ZN(npu_inst_pe_1_4_3_n46) );
  NOR2_X1 npu_inst_pe_1_4_3_U18 ( .A1(npu_inst_pe_1_4_3_n40), .A2(
        npu_inst_pe_1_4_3_n3), .ZN(npu_inst_pe_1_4_3_n38) );
  NOR2_X1 npu_inst_pe_1_4_3_U17 ( .A1(npu_inst_pe_1_4_3_n44), .A2(
        npu_inst_pe_1_4_3_n3), .ZN(npu_inst_pe_1_4_3_n42) );
  BUF_X1 npu_inst_pe_1_4_3_U16 ( .A(npu_inst_n99), .Z(npu_inst_pe_1_4_3_n8) );
  BUF_X1 npu_inst_pe_1_4_3_U15 ( .A(npu_inst_pe_1_4_3_n12), .Z(
        npu_inst_pe_1_4_3_n11) );
  BUF_X1 npu_inst_pe_1_4_3_U14 ( .A(npu_inst_pe_1_4_3_n12), .Z(
        npu_inst_pe_1_4_3_n10) );
  BUF_X1 npu_inst_pe_1_4_3_U13 ( .A(npu_inst_pe_1_4_3_n12), .Z(
        npu_inst_pe_1_4_3_n9) );
  INV_X1 npu_inst_pe_1_4_3_U12 ( .A(npu_inst_pe_1_4_3_n38), .ZN(
        npu_inst_pe_1_4_3_n118) );
  INV_X1 npu_inst_pe_1_4_3_U11 ( .A(npu_inst_pe_1_4_3_n58), .ZN(
        npu_inst_pe_1_4_3_n114) );
  INV_X1 npu_inst_pe_1_4_3_U10 ( .A(npu_inst_pe_1_4_3_n54), .ZN(
        npu_inst_pe_1_4_3_n115) );
  INV_X1 npu_inst_pe_1_4_3_U9 ( .A(npu_inst_pe_1_4_3_n50), .ZN(
        npu_inst_pe_1_4_3_n116) );
  INV_X1 npu_inst_pe_1_4_3_U8 ( .A(npu_inst_pe_1_4_3_n46), .ZN(
        npu_inst_pe_1_4_3_n117) );
  INV_X1 npu_inst_pe_1_4_3_U7 ( .A(npu_inst_pe_1_4_3_n42), .ZN(
        npu_inst_pe_1_4_3_n119) );
  BUF_X1 npu_inst_pe_1_4_3_U6 ( .A(npu_inst_n21), .Z(npu_inst_pe_1_4_3_n2) );
  BUF_X1 npu_inst_pe_1_4_3_U5 ( .A(npu_inst_n21), .Z(npu_inst_pe_1_4_3_n1) );
  NOR2_X1 npu_inst_pe_1_4_3_U4 ( .A1(npu_inst_pe_1_4_3_int_q_weight_0_), .A2(
        npu_inst_pe_1_4_3_n1), .ZN(npu_inst_pe_1_4_3_n76) );
  NOR2_X1 npu_inst_pe_1_4_3_U3 ( .A1(npu_inst_pe_1_4_3_n27), .A2(
        npu_inst_pe_1_4_3_n1), .ZN(npu_inst_pe_1_4_3_n77) );
  FA_X1 npu_inst_pe_1_4_3_sub_77_U2_1 ( .A(npu_inst_pe_1_4_3_int_q_acc_1_), 
        .B(npu_inst_pe_1_4_3_n14), .CI(npu_inst_pe_1_4_3_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_4_3_sub_77_carry_2_), .S(npu_inst_pe_1_4_3_N66) );
  FA_X1 npu_inst_pe_1_4_3_add_79_U1_1 ( .A(npu_inst_pe_1_4_3_int_q_acc_1_), 
        .B(npu_inst_pe_1_4_3_int_data_1_), .CI(
        npu_inst_pe_1_4_3_add_79_carry_1_), .CO(
        npu_inst_pe_1_4_3_add_79_carry_2_), .S(npu_inst_pe_1_4_3_N74) );
  NAND3_X1 npu_inst_pe_1_4_3_U109 ( .A1(npu_inst_pe_1_4_3_n5), .A2(
        npu_inst_pe_1_4_3_n7), .A3(npu_inst_pe_1_4_3_n8), .ZN(
        npu_inst_pe_1_4_3_n44) );
  NAND3_X1 npu_inst_pe_1_4_3_U108 ( .A1(npu_inst_pe_1_4_3_n4), .A2(
        npu_inst_pe_1_4_3_n7), .A3(npu_inst_pe_1_4_3_n8), .ZN(
        npu_inst_pe_1_4_3_n40) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_4_3_n34), .CK(
        npu_inst_pe_1_4_3_net3488), .RN(npu_inst_pe_1_4_3_n9), .Q(
        npu_inst_pe_1_4_3_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_4_3_n35), .CK(
        npu_inst_pe_1_4_3_net3488), .RN(npu_inst_pe_1_4_3_n9), .Q(
        npu_inst_pe_1_4_3_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_4_3_n36), .CK(
        npu_inst_pe_1_4_3_net3488), .RN(npu_inst_pe_1_4_3_n9), .Q(
        npu_inst_pe_1_4_3_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_4_3_n98), .CK(
        npu_inst_pe_1_4_3_net3488), .RN(npu_inst_pe_1_4_3_n9), .Q(
        npu_inst_pe_1_4_3_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_4_3_n99), .CK(
        npu_inst_pe_1_4_3_net3488), .RN(npu_inst_pe_1_4_3_n9), .Q(
        npu_inst_pe_1_4_3_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_4_3_n100), 
        .CK(npu_inst_pe_1_4_3_net3488), .RN(npu_inst_pe_1_4_3_n9), .Q(
        npu_inst_pe_1_4_3_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_4_3_n33), .CK(
        npu_inst_pe_1_4_3_net3488), .RN(npu_inst_pe_1_4_3_n9), .Q(
        npu_inst_pe_1_4_3_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_4_3_n101), 
        .CK(npu_inst_pe_1_4_3_net3488), .RN(npu_inst_pe_1_4_3_n9), .Q(
        npu_inst_pe_1_4_3_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_weight_reg_0_ ( .D(npu_inst_n110), .CK(
        npu_inst_pe_1_4_3_net3494), .RN(npu_inst_pe_1_4_3_n9), .Q(
        npu_inst_pe_1_4_3_int_q_weight_0_), .QN(npu_inst_pe_1_4_3_n27) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_weight_reg_1_ ( .D(npu_inst_n116), .CK(
        npu_inst_pe_1_4_3_net3494), .RN(npu_inst_pe_1_4_3_n9), .Q(
        npu_inst_pe_1_4_3_int_q_weight_1_), .QN(npu_inst_pe_1_4_3_n26) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_4_3_n113), 
        .CK(npu_inst_pe_1_4_3_net3494), .RN(npu_inst_pe_1_4_3_n9), .Q(
        npu_inst_pe_1_4_3_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_4_3_n107), 
        .CK(npu_inst_pe_1_4_3_net3494), .RN(npu_inst_pe_1_4_3_n9), .Q(
        npu_inst_pe_1_4_3_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_4_3_n112), 
        .CK(npu_inst_pe_1_4_3_net3494), .RN(npu_inst_pe_1_4_3_n10), .Q(
        npu_inst_pe_1_4_3_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_4_3_n106), 
        .CK(npu_inst_pe_1_4_3_net3494), .RN(npu_inst_pe_1_4_3_n10), .Q(
        npu_inst_pe_1_4_3_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_4_3_n111), 
        .CK(npu_inst_pe_1_4_3_net3494), .RN(npu_inst_pe_1_4_3_n10), .Q(
        npu_inst_pe_1_4_3_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_4_3_n105), 
        .CK(npu_inst_pe_1_4_3_net3494), .RN(npu_inst_pe_1_4_3_n10), .Q(
        npu_inst_pe_1_4_3_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_4_3_n110), 
        .CK(npu_inst_pe_1_4_3_net3494), .RN(npu_inst_pe_1_4_3_n10), .Q(
        npu_inst_pe_1_4_3_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_4_3_n104), 
        .CK(npu_inst_pe_1_4_3_net3494), .RN(npu_inst_pe_1_4_3_n10), .Q(
        npu_inst_pe_1_4_3_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_4_3_n109), 
        .CK(npu_inst_pe_1_4_3_net3494), .RN(npu_inst_pe_1_4_3_n10), .Q(
        npu_inst_pe_1_4_3_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_4_3_n103), 
        .CK(npu_inst_pe_1_4_3_net3494), .RN(npu_inst_pe_1_4_3_n10), .Q(
        npu_inst_pe_1_4_3_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_4_3_n108), 
        .CK(npu_inst_pe_1_4_3_net3494), .RN(npu_inst_pe_1_4_3_n10), .Q(
        npu_inst_pe_1_4_3_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_4_3_n102), 
        .CK(npu_inst_pe_1_4_3_net3494), .RN(npu_inst_pe_1_4_3_n10), .Q(
        npu_inst_pe_1_4_3_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_4_3_n86), 
        .CK(npu_inst_pe_1_4_3_net3494), .RN(npu_inst_pe_1_4_3_n10), .Q(
        npu_inst_pe_1_4_3_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_4_3_n87), 
        .CK(npu_inst_pe_1_4_3_net3494), .RN(npu_inst_pe_1_4_3_n10), .Q(
        npu_inst_pe_1_4_3_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_4_3_n88), 
        .CK(npu_inst_pe_1_4_3_net3494), .RN(npu_inst_pe_1_4_3_n11), .Q(
        npu_inst_pe_1_4_3_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_4_3_n89), 
        .CK(npu_inst_pe_1_4_3_net3494), .RN(npu_inst_pe_1_4_3_n11), .Q(
        npu_inst_pe_1_4_3_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_4_3_n90), 
        .CK(npu_inst_pe_1_4_3_net3494), .RN(npu_inst_pe_1_4_3_n11), .Q(
        npu_inst_pe_1_4_3_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_4_3_n91), 
        .CK(npu_inst_pe_1_4_3_net3494), .RN(npu_inst_pe_1_4_3_n11), .Q(
        npu_inst_pe_1_4_3_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_4_3_n92), 
        .CK(npu_inst_pe_1_4_3_net3494), .RN(npu_inst_pe_1_4_3_n11), .Q(
        npu_inst_pe_1_4_3_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_4_3_n93), 
        .CK(npu_inst_pe_1_4_3_net3494), .RN(npu_inst_pe_1_4_3_n11), .Q(
        npu_inst_pe_1_4_3_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_4_3_n94), 
        .CK(npu_inst_pe_1_4_3_net3494), .RN(npu_inst_pe_1_4_3_n11), .Q(
        npu_inst_pe_1_4_3_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_4_3_n95), 
        .CK(npu_inst_pe_1_4_3_net3494), .RN(npu_inst_pe_1_4_3_n11), .Q(
        npu_inst_pe_1_4_3_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_4_3_n96), 
        .CK(npu_inst_pe_1_4_3_net3494), .RN(npu_inst_pe_1_4_3_n11), .Q(
        npu_inst_pe_1_4_3_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_4_3_n97), 
        .CK(npu_inst_pe_1_4_3_net3494), .RN(npu_inst_pe_1_4_3_n11), .Q(
        npu_inst_pe_1_4_3_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_4_3_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_4_3_N84), .SE(1'b0), .GCK(npu_inst_pe_1_4_3_net3488) );
  CLKGATETST_X1 npu_inst_pe_1_4_3_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n63), .SE(1'b0), .GCK(npu_inst_pe_1_4_3_net3494) );
  MUX2_X1 npu_inst_pe_1_4_4_U162 ( .A(npu_inst_pe_1_4_4_n32), .B(
        npu_inst_pe_1_4_4_n29), .S(npu_inst_pe_1_4_4_n8), .Z(
        npu_inst_pe_1_4_4_N93) );
  MUX2_X1 npu_inst_pe_1_4_4_U161 ( .A(npu_inst_pe_1_4_4_n31), .B(
        npu_inst_pe_1_4_4_n30), .S(npu_inst_pe_1_4_4_n6), .Z(
        npu_inst_pe_1_4_4_n32) );
  MUX2_X1 npu_inst_pe_1_4_4_U160 ( .A(npu_inst_pe_1_4_4_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_4_4_int_q_reg_v_1__0_), .S(npu_inst_pe_1_4_4_n4), .Z(
        npu_inst_pe_1_4_4_n31) );
  MUX2_X1 npu_inst_pe_1_4_4_U159 ( .A(npu_inst_pe_1_4_4_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_4_4_int_q_reg_v_3__0_), .S(npu_inst_pe_1_4_4_n4), .Z(
        npu_inst_pe_1_4_4_n30) );
  MUX2_X1 npu_inst_pe_1_4_4_U158 ( .A(npu_inst_pe_1_4_4_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_4_4_int_q_reg_v_5__0_), .S(npu_inst_pe_1_4_4_n4), .Z(
        npu_inst_pe_1_4_4_n29) );
  MUX2_X1 npu_inst_pe_1_4_4_U157 ( .A(npu_inst_pe_1_4_4_n28), .B(
        npu_inst_pe_1_4_4_n23), .S(npu_inst_pe_1_4_4_n8), .Z(
        npu_inst_pe_1_4_4_N94) );
  MUX2_X1 npu_inst_pe_1_4_4_U156 ( .A(npu_inst_pe_1_4_4_n25), .B(
        npu_inst_pe_1_4_4_n24), .S(npu_inst_pe_1_4_4_n6), .Z(
        npu_inst_pe_1_4_4_n28) );
  MUX2_X1 npu_inst_pe_1_4_4_U155 ( .A(npu_inst_pe_1_4_4_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_4_4_int_q_reg_v_1__1_), .S(npu_inst_pe_1_4_4_n4), .Z(
        npu_inst_pe_1_4_4_n25) );
  MUX2_X1 npu_inst_pe_1_4_4_U154 ( .A(npu_inst_pe_1_4_4_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_4_4_int_q_reg_v_3__1_), .S(npu_inst_pe_1_4_4_n4), .Z(
        npu_inst_pe_1_4_4_n24) );
  MUX2_X1 npu_inst_pe_1_4_4_U153 ( .A(npu_inst_pe_1_4_4_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_4_4_int_q_reg_v_5__1_), .S(npu_inst_pe_1_4_4_n4), .Z(
        npu_inst_pe_1_4_4_n23) );
  MUX2_X1 npu_inst_pe_1_4_4_U152 ( .A(npu_inst_pe_1_4_4_n22), .B(
        npu_inst_pe_1_4_4_n19), .S(npu_inst_pe_1_4_4_n8), .Z(
        npu_inst_int_data_x_4__4__1_) );
  MUX2_X1 npu_inst_pe_1_4_4_U151 ( .A(npu_inst_pe_1_4_4_n21), .B(
        npu_inst_pe_1_4_4_n20), .S(npu_inst_pe_1_4_4_n6), .Z(
        npu_inst_pe_1_4_4_n22) );
  MUX2_X1 npu_inst_pe_1_4_4_U150 ( .A(npu_inst_pe_1_4_4_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_4_4_int_q_reg_h_1__1_), .S(npu_inst_pe_1_4_4_n4), .Z(
        npu_inst_pe_1_4_4_n21) );
  MUX2_X1 npu_inst_pe_1_4_4_U149 ( .A(npu_inst_pe_1_4_4_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_4_4_int_q_reg_h_3__1_), .S(npu_inst_pe_1_4_4_n4), .Z(
        npu_inst_pe_1_4_4_n20) );
  MUX2_X1 npu_inst_pe_1_4_4_U148 ( .A(npu_inst_pe_1_4_4_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_4_4_int_q_reg_h_5__1_), .S(npu_inst_pe_1_4_4_n4), .Z(
        npu_inst_pe_1_4_4_n19) );
  MUX2_X1 npu_inst_pe_1_4_4_U147 ( .A(npu_inst_pe_1_4_4_n18), .B(
        npu_inst_pe_1_4_4_n15), .S(npu_inst_pe_1_4_4_n8), .Z(
        npu_inst_int_data_x_4__4__0_) );
  MUX2_X1 npu_inst_pe_1_4_4_U146 ( .A(npu_inst_pe_1_4_4_n17), .B(
        npu_inst_pe_1_4_4_n16), .S(npu_inst_pe_1_4_4_n6), .Z(
        npu_inst_pe_1_4_4_n18) );
  MUX2_X1 npu_inst_pe_1_4_4_U145 ( .A(npu_inst_pe_1_4_4_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_4_4_int_q_reg_h_1__0_), .S(npu_inst_pe_1_4_4_n4), .Z(
        npu_inst_pe_1_4_4_n17) );
  MUX2_X1 npu_inst_pe_1_4_4_U144 ( .A(npu_inst_pe_1_4_4_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_4_4_int_q_reg_h_3__0_), .S(npu_inst_pe_1_4_4_n4), .Z(
        npu_inst_pe_1_4_4_n16) );
  MUX2_X1 npu_inst_pe_1_4_4_U143 ( .A(npu_inst_pe_1_4_4_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_4_4_int_q_reg_h_5__0_), .S(npu_inst_pe_1_4_4_n4), .Z(
        npu_inst_pe_1_4_4_n15) );
  XOR2_X1 npu_inst_pe_1_4_4_U142 ( .A(npu_inst_pe_1_4_4_int_data_0_), .B(
        npu_inst_pe_1_4_4_int_q_acc_0_), .Z(npu_inst_pe_1_4_4_N73) );
  AND2_X1 npu_inst_pe_1_4_4_U141 ( .A1(npu_inst_pe_1_4_4_int_q_acc_0_), .A2(
        npu_inst_pe_1_4_4_int_data_0_), .ZN(npu_inst_pe_1_4_4_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_4_4_U140 ( .A(npu_inst_pe_1_4_4_int_q_acc_0_), .B(
        npu_inst_pe_1_4_4_n13), .ZN(npu_inst_pe_1_4_4_N65) );
  OR2_X1 npu_inst_pe_1_4_4_U139 ( .A1(npu_inst_pe_1_4_4_n13), .A2(
        npu_inst_pe_1_4_4_int_q_acc_0_), .ZN(npu_inst_pe_1_4_4_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_4_4_U138 ( .A(npu_inst_pe_1_4_4_int_q_acc_2_), .B(
        npu_inst_pe_1_4_4_add_79_carry_2_), .Z(npu_inst_pe_1_4_4_N75) );
  AND2_X1 npu_inst_pe_1_4_4_U137 ( .A1(npu_inst_pe_1_4_4_add_79_carry_2_), 
        .A2(npu_inst_pe_1_4_4_int_q_acc_2_), .ZN(
        npu_inst_pe_1_4_4_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_4_4_U136 ( .A(npu_inst_pe_1_4_4_int_q_acc_3_), .B(
        npu_inst_pe_1_4_4_add_79_carry_3_), .Z(npu_inst_pe_1_4_4_N76) );
  AND2_X1 npu_inst_pe_1_4_4_U135 ( .A1(npu_inst_pe_1_4_4_add_79_carry_3_), 
        .A2(npu_inst_pe_1_4_4_int_q_acc_3_), .ZN(
        npu_inst_pe_1_4_4_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_4_4_U134 ( .A(npu_inst_pe_1_4_4_int_q_acc_4_), .B(
        npu_inst_pe_1_4_4_add_79_carry_4_), .Z(npu_inst_pe_1_4_4_N77) );
  AND2_X1 npu_inst_pe_1_4_4_U133 ( .A1(npu_inst_pe_1_4_4_add_79_carry_4_), 
        .A2(npu_inst_pe_1_4_4_int_q_acc_4_), .ZN(
        npu_inst_pe_1_4_4_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_4_4_U132 ( .A(npu_inst_pe_1_4_4_int_q_acc_5_), .B(
        npu_inst_pe_1_4_4_add_79_carry_5_), .Z(npu_inst_pe_1_4_4_N78) );
  AND2_X1 npu_inst_pe_1_4_4_U131 ( .A1(npu_inst_pe_1_4_4_add_79_carry_5_), 
        .A2(npu_inst_pe_1_4_4_int_q_acc_5_), .ZN(
        npu_inst_pe_1_4_4_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_4_4_U130 ( .A(npu_inst_pe_1_4_4_int_q_acc_6_), .B(
        npu_inst_pe_1_4_4_add_79_carry_6_), .Z(npu_inst_pe_1_4_4_N79) );
  AND2_X1 npu_inst_pe_1_4_4_U129 ( .A1(npu_inst_pe_1_4_4_add_79_carry_6_), 
        .A2(npu_inst_pe_1_4_4_int_q_acc_6_), .ZN(
        npu_inst_pe_1_4_4_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_4_4_U128 ( .A(npu_inst_pe_1_4_4_int_q_acc_7_), .B(
        npu_inst_pe_1_4_4_add_79_carry_7_), .Z(npu_inst_pe_1_4_4_N80) );
  XNOR2_X1 npu_inst_pe_1_4_4_U127 ( .A(npu_inst_pe_1_4_4_sub_77_carry_2_), .B(
        npu_inst_pe_1_4_4_int_q_acc_2_), .ZN(npu_inst_pe_1_4_4_N67) );
  OR2_X1 npu_inst_pe_1_4_4_U126 ( .A1(npu_inst_pe_1_4_4_int_q_acc_2_), .A2(
        npu_inst_pe_1_4_4_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_4_4_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_4_4_U125 ( .A(npu_inst_pe_1_4_4_sub_77_carry_3_), .B(
        npu_inst_pe_1_4_4_int_q_acc_3_), .ZN(npu_inst_pe_1_4_4_N68) );
  OR2_X1 npu_inst_pe_1_4_4_U124 ( .A1(npu_inst_pe_1_4_4_int_q_acc_3_), .A2(
        npu_inst_pe_1_4_4_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_4_4_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_4_4_U123 ( .A(npu_inst_pe_1_4_4_sub_77_carry_4_), .B(
        npu_inst_pe_1_4_4_int_q_acc_4_), .ZN(npu_inst_pe_1_4_4_N69) );
  OR2_X1 npu_inst_pe_1_4_4_U122 ( .A1(npu_inst_pe_1_4_4_int_q_acc_4_), .A2(
        npu_inst_pe_1_4_4_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_4_4_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_4_4_U121 ( .A(npu_inst_pe_1_4_4_sub_77_carry_5_), .B(
        npu_inst_pe_1_4_4_int_q_acc_5_), .ZN(npu_inst_pe_1_4_4_N70) );
  OR2_X1 npu_inst_pe_1_4_4_U120 ( .A1(npu_inst_pe_1_4_4_int_q_acc_5_), .A2(
        npu_inst_pe_1_4_4_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_4_4_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_4_4_U119 ( .A(npu_inst_pe_1_4_4_sub_77_carry_6_), .B(
        npu_inst_pe_1_4_4_int_q_acc_6_), .ZN(npu_inst_pe_1_4_4_N71) );
  OR2_X1 npu_inst_pe_1_4_4_U118 ( .A1(npu_inst_pe_1_4_4_int_q_acc_6_), .A2(
        npu_inst_pe_1_4_4_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_4_4_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_4_4_U117 ( .A(npu_inst_pe_1_4_4_int_q_acc_7_), .B(
        npu_inst_pe_1_4_4_sub_77_carry_7_), .ZN(npu_inst_pe_1_4_4_N72) );
  INV_X1 npu_inst_pe_1_4_4_U116 ( .A(npu_inst_n77), .ZN(npu_inst_pe_1_4_4_n7)
         );
  INV_X1 npu_inst_pe_1_4_4_U115 ( .A(npu_inst_pe_1_4_4_n7), .ZN(
        npu_inst_pe_1_4_4_n6) );
  INV_X1 npu_inst_pe_1_4_4_U114 ( .A(npu_inst_n55), .ZN(npu_inst_pe_1_4_4_n3)
         );
  AOI22_X1 npu_inst_pe_1_4_4_U113 ( .A1(npu_inst_int_data_y_5__4__0_), .A2(
        npu_inst_pe_1_4_4_n58), .B1(npu_inst_pe_1_4_4_n114), .B2(
        npu_inst_pe_1_4_4_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_4_4_n57) );
  INV_X1 npu_inst_pe_1_4_4_U112 ( .A(npu_inst_pe_1_4_4_n57), .ZN(
        npu_inst_pe_1_4_4_n108) );
  AOI22_X1 npu_inst_pe_1_4_4_U111 ( .A1(npu_inst_int_data_y_5__4__0_), .A2(
        npu_inst_pe_1_4_4_n54), .B1(npu_inst_pe_1_4_4_n115), .B2(
        npu_inst_pe_1_4_4_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_4_4_n53) );
  INV_X1 npu_inst_pe_1_4_4_U110 ( .A(npu_inst_pe_1_4_4_n53), .ZN(
        npu_inst_pe_1_4_4_n109) );
  AOI22_X1 npu_inst_pe_1_4_4_U107 ( .A1(npu_inst_int_data_y_5__4__0_), .A2(
        npu_inst_pe_1_4_4_n50), .B1(npu_inst_pe_1_4_4_n116), .B2(
        npu_inst_pe_1_4_4_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_4_4_n49) );
  INV_X1 npu_inst_pe_1_4_4_U106 ( .A(npu_inst_pe_1_4_4_n49), .ZN(
        npu_inst_pe_1_4_4_n110) );
  AOI22_X1 npu_inst_pe_1_4_4_U105 ( .A1(npu_inst_int_data_y_5__4__0_), .A2(
        npu_inst_pe_1_4_4_n46), .B1(npu_inst_pe_1_4_4_n117), .B2(
        npu_inst_pe_1_4_4_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_4_4_n45) );
  INV_X1 npu_inst_pe_1_4_4_U104 ( .A(npu_inst_pe_1_4_4_n45), .ZN(
        npu_inst_pe_1_4_4_n111) );
  AOI22_X1 npu_inst_pe_1_4_4_U103 ( .A1(npu_inst_int_data_y_5__4__0_), .A2(
        npu_inst_pe_1_4_4_n42), .B1(npu_inst_pe_1_4_4_n119), .B2(
        npu_inst_pe_1_4_4_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_4_4_n41) );
  INV_X1 npu_inst_pe_1_4_4_U102 ( .A(npu_inst_pe_1_4_4_n41), .ZN(
        npu_inst_pe_1_4_4_n112) );
  AOI22_X1 npu_inst_pe_1_4_4_U101 ( .A1(npu_inst_int_data_y_5__4__1_), .A2(
        npu_inst_pe_1_4_4_n58), .B1(npu_inst_pe_1_4_4_n114), .B2(
        npu_inst_pe_1_4_4_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_4_4_n59) );
  INV_X1 npu_inst_pe_1_4_4_U100 ( .A(npu_inst_pe_1_4_4_n59), .ZN(
        npu_inst_pe_1_4_4_n102) );
  AOI22_X1 npu_inst_pe_1_4_4_U99 ( .A1(npu_inst_int_data_y_5__4__1_), .A2(
        npu_inst_pe_1_4_4_n54), .B1(npu_inst_pe_1_4_4_n115), .B2(
        npu_inst_pe_1_4_4_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_4_4_n55) );
  INV_X1 npu_inst_pe_1_4_4_U98 ( .A(npu_inst_pe_1_4_4_n55), .ZN(
        npu_inst_pe_1_4_4_n103) );
  AOI22_X1 npu_inst_pe_1_4_4_U97 ( .A1(npu_inst_int_data_y_5__4__1_), .A2(
        npu_inst_pe_1_4_4_n50), .B1(npu_inst_pe_1_4_4_n116), .B2(
        npu_inst_pe_1_4_4_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_4_4_n51) );
  INV_X1 npu_inst_pe_1_4_4_U96 ( .A(npu_inst_pe_1_4_4_n51), .ZN(
        npu_inst_pe_1_4_4_n104) );
  AOI22_X1 npu_inst_pe_1_4_4_U95 ( .A1(npu_inst_int_data_y_5__4__1_), .A2(
        npu_inst_pe_1_4_4_n46), .B1(npu_inst_pe_1_4_4_n117), .B2(
        npu_inst_pe_1_4_4_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_4_4_n47) );
  INV_X1 npu_inst_pe_1_4_4_U94 ( .A(npu_inst_pe_1_4_4_n47), .ZN(
        npu_inst_pe_1_4_4_n105) );
  AOI22_X1 npu_inst_pe_1_4_4_U93 ( .A1(npu_inst_int_data_y_5__4__1_), .A2(
        npu_inst_pe_1_4_4_n42), .B1(npu_inst_pe_1_4_4_n119), .B2(
        npu_inst_pe_1_4_4_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_4_4_n43) );
  INV_X1 npu_inst_pe_1_4_4_U92 ( .A(npu_inst_pe_1_4_4_n43), .ZN(
        npu_inst_pe_1_4_4_n106) );
  AOI22_X1 npu_inst_pe_1_4_4_U91 ( .A1(npu_inst_pe_1_4_4_n38), .A2(
        npu_inst_int_data_y_5__4__1_), .B1(npu_inst_pe_1_4_4_n118), .B2(
        npu_inst_pe_1_4_4_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_4_4_n39) );
  INV_X1 npu_inst_pe_1_4_4_U90 ( .A(npu_inst_pe_1_4_4_n39), .ZN(
        npu_inst_pe_1_4_4_n107) );
  AOI22_X1 npu_inst_pe_1_4_4_U89 ( .A1(npu_inst_pe_1_4_4_n38), .A2(
        npu_inst_int_data_y_5__4__0_), .B1(npu_inst_pe_1_4_4_n118), .B2(
        npu_inst_pe_1_4_4_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_4_4_n37) );
  INV_X1 npu_inst_pe_1_4_4_U88 ( .A(npu_inst_pe_1_4_4_n37), .ZN(
        npu_inst_pe_1_4_4_n113) );
  NOR3_X1 npu_inst_pe_1_4_4_U87 ( .A1(npu_inst_pe_1_4_4_n26), .A2(npu_inst_n55), .A3(npu_inst_int_ckg[27]), .ZN(npu_inst_pe_1_4_4_n85) );
  OR2_X1 npu_inst_pe_1_4_4_U86 ( .A1(npu_inst_pe_1_4_4_n85), .A2(
        npu_inst_pe_1_4_4_n2), .ZN(npu_inst_pe_1_4_4_N84) );
  NAND2_X1 npu_inst_pe_1_4_4_U85 ( .A1(npu_inst_pe_1_4_4_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_4_4_n60), .ZN(npu_inst_pe_1_4_4_n74) );
  OAI21_X1 npu_inst_pe_1_4_4_U84 ( .B1(npu_inst_pe_1_4_4_n63), .B2(
        npu_inst_pe_1_4_4_n60), .A(npu_inst_pe_1_4_4_n74), .ZN(
        npu_inst_pe_1_4_4_n97) );
  NAND2_X1 npu_inst_pe_1_4_4_U83 ( .A1(npu_inst_pe_1_4_4_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_4_4_n60), .ZN(npu_inst_pe_1_4_4_n73) );
  OAI21_X1 npu_inst_pe_1_4_4_U82 ( .B1(npu_inst_pe_1_4_4_n61), .B2(
        npu_inst_pe_1_4_4_n60), .A(npu_inst_pe_1_4_4_n73), .ZN(
        npu_inst_pe_1_4_4_n96) );
  NAND2_X1 npu_inst_pe_1_4_4_U81 ( .A1(npu_inst_pe_1_4_4_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_4_4_n56), .ZN(npu_inst_pe_1_4_4_n72) );
  OAI21_X1 npu_inst_pe_1_4_4_U80 ( .B1(npu_inst_pe_1_4_4_n63), .B2(
        npu_inst_pe_1_4_4_n56), .A(npu_inst_pe_1_4_4_n72), .ZN(
        npu_inst_pe_1_4_4_n95) );
  NAND2_X1 npu_inst_pe_1_4_4_U79 ( .A1(npu_inst_pe_1_4_4_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_4_4_n56), .ZN(npu_inst_pe_1_4_4_n71) );
  OAI21_X1 npu_inst_pe_1_4_4_U78 ( .B1(npu_inst_pe_1_4_4_n61), .B2(
        npu_inst_pe_1_4_4_n56), .A(npu_inst_pe_1_4_4_n71), .ZN(
        npu_inst_pe_1_4_4_n94) );
  NAND2_X1 npu_inst_pe_1_4_4_U77 ( .A1(npu_inst_pe_1_4_4_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_4_4_n52), .ZN(npu_inst_pe_1_4_4_n70) );
  OAI21_X1 npu_inst_pe_1_4_4_U76 ( .B1(npu_inst_pe_1_4_4_n63), .B2(
        npu_inst_pe_1_4_4_n52), .A(npu_inst_pe_1_4_4_n70), .ZN(
        npu_inst_pe_1_4_4_n93) );
  NAND2_X1 npu_inst_pe_1_4_4_U75 ( .A1(npu_inst_pe_1_4_4_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_4_4_n52), .ZN(npu_inst_pe_1_4_4_n69) );
  OAI21_X1 npu_inst_pe_1_4_4_U74 ( .B1(npu_inst_pe_1_4_4_n61), .B2(
        npu_inst_pe_1_4_4_n52), .A(npu_inst_pe_1_4_4_n69), .ZN(
        npu_inst_pe_1_4_4_n92) );
  NAND2_X1 npu_inst_pe_1_4_4_U73 ( .A1(npu_inst_pe_1_4_4_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_4_4_n48), .ZN(npu_inst_pe_1_4_4_n68) );
  OAI21_X1 npu_inst_pe_1_4_4_U72 ( .B1(npu_inst_pe_1_4_4_n63), .B2(
        npu_inst_pe_1_4_4_n48), .A(npu_inst_pe_1_4_4_n68), .ZN(
        npu_inst_pe_1_4_4_n91) );
  NAND2_X1 npu_inst_pe_1_4_4_U71 ( .A1(npu_inst_pe_1_4_4_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_4_4_n48), .ZN(npu_inst_pe_1_4_4_n67) );
  OAI21_X1 npu_inst_pe_1_4_4_U70 ( .B1(npu_inst_pe_1_4_4_n61), .B2(
        npu_inst_pe_1_4_4_n48), .A(npu_inst_pe_1_4_4_n67), .ZN(
        npu_inst_pe_1_4_4_n90) );
  NAND2_X1 npu_inst_pe_1_4_4_U69 ( .A1(npu_inst_pe_1_4_4_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_4_4_n44), .ZN(npu_inst_pe_1_4_4_n66) );
  OAI21_X1 npu_inst_pe_1_4_4_U68 ( .B1(npu_inst_pe_1_4_4_n63), .B2(
        npu_inst_pe_1_4_4_n44), .A(npu_inst_pe_1_4_4_n66), .ZN(
        npu_inst_pe_1_4_4_n89) );
  NAND2_X1 npu_inst_pe_1_4_4_U67 ( .A1(npu_inst_pe_1_4_4_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_4_4_n44), .ZN(npu_inst_pe_1_4_4_n65) );
  OAI21_X1 npu_inst_pe_1_4_4_U66 ( .B1(npu_inst_pe_1_4_4_n61), .B2(
        npu_inst_pe_1_4_4_n44), .A(npu_inst_pe_1_4_4_n65), .ZN(
        npu_inst_pe_1_4_4_n88) );
  NAND2_X1 npu_inst_pe_1_4_4_U65 ( .A1(npu_inst_pe_1_4_4_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_4_4_n40), .ZN(npu_inst_pe_1_4_4_n64) );
  OAI21_X1 npu_inst_pe_1_4_4_U64 ( .B1(npu_inst_pe_1_4_4_n63), .B2(
        npu_inst_pe_1_4_4_n40), .A(npu_inst_pe_1_4_4_n64), .ZN(
        npu_inst_pe_1_4_4_n87) );
  NAND2_X1 npu_inst_pe_1_4_4_U63 ( .A1(npu_inst_pe_1_4_4_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_4_4_n40), .ZN(npu_inst_pe_1_4_4_n62) );
  OAI21_X1 npu_inst_pe_1_4_4_U62 ( .B1(npu_inst_pe_1_4_4_n61), .B2(
        npu_inst_pe_1_4_4_n40), .A(npu_inst_pe_1_4_4_n62), .ZN(
        npu_inst_pe_1_4_4_n86) );
  AND2_X1 npu_inst_pe_1_4_4_U61 ( .A1(npu_inst_pe_1_4_4_N93), .A2(npu_inst_n55), .ZN(npu_inst_int_data_y_4__4__0_) );
  AND2_X1 npu_inst_pe_1_4_4_U60 ( .A1(npu_inst_n55), .A2(npu_inst_pe_1_4_4_N94), .ZN(npu_inst_int_data_y_4__4__1_) );
  AND2_X1 npu_inst_pe_1_4_4_U59 ( .A1(npu_inst_pe_1_4_4_int_q_acc_0_), .A2(
        npu_inst_pe_1_4_4_n1), .ZN(npu_inst_int_data_res_4__4__0_) );
  AND2_X1 npu_inst_pe_1_4_4_U58 ( .A1(npu_inst_pe_1_4_4_n2), .A2(
        npu_inst_pe_1_4_4_int_q_acc_7_), .ZN(npu_inst_int_data_res_4__4__7_)
         );
  AND2_X1 npu_inst_pe_1_4_4_U57 ( .A1(npu_inst_pe_1_4_4_int_q_acc_1_), .A2(
        npu_inst_pe_1_4_4_n1), .ZN(npu_inst_int_data_res_4__4__1_) );
  AND2_X1 npu_inst_pe_1_4_4_U56 ( .A1(npu_inst_pe_1_4_4_int_q_acc_2_), .A2(
        npu_inst_pe_1_4_4_n1), .ZN(npu_inst_int_data_res_4__4__2_) );
  AND2_X1 npu_inst_pe_1_4_4_U55 ( .A1(npu_inst_pe_1_4_4_int_q_acc_3_), .A2(
        npu_inst_pe_1_4_4_n2), .ZN(npu_inst_int_data_res_4__4__3_) );
  AND2_X1 npu_inst_pe_1_4_4_U54 ( .A1(npu_inst_pe_1_4_4_int_q_acc_4_), .A2(
        npu_inst_pe_1_4_4_n2), .ZN(npu_inst_int_data_res_4__4__4_) );
  AND2_X1 npu_inst_pe_1_4_4_U53 ( .A1(npu_inst_pe_1_4_4_int_q_acc_5_), .A2(
        npu_inst_pe_1_4_4_n2), .ZN(npu_inst_int_data_res_4__4__5_) );
  AND2_X1 npu_inst_pe_1_4_4_U52 ( .A1(npu_inst_pe_1_4_4_int_q_acc_6_), .A2(
        npu_inst_pe_1_4_4_n2), .ZN(npu_inst_int_data_res_4__4__6_) );
  AOI222_X1 npu_inst_pe_1_4_4_U51 ( .A1(npu_inst_int_data_res_5__4__0_), .A2(
        npu_inst_pe_1_4_4_n1), .B1(npu_inst_pe_1_4_4_N73), .B2(
        npu_inst_pe_1_4_4_n76), .C1(npu_inst_pe_1_4_4_N65), .C2(
        npu_inst_pe_1_4_4_n77), .ZN(npu_inst_pe_1_4_4_n84) );
  INV_X1 npu_inst_pe_1_4_4_U50 ( .A(npu_inst_pe_1_4_4_n84), .ZN(
        npu_inst_pe_1_4_4_n101) );
  AOI222_X1 npu_inst_pe_1_4_4_U49 ( .A1(npu_inst_int_data_res_5__4__7_), .A2(
        npu_inst_pe_1_4_4_n1), .B1(npu_inst_pe_1_4_4_N80), .B2(
        npu_inst_pe_1_4_4_n76), .C1(npu_inst_pe_1_4_4_N72), .C2(
        npu_inst_pe_1_4_4_n77), .ZN(npu_inst_pe_1_4_4_n75) );
  INV_X1 npu_inst_pe_1_4_4_U48 ( .A(npu_inst_pe_1_4_4_n75), .ZN(
        npu_inst_pe_1_4_4_n33) );
  AOI222_X1 npu_inst_pe_1_4_4_U47 ( .A1(npu_inst_int_data_res_5__4__1_), .A2(
        npu_inst_pe_1_4_4_n1), .B1(npu_inst_pe_1_4_4_N74), .B2(
        npu_inst_pe_1_4_4_n76), .C1(npu_inst_pe_1_4_4_N66), .C2(
        npu_inst_pe_1_4_4_n77), .ZN(npu_inst_pe_1_4_4_n83) );
  INV_X1 npu_inst_pe_1_4_4_U46 ( .A(npu_inst_pe_1_4_4_n83), .ZN(
        npu_inst_pe_1_4_4_n100) );
  AOI222_X1 npu_inst_pe_1_4_4_U45 ( .A1(npu_inst_int_data_res_5__4__2_), .A2(
        npu_inst_pe_1_4_4_n1), .B1(npu_inst_pe_1_4_4_N75), .B2(
        npu_inst_pe_1_4_4_n76), .C1(npu_inst_pe_1_4_4_N67), .C2(
        npu_inst_pe_1_4_4_n77), .ZN(npu_inst_pe_1_4_4_n82) );
  INV_X1 npu_inst_pe_1_4_4_U44 ( .A(npu_inst_pe_1_4_4_n82), .ZN(
        npu_inst_pe_1_4_4_n99) );
  AOI222_X1 npu_inst_pe_1_4_4_U43 ( .A1(npu_inst_int_data_res_5__4__3_), .A2(
        npu_inst_pe_1_4_4_n1), .B1(npu_inst_pe_1_4_4_N76), .B2(
        npu_inst_pe_1_4_4_n76), .C1(npu_inst_pe_1_4_4_N68), .C2(
        npu_inst_pe_1_4_4_n77), .ZN(npu_inst_pe_1_4_4_n81) );
  INV_X1 npu_inst_pe_1_4_4_U42 ( .A(npu_inst_pe_1_4_4_n81), .ZN(
        npu_inst_pe_1_4_4_n98) );
  AOI222_X1 npu_inst_pe_1_4_4_U41 ( .A1(npu_inst_int_data_res_5__4__4_), .A2(
        npu_inst_pe_1_4_4_n1), .B1(npu_inst_pe_1_4_4_N77), .B2(
        npu_inst_pe_1_4_4_n76), .C1(npu_inst_pe_1_4_4_N69), .C2(
        npu_inst_pe_1_4_4_n77), .ZN(npu_inst_pe_1_4_4_n80) );
  INV_X1 npu_inst_pe_1_4_4_U40 ( .A(npu_inst_pe_1_4_4_n80), .ZN(
        npu_inst_pe_1_4_4_n36) );
  AOI222_X1 npu_inst_pe_1_4_4_U39 ( .A1(npu_inst_int_data_res_5__4__5_), .A2(
        npu_inst_pe_1_4_4_n1), .B1(npu_inst_pe_1_4_4_N78), .B2(
        npu_inst_pe_1_4_4_n76), .C1(npu_inst_pe_1_4_4_N70), .C2(
        npu_inst_pe_1_4_4_n77), .ZN(npu_inst_pe_1_4_4_n79) );
  INV_X1 npu_inst_pe_1_4_4_U38 ( .A(npu_inst_pe_1_4_4_n79), .ZN(
        npu_inst_pe_1_4_4_n35) );
  AOI222_X1 npu_inst_pe_1_4_4_U37 ( .A1(npu_inst_int_data_res_5__4__6_), .A2(
        npu_inst_pe_1_4_4_n1), .B1(npu_inst_pe_1_4_4_N79), .B2(
        npu_inst_pe_1_4_4_n76), .C1(npu_inst_pe_1_4_4_N71), .C2(
        npu_inst_pe_1_4_4_n77), .ZN(npu_inst_pe_1_4_4_n78) );
  INV_X1 npu_inst_pe_1_4_4_U36 ( .A(npu_inst_pe_1_4_4_n78), .ZN(
        npu_inst_pe_1_4_4_n34) );
  INV_X1 npu_inst_pe_1_4_4_U35 ( .A(npu_inst_pe_1_4_4_int_data_1_), .ZN(
        npu_inst_pe_1_4_4_n14) );
  AND2_X1 npu_inst_pe_1_4_4_U34 ( .A1(npu_inst_int_data_x_4__4__1_), .A2(
        npu_inst_pe_1_4_4_int_q_weight_1_), .ZN(npu_inst_pe_1_4_4_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_4_4_U33 ( .A1(npu_inst_int_data_x_4__4__0_), .A2(
        npu_inst_pe_1_4_4_int_q_weight_1_), .ZN(npu_inst_pe_1_4_4_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_4_4_U32 ( .A1(npu_inst_n55), .A2(
        npu_inst_int_data_y_5__4__1_), .B1(npu_inst_pe_1_4_4_n3), .B2(
        npu_inst_int_data_x_4__5__1_), .ZN(npu_inst_pe_1_4_4_n63) );
  AOI22_X1 npu_inst_pe_1_4_4_U31 ( .A1(npu_inst_n55), .A2(
        npu_inst_int_data_y_5__4__0_), .B1(npu_inst_pe_1_4_4_n3), .B2(
        npu_inst_int_data_x_4__5__0_), .ZN(npu_inst_pe_1_4_4_n61) );
  INV_X1 npu_inst_pe_1_4_4_U30 ( .A(npu_inst_pe_1_4_4_int_data_0_), .ZN(
        npu_inst_pe_1_4_4_n13) );
  INV_X1 npu_inst_pe_1_4_4_U29 ( .A(npu_inst_n69), .ZN(npu_inst_pe_1_4_4_n5)
         );
  OR3_X1 npu_inst_pe_1_4_4_U28 ( .A1(npu_inst_pe_1_4_4_n6), .A2(
        npu_inst_pe_1_4_4_n8), .A3(npu_inst_pe_1_4_4_n5), .ZN(
        npu_inst_pe_1_4_4_n56) );
  OR3_X1 npu_inst_pe_1_4_4_U27 ( .A1(npu_inst_pe_1_4_4_n5), .A2(
        npu_inst_pe_1_4_4_n8), .A3(npu_inst_pe_1_4_4_n7), .ZN(
        npu_inst_pe_1_4_4_n48) );
  INV_X1 npu_inst_pe_1_4_4_U26 ( .A(npu_inst_pe_1_4_4_n5), .ZN(
        npu_inst_pe_1_4_4_n4) );
  INV_X1 npu_inst_pe_1_4_4_U25 ( .A(npu_inst_n124), .ZN(npu_inst_pe_1_4_4_n12)
         );
  OR3_X1 npu_inst_pe_1_4_4_U24 ( .A1(npu_inst_pe_1_4_4_n4), .A2(
        npu_inst_pe_1_4_4_n8), .A3(npu_inst_pe_1_4_4_n7), .ZN(
        npu_inst_pe_1_4_4_n52) );
  OR3_X1 npu_inst_pe_1_4_4_U23 ( .A1(npu_inst_pe_1_4_4_n6), .A2(
        npu_inst_pe_1_4_4_n8), .A3(npu_inst_pe_1_4_4_n4), .ZN(
        npu_inst_pe_1_4_4_n60) );
  NOR2_X1 npu_inst_pe_1_4_4_U22 ( .A1(npu_inst_pe_1_4_4_n60), .A2(
        npu_inst_pe_1_4_4_n3), .ZN(npu_inst_pe_1_4_4_n58) );
  NOR2_X1 npu_inst_pe_1_4_4_U21 ( .A1(npu_inst_pe_1_4_4_n56), .A2(
        npu_inst_pe_1_4_4_n3), .ZN(npu_inst_pe_1_4_4_n54) );
  NOR2_X1 npu_inst_pe_1_4_4_U20 ( .A1(npu_inst_pe_1_4_4_n52), .A2(
        npu_inst_pe_1_4_4_n3), .ZN(npu_inst_pe_1_4_4_n50) );
  NOR2_X1 npu_inst_pe_1_4_4_U19 ( .A1(npu_inst_pe_1_4_4_n48), .A2(
        npu_inst_pe_1_4_4_n3), .ZN(npu_inst_pe_1_4_4_n46) );
  NOR2_X1 npu_inst_pe_1_4_4_U18 ( .A1(npu_inst_pe_1_4_4_n40), .A2(
        npu_inst_pe_1_4_4_n3), .ZN(npu_inst_pe_1_4_4_n38) );
  NOR2_X1 npu_inst_pe_1_4_4_U17 ( .A1(npu_inst_pe_1_4_4_n44), .A2(
        npu_inst_pe_1_4_4_n3), .ZN(npu_inst_pe_1_4_4_n42) );
  BUF_X1 npu_inst_pe_1_4_4_U16 ( .A(npu_inst_n98), .Z(npu_inst_pe_1_4_4_n8) );
  BUF_X1 npu_inst_pe_1_4_4_U15 ( .A(npu_inst_pe_1_4_4_n12), .Z(
        npu_inst_pe_1_4_4_n11) );
  BUF_X1 npu_inst_pe_1_4_4_U14 ( .A(npu_inst_pe_1_4_4_n12), .Z(
        npu_inst_pe_1_4_4_n10) );
  BUF_X1 npu_inst_pe_1_4_4_U13 ( .A(npu_inst_pe_1_4_4_n12), .Z(
        npu_inst_pe_1_4_4_n9) );
  INV_X1 npu_inst_pe_1_4_4_U12 ( .A(npu_inst_pe_1_4_4_n38), .ZN(
        npu_inst_pe_1_4_4_n118) );
  INV_X1 npu_inst_pe_1_4_4_U11 ( .A(npu_inst_pe_1_4_4_n58), .ZN(
        npu_inst_pe_1_4_4_n114) );
  INV_X1 npu_inst_pe_1_4_4_U10 ( .A(npu_inst_pe_1_4_4_n54), .ZN(
        npu_inst_pe_1_4_4_n115) );
  INV_X1 npu_inst_pe_1_4_4_U9 ( .A(npu_inst_pe_1_4_4_n50), .ZN(
        npu_inst_pe_1_4_4_n116) );
  INV_X1 npu_inst_pe_1_4_4_U8 ( .A(npu_inst_pe_1_4_4_n46), .ZN(
        npu_inst_pe_1_4_4_n117) );
  INV_X1 npu_inst_pe_1_4_4_U7 ( .A(npu_inst_pe_1_4_4_n42), .ZN(
        npu_inst_pe_1_4_4_n119) );
  BUF_X1 npu_inst_pe_1_4_4_U6 ( .A(npu_inst_n20), .Z(npu_inst_pe_1_4_4_n2) );
  BUF_X1 npu_inst_pe_1_4_4_U5 ( .A(npu_inst_n20), .Z(npu_inst_pe_1_4_4_n1) );
  NOR2_X1 npu_inst_pe_1_4_4_U4 ( .A1(npu_inst_pe_1_4_4_int_q_weight_0_), .A2(
        npu_inst_pe_1_4_4_n1), .ZN(npu_inst_pe_1_4_4_n76) );
  NOR2_X1 npu_inst_pe_1_4_4_U3 ( .A1(npu_inst_pe_1_4_4_n27), .A2(
        npu_inst_pe_1_4_4_n1), .ZN(npu_inst_pe_1_4_4_n77) );
  FA_X1 npu_inst_pe_1_4_4_sub_77_U2_1 ( .A(npu_inst_pe_1_4_4_int_q_acc_1_), 
        .B(npu_inst_pe_1_4_4_n14), .CI(npu_inst_pe_1_4_4_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_4_4_sub_77_carry_2_), .S(npu_inst_pe_1_4_4_N66) );
  FA_X1 npu_inst_pe_1_4_4_add_79_U1_1 ( .A(npu_inst_pe_1_4_4_int_q_acc_1_), 
        .B(npu_inst_pe_1_4_4_int_data_1_), .CI(
        npu_inst_pe_1_4_4_add_79_carry_1_), .CO(
        npu_inst_pe_1_4_4_add_79_carry_2_), .S(npu_inst_pe_1_4_4_N74) );
  NAND3_X1 npu_inst_pe_1_4_4_U109 ( .A1(npu_inst_pe_1_4_4_n5), .A2(
        npu_inst_pe_1_4_4_n7), .A3(npu_inst_pe_1_4_4_n8), .ZN(
        npu_inst_pe_1_4_4_n44) );
  NAND3_X1 npu_inst_pe_1_4_4_U108 ( .A1(npu_inst_pe_1_4_4_n4), .A2(
        npu_inst_pe_1_4_4_n7), .A3(npu_inst_pe_1_4_4_n8), .ZN(
        npu_inst_pe_1_4_4_n40) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_4_4_n34), .CK(
        npu_inst_pe_1_4_4_net3465), .RN(npu_inst_pe_1_4_4_n9), .Q(
        npu_inst_pe_1_4_4_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_4_4_n35), .CK(
        npu_inst_pe_1_4_4_net3465), .RN(npu_inst_pe_1_4_4_n9), .Q(
        npu_inst_pe_1_4_4_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_4_4_n36), .CK(
        npu_inst_pe_1_4_4_net3465), .RN(npu_inst_pe_1_4_4_n9), .Q(
        npu_inst_pe_1_4_4_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_4_4_n98), .CK(
        npu_inst_pe_1_4_4_net3465), .RN(npu_inst_pe_1_4_4_n9), .Q(
        npu_inst_pe_1_4_4_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_4_4_n99), .CK(
        npu_inst_pe_1_4_4_net3465), .RN(npu_inst_pe_1_4_4_n9), .Q(
        npu_inst_pe_1_4_4_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_4_4_n100), 
        .CK(npu_inst_pe_1_4_4_net3465), .RN(npu_inst_pe_1_4_4_n9), .Q(
        npu_inst_pe_1_4_4_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_4_4_n33), .CK(
        npu_inst_pe_1_4_4_net3465), .RN(npu_inst_pe_1_4_4_n9), .Q(
        npu_inst_pe_1_4_4_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_4_4_n101), 
        .CK(npu_inst_pe_1_4_4_net3465), .RN(npu_inst_pe_1_4_4_n9), .Q(
        npu_inst_pe_1_4_4_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_weight_reg_0_ ( .D(npu_inst_n110), .CK(
        npu_inst_pe_1_4_4_net3471), .RN(npu_inst_pe_1_4_4_n9), .Q(
        npu_inst_pe_1_4_4_int_q_weight_0_), .QN(npu_inst_pe_1_4_4_n27) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_weight_reg_1_ ( .D(npu_inst_n116), .CK(
        npu_inst_pe_1_4_4_net3471), .RN(npu_inst_pe_1_4_4_n9), .Q(
        npu_inst_pe_1_4_4_int_q_weight_1_), .QN(npu_inst_pe_1_4_4_n26) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_4_4_n113), 
        .CK(npu_inst_pe_1_4_4_net3471), .RN(npu_inst_pe_1_4_4_n9), .Q(
        npu_inst_pe_1_4_4_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_4_4_n107), 
        .CK(npu_inst_pe_1_4_4_net3471), .RN(npu_inst_pe_1_4_4_n9), .Q(
        npu_inst_pe_1_4_4_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_4_4_n112), 
        .CK(npu_inst_pe_1_4_4_net3471), .RN(npu_inst_pe_1_4_4_n10), .Q(
        npu_inst_pe_1_4_4_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_4_4_n106), 
        .CK(npu_inst_pe_1_4_4_net3471), .RN(npu_inst_pe_1_4_4_n10), .Q(
        npu_inst_pe_1_4_4_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_4_4_n111), 
        .CK(npu_inst_pe_1_4_4_net3471), .RN(npu_inst_pe_1_4_4_n10), .Q(
        npu_inst_pe_1_4_4_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_4_4_n105), 
        .CK(npu_inst_pe_1_4_4_net3471), .RN(npu_inst_pe_1_4_4_n10), .Q(
        npu_inst_pe_1_4_4_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_4_4_n110), 
        .CK(npu_inst_pe_1_4_4_net3471), .RN(npu_inst_pe_1_4_4_n10), .Q(
        npu_inst_pe_1_4_4_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_4_4_n104), 
        .CK(npu_inst_pe_1_4_4_net3471), .RN(npu_inst_pe_1_4_4_n10), .Q(
        npu_inst_pe_1_4_4_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_4_4_n109), 
        .CK(npu_inst_pe_1_4_4_net3471), .RN(npu_inst_pe_1_4_4_n10), .Q(
        npu_inst_pe_1_4_4_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_4_4_n103), 
        .CK(npu_inst_pe_1_4_4_net3471), .RN(npu_inst_pe_1_4_4_n10), .Q(
        npu_inst_pe_1_4_4_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_4_4_n108), 
        .CK(npu_inst_pe_1_4_4_net3471), .RN(npu_inst_pe_1_4_4_n10), .Q(
        npu_inst_pe_1_4_4_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_4_4_n102), 
        .CK(npu_inst_pe_1_4_4_net3471), .RN(npu_inst_pe_1_4_4_n10), .Q(
        npu_inst_pe_1_4_4_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_4_4_n86), 
        .CK(npu_inst_pe_1_4_4_net3471), .RN(npu_inst_pe_1_4_4_n10), .Q(
        npu_inst_pe_1_4_4_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_4_4_n87), 
        .CK(npu_inst_pe_1_4_4_net3471), .RN(npu_inst_pe_1_4_4_n10), .Q(
        npu_inst_pe_1_4_4_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_4_4_n88), 
        .CK(npu_inst_pe_1_4_4_net3471), .RN(npu_inst_pe_1_4_4_n11), .Q(
        npu_inst_pe_1_4_4_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_4_4_n89), 
        .CK(npu_inst_pe_1_4_4_net3471), .RN(npu_inst_pe_1_4_4_n11), .Q(
        npu_inst_pe_1_4_4_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_4_4_n90), 
        .CK(npu_inst_pe_1_4_4_net3471), .RN(npu_inst_pe_1_4_4_n11), .Q(
        npu_inst_pe_1_4_4_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_4_4_n91), 
        .CK(npu_inst_pe_1_4_4_net3471), .RN(npu_inst_pe_1_4_4_n11), .Q(
        npu_inst_pe_1_4_4_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_4_4_n92), 
        .CK(npu_inst_pe_1_4_4_net3471), .RN(npu_inst_pe_1_4_4_n11), .Q(
        npu_inst_pe_1_4_4_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_4_4_n93), 
        .CK(npu_inst_pe_1_4_4_net3471), .RN(npu_inst_pe_1_4_4_n11), .Q(
        npu_inst_pe_1_4_4_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_4_4_n94), 
        .CK(npu_inst_pe_1_4_4_net3471), .RN(npu_inst_pe_1_4_4_n11), .Q(
        npu_inst_pe_1_4_4_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_4_4_n95), 
        .CK(npu_inst_pe_1_4_4_net3471), .RN(npu_inst_pe_1_4_4_n11), .Q(
        npu_inst_pe_1_4_4_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_4_4_n96), 
        .CK(npu_inst_pe_1_4_4_net3471), .RN(npu_inst_pe_1_4_4_n11), .Q(
        npu_inst_pe_1_4_4_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_4_4_n97), 
        .CK(npu_inst_pe_1_4_4_net3471), .RN(npu_inst_pe_1_4_4_n11), .Q(
        npu_inst_pe_1_4_4_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_4_4_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_4_4_N84), .SE(1'b0), .GCK(npu_inst_pe_1_4_4_net3465) );
  CLKGATETST_X1 npu_inst_pe_1_4_4_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n63), .SE(1'b0), .GCK(npu_inst_pe_1_4_4_net3471) );
  MUX2_X1 npu_inst_pe_1_4_5_U162 ( .A(npu_inst_pe_1_4_5_n32), .B(
        npu_inst_pe_1_4_5_n29), .S(npu_inst_pe_1_4_5_n8), .Z(
        npu_inst_pe_1_4_5_N93) );
  MUX2_X1 npu_inst_pe_1_4_5_U161 ( .A(npu_inst_pe_1_4_5_n31), .B(
        npu_inst_pe_1_4_5_n30), .S(npu_inst_pe_1_4_5_n6), .Z(
        npu_inst_pe_1_4_5_n32) );
  MUX2_X1 npu_inst_pe_1_4_5_U160 ( .A(npu_inst_pe_1_4_5_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_4_5_int_q_reg_v_1__0_), .S(npu_inst_pe_1_4_5_n4), .Z(
        npu_inst_pe_1_4_5_n31) );
  MUX2_X1 npu_inst_pe_1_4_5_U159 ( .A(npu_inst_pe_1_4_5_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_4_5_int_q_reg_v_3__0_), .S(npu_inst_pe_1_4_5_n4), .Z(
        npu_inst_pe_1_4_5_n30) );
  MUX2_X1 npu_inst_pe_1_4_5_U158 ( .A(npu_inst_pe_1_4_5_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_4_5_int_q_reg_v_5__0_), .S(npu_inst_pe_1_4_5_n4), .Z(
        npu_inst_pe_1_4_5_n29) );
  MUX2_X1 npu_inst_pe_1_4_5_U157 ( .A(npu_inst_pe_1_4_5_n28), .B(
        npu_inst_pe_1_4_5_n23), .S(npu_inst_pe_1_4_5_n8), .Z(
        npu_inst_pe_1_4_5_N94) );
  MUX2_X1 npu_inst_pe_1_4_5_U156 ( .A(npu_inst_pe_1_4_5_n25), .B(
        npu_inst_pe_1_4_5_n24), .S(npu_inst_pe_1_4_5_n6), .Z(
        npu_inst_pe_1_4_5_n28) );
  MUX2_X1 npu_inst_pe_1_4_5_U155 ( .A(npu_inst_pe_1_4_5_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_4_5_int_q_reg_v_1__1_), .S(npu_inst_pe_1_4_5_n4), .Z(
        npu_inst_pe_1_4_5_n25) );
  MUX2_X1 npu_inst_pe_1_4_5_U154 ( .A(npu_inst_pe_1_4_5_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_4_5_int_q_reg_v_3__1_), .S(npu_inst_pe_1_4_5_n4), .Z(
        npu_inst_pe_1_4_5_n24) );
  MUX2_X1 npu_inst_pe_1_4_5_U153 ( .A(npu_inst_pe_1_4_5_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_4_5_int_q_reg_v_5__1_), .S(npu_inst_pe_1_4_5_n4), .Z(
        npu_inst_pe_1_4_5_n23) );
  MUX2_X1 npu_inst_pe_1_4_5_U152 ( .A(npu_inst_pe_1_4_5_n22), .B(
        npu_inst_pe_1_4_5_n19), .S(npu_inst_pe_1_4_5_n8), .Z(
        npu_inst_int_data_x_4__5__1_) );
  MUX2_X1 npu_inst_pe_1_4_5_U151 ( .A(npu_inst_pe_1_4_5_n21), .B(
        npu_inst_pe_1_4_5_n20), .S(npu_inst_pe_1_4_5_n6), .Z(
        npu_inst_pe_1_4_5_n22) );
  MUX2_X1 npu_inst_pe_1_4_5_U150 ( .A(npu_inst_pe_1_4_5_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_4_5_int_q_reg_h_1__1_), .S(npu_inst_pe_1_4_5_n4), .Z(
        npu_inst_pe_1_4_5_n21) );
  MUX2_X1 npu_inst_pe_1_4_5_U149 ( .A(npu_inst_pe_1_4_5_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_4_5_int_q_reg_h_3__1_), .S(npu_inst_pe_1_4_5_n4), .Z(
        npu_inst_pe_1_4_5_n20) );
  MUX2_X1 npu_inst_pe_1_4_5_U148 ( .A(npu_inst_pe_1_4_5_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_4_5_int_q_reg_h_5__1_), .S(npu_inst_pe_1_4_5_n4), .Z(
        npu_inst_pe_1_4_5_n19) );
  MUX2_X1 npu_inst_pe_1_4_5_U147 ( .A(npu_inst_pe_1_4_5_n18), .B(
        npu_inst_pe_1_4_5_n15), .S(npu_inst_pe_1_4_5_n8), .Z(
        npu_inst_int_data_x_4__5__0_) );
  MUX2_X1 npu_inst_pe_1_4_5_U146 ( .A(npu_inst_pe_1_4_5_n17), .B(
        npu_inst_pe_1_4_5_n16), .S(npu_inst_pe_1_4_5_n6), .Z(
        npu_inst_pe_1_4_5_n18) );
  MUX2_X1 npu_inst_pe_1_4_5_U145 ( .A(npu_inst_pe_1_4_5_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_4_5_int_q_reg_h_1__0_), .S(npu_inst_pe_1_4_5_n4), .Z(
        npu_inst_pe_1_4_5_n17) );
  MUX2_X1 npu_inst_pe_1_4_5_U144 ( .A(npu_inst_pe_1_4_5_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_4_5_int_q_reg_h_3__0_), .S(npu_inst_pe_1_4_5_n4), .Z(
        npu_inst_pe_1_4_5_n16) );
  MUX2_X1 npu_inst_pe_1_4_5_U143 ( .A(npu_inst_pe_1_4_5_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_4_5_int_q_reg_h_5__0_), .S(npu_inst_pe_1_4_5_n4), .Z(
        npu_inst_pe_1_4_5_n15) );
  XOR2_X1 npu_inst_pe_1_4_5_U142 ( .A(npu_inst_pe_1_4_5_int_data_0_), .B(
        npu_inst_pe_1_4_5_int_q_acc_0_), .Z(npu_inst_pe_1_4_5_N73) );
  AND2_X1 npu_inst_pe_1_4_5_U141 ( .A1(npu_inst_pe_1_4_5_int_q_acc_0_), .A2(
        npu_inst_pe_1_4_5_int_data_0_), .ZN(npu_inst_pe_1_4_5_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_4_5_U140 ( .A(npu_inst_pe_1_4_5_int_q_acc_0_), .B(
        npu_inst_pe_1_4_5_n13), .ZN(npu_inst_pe_1_4_5_N65) );
  OR2_X1 npu_inst_pe_1_4_5_U139 ( .A1(npu_inst_pe_1_4_5_n13), .A2(
        npu_inst_pe_1_4_5_int_q_acc_0_), .ZN(npu_inst_pe_1_4_5_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_4_5_U138 ( .A(npu_inst_pe_1_4_5_int_q_acc_2_), .B(
        npu_inst_pe_1_4_5_add_79_carry_2_), .Z(npu_inst_pe_1_4_5_N75) );
  AND2_X1 npu_inst_pe_1_4_5_U137 ( .A1(npu_inst_pe_1_4_5_add_79_carry_2_), 
        .A2(npu_inst_pe_1_4_5_int_q_acc_2_), .ZN(
        npu_inst_pe_1_4_5_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_4_5_U136 ( .A(npu_inst_pe_1_4_5_int_q_acc_3_), .B(
        npu_inst_pe_1_4_5_add_79_carry_3_), .Z(npu_inst_pe_1_4_5_N76) );
  AND2_X1 npu_inst_pe_1_4_5_U135 ( .A1(npu_inst_pe_1_4_5_add_79_carry_3_), 
        .A2(npu_inst_pe_1_4_5_int_q_acc_3_), .ZN(
        npu_inst_pe_1_4_5_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_4_5_U134 ( .A(npu_inst_pe_1_4_5_int_q_acc_4_), .B(
        npu_inst_pe_1_4_5_add_79_carry_4_), .Z(npu_inst_pe_1_4_5_N77) );
  AND2_X1 npu_inst_pe_1_4_5_U133 ( .A1(npu_inst_pe_1_4_5_add_79_carry_4_), 
        .A2(npu_inst_pe_1_4_5_int_q_acc_4_), .ZN(
        npu_inst_pe_1_4_5_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_4_5_U132 ( .A(npu_inst_pe_1_4_5_int_q_acc_5_), .B(
        npu_inst_pe_1_4_5_add_79_carry_5_), .Z(npu_inst_pe_1_4_5_N78) );
  AND2_X1 npu_inst_pe_1_4_5_U131 ( .A1(npu_inst_pe_1_4_5_add_79_carry_5_), 
        .A2(npu_inst_pe_1_4_5_int_q_acc_5_), .ZN(
        npu_inst_pe_1_4_5_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_4_5_U130 ( .A(npu_inst_pe_1_4_5_int_q_acc_6_), .B(
        npu_inst_pe_1_4_5_add_79_carry_6_), .Z(npu_inst_pe_1_4_5_N79) );
  AND2_X1 npu_inst_pe_1_4_5_U129 ( .A1(npu_inst_pe_1_4_5_add_79_carry_6_), 
        .A2(npu_inst_pe_1_4_5_int_q_acc_6_), .ZN(
        npu_inst_pe_1_4_5_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_4_5_U128 ( .A(npu_inst_pe_1_4_5_int_q_acc_7_), .B(
        npu_inst_pe_1_4_5_add_79_carry_7_), .Z(npu_inst_pe_1_4_5_N80) );
  XNOR2_X1 npu_inst_pe_1_4_5_U127 ( .A(npu_inst_pe_1_4_5_sub_77_carry_2_), .B(
        npu_inst_pe_1_4_5_int_q_acc_2_), .ZN(npu_inst_pe_1_4_5_N67) );
  OR2_X1 npu_inst_pe_1_4_5_U126 ( .A1(npu_inst_pe_1_4_5_int_q_acc_2_), .A2(
        npu_inst_pe_1_4_5_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_4_5_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_4_5_U125 ( .A(npu_inst_pe_1_4_5_sub_77_carry_3_), .B(
        npu_inst_pe_1_4_5_int_q_acc_3_), .ZN(npu_inst_pe_1_4_5_N68) );
  OR2_X1 npu_inst_pe_1_4_5_U124 ( .A1(npu_inst_pe_1_4_5_int_q_acc_3_), .A2(
        npu_inst_pe_1_4_5_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_4_5_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_4_5_U123 ( .A(npu_inst_pe_1_4_5_sub_77_carry_4_), .B(
        npu_inst_pe_1_4_5_int_q_acc_4_), .ZN(npu_inst_pe_1_4_5_N69) );
  OR2_X1 npu_inst_pe_1_4_5_U122 ( .A1(npu_inst_pe_1_4_5_int_q_acc_4_), .A2(
        npu_inst_pe_1_4_5_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_4_5_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_4_5_U121 ( .A(npu_inst_pe_1_4_5_sub_77_carry_5_), .B(
        npu_inst_pe_1_4_5_int_q_acc_5_), .ZN(npu_inst_pe_1_4_5_N70) );
  OR2_X1 npu_inst_pe_1_4_5_U120 ( .A1(npu_inst_pe_1_4_5_int_q_acc_5_), .A2(
        npu_inst_pe_1_4_5_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_4_5_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_4_5_U119 ( .A(npu_inst_pe_1_4_5_sub_77_carry_6_), .B(
        npu_inst_pe_1_4_5_int_q_acc_6_), .ZN(npu_inst_pe_1_4_5_N71) );
  OR2_X1 npu_inst_pe_1_4_5_U118 ( .A1(npu_inst_pe_1_4_5_int_q_acc_6_), .A2(
        npu_inst_pe_1_4_5_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_4_5_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_4_5_U117 ( .A(npu_inst_pe_1_4_5_int_q_acc_7_), .B(
        npu_inst_pe_1_4_5_sub_77_carry_7_), .ZN(npu_inst_pe_1_4_5_N72) );
  INV_X1 npu_inst_pe_1_4_5_U116 ( .A(npu_inst_n77), .ZN(npu_inst_pe_1_4_5_n7)
         );
  INV_X1 npu_inst_pe_1_4_5_U115 ( .A(npu_inst_pe_1_4_5_n7), .ZN(
        npu_inst_pe_1_4_5_n6) );
  INV_X1 npu_inst_pe_1_4_5_U114 ( .A(npu_inst_n55), .ZN(npu_inst_pe_1_4_5_n3)
         );
  AOI22_X1 npu_inst_pe_1_4_5_U113 ( .A1(npu_inst_int_data_y_5__5__0_), .A2(
        npu_inst_pe_1_4_5_n58), .B1(npu_inst_pe_1_4_5_n114), .B2(
        npu_inst_pe_1_4_5_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_4_5_n57) );
  INV_X1 npu_inst_pe_1_4_5_U112 ( .A(npu_inst_pe_1_4_5_n57), .ZN(
        npu_inst_pe_1_4_5_n108) );
  AOI22_X1 npu_inst_pe_1_4_5_U111 ( .A1(npu_inst_int_data_y_5__5__0_), .A2(
        npu_inst_pe_1_4_5_n54), .B1(npu_inst_pe_1_4_5_n115), .B2(
        npu_inst_pe_1_4_5_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_4_5_n53) );
  INV_X1 npu_inst_pe_1_4_5_U110 ( .A(npu_inst_pe_1_4_5_n53), .ZN(
        npu_inst_pe_1_4_5_n109) );
  AOI22_X1 npu_inst_pe_1_4_5_U107 ( .A1(npu_inst_int_data_y_5__5__0_), .A2(
        npu_inst_pe_1_4_5_n50), .B1(npu_inst_pe_1_4_5_n116), .B2(
        npu_inst_pe_1_4_5_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_4_5_n49) );
  INV_X1 npu_inst_pe_1_4_5_U106 ( .A(npu_inst_pe_1_4_5_n49), .ZN(
        npu_inst_pe_1_4_5_n110) );
  AOI22_X1 npu_inst_pe_1_4_5_U105 ( .A1(npu_inst_int_data_y_5__5__0_), .A2(
        npu_inst_pe_1_4_5_n46), .B1(npu_inst_pe_1_4_5_n117), .B2(
        npu_inst_pe_1_4_5_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_4_5_n45) );
  INV_X1 npu_inst_pe_1_4_5_U104 ( .A(npu_inst_pe_1_4_5_n45), .ZN(
        npu_inst_pe_1_4_5_n111) );
  AOI22_X1 npu_inst_pe_1_4_5_U103 ( .A1(npu_inst_int_data_y_5__5__0_), .A2(
        npu_inst_pe_1_4_5_n42), .B1(npu_inst_pe_1_4_5_n119), .B2(
        npu_inst_pe_1_4_5_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_4_5_n41) );
  INV_X1 npu_inst_pe_1_4_5_U102 ( .A(npu_inst_pe_1_4_5_n41), .ZN(
        npu_inst_pe_1_4_5_n112) );
  AOI22_X1 npu_inst_pe_1_4_5_U101 ( .A1(npu_inst_int_data_y_5__5__1_), .A2(
        npu_inst_pe_1_4_5_n58), .B1(npu_inst_pe_1_4_5_n114), .B2(
        npu_inst_pe_1_4_5_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_4_5_n59) );
  INV_X1 npu_inst_pe_1_4_5_U100 ( .A(npu_inst_pe_1_4_5_n59), .ZN(
        npu_inst_pe_1_4_5_n102) );
  AOI22_X1 npu_inst_pe_1_4_5_U99 ( .A1(npu_inst_int_data_y_5__5__1_), .A2(
        npu_inst_pe_1_4_5_n54), .B1(npu_inst_pe_1_4_5_n115), .B2(
        npu_inst_pe_1_4_5_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_4_5_n55) );
  INV_X1 npu_inst_pe_1_4_5_U98 ( .A(npu_inst_pe_1_4_5_n55), .ZN(
        npu_inst_pe_1_4_5_n103) );
  AOI22_X1 npu_inst_pe_1_4_5_U97 ( .A1(npu_inst_int_data_y_5__5__1_), .A2(
        npu_inst_pe_1_4_5_n50), .B1(npu_inst_pe_1_4_5_n116), .B2(
        npu_inst_pe_1_4_5_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_4_5_n51) );
  INV_X1 npu_inst_pe_1_4_5_U96 ( .A(npu_inst_pe_1_4_5_n51), .ZN(
        npu_inst_pe_1_4_5_n104) );
  AOI22_X1 npu_inst_pe_1_4_5_U95 ( .A1(npu_inst_int_data_y_5__5__1_), .A2(
        npu_inst_pe_1_4_5_n46), .B1(npu_inst_pe_1_4_5_n117), .B2(
        npu_inst_pe_1_4_5_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_4_5_n47) );
  INV_X1 npu_inst_pe_1_4_5_U94 ( .A(npu_inst_pe_1_4_5_n47), .ZN(
        npu_inst_pe_1_4_5_n105) );
  AOI22_X1 npu_inst_pe_1_4_5_U93 ( .A1(npu_inst_int_data_y_5__5__1_), .A2(
        npu_inst_pe_1_4_5_n42), .B1(npu_inst_pe_1_4_5_n119), .B2(
        npu_inst_pe_1_4_5_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_4_5_n43) );
  INV_X1 npu_inst_pe_1_4_5_U92 ( .A(npu_inst_pe_1_4_5_n43), .ZN(
        npu_inst_pe_1_4_5_n106) );
  AOI22_X1 npu_inst_pe_1_4_5_U91 ( .A1(npu_inst_pe_1_4_5_n38), .A2(
        npu_inst_int_data_y_5__5__1_), .B1(npu_inst_pe_1_4_5_n118), .B2(
        npu_inst_pe_1_4_5_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_4_5_n39) );
  INV_X1 npu_inst_pe_1_4_5_U90 ( .A(npu_inst_pe_1_4_5_n39), .ZN(
        npu_inst_pe_1_4_5_n107) );
  AOI22_X1 npu_inst_pe_1_4_5_U89 ( .A1(npu_inst_pe_1_4_5_n38), .A2(
        npu_inst_int_data_y_5__5__0_), .B1(npu_inst_pe_1_4_5_n118), .B2(
        npu_inst_pe_1_4_5_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_4_5_n37) );
  INV_X1 npu_inst_pe_1_4_5_U88 ( .A(npu_inst_pe_1_4_5_n37), .ZN(
        npu_inst_pe_1_4_5_n113) );
  NAND2_X1 npu_inst_pe_1_4_5_U87 ( .A1(npu_inst_pe_1_4_5_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_4_5_n60), .ZN(npu_inst_pe_1_4_5_n74) );
  OAI21_X1 npu_inst_pe_1_4_5_U86 ( .B1(npu_inst_pe_1_4_5_n63), .B2(
        npu_inst_pe_1_4_5_n60), .A(npu_inst_pe_1_4_5_n74), .ZN(
        npu_inst_pe_1_4_5_n97) );
  NAND2_X1 npu_inst_pe_1_4_5_U85 ( .A1(npu_inst_pe_1_4_5_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_4_5_n60), .ZN(npu_inst_pe_1_4_5_n73) );
  OAI21_X1 npu_inst_pe_1_4_5_U84 ( .B1(npu_inst_pe_1_4_5_n61), .B2(
        npu_inst_pe_1_4_5_n60), .A(npu_inst_pe_1_4_5_n73), .ZN(
        npu_inst_pe_1_4_5_n96) );
  NAND2_X1 npu_inst_pe_1_4_5_U83 ( .A1(npu_inst_pe_1_4_5_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_4_5_n56), .ZN(npu_inst_pe_1_4_5_n72) );
  OAI21_X1 npu_inst_pe_1_4_5_U82 ( .B1(npu_inst_pe_1_4_5_n63), .B2(
        npu_inst_pe_1_4_5_n56), .A(npu_inst_pe_1_4_5_n72), .ZN(
        npu_inst_pe_1_4_5_n95) );
  NAND2_X1 npu_inst_pe_1_4_5_U81 ( .A1(npu_inst_pe_1_4_5_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_4_5_n56), .ZN(npu_inst_pe_1_4_5_n71) );
  OAI21_X1 npu_inst_pe_1_4_5_U80 ( .B1(npu_inst_pe_1_4_5_n61), .B2(
        npu_inst_pe_1_4_5_n56), .A(npu_inst_pe_1_4_5_n71), .ZN(
        npu_inst_pe_1_4_5_n94) );
  NAND2_X1 npu_inst_pe_1_4_5_U79 ( .A1(npu_inst_pe_1_4_5_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_4_5_n52), .ZN(npu_inst_pe_1_4_5_n70) );
  OAI21_X1 npu_inst_pe_1_4_5_U78 ( .B1(npu_inst_pe_1_4_5_n63), .B2(
        npu_inst_pe_1_4_5_n52), .A(npu_inst_pe_1_4_5_n70), .ZN(
        npu_inst_pe_1_4_5_n93) );
  NAND2_X1 npu_inst_pe_1_4_5_U77 ( .A1(npu_inst_pe_1_4_5_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_4_5_n52), .ZN(npu_inst_pe_1_4_5_n69) );
  OAI21_X1 npu_inst_pe_1_4_5_U76 ( .B1(npu_inst_pe_1_4_5_n61), .B2(
        npu_inst_pe_1_4_5_n52), .A(npu_inst_pe_1_4_5_n69), .ZN(
        npu_inst_pe_1_4_5_n92) );
  NAND2_X1 npu_inst_pe_1_4_5_U75 ( .A1(npu_inst_pe_1_4_5_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_4_5_n48), .ZN(npu_inst_pe_1_4_5_n68) );
  OAI21_X1 npu_inst_pe_1_4_5_U74 ( .B1(npu_inst_pe_1_4_5_n63), .B2(
        npu_inst_pe_1_4_5_n48), .A(npu_inst_pe_1_4_5_n68), .ZN(
        npu_inst_pe_1_4_5_n91) );
  NAND2_X1 npu_inst_pe_1_4_5_U73 ( .A1(npu_inst_pe_1_4_5_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_4_5_n48), .ZN(npu_inst_pe_1_4_5_n67) );
  OAI21_X1 npu_inst_pe_1_4_5_U72 ( .B1(npu_inst_pe_1_4_5_n61), .B2(
        npu_inst_pe_1_4_5_n48), .A(npu_inst_pe_1_4_5_n67), .ZN(
        npu_inst_pe_1_4_5_n90) );
  NAND2_X1 npu_inst_pe_1_4_5_U71 ( .A1(npu_inst_pe_1_4_5_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_4_5_n44), .ZN(npu_inst_pe_1_4_5_n66) );
  OAI21_X1 npu_inst_pe_1_4_5_U70 ( .B1(npu_inst_pe_1_4_5_n63), .B2(
        npu_inst_pe_1_4_5_n44), .A(npu_inst_pe_1_4_5_n66), .ZN(
        npu_inst_pe_1_4_5_n89) );
  NAND2_X1 npu_inst_pe_1_4_5_U69 ( .A1(npu_inst_pe_1_4_5_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_4_5_n44), .ZN(npu_inst_pe_1_4_5_n65) );
  OAI21_X1 npu_inst_pe_1_4_5_U68 ( .B1(npu_inst_pe_1_4_5_n61), .B2(
        npu_inst_pe_1_4_5_n44), .A(npu_inst_pe_1_4_5_n65), .ZN(
        npu_inst_pe_1_4_5_n88) );
  NAND2_X1 npu_inst_pe_1_4_5_U67 ( .A1(npu_inst_pe_1_4_5_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_4_5_n40), .ZN(npu_inst_pe_1_4_5_n64) );
  OAI21_X1 npu_inst_pe_1_4_5_U66 ( .B1(npu_inst_pe_1_4_5_n63), .B2(
        npu_inst_pe_1_4_5_n40), .A(npu_inst_pe_1_4_5_n64), .ZN(
        npu_inst_pe_1_4_5_n87) );
  NAND2_X1 npu_inst_pe_1_4_5_U65 ( .A1(npu_inst_pe_1_4_5_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_4_5_n40), .ZN(npu_inst_pe_1_4_5_n62) );
  OAI21_X1 npu_inst_pe_1_4_5_U64 ( .B1(npu_inst_pe_1_4_5_n61), .B2(
        npu_inst_pe_1_4_5_n40), .A(npu_inst_pe_1_4_5_n62), .ZN(
        npu_inst_pe_1_4_5_n86) );
  AND2_X1 npu_inst_pe_1_4_5_U63 ( .A1(npu_inst_pe_1_4_5_N93), .A2(npu_inst_n55), .ZN(npu_inst_int_data_y_4__5__0_) );
  AND2_X1 npu_inst_pe_1_4_5_U62 ( .A1(npu_inst_n55), .A2(npu_inst_pe_1_4_5_N94), .ZN(npu_inst_int_data_y_4__5__1_) );
  NOR3_X1 npu_inst_pe_1_4_5_U61 ( .A1(npu_inst_pe_1_4_5_n26), .A2(npu_inst_n55), .A3(npu_inst_int_ckg[26]), .ZN(npu_inst_pe_1_4_5_n85) );
  OR2_X1 npu_inst_pe_1_4_5_U60 ( .A1(npu_inst_pe_1_4_5_n85), .A2(
        npu_inst_pe_1_4_5_n2), .ZN(npu_inst_pe_1_4_5_N84) );
  AND2_X1 npu_inst_pe_1_4_5_U59 ( .A1(npu_inst_pe_1_4_5_int_q_acc_0_), .A2(
        npu_inst_pe_1_4_5_n1), .ZN(npu_inst_int_data_res_4__5__0_) );
  AND2_X1 npu_inst_pe_1_4_5_U58 ( .A1(npu_inst_pe_1_4_5_n2), .A2(
        npu_inst_pe_1_4_5_int_q_acc_7_), .ZN(npu_inst_int_data_res_4__5__7_)
         );
  AND2_X1 npu_inst_pe_1_4_5_U57 ( .A1(npu_inst_pe_1_4_5_int_q_acc_1_), .A2(
        npu_inst_pe_1_4_5_n1), .ZN(npu_inst_int_data_res_4__5__1_) );
  AND2_X1 npu_inst_pe_1_4_5_U56 ( .A1(npu_inst_pe_1_4_5_int_q_acc_2_), .A2(
        npu_inst_pe_1_4_5_n1), .ZN(npu_inst_int_data_res_4__5__2_) );
  AND2_X1 npu_inst_pe_1_4_5_U55 ( .A1(npu_inst_pe_1_4_5_int_q_acc_3_), .A2(
        npu_inst_pe_1_4_5_n2), .ZN(npu_inst_int_data_res_4__5__3_) );
  AND2_X1 npu_inst_pe_1_4_5_U54 ( .A1(npu_inst_pe_1_4_5_int_q_acc_4_), .A2(
        npu_inst_pe_1_4_5_n2), .ZN(npu_inst_int_data_res_4__5__4_) );
  AND2_X1 npu_inst_pe_1_4_5_U53 ( .A1(npu_inst_pe_1_4_5_int_q_acc_5_), .A2(
        npu_inst_pe_1_4_5_n2), .ZN(npu_inst_int_data_res_4__5__5_) );
  AND2_X1 npu_inst_pe_1_4_5_U52 ( .A1(npu_inst_pe_1_4_5_int_q_acc_6_), .A2(
        npu_inst_pe_1_4_5_n2), .ZN(npu_inst_int_data_res_4__5__6_) );
  AOI222_X1 npu_inst_pe_1_4_5_U51 ( .A1(npu_inst_int_data_res_5__5__0_), .A2(
        npu_inst_pe_1_4_5_n1), .B1(npu_inst_pe_1_4_5_N73), .B2(
        npu_inst_pe_1_4_5_n76), .C1(npu_inst_pe_1_4_5_N65), .C2(
        npu_inst_pe_1_4_5_n77), .ZN(npu_inst_pe_1_4_5_n84) );
  INV_X1 npu_inst_pe_1_4_5_U50 ( .A(npu_inst_pe_1_4_5_n84), .ZN(
        npu_inst_pe_1_4_5_n101) );
  AOI222_X1 npu_inst_pe_1_4_5_U49 ( .A1(npu_inst_int_data_res_5__5__7_), .A2(
        npu_inst_pe_1_4_5_n1), .B1(npu_inst_pe_1_4_5_N80), .B2(
        npu_inst_pe_1_4_5_n76), .C1(npu_inst_pe_1_4_5_N72), .C2(
        npu_inst_pe_1_4_5_n77), .ZN(npu_inst_pe_1_4_5_n75) );
  INV_X1 npu_inst_pe_1_4_5_U48 ( .A(npu_inst_pe_1_4_5_n75), .ZN(
        npu_inst_pe_1_4_5_n33) );
  AOI222_X1 npu_inst_pe_1_4_5_U47 ( .A1(npu_inst_int_data_res_5__5__1_), .A2(
        npu_inst_pe_1_4_5_n1), .B1(npu_inst_pe_1_4_5_N74), .B2(
        npu_inst_pe_1_4_5_n76), .C1(npu_inst_pe_1_4_5_N66), .C2(
        npu_inst_pe_1_4_5_n77), .ZN(npu_inst_pe_1_4_5_n83) );
  INV_X1 npu_inst_pe_1_4_5_U46 ( .A(npu_inst_pe_1_4_5_n83), .ZN(
        npu_inst_pe_1_4_5_n100) );
  AOI222_X1 npu_inst_pe_1_4_5_U45 ( .A1(npu_inst_int_data_res_5__5__2_), .A2(
        npu_inst_pe_1_4_5_n1), .B1(npu_inst_pe_1_4_5_N75), .B2(
        npu_inst_pe_1_4_5_n76), .C1(npu_inst_pe_1_4_5_N67), .C2(
        npu_inst_pe_1_4_5_n77), .ZN(npu_inst_pe_1_4_5_n82) );
  INV_X1 npu_inst_pe_1_4_5_U44 ( .A(npu_inst_pe_1_4_5_n82), .ZN(
        npu_inst_pe_1_4_5_n99) );
  AOI222_X1 npu_inst_pe_1_4_5_U43 ( .A1(npu_inst_int_data_res_5__5__3_), .A2(
        npu_inst_pe_1_4_5_n1), .B1(npu_inst_pe_1_4_5_N76), .B2(
        npu_inst_pe_1_4_5_n76), .C1(npu_inst_pe_1_4_5_N68), .C2(
        npu_inst_pe_1_4_5_n77), .ZN(npu_inst_pe_1_4_5_n81) );
  INV_X1 npu_inst_pe_1_4_5_U42 ( .A(npu_inst_pe_1_4_5_n81), .ZN(
        npu_inst_pe_1_4_5_n98) );
  AOI222_X1 npu_inst_pe_1_4_5_U41 ( .A1(npu_inst_int_data_res_5__5__4_), .A2(
        npu_inst_pe_1_4_5_n1), .B1(npu_inst_pe_1_4_5_N77), .B2(
        npu_inst_pe_1_4_5_n76), .C1(npu_inst_pe_1_4_5_N69), .C2(
        npu_inst_pe_1_4_5_n77), .ZN(npu_inst_pe_1_4_5_n80) );
  INV_X1 npu_inst_pe_1_4_5_U40 ( .A(npu_inst_pe_1_4_5_n80), .ZN(
        npu_inst_pe_1_4_5_n36) );
  AOI222_X1 npu_inst_pe_1_4_5_U39 ( .A1(npu_inst_int_data_res_5__5__5_), .A2(
        npu_inst_pe_1_4_5_n1), .B1(npu_inst_pe_1_4_5_N78), .B2(
        npu_inst_pe_1_4_5_n76), .C1(npu_inst_pe_1_4_5_N70), .C2(
        npu_inst_pe_1_4_5_n77), .ZN(npu_inst_pe_1_4_5_n79) );
  INV_X1 npu_inst_pe_1_4_5_U38 ( .A(npu_inst_pe_1_4_5_n79), .ZN(
        npu_inst_pe_1_4_5_n35) );
  AOI222_X1 npu_inst_pe_1_4_5_U37 ( .A1(npu_inst_int_data_res_5__5__6_), .A2(
        npu_inst_pe_1_4_5_n1), .B1(npu_inst_pe_1_4_5_N79), .B2(
        npu_inst_pe_1_4_5_n76), .C1(npu_inst_pe_1_4_5_N71), .C2(
        npu_inst_pe_1_4_5_n77), .ZN(npu_inst_pe_1_4_5_n78) );
  INV_X1 npu_inst_pe_1_4_5_U36 ( .A(npu_inst_pe_1_4_5_n78), .ZN(
        npu_inst_pe_1_4_5_n34) );
  INV_X1 npu_inst_pe_1_4_5_U35 ( .A(npu_inst_pe_1_4_5_int_data_1_), .ZN(
        npu_inst_pe_1_4_5_n14) );
  AND2_X1 npu_inst_pe_1_4_5_U34 ( .A1(npu_inst_int_data_x_4__5__1_), .A2(
        npu_inst_pe_1_4_5_int_q_weight_1_), .ZN(npu_inst_pe_1_4_5_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_4_5_U33 ( .A1(npu_inst_int_data_x_4__5__0_), .A2(
        npu_inst_pe_1_4_5_int_q_weight_1_), .ZN(npu_inst_pe_1_4_5_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_4_5_U32 ( .A1(npu_inst_n55), .A2(
        npu_inst_int_data_y_5__5__1_), .B1(npu_inst_pe_1_4_5_n3), .B2(
        npu_inst_int_data_x_4__6__1_), .ZN(npu_inst_pe_1_4_5_n63) );
  AOI22_X1 npu_inst_pe_1_4_5_U31 ( .A1(npu_inst_n55), .A2(
        npu_inst_int_data_y_5__5__0_), .B1(npu_inst_pe_1_4_5_n3), .B2(
        npu_inst_int_data_x_4__6__0_), .ZN(npu_inst_pe_1_4_5_n61) );
  INV_X1 npu_inst_pe_1_4_5_U30 ( .A(npu_inst_pe_1_4_5_int_data_0_), .ZN(
        npu_inst_pe_1_4_5_n13) );
  INV_X1 npu_inst_pe_1_4_5_U29 ( .A(npu_inst_n69), .ZN(npu_inst_pe_1_4_5_n5)
         );
  OR3_X1 npu_inst_pe_1_4_5_U28 ( .A1(npu_inst_pe_1_4_5_n6), .A2(
        npu_inst_pe_1_4_5_n8), .A3(npu_inst_pe_1_4_5_n5), .ZN(
        npu_inst_pe_1_4_5_n56) );
  OR3_X1 npu_inst_pe_1_4_5_U27 ( .A1(npu_inst_pe_1_4_5_n5), .A2(
        npu_inst_pe_1_4_5_n8), .A3(npu_inst_pe_1_4_5_n7), .ZN(
        npu_inst_pe_1_4_5_n48) );
  INV_X1 npu_inst_pe_1_4_5_U26 ( .A(npu_inst_pe_1_4_5_n5), .ZN(
        npu_inst_pe_1_4_5_n4) );
  INV_X1 npu_inst_pe_1_4_5_U25 ( .A(npu_inst_n124), .ZN(npu_inst_pe_1_4_5_n12)
         );
  OR3_X1 npu_inst_pe_1_4_5_U24 ( .A1(npu_inst_pe_1_4_5_n4), .A2(
        npu_inst_pe_1_4_5_n8), .A3(npu_inst_pe_1_4_5_n7), .ZN(
        npu_inst_pe_1_4_5_n52) );
  OR3_X1 npu_inst_pe_1_4_5_U23 ( .A1(npu_inst_pe_1_4_5_n6), .A2(
        npu_inst_pe_1_4_5_n8), .A3(npu_inst_pe_1_4_5_n4), .ZN(
        npu_inst_pe_1_4_5_n60) );
  NOR2_X1 npu_inst_pe_1_4_5_U22 ( .A1(npu_inst_pe_1_4_5_n60), .A2(
        npu_inst_pe_1_4_5_n3), .ZN(npu_inst_pe_1_4_5_n58) );
  NOR2_X1 npu_inst_pe_1_4_5_U21 ( .A1(npu_inst_pe_1_4_5_n56), .A2(
        npu_inst_pe_1_4_5_n3), .ZN(npu_inst_pe_1_4_5_n54) );
  NOR2_X1 npu_inst_pe_1_4_5_U20 ( .A1(npu_inst_pe_1_4_5_n52), .A2(
        npu_inst_pe_1_4_5_n3), .ZN(npu_inst_pe_1_4_5_n50) );
  NOR2_X1 npu_inst_pe_1_4_5_U19 ( .A1(npu_inst_pe_1_4_5_n48), .A2(
        npu_inst_pe_1_4_5_n3), .ZN(npu_inst_pe_1_4_5_n46) );
  NOR2_X1 npu_inst_pe_1_4_5_U18 ( .A1(npu_inst_pe_1_4_5_n40), .A2(
        npu_inst_pe_1_4_5_n3), .ZN(npu_inst_pe_1_4_5_n38) );
  NOR2_X1 npu_inst_pe_1_4_5_U17 ( .A1(npu_inst_pe_1_4_5_n44), .A2(
        npu_inst_pe_1_4_5_n3), .ZN(npu_inst_pe_1_4_5_n42) );
  BUF_X1 npu_inst_pe_1_4_5_U16 ( .A(npu_inst_n98), .Z(npu_inst_pe_1_4_5_n8) );
  BUF_X1 npu_inst_pe_1_4_5_U15 ( .A(npu_inst_pe_1_4_5_n12), .Z(
        npu_inst_pe_1_4_5_n11) );
  BUF_X1 npu_inst_pe_1_4_5_U14 ( .A(npu_inst_pe_1_4_5_n12), .Z(
        npu_inst_pe_1_4_5_n10) );
  BUF_X1 npu_inst_pe_1_4_5_U13 ( .A(npu_inst_pe_1_4_5_n12), .Z(
        npu_inst_pe_1_4_5_n9) );
  INV_X1 npu_inst_pe_1_4_5_U12 ( .A(npu_inst_pe_1_4_5_n38), .ZN(
        npu_inst_pe_1_4_5_n118) );
  INV_X1 npu_inst_pe_1_4_5_U11 ( .A(npu_inst_pe_1_4_5_n58), .ZN(
        npu_inst_pe_1_4_5_n114) );
  INV_X1 npu_inst_pe_1_4_5_U10 ( .A(npu_inst_pe_1_4_5_n54), .ZN(
        npu_inst_pe_1_4_5_n115) );
  INV_X1 npu_inst_pe_1_4_5_U9 ( .A(npu_inst_pe_1_4_5_n50), .ZN(
        npu_inst_pe_1_4_5_n116) );
  INV_X1 npu_inst_pe_1_4_5_U8 ( .A(npu_inst_pe_1_4_5_n46), .ZN(
        npu_inst_pe_1_4_5_n117) );
  INV_X1 npu_inst_pe_1_4_5_U7 ( .A(npu_inst_pe_1_4_5_n42), .ZN(
        npu_inst_pe_1_4_5_n119) );
  BUF_X1 npu_inst_pe_1_4_5_U6 ( .A(npu_inst_n20), .Z(npu_inst_pe_1_4_5_n2) );
  BUF_X1 npu_inst_pe_1_4_5_U5 ( .A(npu_inst_n20), .Z(npu_inst_pe_1_4_5_n1) );
  NOR2_X1 npu_inst_pe_1_4_5_U4 ( .A1(npu_inst_pe_1_4_5_int_q_weight_0_), .A2(
        npu_inst_pe_1_4_5_n1), .ZN(npu_inst_pe_1_4_5_n76) );
  NOR2_X1 npu_inst_pe_1_4_5_U3 ( .A1(npu_inst_pe_1_4_5_n27), .A2(
        npu_inst_pe_1_4_5_n1), .ZN(npu_inst_pe_1_4_5_n77) );
  FA_X1 npu_inst_pe_1_4_5_sub_77_U2_1 ( .A(npu_inst_pe_1_4_5_int_q_acc_1_), 
        .B(npu_inst_pe_1_4_5_n14), .CI(npu_inst_pe_1_4_5_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_4_5_sub_77_carry_2_), .S(npu_inst_pe_1_4_5_N66) );
  FA_X1 npu_inst_pe_1_4_5_add_79_U1_1 ( .A(npu_inst_pe_1_4_5_int_q_acc_1_), 
        .B(npu_inst_pe_1_4_5_int_data_1_), .CI(
        npu_inst_pe_1_4_5_add_79_carry_1_), .CO(
        npu_inst_pe_1_4_5_add_79_carry_2_), .S(npu_inst_pe_1_4_5_N74) );
  NAND3_X1 npu_inst_pe_1_4_5_U109 ( .A1(npu_inst_pe_1_4_5_n5), .A2(
        npu_inst_pe_1_4_5_n7), .A3(npu_inst_pe_1_4_5_n8), .ZN(
        npu_inst_pe_1_4_5_n44) );
  NAND3_X1 npu_inst_pe_1_4_5_U108 ( .A1(npu_inst_pe_1_4_5_n4), .A2(
        npu_inst_pe_1_4_5_n7), .A3(npu_inst_pe_1_4_5_n8), .ZN(
        npu_inst_pe_1_4_5_n40) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_4_5_n34), .CK(
        npu_inst_pe_1_4_5_net3442), .RN(npu_inst_pe_1_4_5_n9), .Q(
        npu_inst_pe_1_4_5_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_4_5_n35), .CK(
        npu_inst_pe_1_4_5_net3442), .RN(npu_inst_pe_1_4_5_n9), .Q(
        npu_inst_pe_1_4_5_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_4_5_n36), .CK(
        npu_inst_pe_1_4_5_net3442), .RN(npu_inst_pe_1_4_5_n9), .Q(
        npu_inst_pe_1_4_5_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_4_5_n98), .CK(
        npu_inst_pe_1_4_5_net3442), .RN(npu_inst_pe_1_4_5_n9), .Q(
        npu_inst_pe_1_4_5_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_4_5_n99), .CK(
        npu_inst_pe_1_4_5_net3442), .RN(npu_inst_pe_1_4_5_n9), .Q(
        npu_inst_pe_1_4_5_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_4_5_n100), 
        .CK(npu_inst_pe_1_4_5_net3442), .RN(npu_inst_pe_1_4_5_n9), .Q(
        npu_inst_pe_1_4_5_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_4_5_n33), .CK(
        npu_inst_pe_1_4_5_net3442), .RN(npu_inst_pe_1_4_5_n9), .Q(
        npu_inst_pe_1_4_5_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_4_5_n101), 
        .CK(npu_inst_pe_1_4_5_net3442), .RN(npu_inst_pe_1_4_5_n9), .Q(
        npu_inst_pe_1_4_5_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_weight_reg_0_ ( .D(npu_inst_n110), .CK(
        npu_inst_pe_1_4_5_net3448), .RN(npu_inst_pe_1_4_5_n9), .Q(
        npu_inst_pe_1_4_5_int_q_weight_0_), .QN(npu_inst_pe_1_4_5_n27) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_weight_reg_1_ ( .D(npu_inst_n116), .CK(
        npu_inst_pe_1_4_5_net3448), .RN(npu_inst_pe_1_4_5_n9), .Q(
        npu_inst_pe_1_4_5_int_q_weight_1_), .QN(npu_inst_pe_1_4_5_n26) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_4_5_n113), 
        .CK(npu_inst_pe_1_4_5_net3448), .RN(npu_inst_pe_1_4_5_n9), .Q(
        npu_inst_pe_1_4_5_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_4_5_n107), 
        .CK(npu_inst_pe_1_4_5_net3448), .RN(npu_inst_pe_1_4_5_n9), .Q(
        npu_inst_pe_1_4_5_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_4_5_n112), 
        .CK(npu_inst_pe_1_4_5_net3448), .RN(npu_inst_pe_1_4_5_n10), .Q(
        npu_inst_pe_1_4_5_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_4_5_n106), 
        .CK(npu_inst_pe_1_4_5_net3448), .RN(npu_inst_pe_1_4_5_n10), .Q(
        npu_inst_pe_1_4_5_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_4_5_n111), 
        .CK(npu_inst_pe_1_4_5_net3448), .RN(npu_inst_pe_1_4_5_n10), .Q(
        npu_inst_pe_1_4_5_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_4_5_n105), 
        .CK(npu_inst_pe_1_4_5_net3448), .RN(npu_inst_pe_1_4_5_n10), .Q(
        npu_inst_pe_1_4_5_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_4_5_n110), 
        .CK(npu_inst_pe_1_4_5_net3448), .RN(npu_inst_pe_1_4_5_n10), .Q(
        npu_inst_pe_1_4_5_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_4_5_n104), 
        .CK(npu_inst_pe_1_4_5_net3448), .RN(npu_inst_pe_1_4_5_n10), .Q(
        npu_inst_pe_1_4_5_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_4_5_n109), 
        .CK(npu_inst_pe_1_4_5_net3448), .RN(npu_inst_pe_1_4_5_n10), .Q(
        npu_inst_pe_1_4_5_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_4_5_n103), 
        .CK(npu_inst_pe_1_4_5_net3448), .RN(npu_inst_pe_1_4_5_n10), .Q(
        npu_inst_pe_1_4_5_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_4_5_n108), 
        .CK(npu_inst_pe_1_4_5_net3448), .RN(npu_inst_pe_1_4_5_n10), .Q(
        npu_inst_pe_1_4_5_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_4_5_n102), 
        .CK(npu_inst_pe_1_4_5_net3448), .RN(npu_inst_pe_1_4_5_n10), .Q(
        npu_inst_pe_1_4_5_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_4_5_n86), 
        .CK(npu_inst_pe_1_4_5_net3448), .RN(npu_inst_pe_1_4_5_n10), .Q(
        npu_inst_pe_1_4_5_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_4_5_n87), 
        .CK(npu_inst_pe_1_4_5_net3448), .RN(npu_inst_pe_1_4_5_n10), .Q(
        npu_inst_pe_1_4_5_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_4_5_n88), 
        .CK(npu_inst_pe_1_4_5_net3448), .RN(npu_inst_pe_1_4_5_n11), .Q(
        npu_inst_pe_1_4_5_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_4_5_n89), 
        .CK(npu_inst_pe_1_4_5_net3448), .RN(npu_inst_pe_1_4_5_n11), .Q(
        npu_inst_pe_1_4_5_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_4_5_n90), 
        .CK(npu_inst_pe_1_4_5_net3448), .RN(npu_inst_pe_1_4_5_n11), .Q(
        npu_inst_pe_1_4_5_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_4_5_n91), 
        .CK(npu_inst_pe_1_4_5_net3448), .RN(npu_inst_pe_1_4_5_n11), .Q(
        npu_inst_pe_1_4_5_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_4_5_n92), 
        .CK(npu_inst_pe_1_4_5_net3448), .RN(npu_inst_pe_1_4_5_n11), .Q(
        npu_inst_pe_1_4_5_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_4_5_n93), 
        .CK(npu_inst_pe_1_4_5_net3448), .RN(npu_inst_pe_1_4_5_n11), .Q(
        npu_inst_pe_1_4_5_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_4_5_n94), 
        .CK(npu_inst_pe_1_4_5_net3448), .RN(npu_inst_pe_1_4_5_n11), .Q(
        npu_inst_pe_1_4_5_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_4_5_n95), 
        .CK(npu_inst_pe_1_4_5_net3448), .RN(npu_inst_pe_1_4_5_n11), .Q(
        npu_inst_pe_1_4_5_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_4_5_n96), 
        .CK(npu_inst_pe_1_4_5_net3448), .RN(npu_inst_pe_1_4_5_n11), .Q(
        npu_inst_pe_1_4_5_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_4_5_n97), 
        .CK(npu_inst_pe_1_4_5_net3448), .RN(npu_inst_pe_1_4_5_n11), .Q(
        npu_inst_pe_1_4_5_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_4_5_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_4_5_N84), .SE(1'b0), .GCK(npu_inst_pe_1_4_5_net3442) );
  CLKGATETST_X1 npu_inst_pe_1_4_5_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n63), .SE(1'b0), .GCK(npu_inst_pe_1_4_5_net3448) );
  MUX2_X1 npu_inst_pe_1_4_6_U162 ( .A(npu_inst_pe_1_4_6_n32), .B(
        npu_inst_pe_1_4_6_n29), .S(npu_inst_pe_1_4_6_n8), .Z(
        npu_inst_pe_1_4_6_N93) );
  MUX2_X1 npu_inst_pe_1_4_6_U161 ( .A(npu_inst_pe_1_4_6_n31), .B(
        npu_inst_pe_1_4_6_n30), .S(npu_inst_pe_1_4_6_n6), .Z(
        npu_inst_pe_1_4_6_n32) );
  MUX2_X1 npu_inst_pe_1_4_6_U160 ( .A(npu_inst_pe_1_4_6_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_4_6_int_q_reg_v_1__0_), .S(npu_inst_pe_1_4_6_n4), .Z(
        npu_inst_pe_1_4_6_n31) );
  MUX2_X1 npu_inst_pe_1_4_6_U159 ( .A(npu_inst_pe_1_4_6_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_4_6_int_q_reg_v_3__0_), .S(npu_inst_pe_1_4_6_n4), .Z(
        npu_inst_pe_1_4_6_n30) );
  MUX2_X1 npu_inst_pe_1_4_6_U158 ( .A(npu_inst_pe_1_4_6_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_4_6_int_q_reg_v_5__0_), .S(npu_inst_pe_1_4_6_n4), .Z(
        npu_inst_pe_1_4_6_n29) );
  MUX2_X1 npu_inst_pe_1_4_6_U157 ( .A(npu_inst_pe_1_4_6_n28), .B(
        npu_inst_pe_1_4_6_n23), .S(npu_inst_pe_1_4_6_n8), .Z(
        npu_inst_pe_1_4_6_N94) );
  MUX2_X1 npu_inst_pe_1_4_6_U156 ( .A(npu_inst_pe_1_4_6_n25), .B(
        npu_inst_pe_1_4_6_n24), .S(npu_inst_pe_1_4_6_n6), .Z(
        npu_inst_pe_1_4_6_n28) );
  MUX2_X1 npu_inst_pe_1_4_6_U155 ( .A(npu_inst_pe_1_4_6_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_4_6_int_q_reg_v_1__1_), .S(npu_inst_pe_1_4_6_n4), .Z(
        npu_inst_pe_1_4_6_n25) );
  MUX2_X1 npu_inst_pe_1_4_6_U154 ( .A(npu_inst_pe_1_4_6_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_4_6_int_q_reg_v_3__1_), .S(npu_inst_pe_1_4_6_n4), .Z(
        npu_inst_pe_1_4_6_n24) );
  MUX2_X1 npu_inst_pe_1_4_6_U153 ( .A(npu_inst_pe_1_4_6_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_4_6_int_q_reg_v_5__1_), .S(npu_inst_pe_1_4_6_n4), .Z(
        npu_inst_pe_1_4_6_n23) );
  MUX2_X1 npu_inst_pe_1_4_6_U152 ( .A(npu_inst_pe_1_4_6_n22), .B(
        npu_inst_pe_1_4_6_n19), .S(npu_inst_pe_1_4_6_n8), .Z(
        npu_inst_int_data_x_4__6__1_) );
  MUX2_X1 npu_inst_pe_1_4_6_U151 ( .A(npu_inst_pe_1_4_6_n21), .B(
        npu_inst_pe_1_4_6_n20), .S(npu_inst_pe_1_4_6_n6), .Z(
        npu_inst_pe_1_4_6_n22) );
  MUX2_X1 npu_inst_pe_1_4_6_U150 ( .A(npu_inst_pe_1_4_6_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_4_6_int_q_reg_h_1__1_), .S(npu_inst_pe_1_4_6_n4), .Z(
        npu_inst_pe_1_4_6_n21) );
  MUX2_X1 npu_inst_pe_1_4_6_U149 ( .A(npu_inst_pe_1_4_6_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_4_6_int_q_reg_h_3__1_), .S(npu_inst_pe_1_4_6_n4), .Z(
        npu_inst_pe_1_4_6_n20) );
  MUX2_X1 npu_inst_pe_1_4_6_U148 ( .A(npu_inst_pe_1_4_6_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_4_6_int_q_reg_h_5__1_), .S(npu_inst_pe_1_4_6_n4), .Z(
        npu_inst_pe_1_4_6_n19) );
  MUX2_X1 npu_inst_pe_1_4_6_U147 ( .A(npu_inst_pe_1_4_6_n18), .B(
        npu_inst_pe_1_4_6_n15), .S(npu_inst_pe_1_4_6_n8), .Z(
        npu_inst_int_data_x_4__6__0_) );
  MUX2_X1 npu_inst_pe_1_4_6_U146 ( .A(npu_inst_pe_1_4_6_n17), .B(
        npu_inst_pe_1_4_6_n16), .S(npu_inst_pe_1_4_6_n6), .Z(
        npu_inst_pe_1_4_6_n18) );
  MUX2_X1 npu_inst_pe_1_4_6_U145 ( .A(npu_inst_pe_1_4_6_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_4_6_int_q_reg_h_1__0_), .S(npu_inst_pe_1_4_6_n4), .Z(
        npu_inst_pe_1_4_6_n17) );
  MUX2_X1 npu_inst_pe_1_4_6_U144 ( .A(npu_inst_pe_1_4_6_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_4_6_int_q_reg_h_3__0_), .S(npu_inst_pe_1_4_6_n4), .Z(
        npu_inst_pe_1_4_6_n16) );
  MUX2_X1 npu_inst_pe_1_4_6_U143 ( .A(npu_inst_pe_1_4_6_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_4_6_int_q_reg_h_5__0_), .S(npu_inst_pe_1_4_6_n4), .Z(
        npu_inst_pe_1_4_6_n15) );
  XOR2_X1 npu_inst_pe_1_4_6_U142 ( .A(npu_inst_pe_1_4_6_int_data_0_), .B(
        npu_inst_pe_1_4_6_int_q_acc_0_), .Z(npu_inst_pe_1_4_6_N73) );
  AND2_X1 npu_inst_pe_1_4_6_U141 ( .A1(npu_inst_pe_1_4_6_int_q_acc_0_), .A2(
        npu_inst_pe_1_4_6_int_data_0_), .ZN(npu_inst_pe_1_4_6_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_4_6_U140 ( .A(npu_inst_pe_1_4_6_int_q_acc_0_), .B(
        npu_inst_pe_1_4_6_n13), .ZN(npu_inst_pe_1_4_6_N65) );
  OR2_X1 npu_inst_pe_1_4_6_U139 ( .A1(npu_inst_pe_1_4_6_n13), .A2(
        npu_inst_pe_1_4_6_int_q_acc_0_), .ZN(npu_inst_pe_1_4_6_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_4_6_U138 ( .A(npu_inst_pe_1_4_6_int_q_acc_2_), .B(
        npu_inst_pe_1_4_6_add_79_carry_2_), .Z(npu_inst_pe_1_4_6_N75) );
  AND2_X1 npu_inst_pe_1_4_6_U137 ( .A1(npu_inst_pe_1_4_6_add_79_carry_2_), 
        .A2(npu_inst_pe_1_4_6_int_q_acc_2_), .ZN(
        npu_inst_pe_1_4_6_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_4_6_U136 ( .A(npu_inst_pe_1_4_6_int_q_acc_3_), .B(
        npu_inst_pe_1_4_6_add_79_carry_3_), .Z(npu_inst_pe_1_4_6_N76) );
  AND2_X1 npu_inst_pe_1_4_6_U135 ( .A1(npu_inst_pe_1_4_6_add_79_carry_3_), 
        .A2(npu_inst_pe_1_4_6_int_q_acc_3_), .ZN(
        npu_inst_pe_1_4_6_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_4_6_U134 ( .A(npu_inst_pe_1_4_6_int_q_acc_4_), .B(
        npu_inst_pe_1_4_6_add_79_carry_4_), .Z(npu_inst_pe_1_4_6_N77) );
  AND2_X1 npu_inst_pe_1_4_6_U133 ( .A1(npu_inst_pe_1_4_6_add_79_carry_4_), 
        .A2(npu_inst_pe_1_4_6_int_q_acc_4_), .ZN(
        npu_inst_pe_1_4_6_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_4_6_U132 ( .A(npu_inst_pe_1_4_6_int_q_acc_5_), .B(
        npu_inst_pe_1_4_6_add_79_carry_5_), .Z(npu_inst_pe_1_4_6_N78) );
  AND2_X1 npu_inst_pe_1_4_6_U131 ( .A1(npu_inst_pe_1_4_6_add_79_carry_5_), 
        .A2(npu_inst_pe_1_4_6_int_q_acc_5_), .ZN(
        npu_inst_pe_1_4_6_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_4_6_U130 ( .A(npu_inst_pe_1_4_6_int_q_acc_6_), .B(
        npu_inst_pe_1_4_6_add_79_carry_6_), .Z(npu_inst_pe_1_4_6_N79) );
  AND2_X1 npu_inst_pe_1_4_6_U129 ( .A1(npu_inst_pe_1_4_6_add_79_carry_6_), 
        .A2(npu_inst_pe_1_4_6_int_q_acc_6_), .ZN(
        npu_inst_pe_1_4_6_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_4_6_U128 ( .A(npu_inst_pe_1_4_6_int_q_acc_7_), .B(
        npu_inst_pe_1_4_6_add_79_carry_7_), .Z(npu_inst_pe_1_4_6_N80) );
  XNOR2_X1 npu_inst_pe_1_4_6_U127 ( .A(npu_inst_pe_1_4_6_sub_77_carry_2_), .B(
        npu_inst_pe_1_4_6_int_q_acc_2_), .ZN(npu_inst_pe_1_4_6_N67) );
  OR2_X1 npu_inst_pe_1_4_6_U126 ( .A1(npu_inst_pe_1_4_6_int_q_acc_2_), .A2(
        npu_inst_pe_1_4_6_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_4_6_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_4_6_U125 ( .A(npu_inst_pe_1_4_6_sub_77_carry_3_), .B(
        npu_inst_pe_1_4_6_int_q_acc_3_), .ZN(npu_inst_pe_1_4_6_N68) );
  OR2_X1 npu_inst_pe_1_4_6_U124 ( .A1(npu_inst_pe_1_4_6_int_q_acc_3_), .A2(
        npu_inst_pe_1_4_6_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_4_6_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_4_6_U123 ( .A(npu_inst_pe_1_4_6_sub_77_carry_4_), .B(
        npu_inst_pe_1_4_6_int_q_acc_4_), .ZN(npu_inst_pe_1_4_6_N69) );
  OR2_X1 npu_inst_pe_1_4_6_U122 ( .A1(npu_inst_pe_1_4_6_int_q_acc_4_), .A2(
        npu_inst_pe_1_4_6_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_4_6_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_4_6_U121 ( .A(npu_inst_pe_1_4_6_sub_77_carry_5_), .B(
        npu_inst_pe_1_4_6_int_q_acc_5_), .ZN(npu_inst_pe_1_4_6_N70) );
  OR2_X1 npu_inst_pe_1_4_6_U120 ( .A1(npu_inst_pe_1_4_6_int_q_acc_5_), .A2(
        npu_inst_pe_1_4_6_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_4_6_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_4_6_U119 ( .A(npu_inst_pe_1_4_6_sub_77_carry_6_), .B(
        npu_inst_pe_1_4_6_int_q_acc_6_), .ZN(npu_inst_pe_1_4_6_N71) );
  OR2_X1 npu_inst_pe_1_4_6_U118 ( .A1(npu_inst_pe_1_4_6_int_q_acc_6_), .A2(
        npu_inst_pe_1_4_6_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_4_6_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_4_6_U117 ( .A(npu_inst_pe_1_4_6_int_q_acc_7_), .B(
        npu_inst_pe_1_4_6_sub_77_carry_7_), .ZN(npu_inst_pe_1_4_6_N72) );
  INV_X1 npu_inst_pe_1_4_6_U116 ( .A(npu_inst_n77), .ZN(npu_inst_pe_1_4_6_n7)
         );
  INV_X1 npu_inst_pe_1_4_6_U115 ( .A(npu_inst_pe_1_4_6_n7), .ZN(
        npu_inst_pe_1_4_6_n6) );
  INV_X1 npu_inst_pe_1_4_6_U114 ( .A(npu_inst_n55), .ZN(npu_inst_pe_1_4_6_n3)
         );
  AOI22_X1 npu_inst_pe_1_4_6_U113 ( .A1(npu_inst_int_data_y_5__6__0_), .A2(
        npu_inst_pe_1_4_6_n58), .B1(npu_inst_pe_1_4_6_n114), .B2(
        npu_inst_pe_1_4_6_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_4_6_n57) );
  INV_X1 npu_inst_pe_1_4_6_U112 ( .A(npu_inst_pe_1_4_6_n57), .ZN(
        npu_inst_pe_1_4_6_n108) );
  AOI22_X1 npu_inst_pe_1_4_6_U111 ( .A1(npu_inst_int_data_y_5__6__0_), .A2(
        npu_inst_pe_1_4_6_n54), .B1(npu_inst_pe_1_4_6_n115), .B2(
        npu_inst_pe_1_4_6_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_4_6_n53) );
  INV_X1 npu_inst_pe_1_4_6_U110 ( .A(npu_inst_pe_1_4_6_n53), .ZN(
        npu_inst_pe_1_4_6_n109) );
  AOI22_X1 npu_inst_pe_1_4_6_U107 ( .A1(npu_inst_int_data_y_5__6__0_), .A2(
        npu_inst_pe_1_4_6_n50), .B1(npu_inst_pe_1_4_6_n116), .B2(
        npu_inst_pe_1_4_6_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_4_6_n49) );
  INV_X1 npu_inst_pe_1_4_6_U106 ( .A(npu_inst_pe_1_4_6_n49), .ZN(
        npu_inst_pe_1_4_6_n110) );
  AOI22_X1 npu_inst_pe_1_4_6_U105 ( .A1(npu_inst_int_data_y_5__6__0_), .A2(
        npu_inst_pe_1_4_6_n46), .B1(npu_inst_pe_1_4_6_n117), .B2(
        npu_inst_pe_1_4_6_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_4_6_n45) );
  INV_X1 npu_inst_pe_1_4_6_U104 ( .A(npu_inst_pe_1_4_6_n45), .ZN(
        npu_inst_pe_1_4_6_n111) );
  AOI22_X1 npu_inst_pe_1_4_6_U103 ( .A1(npu_inst_int_data_y_5__6__0_), .A2(
        npu_inst_pe_1_4_6_n42), .B1(npu_inst_pe_1_4_6_n119), .B2(
        npu_inst_pe_1_4_6_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_4_6_n41) );
  INV_X1 npu_inst_pe_1_4_6_U102 ( .A(npu_inst_pe_1_4_6_n41), .ZN(
        npu_inst_pe_1_4_6_n112) );
  AOI22_X1 npu_inst_pe_1_4_6_U101 ( .A1(npu_inst_int_data_y_5__6__1_), .A2(
        npu_inst_pe_1_4_6_n58), .B1(npu_inst_pe_1_4_6_n114), .B2(
        npu_inst_pe_1_4_6_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_4_6_n59) );
  INV_X1 npu_inst_pe_1_4_6_U100 ( .A(npu_inst_pe_1_4_6_n59), .ZN(
        npu_inst_pe_1_4_6_n102) );
  AOI22_X1 npu_inst_pe_1_4_6_U99 ( .A1(npu_inst_int_data_y_5__6__1_), .A2(
        npu_inst_pe_1_4_6_n54), .B1(npu_inst_pe_1_4_6_n115), .B2(
        npu_inst_pe_1_4_6_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_4_6_n55) );
  INV_X1 npu_inst_pe_1_4_6_U98 ( .A(npu_inst_pe_1_4_6_n55), .ZN(
        npu_inst_pe_1_4_6_n103) );
  AOI22_X1 npu_inst_pe_1_4_6_U97 ( .A1(npu_inst_int_data_y_5__6__1_), .A2(
        npu_inst_pe_1_4_6_n50), .B1(npu_inst_pe_1_4_6_n116), .B2(
        npu_inst_pe_1_4_6_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_4_6_n51) );
  INV_X1 npu_inst_pe_1_4_6_U96 ( .A(npu_inst_pe_1_4_6_n51), .ZN(
        npu_inst_pe_1_4_6_n104) );
  AOI22_X1 npu_inst_pe_1_4_6_U95 ( .A1(npu_inst_int_data_y_5__6__1_), .A2(
        npu_inst_pe_1_4_6_n46), .B1(npu_inst_pe_1_4_6_n117), .B2(
        npu_inst_pe_1_4_6_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_4_6_n47) );
  INV_X1 npu_inst_pe_1_4_6_U94 ( .A(npu_inst_pe_1_4_6_n47), .ZN(
        npu_inst_pe_1_4_6_n105) );
  AOI22_X1 npu_inst_pe_1_4_6_U93 ( .A1(npu_inst_int_data_y_5__6__1_), .A2(
        npu_inst_pe_1_4_6_n42), .B1(npu_inst_pe_1_4_6_n119), .B2(
        npu_inst_pe_1_4_6_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_4_6_n43) );
  INV_X1 npu_inst_pe_1_4_6_U92 ( .A(npu_inst_pe_1_4_6_n43), .ZN(
        npu_inst_pe_1_4_6_n106) );
  AOI22_X1 npu_inst_pe_1_4_6_U91 ( .A1(npu_inst_pe_1_4_6_n38), .A2(
        npu_inst_int_data_y_5__6__1_), .B1(npu_inst_pe_1_4_6_n118), .B2(
        npu_inst_pe_1_4_6_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_4_6_n39) );
  INV_X1 npu_inst_pe_1_4_6_U90 ( .A(npu_inst_pe_1_4_6_n39), .ZN(
        npu_inst_pe_1_4_6_n107) );
  AOI22_X1 npu_inst_pe_1_4_6_U89 ( .A1(npu_inst_pe_1_4_6_n38), .A2(
        npu_inst_int_data_y_5__6__0_), .B1(npu_inst_pe_1_4_6_n118), .B2(
        npu_inst_pe_1_4_6_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_4_6_n37) );
  INV_X1 npu_inst_pe_1_4_6_U88 ( .A(npu_inst_pe_1_4_6_n37), .ZN(
        npu_inst_pe_1_4_6_n113) );
  NAND2_X1 npu_inst_pe_1_4_6_U87 ( .A1(npu_inst_pe_1_4_6_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_4_6_n60), .ZN(npu_inst_pe_1_4_6_n74) );
  OAI21_X1 npu_inst_pe_1_4_6_U86 ( .B1(npu_inst_pe_1_4_6_n63), .B2(
        npu_inst_pe_1_4_6_n60), .A(npu_inst_pe_1_4_6_n74), .ZN(
        npu_inst_pe_1_4_6_n97) );
  NAND2_X1 npu_inst_pe_1_4_6_U85 ( .A1(npu_inst_pe_1_4_6_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_4_6_n60), .ZN(npu_inst_pe_1_4_6_n73) );
  OAI21_X1 npu_inst_pe_1_4_6_U84 ( .B1(npu_inst_pe_1_4_6_n61), .B2(
        npu_inst_pe_1_4_6_n60), .A(npu_inst_pe_1_4_6_n73), .ZN(
        npu_inst_pe_1_4_6_n96) );
  NAND2_X1 npu_inst_pe_1_4_6_U83 ( .A1(npu_inst_pe_1_4_6_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_4_6_n56), .ZN(npu_inst_pe_1_4_6_n72) );
  OAI21_X1 npu_inst_pe_1_4_6_U82 ( .B1(npu_inst_pe_1_4_6_n63), .B2(
        npu_inst_pe_1_4_6_n56), .A(npu_inst_pe_1_4_6_n72), .ZN(
        npu_inst_pe_1_4_6_n95) );
  NAND2_X1 npu_inst_pe_1_4_6_U81 ( .A1(npu_inst_pe_1_4_6_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_4_6_n56), .ZN(npu_inst_pe_1_4_6_n71) );
  OAI21_X1 npu_inst_pe_1_4_6_U80 ( .B1(npu_inst_pe_1_4_6_n61), .B2(
        npu_inst_pe_1_4_6_n56), .A(npu_inst_pe_1_4_6_n71), .ZN(
        npu_inst_pe_1_4_6_n94) );
  NAND2_X1 npu_inst_pe_1_4_6_U79 ( .A1(npu_inst_pe_1_4_6_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_4_6_n52), .ZN(npu_inst_pe_1_4_6_n70) );
  OAI21_X1 npu_inst_pe_1_4_6_U78 ( .B1(npu_inst_pe_1_4_6_n63), .B2(
        npu_inst_pe_1_4_6_n52), .A(npu_inst_pe_1_4_6_n70), .ZN(
        npu_inst_pe_1_4_6_n93) );
  NAND2_X1 npu_inst_pe_1_4_6_U77 ( .A1(npu_inst_pe_1_4_6_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_4_6_n52), .ZN(npu_inst_pe_1_4_6_n69) );
  OAI21_X1 npu_inst_pe_1_4_6_U76 ( .B1(npu_inst_pe_1_4_6_n61), .B2(
        npu_inst_pe_1_4_6_n52), .A(npu_inst_pe_1_4_6_n69), .ZN(
        npu_inst_pe_1_4_6_n92) );
  NAND2_X1 npu_inst_pe_1_4_6_U75 ( .A1(npu_inst_pe_1_4_6_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_4_6_n48), .ZN(npu_inst_pe_1_4_6_n68) );
  OAI21_X1 npu_inst_pe_1_4_6_U74 ( .B1(npu_inst_pe_1_4_6_n63), .B2(
        npu_inst_pe_1_4_6_n48), .A(npu_inst_pe_1_4_6_n68), .ZN(
        npu_inst_pe_1_4_6_n91) );
  NAND2_X1 npu_inst_pe_1_4_6_U73 ( .A1(npu_inst_pe_1_4_6_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_4_6_n48), .ZN(npu_inst_pe_1_4_6_n67) );
  OAI21_X1 npu_inst_pe_1_4_6_U72 ( .B1(npu_inst_pe_1_4_6_n61), .B2(
        npu_inst_pe_1_4_6_n48), .A(npu_inst_pe_1_4_6_n67), .ZN(
        npu_inst_pe_1_4_6_n90) );
  NAND2_X1 npu_inst_pe_1_4_6_U71 ( .A1(npu_inst_pe_1_4_6_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_4_6_n44), .ZN(npu_inst_pe_1_4_6_n66) );
  OAI21_X1 npu_inst_pe_1_4_6_U70 ( .B1(npu_inst_pe_1_4_6_n63), .B2(
        npu_inst_pe_1_4_6_n44), .A(npu_inst_pe_1_4_6_n66), .ZN(
        npu_inst_pe_1_4_6_n89) );
  NAND2_X1 npu_inst_pe_1_4_6_U69 ( .A1(npu_inst_pe_1_4_6_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_4_6_n44), .ZN(npu_inst_pe_1_4_6_n65) );
  OAI21_X1 npu_inst_pe_1_4_6_U68 ( .B1(npu_inst_pe_1_4_6_n61), .B2(
        npu_inst_pe_1_4_6_n44), .A(npu_inst_pe_1_4_6_n65), .ZN(
        npu_inst_pe_1_4_6_n88) );
  NAND2_X1 npu_inst_pe_1_4_6_U67 ( .A1(npu_inst_pe_1_4_6_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_4_6_n40), .ZN(npu_inst_pe_1_4_6_n64) );
  OAI21_X1 npu_inst_pe_1_4_6_U66 ( .B1(npu_inst_pe_1_4_6_n63), .B2(
        npu_inst_pe_1_4_6_n40), .A(npu_inst_pe_1_4_6_n64), .ZN(
        npu_inst_pe_1_4_6_n87) );
  NAND2_X1 npu_inst_pe_1_4_6_U65 ( .A1(npu_inst_pe_1_4_6_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_4_6_n40), .ZN(npu_inst_pe_1_4_6_n62) );
  OAI21_X1 npu_inst_pe_1_4_6_U64 ( .B1(npu_inst_pe_1_4_6_n61), .B2(
        npu_inst_pe_1_4_6_n40), .A(npu_inst_pe_1_4_6_n62), .ZN(
        npu_inst_pe_1_4_6_n86) );
  AND2_X1 npu_inst_pe_1_4_6_U63 ( .A1(npu_inst_pe_1_4_6_N93), .A2(npu_inst_n55), .ZN(npu_inst_int_data_y_4__6__0_) );
  AND2_X1 npu_inst_pe_1_4_6_U62 ( .A1(npu_inst_n55), .A2(npu_inst_pe_1_4_6_N94), .ZN(npu_inst_int_data_y_4__6__1_) );
  NOR3_X1 npu_inst_pe_1_4_6_U61 ( .A1(npu_inst_pe_1_4_6_n26), .A2(npu_inst_n55), .A3(npu_inst_int_ckg[25]), .ZN(npu_inst_pe_1_4_6_n85) );
  OR2_X1 npu_inst_pe_1_4_6_U60 ( .A1(npu_inst_pe_1_4_6_n85), .A2(
        npu_inst_pe_1_4_6_n2), .ZN(npu_inst_pe_1_4_6_N84) );
  AND2_X1 npu_inst_pe_1_4_6_U59 ( .A1(npu_inst_pe_1_4_6_int_q_acc_0_), .A2(
        npu_inst_pe_1_4_6_n1), .ZN(npu_inst_int_data_res_4__6__0_) );
  AND2_X1 npu_inst_pe_1_4_6_U58 ( .A1(npu_inst_pe_1_4_6_n2), .A2(
        npu_inst_pe_1_4_6_int_q_acc_7_), .ZN(npu_inst_int_data_res_4__6__7_)
         );
  AND2_X1 npu_inst_pe_1_4_6_U57 ( .A1(npu_inst_pe_1_4_6_int_q_acc_1_), .A2(
        npu_inst_pe_1_4_6_n1), .ZN(npu_inst_int_data_res_4__6__1_) );
  AND2_X1 npu_inst_pe_1_4_6_U56 ( .A1(npu_inst_pe_1_4_6_int_q_acc_2_), .A2(
        npu_inst_pe_1_4_6_n1), .ZN(npu_inst_int_data_res_4__6__2_) );
  AND2_X1 npu_inst_pe_1_4_6_U55 ( .A1(npu_inst_pe_1_4_6_int_q_acc_3_), .A2(
        npu_inst_pe_1_4_6_n2), .ZN(npu_inst_int_data_res_4__6__3_) );
  AND2_X1 npu_inst_pe_1_4_6_U54 ( .A1(npu_inst_pe_1_4_6_int_q_acc_4_), .A2(
        npu_inst_pe_1_4_6_n2), .ZN(npu_inst_int_data_res_4__6__4_) );
  AND2_X1 npu_inst_pe_1_4_6_U53 ( .A1(npu_inst_pe_1_4_6_int_q_acc_5_), .A2(
        npu_inst_pe_1_4_6_n2), .ZN(npu_inst_int_data_res_4__6__5_) );
  AND2_X1 npu_inst_pe_1_4_6_U52 ( .A1(npu_inst_pe_1_4_6_int_q_acc_6_), .A2(
        npu_inst_pe_1_4_6_n2), .ZN(npu_inst_int_data_res_4__6__6_) );
  AOI222_X1 npu_inst_pe_1_4_6_U51 ( .A1(npu_inst_int_data_res_5__6__0_), .A2(
        npu_inst_pe_1_4_6_n1), .B1(npu_inst_pe_1_4_6_N73), .B2(
        npu_inst_pe_1_4_6_n76), .C1(npu_inst_pe_1_4_6_N65), .C2(
        npu_inst_pe_1_4_6_n77), .ZN(npu_inst_pe_1_4_6_n84) );
  INV_X1 npu_inst_pe_1_4_6_U50 ( .A(npu_inst_pe_1_4_6_n84), .ZN(
        npu_inst_pe_1_4_6_n101) );
  AOI222_X1 npu_inst_pe_1_4_6_U49 ( .A1(npu_inst_int_data_res_5__6__7_), .A2(
        npu_inst_pe_1_4_6_n1), .B1(npu_inst_pe_1_4_6_N80), .B2(
        npu_inst_pe_1_4_6_n76), .C1(npu_inst_pe_1_4_6_N72), .C2(
        npu_inst_pe_1_4_6_n77), .ZN(npu_inst_pe_1_4_6_n75) );
  INV_X1 npu_inst_pe_1_4_6_U48 ( .A(npu_inst_pe_1_4_6_n75), .ZN(
        npu_inst_pe_1_4_6_n33) );
  AOI222_X1 npu_inst_pe_1_4_6_U47 ( .A1(npu_inst_int_data_res_5__6__1_), .A2(
        npu_inst_pe_1_4_6_n1), .B1(npu_inst_pe_1_4_6_N74), .B2(
        npu_inst_pe_1_4_6_n76), .C1(npu_inst_pe_1_4_6_N66), .C2(
        npu_inst_pe_1_4_6_n77), .ZN(npu_inst_pe_1_4_6_n83) );
  INV_X1 npu_inst_pe_1_4_6_U46 ( .A(npu_inst_pe_1_4_6_n83), .ZN(
        npu_inst_pe_1_4_6_n100) );
  AOI222_X1 npu_inst_pe_1_4_6_U45 ( .A1(npu_inst_int_data_res_5__6__2_), .A2(
        npu_inst_pe_1_4_6_n1), .B1(npu_inst_pe_1_4_6_N75), .B2(
        npu_inst_pe_1_4_6_n76), .C1(npu_inst_pe_1_4_6_N67), .C2(
        npu_inst_pe_1_4_6_n77), .ZN(npu_inst_pe_1_4_6_n82) );
  INV_X1 npu_inst_pe_1_4_6_U44 ( .A(npu_inst_pe_1_4_6_n82), .ZN(
        npu_inst_pe_1_4_6_n99) );
  AOI222_X1 npu_inst_pe_1_4_6_U43 ( .A1(npu_inst_int_data_res_5__6__3_), .A2(
        npu_inst_pe_1_4_6_n1), .B1(npu_inst_pe_1_4_6_N76), .B2(
        npu_inst_pe_1_4_6_n76), .C1(npu_inst_pe_1_4_6_N68), .C2(
        npu_inst_pe_1_4_6_n77), .ZN(npu_inst_pe_1_4_6_n81) );
  INV_X1 npu_inst_pe_1_4_6_U42 ( .A(npu_inst_pe_1_4_6_n81), .ZN(
        npu_inst_pe_1_4_6_n98) );
  AOI222_X1 npu_inst_pe_1_4_6_U41 ( .A1(npu_inst_int_data_res_5__6__4_), .A2(
        npu_inst_pe_1_4_6_n1), .B1(npu_inst_pe_1_4_6_N77), .B2(
        npu_inst_pe_1_4_6_n76), .C1(npu_inst_pe_1_4_6_N69), .C2(
        npu_inst_pe_1_4_6_n77), .ZN(npu_inst_pe_1_4_6_n80) );
  INV_X1 npu_inst_pe_1_4_6_U40 ( .A(npu_inst_pe_1_4_6_n80), .ZN(
        npu_inst_pe_1_4_6_n36) );
  AOI222_X1 npu_inst_pe_1_4_6_U39 ( .A1(npu_inst_int_data_res_5__6__5_), .A2(
        npu_inst_pe_1_4_6_n1), .B1(npu_inst_pe_1_4_6_N78), .B2(
        npu_inst_pe_1_4_6_n76), .C1(npu_inst_pe_1_4_6_N70), .C2(
        npu_inst_pe_1_4_6_n77), .ZN(npu_inst_pe_1_4_6_n79) );
  INV_X1 npu_inst_pe_1_4_6_U38 ( .A(npu_inst_pe_1_4_6_n79), .ZN(
        npu_inst_pe_1_4_6_n35) );
  AOI222_X1 npu_inst_pe_1_4_6_U37 ( .A1(npu_inst_int_data_res_5__6__6_), .A2(
        npu_inst_pe_1_4_6_n1), .B1(npu_inst_pe_1_4_6_N79), .B2(
        npu_inst_pe_1_4_6_n76), .C1(npu_inst_pe_1_4_6_N71), .C2(
        npu_inst_pe_1_4_6_n77), .ZN(npu_inst_pe_1_4_6_n78) );
  INV_X1 npu_inst_pe_1_4_6_U36 ( .A(npu_inst_pe_1_4_6_n78), .ZN(
        npu_inst_pe_1_4_6_n34) );
  INV_X1 npu_inst_pe_1_4_6_U35 ( .A(npu_inst_pe_1_4_6_int_data_1_), .ZN(
        npu_inst_pe_1_4_6_n14) );
  AND2_X1 npu_inst_pe_1_4_6_U34 ( .A1(npu_inst_int_data_x_4__6__1_), .A2(
        npu_inst_pe_1_4_6_int_q_weight_1_), .ZN(npu_inst_pe_1_4_6_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_4_6_U33 ( .A1(npu_inst_int_data_x_4__6__0_), .A2(
        npu_inst_pe_1_4_6_int_q_weight_1_), .ZN(npu_inst_pe_1_4_6_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_4_6_U32 ( .A1(npu_inst_n55), .A2(
        npu_inst_int_data_y_5__6__1_), .B1(npu_inst_pe_1_4_6_n3), .B2(
        npu_inst_int_data_x_4__7__1_), .ZN(npu_inst_pe_1_4_6_n63) );
  AOI22_X1 npu_inst_pe_1_4_6_U31 ( .A1(npu_inst_n55), .A2(
        npu_inst_int_data_y_5__6__0_), .B1(npu_inst_pe_1_4_6_n3), .B2(
        npu_inst_int_data_x_4__7__0_), .ZN(npu_inst_pe_1_4_6_n61) );
  INV_X1 npu_inst_pe_1_4_6_U30 ( .A(npu_inst_pe_1_4_6_int_data_0_), .ZN(
        npu_inst_pe_1_4_6_n13) );
  INV_X1 npu_inst_pe_1_4_6_U29 ( .A(npu_inst_n69), .ZN(npu_inst_pe_1_4_6_n5)
         );
  OR3_X1 npu_inst_pe_1_4_6_U28 ( .A1(npu_inst_pe_1_4_6_n6), .A2(
        npu_inst_pe_1_4_6_n8), .A3(npu_inst_pe_1_4_6_n5), .ZN(
        npu_inst_pe_1_4_6_n56) );
  OR3_X1 npu_inst_pe_1_4_6_U27 ( .A1(npu_inst_pe_1_4_6_n5), .A2(
        npu_inst_pe_1_4_6_n8), .A3(npu_inst_pe_1_4_6_n7), .ZN(
        npu_inst_pe_1_4_6_n48) );
  INV_X1 npu_inst_pe_1_4_6_U26 ( .A(npu_inst_pe_1_4_6_n5), .ZN(
        npu_inst_pe_1_4_6_n4) );
  INV_X1 npu_inst_pe_1_4_6_U25 ( .A(npu_inst_n124), .ZN(npu_inst_pe_1_4_6_n12)
         );
  OR3_X1 npu_inst_pe_1_4_6_U24 ( .A1(npu_inst_pe_1_4_6_n4), .A2(
        npu_inst_pe_1_4_6_n8), .A3(npu_inst_pe_1_4_6_n7), .ZN(
        npu_inst_pe_1_4_6_n52) );
  OR3_X1 npu_inst_pe_1_4_6_U23 ( .A1(npu_inst_pe_1_4_6_n6), .A2(
        npu_inst_pe_1_4_6_n8), .A3(npu_inst_pe_1_4_6_n4), .ZN(
        npu_inst_pe_1_4_6_n60) );
  NOR2_X1 npu_inst_pe_1_4_6_U22 ( .A1(npu_inst_pe_1_4_6_n60), .A2(
        npu_inst_pe_1_4_6_n3), .ZN(npu_inst_pe_1_4_6_n58) );
  NOR2_X1 npu_inst_pe_1_4_6_U21 ( .A1(npu_inst_pe_1_4_6_n56), .A2(
        npu_inst_pe_1_4_6_n3), .ZN(npu_inst_pe_1_4_6_n54) );
  NOR2_X1 npu_inst_pe_1_4_6_U20 ( .A1(npu_inst_pe_1_4_6_n52), .A2(
        npu_inst_pe_1_4_6_n3), .ZN(npu_inst_pe_1_4_6_n50) );
  NOR2_X1 npu_inst_pe_1_4_6_U19 ( .A1(npu_inst_pe_1_4_6_n48), .A2(
        npu_inst_pe_1_4_6_n3), .ZN(npu_inst_pe_1_4_6_n46) );
  NOR2_X1 npu_inst_pe_1_4_6_U18 ( .A1(npu_inst_pe_1_4_6_n40), .A2(
        npu_inst_pe_1_4_6_n3), .ZN(npu_inst_pe_1_4_6_n38) );
  NOR2_X1 npu_inst_pe_1_4_6_U17 ( .A1(npu_inst_pe_1_4_6_n44), .A2(
        npu_inst_pe_1_4_6_n3), .ZN(npu_inst_pe_1_4_6_n42) );
  BUF_X1 npu_inst_pe_1_4_6_U16 ( .A(npu_inst_n98), .Z(npu_inst_pe_1_4_6_n8) );
  BUF_X1 npu_inst_pe_1_4_6_U15 ( .A(npu_inst_pe_1_4_6_n12), .Z(
        npu_inst_pe_1_4_6_n11) );
  BUF_X1 npu_inst_pe_1_4_6_U14 ( .A(npu_inst_pe_1_4_6_n12), .Z(
        npu_inst_pe_1_4_6_n10) );
  BUF_X1 npu_inst_pe_1_4_6_U13 ( .A(npu_inst_pe_1_4_6_n12), .Z(
        npu_inst_pe_1_4_6_n9) );
  INV_X1 npu_inst_pe_1_4_6_U12 ( .A(npu_inst_pe_1_4_6_n38), .ZN(
        npu_inst_pe_1_4_6_n118) );
  INV_X1 npu_inst_pe_1_4_6_U11 ( .A(npu_inst_pe_1_4_6_n58), .ZN(
        npu_inst_pe_1_4_6_n114) );
  INV_X1 npu_inst_pe_1_4_6_U10 ( .A(npu_inst_pe_1_4_6_n54), .ZN(
        npu_inst_pe_1_4_6_n115) );
  INV_X1 npu_inst_pe_1_4_6_U9 ( .A(npu_inst_pe_1_4_6_n50), .ZN(
        npu_inst_pe_1_4_6_n116) );
  INV_X1 npu_inst_pe_1_4_6_U8 ( .A(npu_inst_pe_1_4_6_n46), .ZN(
        npu_inst_pe_1_4_6_n117) );
  INV_X1 npu_inst_pe_1_4_6_U7 ( .A(npu_inst_pe_1_4_6_n42), .ZN(
        npu_inst_pe_1_4_6_n119) );
  BUF_X1 npu_inst_pe_1_4_6_U6 ( .A(npu_inst_n19), .Z(npu_inst_pe_1_4_6_n2) );
  BUF_X1 npu_inst_pe_1_4_6_U5 ( .A(npu_inst_n19), .Z(npu_inst_pe_1_4_6_n1) );
  NOR2_X1 npu_inst_pe_1_4_6_U4 ( .A1(npu_inst_pe_1_4_6_int_q_weight_0_), .A2(
        npu_inst_pe_1_4_6_n1), .ZN(npu_inst_pe_1_4_6_n76) );
  NOR2_X1 npu_inst_pe_1_4_6_U3 ( .A1(npu_inst_pe_1_4_6_n27), .A2(
        npu_inst_pe_1_4_6_n1), .ZN(npu_inst_pe_1_4_6_n77) );
  FA_X1 npu_inst_pe_1_4_6_sub_77_U2_1 ( .A(npu_inst_pe_1_4_6_int_q_acc_1_), 
        .B(npu_inst_pe_1_4_6_n14), .CI(npu_inst_pe_1_4_6_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_4_6_sub_77_carry_2_), .S(npu_inst_pe_1_4_6_N66) );
  FA_X1 npu_inst_pe_1_4_6_add_79_U1_1 ( .A(npu_inst_pe_1_4_6_int_q_acc_1_), 
        .B(npu_inst_pe_1_4_6_int_data_1_), .CI(
        npu_inst_pe_1_4_6_add_79_carry_1_), .CO(
        npu_inst_pe_1_4_6_add_79_carry_2_), .S(npu_inst_pe_1_4_6_N74) );
  NAND3_X1 npu_inst_pe_1_4_6_U109 ( .A1(npu_inst_pe_1_4_6_n5), .A2(
        npu_inst_pe_1_4_6_n7), .A3(npu_inst_pe_1_4_6_n8), .ZN(
        npu_inst_pe_1_4_6_n44) );
  NAND3_X1 npu_inst_pe_1_4_6_U108 ( .A1(npu_inst_pe_1_4_6_n4), .A2(
        npu_inst_pe_1_4_6_n7), .A3(npu_inst_pe_1_4_6_n8), .ZN(
        npu_inst_pe_1_4_6_n40) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_4_6_n34), .CK(
        npu_inst_pe_1_4_6_net3419), .RN(npu_inst_pe_1_4_6_n9), .Q(
        npu_inst_pe_1_4_6_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_4_6_n35), .CK(
        npu_inst_pe_1_4_6_net3419), .RN(npu_inst_pe_1_4_6_n9), .Q(
        npu_inst_pe_1_4_6_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_4_6_n36), .CK(
        npu_inst_pe_1_4_6_net3419), .RN(npu_inst_pe_1_4_6_n9), .Q(
        npu_inst_pe_1_4_6_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_4_6_n98), .CK(
        npu_inst_pe_1_4_6_net3419), .RN(npu_inst_pe_1_4_6_n9), .Q(
        npu_inst_pe_1_4_6_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_4_6_n99), .CK(
        npu_inst_pe_1_4_6_net3419), .RN(npu_inst_pe_1_4_6_n9), .Q(
        npu_inst_pe_1_4_6_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_4_6_n100), 
        .CK(npu_inst_pe_1_4_6_net3419), .RN(npu_inst_pe_1_4_6_n9), .Q(
        npu_inst_pe_1_4_6_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_4_6_n33), .CK(
        npu_inst_pe_1_4_6_net3419), .RN(npu_inst_pe_1_4_6_n9), .Q(
        npu_inst_pe_1_4_6_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_4_6_n101), 
        .CK(npu_inst_pe_1_4_6_net3419), .RN(npu_inst_pe_1_4_6_n9), .Q(
        npu_inst_pe_1_4_6_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_weight_reg_0_ ( .D(npu_inst_n110), .CK(
        npu_inst_pe_1_4_6_net3425), .RN(npu_inst_pe_1_4_6_n9), .Q(
        npu_inst_pe_1_4_6_int_q_weight_0_), .QN(npu_inst_pe_1_4_6_n27) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_weight_reg_1_ ( .D(npu_inst_n116), .CK(
        npu_inst_pe_1_4_6_net3425), .RN(npu_inst_pe_1_4_6_n9), .Q(
        npu_inst_pe_1_4_6_int_q_weight_1_), .QN(npu_inst_pe_1_4_6_n26) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_4_6_n113), 
        .CK(npu_inst_pe_1_4_6_net3425), .RN(npu_inst_pe_1_4_6_n9), .Q(
        npu_inst_pe_1_4_6_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_4_6_n107), 
        .CK(npu_inst_pe_1_4_6_net3425), .RN(npu_inst_pe_1_4_6_n9), .Q(
        npu_inst_pe_1_4_6_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_4_6_n112), 
        .CK(npu_inst_pe_1_4_6_net3425), .RN(npu_inst_pe_1_4_6_n10), .Q(
        npu_inst_pe_1_4_6_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_4_6_n106), 
        .CK(npu_inst_pe_1_4_6_net3425), .RN(npu_inst_pe_1_4_6_n10), .Q(
        npu_inst_pe_1_4_6_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_4_6_n111), 
        .CK(npu_inst_pe_1_4_6_net3425), .RN(npu_inst_pe_1_4_6_n10), .Q(
        npu_inst_pe_1_4_6_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_4_6_n105), 
        .CK(npu_inst_pe_1_4_6_net3425), .RN(npu_inst_pe_1_4_6_n10), .Q(
        npu_inst_pe_1_4_6_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_4_6_n110), 
        .CK(npu_inst_pe_1_4_6_net3425), .RN(npu_inst_pe_1_4_6_n10), .Q(
        npu_inst_pe_1_4_6_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_4_6_n104), 
        .CK(npu_inst_pe_1_4_6_net3425), .RN(npu_inst_pe_1_4_6_n10), .Q(
        npu_inst_pe_1_4_6_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_4_6_n109), 
        .CK(npu_inst_pe_1_4_6_net3425), .RN(npu_inst_pe_1_4_6_n10), .Q(
        npu_inst_pe_1_4_6_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_4_6_n103), 
        .CK(npu_inst_pe_1_4_6_net3425), .RN(npu_inst_pe_1_4_6_n10), .Q(
        npu_inst_pe_1_4_6_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_4_6_n108), 
        .CK(npu_inst_pe_1_4_6_net3425), .RN(npu_inst_pe_1_4_6_n10), .Q(
        npu_inst_pe_1_4_6_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_4_6_n102), 
        .CK(npu_inst_pe_1_4_6_net3425), .RN(npu_inst_pe_1_4_6_n10), .Q(
        npu_inst_pe_1_4_6_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_4_6_n86), 
        .CK(npu_inst_pe_1_4_6_net3425), .RN(npu_inst_pe_1_4_6_n10), .Q(
        npu_inst_pe_1_4_6_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_4_6_n87), 
        .CK(npu_inst_pe_1_4_6_net3425), .RN(npu_inst_pe_1_4_6_n10), .Q(
        npu_inst_pe_1_4_6_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_4_6_n88), 
        .CK(npu_inst_pe_1_4_6_net3425), .RN(npu_inst_pe_1_4_6_n11), .Q(
        npu_inst_pe_1_4_6_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_4_6_n89), 
        .CK(npu_inst_pe_1_4_6_net3425), .RN(npu_inst_pe_1_4_6_n11), .Q(
        npu_inst_pe_1_4_6_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_4_6_n90), 
        .CK(npu_inst_pe_1_4_6_net3425), .RN(npu_inst_pe_1_4_6_n11), .Q(
        npu_inst_pe_1_4_6_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_4_6_n91), 
        .CK(npu_inst_pe_1_4_6_net3425), .RN(npu_inst_pe_1_4_6_n11), .Q(
        npu_inst_pe_1_4_6_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_4_6_n92), 
        .CK(npu_inst_pe_1_4_6_net3425), .RN(npu_inst_pe_1_4_6_n11), .Q(
        npu_inst_pe_1_4_6_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_4_6_n93), 
        .CK(npu_inst_pe_1_4_6_net3425), .RN(npu_inst_pe_1_4_6_n11), .Q(
        npu_inst_pe_1_4_6_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_4_6_n94), 
        .CK(npu_inst_pe_1_4_6_net3425), .RN(npu_inst_pe_1_4_6_n11), .Q(
        npu_inst_pe_1_4_6_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_4_6_n95), 
        .CK(npu_inst_pe_1_4_6_net3425), .RN(npu_inst_pe_1_4_6_n11), .Q(
        npu_inst_pe_1_4_6_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_4_6_n96), 
        .CK(npu_inst_pe_1_4_6_net3425), .RN(npu_inst_pe_1_4_6_n11), .Q(
        npu_inst_pe_1_4_6_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_4_6_n97), 
        .CK(npu_inst_pe_1_4_6_net3425), .RN(npu_inst_pe_1_4_6_n11), .Q(
        npu_inst_pe_1_4_6_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_4_6_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_4_6_N84), .SE(1'b0), .GCK(npu_inst_pe_1_4_6_net3419) );
  CLKGATETST_X1 npu_inst_pe_1_4_6_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n63), .SE(1'b0), .GCK(npu_inst_pe_1_4_6_net3425) );
  MUX2_X1 npu_inst_pe_1_4_7_U162 ( .A(npu_inst_pe_1_4_7_n32), .B(
        npu_inst_pe_1_4_7_n29), .S(npu_inst_pe_1_4_7_n8), .Z(
        npu_inst_pe_1_4_7_N93) );
  MUX2_X1 npu_inst_pe_1_4_7_U161 ( .A(npu_inst_pe_1_4_7_n31), .B(
        npu_inst_pe_1_4_7_n30), .S(npu_inst_pe_1_4_7_n6), .Z(
        npu_inst_pe_1_4_7_n32) );
  MUX2_X1 npu_inst_pe_1_4_7_U160 ( .A(npu_inst_pe_1_4_7_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_4_7_int_q_reg_v_1__0_), .S(npu_inst_pe_1_4_7_n4), .Z(
        npu_inst_pe_1_4_7_n31) );
  MUX2_X1 npu_inst_pe_1_4_7_U159 ( .A(npu_inst_pe_1_4_7_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_4_7_int_q_reg_v_3__0_), .S(npu_inst_pe_1_4_7_n4), .Z(
        npu_inst_pe_1_4_7_n30) );
  MUX2_X1 npu_inst_pe_1_4_7_U158 ( .A(npu_inst_pe_1_4_7_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_4_7_int_q_reg_v_5__0_), .S(npu_inst_pe_1_4_7_n4), .Z(
        npu_inst_pe_1_4_7_n29) );
  MUX2_X1 npu_inst_pe_1_4_7_U157 ( .A(npu_inst_pe_1_4_7_n28), .B(
        npu_inst_pe_1_4_7_n23), .S(npu_inst_pe_1_4_7_n8), .Z(
        npu_inst_pe_1_4_7_N94) );
  MUX2_X1 npu_inst_pe_1_4_7_U156 ( .A(npu_inst_pe_1_4_7_n25), .B(
        npu_inst_pe_1_4_7_n24), .S(npu_inst_pe_1_4_7_n6), .Z(
        npu_inst_pe_1_4_7_n28) );
  MUX2_X1 npu_inst_pe_1_4_7_U155 ( .A(npu_inst_pe_1_4_7_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_4_7_int_q_reg_v_1__1_), .S(npu_inst_pe_1_4_7_n4), .Z(
        npu_inst_pe_1_4_7_n25) );
  MUX2_X1 npu_inst_pe_1_4_7_U154 ( .A(npu_inst_pe_1_4_7_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_4_7_int_q_reg_v_3__1_), .S(npu_inst_pe_1_4_7_n4), .Z(
        npu_inst_pe_1_4_7_n24) );
  MUX2_X1 npu_inst_pe_1_4_7_U153 ( .A(npu_inst_pe_1_4_7_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_4_7_int_q_reg_v_5__1_), .S(npu_inst_pe_1_4_7_n4), .Z(
        npu_inst_pe_1_4_7_n23) );
  MUX2_X1 npu_inst_pe_1_4_7_U152 ( .A(npu_inst_pe_1_4_7_n22), .B(
        npu_inst_pe_1_4_7_n19), .S(npu_inst_pe_1_4_7_n8), .Z(
        npu_inst_int_data_x_4__7__1_) );
  MUX2_X1 npu_inst_pe_1_4_7_U151 ( .A(npu_inst_pe_1_4_7_n21), .B(
        npu_inst_pe_1_4_7_n20), .S(npu_inst_pe_1_4_7_n6), .Z(
        npu_inst_pe_1_4_7_n22) );
  MUX2_X1 npu_inst_pe_1_4_7_U150 ( .A(npu_inst_pe_1_4_7_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_4_7_int_q_reg_h_1__1_), .S(npu_inst_pe_1_4_7_n4), .Z(
        npu_inst_pe_1_4_7_n21) );
  MUX2_X1 npu_inst_pe_1_4_7_U149 ( .A(npu_inst_pe_1_4_7_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_4_7_int_q_reg_h_3__1_), .S(npu_inst_pe_1_4_7_n4), .Z(
        npu_inst_pe_1_4_7_n20) );
  MUX2_X1 npu_inst_pe_1_4_7_U148 ( .A(npu_inst_pe_1_4_7_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_4_7_int_q_reg_h_5__1_), .S(npu_inst_pe_1_4_7_n4), .Z(
        npu_inst_pe_1_4_7_n19) );
  MUX2_X1 npu_inst_pe_1_4_7_U147 ( .A(npu_inst_pe_1_4_7_n18), .B(
        npu_inst_pe_1_4_7_n15), .S(npu_inst_pe_1_4_7_n8), .Z(
        npu_inst_int_data_x_4__7__0_) );
  MUX2_X1 npu_inst_pe_1_4_7_U146 ( .A(npu_inst_pe_1_4_7_n17), .B(
        npu_inst_pe_1_4_7_n16), .S(npu_inst_pe_1_4_7_n6), .Z(
        npu_inst_pe_1_4_7_n18) );
  MUX2_X1 npu_inst_pe_1_4_7_U145 ( .A(npu_inst_pe_1_4_7_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_4_7_int_q_reg_h_1__0_), .S(npu_inst_pe_1_4_7_n4), .Z(
        npu_inst_pe_1_4_7_n17) );
  MUX2_X1 npu_inst_pe_1_4_7_U144 ( .A(npu_inst_pe_1_4_7_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_4_7_int_q_reg_h_3__0_), .S(npu_inst_pe_1_4_7_n4), .Z(
        npu_inst_pe_1_4_7_n16) );
  MUX2_X1 npu_inst_pe_1_4_7_U143 ( .A(npu_inst_pe_1_4_7_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_4_7_int_q_reg_h_5__0_), .S(npu_inst_pe_1_4_7_n4), .Z(
        npu_inst_pe_1_4_7_n15) );
  XOR2_X1 npu_inst_pe_1_4_7_U142 ( .A(npu_inst_pe_1_4_7_int_data_0_), .B(
        npu_inst_pe_1_4_7_int_q_acc_0_), .Z(npu_inst_pe_1_4_7_N73) );
  AND2_X1 npu_inst_pe_1_4_7_U141 ( .A1(npu_inst_pe_1_4_7_int_q_acc_0_), .A2(
        npu_inst_pe_1_4_7_int_data_0_), .ZN(npu_inst_pe_1_4_7_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_4_7_U140 ( .A(npu_inst_pe_1_4_7_int_q_acc_0_), .B(
        npu_inst_pe_1_4_7_n13), .ZN(npu_inst_pe_1_4_7_N65) );
  OR2_X1 npu_inst_pe_1_4_7_U139 ( .A1(npu_inst_pe_1_4_7_n13), .A2(
        npu_inst_pe_1_4_7_int_q_acc_0_), .ZN(npu_inst_pe_1_4_7_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_4_7_U138 ( .A(npu_inst_pe_1_4_7_int_q_acc_2_), .B(
        npu_inst_pe_1_4_7_add_79_carry_2_), .Z(npu_inst_pe_1_4_7_N75) );
  AND2_X1 npu_inst_pe_1_4_7_U137 ( .A1(npu_inst_pe_1_4_7_add_79_carry_2_), 
        .A2(npu_inst_pe_1_4_7_int_q_acc_2_), .ZN(
        npu_inst_pe_1_4_7_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_4_7_U136 ( .A(npu_inst_pe_1_4_7_int_q_acc_3_), .B(
        npu_inst_pe_1_4_7_add_79_carry_3_), .Z(npu_inst_pe_1_4_7_N76) );
  AND2_X1 npu_inst_pe_1_4_7_U135 ( .A1(npu_inst_pe_1_4_7_add_79_carry_3_), 
        .A2(npu_inst_pe_1_4_7_int_q_acc_3_), .ZN(
        npu_inst_pe_1_4_7_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_4_7_U134 ( .A(npu_inst_pe_1_4_7_int_q_acc_4_), .B(
        npu_inst_pe_1_4_7_add_79_carry_4_), .Z(npu_inst_pe_1_4_7_N77) );
  AND2_X1 npu_inst_pe_1_4_7_U133 ( .A1(npu_inst_pe_1_4_7_add_79_carry_4_), 
        .A2(npu_inst_pe_1_4_7_int_q_acc_4_), .ZN(
        npu_inst_pe_1_4_7_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_4_7_U132 ( .A(npu_inst_pe_1_4_7_int_q_acc_5_), .B(
        npu_inst_pe_1_4_7_add_79_carry_5_), .Z(npu_inst_pe_1_4_7_N78) );
  AND2_X1 npu_inst_pe_1_4_7_U131 ( .A1(npu_inst_pe_1_4_7_add_79_carry_5_), 
        .A2(npu_inst_pe_1_4_7_int_q_acc_5_), .ZN(
        npu_inst_pe_1_4_7_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_4_7_U130 ( .A(npu_inst_pe_1_4_7_int_q_acc_6_), .B(
        npu_inst_pe_1_4_7_add_79_carry_6_), .Z(npu_inst_pe_1_4_7_N79) );
  AND2_X1 npu_inst_pe_1_4_7_U129 ( .A1(npu_inst_pe_1_4_7_add_79_carry_6_), 
        .A2(npu_inst_pe_1_4_7_int_q_acc_6_), .ZN(
        npu_inst_pe_1_4_7_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_4_7_U128 ( .A(npu_inst_pe_1_4_7_int_q_acc_7_), .B(
        npu_inst_pe_1_4_7_add_79_carry_7_), .Z(npu_inst_pe_1_4_7_N80) );
  XNOR2_X1 npu_inst_pe_1_4_7_U127 ( .A(npu_inst_pe_1_4_7_sub_77_carry_2_), .B(
        npu_inst_pe_1_4_7_int_q_acc_2_), .ZN(npu_inst_pe_1_4_7_N67) );
  OR2_X1 npu_inst_pe_1_4_7_U126 ( .A1(npu_inst_pe_1_4_7_int_q_acc_2_), .A2(
        npu_inst_pe_1_4_7_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_4_7_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_4_7_U125 ( .A(npu_inst_pe_1_4_7_sub_77_carry_3_), .B(
        npu_inst_pe_1_4_7_int_q_acc_3_), .ZN(npu_inst_pe_1_4_7_N68) );
  OR2_X1 npu_inst_pe_1_4_7_U124 ( .A1(npu_inst_pe_1_4_7_int_q_acc_3_), .A2(
        npu_inst_pe_1_4_7_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_4_7_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_4_7_U123 ( .A(npu_inst_pe_1_4_7_sub_77_carry_4_), .B(
        npu_inst_pe_1_4_7_int_q_acc_4_), .ZN(npu_inst_pe_1_4_7_N69) );
  OR2_X1 npu_inst_pe_1_4_7_U122 ( .A1(npu_inst_pe_1_4_7_int_q_acc_4_), .A2(
        npu_inst_pe_1_4_7_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_4_7_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_4_7_U121 ( .A(npu_inst_pe_1_4_7_sub_77_carry_5_), .B(
        npu_inst_pe_1_4_7_int_q_acc_5_), .ZN(npu_inst_pe_1_4_7_N70) );
  OR2_X1 npu_inst_pe_1_4_7_U120 ( .A1(npu_inst_pe_1_4_7_int_q_acc_5_), .A2(
        npu_inst_pe_1_4_7_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_4_7_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_4_7_U119 ( .A(npu_inst_pe_1_4_7_sub_77_carry_6_), .B(
        npu_inst_pe_1_4_7_int_q_acc_6_), .ZN(npu_inst_pe_1_4_7_N71) );
  OR2_X1 npu_inst_pe_1_4_7_U118 ( .A1(npu_inst_pe_1_4_7_int_q_acc_6_), .A2(
        npu_inst_pe_1_4_7_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_4_7_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_4_7_U117 ( .A(npu_inst_pe_1_4_7_int_q_acc_7_), .B(
        npu_inst_pe_1_4_7_sub_77_carry_7_), .ZN(npu_inst_pe_1_4_7_N72) );
  INV_X1 npu_inst_pe_1_4_7_U116 ( .A(npu_inst_n77), .ZN(npu_inst_pe_1_4_7_n7)
         );
  INV_X1 npu_inst_pe_1_4_7_U115 ( .A(npu_inst_pe_1_4_7_n7), .ZN(
        npu_inst_pe_1_4_7_n6) );
  INV_X1 npu_inst_pe_1_4_7_U114 ( .A(npu_inst_n55), .ZN(npu_inst_pe_1_4_7_n3)
         );
  AOI22_X1 npu_inst_pe_1_4_7_U113 ( .A1(npu_inst_int_data_y_5__7__0_), .A2(
        npu_inst_pe_1_4_7_n58), .B1(npu_inst_pe_1_4_7_n114), .B2(
        npu_inst_pe_1_4_7_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_4_7_n57) );
  INV_X1 npu_inst_pe_1_4_7_U112 ( .A(npu_inst_pe_1_4_7_n57), .ZN(
        npu_inst_pe_1_4_7_n108) );
  AOI22_X1 npu_inst_pe_1_4_7_U111 ( .A1(npu_inst_int_data_y_5__7__0_), .A2(
        npu_inst_pe_1_4_7_n54), .B1(npu_inst_pe_1_4_7_n115), .B2(
        npu_inst_pe_1_4_7_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_4_7_n53) );
  INV_X1 npu_inst_pe_1_4_7_U110 ( .A(npu_inst_pe_1_4_7_n53), .ZN(
        npu_inst_pe_1_4_7_n109) );
  AOI22_X1 npu_inst_pe_1_4_7_U107 ( .A1(npu_inst_int_data_y_5__7__0_), .A2(
        npu_inst_pe_1_4_7_n50), .B1(npu_inst_pe_1_4_7_n116), .B2(
        npu_inst_pe_1_4_7_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_4_7_n49) );
  INV_X1 npu_inst_pe_1_4_7_U106 ( .A(npu_inst_pe_1_4_7_n49), .ZN(
        npu_inst_pe_1_4_7_n110) );
  AOI22_X1 npu_inst_pe_1_4_7_U105 ( .A1(npu_inst_int_data_y_5__7__0_), .A2(
        npu_inst_pe_1_4_7_n46), .B1(npu_inst_pe_1_4_7_n117), .B2(
        npu_inst_pe_1_4_7_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_4_7_n45) );
  INV_X1 npu_inst_pe_1_4_7_U104 ( .A(npu_inst_pe_1_4_7_n45), .ZN(
        npu_inst_pe_1_4_7_n111) );
  AOI22_X1 npu_inst_pe_1_4_7_U103 ( .A1(npu_inst_int_data_y_5__7__0_), .A2(
        npu_inst_pe_1_4_7_n42), .B1(npu_inst_pe_1_4_7_n119), .B2(
        npu_inst_pe_1_4_7_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_4_7_n41) );
  INV_X1 npu_inst_pe_1_4_7_U102 ( .A(npu_inst_pe_1_4_7_n41), .ZN(
        npu_inst_pe_1_4_7_n112) );
  AOI22_X1 npu_inst_pe_1_4_7_U101 ( .A1(npu_inst_int_data_y_5__7__1_), .A2(
        npu_inst_pe_1_4_7_n58), .B1(npu_inst_pe_1_4_7_n114), .B2(
        npu_inst_pe_1_4_7_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_4_7_n59) );
  INV_X1 npu_inst_pe_1_4_7_U100 ( .A(npu_inst_pe_1_4_7_n59), .ZN(
        npu_inst_pe_1_4_7_n102) );
  AOI22_X1 npu_inst_pe_1_4_7_U99 ( .A1(npu_inst_int_data_y_5__7__1_), .A2(
        npu_inst_pe_1_4_7_n54), .B1(npu_inst_pe_1_4_7_n115), .B2(
        npu_inst_pe_1_4_7_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_4_7_n55) );
  INV_X1 npu_inst_pe_1_4_7_U98 ( .A(npu_inst_pe_1_4_7_n55), .ZN(
        npu_inst_pe_1_4_7_n103) );
  AOI22_X1 npu_inst_pe_1_4_7_U97 ( .A1(npu_inst_int_data_y_5__7__1_), .A2(
        npu_inst_pe_1_4_7_n50), .B1(npu_inst_pe_1_4_7_n116), .B2(
        npu_inst_pe_1_4_7_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_4_7_n51) );
  INV_X1 npu_inst_pe_1_4_7_U96 ( .A(npu_inst_pe_1_4_7_n51), .ZN(
        npu_inst_pe_1_4_7_n104) );
  AOI22_X1 npu_inst_pe_1_4_7_U95 ( .A1(npu_inst_int_data_y_5__7__1_), .A2(
        npu_inst_pe_1_4_7_n46), .B1(npu_inst_pe_1_4_7_n117), .B2(
        npu_inst_pe_1_4_7_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_4_7_n47) );
  INV_X1 npu_inst_pe_1_4_7_U94 ( .A(npu_inst_pe_1_4_7_n47), .ZN(
        npu_inst_pe_1_4_7_n105) );
  AOI22_X1 npu_inst_pe_1_4_7_U93 ( .A1(npu_inst_int_data_y_5__7__1_), .A2(
        npu_inst_pe_1_4_7_n42), .B1(npu_inst_pe_1_4_7_n119), .B2(
        npu_inst_pe_1_4_7_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_4_7_n43) );
  INV_X1 npu_inst_pe_1_4_7_U92 ( .A(npu_inst_pe_1_4_7_n43), .ZN(
        npu_inst_pe_1_4_7_n106) );
  AOI22_X1 npu_inst_pe_1_4_7_U91 ( .A1(npu_inst_pe_1_4_7_n38), .A2(
        npu_inst_int_data_y_5__7__1_), .B1(npu_inst_pe_1_4_7_n118), .B2(
        npu_inst_pe_1_4_7_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_4_7_n39) );
  INV_X1 npu_inst_pe_1_4_7_U90 ( .A(npu_inst_pe_1_4_7_n39), .ZN(
        npu_inst_pe_1_4_7_n107) );
  AOI22_X1 npu_inst_pe_1_4_7_U89 ( .A1(npu_inst_pe_1_4_7_n38), .A2(
        npu_inst_int_data_y_5__7__0_), .B1(npu_inst_pe_1_4_7_n118), .B2(
        npu_inst_pe_1_4_7_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_4_7_n37) );
  INV_X1 npu_inst_pe_1_4_7_U88 ( .A(npu_inst_pe_1_4_7_n37), .ZN(
        npu_inst_pe_1_4_7_n113) );
  AND2_X1 npu_inst_pe_1_4_7_U87 ( .A1(npu_inst_pe_1_4_7_N93), .A2(npu_inst_n55), .ZN(npu_inst_int_data_y_4__7__0_) );
  AND2_X1 npu_inst_pe_1_4_7_U86 ( .A1(npu_inst_n55), .A2(npu_inst_pe_1_4_7_N94), .ZN(npu_inst_int_data_y_4__7__1_) );
  NOR3_X1 npu_inst_pe_1_4_7_U85 ( .A1(npu_inst_pe_1_4_7_n26), .A2(npu_inst_n55), .A3(npu_inst_int_ckg[24]), .ZN(npu_inst_pe_1_4_7_n85) );
  OR2_X1 npu_inst_pe_1_4_7_U84 ( .A1(npu_inst_pe_1_4_7_n85), .A2(
        npu_inst_pe_1_4_7_n2), .ZN(npu_inst_pe_1_4_7_N84) );
  AND2_X1 npu_inst_pe_1_4_7_U83 ( .A1(npu_inst_pe_1_4_7_int_q_acc_0_), .A2(
        npu_inst_pe_1_4_7_n1), .ZN(npu_inst_int_data_res_4__7__0_) );
  AND2_X1 npu_inst_pe_1_4_7_U82 ( .A1(npu_inst_pe_1_4_7_n2), .A2(
        npu_inst_pe_1_4_7_int_q_acc_7_), .ZN(npu_inst_int_data_res_4__7__7_)
         );
  AND2_X1 npu_inst_pe_1_4_7_U81 ( .A1(npu_inst_pe_1_4_7_int_q_acc_1_), .A2(
        npu_inst_pe_1_4_7_n1), .ZN(npu_inst_int_data_res_4__7__1_) );
  AND2_X1 npu_inst_pe_1_4_7_U80 ( .A1(npu_inst_pe_1_4_7_int_q_acc_2_), .A2(
        npu_inst_pe_1_4_7_n1), .ZN(npu_inst_int_data_res_4__7__2_) );
  AND2_X1 npu_inst_pe_1_4_7_U79 ( .A1(npu_inst_pe_1_4_7_int_q_acc_3_), .A2(
        npu_inst_pe_1_4_7_n2), .ZN(npu_inst_int_data_res_4__7__3_) );
  AND2_X1 npu_inst_pe_1_4_7_U78 ( .A1(npu_inst_pe_1_4_7_int_q_acc_4_), .A2(
        npu_inst_pe_1_4_7_n2), .ZN(npu_inst_int_data_res_4__7__4_) );
  AND2_X1 npu_inst_pe_1_4_7_U77 ( .A1(npu_inst_pe_1_4_7_int_q_acc_5_), .A2(
        npu_inst_pe_1_4_7_n2), .ZN(npu_inst_int_data_res_4__7__5_) );
  AND2_X1 npu_inst_pe_1_4_7_U76 ( .A1(npu_inst_pe_1_4_7_int_q_acc_6_), .A2(
        npu_inst_pe_1_4_7_n2), .ZN(npu_inst_int_data_res_4__7__6_) );
  AOI222_X1 npu_inst_pe_1_4_7_U75 ( .A1(npu_inst_int_data_res_5__7__0_), .A2(
        npu_inst_pe_1_4_7_n1), .B1(npu_inst_pe_1_4_7_N73), .B2(
        npu_inst_pe_1_4_7_n76), .C1(npu_inst_pe_1_4_7_N65), .C2(
        npu_inst_pe_1_4_7_n77), .ZN(npu_inst_pe_1_4_7_n84) );
  INV_X1 npu_inst_pe_1_4_7_U74 ( .A(npu_inst_pe_1_4_7_n84), .ZN(
        npu_inst_pe_1_4_7_n101) );
  AOI222_X1 npu_inst_pe_1_4_7_U73 ( .A1(npu_inst_int_data_res_5__7__7_), .A2(
        npu_inst_pe_1_4_7_n1), .B1(npu_inst_pe_1_4_7_N80), .B2(
        npu_inst_pe_1_4_7_n76), .C1(npu_inst_pe_1_4_7_N72), .C2(
        npu_inst_pe_1_4_7_n77), .ZN(npu_inst_pe_1_4_7_n75) );
  INV_X1 npu_inst_pe_1_4_7_U72 ( .A(npu_inst_pe_1_4_7_n75), .ZN(
        npu_inst_pe_1_4_7_n33) );
  AOI222_X1 npu_inst_pe_1_4_7_U71 ( .A1(npu_inst_int_data_res_5__7__1_), .A2(
        npu_inst_pe_1_4_7_n1), .B1(npu_inst_pe_1_4_7_N74), .B2(
        npu_inst_pe_1_4_7_n76), .C1(npu_inst_pe_1_4_7_N66), .C2(
        npu_inst_pe_1_4_7_n77), .ZN(npu_inst_pe_1_4_7_n83) );
  INV_X1 npu_inst_pe_1_4_7_U70 ( .A(npu_inst_pe_1_4_7_n83), .ZN(
        npu_inst_pe_1_4_7_n100) );
  AOI222_X1 npu_inst_pe_1_4_7_U69 ( .A1(npu_inst_int_data_res_5__7__2_), .A2(
        npu_inst_pe_1_4_7_n1), .B1(npu_inst_pe_1_4_7_N75), .B2(
        npu_inst_pe_1_4_7_n76), .C1(npu_inst_pe_1_4_7_N67), .C2(
        npu_inst_pe_1_4_7_n77), .ZN(npu_inst_pe_1_4_7_n82) );
  INV_X1 npu_inst_pe_1_4_7_U68 ( .A(npu_inst_pe_1_4_7_n82), .ZN(
        npu_inst_pe_1_4_7_n99) );
  AOI222_X1 npu_inst_pe_1_4_7_U67 ( .A1(npu_inst_int_data_res_5__7__3_), .A2(
        npu_inst_pe_1_4_7_n1), .B1(npu_inst_pe_1_4_7_N76), .B2(
        npu_inst_pe_1_4_7_n76), .C1(npu_inst_pe_1_4_7_N68), .C2(
        npu_inst_pe_1_4_7_n77), .ZN(npu_inst_pe_1_4_7_n81) );
  INV_X1 npu_inst_pe_1_4_7_U66 ( .A(npu_inst_pe_1_4_7_n81), .ZN(
        npu_inst_pe_1_4_7_n98) );
  AOI222_X1 npu_inst_pe_1_4_7_U65 ( .A1(npu_inst_int_data_res_5__7__4_), .A2(
        npu_inst_pe_1_4_7_n1), .B1(npu_inst_pe_1_4_7_N77), .B2(
        npu_inst_pe_1_4_7_n76), .C1(npu_inst_pe_1_4_7_N69), .C2(
        npu_inst_pe_1_4_7_n77), .ZN(npu_inst_pe_1_4_7_n80) );
  INV_X1 npu_inst_pe_1_4_7_U64 ( .A(npu_inst_pe_1_4_7_n80), .ZN(
        npu_inst_pe_1_4_7_n36) );
  AOI222_X1 npu_inst_pe_1_4_7_U63 ( .A1(npu_inst_int_data_res_5__7__5_), .A2(
        npu_inst_pe_1_4_7_n1), .B1(npu_inst_pe_1_4_7_N78), .B2(
        npu_inst_pe_1_4_7_n76), .C1(npu_inst_pe_1_4_7_N70), .C2(
        npu_inst_pe_1_4_7_n77), .ZN(npu_inst_pe_1_4_7_n79) );
  INV_X1 npu_inst_pe_1_4_7_U62 ( .A(npu_inst_pe_1_4_7_n79), .ZN(
        npu_inst_pe_1_4_7_n35) );
  AOI222_X1 npu_inst_pe_1_4_7_U61 ( .A1(npu_inst_int_data_res_5__7__6_), .A2(
        npu_inst_pe_1_4_7_n1), .B1(npu_inst_pe_1_4_7_N79), .B2(
        npu_inst_pe_1_4_7_n76), .C1(npu_inst_pe_1_4_7_N71), .C2(
        npu_inst_pe_1_4_7_n77), .ZN(npu_inst_pe_1_4_7_n78) );
  INV_X1 npu_inst_pe_1_4_7_U60 ( .A(npu_inst_pe_1_4_7_n78), .ZN(
        npu_inst_pe_1_4_7_n34) );
  INV_X1 npu_inst_pe_1_4_7_U59 ( .A(npu_inst_pe_1_4_7_int_data_1_), .ZN(
        npu_inst_pe_1_4_7_n14) );
  AND2_X1 npu_inst_pe_1_4_7_U58 ( .A1(npu_inst_int_data_x_4__7__1_), .A2(
        npu_inst_pe_1_4_7_int_q_weight_1_), .ZN(npu_inst_pe_1_4_7_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_4_7_U57 ( .A1(npu_inst_int_data_x_4__7__0_), .A2(
        npu_inst_pe_1_4_7_int_q_weight_1_), .ZN(npu_inst_pe_1_4_7_int_data_0_)
         );
  NAND2_X1 npu_inst_pe_1_4_7_U56 ( .A1(npu_inst_pe_1_4_7_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_4_7_n60), .ZN(npu_inst_pe_1_4_7_n74) );
  OAI21_X1 npu_inst_pe_1_4_7_U55 ( .B1(npu_inst_pe_1_4_7_n63), .B2(
        npu_inst_pe_1_4_7_n60), .A(npu_inst_pe_1_4_7_n74), .ZN(
        npu_inst_pe_1_4_7_n97) );
  NAND2_X1 npu_inst_pe_1_4_7_U54 ( .A1(npu_inst_pe_1_4_7_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_4_7_n60), .ZN(npu_inst_pe_1_4_7_n73) );
  OAI21_X1 npu_inst_pe_1_4_7_U53 ( .B1(npu_inst_pe_1_4_7_n61), .B2(
        npu_inst_pe_1_4_7_n60), .A(npu_inst_pe_1_4_7_n73), .ZN(
        npu_inst_pe_1_4_7_n96) );
  NAND2_X1 npu_inst_pe_1_4_7_U52 ( .A1(npu_inst_pe_1_4_7_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_4_7_n56), .ZN(npu_inst_pe_1_4_7_n72) );
  OAI21_X1 npu_inst_pe_1_4_7_U51 ( .B1(npu_inst_pe_1_4_7_n63), .B2(
        npu_inst_pe_1_4_7_n56), .A(npu_inst_pe_1_4_7_n72), .ZN(
        npu_inst_pe_1_4_7_n95) );
  NAND2_X1 npu_inst_pe_1_4_7_U50 ( .A1(npu_inst_pe_1_4_7_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_4_7_n56), .ZN(npu_inst_pe_1_4_7_n71) );
  OAI21_X1 npu_inst_pe_1_4_7_U49 ( .B1(npu_inst_pe_1_4_7_n61), .B2(
        npu_inst_pe_1_4_7_n56), .A(npu_inst_pe_1_4_7_n71), .ZN(
        npu_inst_pe_1_4_7_n94) );
  NAND2_X1 npu_inst_pe_1_4_7_U48 ( .A1(npu_inst_pe_1_4_7_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_4_7_n52), .ZN(npu_inst_pe_1_4_7_n70) );
  OAI21_X1 npu_inst_pe_1_4_7_U47 ( .B1(npu_inst_pe_1_4_7_n63), .B2(
        npu_inst_pe_1_4_7_n52), .A(npu_inst_pe_1_4_7_n70), .ZN(
        npu_inst_pe_1_4_7_n93) );
  NAND2_X1 npu_inst_pe_1_4_7_U46 ( .A1(npu_inst_pe_1_4_7_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_4_7_n52), .ZN(npu_inst_pe_1_4_7_n69) );
  OAI21_X1 npu_inst_pe_1_4_7_U45 ( .B1(npu_inst_pe_1_4_7_n61), .B2(
        npu_inst_pe_1_4_7_n52), .A(npu_inst_pe_1_4_7_n69), .ZN(
        npu_inst_pe_1_4_7_n92) );
  NAND2_X1 npu_inst_pe_1_4_7_U44 ( .A1(npu_inst_pe_1_4_7_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_4_7_n48), .ZN(npu_inst_pe_1_4_7_n68) );
  OAI21_X1 npu_inst_pe_1_4_7_U43 ( .B1(npu_inst_pe_1_4_7_n63), .B2(
        npu_inst_pe_1_4_7_n48), .A(npu_inst_pe_1_4_7_n68), .ZN(
        npu_inst_pe_1_4_7_n91) );
  NAND2_X1 npu_inst_pe_1_4_7_U42 ( .A1(npu_inst_pe_1_4_7_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_4_7_n48), .ZN(npu_inst_pe_1_4_7_n67) );
  OAI21_X1 npu_inst_pe_1_4_7_U41 ( .B1(npu_inst_pe_1_4_7_n61), .B2(
        npu_inst_pe_1_4_7_n48), .A(npu_inst_pe_1_4_7_n67), .ZN(
        npu_inst_pe_1_4_7_n90) );
  NAND2_X1 npu_inst_pe_1_4_7_U40 ( .A1(npu_inst_pe_1_4_7_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_4_7_n44), .ZN(npu_inst_pe_1_4_7_n66) );
  OAI21_X1 npu_inst_pe_1_4_7_U39 ( .B1(npu_inst_pe_1_4_7_n63), .B2(
        npu_inst_pe_1_4_7_n44), .A(npu_inst_pe_1_4_7_n66), .ZN(
        npu_inst_pe_1_4_7_n89) );
  NAND2_X1 npu_inst_pe_1_4_7_U38 ( .A1(npu_inst_pe_1_4_7_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_4_7_n44), .ZN(npu_inst_pe_1_4_7_n65) );
  OAI21_X1 npu_inst_pe_1_4_7_U37 ( .B1(npu_inst_pe_1_4_7_n61), .B2(
        npu_inst_pe_1_4_7_n44), .A(npu_inst_pe_1_4_7_n65), .ZN(
        npu_inst_pe_1_4_7_n88) );
  NAND2_X1 npu_inst_pe_1_4_7_U36 ( .A1(npu_inst_pe_1_4_7_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_4_7_n40), .ZN(npu_inst_pe_1_4_7_n64) );
  OAI21_X1 npu_inst_pe_1_4_7_U35 ( .B1(npu_inst_pe_1_4_7_n63), .B2(
        npu_inst_pe_1_4_7_n40), .A(npu_inst_pe_1_4_7_n64), .ZN(
        npu_inst_pe_1_4_7_n87) );
  NAND2_X1 npu_inst_pe_1_4_7_U34 ( .A1(npu_inst_pe_1_4_7_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_4_7_n40), .ZN(npu_inst_pe_1_4_7_n62) );
  OAI21_X1 npu_inst_pe_1_4_7_U33 ( .B1(npu_inst_pe_1_4_7_n61), .B2(
        npu_inst_pe_1_4_7_n40), .A(npu_inst_pe_1_4_7_n62), .ZN(
        npu_inst_pe_1_4_7_n86) );
  INV_X1 npu_inst_pe_1_4_7_U32 ( .A(npu_inst_pe_1_4_7_int_data_0_), .ZN(
        npu_inst_pe_1_4_7_n13) );
  INV_X1 npu_inst_pe_1_4_7_U31 ( .A(npu_inst_n69), .ZN(npu_inst_pe_1_4_7_n5)
         );
  AOI22_X1 npu_inst_pe_1_4_7_U30 ( .A1(npu_inst_n55), .A2(
        npu_inst_int_data_y_5__7__1_), .B1(npu_inst_pe_1_4_7_n3), .B2(
        int_i_data_h_npu5[1]), .ZN(npu_inst_pe_1_4_7_n63) );
  AOI22_X1 npu_inst_pe_1_4_7_U29 ( .A1(npu_inst_n55), .A2(
        npu_inst_int_data_y_5__7__0_), .B1(npu_inst_pe_1_4_7_n3), .B2(
        int_i_data_h_npu5[0]), .ZN(npu_inst_pe_1_4_7_n61) );
  OR3_X1 npu_inst_pe_1_4_7_U28 ( .A1(npu_inst_pe_1_4_7_n6), .A2(
        npu_inst_pe_1_4_7_n8), .A3(npu_inst_pe_1_4_7_n5), .ZN(
        npu_inst_pe_1_4_7_n56) );
  OR3_X1 npu_inst_pe_1_4_7_U27 ( .A1(npu_inst_pe_1_4_7_n5), .A2(
        npu_inst_pe_1_4_7_n8), .A3(npu_inst_pe_1_4_7_n7), .ZN(
        npu_inst_pe_1_4_7_n48) );
  INV_X1 npu_inst_pe_1_4_7_U26 ( .A(npu_inst_pe_1_4_7_n5), .ZN(
        npu_inst_pe_1_4_7_n4) );
  INV_X1 npu_inst_pe_1_4_7_U25 ( .A(npu_inst_n124), .ZN(npu_inst_pe_1_4_7_n12)
         );
  OR3_X1 npu_inst_pe_1_4_7_U24 ( .A1(npu_inst_pe_1_4_7_n4), .A2(
        npu_inst_pe_1_4_7_n8), .A3(npu_inst_pe_1_4_7_n7), .ZN(
        npu_inst_pe_1_4_7_n52) );
  OR3_X1 npu_inst_pe_1_4_7_U23 ( .A1(npu_inst_pe_1_4_7_n6), .A2(
        npu_inst_pe_1_4_7_n8), .A3(npu_inst_pe_1_4_7_n4), .ZN(
        npu_inst_pe_1_4_7_n60) );
  NOR2_X1 npu_inst_pe_1_4_7_U22 ( .A1(npu_inst_pe_1_4_7_n60), .A2(
        npu_inst_pe_1_4_7_n3), .ZN(npu_inst_pe_1_4_7_n58) );
  NOR2_X1 npu_inst_pe_1_4_7_U21 ( .A1(npu_inst_pe_1_4_7_n56), .A2(
        npu_inst_pe_1_4_7_n3), .ZN(npu_inst_pe_1_4_7_n54) );
  NOR2_X1 npu_inst_pe_1_4_7_U20 ( .A1(npu_inst_pe_1_4_7_n52), .A2(
        npu_inst_pe_1_4_7_n3), .ZN(npu_inst_pe_1_4_7_n50) );
  NOR2_X1 npu_inst_pe_1_4_7_U19 ( .A1(npu_inst_pe_1_4_7_n48), .A2(
        npu_inst_pe_1_4_7_n3), .ZN(npu_inst_pe_1_4_7_n46) );
  NOR2_X1 npu_inst_pe_1_4_7_U18 ( .A1(npu_inst_pe_1_4_7_n40), .A2(
        npu_inst_pe_1_4_7_n3), .ZN(npu_inst_pe_1_4_7_n38) );
  NOR2_X1 npu_inst_pe_1_4_7_U17 ( .A1(npu_inst_pe_1_4_7_n44), .A2(
        npu_inst_pe_1_4_7_n3), .ZN(npu_inst_pe_1_4_7_n42) );
  BUF_X1 npu_inst_pe_1_4_7_U16 ( .A(npu_inst_n98), .Z(npu_inst_pe_1_4_7_n8) );
  BUF_X1 npu_inst_pe_1_4_7_U15 ( .A(npu_inst_pe_1_4_7_n12), .Z(
        npu_inst_pe_1_4_7_n11) );
  BUF_X1 npu_inst_pe_1_4_7_U14 ( .A(npu_inst_pe_1_4_7_n12), .Z(
        npu_inst_pe_1_4_7_n10) );
  BUF_X1 npu_inst_pe_1_4_7_U13 ( .A(npu_inst_pe_1_4_7_n12), .Z(
        npu_inst_pe_1_4_7_n9) );
  INV_X1 npu_inst_pe_1_4_7_U12 ( .A(npu_inst_pe_1_4_7_n38), .ZN(
        npu_inst_pe_1_4_7_n118) );
  INV_X1 npu_inst_pe_1_4_7_U11 ( .A(npu_inst_pe_1_4_7_n58), .ZN(
        npu_inst_pe_1_4_7_n114) );
  INV_X1 npu_inst_pe_1_4_7_U10 ( .A(npu_inst_pe_1_4_7_n54), .ZN(
        npu_inst_pe_1_4_7_n115) );
  INV_X1 npu_inst_pe_1_4_7_U9 ( .A(npu_inst_pe_1_4_7_n50), .ZN(
        npu_inst_pe_1_4_7_n116) );
  INV_X1 npu_inst_pe_1_4_7_U8 ( .A(npu_inst_pe_1_4_7_n46), .ZN(
        npu_inst_pe_1_4_7_n117) );
  INV_X1 npu_inst_pe_1_4_7_U7 ( .A(npu_inst_pe_1_4_7_n42), .ZN(
        npu_inst_pe_1_4_7_n119) );
  BUF_X1 npu_inst_pe_1_4_7_U6 ( .A(npu_inst_n19), .Z(npu_inst_pe_1_4_7_n2) );
  BUF_X1 npu_inst_pe_1_4_7_U5 ( .A(npu_inst_n19), .Z(npu_inst_pe_1_4_7_n1) );
  NOR2_X1 npu_inst_pe_1_4_7_U4 ( .A1(npu_inst_pe_1_4_7_int_q_weight_0_), .A2(
        npu_inst_pe_1_4_7_n1), .ZN(npu_inst_pe_1_4_7_n76) );
  NOR2_X1 npu_inst_pe_1_4_7_U3 ( .A1(npu_inst_pe_1_4_7_n27), .A2(
        npu_inst_pe_1_4_7_n1), .ZN(npu_inst_pe_1_4_7_n77) );
  FA_X1 npu_inst_pe_1_4_7_sub_77_U2_1 ( .A(npu_inst_pe_1_4_7_int_q_acc_1_), 
        .B(npu_inst_pe_1_4_7_n14), .CI(npu_inst_pe_1_4_7_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_4_7_sub_77_carry_2_), .S(npu_inst_pe_1_4_7_N66) );
  FA_X1 npu_inst_pe_1_4_7_add_79_U1_1 ( .A(npu_inst_pe_1_4_7_int_q_acc_1_), 
        .B(npu_inst_pe_1_4_7_int_data_1_), .CI(
        npu_inst_pe_1_4_7_add_79_carry_1_), .CO(
        npu_inst_pe_1_4_7_add_79_carry_2_), .S(npu_inst_pe_1_4_7_N74) );
  NAND3_X1 npu_inst_pe_1_4_7_U109 ( .A1(npu_inst_pe_1_4_7_n5), .A2(
        npu_inst_pe_1_4_7_n7), .A3(npu_inst_pe_1_4_7_n8), .ZN(
        npu_inst_pe_1_4_7_n44) );
  NAND3_X1 npu_inst_pe_1_4_7_U108 ( .A1(npu_inst_pe_1_4_7_n4), .A2(
        npu_inst_pe_1_4_7_n7), .A3(npu_inst_pe_1_4_7_n8), .ZN(
        npu_inst_pe_1_4_7_n40) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_4_7_n34), .CK(
        npu_inst_pe_1_4_7_net3396), .RN(npu_inst_pe_1_4_7_n9), .Q(
        npu_inst_pe_1_4_7_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_4_7_n35), .CK(
        npu_inst_pe_1_4_7_net3396), .RN(npu_inst_pe_1_4_7_n9), .Q(
        npu_inst_pe_1_4_7_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_4_7_n36), .CK(
        npu_inst_pe_1_4_7_net3396), .RN(npu_inst_pe_1_4_7_n9), .Q(
        npu_inst_pe_1_4_7_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_4_7_n98), .CK(
        npu_inst_pe_1_4_7_net3396), .RN(npu_inst_pe_1_4_7_n9), .Q(
        npu_inst_pe_1_4_7_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_4_7_n99), .CK(
        npu_inst_pe_1_4_7_net3396), .RN(npu_inst_pe_1_4_7_n9), .Q(
        npu_inst_pe_1_4_7_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_4_7_n100), 
        .CK(npu_inst_pe_1_4_7_net3396), .RN(npu_inst_pe_1_4_7_n9), .Q(
        npu_inst_pe_1_4_7_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_4_7_n33), .CK(
        npu_inst_pe_1_4_7_net3396), .RN(npu_inst_pe_1_4_7_n9), .Q(
        npu_inst_pe_1_4_7_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_4_7_n101), 
        .CK(npu_inst_pe_1_4_7_net3396), .RN(npu_inst_pe_1_4_7_n9), .Q(
        npu_inst_pe_1_4_7_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_weight_reg_0_ ( .D(npu_inst_n110), .CK(
        npu_inst_pe_1_4_7_net3402), .RN(npu_inst_pe_1_4_7_n9), .Q(
        npu_inst_pe_1_4_7_int_q_weight_0_), .QN(npu_inst_pe_1_4_7_n27) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_weight_reg_1_ ( .D(npu_inst_n116), .CK(
        npu_inst_pe_1_4_7_net3402), .RN(npu_inst_pe_1_4_7_n9), .Q(
        npu_inst_pe_1_4_7_int_q_weight_1_), .QN(npu_inst_pe_1_4_7_n26) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_4_7_n113), 
        .CK(npu_inst_pe_1_4_7_net3402), .RN(npu_inst_pe_1_4_7_n9), .Q(
        npu_inst_pe_1_4_7_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_4_7_n107), 
        .CK(npu_inst_pe_1_4_7_net3402), .RN(npu_inst_pe_1_4_7_n9), .Q(
        npu_inst_pe_1_4_7_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_4_7_n112), 
        .CK(npu_inst_pe_1_4_7_net3402), .RN(npu_inst_pe_1_4_7_n10), .Q(
        npu_inst_pe_1_4_7_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_4_7_n106), 
        .CK(npu_inst_pe_1_4_7_net3402), .RN(npu_inst_pe_1_4_7_n10), .Q(
        npu_inst_pe_1_4_7_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_4_7_n111), 
        .CK(npu_inst_pe_1_4_7_net3402), .RN(npu_inst_pe_1_4_7_n10), .Q(
        npu_inst_pe_1_4_7_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_4_7_n105), 
        .CK(npu_inst_pe_1_4_7_net3402), .RN(npu_inst_pe_1_4_7_n10), .Q(
        npu_inst_pe_1_4_7_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_4_7_n110), 
        .CK(npu_inst_pe_1_4_7_net3402), .RN(npu_inst_pe_1_4_7_n10), .Q(
        npu_inst_pe_1_4_7_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_4_7_n104), 
        .CK(npu_inst_pe_1_4_7_net3402), .RN(npu_inst_pe_1_4_7_n10), .Q(
        npu_inst_pe_1_4_7_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_4_7_n109), 
        .CK(npu_inst_pe_1_4_7_net3402), .RN(npu_inst_pe_1_4_7_n10), .Q(
        npu_inst_pe_1_4_7_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_4_7_n103), 
        .CK(npu_inst_pe_1_4_7_net3402), .RN(npu_inst_pe_1_4_7_n10), .Q(
        npu_inst_pe_1_4_7_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_4_7_n108), 
        .CK(npu_inst_pe_1_4_7_net3402), .RN(npu_inst_pe_1_4_7_n10), .Q(
        npu_inst_pe_1_4_7_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_4_7_n102), 
        .CK(npu_inst_pe_1_4_7_net3402), .RN(npu_inst_pe_1_4_7_n10), .Q(
        npu_inst_pe_1_4_7_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_4_7_n86), 
        .CK(npu_inst_pe_1_4_7_net3402), .RN(npu_inst_pe_1_4_7_n10), .Q(
        npu_inst_pe_1_4_7_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_4_7_n87), 
        .CK(npu_inst_pe_1_4_7_net3402), .RN(npu_inst_pe_1_4_7_n10), .Q(
        npu_inst_pe_1_4_7_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_4_7_n88), 
        .CK(npu_inst_pe_1_4_7_net3402), .RN(npu_inst_pe_1_4_7_n11), .Q(
        npu_inst_pe_1_4_7_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_4_7_n89), 
        .CK(npu_inst_pe_1_4_7_net3402), .RN(npu_inst_pe_1_4_7_n11), .Q(
        npu_inst_pe_1_4_7_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_4_7_n90), 
        .CK(npu_inst_pe_1_4_7_net3402), .RN(npu_inst_pe_1_4_7_n11), .Q(
        npu_inst_pe_1_4_7_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_4_7_n91), 
        .CK(npu_inst_pe_1_4_7_net3402), .RN(npu_inst_pe_1_4_7_n11), .Q(
        npu_inst_pe_1_4_7_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_4_7_n92), 
        .CK(npu_inst_pe_1_4_7_net3402), .RN(npu_inst_pe_1_4_7_n11), .Q(
        npu_inst_pe_1_4_7_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_4_7_n93), 
        .CK(npu_inst_pe_1_4_7_net3402), .RN(npu_inst_pe_1_4_7_n11), .Q(
        npu_inst_pe_1_4_7_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_4_7_n94), 
        .CK(npu_inst_pe_1_4_7_net3402), .RN(npu_inst_pe_1_4_7_n11), .Q(
        npu_inst_pe_1_4_7_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_4_7_n95), 
        .CK(npu_inst_pe_1_4_7_net3402), .RN(npu_inst_pe_1_4_7_n11), .Q(
        npu_inst_pe_1_4_7_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_4_7_n96), 
        .CK(npu_inst_pe_1_4_7_net3402), .RN(npu_inst_pe_1_4_7_n11), .Q(
        npu_inst_pe_1_4_7_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_4_7_n97), 
        .CK(npu_inst_pe_1_4_7_net3402), .RN(npu_inst_pe_1_4_7_n11), .Q(
        npu_inst_pe_1_4_7_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_4_7_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_4_7_N84), .SE(1'b0), .GCK(npu_inst_pe_1_4_7_net3396) );
  CLKGATETST_X1 npu_inst_pe_1_4_7_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n63), .SE(1'b0), .GCK(npu_inst_pe_1_4_7_net3402) );
  MUX2_X1 npu_inst_pe_1_5_0_U161 ( .A(npu_inst_pe_1_5_0_n31), .B(
        npu_inst_pe_1_5_0_n28), .S(npu_inst_pe_1_5_0_n7), .Z(
        npu_inst_pe_1_5_0_N93) );
  MUX2_X1 npu_inst_pe_1_5_0_U160 ( .A(npu_inst_pe_1_5_0_n30), .B(
        npu_inst_pe_1_5_0_n29), .S(npu_inst_n76), .Z(npu_inst_pe_1_5_0_n31) );
  MUX2_X1 npu_inst_pe_1_5_0_U159 ( .A(npu_inst_pe_1_5_0_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_5_0_int_q_reg_v_1__0_), .S(npu_inst_pe_1_5_0_n4), .Z(
        npu_inst_pe_1_5_0_n30) );
  MUX2_X1 npu_inst_pe_1_5_0_U158 ( .A(npu_inst_pe_1_5_0_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_5_0_int_q_reg_v_3__0_), .S(npu_inst_pe_1_5_0_n4), .Z(
        npu_inst_pe_1_5_0_n29) );
  MUX2_X1 npu_inst_pe_1_5_0_U157 ( .A(npu_inst_pe_1_5_0_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_5_0_int_q_reg_v_5__0_), .S(npu_inst_pe_1_5_0_n4), .Z(
        npu_inst_pe_1_5_0_n28) );
  MUX2_X1 npu_inst_pe_1_5_0_U156 ( .A(npu_inst_pe_1_5_0_n25), .B(
        npu_inst_pe_1_5_0_n22), .S(npu_inst_pe_1_5_0_n7), .Z(
        npu_inst_pe_1_5_0_N94) );
  MUX2_X1 npu_inst_pe_1_5_0_U155 ( .A(npu_inst_pe_1_5_0_n24), .B(
        npu_inst_pe_1_5_0_n23), .S(npu_inst_n76), .Z(npu_inst_pe_1_5_0_n25) );
  MUX2_X1 npu_inst_pe_1_5_0_U154 ( .A(npu_inst_pe_1_5_0_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_5_0_int_q_reg_v_1__1_), .S(npu_inst_pe_1_5_0_n4), .Z(
        npu_inst_pe_1_5_0_n24) );
  MUX2_X1 npu_inst_pe_1_5_0_U153 ( .A(npu_inst_pe_1_5_0_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_5_0_int_q_reg_v_3__1_), .S(npu_inst_pe_1_5_0_n4), .Z(
        npu_inst_pe_1_5_0_n23) );
  MUX2_X1 npu_inst_pe_1_5_0_U152 ( .A(npu_inst_pe_1_5_0_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_5_0_int_q_reg_v_5__1_), .S(npu_inst_pe_1_5_0_n4), .Z(
        npu_inst_pe_1_5_0_n22) );
  MUX2_X1 npu_inst_pe_1_5_0_U151 ( .A(npu_inst_pe_1_5_0_n21), .B(
        npu_inst_pe_1_5_0_n18), .S(npu_inst_pe_1_5_0_n7), .Z(
        npu_inst_pe_1_5_0_o_data_h_1_) );
  MUX2_X1 npu_inst_pe_1_5_0_U150 ( .A(npu_inst_pe_1_5_0_n20), .B(
        npu_inst_pe_1_5_0_n19), .S(npu_inst_n76), .Z(npu_inst_pe_1_5_0_n21) );
  MUX2_X1 npu_inst_pe_1_5_0_U149 ( .A(npu_inst_pe_1_5_0_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_5_0_int_q_reg_h_1__1_), .S(npu_inst_pe_1_5_0_n4), .Z(
        npu_inst_pe_1_5_0_n20) );
  MUX2_X1 npu_inst_pe_1_5_0_U148 ( .A(npu_inst_pe_1_5_0_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_5_0_int_q_reg_h_3__1_), .S(npu_inst_pe_1_5_0_n4), .Z(
        npu_inst_pe_1_5_0_n19) );
  MUX2_X1 npu_inst_pe_1_5_0_U147 ( .A(npu_inst_pe_1_5_0_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_5_0_int_q_reg_h_5__1_), .S(npu_inst_pe_1_5_0_n4), .Z(
        npu_inst_pe_1_5_0_n18) );
  MUX2_X1 npu_inst_pe_1_5_0_U146 ( .A(npu_inst_pe_1_5_0_n17), .B(
        npu_inst_pe_1_5_0_n14), .S(npu_inst_pe_1_5_0_n7), .Z(
        npu_inst_pe_1_5_0_o_data_h_0_) );
  MUX2_X1 npu_inst_pe_1_5_0_U145 ( .A(npu_inst_pe_1_5_0_n16), .B(
        npu_inst_pe_1_5_0_n15), .S(npu_inst_n76), .Z(npu_inst_pe_1_5_0_n17) );
  MUX2_X1 npu_inst_pe_1_5_0_U144 ( .A(npu_inst_pe_1_5_0_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_5_0_int_q_reg_h_1__0_), .S(npu_inst_pe_1_5_0_n4), .Z(
        npu_inst_pe_1_5_0_n16) );
  MUX2_X1 npu_inst_pe_1_5_0_U143 ( .A(npu_inst_pe_1_5_0_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_5_0_int_q_reg_h_3__0_), .S(npu_inst_pe_1_5_0_n4), .Z(
        npu_inst_pe_1_5_0_n15) );
  MUX2_X1 npu_inst_pe_1_5_0_U142 ( .A(npu_inst_pe_1_5_0_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_5_0_int_q_reg_h_5__0_), .S(npu_inst_pe_1_5_0_n4), .Z(
        npu_inst_pe_1_5_0_n14) );
  XOR2_X1 npu_inst_pe_1_5_0_U141 ( .A(npu_inst_pe_1_5_0_int_data_0_), .B(
        npu_inst_pe_1_5_0_int_q_acc_0_), .Z(npu_inst_pe_1_5_0_N73) );
  AND2_X1 npu_inst_pe_1_5_0_U140 ( .A1(npu_inst_pe_1_5_0_int_q_acc_0_), .A2(
        npu_inst_pe_1_5_0_int_data_0_), .ZN(npu_inst_pe_1_5_0_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_5_0_U139 ( .A(npu_inst_pe_1_5_0_int_q_acc_0_), .B(
        npu_inst_pe_1_5_0_n12), .ZN(npu_inst_pe_1_5_0_N65) );
  OR2_X1 npu_inst_pe_1_5_0_U138 ( .A1(npu_inst_pe_1_5_0_n12), .A2(
        npu_inst_pe_1_5_0_int_q_acc_0_), .ZN(npu_inst_pe_1_5_0_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_5_0_U137 ( .A(npu_inst_pe_1_5_0_int_q_acc_2_), .B(
        npu_inst_pe_1_5_0_add_79_carry_2_), .Z(npu_inst_pe_1_5_0_N75) );
  AND2_X1 npu_inst_pe_1_5_0_U136 ( .A1(npu_inst_pe_1_5_0_add_79_carry_2_), 
        .A2(npu_inst_pe_1_5_0_int_q_acc_2_), .ZN(
        npu_inst_pe_1_5_0_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_5_0_U135 ( .A(npu_inst_pe_1_5_0_int_q_acc_3_), .B(
        npu_inst_pe_1_5_0_add_79_carry_3_), .Z(npu_inst_pe_1_5_0_N76) );
  AND2_X1 npu_inst_pe_1_5_0_U134 ( .A1(npu_inst_pe_1_5_0_add_79_carry_3_), 
        .A2(npu_inst_pe_1_5_0_int_q_acc_3_), .ZN(
        npu_inst_pe_1_5_0_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_5_0_U133 ( .A(npu_inst_pe_1_5_0_int_q_acc_4_), .B(
        npu_inst_pe_1_5_0_add_79_carry_4_), .Z(npu_inst_pe_1_5_0_N77) );
  AND2_X1 npu_inst_pe_1_5_0_U132 ( .A1(npu_inst_pe_1_5_0_add_79_carry_4_), 
        .A2(npu_inst_pe_1_5_0_int_q_acc_4_), .ZN(
        npu_inst_pe_1_5_0_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_5_0_U131 ( .A(npu_inst_pe_1_5_0_int_q_acc_5_), .B(
        npu_inst_pe_1_5_0_add_79_carry_5_), .Z(npu_inst_pe_1_5_0_N78) );
  AND2_X1 npu_inst_pe_1_5_0_U130 ( .A1(npu_inst_pe_1_5_0_add_79_carry_5_), 
        .A2(npu_inst_pe_1_5_0_int_q_acc_5_), .ZN(
        npu_inst_pe_1_5_0_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_5_0_U129 ( .A(npu_inst_pe_1_5_0_int_q_acc_6_), .B(
        npu_inst_pe_1_5_0_add_79_carry_6_), .Z(npu_inst_pe_1_5_0_N79) );
  AND2_X1 npu_inst_pe_1_5_0_U128 ( .A1(npu_inst_pe_1_5_0_add_79_carry_6_), 
        .A2(npu_inst_pe_1_5_0_int_q_acc_6_), .ZN(
        npu_inst_pe_1_5_0_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_5_0_U127 ( .A(npu_inst_pe_1_5_0_int_q_acc_7_), .B(
        npu_inst_pe_1_5_0_add_79_carry_7_), .Z(npu_inst_pe_1_5_0_N80) );
  XNOR2_X1 npu_inst_pe_1_5_0_U126 ( .A(npu_inst_pe_1_5_0_sub_77_carry_2_), .B(
        npu_inst_pe_1_5_0_int_q_acc_2_), .ZN(npu_inst_pe_1_5_0_N67) );
  OR2_X1 npu_inst_pe_1_5_0_U125 ( .A1(npu_inst_pe_1_5_0_int_q_acc_2_), .A2(
        npu_inst_pe_1_5_0_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_5_0_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_5_0_U124 ( .A(npu_inst_pe_1_5_0_sub_77_carry_3_), .B(
        npu_inst_pe_1_5_0_int_q_acc_3_), .ZN(npu_inst_pe_1_5_0_N68) );
  OR2_X1 npu_inst_pe_1_5_0_U123 ( .A1(npu_inst_pe_1_5_0_int_q_acc_3_), .A2(
        npu_inst_pe_1_5_0_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_5_0_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_5_0_U122 ( .A(npu_inst_pe_1_5_0_sub_77_carry_4_), .B(
        npu_inst_pe_1_5_0_int_q_acc_4_), .ZN(npu_inst_pe_1_5_0_N69) );
  OR2_X1 npu_inst_pe_1_5_0_U121 ( .A1(npu_inst_pe_1_5_0_int_q_acc_4_), .A2(
        npu_inst_pe_1_5_0_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_5_0_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_5_0_U120 ( .A(npu_inst_pe_1_5_0_sub_77_carry_5_), .B(
        npu_inst_pe_1_5_0_int_q_acc_5_), .ZN(npu_inst_pe_1_5_0_N70) );
  OR2_X1 npu_inst_pe_1_5_0_U119 ( .A1(npu_inst_pe_1_5_0_int_q_acc_5_), .A2(
        npu_inst_pe_1_5_0_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_5_0_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_5_0_U118 ( .A(npu_inst_pe_1_5_0_sub_77_carry_6_), .B(
        npu_inst_pe_1_5_0_int_q_acc_6_), .ZN(npu_inst_pe_1_5_0_N71) );
  OR2_X1 npu_inst_pe_1_5_0_U117 ( .A1(npu_inst_pe_1_5_0_int_q_acc_6_), .A2(
        npu_inst_pe_1_5_0_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_5_0_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_5_0_U116 ( .A(npu_inst_pe_1_5_0_int_q_acc_7_), .B(
        npu_inst_pe_1_5_0_sub_77_carry_7_), .ZN(npu_inst_pe_1_5_0_N72) );
  INV_X1 npu_inst_pe_1_5_0_U115 ( .A(npu_inst_n76), .ZN(npu_inst_pe_1_5_0_n6)
         );
  INV_X1 npu_inst_pe_1_5_0_U114 ( .A(npu_inst_n55), .ZN(npu_inst_pe_1_5_0_n3)
         );
  AOI22_X1 npu_inst_pe_1_5_0_U113 ( .A1(npu_inst_int_data_y_6__0__0_), .A2(
        npu_inst_pe_1_5_0_n58), .B1(npu_inst_pe_1_5_0_n113), .B2(
        npu_inst_pe_1_5_0_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_5_0_n57) );
  INV_X1 npu_inst_pe_1_5_0_U112 ( .A(npu_inst_pe_1_5_0_n57), .ZN(
        npu_inst_pe_1_5_0_n107) );
  AOI22_X1 npu_inst_pe_1_5_0_U111 ( .A1(npu_inst_int_data_y_6__0__0_), .A2(
        npu_inst_pe_1_5_0_n54), .B1(npu_inst_pe_1_5_0_n114), .B2(
        npu_inst_pe_1_5_0_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_5_0_n53) );
  INV_X1 npu_inst_pe_1_5_0_U110 ( .A(npu_inst_pe_1_5_0_n53), .ZN(
        npu_inst_pe_1_5_0_n108) );
  AOI22_X1 npu_inst_pe_1_5_0_U107 ( .A1(npu_inst_int_data_y_6__0__0_), .A2(
        npu_inst_pe_1_5_0_n50), .B1(npu_inst_pe_1_5_0_n115), .B2(
        npu_inst_pe_1_5_0_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_5_0_n49) );
  INV_X1 npu_inst_pe_1_5_0_U106 ( .A(npu_inst_pe_1_5_0_n49), .ZN(
        npu_inst_pe_1_5_0_n109) );
  AOI22_X1 npu_inst_pe_1_5_0_U105 ( .A1(npu_inst_int_data_y_6__0__0_), .A2(
        npu_inst_pe_1_5_0_n46), .B1(npu_inst_pe_1_5_0_n116), .B2(
        npu_inst_pe_1_5_0_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_5_0_n45) );
  INV_X1 npu_inst_pe_1_5_0_U104 ( .A(npu_inst_pe_1_5_0_n45), .ZN(
        npu_inst_pe_1_5_0_n110) );
  AOI22_X1 npu_inst_pe_1_5_0_U103 ( .A1(npu_inst_int_data_y_6__0__0_), .A2(
        npu_inst_pe_1_5_0_n42), .B1(npu_inst_pe_1_5_0_n118), .B2(
        npu_inst_pe_1_5_0_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_5_0_n41) );
  INV_X1 npu_inst_pe_1_5_0_U102 ( .A(npu_inst_pe_1_5_0_n41), .ZN(
        npu_inst_pe_1_5_0_n111) );
  AOI22_X1 npu_inst_pe_1_5_0_U101 ( .A1(npu_inst_int_data_y_6__0__1_), .A2(
        npu_inst_pe_1_5_0_n58), .B1(npu_inst_pe_1_5_0_n113), .B2(
        npu_inst_pe_1_5_0_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_5_0_n59) );
  INV_X1 npu_inst_pe_1_5_0_U100 ( .A(npu_inst_pe_1_5_0_n59), .ZN(
        npu_inst_pe_1_5_0_n101) );
  AOI22_X1 npu_inst_pe_1_5_0_U99 ( .A1(npu_inst_int_data_y_6__0__1_), .A2(
        npu_inst_pe_1_5_0_n54), .B1(npu_inst_pe_1_5_0_n114), .B2(
        npu_inst_pe_1_5_0_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_5_0_n55) );
  INV_X1 npu_inst_pe_1_5_0_U98 ( .A(npu_inst_pe_1_5_0_n55), .ZN(
        npu_inst_pe_1_5_0_n102) );
  AOI22_X1 npu_inst_pe_1_5_0_U97 ( .A1(npu_inst_int_data_y_6__0__1_), .A2(
        npu_inst_pe_1_5_0_n50), .B1(npu_inst_pe_1_5_0_n115), .B2(
        npu_inst_pe_1_5_0_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_5_0_n51) );
  INV_X1 npu_inst_pe_1_5_0_U96 ( .A(npu_inst_pe_1_5_0_n51), .ZN(
        npu_inst_pe_1_5_0_n103) );
  AOI22_X1 npu_inst_pe_1_5_0_U95 ( .A1(npu_inst_int_data_y_6__0__1_), .A2(
        npu_inst_pe_1_5_0_n46), .B1(npu_inst_pe_1_5_0_n116), .B2(
        npu_inst_pe_1_5_0_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_5_0_n47) );
  INV_X1 npu_inst_pe_1_5_0_U94 ( .A(npu_inst_pe_1_5_0_n47), .ZN(
        npu_inst_pe_1_5_0_n104) );
  AOI22_X1 npu_inst_pe_1_5_0_U93 ( .A1(npu_inst_int_data_y_6__0__1_), .A2(
        npu_inst_pe_1_5_0_n42), .B1(npu_inst_pe_1_5_0_n118), .B2(
        npu_inst_pe_1_5_0_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_5_0_n43) );
  INV_X1 npu_inst_pe_1_5_0_U92 ( .A(npu_inst_pe_1_5_0_n43), .ZN(
        npu_inst_pe_1_5_0_n105) );
  AOI22_X1 npu_inst_pe_1_5_0_U91 ( .A1(npu_inst_pe_1_5_0_n38), .A2(
        npu_inst_int_data_y_6__0__1_), .B1(npu_inst_pe_1_5_0_n117), .B2(
        npu_inst_pe_1_5_0_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_5_0_n39) );
  INV_X1 npu_inst_pe_1_5_0_U90 ( .A(npu_inst_pe_1_5_0_n39), .ZN(
        npu_inst_pe_1_5_0_n106) );
  AOI22_X1 npu_inst_pe_1_5_0_U89 ( .A1(npu_inst_pe_1_5_0_n38), .A2(
        npu_inst_int_data_y_6__0__0_), .B1(npu_inst_pe_1_5_0_n117), .B2(
        npu_inst_pe_1_5_0_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_5_0_n37) );
  INV_X1 npu_inst_pe_1_5_0_U88 ( .A(npu_inst_pe_1_5_0_n37), .ZN(
        npu_inst_pe_1_5_0_n112) );
  NAND2_X1 npu_inst_pe_1_5_0_U87 ( .A1(npu_inst_pe_1_5_0_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_5_0_n60), .ZN(npu_inst_pe_1_5_0_n74) );
  OAI21_X1 npu_inst_pe_1_5_0_U86 ( .B1(npu_inst_pe_1_5_0_n63), .B2(
        npu_inst_pe_1_5_0_n60), .A(npu_inst_pe_1_5_0_n74), .ZN(
        npu_inst_pe_1_5_0_n97) );
  NAND2_X1 npu_inst_pe_1_5_0_U85 ( .A1(npu_inst_pe_1_5_0_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_5_0_n60), .ZN(npu_inst_pe_1_5_0_n73) );
  OAI21_X1 npu_inst_pe_1_5_0_U84 ( .B1(npu_inst_pe_1_5_0_n61), .B2(
        npu_inst_pe_1_5_0_n60), .A(npu_inst_pe_1_5_0_n73), .ZN(
        npu_inst_pe_1_5_0_n96) );
  NAND2_X1 npu_inst_pe_1_5_0_U83 ( .A1(npu_inst_pe_1_5_0_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_5_0_n56), .ZN(npu_inst_pe_1_5_0_n72) );
  OAI21_X1 npu_inst_pe_1_5_0_U82 ( .B1(npu_inst_pe_1_5_0_n63), .B2(
        npu_inst_pe_1_5_0_n56), .A(npu_inst_pe_1_5_0_n72), .ZN(
        npu_inst_pe_1_5_0_n95) );
  NAND2_X1 npu_inst_pe_1_5_0_U81 ( .A1(npu_inst_pe_1_5_0_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_5_0_n56), .ZN(npu_inst_pe_1_5_0_n71) );
  OAI21_X1 npu_inst_pe_1_5_0_U80 ( .B1(npu_inst_pe_1_5_0_n61), .B2(
        npu_inst_pe_1_5_0_n56), .A(npu_inst_pe_1_5_0_n71), .ZN(
        npu_inst_pe_1_5_0_n94) );
  NAND2_X1 npu_inst_pe_1_5_0_U79 ( .A1(npu_inst_pe_1_5_0_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_5_0_n52), .ZN(npu_inst_pe_1_5_0_n70) );
  OAI21_X1 npu_inst_pe_1_5_0_U78 ( .B1(npu_inst_pe_1_5_0_n63), .B2(
        npu_inst_pe_1_5_0_n52), .A(npu_inst_pe_1_5_0_n70), .ZN(
        npu_inst_pe_1_5_0_n93) );
  NAND2_X1 npu_inst_pe_1_5_0_U77 ( .A1(npu_inst_pe_1_5_0_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_5_0_n52), .ZN(npu_inst_pe_1_5_0_n69) );
  OAI21_X1 npu_inst_pe_1_5_0_U76 ( .B1(npu_inst_pe_1_5_0_n61), .B2(
        npu_inst_pe_1_5_0_n52), .A(npu_inst_pe_1_5_0_n69), .ZN(
        npu_inst_pe_1_5_0_n92) );
  NAND2_X1 npu_inst_pe_1_5_0_U75 ( .A1(npu_inst_pe_1_5_0_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_5_0_n48), .ZN(npu_inst_pe_1_5_0_n68) );
  OAI21_X1 npu_inst_pe_1_5_0_U74 ( .B1(npu_inst_pe_1_5_0_n63), .B2(
        npu_inst_pe_1_5_0_n48), .A(npu_inst_pe_1_5_0_n68), .ZN(
        npu_inst_pe_1_5_0_n91) );
  NAND2_X1 npu_inst_pe_1_5_0_U73 ( .A1(npu_inst_pe_1_5_0_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_5_0_n48), .ZN(npu_inst_pe_1_5_0_n67) );
  OAI21_X1 npu_inst_pe_1_5_0_U72 ( .B1(npu_inst_pe_1_5_0_n61), .B2(
        npu_inst_pe_1_5_0_n48), .A(npu_inst_pe_1_5_0_n67), .ZN(
        npu_inst_pe_1_5_0_n90) );
  NAND2_X1 npu_inst_pe_1_5_0_U71 ( .A1(npu_inst_pe_1_5_0_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_5_0_n44), .ZN(npu_inst_pe_1_5_0_n66) );
  OAI21_X1 npu_inst_pe_1_5_0_U70 ( .B1(npu_inst_pe_1_5_0_n63), .B2(
        npu_inst_pe_1_5_0_n44), .A(npu_inst_pe_1_5_0_n66), .ZN(
        npu_inst_pe_1_5_0_n89) );
  NAND2_X1 npu_inst_pe_1_5_0_U69 ( .A1(npu_inst_pe_1_5_0_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_5_0_n44), .ZN(npu_inst_pe_1_5_0_n65) );
  OAI21_X1 npu_inst_pe_1_5_0_U68 ( .B1(npu_inst_pe_1_5_0_n61), .B2(
        npu_inst_pe_1_5_0_n44), .A(npu_inst_pe_1_5_0_n65), .ZN(
        npu_inst_pe_1_5_0_n88) );
  NAND2_X1 npu_inst_pe_1_5_0_U67 ( .A1(npu_inst_pe_1_5_0_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_5_0_n40), .ZN(npu_inst_pe_1_5_0_n64) );
  OAI21_X1 npu_inst_pe_1_5_0_U66 ( .B1(npu_inst_pe_1_5_0_n63), .B2(
        npu_inst_pe_1_5_0_n40), .A(npu_inst_pe_1_5_0_n64), .ZN(
        npu_inst_pe_1_5_0_n87) );
  NAND2_X1 npu_inst_pe_1_5_0_U65 ( .A1(npu_inst_pe_1_5_0_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_5_0_n40), .ZN(npu_inst_pe_1_5_0_n62) );
  OAI21_X1 npu_inst_pe_1_5_0_U64 ( .B1(npu_inst_pe_1_5_0_n61), .B2(
        npu_inst_pe_1_5_0_n40), .A(npu_inst_pe_1_5_0_n62), .ZN(
        npu_inst_pe_1_5_0_n86) );
  AND2_X1 npu_inst_pe_1_5_0_U63 ( .A1(npu_inst_pe_1_5_0_N93), .A2(npu_inst_n55), .ZN(npu_inst_int_data_y_5__0__0_) );
  AND2_X1 npu_inst_pe_1_5_0_U62 ( .A1(npu_inst_n55), .A2(npu_inst_pe_1_5_0_N94), .ZN(npu_inst_int_data_y_5__0__1_) );
  NOR3_X1 npu_inst_pe_1_5_0_U61 ( .A1(npu_inst_pe_1_5_0_n26), .A2(npu_inst_n55), .A3(npu_inst_int_ckg[23]), .ZN(npu_inst_pe_1_5_0_n85) );
  OR2_X1 npu_inst_pe_1_5_0_U60 ( .A1(npu_inst_pe_1_5_0_n85), .A2(
        npu_inst_pe_1_5_0_n2), .ZN(npu_inst_pe_1_5_0_N84) );
  AND2_X1 npu_inst_pe_1_5_0_U59 ( .A1(npu_inst_pe_1_5_0_int_q_acc_0_), .A2(
        npu_inst_pe_1_5_0_n1), .ZN(npu_inst_int_data_res_5__0__0_) );
  AND2_X1 npu_inst_pe_1_5_0_U58 ( .A1(npu_inst_pe_1_5_0_n2), .A2(
        npu_inst_pe_1_5_0_int_q_acc_7_), .ZN(npu_inst_int_data_res_5__0__7_)
         );
  AND2_X1 npu_inst_pe_1_5_0_U57 ( .A1(npu_inst_pe_1_5_0_int_q_acc_1_), .A2(
        npu_inst_pe_1_5_0_n1), .ZN(npu_inst_int_data_res_5__0__1_) );
  AND2_X1 npu_inst_pe_1_5_0_U56 ( .A1(npu_inst_pe_1_5_0_int_q_acc_2_), .A2(
        npu_inst_pe_1_5_0_n1), .ZN(npu_inst_int_data_res_5__0__2_) );
  AND2_X1 npu_inst_pe_1_5_0_U55 ( .A1(npu_inst_pe_1_5_0_int_q_acc_3_), .A2(
        npu_inst_pe_1_5_0_n2), .ZN(npu_inst_int_data_res_5__0__3_) );
  AND2_X1 npu_inst_pe_1_5_0_U54 ( .A1(npu_inst_pe_1_5_0_int_q_acc_4_), .A2(
        npu_inst_pe_1_5_0_n2), .ZN(npu_inst_int_data_res_5__0__4_) );
  AND2_X1 npu_inst_pe_1_5_0_U53 ( .A1(npu_inst_pe_1_5_0_int_q_acc_5_), .A2(
        npu_inst_pe_1_5_0_n2), .ZN(npu_inst_int_data_res_5__0__5_) );
  AND2_X1 npu_inst_pe_1_5_0_U52 ( .A1(npu_inst_pe_1_5_0_int_q_acc_6_), .A2(
        npu_inst_pe_1_5_0_n2), .ZN(npu_inst_int_data_res_5__0__6_) );
  AOI222_X1 npu_inst_pe_1_5_0_U51 ( .A1(npu_inst_int_data_res_6__0__0_), .A2(
        npu_inst_pe_1_5_0_n1), .B1(npu_inst_pe_1_5_0_N73), .B2(
        npu_inst_pe_1_5_0_n76), .C1(npu_inst_pe_1_5_0_N65), .C2(
        npu_inst_pe_1_5_0_n77), .ZN(npu_inst_pe_1_5_0_n84) );
  INV_X1 npu_inst_pe_1_5_0_U50 ( .A(npu_inst_pe_1_5_0_n84), .ZN(
        npu_inst_pe_1_5_0_n100) );
  AOI222_X1 npu_inst_pe_1_5_0_U49 ( .A1(npu_inst_int_data_res_6__0__7_), .A2(
        npu_inst_pe_1_5_0_n1), .B1(npu_inst_pe_1_5_0_N80), .B2(
        npu_inst_pe_1_5_0_n76), .C1(npu_inst_pe_1_5_0_N72), .C2(
        npu_inst_pe_1_5_0_n77), .ZN(npu_inst_pe_1_5_0_n75) );
  INV_X1 npu_inst_pe_1_5_0_U48 ( .A(npu_inst_pe_1_5_0_n75), .ZN(
        npu_inst_pe_1_5_0_n32) );
  AOI222_X1 npu_inst_pe_1_5_0_U47 ( .A1(npu_inst_int_data_res_6__0__1_), .A2(
        npu_inst_pe_1_5_0_n1), .B1(npu_inst_pe_1_5_0_N74), .B2(
        npu_inst_pe_1_5_0_n76), .C1(npu_inst_pe_1_5_0_N66), .C2(
        npu_inst_pe_1_5_0_n77), .ZN(npu_inst_pe_1_5_0_n83) );
  INV_X1 npu_inst_pe_1_5_0_U46 ( .A(npu_inst_pe_1_5_0_n83), .ZN(
        npu_inst_pe_1_5_0_n99) );
  AOI222_X1 npu_inst_pe_1_5_0_U45 ( .A1(npu_inst_int_data_res_6__0__2_), .A2(
        npu_inst_pe_1_5_0_n1), .B1(npu_inst_pe_1_5_0_N75), .B2(
        npu_inst_pe_1_5_0_n76), .C1(npu_inst_pe_1_5_0_N67), .C2(
        npu_inst_pe_1_5_0_n77), .ZN(npu_inst_pe_1_5_0_n82) );
  INV_X1 npu_inst_pe_1_5_0_U44 ( .A(npu_inst_pe_1_5_0_n82), .ZN(
        npu_inst_pe_1_5_0_n98) );
  AOI222_X1 npu_inst_pe_1_5_0_U43 ( .A1(npu_inst_int_data_res_6__0__3_), .A2(
        npu_inst_pe_1_5_0_n1), .B1(npu_inst_pe_1_5_0_N76), .B2(
        npu_inst_pe_1_5_0_n76), .C1(npu_inst_pe_1_5_0_N68), .C2(
        npu_inst_pe_1_5_0_n77), .ZN(npu_inst_pe_1_5_0_n81) );
  INV_X1 npu_inst_pe_1_5_0_U42 ( .A(npu_inst_pe_1_5_0_n81), .ZN(
        npu_inst_pe_1_5_0_n36) );
  AOI222_X1 npu_inst_pe_1_5_0_U41 ( .A1(npu_inst_int_data_res_6__0__4_), .A2(
        npu_inst_pe_1_5_0_n1), .B1(npu_inst_pe_1_5_0_N77), .B2(
        npu_inst_pe_1_5_0_n76), .C1(npu_inst_pe_1_5_0_N69), .C2(
        npu_inst_pe_1_5_0_n77), .ZN(npu_inst_pe_1_5_0_n80) );
  INV_X1 npu_inst_pe_1_5_0_U40 ( .A(npu_inst_pe_1_5_0_n80), .ZN(
        npu_inst_pe_1_5_0_n35) );
  AOI222_X1 npu_inst_pe_1_5_0_U39 ( .A1(npu_inst_int_data_res_6__0__5_), .A2(
        npu_inst_pe_1_5_0_n1), .B1(npu_inst_pe_1_5_0_N78), .B2(
        npu_inst_pe_1_5_0_n76), .C1(npu_inst_pe_1_5_0_N70), .C2(
        npu_inst_pe_1_5_0_n77), .ZN(npu_inst_pe_1_5_0_n79) );
  INV_X1 npu_inst_pe_1_5_0_U38 ( .A(npu_inst_pe_1_5_0_n79), .ZN(
        npu_inst_pe_1_5_0_n34) );
  AOI222_X1 npu_inst_pe_1_5_0_U37 ( .A1(npu_inst_int_data_res_6__0__6_), .A2(
        npu_inst_pe_1_5_0_n1), .B1(npu_inst_pe_1_5_0_N79), .B2(
        npu_inst_pe_1_5_0_n76), .C1(npu_inst_pe_1_5_0_N71), .C2(
        npu_inst_pe_1_5_0_n77), .ZN(npu_inst_pe_1_5_0_n78) );
  INV_X1 npu_inst_pe_1_5_0_U36 ( .A(npu_inst_pe_1_5_0_n78), .ZN(
        npu_inst_pe_1_5_0_n33) );
  AND2_X1 npu_inst_pe_1_5_0_U35 ( .A1(npu_inst_pe_1_5_0_o_data_h_1_), .A2(
        npu_inst_pe_1_5_0_int_q_weight_1_), .ZN(npu_inst_pe_1_5_0_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_5_0_U34 ( .A1(npu_inst_pe_1_5_0_o_data_h_0_), .A2(
        npu_inst_pe_1_5_0_int_q_weight_1_), .ZN(npu_inst_pe_1_5_0_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_5_0_U33 ( .A(npu_inst_pe_1_5_0_int_data_1_), .ZN(
        npu_inst_pe_1_5_0_n13) );
  AOI22_X1 npu_inst_pe_1_5_0_U32 ( .A1(npu_inst_n55), .A2(
        npu_inst_int_data_y_6__0__1_), .B1(npu_inst_pe_1_5_0_n3), .B2(
        npu_inst_int_data_x_5__1__1_), .ZN(npu_inst_pe_1_5_0_n63) );
  AOI22_X1 npu_inst_pe_1_5_0_U31 ( .A1(npu_inst_n55), .A2(
        npu_inst_int_data_y_6__0__0_), .B1(npu_inst_pe_1_5_0_n3), .B2(
        npu_inst_int_data_x_5__1__0_), .ZN(npu_inst_pe_1_5_0_n61) );
  INV_X1 npu_inst_pe_1_5_0_U30 ( .A(npu_inst_pe_1_5_0_int_data_0_), .ZN(
        npu_inst_pe_1_5_0_n12) );
  INV_X1 npu_inst_pe_1_5_0_U29 ( .A(npu_inst_n68), .ZN(npu_inst_pe_1_5_0_n5)
         );
  OR3_X1 npu_inst_pe_1_5_0_U28 ( .A1(npu_inst_n76), .A2(npu_inst_pe_1_5_0_n7), 
        .A3(npu_inst_pe_1_5_0_n5), .ZN(npu_inst_pe_1_5_0_n56) );
  OR3_X1 npu_inst_pe_1_5_0_U27 ( .A1(npu_inst_pe_1_5_0_n5), .A2(
        npu_inst_pe_1_5_0_n7), .A3(npu_inst_pe_1_5_0_n6), .ZN(
        npu_inst_pe_1_5_0_n48) );
  INV_X1 npu_inst_pe_1_5_0_U26 ( .A(npu_inst_pe_1_5_0_n5), .ZN(
        npu_inst_pe_1_5_0_n4) );
  INV_X1 npu_inst_pe_1_5_0_U25 ( .A(npu_inst_n123), .ZN(npu_inst_pe_1_5_0_n11)
         );
  OR3_X1 npu_inst_pe_1_5_0_U24 ( .A1(npu_inst_pe_1_5_0_n4), .A2(
        npu_inst_pe_1_5_0_n7), .A3(npu_inst_pe_1_5_0_n6), .ZN(
        npu_inst_pe_1_5_0_n52) );
  OR3_X1 npu_inst_pe_1_5_0_U23 ( .A1(npu_inst_n76), .A2(npu_inst_pe_1_5_0_n7), 
        .A3(npu_inst_pe_1_5_0_n4), .ZN(npu_inst_pe_1_5_0_n60) );
  NOR2_X1 npu_inst_pe_1_5_0_U22 ( .A1(npu_inst_pe_1_5_0_n60), .A2(
        npu_inst_pe_1_5_0_n3), .ZN(npu_inst_pe_1_5_0_n58) );
  NOR2_X1 npu_inst_pe_1_5_0_U21 ( .A1(npu_inst_pe_1_5_0_n56), .A2(
        npu_inst_pe_1_5_0_n3), .ZN(npu_inst_pe_1_5_0_n54) );
  NOR2_X1 npu_inst_pe_1_5_0_U20 ( .A1(npu_inst_pe_1_5_0_n52), .A2(
        npu_inst_pe_1_5_0_n3), .ZN(npu_inst_pe_1_5_0_n50) );
  NOR2_X1 npu_inst_pe_1_5_0_U19 ( .A1(npu_inst_pe_1_5_0_n48), .A2(
        npu_inst_pe_1_5_0_n3), .ZN(npu_inst_pe_1_5_0_n46) );
  NOR2_X1 npu_inst_pe_1_5_0_U18 ( .A1(npu_inst_pe_1_5_0_n40), .A2(
        npu_inst_pe_1_5_0_n3), .ZN(npu_inst_pe_1_5_0_n38) );
  NOR2_X1 npu_inst_pe_1_5_0_U17 ( .A1(npu_inst_pe_1_5_0_n44), .A2(
        npu_inst_pe_1_5_0_n3), .ZN(npu_inst_pe_1_5_0_n42) );
  BUF_X1 npu_inst_pe_1_5_0_U16 ( .A(npu_inst_n97), .Z(npu_inst_pe_1_5_0_n7) );
  BUF_X1 npu_inst_pe_1_5_0_U15 ( .A(npu_inst_pe_1_5_0_n11), .Z(
        npu_inst_pe_1_5_0_n10) );
  BUF_X1 npu_inst_pe_1_5_0_U14 ( .A(npu_inst_pe_1_5_0_n11), .Z(
        npu_inst_pe_1_5_0_n9) );
  BUF_X1 npu_inst_pe_1_5_0_U13 ( .A(npu_inst_pe_1_5_0_n11), .Z(
        npu_inst_pe_1_5_0_n8) );
  INV_X1 npu_inst_pe_1_5_0_U12 ( .A(npu_inst_pe_1_5_0_n38), .ZN(
        npu_inst_pe_1_5_0_n117) );
  INV_X1 npu_inst_pe_1_5_0_U11 ( .A(npu_inst_pe_1_5_0_n58), .ZN(
        npu_inst_pe_1_5_0_n113) );
  INV_X1 npu_inst_pe_1_5_0_U10 ( .A(npu_inst_pe_1_5_0_n54), .ZN(
        npu_inst_pe_1_5_0_n114) );
  INV_X1 npu_inst_pe_1_5_0_U9 ( .A(npu_inst_pe_1_5_0_n50), .ZN(
        npu_inst_pe_1_5_0_n115) );
  INV_X1 npu_inst_pe_1_5_0_U8 ( .A(npu_inst_pe_1_5_0_n46), .ZN(
        npu_inst_pe_1_5_0_n116) );
  INV_X1 npu_inst_pe_1_5_0_U7 ( .A(npu_inst_pe_1_5_0_n42), .ZN(
        npu_inst_pe_1_5_0_n118) );
  BUF_X1 npu_inst_pe_1_5_0_U6 ( .A(npu_inst_n18), .Z(npu_inst_pe_1_5_0_n2) );
  BUF_X1 npu_inst_pe_1_5_0_U5 ( .A(npu_inst_n18), .Z(npu_inst_pe_1_5_0_n1) );
  NOR2_X1 npu_inst_pe_1_5_0_U4 ( .A1(npu_inst_pe_1_5_0_int_q_weight_0_), .A2(
        npu_inst_pe_1_5_0_n1), .ZN(npu_inst_pe_1_5_0_n76) );
  NOR2_X1 npu_inst_pe_1_5_0_U3 ( .A1(npu_inst_pe_1_5_0_n27), .A2(
        npu_inst_pe_1_5_0_n1), .ZN(npu_inst_pe_1_5_0_n77) );
  FA_X1 npu_inst_pe_1_5_0_sub_77_U2_1 ( .A(npu_inst_pe_1_5_0_int_q_acc_1_), 
        .B(npu_inst_pe_1_5_0_n13), .CI(npu_inst_pe_1_5_0_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_5_0_sub_77_carry_2_), .S(npu_inst_pe_1_5_0_N66) );
  FA_X1 npu_inst_pe_1_5_0_add_79_U1_1 ( .A(npu_inst_pe_1_5_0_int_q_acc_1_), 
        .B(npu_inst_pe_1_5_0_int_data_1_), .CI(
        npu_inst_pe_1_5_0_add_79_carry_1_), .CO(
        npu_inst_pe_1_5_0_add_79_carry_2_), .S(npu_inst_pe_1_5_0_N74) );
  NAND3_X1 npu_inst_pe_1_5_0_U109 ( .A1(npu_inst_pe_1_5_0_n5), .A2(
        npu_inst_pe_1_5_0_n6), .A3(npu_inst_pe_1_5_0_n7), .ZN(
        npu_inst_pe_1_5_0_n44) );
  NAND3_X1 npu_inst_pe_1_5_0_U108 ( .A1(npu_inst_pe_1_5_0_n4), .A2(
        npu_inst_pe_1_5_0_n6), .A3(npu_inst_pe_1_5_0_n7), .ZN(
        npu_inst_pe_1_5_0_n40) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_5_0_n33), .CK(
        npu_inst_pe_1_5_0_net3373), .RN(npu_inst_pe_1_5_0_n8), .Q(
        npu_inst_pe_1_5_0_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_5_0_n34), .CK(
        npu_inst_pe_1_5_0_net3373), .RN(npu_inst_pe_1_5_0_n8), .Q(
        npu_inst_pe_1_5_0_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_5_0_n35), .CK(
        npu_inst_pe_1_5_0_net3373), .RN(npu_inst_pe_1_5_0_n8), .Q(
        npu_inst_pe_1_5_0_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_5_0_n36), .CK(
        npu_inst_pe_1_5_0_net3373), .RN(npu_inst_pe_1_5_0_n8), .Q(
        npu_inst_pe_1_5_0_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_5_0_n98), .CK(
        npu_inst_pe_1_5_0_net3373), .RN(npu_inst_pe_1_5_0_n8), .Q(
        npu_inst_pe_1_5_0_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_5_0_n99), .CK(
        npu_inst_pe_1_5_0_net3373), .RN(npu_inst_pe_1_5_0_n8), .Q(
        npu_inst_pe_1_5_0_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_5_0_n32), .CK(
        npu_inst_pe_1_5_0_net3373), .RN(npu_inst_pe_1_5_0_n8), .Q(
        npu_inst_pe_1_5_0_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_5_0_n100), 
        .CK(npu_inst_pe_1_5_0_net3373), .RN(npu_inst_pe_1_5_0_n8), .Q(
        npu_inst_pe_1_5_0_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_weight_reg_0_ ( .D(npu_inst_n109), .CK(
        npu_inst_pe_1_5_0_net3379), .RN(npu_inst_pe_1_5_0_n8), .Q(
        npu_inst_pe_1_5_0_int_q_weight_0_), .QN(npu_inst_pe_1_5_0_n27) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_weight_reg_1_ ( .D(npu_inst_n115), .CK(
        npu_inst_pe_1_5_0_net3379), .RN(npu_inst_pe_1_5_0_n8), .Q(
        npu_inst_pe_1_5_0_int_q_weight_1_), .QN(npu_inst_pe_1_5_0_n26) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_5_0_n112), 
        .CK(npu_inst_pe_1_5_0_net3379), .RN(npu_inst_pe_1_5_0_n8), .Q(
        npu_inst_pe_1_5_0_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_5_0_n106), 
        .CK(npu_inst_pe_1_5_0_net3379), .RN(npu_inst_pe_1_5_0_n8), .Q(
        npu_inst_pe_1_5_0_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_5_0_n111), 
        .CK(npu_inst_pe_1_5_0_net3379), .RN(npu_inst_pe_1_5_0_n9), .Q(
        npu_inst_pe_1_5_0_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_5_0_n105), 
        .CK(npu_inst_pe_1_5_0_net3379), .RN(npu_inst_pe_1_5_0_n9), .Q(
        npu_inst_pe_1_5_0_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_5_0_n110), 
        .CK(npu_inst_pe_1_5_0_net3379), .RN(npu_inst_pe_1_5_0_n9), .Q(
        npu_inst_pe_1_5_0_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_5_0_n104), 
        .CK(npu_inst_pe_1_5_0_net3379), .RN(npu_inst_pe_1_5_0_n9), .Q(
        npu_inst_pe_1_5_0_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_5_0_n109), 
        .CK(npu_inst_pe_1_5_0_net3379), .RN(npu_inst_pe_1_5_0_n9), .Q(
        npu_inst_pe_1_5_0_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_5_0_n103), 
        .CK(npu_inst_pe_1_5_0_net3379), .RN(npu_inst_pe_1_5_0_n9), .Q(
        npu_inst_pe_1_5_0_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_5_0_n108), 
        .CK(npu_inst_pe_1_5_0_net3379), .RN(npu_inst_pe_1_5_0_n9), .Q(
        npu_inst_pe_1_5_0_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_5_0_n102), 
        .CK(npu_inst_pe_1_5_0_net3379), .RN(npu_inst_pe_1_5_0_n9), .Q(
        npu_inst_pe_1_5_0_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_5_0_n107), 
        .CK(npu_inst_pe_1_5_0_net3379), .RN(npu_inst_pe_1_5_0_n9), .Q(
        npu_inst_pe_1_5_0_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_5_0_n101), 
        .CK(npu_inst_pe_1_5_0_net3379), .RN(npu_inst_pe_1_5_0_n9), .Q(
        npu_inst_pe_1_5_0_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_5_0_n86), 
        .CK(npu_inst_pe_1_5_0_net3379), .RN(npu_inst_pe_1_5_0_n9), .Q(
        npu_inst_pe_1_5_0_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_5_0_n87), 
        .CK(npu_inst_pe_1_5_0_net3379), .RN(npu_inst_pe_1_5_0_n9), .Q(
        npu_inst_pe_1_5_0_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_5_0_n88), 
        .CK(npu_inst_pe_1_5_0_net3379), .RN(npu_inst_pe_1_5_0_n10), .Q(
        npu_inst_pe_1_5_0_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_5_0_n89), 
        .CK(npu_inst_pe_1_5_0_net3379), .RN(npu_inst_pe_1_5_0_n10), .Q(
        npu_inst_pe_1_5_0_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_5_0_n90), 
        .CK(npu_inst_pe_1_5_0_net3379), .RN(npu_inst_pe_1_5_0_n10), .Q(
        npu_inst_pe_1_5_0_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_5_0_n91), 
        .CK(npu_inst_pe_1_5_0_net3379), .RN(npu_inst_pe_1_5_0_n10), .Q(
        npu_inst_pe_1_5_0_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_5_0_n92), 
        .CK(npu_inst_pe_1_5_0_net3379), .RN(npu_inst_pe_1_5_0_n10), .Q(
        npu_inst_pe_1_5_0_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_5_0_n93), 
        .CK(npu_inst_pe_1_5_0_net3379), .RN(npu_inst_pe_1_5_0_n10), .Q(
        npu_inst_pe_1_5_0_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_5_0_n94), 
        .CK(npu_inst_pe_1_5_0_net3379), .RN(npu_inst_pe_1_5_0_n10), .Q(
        npu_inst_pe_1_5_0_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_5_0_n95), 
        .CK(npu_inst_pe_1_5_0_net3379), .RN(npu_inst_pe_1_5_0_n10), .Q(
        npu_inst_pe_1_5_0_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_5_0_n96), 
        .CK(npu_inst_pe_1_5_0_net3379), .RN(npu_inst_pe_1_5_0_n10), .Q(
        npu_inst_pe_1_5_0_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_5_0_n97), 
        .CK(npu_inst_pe_1_5_0_net3379), .RN(npu_inst_pe_1_5_0_n10), .Q(
        npu_inst_pe_1_5_0_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_5_0_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_5_0_N84), .SE(1'b0), .GCK(npu_inst_pe_1_5_0_net3373) );
  CLKGATETST_X1 npu_inst_pe_1_5_0_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n63), .SE(1'b0), .GCK(npu_inst_pe_1_5_0_net3379) );
  MUX2_X1 npu_inst_pe_1_5_1_U162 ( .A(npu_inst_pe_1_5_1_n32), .B(
        npu_inst_pe_1_5_1_n29), .S(npu_inst_pe_1_5_1_n8), .Z(
        npu_inst_pe_1_5_1_N93) );
  MUX2_X1 npu_inst_pe_1_5_1_U161 ( .A(npu_inst_pe_1_5_1_n31), .B(
        npu_inst_pe_1_5_1_n30), .S(npu_inst_pe_1_5_1_n6), .Z(
        npu_inst_pe_1_5_1_n32) );
  MUX2_X1 npu_inst_pe_1_5_1_U160 ( .A(npu_inst_pe_1_5_1_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_5_1_int_q_reg_v_1__0_), .S(npu_inst_pe_1_5_1_n4), .Z(
        npu_inst_pe_1_5_1_n31) );
  MUX2_X1 npu_inst_pe_1_5_1_U159 ( .A(npu_inst_pe_1_5_1_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_5_1_int_q_reg_v_3__0_), .S(npu_inst_pe_1_5_1_n4), .Z(
        npu_inst_pe_1_5_1_n30) );
  MUX2_X1 npu_inst_pe_1_5_1_U158 ( .A(npu_inst_pe_1_5_1_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_5_1_int_q_reg_v_5__0_), .S(npu_inst_pe_1_5_1_n4), .Z(
        npu_inst_pe_1_5_1_n29) );
  MUX2_X1 npu_inst_pe_1_5_1_U157 ( .A(npu_inst_pe_1_5_1_n28), .B(
        npu_inst_pe_1_5_1_n23), .S(npu_inst_pe_1_5_1_n8), .Z(
        npu_inst_pe_1_5_1_N94) );
  MUX2_X1 npu_inst_pe_1_5_1_U156 ( .A(npu_inst_pe_1_5_1_n25), .B(
        npu_inst_pe_1_5_1_n24), .S(npu_inst_pe_1_5_1_n6), .Z(
        npu_inst_pe_1_5_1_n28) );
  MUX2_X1 npu_inst_pe_1_5_1_U155 ( .A(npu_inst_pe_1_5_1_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_5_1_int_q_reg_v_1__1_), .S(npu_inst_pe_1_5_1_n4), .Z(
        npu_inst_pe_1_5_1_n25) );
  MUX2_X1 npu_inst_pe_1_5_1_U154 ( .A(npu_inst_pe_1_5_1_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_5_1_int_q_reg_v_3__1_), .S(npu_inst_pe_1_5_1_n4), .Z(
        npu_inst_pe_1_5_1_n24) );
  MUX2_X1 npu_inst_pe_1_5_1_U153 ( .A(npu_inst_pe_1_5_1_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_5_1_int_q_reg_v_5__1_), .S(npu_inst_pe_1_5_1_n4), .Z(
        npu_inst_pe_1_5_1_n23) );
  MUX2_X1 npu_inst_pe_1_5_1_U152 ( .A(npu_inst_pe_1_5_1_n22), .B(
        npu_inst_pe_1_5_1_n19), .S(npu_inst_pe_1_5_1_n8), .Z(
        npu_inst_int_data_x_5__1__1_) );
  MUX2_X1 npu_inst_pe_1_5_1_U151 ( .A(npu_inst_pe_1_5_1_n21), .B(
        npu_inst_pe_1_5_1_n20), .S(npu_inst_pe_1_5_1_n6), .Z(
        npu_inst_pe_1_5_1_n22) );
  MUX2_X1 npu_inst_pe_1_5_1_U150 ( .A(npu_inst_pe_1_5_1_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_5_1_int_q_reg_h_1__1_), .S(npu_inst_pe_1_5_1_n4), .Z(
        npu_inst_pe_1_5_1_n21) );
  MUX2_X1 npu_inst_pe_1_5_1_U149 ( .A(npu_inst_pe_1_5_1_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_5_1_int_q_reg_h_3__1_), .S(npu_inst_pe_1_5_1_n4), .Z(
        npu_inst_pe_1_5_1_n20) );
  MUX2_X1 npu_inst_pe_1_5_1_U148 ( .A(npu_inst_pe_1_5_1_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_5_1_int_q_reg_h_5__1_), .S(npu_inst_pe_1_5_1_n4), .Z(
        npu_inst_pe_1_5_1_n19) );
  MUX2_X1 npu_inst_pe_1_5_1_U147 ( .A(npu_inst_pe_1_5_1_n18), .B(
        npu_inst_pe_1_5_1_n15), .S(npu_inst_pe_1_5_1_n8), .Z(
        npu_inst_int_data_x_5__1__0_) );
  MUX2_X1 npu_inst_pe_1_5_1_U146 ( .A(npu_inst_pe_1_5_1_n17), .B(
        npu_inst_pe_1_5_1_n16), .S(npu_inst_pe_1_5_1_n6), .Z(
        npu_inst_pe_1_5_1_n18) );
  MUX2_X1 npu_inst_pe_1_5_1_U145 ( .A(npu_inst_pe_1_5_1_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_5_1_int_q_reg_h_1__0_), .S(npu_inst_pe_1_5_1_n4), .Z(
        npu_inst_pe_1_5_1_n17) );
  MUX2_X1 npu_inst_pe_1_5_1_U144 ( .A(npu_inst_pe_1_5_1_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_5_1_int_q_reg_h_3__0_), .S(npu_inst_pe_1_5_1_n4), .Z(
        npu_inst_pe_1_5_1_n16) );
  MUX2_X1 npu_inst_pe_1_5_1_U143 ( .A(npu_inst_pe_1_5_1_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_5_1_int_q_reg_h_5__0_), .S(npu_inst_pe_1_5_1_n4), .Z(
        npu_inst_pe_1_5_1_n15) );
  XOR2_X1 npu_inst_pe_1_5_1_U142 ( .A(npu_inst_pe_1_5_1_int_data_0_), .B(
        npu_inst_pe_1_5_1_int_q_acc_0_), .Z(npu_inst_pe_1_5_1_N73) );
  AND2_X1 npu_inst_pe_1_5_1_U141 ( .A1(npu_inst_pe_1_5_1_int_q_acc_0_), .A2(
        npu_inst_pe_1_5_1_int_data_0_), .ZN(npu_inst_pe_1_5_1_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_5_1_U140 ( .A(npu_inst_pe_1_5_1_int_q_acc_0_), .B(
        npu_inst_pe_1_5_1_n13), .ZN(npu_inst_pe_1_5_1_N65) );
  OR2_X1 npu_inst_pe_1_5_1_U139 ( .A1(npu_inst_pe_1_5_1_n13), .A2(
        npu_inst_pe_1_5_1_int_q_acc_0_), .ZN(npu_inst_pe_1_5_1_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_5_1_U138 ( .A(npu_inst_pe_1_5_1_int_q_acc_2_), .B(
        npu_inst_pe_1_5_1_add_79_carry_2_), .Z(npu_inst_pe_1_5_1_N75) );
  AND2_X1 npu_inst_pe_1_5_1_U137 ( .A1(npu_inst_pe_1_5_1_add_79_carry_2_), 
        .A2(npu_inst_pe_1_5_1_int_q_acc_2_), .ZN(
        npu_inst_pe_1_5_1_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_5_1_U136 ( .A(npu_inst_pe_1_5_1_int_q_acc_3_), .B(
        npu_inst_pe_1_5_1_add_79_carry_3_), .Z(npu_inst_pe_1_5_1_N76) );
  AND2_X1 npu_inst_pe_1_5_1_U135 ( .A1(npu_inst_pe_1_5_1_add_79_carry_3_), 
        .A2(npu_inst_pe_1_5_1_int_q_acc_3_), .ZN(
        npu_inst_pe_1_5_1_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_5_1_U134 ( .A(npu_inst_pe_1_5_1_int_q_acc_4_), .B(
        npu_inst_pe_1_5_1_add_79_carry_4_), .Z(npu_inst_pe_1_5_1_N77) );
  AND2_X1 npu_inst_pe_1_5_1_U133 ( .A1(npu_inst_pe_1_5_1_add_79_carry_4_), 
        .A2(npu_inst_pe_1_5_1_int_q_acc_4_), .ZN(
        npu_inst_pe_1_5_1_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_5_1_U132 ( .A(npu_inst_pe_1_5_1_int_q_acc_5_), .B(
        npu_inst_pe_1_5_1_add_79_carry_5_), .Z(npu_inst_pe_1_5_1_N78) );
  AND2_X1 npu_inst_pe_1_5_1_U131 ( .A1(npu_inst_pe_1_5_1_add_79_carry_5_), 
        .A2(npu_inst_pe_1_5_1_int_q_acc_5_), .ZN(
        npu_inst_pe_1_5_1_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_5_1_U130 ( .A(npu_inst_pe_1_5_1_int_q_acc_6_), .B(
        npu_inst_pe_1_5_1_add_79_carry_6_), .Z(npu_inst_pe_1_5_1_N79) );
  AND2_X1 npu_inst_pe_1_5_1_U129 ( .A1(npu_inst_pe_1_5_1_add_79_carry_6_), 
        .A2(npu_inst_pe_1_5_1_int_q_acc_6_), .ZN(
        npu_inst_pe_1_5_1_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_5_1_U128 ( .A(npu_inst_pe_1_5_1_int_q_acc_7_), .B(
        npu_inst_pe_1_5_1_add_79_carry_7_), .Z(npu_inst_pe_1_5_1_N80) );
  XNOR2_X1 npu_inst_pe_1_5_1_U127 ( .A(npu_inst_pe_1_5_1_sub_77_carry_2_), .B(
        npu_inst_pe_1_5_1_int_q_acc_2_), .ZN(npu_inst_pe_1_5_1_N67) );
  OR2_X1 npu_inst_pe_1_5_1_U126 ( .A1(npu_inst_pe_1_5_1_int_q_acc_2_), .A2(
        npu_inst_pe_1_5_1_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_5_1_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_5_1_U125 ( .A(npu_inst_pe_1_5_1_sub_77_carry_3_), .B(
        npu_inst_pe_1_5_1_int_q_acc_3_), .ZN(npu_inst_pe_1_5_1_N68) );
  OR2_X1 npu_inst_pe_1_5_1_U124 ( .A1(npu_inst_pe_1_5_1_int_q_acc_3_), .A2(
        npu_inst_pe_1_5_1_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_5_1_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_5_1_U123 ( .A(npu_inst_pe_1_5_1_sub_77_carry_4_), .B(
        npu_inst_pe_1_5_1_int_q_acc_4_), .ZN(npu_inst_pe_1_5_1_N69) );
  OR2_X1 npu_inst_pe_1_5_1_U122 ( .A1(npu_inst_pe_1_5_1_int_q_acc_4_), .A2(
        npu_inst_pe_1_5_1_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_5_1_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_5_1_U121 ( .A(npu_inst_pe_1_5_1_sub_77_carry_5_), .B(
        npu_inst_pe_1_5_1_int_q_acc_5_), .ZN(npu_inst_pe_1_5_1_N70) );
  OR2_X1 npu_inst_pe_1_5_1_U120 ( .A1(npu_inst_pe_1_5_1_int_q_acc_5_), .A2(
        npu_inst_pe_1_5_1_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_5_1_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_5_1_U119 ( .A(npu_inst_pe_1_5_1_sub_77_carry_6_), .B(
        npu_inst_pe_1_5_1_int_q_acc_6_), .ZN(npu_inst_pe_1_5_1_N71) );
  OR2_X1 npu_inst_pe_1_5_1_U118 ( .A1(npu_inst_pe_1_5_1_int_q_acc_6_), .A2(
        npu_inst_pe_1_5_1_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_5_1_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_5_1_U117 ( .A(npu_inst_pe_1_5_1_int_q_acc_7_), .B(
        npu_inst_pe_1_5_1_sub_77_carry_7_), .ZN(npu_inst_pe_1_5_1_N72) );
  INV_X1 npu_inst_pe_1_5_1_U116 ( .A(npu_inst_n76), .ZN(npu_inst_pe_1_5_1_n7)
         );
  INV_X1 npu_inst_pe_1_5_1_U115 ( .A(npu_inst_pe_1_5_1_n7), .ZN(
        npu_inst_pe_1_5_1_n6) );
  INV_X1 npu_inst_pe_1_5_1_U114 ( .A(npu_inst_n55), .ZN(npu_inst_pe_1_5_1_n3)
         );
  AOI22_X1 npu_inst_pe_1_5_1_U113 ( .A1(npu_inst_int_data_y_6__1__0_), .A2(
        npu_inst_pe_1_5_1_n58), .B1(npu_inst_pe_1_5_1_n114), .B2(
        npu_inst_pe_1_5_1_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_5_1_n57) );
  INV_X1 npu_inst_pe_1_5_1_U112 ( .A(npu_inst_pe_1_5_1_n57), .ZN(
        npu_inst_pe_1_5_1_n108) );
  AOI22_X1 npu_inst_pe_1_5_1_U111 ( .A1(npu_inst_int_data_y_6__1__0_), .A2(
        npu_inst_pe_1_5_1_n54), .B1(npu_inst_pe_1_5_1_n115), .B2(
        npu_inst_pe_1_5_1_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_5_1_n53) );
  INV_X1 npu_inst_pe_1_5_1_U110 ( .A(npu_inst_pe_1_5_1_n53), .ZN(
        npu_inst_pe_1_5_1_n109) );
  AOI22_X1 npu_inst_pe_1_5_1_U107 ( .A1(npu_inst_int_data_y_6__1__0_), .A2(
        npu_inst_pe_1_5_1_n50), .B1(npu_inst_pe_1_5_1_n116), .B2(
        npu_inst_pe_1_5_1_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_5_1_n49) );
  INV_X1 npu_inst_pe_1_5_1_U106 ( .A(npu_inst_pe_1_5_1_n49), .ZN(
        npu_inst_pe_1_5_1_n110) );
  AOI22_X1 npu_inst_pe_1_5_1_U105 ( .A1(npu_inst_int_data_y_6__1__0_), .A2(
        npu_inst_pe_1_5_1_n46), .B1(npu_inst_pe_1_5_1_n117), .B2(
        npu_inst_pe_1_5_1_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_5_1_n45) );
  INV_X1 npu_inst_pe_1_5_1_U104 ( .A(npu_inst_pe_1_5_1_n45), .ZN(
        npu_inst_pe_1_5_1_n111) );
  AOI22_X1 npu_inst_pe_1_5_1_U103 ( .A1(npu_inst_int_data_y_6__1__0_), .A2(
        npu_inst_pe_1_5_1_n42), .B1(npu_inst_pe_1_5_1_n119), .B2(
        npu_inst_pe_1_5_1_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_5_1_n41) );
  INV_X1 npu_inst_pe_1_5_1_U102 ( .A(npu_inst_pe_1_5_1_n41), .ZN(
        npu_inst_pe_1_5_1_n112) );
  AOI22_X1 npu_inst_pe_1_5_1_U101 ( .A1(npu_inst_int_data_y_6__1__1_), .A2(
        npu_inst_pe_1_5_1_n58), .B1(npu_inst_pe_1_5_1_n114), .B2(
        npu_inst_pe_1_5_1_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_5_1_n59) );
  INV_X1 npu_inst_pe_1_5_1_U100 ( .A(npu_inst_pe_1_5_1_n59), .ZN(
        npu_inst_pe_1_5_1_n102) );
  AOI22_X1 npu_inst_pe_1_5_1_U99 ( .A1(npu_inst_int_data_y_6__1__1_), .A2(
        npu_inst_pe_1_5_1_n54), .B1(npu_inst_pe_1_5_1_n115), .B2(
        npu_inst_pe_1_5_1_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_5_1_n55) );
  INV_X1 npu_inst_pe_1_5_1_U98 ( .A(npu_inst_pe_1_5_1_n55), .ZN(
        npu_inst_pe_1_5_1_n103) );
  AOI22_X1 npu_inst_pe_1_5_1_U97 ( .A1(npu_inst_int_data_y_6__1__1_), .A2(
        npu_inst_pe_1_5_1_n50), .B1(npu_inst_pe_1_5_1_n116), .B2(
        npu_inst_pe_1_5_1_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_5_1_n51) );
  INV_X1 npu_inst_pe_1_5_1_U96 ( .A(npu_inst_pe_1_5_1_n51), .ZN(
        npu_inst_pe_1_5_1_n104) );
  AOI22_X1 npu_inst_pe_1_5_1_U95 ( .A1(npu_inst_int_data_y_6__1__1_), .A2(
        npu_inst_pe_1_5_1_n46), .B1(npu_inst_pe_1_5_1_n117), .B2(
        npu_inst_pe_1_5_1_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_5_1_n47) );
  INV_X1 npu_inst_pe_1_5_1_U94 ( .A(npu_inst_pe_1_5_1_n47), .ZN(
        npu_inst_pe_1_5_1_n105) );
  AOI22_X1 npu_inst_pe_1_5_1_U93 ( .A1(npu_inst_int_data_y_6__1__1_), .A2(
        npu_inst_pe_1_5_1_n42), .B1(npu_inst_pe_1_5_1_n119), .B2(
        npu_inst_pe_1_5_1_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_5_1_n43) );
  INV_X1 npu_inst_pe_1_5_1_U92 ( .A(npu_inst_pe_1_5_1_n43), .ZN(
        npu_inst_pe_1_5_1_n106) );
  AOI22_X1 npu_inst_pe_1_5_1_U91 ( .A1(npu_inst_pe_1_5_1_n38), .A2(
        npu_inst_int_data_y_6__1__1_), .B1(npu_inst_pe_1_5_1_n118), .B2(
        npu_inst_pe_1_5_1_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_5_1_n39) );
  INV_X1 npu_inst_pe_1_5_1_U90 ( .A(npu_inst_pe_1_5_1_n39), .ZN(
        npu_inst_pe_1_5_1_n107) );
  AOI22_X1 npu_inst_pe_1_5_1_U89 ( .A1(npu_inst_pe_1_5_1_n38), .A2(
        npu_inst_int_data_y_6__1__0_), .B1(npu_inst_pe_1_5_1_n118), .B2(
        npu_inst_pe_1_5_1_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_5_1_n37) );
  INV_X1 npu_inst_pe_1_5_1_U88 ( .A(npu_inst_pe_1_5_1_n37), .ZN(
        npu_inst_pe_1_5_1_n113) );
  NAND2_X1 npu_inst_pe_1_5_1_U87 ( .A1(npu_inst_pe_1_5_1_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_5_1_n60), .ZN(npu_inst_pe_1_5_1_n74) );
  OAI21_X1 npu_inst_pe_1_5_1_U86 ( .B1(npu_inst_pe_1_5_1_n63), .B2(
        npu_inst_pe_1_5_1_n60), .A(npu_inst_pe_1_5_1_n74), .ZN(
        npu_inst_pe_1_5_1_n97) );
  NAND2_X1 npu_inst_pe_1_5_1_U85 ( .A1(npu_inst_pe_1_5_1_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_5_1_n60), .ZN(npu_inst_pe_1_5_1_n73) );
  OAI21_X1 npu_inst_pe_1_5_1_U84 ( .B1(npu_inst_pe_1_5_1_n61), .B2(
        npu_inst_pe_1_5_1_n60), .A(npu_inst_pe_1_5_1_n73), .ZN(
        npu_inst_pe_1_5_1_n96) );
  NAND2_X1 npu_inst_pe_1_5_1_U83 ( .A1(npu_inst_pe_1_5_1_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_5_1_n56), .ZN(npu_inst_pe_1_5_1_n72) );
  OAI21_X1 npu_inst_pe_1_5_1_U82 ( .B1(npu_inst_pe_1_5_1_n63), .B2(
        npu_inst_pe_1_5_1_n56), .A(npu_inst_pe_1_5_1_n72), .ZN(
        npu_inst_pe_1_5_1_n95) );
  NAND2_X1 npu_inst_pe_1_5_1_U81 ( .A1(npu_inst_pe_1_5_1_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_5_1_n56), .ZN(npu_inst_pe_1_5_1_n71) );
  OAI21_X1 npu_inst_pe_1_5_1_U80 ( .B1(npu_inst_pe_1_5_1_n61), .B2(
        npu_inst_pe_1_5_1_n56), .A(npu_inst_pe_1_5_1_n71), .ZN(
        npu_inst_pe_1_5_1_n94) );
  NAND2_X1 npu_inst_pe_1_5_1_U79 ( .A1(npu_inst_pe_1_5_1_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_5_1_n52), .ZN(npu_inst_pe_1_5_1_n70) );
  OAI21_X1 npu_inst_pe_1_5_1_U78 ( .B1(npu_inst_pe_1_5_1_n63), .B2(
        npu_inst_pe_1_5_1_n52), .A(npu_inst_pe_1_5_1_n70), .ZN(
        npu_inst_pe_1_5_1_n93) );
  NAND2_X1 npu_inst_pe_1_5_1_U77 ( .A1(npu_inst_pe_1_5_1_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_5_1_n52), .ZN(npu_inst_pe_1_5_1_n69) );
  OAI21_X1 npu_inst_pe_1_5_1_U76 ( .B1(npu_inst_pe_1_5_1_n61), .B2(
        npu_inst_pe_1_5_1_n52), .A(npu_inst_pe_1_5_1_n69), .ZN(
        npu_inst_pe_1_5_1_n92) );
  NAND2_X1 npu_inst_pe_1_5_1_U75 ( .A1(npu_inst_pe_1_5_1_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_5_1_n48), .ZN(npu_inst_pe_1_5_1_n68) );
  OAI21_X1 npu_inst_pe_1_5_1_U74 ( .B1(npu_inst_pe_1_5_1_n63), .B2(
        npu_inst_pe_1_5_1_n48), .A(npu_inst_pe_1_5_1_n68), .ZN(
        npu_inst_pe_1_5_1_n91) );
  NAND2_X1 npu_inst_pe_1_5_1_U73 ( .A1(npu_inst_pe_1_5_1_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_5_1_n48), .ZN(npu_inst_pe_1_5_1_n67) );
  OAI21_X1 npu_inst_pe_1_5_1_U72 ( .B1(npu_inst_pe_1_5_1_n61), .B2(
        npu_inst_pe_1_5_1_n48), .A(npu_inst_pe_1_5_1_n67), .ZN(
        npu_inst_pe_1_5_1_n90) );
  NAND2_X1 npu_inst_pe_1_5_1_U71 ( .A1(npu_inst_pe_1_5_1_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_5_1_n44), .ZN(npu_inst_pe_1_5_1_n66) );
  OAI21_X1 npu_inst_pe_1_5_1_U70 ( .B1(npu_inst_pe_1_5_1_n63), .B2(
        npu_inst_pe_1_5_1_n44), .A(npu_inst_pe_1_5_1_n66), .ZN(
        npu_inst_pe_1_5_1_n89) );
  NAND2_X1 npu_inst_pe_1_5_1_U69 ( .A1(npu_inst_pe_1_5_1_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_5_1_n44), .ZN(npu_inst_pe_1_5_1_n65) );
  OAI21_X1 npu_inst_pe_1_5_1_U68 ( .B1(npu_inst_pe_1_5_1_n61), .B2(
        npu_inst_pe_1_5_1_n44), .A(npu_inst_pe_1_5_1_n65), .ZN(
        npu_inst_pe_1_5_1_n88) );
  NAND2_X1 npu_inst_pe_1_5_1_U67 ( .A1(npu_inst_pe_1_5_1_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_5_1_n40), .ZN(npu_inst_pe_1_5_1_n64) );
  OAI21_X1 npu_inst_pe_1_5_1_U66 ( .B1(npu_inst_pe_1_5_1_n63), .B2(
        npu_inst_pe_1_5_1_n40), .A(npu_inst_pe_1_5_1_n64), .ZN(
        npu_inst_pe_1_5_1_n87) );
  NAND2_X1 npu_inst_pe_1_5_1_U65 ( .A1(npu_inst_pe_1_5_1_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_5_1_n40), .ZN(npu_inst_pe_1_5_1_n62) );
  OAI21_X1 npu_inst_pe_1_5_1_U64 ( .B1(npu_inst_pe_1_5_1_n61), .B2(
        npu_inst_pe_1_5_1_n40), .A(npu_inst_pe_1_5_1_n62), .ZN(
        npu_inst_pe_1_5_1_n86) );
  AND2_X1 npu_inst_pe_1_5_1_U63 ( .A1(npu_inst_pe_1_5_1_N93), .A2(npu_inst_n55), .ZN(npu_inst_int_data_y_5__1__0_) );
  AND2_X1 npu_inst_pe_1_5_1_U62 ( .A1(npu_inst_n55), .A2(npu_inst_pe_1_5_1_N94), .ZN(npu_inst_int_data_y_5__1__1_) );
  NOR3_X1 npu_inst_pe_1_5_1_U61 ( .A1(npu_inst_pe_1_5_1_n26), .A2(npu_inst_n55), .A3(npu_inst_int_ckg[22]), .ZN(npu_inst_pe_1_5_1_n85) );
  OR2_X1 npu_inst_pe_1_5_1_U60 ( .A1(npu_inst_pe_1_5_1_n85), .A2(
        npu_inst_pe_1_5_1_n2), .ZN(npu_inst_pe_1_5_1_N84) );
  AND2_X1 npu_inst_pe_1_5_1_U59 ( .A1(npu_inst_pe_1_5_1_int_q_acc_0_), .A2(
        npu_inst_pe_1_5_1_n1), .ZN(npu_inst_int_data_res_5__1__0_) );
  AND2_X1 npu_inst_pe_1_5_1_U58 ( .A1(npu_inst_pe_1_5_1_n2), .A2(
        npu_inst_pe_1_5_1_int_q_acc_7_), .ZN(npu_inst_int_data_res_5__1__7_)
         );
  AND2_X1 npu_inst_pe_1_5_1_U57 ( .A1(npu_inst_pe_1_5_1_int_q_acc_1_), .A2(
        npu_inst_pe_1_5_1_n1), .ZN(npu_inst_int_data_res_5__1__1_) );
  AND2_X1 npu_inst_pe_1_5_1_U56 ( .A1(npu_inst_pe_1_5_1_int_q_acc_2_), .A2(
        npu_inst_pe_1_5_1_n1), .ZN(npu_inst_int_data_res_5__1__2_) );
  AND2_X1 npu_inst_pe_1_5_1_U55 ( .A1(npu_inst_pe_1_5_1_int_q_acc_3_), .A2(
        npu_inst_pe_1_5_1_n2), .ZN(npu_inst_int_data_res_5__1__3_) );
  AND2_X1 npu_inst_pe_1_5_1_U54 ( .A1(npu_inst_pe_1_5_1_int_q_acc_4_), .A2(
        npu_inst_pe_1_5_1_n2), .ZN(npu_inst_int_data_res_5__1__4_) );
  AND2_X1 npu_inst_pe_1_5_1_U53 ( .A1(npu_inst_pe_1_5_1_int_q_acc_5_), .A2(
        npu_inst_pe_1_5_1_n2), .ZN(npu_inst_int_data_res_5__1__5_) );
  AND2_X1 npu_inst_pe_1_5_1_U52 ( .A1(npu_inst_pe_1_5_1_int_q_acc_6_), .A2(
        npu_inst_pe_1_5_1_n2), .ZN(npu_inst_int_data_res_5__1__6_) );
  AOI222_X1 npu_inst_pe_1_5_1_U51 ( .A1(npu_inst_int_data_res_6__1__0_), .A2(
        npu_inst_pe_1_5_1_n1), .B1(npu_inst_pe_1_5_1_N73), .B2(
        npu_inst_pe_1_5_1_n76), .C1(npu_inst_pe_1_5_1_N65), .C2(
        npu_inst_pe_1_5_1_n77), .ZN(npu_inst_pe_1_5_1_n84) );
  INV_X1 npu_inst_pe_1_5_1_U50 ( .A(npu_inst_pe_1_5_1_n84), .ZN(
        npu_inst_pe_1_5_1_n101) );
  AOI222_X1 npu_inst_pe_1_5_1_U49 ( .A1(npu_inst_int_data_res_6__1__7_), .A2(
        npu_inst_pe_1_5_1_n1), .B1(npu_inst_pe_1_5_1_N80), .B2(
        npu_inst_pe_1_5_1_n76), .C1(npu_inst_pe_1_5_1_N72), .C2(
        npu_inst_pe_1_5_1_n77), .ZN(npu_inst_pe_1_5_1_n75) );
  INV_X1 npu_inst_pe_1_5_1_U48 ( .A(npu_inst_pe_1_5_1_n75), .ZN(
        npu_inst_pe_1_5_1_n33) );
  AOI222_X1 npu_inst_pe_1_5_1_U47 ( .A1(npu_inst_int_data_res_6__1__1_), .A2(
        npu_inst_pe_1_5_1_n1), .B1(npu_inst_pe_1_5_1_N74), .B2(
        npu_inst_pe_1_5_1_n76), .C1(npu_inst_pe_1_5_1_N66), .C2(
        npu_inst_pe_1_5_1_n77), .ZN(npu_inst_pe_1_5_1_n83) );
  INV_X1 npu_inst_pe_1_5_1_U46 ( .A(npu_inst_pe_1_5_1_n83), .ZN(
        npu_inst_pe_1_5_1_n100) );
  AOI222_X1 npu_inst_pe_1_5_1_U45 ( .A1(npu_inst_int_data_res_6__1__2_), .A2(
        npu_inst_pe_1_5_1_n1), .B1(npu_inst_pe_1_5_1_N75), .B2(
        npu_inst_pe_1_5_1_n76), .C1(npu_inst_pe_1_5_1_N67), .C2(
        npu_inst_pe_1_5_1_n77), .ZN(npu_inst_pe_1_5_1_n82) );
  INV_X1 npu_inst_pe_1_5_1_U44 ( .A(npu_inst_pe_1_5_1_n82), .ZN(
        npu_inst_pe_1_5_1_n99) );
  AOI222_X1 npu_inst_pe_1_5_1_U43 ( .A1(npu_inst_int_data_res_6__1__3_), .A2(
        npu_inst_pe_1_5_1_n1), .B1(npu_inst_pe_1_5_1_N76), .B2(
        npu_inst_pe_1_5_1_n76), .C1(npu_inst_pe_1_5_1_N68), .C2(
        npu_inst_pe_1_5_1_n77), .ZN(npu_inst_pe_1_5_1_n81) );
  INV_X1 npu_inst_pe_1_5_1_U42 ( .A(npu_inst_pe_1_5_1_n81), .ZN(
        npu_inst_pe_1_5_1_n98) );
  AOI222_X1 npu_inst_pe_1_5_1_U41 ( .A1(npu_inst_int_data_res_6__1__4_), .A2(
        npu_inst_pe_1_5_1_n1), .B1(npu_inst_pe_1_5_1_N77), .B2(
        npu_inst_pe_1_5_1_n76), .C1(npu_inst_pe_1_5_1_N69), .C2(
        npu_inst_pe_1_5_1_n77), .ZN(npu_inst_pe_1_5_1_n80) );
  INV_X1 npu_inst_pe_1_5_1_U40 ( .A(npu_inst_pe_1_5_1_n80), .ZN(
        npu_inst_pe_1_5_1_n36) );
  AOI222_X1 npu_inst_pe_1_5_1_U39 ( .A1(npu_inst_int_data_res_6__1__5_), .A2(
        npu_inst_pe_1_5_1_n1), .B1(npu_inst_pe_1_5_1_N78), .B2(
        npu_inst_pe_1_5_1_n76), .C1(npu_inst_pe_1_5_1_N70), .C2(
        npu_inst_pe_1_5_1_n77), .ZN(npu_inst_pe_1_5_1_n79) );
  INV_X1 npu_inst_pe_1_5_1_U38 ( .A(npu_inst_pe_1_5_1_n79), .ZN(
        npu_inst_pe_1_5_1_n35) );
  AOI222_X1 npu_inst_pe_1_5_1_U37 ( .A1(npu_inst_int_data_res_6__1__6_), .A2(
        npu_inst_pe_1_5_1_n1), .B1(npu_inst_pe_1_5_1_N79), .B2(
        npu_inst_pe_1_5_1_n76), .C1(npu_inst_pe_1_5_1_N71), .C2(
        npu_inst_pe_1_5_1_n77), .ZN(npu_inst_pe_1_5_1_n78) );
  INV_X1 npu_inst_pe_1_5_1_U36 ( .A(npu_inst_pe_1_5_1_n78), .ZN(
        npu_inst_pe_1_5_1_n34) );
  INV_X1 npu_inst_pe_1_5_1_U35 ( .A(npu_inst_pe_1_5_1_int_data_1_), .ZN(
        npu_inst_pe_1_5_1_n14) );
  AND2_X1 npu_inst_pe_1_5_1_U34 ( .A1(npu_inst_int_data_x_5__1__1_), .A2(
        npu_inst_pe_1_5_1_int_q_weight_1_), .ZN(npu_inst_pe_1_5_1_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_5_1_U33 ( .A1(npu_inst_int_data_x_5__1__0_), .A2(
        npu_inst_pe_1_5_1_int_q_weight_1_), .ZN(npu_inst_pe_1_5_1_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_5_1_U32 ( .A1(npu_inst_n55), .A2(
        npu_inst_int_data_y_6__1__1_), .B1(npu_inst_pe_1_5_1_n3), .B2(
        npu_inst_int_data_x_5__2__1_), .ZN(npu_inst_pe_1_5_1_n63) );
  AOI22_X1 npu_inst_pe_1_5_1_U31 ( .A1(npu_inst_n55), .A2(
        npu_inst_int_data_y_6__1__0_), .B1(npu_inst_pe_1_5_1_n3), .B2(
        npu_inst_int_data_x_5__2__0_), .ZN(npu_inst_pe_1_5_1_n61) );
  INV_X1 npu_inst_pe_1_5_1_U30 ( .A(npu_inst_pe_1_5_1_int_data_0_), .ZN(
        npu_inst_pe_1_5_1_n13) );
  INV_X1 npu_inst_pe_1_5_1_U29 ( .A(npu_inst_n68), .ZN(npu_inst_pe_1_5_1_n5)
         );
  OR3_X1 npu_inst_pe_1_5_1_U28 ( .A1(npu_inst_pe_1_5_1_n6), .A2(
        npu_inst_pe_1_5_1_n8), .A3(npu_inst_pe_1_5_1_n5), .ZN(
        npu_inst_pe_1_5_1_n56) );
  OR3_X1 npu_inst_pe_1_5_1_U27 ( .A1(npu_inst_pe_1_5_1_n5), .A2(
        npu_inst_pe_1_5_1_n8), .A3(npu_inst_pe_1_5_1_n7), .ZN(
        npu_inst_pe_1_5_1_n48) );
  INV_X1 npu_inst_pe_1_5_1_U26 ( .A(npu_inst_pe_1_5_1_n5), .ZN(
        npu_inst_pe_1_5_1_n4) );
  INV_X1 npu_inst_pe_1_5_1_U25 ( .A(npu_inst_n123), .ZN(npu_inst_pe_1_5_1_n12)
         );
  OR3_X1 npu_inst_pe_1_5_1_U24 ( .A1(npu_inst_pe_1_5_1_n4), .A2(
        npu_inst_pe_1_5_1_n8), .A3(npu_inst_pe_1_5_1_n7), .ZN(
        npu_inst_pe_1_5_1_n52) );
  OR3_X1 npu_inst_pe_1_5_1_U23 ( .A1(npu_inst_pe_1_5_1_n6), .A2(
        npu_inst_pe_1_5_1_n8), .A3(npu_inst_pe_1_5_1_n4), .ZN(
        npu_inst_pe_1_5_1_n60) );
  NOR2_X1 npu_inst_pe_1_5_1_U22 ( .A1(npu_inst_pe_1_5_1_n60), .A2(
        npu_inst_pe_1_5_1_n3), .ZN(npu_inst_pe_1_5_1_n58) );
  NOR2_X1 npu_inst_pe_1_5_1_U21 ( .A1(npu_inst_pe_1_5_1_n56), .A2(
        npu_inst_pe_1_5_1_n3), .ZN(npu_inst_pe_1_5_1_n54) );
  NOR2_X1 npu_inst_pe_1_5_1_U20 ( .A1(npu_inst_pe_1_5_1_n52), .A2(
        npu_inst_pe_1_5_1_n3), .ZN(npu_inst_pe_1_5_1_n50) );
  NOR2_X1 npu_inst_pe_1_5_1_U19 ( .A1(npu_inst_pe_1_5_1_n48), .A2(
        npu_inst_pe_1_5_1_n3), .ZN(npu_inst_pe_1_5_1_n46) );
  NOR2_X1 npu_inst_pe_1_5_1_U18 ( .A1(npu_inst_pe_1_5_1_n40), .A2(
        npu_inst_pe_1_5_1_n3), .ZN(npu_inst_pe_1_5_1_n38) );
  NOR2_X1 npu_inst_pe_1_5_1_U17 ( .A1(npu_inst_pe_1_5_1_n44), .A2(
        npu_inst_pe_1_5_1_n3), .ZN(npu_inst_pe_1_5_1_n42) );
  BUF_X1 npu_inst_pe_1_5_1_U16 ( .A(npu_inst_n97), .Z(npu_inst_pe_1_5_1_n8) );
  BUF_X1 npu_inst_pe_1_5_1_U15 ( .A(npu_inst_pe_1_5_1_n12), .Z(
        npu_inst_pe_1_5_1_n11) );
  BUF_X1 npu_inst_pe_1_5_1_U14 ( .A(npu_inst_pe_1_5_1_n12), .Z(
        npu_inst_pe_1_5_1_n10) );
  BUF_X1 npu_inst_pe_1_5_1_U13 ( .A(npu_inst_pe_1_5_1_n12), .Z(
        npu_inst_pe_1_5_1_n9) );
  INV_X1 npu_inst_pe_1_5_1_U12 ( .A(npu_inst_pe_1_5_1_n38), .ZN(
        npu_inst_pe_1_5_1_n118) );
  INV_X1 npu_inst_pe_1_5_1_U11 ( .A(npu_inst_pe_1_5_1_n58), .ZN(
        npu_inst_pe_1_5_1_n114) );
  INV_X1 npu_inst_pe_1_5_1_U10 ( .A(npu_inst_pe_1_5_1_n54), .ZN(
        npu_inst_pe_1_5_1_n115) );
  INV_X1 npu_inst_pe_1_5_1_U9 ( .A(npu_inst_pe_1_5_1_n50), .ZN(
        npu_inst_pe_1_5_1_n116) );
  INV_X1 npu_inst_pe_1_5_1_U8 ( .A(npu_inst_pe_1_5_1_n46), .ZN(
        npu_inst_pe_1_5_1_n117) );
  INV_X1 npu_inst_pe_1_5_1_U7 ( .A(npu_inst_pe_1_5_1_n42), .ZN(
        npu_inst_pe_1_5_1_n119) );
  BUF_X1 npu_inst_pe_1_5_1_U6 ( .A(npu_inst_n18), .Z(npu_inst_pe_1_5_1_n2) );
  BUF_X1 npu_inst_pe_1_5_1_U5 ( .A(npu_inst_n18), .Z(npu_inst_pe_1_5_1_n1) );
  NOR2_X1 npu_inst_pe_1_5_1_U4 ( .A1(npu_inst_pe_1_5_1_int_q_weight_0_), .A2(
        npu_inst_pe_1_5_1_n1), .ZN(npu_inst_pe_1_5_1_n76) );
  NOR2_X1 npu_inst_pe_1_5_1_U3 ( .A1(npu_inst_pe_1_5_1_n27), .A2(
        npu_inst_pe_1_5_1_n1), .ZN(npu_inst_pe_1_5_1_n77) );
  FA_X1 npu_inst_pe_1_5_1_sub_77_U2_1 ( .A(npu_inst_pe_1_5_1_int_q_acc_1_), 
        .B(npu_inst_pe_1_5_1_n14), .CI(npu_inst_pe_1_5_1_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_5_1_sub_77_carry_2_), .S(npu_inst_pe_1_5_1_N66) );
  FA_X1 npu_inst_pe_1_5_1_add_79_U1_1 ( .A(npu_inst_pe_1_5_1_int_q_acc_1_), 
        .B(npu_inst_pe_1_5_1_int_data_1_), .CI(
        npu_inst_pe_1_5_1_add_79_carry_1_), .CO(
        npu_inst_pe_1_5_1_add_79_carry_2_), .S(npu_inst_pe_1_5_1_N74) );
  NAND3_X1 npu_inst_pe_1_5_1_U109 ( .A1(npu_inst_pe_1_5_1_n5), .A2(
        npu_inst_pe_1_5_1_n7), .A3(npu_inst_pe_1_5_1_n8), .ZN(
        npu_inst_pe_1_5_1_n44) );
  NAND3_X1 npu_inst_pe_1_5_1_U108 ( .A1(npu_inst_pe_1_5_1_n4), .A2(
        npu_inst_pe_1_5_1_n7), .A3(npu_inst_pe_1_5_1_n8), .ZN(
        npu_inst_pe_1_5_1_n40) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_5_1_n34), .CK(
        npu_inst_pe_1_5_1_net3350), .RN(npu_inst_pe_1_5_1_n9), .Q(
        npu_inst_pe_1_5_1_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_5_1_n35), .CK(
        npu_inst_pe_1_5_1_net3350), .RN(npu_inst_pe_1_5_1_n9), .Q(
        npu_inst_pe_1_5_1_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_5_1_n36), .CK(
        npu_inst_pe_1_5_1_net3350), .RN(npu_inst_pe_1_5_1_n9), .Q(
        npu_inst_pe_1_5_1_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_5_1_n98), .CK(
        npu_inst_pe_1_5_1_net3350), .RN(npu_inst_pe_1_5_1_n9), .Q(
        npu_inst_pe_1_5_1_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_5_1_n99), .CK(
        npu_inst_pe_1_5_1_net3350), .RN(npu_inst_pe_1_5_1_n9), .Q(
        npu_inst_pe_1_5_1_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_5_1_n100), 
        .CK(npu_inst_pe_1_5_1_net3350), .RN(npu_inst_pe_1_5_1_n9), .Q(
        npu_inst_pe_1_5_1_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_5_1_n33), .CK(
        npu_inst_pe_1_5_1_net3350), .RN(npu_inst_pe_1_5_1_n9), .Q(
        npu_inst_pe_1_5_1_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_5_1_n101), 
        .CK(npu_inst_pe_1_5_1_net3350), .RN(npu_inst_pe_1_5_1_n9), .Q(
        npu_inst_pe_1_5_1_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_weight_reg_0_ ( .D(npu_inst_n109), .CK(
        npu_inst_pe_1_5_1_net3356), .RN(npu_inst_pe_1_5_1_n9), .Q(
        npu_inst_pe_1_5_1_int_q_weight_0_), .QN(npu_inst_pe_1_5_1_n27) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_weight_reg_1_ ( .D(npu_inst_n115), .CK(
        npu_inst_pe_1_5_1_net3356), .RN(npu_inst_pe_1_5_1_n9), .Q(
        npu_inst_pe_1_5_1_int_q_weight_1_), .QN(npu_inst_pe_1_5_1_n26) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_5_1_n113), 
        .CK(npu_inst_pe_1_5_1_net3356), .RN(npu_inst_pe_1_5_1_n9), .Q(
        npu_inst_pe_1_5_1_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_5_1_n107), 
        .CK(npu_inst_pe_1_5_1_net3356), .RN(npu_inst_pe_1_5_1_n9), .Q(
        npu_inst_pe_1_5_1_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_5_1_n112), 
        .CK(npu_inst_pe_1_5_1_net3356), .RN(npu_inst_pe_1_5_1_n10), .Q(
        npu_inst_pe_1_5_1_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_5_1_n106), 
        .CK(npu_inst_pe_1_5_1_net3356), .RN(npu_inst_pe_1_5_1_n10), .Q(
        npu_inst_pe_1_5_1_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_5_1_n111), 
        .CK(npu_inst_pe_1_5_1_net3356), .RN(npu_inst_pe_1_5_1_n10), .Q(
        npu_inst_pe_1_5_1_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_5_1_n105), 
        .CK(npu_inst_pe_1_5_1_net3356), .RN(npu_inst_pe_1_5_1_n10), .Q(
        npu_inst_pe_1_5_1_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_5_1_n110), 
        .CK(npu_inst_pe_1_5_1_net3356), .RN(npu_inst_pe_1_5_1_n10), .Q(
        npu_inst_pe_1_5_1_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_5_1_n104), 
        .CK(npu_inst_pe_1_5_1_net3356), .RN(npu_inst_pe_1_5_1_n10), .Q(
        npu_inst_pe_1_5_1_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_5_1_n109), 
        .CK(npu_inst_pe_1_5_1_net3356), .RN(npu_inst_pe_1_5_1_n10), .Q(
        npu_inst_pe_1_5_1_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_5_1_n103), 
        .CK(npu_inst_pe_1_5_1_net3356), .RN(npu_inst_pe_1_5_1_n10), .Q(
        npu_inst_pe_1_5_1_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_5_1_n108), 
        .CK(npu_inst_pe_1_5_1_net3356), .RN(npu_inst_pe_1_5_1_n10), .Q(
        npu_inst_pe_1_5_1_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_5_1_n102), 
        .CK(npu_inst_pe_1_5_1_net3356), .RN(npu_inst_pe_1_5_1_n10), .Q(
        npu_inst_pe_1_5_1_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_5_1_n86), 
        .CK(npu_inst_pe_1_5_1_net3356), .RN(npu_inst_pe_1_5_1_n10), .Q(
        npu_inst_pe_1_5_1_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_5_1_n87), 
        .CK(npu_inst_pe_1_5_1_net3356), .RN(npu_inst_pe_1_5_1_n10), .Q(
        npu_inst_pe_1_5_1_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_5_1_n88), 
        .CK(npu_inst_pe_1_5_1_net3356), .RN(npu_inst_pe_1_5_1_n11), .Q(
        npu_inst_pe_1_5_1_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_5_1_n89), 
        .CK(npu_inst_pe_1_5_1_net3356), .RN(npu_inst_pe_1_5_1_n11), .Q(
        npu_inst_pe_1_5_1_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_5_1_n90), 
        .CK(npu_inst_pe_1_5_1_net3356), .RN(npu_inst_pe_1_5_1_n11), .Q(
        npu_inst_pe_1_5_1_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_5_1_n91), 
        .CK(npu_inst_pe_1_5_1_net3356), .RN(npu_inst_pe_1_5_1_n11), .Q(
        npu_inst_pe_1_5_1_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_5_1_n92), 
        .CK(npu_inst_pe_1_5_1_net3356), .RN(npu_inst_pe_1_5_1_n11), .Q(
        npu_inst_pe_1_5_1_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_5_1_n93), 
        .CK(npu_inst_pe_1_5_1_net3356), .RN(npu_inst_pe_1_5_1_n11), .Q(
        npu_inst_pe_1_5_1_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_5_1_n94), 
        .CK(npu_inst_pe_1_5_1_net3356), .RN(npu_inst_pe_1_5_1_n11), .Q(
        npu_inst_pe_1_5_1_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_5_1_n95), 
        .CK(npu_inst_pe_1_5_1_net3356), .RN(npu_inst_pe_1_5_1_n11), .Q(
        npu_inst_pe_1_5_1_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_5_1_n96), 
        .CK(npu_inst_pe_1_5_1_net3356), .RN(npu_inst_pe_1_5_1_n11), .Q(
        npu_inst_pe_1_5_1_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_5_1_n97), 
        .CK(npu_inst_pe_1_5_1_net3356), .RN(npu_inst_pe_1_5_1_n11), .Q(
        npu_inst_pe_1_5_1_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_5_1_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_5_1_N84), .SE(1'b0), .GCK(npu_inst_pe_1_5_1_net3350) );
  CLKGATETST_X1 npu_inst_pe_1_5_1_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n63), .SE(1'b0), .GCK(npu_inst_pe_1_5_1_net3356) );
  MUX2_X1 npu_inst_pe_1_5_2_U162 ( .A(npu_inst_pe_1_5_2_n32), .B(
        npu_inst_pe_1_5_2_n29), .S(npu_inst_pe_1_5_2_n8), .Z(
        npu_inst_pe_1_5_2_N93) );
  MUX2_X1 npu_inst_pe_1_5_2_U161 ( .A(npu_inst_pe_1_5_2_n31), .B(
        npu_inst_pe_1_5_2_n30), .S(npu_inst_pe_1_5_2_n6), .Z(
        npu_inst_pe_1_5_2_n32) );
  MUX2_X1 npu_inst_pe_1_5_2_U160 ( .A(npu_inst_pe_1_5_2_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_5_2_int_q_reg_v_1__0_), .S(npu_inst_pe_1_5_2_n4), .Z(
        npu_inst_pe_1_5_2_n31) );
  MUX2_X1 npu_inst_pe_1_5_2_U159 ( .A(npu_inst_pe_1_5_2_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_5_2_int_q_reg_v_3__0_), .S(npu_inst_pe_1_5_2_n4), .Z(
        npu_inst_pe_1_5_2_n30) );
  MUX2_X1 npu_inst_pe_1_5_2_U158 ( .A(npu_inst_pe_1_5_2_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_5_2_int_q_reg_v_5__0_), .S(npu_inst_pe_1_5_2_n4), .Z(
        npu_inst_pe_1_5_2_n29) );
  MUX2_X1 npu_inst_pe_1_5_2_U157 ( .A(npu_inst_pe_1_5_2_n28), .B(
        npu_inst_pe_1_5_2_n23), .S(npu_inst_pe_1_5_2_n8), .Z(
        npu_inst_pe_1_5_2_N94) );
  MUX2_X1 npu_inst_pe_1_5_2_U156 ( .A(npu_inst_pe_1_5_2_n25), .B(
        npu_inst_pe_1_5_2_n24), .S(npu_inst_pe_1_5_2_n6), .Z(
        npu_inst_pe_1_5_2_n28) );
  MUX2_X1 npu_inst_pe_1_5_2_U155 ( .A(npu_inst_pe_1_5_2_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_5_2_int_q_reg_v_1__1_), .S(npu_inst_pe_1_5_2_n4), .Z(
        npu_inst_pe_1_5_2_n25) );
  MUX2_X1 npu_inst_pe_1_5_2_U154 ( .A(npu_inst_pe_1_5_2_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_5_2_int_q_reg_v_3__1_), .S(npu_inst_pe_1_5_2_n4), .Z(
        npu_inst_pe_1_5_2_n24) );
  MUX2_X1 npu_inst_pe_1_5_2_U153 ( .A(npu_inst_pe_1_5_2_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_5_2_int_q_reg_v_5__1_), .S(npu_inst_pe_1_5_2_n4), .Z(
        npu_inst_pe_1_5_2_n23) );
  MUX2_X1 npu_inst_pe_1_5_2_U152 ( .A(npu_inst_pe_1_5_2_n22), .B(
        npu_inst_pe_1_5_2_n19), .S(npu_inst_pe_1_5_2_n8), .Z(
        npu_inst_int_data_x_5__2__1_) );
  MUX2_X1 npu_inst_pe_1_5_2_U151 ( .A(npu_inst_pe_1_5_2_n21), .B(
        npu_inst_pe_1_5_2_n20), .S(npu_inst_pe_1_5_2_n6), .Z(
        npu_inst_pe_1_5_2_n22) );
  MUX2_X1 npu_inst_pe_1_5_2_U150 ( .A(npu_inst_pe_1_5_2_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_5_2_int_q_reg_h_1__1_), .S(npu_inst_pe_1_5_2_n4), .Z(
        npu_inst_pe_1_5_2_n21) );
  MUX2_X1 npu_inst_pe_1_5_2_U149 ( .A(npu_inst_pe_1_5_2_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_5_2_int_q_reg_h_3__1_), .S(npu_inst_pe_1_5_2_n4), .Z(
        npu_inst_pe_1_5_2_n20) );
  MUX2_X1 npu_inst_pe_1_5_2_U148 ( .A(npu_inst_pe_1_5_2_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_5_2_int_q_reg_h_5__1_), .S(npu_inst_pe_1_5_2_n4), .Z(
        npu_inst_pe_1_5_2_n19) );
  MUX2_X1 npu_inst_pe_1_5_2_U147 ( .A(npu_inst_pe_1_5_2_n18), .B(
        npu_inst_pe_1_5_2_n15), .S(npu_inst_pe_1_5_2_n8), .Z(
        npu_inst_int_data_x_5__2__0_) );
  MUX2_X1 npu_inst_pe_1_5_2_U146 ( .A(npu_inst_pe_1_5_2_n17), .B(
        npu_inst_pe_1_5_2_n16), .S(npu_inst_pe_1_5_2_n6), .Z(
        npu_inst_pe_1_5_2_n18) );
  MUX2_X1 npu_inst_pe_1_5_2_U145 ( .A(npu_inst_pe_1_5_2_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_5_2_int_q_reg_h_1__0_), .S(npu_inst_pe_1_5_2_n4), .Z(
        npu_inst_pe_1_5_2_n17) );
  MUX2_X1 npu_inst_pe_1_5_2_U144 ( .A(npu_inst_pe_1_5_2_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_5_2_int_q_reg_h_3__0_), .S(npu_inst_pe_1_5_2_n4), .Z(
        npu_inst_pe_1_5_2_n16) );
  MUX2_X1 npu_inst_pe_1_5_2_U143 ( .A(npu_inst_pe_1_5_2_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_5_2_int_q_reg_h_5__0_), .S(npu_inst_pe_1_5_2_n4), .Z(
        npu_inst_pe_1_5_2_n15) );
  XOR2_X1 npu_inst_pe_1_5_2_U142 ( .A(npu_inst_pe_1_5_2_int_data_0_), .B(
        npu_inst_pe_1_5_2_int_q_acc_0_), .Z(npu_inst_pe_1_5_2_N73) );
  AND2_X1 npu_inst_pe_1_5_2_U141 ( .A1(npu_inst_pe_1_5_2_int_q_acc_0_), .A2(
        npu_inst_pe_1_5_2_int_data_0_), .ZN(npu_inst_pe_1_5_2_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_5_2_U140 ( .A(npu_inst_pe_1_5_2_int_q_acc_0_), .B(
        npu_inst_pe_1_5_2_n13), .ZN(npu_inst_pe_1_5_2_N65) );
  OR2_X1 npu_inst_pe_1_5_2_U139 ( .A1(npu_inst_pe_1_5_2_n13), .A2(
        npu_inst_pe_1_5_2_int_q_acc_0_), .ZN(npu_inst_pe_1_5_2_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_5_2_U138 ( .A(npu_inst_pe_1_5_2_int_q_acc_2_), .B(
        npu_inst_pe_1_5_2_add_79_carry_2_), .Z(npu_inst_pe_1_5_2_N75) );
  AND2_X1 npu_inst_pe_1_5_2_U137 ( .A1(npu_inst_pe_1_5_2_add_79_carry_2_), 
        .A2(npu_inst_pe_1_5_2_int_q_acc_2_), .ZN(
        npu_inst_pe_1_5_2_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_5_2_U136 ( .A(npu_inst_pe_1_5_2_int_q_acc_3_), .B(
        npu_inst_pe_1_5_2_add_79_carry_3_), .Z(npu_inst_pe_1_5_2_N76) );
  AND2_X1 npu_inst_pe_1_5_2_U135 ( .A1(npu_inst_pe_1_5_2_add_79_carry_3_), 
        .A2(npu_inst_pe_1_5_2_int_q_acc_3_), .ZN(
        npu_inst_pe_1_5_2_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_5_2_U134 ( .A(npu_inst_pe_1_5_2_int_q_acc_4_), .B(
        npu_inst_pe_1_5_2_add_79_carry_4_), .Z(npu_inst_pe_1_5_2_N77) );
  AND2_X1 npu_inst_pe_1_5_2_U133 ( .A1(npu_inst_pe_1_5_2_add_79_carry_4_), 
        .A2(npu_inst_pe_1_5_2_int_q_acc_4_), .ZN(
        npu_inst_pe_1_5_2_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_5_2_U132 ( .A(npu_inst_pe_1_5_2_int_q_acc_5_), .B(
        npu_inst_pe_1_5_2_add_79_carry_5_), .Z(npu_inst_pe_1_5_2_N78) );
  AND2_X1 npu_inst_pe_1_5_2_U131 ( .A1(npu_inst_pe_1_5_2_add_79_carry_5_), 
        .A2(npu_inst_pe_1_5_2_int_q_acc_5_), .ZN(
        npu_inst_pe_1_5_2_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_5_2_U130 ( .A(npu_inst_pe_1_5_2_int_q_acc_6_), .B(
        npu_inst_pe_1_5_2_add_79_carry_6_), .Z(npu_inst_pe_1_5_2_N79) );
  AND2_X1 npu_inst_pe_1_5_2_U129 ( .A1(npu_inst_pe_1_5_2_add_79_carry_6_), 
        .A2(npu_inst_pe_1_5_2_int_q_acc_6_), .ZN(
        npu_inst_pe_1_5_2_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_5_2_U128 ( .A(npu_inst_pe_1_5_2_int_q_acc_7_), .B(
        npu_inst_pe_1_5_2_add_79_carry_7_), .Z(npu_inst_pe_1_5_2_N80) );
  XNOR2_X1 npu_inst_pe_1_5_2_U127 ( .A(npu_inst_pe_1_5_2_sub_77_carry_2_), .B(
        npu_inst_pe_1_5_2_int_q_acc_2_), .ZN(npu_inst_pe_1_5_2_N67) );
  OR2_X1 npu_inst_pe_1_5_2_U126 ( .A1(npu_inst_pe_1_5_2_int_q_acc_2_), .A2(
        npu_inst_pe_1_5_2_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_5_2_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_5_2_U125 ( .A(npu_inst_pe_1_5_2_sub_77_carry_3_), .B(
        npu_inst_pe_1_5_2_int_q_acc_3_), .ZN(npu_inst_pe_1_5_2_N68) );
  OR2_X1 npu_inst_pe_1_5_2_U124 ( .A1(npu_inst_pe_1_5_2_int_q_acc_3_), .A2(
        npu_inst_pe_1_5_2_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_5_2_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_5_2_U123 ( .A(npu_inst_pe_1_5_2_sub_77_carry_4_), .B(
        npu_inst_pe_1_5_2_int_q_acc_4_), .ZN(npu_inst_pe_1_5_2_N69) );
  OR2_X1 npu_inst_pe_1_5_2_U122 ( .A1(npu_inst_pe_1_5_2_int_q_acc_4_), .A2(
        npu_inst_pe_1_5_2_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_5_2_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_5_2_U121 ( .A(npu_inst_pe_1_5_2_sub_77_carry_5_), .B(
        npu_inst_pe_1_5_2_int_q_acc_5_), .ZN(npu_inst_pe_1_5_2_N70) );
  OR2_X1 npu_inst_pe_1_5_2_U120 ( .A1(npu_inst_pe_1_5_2_int_q_acc_5_), .A2(
        npu_inst_pe_1_5_2_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_5_2_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_5_2_U119 ( .A(npu_inst_pe_1_5_2_sub_77_carry_6_), .B(
        npu_inst_pe_1_5_2_int_q_acc_6_), .ZN(npu_inst_pe_1_5_2_N71) );
  OR2_X1 npu_inst_pe_1_5_2_U118 ( .A1(npu_inst_pe_1_5_2_int_q_acc_6_), .A2(
        npu_inst_pe_1_5_2_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_5_2_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_5_2_U117 ( .A(npu_inst_pe_1_5_2_int_q_acc_7_), .B(
        npu_inst_pe_1_5_2_sub_77_carry_7_), .ZN(npu_inst_pe_1_5_2_N72) );
  INV_X1 npu_inst_pe_1_5_2_U116 ( .A(npu_inst_n76), .ZN(npu_inst_pe_1_5_2_n7)
         );
  INV_X1 npu_inst_pe_1_5_2_U115 ( .A(npu_inst_pe_1_5_2_n7), .ZN(
        npu_inst_pe_1_5_2_n6) );
  INV_X1 npu_inst_pe_1_5_2_U114 ( .A(npu_inst_n55), .ZN(npu_inst_pe_1_5_2_n3)
         );
  AOI22_X1 npu_inst_pe_1_5_2_U113 ( .A1(npu_inst_int_data_y_6__2__0_), .A2(
        npu_inst_pe_1_5_2_n58), .B1(npu_inst_pe_1_5_2_n114), .B2(
        npu_inst_pe_1_5_2_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_5_2_n57) );
  INV_X1 npu_inst_pe_1_5_2_U112 ( .A(npu_inst_pe_1_5_2_n57), .ZN(
        npu_inst_pe_1_5_2_n108) );
  AOI22_X1 npu_inst_pe_1_5_2_U111 ( .A1(npu_inst_int_data_y_6__2__0_), .A2(
        npu_inst_pe_1_5_2_n54), .B1(npu_inst_pe_1_5_2_n115), .B2(
        npu_inst_pe_1_5_2_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_5_2_n53) );
  INV_X1 npu_inst_pe_1_5_2_U110 ( .A(npu_inst_pe_1_5_2_n53), .ZN(
        npu_inst_pe_1_5_2_n109) );
  AOI22_X1 npu_inst_pe_1_5_2_U107 ( .A1(npu_inst_int_data_y_6__2__0_), .A2(
        npu_inst_pe_1_5_2_n50), .B1(npu_inst_pe_1_5_2_n116), .B2(
        npu_inst_pe_1_5_2_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_5_2_n49) );
  INV_X1 npu_inst_pe_1_5_2_U106 ( .A(npu_inst_pe_1_5_2_n49), .ZN(
        npu_inst_pe_1_5_2_n110) );
  AOI22_X1 npu_inst_pe_1_5_2_U105 ( .A1(npu_inst_int_data_y_6__2__0_), .A2(
        npu_inst_pe_1_5_2_n46), .B1(npu_inst_pe_1_5_2_n117), .B2(
        npu_inst_pe_1_5_2_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_5_2_n45) );
  INV_X1 npu_inst_pe_1_5_2_U104 ( .A(npu_inst_pe_1_5_2_n45), .ZN(
        npu_inst_pe_1_5_2_n111) );
  AOI22_X1 npu_inst_pe_1_5_2_U103 ( .A1(npu_inst_int_data_y_6__2__0_), .A2(
        npu_inst_pe_1_5_2_n42), .B1(npu_inst_pe_1_5_2_n119), .B2(
        npu_inst_pe_1_5_2_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_5_2_n41) );
  INV_X1 npu_inst_pe_1_5_2_U102 ( .A(npu_inst_pe_1_5_2_n41), .ZN(
        npu_inst_pe_1_5_2_n112) );
  AOI22_X1 npu_inst_pe_1_5_2_U101 ( .A1(npu_inst_int_data_y_6__2__1_), .A2(
        npu_inst_pe_1_5_2_n58), .B1(npu_inst_pe_1_5_2_n114), .B2(
        npu_inst_pe_1_5_2_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_5_2_n59) );
  INV_X1 npu_inst_pe_1_5_2_U100 ( .A(npu_inst_pe_1_5_2_n59), .ZN(
        npu_inst_pe_1_5_2_n102) );
  AOI22_X1 npu_inst_pe_1_5_2_U99 ( .A1(npu_inst_int_data_y_6__2__1_), .A2(
        npu_inst_pe_1_5_2_n54), .B1(npu_inst_pe_1_5_2_n115), .B2(
        npu_inst_pe_1_5_2_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_5_2_n55) );
  INV_X1 npu_inst_pe_1_5_2_U98 ( .A(npu_inst_pe_1_5_2_n55), .ZN(
        npu_inst_pe_1_5_2_n103) );
  AOI22_X1 npu_inst_pe_1_5_2_U97 ( .A1(npu_inst_int_data_y_6__2__1_), .A2(
        npu_inst_pe_1_5_2_n50), .B1(npu_inst_pe_1_5_2_n116), .B2(
        npu_inst_pe_1_5_2_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_5_2_n51) );
  INV_X1 npu_inst_pe_1_5_2_U96 ( .A(npu_inst_pe_1_5_2_n51), .ZN(
        npu_inst_pe_1_5_2_n104) );
  AOI22_X1 npu_inst_pe_1_5_2_U95 ( .A1(npu_inst_int_data_y_6__2__1_), .A2(
        npu_inst_pe_1_5_2_n46), .B1(npu_inst_pe_1_5_2_n117), .B2(
        npu_inst_pe_1_5_2_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_5_2_n47) );
  INV_X1 npu_inst_pe_1_5_2_U94 ( .A(npu_inst_pe_1_5_2_n47), .ZN(
        npu_inst_pe_1_5_2_n105) );
  AOI22_X1 npu_inst_pe_1_5_2_U93 ( .A1(npu_inst_int_data_y_6__2__1_), .A2(
        npu_inst_pe_1_5_2_n42), .B1(npu_inst_pe_1_5_2_n119), .B2(
        npu_inst_pe_1_5_2_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_5_2_n43) );
  INV_X1 npu_inst_pe_1_5_2_U92 ( .A(npu_inst_pe_1_5_2_n43), .ZN(
        npu_inst_pe_1_5_2_n106) );
  AOI22_X1 npu_inst_pe_1_5_2_U91 ( .A1(npu_inst_pe_1_5_2_n38), .A2(
        npu_inst_int_data_y_6__2__1_), .B1(npu_inst_pe_1_5_2_n118), .B2(
        npu_inst_pe_1_5_2_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_5_2_n39) );
  INV_X1 npu_inst_pe_1_5_2_U90 ( .A(npu_inst_pe_1_5_2_n39), .ZN(
        npu_inst_pe_1_5_2_n107) );
  AOI22_X1 npu_inst_pe_1_5_2_U89 ( .A1(npu_inst_pe_1_5_2_n38), .A2(
        npu_inst_int_data_y_6__2__0_), .B1(npu_inst_pe_1_5_2_n118), .B2(
        npu_inst_pe_1_5_2_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_5_2_n37) );
  INV_X1 npu_inst_pe_1_5_2_U88 ( .A(npu_inst_pe_1_5_2_n37), .ZN(
        npu_inst_pe_1_5_2_n113) );
  NAND2_X1 npu_inst_pe_1_5_2_U87 ( .A1(npu_inst_pe_1_5_2_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_5_2_n60), .ZN(npu_inst_pe_1_5_2_n74) );
  OAI21_X1 npu_inst_pe_1_5_2_U86 ( .B1(npu_inst_pe_1_5_2_n63), .B2(
        npu_inst_pe_1_5_2_n60), .A(npu_inst_pe_1_5_2_n74), .ZN(
        npu_inst_pe_1_5_2_n97) );
  NAND2_X1 npu_inst_pe_1_5_2_U85 ( .A1(npu_inst_pe_1_5_2_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_5_2_n60), .ZN(npu_inst_pe_1_5_2_n73) );
  OAI21_X1 npu_inst_pe_1_5_2_U84 ( .B1(npu_inst_pe_1_5_2_n61), .B2(
        npu_inst_pe_1_5_2_n60), .A(npu_inst_pe_1_5_2_n73), .ZN(
        npu_inst_pe_1_5_2_n96) );
  NAND2_X1 npu_inst_pe_1_5_2_U83 ( .A1(npu_inst_pe_1_5_2_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_5_2_n56), .ZN(npu_inst_pe_1_5_2_n72) );
  OAI21_X1 npu_inst_pe_1_5_2_U82 ( .B1(npu_inst_pe_1_5_2_n63), .B2(
        npu_inst_pe_1_5_2_n56), .A(npu_inst_pe_1_5_2_n72), .ZN(
        npu_inst_pe_1_5_2_n95) );
  NAND2_X1 npu_inst_pe_1_5_2_U81 ( .A1(npu_inst_pe_1_5_2_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_5_2_n56), .ZN(npu_inst_pe_1_5_2_n71) );
  OAI21_X1 npu_inst_pe_1_5_2_U80 ( .B1(npu_inst_pe_1_5_2_n61), .B2(
        npu_inst_pe_1_5_2_n56), .A(npu_inst_pe_1_5_2_n71), .ZN(
        npu_inst_pe_1_5_2_n94) );
  NAND2_X1 npu_inst_pe_1_5_2_U79 ( .A1(npu_inst_pe_1_5_2_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_5_2_n52), .ZN(npu_inst_pe_1_5_2_n70) );
  OAI21_X1 npu_inst_pe_1_5_2_U78 ( .B1(npu_inst_pe_1_5_2_n63), .B2(
        npu_inst_pe_1_5_2_n52), .A(npu_inst_pe_1_5_2_n70), .ZN(
        npu_inst_pe_1_5_2_n93) );
  NAND2_X1 npu_inst_pe_1_5_2_U77 ( .A1(npu_inst_pe_1_5_2_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_5_2_n52), .ZN(npu_inst_pe_1_5_2_n69) );
  OAI21_X1 npu_inst_pe_1_5_2_U76 ( .B1(npu_inst_pe_1_5_2_n61), .B2(
        npu_inst_pe_1_5_2_n52), .A(npu_inst_pe_1_5_2_n69), .ZN(
        npu_inst_pe_1_5_2_n92) );
  NAND2_X1 npu_inst_pe_1_5_2_U75 ( .A1(npu_inst_pe_1_5_2_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_5_2_n48), .ZN(npu_inst_pe_1_5_2_n68) );
  OAI21_X1 npu_inst_pe_1_5_2_U74 ( .B1(npu_inst_pe_1_5_2_n63), .B2(
        npu_inst_pe_1_5_2_n48), .A(npu_inst_pe_1_5_2_n68), .ZN(
        npu_inst_pe_1_5_2_n91) );
  NAND2_X1 npu_inst_pe_1_5_2_U73 ( .A1(npu_inst_pe_1_5_2_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_5_2_n48), .ZN(npu_inst_pe_1_5_2_n67) );
  OAI21_X1 npu_inst_pe_1_5_2_U72 ( .B1(npu_inst_pe_1_5_2_n61), .B2(
        npu_inst_pe_1_5_2_n48), .A(npu_inst_pe_1_5_2_n67), .ZN(
        npu_inst_pe_1_5_2_n90) );
  NAND2_X1 npu_inst_pe_1_5_2_U71 ( .A1(npu_inst_pe_1_5_2_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_5_2_n44), .ZN(npu_inst_pe_1_5_2_n66) );
  OAI21_X1 npu_inst_pe_1_5_2_U70 ( .B1(npu_inst_pe_1_5_2_n63), .B2(
        npu_inst_pe_1_5_2_n44), .A(npu_inst_pe_1_5_2_n66), .ZN(
        npu_inst_pe_1_5_2_n89) );
  NAND2_X1 npu_inst_pe_1_5_2_U69 ( .A1(npu_inst_pe_1_5_2_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_5_2_n44), .ZN(npu_inst_pe_1_5_2_n65) );
  OAI21_X1 npu_inst_pe_1_5_2_U68 ( .B1(npu_inst_pe_1_5_2_n61), .B2(
        npu_inst_pe_1_5_2_n44), .A(npu_inst_pe_1_5_2_n65), .ZN(
        npu_inst_pe_1_5_2_n88) );
  NAND2_X1 npu_inst_pe_1_5_2_U67 ( .A1(npu_inst_pe_1_5_2_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_5_2_n40), .ZN(npu_inst_pe_1_5_2_n64) );
  OAI21_X1 npu_inst_pe_1_5_2_U66 ( .B1(npu_inst_pe_1_5_2_n63), .B2(
        npu_inst_pe_1_5_2_n40), .A(npu_inst_pe_1_5_2_n64), .ZN(
        npu_inst_pe_1_5_2_n87) );
  NAND2_X1 npu_inst_pe_1_5_2_U65 ( .A1(npu_inst_pe_1_5_2_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_5_2_n40), .ZN(npu_inst_pe_1_5_2_n62) );
  OAI21_X1 npu_inst_pe_1_5_2_U64 ( .B1(npu_inst_pe_1_5_2_n61), .B2(
        npu_inst_pe_1_5_2_n40), .A(npu_inst_pe_1_5_2_n62), .ZN(
        npu_inst_pe_1_5_2_n86) );
  AND2_X1 npu_inst_pe_1_5_2_U63 ( .A1(npu_inst_pe_1_5_2_N93), .A2(npu_inst_n55), .ZN(npu_inst_int_data_y_5__2__0_) );
  AND2_X1 npu_inst_pe_1_5_2_U62 ( .A1(npu_inst_n55), .A2(npu_inst_pe_1_5_2_N94), .ZN(npu_inst_int_data_y_5__2__1_) );
  NOR3_X1 npu_inst_pe_1_5_2_U61 ( .A1(npu_inst_pe_1_5_2_n26), .A2(npu_inst_n55), .A3(npu_inst_int_ckg[21]), .ZN(npu_inst_pe_1_5_2_n85) );
  OR2_X1 npu_inst_pe_1_5_2_U60 ( .A1(npu_inst_pe_1_5_2_n85), .A2(
        npu_inst_pe_1_5_2_n2), .ZN(npu_inst_pe_1_5_2_N84) );
  AND2_X1 npu_inst_pe_1_5_2_U59 ( .A1(npu_inst_pe_1_5_2_int_q_acc_0_), .A2(
        npu_inst_pe_1_5_2_n1), .ZN(npu_inst_int_data_res_5__2__0_) );
  AND2_X1 npu_inst_pe_1_5_2_U58 ( .A1(npu_inst_pe_1_5_2_n2), .A2(
        npu_inst_pe_1_5_2_int_q_acc_7_), .ZN(npu_inst_int_data_res_5__2__7_)
         );
  AND2_X1 npu_inst_pe_1_5_2_U57 ( .A1(npu_inst_pe_1_5_2_int_q_acc_1_), .A2(
        npu_inst_pe_1_5_2_n1), .ZN(npu_inst_int_data_res_5__2__1_) );
  AND2_X1 npu_inst_pe_1_5_2_U56 ( .A1(npu_inst_pe_1_5_2_int_q_acc_2_), .A2(
        npu_inst_pe_1_5_2_n1), .ZN(npu_inst_int_data_res_5__2__2_) );
  AND2_X1 npu_inst_pe_1_5_2_U55 ( .A1(npu_inst_pe_1_5_2_int_q_acc_3_), .A2(
        npu_inst_pe_1_5_2_n2), .ZN(npu_inst_int_data_res_5__2__3_) );
  AND2_X1 npu_inst_pe_1_5_2_U54 ( .A1(npu_inst_pe_1_5_2_int_q_acc_4_), .A2(
        npu_inst_pe_1_5_2_n2), .ZN(npu_inst_int_data_res_5__2__4_) );
  AND2_X1 npu_inst_pe_1_5_2_U53 ( .A1(npu_inst_pe_1_5_2_int_q_acc_5_), .A2(
        npu_inst_pe_1_5_2_n2), .ZN(npu_inst_int_data_res_5__2__5_) );
  AND2_X1 npu_inst_pe_1_5_2_U52 ( .A1(npu_inst_pe_1_5_2_int_q_acc_6_), .A2(
        npu_inst_pe_1_5_2_n2), .ZN(npu_inst_int_data_res_5__2__6_) );
  AOI222_X1 npu_inst_pe_1_5_2_U51 ( .A1(npu_inst_int_data_res_6__2__0_), .A2(
        npu_inst_pe_1_5_2_n1), .B1(npu_inst_pe_1_5_2_N73), .B2(
        npu_inst_pe_1_5_2_n76), .C1(npu_inst_pe_1_5_2_N65), .C2(
        npu_inst_pe_1_5_2_n77), .ZN(npu_inst_pe_1_5_2_n84) );
  INV_X1 npu_inst_pe_1_5_2_U50 ( .A(npu_inst_pe_1_5_2_n84), .ZN(
        npu_inst_pe_1_5_2_n101) );
  AOI222_X1 npu_inst_pe_1_5_2_U49 ( .A1(npu_inst_int_data_res_6__2__7_), .A2(
        npu_inst_pe_1_5_2_n1), .B1(npu_inst_pe_1_5_2_N80), .B2(
        npu_inst_pe_1_5_2_n76), .C1(npu_inst_pe_1_5_2_N72), .C2(
        npu_inst_pe_1_5_2_n77), .ZN(npu_inst_pe_1_5_2_n75) );
  INV_X1 npu_inst_pe_1_5_2_U48 ( .A(npu_inst_pe_1_5_2_n75), .ZN(
        npu_inst_pe_1_5_2_n33) );
  AOI222_X1 npu_inst_pe_1_5_2_U47 ( .A1(npu_inst_int_data_res_6__2__1_), .A2(
        npu_inst_pe_1_5_2_n1), .B1(npu_inst_pe_1_5_2_N74), .B2(
        npu_inst_pe_1_5_2_n76), .C1(npu_inst_pe_1_5_2_N66), .C2(
        npu_inst_pe_1_5_2_n77), .ZN(npu_inst_pe_1_5_2_n83) );
  INV_X1 npu_inst_pe_1_5_2_U46 ( .A(npu_inst_pe_1_5_2_n83), .ZN(
        npu_inst_pe_1_5_2_n100) );
  AOI222_X1 npu_inst_pe_1_5_2_U45 ( .A1(npu_inst_int_data_res_6__2__2_), .A2(
        npu_inst_pe_1_5_2_n1), .B1(npu_inst_pe_1_5_2_N75), .B2(
        npu_inst_pe_1_5_2_n76), .C1(npu_inst_pe_1_5_2_N67), .C2(
        npu_inst_pe_1_5_2_n77), .ZN(npu_inst_pe_1_5_2_n82) );
  INV_X1 npu_inst_pe_1_5_2_U44 ( .A(npu_inst_pe_1_5_2_n82), .ZN(
        npu_inst_pe_1_5_2_n99) );
  AOI222_X1 npu_inst_pe_1_5_2_U43 ( .A1(npu_inst_int_data_res_6__2__3_), .A2(
        npu_inst_pe_1_5_2_n1), .B1(npu_inst_pe_1_5_2_N76), .B2(
        npu_inst_pe_1_5_2_n76), .C1(npu_inst_pe_1_5_2_N68), .C2(
        npu_inst_pe_1_5_2_n77), .ZN(npu_inst_pe_1_5_2_n81) );
  INV_X1 npu_inst_pe_1_5_2_U42 ( .A(npu_inst_pe_1_5_2_n81), .ZN(
        npu_inst_pe_1_5_2_n98) );
  AOI222_X1 npu_inst_pe_1_5_2_U41 ( .A1(npu_inst_int_data_res_6__2__4_), .A2(
        npu_inst_pe_1_5_2_n1), .B1(npu_inst_pe_1_5_2_N77), .B2(
        npu_inst_pe_1_5_2_n76), .C1(npu_inst_pe_1_5_2_N69), .C2(
        npu_inst_pe_1_5_2_n77), .ZN(npu_inst_pe_1_5_2_n80) );
  INV_X1 npu_inst_pe_1_5_2_U40 ( .A(npu_inst_pe_1_5_2_n80), .ZN(
        npu_inst_pe_1_5_2_n36) );
  AOI222_X1 npu_inst_pe_1_5_2_U39 ( .A1(npu_inst_int_data_res_6__2__5_), .A2(
        npu_inst_pe_1_5_2_n1), .B1(npu_inst_pe_1_5_2_N78), .B2(
        npu_inst_pe_1_5_2_n76), .C1(npu_inst_pe_1_5_2_N70), .C2(
        npu_inst_pe_1_5_2_n77), .ZN(npu_inst_pe_1_5_2_n79) );
  INV_X1 npu_inst_pe_1_5_2_U38 ( .A(npu_inst_pe_1_5_2_n79), .ZN(
        npu_inst_pe_1_5_2_n35) );
  AOI222_X1 npu_inst_pe_1_5_2_U37 ( .A1(npu_inst_int_data_res_6__2__6_), .A2(
        npu_inst_pe_1_5_2_n1), .B1(npu_inst_pe_1_5_2_N79), .B2(
        npu_inst_pe_1_5_2_n76), .C1(npu_inst_pe_1_5_2_N71), .C2(
        npu_inst_pe_1_5_2_n77), .ZN(npu_inst_pe_1_5_2_n78) );
  INV_X1 npu_inst_pe_1_5_2_U36 ( .A(npu_inst_pe_1_5_2_n78), .ZN(
        npu_inst_pe_1_5_2_n34) );
  INV_X1 npu_inst_pe_1_5_2_U35 ( .A(npu_inst_pe_1_5_2_int_data_1_), .ZN(
        npu_inst_pe_1_5_2_n14) );
  AND2_X1 npu_inst_pe_1_5_2_U34 ( .A1(npu_inst_int_data_x_5__2__1_), .A2(
        npu_inst_pe_1_5_2_int_q_weight_1_), .ZN(npu_inst_pe_1_5_2_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_5_2_U33 ( .A1(npu_inst_int_data_x_5__2__0_), .A2(
        npu_inst_pe_1_5_2_int_q_weight_1_), .ZN(npu_inst_pe_1_5_2_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_5_2_U32 ( .A1(npu_inst_n55), .A2(
        npu_inst_int_data_y_6__2__1_), .B1(npu_inst_pe_1_5_2_n3), .B2(
        npu_inst_int_data_x_5__3__1_), .ZN(npu_inst_pe_1_5_2_n63) );
  AOI22_X1 npu_inst_pe_1_5_2_U31 ( .A1(npu_inst_n55), .A2(
        npu_inst_int_data_y_6__2__0_), .B1(npu_inst_pe_1_5_2_n3), .B2(
        npu_inst_int_data_x_5__3__0_), .ZN(npu_inst_pe_1_5_2_n61) );
  INV_X1 npu_inst_pe_1_5_2_U30 ( .A(npu_inst_pe_1_5_2_int_data_0_), .ZN(
        npu_inst_pe_1_5_2_n13) );
  INV_X1 npu_inst_pe_1_5_2_U29 ( .A(npu_inst_n68), .ZN(npu_inst_pe_1_5_2_n5)
         );
  OR3_X1 npu_inst_pe_1_5_2_U28 ( .A1(npu_inst_pe_1_5_2_n6), .A2(
        npu_inst_pe_1_5_2_n8), .A3(npu_inst_pe_1_5_2_n5), .ZN(
        npu_inst_pe_1_5_2_n56) );
  OR3_X1 npu_inst_pe_1_5_2_U27 ( .A1(npu_inst_pe_1_5_2_n5), .A2(
        npu_inst_pe_1_5_2_n8), .A3(npu_inst_pe_1_5_2_n7), .ZN(
        npu_inst_pe_1_5_2_n48) );
  INV_X1 npu_inst_pe_1_5_2_U26 ( .A(npu_inst_pe_1_5_2_n5), .ZN(
        npu_inst_pe_1_5_2_n4) );
  INV_X1 npu_inst_pe_1_5_2_U25 ( .A(npu_inst_n123), .ZN(npu_inst_pe_1_5_2_n12)
         );
  OR3_X1 npu_inst_pe_1_5_2_U24 ( .A1(npu_inst_pe_1_5_2_n4), .A2(
        npu_inst_pe_1_5_2_n8), .A3(npu_inst_pe_1_5_2_n7), .ZN(
        npu_inst_pe_1_5_2_n52) );
  OR3_X1 npu_inst_pe_1_5_2_U23 ( .A1(npu_inst_pe_1_5_2_n6), .A2(
        npu_inst_pe_1_5_2_n8), .A3(npu_inst_pe_1_5_2_n4), .ZN(
        npu_inst_pe_1_5_2_n60) );
  NOR2_X1 npu_inst_pe_1_5_2_U22 ( .A1(npu_inst_pe_1_5_2_n60), .A2(
        npu_inst_pe_1_5_2_n3), .ZN(npu_inst_pe_1_5_2_n58) );
  NOR2_X1 npu_inst_pe_1_5_2_U21 ( .A1(npu_inst_pe_1_5_2_n56), .A2(
        npu_inst_pe_1_5_2_n3), .ZN(npu_inst_pe_1_5_2_n54) );
  NOR2_X1 npu_inst_pe_1_5_2_U20 ( .A1(npu_inst_pe_1_5_2_n52), .A2(
        npu_inst_pe_1_5_2_n3), .ZN(npu_inst_pe_1_5_2_n50) );
  NOR2_X1 npu_inst_pe_1_5_2_U19 ( .A1(npu_inst_pe_1_5_2_n48), .A2(
        npu_inst_pe_1_5_2_n3), .ZN(npu_inst_pe_1_5_2_n46) );
  NOR2_X1 npu_inst_pe_1_5_2_U18 ( .A1(npu_inst_pe_1_5_2_n40), .A2(
        npu_inst_pe_1_5_2_n3), .ZN(npu_inst_pe_1_5_2_n38) );
  NOR2_X1 npu_inst_pe_1_5_2_U17 ( .A1(npu_inst_pe_1_5_2_n44), .A2(
        npu_inst_pe_1_5_2_n3), .ZN(npu_inst_pe_1_5_2_n42) );
  BUF_X1 npu_inst_pe_1_5_2_U16 ( .A(npu_inst_n97), .Z(npu_inst_pe_1_5_2_n8) );
  BUF_X1 npu_inst_pe_1_5_2_U15 ( .A(npu_inst_pe_1_5_2_n12), .Z(
        npu_inst_pe_1_5_2_n11) );
  BUF_X1 npu_inst_pe_1_5_2_U14 ( .A(npu_inst_pe_1_5_2_n12), .Z(
        npu_inst_pe_1_5_2_n10) );
  BUF_X1 npu_inst_pe_1_5_2_U13 ( .A(npu_inst_pe_1_5_2_n12), .Z(
        npu_inst_pe_1_5_2_n9) );
  INV_X1 npu_inst_pe_1_5_2_U12 ( .A(npu_inst_pe_1_5_2_n38), .ZN(
        npu_inst_pe_1_5_2_n118) );
  INV_X1 npu_inst_pe_1_5_2_U11 ( .A(npu_inst_pe_1_5_2_n58), .ZN(
        npu_inst_pe_1_5_2_n114) );
  INV_X1 npu_inst_pe_1_5_2_U10 ( .A(npu_inst_pe_1_5_2_n54), .ZN(
        npu_inst_pe_1_5_2_n115) );
  INV_X1 npu_inst_pe_1_5_2_U9 ( .A(npu_inst_pe_1_5_2_n50), .ZN(
        npu_inst_pe_1_5_2_n116) );
  INV_X1 npu_inst_pe_1_5_2_U8 ( .A(npu_inst_pe_1_5_2_n46), .ZN(
        npu_inst_pe_1_5_2_n117) );
  INV_X1 npu_inst_pe_1_5_2_U7 ( .A(npu_inst_pe_1_5_2_n42), .ZN(
        npu_inst_pe_1_5_2_n119) );
  BUF_X1 npu_inst_pe_1_5_2_U6 ( .A(npu_inst_n17), .Z(npu_inst_pe_1_5_2_n2) );
  BUF_X1 npu_inst_pe_1_5_2_U5 ( .A(npu_inst_n17), .Z(npu_inst_pe_1_5_2_n1) );
  NOR2_X1 npu_inst_pe_1_5_2_U4 ( .A1(npu_inst_pe_1_5_2_int_q_weight_0_), .A2(
        npu_inst_pe_1_5_2_n1), .ZN(npu_inst_pe_1_5_2_n76) );
  NOR2_X1 npu_inst_pe_1_5_2_U3 ( .A1(npu_inst_pe_1_5_2_n27), .A2(
        npu_inst_pe_1_5_2_n1), .ZN(npu_inst_pe_1_5_2_n77) );
  FA_X1 npu_inst_pe_1_5_2_sub_77_U2_1 ( .A(npu_inst_pe_1_5_2_int_q_acc_1_), 
        .B(npu_inst_pe_1_5_2_n14), .CI(npu_inst_pe_1_5_2_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_5_2_sub_77_carry_2_), .S(npu_inst_pe_1_5_2_N66) );
  FA_X1 npu_inst_pe_1_5_2_add_79_U1_1 ( .A(npu_inst_pe_1_5_2_int_q_acc_1_), 
        .B(npu_inst_pe_1_5_2_int_data_1_), .CI(
        npu_inst_pe_1_5_2_add_79_carry_1_), .CO(
        npu_inst_pe_1_5_2_add_79_carry_2_), .S(npu_inst_pe_1_5_2_N74) );
  NAND3_X1 npu_inst_pe_1_5_2_U109 ( .A1(npu_inst_pe_1_5_2_n5), .A2(
        npu_inst_pe_1_5_2_n7), .A3(npu_inst_pe_1_5_2_n8), .ZN(
        npu_inst_pe_1_5_2_n44) );
  NAND3_X1 npu_inst_pe_1_5_2_U108 ( .A1(npu_inst_pe_1_5_2_n4), .A2(
        npu_inst_pe_1_5_2_n7), .A3(npu_inst_pe_1_5_2_n8), .ZN(
        npu_inst_pe_1_5_2_n40) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_5_2_n34), .CK(
        npu_inst_pe_1_5_2_net3327), .RN(npu_inst_pe_1_5_2_n9), .Q(
        npu_inst_pe_1_5_2_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_5_2_n35), .CK(
        npu_inst_pe_1_5_2_net3327), .RN(npu_inst_pe_1_5_2_n9), .Q(
        npu_inst_pe_1_5_2_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_5_2_n36), .CK(
        npu_inst_pe_1_5_2_net3327), .RN(npu_inst_pe_1_5_2_n9), .Q(
        npu_inst_pe_1_5_2_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_5_2_n98), .CK(
        npu_inst_pe_1_5_2_net3327), .RN(npu_inst_pe_1_5_2_n9), .Q(
        npu_inst_pe_1_5_2_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_5_2_n99), .CK(
        npu_inst_pe_1_5_2_net3327), .RN(npu_inst_pe_1_5_2_n9), .Q(
        npu_inst_pe_1_5_2_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_5_2_n100), 
        .CK(npu_inst_pe_1_5_2_net3327), .RN(npu_inst_pe_1_5_2_n9), .Q(
        npu_inst_pe_1_5_2_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_5_2_n33), .CK(
        npu_inst_pe_1_5_2_net3327), .RN(npu_inst_pe_1_5_2_n9), .Q(
        npu_inst_pe_1_5_2_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_5_2_n101), 
        .CK(npu_inst_pe_1_5_2_net3327), .RN(npu_inst_pe_1_5_2_n9), .Q(
        npu_inst_pe_1_5_2_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_weight_reg_0_ ( .D(npu_inst_n109), .CK(
        npu_inst_pe_1_5_2_net3333), .RN(npu_inst_pe_1_5_2_n9), .Q(
        npu_inst_pe_1_5_2_int_q_weight_0_), .QN(npu_inst_pe_1_5_2_n27) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_weight_reg_1_ ( .D(npu_inst_n115), .CK(
        npu_inst_pe_1_5_2_net3333), .RN(npu_inst_pe_1_5_2_n9), .Q(
        npu_inst_pe_1_5_2_int_q_weight_1_), .QN(npu_inst_pe_1_5_2_n26) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_5_2_n113), 
        .CK(npu_inst_pe_1_5_2_net3333), .RN(npu_inst_pe_1_5_2_n9), .Q(
        npu_inst_pe_1_5_2_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_5_2_n107), 
        .CK(npu_inst_pe_1_5_2_net3333), .RN(npu_inst_pe_1_5_2_n9), .Q(
        npu_inst_pe_1_5_2_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_5_2_n112), 
        .CK(npu_inst_pe_1_5_2_net3333), .RN(npu_inst_pe_1_5_2_n10), .Q(
        npu_inst_pe_1_5_2_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_5_2_n106), 
        .CK(npu_inst_pe_1_5_2_net3333), .RN(npu_inst_pe_1_5_2_n10), .Q(
        npu_inst_pe_1_5_2_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_5_2_n111), 
        .CK(npu_inst_pe_1_5_2_net3333), .RN(npu_inst_pe_1_5_2_n10), .Q(
        npu_inst_pe_1_5_2_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_5_2_n105), 
        .CK(npu_inst_pe_1_5_2_net3333), .RN(npu_inst_pe_1_5_2_n10), .Q(
        npu_inst_pe_1_5_2_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_5_2_n110), 
        .CK(npu_inst_pe_1_5_2_net3333), .RN(npu_inst_pe_1_5_2_n10), .Q(
        npu_inst_pe_1_5_2_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_5_2_n104), 
        .CK(npu_inst_pe_1_5_2_net3333), .RN(npu_inst_pe_1_5_2_n10), .Q(
        npu_inst_pe_1_5_2_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_5_2_n109), 
        .CK(npu_inst_pe_1_5_2_net3333), .RN(npu_inst_pe_1_5_2_n10), .Q(
        npu_inst_pe_1_5_2_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_5_2_n103), 
        .CK(npu_inst_pe_1_5_2_net3333), .RN(npu_inst_pe_1_5_2_n10), .Q(
        npu_inst_pe_1_5_2_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_5_2_n108), 
        .CK(npu_inst_pe_1_5_2_net3333), .RN(npu_inst_pe_1_5_2_n10), .Q(
        npu_inst_pe_1_5_2_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_5_2_n102), 
        .CK(npu_inst_pe_1_5_2_net3333), .RN(npu_inst_pe_1_5_2_n10), .Q(
        npu_inst_pe_1_5_2_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_5_2_n86), 
        .CK(npu_inst_pe_1_5_2_net3333), .RN(npu_inst_pe_1_5_2_n10), .Q(
        npu_inst_pe_1_5_2_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_5_2_n87), 
        .CK(npu_inst_pe_1_5_2_net3333), .RN(npu_inst_pe_1_5_2_n10), .Q(
        npu_inst_pe_1_5_2_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_5_2_n88), 
        .CK(npu_inst_pe_1_5_2_net3333), .RN(npu_inst_pe_1_5_2_n11), .Q(
        npu_inst_pe_1_5_2_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_5_2_n89), 
        .CK(npu_inst_pe_1_5_2_net3333), .RN(npu_inst_pe_1_5_2_n11), .Q(
        npu_inst_pe_1_5_2_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_5_2_n90), 
        .CK(npu_inst_pe_1_5_2_net3333), .RN(npu_inst_pe_1_5_2_n11), .Q(
        npu_inst_pe_1_5_2_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_5_2_n91), 
        .CK(npu_inst_pe_1_5_2_net3333), .RN(npu_inst_pe_1_5_2_n11), .Q(
        npu_inst_pe_1_5_2_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_5_2_n92), 
        .CK(npu_inst_pe_1_5_2_net3333), .RN(npu_inst_pe_1_5_2_n11), .Q(
        npu_inst_pe_1_5_2_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_5_2_n93), 
        .CK(npu_inst_pe_1_5_2_net3333), .RN(npu_inst_pe_1_5_2_n11), .Q(
        npu_inst_pe_1_5_2_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_5_2_n94), 
        .CK(npu_inst_pe_1_5_2_net3333), .RN(npu_inst_pe_1_5_2_n11), .Q(
        npu_inst_pe_1_5_2_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_5_2_n95), 
        .CK(npu_inst_pe_1_5_2_net3333), .RN(npu_inst_pe_1_5_2_n11), .Q(
        npu_inst_pe_1_5_2_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_5_2_n96), 
        .CK(npu_inst_pe_1_5_2_net3333), .RN(npu_inst_pe_1_5_2_n11), .Q(
        npu_inst_pe_1_5_2_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_5_2_n97), 
        .CK(npu_inst_pe_1_5_2_net3333), .RN(npu_inst_pe_1_5_2_n11), .Q(
        npu_inst_pe_1_5_2_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_5_2_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_5_2_N84), .SE(1'b0), .GCK(npu_inst_pe_1_5_2_net3327) );
  CLKGATETST_X1 npu_inst_pe_1_5_2_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n62), .SE(1'b0), .GCK(npu_inst_pe_1_5_2_net3333) );
  MUX2_X1 npu_inst_pe_1_5_3_U162 ( .A(npu_inst_pe_1_5_3_n32), .B(
        npu_inst_pe_1_5_3_n29), .S(npu_inst_pe_1_5_3_n8), .Z(
        npu_inst_pe_1_5_3_N93) );
  MUX2_X1 npu_inst_pe_1_5_3_U161 ( .A(npu_inst_pe_1_5_3_n31), .B(
        npu_inst_pe_1_5_3_n30), .S(npu_inst_pe_1_5_3_n6), .Z(
        npu_inst_pe_1_5_3_n32) );
  MUX2_X1 npu_inst_pe_1_5_3_U160 ( .A(npu_inst_pe_1_5_3_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_5_3_int_q_reg_v_1__0_), .S(npu_inst_pe_1_5_3_n4), .Z(
        npu_inst_pe_1_5_3_n31) );
  MUX2_X1 npu_inst_pe_1_5_3_U159 ( .A(npu_inst_pe_1_5_3_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_5_3_int_q_reg_v_3__0_), .S(npu_inst_pe_1_5_3_n4), .Z(
        npu_inst_pe_1_5_3_n30) );
  MUX2_X1 npu_inst_pe_1_5_3_U158 ( .A(npu_inst_pe_1_5_3_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_5_3_int_q_reg_v_5__0_), .S(npu_inst_pe_1_5_3_n4), .Z(
        npu_inst_pe_1_5_3_n29) );
  MUX2_X1 npu_inst_pe_1_5_3_U157 ( .A(npu_inst_pe_1_5_3_n28), .B(
        npu_inst_pe_1_5_3_n23), .S(npu_inst_pe_1_5_3_n8), .Z(
        npu_inst_pe_1_5_3_N94) );
  MUX2_X1 npu_inst_pe_1_5_3_U156 ( .A(npu_inst_pe_1_5_3_n25), .B(
        npu_inst_pe_1_5_3_n24), .S(npu_inst_pe_1_5_3_n6), .Z(
        npu_inst_pe_1_5_3_n28) );
  MUX2_X1 npu_inst_pe_1_5_3_U155 ( .A(npu_inst_pe_1_5_3_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_5_3_int_q_reg_v_1__1_), .S(npu_inst_pe_1_5_3_n4), .Z(
        npu_inst_pe_1_5_3_n25) );
  MUX2_X1 npu_inst_pe_1_5_3_U154 ( .A(npu_inst_pe_1_5_3_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_5_3_int_q_reg_v_3__1_), .S(npu_inst_pe_1_5_3_n4), .Z(
        npu_inst_pe_1_5_3_n24) );
  MUX2_X1 npu_inst_pe_1_5_3_U153 ( .A(npu_inst_pe_1_5_3_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_5_3_int_q_reg_v_5__1_), .S(npu_inst_pe_1_5_3_n4), .Z(
        npu_inst_pe_1_5_3_n23) );
  MUX2_X1 npu_inst_pe_1_5_3_U152 ( .A(npu_inst_pe_1_5_3_n22), .B(
        npu_inst_pe_1_5_3_n19), .S(npu_inst_pe_1_5_3_n8), .Z(
        npu_inst_int_data_x_5__3__1_) );
  MUX2_X1 npu_inst_pe_1_5_3_U151 ( .A(npu_inst_pe_1_5_3_n21), .B(
        npu_inst_pe_1_5_3_n20), .S(npu_inst_pe_1_5_3_n6), .Z(
        npu_inst_pe_1_5_3_n22) );
  MUX2_X1 npu_inst_pe_1_5_3_U150 ( .A(npu_inst_pe_1_5_3_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_5_3_int_q_reg_h_1__1_), .S(npu_inst_pe_1_5_3_n4), .Z(
        npu_inst_pe_1_5_3_n21) );
  MUX2_X1 npu_inst_pe_1_5_3_U149 ( .A(npu_inst_pe_1_5_3_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_5_3_int_q_reg_h_3__1_), .S(npu_inst_pe_1_5_3_n4), .Z(
        npu_inst_pe_1_5_3_n20) );
  MUX2_X1 npu_inst_pe_1_5_3_U148 ( .A(npu_inst_pe_1_5_3_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_5_3_int_q_reg_h_5__1_), .S(npu_inst_pe_1_5_3_n4), .Z(
        npu_inst_pe_1_5_3_n19) );
  MUX2_X1 npu_inst_pe_1_5_3_U147 ( .A(npu_inst_pe_1_5_3_n18), .B(
        npu_inst_pe_1_5_3_n15), .S(npu_inst_pe_1_5_3_n8), .Z(
        npu_inst_int_data_x_5__3__0_) );
  MUX2_X1 npu_inst_pe_1_5_3_U146 ( .A(npu_inst_pe_1_5_3_n17), .B(
        npu_inst_pe_1_5_3_n16), .S(npu_inst_pe_1_5_3_n6), .Z(
        npu_inst_pe_1_5_3_n18) );
  MUX2_X1 npu_inst_pe_1_5_3_U145 ( .A(npu_inst_pe_1_5_3_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_5_3_int_q_reg_h_1__0_), .S(npu_inst_pe_1_5_3_n4), .Z(
        npu_inst_pe_1_5_3_n17) );
  MUX2_X1 npu_inst_pe_1_5_3_U144 ( .A(npu_inst_pe_1_5_3_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_5_3_int_q_reg_h_3__0_), .S(npu_inst_pe_1_5_3_n4), .Z(
        npu_inst_pe_1_5_3_n16) );
  MUX2_X1 npu_inst_pe_1_5_3_U143 ( .A(npu_inst_pe_1_5_3_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_5_3_int_q_reg_h_5__0_), .S(npu_inst_pe_1_5_3_n4), .Z(
        npu_inst_pe_1_5_3_n15) );
  XOR2_X1 npu_inst_pe_1_5_3_U142 ( .A(npu_inst_pe_1_5_3_int_data_0_), .B(
        npu_inst_pe_1_5_3_int_q_acc_0_), .Z(npu_inst_pe_1_5_3_N73) );
  AND2_X1 npu_inst_pe_1_5_3_U141 ( .A1(npu_inst_pe_1_5_3_int_q_acc_0_), .A2(
        npu_inst_pe_1_5_3_int_data_0_), .ZN(npu_inst_pe_1_5_3_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_5_3_U140 ( .A(npu_inst_pe_1_5_3_int_q_acc_0_), .B(
        npu_inst_pe_1_5_3_n13), .ZN(npu_inst_pe_1_5_3_N65) );
  OR2_X1 npu_inst_pe_1_5_3_U139 ( .A1(npu_inst_pe_1_5_3_n13), .A2(
        npu_inst_pe_1_5_3_int_q_acc_0_), .ZN(npu_inst_pe_1_5_3_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_5_3_U138 ( .A(npu_inst_pe_1_5_3_int_q_acc_2_), .B(
        npu_inst_pe_1_5_3_add_79_carry_2_), .Z(npu_inst_pe_1_5_3_N75) );
  AND2_X1 npu_inst_pe_1_5_3_U137 ( .A1(npu_inst_pe_1_5_3_add_79_carry_2_), 
        .A2(npu_inst_pe_1_5_3_int_q_acc_2_), .ZN(
        npu_inst_pe_1_5_3_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_5_3_U136 ( .A(npu_inst_pe_1_5_3_int_q_acc_3_), .B(
        npu_inst_pe_1_5_3_add_79_carry_3_), .Z(npu_inst_pe_1_5_3_N76) );
  AND2_X1 npu_inst_pe_1_5_3_U135 ( .A1(npu_inst_pe_1_5_3_add_79_carry_3_), 
        .A2(npu_inst_pe_1_5_3_int_q_acc_3_), .ZN(
        npu_inst_pe_1_5_3_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_5_3_U134 ( .A(npu_inst_pe_1_5_3_int_q_acc_4_), .B(
        npu_inst_pe_1_5_3_add_79_carry_4_), .Z(npu_inst_pe_1_5_3_N77) );
  AND2_X1 npu_inst_pe_1_5_3_U133 ( .A1(npu_inst_pe_1_5_3_add_79_carry_4_), 
        .A2(npu_inst_pe_1_5_3_int_q_acc_4_), .ZN(
        npu_inst_pe_1_5_3_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_5_3_U132 ( .A(npu_inst_pe_1_5_3_int_q_acc_5_), .B(
        npu_inst_pe_1_5_3_add_79_carry_5_), .Z(npu_inst_pe_1_5_3_N78) );
  AND2_X1 npu_inst_pe_1_5_3_U131 ( .A1(npu_inst_pe_1_5_3_add_79_carry_5_), 
        .A2(npu_inst_pe_1_5_3_int_q_acc_5_), .ZN(
        npu_inst_pe_1_5_3_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_5_3_U130 ( .A(npu_inst_pe_1_5_3_int_q_acc_6_), .B(
        npu_inst_pe_1_5_3_add_79_carry_6_), .Z(npu_inst_pe_1_5_3_N79) );
  AND2_X1 npu_inst_pe_1_5_3_U129 ( .A1(npu_inst_pe_1_5_3_add_79_carry_6_), 
        .A2(npu_inst_pe_1_5_3_int_q_acc_6_), .ZN(
        npu_inst_pe_1_5_3_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_5_3_U128 ( .A(npu_inst_pe_1_5_3_int_q_acc_7_), .B(
        npu_inst_pe_1_5_3_add_79_carry_7_), .Z(npu_inst_pe_1_5_3_N80) );
  XNOR2_X1 npu_inst_pe_1_5_3_U127 ( .A(npu_inst_pe_1_5_3_sub_77_carry_2_), .B(
        npu_inst_pe_1_5_3_int_q_acc_2_), .ZN(npu_inst_pe_1_5_3_N67) );
  OR2_X1 npu_inst_pe_1_5_3_U126 ( .A1(npu_inst_pe_1_5_3_int_q_acc_2_), .A2(
        npu_inst_pe_1_5_3_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_5_3_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_5_3_U125 ( .A(npu_inst_pe_1_5_3_sub_77_carry_3_), .B(
        npu_inst_pe_1_5_3_int_q_acc_3_), .ZN(npu_inst_pe_1_5_3_N68) );
  OR2_X1 npu_inst_pe_1_5_3_U124 ( .A1(npu_inst_pe_1_5_3_int_q_acc_3_), .A2(
        npu_inst_pe_1_5_3_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_5_3_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_5_3_U123 ( .A(npu_inst_pe_1_5_3_sub_77_carry_4_), .B(
        npu_inst_pe_1_5_3_int_q_acc_4_), .ZN(npu_inst_pe_1_5_3_N69) );
  OR2_X1 npu_inst_pe_1_5_3_U122 ( .A1(npu_inst_pe_1_5_3_int_q_acc_4_), .A2(
        npu_inst_pe_1_5_3_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_5_3_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_5_3_U121 ( .A(npu_inst_pe_1_5_3_sub_77_carry_5_), .B(
        npu_inst_pe_1_5_3_int_q_acc_5_), .ZN(npu_inst_pe_1_5_3_N70) );
  OR2_X1 npu_inst_pe_1_5_3_U120 ( .A1(npu_inst_pe_1_5_3_int_q_acc_5_), .A2(
        npu_inst_pe_1_5_3_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_5_3_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_5_3_U119 ( .A(npu_inst_pe_1_5_3_sub_77_carry_6_), .B(
        npu_inst_pe_1_5_3_int_q_acc_6_), .ZN(npu_inst_pe_1_5_3_N71) );
  OR2_X1 npu_inst_pe_1_5_3_U118 ( .A1(npu_inst_pe_1_5_3_int_q_acc_6_), .A2(
        npu_inst_pe_1_5_3_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_5_3_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_5_3_U117 ( .A(npu_inst_pe_1_5_3_int_q_acc_7_), .B(
        npu_inst_pe_1_5_3_sub_77_carry_7_), .ZN(npu_inst_pe_1_5_3_N72) );
  INV_X1 npu_inst_pe_1_5_3_U116 ( .A(npu_inst_n76), .ZN(npu_inst_pe_1_5_3_n7)
         );
  INV_X1 npu_inst_pe_1_5_3_U115 ( .A(npu_inst_pe_1_5_3_n7), .ZN(
        npu_inst_pe_1_5_3_n6) );
  INV_X1 npu_inst_pe_1_5_3_U114 ( .A(npu_inst_n54), .ZN(npu_inst_pe_1_5_3_n3)
         );
  AOI22_X1 npu_inst_pe_1_5_3_U113 ( .A1(npu_inst_int_data_y_6__3__0_), .A2(
        npu_inst_pe_1_5_3_n58), .B1(npu_inst_pe_1_5_3_n114), .B2(
        npu_inst_pe_1_5_3_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_5_3_n57) );
  INV_X1 npu_inst_pe_1_5_3_U112 ( .A(npu_inst_pe_1_5_3_n57), .ZN(
        npu_inst_pe_1_5_3_n108) );
  AOI22_X1 npu_inst_pe_1_5_3_U111 ( .A1(npu_inst_int_data_y_6__3__0_), .A2(
        npu_inst_pe_1_5_3_n54), .B1(npu_inst_pe_1_5_3_n115), .B2(
        npu_inst_pe_1_5_3_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_5_3_n53) );
  INV_X1 npu_inst_pe_1_5_3_U110 ( .A(npu_inst_pe_1_5_3_n53), .ZN(
        npu_inst_pe_1_5_3_n109) );
  AOI22_X1 npu_inst_pe_1_5_3_U107 ( .A1(npu_inst_int_data_y_6__3__0_), .A2(
        npu_inst_pe_1_5_3_n50), .B1(npu_inst_pe_1_5_3_n116), .B2(
        npu_inst_pe_1_5_3_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_5_3_n49) );
  INV_X1 npu_inst_pe_1_5_3_U106 ( .A(npu_inst_pe_1_5_3_n49), .ZN(
        npu_inst_pe_1_5_3_n110) );
  AOI22_X1 npu_inst_pe_1_5_3_U105 ( .A1(npu_inst_int_data_y_6__3__0_), .A2(
        npu_inst_pe_1_5_3_n46), .B1(npu_inst_pe_1_5_3_n117), .B2(
        npu_inst_pe_1_5_3_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_5_3_n45) );
  INV_X1 npu_inst_pe_1_5_3_U104 ( .A(npu_inst_pe_1_5_3_n45), .ZN(
        npu_inst_pe_1_5_3_n111) );
  AOI22_X1 npu_inst_pe_1_5_3_U103 ( .A1(npu_inst_int_data_y_6__3__0_), .A2(
        npu_inst_pe_1_5_3_n42), .B1(npu_inst_pe_1_5_3_n119), .B2(
        npu_inst_pe_1_5_3_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_5_3_n41) );
  INV_X1 npu_inst_pe_1_5_3_U102 ( .A(npu_inst_pe_1_5_3_n41), .ZN(
        npu_inst_pe_1_5_3_n112) );
  AOI22_X1 npu_inst_pe_1_5_3_U101 ( .A1(npu_inst_int_data_y_6__3__1_), .A2(
        npu_inst_pe_1_5_3_n58), .B1(npu_inst_pe_1_5_3_n114), .B2(
        npu_inst_pe_1_5_3_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_5_3_n59) );
  INV_X1 npu_inst_pe_1_5_3_U100 ( .A(npu_inst_pe_1_5_3_n59), .ZN(
        npu_inst_pe_1_5_3_n102) );
  AOI22_X1 npu_inst_pe_1_5_3_U99 ( .A1(npu_inst_int_data_y_6__3__1_), .A2(
        npu_inst_pe_1_5_3_n54), .B1(npu_inst_pe_1_5_3_n115), .B2(
        npu_inst_pe_1_5_3_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_5_3_n55) );
  INV_X1 npu_inst_pe_1_5_3_U98 ( .A(npu_inst_pe_1_5_3_n55), .ZN(
        npu_inst_pe_1_5_3_n103) );
  AOI22_X1 npu_inst_pe_1_5_3_U97 ( .A1(npu_inst_int_data_y_6__3__1_), .A2(
        npu_inst_pe_1_5_3_n50), .B1(npu_inst_pe_1_5_3_n116), .B2(
        npu_inst_pe_1_5_3_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_5_3_n51) );
  INV_X1 npu_inst_pe_1_5_3_U96 ( .A(npu_inst_pe_1_5_3_n51), .ZN(
        npu_inst_pe_1_5_3_n104) );
  AOI22_X1 npu_inst_pe_1_5_3_U95 ( .A1(npu_inst_int_data_y_6__3__1_), .A2(
        npu_inst_pe_1_5_3_n46), .B1(npu_inst_pe_1_5_3_n117), .B2(
        npu_inst_pe_1_5_3_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_5_3_n47) );
  INV_X1 npu_inst_pe_1_5_3_U94 ( .A(npu_inst_pe_1_5_3_n47), .ZN(
        npu_inst_pe_1_5_3_n105) );
  AOI22_X1 npu_inst_pe_1_5_3_U93 ( .A1(npu_inst_int_data_y_6__3__1_), .A2(
        npu_inst_pe_1_5_3_n42), .B1(npu_inst_pe_1_5_3_n119), .B2(
        npu_inst_pe_1_5_3_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_5_3_n43) );
  INV_X1 npu_inst_pe_1_5_3_U92 ( .A(npu_inst_pe_1_5_3_n43), .ZN(
        npu_inst_pe_1_5_3_n106) );
  AOI22_X1 npu_inst_pe_1_5_3_U91 ( .A1(npu_inst_pe_1_5_3_n38), .A2(
        npu_inst_int_data_y_6__3__1_), .B1(npu_inst_pe_1_5_3_n118), .B2(
        npu_inst_pe_1_5_3_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_5_3_n39) );
  INV_X1 npu_inst_pe_1_5_3_U90 ( .A(npu_inst_pe_1_5_3_n39), .ZN(
        npu_inst_pe_1_5_3_n107) );
  AOI22_X1 npu_inst_pe_1_5_3_U89 ( .A1(npu_inst_pe_1_5_3_n38), .A2(
        npu_inst_int_data_y_6__3__0_), .B1(npu_inst_pe_1_5_3_n118), .B2(
        npu_inst_pe_1_5_3_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_5_3_n37) );
  INV_X1 npu_inst_pe_1_5_3_U88 ( .A(npu_inst_pe_1_5_3_n37), .ZN(
        npu_inst_pe_1_5_3_n113) );
  NAND2_X1 npu_inst_pe_1_5_3_U87 ( .A1(npu_inst_pe_1_5_3_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_5_3_n60), .ZN(npu_inst_pe_1_5_3_n74) );
  OAI21_X1 npu_inst_pe_1_5_3_U86 ( .B1(npu_inst_pe_1_5_3_n63), .B2(
        npu_inst_pe_1_5_3_n60), .A(npu_inst_pe_1_5_3_n74), .ZN(
        npu_inst_pe_1_5_3_n97) );
  NAND2_X1 npu_inst_pe_1_5_3_U85 ( .A1(npu_inst_pe_1_5_3_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_5_3_n60), .ZN(npu_inst_pe_1_5_3_n73) );
  OAI21_X1 npu_inst_pe_1_5_3_U84 ( .B1(npu_inst_pe_1_5_3_n61), .B2(
        npu_inst_pe_1_5_3_n60), .A(npu_inst_pe_1_5_3_n73), .ZN(
        npu_inst_pe_1_5_3_n96) );
  NAND2_X1 npu_inst_pe_1_5_3_U83 ( .A1(npu_inst_pe_1_5_3_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_5_3_n56), .ZN(npu_inst_pe_1_5_3_n72) );
  OAI21_X1 npu_inst_pe_1_5_3_U82 ( .B1(npu_inst_pe_1_5_3_n63), .B2(
        npu_inst_pe_1_5_3_n56), .A(npu_inst_pe_1_5_3_n72), .ZN(
        npu_inst_pe_1_5_3_n95) );
  NAND2_X1 npu_inst_pe_1_5_3_U81 ( .A1(npu_inst_pe_1_5_3_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_5_3_n56), .ZN(npu_inst_pe_1_5_3_n71) );
  OAI21_X1 npu_inst_pe_1_5_3_U80 ( .B1(npu_inst_pe_1_5_3_n61), .B2(
        npu_inst_pe_1_5_3_n56), .A(npu_inst_pe_1_5_3_n71), .ZN(
        npu_inst_pe_1_5_3_n94) );
  NAND2_X1 npu_inst_pe_1_5_3_U79 ( .A1(npu_inst_pe_1_5_3_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_5_3_n52), .ZN(npu_inst_pe_1_5_3_n70) );
  OAI21_X1 npu_inst_pe_1_5_3_U78 ( .B1(npu_inst_pe_1_5_3_n63), .B2(
        npu_inst_pe_1_5_3_n52), .A(npu_inst_pe_1_5_3_n70), .ZN(
        npu_inst_pe_1_5_3_n93) );
  NAND2_X1 npu_inst_pe_1_5_3_U77 ( .A1(npu_inst_pe_1_5_3_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_5_3_n52), .ZN(npu_inst_pe_1_5_3_n69) );
  OAI21_X1 npu_inst_pe_1_5_3_U76 ( .B1(npu_inst_pe_1_5_3_n61), .B2(
        npu_inst_pe_1_5_3_n52), .A(npu_inst_pe_1_5_3_n69), .ZN(
        npu_inst_pe_1_5_3_n92) );
  NAND2_X1 npu_inst_pe_1_5_3_U75 ( .A1(npu_inst_pe_1_5_3_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_5_3_n48), .ZN(npu_inst_pe_1_5_3_n68) );
  OAI21_X1 npu_inst_pe_1_5_3_U74 ( .B1(npu_inst_pe_1_5_3_n63), .B2(
        npu_inst_pe_1_5_3_n48), .A(npu_inst_pe_1_5_3_n68), .ZN(
        npu_inst_pe_1_5_3_n91) );
  NAND2_X1 npu_inst_pe_1_5_3_U73 ( .A1(npu_inst_pe_1_5_3_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_5_3_n48), .ZN(npu_inst_pe_1_5_3_n67) );
  OAI21_X1 npu_inst_pe_1_5_3_U72 ( .B1(npu_inst_pe_1_5_3_n61), .B2(
        npu_inst_pe_1_5_3_n48), .A(npu_inst_pe_1_5_3_n67), .ZN(
        npu_inst_pe_1_5_3_n90) );
  NAND2_X1 npu_inst_pe_1_5_3_U71 ( .A1(npu_inst_pe_1_5_3_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_5_3_n44), .ZN(npu_inst_pe_1_5_3_n66) );
  OAI21_X1 npu_inst_pe_1_5_3_U70 ( .B1(npu_inst_pe_1_5_3_n63), .B2(
        npu_inst_pe_1_5_3_n44), .A(npu_inst_pe_1_5_3_n66), .ZN(
        npu_inst_pe_1_5_3_n89) );
  NAND2_X1 npu_inst_pe_1_5_3_U69 ( .A1(npu_inst_pe_1_5_3_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_5_3_n44), .ZN(npu_inst_pe_1_5_3_n65) );
  OAI21_X1 npu_inst_pe_1_5_3_U68 ( .B1(npu_inst_pe_1_5_3_n61), .B2(
        npu_inst_pe_1_5_3_n44), .A(npu_inst_pe_1_5_3_n65), .ZN(
        npu_inst_pe_1_5_3_n88) );
  NAND2_X1 npu_inst_pe_1_5_3_U67 ( .A1(npu_inst_pe_1_5_3_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_5_3_n40), .ZN(npu_inst_pe_1_5_3_n64) );
  OAI21_X1 npu_inst_pe_1_5_3_U66 ( .B1(npu_inst_pe_1_5_3_n63), .B2(
        npu_inst_pe_1_5_3_n40), .A(npu_inst_pe_1_5_3_n64), .ZN(
        npu_inst_pe_1_5_3_n87) );
  NAND2_X1 npu_inst_pe_1_5_3_U65 ( .A1(npu_inst_pe_1_5_3_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_5_3_n40), .ZN(npu_inst_pe_1_5_3_n62) );
  OAI21_X1 npu_inst_pe_1_5_3_U64 ( .B1(npu_inst_pe_1_5_3_n61), .B2(
        npu_inst_pe_1_5_3_n40), .A(npu_inst_pe_1_5_3_n62), .ZN(
        npu_inst_pe_1_5_3_n86) );
  AND2_X1 npu_inst_pe_1_5_3_U63 ( .A1(npu_inst_pe_1_5_3_N93), .A2(npu_inst_n54), .ZN(npu_inst_int_data_y_5__3__0_) );
  AND2_X1 npu_inst_pe_1_5_3_U62 ( .A1(npu_inst_n54), .A2(npu_inst_pe_1_5_3_N94), .ZN(npu_inst_int_data_y_5__3__1_) );
  NOR3_X1 npu_inst_pe_1_5_3_U61 ( .A1(npu_inst_pe_1_5_3_n26), .A2(npu_inst_n54), .A3(npu_inst_int_ckg[20]), .ZN(npu_inst_pe_1_5_3_n85) );
  OR2_X1 npu_inst_pe_1_5_3_U60 ( .A1(npu_inst_pe_1_5_3_n85), .A2(
        npu_inst_pe_1_5_3_n2), .ZN(npu_inst_pe_1_5_3_N84) );
  AND2_X1 npu_inst_pe_1_5_3_U59 ( .A1(npu_inst_pe_1_5_3_int_q_acc_0_), .A2(
        npu_inst_pe_1_5_3_n1), .ZN(npu_inst_int_data_res_5__3__0_) );
  AND2_X1 npu_inst_pe_1_5_3_U58 ( .A1(npu_inst_pe_1_5_3_n2), .A2(
        npu_inst_pe_1_5_3_int_q_acc_7_), .ZN(npu_inst_int_data_res_5__3__7_)
         );
  AND2_X1 npu_inst_pe_1_5_3_U57 ( .A1(npu_inst_pe_1_5_3_int_q_acc_1_), .A2(
        npu_inst_pe_1_5_3_n1), .ZN(npu_inst_int_data_res_5__3__1_) );
  AND2_X1 npu_inst_pe_1_5_3_U56 ( .A1(npu_inst_pe_1_5_3_int_q_acc_2_), .A2(
        npu_inst_pe_1_5_3_n1), .ZN(npu_inst_int_data_res_5__3__2_) );
  AND2_X1 npu_inst_pe_1_5_3_U55 ( .A1(npu_inst_pe_1_5_3_int_q_acc_3_), .A2(
        npu_inst_pe_1_5_3_n2), .ZN(npu_inst_int_data_res_5__3__3_) );
  AND2_X1 npu_inst_pe_1_5_3_U54 ( .A1(npu_inst_pe_1_5_3_int_q_acc_4_), .A2(
        npu_inst_pe_1_5_3_n2), .ZN(npu_inst_int_data_res_5__3__4_) );
  AND2_X1 npu_inst_pe_1_5_3_U53 ( .A1(npu_inst_pe_1_5_3_int_q_acc_5_), .A2(
        npu_inst_pe_1_5_3_n2), .ZN(npu_inst_int_data_res_5__3__5_) );
  AND2_X1 npu_inst_pe_1_5_3_U52 ( .A1(npu_inst_pe_1_5_3_int_q_acc_6_), .A2(
        npu_inst_pe_1_5_3_n2), .ZN(npu_inst_int_data_res_5__3__6_) );
  AOI222_X1 npu_inst_pe_1_5_3_U51 ( .A1(npu_inst_int_data_res_6__3__0_), .A2(
        npu_inst_pe_1_5_3_n1), .B1(npu_inst_pe_1_5_3_N73), .B2(
        npu_inst_pe_1_5_3_n76), .C1(npu_inst_pe_1_5_3_N65), .C2(
        npu_inst_pe_1_5_3_n77), .ZN(npu_inst_pe_1_5_3_n84) );
  INV_X1 npu_inst_pe_1_5_3_U50 ( .A(npu_inst_pe_1_5_3_n84), .ZN(
        npu_inst_pe_1_5_3_n101) );
  AOI222_X1 npu_inst_pe_1_5_3_U49 ( .A1(npu_inst_int_data_res_6__3__7_), .A2(
        npu_inst_pe_1_5_3_n1), .B1(npu_inst_pe_1_5_3_N80), .B2(
        npu_inst_pe_1_5_3_n76), .C1(npu_inst_pe_1_5_3_N72), .C2(
        npu_inst_pe_1_5_3_n77), .ZN(npu_inst_pe_1_5_3_n75) );
  INV_X1 npu_inst_pe_1_5_3_U48 ( .A(npu_inst_pe_1_5_3_n75), .ZN(
        npu_inst_pe_1_5_3_n33) );
  AOI222_X1 npu_inst_pe_1_5_3_U47 ( .A1(npu_inst_int_data_res_6__3__1_), .A2(
        npu_inst_pe_1_5_3_n1), .B1(npu_inst_pe_1_5_3_N74), .B2(
        npu_inst_pe_1_5_3_n76), .C1(npu_inst_pe_1_5_3_N66), .C2(
        npu_inst_pe_1_5_3_n77), .ZN(npu_inst_pe_1_5_3_n83) );
  INV_X1 npu_inst_pe_1_5_3_U46 ( .A(npu_inst_pe_1_5_3_n83), .ZN(
        npu_inst_pe_1_5_3_n100) );
  AOI222_X1 npu_inst_pe_1_5_3_U45 ( .A1(npu_inst_int_data_res_6__3__2_), .A2(
        npu_inst_pe_1_5_3_n1), .B1(npu_inst_pe_1_5_3_N75), .B2(
        npu_inst_pe_1_5_3_n76), .C1(npu_inst_pe_1_5_3_N67), .C2(
        npu_inst_pe_1_5_3_n77), .ZN(npu_inst_pe_1_5_3_n82) );
  INV_X1 npu_inst_pe_1_5_3_U44 ( .A(npu_inst_pe_1_5_3_n82), .ZN(
        npu_inst_pe_1_5_3_n99) );
  AOI222_X1 npu_inst_pe_1_5_3_U43 ( .A1(npu_inst_int_data_res_6__3__3_), .A2(
        npu_inst_pe_1_5_3_n1), .B1(npu_inst_pe_1_5_3_N76), .B2(
        npu_inst_pe_1_5_3_n76), .C1(npu_inst_pe_1_5_3_N68), .C2(
        npu_inst_pe_1_5_3_n77), .ZN(npu_inst_pe_1_5_3_n81) );
  INV_X1 npu_inst_pe_1_5_3_U42 ( .A(npu_inst_pe_1_5_3_n81), .ZN(
        npu_inst_pe_1_5_3_n98) );
  AOI222_X1 npu_inst_pe_1_5_3_U41 ( .A1(npu_inst_int_data_res_6__3__4_), .A2(
        npu_inst_pe_1_5_3_n1), .B1(npu_inst_pe_1_5_3_N77), .B2(
        npu_inst_pe_1_5_3_n76), .C1(npu_inst_pe_1_5_3_N69), .C2(
        npu_inst_pe_1_5_3_n77), .ZN(npu_inst_pe_1_5_3_n80) );
  INV_X1 npu_inst_pe_1_5_3_U40 ( .A(npu_inst_pe_1_5_3_n80), .ZN(
        npu_inst_pe_1_5_3_n36) );
  AOI222_X1 npu_inst_pe_1_5_3_U39 ( .A1(npu_inst_int_data_res_6__3__5_), .A2(
        npu_inst_pe_1_5_3_n1), .B1(npu_inst_pe_1_5_3_N78), .B2(
        npu_inst_pe_1_5_3_n76), .C1(npu_inst_pe_1_5_3_N70), .C2(
        npu_inst_pe_1_5_3_n77), .ZN(npu_inst_pe_1_5_3_n79) );
  INV_X1 npu_inst_pe_1_5_3_U38 ( .A(npu_inst_pe_1_5_3_n79), .ZN(
        npu_inst_pe_1_5_3_n35) );
  AOI222_X1 npu_inst_pe_1_5_3_U37 ( .A1(npu_inst_int_data_res_6__3__6_), .A2(
        npu_inst_pe_1_5_3_n1), .B1(npu_inst_pe_1_5_3_N79), .B2(
        npu_inst_pe_1_5_3_n76), .C1(npu_inst_pe_1_5_3_N71), .C2(
        npu_inst_pe_1_5_3_n77), .ZN(npu_inst_pe_1_5_3_n78) );
  INV_X1 npu_inst_pe_1_5_3_U36 ( .A(npu_inst_pe_1_5_3_n78), .ZN(
        npu_inst_pe_1_5_3_n34) );
  INV_X1 npu_inst_pe_1_5_3_U35 ( .A(npu_inst_pe_1_5_3_int_data_1_), .ZN(
        npu_inst_pe_1_5_3_n14) );
  AND2_X1 npu_inst_pe_1_5_3_U34 ( .A1(npu_inst_int_data_x_5__3__1_), .A2(
        npu_inst_pe_1_5_3_int_q_weight_1_), .ZN(npu_inst_pe_1_5_3_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_5_3_U33 ( .A1(npu_inst_int_data_x_5__3__0_), .A2(
        npu_inst_pe_1_5_3_int_q_weight_1_), .ZN(npu_inst_pe_1_5_3_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_5_3_U32 ( .A1(npu_inst_n54), .A2(
        npu_inst_int_data_y_6__3__1_), .B1(npu_inst_pe_1_5_3_n3), .B2(
        npu_inst_int_data_x_5__4__1_), .ZN(npu_inst_pe_1_5_3_n63) );
  AOI22_X1 npu_inst_pe_1_5_3_U31 ( .A1(npu_inst_n54), .A2(
        npu_inst_int_data_y_6__3__0_), .B1(npu_inst_pe_1_5_3_n3), .B2(
        npu_inst_int_data_x_5__4__0_), .ZN(npu_inst_pe_1_5_3_n61) );
  INV_X1 npu_inst_pe_1_5_3_U30 ( .A(npu_inst_pe_1_5_3_int_data_0_), .ZN(
        npu_inst_pe_1_5_3_n13) );
  INV_X1 npu_inst_pe_1_5_3_U29 ( .A(npu_inst_n68), .ZN(npu_inst_pe_1_5_3_n5)
         );
  OR3_X1 npu_inst_pe_1_5_3_U28 ( .A1(npu_inst_pe_1_5_3_n6), .A2(
        npu_inst_pe_1_5_3_n8), .A3(npu_inst_pe_1_5_3_n5), .ZN(
        npu_inst_pe_1_5_3_n56) );
  OR3_X1 npu_inst_pe_1_5_3_U27 ( .A1(npu_inst_pe_1_5_3_n5), .A2(
        npu_inst_pe_1_5_3_n8), .A3(npu_inst_pe_1_5_3_n7), .ZN(
        npu_inst_pe_1_5_3_n48) );
  INV_X1 npu_inst_pe_1_5_3_U26 ( .A(npu_inst_pe_1_5_3_n5), .ZN(
        npu_inst_pe_1_5_3_n4) );
  INV_X1 npu_inst_pe_1_5_3_U25 ( .A(npu_inst_n123), .ZN(npu_inst_pe_1_5_3_n12)
         );
  OR3_X1 npu_inst_pe_1_5_3_U24 ( .A1(npu_inst_pe_1_5_3_n4), .A2(
        npu_inst_pe_1_5_3_n8), .A3(npu_inst_pe_1_5_3_n7), .ZN(
        npu_inst_pe_1_5_3_n52) );
  OR3_X1 npu_inst_pe_1_5_3_U23 ( .A1(npu_inst_pe_1_5_3_n6), .A2(
        npu_inst_pe_1_5_3_n8), .A3(npu_inst_pe_1_5_3_n4), .ZN(
        npu_inst_pe_1_5_3_n60) );
  NOR2_X1 npu_inst_pe_1_5_3_U22 ( .A1(npu_inst_pe_1_5_3_n60), .A2(
        npu_inst_pe_1_5_3_n3), .ZN(npu_inst_pe_1_5_3_n58) );
  NOR2_X1 npu_inst_pe_1_5_3_U21 ( .A1(npu_inst_pe_1_5_3_n56), .A2(
        npu_inst_pe_1_5_3_n3), .ZN(npu_inst_pe_1_5_3_n54) );
  NOR2_X1 npu_inst_pe_1_5_3_U20 ( .A1(npu_inst_pe_1_5_3_n52), .A2(
        npu_inst_pe_1_5_3_n3), .ZN(npu_inst_pe_1_5_3_n50) );
  NOR2_X1 npu_inst_pe_1_5_3_U19 ( .A1(npu_inst_pe_1_5_3_n48), .A2(
        npu_inst_pe_1_5_3_n3), .ZN(npu_inst_pe_1_5_3_n46) );
  NOR2_X1 npu_inst_pe_1_5_3_U18 ( .A1(npu_inst_pe_1_5_3_n40), .A2(
        npu_inst_pe_1_5_3_n3), .ZN(npu_inst_pe_1_5_3_n38) );
  NOR2_X1 npu_inst_pe_1_5_3_U17 ( .A1(npu_inst_pe_1_5_3_n44), .A2(
        npu_inst_pe_1_5_3_n3), .ZN(npu_inst_pe_1_5_3_n42) );
  BUF_X1 npu_inst_pe_1_5_3_U16 ( .A(npu_inst_n97), .Z(npu_inst_pe_1_5_3_n8) );
  BUF_X1 npu_inst_pe_1_5_3_U15 ( .A(npu_inst_pe_1_5_3_n12), .Z(
        npu_inst_pe_1_5_3_n11) );
  BUF_X1 npu_inst_pe_1_5_3_U14 ( .A(npu_inst_pe_1_5_3_n12), .Z(
        npu_inst_pe_1_5_3_n10) );
  BUF_X1 npu_inst_pe_1_5_3_U13 ( .A(npu_inst_pe_1_5_3_n12), .Z(
        npu_inst_pe_1_5_3_n9) );
  INV_X1 npu_inst_pe_1_5_3_U12 ( .A(npu_inst_pe_1_5_3_n38), .ZN(
        npu_inst_pe_1_5_3_n118) );
  INV_X1 npu_inst_pe_1_5_3_U11 ( .A(npu_inst_pe_1_5_3_n58), .ZN(
        npu_inst_pe_1_5_3_n114) );
  INV_X1 npu_inst_pe_1_5_3_U10 ( .A(npu_inst_pe_1_5_3_n54), .ZN(
        npu_inst_pe_1_5_3_n115) );
  INV_X1 npu_inst_pe_1_5_3_U9 ( .A(npu_inst_pe_1_5_3_n50), .ZN(
        npu_inst_pe_1_5_3_n116) );
  INV_X1 npu_inst_pe_1_5_3_U8 ( .A(npu_inst_pe_1_5_3_n46), .ZN(
        npu_inst_pe_1_5_3_n117) );
  INV_X1 npu_inst_pe_1_5_3_U7 ( .A(npu_inst_pe_1_5_3_n42), .ZN(
        npu_inst_pe_1_5_3_n119) );
  BUF_X1 npu_inst_pe_1_5_3_U6 ( .A(npu_inst_n17), .Z(npu_inst_pe_1_5_3_n2) );
  BUF_X1 npu_inst_pe_1_5_3_U5 ( .A(npu_inst_n17), .Z(npu_inst_pe_1_5_3_n1) );
  NOR2_X1 npu_inst_pe_1_5_3_U4 ( .A1(npu_inst_pe_1_5_3_int_q_weight_0_), .A2(
        npu_inst_pe_1_5_3_n1), .ZN(npu_inst_pe_1_5_3_n76) );
  NOR2_X1 npu_inst_pe_1_5_3_U3 ( .A1(npu_inst_pe_1_5_3_n27), .A2(
        npu_inst_pe_1_5_3_n1), .ZN(npu_inst_pe_1_5_3_n77) );
  FA_X1 npu_inst_pe_1_5_3_sub_77_U2_1 ( .A(npu_inst_pe_1_5_3_int_q_acc_1_), 
        .B(npu_inst_pe_1_5_3_n14), .CI(npu_inst_pe_1_5_3_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_5_3_sub_77_carry_2_), .S(npu_inst_pe_1_5_3_N66) );
  FA_X1 npu_inst_pe_1_5_3_add_79_U1_1 ( .A(npu_inst_pe_1_5_3_int_q_acc_1_), 
        .B(npu_inst_pe_1_5_3_int_data_1_), .CI(
        npu_inst_pe_1_5_3_add_79_carry_1_), .CO(
        npu_inst_pe_1_5_3_add_79_carry_2_), .S(npu_inst_pe_1_5_3_N74) );
  NAND3_X1 npu_inst_pe_1_5_3_U109 ( .A1(npu_inst_pe_1_5_3_n5), .A2(
        npu_inst_pe_1_5_3_n7), .A3(npu_inst_pe_1_5_3_n8), .ZN(
        npu_inst_pe_1_5_3_n44) );
  NAND3_X1 npu_inst_pe_1_5_3_U108 ( .A1(npu_inst_pe_1_5_3_n4), .A2(
        npu_inst_pe_1_5_3_n7), .A3(npu_inst_pe_1_5_3_n8), .ZN(
        npu_inst_pe_1_5_3_n40) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_5_3_n34), .CK(
        npu_inst_pe_1_5_3_net3304), .RN(npu_inst_pe_1_5_3_n9), .Q(
        npu_inst_pe_1_5_3_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_5_3_n35), .CK(
        npu_inst_pe_1_5_3_net3304), .RN(npu_inst_pe_1_5_3_n9), .Q(
        npu_inst_pe_1_5_3_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_5_3_n36), .CK(
        npu_inst_pe_1_5_3_net3304), .RN(npu_inst_pe_1_5_3_n9), .Q(
        npu_inst_pe_1_5_3_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_5_3_n98), .CK(
        npu_inst_pe_1_5_3_net3304), .RN(npu_inst_pe_1_5_3_n9), .Q(
        npu_inst_pe_1_5_3_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_5_3_n99), .CK(
        npu_inst_pe_1_5_3_net3304), .RN(npu_inst_pe_1_5_3_n9), .Q(
        npu_inst_pe_1_5_3_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_5_3_n100), 
        .CK(npu_inst_pe_1_5_3_net3304), .RN(npu_inst_pe_1_5_3_n9), .Q(
        npu_inst_pe_1_5_3_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_5_3_n33), .CK(
        npu_inst_pe_1_5_3_net3304), .RN(npu_inst_pe_1_5_3_n9), .Q(
        npu_inst_pe_1_5_3_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_5_3_n101), 
        .CK(npu_inst_pe_1_5_3_net3304), .RN(npu_inst_pe_1_5_3_n9), .Q(
        npu_inst_pe_1_5_3_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_weight_reg_0_ ( .D(npu_inst_n109), .CK(
        npu_inst_pe_1_5_3_net3310), .RN(npu_inst_pe_1_5_3_n9), .Q(
        npu_inst_pe_1_5_3_int_q_weight_0_), .QN(npu_inst_pe_1_5_3_n27) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_weight_reg_1_ ( .D(npu_inst_n115), .CK(
        npu_inst_pe_1_5_3_net3310), .RN(npu_inst_pe_1_5_3_n9), .Q(
        npu_inst_pe_1_5_3_int_q_weight_1_), .QN(npu_inst_pe_1_5_3_n26) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_5_3_n113), 
        .CK(npu_inst_pe_1_5_3_net3310), .RN(npu_inst_pe_1_5_3_n9), .Q(
        npu_inst_pe_1_5_3_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_5_3_n107), 
        .CK(npu_inst_pe_1_5_3_net3310), .RN(npu_inst_pe_1_5_3_n9), .Q(
        npu_inst_pe_1_5_3_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_5_3_n112), 
        .CK(npu_inst_pe_1_5_3_net3310), .RN(npu_inst_pe_1_5_3_n10), .Q(
        npu_inst_pe_1_5_3_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_5_3_n106), 
        .CK(npu_inst_pe_1_5_3_net3310), .RN(npu_inst_pe_1_5_3_n10), .Q(
        npu_inst_pe_1_5_3_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_5_3_n111), 
        .CK(npu_inst_pe_1_5_3_net3310), .RN(npu_inst_pe_1_5_3_n10), .Q(
        npu_inst_pe_1_5_3_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_5_3_n105), 
        .CK(npu_inst_pe_1_5_3_net3310), .RN(npu_inst_pe_1_5_3_n10), .Q(
        npu_inst_pe_1_5_3_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_5_3_n110), 
        .CK(npu_inst_pe_1_5_3_net3310), .RN(npu_inst_pe_1_5_3_n10), .Q(
        npu_inst_pe_1_5_3_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_5_3_n104), 
        .CK(npu_inst_pe_1_5_3_net3310), .RN(npu_inst_pe_1_5_3_n10), .Q(
        npu_inst_pe_1_5_3_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_5_3_n109), 
        .CK(npu_inst_pe_1_5_3_net3310), .RN(npu_inst_pe_1_5_3_n10), .Q(
        npu_inst_pe_1_5_3_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_5_3_n103), 
        .CK(npu_inst_pe_1_5_3_net3310), .RN(npu_inst_pe_1_5_3_n10), .Q(
        npu_inst_pe_1_5_3_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_5_3_n108), 
        .CK(npu_inst_pe_1_5_3_net3310), .RN(npu_inst_pe_1_5_3_n10), .Q(
        npu_inst_pe_1_5_3_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_5_3_n102), 
        .CK(npu_inst_pe_1_5_3_net3310), .RN(npu_inst_pe_1_5_3_n10), .Q(
        npu_inst_pe_1_5_3_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_5_3_n86), 
        .CK(npu_inst_pe_1_5_3_net3310), .RN(npu_inst_pe_1_5_3_n10), .Q(
        npu_inst_pe_1_5_3_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_5_3_n87), 
        .CK(npu_inst_pe_1_5_3_net3310), .RN(npu_inst_pe_1_5_3_n10), .Q(
        npu_inst_pe_1_5_3_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_5_3_n88), 
        .CK(npu_inst_pe_1_5_3_net3310), .RN(npu_inst_pe_1_5_3_n11), .Q(
        npu_inst_pe_1_5_3_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_5_3_n89), 
        .CK(npu_inst_pe_1_5_3_net3310), .RN(npu_inst_pe_1_5_3_n11), .Q(
        npu_inst_pe_1_5_3_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_5_3_n90), 
        .CK(npu_inst_pe_1_5_3_net3310), .RN(npu_inst_pe_1_5_3_n11), .Q(
        npu_inst_pe_1_5_3_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_5_3_n91), 
        .CK(npu_inst_pe_1_5_3_net3310), .RN(npu_inst_pe_1_5_3_n11), .Q(
        npu_inst_pe_1_5_3_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_5_3_n92), 
        .CK(npu_inst_pe_1_5_3_net3310), .RN(npu_inst_pe_1_5_3_n11), .Q(
        npu_inst_pe_1_5_3_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_5_3_n93), 
        .CK(npu_inst_pe_1_5_3_net3310), .RN(npu_inst_pe_1_5_3_n11), .Q(
        npu_inst_pe_1_5_3_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_5_3_n94), 
        .CK(npu_inst_pe_1_5_3_net3310), .RN(npu_inst_pe_1_5_3_n11), .Q(
        npu_inst_pe_1_5_3_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_5_3_n95), 
        .CK(npu_inst_pe_1_5_3_net3310), .RN(npu_inst_pe_1_5_3_n11), .Q(
        npu_inst_pe_1_5_3_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_5_3_n96), 
        .CK(npu_inst_pe_1_5_3_net3310), .RN(npu_inst_pe_1_5_3_n11), .Q(
        npu_inst_pe_1_5_3_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_5_3_n97), 
        .CK(npu_inst_pe_1_5_3_net3310), .RN(npu_inst_pe_1_5_3_n11), .Q(
        npu_inst_pe_1_5_3_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_5_3_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_5_3_N84), .SE(1'b0), .GCK(npu_inst_pe_1_5_3_net3304) );
  CLKGATETST_X1 npu_inst_pe_1_5_3_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n62), .SE(1'b0), .GCK(npu_inst_pe_1_5_3_net3310) );
  MUX2_X1 npu_inst_pe_1_5_4_U162 ( .A(npu_inst_pe_1_5_4_n32), .B(
        npu_inst_pe_1_5_4_n29), .S(npu_inst_pe_1_5_4_n8), .Z(
        npu_inst_pe_1_5_4_N93) );
  MUX2_X1 npu_inst_pe_1_5_4_U161 ( .A(npu_inst_pe_1_5_4_n31), .B(
        npu_inst_pe_1_5_4_n30), .S(npu_inst_pe_1_5_4_n6), .Z(
        npu_inst_pe_1_5_4_n32) );
  MUX2_X1 npu_inst_pe_1_5_4_U160 ( .A(npu_inst_pe_1_5_4_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_5_4_int_q_reg_v_1__0_), .S(npu_inst_pe_1_5_4_n4), .Z(
        npu_inst_pe_1_5_4_n31) );
  MUX2_X1 npu_inst_pe_1_5_4_U159 ( .A(npu_inst_pe_1_5_4_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_5_4_int_q_reg_v_3__0_), .S(npu_inst_pe_1_5_4_n4), .Z(
        npu_inst_pe_1_5_4_n30) );
  MUX2_X1 npu_inst_pe_1_5_4_U158 ( .A(npu_inst_pe_1_5_4_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_5_4_int_q_reg_v_5__0_), .S(npu_inst_pe_1_5_4_n4), .Z(
        npu_inst_pe_1_5_4_n29) );
  MUX2_X1 npu_inst_pe_1_5_4_U157 ( .A(npu_inst_pe_1_5_4_n28), .B(
        npu_inst_pe_1_5_4_n23), .S(npu_inst_pe_1_5_4_n8), .Z(
        npu_inst_pe_1_5_4_N94) );
  MUX2_X1 npu_inst_pe_1_5_4_U156 ( .A(npu_inst_pe_1_5_4_n25), .B(
        npu_inst_pe_1_5_4_n24), .S(npu_inst_pe_1_5_4_n6), .Z(
        npu_inst_pe_1_5_4_n28) );
  MUX2_X1 npu_inst_pe_1_5_4_U155 ( .A(npu_inst_pe_1_5_4_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_5_4_int_q_reg_v_1__1_), .S(npu_inst_pe_1_5_4_n4), .Z(
        npu_inst_pe_1_5_4_n25) );
  MUX2_X1 npu_inst_pe_1_5_4_U154 ( .A(npu_inst_pe_1_5_4_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_5_4_int_q_reg_v_3__1_), .S(npu_inst_pe_1_5_4_n4), .Z(
        npu_inst_pe_1_5_4_n24) );
  MUX2_X1 npu_inst_pe_1_5_4_U153 ( .A(npu_inst_pe_1_5_4_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_5_4_int_q_reg_v_5__1_), .S(npu_inst_pe_1_5_4_n4), .Z(
        npu_inst_pe_1_5_4_n23) );
  MUX2_X1 npu_inst_pe_1_5_4_U152 ( .A(npu_inst_pe_1_5_4_n22), .B(
        npu_inst_pe_1_5_4_n19), .S(npu_inst_pe_1_5_4_n8), .Z(
        npu_inst_int_data_x_5__4__1_) );
  MUX2_X1 npu_inst_pe_1_5_4_U151 ( .A(npu_inst_pe_1_5_4_n21), .B(
        npu_inst_pe_1_5_4_n20), .S(npu_inst_pe_1_5_4_n6), .Z(
        npu_inst_pe_1_5_4_n22) );
  MUX2_X1 npu_inst_pe_1_5_4_U150 ( .A(npu_inst_pe_1_5_4_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_5_4_int_q_reg_h_1__1_), .S(npu_inst_pe_1_5_4_n4), .Z(
        npu_inst_pe_1_5_4_n21) );
  MUX2_X1 npu_inst_pe_1_5_4_U149 ( .A(npu_inst_pe_1_5_4_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_5_4_int_q_reg_h_3__1_), .S(npu_inst_pe_1_5_4_n4), .Z(
        npu_inst_pe_1_5_4_n20) );
  MUX2_X1 npu_inst_pe_1_5_4_U148 ( .A(npu_inst_pe_1_5_4_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_5_4_int_q_reg_h_5__1_), .S(npu_inst_pe_1_5_4_n4), .Z(
        npu_inst_pe_1_5_4_n19) );
  MUX2_X1 npu_inst_pe_1_5_4_U147 ( .A(npu_inst_pe_1_5_4_n18), .B(
        npu_inst_pe_1_5_4_n15), .S(npu_inst_pe_1_5_4_n8), .Z(
        npu_inst_int_data_x_5__4__0_) );
  MUX2_X1 npu_inst_pe_1_5_4_U146 ( .A(npu_inst_pe_1_5_4_n17), .B(
        npu_inst_pe_1_5_4_n16), .S(npu_inst_pe_1_5_4_n6), .Z(
        npu_inst_pe_1_5_4_n18) );
  MUX2_X1 npu_inst_pe_1_5_4_U145 ( .A(npu_inst_pe_1_5_4_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_5_4_int_q_reg_h_1__0_), .S(npu_inst_pe_1_5_4_n4), .Z(
        npu_inst_pe_1_5_4_n17) );
  MUX2_X1 npu_inst_pe_1_5_4_U144 ( .A(npu_inst_pe_1_5_4_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_5_4_int_q_reg_h_3__0_), .S(npu_inst_pe_1_5_4_n4), .Z(
        npu_inst_pe_1_5_4_n16) );
  MUX2_X1 npu_inst_pe_1_5_4_U143 ( .A(npu_inst_pe_1_5_4_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_5_4_int_q_reg_h_5__0_), .S(npu_inst_pe_1_5_4_n4), .Z(
        npu_inst_pe_1_5_4_n15) );
  XOR2_X1 npu_inst_pe_1_5_4_U142 ( .A(npu_inst_pe_1_5_4_int_data_0_), .B(
        npu_inst_pe_1_5_4_int_q_acc_0_), .Z(npu_inst_pe_1_5_4_N73) );
  AND2_X1 npu_inst_pe_1_5_4_U141 ( .A1(npu_inst_pe_1_5_4_int_q_acc_0_), .A2(
        npu_inst_pe_1_5_4_int_data_0_), .ZN(npu_inst_pe_1_5_4_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_5_4_U140 ( .A(npu_inst_pe_1_5_4_int_q_acc_0_), .B(
        npu_inst_pe_1_5_4_n13), .ZN(npu_inst_pe_1_5_4_N65) );
  OR2_X1 npu_inst_pe_1_5_4_U139 ( .A1(npu_inst_pe_1_5_4_n13), .A2(
        npu_inst_pe_1_5_4_int_q_acc_0_), .ZN(npu_inst_pe_1_5_4_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_5_4_U138 ( .A(npu_inst_pe_1_5_4_int_q_acc_2_), .B(
        npu_inst_pe_1_5_4_add_79_carry_2_), .Z(npu_inst_pe_1_5_4_N75) );
  AND2_X1 npu_inst_pe_1_5_4_U137 ( .A1(npu_inst_pe_1_5_4_add_79_carry_2_), 
        .A2(npu_inst_pe_1_5_4_int_q_acc_2_), .ZN(
        npu_inst_pe_1_5_4_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_5_4_U136 ( .A(npu_inst_pe_1_5_4_int_q_acc_3_), .B(
        npu_inst_pe_1_5_4_add_79_carry_3_), .Z(npu_inst_pe_1_5_4_N76) );
  AND2_X1 npu_inst_pe_1_5_4_U135 ( .A1(npu_inst_pe_1_5_4_add_79_carry_3_), 
        .A2(npu_inst_pe_1_5_4_int_q_acc_3_), .ZN(
        npu_inst_pe_1_5_4_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_5_4_U134 ( .A(npu_inst_pe_1_5_4_int_q_acc_4_), .B(
        npu_inst_pe_1_5_4_add_79_carry_4_), .Z(npu_inst_pe_1_5_4_N77) );
  AND2_X1 npu_inst_pe_1_5_4_U133 ( .A1(npu_inst_pe_1_5_4_add_79_carry_4_), 
        .A2(npu_inst_pe_1_5_4_int_q_acc_4_), .ZN(
        npu_inst_pe_1_5_4_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_5_4_U132 ( .A(npu_inst_pe_1_5_4_int_q_acc_5_), .B(
        npu_inst_pe_1_5_4_add_79_carry_5_), .Z(npu_inst_pe_1_5_4_N78) );
  AND2_X1 npu_inst_pe_1_5_4_U131 ( .A1(npu_inst_pe_1_5_4_add_79_carry_5_), 
        .A2(npu_inst_pe_1_5_4_int_q_acc_5_), .ZN(
        npu_inst_pe_1_5_4_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_5_4_U130 ( .A(npu_inst_pe_1_5_4_int_q_acc_6_), .B(
        npu_inst_pe_1_5_4_add_79_carry_6_), .Z(npu_inst_pe_1_5_4_N79) );
  AND2_X1 npu_inst_pe_1_5_4_U129 ( .A1(npu_inst_pe_1_5_4_add_79_carry_6_), 
        .A2(npu_inst_pe_1_5_4_int_q_acc_6_), .ZN(
        npu_inst_pe_1_5_4_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_5_4_U128 ( .A(npu_inst_pe_1_5_4_int_q_acc_7_), .B(
        npu_inst_pe_1_5_4_add_79_carry_7_), .Z(npu_inst_pe_1_5_4_N80) );
  XNOR2_X1 npu_inst_pe_1_5_4_U127 ( .A(npu_inst_pe_1_5_4_sub_77_carry_2_), .B(
        npu_inst_pe_1_5_4_int_q_acc_2_), .ZN(npu_inst_pe_1_5_4_N67) );
  OR2_X1 npu_inst_pe_1_5_4_U126 ( .A1(npu_inst_pe_1_5_4_int_q_acc_2_), .A2(
        npu_inst_pe_1_5_4_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_5_4_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_5_4_U125 ( .A(npu_inst_pe_1_5_4_sub_77_carry_3_), .B(
        npu_inst_pe_1_5_4_int_q_acc_3_), .ZN(npu_inst_pe_1_5_4_N68) );
  OR2_X1 npu_inst_pe_1_5_4_U124 ( .A1(npu_inst_pe_1_5_4_int_q_acc_3_), .A2(
        npu_inst_pe_1_5_4_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_5_4_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_5_4_U123 ( .A(npu_inst_pe_1_5_4_sub_77_carry_4_), .B(
        npu_inst_pe_1_5_4_int_q_acc_4_), .ZN(npu_inst_pe_1_5_4_N69) );
  OR2_X1 npu_inst_pe_1_5_4_U122 ( .A1(npu_inst_pe_1_5_4_int_q_acc_4_), .A2(
        npu_inst_pe_1_5_4_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_5_4_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_5_4_U121 ( .A(npu_inst_pe_1_5_4_sub_77_carry_5_), .B(
        npu_inst_pe_1_5_4_int_q_acc_5_), .ZN(npu_inst_pe_1_5_4_N70) );
  OR2_X1 npu_inst_pe_1_5_4_U120 ( .A1(npu_inst_pe_1_5_4_int_q_acc_5_), .A2(
        npu_inst_pe_1_5_4_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_5_4_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_5_4_U119 ( .A(npu_inst_pe_1_5_4_sub_77_carry_6_), .B(
        npu_inst_pe_1_5_4_int_q_acc_6_), .ZN(npu_inst_pe_1_5_4_N71) );
  OR2_X1 npu_inst_pe_1_5_4_U118 ( .A1(npu_inst_pe_1_5_4_int_q_acc_6_), .A2(
        npu_inst_pe_1_5_4_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_5_4_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_5_4_U117 ( .A(npu_inst_pe_1_5_4_int_q_acc_7_), .B(
        npu_inst_pe_1_5_4_sub_77_carry_7_), .ZN(npu_inst_pe_1_5_4_N72) );
  INV_X1 npu_inst_pe_1_5_4_U116 ( .A(npu_inst_n76), .ZN(npu_inst_pe_1_5_4_n7)
         );
  INV_X1 npu_inst_pe_1_5_4_U115 ( .A(npu_inst_pe_1_5_4_n7), .ZN(
        npu_inst_pe_1_5_4_n6) );
  INV_X1 npu_inst_pe_1_5_4_U114 ( .A(npu_inst_n54), .ZN(npu_inst_pe_1_5_4_n3)
         );
  AOI22_X1 npu_inst_pe_1_5_4_U113 ( .A1(npu_inst_int_data_y_6__4__0_), .A2(
        npu_inst_pe_1_5_4_n58), .B1(npu_inst_pe_1_5_4_n114), .B2(
        npu_inst_pe_1_5_4_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_5_4_n57) );
  INV_X1 npu_inst_pe_1_5_4_U112 ( .A(npu_inst_pe_1_5_4_n57), .ZN(
        npu_inst_pe_1_5_4_n108) );
  AOI22_X1 npu_inst_pe_1_5_4_U111 ( .A1(npu_inst_int_data_y_6__4__0_), .A2(
        npu_inst_pe_1_5_4_n54), .B1(npu_inst_pe_1_5_4_n115), .B2(
        npu_inst_pe_1_5_4_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_5_4_n53) );
  INV_X1 npu_inst_pe_1_5_4_U110 ( .A(npu_inst_pe_1_5_4_n53), .ZN(
        npu_inst_pe_1_5_4_n109) );
  AOI22_X1 npu_inst_pe_1_5_4_U107 ( .A1(npu_inst_int_data_y_6__4__0_), .A2(
        npu_inst_pe_1_5_4_n50), .B1(npu_inst_pe_1_5_4_n116), .B2(
        npu_inst_pe_1_5_4_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_5_4_n49) );
  INV_X1 npu_inst_pe_1_5_4_U106 ( .A(npu_inst_pe_1_5_4_n49), .ZN(
        npu_inst_pe_1_5_4_n110) );
  AOI22_X1 npu_inst_pe_1_5_4_U105 ( .A1(npu_inst_int_data_y_6__4__0_), .A2(
        npu_inst_pe_1_5_4_n46), .B1(npu_inst_pe_1_5_4_n117), .B2(
        npu_inst_pe_1_5_4_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_5_4_n45) );
  INV_X1 npu_inst_pe_1_5_4_U104 ( .A(npu_inst_pe_1_5_4_n45), .ZN(
        npu_inst_pe_1_5_4_n111) );
  AOI22_X1 npu_inst_pe_1_5_4_U103 ( .A1(npu_inst_int_data_y_6__4__0_), .A2(
        npu_inst_pe_1_5_4_n42), .B1(npu_inst_pe_1_5_4_n119), .B2(
        npu_inst_pe_1_5_4_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_5_4_n41) );
  INV_X1 npu_inst_pe_1_5_4_U102 ( .A(npu_inst_pe_1_5_4_n41), .ZN(
        npu_inst_pe_1_5_4_n112) );
  AOI22_X1 npu_inst_pe_1_5_4_U101 ( .A1(npu_inst_int_data_y_6__4__1_), .A2(
        npu_inst_pe_1_5_4_n58), .B1(npu_inst_pe_1_5_4_n114), .B2(
        npu_inst_pe_1_5_4_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_5_4_n59) );
  INV_X1 npu_inst_pe_1_5_4_U100 ( .A(npu_inst_pe_1_5_4_n59), .ZN(
        npu_inst_pe_1_5_4_n102) );
  AOI22_X1 npu_inst_pe_1_5_4_U99 ( .A1(npu_inst_int_data_y_6__4__1_), .A2(
        npu_inst_pe_1_5_4_n54), .B1(npu_inst_pe_1_5_4_n115), .B2(
        npu_inst_pe_1_5_4_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_5_4_n55) );
  INV_X1 npu_inst_pe_1_5_4_U98 ( .A(npu_inst_pe_1_5_4_n55), .ZN(
        npu_inst_pe_1_5_4_n103) );
  AOI22_X1 npu_inst_pe_1_5_4_U97 ( .A1(npu_inst_int_data_y_6__4__1_), .A2(
        npu_inst_pe_1_5_4_n50), .B1(npu_inst_pe_1_5_4_n116), .B2(
        npu_inst_pe_1_5_4_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_5_4_n51) );
  INV_X1 npu_inst_pe_1_5_4_U96 ( .A(npu_inst_pe_1_5_4_n51), .ZN(
        npu_inst_pe_1_5_4_n104) );
  AOI22_X1 npu_inst_pe_1_5_4_U95 ( .A1(npu_inst_int_data_y_6__4__1_), .A2(
        npu_inst_pe_1_5_4_n46), .B1(npu_inst_pe_1_5_4_n117), .B2(
        npu_inst_pe_1_5_4_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_5_4_n47) );
  INV_X1 npu_inst_pe_1_5_4_U94 ( .A(npu_inst_pe_1_5_4_n47), .ZN(
        npu_inst_pe_1_5_4_n105) );
  AOI22_X1 npu_inst_pe_1_5_4_U93 ( .A1(npu_inst_int_data_y_6__4__1_), .A2(
        npu_inst_pe_1_5_4_n42), .B1(npu_inst_pe_1_5_4_n119), .B2(
        npu_inst_pe_1_5_4_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_5_4_n43) );
  INV_X1 npu_inst_pe_1_5_4_U92 ( .A(npu_inst_pe_1_5_4_n43), .ZN(
        npu_inst_pe_1_5_4_n106) );
  AOI22_X1 npu_inst_pe_1_5_4_U91 ( .A1(npu_inst_pe_1_5_4_n38), .A2(
        npu_inst_int_data_y_6__4__1_), .B1(npu_inst_pe_1_5_4_n118), .B2(
        npu_inst_pe_1_5_4_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_5_4_n39) );
  INV_X1 npu_inst_pe_1_5_4_U90 ( .A(npu_inst_pe_1_5_4_n39), .ZN(
        npu_inst_pe_1_5_4_n107) );
  AOI22_X1 npu_inst_pe_1_5_4_U89 ( .A1(npu_inst_pe_1_5_4_n38), .A2(
        npu_inst_int_data_y_6__4__0_), .B1(npu_inst_pe_1_5_4_n118), .B2(
        npu_inst_pe_1_5_4_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_5_4_n37) );
  INV_X1 npu_inst_pe_1_5_4_U88 ( .A(npu_inst_pe_1_5_4_n37), .ZN(
        npu_inst_pe_1_5_4_n113) );
  NAND2_X1 npu_inst_pe_1_5_4_U87 ( .A1(npu_inst_pe_1_5_4_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_5_4_n60), .ZN(npu_inst_pe_1_5_4_n74) );
  OAI21_X1 npu_inst_pe_1_5_4_U86 ( .B1(npu_inst_pe_1_5_4_n63), .B2(
        npu_inst_pe_1_5_4_n60), .A(npu_inst_pe_1_5_4_n74), .ZN(
        npu_inst_pe_1_5_4_n97) );
  NAND2_X1 npu_inst_pe_1_5_4_U85 ( .A1(npu_inst_pe_1_5_4_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_5_4_n60), .ZN(npu_inst_pe_1_5_4_n73) );
  OAI21_X1 npu_inst_pe_1_5_4_U84 ( .B1(npu_inst_pe_1_5_4_n61), .B2(
        npu_inst_pe_1_5_4_n60), .A(npu_inst_pe_1_5_4_n73), .ZN(
        npu_inst_pe_1_5_4_n96) );
  NAND2_X1 npu_inst_pe_1_5_4_U83 ( .A1(npu_inst_pe_1_5_4_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_5_4_n56), .ZN(npu_inst_pe_1_5_4_n72) );
  OAI21_X1 npu_inst_pe_1_5_4_U82 ( .B1(npu_inst_pe_1_5_4_n63), .B2(
        npu_inst_pe_1_5_4_n56), .A(npu_inst_pe_1_5_4_n72), .ZN(
        npu_inst_pe_1_5_4_n95) );
  NAND2_X1 npu_inst_pe_1_5_4_U81 ( .A1(npu_inst_pe_1_5_4_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_5_4_n56), .ZN(npu_inst_pe_1_5_4_n71) );
  OAI21_X1 npu_inst_pe_1_5_4_U80 ( .B1(npu_inst_pe_1_5_4_n61), .B2(
        npu_inst_pe_1_5_4_n56), .A(npu_inst_pe_1_5_4_n71), .ZN(
        npu_inst_pe_1_5_4_n94) );
  NAND2_X1 npu_inst_pe_1_5_4_U79 ( .A1(npu_inst_pe_1_5_4_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_5_4_n52), .ZN(npu_inst_pe_1_5_4_n70) );
  OAI21_X1 npu_inst_pe_1_5_4_U78 ( .B1(npu_inst_pe_1_5_4_n63), .B2(
        npu_inst_pe_1_5_4_n52), .A(npu_inst_pe_1_5_4_n70), .ZN(
        npu_inst_pe_1_5_4_n93) );
  NAND2_X1 npu_inst_pe_1_5_4_U77 ( .A1(npu_inst_pe_1_5_4_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_5_4_n52), .ZN(npu_inst_pe_1_5_4_n69) );
  OAI21_X1 npu_inst_pe_1_5_4_U76 ( .B1(npu_inst_pe_1_5_4_n61), .B2(
        npu_inst_pe_1_5_4_n52), .A(npu_inst_pe_1_5_4_n69), .ZN(
        npu_inst_pe_1_5_4_n92) );
  NAND2_X1 npu_inst_pe_1_5_4_U75 ( .A1(npu_inst_pe_1_5_4_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_5_4_n48), .ZN(npu_inst_pe_1_5_4_n68) );
  OAI21_X1 npu_inst_pe_1_5_4_U74 ( .B1(npu_inst_pe_1_5_4_n63), .B2(
        npu_inst_pe_1_5_4_n48), .A(npu_inst_pe_1_5_4_n68), .ZN(
        npu_inst_pe_1_5_4_n91) );
  NAND2_X1 npu_inst_pe_1_5_4_U73 ( .A1(npu_inst_pe_1_5_4_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_5_4_n48), .ZN(npu_inst_pe_1_5_4_n67) );
  OAI21_X1 npu_inst_pe_1_5_4_U72 ( .B1(npu_inst_pe_1_5_4_n61), .B2(
        npu_inst_pe_1_5_4_n48), .A(npu_inst_pe_1_5_4_n67), .ZN(
        npu_inst_pe_1_5_4_n90) );
  NAND2_X1 npu_inst_pe_1_5_4_U71 ( .A1(npu_inst_pe_1_5_4_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_5_4_n44), .ZN(npu_inst_pe_1_5_4_n66) );
  OAI21_X1 npu_inst_pe_1_5_4_U70 ( .B1(npu_inst_pe_1_5_4_n63), .B2(
        npu_inst_pe_1_5_4_n44), .A(npu_inst_pe_1_5_4_n66), .ZN(
        npu_inst_pe_1_5_4_n89) );
  NAND2_X1 npu_inst_pe_1_5_4_U69 ( .A1(npu_inst_pe_1_5_4_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_5_4_n44), .ZN(npu_inst_pe_1_5_4_n65) );
  OAI21_X1 npu_inst_pe_1_5_4_U68 ( .B1(npu_inst_pe_1_5_4_n61), .B2(
        npu_inst_pe_1_5_4_n44), .A(npu_inst_pe_1_5_4_n65), .ZN(
        npu_inst_pe_1_5_4_n88) );
  NAND2_X1 npu_inst_pe_1_5_4_U67 ( .A1(npu_inst_pe_1_5_4_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_5_4_n40), .ZN(npu_inst_pe_1_5_4_n64) );
  OAI21_X1 npu_inst_pe_1_5_4_U66 ( .B1(npu_inst_pe_1_5_4_n63), .B2(
        npu_inst_pe_1_5_4_n40), .A(npu_inst_pe_1_5_4_n64), .ZN(
        npu_inst_pe_1_5_4_n87) );
  NAND2_X1 npu_inst_pe_1_5_4_U65 ( .A1(npu_inst_pe_1_5_4_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_5_4_n40), .ZN(npu_inst_pe_1_5_4_n62) );
  OAI21_X1 npu_inst_pe_1_5_4_U64 ( .B1(npu_inst_pe_1_5_4_n61), .B2(
        npu_inst_pe_1_5_4_n40), .A(npu_inst_pe_1_5_4_n62), .ZN(
        npu_inst_pe_1_5_4_n86) );
  AND2_X1 npu_inst_pe_1_5_4_U63 ( .A1(npu_inst_pe_1_5_4_N93), .A2(npu_inst_n54), .ZN(npu_inst_int_data_y_5__4__0_) );
  AND2_X1 npu_inst_pe_1_5_4_U62 ( .A1(npu_inst_n54), .A2(npu_inst_pe_1_5_4_N94), .ZN(npu_inst_int_data_y_5__4__1_) );
  NOR3_X1 npu_inst_pe_1_5_4_U61 ( .A1(npu_inst_pe_1_5_4_n26), .A2(npu_inst_n54), .A3(npu_inst_int_ckg[19]), .ZN(npu_inst_pe_1_5_4_n85) );
  OR2_X1 npu_inst_pe_1_5_4_U60 ( .A1(npu_inst_pe_1_5_4_n85), .A2(
        npu_inst_pe_1_5_4_n2), .ZN(npu_inst_pe_1_5_4_N84) );
  AND2_X1 npu_inst_pe_1_5_4_U59 ( .A1(npu_inst_pe_1_5_4_int_q_acc_0_), .A2(
        npu_inst_pe_1_5_4_n1), .ZN(npu_inst_int_data_res_5__4__0_) );
  AND2_X1 npu_inst_pe_1_5_4_U58 ( .A1(npu_inst_pe_1_5_4_n2), .A2(
        npu_inst_pe_1_5_4_int_q_acc_7_), .ZN(npu_inst_int_data_res_5__4__7_)
         );
  AND2_X1 npu_inst_pe_1_5_4_U57 ( .A1(npu_inst_pe_1_5_4_int_q_acc_1_), .A2(
        npu_inst_pe_1_5_4_n1), .ZN(npu_inst_int_data_res_5__4__1_) );
  AND2_X1 npu_inst_pe_1_5_4_U56 ( .A1(npu_inst_pe_1_5_4_int_q_acc_2_), .A2(
        npu_inst_pe_1_5_4_n1), .ZN(npu_inst_int_data_res_5__4__2_) );
  AND2_X1 npu_inst_pe_1_5_4_U55 ( .A1(npu_inst_pe_1_5_4_int_q_acc_3_), .A2(
        npu_inst_pe_1_5_4_n2), .ZN(npu_inst_int_data_res_5__4__3_) );
  AND2_X1 npu_inst_pe_1_5_4_U54 ( .A1(npu_inst_pe_1_5_4_int_q_acc_4_), .A2(
        npu_inst_pe_1_5_4_n2), .ZN(npu_inst_int_data_res_5__4__4_) );
  AND2_X1 npu_inst_pe_1_5_4_U53 ( .A1(npu_inst_pe_1_5_4_int_q_acc_5_), .A2(
        npu_inst_pe_1_5_4_n2), .ZN(npu_inst_int_data_res_5__4__5_) );
  AND2_X1 npu_inst_pe_1_5_4_U52 ( .A1(npu_inst_pe_1_5_4_int_q_acc_6_), .A2(
        npu_inst_pe_1_5_4_n2), .ZN(npu_inst_int_data_res_5__4__6_) );
  AOI222_X1 npu_inst_pe_1_5_4_U51 ( .A1(npu_inst_int_data_res_6__4__0_), .A2(
        npu_inst_pe_1_5_4_n1), .B1(npu_inst_pe_1_5_4_N73), .B2(
        npu_inst_pe_1_5_4_n76), .C1(npu_inst_pe_1_5_4_N65), .C2(
        npu_inst_pe_1_5_4_n77), .ZN(npu_inst_pe_1_5_4_n84) );
  INV_X1 npu_inst_pe_1_5_4_U50 ( .A(npu_inst_pe_1_5_4_n84), .ZN(
        npu_inst_pe_1_5_4_n101) );
  AOI222_X1 npu_inst_pe_1_5_4_U49 ( .A1(npu_inst_int_data_res_6__4__7_), .A2(
        npu_inst_pe_1_5_4_n1), .B1(npu_inst_pe_1_5_4_N80), .B2(
        npu_inst_pe_1_5_4_n76), .C1(npu_inst_pe_1_5_4_N72), .C2(
        npu_inst_pe_1_5_4_n77), .ZN(npu_inst_pe_1_5_4_n75) );
  INV_X1 npu_inst_pe_1_5_4_U48 ( .A(npu_inst_pe_1_5_4_n75), .ZN(
        npu_inst_pe_1_5_4_n33) );
  AOI222_X1 npu_inst_pe_1_5_4_U47 ( .A1(npu_inst_int_data_res_6__4__1_), .A2(
        npu_inst_pe_1_5_4_n1), .B1(npu_inst_pe_1_5_4_N74), .B2(
        npu_inst_pe_1_5_4_n76), .C1(npu_inst_pe_1_5_4_N66), .C2(
        npu_inst_pe_1_5_4_n77), .ZN(npu_inst_pe_1_5_4_n83) );
  INV_X1 npu_inst_pe_1_5_4_U46 ( .A(npu_inst_pe_1_5_4_n83), .ZN(
        npu_inst_pe_1_5_4_n100) );
  AOI222_X1 npu_inst_pe_1_5_4_U45 ( .A1(npu_inst_int_data_res_6__4__2_), .A2(
        npu_inst_pe_1_5_4_n1), .B1(npu_inst_pe_1_5_4_N75), .B2(
        npu_inst_pe_1_5_4_n76), .C1(npu_inst_pe_1_5_4_N67), .C2(
        npu_inst_pe_1_5_4_n77), .ZN(npu_inst_pe_1_5_4_n82) );
  INV_X1 npu_inst_pe_1_5_4_U44 ( .A(npu_inst_pe_1_5_4_n82), .ZN(
        npu_inst_pe_1_5_4_n99) );
  AOI222_X1 npu_inst_pe_1_5_4_U43 ( .A1(npu_inst_int_data_res_6__4__3_), .A2(
        npu_inst_pe_1_5_4_n1), .B1(npu_inst_pe_1_5_4_N76), .B2(
        npu_inst_pe_1_5_4_n76), .C1(npu_inst_pe_1_5_4_N68), .C2(
        npu_inst_pe_1_5_4_n77), .ZN(npu_inst_pe_1_5_4_n81) );
  INV_X1 npu_inst_pe_1_5_4_U42 ( .A(npu_inst_pe_1_5_4_n81), .ZN(
        npu_inst_pe_1_5_4_n98) );
  AOI222_X1 npu_inst_pe_1_5_4_U41 ( .A1(npu_inst_int_data_res_6__4__4_), .A2(
        npu_inst_pe_1_5_4_n1), .B1(npu_inst_pe_1_5_4_N77), .B2(
        npu_inst_pe_1_5_4_n76), .C1(npu_inst_pe_1_5_4_N69), .C2(
        npu_inst_pe_1_5_4_n77), .ZN(npu_inst_pe_1_5_4_n80) );
  INV_X1 npu_inst_pe_1_5_4_U40 ( .A(npu_inst_pe_1_5_4_n80), .ZN(
        npu_inst_pe_1_5_4_n36) );
  AOI222_X1 npu_inst_pe_1_5_4_U39 ( .A1(npu_inst_int_data_res_6__4__5_), .A2(
        npu_inst_pe_1_5_4_n1), .B1(npu_inst_pe_1_5_4_N78), .B2(
        npu_inst_pe_1_5_4_n76), .C1(npu_inst_pe_1_5_4_N70), .C2(
        npu_inst_pe_1_5_4_n77), .ZN(npu_inst_pe_1_5_4_n79) );
  INV_X1 npu_inst_pe_1_5_4_U38 ( .A(npu_inst_pe_1_5_4_n79), .ZN(
        npu_inst_pe_1_5_4_n35) );
  AOI222_X1 npu_inst_pe_1_5_4_U37 ( .A1(npu_inst_int_data_res_6__4__6_), .A2(
        npu_inst_pe_1_5_4_n1), .B1(npu_inst_pe_1_5_4_N79), .B2(
        npu_inst_pe_1_5_4_n76), .C1(npu_inst_pe_1_5_4_N71), .C2(
        npu_inst_pe_1_5_4_n77), .ZN(npu_inst_pe_1_5_4_n78) );
  INV_X1 npu_inst_pe_1_5_4_U36 ( .A(npu_inst_pe_1_5_4_n78), .ZN(
        npu_inst_pe_1_5_4_n34) );
  INV_X1 npu_inst_pe_1_5_4_U35 ( .A(npu_inst_pe_1_5_4_int_data_1_), .ZN(
        npu_inst_pe_1_5_4_n14) );
  AND2_X1 npu_inst_pe_1_5_4_U34 ( .A1(npu_inst_int_data_x_5__4__1_), .A2(
        npu_inst_pe_1_5_4_int_q_weight_1_), .ZN(npu_inst_pe_1_5_4_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_5_4_U33 ( .A1(npu_inst_int_data_x_5__4__0_), .A2(
        npu_inst_pe_1_5_4_int_q_weight_1_), .ZN(npu_inst_pe_1_5_4_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_5_4_U32 ( .A1(npu_inst_n54), .A2(
        npu_inst_int_data_y_6__4__1_), .B1(npu_inst_pe_1_5_4_n3), .B2(
        npu_inst_int_data_x_5__5__1_), .ZN(npu_inst_pe_1_5_4_n63) );
  AOI22_X1 npu_inst_pe_1_5_4_U31 ( .A1(npu_inst_n54), .A2(
        npu_inst_int_data_y_6__4__0_), .B1(npu_inst_pe_1_5_4_n3), .B2(
        npu_inst_int_data_x_5__5__0_), .ZN(npu_inst_pe_1_5_4_n61) );
  INV_X1 npu_inst_pe_1_5_4_U30 ( .A(npu_inst_pe_1_5_4_int_data_0_), .ZN(
        npu_inst_pe_1_5_4_n13) );
  INV_X1 npu_inst_pe_1_5_4_U29 ( .A(npu_inst_n68), .ZN(npu_inst_pe_1_5_4_n5)
         );
  OR3_X1 npu_inst_pe_1_5_4_U28 ( .A1(npu_inst_pe_1_5_4_n6), .A2(
        npu_inst_pe_1_5_4_n8), .A3(npu_inst_pe_1_5_4_n5), .ZN(
        npu_inst_pe_1_5_4_n56) );
  OR3_X1 npu_inst_pe_1_5_4_U27 ( .A1(npu_inst_pe_1_5_4_n5), .A2(
        npu_inst_pe_1_5_4_n8), .A3(npu_inst_pe_1_5_4_n7), .ZN(
        npu_inst_pe_1_5_4_n48) );
  INV_X1 npu_inst_pe_1_5_4_U26 ( .A(npu_inst_pe_1_5_4_n5), .ZN(
        npu_inst_pe_1_5_4_n4) );
  INV_X1 npu_inst_pe_1_5_4_U25 ( .A(npu_inst_n123), .ZN(npu_inst_pe_1_5_4_n12)
         );
  OR3_X1 npu_inst_pe_1_5_4_U24 ( .A1(npu_inst_pe_1_5_4_n4), .A2(
        npu_inst_pe_1_5_4_n8), .A3(npu_inst_pe_1_5_4_n7), .ZN(
        npu_inst_pe_1_5_4_n52) );
  OR3_X1 npu_inst_pe_1_5_4_U23 ( .A1(npu_inst_pe_1_5_4_n6), .A2(
        npu_inst_pe_1_5_4_n8), .A3(npu_inst_pe_1_5_4_n4), .ZN(
        npu_inst_pe_1_5_4_n60) );
  NOR2_X1 npu_inst_pe_1_5_4_U22 ( .A1(npu_inst_pe_1_5_4_n60), .A2(
        npu_inst_pe_1_5_4_n3), .ZN(npu_inst_pe_1_5_4_n58) );
  NOR2_X1 npu_inst_pe_1_5_4_U21 ( .A1(npu_inst_pe_1_5_4_n56), .A2(
        npu_inst_pe_1_5_4_n3), .ZN(npu_inst_pe_1_5_4_n54) );
  NOR2_X1 npu_inst_pe_1_5_4_U20 ( .A1(npu_inst_pe_1_5_4_n52), .A2(
        npu_inst_pe_1_5_4_n3), .ZN(npu_inst_pe_1_5_4_n50) );
  NOR2_X1 npu_inst_pe_1_5_4_U19 ( .A1(npu_inst_pe_1_5_4_n48), .A2(
        npu_inst_pe_1_5_4_n3), .ZN(npu_inst_pe_1_5_4_n46) );
  NOR2_X1 npu_inst_pe_1_5_4_U18 ( .A1(npu_inst_pe_1_5_4_n40), .A2(
        npu_inst_pe_1_5_4_n3), .ZN(npu_inst_pe_1_5_4_n38) );
  NOR2_X1 npu_inst_pe_1_5_4_U17 ( .A1(npu_inst_pe_1_5_4_n44), .A2(
        npu_inst_pe_1_5_4_n3), .ZN(npu_inst_pe_1_5_4_n42) );
  BUF_X1 npu_inst_pe_1_5_4_U16 ( .A(npu_inst_n96), .Z(npu_inst_pe_1_5_4_n8) );
  BUF_X1 npu_inst_pe_1_5_4_U15 ( .A(npu_inst_pe_1_5_4_n12), .Z(
        npu_inst_pe_1_5_4_n11) );
  BUF_X1 npu_inst_pe_1_5_4_U14 ( .A(npu_inst_pe_1_5_4_n12), .Z(
        npu_inst_pe_1_5_4_n10) );
  BUF_X1 npu_inst_pe_1_5_4_U13 ( .A(npu_inst_pe_1_5_4_n12), .Z(
        npu_inst_pe_1_5_4_n9) );
  INV_X1 npu_inst_pe_1_5_4_U12 ( .A(npu_inst_pe_1_5_4_n38), .ZN(
        npu_inst_pe_1_5_4_n118) );
  INV_X1 npu_inst_pe_1_5_4_U11 ( .A(npu_inst_pe_1_5_4_n58), .ZN(
        npu_inst_pe_1_5_4_n114) );
  INV_X1 npu_inst_pe_1_5_4_U10 ( .A(npu_inst_pe_1_5_4_n54), .ZN(
        npu_inst_pe_1_5_4_n115) );
  INV_X1 npu_inst_pe_1_5_4_U9 ( .A(npu_inst_pe_1_5_4_n50), .ZN(
        npu_inst_pe_1_5_4_n116) );
  INV_X1 npu_inst_pe_1_5_4_U8 ( .A(npu_inst_pe_1_5_4_n46), .ZN(
        npu_inst_pe_1_5_4_n117) );
  INV_X1 npu_inst_pe_1_5_4_U7 ( .A(npu_inst_pe_1_5_4_n42), .ZN(
        npu_inst_pe_1_5_4_n119) );
  BUF_X1 npu_inst_pe_1_5_4_U6 ( .A(npu_inst_n16), .Z(npu_inst_pe_1_5_4_n2) );
  BUF_X1 npu_inst_pe_1_5_4_U5 ( .A(npu_inst_n16), .Z(npu_inst_pe_1_5_4_n1) );
  NOR2_X1 npu_inst_pe_1_5_4_U4 ( .A1(npu_inst_pe_1_5_4_int_q_weight_0_), .A2(
        npu_inst_pe_1_5_4_n1), .ZN(npu_inst_pe_1_5_4_n76) );
  NOR2_X1 npu_inst_pe_1_5_4_U3 ( .A1(npu_inst_pe_1_5_4_n27), .A2(
        npu_inst_pe_1_5_4_n1), .ZN(npu_inst_pe_1_5_4_n77) );
  FA_X1 npu_inst_pe_1_5_4_sub_77_U2_1 ( .A(npu_inst_pe_1_5_4_int_q_acc_1_), 
        .B(npu_inst_pe_1_5_4_n14), .CI(npu_inst_pe_1_5_4_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_5_4_sub_77_carry_2_), .S(npu_inst_pe_1_5_4_N66) );
  FA_X1 npu_inst_pe_1_5_4_add_79_U1_1 ( .A(npu_inst_pe_1_5_4_int_q_acc_1_), 
        .B(npu_inst_pe_1_5_4_int_data_1_), .CI(
        npu_inst_pe_1_5_4_add_79_carry_1_), .CO(
        npu_inst_pe_1_5_4_add_79_carry_2_), .S(npu_inst_pe_1_5_4_N74) );
  NAND3_X1 npu_inst_pe_1_5_4_U109 ( .A1(npu_inst_pe_1_5_4_n5), .A2(
        npu_inst_pe_1_5_4_n7), .A3(npu_inst_pe_1_5_4_n8), .ZN(
        npu_inst_pe_1_5_4_n44) );
  NAND3_X1 npu_inst_pe_1_5_4_U108 ( .A1(npu_inst_pe_1_5_4_n4), .A2(
        npu_inst_pe_1_5_4_n7), .A3(npu_inst_pe_1_5_4_n8), .ZN(
        npu_inst_pe_1_5_4_n40) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_5_4_n34), .CK(
        npu_inst_pe_1_5_4_net3281), .RN(npu_inst_pe_1_5_4_n9), .Q(
        npu_inst_pe_1_5_4_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_5_4_n35), .CK(
        npu_inst_pe_1_5_4_net3281), .RN(npu_inst_pe_1_5_4_n9), .Q(
        npu_inst_pe_1_5_4_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_5_4_n36), .CK(
        npu_inst_pe_1_5_4_net3281), .RN(npu_inst_pe_1_5_4_n9), .Q(
        npu_inst_pe_1_5_4_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_5_4_n98), .CK(
        npu_inst_pe_1_5_4_net3281), .RN(npu_inst_pe_1_5_4_n9), .Q(
        npu_inst_pe_1_5_4_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_5_4_n99), .CK(
        npu_inst_pe_1_5_4_net3281), .RN(npu_inst_pe_1_5_4_n9), .Q(
        npu_inst_pe_1_5_4_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_5_4_n100), 
        .CK(npu_inst_pe_1_5_4_net3281), .RN(npu_inst_pe_1_5_4_n9), .Q(
        npu_inst_pe_1_5_4_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_5_4_n33), .CK(
        npu_inst_pe_1_5_4_net3281), .RN(npu_inst_pe_1_5_4_n9), .Q(
        npu_inst_pe_1_5_4_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_5_4_n101), 
        .CK(npu_inst_pe_1_5_4_net3281), .RN(npu_inst_pe_1_5_4_n9), .Q(
        npu_inst_pe_1_5_4_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_weight_reg_0_ ( .D(npu_inst_n109), .CK(
        npu_inst_pe_1_5_4_net3287), .RN(npu_inst_pe_1_5_4_n9), .Q(
        npu_inst_pe_1_5_4_int_q_weight_0_), .QN(npu_inst_pe_1_5_4_n27) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_weight_reg_1_ ( .D(npu_inst_n115), .CK(
        npu_inst_pe_1_5_4_net3287), .RN(npu_inst_pe_1_5_4_n9), .Q(
        npu_inst_pe_1_5_4_int_q_weight_1_), .QN(npu_inst_pe_1_5_4_n26) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_5_4_n113), 
        .CK(npu_inst_pe_1_5_4_net3287), .RN(npu_inst_pe_1_5_4_n9), .Q(
        npu_inst_pe_1_5_4_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_5_4_n107), 
        .CK(npu_inst_pe_1_5_4_net3287), .RN(npu_inst_pe_1_5_4_n9), .Q(
        npu_inst_pe_1_5_4_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_5_4_n112), 
        .CK(npu_inst_pe_1_5_4_net3287), .RN(npu_inst_pe_1_5_4_n10), .Q(
        npu_inst_pe_1_5_4_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_5_4_n106), 
        .CK(npu_inst_pe_1_5_4_net3287), .RN(npu_inst_pe_1_5_4_n10), .Q(
        npu_inst_pe_1_5_4_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_5_4_n111), 
        .CK(npu_inst_pe_1_5_4_net3287), .RN(npu_inst_pe_1_5_4_n10), .Q(
        npu_inst_pe_1_5_4_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_5_4_n105), 
        .CK(npu_inst_pe_1_5_4_net3287), .RN(npu_inst_pe_1_5_4_n10), .Q(
        npu_inst_pe_1_5_4_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_5_4_n110), 
        .CK(npu_inst_pe_1_5_4_net3287), .RN(npu_inst_pe_1_5_4_n10), .Q(
        npu_inst_pe_1_5_4_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_5_4_n104), 
        .CK(npu_inst_pe_1_5_4_net3287), .RN(npu_inst_pe_1_5_4_n10), .Q(
        npu_inst_pe_1_5_4_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_5_4_n109), 
        .CK(npu_inst_pe_1_5_4_net3287), .RN(npu_inst_pe_1_5_4_n10), .Q(
        npu_inst_pe_1_5_4_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_5_4_n103), 
        .CK(npu_inst_pe_1_5_4_net3287), .RN(npu_inst_pe_1_5_4_n10), .Q(
        npu_inst_pe_1_5_4_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_5_4_n108), 
        .CK(npu_inst_pe_1_5_4_net3287), .RN(npu_inst_pe_1_5_4_n10), .Q(
        npu_inst_pe_1_5_4_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_5_4_n102), 
        .CK(npu_inst_pe_1_5_4_net3287), .RN(npu_inst_pe_1_5_4_n10), .Q(
        npu_inst_pe_1_5_4_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_5_4_n86), 
        .CK(npu_inst_pe_1_5_4_net3287), .RN(npu_inst_pe_1_5_4_n10), .Q(
        npu_inst_pe_1_5_4_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_5_4_n87), 
        .CK(npu_inst_pe_1_5_4_net3287), .RN(npu_inst_pe_1_5_4_n10), .Q(
        npu_inst_pe_1_5_4_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_5_4_n88), 
        .CK(npu_inst_pe_1_5_4_net3287), .RN(npu_inst_pe_1_5_4_n11), .Q(
        npu_inst_pe_1_5_4_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_5_4_n89), 
        .CK(npu_inst_pe_1_5_4_net3287), .RN(npu_inst_pe_1_5_4_n11), .Q(
        npu_inst_pe_1_5_4_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_5_4_n90), 
        .CK(npu_inst_pe_1_5_4_net3287), .RN(npu_inst_pe_1_5_4_n11), .Q(
        npu_inst_pe_1_5_4_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_5_4_n91), 
        .CK(npu_inst_pe_1_5_4_net3287), .RN(npu_inst_pe_1_5_4_n11), .Q(
        npu_inst_pe_1_5_4_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_5_4_n92), 
        .CK(npu_inst_pe_1_5_4_net3287), .RN(npu_inst_pe_1_5_4_n11), .Q(
        npu_inst_pe_1_5_4_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_5_4_n93), 
        .CK(npu_inst_pe_1_5_4_net3287), .RN(npu_inst_pe_1_5_4_n11), .Q(
        npu_inst_pe_1_5_4_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_5_4_n94), 
        .CK(npu_inst_pe_1_5_4_net3287), .RN(npu_inst_pe_1_5_4_n11), .Q(
        npu_inst_pe_1_5_4_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_5_4_n95), 
        .CK(npu_inst_pe_1_5_4_net3287), .RN(npu_inst_pe_1_5_4_n11), .Q(
        npu_inst_pe_1_5_4_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_5_4_n96), 
        .CK(npu_inst_pe_1_5_4_net3287), .RN(npu_inst_pe_1_5_4_n11), .Q(
        npu_inst_pe_1_5_4_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_5_4_n97), 
        .CK(npu_inst_pe_1_5_4_net3287), .RN(npu_inst_pe_1_5_4_n11), .Q(
        npu_inst_pe_1_5_4_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_5_4_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_5_4_N84), .SE(1'b0), .GCK(npu_inst_pe_1_5_4_net3281) );
  CLKGATETST_X1 npu_inst_pe_1_5_4_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n62), .SE(1'b0), .GCK(npu_inst_pe_1_5_4_net3287) );
  MUX2_X1 npu_inst_pe_1_5_5_U162 ( .A(npu_inst_pe_1_5_5_n32), .B(
        npu_inst_pe_1_5_5_n29), .S(npu_inst_pe_1_5_5_n8), .Z(
        npu_inst_pe_1_5_5_N93) );
  MUX2_X1 npu_inst_pe_1_5_5_U161 ( .A(npu_inst_pe_1_5_5_n31), .B(
        npu_inst_pe_1_5_5_n30), .S(npu_inst_pe_1_5_5_n6), .Z(
        npu_inst_pe_1_5_5_n32) );
  MUX2_X1 npu_inst_pe_1_5_5_U160 ( .A(npu_inst_pe_1_5_5_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_5_5_int_q_reg_v_1__0_), .S(npu_inst_pe_1_5_5_n4), .Z(
        npu_inst_pe_1_5_5_n31) );
  MUX2_X1 npu_inst_pe_1_5_5_U159 ( .A(npu_inst_pe_1_5_5_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_5_5_int_q_reg_v_3__0_), .S(npu_inst_pe_1_5_5_n4), .Z(
        npu_inst_pe_1_5_5_n30) );
  MUX2_X1 npu_inst_pe_1_5_5_U158 ( .A(npu_inst_pe_1_5_5_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_5_5_int_q_reg_v_5__0_), .S(npu_inst_pe_1_5_5_n4), .Z(
        npu_inst_pe_1_5_5_n29) );
  MUX2_X1 npu_inst_pe_1_5_5_U157 ( .A(npu_inst_pe_1_5_5_n28), .B(
        npu_inst_pe_1_5_5_n23), .S(npu_inst_pe_1_5_5_n8), .Z(
        npu_inst_pe_1_5_5_N94) );
  MUX2_X1 npu_inst_pe_1_5_5_U156 ( .A(npu_inst_pe_1_5_5_n25), .B(
        npu_inst_pe_1_5_5_n24), .S(npu_inst_pe_1_5_5_n6), .Z(
        npu_inst_pe_1_5_5_n28) );
  MUX2_X1 npu_inst_pe_1_5_5_U155 ( .A(npu_inst_pe_1_5_5_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_5_5_int_q_reg_v_1__1_), .S(npu_inst_pe_1_5_5_n4), .Z(
        npu_inst_pe_1_5_5_n25) );
  MUX2_X1 npu_inst_pe_1_5_5_U154 ( .A(npu_inst_pe_1_5_5_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_5_5_int_q_reg_v_3__1_), .S(npu_inst_pe_1_5_5_n4), .Z(
        npu_inst_pe_1_5_5_n24) );
  MUX2_X1 npu_inst_pe_1_5_5_U153 ( .A(npu_inst_pe_1_5_5_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_5_5_int_q_reg_v_5__1_), .S(npu_inst_pe_1_5_5_n4), .Z(
        npu_inst_pe_1_5_5_n23) );
  MUX2_X1 npu_inst_pe_1_5_5_U152 ( .A(npu_inst_pe_1_5_5_n22), .B(
        npu_inst_pe_1_5_5_n19), .S(npu_inst_pe_1_5_5_n8), .Z(
        npu_inst_int_data_x_5__5__1_) );
  MUX2_X1 npu_inst_pe_1_5_5_U151 ( .A(npu_inst_pe_1_5_5_n21), .B(
        npu_inst_pe_1_5_5_n20), .S(npu_inst_pe_1_5_5_n6), .Z(
        npu_inst_pe_1_5_5_n22) );
  MUX2_X1 npu_inst_pe_1_5_5_U150 ( .A(npu_inst_pe_1_5_5_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_5_5_int_q_reg_h_1__1_), .S(npu_inst_pe_1_5_5_n4), .Z(
        npu_inst_pe_1_5_5_n21) );
  MUX2_X1 npu_inst_pe_1_5_5_U149 ( .A(npu_inst_pe_1_5_5_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_5_5_int_q_reg_h_3__1_), .S(npu_inst_pe_1_5_5_n4), .Z(
        npu_inst_pe_1_5_5_n20) );
  MUX2_X1 npu_inst_pe_1_5_5_U148 ( .A(npu_inst_pe_1_5_5_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_5_5_int_q_reg_h_5__1_), .S(npu_inst_pe_1_5_5_n4), .Z(
        npu_inst_pe_1_5_5_n19) );
  MUX2_X1 npu_inst_pe_1_5_5_U147 ( .A(npu_inst_pe_1_5_5_n18), .B(
        npu_inst_pe_1_5_5_n15), .S(npu_inst_pe_1_5_5_n8), .Z(
        npu_inst_int_data_x_5__5__0_) );
  MUX2_X1 npu_inst_pe_1_5_5_U146 ( .A(npu_inst_pe_1_5_5_n17), .B(
        npu_inst_pe_1_5_5_n16), .S(npu_inst_pe_1_5_5_n6), .Z(
        npu_inst_pe_1_5_5_n18) );
  MUX2_X1 npu_inst_pe_1_5_5_U145 ( .A(npu_inst_pe_1_5_5_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_5_5_int_q_reg_h_1__0_), .S(npu_inst_pe_1_5_5_n4), .Z(
        npu_inst_pe_1_5_5_n17) );
  MUX2_X1 npu_inst_pe_1_5_5_U144 ( .A(npu_inst_pe_1_5_5_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_5_5_int_q_reg_h_3__0_), .S(npu_inst_pe_1_5_5_n4), .Z(
        npu_inst_pe_1_5_5_n16) );
  MUX2_X1 npu_inst_pe_1_5_5_U143 ( .A(npu_inst_pe_1_5_5_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_5_5_int_q_reg_h_5__0_), .S(npu_inst_pe_1_5_5_n4), .Z(
        npu_inst_pe_1_5_5_n15) );
  XOR2_X1 npu_inst_pe_1_5_5_U142 ( .A(npu_inst_pe_1_5_5_int_data_0_), .B(
        npu_inst_pe_1_5_5_int_q_acc_0_), .Z(npu_inst_pe_1_5_5_N73) );
  AND2_X1 npu_inst_pe_1_5_5_U141 ( .A1(npu_inst_pe_1_5_5_int_q_acc_0_), .A2(
        npu_inst_pe_1_5_5_int_data_0_), .ZN(npu_inst_pe_1_5_5_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_5_5_U140 ( .A(npu_inst_pe_1_5_5_int_q_acc_0_), .B(
        npu_inst_pe_1_5_5_n13), .ZN(npu_inst_pe_1_5_5_N65) );
  OR2_X1 npu_inst_pe_1_5_5_U139 ( .A1(npu_inst_pe_1_5_5_n13), .A2(
        npu_inst_pe_1_5_5_int_q_acc_0_), .ZN(npu_inst_pe_1_5_5_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_5_5_U138 ( .A(npu_inst_pe_1_5_5_int_q_acc_2_), .B(
        npu_inst_pe_1_5_5_add_79_carry_2_), .Z(npu_inst_pe_1_5_5_N75) );
  AND2_X1 npu_inst_pe_1_5_5_U137 ( .A1(npu_inst_pe_1_5_5_add_79_carry_2_), 
        .A2(npu_inst_pe_1_5_5_int_q_acc_2_), .ZN(
        npu_inst_pe_1_5_5_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_5_5_U136 ( .A(npu_inst_pe_1_5_5_int_q_acc_3_), .B(
        npu_inst_pe_1_5_5_add_79_carry_3_), .Z(npu_inst_pe_1_5_5_N76) );
  AND2_X1 npu_inst_pe_1_5_5_U135 ( .A1(npu_inst_pe_1_5_5_add_79_carry_3_), 
        .A2(npu_inst_pe_1_5_5_int_q_acc_3_), .ZN(
        npu_inst_pe_1_5_5_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_5_5_U134 ( .A(npu_inst_pe_1_5_5_int_q_acc_4_), .B(
        npu_inst_pe_1_5_5_add_79_carry_4_), .Z(npu_inst_pe_1_5_5_N77) );
  AND2_X1 npu_inst_pe_1_5_5_U133 ( .A1(npu_inst_pe_1_5_5_add_79_carry_4_), 
        .A2(npu_inst_pe_1_5_5_int_q_acc_4_), .ZN(
        npu_inst_pe_1_5_5_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_5_5_U132 ( .A(npu_inst_pe_1_5_5_int_q_acc_5_), .B(
        npu_inst_pe_1_5_5_add_79_carry_5_), .Z(npu_inst_pe_1_5_5_N78) );
  AND2_X1 npu_inst_pe_1_5_5_U131 ( .A1(npu_inst_pe_1_5_5_add_79_carry_5_), 
        .A2(npu_inst_pe_1_5_5_int_q_acc_5_), .ZN(
        npu_inst_pe_1_5_5_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_5_5_U130 ( .A(npu_inst_pe_1_5_5_int_q_acc_6_), .B(
        npu_inst_pe_1_5_5_add_79_carry_6_), .Z(npu_inst_pe_1_5_5_N79) );
  AND2_X1 npu_inst_pe_1_5_5_U129 ( .A1(npu_inst_pe_1_5_5_add_79_carry_6_), 
        .A2(npu_inst_pe_1_5_5_int_q_acc_6_), .ZN(
        npu_inst_pe_1_5_5_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_5_5_U128 ( .A(npu_inst_pe_1_5_5_int_q_acc_7_), .B(
        npu_inst_pe_1_5_5_add_79_carry_7_), .Z(npu_inst_pe_1_5_5_N80) );
  XNOR2_X1 npu_inst_pe_1_5_5_U127 ( .A(npu_inst_pe_1_5_5_sub_77_carry_2_), .B(
        npu_inst_pe_1_5_5_int_q_acc_2_), .ZN(npu_inst_pe_1_5_5_N67) );
  OR2_X1 npu_inst_pe_1_5_5_U126 ( .A1(npu_inst_pe_1_5_5_int_q_acc_2_), .A2(
        npu_inst_pe_1_5_5_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_5_5_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_5_5_U125 ( .A(npu_inst_pe_1_5_5_sub_77_carry_3_), .B(
        npu_inst_pe_1_5_5_int_q_acc_3_), .ZN(npu_inst_pe_1_5_5_N68) );
  OR2_X1 npu_inst_pe_1_5_5_U124 ( .A1(npu_inst_pe_1_5_5_int_q_acc_3_), .A2(
        npu_inst_pe_1_5_5_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_5_5_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_5_5_U123 ( .A(npu_inst_pe_1_5_5_sub_77_carry_4_), .B(
        npu_inst_pe_1_5_5_int_q_acc_4_), .ZN(npu_inst_pe_1_5_5_N69) );
  OR2_X1 npu_inst_pe_1_5_5_U122 ( .A1(npu_inst_pe_1_5_5_int_q_acc_4_), .A2(
        npu_inst_pe_1_5_5_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_5_5_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_5_5_U121 ( .A(npu_inst_pe_1_5_5_sub_77_carry_5_), .B(
        npu_inst_pe_1_5_5_int_q_acc_5_), .ZN(npu_inst_pe_1_5_5_N70) );
  OR2_X1 npu_inst_pe_1_5_5_U120 ( .A1(npu_inst_pe_1_5_5_int_q_acc_5_), .A2(
        npu_inst_pe_1_5_5_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_5_5_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_5_5_U119 ( .A(npu_inst_pe_1_5_5_sub_77_carry_6_), .B(
        npu_inst_pe_1_5_5_int_q_acc_6_), .ZN(npu_inst_pe_1_5_5_N71) );
  OR2_X1 npu_inst_pe_1_5_5_U118 ( .A1(npu_inst_pe_1_5_5_int_q_acc_6_), .A2(
        npu_inst_pe_1_5_5_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_5_5_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_5_5_U117 ( .A(npu_inst_pe_1_5_5_int_q_acc_7_), .B(
        npu_inst_pe_1_5_5_sub_77_carry_7_), .ZN(npu_inst_pe_1_5_5_N72) );
  INV_X1 npu_inst_pe_1_5_5_U116 ( .A(npu_inst_n76), .ZN(npu_inst_pe_1_5_5_n7)
         );
  INV_X1 npu_inst_pe_1_5_5_U115 ( .A(npu_inst_pe_1_5_5_n7), .ZN(
        npu_inst_pe_1_5_5_n6) );
  INV_X1 npu_inst_pe_1_5_5_U114 ( .A(npu_inst_n54), .ZN(npu_inst_pe_1_5_5_n3)
         );
  AOI22_X1 npu_inst_pe_1_5_5_U113 ( .A1(npu_inst_int_data_y_6__5__0_), .A2(
        npu_inst_pe_1_5_5_n58), .B1(npu_inst_pe_1_5_5_n114), .B2(
        npu_inst_pe_1_5_5_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_5_5_n57) );
  INV_X1 npu_inst_pe_1_5_5_U112 ( .A(npu_inst_pe_1_5_5_n57), .ZN(
        npu_inst_pe_1_5_5_n108) );
  AOI22_X1 npu_inst_pe_1_5_5_U111 ( .A1(npu_inst_int_data_y_6__5__0_), .A2(
        npu_inst_pe_1_5_5_n54), .B1(npu_inst_pe_1_5_5_n115), .B2(
        npu_inst_pe_1_5_5_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_5_5_n53) );
  INV_X1 npu_inst_pe_1_5_5_U110 ( .A(npu_inst_pe_1_5_5_n53), .ZN(
        npu_inst_pe_1_5_5_n109) );
  AOI22_X1 npu_inst_pe_1_5_5_U107 ( .A1(npu_inst_int_data_y_6__5__0_), .A2(
        npu_inst_pe_1_5_5_n50), .B1(npu_inst_pe_1_5_5_n116), .B2(
        npu_inst_pe_1_5_5_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_5_5_n49) );
  INV_X1 npu_inst_pe_1_5_5_U106 ( .A(npu_inst_pe_1_5_5_n49), .ZN(
        npu_inst_pe_1_5_5_n110) );
  AOI22_X1 npu_inst_pe_1_5_5_U105 ( .A1(npu_inst_int_data_y_6__5__0_), .A2(
        npu_inst_pe_1_5_5_n46), .B1(npu_inst_pe_1_5_5_n117), .B2(
        npu_inst_pe_1_5_5_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_5_5_n45) );
  INV_X1 npu_inst_pe_1_5_5_U104 ( .A(npu_inst_pe_1_5_5_n45), .ZN(
        npu_inst_pe_1_5_5_n111) );
  AOI22_X1 npu_inst_pe_1_5_5_U103 ( .A1(npu_inst_int_data_y_6__5__0_), .A2(
        npu_inst_pe_1_5_5_n42), .B1(npu_inst_pe_1_5_5_n119), .B2(
        npu_inst_pe_1_5_5_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_5_5_n41) );
  INV_X1 npu_inst_pe_1_5_5_U102 ( .A(npu_inst_pe_1_5_5_n41), .ZN(
        npu_inst_pe_1_5_5_n112) );
  AOI22_X1 npu_inst_pe_1_5_5_U101 ( .A1(npu_inst_int_data_y_6__5__1_), .A2(
        npu_inst_pe_1_5_5_n58), .B1(npu_inst_pe_1_5_5_n114), .B2(
        npu_inst_pe_1_5_5_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_5_5_n59) );
  INV_X1 npu_inst_pe_1_5_5_U100 ( .A(npu_inst_pe_1_5_5_n59), .ZN(
        npu_inst_pe_1_5_5_n102) );
  AOI22_X1 npu_inst_pe_1_5_5_U99 ( .A1(npu_inst_int_data_y_6__5__1_), .A2(
        npu_inst_pe_1_5_5_n54), .B1(npu_inst_pe_1_5_5_n115), .B2(
        npu_inst_pe_1_5_5_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_5_5_n55) );
  INV_X1 npu_inst_pe_1_5_5_U98 ( .A(npu_inst_pe_1_5_5_n55), .ZN(
        npu_inst_pe_1_5_5_n103) );
  AOI22_X1 npu_inst_pe_1_5_5_U97 ( .A1(npu_inst_int_data_y_6__5__1_), .A2(
        npu_inst_pe_1_5_5_n50), .B1(npu_inst_pe_1_5_5_n116), .B2(
        npu_inst_pe_1_5_5_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_5_5_n51) );
  INV_X1 npu_inst_pe_1_5_5_U96 ( .A(npu_inst_pe_1_5_5_n51), .ZN(
        npu_inst_pe_1_5_5_n104) );
  AOI22_X1 npu_inst_pe_1_5_5_U95 ( .A1(npu_inst_int_data_y_6__5__1_), .A2(
        npu_inst_pe_1_5_5_n46), .B1(npu_inst_pe_1_5_5_n117), .B2(
        npu_inst_pe_1_5_5_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_5_5_n47) );
  INV_X1 npu_inst_pe_1_5_5_U94 ( .A(npu_inst_pe_1_5_5_n47), .ZN(
        npu_inst_pe_1_5_5_n105) );
  AOI22_X1 npu_inst_pe_1_5_5_U93 ( .A1(npu_inst_int_data_y_6__5__1_), .A2(
        npu_inst_pe_1_5_5_n42), .B1(npu_inst_pe_1_5_5_n119), .B2(
        npu_inst_pe_1_5_5_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_5_5_n43) );
  INV_X1 npu_inst_pe_1_5_5_U92 ( .A(npu_inst_pe_1_5_5_n43), .ZN(
        npu_inst_pe_1_5_5_n106) );
  AOI22_X1 npu_inst_pe_1_5_5_U91 ( .A1(npu_inst_pe_1_5_5_n38), .A2(
        npu_inst_int_data_y_6__5__1_), .B1(npu_inst_pe_1_5_5_n118), .B2(
        npu_inst_pe_1_5_5_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_5_5_n39) );
  INV_X1 npu_inst_pe_1_5_5_U90 ( .A(npu_inst_pe_1_5_5_n39), .ZN(
        npu_inst_pe_1_5_5_n107) );
  AOI22_X1 npu_inst_pe_1_5_5_U89 ( .A1(npu_inst_pe_1_5_5_n38), .A2(
        npu_inst_int_data_y_6__5__0_), .B1(npu_inst_pe_1_5_5_n118), .B2(
        npu_inst_pe_1_5_5_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_5_5_n37) );
  INV_X1 npu_inst_pe_1_5_5_U88 ( .A(npu_inst_pe_1_5_5_n37), .ZN(
        npu_inst_pe_1_5_5_n113) );
  NAND2_X1 npu_inst_pe_1_5_5_U87 ( .A1(npu_inst_pe_1_5_5_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_5_5_n60), .ZN(npu_inst_pe_1_5_5_n74) );
  OAI21_X1 npu_inst_pe_1_5_5_U86 ( .B1(npu_inst_pe_1_5_5_n63), .B2(
        npu_inst_pe_1_5_5_n60), .A(npu_inst_pe_1_5_5_n74), .ZN(
        npu_inst_pe_1_5_5_n97) );
  NAND2_X1 npu_inst_pe_1_5_5_U85 ( .A1(npu_inst_pe_1_5_5_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_5_5_n60), .ZN(npu_inst_pe_1_5_5_n73) );
  OAI21_X1 npu_inst_pe_1_5_5_U84 ( .B1(npu_inst_pe_1_5_5_n61), .B2(
        npu_inst_pe_1_5_5_n60), .A(npu_inst_pe_1_5_5_n73), .ZN(
        npu_inst_pe_1_5_5_n96) );
  NAND2_X1 npu_inst_pe_1_5_5_U83 ( .A1(npu_inst_pe_1_5_5_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_5_5_n56), .ZN(npu_inst_pe_1_5_5_n72) );
  OAI21_X1 npu_inst_pe_1_5_5_U82 ( .B1(npu_inst_pe_1_5_5_n63), .B2(
        npu_inst_pe_1_5_5_n56), .A(npu_inst_pe_1_5_5_n72), .ZN(
        npu_inst_pe_1_5_5_n95) );
  NAND2_X1 npu_inst_pe_1_5_5_U81 ( .A1(npu_inst_pe_1_5_5_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_5_5_n56), .ZN(npu_inst_pe_1_5_5_n71) );
  OAI21_X1 npu_inst_pe_1_5_5_U80 ( .B1(npu_inst_pe_1_5_5_n61), .B2(
        npu_inst_pe_1_5_5_n56), .A(npu_inst_pe_1_5_5_n71), .ZN(
        npu_inst_pe_1_5_5_n94) );
  NAND2_X1 npu_inst_pe_1_5_5_U79 ( .A1(npu_inst_pe_1_5_5_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_5_5_n52), .ZN(npu_inst_pe_1_5_5_n70) );
  OAI21_X1 npu_inst_pe_1_5_5_U78 ( .B1(npu_inst_pe_1_5_5_n63), .B2(
        npu_inst_pe_1_5_5_n52), .A(npu_inst_pe_1_5_5_n70), .ZN(
        npu_inst_pe_1_5_5_n93) );
  NAND2_X1 npu_inst_pe_1_5_5_U77 ( .A1(npu_inst_pe_1_5_5_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_5_5_n52), .ZN(npu_inst_pe_1_5_5_n69) );
  OAI21_X1 npu_inst_pe_1_5_5_U76 ( .B1(npu_inst_pe_1_5_5_n61), .B2(
        npu_inst_pe_1_5_5_n52), .A(npu_inst_pe_1_5_5_n69), .ZN(
        npu_inst_pe_1_5_5_n92) );
  NAND2_X1 npu_inst_pe_1_5_5_U75 ( .A1(npu_inst_pe_1_5_5_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_5_5_n48), .ZN(npu_inst_pe_1_5_5_n68) );
  OAI21_X1 npu_inst_pe_1_5_5_U74 ( .B1(npu_inst_pe_1_5_5_n63), .B2(
        npu_inst_pe_1_5_5_n48), .A(npu_inst_pe_1_5_5_n68), .ZN(
        npu_inst_pe_1_5_5_n91) );
  NAND2_X1 npu_inst_pe_1_5_5_U73 ( .A1(npu_inst_pe_1_5_5_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_5_5_n48), .ZN(npu_inst_pe_1_5_5_n67) );
  OAI21_X1 npu_inst_pe_1_5_5_U72 ( .B1(npu_inst_pe_1_5_5_n61), .B2(
        npu_inst_pe_1_5_5_n48), .A(npu_inst_pe_1_5_5_n67), .ZN(
        npu_inst_pe_1_5_5_n90) );
  NAND2_X1 npu_inst_pe_1_5_5_U71 ( .A1(npu_inst_pe_1_5_5_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_5_5_n44), .ZN(npu_inst_pe_1_5_5_n66) );
  OAI21_X1 npu_inst_pe_1_5_5_U70 ( .B1(npu_inst_pe_1_5_5_n63), .B2(
        npu_inst_pe_1_5_5_n44), .A(npu_inst_pe_1_5_5_n66), .ZN(
        npu_inst_pe_1_5_5_n89) );
  NAND2_X1 npu_inst_pe_1_5_5_U69 ( .A1(npu_inst_pe_1_5_5_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_5_5_n44), .ZN(npu_inst_pe_1_5_5_n65) );
  OAI21_X1 npu_inst_pe_1_5_5_U68 ( .B1(npu_inst_pe_1_5_5_n61), .B2(
        npu_inst_pe_1_5_5_n44), .A(npu_inst_pe_1_5_5_n65), .ZN(
        npu_inst_pe_1_5_5_n88) );
  NAND2_X1 npu_inst_pe_1_5_5_U67 ( .A1(npu_inst_pe_1_5_5_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_5_5_n40), .ZN(npu_inst_pe_1_5_5_n64) );
  OAI21_X1 npu_inst_pe_1_5_5_U66 ( .B1(npu_inst_pe_1_5_5_n63), .B2(
        npu_inst_pe_1_5_5_n40), .A(npu_inst_pe_1_5_5_n64), .ZN(
        npu_inst_pe_1_5_5_n87) );
  NAND2_X1 npu_inst_pe_1_5_5_U65 ( .A1(npu_inst_pe_1_5_5_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_5_5_n40), .ZN(npu_inst_pe_1_5_5_n62) );
  OAI21_X1 npu_inst_pe_1_5_5_U64 ( .B1(npu_inst_pe_1_5_5_n61), .B2(
        npu_inst_pe_1_5_5_n40), .A(npu_inst_pe_1_5_5_n62), .ZN(
        npu_inst_pe_1_5_5_n86) );
  AND2_X1 npu_inst_pe_1_5_5_U63 ( .A1(npu_inst_pe_1_5_5_N93), .A2(npu_inst_n54), .ZN(npu_inst_int_data_y_5__5__0_) );
  AND2_X1 npu_inst_pe_1_5_5_U62 ( .A1(npu_inst_n54), .A2(npu_inst_pe_1_5_5_N94), .ZN(npu_inst_int_data_y_5__5__1_) );
  NOR3_X1 npu_inst_pe_1_5_5_U61 ( .A1(npu_inst_pe_1_5_5_n26), .A2(npu_inst_n54), .A3(npu_inst_int_ckg[18]), .ZN(npu_inst_pe_1_5_5_n85) );
  OR2_X1 npu_inst_pe_1_5_5_U60 ( .A1(npu_inst_pe_1_5_5_n85), .A2(
        npu_inst_pe_1_5_5_n2), .ZN(npu_inst_pe_1_5_5_N84) );
  AND2_X1 npu_inst_pe_1_5_5_U59 ( .A1(npu_inst_pe_1_5_5_int_q_acc_0_), .A2(
        npu_inst_pe_1_5_5_n1), .ZN(npu_inst_int_data_res_5__5__0_) );
  AND2_X1 npu_inst_pe_1_5_5_U58 ( .A1(npu_inst_pe_1_5_5_n2), .A2(
        npu_inst_pe_1_5_5_int_q_acc_7_), .ZN(npu_inst_int_data_res_5__5__7_)
         );
  AND2_X1 npu_inst_pe_1_5_5_U57 ( .A1(npu_inst_pe_1_5_5_int_q_acc_1_), .A2(
        npu_inst_pe_1_5_5_n1), .ZN(npu_inst_int_data_res_5__5__1_) );
  AND2_X1 npu_inst_pe_1_5_5_U56 ( .A1(npu_inst_pe_1_5_5_int_q_acc_2_), .A2(
        npu_inst_pe_1_5_5_n1), .ZN(npu_inst_int_data_res_5__5__2_) );
  AND2_X1 npu_inst_pe_1_5_5_U55 ( .A1(npu_inst_pe_1_5_5_int_q_acc_3_), .A2(
        npu_inst_pe_1_5_5_n2), .ZN(npu_inst_int_data_res_5__5__3_) );
  AND2_X1 npu_inst_pe_1_5_5_U54 ( .A1(npu_inst_pe_1_5_5_int_q_acc_4_), .A2(
        npu_inst_pe_1_5_5_n2), .ZN(npu_inst_int_data_res_5__5__4_) );
  AND2_X1 npu_inst_pe_1_5_5_U53 ( .A1(npu_inst_pe_1_5_5_int_q_acc_5_), .A2(
        npu_inst_pe_1_5_5_n2), .ZN(npu_inst_int_data_res_5__5__5_) );
  AND2_X1 npu_inst_pe_1_5_5_U52 ( .A1(npu_inst_pe_1_5_5_int_q_acc_6_), .A2(
        npu_inst_pe_1_5_5_n2), .ZN(npu_inst_int_data_res_5__5__6_) );
  AOI222_X1 npu_inst_pe_1_5_5_U51 ( .A1(npu_inst_int_data_res_6__5__0_), .A2(
        npu_inst_pe_1_5_5_n1), .B1(npu_inst_pe_1_5_5_N73), .B2(
        npu_inst_pe_1_5_5_n76), .C1(npu_inst_pe_1_5_5_N65), .C2(
        npu_inst_pe_1_5_5_n77), .ZN(npu_inst_pe_1_5_5_n84) );
  INV_X1 npu_inst_pe_1_5_5_U50 ( .A(npu_inst_pe_1_5_5_n84), .ZN(
        npu_inst_pe_1_5_5_n101) );
  AOI222_X1 npu_inst_pe_1_5_5_U49 ( .A1(npu_inst_int_data_res_6__5__7_), .A2(
        npu_inst_pe_1_5_5_n1), .B1(npu_inst_pe_1_5_5_N80), .B2(
        npu_inst_pe_1_5_5_n76), .C1(npu_inst_pe_1_5_5_N72), .C2(
        npu_inst_pe_1_5_5_n77), .ZN(npu_inst_pe_1_5_5_n75) );
  INV_X1 npu_inst_pe_1_5_5_U48 ( .A(npu_inst_pe_1_5_5_n75), .ZN(
        npu_inst_pe_1_5_5_n33) );
  AOI222_X1 npu_inst_pe_1_5_5_U47 ( .A1(npu_inst_int_data_res_6__5__1_), .A2(
        npu_inst_pe_1_5_5_n1), .B1(npu_inst_pe_1_5_5_N74), .B2(
        npu_inst_pe_1_5_5_n76), .C1(npu_inst_pe_1_5_5_N66), .C2(
        npu_inst_pe_1_5_5_n77), .ZN(npu_inst_pe_1_5_5_n83) );
  INV_X1 npu_inst_pe_1_5_5_U46 ( .A(npu_inst_pe_1_5_5_n83), .ZN(
        npu_inst_pe_1_5_5_n100) );
  AOI222_X1 npu_inst_pe_1_5_5_U45 ( .A1(npu_inst_int_data_res_6__5__2_), .A2(
        npu_inst_pe_1_5_5_n1), .B1(npu_inst_pe_1_5_5_N75), .B2(
        npu_inst_pe_1_5_5_n76), .C1(npu_inst_pe_1_5_5_N67), .C2(
        npu_inst_pe_1_5_5_n77), .ZN(npu_inst_pe_1_5_5_n82) );
  INV_X1 npu_inst_pe_1_5_5_U44 ( .A(npu_inst_pe_1_5_5_n82), .ZN(
        npu_inst_pe_1_5_5_n99) );
  AOI222_X1 npu_inst_pe_1_5_5_U43 ( .A1(npu_inst_int_data_res_6__5__3_), .A2(
        npu_inst_pe_1_5_5_n1), .B1(npu_inst_pe_1_5_5_N76), .B2(
        npu_inst_pe_1_5_5_n76), .C1(npu_inst_pe_1_5_5_N68), .C2(
        npu_inst_pe_1_5_5_n77), .ZN(npu_inst_pe_1_5_5_n81) );
  INV_X1 npu_inst_pe_1_5_5_U42 ( .A(npu_inst_pe_1_5_5_n81), .ZN(
        npu_inst_pe_1_5_5_n98) );
  AOI222_X1 npu_inst_pe_1_5_5_U41 ( .A1(npu_inst_int_data_res_6__5__4_), .A2(
        npu_inst_pe_1_5_5_n1), .B1(npu_inst_pe_1_5_5_N77), .B2(
        npu_inst_pe_1_5_5_n76), .C1(npu_inst_pe_1_5_5_N69), .C2(
        npu_inst_pe_1_5_5_n77), .ZN(npu_inst_pe_1_5_5_n80) );
  INV_X1 npu_inst_pe_1_5_5_U40 ( .A(npu_inst_pe_1_5_5_n80), .ZN(
        npu_inst_pe_1_5_5_n36) );
  AOI222_X1 npu_inst_pe_1_5_5_U39 ( .A1(npu_inst_int_data_res_6__5__5_), .A2(
        npu_inst_pe_1_5_5_n1), .B1(npu_inst_pe_1_5_5_N78), .B2(
        npu_inst_pe_1_5_5_n76), .C1(npu_inst_pe_1_5_5_N70), .C2(
        npu_inst_pe_1_5_5_n77), .ZN(npu_inst_pe_1_5_5_n79) );
  INV_X1 npu_inst_pe_1_5_5_U38 ( .A(npu_inst_pe_1_5_5_n79), .ZN(
        npu_inst_pe_1_5_5_n35) );
  AOI222_X1 npu_inst_pe_1_5_5_U37 ( .A1(npu_inst_int_data_res_6__5__6_), .A2(
        npu_inst_pe_1_5_5_n1), .B1(npu_inst_pe_1_5_5_N79), .B2(
        npu_inst_pe_1_5_5_n76), .C1(npu_inst_pe_1_5_5_N71), .C2(
        npu_inst_pe_1_5_5_n77), .ZN(npu_inst_pe_1_5_5_n78) );
  INV_X1 npu_inst_pe_1_5_5_U36 ( .A(npu_inst_pe_1_5_5_n78), .ZN(
        npu_inst_pe_1_5_5_n34) );
  INV_X1 npu_inst_pe_1_5_5_U35 ( .A(npu_inst_pe_1_5_5_int_data_1_), .ZN(
        npu_inst_pe_1_5_5_n14) );
  AND2_X1 npu_inst_pe_1_5_5_U34 ( .A1(npu_inst_int_data_x_5__5__1_), .A2(
        npu_inst_pe_1_5_5_int_q_weight_1_), .ZN(npu_inst_pe_1_5_5_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_5_5_U33 ( .A1(npu_inst_int_data_x_5__5__0_), .A2(
        npu_inst_pe_1_5_5_int_q_weight_1_), .ZN(npu_inst_pe_1_5_5_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_5_5_U32 ( .A1(npu_inst_n54), .A2(
        npu_inst_int_data_y_6__5__1_), .B1(npu_inst_pe_1_5_5_n3), .B2(
        npu_inst_int_data_x_5__6__1_), .ZN(npu_inst_pe_1_5_5_n63) );
  AOI22_X1 npu_inst_pe_1_5_5_U31 ( .A1(npu_inst_n54), .A2(
        npu_inst_int_data_y_6__5__0_), .B1(npu_inst_pe_1_5_5_n3), .B2(
        npu_inst_int_data_x_5__6__0_), .ZN(npu_inst_pe_1_5_5_n61) );
  INV_X1 npu_inst_pe_1_5_5_U30 ( .A(npu_inst_pe_1_5_5_int_data_0_), .ZN(
        npu_inst_pe_1_5_5_n13) );
  INV_X1 npu_inst_pe_1_5_5_U29 ( .A(npu_inst_n68), .ZN(npu_inst_pe_1_5_5_n5)
         );
  OR3_X1 npu_inst_pe_1_5_5_U28 ( .A1(npu_inst_pe_1_5_5_n6), .A2(
        npu_inst_pe_1_5_5_n8), .A3(npu_inst_pe_1_5_5_n5), .ZN(
        npu_inst_pe_1_5_5_n56) );
  OR3_X1 npu_inst_pe_1_5_5_U27 ( .A1(npu_inst_pe_1_5_5_n5), .A2(
        npu_inst_pe_1_5_5_n8), .A3(npu_inst_pe_1_5_5_n7), .ZN(
        npu_inst_pe_1_5_5_n48) );
  INV_X1 npu_inst_pe_1_5_5_U26 ( .A(npu_inst_pe_1_5_5_n5), .ZN(
        npu_inst_pe_1_5_5_n4) );
  INV_X1 npu_inst_pe_1_5_5_U25 ( .A(npu_inst_n123), .ZN(npu_inst_pe_1_5_5_n12)
         );
  OR3_X1 npu_inst_pe_1_5_5_U24 ( .A1(npu_inst_pe_1_5_5_n4), .A2(
        npu_inst_pe_1_5_5_n8), .A3(npu_inst_pe_1_5_5_n7), .ZN(
        npu_inst_pe_1_5_5_n52) );
  OR3_X1 npu_inst_pe_1_5_5_U23 ( .A1(npu_inst_pe_1_5_5_n6), .A2(
        npu_inst_pe_1_5_5_n8), .A3(npu_inst_pe_1_5_5_n4), .ZN(
        npu_inst_pe_1_5_5_n60) );
  NOR2_X1 npu_inst_pe_1_5_5_U22 ( .A1(npu_inst_pe_1_5_5_n60), .A2(
        npu_inst_pe_1_5_5_n3), .ZN(npu_inst_pe_1_5_5_n58) );
  NOR2_X1 npu_inst_pe_1_5_5_U21 ( .A1(npu_inst_pe_1_5_5_n56), .A2(
        npu_inst_pe_1_5_5_n3), .ZN(npu_inst_pe_1_5_5_n54) );
  NOR2_X1 npu_inst_pe_1_5_5_U20 ( .A1(npu_inst_pe_1_5_5_n52), .A2(
        npu_inst_pe_1_5_5_n3), .ZN(npu_inst_pe_1_5_5_n50) );
  NOR2_X1 npu_inst_pe_1_5_5_U19 ( .A1(npu_inst_pe_1_5_5_n48), .A2(
        npu_inst_pe_1_5_5_n3), .ZN(npu_inst_pe_1_5_5_n46) );
  NOR2_X1 npu_inst_pe_1_5_5_U18 ( .A1(npu_inst_pe_1_5_5_n40), .A2(
        npu_inst_pe_1_5_5_n3), .ZN(npu_inst_pe_1_5_5_n38) );
  NOR2_X1 npu_inst_pe_1_5_5_U17 ( .A1(npu_inst_pe_1_5_5_n44), .A2(
        npu_inst_pe_1_5_5_n3), .ZN(npu_inst_pe_1_5_5_n42) );
  BUF_X1 npu_inst_pe_1_5_5_U16 ( .A(npu_inst_n96), .Z(npu_inst_pe_1_5_5_n8) );
  BUF_X1 npu_inst_pe_1_5_5_U15 ( .A(npu_inst_pe_1_5_5_n12), .Z(
        npu_inst_pe_1_5_5_n11) );
  BUF_X1 npu_inst_pe_1_5_5_U14 ( .A(npu_inst_pe_1_5_5_n12), .Z(
        npu_inst_pe_1_5_5_n10) );
  BUF_X1 npu_inst_pe_1_5_5_U13 ( .A(npu_inst_pe_1_5_5_n12), .Z(
        npu_inst_pe_1_5_5_n9) );
  INV_X1 npu_inst_pe_1_5_5_U12 ( .A(npu_inst_pe_1_5_5_n38), .ZN(
        npu_inst_pe_1_5_5_n118) );
  INV_X1 npu_inst_pe_1_5_5_U11 ( .A(npu_inst_pe_1_5_5_n58), .ZN(
        npu_inst_pe_1_5_5_n114) );
  INV_X1 npu_inst_pe_1_5_5_U10 ( .A(npu_inst_pe_1_5_5_n54), .ZN(
        npu_inst_pe_1_5_5_n115) );
  INV_X1 npu_inst_pe_1_5_5_U9 ( .A(npu_inst_pe_1_5_5_n50), .ZN(
        npu_inst_pe_1_5_5_n116) );
  INV_X1 npu_inst_pe_1_5_5_U8 ( .A(npu_inst_pe_1_5_5_n46), .ZN(
        npu_inst_pe_1_5_5_n117) );
  INV_X1 npu_inst_pe_1_5_5_U7 ( .A(npu_inst_pe_1_5_5_n42), .ZN(
        npu_inst_pe_1_5_5_n119) );
  BUF_X1 npu_inst_pe_1_5_5_U6 ( .A(npu_inst_n16), .Z(npu_inst_pe_1_5_5_n2) );
  BUF_X1 npu_inst_pe_1_5_5_U5 ( .A(npu_inst_n16), .Z(npu_inst_pe_1_5_5_n1) );
  NOR2_X1 npu_inst_pe_1_5_5_U4 ( .A1(npu_inst_pe_1_5_5_int_q_weight_0_), .A2(
        npu_inst_pe_1_5_5_n1), .ZN(npu_inst_pe_1_5_5_n76) );
  NOR2_X1 npu_inst_pe_1_5_5_U3 ( .A1(npu_inst_pe_1_5_5_n27), .A2(
        npu_inst_pe_1_5_5_n1), .ZN(npu_inst_pe_1_5_5_n77) );
  FA_X1 npu_inst_pe_1_5_5_sub_77_U2_1 ( .A(npu_inst_pe_1_5_5_int_q_acc_1_), 
        .B(npu_inst_pe_1_5_5_n14), .CI(npu_inst_pe_1_5_5_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_5_5_sub_77_carry_2_), .S(npu_inst_pe_1_5_5_N66) );
  FA_X1 npu_inst_pe_1_5_5_add_79_U1_1 ( .A(npu_inst_pe_1_5_5_int_q_acc_1_), 
        .B(npu_inst_pe_1_5_5_int_data_1_), .CI(
        npu_inst_pe_1_5_5_add_79_carry_1_), .CO(
        npu_inst_pe_1_5_5_add_79_carry_2_), .S(npu_inst_pe_1_5_5_N74) );
  NAND3_X1 npu_inst_pe_1_5_5_U109 ( .A1(npu_inst_pe_1_5_5_n5), .A2(
        npu_inst_pe_1_5_5_n7), .A3(npu_inst_pe_1_5_5_n8), .ZN(
        npu_inst_pe_1_5_5_n44) );
  NAND3_X1 npu_inst_pe_1_5_5_U108 ( .A1(npu_inst_pe_1_5_5_n4), .A2(
        npu_inst_pe_1_5_5_n7), .A3(npu_inst_pe_1_5_5_n8), .ZN(
        npu_inst_pe_1_5_5_n40) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_5_5_n34), .CK(
        npu_inst_pe_1_5_5_net3258), .RN(npu_inst_pe_1_5_5_n9), .Q(
        npu_inst_pe_1_5_5_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_5_5_n35), .CK(
        npu_inst_pe_1_5_5_net3258), .RN(npu_inst_pe_1_5_5_n9), .Q(
        npu_inst_pe_1_5_5_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_5_5_n36), .CK(
        npu_inst_pe_1_5_5_net3258), .RN(npu_inst_pe_1_5_5_n9), .Q(
        npu_inst_pe_1_5_5_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_5_5_n98), .CK(
        npu_inst_pe_1_5_5_net3258), .RN(npu_inst_pe_1_5_5_n9), .Q(
        npu_inst_pe_1_5_5_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_5_5_n99), .CK(
        npu_inst_pe_1_5_5_net3258), .RN(npu_inst_pe_1_5_5_n9), .Q(
        npu_inst_pe_1_5_5_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_5_5_n100), 
        .CK(npu_inst_pe_1_5_5_net3258), .RN(npu_inst_pe_1_5_5_n9), .Q(
        npu_inst_pe_1_5_5_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_5_5_n33), .CK(
        npu_inst_pe_1_5_5_net3258), .RN(npu_inst_pe_1_5_5_n9), .Q(
        npu_inst_pe_1_5_5_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_5_5_n101), 
        .CK(npu_inst_pe_1_5_5_net3258), .RN(npu_inst_pe_1_5_5_n9), .Q(
        npu_inst_pe_1_5_5_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_weight_reg_0_ ( .D(npu_inst_n109), .CK(
        npu_inst_pe_1_5_5_net3264), .RN(npu_inst_pe_1_5_5_n9), .Q(
        npu_inst_pe_1_5_5_int_q_weight_0_), .QN(npu_inst_pe_1_5_5_n27) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_weight_reg_1_ ( .D(npu_inst_n115), .CK(
        npu_inst_pe_1_5_5_net3264), .RN(npu_inst_pe_1_5_5_n9), .Q(
        npu_inst_pe_1_5_5_int_q_weight_1_), .QN(npu_inst_pe_1_5_5_n26) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_5_5_n113), 
        .CK(npu_inst_pe_1_5_5_net3264), .RN(npu_inst_pe_1_5_5_n9), .Q(
        npu_inst_pe_1_5_5_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_5_5_n107), 
        .CK(npu_inst_pe_1_5_5_net3264), .RN(npu_inst_pe_1_5_5_n9), .Q(
        npu_inst_pe_1_5_5_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_5_5_n112), 
        .CK(npu_inst_pe_1_5_5_net3264), .RN(npu_inst_pe_1_5_5_n10), .Q(
        npu_inst_pe_1_5_5_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_5_5_n106), 
        .CK(npu_inst_pe_1_5_5_net3264), .RN(npu_inst_pe_1_5_5_n10), .Q(
        npu_inst_pe_1_5_5_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_5_5_n111), 
        .CK(npu_inst_pe_1_5_5_net3264), .RN(npu_inst_pe_1_5_5_n10), .Q(
        npu_inst_pe_1_5_5_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_5_5_n105), 
        .CK(npu_inst_pe_1_5_5_net3264), .RN(npu_inst_pe_1_5_5_n10), .Q(
        npu_inst_pe_1_5_5_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_5_5_n110), 
        .CK(npu_inst_pe_1_5_5_net3264), .RN(npu_inst_pe_1_5_5_n10), .Q(
        npu_inst_pe_1_5_5_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_5_5_n104), 
        .CK(npu_inst_pe_1_5_5_net3264), .RN(npu_inst_pe_1_5_5_n10), .Q(
        npu_inst_pe_1_5_5_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_5_5_n109), 
        .CK(npu_inst_pe_1_5_5_net3264), .RN(npu_inst_pe_1_5_5_n10), .Q(
        npu_inst_pe_1_5_5_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_5_5_n103), 
        .CK(npu_inst_pe_1_5_5_net3264), .RN(npu_inst_pe_1_5_5_n10), .Q(
        npu_inst_pe_1_5_5_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_5_5_n108), 
        .CK(npu_inst_pe_1_5_5_net3264), .RN(npu_inst_pe_1_5_5_n10), .Q(
        npu_inst_pe_1_5_5_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_5_5_n102), 
        .CK(npu_inst_pe_1_5_5_net3264), .RN(npu_inst_pe_1_5_5_n10), .Q(
        npu_inst_pe_1_5_5_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_5_5_n86), 
        .CK(npu_inst_pe_1_5_5_net3264), .RN(npu_inst_pe_1_5_5_n10), .Q(
        npu_inst_pe_1_5_5_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_5_5_n87), 
        .CK(npu_inst_pe_1_5_5_net3264), .RN(npu_inst_pe_1_5_5_n10), .Q(
        npu_inst_pe_1_5_5_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_5_5_n88), 
        .CK(npu_inst_pe_1_5_5_net3264), .RN(npu_inst_pe_1_5_5_n11), .Q(
        npu_inst_pe_1_5_5_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_5_5_n89), 
        .CK(npu_inst_pe_1_5_5_net3264), .RN(npu_inst_pe_1_5_5_n11), .Q(
        npu_inst_pe_1_5_5_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_5_5_n90), 
        .CK(npu_inst_pe_1_5_5_net3264), .RN(npu_inst_pe_1_5_5_n11), .Q(
        npu_inst_pe_1_5_5_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_5_5_n91), 
        .CK(npu_inst_pe_1_5_5_net3264), .RN(npu_inst_pe_1_5_5_n11), .Q(
        npu_inst_pe_1_5_5_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_5_5_n92), 
        .CK(npu_inst_pe_1_5_5_net3264), .RN(npu_inst_pe_1_5_5_n11), .Q(
        npu_inst_pe_1_5_5_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_5_5_n93), 
        .CK(npu_inst_pe_1_5_5_net3264), .RN(npu_inst_pe_1_5_5_n11), .Q(
        npu_inst_pe_1_5_5_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_5_5_n94), 
        .CK(npu_inst_pe_1_5_5_net3264), .RN(npu_inst_pe_1_5_5_n11), .Q(
        npu_inst_pe_1_5_5_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_5_5_n95), 
        .CK(npu_inst_pe_1_5_5_net3264), .RN(npu_inst_pe_1_5_5_n11), .Q(
        npu_inst_pe_1_5_5_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_5_5_n96), 
        .CK(npu_inst_pe_1_5_5_net3264), .RN(npu_inst_pe_1_5_5_n11), .Q(
        npu_inst_pe_1_5_5_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_5_5_n97), 
        .CK(npu_inst_pe_1_5_5_net3264), .RN(npu_inst_pe_1_5_5_n11), .Q(
        npu_inst_pe_1_5_5_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_5_5_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_5_5_N84), .SE(1'b0), .GCK(npu_inst_pe_1_5_5_net3258) );
  CLKGATETST_X1 npu_inst_pe_1_5_5_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n62), .SE(1'b0), .GCK(npu_inst_pe_1_5_5_net3264) );
  MUX2_X1 npu_inst_pe_1_5_6_U162 ( .A(npu_inst_pe_1_5_6_n32), .B(
        npu_inst_pe_1_5_6_n29), .S(npu_inst_pe_1_5_6_n8), .Z(
        npu_inst_pe_1_5_6_N93) );
  MUX2_X1 npu_inst_pe_1_5_6_U161 ( .A(npu_inst_pe_1_5_6_n31), .B(
        npu_inst_pe_1_5_6_n30), .S(npu_inst_pe_1_5_6_n6), .Z(
        npu_inst_pe_1_5_6_n32) );
  MUX2_X1 npu_inst_pe_1_5_6_U160 ( .A(npu_inst_pe_1_5_6_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_5_6_int_q_reg_v_1__0_), .S(npu_inst_pe_1_5_6_n4), .Z(
        npu_inst_pe_1_5_6_n31) );
  MUX2_X1 npu_inst_pe_1_5_6_U159 ( .A(npu_inst_pe_1_5_6_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_5_6_int_q_reg_v_3__0_), .S(npu_inst_pe_1_5_6_n4), .Z(
        npu_inst_pe_1_5_6_n30) );
  MUX2_X1 npu_inst_pe_1_5_6_U158 ( .A(npu_inst_pe_1_5_6_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_5_6_int_q_reg_v_5__0_), .S(npu_inst_pe_1_5_6_n4), .Z(
        npu_inst_pe_1_5_6_n29) );
  MUX2_X1 npu_inst_pe_1_5_6_U157 ( .A(npu_inst_pe_1_5_6_n28), .B(
        npu_inst_pe_1_5_6_n23), .S(npu_inst_pe_1_5_6_n8), .Z(
        npu_inst_pe_1_5_6_N94) );
  MUX2_X1 npu_inst_pe_1_5_6_U156 ( .A(npu_inst_pe_1_5_6_n25), .B(
        npu_inst_pe_1_5_6_n24), .S(npu_inst_pe_1_5_6_n6), .Z(
        npu_inst_pe_1_5_6_n28) );
  MUX2_X1 npu_inst_pe_1_5_6_U155 ( .A(npu_inst_pe_1_5_6_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_5_6_int_q_reg_v_1__1_), .S(npu_inst_pe_1_5_6_n4), .Z(
        npu_inst_pe_1_5_6_n25) );
  MUX2_X1 npu_inst_pe_1_5_6_U154 ( .A(npu_inst_pe_1_5_6_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_5_6_int_q_reg_v_3__1_), .S(npu_inst_pe_1_5_6_n4), .Z(
        npu_inst_pe_1_5_6_n24) );
  MUX2_X1 npu_inst_pe_1_5_6_U153 ( .A(npu_inst_pe_1_5_6_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_5_6_int_q_reg_v_5__1_), .S(npu_inst_pe_1_5_6_n4), .Z(
        npu_inst_pe_1_5_6_n23) );
  MUX2_X1 npu_inst_pe_1_5_6_U152 ( .A(npu_inst_pe_1_5_6_n22), .B(
        npu_inst_pe_1_5_6_n19), .S(npu_inst_pe_1_5_6_n8), .Z(
        npu_inst_int_data_x_5__6__1_) );
  MUX2_X1 npu_inst_pe_1_5_6_U151 ( .A(npu_inst_pe_1_5_6_n21), .B(
        npu_inst_pe_1_5_6_n20), .S(npu_inst_pe_1_5_6_n6), .Z(
        npu_inst_pe_1_5_6_n22) );
  MUX2_X1 npu_inst_pe_1_5_6_U150 ( .A(npu_inst_pe_1_5_6_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_5_6_int_q_reg_h_1__1_), .S(npu_inst_pe_1_5_6_n4), .Z(
        npu_inst_pe_1_5_6_n21) );
  MUX2_X1 npu_inst_pe_1_5_6_U149 ( .A(npu_inst_pe_1_5_6_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_5_6_int_q_reg_h_3__1_), .S(npu_inst_pe_1_5_6_n4), .Z(
        npu_inst_pe_1_5_6_n20) );
  MUX2_X1 npu_inst_pe_1_5_6_U148 ( .A(npu_inst_pe_1_5_6_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_5_6_int_q_reg_h_5__1_), .S(npu_inst_pe_1_5_6_n4), .Z(
        npu_inst_pe_1_5_6_n19) );
  MUX2_X1 npu_inst_pe_1_5_6_U147 ( .A(npu_inst_pe_1_5_6_n18), .B(
        npu_inst_pe_1_5_6_n15), .S(npu_inst_pe_1_5_6_n8), .Z(
        npu_inst_int_data_x_5__6__0_) );
  MUX2_X1 npu_inst_pe_1_5_6_U146 ( .A(npu_inst_pe_1_5_6_n17), .B(
        npu_inst_pe_1_5_6_n16), .S(npu_inst_pe_1_5_6_n6), .Z(
        npu_inst_pe_1_5_6_n18) );
  MUX2_X1 npu_inst_pe_1_5_6_U145 ( .A(npu_inst_pe_1_5_6_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_5_6_int_q_reg_h_1__0_), .S(npu_inst_pe_1_5_6_n4), .Z(
        npu_inst_pe_1_5_6_n17) );
  MUX2_X1 npu_inst_pe_1_5_6_U144 ( .A(npu_inst_pe_1_5_6_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_5_6_int_q_reg_h_3__0_), .S(npu_inst_pe_1_5_6_n4), .Z(
        npu_inst_pe_1_5_6_n16) );
  MUX2_X1 npu_inst_pe_1_5_6_U143 ( .A(npu_inst_pe_1_5_6_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_5_6_int_q_reg_h_5__0_), .S(npu_inst_pe_1_5_6_n4), .Z(
        npu_inst_pe_1_5_6_n15) );
  XOR2_X1 npu_inst_pe_1_5_6_U142 ( .A(npu_inst_pe_1_5_6_int_data_0_), .B(
        npu_inst_pe_1_5_6_int_q_acc_0_), .Z(npu_inst_pe_1_5_6_N73) );
  AND2_X1 npu_inst_pe_1_5_6_U141 ( .A1(npu_inst_pe_1_5_6_int_q_acc_0_), .A2(
        npu_inst_pe_1_5_6_int_data_0_), .ZN(npu_inst_pe_1_5_6_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_5_6_U140 ( .A(npu_inst_pe_1_5_6_int_q_acc_0_), .B(
        npu_inst_pe_1_5_6_n13), .ZN(npu_inst_pe_1_5_6_N65) );
  OR2_X1 npu_inst_pe_1_5_6_U139 ( .A1(npu_inst_pe_1_5_6_n13), .A2(
        npu_inst_pe_1_5_6_int_q_acc_0_), .ZN(npu_inst_pe_1_5_6_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_5_6_U138 ( .A(npu_inst_pe_1_5_6_int_q_acc_2_), .B(
        npu_inst_pe_1_5_6_add_79_carry_2_), .Z(npu_inst_pe_1_5_6_N75) );
  AND2_X1 npu_inst_pe_1_5_6_U137 ( .A1(npu_inst_pe_1_5_6_add_79_carry_2_), 
        .A2(npu_inst_pe_1_5_6_int_q_acc_2_), .ZN(
        npu_inst_pe_1_5_6_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_5_6_U136 ( .A(npu_inst_pe_1_5_6_int_q_acc_3_), .B(
        npu_inst_pe_1_5_6_add_79_carry_3_), .Z(npu_inst_pe_1_5_6_N76) );
  AND2_X1 npu_inst_pe_1_5_6_U135 ( .A1(npu_inst_pe_1_5_6_add_79_carry_3_), 
        .A2(npu_inst_pe_1_5_6_int_q_acc_3_), .ZN(
        npu_inst_pe_1_5_6_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_5_6_U134 ( .A(npu_inst_pe_1_5_6_int_q_acc_4_), .B(
        npu_inst_pe_1_5_6_add_79_carry_4_), .Z(npu_inst_pe_1_5_6_N77) );
  AND2_X1 npu_inst_pe_1_5_6_U133 ( .A1(npu_inst_pe_1_5_6_add_79_carry_4_), 
        .A2(npu_inst_pe_1_5_6_int_q_acc_4_), .ZN(
        npu_inst_pe_1_5_6_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_5_6_U132 ( .A(npu_inst_pe_1_5_6_int_q_acc_5_), .B(
        npu_inst_pe_1_5_6_add_79_carry_5_), .Z(npu_inst_pe_1_5_6_N78) );
  AND2_X1 npu_inst_pe_1_5_6_U131 ( .A1(npu_inst_pe_1_5_6_add_79_carry_5_), 
        .A2(npu_inst_pe_1_5_6_int_q_acc_5_), .ZN(
        npu_inst_pe_1_5_6_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_5_6_U130 ( .A(npu_inst_pe_1_5_6_int_q_acc_6_), .B(
        npu_inst_pe_1_5_6_add_79_carry_6_), .Z(npu_inst_pe_1_5_6_N79) );
  AND2_X1 npu_inst_pe_1_5_6_U129 ( .A1(npu_inst_pe_1_5_6_add_79_carry_6_), 
        .A2(npu_inst_pe_1_5_6_int_q_acc_6_), .ZN(
        npu_inst_pe_1_5_6_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_5_6_U128 ( .A(npu_inst_pe_1_5_6_int_q_acc_7_), .B(
        npu_inst_pe_1_5_6_add_79_carry_7_), .Z(npu_inst_pe_1_5_6_N80) );
  XNOR2_X1 npu_inst_pe_1_5_6_U127 ( .A(npu_inst_pe_1_5_6_sub_77_carry_2_), .B(
        npu_inst_pe_1_5_6_int_q_acc_2_), .ZN(npu_inst_pe_1_5_6_N67) );
  OR2_X1 npu_inst_pe_1_5_6_U126 ( .A1(npu_inst_pe_1_5_6_int_q_acc_2_), .A2(
        npu_inst_pe_1_5_6_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_5_6_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_5_6_U125 ( .A(npu_inst_pe_1_5_6_sub_77_carry_3_), .B(
        npu_inst_pe_1_5_6_int_q_acc_3_), .ZN(npu_inst_pe_1_5_6_N68) );
  OR2_X1 npu_inst_pe_1_5_6_U124 ( .A1(npu_inst_pe_1_5_6_int_q_acc_3_), .A2(
        npu_inst_pe_1_5_6_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_5_6_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_5_6_U123 ( .A(npu_inst_pe_1_5_6_sub_77_carry_4_), .B(
        npu_inst_pe_1_5_6_int_q_acc_4_), .ZN(npu_inst_pe_1_5_6_N69) );
  OR2_X1 npu_inst_pe_1_5_6_U122 ( .A1(npu_inst_pe_1_5_6_int_q_acc_4_), .A2(
        npu_inst_pe_1_5_6_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_5_6_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_5_6_U121 ( .A(npu_inst_pe_1_5_6_sub_77_carry_5_), .B(
        npu_inst_pe_1_5_6_int_q_acc_5_), .ZN(npu_inst_pe_1_5_6_N70) );
  OR2_X1 npu_inst_pe_1_5_6_U120 ( .A1(npu_inst_pe_1_5_6_int_q_acc_5_), .A2(
        npu_inst_pe_1_5_6_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_5_6_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_5_6_U119 ( .A(npu_inst_pe_1_5_6_sub_77_carry_6_), .B(
        npu_inst_pe_1_5_6_int_q_acc_6_), .ZN(npu_inst_pe_1_5_6_N71) );
  OR2_X1 npu_inst_pe_1_5_6_U118 ( .A1(npu_inst_pe_1_5_6_int_q_acc_6_), .A2(
        npu_inst_pe_1_5_6_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_5_6_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_5_6_U117 ( .A(npu_inst_pe_1_5_6_int_q_acc_7_), .B(
        npu_inst_pe_1_5_6_sub_77_carry_7_), .ZN(npu_inst_pe_1_5_6_N72) );
  INV_X1 npu_inst_pe_1_5_6_U116 ( .A(npu_inst_n76), .ZN(npu_inst_pe_1_5_6_n7)
         );
  INV_X1 npu_inst_pe_1_5_6_U115 ( .A(npu_inst_pe_1_5_6_n7), .ZN(
        npu_inst_pe_1_5_6_n6) );
  INV_X1 npu_inst_pe_1_5_6_U114 ( .A(npu_inst_n54), .ZN(npu_inst_pe_1_5_6_n3)
         );
  AOI22_X1 npu_inst_pe_1_5_6_U113 ( .A1(npu_inst_int_data_y_6__6__0_), .A2(
        npu_inst_pe_1_5_6_n58), .B1(npu_inst_pe_1_5_6_n114), .B2(
        npu_inst_pe_1_5_6_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_5_6_n57) );
  INV_X1 npu_inst_pe_1_5_6_U112 ( .A(npu_inst_pe_1_5_6_n57), .ZN(
        npu_inst_pe_1_5_6_n108) );
  AOI22_X1 npu_inst_pe_1_5_6_U111 ( .A1(npu_inst_int_data_y_6__6__0_), .A2(
        npu_inst_pe_1_5_6_n54), .B1(npu_inst_pe_1_5_6_n115), .B2(
        npu_inst_pe_1_5_6_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_5_6_n53) );
  INV_X1 npu_inst_pe_1_5_6_U110 ( .A(npu_inst_pe_1_5_6_n53), .ZN(
        npu_inst_pe_1_5_6_n109) );
  AOI22_X1 npu_inst_pe_1_5_6_U107 ( .A1(npu_inst_int_data_y_6__6__0_), .A2(
        npu_inst_pe_1_5_6_n50), .B1(npu_inst_pe_1_5_6_n116), .B2(
        npu_inst_pe_1_5_6_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_5_6_n49) );
  INV_X1 npu_inst_pe_1_5_6_U106 ( .A(npu_inst_pe_1_5_6_n49), .ZN(
        npu_inst_pe_1_5_6_n110) );
  AOI22_X1 npu_inst_pe_1_5_6_U105 ( .A1(npu_inst_int_data_y_6__6__0_), .A2(
        npu_inst_pe_1_5_6_n46), .B1(npu_inst_pe_1_5_6_n117), .B2(
        npu_inst_pe_1_5_6_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_5_6_n45) );
  INV_X1 npu_inst_pe_1_5_6_U104 ( .A(npu_inst_pe_1_5_6_n45), .ZN(
        npu_inst_pe_1_5_6_n111) );
  AOI22_X1 npu_inst_pe_1_5_6_U103 ( .A1(npu_inst_int_data_y_6__6__0_), .A2(
        npu_inst_pe_1_5_6_n42), .B1(npu_inst_pe_1_5_6_n119), .B2(
        npu_inst_pe_1_5_6_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_5_6_n41) );
  INV_X1 npu_inst_pe_1_5_6_U102 ( .A(npu_inst_pe_1_5_6_n41), .ZN(
        npu_inst_pe_1_5_6_n112) );
  AOI22_X1 npu_inst_pe_1_5_6_U101 ( .A1(npu_inst_int_data_y_6__6__1_), .A2(
        npu_inst_pe_1_5_6_n58), .B1(npu_inst_pe_1_5_6_n114), .B2(
        npu_inst_pe_1_5_6_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_5_6_n59) );
  INV_X1 npu_inst_pe_1_5_6_U100 ( .A(npu_inst_pe_1_5_6_n59), .ZN(
        npu_inst_pe_1_5_6_n102) );
  AOI22_X1 npu_inst_pe_1_5_6_U99 ( .A1(npu_inst_int_data_y_6__6__1_), .A2(
        npu_inst_pe_1_5_6_n54), .B1(npu_inst_pe_1_5_6_n115), .B2(
        npu_inst_pe_1_5_6_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_5_6_n55) );
  INV_X1 npu_inst_pe_1_5_6_U98 ( .A(npu_inst_pe_1_5_6_n55), .ZN(
        npu_inst_pe_1_5_6_n103) );
  AOI22_X1 npu_inst_pe_1_5_6_U97 ( .A1(npu_inst_int_data_y_6__6__1_), .A2(
        npu_inst_pe_1_5_6_n50), .B1(npu_inst_pe_1_5_6_n116), .B2(
        npu_inst_pe_1_5_6_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_5_6_n51) );
  INV_X1 npu_inst_pe_1_5_6_U96 ( .A(npu_inst_pe_1_5_6_n51), .ZN(
        npu_inst_pe_1_5_6_n104) );
  AOI22_X1 npu_inst_pe_1_5_6_U95 ( .A1(npu_inst_int_data_y_6__6__1_), .A2(
        npu_inst_pe_1_5_6_n46), .B1(npu_inst_pe_1_5_6_n117), .B2(
        npu_inst_pe_1_5_6_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_5_6_n47) );
  INV_X1 npu_inst_pe_1_5_6_U94 ( .A(npu_inst_pe_1_5_6_n47), .ZN(
        npu_inst_pe_1_5_6_n105) );
  AOI22_X1 npu_inst_pe_1_5_6_U93 ( .A1(npu_inst_int_data_y_6__6__1_), .A2(
        npu_inst_pe_1_5_6_n42), .B1(npu_inst_pe_1_5_6_n119), .B2(
        npu_inst_pe_1_5_6_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_5_6_n43) );
  INV_X1 npu_inst_pe_1_5_6_U92 ( .A(npu_inst_pe_1_5_6_n43), .ZN(
        npu_inst_pe_1_5_6_n106) );
  AOI22_X1 npu_inst_pe_1_5_6_U91 ( .A1(npu_inst_pe_1_5_6_n38), .A2(
        npu_inst_int_data_y_6__6__1_), .B1(npu_inst_pe_1_5_6_n118), .B2(
        npu_inst_pe_1_5_6_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_5_6_n39) );
  INV_X1 npu_inst_pe_1_5_6_U90 ( .A(npu_inst_pe_1_5_6_n39), .ZN(
        npu_inst_pe_1_5_6_n107) );
  AOI22_X1 npu_inst_pe_1_5_6_U89 ( .A1(npu_inst_pe_1_5_6_n38), .A2(
        npu_inst_int_data_y_6__6__0_), .B1(npu_inst_pe_1_5_6_n118), .B2(
        npu_inst_pe_1_5_6_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_5_6_n37) );
  INV_X1 npu_inst_pe_1_5_6_U88 ( .A(npu_inst_pe_1_5_6_n37), .ZN(
        npu_inst_pe_1_5_6_n113) );
  NAND2_X1 npu_inst_pe_1_5_6_U87 ( .A1(npu_inst_pe_1_5_6_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_5_6_n60), .ZN(npu_inst_pe_1_5_6_n74) );
  OAI21_X1 npu_inst_pe_1_5_6_U86 ( .B1(npu_inst_pe_1_5_6_n63), .B2(
        npu_inst_pe_1_5_6_n60), .A(npu_inst_pe_1_5_6_n74), .ZN(
        npu_inst_pe_1_5_6_n97) );
  NAND2_X1 npu_inst_pe_1_5_6_U85 ( .A1(npu_inst_pe_1_5_6_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_5_6_n60), .ZN(npu_inst_pe_1_5_6_n73) );
  OAI21_X1 npu_inst_pe_1_5_6_U84 ( .B1(npu_inst_pe_1_5_6_n61), .B2(
        npu_inst_pe_1_5_6_n60), .A(npu_inst_pe_1_5_6_n73), .ZN(
        npu_inst_pe_1_5_6_n96) );
  NAND2_X1 npu_inst_pe_1_5_6_U83 ( .A1(npu_inst_pe_1_5_6_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_5_6_n56), .ZN(npu_inst_pe_1_5_6_n72) );
  OAI21_X1 npu_inst_pe_1_5_6_U82 ( .B1(npu_inst_pe_1_5_6_n63), .B2(
        npu_inst_pe_1_5_6_n56), .A(npu_inst_pe_1_5_6_n72), .ZN(
        npu_inst_pe_1_5_6_n95) );
  NAND2_X1 npu_inst_pe_1_5_6_U81 ( .A1(npu_inst_pe_1_5_6_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_5_6_n56), .ZN(npu_inst_pe_1_5_6_n71) );
  OAI21_X1 npu_inst_pe_1_5_6_U80 ( .B1(npu_inst_pe_1_5_6_n61), .B2(
        npu_inst_pe_1_5_6_n56), .A(npu_inst_pe_1_5_6_n71), .ZN(
        npu_inst_pe_1_5_6_n94) );
  NAND2_X1 npu_inst_pe_1_5_6_U79 ( .A1(npu_inst_pe_1_5_6_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_5_6_n52), .ZN(npu_inst_pe_1_5_6_n70) );
  OAI21_X1 npu_inst_pe_1_5_6_U78 ( .B1(npu_inst_pe_1_5_6_n63), .B2(
        npu_inst_pe_1_5_6_n52), .A(npu_inst_pe_1_5_6_n70), .ZN(
        npu_inst_pe_1_5_6_n93) );
  NAND2_X1 npu_inst_pe_1_5_6_U77 ( .A1(npu_inst_pe_1_5_6_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_5_6_n52), .ZN(npu_inst_pe_1_5_6_n69) );
  OAI21_X1 npu_inst_pe_1_5_6_U76 ( .B1(npu_inst_pe_1_5_6_n61), .B2(
        npu_inst_pe_1_5_6_n52), .A(npu_inst_pe_1_5_6_n69), .ZN(
        npu_inst_pe_1_5_6_n92) );
  NAND2_X1 npu_inst_pe_1_5_6_U75 ( .A1(npu_inst_pe_1_5_6_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_5_6_n48), .ZN(npu_inst_pe_1_5_6_n68) );
  OAI21_X1 npu_inst_pe_1_5_6_U74 ( .B1(npu_inst_pe_1_5_6_n63), .B2(
        npu_inst_pe_1_5_6_n48), .A(npu_inst_pe_1_5_6_n68), .ZN(
        npu_inst_pe_1_5_6_n91) );
  NAND2_X1 npu_inst_pe_1_5_6_U73 ( .A1(npu_inst_pe_1_5_6_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_5_6_n48), .ZN(npu_inst_pe_1_5_6_n67) );
  OAI21_X1 npu_inst_pe_1_5_6_U72 ( .B1(npu_inst_pe_1_5_6_n61), .B2(
        npu_inst_pe_1_5_6_n48), .A(npu_inst_pe_1_5_6_n67), .ZN(
        npu_inst_pe_1_5_6_n90) );
  NAND2_X1 npu_inst_pe_1_5_6_U71 ( .A1(npu_inst_pe_1_5_6_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_5_6_n44), .ZN(npu_inst_pe_1_5_6_n66) );
  OAI21_X1 npu_inst_pe_1_5_6_U70 ( .B1(npu_inst_pe_1_5_6_n63), .B2(
        npu_inst_pe_1_5_6_n44), .A(npu_inst_pe_1_5_6_n66), .ZN(
        npu_inst_pe_1_5_6_n89) );
  NAND2_X1 npu_inst_pe_1_5_6_U69 ( .A1(npu_inst_pe_1_5_6_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_5_6_n44), .ZN(npu_inst_pe_1_5_6_n65) );
  OAI21_X1 npu_inst_pe_1_5_6_U68 ( .B1(npu_inst_pe_1_5_6_n61), .B2(
        npu_inst_pe_1_5_6_n44), .A(npu_inst_pe_1_5_6_n65), .ZN(
        npu_inst_pe_1_5_6_n88) );
  NAND2_X1 npu_inst_pe_1_5_6_U67 ( .A1(npu_inst_pe_1_5_6_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_5_6_n40), .ZN(npu_inst_pe_1_5_6_n64) );
  OAI21_X1 npu_inst_pe_1_5_6_U66 ( .B1(npu_inst_pe_1_5_6_n63), .B2(
        npu_inst_pe_1_5_6_n40), .A(npu_inst_pe_1_5_6_n64), .ZN(
        npu_inst_pe_1_5_6_n87) );
  NAND2_X1 npu_inst_pe_1_5_6_U65 ( .A1(npu_inst_pe_1_5_6_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_5_6_n40), .ZN(npu_inst_pe_1_5_6_n62) );
  OAI21_X1 npu_inst_pe_1_5_6_U64 ( .B1(npu_inst_pe_1_5_6_n61), .B2(
        npu_inst_pe_1_5_6_n40), .A(npu_inst_pe_1_5_6_n62), .ZN(
        npu_inst_pe_1_5_6_n86) );
  AND2_X1 npu_inst_pe_1_5_6_U63 ( .A1(npu_inst_pe_1_5_6_N93), .A2(npu_inst_n54), .ZN(npu_inst_int_data_y_5__6__0_) );
  AND2_X1 npu_inst_pe_1_5_6_U62 ( .A1(npu_inst_n54), .A2(npu_inst_pe_1_5_6_N94), .ZN(npu_inst_int_data_y_5__6__1_) );
  NOR3_X1 npu_inst_pe_1_5_6_U61 ( .A1(npu_inst_pe_1_5_6_n26), .A2(npu_inst_n54), .A3(npu_inst_int_ckg[17]), .ZN(npu_inst_pe_1_5_6_n85) );
  OR2_X1 npu_inst_pe_1_5_6_U60 ( .A1(npu_inst_pe_1_5_6_n85), .A2(
        npu_inst_pe_1_5_6_n2), .ZN(npu_inst_pe_1_5_6_N84) );
  AND2_X1 npu_inst_pe_1_5_6_U59 ( .A1(npu_inst_pe_1_5_6_int_q_acc_0_), .A2(
        npu_inst_pe_1_5_6_n1), .ZN(npu_inst_int_data_res_5__6__0_) );
  AND2_X1 npu_inst_pe_1_5_6_U58 ( .A1(npu_inst_pe_1_5_6_n2), .A2(
        npu_inst_pe_1_5_6_int_q_acc_7_), .ZN(npu_inst_int_data_res_5__6__7_)
         );
  AND2_X1 npu_inst_pe_1_5_6_U57 ( .A1(npu_inst_pe_1_5_6_int_q_acc_1_), .A2(
        npu_inst_pe_1_5_6_n1), .ZN(npu_inst_int_data_res_5__6__1_) );
  AND2_X1 npu_inst_pe_1_5_6_U56 ( .A1(npu_inst_pe_1_5_6_int_q_acc_2_), .A2(
        npu_inst_pe_1_5_6_n1), .ZN(npu_inst_int_data_res_5__6__2_) );
  AND2_X1 npu_inst_pe_1_5_6_U55 ( .A1(npu_inst_pe_1_5_6_int_q_acc_3_), .A2(
        npu_inst_pe_1_5_6_n2), .ZN(npu_inst_int_data_res_5__6__3_) );
  AND2_X1 npu_inst_pe_1_5_6_U54 ( .A1(npu_inst_pe_1_5_6_int_q_acc_4_), .A2(
        npu_inst_pe_1_5_6_n2), .ZN(npu_inst_int_data_res_5__6__4_) );
  AND2_X1 npu_inst_pe_1_5_6_U53 ( .A1(npu_inst_pe_1_5_6_int_q_acc_5_), .A2(
        npu_inst_pe_1_5_6_n2), .ZN(npu_inst_int_data_res_5__6__5_) );
  AND2_X1 npu_inst_pe_1_5_6_U52 ( .A1(npu_inst_pe_1_5_6_int_q_acc_6_), .A2(
        npu_inst_pe_1_5_6_n2), .ZN(npu_inst_int_data_res_5__6__6_) );
  AOI222_X1 npu_inst_pe_1_5_6_U51 ( .A1(npu_inst_int_data_res_6__6__0_), .A2(
        npu_inst_pe_1_5_6_n1), .B1(npu_inst_pe_1_5_6_N73), .B2(
        npu_inst_pe_1_5_6_n76), .C1(npu_inst_pe_1_5_6_N65), .C2(
        npu_inst_pe_1_5_6_n77), .ZN(npu_inst_pe_1_5_6_n84) );
  INV_X1 npu_inst_pe_1_5_6_U50 ( .A(npu_inst_pe_1_5_6_n84), .ZN(
        npu_inst_pe_1_5_6_n101) );
  AOI222_X1 npu_inst_pe_1_5_6_U49 ( .A1(npu_inst_int_data_res_6__6__7_), .A2(
        npu_inst_pe_1_5_6_n1), .B1(npu_inst_pe_1_5_6_N80), .B2(
        npu_inst_pe_1_5_6_n76), .C1(npu_inst_pe_1_5_6_N72), .C2(
        npu_inst_pe_1_5_6_n77), .ZN(npu_inst_pe_1_5_6_n75) );
  INV_X1 npu_inst_pe_1_5_6_U48 ( .A(npu_inst_pe_1_5_6_n75), .ZN(
        npu_inst_pe_1_5_6_n33) );
  AOI222_X1 npu_inst_pe_1_5_6_U47 ( .A1(npu_inst_int_data_res_6__6__1_), .A2(
        npu_inst_pe_1_5_6_n1), .B1(npu_inst_pe_1_5_6_N74), .B2(
        npu_inst_pe_1_5_6_n76), .C1(npu_inst_pe_1_5_6_N66), .C2(
        npu_inst_pe_1_5_6_n77), .ZN(npu_inst_pe_1_5_6_n83) );
  INV_X1 npu_inst_pe_1_5_6_U46 ( .A(npu_inst_pe_1_5_6_n83), .ZN(
        npu_inst_pe_1_5_6_n100) );
  AOI222_X1 npu_inst_pe_1_5_6_U45 ( .A1(npu_inst_int_data_res_6__6__2_), .A2(
        npu_inst_pe_1_5_6_n1), .B1(npu_inst_pe_1_5_6_N75), .B2(
        npu_inst_pe_1_5_6_n76), .C1(npu_inst_pe_1_5_6_N67), .C2(
        npu_inst_pe_1_5_6_n77), .ZN(npu_inst_pe_1_5_6_n82) );
  INV_X1 npu_inst_pe_1_5_6_U44 ( .A(npu_inst_pe_1_5_6_n82), .ZN(
        npu_inst_pe_1_5_6_n99) );
  AOI222_X1 npu_inst_pe_1_5_6_U43 ( .A1(npu_inst_int_data_res_6__6__3_), .A2(
        npu_inst_pe_1_5_6_n1), .B1(npu_inst_pe_1_5_6_N76), .B2(
        npu_inst_pe_1_5_6_n76), .C1(npu_inst_pe_1_5_6_N68), .C2(
        npu_inst_pe_1_5_6_n77), .ZN(npu_inst_pe_1_5_6_n81) );
  INV_X1 npu_inst_pe_1_5_6_U42 ( .A(npu_inst_pe_1_5_6_n81), .ZN(
        npu_inst_pe_1_5_6_n98) );
  AOI222_X1 npu_inst_pe_1_5_6_U41 ( .A1(npu_inst_int_data_res_6__6__4_), .A2(
        npu_inst_pe_1_5_6_n1), .B1(npu_inst_pe_1_5_6_N77), .B2(
        npu_inst_pe_1_5_6_n76), .C1(npu_inst_pe_1_5_6_N69), .C2(
        npu_inst_pe_1_5_6_n77), .ZN(npu_inst_pe_1_5_6_n80) );
  INV_X1 npu_inst_pe_1_5_6_U40 ( .A(npu_inst_pe_1_5_6_n80), .ZN(
        npu_inst_pe_1_5_6_n36) );
  AOI222_X1 npu_inst_pe_1_5_6_U39 ( .A1(npu_inst_int_data_res_6__6__5_), .A2(
        npu_inst_pe_1_5_6_n1), .B1(npu_inst_pe_1_5_6_N78), .B2(
        npu_inst_pe_1_5_6_n76), .C1(npu_inst_pe_1_5_6_N70), .C2(
        npu_inst_pe_1_5_6_n77), .ZN(npu_inst_pe_1_5_6_n79) );
  INV_X1 npu_inst_pe_1_5_6_U38 ( .A(npu_inst_pe_1_5_6_n79), .ZN(
        npu_inst_pe_1_5_6_n35) );
  AOI222_X1 npu_inst_pe_1_5_6_U37 ( .A1(npu_inst_int_data_res_6__6__6_), .A2(
        npu_inst_pe_1_5_6_n1), .B1(npu_inst_pe_1_5_6_N79), .B2(
        npu_inst_pe_1_5_6_n76), .C1(npu_inst_pe_1_5_6_N71), .C2(
        npu_inst_pe_1_5_6_n77), .ZN(npu_inst_pe_1_5_6_n78) );
  INV_X1 npu_inst_pe_1_5_6_U36 ( .A(npu_inst_pe_1_5_6_n78), .ZN(
        npu_inst_pe_1_5_6_n34) );
  INV_X1 npu_inst_pe_1_5_6_U35 ( .A(npu_inst_pe_1_5_6_int_data_1_), .ZN(
        npu_inst_pe_1_5_6_n14) );
  AND2_X1 npu_inst_pe_1_5_6_U34 ( .A1(npu_inst_int_data_x_5__6__1_), .A2(
        npu_inst_pe_1_5_6_int_q_weight_1_), .ZN(npu_inst_pe_1_5_6_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_5_6_U33 ( .A1(npu_inst_int_data_x_5__6__0_), .A2(
        npu_inst_pe_1_5_6_int_q_weight_1_), .ZN(npu_inst_pe_1_5_6_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_5_6_U32 ( .A1(npu_inst_n54), .A2(
        npu_inst_int_data_y_6__6__1_), .B1(npu_inst_pe_1_5_6_n3), .B2(
        npu_inst_int_data_x_5__7__1_), .ZN(npu_inst_pe_1_5_6_n63) );
  AOI22_X1 npu_inst_pe_1_5_6_U31 ( .A1(npu_inst_n54), .A2(
        npu_inst_int_data_y_6__6__0_), .B1(npu_inst_pe_1_5_6_n3), .B2(
        npu_inst_int_data_x_5__7__0_), .ZN(npu_inst_pe_1_5_6_n61) );
  INV_X1 npu_inst_pe_1_5_6_U30 ( .A(npu_inst_pe_1_5_6_int_data_0_), .ZN(
        npu_inst_pe_1_5_6_n13) );
  INV_X1 npu_inst_pe_1_5_6_U29 ( .A(npu_inst_n68), .ZN(npu_inst_pe_1_5_6_n5)
         );
  OR3_X1 npu_inst_pe_1_5_6_U28 ( .A1(npu_inst_pe_1_5_6_n6), .A2(
        npu_inst_pe_1_5_6_n8), .A3(npu_inst_pe_1_5_6_n5), .ZN(
        npu_inst_pe_1_5_6_n56) );
  OR3_X1 npu_inst_pe_1_5_6_U27 ( .A1(npu_inst_pe_1_5_6_n5), .A2(
        npu_inst_pe_1_5_6_n8), .A3(npu_inst_pe_1_5_6_n7), .ZN(
        npu_inst_pe_1_5_6_n48) );
  INV_X1 npu_inst_pe_1_5_6_U26 ( .A(npu_inst_pe_1_5_6_n5), .ZN(
        npu_inst_pe_1_5_6_n4) );
  INV_X1 npu_inst_pe_1_5_6_U25 ( .A(npu_inst_n123), .ZN(npu_inst_pe_1_5_6_n12)
         );
  OR3_X1 npu_inst_pe_1_5_6_U24 ( .A1(npu_inst_pe_1_5_6_n4), .A2(
        npu_inst_pe_1_5_6_n8), .A3(npu_inst_pe_1_5_6_n7), .ZN(
        npu_inst_pe_1_5_6_n52) );
  OR3_X1 npu_inst_pe_1_5_6_U23 ( .A1(npu_inst_pe_1_5_6_n6), .A2(
        npu_inst_pe_1_5_6_n8), .A3(npu_inst_pe_1_5_6_n4), .ZN(
        npu_inst_pe_1_5_6_n60) );
  NOR2_X1 npu_inst_pe_1_5_6_U22 ( .A1(npu_inst_pe_1_5_6_n60), .A2(
        npu_inst_pe_1_5_6_n3), .ZN(npu_inst_pe_1_5_6_n58) );
  NOR2_X1 npu_inst_pe_1_5_6_U21 ( .A1(npu_inst_pe_1_5_6_n56), .A2(
        npu_inst_pe_1_5_6_n3), .ZN(npu_inst_pe_1_5_6_n54) );
  NOR2_X1 npu_inst_pe_1_5_6_U20 ( .A1(npu_inst_pe_1_5_6_n52), .A2(
        npu_inst_pe_1_5_6_n3), .ZN(npu_inst_pe_1_5_6_n50) );
  NOR2_X1 npu_inst_pe_1_5_6_U19 ( .A1(npu_inst_pe_1_5_6_n48), .A2(
        npu_inst_pe_1_5_6_n3), .ZN(npu_inst_pe_1_5_6_n46) );
  NOR2_X1 npu_inst_pe_1_5_6_U18 ( .A1(npu_inst_pe_1_5_6_n40), .A2(
        npu_inst_pe_1_5_6_n3), .ZN(npu_inst_pe_1_5_6_n38) );
  NOR2_X1 npu_inst_pe_1_5_6_U17 ( .A1(npu_inst_pe_1_5_6_n44), .A2(
        npu_inst_pe_1_5_6_n3), .ZN(npu_inst_pe_1_5_6_n42) );
  BUF_X1 npu_inst_pe_1_5_6_U16 ( .A(npu_inst_n96), .Z(npu_inst_pe_1_5_6_n8) );
  BUF_X1 npu_inst_pe_1_5_6_U15 ( .A(npu_inst_pe_1_5_6_n12), .Z(
        npu_inst_pe_1_5_6_n11) );
  BUF_X1 npu_inst_pe_1_5_6_U14 ( .A(npu_inst_pe_1_5_6_n12), .Z(
        npu_inst_pe_1_5_6_n10) );
  BUF_X1 npu_inst_pe_1_5_6_U13 ( .A(npu_inst_pe_1_5_6_n12), .Z(
        npu_inst_pe_1_5_6_n9) );
  INV_X1 npu_inst_pe_1_5_6_U12 ( .A(npu_inst_pe_1_5_6_n38), .ZN(
        npu_inst_pe_1_5_6_n118) );
  INV_X1 npu_inst_pe_1_5_6_U11 ( .A(npu_inst_pe_1_5_6_n58), .ZN(
        npu_inst_pe_1_5_6_n114) );
  INV_X1 npu_inst_pe_1_5_6_U10 ( .A(npu_inst_pe_1_5_6_n54), .ZN(
        npu_inst_pe_1_5_6_n115) );
  INV_X1 npu_inst_pe_1_5_6_U9 ( .A(npu_inst_pe_1_5_6_n50), .ZN(
        npu_inst_pe_1_5_6_n116) );
  INV_X1 npu_inst_pe_1_5_6_U8 ( .A(npu_inst_pe_1_5_6_n46), .ZN(
        npu_inst_pe_1_5_6_n117) );
  INV_X1 npu_inst_pe_1_5_6_U7 ( .A(npu_inst_pe_1_5_6_n42), .ZN(
        npu_inst_pe_1_5_6_n119) );
  BUF_X1 npu_inst_pe_1_5_6_U6 ( .A(npu_inst_n15), .Z(npu_inst_pe_1_5_6_n2) );
  BUF_X1 npu_inst_pe_1_5_6_U5 ( .A(npu_inst_n15), .Z(npu_inst_pe_1_5_6_n1) );
  NOR2_X1 npu_inst_pe_1_5_6_U4 ( .A1(npu_inst_pe_1_5_6_int_q_weight_0_), .A2(
        npu_inst_pe_1_5_6_n1), .ZN(npu_inst_pe_1_5_6_n76) );
  NOR2_X1 npu_inst_pe_1_5_6_U3 ( .A1(npu_inst_pe_1_5_6_n27), .A2(
        npu_inst_pe_1_5_6_n1), .ZN(npu_inst_pe_1_5_6_n77) );
  FA_X1 npu_inst_pe_1_5_6_sub_77_U2_1 ( .A(npu_inst_pe_1_5_6_int_q_acc_1_), 
        .B(npu_inst_pe_1_5_6_n14), .CI(npu_inst_pe_1_5_6_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_5_6_sub_77_carry_2_), .S(npu_inst_pe_1_5_6_N66) );
  FA_X1 npu_inst_pe_1_5_6_add_79_U1_1 ( .A(npu_inst_pe_1_5_6_int_q_acc_1_), 
        .B(npu_inst_pe_1_5_6_int_data_1_), .CI(
        npu_inst_pe_1_5_6_add_79_carry_1_), .CO(
        npu_inst_pe_1_5_6_add_79_carry_2_), .S(npu_inst_pe_1_5_6_N74) );
  NAND3_X1 npu_inst_pe_1_5_6_U109 ( .A1(npu_inst_pe_1_5_6_n5), .A2(
        npu_inst_pe_1_5_6_n7), .A3(npu_inst_pe_1_5_6_n8), .ZN(
        npu_inst_pe_1_5_6_n44) );
  NAND3_X1 npu_inst_pe_1_5_6_U108 ( .A1(npu_inst_pe_1_5_6_n4), .A2(
        npu_inst_pe_1_5_6_n7), .A3(npu_inst_pe_1_5_6_n8), .ZN(
        npu_inst_pe_1_5_6_n40) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_5_6_n34), .CK(
        npu_inst_pe_1_5_6_net3235), .RN(npu_inst_pe_1_5_6_n9), .Q(
        npu_inst_pe_1_5_6_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_5_6_n35), .CK(
        npu_inst_pe_1_5_6_net3235), .RN(npu_inst_pe_1_5_6_n9), .Q(
        npu_inst_pe_1_5_6_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_5_6_n36), .CK(
        npu_inst_pe_1_5_6_net3235), .RN(npu_inst_pe_1_5_6_n9), .Q(
        npu_inst_pe_1_5_6_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_5_6_n98), .CK(
        npu_inst_pe_1_5_6_net3235), .RN(npu_inst_pe_1_5_6_n9), .Q(
        npu_inst_pe_1_5_6_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_5_6_n99), .CK(
        npu_inst_pe_1_5_6_net3235), .RN(npu_inst_pe_1_5_6_n9), .Q(
        npu_inst_pe_1_5_6_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_5_6_n100), 
        .CK(npu_inst_pe_1_5_6_net3235), .RN(npu_inst_pe_1_5_6_n9), .Q(
        npu_inst_pe_1_5_6_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_5_6_n33), .CK(
        npu_inst_pe_1_5_6_net3235), .RN(npu_inst_pe_1_5_6_n9), .Q(
        npu_inst_pe_1_5_6_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_5_6_n101), 
        .CK(npu_inst_pe_1_5_6_net3235), .RN(npu_inst_pe_1_5_6_n9), .Q(
        npu_inst_pe_1_5_6_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_weight_reg_0_ ( .D(npu_inst_n109), .CK(
        npu_inst_pe_1_5_6_net3241), .RN(npu_inst_pe_1_5_6_n9), .Q(
        npu_inst_pe_1_5_6_int_q_weight_0_), .QN(npu_inst_pe_1_5_6_n27) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_weight_reg_1_ ( .D(npu_inst_n115), .CK(
        npu_inst_pe_1_5_6_net3241), .RN(npu_inst_pe_1_5_6_n9), .Q(
        npu_inst_pe_1_5_6_int_q_weight_1_), .QN(npu_inst_pe_1_5_6_n26) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_5_6_n113), 
        .CK(npu_inst_pe_1_5_6_net3241), .RN(npu_inst_pe_1_5_6_n9), .Q(
        npu_inst_pe_1_5_6_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_5_6_n107), 
        .CK(npu_inst_pe_1_5_6_net3241), .RN(npu_inst_pe_1_5_6_n9), .Q(
        npu_inst_pe_1_5_6_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_5_6_n112), 
        .CK(npu_inst_pe_1_5_6_net3241), .RN(npu_inst_pe_1_5_6_n10), .Q(
        npu_inst_pe_1_5_6_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_5_6_n106), 
        .CK(npu_inst_pe_1_5_6_net3241), .RN(npu_inst_pe_1_5_6_n10), .Q(
        npu_inst_pe_1_5_6_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_5_6_n111), 
        .CK(npu_inst_pe_1_5_6_net3241), .RN(npu_inst_pe_1_5_6_n10), .Q(
        npu_inst_pe_1_5_6_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_5_6_n105), 
        .CK(npu_inst_pe_1_5_6_net3241), .RN(npu_inst_pe_1_5_6_n10), .Q(
        npu_inst_pe_1_5_6_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_5_6_n110), 
        .CK(npu_inst_pe_1_5_6_net3241), .RN(npu_inst_pe_1_5_6_n10), .Q(
        npu_inst_pe_1_5_6_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_5_6_n104), 
        .CK(npu_inst_pe_1_5_6_net3241), .RN(npu_inst_pe_1_5_6_n10), .Q(
        npu_inst_pe_1_5_6_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_5_6_n109), 
        .CK(npu_inst_pe_1_5_6_net3241), .RN(npu_inst_pe_1_5_6_n10), .Q(
        npu_inst_pe_1_5_6_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_5_6_n103), 
        .CK(npu_inst_pe_1_5_6_net3241), .RN(npu_inst_pe_1_5_6_n10), .Q(
        npu_inst_pe_1_5_6_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_5_6_n108), 
        .CK(npu_inst_pe_1_5_6_net3241), .RN(npu_inst_pe_1_5_6_n10), .Q(
        npu_inst_pe_1_5_6_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_5_6_n102), 
        .CK(npu_inst_pe_1_5_6_net3241), .RN(npu_inst_pe_1_5_6_n10), .Q(
        npu_inst_pe_1_5_6_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_5_6_n86), 
        .CK(npu_inst_pe_1_5_6_net3241), .RN(npu_inst_pe_1_5_6_n10), .Q(
        npu_inst_pe_1_5_6_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_5_6_n87), 
        .CK(npu_inst_pe_1_5_6_net3241), .RN(npu_inst_pe_1_5_6_n10), .Q(
        npu_inst_pe_1_5_6_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_5_6_n88), 
        .CK(npu_inst_pe_1_5_6_net3241), .RN(npu_inst_pe_1_5_6_n11), .Q(
        npu_inst_pe_1_5_6_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_5_6_n89), 
        .CK(npu_inst_pe_1_5_6_net3241), .RN(npu_inst_pe_1_5_6_n11), .Q(
        npu_inst_pe_1_5_6_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_5_6_n90), 
        .CK(npu_inst_pe_1_5_6_net3241), .RN(npu_inst_pe_1_5_6_n11), .Q(
        npu_inst_pe_1_5_6_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_5_6_n91), 
        .CK(npu_inst_pe_1_5_6_net3241), .RN(npu_inst_pe_1_5_6_n11), .Q(
        npu_inst_pe_1_5_6_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_5_6_n92), 
        .CK(npu_inst_pe_1_5_6_net3241), .RN(npu_inst_pe_1_5_6_n11), .Q(
        npu_inst_pe_1_5_6_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_5_6_n93), 
        .CK(npu_inst_pe_1_5_6_net3241), .RN(npu_inst_pe_1_5_6_n11), .Q(
        npu_inst_pe_1_5_6_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_5_6_n94), 
        .CK(npu_inst_pe_1_5_6_net3241), .RN(npu_inst_pe_1_5_6_n11), .Q(
        npu_inst_pe_1_5_6_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_5_6_n95), 
        .CK(npu_inst_pe_1_5_6_net3241), .RN(npu_inst_pe_1_5_6_n11), .Q(
        npu_inst_pe_1_5_6_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_5_6_n96), 
        .CK(npu_inst_pe_1_5_6_net3241), .RN(npu_inst_pe_1_5_6_n11), .Q(
        npu_inst_pe_1_5_6_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_5_6_n97), 
        .CK(npu_inst_pe_1_5_6_net3241), .RN(npu_inst_pe_1_5_6_n11), .Q(
        npu_inst_pe_1_5_6_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_5_6_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_5_6_N84), .SE(1'b0), .GCK(npu_inst_pe_1_5_6_net3235) );
  CLKGATETST_X1 npu_inst_pe_1_5_6_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n62), .SE(1'b0), .GCK(npu_inst_pe_1_5_6_net3241) );
  MUX2_X1 npu_inst_pe_1_5_7_U162 ( .A(npu_inst_pe_1_5_7_n32), .B(
        npu_inst_pe_1_5_7_n29), .S(npu_inst_pe_1_5_7_n8), .Z(
        npu_inst_pe_1_5_7_N93) );
  MUX2_X1 npu_inst_pe_1_5_7_U161 ( .A(npu_inst_pe_1_5_7_n31), .B(
        npu_inst_pe_1_5_7_n30), .S(npu_inst_pe_1_5_7_n6), .Z(
        npu_inst_pe_1_5_7_n32) );
  MUX2_X1 npu_inst_pe_1_5_7_U160 ( .A(npu_inst_pe_1_5_7_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_5_7_int_q_reg_v_1__0_), .S(npu_inst_pe_1_5_7_n4), .Z(
        npu_inst_pe_1_5_7_n31) );
  MUX2_X1 npu_inst_pe_1_5_7_U159 ( .A(npu_inst_pe_1_5_7_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_5_7_int_q_reg_v_3__0_), .S(npu_inst_pe_1_5_7_n4), .Z(
        npu_inst_pe_1_5_7_n30) );
  MUX2_X1 npu_inst_pe_1_5_7_U158 ( .A(npu_inst_pe_1_5_7_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_5_7_int_q_reg_v_5__0_), .S(npu_inst_pe_1_5_7_n4), .Z(
        npu_inst_pe_1_5_7_n29) );
  MUX2_X1 npu_inst_pe_1_5_7_U157 ( .A(npu_inst_pe_1_5_7_n28), .B(
        npu_inst_pe_1_5_7_n23), .S(npu_inst_pe_1_5_7_n8), .Z(
        npu_inst_pe_1_5_7_N94) );
  MUX2_X1 npu_inst_pe_1_5_7_U156 ( .A(npu_inst_pe_1_5_7_n25), .B(
        npu_inst_pe_1_5_7_n24), .S(npu_inst_pe_1_5_7_n6), .Z(
        npu_inst_pe_1_5_7_n28) );
  MUX2_X1 npu_inst_pe_1_5_7_U155 ( .A(npu_inst_pe_1_5_7_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_5_7_int_q_reg_v_1__1_), .S(npu_inst_pe_1_5_7_n4), .Z(
        npu_inst_pe_1_5_7_n25) );
  MUX2_X1 npu_inst_pe_1_5_7_U154 ( .A(npu_inst_pe_1_5_7_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_5_7_int_q_reg_v_3__1_), .S(npu_inst_pe_1_5_7_n4), .Z(
        npu_inst_pe_1_5_7_n24) );
  MUX2_X1 npu_inst_pe_1_5_7_U153 ( .A(npu_inst_pe_1_5_7_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_5_7_int_q_reg_v_5__1_), .S(npu_inst_pe_1_5_7_n4), .Z(
        npu_inst_pe_1_5_7_n23) );
  MUX2_X1 npu_inst_pe_1_5_7_U152 ( .A(npu_inst_pe_1_5_7_n22), .B(
        npu_inst_pe_1_5_7_n19), .S(npu_inst_pe_1_5_7_n8), .Z(
        npu_inst_int_data_x_5__7__1_) );
  MUX2_X1 npu_inst_pe_1_5_7_U151 ( .A(npu_inst_pe_1_5_7_n21), .B(
        npu_inst_pe_1_5_7_n20), .S(npu_inst_pe_1_5_7_n6), .Z(
        npu_inst_pe_1_5_7_n22) );
  MUX2_X1 npu_inst_pe_1_5_7_U150 ( .A(npu_inst_pe_1_5_7_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_5_7_int_q_reg_h_1__1_), .S(npu_inst_pe_1_5_7_n4), .Z(
        npu_inst_pe_1_5_7_n21) );
  MUX2_X1 npu_inst_pe_1_5_7_U149 ( .A(npu_inst_pe_1_5_7_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_5_7_int_q_reg_h_3__1_), .S(npu_inst_pe_1_5_7_n4), .Z(
        npu_inst_pe_1_5_7_n20) );
  MUX2_X1 npu_inst_pe_1_5_7_U148 ( .A(npu_inst_pe_1_5_7_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_5_7_int_q_reg_h_5__1_), .S(npu_inst_pe_1_5_7_n4), .Z(
        npu_inst_pe_1_5_7_n19) );
  MUX2_X1 npu_inst_pe_1_5_7_U147 ( .A(npu_inst_pe_1_5_7_n18), .B(
        npu_inst_pe_1_5_7_n15), .S(npu_inst_pe_1_5_7_n8), .Z(
        npu_inst_int_data_x_5__7__0_) );
  MUX2_X1 npu_inst_pe_1_5_7_U146 ( .A(npu_inst_pe_1_5_7_n17), .B(
        npu_inst_pe_1_5_7_n16), .S(npu_inst_pe_1_5_7_n6), .Z(
        npu_inst_pe_1_5_7_n18) );
  MUX2_X1 npu_inst_pe_1_5_7_U145 ( .A(npu_inst_pe_1_5_7_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_5_7_int_q_reg_h_1__0_), .S(npu_inst_pe_1_5_7_n4), .Z(
        npu_inst_pe_1_5_7_n17) );
  MUX2_X1 npu_inst_pe_1_5_7_U144 ( .A(npu_inst_pe_1_5_7_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_5_7_int_q_reg_h_3__0_), .S(npu_inst_pe_1_5_7_n4), .Z(
        npu_inst_pe_1_5_7_n16) );
  MUX2_X1 npu_inst_pe_1_5_7_U143 ( .A(npu_inst_pe_1_5_7_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_5_7_int_q_reg_h_5__0_), .S(npu_inst_pe_1_5_7_n4), .Z(
        npu_inst_pe_1_5_7_n15) );
  XOR2_X1 npu_inst_pe_1_5_7_U142 ( .A(npu_inst_pe_1_5_7_int_data_0_), .B(
        npu_inst_pe_1_5_7_int_q_acc_0_), .Z(npu_inst_pe_1_5_7_N73) );
  AND2_X1 npu_inst_pe_1_5_7_U141 ( .A1(npu_inst_pe_1_5_7_int_q_acc_0_), .A2(
        npu_inst_pe_1_5_7_int_data_0_), .ZN(npu_inst_pe_1_5_7_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_5_7_U140 ( .A(npu_inst_pe_1_5_7_int_q_acc_0_), .B(
        npu_inst_pe_1_5_7_n13), .ZN(npu_inst_pe_1_5_7_N65) );
  OR2_X1 npu_inst_pe_1_5_7_U139 ( .A1(npu_inst_pe_1_5_7_n13), .A2(
        npu_inst_pe_1_5_7_int_q_acc_0_), .ZN(npu_inst_pe_1_5_7_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_5_7_U138 ( .A(npu_inst_pe_1_5_7_int_q_acc_2_), .B(
        npu_inst_pe_1_5_7_add_79_carry_2_), .Z(npu_inst_pe_1_5_7_N75) );
  AND2_X1 npu_inst_pe_1_5_7_U137 ( .A1(npu_inst_pe_1_5_7_add_79_carry_2_), 
        .A2(npu_inst_pe_1_5_7_int_q_acc_2_), .ZN(
        npu_inst_pe_1_5_7_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_5_7_U136 ( .A(npu_inst_pe_1_5_7_int_q_acc_3_), .B(
        npu_inst_pe_1_5_7_add_79_carry_3_), .Z(npu_inst_pe_1_5_7_N76) );
  AND2_X1 npu_inst_pe_1_5_7_U135 ( .A1(npu_inst_pe_1_5_7_add_79_carry_3_), 
        .A2(npu_inst_pe_1_5_7_int_q_acc_3_), .ZN(
        npu_inst_pe_1_5_7_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_5_7_U134 ( .A(npu_inst_pe_1_5_7_int_q_acc_4_), .B(
        npu_inst_pe_1_5_7_add_79_carry_4_), .Z(npu_inst_pe_1_5_7_N77) );
  AND2_X1 npu_inst_pe_1_5_7_U133 ( .A1(npu_inst_pe_1_5_7_add_79_carry_4_), 
        .A2(npu_inst_pe_1_5_7_int_q_acc_4_), .ZN(
        npu_inst_pe_1_5_7_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_5_7_U132 ( .A(npu_inst_pe_1_5_7_int_q_acc_5_), .B(
        npu_inst_pe_1_5_7_add_79_carry_5_), .Z(npu_inst_pe_1_5_7_N78) );
  AND2_X1 npu_inst_pe_1_5_7_U131 ( .A1(npu_inst_pe_1_5_7_add_79_carry_5_), 
        .A2(npu_inst_pe_1_5_7_int_q_acc_5_), .ZN(
        npu_inst_pe_1_5_7_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_5_7_U130 ( .A(npu_inst_pe_1_5_7_int_q_acc_6_), .B(
        npu_inst_pe_1_5_7_add_79_carry_6_), .Z(npu_inst_pe_1_5_7_N79) );
  AND2_X1 npu_inst_pe_1_5_7_U129 ( .A1(npu_inst_pe_1_5_7_add_79_carry_6_), 
        .A2(npu_inst_pe_1_5_7_int_q_acc_6_), .ZN(
        npu_inst_pe_1_5_7_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_5_7_U128 ( .A(npu_inst_pe_1_5_7_int_q_acc_7_), .B(
        npu_inst_pe_1_5_7_add_79_carry_7_), .Z(npu_inst_pe_1_5_7_N80) );
  XNOR2_X1 npu_inst_pe_1_5_7_U127 ( .A(npu_inst_pe_1_5_7_sub_77_carry_2_), .B(
        npu_inst_pe_1_5_7_int_q_acc_2_), .ZN(npu_inst_pe_1_5_7_N67) );
  OR2_X1 npu_inst_pe_1_5_7_U126 ( .A1(npu_inst_pe_1_5_7_int_q_acc_2_), .A2(
        npu_inst_pe_1_5_7_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_5_7_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_5_7_U125 ( .A(npu_inst_pe_1_5_7_sub_77_carry_3_), .B(
        npu_inst_pe_1_5_7_int_q_acc_3_), .ZN(npu_inst_pe_1_5_7_N68) );
  OR2_X1 npu_inst_pe_1_5_7_U124 ( .A1(npu_inst_pe_1_5_7_int_q_acc_3_), .A2(
        npu_inst_pe_1_5_7_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_5_7_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_5_7_U123 ( .A(npu_inst_pe_1_5_7_sub_77_carry_4_), .B(
        npu_inst_pe_1_5_7_int_q_acc_4_), .ZN(npu_inst_pe_1_5_7_N69) );
  OR2_X1 npu_inst_pe_1_5_7_U122 ( .A1(npu_inst_pe_1_5_7_int_q_acc_4_), .A2(
        npu_inst_pe_1_5_7_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_5_7_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_5_7_U121 ( .A(npu_inst_pe_1_5_7_sub_77_carry_5_), .B(
        npu_inst_pe_1_5_7_int_q_acc_5_), .ZN(npu_inst_pe_1_5_7_N70) );
  OR2_X1 npu_inst_pe_1_5_7_U120 ( .A1(npu_inst_pe_1_5_7_int_q_acc_5_), .A2(
        npu_inst_pe_1_5_7_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_5_7_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_5_7_U119 ( .A(npu_inst_pe_1_5_7_sub_77_carry_6_), .B(
        npu_inst_pe_1_5_7_int_q_acc_6_), .ZN(npu_inst_pe_1_5_7_N71) );
  OR2_X1 npu_inst_pe_1_5_7_U118 ( .A1(npu_inst_pe_1_5_7_int_q_acc_6_), .A2(
        npu_inst_pe_1_5_7_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_5_7_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_5_7_U117 ( .A(npu_inst_pe_1_5_7_int_q_acc_7_), .B(
        npu_inst_pe_1_5_7_sub_77_carry_7_), .ZN(npu_inst_pe_1_5_7_N72) );
  INV_X1 npu_inst_pe_1_5_7_U116 ( .A(npu_inst_n76), .ZN(npu_inst_pe_1_5_7_n7)
         );
  INV_X1 npu_inst_pe_1_5_7_U115 ( .A(npu_inst_pe_1_5_7_n7), .ZN(
        npu_inst_pe_1_5_7_n6) );
  INV_X1 npu_inst_pe_1_5_7_U114 ( .A(npu_inst_n54), .ZN(npu_inst_pe_1_5_7_n3)
         );
  AOI22_X1 npu_inst_pe_1_5_7_U113 ( .A1(npu_inst_int_data_y_6__7__0_), .A2(
        npu_inst_pe_1_5_7_n58), .B1(npu_inst_pe_1_5_7_n114), .B2(
        npu_inst_pe_1_5_7_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_5_7_n57) );
  INV_X1 npu_inst_pe_1_5_7_U112 ( .A(npu_inst_pe_1_5_7_n57), .ZN(
        npu_inst_pe_1_5_7_n108) );
  AOI22_X1 npu_inst_pe_1_5_7_U111 ( .A1(npu_inst_int_data_y_6__7__0_), .A2(
        npu_inst_pe_1_5_7_n54), .B1(npu_inst_pe_1_5_7_n115), .B2(
        npu_inst_pe_1_5_7_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_5_7_n53) );
  INV_X1 npu_inst_pe_1_5_7_U110 ( .A(npu_inst_pe_1_5_7_n53), .ZN(
        npu_inst_pe_1_5_7_n109) );
  AOI22_X1 npu_inst_pe_1_5_7_U107 ( .A1(npu_inst_int_data_y_6__7__0_), .A2(
        npu_inst_pe_1_5_7_n50), .B1(npu_inst_pe_1_5_7_n116), .B2(
        npu_inst_pe_1_5_7_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_5_7_n49) );
  INV_X1 npu_inst_pe_1_5_7_U106 ( .A(npu_inst_pe_1_5_7_n49), .ZN(
        npu_inst_pe_1_5_7_n110) );
  AOI22_X1 npu_inst_pe_1_5_7_U105 ( .A1(npu_inst_int_data_y_6__7__0_), .A2(
        npu_inst_pe_1_5_7_n46), .B1(npu_inst_pe_1_5_7_n117), .B2(
        npu_inst_pe_1_5_7_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_5_7_n45) );
  INV_X1 npu_inst_pe_1_5_7_U104 ( .A(npu_inst_pe_1_5_7_n45), .ZN(
        npu_inst_pe_1_5_7_n111) );
  AOI22_X1 npu_inst_pe_1_5_7_U103 ( .A1(npu_inst_int_data_y_6__7__0_), .A2(
        npu_inst_pe_1_5_7_n42), .B1(npu_inst_pe_1_5_7_n119), .B2(
        npu_inst_pe_1_5_7_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_5_7_n41) );
  INV_X1 npu_inst_pe_1_5_7_U102 ( .A(npu_inst_pe_1_5_7_n41), .ZN(
        npu_inst_pe_1_5_7_n112) );
  AOI22_X1 npu_inst_pe_1_5_7_U101 ( .A1(npu_inst_int_data_y_6__7__1_), .A2(
        npu_inst_pe_1_5_7_n58), .B1(npu_inst_pe_1_5_7_n114), .B2(
        npu_inst_pe_1_5_7_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_5_7_n59) );
  INV_X1 npu_inst_pe_1_5_7_U100 ( .A(npu_inst_pe_1_5_7_n59), .ZN(
        npu_inst_pe_1_5_7_n102) );
  AOI22_X1 npu_inst_pe_1_5_7_U99 ( .A1(npu_inst_int_data_y_6__7__1_), .A2(
        npu_inst_pe_1_5_7_n54), .B1(npu_inst_pe_1_5_7_n115), .B2(
        npu_inst_pe_1_5_7_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_5_7_n55) );
  INV_X1 npu_inst_pe_1_5_7_U98 ( .A(npu_inst_pe_1_5_7_n55), .ZN(
        npu_inst_pe_1_5_7_n103) );
  AOI22_X1 npu_inst_pe_1_5_7_U97 ( .A1(npu_inst_int_data_y_6__7__1_), .A2(
        npu_inst_pe_1_5_7_n50), .B1(npu_inst_pe_1_5_7_n116), .B2(
        npu_inst_pe_1_5_7_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_5_7_n51) );
  INV_X1 npu_inst_pe_1_5_7_U96 ( .A(npu_inst_pe_1_5_7_n51), .ZN(
        npu_inst_pe_1_5_7_n104) );
  AOI22_X1 npu_inst_pe_1_5_7_U95 ( .A1(npu_inst_int_data_y_6__7__1_), .A2(
        npu_inst_pe_1_5_7_n46), .B1(npu_inst_pe_1_5_7_n117), .B2(
        npu_inst_pe_1_5_7_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_5_7_n47) );
  INV_X1 npu_inst_pe_1_5_7_U94 ( .A(npu_inst_pe_1_5_7_n47), .ZN(
        npu_inst_pe_1_5_7_n105) );
  AOI22_X1 npu_inst_pe_1_5_7_U93 ( .A1(npu_inst_int_data_y_6__7__1_), .A2(
        npu_inst_pe_1_5_7_n42), .B1(npu_inst_pe_1_5_7_n119), .B2(
        npu_inst_pe_1_5_7_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_5_7_n43) );
  INV_X1 npu_inst_pe_1_5_7_U92 ( .A(npu_inst_pe_1_5_7_n43), .ZN(
        npu_inst_pe_1_5_7_n106) );
  AOI22_X1 npu_inst_pe_1_5_7_U91 ( .A1(npu_inst_pe_1_5_7_n38), .A2(
        npu_inst_int_data_y_6__7__1_), .B1(npu_inst_pe_1_5_7_n118), .B2(
        npu_inst_pe_1_5_7_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_5_7_n39) );
  INV_X1 npu_inst_pe_1_5_7_U90 ( .A(npu_inst_pe_1_5_7_n39), .ZN(
        npu_inst_pe_1_5_7_n107) );
  AOI22_X1 npu_inst_pe_1_5_7_U89 ( .A1(npu_inst_pe_1_5_7_n38), .A2(
        npu_inst_int_data_y_6__7__0_), .B1(npu_inst_pe_1_5_7_n118), .B2(
        npu_inst_pe_1_5_7_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_5_7_n37) );
  INV_X1 npu_inst_pe_1_5_7_U88 ( .A(npu_inst_pe_1_5_7_n37), .ZN(
        npu_inst_pe_1_5_7_n113) );
  AND2_X1 npu_inst_pe_1_5_7_U87 ( .A1(npu_inst_pe_1_5_7_N93), .A2(npu_inst_n54), .ZN(npu_inst_int_data_y_5__7__0_) );
  AND2_X1 npu_inst_pe_1_5_7_U86 ( .A1(npu_inst_n54), .A2(npu_inst_pe_1_5_7_N94), .ZN(npu_inst_int_data_y_5__7__1_) );
  NOR3_X1 npu_inst_pe_1_5_7_U85 ( .A1(npu_inst_pe_1_5_7_n26), .A2(npu_inst_n54), .A3(npu_inst_int_ckg[16]), .ZN(npu_inst_pe_1_5_7_n85) );
  OR2_X1 npu_inst_pe_1_5_7_U84 ( .A1(npu_inst_pe_1_5_7_n85), .A2(
        npu_inst_pe_1_5_7_n2), .ZN(npu_inst_pe_1_5_7_N84) );
  AND2_X1 npu_inst_pe_1_5_7_U83 ( .A1(npu_inst_pe_1_5_7_int_q_acc_0_), .A2(
        npu_inst_pe_1_5_7_n1), .ZN(npu_inst_int_data_res_5__7__0_) );
  AND2_X1 npu_inst_pe_1_5_7_U82 ( .A1(npu_inst_pe_1_5_7_n2), .A2(
        npu_inst_pe_1_5_7_int_q_acc_7_), .ZN(npu_inst_int_data_res_5__7__7_)
         );
  AND2_X1 npu_inst_pe_1_5_7_U81 ( .A1(npu_inst_pe_1_5_7_int_q_acc_1_), .A2(
        npu_inst_pe_1_5_7_n1), .ZN(npu_inst_int_data_res_5__7__1_) );
  AND2_X1 npu_inst_pe_1_5_7_U80 ( .A1(npu_inst_pe_1_5_7_int_q_acc_2_), .A2(
        npu_inst_pe_1_5_7_n1), .ZN(npu_inst_int_data_res_5__7__2_) );
  AND2_X1 npu_inst_pe_1_5_7_U79 ( .A1(npu_inst_pe_1_5_7_int_q_acc_3_), .A2(
        npu_inst_pe_1_5_7_n2), .ZN(npu_inst_int_data_res_5__7__3_) );
  AND2_X1 npu_inst_pe_1_5_7_U78 ( .A1(npu_inst_pe_1_5_7_int_q_acc_4_), .A2(
        npu_inst_pe_1_5_7_n2), .ZN(npu_inst_int_data_res_5__7__4_) );
  AND2_X1 npu_inst_pe_1_5_7_U77 ( .A1(npu_inst_pe_1_5_7_int_q_acc_5_), .A2(
        npu_inst_pe_1_5_7_n2), .ZN(npu_inst_int_data_res_5__7__5_) );
  AND2_X1 npu_inst_pe_1_5_7_U76 ( .A1(npu_inst_pe_1_5_7_int_q_acc_6_), .A2(
        npu_inst_pe_1_5_7_n2), .ZN(npu_inst_int_data_res_5__7__6_) );
  AOI222_X1 npu_inst_pe_1_5_7_U75 ( .A1(npu_inst_int_data_res_6__7__0_), .A2(
        npu_inst_pe_1_5_7_n1), .B1(npu_inst_pe_1_5_7_N73), .B2(
        npu_inst_pe_1_5_7_n76), .C1(npu_inst_pe_1_5_7_N65), .C2(
        npu_inst_pe_1_5_7_n77), .ZN(npu_inst_pe_1_5_7_n84) );
  INV_X1 npu_inst_pe_1_5_7_U74 ( .A(npu_inst_pe_1_5_7_n84), .ZN(
        npu_inst_pe_1_5_7_n101) );
  AOI222_X1 npu_inst_pe_1_5_7_U73 ( .A1(npu_inst_int_data_res_6__7__7_), .A2(
        npu_inst_pe_1_5_7_n1), .B1(npu_inst_pe_1_5_7_N80), .B2(
        npu_inst_pe_1_5_7_n76), .C1(npu_inst_pe_1_5_7_N72), .C2(
        npu_inst_pe_1_5_7_n77), .ZN(npu_inst_pe_1_5_7_n75) );
  INV_X1 npu_inst_pe_1_5_7_U72 ( .A(npu_inst_pe_1_5_7_n75), .ZN(
        npu_inst_pe_1_5_7_n33) );
  AOI222_X1 npu_inst_pe_1_5_7_U71 ( .A1(npu_inst_int_data_res_6__7__1_), .A2(
        npu_inst_pe_1_5_7_n1), .B1(npu_inst_pe_1_5_7_N74), .B2(
        npu_inst_pe_1_5_7_n76), .C1(npu_inst_pe_1_5_7_N66), .C2(
        npu_inst_pe_1_5_7_n77), .ZN(npu_inst_pe_1_5_7_n83) );
  INV_X1 npu_inst_pe_1_5_7_U70 ( .A(npu_inst_pe_1_5_7_n83), .ZN(
        npu_inst_pe_1_5_7_n100) );
  AOI222_X1 npu_inst_pe_1_5_7_U69 ( .A1(npu_inst_int_data_res_6__7__2_), .A2(
        npu_inst_pe_1_5_7_n1), .B1(npu_inst_pe_1_5_7_N75), .B2(
        npu_inst_pe_1_5_7_n76), .C1(npu_inst_pe_1_5_7_N67), .C2(
        npu_inst_pe_1_5_7_n77), .ZN(npu_inst_pe_1_5_7_n82) );
  INV_X1 npu_inst_pe_1_5_7_U68 ( .A(npu_inst_pe_1_5_7_n82), .ZN(
        npu_inst_pe_1_5_7_n99) );
  AOI222_X1 npu_inst_pe_1_5_7_U67 ( .A1(npu_inst_int_data_res_6__7__3_), .A2(
        npu_inst_pe_1_5_7_n1), .B1(npu_inst_pe_1_5_7_N76), .B2(
        npu_inst_pe_1_5_7_n76), .C1(npu_inst_pe_1_5_7_N68), .C2(
        npu_inst_pe_1_5_7_n77), .ZN(npu_inst_pe_1_5_7_n81) );
  INV_X1 npu_inst_pe_1_5_7_U66 ( .A(npu_inst_pe_1_5_7_n81), .ZN(
        npu_inst_pe_1_5_7_n98) );
  AOI222_X1 npu_inst_pe_1_5_7_U65 ( .A1(npu_inst_int_data_res_6__7__4_), .A2(
        npu_inst_pe_1_5_7_n1), .B1(npu_inst_pe_1_5_7_N77), .B2(
        npu_inst_pe_1_5_7_n76), .C1(npu_inst_pe_1_5_7_N69), .C2(
        npu_inst_pe_1_5_7_n77), .ZN(npu_inst_pe_1_5_7_n80) );
  INV_X1 npu_inst_pe_1_5_7_U64 ( .A(npu_inst_pe_1_5_7_n80), .ZN(
        npu_inst_pe_1_5_7_n36) );
  AOI222_X1 npu_inst_pe_1_5_7_U63 ( .A1(npu_inst_int_data_res_6__7__5_), .A2(
        npu_inst_pe_1_5_7_n1), .B1(npu_inst_pe_1_5_7_N78), .B2(
        npu_inst_pe_1_5_7_n76), .C1(npu_inst_pe_1_5_7_N70), .C2(
        npu_inst_pe_1_5_7_n77), .ZN(npu_inst_pe_1_5_7_n79) );
  INV_X1 npu_inst_pe_1_5_7_U62 ( .A(npu_inst_pe_1_5_7_n79), .ZN(
        npu_inst_pe_1_5_7_n35) );
  AOI222_X1 npu_inst_pe_1_5_7_U61 ( .A1(npu_inst_int_data_res_6__7__6_), .A2(
        npu_inst_pe_1_5_7_n1), .B1(npu_inst_pe_1_5_7_N79), .B2(
        npu_inst_pe_1_5_7_n76), .C1(npu_inst_pe_1_5_7_N71), .C2(
        npu_inst_pe_1_5_7_n77), .ZN(npu_inst_pe_1_5_7_n78) );
  INV_X1 npu_inst_pe_1_5_7_U60 ( .A(npu_inst_pe_1_5_7_n78), .ZN(
        npu_inst_pe_1_5_7_n34) );
  INV_X1 npu_inst_pe_1_5_7_U59 ( .A(npu_inst_pe_1_5_7_int_data_1_), .ZN(
        npu_inst_pe_1_5_7_n14) );
  AND2_X1 npu_inst_pe_1_5_7_U58 ( .A1(npu_inst_int_data_x_5__7__1_), .A2(
        npu_inst_pe_1_5_7_int_q_weight_1_), .ZN(npu_inst_pe_1_5_7_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_5_7_U57 ( .A1(npu_inst_int_data_x_5__7__0_), .A2(
        npu_inst_pe_1_5_7_int_q_weight_1_), .ZN(npu_inst_pe_1_5_7_int_data_0_)
         );
  NAND2_X1 npu_inst_pe_1_5_7_U56 ( .A1(npu_inst_pe_1_5_7_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_5_7_n60), .ZN(npu_inst_pe_1_5_7_n74) );
  OAI21_X1 npu_inst_pe_1_5_7_U55 ( .B1(npu_inst_pe_1_5_7_n63), .B2(
        npu_inst_pe_1_5_7_n60), .A(npu_inst_pe_1_5_7_n74), .ZN(
        npu_inst_pe_1_5_7_n97) );
  NAND2_X1 npu_inst_pe_1_5_7_U54 ( .A1(npu_inst_pe_1_5_7_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_5_7_n60), .ZN(npu_inst_pe_1_5_7_n73) );
  OAI21_X1 npu_inst_pe_1_5_7_U53 ( .B1(npu_inst_pe_1_5_7_n61), .B2(
        npu_inst_pe_1_5_7_n60), .A(npu_inst_pe_1_5_7_n73), .ZN(
        npu_inst_pe_1_5_7_n96) );
  NAND2_X1 npu_inst_pe_1_5_7_U52 ( .A1(npu_inst_pe_1_5_7_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_5_7_n56), .ZN(npu_inst_pe_1_5_7_n72) );
  OAI21_X1 npu_inst_pe_1_5_7_U51 ( .B1(npu_inst_pe_1_5_7_n63), .B2(
        npu_inst_pe_1_5_7_n56), .A(npu_inst_pe_1_5_7_n72), .ZN(
        npu_inst_pe_1_5_7_n95) );
  NAND2_X1 npu_inst_pe_1_5_7_U50 ( .A1(npu_inst_pe_1_5_7_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_5_7_n56), .ZN(npu_inst_pe_1_5_7_n71) );
  OAI21_X1 npu_inst_pe_1_5_7_U49 ( .B1(npu_inst_pe_1_5_7_n61), .B2(
        npu_inst_pe_1_5_7_n56), .A(npu_inst_pe_1_5_7_n71), .ZN(
        npu_inst_pe_1_5_7_n94) );
  NAND2_X1 npu_inst_pe_1_5_7_U48 ( .A1(npu_inst_pe_1_5_7_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_5_7_n52), .ZN(npu_inst_pe_1_5_7_n70) );
  OAI21_X1 npu_inst_pe_1_5_7_U47 ( .B1(npu_inst_pe_1_5_7_n63), .B2(
        npu_inst_pe_1_5_7_n52), .A(npu_inst_pe_1_5_7_n70), .ZN(
        npu_inst_pe_1_5_7_n93) );
  NAND2_X1 npu_inst_pe_1_5_7_U46 ( .A1(npu_inst_pe_1_5_7_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_5_7_n52), .ZN(npu_inst_pe_1_5_7_n69) );
  OAI21_X1 npu_inst_pe_1_5_7_U45 ( .B1(npu_inst_pe_1_5_7_n61), .B2(
        npu_inst_pe_1_5_7_n52), .A(npu_inst_pe_1_5_7_n69), .ZN(
        npu_inst_pe_1_5_7_n92) );
  NAND2_X1 npu_inst_pe_1_5_7_U44 ( .A1(npu_inst_pe_1_5_7_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_5_7_n48), .ZN(npu_inst_pe_1_5_7_n68) );
  OAI21_X1 npu_inst_pe_1_5_7_U43 ( .B1(npu_inst_pe_1_5_7_n63), .B2(
        npu_inst_pe_1_5_7_n48), .A(npu_inst_pe_1_5_7_n68), .ZN(
        npu_inst_pe_1_5_7_n91) );
  NAND2_X1 npu_inst_pe_1_5_7_U42 ( .A1(npu_inst_pe_1_5_7_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_5_7_n48), .ZN(npu_inst_pe_1_5_7_n67) );
  OAI21_X1 npu_inst_pe_1_5_7_U41 ( .B1(npu_inst_pe_1_5_7_n61), .B2(
        npu_inst_pe_1_5_7_n48), .A(npu_inst_pe_1_5_7_n67), .ZN(
        npu_inst_pe_1_5_7_n90) );
  NAND2_X1 npu_inst_pe_1_5_7_U40 ( .A1(npu_inst_pe_1_5_7_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_5_7_n44), .ZN(npu_inst_pe_1_5_7_n66) );
  OAI21_X1 npu_inst_pe_1_5_7_U39 ( .B1(npu_inst_pe_1_5_7_n63), .B2(
        npu_inst_pe_1_5_7_n44), .A(npu_inst_pe_1_5_7_n66), .ZN(
        npu_inst_pe_1_5_7_n89) );
  NAND2_X1 npu_inst_pe_1_5_7_U38 ( .A1(npu_inst_pe_1_5_7_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_5_7_n44), .ZN(npu_inst_pe_1_5_7_n65) );
  OAI21_X1 npu_inst_pe_1_5_7_U37 ( .B1(npu_inst_pe_1_5_7_n61), .B2(
        npu_inst_pe_1_5_7_n44), .A(npu_inst_pe_1_5_7_n65), .ZN(
        npu_inst_pe_1_5_7_n88) );
  NAND2_X1 npu_inst_pe_1_5_7_U36 ( .A1(npu_inst_pe_1_5_7_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_5_7_n40), .ZN(npu_inst_pe_1_5_7_n64) );
  OAI21_X1 npu_inst_pe_1_5_7_U35 ( .B1(npu_inst_pe_1_5_7_n63), .B2(
        npu_inst_pe_1_5_7_n40), .A(npu_inst_pe_1_5_7_n64), .ZN(
        npu_inst_pe_1_5_7_n87) );
  NAND2_X1 npu_inst_pe_1_5_7_U34 ( .A1(npu_inst_pe_1_5_7_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_5_7_n40), .ZN(npu_inst_pe_1_5_7_n62) );
  OAI21_X1 npu_inst_pe_1_5_7_U33 ( .B1(npu_inst_pe_1_5_7_n61), .B2(
        npu_inst_pe_1_5_7_n40), .A(npu_inst_pe_1_5_7_n62), .ZN(
        npu_inst_pe_1_5_7_n86) );
  INV_X1 npu_inst_pe_1_5_7_U32 ( .A(npu_inst_pe_1_5_7_int_data_0_), .ZN(
        npu_inst_pe_1_5_7_n13) );
  INV_X1 npu_inst_pe_1_5_7_U31 ( .A(npu_inst_n68), .ZN(npu_inst_pe_1_5_7_n5)
         );
  AOI22_X1 npu_inst_pe_1_5_7_U30 ( .A1(npu_inst_n54), .A2(
        npu_inst_int_data_y_6__7__1_), .B1(npu_inst_pe_1_5_7_n3), .B2(
        int_i_data_h_npu6[1]), .ZN(npu_inst_pe_1_5_7_n63) );
  AOI22_X1 npu_inst_pe_1_5_7_U29 ( .A1(npu_inst_n54), .A2(
        npu_inst_int_data_y_6__7__0_), .B1(npu_inst_pe_1_5_7_n3), .B2(
        int_i_data_h_npu6[0]), .ZN(npu_inst_pe_1_5_7_n61) );
  OR3_X1 npu_inst_pe_1_5_7_U28 ( .A1(npu_inst_pe_1_5_7_n6), .A2(
        npu_inst_pe_1_5_7_n8), .A3(npu_inst_pe_1_5_7_n5), .ZN(
        npu_inst_pe_1_5_7_n56) );
  OR3_X1 npu_inst_pe_1_5_7_U27 ( .A1(npu_inst_pe_1_5_7_n5), .A2(
        npu_inst_pe_1_5_7_n8), .A3(npu_inst_pe_1_5_7_n7), .ZN(
        npu_inst_pe_1_5_7_n48) );
  INV_X1 npu_inst_pe_1_5_7_U26 ( .A(npu_inst_pe_1_5_7_n5), .ZN(
        npu_inst_pe_1_5_7_n4) );
  INV_X1 npu_inst_pe_1_5_7_U25 ( .A(npu_inst_n123), .ZN(npu_inst_pe_1_5_7_n12)
         );
  OR3_X1 npu_inst_pe_1_5_7_U24 ( .A1(npu_inst_pe_1_5_7_n4), .A2(
        npu_inst_pe_1_5_7_n8), .A3(npu_inst_pe_1_5_7_n7), .ZN(
        npu_inst_pe_1_5_7_n52) );
  OR3_X1 npu_inst_pe_1_5_7_U23 ( .A1(npu_inst_pe_1_5_7_n6), .A2(
        npu_inst_pe_1_5_7_n8), .A3(npu_inst_pe_1_5_7_n4), .ZN(
        npu_inst_pe_1_5_7_n60) );
  NOR2_X1 npu_inst_pe_1_5_7_U22 ( .A1(npu_inst_pe_1_5_7_n60), .A2(
        npu_inst_pe_1_5_7_n3), .ZN(npu_inst_pe_1_5_7_n58) );
  NOR2_X1 npu_inst_pe_1_5_7_U21 ( .A1(npu_inst_pe_1_5_7_n56), .A2(
        npu_inst_pe_1_5_7_n3), .ZN(npu_inst_pe_1_5_7_n54) );
  NOR2_X1 npu_inst_pe_1_5_7_U20 ( .A1(npu_inst_pe_1_5_7_n52), .A2(
        npu_inst_pe_1_5_7_n3), .ZN(npu_inst_pe_1_5_7_n50) );
  NOR2_X1 npu_inst_pe_1_5_7_U19 ( .A1(npu_inst_pe_1_5_7_n48), .A2(
        npu_inst_pe_1_5_7_n3), .ZN(npu_inst_pe_1_5_7_n46) );
  NOR2_X1 npu_inst_pe_1_5_7_U18 ( .A1(npu_inst_pe_1_5_7_n40), .A2(
        npu_inst_pe_1_5_7_n3), .ZN(npu_inst_pe_1_5_7_n38) );
  NOR2_X1 npu_inst_pe_1_5_7_U17 ( .A1(npu_inst_pe_1_5_7_n44), .A2(
        npu_inst_pe_1_5_7_n3), .ZN(npu_inst_pe_1_5_7_n42) );
  BUF_X1 npu_inst_pe_1_5_7_U16 ( .A(npu_inst_n96), .Z(npu_inst_pe_1_5_7_n8) );
  BUF_X1 npu_inst_pe_1_5_7_U15 ( .A(npu_inst_pe_1_5_7_n12), .Z(
        npu_inst_pe_1_5_7_n11) );
  BUF_X1 npu_inst_pe_1_5_7_U14 ( .A(npu_inst_pe_1_5_7_n12), .Z(
        npu_inst_pe_1_5_7_n10) );
  BUF_X1 npu_inst_pe_1_5_7_U13 ( .A(npu_inst_pe_1_5_7_n12), .Z(
        npu_inst_pe_1_5_7_n9) );
  INV_X1 npu_inst_pe_1_5_7_U12 ( .A(npu_inst_pe_1_5_7_n38), .ZN(
        npu_inst_pe_1_5_7_n118) );
  INV_X1 npu_inst_pe_1_5_7_U11 ( .A(npu_inst_pe_1_5_7_n58), .ZN(
        npu_inst_pe_1_5_7_n114) );
  INV_X1 npu_inst_pe_1_5_7_U10 ( .A(npu_inst_pe_1_5_7_n54), .ZN(
        npu_inst_pe_1_5_7_n115) );
  INV_X1 npu_inst_pe_1_5_7_U9 ( .A(npu_inst_pe_1_5_7_n50), .ZN(
        npu_inst_pe_1_5_7_n116) );
  INV_X1 npu_inst_pe_1_5_7_U8 ( .A(npu_inst_pe_1_5_7_n46), .ZN(
        npu_inst_pe_1_5_7_n117) );
  INV_X1 npu_inst_pe_1_5_7_U7 ( .A(npu_inst_pe_1_5_7_n42), .ZN(
        npu_inst_pe_1_5_7_n119) );
  BUF_X1 npu_inst_pe_1_5_7_U6 ( .A(npu_inst_n15), .Z(npu_inst_pe_1_5_7_n2) );
  BUF_X1 npu_inst_pe_1_5_7_U5 ( .A(npu_inst_n15), .Z(npu_inst_pe_1_5_7_n1) );
  NOR2_X1 npu_inst_pe_1_5_7_U4 ( .A1(npu_inst_pe_1_5_7_int_q_weight_0_), .A2(
        npu_inst_pe_1_5_7_n1), .ZN(npu_inst_pe_1_5_7_n76) );
  NOR2_X1 npu_inst_pe_1_5_7_U3 ( .A1(npu_inst_pe_1_5_7_n27), .A2(
        npu_inst_pe_1_5_7_n1), .ZN(npu_inst_pe_1_5_7_n77) );
  FA_X1 npu_inst_pe_1_5_7_sub_77_U2_1 ( .A(npu_inst_pe_1_5_7_int_q_acc_1_), 
        .B(npu_inst_pe_1_5_7_n14), .CI(npu_inst_pe_1_5_7_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_5_7_sub_77_carry_2_), .S(npu_inst_pe_1_5_7_N66) );
  FA_X1 npu_inst_pe_1_5_7_add_79_U1_1 ( .A(npu_inst_pe_1_5_7_int_q_acc_1_), 
        .B(npu_inst_pe_1_5_7_int_data_1_), .CI(
        npu_inst_pe_1_5_7_add_79_carry_1_), .CO(
        npu_inst_pe_1_5_7_add_79_carry_2_), .S(npu_inst_pe_1_5_7_N74) );
  NAND3_X1 npu_inst_pe_1_5_7_U109 ( .A1(npu_inst_pe_1_5_7_n5), .A2(
        npu_inst_pe_1_5_7_n7), .A3(npu_inst_pe_1_5_7_n8), .ZN(
        npu_inst_pe_1_5_7_n44) );
  NAND3_X1 npu_inst_pe_1_5_7_U108 ( .A1(npu_inst_pe_1_5_7_n4), .A2(
        npu_inst_pe_1_5_7_n7), .A3(npu_inst_pe_1_5_7_n8), .ZN(
        npu_inst_pe_1_5_7_n40) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_5_7_n34), .CK(
        npu_inst_pe_1_5_7_net3212), .RN(npu_inst_pe_1_5_7_n9), .Q(
        npu_inst_pe_1_5_7_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_5_7_n35), .CK(
        npu_inst_pe_1_5_7_net3212), .RN(npu_inst_pe_1_5_7_n9), .Q(
        npu_inst_pe_1_5_7_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_5_7_n36), .CK(
        npu_inst_pe_1_5_7_net3212), .RN(npu_inst_pe_1_5_7_n9), .Q(
        npu_inst_pe_1_5_7_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_5_7_n98), .CK(
        npu_inst_pe_1_5_7_net3212), .RN(npu_inst_pe_1_5_7_n9), .Q(
        npu_inst_pe_1_5_7_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_5_7_n99), .CK(
        npu_inst_pe_1_5_7_net3212), .RN(npu_inst_pe_1_5_7_n9), .Q(
        npu_inst_pe_1_5_7_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_5_7_n100), 
        .CK(npu_inst_pe_1_5_7_net3212), .RN(npu_inst_pe_1_5_7_n9), .Q(
        npu_inst_pe_1_5_7_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_5_7_n33), .CK(
        npu_inst_pe_1_5_7_net3212), .RN(npu_inst_pe_1_5_7_n9), .Q(
        npu_inst_pe_1_5_7_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_5_7_n101), 
        .CK(npu_inst_pe_1_5_7_net3212), .RN(npu_inst_pe_1_5_7_n9), .Q(
        npu_inst_pe_1_5_7_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_weight_reg_0_ ( .D(npu_inst_n109), .CK(
        npu_inst_pe_1_5_7_net3218), .RN(npu_inst_pe_1_5_7_n9), .Q(
        npu_inst_pe_1_5_7_int_q_weight_0_), .QN(npu_inst_pe_1_5_7_n27) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_weight_reg_1_ ( .D(npu_inst_n115), .CK(
        npu_inst_pe_1_5_7_net3218), .RN(npu_inst_pe_1_5_7_n9), .Q(
        npu_inst_pe_1_5_7_int_q_weight_1_), .QN(npu_inst_pe_1_5_7_n26) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_5_7_n113), 
        .CK(npu_inst_pe_1_5_7_net3218), .RN(npu_inst_pe_1_5_7_n9), .Q(
        npu_inst_pe_1_5_7_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_5_7_n107), 
        .CK(npu_inst_pe_1_5_7_net3218), .RN(npu_inst_pe_1_5_7_n9), .Q(
        npu_inst_pe_1_5_7_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_5_7_n112), 
        .CK(npu_inst_pe_1_5_7_net3218), .RN(npu_inst_pe_1_5_7_n10), .Q(
        npu_inst_pe_1_5_7_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_5_7_n106), 
        .CK(npu_inst_pe_1_5_7_net3218), .RN(npu_inst_pe_1_5_7_n10), .Q(
        npu_inst_pe_1_5_7_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_5_7_n111), 
        .CK(npu_inst_pe_1_5_7_net3218), .RN(npu_inst_pe_1_5_7_n10), .Q(
        npu_inst_pe_1_5_7_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_5_7_n105), 
        .CK(npu_inst_pe_1_5_7_net3218), .RN(npu_inst_pe_1_5_7_n10), .Q(
        npu_inst_pe_1_5_7_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_5_7_n110), 
        .CK(npu_inst_pe_1_5_7_net3218), .RN(npu_inst_pe_1_5_7_n10), .Q(
        npu_inst_pe_1_5_7_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_5_7_n104), 
        .CK(npu_inst_pe_1_5_7_net3218), .RN(npu_inst_pe_1_5_7_n10), .Q(
        npu_inst_pe_1_5_7_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_5_7_n109), 
        .CK(npu_inst_pe_1_5_7_net3218), .RN(npu_inst_pe_1_5_7_n10), .Q(
        npu_inst_pe_1_5_7_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_5_7_n103), 
        .CK(npu_inst_pe_1_5_7_net3218), .RN(npu_inst_pe_1_5_7_n10), .Q(
        npu_inst_pe_1_5_7_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_5_7_n108), 
        .CK(npu_inst_pe_1_5_7_net3218), .RN(npu_inst_pe_1_5_7_n10), .Q(
        npu_inst_pe_1_5_7_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_5_7_n102), 
        .CK(npu_inst_pe_1_5_7_net3218), .RN(npu_inst_pe_1_5_7_n10), .Q(
        npu_inst_pe_1_5_7_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_5_7_n86), 
        .CK(npu_inst_pe_1_5_7_net3218), .RN(npu_inst_pe_1_5_7_n10), .Q(
        npu_inst_pe_1_5_7_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_5_7_n87), 
        .CK(npu_inst_pe_1_5_7_net3218), .RN(npu_inst_pe_1_5_7_n10), .Q(
        npu_inst_pe_1_5_7_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_5_7_n88), 
        .CK(npu_inst_pe_1_5_7_net3218), .RN(npu_inst_pe_1_5_7_n11), .Q(
        npu_inst_pe_1_5_7_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_5_7_n89), 
        .CK(npu_inst_pe_1_5_7_net3218), .RN(npu_inst_pe_1_5_7_n11), .Q(
        npu_inst_pe_1_5_7_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_5_7_n90), 
        .CK(npu_inst_pe_1_5_7_net3218), .RN(npu_inst_pe_1_5_7_n11), .Q(
        npu_inst_pe_1_5_7_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_5_7_n91), 
        .CK(npu_inst_pe_1_5_7_net3218), .RN(npu_inst_pe_1_5_7_n11), .Q(
        npu_inst_pe_1_5_7_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_5_7_n92), 
        .CK(npu_inst_pe_1_5_7_net3218), .RN(npu_inst_pe_1_5_7_n11), .Q(
        npu_inst_pe_1_5_7_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_5_7_n93), 
        .CK(npu_inst_pe_1_5_7_net3218), .RN(npu_inst_pe_1_5_7_n11), .Q(
        npu_inst_pe_1_5_7_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_5_7_n94), 
        .CK(npu_inst_pe_1_5_7_net3218), .RN(npu_inst_pe_1_5_7_n11), .Q(
        npu_inst_pe_1_5_7_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_5_7_n95), 
        .CK(npu_inst_pe_1_5_7_net3218), .RN(npu_inst_pe_1_5_7_n11), .Q(
        npu_inst_pe_1_5_7_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_5_7_n96), 
        .CK(npu_inst_pe_1_5_7_net3218), .RN(npu_inst_pe_1_5_7_n11), .Q(
        npu_inst_pe_1_5_7_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_5_7_n97), 
        .CK(npu_inst_pe_1_5_7_net3218), .RN(npu_inst_pe_1_5_7_n11), .Q(
        npu_inst_pe_1_5_7_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_5_7_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_5_7_N84), .SE(1'b0), .GCK(npu_inst_pe_1_5_7_net3212) );
  CLKGATETST_X1 npu_inst_pe_1_5_7_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n62), .SE(1'b0), .GCK(npu_inst_pe_1_5_7_net3218) );
  MUX2_X1 npu_inst_pe_1_6_0_U162 ( .A(npu_inst_pe_1_6_0_n32), .B(
        npu_inst_pe_1_6_0_n29), .S(npu_inst_pe_1_6_0_n8), .Z(
        npu_inst_pe_1_6_0_N93) );
  MUX2_X1 npu_inst_pe_1_6_0_U161 ( .A(npu_inst_pe_1_6_0_n31), .B(
        npu_inst_pe_1_6_0_n30), .S(npu_inst_pe_1_6_0_n6), .Z(
        npu_inst_pe_1_6_0_n32) );
  MUX2_X1 npu_inst_pe_1_6_0_U160 ( .A(npu_inst_pe_1_6_0_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_6_0_int_q_reg_v_1__0_), .S(npu_inst_pe_1_6_0_n4), .Z(
        npu_inst_pe_1_6_0_n31) );
  MUX2_X1 npu_inst_pe_1_6_0_U159 ( .A(npu_inst_pe_1_6_0_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_6_0_int_q_reg_v_3__0_), .S(npu_inst_pe_1_6_0_n4), .Z(
        npu_inst_pe_1_6_0_n30) );
  MUX2_X1 npu_inst_pe_1_6_0_U158 ( .A(npu_inst_pe_1_6_0_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_6_0_int_q_reg_v_5__0_), .S(npu_inst_pe_1_6_0_n4), .Z(
        npu_inst_pe_1_6_0_n29) );
  MUX2_X1 npu_inst_pe_1_6_0_U157 ( .A(npu_inst_pe_1_6_0_n28), .B(
        npu_inst_pe_1_6_0_n23), .S(npu_inst_pe_1_6_0_n8), .Z(
        npu_inst_pe_1_6_0_N94) );
  MUX2_X1 npu_inst_pe_1_6_0_U156 ( .A(npu_inst_pe_1_6_0_n25), .B(
        npu_inst_pe_1_6_0_n24), .S(npu_inst_pe_1_6_0_n6), .Z(
        npu_inst_pe_1_6_0_n28) );
  MUX2_X1 npu_inst_pe_1_6_0_U155 ( .A(npu_inst_pe_1_6_0_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_6_0_int_q_reg_v_1__1_), .S(npu_inst_pe_1_6_0_n4), .Z(
        npu_inst_pe_1_6_0_n25) );
  MUX2_X1 npu_inst_pe_1_6_0_U154 ( .A(npu_inst_pe_1_6_0_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_6_0_int_q_reg_v_3__1_), .S(npu_inst_pe_1_6_0_n4), .Z(
        npu_inst_pe_1_6_0_n24) );
  MUX2_X1 npu_inst_pe_1_6_0_U153 ( .A(npu_inst_pe_1_6_0_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_6_0_int_q_reg_v_5__1_), .S(npu_inst_pe_1_6_0_n4), .Z(
        npu_inst_pe_1_6_0_n23) );
  MUX2_X1 npu_inst_pe_1_6_0_U152 ( .A(npu_inst_pe_1_6_0_n22), .B(
        npu_inst_pe_1_6_0_n19), .S(npu_inst_pe_1_6_0_n8), .Z(
        npu_inst_pe_1_6_0_o_data_h_1_) );
  MUX2_X1 npu_inst_pe_1_6_0_U151 ( .A(npu_inst_pe_1_6_0_n21), .B(
        npu_inst_pe_1_6_0_n20), .S(npu_inst_pe_1_6_0_n6), .Z(
        npu_inst_pe_1_6_0_n22) );
  MUX2_X1 npu_inst_pe_1_6_0_U150 ( .A(npu_inst_pe_1_6_0_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_6_0_int_q_reg_h_1__1_), .S(npu_inst_pe_1_6_0_n4), .Z(
        npu_inst_pe_1_6_0_n21) );
  MUX2_X1 npu_inst_pe_1_6_0_U149 ( .A(npu_inst_pe_1_6_0_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_6_0_int_q_reg_h_3__1_), .S(npu_inst_pe_1_6_0_n4), .Z(
        npu_inst_pe_1_6_0_n20) );
  MUX2_X1 npu_inst_pe_1_6_0_U148 ( .A(npu_inst_pe_1_6_0_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_6_0_int_q_reg_h_5__1_), .S(npu_inst_pe_1_6_0_n4), .Z(
        npu_inst_pe_1_6_0_n19) );
  MUX2_X1 npu_inst_pe_1_6_0_U147 ( .A(npu_inst_pe_1_6_0_n18), .B(
        npu_inst_pe_1_6_0_n15), .S(npu_inst_pe_1_6_0_n8), .Z(
        npu_inst_pe_1_6_0_o_data_h_0_) );
  MUX2_X1 npu_inst_pe_1_6_0_U146 ( .A(npu_inst_pe_1_6_0_n17), .B(
        npu_inst_pe_1_6_0_n16), .S(npu_inst_pe_1_6_0_n6), .Z(
        npu_inst_pe_1_6_0_n18) );
  MUX2_X1 npu_inst_pe_1_6_0_U145 ( .A(npu_inst_pe_1_6_0_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_6_0_int_q_reg_h_1__0_), .S(npu_inst_pe_1_6_0_n4), .Z(
        npu_inst_pe_1_6_0_n17) );
  MUX2_X1 npu_inst_pe_1_6_0_U144 ( .A(npu_inst_pe_1_6_0_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_6_0_int_q_reg_h_3__0_), .S(npu_inst_pe_1_6_0_n4), .Z(
        npu_inst_pe_1_6_0_n16) );
  MUX2_X1 npu_inst_pe_1_6_0_U143 ( .A(npu_inst_pe_1_6_0_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_6_0_int_q_reg_h_5__0_), .S(npu_inst_pe_1_6_0_n4), .Z(
        npu_inst_pe_1_6_0_n15) );
  XOR2_X1 npu_inst_pe_1_6_0_U142 ( .A(npu_inst_pe_1_6_0_int_data_0_), .B(
        npu_inst_pe_1_6_0_int_q_acc_0_), .Z(npu_inst_pe_1_6_0_N73) );
  AND2_X1 npu_inst_pe_1_6_0_U141 ( .A1(npu_inst_pe_1_6_0_int_q_acc_0_), .A2(
        npu_inst_pe_1_6_0_int_data_0_), .ZN(npu_inst_pe_1_6_0_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_6_0_U140 ( .A(npu_inst_pe_1_6_0_int_q_acc_0_), .B(
        npu_inst_pe_1_6_0_n13), .ZN(npu_inst_pe_1_6_0_N65) );
  OR2_X1 npu_inst_pe_1_6_0_U139 ( .A1(npu_inst_pe_1_6_0_n13), .A2(
        npu_inst_pe_1_6_0_int_q_acc_0_), .ZN(npu_inst_pe_1_6_0_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_6_0_U138 ( .A(npu_inst_pe_1_6_0_int_q_acc_2_), .B(
        npu_inst_pe_1_6_0_add_79_carry_2_), .Z(npu_inst_pe_1_6_0_N75) );
  AND2_X1 npu_inst_pe_1_6_0_U137 ( .A1(npu_inst_pe_1_6_0_add_79_carry_2_), 
        .A2(npu_inst_pe_1_6_0_int_q_acc_2_), .ZN(
        npu_inst_pe_1_6_0_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_6_0_U136 ( .A(npu_inst_pe_1_6_0_int_q_acc_3_), .B(
        npu_inst_pe_1_6_0_add_79_carry_3_), .Z(npu_inst_pe_1_6_0_N76) );
  AND2_X1 npu_inst_pe_1_6_0_U135 ( .A1(npu_inst_pe_1_6_0_add_79_carry_3_), 
        .A2(npu_inst_pe_1_6_0_int_q_acc_3_), .ZN(
        npu_inst_pe_1_6_0_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_6_0_U134 ( .A(npu_inst_pe_1_6_0_int_q_acc_4_), .B(
        npu_inst_pe_1_6_0_add_79_carry_4_), .Z(npu_inst_pe_1_6_0_N77) );
  AND2_X1 npu_inst_pe_1_6_0_U133 ( .A1(npu_inst_pe_1_6_0_add_79_carry_4_), 
        .A2(npu_inst_pe_1_6_0_int_q_acc_4_), .ZN(
        npu_inst_pe_1_6_0_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_6_0_U132 ( .A(npu_inst_pe_1_6_0_int_q_acc_5_), .B(
        npu_inst_pe_1_6_0_add_79_carry_5_), .Z(npu_inst_pe_1_6_0_N78) );
  AND2_X1 npu_inst_pe_1_6_0_U131 ( .A1(npu_inst_pe_1_6_0_add_79_carry_5_), 
        .A2(npu_inst_pe_1_6_0_int_q_acc_5_), .ZN(
        npu_inst_pe_1_6_0_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_6_0_U130 ( .A(npu_inst_pe_1_6_0_int_q_acc_6_), .B(
        npu_inst_pe_1_6_0_add_79_carry_6_), .Z(npu_inst_pe_1_6_0_N79) );
  AND2_X1 npu_inst_pe_1_6_0_U129 ( .A1(npu_inst_pe_1_6_0_add_79_carry_6_), 
        .A2(npu_inst_pe_1_6_0_int_q_acc_6_), .ZN(
        npu_inst_pe_1_6_0_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_6_0_U128 ( .A(npu_inst_pe_1_6_0_int_q_acc_7_), .B(
        npu_inst_pe_1_6_0_add_79_carry_7_), .Z(npu_inst_pe_1_6_0_N80) );
  XNOR2_X1 npu_inst_pe_1_6_0_U127 ( .A(npu_inst_pe_1_6_0_sub_77_carry_2_), .B(
        npu_inst_pe_1_6_0_int_q_acc_2_), .ZN(npu_inst_pe_1_6_0_N67) );
  OR2_X1 npu_inst_pe_1_6_0_U126 ( .A1(npu_inst_pe_1_6_0_int_q_acc_2_), .A2(
        npu_inst_pe_1_6_0_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_6_0_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_6_0_U125 ( .A(npu_inst_pe_1_6_0_sub_77_carry_3_), .B(
        npu_inst_pe_1_6_0_int_q_acc_3_), .ZN(npu_inst_pe_1_6_0_N68) );
  OR2_X1 npu_inst_pe_1_6_0_U124 ( .A1(npu_inst_pe_1_6_0_int_q_acc_3_), .A2(
        npu_inst_pe_1_6_0_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_6_0_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_6_0_U123 ( .A(npu_inst_pe_1_6_0_sub_77_carry_4_), .B(
        npu_inst_pe_1_6_0_int_q_acc_4_), .ZN(npu_inst_pe_1_6_0_N69) );
  OR2_X1 npu_inst_pe_1_6_0_U122 ( .A1(npu_inst_pe_1_6_0_int_q_acc_4_), .A2(
        npu_inst_pe_1_6_0_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_6_0_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_6_0_U121 ( .A(npu_inst_pe_1_6_0_sub_77_carry_5_), .B(
        npu_inst_pe_1_6_0_int_q_acc_5_), .ZN(npu_inst_pe_1_6_0_N70) );
  OR2_X1 npu_inst_pe_1_6_0_U120 ( .A1(npu_inst_pe_1_6_0_int_q_acc_5_), .A2(
        npu_inst_pe_1_6_0_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_6_0_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_6_0_U119 ( .A(npu_inst_pe_1_6_0_sub_77_carry_6_), .B(
        npu_inst_pe_1_6_0_int_q_acc_6_), .ZN(npu_inst_pe_1_6_0_N71) );
  OR2_X1 npu_inst_pe_1_6_0_U118 ( .A1(npu_inst_pe_1_6_0_int_q_acc_6_), .A2(
        npu_inst_pe_1_6_0_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_6_0_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_6_0_U117 ( .A(npu_inst_pe_1_6_0_int_q_acc_7_), .B(
        npu_inst_pe_1_6_0_sub_77_carry_7_), .ZN(npu_inst_pe_1_6_0_N72) );
  INV_X1 npu_inst_pe_1_6_0_U116 ( .A(npu_inst_n76), .ZN(npu_inst_pe_1_6_0_n7)
         );
  INV_X1 npu_inst_pe_1_6_0_U115 ( .A(npu_inst_pe_1_6_0_n7), .ZN(
        npu_inst_pe_1_6_0_n6) );
  INV_X1 npu_inst_pe_1_6_0_U114 ( .A(npu_inst_n54), .ZN(npu_inst_pe_1_6_0_n3)
         );
  AOI22_X1 npu_inst_pe_1_6_0_U113 ( .A1(npu_inst_int_data_y_7__0__0_), .A2(
        npu_inst_pe_1_6_0_n58), .B1(npu_inst_pe_1_6_0_n114), .B2(
        npu_inst_pe_1_6_0_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_6_0_n57) );
  INV_X1 npu_inst_pe_1_6_0_U112 ( .A(npu_inst_pe_1_6_0_n57), .ZN(
        npu_inst_pe_1_6_0_n108) );
  AOI22_X1 npu_inst_pe_1_6_0_U111 ( .A1(npu_inst_int_data_y_7__0__0_), .A2(
        npu_inst_pe_1_6_0_n54), .B1(npu_inst_pe_1_6_0_n115), .B2(
        npu_inst_pe_1_6_0_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_6_0_n53) );
  INV_X1 npu_inst_pe_1_6_0_U110 ( .A(npu_inst_pe_1_6_0_n53), .ZN(
        npu_inst_pe_1_6_0_n109) );
  AOI22_X1 npu_inst_pe_1_6_0_U107 ( .A1(npu_inst_int_data_y_7__0__0_), .A2(
        npu_inst_pe_1_6_0_n50), .B1(npu_inst_pe_1_6_0_n116), .B2(
        npu_inst_pe_1_6_0_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_6_0_n49) );
  INV_X1 npu_inst_pe_1_6_0_U106 ( .A(npu_inst_pe_1_6_0_n49), .ZN(
        npu_inst_pe_1_6_0_n110) );
  AOI22_X1 npu_inst_pe_1_6_0_U105 ( .A1(npu_inst_int_data_y_7__0__0_), .A2(
        npu_inst_pe_1_6_0_n46), .B1(npu_inst_pe_1_6_0_n117), .B2(
        npu_inst_pe_1_6_0_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_6_0_n45) );
  INV_X1 npu_inst_pe_1_6_0_U104 ( .A(npu_inst_pe_1_6_0_n45), .ZN(
        npu_inst_pe_1_6_0_n111) );
  AOI22_X1 npu_inst_pe_1_6_0_U103 ( .A1(npu_inst_int_data_y_7__0__0_), .A2(
        npu_inst_pe_1_6_0_n42), .B1(npu_inst_pe_1_6_0_n119), .B2(
        npu_inst_pe_1_6_0_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_6_0_n41) );
  INV_X1 npu_inst_pe_1_6_0_U102 ( .A(npu_inst_pe_1_6_0_n41), .ZN(
        npu_inst_pe_1_6_0_n112) );
  AOI22_X1 npu_inst_pe_1_6_0_U101 ( .A1(npu_inst_int_data_y_7__0__1_), .A2(
        npu_inst_pe_1_6_0_n58), .B1(npu_inst_pe_1_6_0_n114), .B2(
        npu_inst_pe_1_6_0_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_6_0_n59) );
  INV_X1 npu_inst_pe_1_6_0_U100 ( .A(npu_inst_pe_1_6_0_n59), .ZN(
        npu_inst_pe_1_6_0_n102) );
  AOI22_X1 npu_inst_pe_1_6_0_U99 ( .A1(npu_inst_int_data_y_7__0__1_), .A2(
        npu_inst_pe_1_6_0_n54), .B1(npu_inst_pe_1_6_0_n115), .B2(
        npu_inst_pe_1_6_0_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_6_0_n55) );
  INV_X1 npu_inst_pe_1_6_0_U98 ( .A(npu_inst_pe_1_6_0_n55), .ZN(
        npu_inst_pe_1_6_0_n103) );
  AOI22_X1 npu_inst_pe_1_6_0_U97 ( .A1(npu_inst_int_data_y_7__0__1_), .A2(
        npu_inst_pe_1_6_0_n50), .B1(npu_inst_pe_1_6_0_n116), .B2(
        npu_inst_pe_1_6_0_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_6_0_n51) );
  INV_X1 npu_inst_pe_1_6_0_U96 ( .A(npu_inst_pe_1_6_0_n51), .ZN(
        npu_inst_pe_1_6_0_n104) );
  AOI22_X1 npu_inst_pe_1_6_0_U95 ( .A1(npu_inst_int_data_y_7__0__1_), .A2(
        npu_inst_pe_1_6_0_n46), .B1(npu_inst_pe_1_6_0_n117), .B2(
        npu_inst_pe_1_6_0_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_6_0_n47) );
  INV_X1 npu_inst_pe_1_6_0_U94 ( .A(npu_inst_pe_1_6_0_n47), .ZN(
        npu_inst_pe_1_6_0_n105) );
  AOI22_X1 npu_inst_pe_1_6_0_U93 ( .A1(npu_inst_int_data_y_7__0__1_), .A2(
        npu_inst_pe_1_6_0_n42), .B1(npu_inst_pe_1_6_0_n119), .B2(
        npu_inst_pe_1_6_0_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_6_0_n43) );
  INV_X1 npu_inst_pe_1_6_0_U92 ( .A(npu_inst_pe_1_6_0_n43), .ZN(
        npu_inst_pe_1_6_0_n106) );
  AOI22_X1 npu_inst_pe_1_6_0_U91 ( .A1(npu_inst_pe_1_6_0_n38), .A2(
        npu_inst_int_data_y_7__0__1_), .B1(npu_inst_pe_1_6_0_n118), .B2(
        npu_inst_pe_1_6_0_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_6_0_n39) );
  INV_X1 npu_inst_pe_1_6_0_U90 ( .A(npu_inst_pe_1_6_0_n39), .ZN(
        npu_inst_pe_1_6_0_n107) );
  AOI22_X1 npu_inst_pe_1_6_0_U89 ( .A1(npu_inst_pe_1_6_0_n38), .A2(
        npu_inst_int_data_y_7__0__0_), .B1(npu_inst_pe_1_6_0_n118), .B2(
        npu_inst_pe_1_6_0_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_6_0_n37) );
  INV_X1 npu_inst_pe_1_6_0_U88 ( .A(npu_inst_pe_1_6_0_n37), .ZN(
        npu_inst_pe_1_6_0_n113) );
  NAND2_X1 npu_inst_pe_1_6_0_U87 ( .A1(npu_inst_pe_1_6_0_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_6_0_n60), .ZN(npu_inst_pe_1_6_0_n74) );
  OAI21_X1 npu_inst_pe_1_6_0_U86 ( .B1(npu_inst_pe_1_6_0_n63), .B2(
        npu_inst_pe_1_6_0_n60), .A(npu_inst_pe_1_6_0_n74), .ZN(
        npu_inst_pe_1_6_0_n97) );
  NAND2_X1 npu_inst_pe_1_6_0_U85 ( .A1(npu_inst_pe_1_6_0_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_6_0_n60), .ZN(npu_inst_pe_1_6_0_n73) );
  OAI21_X1 npu_inst_pe_1_6_0_U84 ( .B1(npu_inst_pe_1_6_0_n61), .B2(
        npu_inst_pe_1_6_0_n60), .A(npu_inst_pe_1_6_0_n73), .ZN(
        npu_inst_pe_1_6_0_n96) );
  NAND2_X1 npu_inst_pe_1_6_0_U83 ( .A1(npu_inst_pe_1_6_0_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_6_0_n56), .ZN(npu_inst_pe_1_6_0_n72) );
  OAI21_X1 npu_inst_pe_1_6_0_U82 ( .B1(npu_inst_pe_1_6_0_n63), .B2(
        npu_inst_pe_1_6_0_n56), .A(npu_inst_pe_1_6_0_n72), .ZN(
        npu_inst_pe_1_6_0_n95) );
  NAND2_X1 npu_inst_pe_1_6_0_U81 ( .A1(npu_inst_pe_1_6_0_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_6_0_n56), .ZN(npu_inst_pe_1_6_0_n71) );
  OAI21_X1 npu_inst_pe_1_6_0_U80 ( .B1(npu_inst_pe_1_6_0_n61), .B2(
        npu_inst_pe_1_6_0_n56), .A(npu_inst_pe_1_6_0_n71), .ZN(
        npu_inst_pe_1_6_0_n94) );
  NAND2_X1 npu_inst_pe_1_6_0_U79 ( .A1(npu_inst_pe_1_6_0_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_6_0_n52), .ZN(npu_inst_pe_1_6_0_n70) );
  OAI21_X1 npu_inst_pe_1_6_0_U78 ( .B1(npu_inst_pe_1_6_0_n63), .B2(
        npu_inst_pe_1_6_0_n52), .A(npu_inst_pe_1_6_0_n70), .ZN(
        npu_inst_pe_1_6_0_n93) );
  NAND2_X1 npu_inst_pe_1_6_0_U77 ( .A1(npu_inst_pe_1_6_0_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_6_0_n52), .ZN(npu_inst_pe_1_6_0_n69) );
  OAI21_X1 npu_inst_pe_1_6_0_U76 ( .B1(npu_inst_pe_1_6_0_n61), .B2(
        npu_inst_pe_1_6_0_n52), .A(npu_inst_pe_1_6_0_n69), .ZN(
        npu_inst_pe_1_6_0_n92) );
  NAND2_X1 npu_inst_pe_1_6_0_U75 ( .A1(npu_inst_pe_1_6_0_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_6_0_n48), .ZN(npu_inst_pe_1_6_0_n68) );
  OAI21_X1 npu_inst_pe_1_6_0_U74 ( .B1(npu_inst_pe_1_6_0_n63), .B2(
        npu_inst_pe_1_6_0_n48), .A(npu_inst_pe_1_6_0_n68), .ZN(
        npu_inst_pe_1_6_0_n91) );
  NAND2_X1 npu_inst_pe_1_6_0_U73 ( .A1(npu_inst_pe_1_6_0_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_6_0_n48), .ZN(npu_inst_pe_1_6_0_n67) );
  OAI21_X1 npu_inst_pe_1_6_0_U72 ( .B1(npu_inst_pe_1_6_0_n61), .B2(
        npu_inst_pe_1_6_0_n48), .A(npu_inst_pe_1_6_0_n67), .ZN(
        npu_inst_pe_1_6_0_n90) );
  NAND2_X1 npu_inst_pe_1_6_0_U71 ( .A1(npu_inst_pe_1_6_0_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_6_0_n44), .ZN(npu_inst_pe_1_6_0_n66) );
  OAI21_X1 npu_inst_pe_1_6_0_U70 ( .B1(npu_inst_pe_1_6_0_n63), .B2(
        npu_inst_pe_1_6_0_n44), .A(npu_inst_pe_1_6_0_n66), .ZN(
        npu_inst_pe_1_6_0_n89) );
  NAND2_X1 npu_inst_pe_1_6_0_U69 ( .A1(npu_inst_pe_1_6_0_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_6_0_n44), .ZN(npu_inst_pe_1_6_0_n65) );
  OAI21_X1 npu_inst_pe_1_6_0_U68 ( .B1(npu_inst_pe_1_6_0_n61), .B2(
        npu_inst_pe_1_6_0_n44), .A(npu_inst_pe_1_6_0_n65), .ZN(
        npu_inst_pe_1_6_0_n88) );
  NAND2_X1 npu_inst_pe_1_6_0_U67 ( .A1(npu_inst_pe_1_6_0_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_6_0_n40), .ZN(npu_inst_pe_1_6_0_n64) );
  OAI21_X1 npu_inst_pe_1_6_0_U66 ( .B1(npu_inst_pe_1_6_0_n63), .B2(
        npu_inst_pe_1_6_0_n40), .A(npu_inst_pe_1_6_0_n64), .ZN(
        npu_inst_pe_1_6_0_n87) );
  NAND2_X1 npu_inst_pe_1_6_0_U65 ( .A1(npu_inst_pe_1_6_0_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_6_0_n40), .ZN(npu_inst_pe_1_6_0_n62) );
  OAI21_X1 npu_inst_pe_1_6_0_U64 ( .B1(npu_inst_pe_1_6_0_n61), .B2(
        npu_inst_pe_1_6_0_n40), .A(npu_inst_pe_1_6_0_n62), .ZN(
        npu_inst_pe_1_6_0_n86) );
  AND2_X1 npu_inst_pe_1_6_0_U63 ( .A1(npu_inst_pe_1_6_0_N93), .A2(npu_inst_n54), .ZN(npu_inst_int_data_y_6__0__0_) );
  AND2_X1 npu_inst_pe_1_6_0_U62 ( .A1(npu_inst_n54), .A2(npu_inst_pe_1_6_0_N94), .ZN(npu_inst_int_data_y_6__0__1_) );
  NOR3_X1 npu_inst_pe_1_6_0_U61 ( .A1(npu_inst_pe_1_6_0_n26), .A2(npu_inst_n54), .A3(npu_inst_int_ckg[15]), .ZN(npu_inst_pe_1_6_0_n85) );
  OR2_X1 npu_inst_pe_1_6_0_U60 ( .A1(npu_inst_pe_1_6_0_n85), .A2(
        npu_inst_pe_1_6_0_n2), .ZN(npu_inst_pe_1_6_0_N84) );
  AND2_X1 npu_inst_pe_1_6_0_U59 ( .A1(npu_inst_pe_1_6_0_int_q_acc_0_), .A2(
        npu_inst_pe_1_6_0_n1), .ZN(npu_inst_int_data_res_6__0__0_) );
  AND2_X1 npu_inst_pe_1_6_0_U58 ( .A1(npu_inst_pe_1_6_0_n2), .A2(
        npu_inst_pe_1_6_0_int_q_acc_7_), .ZN(npu_inst_int_data_res_6__0__7_)
         );
  AND2_X1 npu_inst_pe_1_6_0_U57 ( .A1(npu_inst_pe_1_6_0_int_q_acc_1_), .A2(
        npu_inst_pe_1_6_0_n1), .ZN(npu_inst_int_data_res_6__0__1_) );
  AND2_X1 npu_inst_pe_1_6_0_U56 ( .A1(npu_inst_pe_1_6_0_int_q_acc_2_), .A2(
        npu_inst_pe_1_6_0_n1), .ZN(npu_inst_int_data_res_6__0__2_) );
  AND2_X1 npu_inst_pe_1_6_0_U55 ( .A1(npu_inst_pe_1_6_0_int_q_acc_3_), .A2(
        npu_inst_pe_1_6_0_n2), .ZN(npu_inst_int_data_res_6__0__3_) );
  AND2_X1 npu_inst_pe_1_6_0_U54 ( .A1(npu_inst_pe_1_6_0_int_q_acc_4_), .A2(
        npu_inst_pe_1_6_0_n2), .ZN(npu_inst_int_data_res_6__0__4_) );
  AND2_X1 npu_inst_pe_1_6_0_U53 ( .A1(npu_inst_pe_1_6_0_int_q_acc_5_), .A2(
        npu_inst_pe_1_6_0_n2), .ZN(npu_inst_int_data_res_6__0__5_) );
  AND2_X1 npu_inst_pe_1_6_0_U52 ( .A1(npu_inst_pe_1_6_0_int_q_acc_6_), .A2(
        npu_inst_pe_1_6_0_n2), .ZN(npu_inst_int_data_res_6__0__6_) );
  AOI222_X1 npu_inst_pe_1_6_0_U51 ( .A1(npu_inst_int_data_res_7__0__0_), .A2(
        npu_inst_pe_1_6_0_n1), .B1(npu_inst_pe_1_6_0_N73), .B2(
        npu_inst_pe_1_6_0_n76), .C1(npu_inst_pe_1_6_0_N65), .C2(
        npu_inst_pe_1_6_0_n77), .ZN(npu_inst_pe_1_6_0_n84) );
  INV_X1 npu_inst_pe_1_6_0_U50 ( .A(npu_inst_pe_1_6_0_n84), .ZN(
        npu_inst_pe_1_6_0_n101) );
  AOI222_X1 npu_inst_pe_1_6_0_U49 ( .A1(npu_inst_int_data_res_7__0__7_), .A2(
        npu_inst_pe_1_6_0_n1), .B1(npu_inst_pe_1_6_0_N80), .B2(
        npu_inst_pe_1_6_0_n76), .C1(npu_inst_pe_1_6_0_N72), .C2(
        npu_inst_pe_1_6_0_n77), .ZN(npu_inst_pe_1_6_0_n75) );
  INV_X1 npu_inst_pe_1_6_0_U48 ( .A(npu_inst_pe_1_6_0_n75), .ZN(
        npu_inst_pe_1_6_0_n33) );
  AOI222_X1 npu_inst_pe_1_6_0_U47 ( .A1(npu_inst_int_data_res_7__0__1_), .A2(
        npu_inst_pe_1_6_0_n1), .B1(npu_inst_pe_1_6_0_N74), .B2(
        npu_inst_pe_1_6_0_n76), .C1(npu_inst_pe_1_6_0_N66), .C2(
        npu_inst_pe_1_6_0_n77), .ZN(npu_inst_pe_1_6_0_n83) );
  INV_X1 npu_inst_pe_1_6_0_U46 ( .A(npu_inst_pe_1_6_0_n83), .ZN(
        npu_inst_pe_1_6_0_n100) );
  AOI222_X1 npu_inst_pe_1_6_0_U45 ( .A1(npu_inst_int_data_res_7__0__2_), .A2(
        npu_inst_pe_1_6_0_n1), .B1(npu_inst_pe_1_6_0_N75), .B2(
        npu_inst_pe_1_6_0_n76), .C1(npu_inst_pe_1_6_0_N67), .C2(
        npu_inst_pe_1_6_0_n77), .ZN(npu_inst_pe_1_6_0_n82) );
  INV_X1 npu_inst_pe_1_6_0_U44 ( .A(npu_inst_pe_1_6_0_n82), .ZN(
        npu_inst_pe_1_6_0_n99) );
  AOI222_X1 npu_inst_pe_1_6_0_U43 ( .A1(npu_inst_int_data_res_7__0__3_), .A2(
        npu_inst_pe_1_6_0_n1), .B1(npu_inst_pe_1_6_0_N76), .B2(
        npu_inst_pe_1_6_0_n76), .C1(npu_inst_pe_1_6_0_N68), .C2(
        npu_inst_pe_1_6_0_n77), .ZN(npu_inst_pe_1_6_0_n81) );
  INV_X1 npu_inst_pe_1_6_0_U42 ( .A(npu_inst_pe_1_6_0_n81), .ZN(
        npu_inst_pe_1_6_0_n98) );
  AOI222_X1 npu_inst_pe_1_6_0_U41 ( .A1(npu_inst_int_data_res_7__0__4_), .A2(
        npu_inst_pe_1_6_0_n1), .B1(npu_inst_pe_1_6_0_N77), .B2(
        npu_inst_pe_1_6_0_n76), .C1(npu_inst_pe_1_6_0_N69), .C2(
        npu_inst_pe_1_6_0_n77), .ZN(npu_inst_pe_1_6_0_n80) );
  INV_X1 npu_inst_pe_1_6_0_U40 ( .A(npu_inst_pe_1_6_0_n80), .ZN(
        npu_inst_pe_1_6_0_n36) );
  AOI222_X1 npu_inst_pe_1_6_0_U39 ( .A1(npu_inst_int_data_res_7__0__5_), .A2(
        npu_inst_pe_1_6_0_n1), .B1(npu_inst_pe_1_6_0_N78), .B2(
        npu_inst_pe_1_6_0_n76), .C1(npu_inst_pe_1_6_0_N70), .C2(
        npu_inst_pe_1_6_0_n77), .ZN(npu_inst_pe_1_6_0_n79) );
  INV_X1 npu_inst_pe_1_6_0_U38 ( .A(npu_inst_pe_1_6_0_n79), .ZN(
        npu_inst_pe_1_6_0_n35) );
  AOI222_X1 npu_inst_pe_1_6_0_U37 ( .A1(npu_inst_int_data_res_7__0__6_), .A2(
        npu_inst_pe_1_6_0_n1), .B1(npu_inst_pe_1_6_0_N79), .B2(
        npu_inst_pe_1_6_0_n76), .C1(npu_inst_pe_1_6_0_N71), .C2(
        npu_inst_pe_1_6_0_n77), .ZN(npu_inst_pe_1_6_0_n78) );
  INV_X1 npu_inst_pe_1_6_0_U36 ( .A(npu_inst_pe_1_6_0_n78), .ZN(
        npu_inst_pe_1_6_0_n34) );
  AND2_X1 npu_inst_pe_1_6_0_U35 ( .A1(npu_inst_pe_1_6_0_o_data_h_1_), .A2(
        npu_inst_pe_1_6_0_int_q_weight_1_), .ZN(npu_inst_pe_1_6_0_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_6_0_U34 ( .A1(npu_inst_pe_1_6_0_o_data_h_0_), .A2(
        npu_inst_pe_1_6_0_int_q_weight_1_), .ZN(npu_inst_pe_1_6_0_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_6_0_U33 ( .A(npu_inst_pe_1_6_0_int_data_1_), .ZN(
        npu_inst_pe_1_6_0_n14) );
  AOI22_X1 npu_inst_pe_1_6_0_U32 ( .A1(npu_inst_n54), .A2(
        npu_inst_int_data_y_7__0__1_), .B1(npu_inst_pe_1_6_0_n3), .B2(
        npu_inst_int_data_x_6__1__1_), .ZN(npu_inst_pe_1_6_0_n63) );
  AOI22_X1 npu_inst_pe_1_6_0_U31 ( .A1(npu_inst_n54), .A2(
        npu_inst_int_data_y_7__0__0_), .B1(npu_inst_pe_1_6_0_n3), .B2(
        npu_inst_int_data_x_6__1__0_), .ZN(npu_inst_pe_1_6_0_n61) );
  INV_X1 npu_inst_pe_1_6_0_U30 ( .A(npu_inst_pe_1_6_0_int_data_0_), .ZN(
        npu_inst_pe_1_6_0_n13) );
  INV_X1 npu_inst_pe_1_6_0_U29 ( .A(npu_inst_n68), .ZN(npu_inst_pe_1_6_0_n5)
         );
  OR3_X1 npu_inst_pe_1_6_0_U28 ( .A1(npu_inst_pe_1_6_0_n6), .A2(
        npu_inst_pe_1_6_0_n8), .A3(npu_inst_pe_1_6_0_n5), .ZN(
        npu_inst_pe_1_6_0_n56) );
  OR3_X1 npu_inst_pe_1_6_0_U27 ( .A1(npu_inst_pe_1_6_0_n5), .A2(
        npu_inst_pe_1_6_0_n8), .A3(npu_inst_pe_1_6_0_n7), .ZN(
        npu_inst_pe_1_6_0_n48) );
  INV_X1 npu_inst_pe_1_6_0_U26 ( .A(npu_inst_pe_1_6_0_n5), .ZN(
        npu_inst_pe_1_6_0_n4) );
  INV_X1 npu_inst_pe_1_6_0_U25 ( .A(npu_inst_n123), .ZN(npu_inst_pe_1_6_0_n12)
         );
  OR3_X1 npu_inst_pe_1_6_0_U24 ( .A1(npu_inst_pe_1_6_0_n4), .A2(
        npu_inst_pe_1_6_0_n8), .A3(npu_inst_pe_1_6_0_n7), .ZN(
        npu_inst_pe_1_6_0_n52) );
  OR3_X1 npu_inst_pe_1_6_0_U23 ( .A1(npu_inst_pe_1_6_0_n6), .A2(
        npu_inst_pe_1_6_0_n8), .A3(npu_inst_pe_1_6_0_n4), .ZN(
        npu_inst_pe_1_6_0_n60) );
  NOR2_X1 npu_inst_pe_1_6_0_U22 ( .A1(npu_inst_pe_1_6_0_n60), .A2(
        npu_inst_pe_1_6_0_n3), .ZN(npu_inst_pe_1_6_0_n58) );
  NOR2_X1 npu_inst_pe_1_6_0_U21 ( .A1(npu_inst_pe_1_6_0_n56), .A2(
        npu_inst_pe_1_6_0_n3), .ZN(npu_inst_pe_1_6_0_n54) );
  NOR2_X1 npu_inst_pe_1_6_0_U20 ( .A1(npu_inst_pe_1_6_0_n52), .A2(
        npu_inst_pe_1_6_0_n3), .ZN(npu_inst_pe_1_6_0_n50) );
  NOR2_X1 npu_inst_pe_1_6_0_U19 ( .A1(npu_inst_pe_1_6_0_n48), .A2(
        npu_inst_pe_1_6_0_n3), .ZN(npu_inst_pe_1_6_0_n46) );
  NOR2_X1 npu_inst_pe_1_6_0_U18 ( .A1(npu_inst_pe_1_6_0_n40), .A2(
        npu_inst_pe_1_6_0_n3), .ZN(npu_inst_pe_1_6_0_n38) );
  NOR2_X1 npu_inst_pe_1_6_0_U17 ( .A1(npu_inst_pe_1_6_0_n44), .A2(
        npu_inst_pe_1_6_0_n3), .ZN(npu_inst_pe_1_6_0_n42) );
  BUF_X1 npu_inst_pe_1_6_0_U16 ( .A(npu_inst_n95), .Z(npu_inst_pe_1_6_0_n8) );
  BUF_X1 npu_inst_pe_1_6_0_U15 ( .A(npu_inst_pe_1_6_0_n12), .Z(
        npu_inst_pe_1_6_0_n11) );
  BUF_X1 npu_inst_pe_1_6_0_U14 ( .A(npu_inst_pe_1_6_0_n12), .Z(
        npu_inst_pe_1_6_0_n10) );
  BUF_X1 npu_inst_pe_1_6_0_U13 ( .A(npu_inst_pe_1_6_0_n12), .Z(
        npu_inst_pe_1_6_0_n9) );
  INV_X1 npu_inst_pe_1_6_0_U12 ( .A(npu_inst_pe_1_6_0_n38), .ZN(
        npu_inst_pe_1_6_0_n118) );
  INV_X1 npu_inst_pe_1_6_0_U11 ( .A(npu_inst_pe_1_6_0_n58), .ZN(
        npu_inst_pe_1_6_0_n114) );
  INV_X1 npu_inst_pe_1_6_0_U10 ( .A(npu_inst_pe_1_6_0_n54), .ZN(
        npu_inst_pe_1_6_0_n115) );
  INV_X1 npu_inst_pe_1_6_0_U9 ( .A(npu_inst_pe_1_6_0_n50), .ZN(
        npu_inst_pe_1_6_0_n116) );
  INV_X1 npu_inst_pe_1_6_0_U8 ( .A(npu_inst_pe_1_6_0_n46), .ZN(
        npu_inst_pe_1_6_0_n117) );
  INV_X1 npu_inst_pe_1_6_0_U7 ( .A(npu_inst_pe_1_6_0_n42), .ZN(
        npu_inst_pe_1_6_0_n119) );
  BUF_X1 npu_inst_pe_1_6_0_U6 ( .A(npu_inst_n14), .Z(npu_inst_pe_1_6_0_n2) );
  BUF_X1 npu_inst_pe_1_6_0_U5 ( .A(npu_inst_n14), .Z(npu_inst_pe_1_6_0_n1) );
  NOR2_X1 npu_inst_pe_1_6_0_U4 ( .A1(npu_inst_pe_1_6_0_int_q_weight_0_), .A2(
        npu_inst_pe_1_6_0_n1), .ZN(npu_inst_pe_1_6_0_n76) );
  NOR2_X1 npu_inst_pe_1_6_0_U3 ( .A1(npu_inst_pe_1_6_0_n27), .A2(
        npu_inst_pe_1_6_0_n1), .ZN(npu_inst_pe_1_6_0_n77) );
  FA_X1 npu_inst_pe_1_6_0_sub_77_U2_1 ( .A(npu_inst_pe_1_6_0_int_q_acc_1_), 
        .B(npu_inst_pe_1_6_0_n14), .CI(npu_inst_pe_1_6_0_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_6_0_sub_77_carry_2_), .S(npu_inst_pe_1_6_0_N66) );
  FA_X1 npu_inst_pe_1_6_0_add_79_U1_1 ( .A(npu_inst_pe_1_6_0_int_q_acc_1_), 
        .B(npu_inst_pe_1_6_0_int_data_1_), .CI(
        npu_inst_pe_1_6_0_add_79_carry_1_), .CO(
        npu_inst_pe_1_6_0_add_79_carry_2_), .S(npu_inst_pe_1_6_0_N74) );
  NAND3_X1 npu_inst_pe_1_6_0_U109 ( .A1(npu_inst_pe_1_6_0_n5), .A2(
        npu_inst_pe_1_6_0_n7), .A3(npu_inst_pe_1_6_0_n8), .ZN(
        npu_inst_pe_1_6_0_n44) );
  NAND3_X1 npu_inst_pe_1_6_0_U108 ( .A1(npu_inst_pe_1_6_0_n4), .A2(
        npu_inst_pe_1_6_0_n7), .A3(npu_inst_pe_1_6_0_n8), .ZN(
        npu_inst_pe_1_6_0_n40) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_6_0_n34), .CK(
        npu_inst_pe_1_6_0_net3189), .RN(npu_inst_pe_1_6_0_n9), .Q(
        npu_inst_pe_1_6_0_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_6_0_n35), .CK(
        npu_inst_pe_1_6_0_net3189), .RN(npu_inst_pe_1_6_0_n9), .Q(
        npu_inst_pe_1_6_0_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_6_0_n36), .CK(
        npu_inst_pe_1_6_0_net3189), .RN(npu_inst_pe_1_6_0_n9), .Q(
        npu_inst_pe_1_6_0_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_6_0_n98), .CK(
        npu_inst_pe_1_6_0_net3189), .RN(npu_inst_pe_1_6_0_n9), .Q(
        npu_inst_pe_1_6_0_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_6_0_n99), .CK(
        npu_inst_pe_1_6_0_net3189), .RN(npu_inst_pe_1_6_0_n9), .Q(
        npu_inst_pe_1_6_0_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_6_0_n100), 
        .CK(npu_inst_pe_1_6_0_net3189), .RN(npu_inst_pe_1_6_0_n9), .Q(
        npu_inst_pe_1_6_0_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_6_0_n33), .CK(
        npu_inst_pe_1_6_0_net3189), .RN(npu_inst_pe_1_6_0_n9), .Q(
        npu_inst_pe_1_6_0_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_6_0_n101), 
        .CK(npu_inst_pe_1_6_0_net3189), .RN(npu_inst_pe_1_6_0_n9), .Q(
        npu_inst_pe_1_6_0_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_weight_reg_0_ ( .D(npu_inst_n109), .CK(
        npu_inst_pe_1_6_0_net3195), .RN(npu_inst_pe_1_6_0_n9), .Q(
        npu_inst_pe_1_6_0_int_q_weight_0_), .QN(npu_inst_pe_1_6_0_n27) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_weight_reg_1_ ( .D(npu_inst_n115), .CK(
        npu_inst_pe_1_6_0_net3195), .RN(npu_inst_pe_1_6_0_n9), .Q(
        npu_inst_pe_1_6_0_int_q_weight_1_), .QN(npu_inst_pe_1_6_0_n26) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_6_0_n113), 
        .CK(npu_inst_pe_1_6_0_net3195), .RN(npu_inst_pe_1_6_0_n9), .Q(
        npu_inst_pe_1_6_0_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_6_0_n107), 
        .CK(npu_inst_pe_1_6_0_net3195), .RN(npu_inst_pe_1_6_0_n9), .Q(
        npu_inst_pe_1_6_0_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_6_0_n112), 
        .CK(npu_inst_pe_1_6_0_net3195), .RN(npu_inst_pe_1_6_0_n10), .Q(
        npu_inst_pe_1_6_0_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_6_0_n106), 
        .CK(npu_inst_pe_1_6_0_net3195), .RN(npu_inst_pe_1_6_0_n10), .Q(
        npu_inst_pe_1_6_0_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_6_0_n111), 
        .CK(npu_inst_pe_1_6_0_net3195), .RN(npu_inst_pe_1_6_0_n10), .Q(
        npu_inst_pe_1_6_0_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_6_0_n105), 
        .CK(npu_inst_pe_1_6_0_net3195), .RN(npu_inst_pe_1_6_0_n10), .Q(
        npu_inst_pe_1_6_0_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_6_0_n110), 
        .CK(npu_inst_pe_1_6_0_net3195), .RN(npu_inst_pe_1_6_0_n10), .Q(
        npu_inst_pe_1_6_0_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_6_0_n104), 
        .CK(npu_inst_pe_1_6_0_net3195), .RN(npu_inst_pe_1_6_0_n10), .Q(
        npu_inst_pe_1_6_0_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_6_0_n109), 
        .CK(npu_inst_pe_1_6_0_net3195), .RN(npu_inst_pe_1_6_0_n10), .Q(
        npu_inst_pe_1_6_0_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_6_0_n103), 
        .CK(npu_inst_pe_1_6_0_net3195), .RN(npu_inst_pe_1_6_0_n10), .Q(
        npu_inst_pe_1_6_0_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_6_0_n108), 
        .CK(npu_inst_pe_1_6_0_net3195), .RN(npu_inst_pe_1_6_0_n10), .Q(
        npu_inst_pe_1_6_0_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_6_0_n102), 
        .CK(npu_inst_pe_1_6_0_net3195), .RN(npu_inst_pe_1_6_0_n10), .Q(
        npu_inst_pe_1_6_0_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_6_0_n86), 
        .CK(npu_inst_pe_1_6_0_net3195), .RN(npu_inst_pe_1_6_0_n10), .Q(
        npu_inst_pe_1_6_0_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_6_0_n87), 
        .CK(npu_inst_pe_1_6_0_net3195), .RN(npu_inst_pe_1_6_0_n10), .Q(
        npu_inst_pe_1_6_0_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_6_0_n88), 
        .CK(npu_inst_pe_1_6_0_net3195), .RN(npu_inst_pe_1_6_0_n11), .Q(
        npu_inst_pe_1_6_0_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_6_0_n89), 
        .CK(npu_inst_pe_1_6_0_net3195), .RN(npu_inst_pe_1_6_0_n11), .Q(
        npu_inst_pe_1_6_0_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_6_0_n90), 
        .CK(npu_inst_pe_1_6_0_net3195), .RN(npu_inst_pe_1_6_0_n11), .Q(
        npu_inst_pe_1_6_0_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_6_0_n91), 
        .CK(npu_inst_pe_1_6_0_net3195), .RN(npu_inst_pe_1_6_0_n11), .Q(
        npu_inst_pe_1_6_0_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_6_0_n92), 
        .CK(npu_inst_pe_1_6_0_net3195), .RN(npu_inst_pe_1_6_0_n11), .Q(
        npu_inst_pe_1_6_0_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_6_0_n93), 
        .CK(npu_inst_pe_1_6_0_net3195), .RN(npu_inst_pe_1_6_0_n11), .Q(
        npu_inst_pe_1_6_0_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_6_0_n94), 
        .CK(npu_inst_pe_1_6_0_net3195), .RN(npu_inst_pe_1_6_0_n11), .Q(
        npu_inst_pe_1_6_0_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_6_0_n95), 
        .CK(npu_inst_pe_1_6_0_net3195), .RN(npu_inst_pe_1_6_0_n11), .Q(
        npu_inst_pe_1_6_0_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_6_0_n96), 
        .CK(npu_inst_pe_1_6_0_net3195), .RN(npu_inst_pe_1_6_0_n11), .Q(
        npu_inst_pe_1_6_0_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_6_0_n97), 
        .CK(npu_inst_pe_1_6_0_net3195), .RN(npu_inst_pe_1_6_0_n11), .Q(
        npu_inst_pe_1_6_0_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_6_0_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_6_0_N84), .SE(1'b0), .GCK(npu_inst_pe_1_6_0_net3189) );
  CLKGATETST_X1 npu_inst_pe_1_6_0_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n62), .SE(1'b0), .GCK(npu_inst_pe_1_6_0_net3195) );
  MUX2_X1 npu_inst_pe_1_6_1_U162 ( .A(npu_inst_pe_1_6_1_n32), .B(
        npu_inst_pe_1_6_1_n29), .S(npu_inst_pe_1_6_1_n8), .Z(
        npu_inst_pe_1_6_1_N93) );
  MUX2_X1 npu_inst_pe_1_6_1_U161 ( .A(npu_inst_pe_1_6_1_n31), .B(
        npu_inst_pe_1_6_1_n30), .S(npu_inst_pe_1_6_1_n6), .Z(
        npu_inst_pe_1_6_1_n32) );
  MUX2_X1 npu_inst_pe_1_6_1_U160 ( .A(npu_inst_pe_1_6_1_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_6_1_int_q_reg_v_1__0_), .S(npu_inst_pe_1_6_1_n4), .Z(
        npu_inst_pe_1_6_1_n31) );
  MUX2_X1 npu_inst_pe_1_6_1_U159 ( .A(npu_inst_pe_1_6_1_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_6_1_int_q_reg_v_3__0_), .S(npu_inst_pe_1_6_1_n4), .Z(
        npu_inst_pe_1_6_1_n30) );
  MUX2_X1 npu_inst_pe_1_6_1_U158 ( .A(npu_inst_pe_1_6_1_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_6_1_int_q_reg_v_5__0_), .S(npu_inst_pe_1_6_1_n4), .Z(
        npu_inst_pe_1_6_1_n29) );
  MUX2_X1 npu_inst_pe_1_6_1_U157 ( .A(npu_inst_pe_1_6_1_n28), .B(
        npu_inst_pe_1_6_1_n23), .S(npu_inst_pe_1_6_1_n8), .Z(
        npu_inst_pe_1_6_1_N94) );
  MUX2_X1 npu_inst_pe_1_6_1_U156 ( .A(npu_inst_pe_1_6_1_n25), .B(
        npu_inst_pe_1_6_1_n24), .S(npu_inst_pe_1_6_1_n6), .Z(
        npu_inst_pe_1_6_1_n28) );
  MUX2_X1 npu_inst_pe_1_6_1_U155 ( .A(npu_inst_pe_1_6_1_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_6_1_int_q_reg_v_1__1_), .S(npu_inst_pe_1_6_1_n4), .Z(
        npu_inst_pe_1_6_1_n25) );
  MUX2_X1 npu_inst_pe_1_6_1_U154 ( .A(npu_inst_pe_1_6_1_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_6_1_int_q_reg_v_3__1_), .S(npu_inst_pe_1_6_1_n4), .Z(
        npu_inst_pe_1_6_1_n24) );
  MUX2_X1 npu_inst_pe_1_6_1_U153 ( .A(npu_inst_pe_1_6_1_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_6_1_int_q_reg_v_5__1_), .S(npu_inst_pe_1_6_1_n4), .Z(
        npu_inst_pe_1_6_1_n23) );
  MUX2_X1 npu_inst_pe_1_6_1_U152 ( .A(npu_inst_pe_1_6_1_n22), .B(
        npu_inst_pe_1_6_1_n19), .S(npu_inst_pe_1_6_1_n8), .Z(
        npu_inst_int_data_x_6__1__1_) );
  MUX2_X1 npu_inst_pe_1_6_1_U151 ( .A(npu_inst_pe_1_6_1_n21), .B(
        npu_inst_pe_1_6_1_n20), .S(npu_inst_pe_1_6_1_n6), .Z(
        npu_inst_pe_1_6_1_n22) );
  MUX2_X1 npu_inst_pe_1_6_1_U150 ( .A(npu_inst_pe_1_6_1_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_6_1_int_q_reg_h_1__1_), .S(npu_inst_pe_1_6_1_n4), .Z(
        npu_inst_pe_1_6_1_n21) );
  MUX2_X1 npu_inst_pe_1_6_1_U149 ( .A(npu_inst_pe_1_6_1_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_6_1_int_q_reg_h_3__1_), .S(npu_inst_pe_1_6_1_n4), .Z(
        npu_inst_pe_1_6_1_n20) );
  MUX2_X1 npu_inst_pe_1_6_1_U148 ( .A(npu_inst_pe_1_6_1_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_6_1_int_q_reg_h_5__1_), .S(npu_inst_pe_1_6_1_n4), .Z(
        npu_inst_pe_1_6_1_n19) );
  MUX2_X1 npu_inst_pe_1_6_1_U147 ( .A(npu_inst_pe_1_6_1_n18), .B(
        npu_inst_pe_1_6_1_n15), .S(npu_inst_pe_1_6_1_n8), .Z(
        npu_inst_int_data_x_6__1__0_) );
  MUX2_X1 npu_inst_pe_1_6_1_U146 ( .A(npu_inst_pe_1_6_1_n17), .B(
        npu_inst_pe_1_6_1_n16), .S(npu_inst_pe_1_6_1_n6), .Z(
        npu_inst_pe_1_6_1_n18) );
  MUX2_X1 npu_inst_pe_1_6_1_U145 ( .A(npu_inst_pe_1_6_1_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_6_1_int_q_reg_h_1__0_), .S(npu_inst_pe_1_6_1_n4), .Z(
        npu_inst_pe_1_6_1_n17) );
  MUX2_X1 npu_inst_pe_1_6_1_U144 ( .A(npu_inst_pe_1_6_1_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_6_1_int_q_reg_h_3__0_), .S(npu_inst_pe_1_6_1_n4), .Z(
        npu_inst_pe_1_6_1_n16) );
  MUX2_X1 npu_inst_pe_1_6_1_U143 ( .A(npu_inst_pe_1_6_1_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_6_1_int_q_reg_h_5__0_), .S(npu_inst_pe_1_6_1_n4), .Z(
        npu_inst_pe_1_6_1_n15) );
  XOR2_X1 npu_inst_pe_1_6_1_U142 ( .A(npu_inst_pe_1_6_1_int_data_0_), .B(
        npu_inst_pe_1_6_1_int_q_acc_0_), .Z(npu_inst_pe_1_6_1_N73) );
  AND2_X1 npu_inst_pe_1_6_1_U141 ( .A1(npu_inst_pe_1_6_1_int_q_acc_0_), .A2(
        npu_inst_pe_1_6_1_int_data_0_), .ZN(npu_inst_pe_1_6_1_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_6_1_U140 ( .A(npu_inst_pe_1_6_1_int_q_acc_0_), .B(
        npu_inst_pe_1_6_1_n13), .ZN(npu_inst_pe_1_6_1_N65) );
  OR2_X1 npu_inst_pe_1_6_1_U139 ( .A1(npu_inst_pe_1_6_1_n13), .A2(
        npu_inst_pe_1_6_1_int_q_acc_0_), .ZN(npu_inst_pe_1_6_1_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_6_1_U138 ( .A(npu_inst_pe_1_6_1_int_q_acc_2_), .B(
        npu_inst_pe_1_6_1_add_79_carry_2_), .Z(npu_inst_pe_1_6_1_N75) );
  AND2_X1 npu_inst_pe_1_6_1_U137 ( .A1(npu_inst_pe_1_6_1_add_79_carry_2_), 
        .A2(npu_inst_pe_1_6_1_int_q_acc_2_), .ZN(
        npu_inst_pe_1_6_1_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_6_1_U136 ( .A(npu_inst_pe_1_6_1_int_q_acc_3_), .B(
        npu_inst_pe_1_6_1_add_79_carry_3_), .Z(npu_inst_pe_1_6_1_N76) );
  AND2_X1 npu_inst_pe_1_6_1_U135 ( .A1(npu_inst_pe_1_6_1_add_79_carry_3_), 
        .A2(npu_inst_pe_1_6_1_int_q_acc_3_), .ZN(
        npu_inst_pe_1_6_1_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_6_1_U134 ( .A(npu_inst_pe_1_6_1_int_q_acc_4_), .B(
        npu_inst_pe_1_6_1_add_79_carry_4_), .Z(npu_inst_pe_1_6_1_N77) );
  AND2_X1 npu_inst_pe_1_6_1_U133 ( .A1(npu_inst_pe_1_6_1_add_79_carry_4_), 
        .A2(npu_inst_pe_1_6_1_int_q_acc_4_), .ZN(
        npu_inst_pe_1_6_1_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_6_1_U132 ( .A(npu_inst_pe_1_6_1_int_q_acc_5_), .B(
        npu_inst_pe_1_6_1_add_79_carry_5_), .Z(npu_inst_pe_1_6_1_N78) );
  AND2_X1 npu_inst_pe_1_6_1_U131 ( .A1(npu_inst_pe_1_6_1_add_79_carry_5_), 
        .A2(npu_inst_pe_1_6_1_int_q_acc_5_), .ZN(
        npu_inst_pe_1_6_1_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_6_1_U130 ( .A(npu_inst_pe_1_6_1_int_q_acc_6_), .B(
        npu_inst_pe_1_6_1_add_79_carry_6_), .Z(npu_inst_pe_1_6_1_N79) );
  AND2_X1 npu_inst_pe_1_6_1_U129 ( .A1(npu_inst_pe_1_6_1_add_79_carry_6_), 
        .A2(npu_inst_pe_1_6_1_int_q_acc_6_), .ZN(
        npu_inst_pe_1_6_1_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_6_1_U128 ( .A(npu_inst_pe_1_6_1_int_q_acc_7_), .B(
        npu_inst_pe_1_6_1_add_79_carry_7_), .Z(npu_inst_pe_1_6_1_N80) );
  XNOR2_X1 npu_inst_pe_1_6_1_U127 ( .A(npu_inst_pe_1_6_1_sub_77_carry_2_), .B(
        npu_inst_pe_1_6_1_int_q_acc_2_), .ZN(npu_inst_pe_1_6_1_N67) );
  OR2_X1 npu_inst_pe_1_6_1_U126 ( .A1(npu_inst_pe_1_6_1_int_q_acc_2_), .A2(
        npu_inst_pe_1_6_1_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_6_1_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_6_1_U125 ( .A(npu_inst_pe_1_6_1_sub_77_carry_3_), .B(
        npu_inst_pe_1_6_1_int_q_acc_3_), .ZN(npu_inst_pe_1_6_1_N68) );
  OR2_X1 npu_inst_pe_1_6_1_U124 ( .A1(npu_inst_pe_1_6_1_int_q_acc_3_), .A2(
        npu_inst_pe_1_6_1_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_6_1_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_6_1_U123 ( .A(npu_inst_pe_1_6_1_sub_77_carry_4_), .B(
        npu_inst_pe_1_6_1_int_q_acc_4_), .ZN(npu_inst_pe_1_6_1_N69) );
  OR2_X1 npu_inst_pe_1_6_1_U122 ( .A1(npu_inst_pe_1_6_1_int_q_acc_4_), .A2(
        npu_inst_pe_1_6_1_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_6_1_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_6_1_U121 ( .A(npu_inst_pe_1_6_1_sub_77_carry_5_), .B(
        npu_inst_pe_1_6_1_int_q_acc_5_), .ZN(npu_inst_pe_1_6_1_N70) );
  OR2_X1 npu_inst_pe_1_6_1_U120 ( .A1(npu_inst_pe_1_6_1_int_q_acc_5_), .A2(
        npu_inst_pe_1_6_1_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_6_1_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_6_1_U119 ( .A(npu_inst_pe_1_6_1_sub_77_carry_6_), .B(
        npu_inst_pe_1_6_1_int_q_acc_6_), .ZN(npu_inst_pe_1_6_1_N71) );
  OR2_X1 npu_inst_pe_1_6_1_U118 ( .A1(npu_inst_pe_1_6_1_int_q_acc_6_), .A2(
        npu_inst_pe_1_6_1_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_6_1_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_6_1_U117 ( .A(npu_inst_pe_1_6_1_int_q_acc_7_), .B(
        npu_inst_pe_1_6_1_sub_77_carry_7_), .ZN(npu_inst_pe_1_6_1_N72) );
  INV_X1 npu_inst_pe_1_6_1_U116 ( .A(npu_inst_n76), .ZN(npu_inst_pe_1_6_1_n7)
         );
  INV_X1 npu_inst_pe_1_6_1_U115 ( .A(npu_inst_pe_1_6_1_n7), .ZN(
        npu_inst_pe_1_6_1_n6) );
  INV_X1 npu_inst_pe_1_6_1_U114 ( .A(npu_inst_n54), .ZN(npu_inst_pe_1_6_1_n3)
         );
  AOI22_X1 npu_inst_pe_1_6_1_U113 ( .A1(npu_inst_int_data_y_7__1__0_), .A2(
        npu_inst_pe_1_6_1_n58), .B1(npu_inst_pe_1_6_1_n114), .B2(
        npu_inst_pe_1_6_1_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_6_1_n57) );
  INV_X1 npu_inst_pe_1_6_1_U112 ( .A(npu_inst_pe_1_6_1_n57), .ZN(
        npu_inst_pe_1_6_1_n108) );
  AOI22_X1 npu_inst_pe_1_6_1_U111 ( .A1(npu_inst_int_data_y_7__1__0_), .A2(
        npu_inst_pe_1_6_1_n54), .B1(npu_inst_pe_1_6_1_n115), .B2(
        npu_inst_pe_1_6_1_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_6_1_n53) );
  INV_X1 npu_inst_pe_1_6_1_U110 ( .A(npu_inst_pe_1_6_1_n53), .ZN(
        npu_inst_pe_1_6_1_n109) );
  AOI22_X1 npu_inst_pe_1_6_1_U107 ( .A1(npu_inst_int_data_y_7__1__0_), .A2(
        npu_inst_pe_1_6_1_n50), .B1(npu_inst_pe_1_6_1_n116), .B2(
        npu_inst_pe_1_6_1_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_6_1_n49) );
  INV_X1 npu_inst_pe_1_6_1_U106 ( .A(npu_inst_pe_1_6_1_n49), .ZN(
        npu_inst_pe_1_6_1_n110) );
  AOI22_X1 npu_inst_pe_1_6_1_U105 ( .A1(npu_inst_int_data_y_7__1__0_), .A2(
        npu_inst_pe_1_6_1_n46), .B1(npu_inst_pe_1_6_1_n117), .B2(
        npu_inst_pe_1_6_1_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_6_1_n45) );
  INV_X1 npu_inst_pe_1_6_1_U104 ( .A(npu_inst_pe_1_6_1_n45), .ZN(
        npu_inst_pe_1_6_1_n111) );
  AOI22_X1 npu_inst_pe_1_6_1_U103 ( .A1(npu_inst_int_data_y_7__1__0_), .A2(
        npu_inst_pe_1_6_1_n42), .B1(npu_inst_pe_1_6_1_n119), .B2(
        npu_inst_pe_1_6_1_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_6_1_n41) );
  INV_X1 npu_inst_pe_1_6_1_U102 ( .A(npu_inst_pe_1_6_1_n41), .ZN(
        npu_inst_pe_1_6_1_n112) );
  AOI22_X1 npu_inst_pe_1_6_1_U101 ( .A1(npu_inst_int_data_y_7__1__1_), .A2(
        npu_inst_pe_1_6_1_n58), .B1(npu_inst_pe_1_6_1_n114), .B2(
        npu_inst_pe_1_6_1_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_6_1_n59) );
  INV_X1 npu_inst_pe_1_6_1_U100 ( .A(npu_inst_pe_1_6_1_n59), .ZN(
        npu_inst_pe_1_6_1_n102) );
  AOI22_X1 npu_inst_pe_1_6_1_U99 ( .A1(npu_inst_int_data_y_7__1__1_), .A2(
        npu_inst_pe_1_6_1_n54), .B1(npu_inst_pe_1_6_1_n115), .B2(
        npu_inst_pe_1_6_1_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_6_1_n55) );
  INV_X1 npu_inst_pe_1_6_1_U98 ( .A(npu_inst_pe_1_6_1_n55), .ZN(
        npu_inst_pe_1_6_1_n103) );
  AOI22_X1 npu_inst_pe_1_6_1_U97 ( .A1(npu_inst_int_data_y_7__1__1_), .A2(
        npu_inst_pe_1_6_1_n50), .B1(npu_inst_pe_1_6_1_n116), .B2(
        npu_inst_pe_1_6_1_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_6_1_n51) );
  INV_X1 npu_inst_pe_1_6_1_U96 ( .A(npu_inst_pe_1_6_1_n51), .ZN(
        npu_inst_pe_1_6_1_n104) );
  AOI22_X1 npu_inst_pe_1_6_1_U95 ( .A1(npu_inst_int_data_y_7__1__1_), .A2(
        npu_inst_pe_1_6_1_n46), .B1(npu_inst_pe_1_6_1_n117), .B2(
        npu_inst_pe_1_6_1_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_6_1_n47) );
  INV_X1 npu_inst_pe_1_6_1_U94 ( .A(npu_inst_pe_1_6_1_n47), .ZN(
        npu_inst_pe_1_6_1_n105) );
  AOI22_X1 npu_inst_pe_1_6_1_U93 ( .A1(npu_inst_int_data_y_7__1__1_), .A2(
        npu_inst_pe_1_6_1_n42), .B1(npu_inst_pe_1_6_1_n119), .B2(
        npu_inst_pe_1_6_1_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_6_1_n43) );
  INV_X1 npu_inst_pe_1_6_1_U92 ( .A(npu_inst_pe_1_6_1_n43), .ZN(
        npu_inst_pe_1_6_1_n106) );
  AOI22_X1 npu_inst_pe_1_6_1_U91 ( .A1(npu_inst_pe_1_6_1_n38), .A2(
        npu_inst_int_data_y_7__1__1_), .B1(npu_inst_pe_1_6_1_n118), .B2(
        npu_inst_pe_1_6_1_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_6_1_n39) );
  INV_X1 npu_inst_pe_1_6_1_U90 ( .A(npu_inst_pe_1_6_1_n39), .ZN(
        npu_inst_pe_1_6_1_n107) );
  AOI22_X1 npu_inst_pe_1_6_1_U89 ( .A1(npu_inst_pe_1_6_1_n38), .A2(
        npu_inst_int_data_y_7__1__0_), .B1(npu_inst_pe_1_6_1_n118), .B2(
        npu_inst_pe_1_6_1_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_6_1_n37) );
  INV_X1 npu_inst_pe_1_6_1_U88 ( .A(npu_inst_pe_1_6_1_n37), .ZN(
        npu_inst_pe_1_6_1_n113) );
  NAND2_X1 npu_inst_pe_1_6_1_U87 ( .A1(npu_inst_pe_1_6_1_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_6_1_n60), .ZN(npu_inst_pe_1_6_1_n74) );
  OAI21_X1 npu_inst_pe_1_6_1_U86 ( .B1(npu_inst_pe_1_6_1_n63), .B2(
        npu_inst_pe_1_6_1_n60), .A(npu_inst_pe_1_6_1_n74), .ZN(
        npu_inst_pe_1_6_1_n97) );
  NAND2_X1 npu_inst_pe_1_6_1_U85 ( .A1(npu_inst_pe_1_6_1_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_6_1_n60), .ZN(npu_inst_pe_1_6_1_n73) );
  OAI21_X1 npu_inst_pe_1_6_1_U84 ( .B1(npu_inst_pe_1_6_1_n61), .B2(
        npu_inst_pe_1_6_1_n60), .A(npu_inst_pe_1_6_1_n73), .ZN(
        npu_inst_pe_1_6_1_n96) );
  NAND2_X1 npu_inst_pe_1_6_1_U83 ( .A1(npu_inst_pe_1_6_1_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_6_1_n56), .ZN(npu_inst_pe_1_6_1_n72) );
  OAI21_X1 npu_inst_pe_1_6_1_U82 ( .B1(npu_inst_pe_1_6_1_n63), .B2(
        npu_inst_pe_1_6_1_n56), .A(npu_inst_pe_1_6_1_n72), .ZN(
        npu_inst_pe_1_6_1_n95) );
  NAND2_X1 npu_inst_pe_1_6_1_U81 ( .A1(npu_inst_pe_1_6_1_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_6_1_n56), .ZN(npu_inst_pe_1_6_1_n71) );
  OAI21_X1 npu_inst_pe_1_6_1_U80 ( .B1(npu_inst_pe_1_6_1_n61), .B2(
        npu_inst_pe_1_6_1_n56), .A(npu_inst_pe_1_6_1_n71), .ZN(
        npu_inst_pe_1_6_1_n94) );
  NAND2_X1 npu_inst_pe_1_6_1_U79 ( .A1(npu_inst_pe_1_6_1_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_6_1_n52), .ZN(npu_inst_pe_1_6_1_n70) );
  OAI21_X1 npu_inst_pe_1_6_1_U78 ( .B1(npu_inst_pe_1_6_1_n63), .B2(
        npu_inst_pe_1_6_1_n52), .A(npu_inst_pe_1_6_1_n70), .ZN(
        npu_inst_pe_1_6_1_n93) );
  NAND2_X1 npu_inst_pe_1_6_1_U77 ( .A1(npu_inst_pe_1_6_1_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_6_1_n52), .ZN(npu_inst_pe_1_6_1_n69) );
  OAI21_X1 npu_inst_pe_1_6_1_U76 ( .B1(npu_inst_pe_1_6_1_n61), .B2(
        npu_inst_pe_1_6_1_n52), .A(npu_inst_pe_1_6_1_n69), .ZN(
        npu_inst_pe_1_6_1_n92) );
  NAND2_X1 npu_inst_pe_1_6_1_U75 ( .A1(npu_inst_pe_1_6_1_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_6_1_n48), .ZN(npu_inst_pe_1_6_1_n68) );
  OAI21_X1 npu_inst_pe_1_6_1_U74 ( .B1(npu_inst_pe_1_6_1_n63), .B2(
        npu_inst_pe_1_6_1_n48), .A(npu_inst_pe_1_6_1_n68), .ZN(
        npu_inst_pe_1_6_1_n91) );
  NAND2_X1 npu_inst_pe_1_6_1_U73 ( .A1(npu_inst_pe_1_6_1_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_6_1_n48), .ZN(npu_inst_pe_1_6_1_n67) );
  OAI21_X1 npu_inst_pe_1_6_1_U72 ( .B1(npu_inst_pe_1_6_1_n61), .B2(
        npu_inst_pe_1_6_1_n48), .A(npu_inst_pe_1_6_1_n67), .ZN(
        npu_inst_pe_1_6_1_n90) );
  NAND2_X1 npu_inst_pe_1_6_1_U71 ( .A1(npu_inst_pe_1_6_1_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_6_1_n44), .ZN(npu_inst_pe_1_6_1_n66) );
  OAI21_X1 npu_inst_pe_1_6_1_U70 ( .B1(npu_inst_pe_1_6_1_n63), .B2(
        npu_inst_pe_1_6_1_n44), .A(npu_inst_pe_1_6_1_n66), .ZN(
        npu_inst_pe_1_6_1_n89) );
  NAND2_X1 npu_inst_pe_1_6_1_U69 ( .A1(npu_inst_pe_1_6_1_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_6_1_n44), .ZN(npu_inst_pe_1_6_1_n65) );
  OAI21_X1 npu_inst_pe_1_6_1_U68 ( .B1(npu_inst_pe_1_6_1_n61), .B2(
        npu_inst_pe_1_6_1_n44), .A(npu_inst_pe_1_6_1_n65), .ZN(
        npu_inst_pe_1_6_1_n88) );
  NAND2_X1 npu_inst_pe_1_6_1_U67 ( .A1(npu_inst_pe_1_6_1_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_6_1_n40), .ZN(npu_inst_pe_1_6_1_n64) );
  OAI21_X1 npu_inst_pe_1_6_1_U66 ( .B1(npu_inst_pe_1_6_1_n63), .B2(
        npu_inst_pe_1_6_1_n40), .A(npu_inst_pe_1_6_1_n64), .ZN(
        npu_inst_pe_1_6_1_n87) );
  NAND2_X1 npu_inst_pe_1_6_1_U65 ( .A1(npu_inst_pe_1_6_1_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_6_1_n40), .ZN(npu_inst_pe_1_6_1_n62) );
  OAI21_X1 npu_inst_pe_1_6_1_U64 ( .B1(npu_inst_pe_1_6_1_n61), .B2(
        npu_inst_pe_1_6_1_n40), .A(npu_inst_pe_1_6_1_n62), .ZN(
        npu_inst_pe_1_6_1_n86) );
  AND2_X1 npu_inst_pe_1_6_1_U63 ( .A1(npu_inst_pe_1_6_1_N93), .A2(npu_inst_n54), .ZN(npu_inst_int_data_y_6__1__0_) );
  AND2_X1 npu_inst_pe_1_6_1_U62 ( .A1(npu_inst_n54), .A2(npu_inst_pe_1_6_1_N94), .ZN(npu_inst_int_data_y_6__1__1_) );
  NOR3_X1 npu_inst_pe_1_6_1_U61 ( .A1(npu_inst_pe_1_6_1_n26), .A2(npu_inst_n54), .A3(npu_inst_int_ckg[14]), .ZN(npu_inst_pe_1_6_1_n85) );
  OR2_X1 npu_inst_pe_1_6_1_U60 ( .A1(npu_inst_pe_1_6_1_n85), .A2(
        npu_inst_pe_1_6_1_n2), .ZN(npu_inst_pe_1_6_1_N84) );
  AND2_X1 npu_inst_pe_1_6_1_U59 ( .A1(npu_inst_pe_1_6_1_int_q_acc_0_), .A2(
        npu_inst_pe_1_6_1_n1), .ZN(npu_inst_int_data_res_6__1__0_) );
  AND2_X1 npu_inst_pe_1_6_1_U58 ( .A1(npu_inst_pe_1_6_1_n2), .A2(
        npu_inst_pe_1_6_1_int_q_acc_7_), .ZN(npu_inst_int_data_res_6__1__7_)
         );
  AND2_X1 npu_inst_pe_1_6_1_U57 ( .A1(npu_inst_pe_1_6_1_int_q_acc_1_), .A2(
        npu_inst_pe_1_6_1_n1), .ZN(npu_inst_int_data_res_6__1__1_) );
  AND2_X1 npu_inst_pe_1_6_1_U56 ( .A1(npu_inst_pe_1_6_1_int_q_acc_2_), .A2(
        npu_inst_pe_1_6_1_n1), .ZN(npu_inst_int_data_res_6__1__2_) );
  AND2_X1 npu_inst_pe_1_6_1_U55 ( .A1(npu_inst_pe_1_6_1_int_q_acc_3_), .A2(
        npu_inst_pe_1_6_1_n2), .ZN(npu_inst_int_data_res_6__1__3_) );
  AND2_X1 npu_inst_pe_1_6_1_U54 ( .A1(npu_inst_pe_1_6_1_int_q_acc_4_), .A2(
        npu_inst_pe_1_6_1_n2), .ZN(npu_inst_int_data_res_6__1__4_) );
  AND2_X1 npu_inst_pe_1_6_1_U53 ( .A1(npu_inst_pe_1_6_1_int_q_acc_5_), .A2(
        npu_inst_pe_1_6_1_n2), .ZN(npu_inst_int_data_res_6__1__5_) );
  AND2_X1 npu_inst_pe_1_6_1_U52 ( .A1(npu_inst_pe_1_6_1_int_q_acc_6_), .A2(
        npu_inst_pe_1_6_1_n2), .ZN(npu_inst_int_data_res_6__1__6_) );
  AOI222_X1 npu_inst_pe_1_6_1_U51 ( .A1(npu_inst_int_data_res_7__1__0_), .A2(
        npu_inst_pe_1_6_1_n1), .B1(npu_inst_pe_1_6_1_N73), .B2(
        npu_inst_pe_1_6_1_n76), .C1(npu_inst_pe_1_6_1_N65), .C2(
        npu_inst_pe_1_6_1_n77), .ZN(npu_inst_pe_1_6_1_n84) );
  INV_X1 npu_inst_pe_1_6_1_U50 ( .A(npu_inst_pe_1_6_1_n84), .ZN(
        npu_inst_pe_1_6_1_n101) );
  AOI222_X1 npu_inst_pe_1_6_1_U49 ( .A1(npu_inst_int_data_res_7__1__7_), .A2(
        npu_inst_pe_1_6_1_n1), .B1(npu_inst_pe_1_6_1_N80), .B2(
        npu_inst_pe_1_6_1_n76), .C1(npu_inst_pe_1_6_1_N72), .C2(
        npu_inst_pe_1_6_1_n77), .ZN(npu_inst_pe_1_6_1_n75) );
  INV_X1 npu_inst_pe_1_6_1_U48 ( .A(npu_inst_pe_1_6_1_n75), .ZN(
        npu_inst_pe_1_6_1_n33) );
  AOI222_X1 npu_inst_pe_1_6_1_U47 ( .A1(npu_inst_int_data_res_7__1__1_), .A2(
        npu_inst_pe_1_6_1_n1), .B1(npu_inst_pe_1_6_1_N74), .B2(
        npu_inst_pe_1_6_1_n76), .C1(npu_inst_pe_1_6_1_N66), .C2(
        npu_inst_pe_1_6_1_n77), .ZN(npu_inst_pe_1_6_1_n83) );
  INV_X1 npu_inst_pe_1_6_1_U46 ( .A(npu_inst_pe_1_6_1_n83), .ZN(
        npu_inst_pe_1_6_1_n100) );
  AOI222_X1 npu_inst_pe_1_6_1_U45 ( .A1(npu_inst_int_data_res_7__1__2_), .A2(
        npu_inst_pe_1_6_1_n1), .B1(npu_inst_pe_1_6_1_N75), .B2(
        npu_inst_pe_1_6_1_n76), .C1(npu_inst_pe_1_6_1_N67), .C2(
        npu_inst_pe_1_6_1_n77), .ZN(npu_inst_pe_1_6_1_n82) );
  INV_X1 npu_inst_pe_1_6_1_U44 ( .A(npu_inst_pe_1_6_1_n82), .ZN(
        npu_inst_pe_1_6_1_n99) );
  AOI222_X1 npu_inst_pe_1_6_1_U43 ( .A1(npu_inst_int_data_res_7__1__3_), .A2(
        npu_inst_pe_1_6_1_n1), .B1(npu_inst_pe_1_6_1_N76), .B2(
        npu_inst_pe_1_6_1_n76), .C1(npu_inst_pe_1_6_1_N68), .C2(
        npu_inst_pe_1_6_1_n77), .ZN(npu_inst_pe_1_6_1_n81) );
  INV_X1 npu_inst_pe_1_6_1_U42 ( .A(npu_inst_pe_1_6_1_n81), .ZN(
        npu_inst_pe_1_6_1_n98) );
  AOI222_X1 npu_inst_pe_1_6_1_U41 ( .A1(npu_inst_int_data_res_7__1__4_), .A2(
        npu_inst_pe_1_6_1_n1), .B1(npu_inst_pe_1_6_1_N77), .B2(
        npu_inst_pe_1_6_1_n76), .C1(npu_inst_pe_1_6_1_N69), .C2(
        npu_inst_pe_1_6_1_n77), .ZN(npu_inst_pe_1_6_1_n80) );
  INV_X1 npu_inst_pe_1_6_1_U40 ( .A(npu_inst_pe_1_6_1_n80), .ZN(
        npu_inst_pe_1_6_1_n36) );
  AOI222_X1 npu_inst_pe_1_6_1_U39 ( .A1(npu_inst_int_data_res_7__1__5_), .A2(
        npu_inst_pe_1_6_1_n1), .B1(npu_inst_pe_1_6_1_N78), .B2(
        npu_inst_pe_1_6_1_n76), .C1(npu_inst_pe_1_6_1_N70), .C2(
        npu_inst_pe_1_6_1_n77), .ZN(npu_inst_pe_1_6_1_n79) );
  INV_X1 npu_inst_pe_1_6_1_U38 ( .A(npu_inst_pe_1_6_1_n79), .ZN(
        npu_inst_pe_1_6_1_n35) );
  AOI222_X1 npu_inst_pe_1_6_1_U37 ( .A1(npu_inst_int_data_res_7__1__6_), .A2(
        npu_inst_pe_1_6_1_n1), .B1(npu_inst_pe_1_6_1_N79), .B2(
        npu_inst_pe_1_6_1_n76), .C1(npu_inst_pe_1_6_1_N71), .C2(
        npu_inst_pe_1_6_1_n77), .ZN(npu_inst_pe_1_6_1_n78) );
  INV_X1 npu_inst_pe_1_6_1_U36 ( .A(npu_inst_pe_1_6_1_n78), .ZN(
        npu_inst_pe_1_6_1_n34) );
  INV_X1 npu_inst_pe_1_6_1_U35 ( .A(npu_inst_pe_1_6_1_int_data_1_), .ZN(
        npu_inst_pe_1_6_1_n14) );
  AND2_X1 npu_inst_pe_1_6_1_U34 ( .A1(npu_inst_int_data_x_6__1__1_), .A2(
        npu_inst_pe_1_6_1_int_q_weight_1_), .ZN(npu_inst_pe_1_6_1_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_6_1_U33 ( .A1(npu_inst_int_data_x_6__1__0_), .A2(
        npu_inst_pe_1_6_1_int_q_weight_1_), .ZN(npu_inst_pe_1_6_1_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_6_1_U32 ( .A1(npu_inst_n54), .A2(
        npu_inst_int_data_y_7__1__1_), .B1(npu_inst_pe_1_6_1_n3), .B2(
        npu_inst_int_data_x_6__2__1_), .ZN(npu_inst_pe_1_6_1_n63) );
  AOI22_X1 npu_inst_pe_1_6_1_U31 ( .A1(npu_inst_n54), .A2(
        npu_inst_int_data_y_7__1__0_), .B1(npu_inst_pe_1_6_1_n3), .B2(
        npu_inst_int_data_x_6__2__0_), .ZN(npu_inst_pe_1_6_1_n61) );
  INV_X1 npu_inst_pe_1_6_1_U30 ( .A(npu_inst_pe_1_6_1_int_data_0_), .ZN(
        npu_inst_pe_1_6_1_n13) );
  INV_X1 npu_inst_pe_1_6_1_U29 ( .A(npu_inst_n68), .ZN(npu_inst_pe_1_6_1_n5)
         );
  OR3_X1 npu_inst_pe_1_6_1_U28 ( .A1(npu_inst_pe_1_6_1_n6), .A2(
        npu_inst_pe_1_6_1_n8), .A3(npu_inst_pe_1_6_1_n5), .ZN(
        npu_inst_pe_1_6_1_n56) );
  OR3_X1 npu_inst_pe_1_6_1_U27 ( .A1(npu_inst_pe_1_6_1_n5), .A2(
        npu_inst_pe_1_6_1_n8), .A3(npu_inst_pe_1_6_1_n7), .ZN(
        npu_inst_pe_1_6_1_n48) );
  INV_X1 npu_inst_pe_1_6_1_U26 ( .A(npu_inst_pe_1_6_1_n5), .ZN(
        npu_inst_pe_1_6_1_n4) );
  INV_X1 npu_inst_pe_1_6_1_U25 ( .A(npu_inst_n123), .ZN(npu_inst_pe_1_6_1_n12)
         );
  OR3_X1 npu_inst_pe_1_6_1_U24 ( .A1(npu_inst_pe_1_6_1_n4), .A2(
        npu_inst_pe_1_6_1_n8), .A3(npu_inst_pe_1_6_1_n7), .ZN(
        npu_inst_pe_1_6_1_n52) );
  OR3_X1 npu_inst_pe_1_6_1_U23 ( .A1(npu_inst_pe_1_6_1_n6), .A2(
        npu_inst_pe_1_6_1_n8), .A3(npu_inst_pe_1_6_1_n4), .ZN(
        npu_inst_pe_1_6_1_n60) );
  NOR2_X1 npu_inst_pe_1_6_1_U22 ( .A1(npu_inst_pe_1_6_1_n60), .A2(
        npu_inst_pe_1_6_1_n3), .ZN(npu_inst_pe_1_6_1_n58) );
  NOR2_X1 npu_inst_pe_1_6_1_U21 ( .A1(npu_inst_pe_1_6_1_n56), .A2(
        npu_inst_pe_1_6_1_n3), .ZN(npu_inst_pe_1_6_1_n54) );
  NOR2_X1 npu_inst_pe_1_6_1_U20 ( .A1(npu_inst_pe_1_6_1_n52), .A2(
        npu_inst_pe_1_6_1_n3), .ZN(npu_inst_pe_1_6_1_n50) );
  NOR2_X1 npu_inst_pe_1_6_1_U19 ( .A1(npu_inst_pe_1_6_1_n48), .A2(
        npu_inst_pe_1_6_1_n3), .ZN(npu_inst_pe_1_6_1_n46) );
  NOR2_X1 npu_inst_pe_1_6_1_U18 ( .A1(npu_inst_pe_1_6_1_n40), .A2(
        npu_inst_pe_1_6_1_n3), .ZN(npu_inst_pe_1_6_1_n38) );
  NOR2_X1 npu_inst_pe_1_6_1_U17 ( .A1(npu_inst_pe_1_6_1_n44), .A2(
        npu_inst_pe_1_6_1_n3), .ZN(npu_inst_pe_1_6_1_n42) );
  BUF_X1 npu_inst_pe_1_6_1_U16 ( .A(npu_inst_n95), .Z(npu_inst_pe_1_6_1_n8) );
  BUF_X1 npu_inst_pe_1_6_1_U15 ( .A(npu_inst_pe_1_6_1_n12), .Z(
        npu_inst_pe_1_6_1_n11) );
  BUF_X1 npu_inst_pe_1_6_1_U14 ( .A(npu_inst_pe_1_6_1_n12), .Z(
        npu_inst_pe_1_6_1_n10) );
  BUF_X1 npu_inst_pe_1_6_1_U13 ( .A(npu_inst_pe_1_6_1_n12), .Z(
        npu_inst_pe_1_6_1_n9) );
  INV_X1 npu_inst_pe_1_6_1_U12 ( .A(npu_inst_pe_1_6_1_n38), .ZN(
        npu_inst_pe_1_6_1_n118) );
  INV_X1 npu_inst_pe_1_6_1_U11 ( .A(npu_inst_pe_1_6_1_n58), .ZN(
        npu_inst_pe_1_6_1_n114) );
  INV_X1 npu_inst_pe_1_6_1_U10 ( .A(npu_inst_pe_1_6_1_n54), .ZN(
        npu_inst_pe_1_6_1_n115) );
  INV_X1 npu_inst_pe_1_6_1_U9 ( .A(npu_inst_pe_1_6_1_n50), .ZN(
        npu_inst_pe_1_6_1_n116) );
  INV_X1 npu_inst_pe_1_6_1_U8 ( .A(npu_inst_pe_1_6_1_n46), .ZN(
        npu_inst_pe_1_6_1_n117) );
  INV_X1 npu_inst_pe_1_6_1_U7 ( .A(npu_inst_pe_1_6_1_n42), .ZN(
        npu_inst_pe_1_6_1_n119) );
  BUF_X1 npu_inst_pe_1_6_1_U6 ( .A(npu_inst_n14), .Z(npu_inst_pe_1_6_1_n2) );
  BUF_X1 npu_inst_pe_1_6_1_U5 ( .A(npu_inst_n14), .Z(npu_inst_pe_1_6_1_n1) );
  NOR2_X1 npu_inst_pe_1_6_1_U4 ( .A1(npu_inst_pe_1_6_1_int_q_weight_0_), .A2(
        npu_inst_pe_1_6_1_n1), .ZN(npu_inst_pe_1_6_1_n76) );
  NOR2_X1 npu_inst_pe_1_6_1_U3 ( .A1(npu_inst_pe_1_6_1_n27), .A2(
        npu_inst_pe_1_6_1_n1), .ZN(npu_inst_pe_1_6_1_n77) );
  FA_X1 npu_inst_pe_1_6_1_sub_77_U2_1 ( .A(npu_inst_pe_1_6_1_int_q_acc_1_), 
        .B(npu_inst_pe_1_6_1_n14), .CI(npu_inst_pe_1_6_1_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_6_1_sub_77_carry_2_), .S(npu_inst_pe_1_6_1_N66) );
  FA_X1 npu_inst_pe_1_6_1_add_79_U1_1 ( .A(npu_inst_pe_1_6_1_int_q_acc_1_), 
        .B(npu_inst_pe_1_6_1_int_data_1_), .CI(
        npu_inst_pe_1_6_1_add_79_carry_1_), .CO(
        npu_inst_pe_1_6_1_add_79_carry_2_), .S(npu_inst_pe_1_6_1_N74) );
  NAND3_X1 npu_inst_pe_1_6_1_U109 ( .A1(npu_inst_pe_1_6_1_n5), .A2(
        npu_inst_pe_1_6_1_n7), .A3(npu_inst_pe_1_6_1_n8), .ZN(
        npu_inst_pe_1_6_1_n44) );
  NAND3_X1 npu_inst_pe_1_6_1_U108 ( .A1(npu_inst_pe_1_6_1_n4), .A2(
        npu_inst_pe_1_6_1_n7), .A3(npu_inst_pe_1_6_1_n8), .ZN(
        npu_inst_pe_1_6_1_n40) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_6_1_n34), .CK(
        npu_inst_pe_1_6_1_net3166), .RN(npu_inst_pe_1_6_1_n9), .Q(
        npu_inst_pe_1_6_1_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_6_1_n35), .CK(
        npu_inst_pe_1_6_1_net3166), .RN(npu_inst_pe_1_6_1_n9), .Q(
        npu_inst_pe_1_6_1_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_6_1_n36), .CK(
        npu_inst_pe_1_6_1_net3166), .RN(npu_inst_pe_1_6_1_n9), .Q(
        npu_inst_pe_1_6_1_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_6_1_n98), .CK(
        npu_inst_pe_1_6_1_net3166), .RN(npu_inst_pe_1_6_1_n9), .Q(
        npu_inst_pe_1_6_1_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_6_1_n99), .CK(
        npu_inst_pe_1_6_1_net3166), .RN(npu_inst_pe_1_6_1_n9), .Q(
        npu_inst_pe_1_6_1_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_6_1_n100), 
        .CK(npu_inst_pe_1_6_1_net3166), .RN(npu_inst_pe_1_6_1_n9), .Q(
        npu_inst_pe_1_6_1_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_6_1_n33), .CK(
        npu_inst_pe_1_6_1_net3166), .RN(npu_inst_pe_1_6_1_n9), .Q(
        npu_inst_pe_1_6_1_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_6_1_n101), 
        .CK(npu_inst_pe_1_6_1_net3166), .RN(npu_inst_pe_1_6_1_n9), .Q(
        npu_inst_pe_1_6_1_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_weight_reg_0_ ( .D(npu_inst_n109), .CK(
        npu_inst_pe_1_6_1_net3172), .RN(npu_inst_pe_1_6_1_n9), .Q(
        npu_inst_pe_1_6_1_int_q_weight_0_), .QN(npu_inst_pe_1_6_1_n27) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_weight_reg_1_ ( .D(npu_inst_n115), .CK(
        npu_inst_pe_1_6_1_net3172), .RN(npu_inst_pe_1_6_1_n9), .Q(
        npu_inst_pe_1_6_1_int_q_weight_1_), .QN(npu_inst_pe_1_6_1_n26) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_6_1_n113), 
        .CK(npu_inst_pe_1_6_1_net3172), .RN(npu_inst_pe_1_6_1_n9), .Q(
        npu_inst_pe_1_6_1_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_6_1_n107), 
        .CK(npu_inst_pe_1_6_1_net3172), .RN(npu_inst_pe_1_6_1_n9), .Q(
        npu_inst_pe_1_6_1_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_6_1_n112), 
        .CK(npu_inst_pe_1_6_1_net3172), .RN(npu_inst_pe_1_6_1_n10), .Q(
        npu_inst_pe_1_6_1_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_6_1_n106), 
        .CK(npu_inst_pe_1_6_1_net3172), .RN(npu_inst_pe_1_6_1_n10), .Q(
        npu_inst_pe_1_6_1_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_6_1_n111), 
        .CK(npu_inst_pe_1_6_1_net3172), .RN(npu_inst_pe_1_6_1_n10), .Q(
        npu_inst_pe_1_6_1_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_6_1_n105), 
        .CK(npu_inst_pe_1_6_1_net3172), .RN(npu_inst_pe_1_6_1_n10), .Q(
        npu_inst_pe_1_6_1_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_6_1_n110), 
        .CK(npu_inst_pe_1_6_1_net3172), .RN(npu_inst_pe_1_6_1_n10), .Q(
        npu_inst_pe_1_6_1_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_6_1_n104), 
        .CK(npu_inst_pe_1_6_1_net3172), .RN(npu_inst_pe_1_6_1_n10), .Q(
        npu_inst_pe_1_6_1_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_6_1_n109), 
        .CK(npu_inst_pe_1_6_1_net3172), .RN(npu_inst_pe_1_6_1_n10), .Q(
        npu_inst_pe_1_6_1_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_6_1_n103), 
        .CK(npu_inst_pe_1_6_1_net3172), .RN(npu_inst_pe_1_6_1_n10), .Q(
        npu_inst_pe_1_6_1_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_6_1_n108), 
        .CK(npu_inst_pe_1_6_1_net3172), .RN(npu_inst_pe_1_6_1_n10), .Q(
        npu_inst_pe_1_6_1_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_6_1_n102), 
        .CK(npu_inst_pe_1_6_1_net3172), .RN(npu_inst_pe_1_6_1_n10), .Q(
        npu_inst_pe_1_6_1_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_6_1_n86), 
        .CK(npu_inst_pe_1_6_1_net3172), .RN(npu_inst_pe_1_6_1_n10), .Q(
        npu_inst_pe_1_6_1_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_6_1_n87), 
        .CK(npu_inst_pe_1_6_1_net3172), .RN(npu_inst_pe_1_6_1_n10), .Q(
        npu_inst_pe_1_6_1_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_6_1_n88), 
        .CK(npu_inst_pe_1_6_1_net3172), .RN(npu_inst_pe_1_6_1_n11), .Q(
        npu_inst_pe_1_6_1_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_6_1_n89), 
        .CK(npu_inst_pe_1_6_1_net3172), .RN(npu_inst_pe_1_6_1_n11), .Q(
        npu_inst_pe_1_6_1_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_6_1_n90), 
        .CK(npu_inst_pe_1_6_1_net3172), .RN(npu_inst_pe_1_6_1_n11), .Q(
        npu_inst_pe_1_6_1_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_6_1_n91), 
        .CK(npu_inst_pe_1_6_1_net3172), .RN(npu_inst_pe_1_6_1_n11), .Q(
        npu_inst_pe_1_6_1_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_6_1_n92), 
        .CK(npu_inst_pe_1_6_1_net3172), .RN(npu_inst_pe_1_6_1_n11), .Q(
        npu_inst_pe_1_6_1_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_6_1_n93), 
        .CK(npu_inst_pe_1_6_1_net3172), .RN(npu_inst_pe_1_6_1_n11), .Q(
        npu_inst_pe_1_6_1_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_6_1_n94), 
        .CK(npu_inst_pe_1_6_1_net3172), .RN(npu_inst_pe_1_6_1_n11), .Q(
        npu_inst_pe_1_6_1_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_6_1_n95), 
        .CK(npu_inst_pe_1_6_1_net3172), .RN(npu_inst_pe_1_6_1_n11), .Q(
        npu_inst_pe_1_6_1_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_6_1_n96), 
        .CK(npu_inst_pe_1_6_1_net3172), .RN(npu_inst_pe_1_6_1_n11), .Q(
        npu_inst_pe_1_6_1_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_6_1_n97), 
        .CK(npu_inst_pe_1_6_1_net3172), .RN(npu_inst_pe_1_6_1_n11), .Q(
        npu_inst_pe_1_6_1_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_6_1_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_6_1_N84), .SE(1'b0), .GCK(npu_inst_pe_1_6_1_net3166) );
  CLKGATETST_X1 npu_inst_pe_1_6_1_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n62), .SE(1'b0), .GCK(npu_inst_pe_1_6_1_net3172) );
  MUX2_X1 npu_inst_pe_1_6_2_U162 ( .A(npu_inst_pe_1_6_2_n32), .B(
        npu_inst_pe_1_6_2_n29), .S(npu_inst_pe_1_6_2_n8), .Z(
        npu_inst_pe_1_6_2_N93) );
  MUX2_X1 npu_inst_pe_1_6_2_U161 ( .A(npu_inst_pe_1_6_2_n31), .B(
        npu_inst_pe_1_6_2_n30), .S(npu_inst_pe_1_6_2_n6), .Z(
        npu_inst_pe_1_6_2_n32) );
  MUX2_X1 npu_inst_pe_1_6_2_U160 ( .A(npu_inst_pe_1_6_2_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_6_2_int_q_reg_v_1__0_), .S(npu_inst_pe_1_6_2_n4), .Z(
        npu_inst_pe_1_6_2_n31) );
  MUX2_X1 npu_inst_pe_1_6_2_U159 ( .A(npu_inst_pe_1_6_2_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_6_2_int_q_reg_v_3__0_), .S(npu_inst_pe_1_6_2_n4), .Z(
        npu_inst_pe_1_6_2_n30) );
  MUX2_X1 npu_inst_pe_1_6_2_U158 ( .A(npu_inst_pe_1_6_2_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_6_2_int_q_reg_v_5__0_), .S(npu_inst_pe_1_6_2_n4), .Z(
        npu_inst_pe_1_6_2_n29) );
  MUX2_X1 npu_inst_pe_1_6_2_U157 ( .A(npu_inst_pe_1_6_2_n28), .B(
        npu_inst_pe_1_6_2_n23), .S(npu_inst_pe_1_6_2_n8), .Z(
        npu_inst_pe_1_6_2_N94) );
  MUX2_X1 npu_inst_pe_1_6_2_U156 ( .A(npu_inst_pe_1_6_2_n25), .B(
        npu_inst_pe_1_6_2_n24), .S(npu_inst_pe_1_6_2_n6), .Z(
        npu_inst_pe_1_6_2_n28) );
  MUX2_X1 npu_inst_pe_1_6_2_U155 ( .A(npu_inst_pe_1_6_2_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_6_2_int_q_reg_v_1__1_), .S(npu_inst_pe_1_6_2_n4), .Z(
        npu_inst_pe_1_6_2_n25) );
  MUX2_X1 npu_inst_pe_1_6_2_U154 ( .A(npu_inst_pe_1_6_2_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_6_2_int_q_reg_v_3__1_), .S(npu_inst_pe_1_6_2_n4), .Z(
        npu_inst_pe_1_6_2_n24) );
  MUX2_X1 npu_inst_pe_1_6_2_U153 ( .A(npu_inst_pe_1_6_2_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_6_2_int_q_reg_v_5__1_), .S(npu_inst_pe_1_6_2_n4), .Z(
        npu_inst_pe_1_6_2_n23) );
  MUX2_X1 npu_inst_pe_1_6_2_U152 ( .A(npu_inst_pe_1_6_2_n22), .B(
        npu_inst_pe_1_6_2_n19), .S(npu_inst_pe_1_6_2_n8), .Z(
        npu_inst_int_data_x_6__2__1_) );
  MUX2_X1 npu_inst_pe_1_6_2_U151 ( .A(npu_inst_pe_1_6_2_n21), .B(
        npu_inst_pe_1_6_2_n20), .S(npu_inst_pe_1_6_2_n6), .Z(
        npu_inst_pe_1_6_2_n22) );
  MUX2_X1 npu_inst_pe_1_6_2_U150 ( .A(npu_inst_pe_1_6_2_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_6_2_int_q_reg_h_1__1_), .S(npu_inst_pe_1_6_2_n4), .Z(
        npu_inst_pe_1_6_2_n21) );
  MUX2_X1 npu_inst_pe_1_6_2_U149 ( .A(npu_inst_pe_1_6_2_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_6_2_int_q_reg_h_3__1_), .S(npu_inst_pe_1_6_2_n4), .Z(
        npu_inst_pe_1_6_2_n20) );
  MUX2_X1 npu_inst_pe_1_6_2_U148 ( .A(npu_inst_pe_1_6_2_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_6_2_int_q_reg_h_5__1_), .S(npu_inst_pe_1_6_2_n4), .Z(
        npu_inst_pe_1_6_2_n19) );
  MUX2_X1 npu_inst_pe_1_6_2_U147 ( .A(npu_inst_pe_1_6_2_n18), .B(
        npu_inst_pe_1_6_2_n15), .S(npu_inst_pe_1_6_2_n8), .Z(
        npu_inst_int_data_x_6__2__0_) );
  MUX2_X1 npu_inst_pe_1_6_2_U146 ( .A(npu_inst_pe_1_6_2_n17), .B(
        npu_inst_pe_1_6_2_n16), .S(npu_inst_pe_1_6_2_n6), .Z(
        npu_inst_pe_1_6_2_n18) );
  MUX2_X1 npu_inst_pe_1_6_2_U145 ( .A(npu_inst_pe_1_6_2_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_6_2_int_q_reg_h_1__0_), .S(npu_inst_pe_1_6_2_n4), .Z(
        npu_inst_pe_1_6_2_n17) );
  MUX2_X1 npu_inst_pe_1_6_2_U144 ( .A(npu_inst_pe_1_6_2_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_6_2_int_q_reg_h_3__0_), .S(npu_inst_pe_1_6_2_n4), .Z(
        npu_inst_pe_1_6_2_n16) );
  MUX2_X1 npu_inst_pe_1_6_2_U143 ( .A(npu_inst_pe_1_6_2_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_6_2_int_q_reg_h_5__0_), .S(npu_inst_pe_1_6_2_n4), .Z(
        npu_inst_pe_1_6_2_n15) );
  XOR2_X1 npu_inst_pe_1_6_2_U142 ( .A(npu_inst_pe_1_6_2_int_data_0_), .B(
        npu_inst_pe_1_6_2_int_q_acc_0_), .Z(npu_inst_pe_1_6_2_N73) );
  AND2_X1 npu_inst_pe_1_6_2_U141 ( .A1(npu_inst_pe_1_6_2_int_q_acc_0_), .A2(
        npu_inst_pe_1_6_2_int_data_0_), .ZN(npu_inst_pe_1_6_2_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_6_2_U140 ( .A(npu_inst_pe_1_6_2_int_q_acc_0_), .B(
        npu_inst_pe_1_6_2_n13), .ZN(npu_inst_pe_1_6_2_N65) );
  OR2_X1 npu_inst_pe_1_6_2_U139 ( .A1(npu_inst_pe_1_6_2_n13), .A2(
        npu_inst_pe_1_6_2_int_q_acc_0_), .ZN(npu_inst_pe_1_6_2_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_6_2_U138 ( .A(npu_inst_pe_1_6_2_int_q_acc_2_), .B(
        npu_inst_pe_1_6_2_add_79_carry_2_), .Z(npu_inst_pe_1_6_2_N75) );
  AND2_X1 npu_inst_pe_1_6_2_U137 ( .A1(npu_inst_pe_1_6_2_add_79_carry_2_), 
        .A2(npu_inst_pe_1_6_2_int_q_acc_2_), .ZN(
        npu_inst_pe_1_6_2_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_6_2_U136 ( .A(npu_inst_pe_1_6_2_int_q_acc_3_), .B(
        npu_inst_pe_1_6_2_add_79_carry_3_), .Z(npu_inst_pe_1_6_2_N76) );
  AND2_X1 npu_inst_pe_1_6_2_U135 ( .A1(npu_inst_pe_1_6_2_add_79_carry_3_), 
        .A2(npu_inst_pe_1_6_2_int_q_acc_3_), .ZN(
        npu_inst_pe_1_6_2_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_6_2_U134 ( .A(npu_inst_pe_1_6_2_int_q_acc_4_), .B(
        npu_inst_pe_1_6_2_add_79_carry_4_), .Z(npu_inst_pe_1_6_2_N77) );
  AND2_X1 npu_inst_pe_1_6_2_U133 ( .A1(npu_inst_pe_1_6_2_add_79_carry_4_), 
        .A2(npu_inst_pe_1_6_2_int_q_acc_4_), .ZN(
        npu_inst_pe_1_6_2_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_6_2_U132 ( .A(npu_inst_pe_1_6_2_int_q_acc_5_), .B(
        npu_inst_pe_1_6_2_add_79_carry_5_), .Z(npu_inst_pe_1_6_2_N78) );
  AND2_X1 npu_inst_pe_1_6_2_U131 ( .A1(npu_inst_pe_1_6_2_add_79_carry_5_), 
        .A2(npu_inst_pe_1_6_2_int_q_acc_5_), .ZN(
        npu_inst_pe_1_6_2_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_6_2_U130 ( .A(npu_inst_pe_1_6_2_int_q_acc_6_), .B(
        npu_inst_pe_1_6_2_add_79_carry_6_), .Z(npu_inst_pe_1_6_2_N79) );
  AND2_X1 npu_inst_pe_1_6_2_U129 ( .A1(npu_inst_pe_1_6_2_add_79_carry_6_), 
        .A2(npu_inst_pe_1_6_2_int_q_acc_6_), .ZN(
        npu_inst_pe_1_6_2_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_6_2_U128 ( .A(npu_inst_pe_1_6_2_int_q_acc_7_), .B(
        npu_inst_pe_1_6_2_add_79_carry_7_), .Z(npu_inst_pe_1_6_2_N80) );
  XNOR2_X1 npu_inst_pe_1_6_2_U127 ( .A(npu_inst_pe_1_6_2_sub_77_carry_2_), .B(
        npu_inst_pe_1_6_2_int_q_acc_2_), .ZN(npu_inst_pe_1_6_2_N67) );
  OR2_X1 npu_inst_pe_1_6_2_U126 ( .A1(npu_inst_pe_1_6_2_int_q_acc_2_), .A2(
        npu_inst_pe_1_6_2_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_6_2_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_6_2_U125 ( .A(npu_inst_pe_1_6_2_sub_77_carry_3_), .B(
        npu_inst_pe_1_6_2_int_q_acc_3_), .ZN(npu_inst_pe_1_6_2_N68) );
  OR2_X1 npu_inst_pe_1_6_2_U124 ( .A1(npu_inst_pe_1_6_2_int_q_acc_3_), .A2(
        npu_inst_pe_1_6_2_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_6_2_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_6_2_U123 ( .A(npu_inst_pe_1_6_2_sub_77_carry_4_), .B(
        npu_inst_pe_1_6_2_int_q_acc_4_), .ZN(npu_inst_pe_1_6_2_N69) );
  OR2_X1 npu_inst_pe_1_6_2_U122 ( .A1(npu_inst_pe_1_6_2_int_q_acc_4_), .A2(
        npu_inst_pe_1_6_2_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_6_2_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_6_2_U121 ( .A(npu_inst_pe_1_6_2_sub_77_carry_5_), .B(
        npu_inst_pe_1_6_2_int_q_acc_5_), .ZN(npu_inst_pe_1_6_2_N70) );
  OR2_X1 npu_inst_pe_1_6_2_U120 ( .A1(npu_inst_pe_1_6_2_int_q_acc_5_), .A2(
        npu_inst_pe_1_6_2_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_6_2_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_6_2_U119 ( .A(npu_inst_pe_1_6_2_sub_77_carry_6_), .B(
        npu_inst_pe_1_6_2_int_q_acc_6_), .ZN(npu_inst_pe_1_6_2_N71) );
  OR2_X1 npu_inst_pe_1_6_2_U118 ( .A1(npu_inst_pe_1_6_2_int_q_acc_6_), .A2(
        npu_inst_pe_1_6_2_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_6_2_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_6_2_U117 ( .A(npu_inst_pe_1_6_2_int_q_acc_7_), .B(
        npu_inst_pe_1_6_2_sub_77_carry_7_), .ZN(npu_inst_pe_1_6_2_N72) );
  INV_X1 npu_inst_pe_1_6_2_U116 ( .A(npu_inst_n76), .ZN(npu_inst_pe_1_6_2_n7)
         );
  INV_X1 npu_inst_pe_1_6_2_U115 ( .A(npu_inst_pe_1_6_2_n7), .ZN(
        npu_inst_pe_1_6_2_n6) );
  INV_X1 npu_inst_pe_1_6_2_U114 ( .A(npu_inst_n53), .ZN(npu_inst_pe_1_6_2_n3)
         );
  AOI22_X1 npu_inst_pe_1_6_2_U113 ( .A1(npu_inst_int_data_y_7__2__0_), .A2(
        npu_inst_pe_1_6_2_n58), .B1(npu_inst_pe_1_6_2_n114), .B2(
        npu_inst_pe_1_6_2_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_6_2_n57) );
  INV_X1 npu_inst_pe_1_6_2_U112 ( .A(npu_inst_pe_1_6_2_n57), .ZN(
        npu_inst_pe_1_6_2_n108) );
  AOI22_X1 npu_inst_pe_1_6_2_U111 ( .A1(npu_inst_int_data_y_7__2__0_), .A2(
        npu_inst_pe_1_6_2_n54), .B1(npu_inst_pe_1_6_2_n115), .B2(
        npu_inst_pe_1_6_2_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_6_2_n53) );
  INV_X1 npu_inst_pe_1_6_2_U110 ( .A(npu_inst_pe_1_6_2_n53), .ZN(
        npu_inst_pe_1_6_2_n109) );
  AOI22_X1 npu_inst_pe_1_6_2_U107 ( .A1(npu_inst_int_data_y_7__2__0_), .A2(
        npu_inst_pe_1_6_2_n50), .B1(npu_inst_pe_1_6_2_n116), .B2(
        npu_inst_pe_1_6_2_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_6_2_n49) );
  INV_X1 npu_inst_pe_1_6_2_U106 ( .A(npu_inst_pe_1_6_2_n49), .ZN(
        npu_inst_pe_1_6_2_n110) );
  AOI22_X1 npu_inst_pe_1_6_2_U105 ( .A1(npu_inst_int_data_y_7__2__0_), .A2(
        npu_inst_pe_1_6_2_n46), .B1(npu_inst_pe_1_6_2_n117), .B2(
        npu_inst_pe_1_6_2_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_6_2_n45) );
  INV_X1 npu_inst_pe_1_6_2_U104 ( .A(npu_inst_pe_1_6_2_n45), .ZN(
        npu_inst_pe_1_6_2_n111) );
  AOI22_X1 npu_inst_pe_1_6_2_U103 ( .A1(npu_inst_int_data_y_7__2__0_), .A2(
        npu_inst_pe_1_6_2_n42), .B1(npu_inst_pe_1_6_2_n119), .B2(
        npu_inst_pe_1_6_2_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_6_2_n41) );
  INV_X1 npu_inst_pe_1_6_2_U102 ( .A(npu_inst_pe_1_6_2_n41), .ZN(
        npu_inst_pe_1_6_2_n112) );
  AOI22_X1 npu_inst_pe_1_6_2_U101 ( .A1(npu_inst_int_data_y_7__2__1_), .A2(
        npu_inst_pe_1_6_2_n58), .B1(npu_inst_pe_1_6_2_n114), .B2(
        npu_inst_pe_1_6_2_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_6_2_n59) );
  INV_X1 npu_inst_pe_1_6_2_U100 ( .A(npu_inst_pe_1_6_2_n59), .ZN(
        npu_inst_pe_1_6_2_n102) );
  AOI22_X1 npu_inst_pe_1_6_2_U99 ( .A1(npu_inst_int_data_y_7__2__1_), .A2(
        npu_inst_pe_1_6_2_n54), .B1(npu_inst_pe_1_6_2_n115), .B2(
        npu_inst_pe_1_6_2_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_6_2_n55) );
  INV_X1 npu_inst_pe_1_6_2_U98 ( .A(npu_inst_pe_1_6_2_n55), .ZN(
        npu_inst_pe_1_6_2_n103) );
  AOI22_X1 npu_inst_pe_1_6_2_U97 ( .A1(npu_inst_int_data_y_7__2__1_), .A2(
        npu_inst_pe_1_6_2_n50), .B1(npu_inst_pe_1_6_2_n116), .B2(
        npu_inst_pe_1_6_2_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_6_2_n51) );
  INV_X1 npu_inst_pe_1_6_2_U96 ( .A(npu_inst_pe_1_6_2_n51), .ZN(
        npu_inst_pe_1_6_2_n104) );
  AOI22_X1 npu_inst_pe_1_6_2_U95 ( .A1(npu_inst_int_data_y_7__2__1_), .A2(
        npu_inst_pe_1_6_2_n46), .B1(npu_inst_pe_1_6_2_n117), .B2(
        npu_inst_pe_1_6_2_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_6_2_n47) );
  INV_X1 npu_inst_pe_1_6_2_U94 ( .A(npu_inst_pe_1_6_2_n47), .ZN(
        npu_inst_pe_1_6_2_n105) );
  AOI22_X1 npu_inst_pe_1_6_2_U93 ( .A1(npu_inst_int_data_y_7__2__1_), .A2(
        npu_inst_pe_1_6_2_n42), .B1(npu_inst_pe_1_6_2_n119), .B2(
        npu_inst_pe_1_6_2_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_6_2_n43) );
  INV_X1 npu_inst_pe_1_6_2_U92 ( .A(npu_inst_pe_1_6_2_n43), .ZN(
        npu_inst_pe_1_6_2_n106) );
  AOI22_X1 npu_inst_pe_1_6_2_U91 ( .A1(npu_inst_pe_1_6_2_n38), .A2(
        npu_inst_int_data_y_7__2__1_), .B1(npu_inst_pe_1_6_2_n118), .B2(
        npu_inst_pe_1_6_2_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_6_2_n39) );
  INV_X1 npu_inst_pe_1_6_2_U90 ( .A(npu_inst_pe_1_6_2_n39), .ZN(
        npu_inst_pe_1_6_2_n107) );
  AOI22_X1 npu_inst_pe_1_6_2_U89 ( .A1(npu_inst_pe_1_6_2_n38), .A2(
        npu_inst_int_data_y_7__2__0_), .B1(npu_inst_pe_1_6_2_n118), .B2(
        npu_inst_pe_1_6_2_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_6_2_n37) );
  INV_X1 npu_inst_pe_1_6_2_U88 ( .A(npu_inst_pe_1_6_2_n37), .ZN(
        npu_inst_pe_1_6_2_n113) );
  NAND2_X1 npu_inst_pe_1_6_2_U87 ( .A1(npu_inst_pe_1_6_2_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_6_2_n60), .ZN(npu_inst_pe_1_6_2_n74) );
  OAI21_X1 npu_inst_pe_1_6_2_U86 ( .B1(npu_inst_pe_1_6_2_n63), .B2(
        npu_inst_pe_1_6_2_n60), .A(npu_inst_pe_1_6_2_n74), .ZN(
        npu_inst_pe_1_6_2_n97) );
  NAND2_X1 npu_inst_pe_1_6_2_U85 ( .A1(npu_inst_pe_1_6_2_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_6_2_n60), .ZN(npu_inst_pe_1_6_2_n73) );
  OAI21_X1 npu_inst_pe_1_6_2_U84 ( .B1(npu_inst_pe_1_6_2_n61), .B2(
        npu_inst_pe_1_6_2_n60), .A(npu_inst_pe_1_6_2_n73), .ZN(
        npu_inst_pe_1_6_2_n96) );
  NAND2_X1 npu_inst_pe_1_6_2_U83 ( .A1(npu_inst_pe_1_6_2_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_6_2_n56), .ZN(npu_inst_pe_1_6_2_n72) );
  OAI21_X1 npu_inst_pe_1_6_2_U82 ( .B1(npu_inst_pe_1_6_2_n63), .B2(
        npu_inst_pe_1_6_2_n56), .A(npu_inst_pe_1_6_2_n72), .ZN(
        npu_inst_pe_1_6_2_n95) );
  NAND2_X1 npu_inst_pe_1_6_2_U81 ( .A1(npu_inst_pe_1_6_2_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_6_2_n56), .ZN(npu_inst_pe_1_6_2_n71) );
  OAI21_X1 npu_inst_pe_1_6_2_U80 ( .B1(npu_inst_pe_1_6_2_n61), .B2(
        npu_inst_pe_1_6_2_n56), .A(npu_inst_pe_1_6_2_n71), .ZN(
        npu_inst_pe_1_6_2_n94) );
  NAND2_X1 npu_inst_pe_1_6_2_U79 ( .A1(npu_inst_pe_1_6_2_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_6_2_n52), .ZN(npu_inst_pe_1_6_2_n70) );
  OAI21_X1 npu_inst_pe_1_6_2_U78 ( .B1(npu_inst_pe_1_6_2_n63), .B2(
        npu_inst_pe_1_6_2_n52), .A(npu_inst_pe_1_6_2_n70), .ZN(
        npu_inst_pe_1_6_2_n93) );
  NAND2_X1 npu_inst_pe_1_6_2_U77 ( .A1(npu_inst_pe_1_6_2_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_6_2_n52), .ZN(npu_inst_pe_1_6_2_n69) );
  OAI21_X1 npu_inst_pe_1_6_2_U76 ( .B1(npu_inst_pe_1_6_2_n61), .B2(
        npu_inst_pe_1_6_2_n52), .A(npu_inst_pe_1_6_2_n69), .ZN(
        npu_inst_pe_1_6_2_n92) );
  NAND2_X1 npu_inst_pe_1_6_2_U75 ( .A1(npu_inst_pe_1_6_2_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_6_2_n48), .ZN(npu_inst_pe_1_6_2_n68) );
  OAI21_X1 npu_inst_pe_1_6_2_U74 ( .B1(npu_inst_pe_1_6_2_n63), .B2(
        npu_inst_pe_1_6_2_n48), .A(npu_inst_pe_1_6_2_n68), .ZN(
        npu_inst_pe_1_6_2_n91) );
  NAND2_X1 npu_inst_pe_1_6_2_U73 ( .A1(npu_inst_pe_1_6_2_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_6_2_n48), .ZN(npu_inst_pe_1_6_2_n67) );
  OAI21_X1 npu_inst_pe_1_6_2_U72 ( .B1(npu_inst_pe_1_6_2_n61), .B2(
        npu_inst_pe_1_6_2_n48), .A(npu_inst_pe_1_6_2_n67), .ZN(
        npu_inst_pe_1_6_2_n90) );
  NAND2_X1 npu_inst_pe_1_6_2_U71 ( .A1(npu_inst_pe_1_6_2_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_6_2_n44), .ZN(npu_inst_pe_1_6_2_n66) );
  OAI21_X1 npu_inst_pe_1_6_2_U70 ( .B1(npu_inst_pe_1_6_2_n63), .B2(
        npu_inst_pe_1_6_2_n44), .A(npu_inst_pe_1_6_2_n66), .ZN(
        npu_inst_pe_1_6_2_n89) );
  NAND2_X1 npu_inst_pe_1_6_2_U69 ( .A1(npu_inst_pe_1_6_2_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_6_2_n44), .ZN(npu_inst_pe_1_6_2_n65) );
  OAI21_X1 npu_inst_pe_1_6_2_U68 ( .B1(npu_inst_pe_1_6_2_n61), .B2(
        npu_inst_pe_1_6_2_n44), .A(npu_inst_pe_1_6_2_n65), .ZN(
        npu_inst_pe_1_6_2_n88) );
  NAND2_X1 npu_inst_pe_1_6_2_U67 ( .A1(npu_inst_pe_1_6_2_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_6_2_n40), .ZN(npu_inst_pe_1_6_2_n64) );
  OAI21_X1 npu_inst_pe_1_6_2_U66 ( .B1(npu_inst_pe_1_6_2_n63), .B2(
        npu_inst_pe_1_6_2_n40), .A(npu_inst_pe_1_6_2_n64), .ZN(
        npu_inst_pe_1_6_2_n87) );
  NAND2_X1 npu_inst_pe_1_6_2_U65 ( .A1(npu_inst_pe_1_6_2_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_6_2_n40), .ZN(npu_inst_pe_1_6_2_n62) );
  OAI21_X1 npu_inst_pe_1_6_2_U64 ( .B1(npu_inst_pe_1_6_2_n61), .B2(
        npu_inst_pe_1_6_2_n40), .A(npu_inst_pe_1_6_2_n62), .ZN(
        npu_inst_pe_1_6_2_n86) );
  AND2_X1 npu_inst_pe_1_6_2_U63 ( .A1(npu_inst_pe_1_6_2_N93), .A2(npu_inst_n53), .ZN(npu_inst_int_data_y_6__2__0_) );
  AND2_X1 npu_inst_pe_1_6_2_U62 ( .A1(npu_inst_n53), .A2(npu_inst_pe_1_6_2_N94), .ZN(npu_inst_int_data_y_6__2__1_) );
  NOR3_X1 npu_inst_pe_1_6_2_U61 ( .A1(npu_inst_pe_1_6_2_n26), .A2(npu_inst_n53), .A3(npu_inst_int_ckg[13]), .ZN(npu_inst_pe_1_6_2_n85) );
  OR2_X1 npu_inst_pe_1_6_2_U60 ( .A1(npu_inst_pe_1_6_2_n85), .A2(
        npu_inst_pe_1_6_2_n2), .ZN(npu_inst_pe_1_6_2_N84) );
  AND2_X1 npu_inst_pe_1_6_2_U59 ( .A1(npu_inst_pe_1_6_2_int_q_acc_0_), .A2(
        npu_inst_pe_1_6_2_n1), .ZN(npu_inst_int_data_res_6__2__0_) );
  AND2_X1 npu_inst_pe_1_6_2_U58 ( .A1(npu_inst_pe_1_6_2_n2), .A2(
        npu_inst_pe_1_6_2_int_q_acc_7_), .ZN(npu_inst_int_data_res_6__2__7_)
         );
  AND2_X1 npu_inst_pe_1_6_2_U57 ( .A1(npu_inst_pe_1_6_2_int_q_acc_1_), .A2(
        npu_inst_pe_1_6_2_n1), .ZN(npu_inst_int_data_res_6__2__1_) );
  AND2_X1 npu_inst_pe_1_6_2_U56 ( .A1(npu_inst_pe_1_6_2_int_q_acc_2_), .A2(
        npu_inst_pe_1_6_2_n1), .ZN(npu_inst_int_data_res_6__2__2_) );
  AND2_X1 npu_inst_pe_1_6_2_U55 ( .A1(npu_inst_pe_1_6_2_int_q_acc_3_), .A2(
        npu_inst_pe_1_6_2_n2), .ZN(npu_inst_int_data_res_6__2__3_) );
  AND2_X1 npu_inst_pe_1_6_2_U54 ( .A1(npu_inst_pe_1_6_2_int_q_acc_4_), .A2(
        npu_inst_pe_1_6_2_n2), .ZN(npu_inst_int_data_res_6__2__4_) );
  AND2_X1 npu_inst_pe_1_6_2_U53 ( .A1(npu_inst_pe_1_6_2_int_q_acc_5_), .A2(
        npu_inst_pe_1_6_2_n2), .ZN(npu_inst_int_data_res_6__2__5_) );
  AND2_X1 npu_inst_pe_1_6_2_U52 ( .A1(npu_inst_pe_1_6_2_int_q_acc_6_), .A2(
        npu_inst_pe_1_6_2_n2), .ZN(npu_inst_int_data_res_6__2__6_) );
  AOI222_X1 npu_inst_pe_1_6_2_U51 ( .A1(npu_inst_int_data_res_7__2__0_), .A2(
        npu_inst_pe_1_6_2_n1), .B1(npu_inst_pe_1_6_2_N73), .B2(
        npu_inst_pe_1_6_2_n76), .C1(npu_inst_pe_1_6_2_N65), .C2(
        npu_inst_pe_1_6_2_n77), .ZN(npu_inst_pe_1_6_2_n84) );
  INV_X1 npu_inst_pe_1_6_2_U50 ( .A(npu_inst_pe_1_6_2_n84), .ZN(
        npu_inst_pe_1_6_2_n101) );
  AOI222_X1 npu_inst_pe_1_6_2_U49 ( .A1(npu_inst_int_data_res_7__2__7_), .A2(
        npu_inst_pe_1_6_2_n1), .B1(npu_inst_pe_1_6_2_N80), .B2(
        npu_inst_pe_1_6_2_n76), .C1(npu_inst_pe_1_6_2_N72), .C2(
        npu_inst_pe_1_6_2_n77), .ZN(npu_inst_pe_1_6_2_n75) );
  INV_X1 npu_inst_pe_1_6_2_U48 ( .A(npu_inst_pe_1_6_2_n75), .ZN(
        npu_inst_pe_1_6_2_n33) );
  AOI222_X1 npu_inst_pe_1_6_2_U47 ( .A1(npu_inst_int_data_res_7__2__1_), .A2(
        npu_inst_pe_1_6_2_n1), .B1(npu_inst_pe_1_6_2_N74), .B2(
        npu_inst_pe_1_6_2_n76), .C1(npu_inst_pe_1_6_2_N66), .C2(
        npu_inst_pe_1_6_2_n77), .ZN(npu_inst_pe_1_6_2_n83) );
  INV_X1 npu_inst_pe_1_6_2_U46 ( .A(npu_inst_pe_1_6_2_n83), .ZN(
        npu_inst_pe_1_6_2_n100) );
  AOI222_X1 npu_inst_pe_1_6_2_U45 ( .A1(npu_inst_int_data_res_7__2__2_), .A2(
        npu_inst_pe_1_6_2_n1), .B1(npu_inst_pe_1_6_2_N75), .B2(
        npu_inst_pe_1_6_2_n76), .C1(npu_inst_pe_1_6_2_N67), .C2(
        npu_inst_pe_1_6_2_n77), .ZN(npu_inst_pe_1_6_2_n82) );
  INV_X1 npu_inst_pe_1_6_2_U44 ( .A(npu_inst_pe_1_6_2_n82), .ZN(
        npu_inst_pe_1_6_2_n99) );
  AOI222_X1 npu_inst_pe_1_6_2_U43 ( .A1(npu_inst_int_data_res_7__2__3_), .A2(
        npu_inst_pe_1_6_2_n1), .B1(npu_inst_pe_1_6_2_N76), .B2(
        npu_inst_pe_1_6_2_n76), .C1(npu_inst_pe_1_6_2_N68), .C2(
        npu_inst_pe_1_6_2_n77), .ZN(npu_inst_pe_1_6_2_n81) );
  INV_X1 npu_inst_pe_1_6_2_U42 ( .A(npu_inst_pe_1_6_2_n81), .ZN(
        npu_inst_pe_1_6_2_n98) );
  AOI222_X1 npu_inst_pe_1_6_2_U41 ( .A1(npu_inst_int_data_res_7__2__4_), .A2(
        npu_inst_pe_1_6_2_n1), .B1(npu_inst_pe_1_6_2_N77), .B2(
        npu_inst_pe_1_6_2_n76), .C1(npu_inst_pe_1_6_2_N69), .C2(
        npu_inst_pe_1_6_2_n77), .ZN(npu_inst_pe_1_6_2_n80) );
  INV_X1 npu_inst_pe_1_6_2_U40 ( .A(npu_inst_pe_1_6_2_n80), .ZN(
        npu_inst_pe_1_6_2_n36) );
  AOI222_X1 npu_inst_pe_1_6_2_U39 ( .A1(npu_inst_int_data_res_7__2__5_), .A2(
        npu_inst_pe_1_6_2_n1), .B1(npu_inst_pe_1_6_2_N78), .B2(
        npu_inst_pe_1_6_2_n76), .C1(npu_inst_pe_1_6_2_N70), .C2(
        npu_inst_pe_1_6_2_n77), .ZN(npu_inst_pe_1_6_2_n79) );
  INV_X1 npu_inst_pe_1_6_2_U38 ( .A(npu_inst_pe_1_6_2_n79), .ZN(
        npu_inst_pe_1_6_2_n35) );
  AOI222_X1 npu_inst_pe_1_6_2_U37 ( .A1(npu_inst_int_data_res_7__2__6_), .A2(
        npu_inst_pe_1_6_2_n1), .B1(npu_inst_pe_1_6_2_N79), .B2(
        npu_inst_pe_1_6_2_n76), .C1(npu_inst_pe_1_6_2_N71), .C2(
        npu_inst_pe_1_6_2_n77), .ZN(npu_inst_pe_1_6_2_n78) );
  INV_X1 npu_inst_pe_1_6_2_U36 ( .A(npu_inst_pe_1_6_2_n78), .ZN(
        npu_inst_pe_1_6_2_n34) );
  INV_X1 npu_inst_pe_1_6_2_U35 ( .A(npu_inst_pe_1_6_2_int_data_1_), .ZN(
        npu_inst_pe_1_6_2_n14) );
  AND2_X1 npu_inst_pe_1_6_2_U34 ( .A1(npu_inst_int_data_x_6__2__1_), .A2(
        npu_inst_pe_1_6_2_int_q_weight_1_), .ZN(npu_inst_pe_1_6_2_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_6_2_U33 ( .A1(npu_inst_int_data_x_6__2__0_), .A2(
        npu_inst_pe_1_6_2_int_q_weight_1_), .ZN(npu_inst_pe_1_6_2_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_6_2_U32 ( .A1(npu_inst_n53), .A2(
        npu_inst_int_data_y_7__2__1_), .B1(npu_inst_pe_1_6_2_n3), .B2(
        npu_inst_int_data_x_6__3__1_), .ZN(npu_inst_pe_1_6_2_n63) );
  AOI22_X1 npu_inst_pe_1_6_2_U31 ( .A1(npu_inst_n53), .A2(
        npu_inst_int_data_y_7__2__0_), .B1(npu_inst_pe_1_6_2_n3), .B2(
        npu_inst_int_data_x_6__3__0_), .ZN(npu_inst_pe_1_6_2_n61) );
  INV_X1 npu_inst_pe_1_6_2_U30 ( .A(npu_inst_pe_1_6_2_int_data_0_), .ZN(
        npu_inst_pe_1_6_2_n13) );
  INV_X1 npu_inst_pe_1_6_2_U29 ( .A(npu_inst_n68), .ZN(npu_inst_pe_1_6_2_n5)
         );
  OR3_X1 npu_inst_pe_1_6_2_U28 ( .A1(npu_inst_pe_1_6_2_n6), .A2(
        npu_inst_pe_1_6_2_n8), .A3(npu_inst_pe_1_6_2_n5), .ZN(
        npu_inst_pe_1_6_2_n56) );
  OR3_X1 npu_inst_pe_1_6_2_U27 ( .A1(npu_inst_pe_1_6_2_n5), .A2(
        npu_inst_pe_1_6_2_n8), .A3(npu_inst_pe_1_6_2_n7), .ZN(
        npu_inst_pe_1_6_2_n48) );
  INV_X1 npu_inst_pe_1_6_2_U26 ( .A(npu_inst_pe_1_6_2_n5), .ZN(
        npu_inst_pe_1_6_2_n4) );
  INV_X1 npu_inst_pe_1_6_2_U25 ( .A(npu_inst_n123), .ZN(npu_inst_pe_1_6_2_n12)
         );
  OR3_X1 npu_inst_pe_1_6_2_U24 ( .A1(npu_inst_pe_1_6_2_n4), .A2(
        npu_inst_pe_1_6_2_n8), .A3(npu_inst_pe_1_6_2_n7), .ZN(
        npu_inst_pe_1_6_2_n52) );
  OR3_X1 npu_inst_pe_1_6_2_U23 ( .A1(npu_inst_pe_1_6_2_n6), .A2(
        npu_inst_pe_1_6_2_n8), .A3(npu_inst_pe_1_6_2_n4), .ZN(
        npu_inst_pe_1_6_2_n60) );
  NOR2_X1 npu_inst_pe_1_6_2_U22 ( .A1(npu_inst_pe_1_6_2_n60), .A2(
        npu_inst_pe_1_6_2_n3), .ZN(npu_inst_pe_1_6_2_n58) );
  NOR2_X1 npu_inst_pe_1_6_2_U21 ( .A1(npu_inst_pe_1_6_2_n56), .A2(
        npu_inst_pe_1_6_2_n3), .ZN(npu_inst_pe_1_6_2_n54) );
  NOR2_X1 npu_inst_pe_1_6_2_U20 ( .A1(npu_inst_pe_1_6_2_n52), .A2(
        npu_inst_pe_1_6_2_n3), .ZN(npu_inst_pe_1_6_2_n50) );
  NOR2_X1 npu_inst_pe_1_6_2_U19 ( .A1(npu_inst_pe_1_6_2_n48), .A2(
        npu_inst_pe_1_6_2_n3), .ZN(npu_inst_pe_1_6_2_n46) );
  NOR2_X1 npu_inst_pe_1_6_2_U18 ( .A1(npu_inst_pe_1_6_2_n40), .A2(
        npu_inst_pe_1_6_2_n3), .ZN(npu_inst_pe_1_6_2_n38) );
  NOR2_X1 npu_inst_pe_1_6_2_U17 ( .A1(npu_inst_pe_1_6_2_n44), .A2(
        npu_inst_pe_1_6_2_n3), .ZN(npu_inst_pe_1_6_2_n42) );
  BUF_X1 npu_inst_pe_1_6_2_U16 ( .A(npu_inst_n95), .Z(npu_inst_pe_1_6_2_n8) );
  BUF_X1 npu_inst_pe_1_6_2_U15 ( .A(npu_inst_pe_1_6_2_n12), .Z(
        npu_inst_pe_1_6_2_n11) );
  BUF_X1 npu_inst_pe_1_6_2_U14 ( .A(npu_inst_pe_1_6_2_n12), .Z(
        npu_inst_pe_1_6_2_n10) );
  BUF_X1 npu_inst_pe_1_6_2_U13 ( .A(npu_inst_pe_1_6_2_n12), .Z(
        npu_inst_pe_1_6_2_n9) );
  INV_X1 npu_inst_pe_1_6_2_U12 ( .A(npu_inst_pe_1_6_2_n38), .ZN(
        npu_inst_pe_1_6_2_n118) );
  INV_X1 npu_inst_pe_1_6_2_U11 ( .A(npu_inst_pe_1_6_2_n58), .ZN(
        npu_inst_pe_1_6_2_n114) );
  INV_X1 npu_inst_pe_1_6_2_U10 ( .A(npu_inst_pe_1_6_2_n54), .ZN(
        npu_inst_pe_1_6_2_n115) );
  INV_X1 npu_inst_pe_1_6_2_U9 ( .A(npu_inst_pe_1_6_2_n50), .ZN(
        npu_inst_pe_1_6_2_n116) );
  INV_X1 npu_inst_pe_1_6_2_U8 ( .A(npu_inst_pe_1_6_2_n46), .ZN(
        npu_inst_pe_1_6_2_n117) );
  INV_X1 npu_inst_pe_1_6_2_U7 ( .A(npu_inst_pe_1_6_2_n42), .ZN(
        npu_inst_pe_1_6_2_n119) );
  BUF_X1 npu_inst_pe_1_6_2_U6 ( .A(npu_inst_n13), .Z(npu_inst_pe_1_6_2_n2) );
  BUF_X1 npu_inst_pe_1_6_2_U5 ( .A(npu_inst_n13), .Z(npu_inst_pe_1_6_2_n1) );
  NOR2_X1 npu_inst_pe_1_6_2_U4 ( .A1(npu_inst_pe_1_6_2_int_q_weight_0_), .A2(
        npu_inst_pe_1_6_2_n1), .ZN(npu_inst_pe_1_6_2_n76) );
  NOR2_X1 npu_inst_pe_1_6_2_U3 ( .A1(npu_inst_pe_1_6_2_n27), .A2(
        npu_inst_pe_1_6_2_n1), .ZN(npu_inst_pe_1_6_2_n77) );
  FA_X1 npu_inst_pe_1_6_2_sub_77_U2_1 ( .A(npu_inst_pe_1_6_2_int_q_acc_1_), 
        .B(npu_inst_pe_1_6_2_n14), .CI(npu_inst_pe_1_6_2_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_6_2_sub_77_carry_2_), .S(npu_inst_pe_1_6_2_N66) );
  FA_X1 npu_inst_pe_1_6_2_add_79_U1_1 ( .A(npu_inst_pe_1_6_2_int_q_acc_1_), 
        .B(npu_inst_pe_1_6_2_int_data_1_), .CI(
        npu_inst_pe_1_6_2_add_79_carry_1_), .CO(
        npu_inst_pe_1_6_2_add_79_carry_2_), .S(npu_inst_pe_1_6_2_N74) );
  NAND3_X1 npu_inst_pe_1_6_2_U109 ( .A1(npu_inst_pe_1_6_2_n5), .A2(
        npu_inst_pe_1_6_2_n7), .A3(npu_inst_pe_1_6_2_n8), .ZN(
        npu_inst_pe_1_6_2_n44) );
  NAND3_X1 npu_inst_pe_1_6_2_U108 ( .A1(npu_inst_pe_1_6_2_n4), .A2(
        npu_inst_pe_1_6_2_n7), .A3(npu_inst_pe_1_6_2_n8), .ZN(
        npu_inst_pe_1_6_2_n40) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_6_2_n34), .CK(
        npu_inst_pe_1_6_2_net3143), .RN(npu_inst_pe_1_6_2_n9), .Q(
        npu_inst_pe_1_6_2_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_6_2_n35), .CK(
        npu_inst_pe_1_6_2_net3143), .RN(npu_inst_pe_1_6_2_n9), .Q(
        npu_inst_pe_1_6_2_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_6_2_n36), .CK(
        npu_inst_pe_1_6_2_net3143), .RN(npu_inst_pe_1_6_2_n9), .Q(
        npu_inst_pe_1_6_2_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_6_2_n98), .CK(
        npu_inst_pe_1_6_2_net3143), .RN(npu_inst_pe_1_6_2_n9), .Q(
        npu_inst_pe_1_6_2_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_6_2_n99), .CK(
        npu_inst_pe_1_6_2_net3143), .RN(npu_inst_pe_1_6_2_n9), .Q(
        npu_inst_pe_1_6_2_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_6_2_n100), 
        .CK(npu_inst_pe_1_6_2_net3143), .RN(npu_inst_pe_1_6_2_n9), .Q(
        npu_inst_pe_1_6_2_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_6_2_n33), .CK(
        npu_inst_pe_1_6_2_net3143), .RN(npu_inst_pe_1_6_2_n9), .Q(
        npu_inst_pe_1_6_2_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_6_2_n101), 
        .CK(npu_inst_pe_1_6_2_net3143), .RN(npu_inst_pe_1_6_2_n9), .Q(
        npu_inst_pe_1_6_2_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_weight_reg_0_ ( .D(npu_inst_n109), .CK(
        npu_inst_pe_1_6_2_net3149), .RN(npu_inst_pe_1_6_2_n9), .Q(
        npu_inst_pe_1_6_2_int_q_weight_0_), .QN(npu_inst_pe_1_6_2_n27) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_weight_reg_1_ ( .D(npu_inst_n115), .CK(
        npu_inst_pe_1_6_2_net3149), .RN(npu_inst_pe_1_6_2_n9), .Q(
        npu_inst_pe_1_6_2_int_q_weight_1_), .QN(npu_inst_pe_1_6_2_n26) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_6_2_n113), 
        .CK(npu_inst_pe_1_6_2_net3149), .RN(npu_inst_pe_1_6_2_n9), .Q(
        npu_inst_pe_1_6_2_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_6_2_n107), 
        .CK(npu_inst_pe_1_6_2_net3149), .RN(npu_inst_pe_1_6_2_n9), .Q(
        npu_inst_pe_1_6_2_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_6_2_n112), 
        .CK(npu_inst_pe_1_6_2_net3149), .RN(npu_inst_pe_1_6_2_n10), .Q(
        npu_inst_pe_1_6_2_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_6_2_n106), 
        .CK(npu_inst_pe_1_6_2_net3149), .RN(npu_inst_pe_1_6_2_n10), .Q(
        npu_inst_pe_1_6_2_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_6_2_n111), 
        .CK(npu_inst_pe_1_6_2_net3149), .RN(npu_inst_pe_1_6_2_n10), .Q(
        npu_inst_pe_1_6_2_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_6_2_n105), 
        .CK(npu_inst_pe_1_6_2_net3149), .RN(npu_inst_pe_1_6_2_n10), .Q(
        npu_inst_pe_1_6_2_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_6_2_n110), 
        .CK(npu_inst_pe_1_6_2_net3149), .RN(npu_inst_pe_1_6_2_n10), .Q(
        npu_inst_pe_1_6_2_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_6_2_n104), 
        .CK(npu_inst_pe_1_6_2_net3149), .RN(npu_inst_pe_1_6_2_n10), .Q(
        npu_inst_pe_1_6_2_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_6_2_n109), 
        .CK(npu_inst_pe_1_6_2_net3149), .RN(npu_inst_pe_1_6_2_n10), .Q(
        npu_inst_pe_1_6_2_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_6_2_n103), 
        .CK(npu_inst_pe_1_6_2_net3149), .RN(npu_inst_pe_1_6_2_n10), .Q(
        npu_inst_pe_1_6_2_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_6_2_n108), 
        .CK(npu_inst_pe_1_6_2_net3149), .RN(npu_inst_pe_1_6_2_n10), .Q(
        npu_inst_pe_1_6_2_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_6_2_n102), 
        .CK(npu_inst_pe_1_6_2_net3149), .RN(npu_inst_pe_1_6_2_n10), .Q(
        npu_inst_pe_1_6_2_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_6_2_n86), 
        .CK(npu_inst_pe_1_6_2_net3149), .RN(npu_inst_pe_1_6_2_n10), .Q(
        npu_inst_pe_1_6_2_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_6_2_n87), 
        .CK(npu_inst_pe_1_6_2_net3149), .RN(npu_inst_pe_1_6_2_n10), .Q(
        npu_inst_pe_1_6_2_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_6_2_n88), 
        .CK(npu_inst_pe_1_6_2_net3149), .RN(npu_inst_pe_1_6_2_n11), .Q(
        npu_inst_pe_1_6_2_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_6_2_n89), 
        .CK(npu_inst_pe_1_6_2_net3149), .RN(npu_inst_pe_1_6_2_n11), .Q(
        npu_inst_pe_1_6_2_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_6_2_n90), 
        .CK(npu_inst_pe_1_6_2_net3149), .RN(npu_inst_pe_1_6_2_n11), .Q(
        npu_inst_pe_1_6_2_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_6_2_n91), 
        .CK(npu_inst_pe_1_6_2_net3149), .RN(npu_inst_pe_1_6_2_n11), .Q(
        npu_inst_pe_1_6_2_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_6_2_n92), 
        .CK(npu_inst_pe_1_6_2_net3149), .RN(npu_inst_pe_1_6_2_n11), .Q(
        npu_inst_pe_1_6_2_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_6_2_n93), 
        .CK(npu_inst_pe_1_6_2_net3149), .RN(npu_inst_pe_1_6_2_n11), .Q(
        npu_inst_pe_1_6_2_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_6_2_n94), 
        .CK(npu_inst_pe_1_6_2_net3149), .RN(npu_inst_pe_1_6_2_n11), .Q(
        npu_inst_pe_1_6_2_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_6_2_n95), 
        .CK(npu_inst_pe_1_6_2_net3149), .RN(npu_inst_pe_1_6_2_n11), .Q(
        npu_inst_pe_1_6_2_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_6_2_n96), 
        .CK(npu_inst_pe_1_6_2_net3149), .RN(npu_inst_pe_1_6_2_n11), .Q(
        npu_inst_pe_1_6_2_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_6_2_n97), 
        .CK(npu_inst_pe_1_6_2_net3149), .RN(npu_inst_pe_1_6_2_n11), .Q(
        npu_inst_pe_1_6_2_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_6_2_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_6_2_N84), .SE(1'b0), .GCK(npu_inst_pe_1_6_2_net3143) );
  CLKGATETST_X1 npu_inst_pe_1_6_2_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n62), .SE(1'b0), .GCK(npu_inst_pe_1_6_2_net3149) );
  MUX2_X1 npu_inst_pe_1_6_3_U162 ( .A(npu_inst_pe_1_6_3_n32), .B(
        npu_inst_pe_1_6_3_n29), .S(npu_inst_pe_1_6_3_n8), .Z(
        npu_inst_pe_1_6_3_N93) );
  MUX2_X1 npu_inst_pe_1_6_3_U161 ( .A(npu_inst_pe_1_6_3_n31), .B(
        npu_inst_pe_1_6_3_n30), .S(npu_inst_pe_1_6_3_n6), .Z(
        npu_inst_pe_1_6_3_n32) );
  MUX2_X1 npu_inst_pe_1_6_3_U160 ( .A(npu_inst_pe_1_6_3_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_6_3_int_q_reg_v_1__0_), .S(npu_inst_pe_1_6_3_n4), .Z(
        npu_inst_pe_1_6_3_n31) );
  MUX2_X1 npu_inst_pe_1_6_3_U159 ( .A(npu_inst_pe_1_6_3_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_6_3_int_q_reg_v_3__0_), .S(npu_inst_pe_1_6_3_n4), .Z(
        npu_inst_pe_1_6_3_n30) );
  MUX2_X1 npu_inst_pe_1_6_3_U158 ( .A(npu_inst_pe_1_6_3_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_6_3_int_q_reg_v_5__0_), .S(npu_inst_pe_1_6_3_n4), .Z(
        npu_inst_pe_1_6_3_n29) );
  MUX2_X1 npu_inst_pe_1_6_3_U157 ( .A(npu_inst_pe_1_6_3_n28), .B(
        npu_inst_pe_1_6_3_n23), .S(npu_inst_pe_1_6_3_n8), .Z(
        npu_inst_pe_1_6_3_N94) );
  MUX2_X1 npu_inst_pe_1_6_3_U156 ( .A(npu_inst_pe_1_6_3_n25), .B(
        npu_inst_pe_1_6_3_n24), .S(npu_inst_pe_1_6_3_n6), .Z(
        npu_inst_pe_1_6_3_n28) );
  MUX2_X1 npu_inst_pe_1_6_3_U155 ( .A(npu_inst_pe_1_6_3_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_6_3_int_q_reg_v_1__1_), .S(npu_inst_pe_1_6_3_n4), .Z(
        npu_inst_pe_1_6_3_n25) );
  MUX2_X1 npu_inst_pe_1_6_3_U154 ( .A(npu_inst_pe_1_6_3_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_6_3_int_q_reg_v_3__1_), .S(npu_inst_pe_1_6_3_n4), .Z(
        npu_inst_pe_1_6_3_n24) );
  MUX2_X1 npu_inst_pe_1_6_3_U153 ( .A(npu_inst_pe_1_6_3_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_6_3_int_q_reg_v_5__1_), .S(npu_inst_pe_1_6_3_n4), .Z(
        npu_inst_pe_1_6_3_n23) );
  MUX2_X1 npu_inst_pe_1_6_3_U152 ( .A(npu_inst_pe_1_6_3_n22), .B(
        npu_inst_pe_1_6_3_n19), .S(npu_inst_pe_1_6_3_n8), .Z(
        npu_inst_int_data_x_6__3__1_) );
  MUX2_X1 npu_inst_pe_1_6_3_U151 ( .A(npu_inst_pe_1_6_3_n21), .B(
        npu_inst_pe_1_6_3_n20), .S(npu_inst_pe_1_6_3_n6), .Z(
        npu_inst_pe_1_6_3_n22) );
  MUX2_X1 npu_inst_pe_1_6_3_U150 ( .A(npu_inst_pe_1_6_3_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_6_3_int_q_reg_h_1__1_), .S(npu_inst_pe_1_6_3_n4), .Z(
        npu_inst_pe_1_6_3_n21) );
  MUX2_X1 npu_inst_pe_1_6_3_U149 ( .A(npu_inst_pe_1_6_3_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_6_3_int_q_reg_h_3__1_), .S(npu_inst_pe_1_6_3_n4), .Z(
        npu_inst_pe_1_6_3_n20) );
  MUX2_X1 npu_inst_pe_1_6_3_U148 ( .A(npu_inst_pe_1_6_3_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_6_3_int_q_reg_h_5__1_), .S(npu_inst_pe_1_6_3_n4), .Z(
        npu_inst_pe_1_6_3_n19) );
  MUX2_X1 npu_inst_pe_1_6_3_U147 ( .A(npu_inst_pe_1_6_3_n18), .B(
        npu_inst_pe_1_6_3_n15), .S(npu_inst_pe_1_6_3_n8), .Z(
        npu_inst_int_data_x_6__3__0_) );
  MUX2_X1 npu_inst_pe_1_6_3_U146 ( .A(npu_inst_pe_1_6_3_n17), .B(
        npu_inst_pe_1_6_3_n16), .S(npu_inst_pe_1_6_3_n6), .Z(
        npu_inst_pe_1_6_3_n18) );
  MUX2_X1 npu_inst_pe_1_6_3_U145 ( .A(npu_inst_pe_1_6_3_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_6_3_int_q_reg_h_1__0_), .S(npu_inst_pe_1_6_3_n4), .Z(
        npu_inst_pe_1_6_3_n17) );
  MUX2_X1 npu_inst_pe_1_6_3_U144 ( .A(npu_inst_pe_1_6_3_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_6_3_int_q_reg_h_3__0_), .S(npu_inst_pe_1_6_3_n4), .Z(
        npu_inst_pe_1_6_3_n16) );
  MUX2_X1 npu_inst_pe_1_6_3_U143 ( .A(npu_inst_pe_1_6_3_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_6_3_int_q_reg_h_5__0_), .S(npu_inst_pe_1_6_3_n4), .Z(
        npu_inst_pe_1_6_3_n15) );
  XOR2_X1 npu_inst_pe_1_6_3_U142 ( .A(npu_inst_pe_1_6_3_int_data_0_), .B(
        npu_inst_pe_1_6_3_int_q_acc_0_), .Z(npu_inst_pe_1_6_3_N73) );
  AND2_X1 npu_inst_pe_1_6_3_U141 ( .A1(npu_inst_pe_1_6_3_int_q_acc_0_), .A2(
        npu_inst_pe_1_6_3_int_data_0_), .ZN(npu_inst_pe_1_6_3_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_6_3_U140 ( .A(npu_inst_pe_1_6_3_int_q_acc_0_), .B(
        npu_inst_pe_1_6_3_n13), .ZN(npu_inst_pe_1_6_3_N65) );
  OR2_X1 npu_inst_pe_1_6_3_U139 ( .A1(npu_inst_pe_1_6_3_n13), .A2(
        npu_inst_pe_1_6_3_int_q_acc_0_), .ZN(npu_inst_pe_1_6_3_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_6_3_U138 ( .A(npu_inst_pe_1_6_3_int_q_acc_2_), .B(
        npu_inst_pe_1_6_3_add_79_carry_2_), .Z(npu_inst_pe_1_6_3_N75) );
  AND2_X1 npu_inst_pe_1_6_3_U137 ( .A1(npu_inst_pe_1_6_3_add_79_carry_2_), 
        .A2(npu_inst_pe_1_6_3_int_q_acc_2_), .ZN(
        npu_inst_pe_1_6_3_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_6_3_U136 ( .A(npu_inst_pe_1_6_3_int_q_acc_3_), .B(
        npu_inst_pe_1_6_3_add_79_carry_3_), .Z(npu_inst_pe_1_6_3_N76) );
  AND2_X1 npu_inst_pe_1_6_3_U135 ( .A1(npu_inst_pe_1_6_3_add_79_carry_3_), 
        .A2(npu_inst_pe_1_6_3_int_q_acc_3_), .ZN(
        npu_inst_pe_1_6_3_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_6_3_U134 ( .A(npu_inst_pe_1_6_3_int_q_acc_4_), .B(
        npu_inst_pe_1_6_3_add_79_carry_4_), .Z(npu_inst_pe_1_6_3_N77) );
  AND2_X1 npu_inst_pe_1_6_3_U133 ( .A1(npu_inst_pe_1_6_3_add_79_carry_4_), 
        .A2(npu_inst_pe_1_6_3_int_q_acc_4_), .ZN(
        npu_inst_pe_1_6_3_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_6_3_U132 ( .A(npu_inst_pe_1_6_3_int_q_acc_5_), .B(
        npu_inst_pe_1_6_3_add_79_carry_5_), .Z(npu_inst_pe_1_6_3_N78) );
  AND2_X1 npu_inst_pe_1_6_3_U131 ( .A1(npu_inst_pe_1_6_3_add_79_carry_5_), 
        .A2(npu_inst_pe_1_6_3_int_q_acc_5_), .ZN(
        npu_inst_pe_1_6_3_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_6_3_U130 ( .A(npu_inst_pe_1_6_3_int_q_acc_6_), .B(
        npu_inst_pe_1_6_3_add_79_carry_6_), .Z(npu_inst_pe_1_6_3_N79) );
  AND2_X1 npu_inst_pe_1_6_3_U129 ( .A1(npu_inst_pe_1_6_3_add_79_carry_6_), 
        .A2(npu_inst_pe_1_6_3_int_q_acc_6_), .ZN(
        npu_inst_pe_1_6_3_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_6_3_U128 ( .A(npu_inst_pe_1_6_3_int_q_acc_7_), .B(
        npu_inst_pe_1_6_3_add_79_carry_7_), .Z(npu_inst_pe_1_6_3_N80) );
  XNOR2_X1 npu_inst_pe_1_6_3_U127 ( .A(npu_inst_pe_1_6_3_sub_77_carry_2_), .B(
        npu_inst_pe_1_6_3_int_q_acc_2_), .ZN(npu_inst_pe_1_6_3_N67) );
  OR2_X1 npu_inst_pe_1_6_3_U126 ( .A1(npu_inst_pe_1_6_3_int_q_acc_2_), .A2(
        npu_inst_pe_1_6_3_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_6_3_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_6_3_U125 ( .A(npu_inst_pe_1_6_3_sub_77_carry_3_), .B(
        npu_inst_pe_1_6_3_int_q_acc_3_), .ZN(npu_inst_pe_1_6_3_N68) );
  OR2_X1 npu_inst_pe_1_6_3_U124 ( .A1(npu_inst_pe_1_6_3_int_q_acc_3_), .A2(
        npu_inst_pe_1_6_3_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_6_3_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_6_3_U123 ( .A(npu_inst_pe_1_6_3_sub_77_carry_4_), .B(
        npu_inst_pe_1_6_3_int_q_acc_4_), .ZN(npu_inst_pe_1_6_3_N69) );
  OR2_X1 npu_inst_pe_1_6_3_U122 ( .A1(npu_inst_pe_1_6_3_int_q_acc_4_), .A2(
        npu_inst_pe_1_6_3_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_6_3_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_6_3_U121 ( .A(npu_inst_pe_1_6_3_sub_77_carry_5_), .B(
        npu_inst_pe_1_6_3_int_q_acc_5_), .ZN(npu_inst_pe_1_6_3_N70) );
  OR2_X1 npu_inst_pe_1_6_3_U120 ( .A1(npu_inst_pe_1_6_3_int_q_acc_5_), .A2(
        npu_inst_pe_1_6_3_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_6_3_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_6_3_U119 ( .A(npu_inst_pe_1_6_3_sub_77_carry_6_), .B(
        npu_inst_pe_1_6_3_int_q_acc_6_), .ZN(npu_inst_pe_1_6_3_N71) );
  OR2_X1 npu_inst_pe_1_6_3_U118 ( .A1(npu_inst_pe_1_6_3_int_q_acc_6_), .A2(
        npu_inst_pe_1_6_3_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_6_3_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_6_3_U117 ( .A(npu_inst_pe_1_6_3_int_q_acc_7_), .B(
        npu_inst_pe_1_6_3_sub_77_carry_7_), .ZN(npu_inst_pe_1_6_3_N72) );
  INV_X1 npu_inst_pe_1_6_3_U116 ( .A(npu_inst_n76), .ZN(npu_inst_pe_1_6_3_n7)
         );
  INV_X1 npu_inst_pe_1_6_3_U115 ( .A(npu_inst_pe_1_6_3_n7), .ZN(
        npu_inst_pe_1_6_3_n6) );
  INV_X1 npu_inst_pe_1_6_3_U114 ( .A(npu_inst_n53), .ZN(npu_inst_pe_1_6_3_n3)
         );
  AOI22_X1 npu_inst_pe_1_6_3_U113 ( .A1(npu_inst_int_data_y_7__3__0_), .A2(
        npu_inst_pe_1_6_3_n58), .B1(npu_inst_pe_1_6_3_n114), .B2(
        npu_inst_pe_1_6_3_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_6_3_n57) );
  INV_X1 npu_inst_pe_1_6_3_U112 ( .A(npu_inst_pe_1_6_3_n57), .ZN(
        npu_inst_pe_1_6_3_n108) );
  AOI22_X1 npu_inst_pe_1_6_3_U111 ( .A1(npu_inst_int_data_y_7__3__0_), .A2(
        npu_inst_pe_1_6_3_n54), .B1(npu_inst_pe_1_6_3_n115), .B2(
        npu_inst_pe_1_6_3_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_6_3_n53) );
  INV_X1 npu_inst_pe_1_6_3_U110 ( .A(npu_inst_pe_1_6_3_n53), .ZN(
        npu_inst_pe_1_6_3_n109) );
  AOI22_X1 npu_inst_pe_1_6_3_U107 ( .A1(npu_inst_int_data_y_7__3__0_), .A2(
        npu_inst_pe_1_6_3_n50), .B1(npu_inst_pe_1_6_3_n116), .B2(
        npu_inst_pe_1_6_3_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_6_3_n49) );
  INV_X1 npu_inst_pe_1_6_3_U106 ( .A(npu_inst_pe_1_6_3_n49), .ZN(
        npu_inst_pe_1_6_3_n110) );
  AOI22_X1 npu_inst_pe_1_6_3_U105 ( .A1(npu_inst_int_data_y_7__3__0_), .A2(
        npu_inst_pe_1_6_3_n46), .B1(npu_inst_pe_1_6_3_n117), .B2(
        npu_inst_pe_1_6_3_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_6_3_n45) );
  INV_X1 npu_inst_pe_1_6_3_U104 ( .A(npu_inst_pe_1_6_3_n45), .ZN(
        npu_inst_pe_1_6_3_n111) );
  AOI22_X1 npu_inst_pe_1_6_3_U103 ( .A1(npu_inst_int_data_y_7__3__0_), .A2(
        npu_inst_pe_1_6_3_n42), .B1(npu_inst_pe_1_6_3_n119), .B2(
        npu_inst_pe_1_6_3_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_6_3_n41) );
  INV_X1 npu_inst_pe_1_6_3_U102 ( .A(npu_inst_pe_1_6_3_n41), .ZN(
        npu_inst_pe_1_6_3_n112) );
  AOI22_X1 npu_inst_pe_1_6_3_U101 ( .A1(npu_inst_int_data_y_7__3__1_), .A2(
        npu_inst_pe_1_6_3_n58), .B1(npu_inst_pe_1_6_3_n114), .B2(
        npu_inst_pe_1_6_3_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_6_3_n59) );
  INV_X1 npu_inst_pe_1_6_3_U100 ( .A(npu_inst_pe_1_6_3_n59), .ZN(
        npu_inst_pe_1_6_3_n102) );
  AOI22_X1 npu_inst_pe_1_6_3_U99 ( .A1(npu_inst_int_data_y_7__3__1_), .A2(
        npu_inst_pe_1_6_3_n54), .B1(npu_inst_pe_1_6_3_n115), .B2(
        npu_inst_pe_1_6_3_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_6_3_n55) );
  INV_X1 npu_inst_pe_1_6_3_U98 ( .A(npu_inst_pe_1_6_3_n55), .ZN(
        npu_inst_pe_1_6_3_n103) );
  AOI22_X1 npu_inst_pe_1_6_3_U97 ( .A1(npu_inst_int_data_y_7__3__1_), .A2(
        npu_inst_pe_1_6_3_n50), .B1(npu_inst_pe_1_6_3_n116), .B2(
        npu_inst_pe_1_6_3_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_6_3_n51) );
  INV_X1 npu_inst_pe_1_6_3_U96 ( .A(npu_inst_pe_1_6_3_n51), .ZN(
        npu_inst_pe_1_6_3_n104) );
  AOI22_X1 npu_inst_pe_1_6_3_U95 ( .A1(npu_inst_int_data_y_7__3__1_), .A2(
        npu_inst_pe_1_6_3_n46), .B1(npu_inst_pe_1_6_3_n117), .B2(
        npu_inst_pe_1_6_3_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_6_3_n47) );
  INV_X1 npu_inst_pe_1_6_3_U94 ( .A(npu_inst_pe_1_6_3_n47), .ZN(
        npu_inst_pe_1_6_3_n105) );
  AOI22_X1 npu_inst_pe_1_6_3_U93 ( .A1(npu_inst_int_data_y_7__3__1_), .A2(
        npu_inst_pe_1_6_3_n42), .B1(npu_inst_pe_1_6_3_n119), .B2(
        npu_inst_pe_1_6_3_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_6_3_n43) );
  INV_X1 npu_inst_pe_1_6_3_U92 ( .A(npu_inst_pe_1_6_3_n43), .ZN(
        npu_inst_pe_1_6_3_n106) );
  AOI22_X1 npu_inst_pe_1_6_3_U91 ( .A1(npu_inst_pe_1_6_3_n38), .A2(
        npu_inst_int_data_y_7__3__1_), .B1(npu_inst_pe_1_6_3_n118), .B2(
        npu_inst_pe_1_6_3_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_6_3_n39) );
  INV_X1 npu_inst_pe_1_6_3_U90 ( .A(npu_inst_pe_1_6_3_n39), .ZN(
        npu_inst_pe_1_6_3_n107) );
  AOI22_X1 npu_inst_pe_1_6_3_U89 ( .A1(npu_inst_pe_1_6_3_n38), .A2(
        npu_inst_int_data_y_7__3__0_), .B1(npu_inst_pe_1_6_3_n118), .B2(
        npu_inst_pe_1_6_3_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_6_3_n37) );
  INV_X1 npu_inst_pe_1_6_3_U88 ( .A(npu_inst_pe_1_6_3_n37), .ZN(
        npu_inst_pe_1_6_3_n113) );
  NAND2_X1 npu_inst_pe_1_6_3_U87 ( .A1(npu_inst_pe_1_6_3_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_6_3_n60), .ZN(npu_inst_pe_1_6_3_n74) );
  OAI21_X1 npu_inst_pe_1_6_3_U86 ( .B1(npu_inst_pe_1_6_3_n63), .B2(
        npu_inst_pe_1_6_3_n60), .A(npu_inst_pe_1_6_3_n74), .ZN(
        npu_inst_pe_1_6_3_n97) );
  NAND2_X1 npu_inst_pe_1_6_3_U85 ( .A1(npu_inst_pe_1_6_3_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_6_3_n60), .ZN(npu_inst_pe_1_6_3_n73) );
  OAI21_X1 npu_inst_pe_1_6_3_U84 ( .B1(npu_inst_pe_1_6_3_n61), .B2(
        npu_inst_pe_1_6_3_n60), .A(npu_inst_pe_1_6_3_n73), .ZN(
        npu_inst_pe_1_6_3_n96) );
  NAND2_X1 npu_inst_pe_1_6_3_U83 ( .A1(npu_inst_pe_1_6_3_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_6_3_n56), .ZN(npu_inst_pe_1_6_3_n72) );
  OAI21_X1 npu_inst_pe_1_6_3_U82 ( .B1(npu_inst_pe_1_6_3_n63), .B2(
        npu_inst_pe_1_6_3_n56), .A(npu_inst_pe_1_6_3_n72), .ZN(
        npu_inst_pe_1_6_3_n95) );
  NAND2_X1 npu_inst_pe_1_6_3_U81 ( .A1(npu_inst_pe_1_6_3_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_6_3_n56), .ZN(npu_inst_pe_1_6_3_n71) );
  OAI21_X1 npu_inst_pe_1_6_3_U80 ( .B1(npu_inst_pe_1_6_3_n61), .B2(
        npu_inst_pe_1_6_3_n56), .A(npu_inst_pe_1_6_3_n71), .ZN(
        npu_inst_pe_1_6_3_n94) );
  NAND2_X1 npu_inst_pe_1_6_3_U79 ( .A1(npu_inst_pe_1_6_3_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_6_3_n52), .ZN(npu_inst_pe_1_6_3_n70) );
  OAI21_X1 npu_inst_pe_1_6_3_U78 ( .B1(npu_inst_pe_1_6_3_n63), .B2(
        npu_inst_pe_1_6_3_n52), .A(npu_inst_pe_1_6_3_n70), .ZN(
        npu_inst_pe_1_6_3_n93) );
  NAND2_X1 npu_inst_pe_1_6_3_U77 ( .A1(npu_inst_pe_1_6_3_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_6_3_n52), .ZN(npu_inst_pe_1_6_3_n69) );
  OAI21_X1 npu_inst_pe_1_6_3_U76 ( .B1(npu_inst_pe_1_6_3_n61), .B2(
        npu_inst_pe_1_6_3_n52), .A(npu_inst_pe_1_6_3_n69), .ZN(
        npu_inst_pe_1_6_3_n92) );
  NAND2_X1 npu_inst_pe_1_6_3_U75 ( .A1(npu_inst_pe_1_6_3_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_6_3_n48), .ZN(npu_inst_pe_1_6_3_n68) );
  OAI21_X1 npu_inst_pe_1_6_3_U74 ( .B1(npu_inst_pe_1_6_3_n63), .B2(
        npu_inst_pe_1_6_3_n48), .A(npu_inst_pe_1_6_3_n68), .ZN(
        npu_inst_pe_1_6_3_n91) );
  NAND2_X1 npu_inst_pe_1_6_3_U73 ( .A1(npu_inst_pe_1_6_3_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_6_3_n48), .ZN(npu_inst_pe_1_6_3_n67) );
  OAI21_X1 npu_inst_pe_1_6_3_U72 ( .B1(npu_inst_pe_1_6_3_n61), .B2(
        npu_inst_pe_1_6_3_n48), .A(npu_inst_pe_1_6_3_n67), .ZN(
        npu_inst_pe_1_6_3_n90) );
  NAND2_X1 npu_inst_pe_1_6_3_U71 ( .A1(npu_inst_pe_1_6_3_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_6_3_n44), .ZN(npu_inst_pe_1_6_3_n66) );
  OAI21_X1 npu_inst_pe_1_6_3_U70 ( .B1(npu_inst_pe_1_6_3_n63), .B2(
        npu_inst_pe_1_6_3_n44), .A(npu_inst_pe_1_6_3_n66), .ZN(
        npu_inst_pe_1_6_3_n89) );
  NAND2_X1 npu_inst_pe_1_6_3_U69 ( .A1(npu_inst_pe_1_6_3_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_6_3_n44), .ZN(npu_inst_pe_1_6_3_n65) );
  OAI21_X1 npu_inst_pe_1_6_3_U68 ( .B1(npu_inst_pe_1_6_3_n61), .B2(
        npu_inst_pe_1_6_3_n44), .A(npu_inst_pe_1_6_3_n65), .ZN(
        npu_inst_pe_1_6_3_n88) );
  NAND2_X1 npu_inst_pe_1_6_3_U67 ( .A1(npu_inst_pe_1_6_3_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_6_3_n40), .ZN(npu_inst_pe_1_6_3_n64) );
  OAI21_X1 npu_inst_pe_1_6_3_U66 ( .B1(npu_inst_pe_1_6_3_n63), .B2(
        npu_inst_pe_1_6_3_n40), .A(npu_inst_pe_1_6_3_n64), .ZN(
        npu_inst_pe_1_6_3_n87) );
  NAND2_X1 npu_inst_pe_1_6_3_U65 ( .A1(npu_inst_pe_1_6_3_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_6_3_n40), .ZN(npu_inst_pe_1_6_3_n62) );
  OAI21_X1 npu_inst_pe_1_6_3_U64 ( .B1(npu_inst_pe_1_6_3_n61), .B2(
        npu_inst_pe_1_6_3_n40), .A(npu_inst_pe_1_6_3_n62), .ZN(
        npu_inst_pe_1_6_3_n86) );
  AND2_X1 npu_inst_pe_1_6_3_U63 ( .A1(npu_inst_pe_1_6_3_N93), .A2(npu_inst_n53), .ZN(npu_inst_int_data_y_6__3__0_) );
  AND2_X1 npu_inst_pe_1_6_3_U62 ( .A1(npu_inst_n53), .A2(npu_inst_pe_1_6_3_N94), .ZN(npu_inst_int_data_y_6__3__1_) );
  NOR3_X1 npu_inst_pe_1_6_3_U61 ( .A1(npu_inst_pe_1_6_3_n26), .A2(npu_inst_n53), .A3(npu_inst_int_ckg[12]), .ZN(npu_inst_pe_1_6_3_n85) );
  OR2_X1 npu_inst_pe_1_6_3_U60 ( .A1(npu_inst_pe_1_6_3_n85), .A2(
        npu_inst_pe_1_6_3_n2), .ZN(npu_inst_pe_1_6_3_N84) );
  AND2_X1 npu_inst_pe_1_6_3_U59 ( .A1(npu_inst_pe_1_6_3_int_q_acc_0_), .A2(
        npu_inst_pe_1_6_3_n1), .ZN(npu_inst_int_data_res_6__3__0_) );
  AND2_X1 npu_inst_pe_1_6_3_U58 ( .A1(npu_inst_pe_1_6_3_n2), .A2(
        npu_inst_pe_1_6_3_int_q_acc_7_), .ZN(npu_inst_int_data_res_6__3__7_)
         );
  AND2_X1 npu_inst_pe_1_6_3_U57 ( .A1(npu_inst_pe_1_6_3_int_q_acc_1_), .A2(
        npu_inst_pe_1_6_3_n1), .ZN(npu_inst_int_data_res_6__3__1_) );
  AND2_X1 npu_inst_pe_1_6_3_U56 ( .A1(npu_inst_pe_1_6_3_int_q_acc_2_), .A2(
        npu_inst_pe_1_6_3_n1), .ZN(npu_inst_int_data_res_6__3__2_) );
  AND2_X1 npu_inst_pe_1_6_3_U55 ( .A1(npu_inst_pe_1_6_3_int_q_acc_3_), .A2(
        npu_inst_pe_1_6_3_n2), .ZN(npu_inst_int_data_res_6__3__3_) );
  AND2_X1 npu_inst_pe_1_6_3_U54 ( .A1(npu_inst_pe_1_6_3_int_q_acc_4_), .A2(
        npu_inst_pe_1_6_3_n2), .ZN(npu_inst_int_data_res_6__3__4_) );
  AND2_X1 npu_inst_pe_1_6_3_U53 ( .A1(npu_inst_pe_1_6_3_int_q_acc_5_), .A2(
        npu_inst_pe_1_6_3_n2), .ZN(npu_inst_int_data_res_6__3__5_) );
  AND2_X1 npu_inst_pe_1_6_3_U52 ( .A1(npu_inst_pe_1_6_3_int_q_acc_6_), .A2(
        npu_inst_pe_1_6_3_n2), .ZN(npu_inst_int_data_res_6__3__6_) );
  AOI222_X1 npu_inst_pe_1_6_3_U51 ( .A1(npu_inst_int_data_res_7__3__0_), .A2(
        npu_inst_pe_1_6_3_n1), .B1(npu_inst_pe_1_6_3_N73), .B2(
        npu_inst_pe_1_6_3_n76), .C1(npu_inst_pe_1_6_3_N65), .C2(
        npu_inst_pe_1_6_3_n77), .ZN(npu_inst_pe_1_6_3_n84) );
  INV_X1 npu_inst_pe_1_6_3_U50 ( .A(npu_inst_pe_1_6_3_n84), .ZN(
        npu_inst_pe_1_6_3_n101) );
  AOI222_X1 npu_inst_pe_1_6_3_U49 ( .A1(npu_inst_int_data_res_7__3__7_), .A2(
        npu_inst_pe_1_6_3_n1), .B1(npu_inst_pe_1_6_3_N80), .B2(
        npu_inst_pe_1_6_3_n76), .C1(npu_inst_pe_1_6_3_N72), .C2(
        npu_inst_pe_1_6_3_n77), .ZN(npu_inst_pe_1_6_3_n75) );
  INV_X1 npu_inst_pe_1_6_3_U48 ( .A(npu_inst_pe_1_6_3_n75), .ZN(
        npu_inst_pe_1_6_3_n33) );
  AOI222_X1 npu_inst_pe_1_6_3_U47 ( .A1(npu_inst_int_data_res_7__3__1_), .A2(
        npu_inst_pe_1_6_3_n1), .B1(npu_inst_pe_1_6_3_N74), .B2(
        npu_inst_pe_1_6_3_n76), .C1(npu_inst_pe_1_6_3_N66), .C2(
        npu_inst_pe_1_6_3_n77), .ZN(npu_inst_pe_1_6_3_n83) );
  INV_X1 npu_inst_pe_1_6_3_U46 ( .A(npu_inst_pe_1_6_3_n83), .ZN(
        npu_inst_pe_1_6_3_n100) );
  AOI222_X1 npu_inst_pe_1_6_3_U45 ( .A1(npu_inst_int_data_res_7__3__2_), .A2(
        npu_inst_pe_1_6_3_n1), .B1(npu_inst_pe_1_6_3_N75), .B2(
        npu_inst_pe_1_6_3_n76), .C1(npu_inst_pe_1_6_3_N67), .C2(
        npu_inst_pe_1_6_3_n77), .ZN(npu_inst_pe_1_6_3_n82) );
  INV_X1 npu_inst_pe_1_6_3_U44 ( .A(npu_inst_pe_1_6_3_n82), .ZN(
        npu_inst_pe_1_6_3_n99) );
  AOI222_X1 npu_inst_pe_1_6_3_U43 ( .A1(npu_inst_int_data_res_7__3__3_), .A2(
        npu_inst_pe_1_6_3_n1), .B1(npu_inst_pe_1_6_3_N76), .B2(
        npu_inst_pe_1_6_3_n76), .C1(npu_inst_pe_1_6_3_N68), .C2(
        npu_inst_pe_1_6_3_n77), .ZN(npu_inst_pe_1_6_3_n81) );
  INV_X1 npu_inst_pe_1_6_3_U42 ( .A(npu_inst_pe_1_6_3_n81), .ZN(
        npu_inst_pe_1_6_3_n98) );
  AOI222_X1 npu_inst_pe_1_6_3_U41 ( .A1(npu_inst_int_data_res_7__3__4_), .A2(
        npu_inst_pe_1_6_3_n1), .B1(npu_inst_pe_1_6_3_N77), .B2(
        npu_inst_pe_1_6_3_n76), .C1(npu_inst_pe_1_6_3_N69), .C2(
        npu_inst_pe_1_6_3_n77), .ZN(npu_inst_pe_1_6_3_n80) );
  INV_X1 npu_inst_pe_1_6_3_U40 ( .A(npu_inst_pe_1_6_3_n80), .ZN(
        npu_inst_pe_1_6_3_n36) );
  AOI222_X1 npu_inst_pe_1_6_3_U39 ( .A1(npu_inst_int_data_res_7__3__5_), .A2(
        npu_inst_pe_1_6_3_n1), .B1(npu_inst_pe_1_6_3_N78), .B2(
        npu_inst_pe_1_6_3_n76), .C1(npu_inst_pe_1_6_3_N70), .C2(
        npu_inst_pe_1_6_3_n77), .ZN(npu_inst_pe_1_6_3_n79) );
  INV_X1 npu_inst_pe_1_6_3_U38 ( .A(npu_inst_pe_1_6_3_n79), .ZN(
        npu_inst_pe_1_6_3_n35) );
  AOI222_X1 npu_inst_pe_1_6_3_U37 ( .A1(npu_inst_int_data_res_7__3__6_), .A2(
        npu_inst_pe_1_6_3_n1), .B1(npu_inst_pe_1_6_3_N79), .B2(
        npu_inst_pe_1_6_3_n76), .C1(npu_inst_pe_1_6_3_N71), .C2(
        npu_inst_pe_1_6_3_n77), .ZN(npu_inst_pe_1_6_3_n78) );
  INV_X1 npu_inst_pe_1_6_3_U36 ( .A(npu_inst_pe_1_6_3_n78), .ZN(
        npu_inst_pe_1_6_3_n34) );
  INV_X1 npu_inst_pe_1_6_3_U35 ( .A(npu_inst_pe_1_6_3_int_data_1_), .ZN(
        npu_inst_pe_1_6_3_n14) );
  AND2_X1 npu_inst_pe_1_6_3_U34 ( .A1(npu_inst_int_data_x_6__3__1_), .A2(
        npu_inst_pe_1_6_3_int_q_weight_1_), .ZN(npu_inst_pe_1_6_3_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_6_3_U33 ( .A1(npu_inst_int_data_x_6__3__0_), .A2(
        npu_inst_pe_1_6_3_int_q_weight_1_), .ZN(npu_inst_pe_1_6_3_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_6_3_U32 ( .A1(npu_inst_n53), .A2(
        npu_inst_int_data_y_7__3__1_), .B1(npu_inst_pe_1_6_3_n3), .B2(
        npu_inst_int_data_x_6__4__1_), .ZN(npu_inst_pe_1_6_3_n63) );
  AOI22_X1 npu_inst_pe_1_6_3_U31 ( .A1(npu_inst_n53), .A2(
        npu_inst_int_data_y_7__3__0_), .B1(npu_inst_pe_1_6_3_n3), .B2(
        npu_inst_int_data_x_6__4__0_), .ZN(npu_inst_pe_1_6_3_n61) );
  INV_X1 npu_inst_pe_1_6_3_U30 ( .A(npu_inst_pe_1_6_3_int_data_0_), .ZN(
        npu_inst_pe_1_6_3_n13) );
  INV_X1 npu_inst_pe_1_6_3_U29 ( .A(npu_inst_n68), .ZN(npu_inst_pe_1_6_3_n5)
         );
  OR3_X1 npu_inst_pe_1_6_3_U28 ( .A1(npu_inst_pe_1_6_3_n6), .A2(
        npu_inst_pe_1_6_3_n8), .A3(npu_inst_pe_1_6_3_n5), .ZN(
        npu_inst_pe_1_6_3_n56) );
  OR3_X1 npu_inst_pe_1_6_3_U27 ( .A1(npu_inst_pe_1_6_3_n5), .A2(
        npu_inst_pe_1_6_3_n8), .A3(npu_inst_pe_1_6_3_n7), .ZN(
        npu_inst_pe_1_6_3_n48) );
  INV_X1 npu_inst_pe_1_6_3_U26 ( .A(npu_inst_pe_1_6_3_n5), .ZN(
        npu_inst_pe_1_6_3_n4) );
  INV_X1 npu_inst_pe_1_6_3_U25 ( .A(npu_inst_n123), .ZN(npu_inst_pe_1_6_3_n12)
         );
  OR3_X1 npu_inst_pe_1_6_3_U24 ( .A1(npu_inst_pe_1_6_3_n4), .A2(
        npu_inst_pe_1_6_3_n8), .A3(npu_inst_pe_1_6_3_n7), .ZN(
        npu_inst_pe_1_6_3_n52) );
  OR3_X1 npu_inst_pe_1_6_3_U23 ( .A1(npu_inst_pe_1_6_3_n6), .A2(
        npu_inst_pe_1_6_3_n8), .A3(npu_inst_pe_1_6_3_n4), .ZN(
        npu_inst_pe_1_6_3_n60) );
  NOR2_X1 npu_inst_pe_1_6_3_U22 ( .A1(npu_inst_pe_1_6_3_n60), .A2(
        npu_inst_pe_1_6_3_n3), .ZN(npu_inst_pe_1_6_3_n58) );
  NOR2_X1 npu_inst_pe_1_6_3_U21 ( .A1(npu_inst_pe_1_6_3_n56), .A2(
        npu_inst_pe_1_6_3_n3), .ZN(npu_inst_pe_1_6_3_n54) );
  NOR2_X1 npu_inst_pe_1_6_3_U20 ( .A1(npu_inst_pe_1_6_3_n52), .A2(
        npu_inst_pe_1_6_3_n3), .ZN(npu_inst_pe_1_6_3_n50) );
  NOR2_X1 npu_inst_pe_1_6_3_U19 ( .A1(npu_inst_pe_1_6_3_n48), .A2(
        npu_inst_pe_1_6_3_n3), .ZN(npu_inst_pe_1_6_3_n46) );
  NOR2_X1 npu_inst_pe_1_6_3_U18 ( .A1(npu_inst_pe_1_6_3_n40), .A2(
        npu_inst_pe_1_6_3_n3), .ZN(npu_inst_pe_1_6_3_n38) );
  NOR2_X1 npu_inst_pe_1_6_3_U17 ( .A1(npu_inst_pe_1_6_3_n44), .A2(
        npu_inst_pe_1_6_3_n3), .ZN(npu_inst_pe_1_6_3_n42) );
  BUF_X1 npu_inst_pe_1_6_3_U16 ( .A(npu_inst_n95), .Z(npu_inst_pe_1_6_3_n8) );
  BUF_X1 npu_inst_pe_1_6_3_U15 ( .A(npu_inst_pe_1_6_3_n12), .Z(
        npu_inst_pe_1_6_3_n11) );
  BUF_X1 npu_inst_pe_1_6_3_U14 ( .A(npu_inst_pe_1_6_3_n12), .Z(
        npu_inst_pe_1_6_3_n10) );
  BUF_X1 npu_inst_pe_1_6_3_U13 ( .A(npu_inst_pe_1_6_3_n12), .Z(
        npu_inst_pe_1_6_3_n9) );
  INV_X1 npu_inst_pe_1_6_3_U12 ( .A(npu_inst_pe_1_6_3_n38), .ZN(
        npu_inst_pe_1_6_3_n118) );
  INV_X1 npu_inst_pe_1_6_3_U11 ( .A(npu_inst_pe_1_6_3_n58), .ZN(
        npu_inst_pe_1_6_3_n114) );
  INV_X1 npu_inst_pe_1_6_3_U10 ( .A(npu_inst_pe_1_6_3_n54), .ZN(
        npu_inst_pe_1_6_3_n115) );
  INV_X1 npu_inst_pe_1_6_3_U9 ( .A(npu_inst_pe_1_6_3_n50), .ZN(
        npu_inst_pe_1_6_3_n116) );
  INV_X1 npu_inst_pe_1_6_3_U8 ( .A(npu_inst_pe_1_6_3_n46), .ZN(
        npu_inst_pe_1_6_3_n117) );
  INV_X1 npu_inst_pe_1_6_3_U7 ( .A(npu_inst_pe_1_6_3_n42), .ZN(
        npu_inst_pe_1_6_3_n119) );
  BUF_X1 npu_inst_pe_1_6_3_U6 ( .A(npu_inst_n13), .Z(npu_inst_pe_1_6_3_n2) );
  BUF_X1 npu_inst_pe_1_6_3_U5 ( .A(npu_inst_n13), .Z(npu_inst_pe_1_6_3_n1) );
  NOR2_X1 npu_inst_pe_1_6_3_U4 ( .A1(npu_inst_pe_1_6_3_int_q_weight_0_), .A2(
        npu_inst_pe_1_6_3_n1), .ZN(npu_inst_pe_1_6_3_n76) );
  NOR2_X1 npu_inst_pe_1_6_3_U3 ( .A1(npu_inst_pe_1_6_3_n27), .A2(
        npu_inst_pe_1_6_3_n1), .ZN(npu_inst_pe_1_6_3_n77) );
  FA_X1 npu_inst_pe_1_6_3_sub_77_U2_1 ( .A(npu_inst_pe_1_6_3_int_q_acc_1_), 
        .B(npu_inst_pe_1_6_3_n14), .CI(npu_inst_pe_1_6_3_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_6_3_sub_77_carry_2_), .S(npu_inst_pe_1_6_3_N66) );
  FA_X1 npu_inst_pe_1_6_3_add_79_U1_1 ( .A(npu_inst_pe_1_6_3_int_q_acc_1_), 
        .B(npu_inst_pe_1_6_3_int_data_1_), .CI(
        npu_inst_pe_1_6_3_add_79_carry_1_), .CO(
        npu_inst_pe_1_6_3_add_79_carry_2_), .S(npu_inst_pe_1_6_3_N74) );
  NAND3_X1 npu_inst_pe_1_6_3_U109 ( .A1(npu_inst_pe_1_6_3_n5), .A2(
        npu_inst_pe_1_6_3_n7), .A3(npu_inst_pe_1_6_3_n8), .ZN(
        npu_inst_pe_1_6_3_n44) );
  NAND3_X1 npu_inst_pe_1_6_3_U108 ( .A1(npu_inst_pe_1_6_3_n4), .A2(
        npu_inst_pe_1_6_3_n7), .A3(npu_inst_pe_1_6_3_n8), .ZN(
        npu_inst_pe_1_6_3_n40) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_6_3_n34), .CK(
        npu_inst_pe_1_6_3_net3120), .RN(npu_inst_pe_1_6_3_n9), .Q(
        npu_inst_pe_1_6_3_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_6_3_n35), .CK(
        npu_inst_pe_1_6_3_net3120), .RN(npu_inst_pe_1_6_3_n9), .Q(
        npu_inst_pe_1_6_3_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_6_3_n36), .CK(
        npu_inst_pe_1_6_3_net3120), .RN(npu_inst_pe_1_6_3_n9), .Q(
        npu_inst_pe_1_6_3_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_6_3_n98), .CK(
        npu_inst_pe_1_6_3_net3120), .RN(npu_inst_pe_1_6_3_n9), .Q(
        npu_inst_pe_1_6_3_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_6_3_n99), .CK(
        npu_inst_pe_1_6_3_net3120), .RN(npu_inst_pe_1_6_3_n9), .Q(
        npu_inst_pe_1_6_3_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_6_3_n100), 
        .CK(npu_inst_pe_1_6_3_net3120), .RN(npu_inst_pe_1_6_3_n9), .Q(
        npu_inst_pe_1_6_3_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_6_3_n33), .CK(
        npu_inst_pe_1_6_3_net3120), .RN(npu_inst_pe_1_6_3_n9), .Q(
        npu_inst_pe_1_6_3_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_6_3_n101), 
        .CK(npu_inst_pe_1_6_3_net3120), .RN(npu_inst_pe_1_6_3_n9), .Q(
        npu_inst_pe_1_6_3_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_weight_reg_0_ ( .D(npu_inst_n109), .CK(
        npu_inst_pe_1_6_3_net3126), .RN(npu_inst_pe_1_6_3_n9), .Q(
        npu_inst_pe_1_6_3_int_q_weight_0_), .QN(npu_inst_pe_1_6_3_n27) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_weight_reg_1_ ( .D(npu_inst_n115), .CK(
        npu_inst_pe_1_6_3_net3126), .RN(npu_inst_pe_1_6_3_n9), .Q(
        npu_inst_pe_1_6_3_int_q_weight_1_), .QN(npu_inst_pe_1_6_3_n26) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_6_3_n113), 
        .CK(npu_inst_pe_1_6_3_net3126), .RN(npu_inst_pe_1_6_3_n9), .Q(
        npu_inst_pe_1_6_3_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_6_3_n107), 
        .CK(npu_inst_pe_1_6_3_net3126), .RN(npu_inst_pe_1_6_3_n9), .Q(
        npu_inst_pe_1_6_3_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_6_3_n112), 
        .CK(npu_inst_pe_1_6_3_net3126), .RN(npu_inst_pe_1_6_3_n10), .Q(
        npu_inst_pe_1_6_3_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_6_3_n106), 
        .CK(npu_inst_pe_1_6_3_net3126), .RN(npu_inst_pe_1_6_3_n10), .Q(
        npu_inst_pe_1_6_3_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_6_3_n111), 
        .CK(npu_inst_pe_1_6_3_net3126), .RN(npu_inst_pe_1_6_3_n10), .Q(
        npu_inst_pe_1_6_3_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_6_3_n105), 
        .CK(npu_inst_pe_1_6_3_net3126), .RN(npu_inst_pe_1_6_3_n10), .Q(
        npu_inst_pe_1_6_3_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_6_3_n110), 
        .CK(npu_inst_pe_1_6_3_net3126), .RN(npu_inst_pe_1_6_3_n10), .Q(
        npu_inst_pe_1_6_3_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_6_3_n104), 
        .CK(npu_inst_pe_1_6_3_net3126), .RN(npu_inst_pe_1_6_3_n10), .Q(
        npu_inst_pe_1_6_3_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_6_3_n109), 
        .CK(npu_inst_pe_1_6_3_net3126), .RN(npu_inst_pe_1_6_3_n10), .Q(
        npu_inst_pe_1_6_3_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_6_3_n103), 
        .CK(npu_inst_pe_1_6_3_net3126), .RN(npu_inst_pe_1_6_3_n10), .Q(
        npu_inst_pe_1_6_3_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_6_3_n108), 
        .CK(npu_inst_pe_1_6_3_net3126), .RN(npu_inst_pe_1_6_3_n10), .Q(
        npu_inst_pe_1_6_3_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_6_3_n102), 
        .CK(npu_inst_pe_1_6_3_net3126), .RN(npu_inst_pe_1_6_3_n10), .Q(
        npu_inst_pe_1_6_3_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_6_3_n86), 
        .CK(npu_inst_pe_1_6_3_net3126), .RN(npu_inst_pe_1_6_3_n10), .Q(
        npu_inst_pe_1_6_3_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_6_3_n87), 
        .CK(npu_inst_pe_1_6_3_net3126), .RN(npu_inst_pe_1_6_3_n10), .Q(
        npu_inst_pe_1_6_3_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_6_3_n88), 
        .CK(npu_inst_pe_1_6_3_net3126), .RN(npu_inst_pe_1_6_3_n11), .Q(
        npu_inst_pe_1_6_3_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_6_3_n89), 
        .CK(npu_inst_pe_1_6_3_net3126), .RN(npu_inst_pe_1_6_3_n11), .Q(
        npu_inst_pe_1_6_3_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_6_3_n90), 
        .CK(npu_inst_pe_1_6_3_net3126), .RN(npu_inst_pe_1_6_3_n11), .Q(
        npu_inst_pe_1_6_3_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_6_3_n91), 
        .CK(npu_inst_pe_1_6_3_net3126), .RN(npu_inst_pe_1_6_3_n11), .Q(
        npu_inst_pe_1_6_3_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_6_3_n92), 
        .CK(npu_inst_pe_1_6_3_net3126), .RN(npu_inst_pe_1_6_3_n11), .Q(
        npu_inst_pe_1_6_3_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_6_3_n93), 
        .CK(npu_inst_pe_1_6_3_net3126), .RN(npu_inst_pe_1_6_3_n11), .Q(
        npu_inst_pe_1_6_3_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_6_3_n94), 
        .CK(npu_inst_pe_1_6_3_net3126), .RN(npu_inst_pe_1_6_3_n11), .Q(
        npu_inst_pe_1_6_3_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_6_3_n95), 
        .CK(npu_inst_pe_1_6_3_net3126), .RN(npu_inst_pe_1_6_3_n11), .Q(
        npu_inst_pe_1_6_3_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_6_3_n96), 
        .CK(npu_inst_pe_1_6_3_net3126), .RN(npu_inst_pe_1_6_3_n11), .Q(
        npu_inst_pe_1_6_3_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_6_3_n97), 
        .CK(npu_inst_pe_1_6_3_net3126), .RN(npu_inst_pe_1_6_3_n11), .Q(
        npu_inst_pe_1_6_3_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_6_3_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_6_3_N84), .SE(1'b0), .GCK(npu_inst_pe_1_6_3_net3120) );
  CLKGATETST_X1 npu_inst_pe_1_6_3_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n62), .SE(1'b0), .GCK(npu_inst_pe_1_6_3_net3126) );
  MUX2_X1 npu_inst_pe_1_6_4_U161 ( .A(npu_inst_pe_1_6_4_n31), .B(
        npu_inst_pe_1_6_4_n28), .S(npu_inst_pe_1_6_4_n7), .Z(
        npu_inst_pe_1_6_4_N93) );
  MUX2_X1 npu_inst_pe_1_6_4_U160 ( .A(npu_inst_pe_1_6_4_n30), .B(
        npu_inst_pe_1_6_4_n29), .S(npu_inst_n75), .Z(npu_inst_pe_1_6_4_n31) );
  MUX2_X1 npu_inst_pe_1_6_4_U159 ( .A(npu_inst_pe_1_6_4_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_6_4_int_q_reg_v_1__0_), .S(npu_inst_pe_1_6_4_n4), .Z(
        npu_inst_pe_1_6_4_n30) );
  MUX2_X1 npu_inst_pe_1_6_4_U158 ( .A(npu_inst_pe_1_6_4_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_6_4_int_q_reg_v_3__0_), .S(npu_inst_pe_1_6_4_n4), .Z(
        npu_inst_pe_1_6_4_n29) );
  MUX2_X1 npu_inst_pe_1_6_4_U157 ( .A(npu_inst_pe_1_6_4_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_6_4_int_q_reg_v_5__0_), .S(npu_inst_pe_1_6_4_n4), .Z(
        npu_inst_pe_1_6_4_n28) );
  MUX2_X1 npu_inst_pe_1_6_4_U156 ( .A(npu_inst_pe_1_6_4_n25), .B(
        npu_inst_pe_1_6_4_n22), .S(npu_inst_pe_1_6_4_n7), .Z(
        npu_inst_pe_1_6_4_N94) );
  MUX2_X1 npu_inst_pe_1_6_4_U155 ( .A(npu_inst_pe_1_6_4_n24), .B(
        npu_inst_pe_1_6_4_n23), .S(npu_inst_n75), .Z(npu_inst_pe_1_6_4_n25) );
  MUX2_X1 npu_inst_pe_1_6_4_U154 ( .A(npu_inst_pe_1_6_4_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_6_4_int_q_reg_v_1__1_), .S(npu_inst_pe_1_6_4_n4), .Z(
        npu_inst_pe_1_6_4_n24) );
  MUX2_X1 npu_inst_pe_1_6_4_U153 ( .A(npu_inst_pe_1_6_4_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_6_4_int_q_reg_v_3__1_), .S(npu_inst_pe_1_6_4_n4), .Z(
        npu_inst_pe_1_6_4_n23) );
  MUX2_X1 npu_inst_pe_1_6_4_U152 ( .A(npu_inst_pe_1_6_4_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_6_4_int_q_reg_v_5__1_), .S(npu_inst_pe_1_6_4_n4), .Z(
        npu_inst_pe_1_6_4_n22) );
  MUX2_X1 npu_inst_pe_1_6_4_U151 ( .A(npu_inst_pe_1_6_4_n21), .B(
        npu_inst_pe_1_6_4_n18), .S(npu_inst_pe_1_6_4_n7), .Z(
        npu_inst_int_data_x_6__4__1_) );
  MUX2_X1 npu_inst_pe_1_6_4_U150 ( .A(npu_inst_pe_1_6_4_n20), .B(
        npu_inst_pe_1_6_4_n19), .S(npu_inst_n75), .Z(npu_inst_pe_1_6_4_n21) );
  MUX2_X1 npu_inst_pe_1_6_4_U149 ( .A(npu_inst_pe_1_6_4_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_6_4_int_q_reg_h_1__1_), .S(npu_inst_pe_1_6_4_n4), .Z(
        npu_inst_pe_1_6_4_n20) );
  MUX2_X1 npu_inst_pe_1_6_4_U148 ( .A(npu_inst_pe_1_6_4_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_6_4_int_q_reg_h_3__1_), .S(npu_inst_pe_1_6_4_n4), .Z(
        npu_inst_pe_1_6_4_n19) );
  MUX2_X1 npu_inst_pe_1_6_4_U147 ( .A(npu_inst_pe_1_6_4_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_6_4_int_q_reg_h_5__1_), .S(npu_inst_pe_1_6_4_n4), .Z(
        npu_inst_pe_1_6_4_n18) );
  MUX2_X1 npu_inst_pe_1_6_4_U146 ( .A(npu_inst_pe_1_6_4_n17), .B(
        npu_inst_pe_1_6_4_n14), .S(npu_inst_pe_1_6_4_n7), .Z(
        npu_inst_int_data_x_6__4__0_) );
  MUX2_X1 npu_inst_pe_1_6_4_U145 ( .A(npu_inst_pe_1_6_4_n16), .B(
        npu_inst_pe_1_6_4_n15), .S(npu_inst_n75), .Z(npu_inst_pe_1_6_4_n17) );
  MUX2_X1 npu_inst_pe_1_6_4_U144 ( .A(npu_inst_pe_1_6_4_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_6_4_int_q_reg_h_1__0_), .S(npu_inst_pe_1_6_4_n4), .Z(
        npu_inst_pe_1_6_4_n16) );
  MUX2_X1 npu_inst_pe_1_6_4_U143 ( .A(npu_inst_pe_1_6_4_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_6_4_int_q_reg_h_3__0_), .S(npu_inst_pe_1_6_4_n4), .Z(
        npu_inst_pe_1_6_4_n15) );
  MUX2_X1 npu_inst_pe_1_6_4_U142 ( .A(npu_inst_pe_1_6_4_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_6_4_int_q_reg_h_5__0_), .S(npu_inst_pe_1_6_4_n4), .Z(
        npu_inst_pe_1_6_4_n14) );
  XOR2_X1 npu_inst_pe_1_6_4_U141 ( .A(npu_inst_pe_1_6_4_int_data_0_), .B(
        npu_inst_pe_1_6_4_int_q_acc_0_), .Z(npu_inst_pe_1_6_4_N73) );
  AND2_X1 npu_inst_pe_1_6_4_U140 ( .A1(npu_inst_pe_1_6_4_int_q_acc_0_), .A2(
        npu_inst_pe_1_6_4_int_data_0_), .ZN(npu_inst_pe_1_6_4_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_6_4_U139 ( .A(npu_inst_pe_1_6_4_int_q_acc_0_), .B(
        npu_inst_pe_1_6_4_n12), .ZN(npu_inst_pe_1_6_4_N65) );
  OR2_X1 npu_inst_pe_1_6_4_U138 ( .A1(npu_inst_pe_1_6_4_n12), .A2(
        npu_inst_pe_1_6_4_int_q_acc_0_), .ZN(npu_inst_pe_1_6_4_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_6_4_U137 ( .A(npu_inst_pe_1_6_4_int_q_acc_2_), .B(
        npu_inst_pe_1_6_4_add_79_carry_2_), .Z(npu_inst_pe_1_6_4_N75) );
  AND2_X1 npu_inst_pe_1_6_4_U136 ( .A1(npu_inst_pe_1_6_4_add_79_carry_2_), 
        .A2(npu_inst_pe_1_6_4_int_q_acc_2_), .ZN(
        npu_inst_pe_1_6_4_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_6_4_U135 ( .A(npu_inst_pe_1_6_4_int_q_acc_3_), .B(
        npu_inst_pe_1_6_4_add_79_carry_3_), .Z(npu_inst_pe_1_6_4_N76) );
  AND2_X1 npu_inst_pe_1_6_4_U134 ( .A1(npu_inst_pe_1_6_4_add_79_carry_3_), 
        .A2(npu_inst_pe_1_6_4_int_q_acc_3_), .ZN(
        npu_inst_pe_1_6_4_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_6_4_U133 ( .A(npu_inst_pe_1_6_4_int_q_acc_4_), .B(
        npu_inst_pe_1_6_4_add_79_carry_4_), .Z(npu_inst_pe_1_6_4_N77) );
  AND2_X1 npu_inst_pe_1_6_4_U132 ( .A1(npu_inst_pe_1_6_4_add_79_carry_4_), 
        .A2(npu_inst_pe_1_6_4_int_q_acc_4_), .ZN(
        npu_inst_pe_1_6_4_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_6_4_U131 ( .A(npu_inst_pe_1_6_4_int_q_acc_5_), .B(
        npu_inst_pe_1_6_4_add_79_carry_5_), .Z(npu_inst_pe_1_6_4_N78) );
  AND2_X1 npu_inst_pe_1_6_4_U130 ( .A1(npu_inst_pe_1_6_4_add_79_carry_5_), 
        .A2(npu_inst_pe_1_6_4_int_q_acc_5_), .ZN(
        npu_inst_pe_1_6_4_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_6_4_U129 ( .A(npu_inst_pe_1_6_4_int_q_acc_6_), .B(
        npu_inst_pe_1_6_4_add_79_carry_6_), .Z(npu_inst_pe_1_6_4_N79) );
  AND2_X1 npu_inst_pe_1_6_4_U128 ( .A1(npu_inst_pe_1_6_4_add_79_carry_6_), 
        .A2(npu_inst_pe_1_6_4_int_q_acc_6_), .ZN(
        npu_inst_pe_1_6_4_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_6_4_U127 ( .A(npu_inst_pe_1_6_4_int_q_acc_7_), .B(
        npu_inst_pe_1_6_4_add_79_carry_7_), .Z(npu_inst_pe_1_6_4_N80) );
  XNOR2_X1 npu_inst_pe_1_6_4_U126 ( .A(npu_inst_pe_1_6_4_sub_77_carry_2_), .B(
        npu_inst_pe_1_6_4_int_q_acc_2_), .ZN(npu_inst_pe_1_6_4_N67) );
  OR2_X1 npu_inst_pe_1_6_4_U125 ( .A1(npu_inst_pe_1_6_4_int_q_acc_2_), .A2(
        npu_inst_pe_1_6_4_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_6_4_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_6_4_U124 ( .A(npu_inst_pe_1_6_4_sub_77_carry_3_), .B(
        npu_inst_pe_1_6_4_int_q_acc_3_), .ZN(npu_inst_pe_1_6_4_N68) );
  OR2_X1 npu_inst_pe_1_6_4_U123 ( .A1(npu_inst_pe_1_6_4_int_q_acc_3_), .A2(
        npu_inst_pe_1_6_4_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_6_4_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_6_4_U122 ( .A(npu_inst_pe_1_6_4_sub_77_carry_4_), .B(
        npu_inst_pe_1_6_4_int_q_acc_4_), .ZN(npu_inst_pe_1_6_4_N69) );
  OR2_X1 npu_inst_pe_1_6_4_U121 ( .A1(npu_inst_pe_1_6_4_int_q_acc_4_), .A2(
        npu_inst_pe_1_6_4_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_6_4_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_6_4_U120 ( .A(npu_inst_pe_1_6_4_sub_77_carry_5_), .B(
        npu_inst_pe_1_6_4_int_q_acc_5_), .ZN(npu_inst_pe_1_6_4_N70) );
  OR2_X1 npu_inst_pe_1_6_4_U119 ( .A1(npu_inst_pe_1_6_4_int_q_acc_5_), .A2(
        npu_inst_pe_1_6_4_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_6_4_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_6_4_U118 ( .A(npu_inst_pe_1_6_4_sub_77_carry_6_), .B(
        npu_inst_pe_1_6_4_int_q_acc_6_), .ZN(npu_inst_pe_1_6_4_N71) );
  OR2_X1 npu_inst_pe_1_6_4_U117 ( .A1(npu_inst_pe_1_6_4_int_q_acc_6_), .A2(
        npu_inst_pe_1_6_4_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_6_4_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_6_4_U116 ( .A(npu_inst_pe_1_6_4_int_q_acc_7_), .B(
        npu_inst_pe_1_6_4_sub_77_carry_7_), .ZN(npu_inst_pe_1_6_4_N72) );
  INV_X1 npu_inst_pe_1_6_4_U115 ( .A(npu_inst_n75), .ZN(npu_inst_pe_1_6_4_n6)
         );
  INV_X1 npu_inst_pe_1_6_4_U114 ( .A(npu_inst_n53), .ZN(npu_inst_pe_1_6_4_n3)
         );
  AOI22_X1 npu_inst_pe_1_6_4_U113 ( .A1(npu_inst_int_data_y_7__4__0_), .A2(
        npu_inst_pe_1_6_4_n58), .B1(npu_inst_pe_1_6_4_n113), .B2(
        npu_inst_pe_1_6_4_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_6_4_n57) );
  INV_X1 npu_inst_pe_1_6_4_U112 ( .A(npu_inst_pe_1_6_4_n57), .ZN(
        npu_inst_pe_1_6_4_n107) );
  AOI22_X1 npu_inst_pe_1_6_4_U111 ( .A1(npu_inst_int_data_y_7__4__0_), .A2(
        npu_inst_pe_1_6_4_n54), .B1(npu_inst_pe_1_6_4_n114), .B2(
        npu_inst_pe_1_6_4_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_6_4_n53) );
  INV_X1 npu_inst_pe_1_6_4_U110 ( .A(npu_inst_pe_1_6_4_n53), .ZN(
        npu_inst_pe_1_6_4_n108) );
  AOI22_X1 npu_inst_pe_1_6_4_U107 ( .A1(npu_inst_int_data_y_7__4__0_), .A2(
        npu_inst_pe_1_6_4_n50), .B1(npu_inst_pe_1_6_4_n115), .B2(
        npu_inst_pe_1_6_4_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_6_4_n49) );
  INV_X1 npu_inst_pe_1_6_4_U106 ( .A(npu_inst_pe_1_6_4_n49), .ZN(
        npu_inst_pe_1_6_4_n109) );
  AOI22_X1 npu_inst_pe_1_6_4_U105 ( .A1(npu_inst_int_data_y_7__4__0_), .A2(
        npu_inst_pe_1_6_4_n46), .B1(npu_inst_pe_1_6_4_n116), .B2(
        npu_inst_pe_1_6_4_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_6_4_n45) );
  INV_X1 npu_inst_pe_1_6_4_U104 ( .A(npu_inst_pe_1_6_4_n45), .ZN(
        npu_inst_pe_1_6_4_n110) );
  AOI22_X1 npu_inst_pe_1_6_4_U103 ( .A1(npu_inst_int_data_y_7__4__0_), .A2(
        npu_inst_pe_1_6_4_n42), .B1(npu_inst_pe_1_6_4_n118), .B2(
        npu_inst_pe_1_6_4_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_6_4_n41) );
  INV_X1 npu_inst_pe_1_6_4_U102 ( .A(npu_inst_pe_1_6_4_n41), .ZN(
        npu_inst_pe_1_6_4_n111) );
  AOI22_X1 npu_inst_pe_1_6_4_U101 ( .A1(npu_inst_int_data_y_7__4__1_), .A2(
        npu_inst_pe_1_6_4_n58), .B1(npu_inst_pe_1_6_4_n113), .B2(
        npu_inst_pe_1_6_4_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_6_4_n59) );
  INV_X1 npu_inst_pe_1_6_4_U100 ( .A(npu_inst_pe_1_6_4_n59), .ZN(
        npu_inst_pe_1_6_4_n101) );
  AOI22_X1 npu_inst_pe_1_6_4_U99 ( .A1(npu_inst_int_data_y_7__4__1_), .A2(
        npu_inst_pe_1_6_4_n54), .B1(npu_inst_pe_1_6_4_n114), .B2(
        npu_inst_pe_1_6_4_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_6_4_n55) );
  INV_X1 npu_inst_pe_1_6_4_U98 ( .A(npu_inst_pe_1_6_4_n55), .ZN(
        npu_inst_pe_1_6_4_n102) );
  AOI22_X1 npu_inst_pe_1_6_4_U97 ( .A1(npu_inst_int_data_y_7__4__1_), .A2(
        npu_inst_pe_1_6_4_n50), .B1(npu_inst_pe_1_6_4_n115), .B2(
        npu_inst_pe_1_6_4_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_6_4_n51) );
  INV_X1 npu_inst_pe_1_6_4_U96 ( .A(npu_inst_pe_1_6_4_n51), .ZN(
        npu_inst_pe_1_6_4_n103) );
  AOI22_X1 npu_inst_pe_1_6_4_U95 ( .A1(npu_inst_int_data_y_7__4__1_), .A2(
        npu_inst_pe_1_6_4_n46), .B1(npu_inst_pe_1_6_4_n116), .B2(
        npu_inst_pe_1_6_4_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_6_4_n47) );
  INV_X1 npu_inst_pe_1_6_4_U94 ( .A(npu_inst_pe_1_6_4_n47), .ZN(
        npu_inst_pe_1_6_4_n104) );
  AOI22_X1 npu_inst_pe_1_6_4_U93 ( .A1(npu_inst_int_data_y_7__4__1_), .A2(
        npu_inst_pe_1_6_4_n42), .B1(npu_inst_pe_1_6_4_n118), .B2(
        npu_inst_pe_1_6_4_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_6_4_n43) );
  INV_X1 npu_inst_pe_1_6_4_U92 ( .A(npu_inst_pe_1_6_4_n43), .ZN(
        npu_inst_pe_1_6_4_n105) );
  AOI22_X1 npu_inst_pe_1_6_4_U91 ( .A1(npu_inst_pe_1_6_4_n38), .A2(
        npu_inst_int_data_y_7__4__1_), .B1(npu_inst_pe_1_6_4_n117), .B2(
        npu_inst_pe_1_6_4_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_6_4_n39) );
  INV_X1 npu_inst_pe_1_6_4_U90 ( .A(npu_inst_pe_1_6_4_n39), .ZN(
        npu_inst_pe_1_6_4_n106) );
  AOI22_X1 npu_inst_pe_1_6_4_U89 ( .A1(npu_inst_pe_1_6_4_n38), .A2(
        npu_inst_int_data_y_7__4__0_), .B1(npu_inst_pe_1_6_4_n117), .B2(
        npu_inst_pe_1_6_4_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_6_4_n37) );
  INV_X1 npu_inst_pe_1_6_4_U88 ( .A(npu_inst_pe_1_6_4_n37), .ZN(
        npu_inst_pe_1_6_4_n112) );
  NAND2_X1 npu_inst_pe_1_6_4_U87 ( .A1(npu_inst_pe_1_6_4_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_6_4_n60), .ZN(npu_inst_pe_1_6_4_n74) );
  OAI21_X1 npu_inst_pe_1_6_4_U86 ( .B1(npu_inst_pe_1_6_4_n63), .B2(
        npu_inst_pe_1_6_4_n60), .A(npu_inst_pe_1_6_4_n74), .ZN(
        npu_inst_pe_1_6_4_n97) );
  NAND2_X1 npu_inst_pe_1_6_4_U85 ( .A1(npu_inst_pe_1_6_4_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_6_4_n60), .ZN(npu_inst_pe_1_6_4_n73) );
  OAI21_X1 npu_inst_pe_1_6_4_U84 ( .B1(npu_inst_pe_1_6_4_n61), .B2(
        npu_inst_pe_1_6_4_n60), .A(npu_inst_pe_1_6_4_n73), .ZN(
        npu_inst_pe_1_6_4_n96) );
  NAND2_X1 npu_inst_pe_1_6_4_U83 ( .A1(npu_inst_pe_1_6_4_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_6_4_n56), .ZN(npu_inst_pe_1_6_4_n72) );
  OAI21_X1 npu_inst_pe_1_6_4_U82 ( .B1(npu_inst_pe_1_6_4_n63), .B2(
        npu_inst_pe_1_6_4_n56), .A(npu_inst_pe_1_6_4_n72), .ZN(
        npu_inst_pe_1_6_4_n95) );
  NAND2_X1 npu_inst_pe_1_6_4_U81 ( .A1(npu_inst_pe_1_6_4_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_6_4_n56), .ZN(npu_inst_pe_1_6_4_n71) );
  OAI21_X1 npu_inst_pe_1_6_4_U80 ( .B1(npu_inst_pe_1_6_4_n61), .B2(
        npu_inst_pe_1_6_4_n56), .A(npu_inst_pe_1_6_4_n71), .ZN(
        npu_inst_pe_1_6_4_n94) );
  NAND2_X1 npu_inst_pe_1_6_4_U79 ( .A1(npu_inst_pe_1_6_4_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_6_4_n52), .ZN(npu_inst_pe_1_6_4_n70) );
  OAI21_X1 npu_inst_pe_1_6_4_U78 ( .B1(npu_inst_pe_1_6_4_n63), .B2(
        npu_inst_pe_1_6_4_n52), .A(npu_inst_pe_1_6_4_n70), .ZN(
        npu_inst_pe_1_6_4_n93) );
  NAND2_X1 npu_inst_pe_1_6_4_U77 ( .A1(npu_inst_pe_1_6_4_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_6_4_n52), .ZN(npu_inst_pe_1_6_4_n69) );
  OAI21_X1 npu_inst_pe_1_6_4_U76 ( .B1(npu_inst_pe_1_6_4_n61), .B2(
        npu_inst_pe_1_6_4_n52), .A(npu_inst_pe_1_6_4_n69), .ZN(
        npu_inst_pe_1_6_4_n92) );
  NAND2_X1 npu_inst_pe_1_6_4_U75 ( .A1(npu_inst_pe_1_6_4_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_6_4_n48), .ZN(npu_inst_pe_1_6_4_n68) );
  OAI21_X1 npu_inst_pe_1_6_4_U74 ( .B1(npu_inst_pe_1_6_4_n63), .B2(
        npu_inst_pe_1_6_4_n48), .A(npu_inst_pe_1_6_4_n68), .ZN(
        npu_inst_pe_1_6_4_n91) );
  NAND2_X1 npu_inst_pe_1_6_4_U73 ( .A1(npu_inst_pe_1_6_4_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_6_4_n48), .ZN(npu_inst_pe_1_6_4_n67) );
  OAI21_X1 npu_inst_pe_1_6_4_U72 ( .B1(npu_inst_pe_1_6_4_n61), .B2(
        npu_inst_pe_1_6_4_n48), .A(npu_inst_pe_1_6_4_n67), .ZN(
        npu_inst_pe_1_6_4_n90) );
  NAND2_X1 npu_inst_pe_1_6_4_U71 ( .A1(npu_inst_pe_1_6_4_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_6_4_n44), .ZN(npu_inst_pe_1_6_4_n66) );
  OAI21_X1 npu_inst_pe_1_6_4_U70 ( .B1(npu_inst_pe_1_6_4_n63), .B2(
        npu_inst_pe_1_6_4_n44), .A(npu_inst_pe_1_6_4_n66), .ZN(
        npu_inst_pe_1_6_4_n89) );
  NAND2_X1 npu_inst_pe_1_6_4_U69 ( .A1(npu_inst_pe_1_6_4_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_6_4_n44), .ZN(npu_inst_pe_1_6_4_n65) );
  OAI21_X1 npu_inst_pe_1_6_4_U68 ( .B1(npu_inst_pe_1_6_4_n61), .B2(
        npu_inst_pe_1_6_4_n44), .A(npu_inst_pe_1_6_4_n65), .ZN(
        npu_inst_pe_1_6_4_n88) );
  NAND2_X1 npu_inst_pe_1_6_4_U67 ( .A1(npu_inst_pe_1_6_4_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_6_4_n40), .ZN(npu_inst_pe_1_6_4_n64) );
  OAI21_X1 npu_inst_pe_1_6_4_U66 ( .B1(npu_inst_pe_1_6_4_n63), .B2(
        npu_inst_pe_1_6_4_n40), .A(npu_inst_pe_1_6_4_n64), .ZN(
        npu_inst_pe_1_6_4_n87) );
  NAND2_X1 npu_inst_pe_1_6_4_U65 ( .A1(npu_inst_pe_1_6_4_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_6_4_n40), .ZN(npu_inst_pe_1_6_4_n62) );
  OAI21_X1 npu_inst_pe_1_6_4_U64 ( .B1(npu_inst_pe_1_6_4_n61), .B2(
        npu_inst_pe_1_6_4_n40), .A(npu_inst_pe_1_6_4_n62), .ZN(
        npu_inst_pe_1_6_4_n86) );
  AND2_X1 npu_inst_pe_1_6_4_U63 ( .A1(npu_inst_pe_1_6_4_N93), .A2(npu_inst_n53), .ZN(npu_inst_int_data_y_6__4__0_) );
  AND2_X1 npu_inst_pe_1_6_4_U62 ( .A1(npu_inst_n53), .A2(npu_inst_pe_1_6_4_N94), .ZN(npu_inst_int_data_y_6__4__1_) );
  NOR3_X1 npu_inst_pe_1_6_4_U61 ( .A1(npu_inst_pe_1_6_4_n26), .A2(npu_inst_n53), .A3(npu_inst_int_ckg[11]), .ZN(npu_inst_pe_1_6_4_n85) );
  OR2_X1 npu_inst_pe_1_6_4_U60 ( .A1(npu_inst_pe_1_6_4_n85), .A2(
        npu_inst_pe_1_6_4_n2), .ZN(npu_inst_pe_1_6_4_N84) );
  AND2_X1 npu_inst_pe_1_6_4_U59 ( .A1(npu_inst_pe_1_6_4_int_q_acc_0_), .A2(
        npu_inst_pe_1_6_4_n1), .ZN(npu_inst_int_data_res_6__4__0_) );
  AND2_X1 npu_inst_pe_1_6_4_U58 ( .A1(npu_inst_pe_1_6_4_n2), .A2(
        npu_inst_pe_1_6_4_int_q_acc_7_), .ZN(npu_inst_int_data_res_6__4__7_)
         );
  AND2_X1 npu_inst_pe_1_6_4_U57 ( .A1(npu_inst_pe_1_6_4_int_q_acc_1_), .A2(
        npu_inst_pe_1_6_4_n1), .ZN(npu_inst_int_data_res_6__4__1_) );
  AND2_X1 npu_inst_pe_1_6_4_U56 ( .A1(npu_inst_pe_1_6_4_int_q_acc_2_), .A2(
        npu_inst_pe_1_6_4_n1), .ZN(npu_inst_int_data_res_6__4__2_) );
  AND2_X1 npu_inst_pe_1_6_4_U55 ( .A1(npu_inst_pe_1_6_4_int_q_acc_3_), .A2(
        npu_inst_pe_1_6_4_n2), .ZN(npu_inst_int_data_res_6__4__3_) );
  AND2_X1 npu_inst_pe_1_6_4_U54 ( .A1(npu_inst_pe_1_6_4_int_q_acc_4_), .A2(
        npu_inst_pe_1_6_4_n2), .ZN(npu_inst_int_data_res_6__4__4_) );
  AND2_X1 npu_inst_pe_1_6_4_U53 ( .A1(npu_inst_pe_1_6_4_int_q_acc_5_), .A2(
        npu_inst_pe_1_6_4_n2), .ZN(npu_inst_int_data_res_6__4__5_) );
  AND2_X1 npu_inst_pe_1_6_4_U52 ( .A1(npu_inst_pe_1_6_4_int_q_acc_6_), .A2(
        npu_inst_pe_1_6_4_n2), .ZN(npu_inst_int_data_res_6__4__6_) );
  AOI222_X1 npu_inst_pe_1_6_4_U51 ( .A1(npu_inst_int_data_res_7__4__0_), .A2(
        npu_inst_pe_1_6_4_n1), .B1(npu_inst_pe_1_6_4_N73), .B2(
        npu_inst_pe_1_6_4_n76), .C1(npu_inst_pe_1_6_4_N65), .C2(
        npu_inst_pe_1_6_4_n77), .ZN(npu_inst_pe_1_6_4_n84) );
  INV_X1 npu_inst_pe_1_6_4_U50 ( .A(npu_inst_pe_1_6_4_n84), .ZN(
        npu_inst_pe_1_6_4_n100) );
  AOI222_X1 npu_inst_pe_1_6_4_U49 ( .A1(npu_inst_int_data_res_7__4__7_), .A2(
        npu_inst_pe_1_6_4_n1), .B1(npu_inst_pe_1_6_4_N80), .B2(
        npu_inst_pe_1_6_4_n76), .C1(npu_inst_pe_1_6_4_N72), .C2(
        npu_inst_pe_1_6_4_n77), .ZN(npu_inst_pe_1_6_4_n75) );
  INV_X1 npu_inst_pe_1_6_4_U48 ( .A(npu_inst_pe_1_6_4_n75), .ZN(
        npu_inst_pe_1_6_4_n32) );
  AOI222_X1 npu_inst_pe_1_6_4_U47 ( .A1(npu_inst_int_data_res_7__4__1_), .A2(
        npu_inst_pe_1_6_4_n1), .B1(npu_inst_pe_1_6_4_N74), .B2(
        npu_inst_pe_1_6_4_n76), .C1(npu_inst_pe_1_6_4_N66), .C2(
        npu_inst_pe_1_6_4_n77), .ZN(npu_inst_pe_1_6_4_n83) );
  INV_X1 npu_inst_pe_1_6_4_U46 ( .A(npu_inst_pe_1_6_4_n83), .ZN(
        npu_inst_pe_1_6_4_n99) );
  AOI222_X1 npu_inst_pe_1_6_4_U45 ( .A1(npu_inst_int_data_res_7__4__2_), .A2(
        npu_inst_pe_1_6_4_n1), .B1(npu_inst_pe_1_6_4_N75), .B2(
        npu_inst_pe_1_6_4_n76), .C1(npu_inst_pe_1_6_4_N67), .C2(
        npu_inst_pe_1_6_4_n77), .ZN(npu_inst_pe_1_6_4_n82) );
  INV_X1 npu_inst_pe_1_6_4_U44 ( .A(npu_inst_pe_1_6_4_n82), .ZN(
        npu_inst_pe_1_6_4_n98) );
  AOI222_X1 npu_inst_pe_1_6_4_U43 ( .A1(npu_inst_int_data_res_7__4__3_), .A2(
        npu_inst_pe_1_6_4_n1), .B1(npu_inst_pe_1_6_4_N76), .B2(
        npu_inst_pe_1_6_4_n76), .C1(npu_inst_pe_1_6_4_N68), .C2(
        npu_inst_pe_1_6_4_n77), .ZN(npu_inst_pe_1_6_4_n81) );
  INV_X1 npu_inst_pe_1_6_4_U42 ( .A(npu_inst_pe_1_6_4_n81), .ZN(
        npu_inst_pe_1_6_4_n36) );
  AOI222_X1 npu_inst_pe_1_6_4_U41 ( .A1(npu_inst_int_data_res_7__4__4_), .A2(
        npu_inst_pe_1_6_4_n1), .B1(npu_inst_pe_1_6_4_N77), .B2(
        npu_inst_pe_1_6_4_n76), .C1(npu_inst_pe_1_6_4_N69), .C2(
        npu_inst_pe_1_6_4_n77), .ZN(npu_inst_pe_1_6_4_n80) );
  INV_X1 npu_inst_pe_1_6_4_U40 ( .A(npu_inst_pe_1_6_4_n80), .ZN(
        npu_inst_pe_1_6_4_n35) );
  AOI222_X1 npu_inst_pe_1_6_4_U39 ( .A1(npu_inst_int_data_res_7__4__5_), .A2(
        npu_inst_pe_1_6_4_n1), .B1(npu_inst_pe_1_6_4_N78), .B2(
        npu_inst_pe_1_6_4_n76), .C1(npu_inst_pe_1_6_4_N70), .C2(
        npu_inst_pe_1_6_4_n77), .ZN(npu_inst_pe_1_6_4_n79) );
  INV_X1 npu_inst_pe_1_6_4_U38 ( .A(npu_inst_pe_1_6_4_n79), .ZN(
        npu_inst_pe_1_6_4_n34) );
  AOI222_X1 npu_inst_pe_1_6_4_U37 ( .A1(npu_inst_int_data_res_7__4__6_), .A2(
        npu_inst_pe_1_6_4_n1), .B1(npu_inst_pe_1_6_4_N79), .B2(
        npu_inst_pe_1_6_4_n76), .C1(npu_inst_pe_1_6_4_N71), .C2(
        npu_inst_pe_1_6_4_n77), .ZN(npu_inst_pe_1_6_4_n78) );
  INV_X1 npu_inst_pe_1_6_4_U36 ( .A(npu_inst_pe_1_6_4_n78), .ZN(
        npu_inst_pe_1_6_4_n33) );
  INV_X1 npu_inst_pe_1_6_4_U35 ( .A(npu_inst_pe_1_6_4_int_data_1_), .ZN(
        npu_inst_pe_1_6_4_n13) );
  AND2_X1 npu_inst_pe_1_6_4_U34 ( .A1(npu_inst_int_data_x_6__4__1_), .A2(
        npu_inst_pe_1_6_4_int_q_weight_1_), .ZN(npu_inst_pe_1_6_4_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_6_4_U33 ( .A1(npu_inst_int_data_x_6__4__0_), .A2(
        npu_inst_pe_1_6_4_int_q_weight_1_), .ZN(npu_inst_pe_1_6_4_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_6_4_U32 ( .A1(npu_inst_n53), .A2(
        npu_inst_int_data_y_7__4__1_), .B1(npu_inst_pe_1_6_4_n3), .B2(
        npu_inst_int_data_x_6__5__1_), .ZN(npu_inst_pe_1_6_4_n63) );
  AOI22_X1 npu_inst_pe_1_6_4_U31 ( .A1(npu_inst_n53), .A2(
        npu_inst_int_data_y_7__4__0_), .B1(npu_inst_pe_1_6_4_n3), .B2(
        npu_inst_int_data_x_6__5__0_), .ZN(npu_inst_pe_1_6_4_n61) );
  INV_X1 npu_inst_pe_1_6_4_U30 ( .A(npu_inst_pe_1_6_4_int_data_0_), .ZN(
        npu_inst_pe_1_6_4_n12) );
  INV_X1 npu_inst_pe_1_6_4_U29 ( .A(npu_inst_n67), .ZN(npu_inst_pe_1_6_4_n5)
         );
  OR3_X1 npu_inst_pe_1_6_4_U28 ( .A1(npu_inst_n75), .A2(npu_inst_pe_1_6_4_n7), 
        .A3(npu_inst_pe_1_6_4_n5), .ZN(npu_inst_pe_1_6_4_n56) );
  OR3_X1 npu_inst_pe_1_6_4_U27 ( .A1(npu_inst_pe_1_6_4_n5), .A2(
        npu_inst_pe_1_6_4_n7), .A3(npu_inst_pe_1_6_4_n6), .ZN(
        npu_inst_pe_1_6_4_n48) );
  INV_X1 npu_inst_pe_1_6_4_U26 ( .A(npu_inst_pe_1_6_4_n5), .ZN(
        npu_inst_pe_1_6_4_n4) );
  INV_X1 npu_inst_pe_1_6_4_U25 ( .A(npu_inst_n122), .ZN(npu_inst_pe_1_6_4_n11)
         );
  OR3_X1 npu_inst_pe_1_6_4_U24 ( .A1(npu_inst_pe_1_6_4_n4), .A2(
        npu_inst_pe_1_6_4_n7), .A3(npu_inst_pe_1_6_4_n6), .ZN(
        npu_inst_pe_1_6_4_n52) );
  OR3_X1 npu_inst_pe_1_6_4_U23 ( .A1(npu_inst_n75), .A2(npu_inst_pe_1_6_4_n7), 
        .A3(npu_inst_pe_1_6_4_n4), .ZN(npu_inst_pe_1_6_4_n60) );
  NOR2_X1 npu_inst_pe_1_6_4_U22 ( .A1(npu_inst_pe_1_6_4_n60), .A2(
        npu_inst_pe_1_6_4_n3), .ZN(npu_inst_pe_1_6_4_n58) );
  NOR2_X1 npu_inst_pe_1_6_4_U21 ( .A1(npu_inst_pe_1_6_4_n56), .A2(
        npu_inst_pe_1_6_4_n3), .ZN(npu_inst_pe_1_6_4_n54) );
  NOR2_X1 npu_inst_pe_1_6_4_U20 ( .A1(npu_inst_pe_1_6_4_n52), .A2(
        npu_inst_pe_1_6_4_n3), .ZN(npu_inst_pe_1_6_4_n50) );
  NOR2_X1 npu_inst_pe_1_6_4_U19 ( .A1(npu_inst_pe_1_6_4_n48), .A2(
        npu_inst_pe_1_6_4_n3), .ZN(npu_inst_pe_1_6_4_n46) );
  NOR2_X1 npu_inst_pe_1_6_4_U18 ( .A1(npu_inst_pe_1_6_4_n40), .A2(
        npu_inst_pe_1_6_4_n3), .ZN(npu_inst_pe_1_6_4_n38) );
  NOR2_X1 npu_inst_pe_1_6_4_U17 ( .A1(npu_inst_pe_1_6_4_n44), .A2(
        npu_inst_pe_1_6_4_n3), .ZN(npu_inst_pe_1_6_4_n42) );
  BUF_X1 npu_inst_pe_1_6_4_U16 ( .A(npu_inst_n94), .Z(npu_inst_pe_1_6_4_n7) );
  BUF_X1 npu_inst_pe_1_6_4_U15 ( .A(npu_inst_pe_1_6_4_n11), .Z(
        npu_inst_pe_1_6_4_n10) );
  BUF_X1 npu_inst_pe_1_6_4_U14 ( .A(npu_inst_pe_1_6_4_n11), .Z(
        npu_inst_pe_1_6_4_n9) );
  BUF_X1 npu_inst_pe_1_6_4_U13 ( .A(npu_inst_pe_1_6_4_n11), .Z(
        npu_inst_pe_1_6_4_n8) );
  INV_X1 npu_inst_pe_1_6_4_U12 ( .A(npu_inst_pe_1_6_4_n38), .ZN(
        npu_inst_pe_1_6_4_n117) );
  INV_X1 npu_inst_pe_1_6_4_U11 ( .A(npu_inst_pe_1_6_4_n58), .ZN(
        npu_inst_pe_1_6_4_n113) );
  INV_X1 npu_inst_pe_1_6_4_U10 ( .A(npu_inst_pe_1_6_4_n54), .ZN(
        npu_inst_pe_1_6_4_n114) );
  INV_X1 npu_inst_pe_1_6_4_U9 ( .A(npu_inst_pe_1_6_4_n50), .ZN(
        npu_inst_pe_1_6_4_n115) );
  INV_X1 npu_inst_pe_1_6_4_U8 ( .A(npu_inst_pe_1_6_4_n46), .ZN(
        npu_inst_pe_1_6_4_n116) );
  INV_X1 npu_inst_pe_1_6_4_U7 ( .A(npu_inst_pe_1_6_4_n42), .ZN(
        npu_inst_pe_1_6_4_n118) );
  BUF_X1 npu_inst_pe_1_6_4_U6 ( .A(npu_inst_n12), .Z(npu_inst_pe_1_6_4_n2) );
  BUF_X1 npu_inst_pe_1_6_4_U5 ( .A(npu_inst_n12), .Z(npu_inst_pe_1_6_4_n1) );
  NOR2_X1 npu_inst_pe_1_6_4_U4 ( .A1(npu_inst_pe_1_6_4_int_q_weight_0_), .A2(
        npu_inst_pe_1_6_4_n1), .ZN(npu_inst_pe_1_6_4_n76) );
  NOR2_X1 npu_inst_pe_1_6_4_U3 ( .A1(npu_inst_pe_1_6_4_n27), .A2(
        npu_inst_pe_1_6_4_n1), .ZN(npu_inst_pe_1_6_4_n77) );
  FA_X1 npu_inst_pe_1_6_4_sub_77_U2_1 ( .A(npu_inst_pe_1_6_4_int_q_acc_1_), 
        .B(npu_inst_pe_1_6_4_n13), .CI(npu_inst_pe_1_6_4_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_6_4_sub_77_carry_2_), .S(npu_inst_pe_1_6_4_N66) );
  FA_X1 npu_inst_pe_1_6_4_add_79_U1_1 ( .A(npu_inst_pe_1_6_4_int_q_acc_1_), 
        .B(npu_inst_pe_1_6_4_int_data_1_), .CI(
        npu_inst_pe_1_6_4_add_79_carry_1_), .CO(
        npu_inst_pe_1_6_4_add_79_carry_2_), .S(npu_inst_pe_1_6_4_N74) );
  NAND3_X1 npu_inst_pe_1_6_4_U109 ( .A1(npu_inst_pe_1_6_4_n5), .A2(
        npu_inst_pe_1_6_4_n6), .A3(npu_inst_pe_1_6_4_n7), .ZN(
        npu_inst_pe_1_6_4_n44) );
  NAND3_X1 npu_inst_pe_1_6_4_U108 ( .A1(npu_inst_pe_1_6_4_n4), .A2(
        npu_inst_pe_1_6_4_n6), .A3(npu_inst_pe_1_6_4_n7), .ZN(
        npu_inst_pe_1_6_4_n40) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_6_4_n33), .CK(
        npu_inst_pe_1_6_4_net3097), .RN(npu_inst_pe_1_6_4_n8), .Q(
        npu_inst_pe_1_6_4_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_6_4_n34), .CK(
        npu_inst_pe_1_6_4_net3097), .RN(npu_inst_pe_1_6_4_n8), .Q(
        npu_inst_pe_1_6_4_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_6_4_n35), .CK(
        npu_inst_pe_1_6_4_net3097), .RN(npu_inst_pe_1_6_4_n8), .Q(
        npu_inst_pe_1_6_4_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_6_4_n36), .CK(
        npu_inst_pe_1_6_4_net3097), .RN(npu_inst_pe_1_6_4_n8), .Q(
        npu_inst_pe_1_6_4_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_6_4_n98), .CK(
        npu_inst_pe_1_6_4_net3097), .RN(npu_inst_pe_1_6_4_n8), .Q(
        npu_inst_pe_1_6_4_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_6_4_n99), .CK(
        npu_inst_pe_1_6_4_net3097), .RN(npu_inst_pe_1_6_4_n8), .Q(
        npu_inst_pe_1_6_4_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_6_4_n32), .CK(
        npu_inst_pe_1_6_4_net3097), .RN(npu_inst_pe_1_6_4_n8), .Q(
        npu_inst_pe_1_6_4_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_6_4_n100), 
        .CK(npu_inst_pe_1_6_4_net3097), .RN(npu_inst_pe_1_6_4_n8), .Q(
        npu_inst_pe_1_6_4_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_weight_reg_0_ ( .D(npu_inst_n108), .CK(
        npu_inst_pe_1_6_4_net3103), .RN(npu_inst_pe_1_6_4_n8), .Q(
        npu_inst_pe_1_6_4_int_q_weight_0_), .QN(npu_inst_pe_1_6_4_n27) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_weight_reg_1_ ( .D(npu_inst_n114), .CK(
        npu_inst_pe_1_6_4_net3103), .RN(npu_inst_pe_1_6_4_n8), .Q(
        npu_inst_pe_1_6_4_int_q_weight_1_), .QN(npu_inst_pe_1_6_4_n26) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_6_4_n112), 
        .CK(npu_inst_pe_1_6_4_net3103), .RN(npu_inst_pe_1_6_4_n8), .Q(
        npu_inst_pe_1_6_4_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_6_4_n106), 
        .CK(npu_inst_pe_1_6_4_net3103), .RN(npu_inst_pe_1_6_4_n8), .Q(
        npu_inst_pe_1_6_4_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_6_4_n111), 
        .CK(npu_inst_pe_1_6_4_net3103), .RN(npu_inst_pe_1_6_4_n9), .Q(
        npu_inst_pe_1_6_4_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_6_4_n105), 
        .CK(npu_inst_pe_1_6_4_net3103), .RN(npu_inst_pe_1_6_4_n9), .Q(
        npu_inst_pe_1_6_4_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_6_4_n110), 
        .CK(npu_inst_pe_1_6_4_net3103), .RN(npu_inst_pe_1_6_4_n9), .Q(
        npu_inst_pe_1_6_4_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_6_4_n104), 
        .CK(npu_inst_pe_1_6_4_net3103), .RN(npu_inst_pe_1_6_4_n9), .Q(
        npu_inst_pe_1_6_4_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_6_4_n109), 
        .CK(npu_inst_pe_1_6_4_net3103), .RN(npu_inst_pe_1_6_4_n9), .Q(
        npu_inst_pe_1_6_4_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_6_4_n103), 
        .CK(npu_inst_pe_1_6_4_net3103), .RN(npu_inst_pe_1_6_4_n9), .Q(
        npu_inst_pe_1_6_4_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_6_4_n108), 
        .CK(npu_inst_pe_1_6_4_net3103), .RN(npu_inst_pe_1_6_4_n9), .Q(
        npu_inst_pe_1_6_4_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_6_4_n102), 
        .CK(npu_inst_pe_1_6_4_net3103), .RN(npu_inst_pe_1_6_4_n9), .Q(
        npu_inst_pe_1_6_4_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_6_4_n107), 
        .CK(npu_inst_pe_1_6_4_net3103), .RN(npu_inst_pe_1_6_4_n9), .Q(
        npu_inst_pe_1_6_4_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_6_4_n101), 
        .CK(npu_inst_pe_1_6_4_net3103), .RN(npu_inst_pe_1_6_4_n9), .Q(
        npu_inst_pe_1_6_4_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_6_4_n86), 
        .CK(npu_inst_pe_1_6_4_net3103), .RN(npu_inst_pe_1_6_4_n9), .Q(
        npu_inst_pe_1_6_4_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_6_4_n87), 
        .CK(npu_inst_pe_1_6_4_net3103), .RN(npu_inst_pe_1_6_4_n9), .Q(
        npu_inst_pe_1_6_4_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_6_4_n88), 
        .CK(npu_inst_pe_1_6_4_net3103), .RN(npu_inst_pe_1_6_4_n10), .Q(
        npu_inst_pe_1_6_4_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_6_4_n89), 
        .CK(npu_inst_pe_1_6_4_net3103), .RN(npu_inst_pe_1_6_4_n10), .Q(
        npu_inst_pe_1_6_4_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_6_4_n90), 
        .CK(npu_inst_pe_1_6_4_net3103), .RN(npu_inst_pe_1_6_4_n10), .Q(
        npu_inst_pe_1_6_4_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_6_4_n91), 
        .CK(npu_inst_pe_1_6_4_net3103), .RN(npu_inst_pe_1_6_4_n10), .Q(
        npu_inst_pe_1_6_4_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_6_4_n92), 
        .CK(npu_inst_pe_1_6_4_net3103), .RN(npu_inst_pe_1_6_4_n10), .Q(
        npu_inst_pe_1_6_4_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_6_4_n93), 
        .CK(npu_inst_pe_1_6_4_net3103), .RN(npu_inst_pe_1_6_4_n10), .Q(
        npu_inst_pe_1_6_4_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_6_4_n94), 
        .CK(npu_inst_pe_1_6_4_net3103), .RN(npu_inst_pe_1_6_4_n10), .Q(
        npu_inst_pe_1_6_4_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_6_4_n95), 
        .CK(npu_inst_pe_1_6_4_net3103), .RN(npu_inst_pe_1_6_4_n10), .Q(
        npu_inst_pe_1_6_4_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_6_4_n96), 
        .CK(npu_inst_pe_1_6_4_net3103), .RN(npu_inst_pe_1_6_4_n10), .Q(
        npu_inst_pe_1_6_4_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_6_4_n97), 
        .CK(npu_inst_pe_1_6_4_net3103), .RN(npu_inst_pe_1_6_4_n10), .Q(
        npu_inst_pe_1_6_4_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_6_4_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_6_4_N84), .SE(1'b0), .GCK(npu_inst_pe_1_6_4_net3097) );
  CLKGATETST_X1 npu_inst_pe_1_6_4_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n62), .SE(1'b0), .GCK(npu_inst_pe_1_6_4_net3103) );
  MUX2_X1 npu_inst_pe_1_6_5_U162 ( .A(npu_inst_pe_1_6_5_n32), .B(
        npu_inst_pe_1_6_5_n29), .S(npu_inst_pe_1_6_5_n8), .Z(
        npu_inst_pe_1_6_5_N93) );
  MUX2_X1 npu_inst_pe_1_6_5_U161 ( .A(npu_inst_pe_1_6_5_n31), .B(
        npu_inst_pe_1_6_5_n30), .S(npu_inst_pe_1_6_5_n6), .Z(
        npu_inst_pe_1_6_5_n32) );
  MUX2_X1 npu_inst_pe_1_6_5_U160 ( .A(npu_inst_pe_1_6_5_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_6_5_int_q_reg_v_1__0_), .S(npu_inst_pe_1_6_5_n4), .Z(
        npu_inst_pe_1_6_5_n31) );
  MUX2_X1 npu_inst_pe_1_6_5_U159 ( .A(npu_inst_pe_1_6_5_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_6_5_int_q_reg_v_3__0_), .S(npu_inst_pe_1_6_5_n4), .Z(
        npu_inst_pe_1_6_5_n30) );
  MUX2_X1 npu_inst_pe_1_6_5_U158 ( .A(npu_inst_pe_1_6_5_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_6_5_int_q_reg_v_5__0_), .S(npu_inst_pe_1_6_5_n4), .Z(
        npu_inst_pe_1_6_5_n29) );
  MUX2_X1 npu_inst_pe_1_6_5_U157 ( .A(npu_inst_pe_1_6_5_n28), .B(
        npu_inst_pe_1_6_5_n23), .S(npu_inst_pe_1_6_5_n8), .Z(
        npu_inst_pe_1_6_5_N94) );
  MUX2_X1 npu_inst_pe_1_6_5_U156 ( .A(npu_inst_pe_1_6_5_n25), .B(
        npu_inst_pe_1_6_5_n24), .S(npu_inst_pe_1_6_5_n6), .Z(
        npu_inst_pe_1_6_5_n28) );
  MUX2_X1 npu_inst_pe_1_6_5_U155 ( .A(npu_inst_pe_1_6_5_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_6_5_int_q_reg_v_1__1_), .S(npu_inst_pe_1_6_5_n4), .Z(
        npu_inst_pe_1_6_5_n25) );
  MUX2_X1 npu_inst_pe_1_6_5_U154 ( .A(npu_inst_pe_1_6_5_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_6_5_int_q_reg_v_3__1_), .S(npu_inst_pe_1_6_5_n4), .Z(
        npu_inst_pe_1_6_5_n24) );
  MUX2_X1 npu_inst_pe_1_6_5_U153 ( .A(npu_inst_pe_1_6_5_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_6_5_int_q_reg_v_5__1_), .S(npu_inst_pe_1_6_5_n4), .Z(
        npu_inst_pe_1_6_5_n23) );
  MUX2_X1 npu_inst_pe_1_6_5_U152 ( .A(npu_inst_pe_1_6_5_n22), .B(
        npu_inst_pe_1_6_5_n19), .S(npu_inst_pe_1_6_5_n8), .Z(
        npu_inst_int_data_x_6__5__1_) );
  MUX2_X1 npu_inst_pe_1_6_5_U151 ( .A(npu_inst_pe_1_6_5_n21), .B(
        npu_inst_pe_1_6_5_n20), .S(npu_inst_pe_1_6_5_n6), .Z(
        npu_inst_pe_1_6_5_n22) );
  MUX2_X1 npu_inst_pe_1_6_5_U150 ( .A(npu_inst_pe_1_6_5_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_6_5_int_q_reg_h_1__1_), .S(npu_inst_pe_1_6_5_n4), .Z(
        npu_inst_pe_1_6_5_n21) );
  MUX2_X1 npu_inst_pe_1_6_5_U149 ( .A(npu_inst_pe_1_6_5_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_6_5_int_q_reg_h_3__1_), .S(npu_inst_pe_1_6_5_n4), .Z(
        npu_inst_pe_1_6_5_n20) );
  MUX2_X1 npu_inst_pe_1_6_5_U148 ( .A(npu_inst_pe_1_6_5_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_6_5_int_q_reg_h_5__1_), .S(npu_inst_pe_1_6_5_n4), .Z(
        npu_inst_pe_1_6_5_n19) );
  MUX2_X1 npu_inst_pe_1_6_5_U147 ( .A(npu_inst_pe_1_6_5_n18), .B(
        npu_inst_pe_1_6_5_n15), .S(npu_inst_pe_1_6_5_n8), .Z(
        npu_inst_int_data_x_6__5__0_) );
  MUX2_X1 npu_inst_pe_1_6_5_U146 ( .A(npu_inst_pe_1_6_5_n17), .B(
        npu_inst_pe_1_6_5_n16), .S(npu_inst_pe_1_6_5_n6), .Z(
        npu_inst_pe_1_6_5_n18) );
  MUX2_X1 npu_inst_pe_1_6_5_U145 ( .A(npu_inst_pe_1_6_5_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_6_5_int_q_reg_h_1__0_), .S(npu_inst_pe_1_6_5_n4), .Z(
        npu_inst_pe_1_6_5_n17) );
  MUX2_X1 npu_inst_pe_1_6_5_U144 ( .A(npu_inst_pe_1_6_5_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_6_5_int_q_reg_h_3__0_), .S(npu_inst_pe_1_6_5_n4), .Z(
        npu_inst_pe_1_6_5_n16) );
  MUX2_X1 npu_inst_pe_1_6_5_U143 ( .A(npu_inst_pe_1_6_5_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_6_5_int_q_reg_h_5__0_), .S(npu_inst_pe_1_6_5_n4), .Z(
        npu_inst_pe_1_6_5_n15) );
  XOR2_X1 npu_inst_pe_1_6_5_U142 ( .A(npu_inst_pe_1_6_5_int_data_0_), .B(
        npu_inst_pe_1_6_5_int_q_acc_0_), .Z(npu_inst_pe_1_6_5_N73) );
  AND2_X1 npu_inst_pe_1_6_5_U141 ( .A1(npu_inst_pe_1_6_5_int_q_acc_0_), .A2(
        npu_inst_pe_1_6_5_int_data_0_), .ZN(npu_inst_pe_1_6_5_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_6_5_U140 ( .A(npu_inst_pe_1_6_5_int_q_acc_0_), .B(
        npu_inst_pe_1_6_5_n13), .ZN(npu_inst_pe_1_6_5_N65) );
  OR2_X1 npu_inst_pe_1_6_5_U139 ( .A1(npu_inst_pe_1_6_5_n13), .A2(
        npu_inst_pe_1_6_5_int_q_acc_0_), .ZN(npu_inst_pe_1_6_5_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_6_5_U138 ( .A(npu_inst_pe_1_6_5_int_q_acc_2_), .B(
        npu_inst_pe_1_6_5_add_79_carry_2_), .Z(npu_inst_pe_1_6_5_N75) );
  AND2_X1 npu_inst_pe_1_6_5_U137 ( .A1(npu_inst_pe_1_6_5_add_79_carry_2_), 
        .A2(npu_inst_pe_1_6_5_int_q_acc_2_), .ZN(
        npu_inst_pe_1_6_5_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_6_5_U136 ( .A(npu_inst_pe_1_6_5_int_q_acc_3_), .B(
        npu_inst_pe_1_6_5_add_79_carry_3_), .Z(npu_inst_pe_1_6_5_N76) );
  AND2_X1 npu_inst_pe_1_6_5_U135 ( .A1(npu_inst_pe_1_6_5_add_79_carry_3_), 
        .A2(npu_inst_pe_1_6_5_int_q_acc_3_), .ZN(
        npu_inst_pe_1_6_5_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_6_5_U134 ( .A(npu_inst_pe_1_6_5_int_q_acc_4_), .B(
        npu_inst_pe_1_6_5_add_79_carry_4_), .Z(npu_inst_pe_1_6_5_N77) );
  AND2_X1 npu_inst_pe_1_6_5_U133 ( .A1(npu_inst_pe_1_6_5_add_79_carry_4_), 
        .A2(npu_inst_pe_1_6_5_int_q_acc_4_), .ZN(
        npu_inst_pe_1_6_5_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_6_5_U132 ( .A(npu_inst_pe_1_6_5_int_q_acc_5_), .B(
        npu_inst_pe_1_6_5_add_79_carry_5_), .Z(npu_inst_pe_1_6_5_N78) );
  AND2_X1 npu_inst_pe_1_6_5_U131 ( .A1(npu_inst_pe_1_6_5_add_79_carry_5_), 
        .A2(npu_inst_pe_1_6_5_int_q_acc_5_), .ZN(
        npu_inst_pe_1_6_5_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_6_5_U130 ( .A(npu_inst_pe_1_6_5_int_q_acc_6_), .B(
        npu_inst_pe_1_6_5_add_79_carry_6_), .Z(npu_inst_pe_1_6_5_N79) );
  AND2_X1 npu_inst_pe_1_6_5_U129 ( .A1(npu_inst_pe_1_6_5_add_79_carry_6_), 
        .A2(npu_inst_pe_1_6_5_int_q_acc_6_), .ZN(
        npu_inst_pe_1_6_5_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_6_5_U128 ( .A(npu_inst_pe_1_6_5_int_q_acc_7_), .B(
        npu_inst_pe_1_6_5_add_79_carry_7_), .Z(npu_inst_pe_1_6_5_N80) );
  XNOR2_X1 npu_inst_pe_1_6_5_U127 ( .A(npu_inst_pe_1_6_5_sub_77_carry_2_), .B(
        npu_inst_pe_1_6_5_int_q_acc_2_), .ZN(npu_inst_pe_1_6_5_N67) );
  OR2_X1 npu_inst_pe_1_6_5_U126 ( .A1(npu_inst_pe_1_6_5_int_q_acc_2_), .A2(
        npu_inst_pe_1_6_5_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_6_5_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_6_5_U125 ( .A(npu_inst_pe_1_6_5_sub_77_carry_3_), .B(
        npu_inst_pe_1_6_5_int_q_acc_3_), .ZN(npu_inst_pe_1_6_5_N68) );
  OR2_X1 npu_inst_pe_1_6_5_U124 ( .A1(npu_inst_pe_1_6_5_int_q_acc_3_), .A2(
        npu_inst_pe_1_6_5_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_6_5_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_6_5_U123 ( .A(npu_inst_pe_1_6_5_sub_77_carry_4_), .B(
        npu_inst_pe_1_6_5_int_q_acc_4_), .ZN(npu_inst_pe_1_6_5_N69) );
  OR2_X1 npu_inst_pe_1_6_5_U122 ( .A1(npu_inst_pe_1_6_5_int_q_acc_4_), .A2(
        npu_inst_pe_1_6_5_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_6_5_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_6_5_U121 ( .A(npu_inst_pe_1_6_5_sub_77_carry_5_), .B(
        npu_inst_pe_1_6_5_int_q_acc_5_), .ZN(npu_inst_pe_1_6_5_N70) );
  OR2_X1 npu_inst_pe_1_6_5_U120 ( .A1(npu_inst_pe_1_6_5_int_q_acc_5_), .A2(
        npu_inst_pe_1_6_5_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_6_5_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_6_5_U119 ( .A(npu_inst_pe_1_6_5_sub_77_carry_6_), .B(
        npu_inst_pe_1_6_5_int_q_acc_6_), .ZN(npu_inst_pe_1_6_5_N71) );
  OR2_X1 npu_inst_pe_1_6_5_U118 ( .A1(npu_inst_pe_1_6_5_int_q_acc_6_), .A2(
        npu_inst_pe_1_6_5_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_6_5_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_6_5_U117 ( .A(npu_inst_pe_1_6_5_int_q_acc_7_), .B(
        npu_inst_pe_1_6_5_sub_77_carry_7_), .ZN(npu_inst_pe_1_6_5_N72) );
  INV_X1 npu_inst_pe_1_6_5_U116 ( .A(npu_inst_n75), .ZN(npu_inst_pe_1_6_5_n7)
         );
  INV_X1 npu_inst_pe_1_6_5_U115 ( .A(npu_inst_pe_1_6_5_n7), .ZN(
        npu_inst_pe_1_6_5_n6) );
  INV_X1 npu_inst_pe_1_6_5_U114 ( .A(npu_inst_n53), .ZN(npu_inst_pe_1_6_5_n3)
         );
  AOI22_X1 npu_inst_pe_1_6_5_U113 ( .A1(npu_inst_int_data_y_7__5__0_), .A2(
        npu_inst_pe_1_6_5_n58), .B1(npu_inst_pe_1_6_5_n114), .B2(
        npu_inst_pe_1_6_5_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_6_5_n57) );
  INV_X1 npu_inst_pe_1_6_5_U112 ( .A(npu_inst_pe_1_6_5_n57), .ZN(
        npu_inst_pe_1_6_5_n108) );
  AOI22_X1 npu_inst_pe_1_6_5_U111 ( .A1(npu_inst_int_data_y_7__5__0_), .A2(
        npu_inst_pe_1_6_5_n54), .B1(npu_inst_pe_1_6_5_n115), .B2(
        npu_inst_pe_1_6_5_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_6_5_n53) );
  INV_X1 npu_inst_pe_1_6_5_U110 ( .A(npu_inst_pe_1_6_5_n53), .ZN(
        npu_inst_pe_1_6_5_n109) );
  AOI22_X1 npu_inst_pe_1_6_5_U107 ( .A1(npu_inst_int_data_y_7__5__0_), .A2(
        npu_inst_pe_1_6_5_n50), .B1(npu_inst_pe_1_6_5_n116), .B2(
        npu_inst_pe_1_6_5_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_6_5_n49) );
  INV_X1 npu_inst_pe_1_6_5_U106 ( .A(npu_inst_pe_1_6_5_n49), .ZN(
        npu_inst_pe_1_6_5_n110) );
  AOI22_X1 npu_inst_pe_1_6_5_U105 ( .A1(npu_inst_int_data_y_7__5__0_), .A2(
        npu_inst_pe_1_6_5_n46), .B1(npu_inst_pe_1_6_5_n117), .B2(
        npu_inst_pe_1_6_5_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_6_5_n45) );
  INV_X1 npu_inst_pe_1_6_5_U104 ( .A(npu_inst_pe_1_6_5_n45), .ZN(
        npu_inst_pe_1_6_5_n111) );
  AOI22_X1 npu_inst_pe_1_6_5_U103 ( .A1(npu_inst_int_data_y_7__5__0_), .A2(
        npu_inst_pe_1_6_5_n42), .B1(npu_inst_pe_1_6_5_n119), .B2(
        npu_inst_pe_1_6_5_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_6_5_n41) );
  INV_X1 npu_inst_pe_1_6_5_U102 ( .A(npu_inst_pe_1_6_5_n41), .ZN(
        npu_inst_pe_1_6_5_n112) );
  AOI22_X1 npu_inst_pe_1_6_5_U101 ( .A1(npu_inst_int_data_y_7__5__1_), .A2(
        npu_inst_pe_1_6_5_n58), .B1(npu_inst_pe_1_6_5_n114), .B2(
        npu_inst_pe_1_6_5_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_6_5_n59) );
  INV_X1 npu_inst_pe_1_6_5_U100 ( .A(npu_inst_pe_1_6_5_n59), .ZN(
        npu_inst_pe_1_6_5_n102) );
  AOI22_X1 npu_inst_pe_1_6_5_U99 ( .A1(npu_inst_int_data_y_7__5__1_), .A2(
        npu_inst_pe_1_6_5_n54), .B1(npu_inst_pe_1_6_5_n115), .B2(
        npu_inst_pe_1_6_5_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_6_5_n55) );
  INV_X1 npu_inst_pe_1_6_5_U98 ( .A(npu_inst_pe_1_6_5_n55), .ZN(
        npu_inst_pe_1_6_5_n103) );
  AOI22_X1 npu_inst_pe_1_6_5_U97 ( .A1(npu_inst_int_data_y_7__5__1_), .A2(
        npu_inst_pe_1_6_5_n50), .B1(npu_inst_pe_1_6_5_n116), .B2(
        npu_inst_pe_1_6_5_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_6_5_n51) );
  INV_X1 npu_inst_pe_1_6_5_U96 ( .A(npu_inst_pe_1_6_5_n51), .ZN(
        npu_inst_pe_1_6_5_n104) );
  AOI22_X1 npu_inst_pe_1_6_5_U95 ( .A1(npu_inst_int_data_y_7__5__1_), .A2(
        npu_inst_pe_1_6_5_n46), .B1(npu_inst_pe_1_6_5_n117), .B2(
        npu_inst_pe_1_6_5_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_6_5_n47) );
  INV_X1 npu_inst_pe_1_6_5_U94 ( .A(npu_inst_pe_1_6_5_n47), .ZN(
        npu_inst_pe_1_6_5_n105) );
  AOI22_X1 npu_inst_pe_1_6_5_U93 ( .A1(npu_inst_int_data_y_7__5__1_), .A2(
        npu_inst_pe_1_6_5_n42), .B1(npu_inst_pe_1_6_5_n119), .B2(
        npu_inst_pe_1_6_5_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_6_5_n43) );
  INV_X1 npu_inst_pe_1_6_5_U92 ( .A(npu_inst_pe_1_6_5_n43), .ZN(
        npu_inst_pe_1_6_5_n106) );
  AOI22_X1 npu_inst_pe_1_6_5_U91 ( .A1(npu_inst_pe_1_6_5_n38), .A2(
        npu_inst_int_data_y_7__5__1_), .B1(npu_inst_pe_1_6_5_n118), .B2(
        npu_inst_pe_1_6_5_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_6_5_n39) );
  INV_X1 npu_inst_pe_1_6_5_U90 ( .A(npu_inst_pe_1_6_5_n39), .ZN(
        npu_inst_pe_1_6_5_n107) );
  AOI22_X1 npu_inst_pe_1_6_5_U89 ( .A1(npu_inst_pe_1_6_5_n38), .A2(
        npu_inst_int_data_y_7__5__0_), .B1(npu_inst_pe_1_6_5_n118), .B2(
        npu_inst_pe_1_6_5_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_6_5_n37) );
  INV_X1 npu_inst_pe_1_6_5_U88 ( .A(npu_inst_pe_1_6_5_n37), .ZN(
        npu_inst_pe_1_6_5_n113) );
  NAND2_X1 npu_inst_pe_1_6_5_U87 ( .A1(npu_inst_pe_1_6_5_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_6_5_n60), .ZN(npu_inst_pe_1_6_5_n74) );
  OAI21_X1 npu_inst_pe_1_6_5_U86 ( .B1(npu_inst_pe_1_6_5_n63), .B2(
        npu_inst_pe_1_6_5_n60), .A(npu_inst_pe_1_6_5_n74), .ZN(
        npu_inst_pe_1_6_5_n97) );
  NAND2_X1 npu_inst_pe_1_6_5_U85 ( .A1(npu_inst_pe_1_6_5_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_6_5_n60), .ZN(npu_inst_pe_1_6_5_n73) );
  OAI21_X1 npu_inst_pe_1_6_5_U84 ( .B1(npu_inst_pe_1_6_5_n61), .B2(
        npu_inst_pe_1_6_5_n60), .A(npu_inst_pe_1_6_5_n73), .ZN(
        npu_inst_pe_1_6_5_n96) );
  NAND2_X1 npu_inst_pe_1_6_5_U83 ( .A1(npu_inst_pe_1_6_5_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_6_5_n56), .ZN(npu_inst_pe_1_6_5_n72) );
  OAI21_X1 npu_inst_pe_1_6_5_U82 ( .B1(npu_inst_pe_1_6_5_n63), .B2(
        npu_inst_pe_1_6_5_n56), .A(npu_inst_pe_1_6_5_n72), .ZN(
        npu_inst_pe_1_6_5_n95) );
  NAND2_X1 npu_inst_pe_1_6_5_U81 ( .A1(npu_inst_pe_1_6_5_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_6_5_n56), .ZN(npu_inst_pe_1_6_5_n71) );
  OAI21_X1 npu_inst_pe_1_6_5_U80 ( .B1(npu_inst_pe_1_6_5_n61), .B2(
        npu_inst_pe_1_6_5_n56), .A(npu_inst_pe_1_6_5_n71), .ZN(
        npu_inst_pe_1_6_5_n94) );
  NAND2_X1 npu_inst_pe_1_6_5_U79 ( .A1(npu_inst_pe_1_6_5_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_6_5_n52), .ZN(npu_inst_pe_1_6_5_n70) );
  OAI21_X1 npu_inst_pe_1_6_5_U78 ( .B1(npu_inst_pe_1_6_5_n63), .B2(
        npu_inst_pe_1_6_5_n52), .A(npu_inst_pe_1_6_5_n70), .ZN(
        npu_inst_pe_1_6_5_n93) );
  NAND2_X1 npu_inst_pe_1_6_5_U77 ( .A1(npu_inst_pe_1_6_5_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_6_5_n52), .ZN(npu_inst_pe_1_6_5_n69) );
  OAI21_X1 npu_inst_pe_1_6_5_U76 ( .B1(npu_inst_pe_1_6_5_n61), .B2(
        npu_inst_pe_1_6_5_n52), .A(npu_inst_pe_1_6_5_n69), .ZN(
        npu_inst_pe_1_6_5_n92) );
  NAND2_X1 npu_inst_pe_1_6_5_U75 ( .A1(npu_inst_pe_1_6_5_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_6_5_n48), .ZN(npu_inst_pe_1_6_5_n68) );
  OAI21_X1 npu_inst_pe_1_6_5_U74 ( .B1(npu_inst_pe_1_6_5_n63), .B2(
        npu_inst_pe_1_6_5_n48), .A(npu_inst_pe_1_6_5_n68), .ZN(
        npu_inst_pe_1_6_5_n91) );
  NAND2_X1 npu_inst_pe_1_6_5_U73 ( .A1(npu_inst_pe_1_6_5_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_6_5_n48), .ZN(npu_inst_pe_1_6_5_n67) );
  OAI21_X1 npu_inst_pe_1_6_5_U72 ( .B1(npu_inst_pe_1_6_5_n61), .B2(
        npu_inst_pe_1_6_5_n48), .A(npu_inst_pe_1_6_5_n67), .ZN(
        npu_inst_pe_1_6_5_n90) );
  NAND2_X1 npu_inst_pe_1_6_5_U71 ( .A1(npu_inst_pe_1_6_5_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_6_5_n44), .ZN(npu_inst_pe_1_6_5_n66) );
  OAI21_X1 npu_inst_pe_1_6_5_U70 ( .B1(npu_inst_pe_1_6_5_n63), .B2(
        npu_inst_pe_1_6_5_n44), .A(npu_inst_pe_1_6_5_n66), .ZN(
        npu_inst_pe_1_6_5_n89) );
  NAND2_X1 npu_inst_pe_1_6_5_U69 ( .A1(npu_inst_pe_1_6_5_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_6_5_n44), .ZN(npu_inst_pe_1_6_5_n65) );
  OAI21_X1 npu_inst_pe_1_6_5_U68 ( .B1(npu_inst_pe_1_6_5_n61), .B2(
        npu_inst_pe_1_6_5_n44), .A(npu_inst_pe_1_6_5_n65), .ZN(
        npu_inst_pe_1_6_5_n88) );
  NAND2_X1 npu_inst_pe_1_6_5_U67 ( .A1(npu_inst_pe_1_6_5_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_6_5_n40), .ZN(npu_inst_pe_1_6_5_n64) );
  OAI21_X1 npu_inst_pe_1_6_5_U66 ( .B1(npu_inst_pe_1_6_5_n63), .B2(
        npu_inst_pe_1_6_5_n40), .A(npu_inst_pe_1_6_5_n64), .ZN(
        npu_inst_pe_1_6_5_n87) );
  NAND2_X1 npu_inst_pe_1_6_5_U65 ( .A1(npu_inst_pe_1_6_5_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_6_5_n40), .ZN(npu_inst_pe_1_6_5_n62) );
  OAI21_X1 npu_inst_pe_1_6_5_U64 ( .B1(npu_inst_pe_1_6_5_n61), .B2(
        npu_inst_pe_1_6_5_n40), .A(npu_inst_pe_1_6_5_n62), .ZN(
        npu_inst_pe_1_6_5_n86) );
  AND2_X1 npu_inst_pe_1_6_5_U63 ( .A1(npu_inst_pe_1_6_5_N93), .A2(npu_inst_n53), .ZN(npu_inst_int_data_y_6__5__0_) );
  AND2_X1 npu_inst_pe_1_6_5_U62 ( .A1(npu_inst_n53), .A2(npu_inst_pe_1_6_5_N94), .ZN(npu_inst_int_data_y_6__5__1_) );
  NOR3_X1 npu_inst_pe_1_6_5_U61 ( .A1(npu_inst_pe_1_6_5_n26), .A2(npu_inst_n53), .A3(npu_inst_int_ckg[10]), .ZN(npu_inst_pe_1_6_5_n85) );
  OR2_X1 npu_inst_pe_1_6_5_U60 ( .A1(npu_inst_pe_1_6_5_n85), .A2(
        npu_inst_pe_1_6_5_n2), .ZN(npu_inst_pe_1_6_5_N84) );
  AND2_X1 npu_inst_pe_1_6_5_U59 ( .A1(npu_inst_pe_1_6_5_int_q_acc_0_), .A2(
        npu_inst_pe_1_6_5_n1), .ZN(npu_inst_int_data_res_6__5__0_) );
  AND2_X1 npu_inst_pe_1_6_5_U58 ( .A1(npu_inst_pe_1_6_5_n2), .A2(
        npu_inst_pe_1_6_5_int_q_acc_7_), .ZN(npu_inst_int_data_res_6__5__7_)
         );
  AND2_X1 npu_inst_pe_1_6_5_U57 ( .A1(npu_inst_pe_1_6_5_int_q_acc_1_), .A2(
        npu_inst_pe_1_6_5_n1), .ZN(npu_inst_int_data_res_6__5__1_) );
  AND2_X1 npu_inst_pe_1_6_5_U56 ( .A1(npu_inst_pe_1_6_5_int_q_acc_2_), .A2(
        npu_inst_pe_1_6_5_n1), .ZN(npu_inst_int_data_res_6__5__2_) );
  AND2_X1 npu_inst_pe_1_6_5_U55 ( .A1(npu_inst_pe_1_6_5_int_q_acc_3_), .A2(
        npu_inst_pe_1_6_5_n2), .ZN(npu_inst_int_data_res_6__5__3_) );
  AND2_X1 npu_inst_pe_1_6_5_U54 ( .A1(npu_inst_pe_1_6_5_int_q_acc_4_), .A2(
        npu_inst_pe_1_6_5_n2), .ZN(npu_inst_int_data_res_6__5__4_) );
  AND2_X1 npu_inst_pe_1_6_5_U53 ( .A1(npu_inst_pe_1_6_5_int_q_acc_5_), .A2(
        npu_inst_pe_1_6_5_n2), .ZN(npu_inst_int_data_res_6__5__5_) );
  AND2_X1 npu_inst_pe_1_6_5_U52 ( .A1(npu_inst_pe_1_6_5_int_q_acc_6_), .A2(
        npu_inst_pe_1_6_5_n2), .ZN(npu_inst_int_data_res_6__5__6_) );
  AOI222_X1 npu_inst_pe_1_6_5_U51 ( .A1(npu_inst_int_data_res_7__5__0_), .A2(
        npu_inst_pe_1_6_5_n1), .B1(npu_inst_pe_1_6_5_N73), .B2(
        npu_inst_pe_1_6_5_n76), .C1(npu_inst_pe_1_6_5_N65), .C2(
        npu_inst_pe_1_6_5_n77), .ZN(npu_inst_pe_1_6_5_n84) );
  INV_X1 npu_inst_pe_1_6_5_U50 ( .A(npu_inst_pe_1_6_5_n84), .ZN(
        npu_inst_pe_1_6_5_n101) );
  AOI222_X1 npu_inst_pe_1_6_5_U49 ( .A1(npu_inst_int_data_res_7__5__7_), .A2(
        npu_inst_pe_1_6_5_n1), .B1(npu_inst_pe_1_6_5_N80), .B2(
        npu_inst_pe_1_6_5_n76), .C1(npu_inst_pe_1_6_5_N72), .C2(
        npu_inst_pe_1_6_5_n77), .ZN(npu_inst_pe_1_6_5_n75) );
  INV_X1 npu_inst_pe_1_6_5_U48 ( .A(npu_inst_pe_1_6_5_n75), .ZN(
        npu_inst_pe_1_6_5_n33) );
  AOI222_X1 npu_inst_pe_1_6_5_U47 ( .A1(npu_inst_int_data_res_7__5__1_), .A2(
        npu_inst_pe_1_6_5_n1), .B1(npu_inst_pe_1_6_5_N74), .B2(
        npu_inst_pe_1_6_5_n76), .C1(npu_inst_pe_1_6_5_N66), .C2(
        npu_inst_pe_1_6_5_n77), .ZN(npu_inst_pe_1_6_5_n83) );
  INV_X1 npu_inst_pe_1_6_5_U46 ( .A(npu_inst_pe_1_6_5_n83), .ZN(
        npu_inst_pe_1_6_5_n100) );
  AOI222_X1 npu_inst_pe_1_6_5_U45 ( .A1(npu_inst_int_data_res_7__5__2_), .A2(
        npu_inst_pe_1_6_5_n1), .B1(npu_inst_pe_1_6_5_N75), .B2(
        npu_inst_pe_1_6_5_n76), .C1(npu_inst_pe_1_6_5_N67), .C2(
        npu_inst_pe_1_6_5_n77), .ZN(npu_inst_pe_1_6_5_n82) );
  INV_X1 npu_inst_pe_1_6_5_U44 ( .A(npu_inst_pe_1_6_5_n82), .ZN(
        npu_inst_pe_1_6_5_n99) );
  AOI222_X1 npu_inst_pe_1_6_5_U43 ( .A1(npu_inst_int_data_res_7__5__3_), .A2(
        npu_inst_pe_1_6_5_n1), .B1(npu_inst_pe_1_6_5_N76), .B2(
        npu_inst_pe_1_6_5_n76), .C1(npu_inst_pe_1_6_5_N68), .C2(
        npu_inst_pe_1_6_5_n77), .ZN(npu_inst_pe_1_6_5_n81) );
  INV_X1 npu_inst_pe_1_6_5_U42 ( .A(npu_inst_pe_1_6_5_n81), .ZN(
        npu_inst_pe_1_6_5_n98) );
  AOI222_X1 npu_inst_pe_1_6_5_U41 ( .A1(npu_inst_int_data_res_7__5__4_), .A2(
        npu_inst_pe_1_6_5_n1), .B1(npu_inst_pe_1_6_5_N77), .B2(
        npu_inst_pe_1_6_5_n76), .C1(npu_inst_pe_1_6_5_N69), .C2(
        npu_inst_pe_1_6_5_n77), .ZN(npu_inst_pe_1_6_5_n80) );
  INV_X1 npu_inst_pe_1_6_5_U40 ( .A(npu_inst_pe_1_6_5_n80), .ZN(
        npu_inst_pe_1_6_5_n36) );
  AOI222_X1 npu_inst_pe_1_6_5_U39 ( .A1(npu_inst_int_data_res_7__5__5_), .A2(
        npu_inst_pe_1_6_5_n1), .B1(npu_inst_pe_1_6_5_N78), .B2(
        npu_inst_pe_1_6_5_n76), .C1(npu_inst_pe_1_6_5_N70), .C2(
        npu_inst_pe_1_6_5_n77), .ZN(npu_inst_pe_1_6_5_n79) );
  INV_X1 npu_inst_pe_1_6_5_U38 ( .A(npu_inst_pe_1_6_5_n79), .ZN(
        npu_inst_pe_1_6_5_n35) );
  AOI222_X1 npu_inst_pe_1_6_5_U37 ( .A1(npu_inst_int_data_res_7__5__6_), .A2(
        npu_inst_pe_1_6_5_n1), .B1(npu_inst_pe_1_6_5_N79), .B2(
        npu_inst_pe_1_6_5_n76), .C1(npu_inst_pe_1_6_5_N71), .C2(
        npu_inst_pe_1_6_5_n77), .ZN(npu_inst_pe_1_6_5_n78) );
  INV_X1 npu_inst_pe_1_6_5_U36 ( .A(npu_inst_pe_1_6_5_n78), .ZN(
        npu_inst_pe_1_6_5_n34) );
  INV_X1 npu_inst_pe_1_6_5_U35 ( .A(npu_inst_pe_1_6_5_int_data_1_), .ZN(
        npu_inst_pe_1_6_5_n14) );
  AND2_X1 npu_inst_pe_1_6_5_U34 ( .A1(npu_inst_int_data_x_6__5__1_), .A2(
        npu_inst_pe_1_6_5_int_q_weight_1_), .ZN(npu_inst_pe_1_6_5_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_6_5_U33 ( .A1(npu_inst_int_data_x_6__5__0_), .A2(
        npu_inst_pe_1_6_5_int_q_weight_1_), .ZN(npu_inst_pe_1_6_5_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_6_5_U32 ( .A1(npu_inst_n53), .A2(
        npu_inst_int_data_y_7__5__1_), .B1(npu_inst_pe_1_6_5_n3), .B2(
        npu_inst_int_data_x_6__6__1_), .ZN(npu_inst_pe_1_6_5_n63) );
  AOI22_X1 npu_inst_pe_1_6_5_U31 ( .A1(npu_inst_n53), .A2(
        npu_inst_int_data_y_7__5__0_), .B1(npu_inst_pe_1_6_5_n3), .B2(
        npu_inst_int_data_x_6__6__0_), .ZN(npu_inst_pe_1_6_5_n61) );
  INV_X1 npu_inst_pe_1_6_5_U30 ( .A(npu_inst_pe_1_6_5_int_data_0_), .ZN(
        npu_inst_pe_1_6_5_n13) );
  INV_X1 npu_inst_pe_1_6_5_U29 ( .A(npu_inst_n67), .ZN(npu_inst_pe_1_6_5_n5)
         );
  OR3_X1 npu_inst_pe_1_6_5_U28 ( .A1(npu_inst_pe_1_6_5_n6), .A2(
        npu_inst_pe_1_6_5_n8), .A3(npu_inst_pe_1_6_5_n5), .ZN(
        npu_inst_pe_1_6_5_n56) );
  OR3_X1 npu_inst_pe_1_6_5_U27 ( .A1(npu_inst_pe_1_6_5_n5), .A2(
        npu_inst_pe_1_6_5_n8), .A3(npu_inst_pe_1_6_5_n7), .ZN(
        npu_inst_pe_1_6_5_n48) );
  INV_X1 npu_inst_pe_1_6_5_U26 ( .A(npu_inst_pe_1_6_5_n5), .ZN(
        npu_inst_pe_1_6_5_n4) );
  INV_X1 npu_inst_pe_1_6_5_U25 ( .A(npu_inst_n122), .ZN(npu_inst_pe_1_6_5_n12)
         );
  OR3_X1 npu_inst_pe_1_6_5_U24 ( .A1(npu_inst_pe_1_6_5_n4), .A2(
        npu_inst_pe_1_6_5_n8), .A3(npu_inst_pe_1_6_5_n7), .ZN(
        npu_inst_pe_1_6_5_n52) );
  OR3_X1 npu_inst_pe_1_6_5_U23 ( .A1(npu_inst_pe_1_6_5_n6), .A2(
        npu_inst_pe_1_6_5_n8), .A3(npu_inst_pe_1_6_5_n4), .ZN(
        npu_inst_pe_1_6_5_n60) );
  NOR2_X1 npu_inst_pe_1_6_5_U22 ( .A1(npu_inst_pe_1_6_5_n60), .A2(
        npu_inst_pe_1_6_5_n3), .ZN(npu_inst_pe_1_6_5_n58) );
  NOR2_X1 npu_inst_pe_1_6_5_U21 ( .A1(npu_inst_pe_1_6_5_n56), .A2(
        npu_inst_pe_1_6_5_n3), .ZN(npu_inst_pe_1_6_5_n54) );
  NOR2_X1 npu_inst_pe_1_6_5_U20 ( .A1(npu_inst_pe_1_6_5_n52), .A2(
        npu_inst_pe_1_6_5_n3), .ZN(npu_inst_pe_1_6_5_n50) );
  NOR2_X1 npu_inst_pe_1_6_5_U19 ( .A1(npu_inst_pe_1_6_5_n48), .A2(
        npu_inst_pe_1_6_5_n3), .ZN(npu_inst_pe_1_6_5_n46) );
  NOR2_X1 npu_inst_pe_1_6_5_U18 ( .A1(npu_inst_pe_1_6_5_n40), .A2(
        npu_inst_pe_1_6_5_n3), .ZN(npu_inst_pe_1_6_5_n38) );
  NOR2_X1 npu_inst_pe_1_6_5_U17 ( .A1(npu_inst_pe_1_6_5_n44), .A2(
        npu_inst_pe_1_6_5_n3), .ZN(npu_inst_pe_1_6_5_n42) );
  BUF_X1 npu_inst_pe_1_6_5_U16 ( .A(npu_inst_n94), .Z(npu_inst_pe_1_6_5_n8) );
  BUF_X1 npu_inst_pe_1_6_5_U15 ( .A(npu_inst_pe_1_6_5_n12), .Z(
        npu_inst_pe_1_6_5_n11) );
  BUF_X1 npu_inst_pe_1_6_5_U14 ( .A(npu_inst_pe_1_6_5_n12), .Z(
        npu_inst_pe_1_6_5_n10) );
  BUF_X1 npu_inst_pe_1_6_5_U13 ( .A(npu_inst_pe_1_6_5_n12), .Z(
        npu_inst_pe_1_6_5_n9) );
  INV_X1 npu_inst_pe_1_6_5_U12 ( .A(npu_inst_pe_1_6_5_n38), .ZN(
        npu_inst_pe_1_6_5_n118) );
  INV_X1 npu_inst_pe_1_6_5_U11 ( .A(npu_inst_pe_1_6_5_n58), .ZN(
        npu_inst_pe_1_6_5_n114) );
  INV_X1 npu_inst_pe_1_6_5_U10 ( .A(npu_inst_pe_1_6_5_n54), .ZN(
        npu_inst_pe_1_6_5_n115) );
  INV_X1 npu_inst_pe_1_6_5_U9 ( .A(npu_inst_pe_1_6_5_n50), .ZN(
        npu_inst_pe_1_6_5_n116) );
  INV_X1 npu_inst_pe_1_6_5_U8 ( .A(npu_inst_pe_1_6_5_n46), .ZN(
        npu_inst_pe_1_6_5_n117) );
  INV_X1 npu_inst_pe_1_6_5_U7 ( .A(npu_inst_pe_1_6_5_n42), .ZN(
        npu_inst_pe_1_6_5_n119) );
  BUF_X1 npu_inst_pe_1_6_5_U6 ( .A(npu_inst_n12), .Z(npu_inst_pe_1_6_5_n2) );
  BUF_X1 npu_inst_pe_1_6_5_U5 ( .A(npu_inst_n12), .Z(npu_inst_pe_1_6_5_n1) );
  NOR2_X1 npu_inst_pe_1_6_5_U4 ( .A1(npu_inst_pe_1_6_5_int_q_weight_0_), .A2(
        npu_inst_pe_1_6_5_n1), .ZN(npu_inst_pe_1_6_5_n76) );
  NOR2_X1 npu_inst_pe_1_6_5_U3 ( .A1(npu_inst_pe_1_6_5_n27), .A2(
        npu_inst_pe_1_6_5_n1), .ZN(npu_inst_pe_1_6_5_n77) );
  FA_X1 npu_inst_pe_1_6_5_sub_77_U2_1 ( .A(npu_inst_pe_1_6_5_int_q_acc_1_), 
        .B(npu_inst_pe_1_6_5_n14), .CI(npu_inst_pe_1_6_5_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_6_5_sub_77_carry_2_), .S(npu_inst_pe_1_6_5_N66) );
  FA_X1 npu_inst_pe_1_6_5_add_79_U1_1 ( .A(npu_inst_pe_1_6_5_int_q_acc_1_), 
        .B(npu_inst_pe_1_6_5_int_data_1_), .CI(
        npu_inst_pe_1_6_5_add_79_carry_1_), .CO(
        npu_inst_pe_1_6_5_add_79_carry_2_), .S(npu_inst_pe_1_6_5_N74) );
  NAND3_X1 npu_inst_pe_1_6_5_U109 ( .A1(npu_inst_pe_1_6_5_n5), .A2(
        npu_inst_pe_1_6_5_n7), .A3(npu_inst_pe_1_6_5_n8), .ZN(
        npu_inst_pe_1_6_5_n44) );
  NAND3_X1 npu_inst_pe_1_6_5_U108 ( .A1(npu_inst_pe_1_6_5_n4), .A2(
        npu_inst_pe_1_6_5_n7), .A3(npu_inst_pe_1_6_5_n8), .ZN(
        npu_inst_pe_1_6_5_n40) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_6_5_n34), .CK(
        npu_inst_pe_1_6_5_net3074), .RN(npu_inst_pe_1_6_5_n9), .Q(
        npu_inst_pe_1_6_5_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_6_5_n35), .CK(
        npu_inst_pe_1_6_5_net3074), .RN(npu_inst_pe_1_6_5_n9), .Q(
        npu_inst_pe_1_6_5_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_6_5_n36), .CK(
        npu_inst_pe_1_6_5_net3074), .RN(npu_inst_pe_1_6_5_n9), .Q(
        npu_inst_pe_1_6_5_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_6_5_n98), .CK(
        npu_inst_pe_1_6_5_net3074), .RN(npu_inst_pe_1_6_5_n9), .Q(
        npu_inst_pe_1_6_5_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_6_5_n99), .CK(
        npu_inst_pe_1_6_5_net3074), .RN(npu_inst_pe_1_6_5_n9), .Q(
        npu_inst_pe_1_6_5_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_6_5_n100), 
        .CK(npu_inst_pe_1_6_5_net3074), .RN(npu_inst_pe_1_6_5_n9), .Q(
        npu_inst_pe_1_6_5_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_6_5_n33), .CK(
        npu_inst_pe_1_6_5_net3074), .RN(npu_inst_pe_1_6_5_n9), .Q(
        npu_inst_pe_1_6_5_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_6_5_n101), 
        .CK(npu_inst_pe_1_6_5_net3074), .RN(npu_inst_pe_1_6_5_n9), .Q(
        npu_inst_pe_1_6_5_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_weight_reg_0_ ( .D(npu_inst_n108), .CK(
        npu_inst_pe_1_6_5_net3080), .RN(npu_inst_pe_1_6_5_n9), .Q(
        npu_inst_pe_1_6_5_int_q_weight_0_), .QN(npu_inst_pe_1_6_5_n27) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_weight_reg_1_ ( .D(npu_inst_n114), .CK(
        npu_inst_pe_1_6_5_net3080), .RN(npu_inst_pe_1_6_5_n9), .Q(
        npu_inst_pe_1_6_5_int_q_weight_1_), .QN(npu_inst_pe_1_6_5_n26) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_6_5_n113), 
        .CK(npu_inst_pe_1_6_5_net3080), .RN(npu_inst_pe_1_6_5_n9), .Q(
        npu_inst_pe_1_6_5_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_6_5_n107), 
        .CK(npu_inst_pe_1_6_5_net3080), .RN(npu_inst_pe_1_6_5_n9), .Q(
        npu_inst_pe_1_6_5_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_6_5_n112), 
        .CK(npu_inst_pe_1_6_5_net3080), .RN(npu_inst_pe_1_6_5_n10), .Q(
        npu_inst_pe_1_6_5_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_6_5_n106), 
        .CK(npu_inst_pe_1_6_5_net3080), .RN(npu_inst_pe_1_6_5_n10), .Q(
        npu_inst_pe_1_6_5_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_6_5_n111), 
        .CK(npu_inst_pe_1_6_5_net3080), .RN(npu_inst_pe_1_6_5_n10), .Q(
        npu_inst_pe_1_6_5_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_6_5_n105), 
        .CK(npu_inst_pe_1_6_5_net3080), .RN(npu_inst_pe_1_6_5_n10), .Q(
        npu_inst_pe_1_6_5_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_6_5_n110), 
        .CK(npu_inst_pe_1_6_5_net3080), .RN(npu_inst_pe_1_6_5_n10), .Q(
        npu_inst_pe_1_6_5_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_6_5_n104), 
        .CK(npu_inst_pe_1_6_5_net3080), .RN(npu_inst_pe_1_6_5_n10), .Q(
        npu_inst_pe_1_6_5_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_6_5_n109), 
        .CK(npu_inst_pe_1_6_5_net3080), .RN(npu_inst_pe_1_6_5_n10), .Q(
        npu_inst_pe_1_6_5_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_6_5_n103), 
        .CK(npu_inst_pe_1_6_5_net3080), .RN(npu_inst_pe_1_6_5_n10), .Q(
        npu_inst_pe_1_6_5_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_6_5_n108), 
        .CK(npu_inst_pe_1_6_5_net3080), .RN(npu_inst_pe_1_6_5_n10), .Q(
        npu_inst_pe_1_6_5_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_6_5_n102), 
        .CK(npu_inst_pe_1_6_5_net3080), .RN(npu_inst_pe_1_6_5_n10), .Q(
        npu_inst_pe_1_6_5_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_6_5_n86), 
        .CK(npu_inst_pe_1_6_5_net3080), .RN(npu_inst_pe_1_6_5_n10), .Q(
        npu_inst_pe_1_6_5_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_6_5_n87), 
        .CK(npu_inst_pe_1_6_5_net3080), .RN(npu_inst_pe_1_6_5_n10), .Q(
        npu_inst_pe_1_6_5_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_6_5_n88), 
        .CK(npu_inst_pe_1_6_5_net3080), .RN(npu_inst_pe_1_6_5_n11), .Q(
        npu_inst_pe_1_6_5_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_6_5_n89), 
        .CK(npu_inst_pe_1_6_5_net3080), .RN(npu_inst_pe_1_6_5_n11), .Q(
        npu_inst_pe_1_6_5_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_6_5_n90), 
        .CK(npu_inst_pe_1_6_5_net3080), .RN(npu_inst_pe_1_6_5_n11), .Q(
        npu_inst_pe_1_6_5_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_6_5_n91), 
        .CK(npu_inst_pe_1_6_5_net3080), .RN(npu_inst_pe_1_6_5_n11), .Q(
        npu_inst_pe_1_6_5_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_6_5_n92), 
        .CK(npu_inst_pe_1_6_5_net3080), .RN(npu_inst_pe_1_6_5_n11), .Q(
        npu_inst_pe_1_6_5_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_6_5_n93), 
        .CK(npu_inst_pe_1_6_5_net3080), .RN(npu_inst_pe_1_6_5_n11), .Q(
        npu_inst_pe_1_6_5_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_6_5_n94), 
        .CK(npu_inst_pe_1_6_5_net3080), .RN(npu_inst_pe_1_6_5_n11), .Q(
        npu_inst_pe_1_6_5_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_6_5_n95), 
        .CK(npu_inst_pe_1_6_5_net3080), .RN(npu_inst_pe_1_6_5_n11), .Q(
        npu_inst_pe_1_6_5_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_6_5_n96), 
        .CK(npu_inst_pe_1_6_5_net3080), .RN(npu_inst_pe_1_6_5_n11), .Q(
        npu_inst_pe_1_6_5_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_6_5_n97), 
        .CK(npu_inst_pe_1_6_5_net3080), .RN(npu_inst_pe_1_6_5_n11), .Q(
        npu_inst_pe_1_6_5_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_6_5_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_6_5_N84), .SE(1'b0), .GCK(npu_inst_pe_1_6_5_net3074) );
  CLKGATETST_X1 npu_inst_pe_1_6_5_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n61), .SE(1'b0), .GCK(npu_inst_pe_1_6_5_net3080) );
  MUX2_X1 npu_inst_pe_1_6_6_U162 ( .A(npu_inst_pe_1_6_6_n32), .B(
        npu_inst_pe_1_6_6_n29), .S(npu_inst_pe_1_6_6_n8), .Z(
        npu_inst_pe_1_6_6_N93) );
  MUX2_X1 npu_inst_pe_1_6_6_U161 ( .A(npu_inst_pe_1_6_6_n31), .B(
        npu_inst_pe_1_6_6_n30), .S(npu_inst_pe_1_6_6_n6), .Z(
        npu_inst_pe_1_6_6_n32) );
  MUX2_X1 npu_inst_pe_1_6_6_U160 ( .A(npu_inst_pe_1_6_6_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_6_6_int_q_reg_v_1__0_), .S(npu_inst_pe_1_6_6_n4), .Z(
        npu_inst_pe_1_6_6_n31) );
  MUX2_X1 npu_inst_pe_1_6_6_U159 ( .A(npu_inst_pe_1_6_6_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_6_6_int_q_reg_v_3__0_), .S(npu_inst_pe_1_6_6_n4), .Z(
        npu_inst_pe_1_6_6_n30) );
  MUX2_X1 npu_inst_pe_1_6_6_U158 ( .A(npu_inst_pe_1_6_6_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_6_6_int_q_reg_v_5__0_), .S(npu_inst_pe_1_6_6_n4), .Z(
        npu_inst_pe_1_6_6_n29) );
  MUX2_X1 npu_inst_pe_1_6_6_U157 ( .A(npu_inst_pe_1_6_6_n28), .B(
        npu_inst_pe_1_6_6_n23), .S(npu_inst_pe_1_6_6_n8), .Z(
        npu_inst_pe_1_6_6_N94) );
  MUX2_X1 npu_inst_pe_1_6_6_U156 ( .A(npu_inst_pe_1_6_6_n25), .B(
        npu_inst_pe_1_6_6_n24), .S(npu_inst_pe_1_6_6_n6), .Z(
        npu_inst_pe_1_6_6_n28) );
  MUX2_X1 npu_inst_pe_1_6_6_U155 ( .A(npu_inst_pe_1_6_6_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_6_6_int_q_reg_v_1__1_), .S(npu_inst_pe_1_6_6_n4), .Z(
        npu_inst_pe_1_6_6_n25) );
  MUX2_X1 npu_inst_pe_1_6_6_U154 ( .A(npu_inst_pe_1_6_6_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_6_6_int_q_reg_v_3__1_), .S(npu_inst_pe_1_6_6_n4), .Z(
        npu_inst_pe_1_6_6_n24) );
  MUX2_X1 npu_inst_pe_1_6_6_U153 ( .A(npu_inst_pe_1_6_6_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_6_6_int_q_reg_v_5__1_), .S(npu_inst_pe_1_6_6_n4), .Z(
        npu_inst_pe_1_6_6_n23) );
  MUX2_X1 npu_inst_pe_1_6_6_U152 ( .A(npu_inst_pe_1_6_6_n22), .B(
        npu_inst_pe_1_6_6_n19), .S(npu_inst_pe_1_6_6_n8), .Z(
        npu_inst_int_data_x_6__6__1_) );
  MUX2_X1 npu_inst_pe_1_6_6_U151 ( .A(npu_inst_pe_1_6_6_n21), .B(
        npu_inst_pe_1_6_6_n20), .S(npu_inst_pe_1_6_6_n6), .Z(
        npu_inst_pe_1_6_6_n22) );
  MUX2_X1 npu_inst_pe_1_6_6_U150 ( .A(npu_inst_pe_1_6_6_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_6_6_int_q_reg_h_1__1_), .S(npu_inst_pe_1_6_6_n4), .Z(
        npu_inst_pe_1_6_6_n21) );
  MUX2_X1 npu_inst_pe_1_6_6_U149 ( .A(npu_inst_pe_1_6_6_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_6_6_int_q_reg_h_3__1_), .S(npu_inst_pe_1_6_6_n4), .Z(
        npu_inst_pe_1_6_6_n20) );
  MUX2_X1 npu_inst_pe_1_6_6_U148 ( .A(npu_inst_pe_1_6_6_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_6_6_int_q_reg_h_5__1_), .S(npu_inst_pe_1_6_6_n4), .Z(
        npu_inst_pe_1_6_6_n19) );
  MUX2_X1 npu_inst_pe_1_6_6_U147 ( .A(npu_inst_pe_1_6_6_n18), .B(
        npu_inst_pe_1_6_6_n15), .S(npu_inst_pe_1_6_6_n8), .Z(
        npu_inst_int_data_x_6__6__0_) );
  MUX2_X1 npu_inst_pe_1_6_6_U146 ( .A(npu_inst_pe_1_6_6_n17), .B(
        npu_inst_pe_1_6_6_n16), .S(npu_inst_pe_1_6_6_n6), .Z(
        npu_inst_pe_1_6_6_n18) );
  MUX2_X1 npu_inst_pe_1_6_6_U145 ( .A(npu_inst_pe_1_6_6_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_6_6_int_q_reg_h_1__0_), .S(npu_inst_pe_1_6_6_n4), .Z(
        npu_inst_pe_1_6_6_n17) );
  MUX2_X1 npu_inst_pe_1_6_6_U144 ( .A(npu_inst_pe_1_6_6_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_6_6_int_q_reg_h_3__0_), .S(npu_inst_pe_1_6_6_n4), .Z(
        npu_inst_pe_1_6_6_n16) );
  MUX2_X1 npu_inst_pe_1_6_6_U143 ( .A(npu_inst_pe_1_6_6_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_6_6_int_q_reg_h_5__0_), .S(npu_inst_pe_1_6_6_n4), .Z(
        npu_inst_pe_1_6_6_n15) );
  XOR2_X1 npu_inst_pe_1_6_6_U142 ( .A(npu_inst_pe_1_6_6_int_data_0_), .B(
        npu_inst_pe_1_6_6_int_q_acc_0_), .Z(npu_inst_pe_1_6_6_N73) );
  AND2_X1 npu_inst_pe_1_6_6_U141 ( .A1(npu_inst_pe_1_6_6_int_q_acc_0_), .A2(
        npu_inst_pe_1_6_6_int_data_0_), .ZN(npu_inst_pe_1_6_6_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_6_6_U140 ( .A(npu_inst_pe_1_6_6_int_q_acc_0_), .B(
        npu_inst_pe_1_6_6_n13), .ZN(npu_inst_pe_1_6_6_N65) );
  OR2_X1 npu_inst_pe_1_6_6_U139 ( .A1(npu_inst_pe_1_6_6_n13), .A2(
        npu_inst_pe_1_6_6_int_q_acc_0_), .ZN(npu_inst_pe_1_6_6_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_6_6_U138 ( .A(npu_inst_pe_1_6_6_int_q_acc_2_), .B(
        npu_inst_pe_1_6_6_add_79_carry_2_), .Z(npu_inst_pe_1_6_6_N75) );
  AND2_X1 npu_inst_pe_1_6_6_U137 ( .A1(npu_inst_pe_1_6_6_add_79_carry_2_), 
        .A2(npu_inst_pe_1_6_6_int_q_acc_2_), .ZN(
        npu_inst_pe_1_6_6_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_6_6_U136 ( .A(npu_inst_pe_1_6_6_int_q_acc_3_), .B(
        npu_inst_pe_1_6_6_add_79_carry_3_), .Z(npu_inst_pe_1_6_6_N76) );
  AND2_X1 npu_inst_pe_1_6_6_U135 ( .A1(npu_inst_pe_1_6_6_add_79_carry_3_), 
        .A2(npu_inst_pe_1_6_6_int_q_acc_3_), .ZN(
        npu_inst_pe_1_6_6_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_6_6_U134 ( .A(npu_inst_pe_1_6_6_int_q_acc_4_), .B(
        npu_inst_pe_1_6_6_add_79_carry_4_), .Z(npu_inst_pe_1_6_6_N77) );
  AND2_X1 npu_inst_pe_1_6_6_U133 ( .A1(npu_inst_pe_1_6_6_add_79_carry_4_), 
        .A2(npu_inst_pe_1_6_6_int_q_acc_4_), .ZN(
        npu_inst_pe_1_6_6_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_6_6_U132 ( .A(npu_inst_pe_1_6_6_int_q_acc_5_), .B(
        npu_inst_pe_1_6_6_add_79_carry_5_), .Z(npu_inst_pe_1_6_6_N78) );
  AND2_X1 npu_inst_pe_1_6_6_U131 ( .A1(npu_inst_pe_1_6_6_add_79_carry_5_), 
        .A2(npu_inst_pe_1_6_6_int_q_acc_5_), .ZN(
        npu_inst_pe_1_6_6_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_6_6_U130 ( .A(npu_inst_pe_1_6_6_int_q_acc_6_), .B(
        npu_inst_pe_1_6_6_add_79_carry_6_), .Z(npu_inst_pe_1_6_6_N79) );
  AND2_X1 npu_inst_pe_1_6_6_U129 ( .A1(npu_inst_pe_1_6_6_add_79_carry_6_), 
        .A2(npu_inst_pe_1_6_6_int_q_acc_6_), .ZN(
        npu_inst_pe_1_6_6_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_6_6_U128 ( .A(npu_inst_pe_1_6_6_int_q_acc_7_), .B(
        npu_inst_pe_1_6_6_add_79_carry_7_), .Z(npu_inst_pe_1_6_6_N80) );
  XNOR2_X1 npu_inst_pe_1_6_6_U127 ( .A(npu_inst_pe_1_6_6_sub_77_carry_2_), .B(
        npu_inst_pe_1_6_6_int_q_acc_2_), .ZN(npu_inst_pe_1_6_6_N67) );
  OR2_X1 npu_inst_pe_1_6_6_U126 ( .A1(npu_inst_pe_1_6_6_int_q_acc_2_), .A2(
        npu_inst_pe_1_6_6_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_6_6_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_6_6_U125 ( .A(npu_inst_pe_1_6_6_sub_77_carry_3_), .B(
        npu_inst_pe_1_6_6_int_q_acc_3_), .ZN(npu_inst_pe_1_6_6_N68) );
  OR2_X1 npu_inst_pe_1_6_6_U124 ( .A1(npu_inst_pe_1_6_6_int_q_acc_3_), .A2(
        npu_inst_pe_1_6_6_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_6_6_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_6_6_U123 ( .A(npu_inst_pe_1_6_6_sub_77_carry_4_), .B(
        npu_inst_pe_1_6_6_int_q_acc_4_), .ZN(npu_inst_pe_1_6_6_N69) );
  OR2_X1 npu_inst_pe_1_6_6_U122 ( .A1(npu_inst_pe_1_6_6_int_q_acc_4_), .A2(
        npu_inst_pe_1_6_6_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_6_6_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_6_6_U121 ( .A(npu_inst_pe_1_6_6_sub_77_carry_5_), .B(
        npu_inst_pe_1_6_6_int_q_acc_5_), .ZN(npu_inst_pe_1_6_6_N70) );
  OR2_X1 npu_inst_pe_1_6_6_U120 ( .A1(npu_inst_pe_1_6_6_int_q_acc_5_), .A2(
        npu_inst_pe_1_6_6_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_6_6_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_6_6_U119 ( .A(npu_inst_pe_1_6_6_sub_77_carry_6_), .B(
        npu_inst_pe_1_6_6_int_q_acc_6_), .ZN(npu_inst_pe_1_6_6_N71) );
  OR2_X1 npu_inst_pe_1_6_6_U118 ( .A1(npu_inst_pe_1_6_6_int_q_acc_6_), .A2(
        npu_inst_pe_1_6_6_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_6_6_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_6_6_U117 ( .A(npu_inst_pe_1_6_6_int_q_acc_7_), .B(
        npu_inst_pe_1_6_6_sub_77_carry_7_), .ZN(npu_inst_pe_1_6_6_N72) );
  INV_X1 npu_inst_pe_1_6_6_U116 ( .A(npu_inst_n75), .ZN(npu_inst_pe_1_6_6_n7)
         );
  INV_X1 npu_inst_pe_1_6_6_U115 ( .A(npu_inst_pe_1_6_6_n7), .ZN(
        npu_inst_pe_1_6_6_n6) );
  INV_X1 npu_inst_pe_1_6_6_U114 ( .A(npu_inst_n53), .ZN(npu_inst_pe_1_6_6_n3)
         );
  AOI22_X1 npu_inst_pe_1_6_6_U113 ( .A1(npu_inst_int_data_y_7__6__0_), .A2(
        npu_inst_pe_1_6_6_n58), .B1(npu_inst_pe_1_6_6_n114), .B2(
        npu_inst_pe_1_6_6_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_6_6_n57) );
  INV_X1 npu_inst_pe_1_6_6_U112 ( .A(npu_inst_pe_1_6_6_n57), .ZN(
        npu_inst_pe_1_6_6_n108) );
  AOI22_X1 npu_inst_pe_1_6_6_U111 ( .A1(npu_inst_int_data_y_7__6__0_), .A2(
        npu_inst_pe_1_6_6_n54), .B1(npu_inst_pe_1_6_6_n115), .B2(
        npu_inst_pe_1_6_6_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_6_6_n53) );
  INV_X1 npu_inst_pe_1_6_6_U110 ( .A(npu_inst_pe_1_6_6_n53), .ZN(
        npu_inst_pe_1_6_6_n109) );
  AOI22_X1 npu_inst_pe_1_6_6_U107 ( .A1(npu_inst_int_data_y_7__6__0_), .A2(
        npu_inst_pe_1_6_6_n50), .B1(npu_inst_pe_1_6_6_n116), .B2(
        npu_inst_pe_1_6_6_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_6_6_n49) );
  INV_X1 npu_inst_pe_1_6_6_U106 ( .A(npu_inst_pe_1_6_6_n49), .ZN(
        npu_inst_pe_1_6_6_n110) );
  AOI22_X1 npu_inst_pe_1_6_6_U105 ( .A1(npu_inst_int_data_y_7__6__0_), .A2(
        npu_inst_pe_1_6_6_n46), .B1(npu_inst_pe_1_6_6_n117), .B2(
        npu_inst_pe_1_6_6_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_6_6_n45) );
  INV_X1 npu_inst_pe_1_6_6_U104 ( .A(npu_inst_pe_1_6_6_n45), .ZN(
        npu_inst_pe_1_6_6_n111) );
  AOI22_X1 npu_inst_pe_1_6_6_U103 ( .A1(npu_inst_int_data_y_7__6__0_), .A2(
        npu_inst_pe_1_6_6_n42), .B1(npu_inst_pe_1_6_6_n119), .B2(
        npu_inst_pe_1_6_6_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_6_6_n41) );
  INV_X1 npu_inst_pe_1_6_6_U102 ( .A(npu_inst_pe_1_6_6_n41), .ZN(
        npu_inst_pe_1_6_6_n112) );
  AOI22_X1 npu_inst_pe_1_6_6_U101 ( .A1(npu_inst_int_data_y_7__6__1_), .A2(
        npu_inst_pe_1_6_6_n58), .B1(npu_inst_pe_1_6_6_n114), .B2(
        npu_inst_pe_1_6_6_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_6_6_n59) );
  INV_X1 npu_inst_pe_1_6_6_U100 ( .A(npu_inst_pe_1_6_6_n59), .ZN(
        npu_inst_pe_1_6_6_n102) );
  AOI22_X1 npu_inst_pe_1_6_6_U99 ( .A1(npu_inst_int_data_y_7__6__1_), .A2(
        npu_inst_pe_1_6_6_n54), .B1(npu_inst_pe_1_6_6_n115), .B2(
        npu_inst_pe_1_6_6_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_6_6_n55) );
  INV_X1 npu_inst_pe_1_6_6_U98 ( .A(npu_inst_pe_1_6_6_n55), .ZN(
        npu_inst_pe_1_6_6_n103) );
  AOI22_X1 npu_inst_pe_1_6_6_U97 ( .A1(npu_inst_int_data_y_7__6__1_), .A2(
        npu_inst_pe_1_6_6_n50), .B1(npu_inst_pe_1_6_6_n116), .B2(
        npu_inst_pe_1_6_6_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_6_6_n51) );
  INV_X1 npu_inst_pe_1_6_6_U96 ( .A(npu_inst_pe_1_6_6_n51), .ZN(
        npu_inst_pe_1_6_6_n104) );
  AOI22_X1 npu_inst_pe_1_6_6_U95 ( .A1(npu_inst_int_data_y_7__6__1_), .A2(
        npu_inst_pe_1_6_6_n46), .B1(npu_inst_pe_1_6_6_n117), .B2(
        npu_inst_pe_1_6_6_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_6_6_n47) );
  INV_X1 npu_inst_pe_1_6_6_U94 ( .A(npu_inst_pe_1_6_6_n47), .ZN(
        npu_inst_pe_1_6_6_n105) );
  AOI22_X1 npu_inst_pe_1_6_6_U93 ( .A1(npu_inst_int_data_y_7__6__1_), .A2(
        npu_inst_pe_1_6_6_n42), .B1(npu_inst_pe_1_6_6_n119), .B2(
        npu_inst_pe_1_6_6_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_6_6_n43) );
  INV_X1 npu_inst_pe_1_6_6_U92 ( .A(npu_inst_pe_1_6_6_n43), .ZN(
        npu_inst_pe_1_6_6_n106) );
  AOI22_X1 npu_inst_pe_1_6_6_U91 ( .A1(npu_inst_pe_1_6_6_n38), .A2(
        npu_inst_int_data_y_7__6__1_), .B1(npu_inst_pe_1_6_6_n118), .B2(
        npu_inst_pe_1_6_6_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_6_6_n39) );
  INV_X1 npu_inst_pe_1_6_6_U90 ( .A(npu_inst_pe_1_6_6_n39), .ZN(
        npu_inst_pe_1_6_6_n107) );
  AOI22_X1 npu_inst_pe_1_6_6_U89 ( .A1(npu_inst_pe_1_6_6_n38), .A2(
        npu_inst_int_data_y_7__6__0_), .B1(npu_inst_pe_1_6_6_n118), .B2(
        npu_inst_pe_1_6_6_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_6_6_n37) );
  INV_X1 npu_inst_pe_1_6_6_U88 ( .A(npu_inst_pe_1_6_6_n37), .ZN(
        npu_inst_pe_1_6_6_n113) );
  NAND2_X1 npu_inst_pe_1_6_6_U87 ( .A1(npu_inst_pe_1_6_6_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_6_6_n60), .ZN(npu_inst_pe_1_6_6_n74) );
  OAI21_X1 npu_inst_pe_1_6_6_U86 ( .B1(npu_inst_pe_1_6_6_n63), .B2(
        npu_inst_pe_1_6_6_n60), .A(npu_inst_pe_1_6_6_n74), .ZN(
        npu_inst_pe_1_6_6_n97) );
  NAND2_X1 npu_inst_pe_1_6_6_U85 ( .A1(npu_inst_pe_1_6_6_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_6_6_n60), .ZN(npu_inst_pe_1_6_6_n73) );
  OAI21_X1 npu_inst_pe_1_6_6_U84 ( .B1(npu_inst_pe_1_6_6_n61), .B2(
        npu_inst_pe_1_6_6_n60), .A(npu_inst_pe_1_6_6_n73), .ZN(
        npu_inst_pe_1_6_6_n96) );
  NAND2_X1 npu_inst_pe_1_6_6_U83 ( .A1(npu_inst_pe_1_6_6_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_6_6_n56), .ZN(npu_inst_pe_1_6_6_n72) );
  OAI21_X1 npu_inst_pe_1_6_6_U82 ( .B1(npu_inst_pe_1_6_6_n63), .B2(
        npu_inst_pe_1_6_6_n56), .A(npu_inst_pe_1_6_6_n72), .ZN(
        npu_inst_pe_1_6_6_n95) );
  NAND2_X1 npu_inst_pe_1_6_6_U81 ( .A1(npu_inst_pe_1_6_6_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_6_6_n56), .ZN(npu_inst_pe_1_6_6_n71) );
  OAI21_X1 npu_inst_pe_1_6_6_U80 ( .B1(npu_inst_pe_1_6_6_n61), .B2(
        npu_inst_pe_1_6_6_n56), .A(npu_inst_pe_1_6_6_n71), .ZN(
        npu_inst_pe_1_6_6_n94) );
  NAND2_X1 npu_inst_pe_1_6_6_U79 ( .A1(npu_inst_pe_1_6_6_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_6_6_n52), .ZN(npu_inst_pe_1_6_6_n70) );
  OAI21_X1 npu_inst_pe_1_6_6_U78 ( .B1(npu_inst_pe_1_6_6_n63), .B2(
        npu_inst_pe_1_6_6_n52), .A(npu_inst_pe_1_6_6_n70), .ZN(
        npu_inst_pe_1_6_6_n93) );
  NAND2_X1 npu_inst_pe_1_6_6_U77 ( .A1(npu_inst_pe_1_6_6_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_6_6_n52), .ZN(npu_inst_pe_1_6_6_n69) );
  OAI21_X1 npu_inst_pe_1_6_6_U76 ( .B1(npu_inst_pe_1_6_6_n61), .B2(
        npu_inst_pe_1_6_6_n52), .A(npu_inst_pe_1_6_6_n69), .ZN(
        npu_inst_pe_1_6_6_n92) );
  NAND2_X1 npu_inst_pe_1_6_6_U75 ( .A1(npu_inst_pe_1_6_6_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_6_6_n48), .ZN(npu_inst_pe_1_6_6_n68) );
  OAI21_X1 npu_inst_pe_1_6_6_U74 ( .B1(npu_inst_pe_1_6_6_n63), .B2(
        npu_inst_pe_1_6_6_n48), .A(npu_inst_pe_1_6_6_n68), .ZN(
        npu_inst_pe_1_6_6_n91) );
  NAND2_X1 npu_inst_pe_1_6_6_U73 ( .A1(npu_inst_pe_1_6_6_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_6_6_n48), .ZN(npu_inst_pe_1_6_6_n67) );
  OAI21_X1 npu_inst_pe_1_6_6_U72 ( .B1(npu_inst_pe_1_6_6_n61), .B2(
        npu_inst_pe_1_6_6_n48), .A(npu_inst_pe_1_6_6_n67), .ZN(
        npu_inst_pe_1_6_6_n90) );
  NAND2_X1 npu_inst_pe_1_6_6_U71 ( .A1(npu_inst_pe_1_6_6_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_6_6_n44), .ZN(npu_inst_pe_1_6_6_n66) );
  OAI21_X1 npu_inst_pe_1_6_6_U70 ( .B1(npu_inst_pe_1_6_6_n63), .B2(
        npu_inst_pe_1_6_6_n44), .A(npu_inst_pe_1_6_6_n66), .ZN(
        npu_inst_pe_1_6_6_n89) );
  NAND2_X1 npu_inst_pe_1_6_6_U69 ( .A1(npu_inst_pe_1_6_6_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_6_6_n44), .ZN(npu_inst_pe_1_6_6_n65) );
  OAI21_X1 npu_inst_pe_1_6_6_U68 ( .B1(npu_inst_pe_1_6_6_n61), .B2(
        npu_inst_pe_1_6_6_n44), .A(npu_inst_pe_1_6_6_n65), .ZN(
        npu_inst_pe_1_6_6_n88) );
  NAND2_X1 npu_inst_pe_1_6_6_U67 ( .A1(npu_inst_pe_1_6_6_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_6_6_n40), .ZN(npu_inst_pe_1_6_6_n64) );
  OAI21_X1 npu_inst_pe_1_6_6_U66 ( .B1(npu_inst_pe_1_6_6_n63), .B2(
        npu_inst_pe_1_6_6_n40), .A(npu_inst_pe_1_6_6_n64), .ZN(
        npu_inst_pe_1_6_6_n87) );
  NAND2_X1 npu_inst_pe_1_6_6_U65 ( .A1(npu_inst_pe_1_6_6_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_6_6_n40), .ZN(npu_inst_pe_1_6_6_n62) );
  OAI21_X1 npu_inst_pe_1_6_6_U64 ( .B1(npu_inst_pe_1_6_6_n61), .B2(
        npu_inst_pe_1_6_6_n40), .A(npu_inst_pe_1_6_6_n62), .ZN(
        npu_inst_pe_1_6_6_n86) );
  AND2_X1 npu_inst_pe_1_6_6_U63 ( .A1(npu_inst_pe_1_6_6_N93), .A2(npu_inst_n53), .ZN(npu_inst_int_data_y_6__6__0_) );
  AND2_X1 npu_inst_pe_1_6_6_U62 ( .A1(npu_inst_n53), .A2(npu_inst_pe_1_6_6_N94), .ZN(npu_inst_int_data_y_6__6__1_) );
  NOR3_X1 npu_inst_pe_1_6_6_U61 ( .A1(npu_inst_pe_1_6_6_n26), .A2(npu_inst_n53), .A3(npu_inst_int_ckg[9]), .ZN(npu_inst_pe_1_6_6_n85) );
  OR2_X1 npu_inst_pe_1_6_6_U60 ( .A1(npu_inst_pe_1_6_6_n85), .A2(
        npu_inst_pe_1_6_6_n2), .ZN(npu_inst_pe_1_6_6_N84) );
  AND2_X1 npu_inst_pe_1_6_6_U59 ( .A1(npu_inst_pe_1_6_6_int_q_acc_0_), .A2(
        npu_inst_pe_1_6_6_n1), .ZN(npu_inst_int_data_res_6__6__0_) );
  AND2_X1 npu_inst_pe_1_6_6_U58 ( .A1(npu_inst_pe_1_6_6_n2), .A2(
        npu_inst_pe_1_6_6_int_q_acc_7_), .ZN(npu_inst_int_data_res_6__6__7_)
         );
  AND2_X1 npu_inst_pe_1_6_6_U57 ( .A1(npu_inst_pe_1_6_6_int_q_acc_1_), .A2(
        npu_inst_pe_1_6_6_n1), .ZN(npu_inst_int_data_res_6__6__1_) );
  AND2_X1 npu_inst_pe_1_6_6_U56 ( .A1(npu_inst_pe_1_6_6_int_q_acc_2_), .A2(
        npu_inst_pe_1_6_6_n1), .ZN(npu_inst_int_data_res_6__6__2_) );
  AND2_X1 npu_inst_pe_1_6_6_U55 ( .A1(npu_inst_pe_1_6_6_int_q_acc_3_), .A2(
        npu_inst_pe_1_6_6_n2), .ZN(npu_inst_int_data_res_6__6__3_) );
  AND2_X1 npu_inst_pe_1_6_6_U54 ( .A1(npu_inst_pe_1_6_6_int_q_acc_4_), .A2(
        npu_inst_pe_1_6_6_n2), .ZN(npu_inst_int_data_res_6__6__4_) );
  AND2_X1 npu_inst_pe_1_6_6_U53 ( .A1(npu_inst_pe_1_6_6_int_q_acc_5_), .A2(
        npu_inst_pe_1_6_6_n2), .ZN(npu_inst_int_data_res_6__6__5_) );
  AND2_X1 npu_inst_pe_1_6_6_U52 ( .A1(npu_inst_pe_1_6_6_int_q_acc_6_), .A2(
        npu_inst_pe_1_6_6_n2), .ZN(npu_inst_int_data_res_6__6__6_) );
  AOI222_X1 npu_inst_pe_1_6_6_U51 ( .A1(npu_inst_int_data_res_7__6__0_), .A2(
        npu_inst_pe_1_6_6_n1), .B1(npu_inst_pe_1_6_6_N73), .B2(
        npu_inst_pe_1_6_6_n76), .C1(npu_inst_pe_1_6_6_N65), .C2(
        npu_inst_pe_1_6_6_n77), .ZN(npu_inst_pe_1_6_6_n84) );
  INV_X1 npu_inst_pe_1_6_6_U50 ( .A(npu_inst_pe_1_6_6_n84), .ZN(
        npu_inst_pe_1_6_6_n101) );
  AOI222_X1 npu_inst_pe_1_6_6_U49 ( .A1(npu_inst_int_data_res_7__6__7_), .A2(
        npu_inst_pe_1_6_6_n1), .B1(npu_inst_pe_1_6_6_N80), .B2(
        npu_inst_pe_1_6_6_n76), .C1(npu_inst_pe_1_6_6_N72), .C2(
        npu_inst_pe_1_6_6_n77), .ZN(npu_inst_pe_1_6_6_n75) );
  INV_X1 npu_inst_pe_1_6_6_U48 ( .A(npu_inst_pe_1_6_6_n75), .ZN(
        npu_inst_pe_1_6_6_n33) );
  AOI222_X1 npu_inst_pe_1_6_6_U47 ( .A1(npu_inst_int_data_res_7__6__1_), .A2(
        npu_inst_pe_1_6_6_n1), .B1(npu_inst_pe_1_6_6_N74), .B2(
        npu_inst_pe_1_6_6_n76), .C1(npu_inst_pe_1_6_6_N66), .C2(
        npu_inst_pe_1_6_6_n77), .ZN(npu_inst_pe_1_6_6_n83) );
  INV_X1 npu_inst_pe_1_6_6_U46 ( .A(npu_inst_pe_1_6_6_n83), .ZN(
        npu_inst_pe_1_6_6_n100) );
  AOI222_X1 npu_inst_pe_1_6_6_U45 ( .A1(npu_inst_int_data_res_7__6__2_), .A2(
        npu_inst_pe_1_6_6_n1), .B1(npu_inst_pe_1_6_6_N75), .B2(
        npu_inst_pe_1_6_6_n76), .C1(npu_inst_pe_1_6_6_N67), .C2(
        npu_inst_pe_1_6_6_n77), .ZN(npu_inst_pe_1_6_6_n82) );
  INV_X1 npu_inst_pe_1_6_6_U44 ( .A(npu_inst_pe_1_6_6_n82), .ZN(
        npu_inst_pe_1_6_6_n99) );
  AOI222_X1 npu_inst_pe_1_6_6_U43 ( .A1(npu_inst_int_data_res_7__6__3_), .A2(
        npu_inst_pe_1_6_6_n1), .B1(npu_inst_pe_1_6_6_N76), .B2(
        npu_inst_pe_1_6_6_n76), .C1(npu_inst_pe_1_6_6_N68), .C2(
        npu_inst_pe_1_6_6_n77), .ZN(npu_inst_pe_1_6_6_n81) );
  INV_X1 npu_inst_pe_1_6_6_U42 ( .A(npu_inst_pe_1_6_6_n81), .ZN(
        npu_inst_pe_1_6_6_n98) );
  AOI222_X1 npu_inst_pe_1_6_6_U41 ( .A1(npu_inst_int_data_res_7__6__4_), .A2(
        npu_inst_pe_1_6_6_n1), .B1(npu_inst_pe_1_6_6_N77), .B2(
        npu_inst_pe_1_6_6_n76), .C1(npu_inst_pe_1_6_6_N69), .C2(
        npu_inst_pe_1_6_6_n77), .ZN(npu_inst_pe_1_6_6_n80) );
  INV_X1 npu_inst_pe_1_6_6_U40 ( .A(npu_inst_pe_1_6_6_n80), .ZN(
        npu_inst_pe_1_6_6_n36) );
  AOI222_X1 npu_inst_pe_1_6_6_U39 ( .A1(npu_inst_int_data_res_7__6__5_), .A2(
        npu_inst_pe_1_6_6_n1), .B1(npu_inst_pe_1_6_6_N78), .B2(
        npu_inst_pe_1_6_6_n76), .C1(npu_inst_pe_1_6_6_N70), .C2(
        npu_inst_pe_1_6_6_n77), .ZN(npu_inst_pe_1_6_6_n79) );
  INV_X1 npu_inst_pe_1_6_6_U38 ( .A(npu_inst_pe_1_6_6_n79), .ZN(
        npu_inst_pe_1_6_6_n35) );
  AOI222_X1 npu_inst_pe_1_6_6_U37 ( .A1(npu_inst_int_data_res_7__6__6_), .A2(
        npu_inst_pe_1_6_6_n1), .B1(npu_inst_pe_1_6_6_N79), .B2(
        npu_inst_pe_1_6_6_n76), .C1(npu_inst_pe_1_6_6_N71), .C2(
        npu_inst_pe_1_6_6_n77), .ZN(npu_inst_pe_1_6_6_n78) );
  INV_X1 npu_inst_pe_1_6_6_U36 ( .A(npu_inst_pe_1_6_6_n78), .ZN(
        npu_inst_pe_1_6_6_n34) );
  INV_X1 npu_inst_pe_1_6_6_U35 ( .A(npu_inst_pe_1_6_6_int_data_1_), .ZN(
        npu_inst_pe_1_6_6_n14) );
  AND2_X1 npu_inst_pe_1_6_6_U34 ( .A1(npu_inst_int_data_x_6__6__1_), .A2(
        npu_inst_pe_1_6_6_int_q_weight_1_), .ZN(npu_inst_pe_1_6_6_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_6_6_U33 ( .A1(npu_inst_int_data_x_6__6__0_), .A2(
        npu_inst_pe_1_6_6_int_q_weight_1_), .ZN(npu_inst_pe_1_6_6_int_data_0_)
         );
  AOI22_X1 npu_inst_pe_1_6_6_U32 ( .A1(npu_inst_n53), .A2(
        npu_inst_int_data_y_7__6__1_), .B1(npu_inst_pe_1_6_6_n3), .B2(
        npu_inst_int_data_x_6__7__1_), .ZN(npu_inst_pe_1_6_6_n63) );
  AOI22_X1 npu_inst_pe_1_6_6_U31 ( .A1(npu_inst_n53), .A2(
        npu_inst_int_data_y_7__6__0_), .B1(npu_inst_pe_1_6_6_n3), .B2(
        npu_inst_int_data_x_6__7__0_), .ZN(npu_inst_pe_1_6_6_n61) );
  INV_X1 npu_inst_pe_1_6_6_U30 ( .A(npu_inst_pe_1_6_6_int_data_0_), .ZN(
        npu_inst_pe_1_6_6_n13) );
  INV_X1 npu_inst_pe_1_6_6_U29 ( .A(npu_inst_n67), .ZN(npu_inst_pe_1_6_6_n5)
         );
  OR3_X1 npu_inst_pe_1_6_6_U28 ( .A1(npu_inst_pe_1_6_6_n6), .A2(
        npu_inst_pe_1_6_6_n8), .A3(npu_inst_pe_1_6_6_n5), .ZN(
        npu_inst_pe_1_6_6_n56) );
  OR3_X1 npu_inst_pe_1_6_6_U27 ( .A1(npu_inst_pe_1_6_6_n5), .A2(
        npu_inst_pe_1_6_6_n8), .A3(npu_inst_pe_1_6_6_n7), .ZN(
        npu_inst_pe_1_6_6_n48) );
  INV_X1 npu_inst_pe_1_6_6_U26 ( .A(npu_inst_pe_1_6_6_n5), .ZN(
        npu_inst_pe_1_6_6_n4) );
  INV_X1 npu_inst_pe_1_6_6_U25 ( .A(npu_inst_n122), .ZN(npu_inst_pe_1_6_6_n12)
         );
  OR3_X1 npu_inst_pe_1_6_6_U24 ( .A1(npu_inst_pe_1_6_6_n4), .A2(
        npu_inst_pe_1_6_6_n8), .A3(npu_inst_pe_1_6_6_n7), .ZN(
        npu_inst_pe_1_6_6_n52) );
  OR3_X1 npu_inst_pe_1_6_6_U23 ( .A1(npu_inst_pe_1_6_6_n6), .A2(
        npu_inst_pe_1_6_6_n8), .A3(npu_inst_pe_1_6_6_n4), .ZN(
        npu_inst_pe_1_6_6_n60) );
  NOR2_X1 npu_inst_pe_1_6_6_U22 ( .A1(npu_inst_pe_1_6_6_n60), .A2(
        npu_inst_pe_1_6_6_n3), .ZN(npu_inst_pe_1_6_6_n58) );
  NOR2_X1 npu_inst_pe_1_6_6_U21 ( .A1(npu_inst_pe_1_6_6_n56), .A2(
        npu_inst_pe_1_6_6_n3), .ZN(npu_inst_pe_1_6_6_n54) );
  NOR2_X1 npu_inst_pe_1_6_6_U20 ( .A1(npu_inst_pe_1_6_6_n52), .A2(
        npu_inst_pe_1_6_6_n3), .ZN(npu_inst_pe_1_6_6_n50) );
  NOR2_X1 npu_inst_pe_1_6_6_U19 ( .A1(npu_inst_pe_1_6_6_n48), .A2(
        npu_inst_pe_1_6_6_n3), .ZN(npu_inst_pe_1_6_6_n46) );
  NOR2_X1 npu_inst_pe_1_6_6_U18 ( .A1(npu_inst_pe_1_6_6_n40), .A2(
        npu_inst_pe_1_6_6_n3), .ZN(npu_inst_pe_1_6_6_n38) );
  NOR2_X1 npu_inst_pe_1_6_6_U17 ( .A1(npu_inst_pe_1_6_6_n44), .A2(
        npu_inst_pe_1_6_6_n3), .ZN(npu_inst_pe_1_6_6_n42) );
  BUF_X1 npu_inst_pe_1_6_6_U16 ( .A(npu_inst_n94), .Z(npu_inst_pe_1_6_6_n8) );
  BUF_X1 npu_inst_pe_1_6_6_U15 ( .A(npu_inst_pe_1_6_6_n12), .Z(
        npu_inst_pe_1_6_6_n11) );
  BUF_X1 npu_inst_pe_1_6_6_U14 ( .A(npu_inst_pe_1_6_6_n12), .Z(
        npu_inst_pe_1_6_6_n10) );
  BUF_X1 npu_inst_pe_1_6_6_U13 ( .A(npu_inst_pe_1_6_6_n12), .Z(
        npu_inst_pe_1_6_6_n9) );
  INV_X1 npu_inst_pe_1_6_6_U12 ( .A(npu_inst_pe_1_6_6_n38), .ZN(
        npu_inst_pe_1_6_6_n118) );
  INV_X1 npu_inst_pe_1_6_6_U11 ( .A(npu_inst_pe_1_6_6_n58), .ZN(
        npu_inst_pe_1_6_6_n114) );
  INV_X1 npu_inst_pe_1_6_6_U10 ( .A(npu_inst_pe_1_6_6_n54), .ZN(
        npu_inst_pe_1_6_6_n115) );
  INV_X1 npu_inst_pe_1_6_6_U9 ( .A(npu_inst_pe_1_6_6_n50), .ZN(
        npu_inst_pe_1_6_6_n116) );
  INV_X1 npu_inst_pe_1_6_6_U8 ( .A(npu_inst_pe_1_6_6_n46), .ZN(
        npu_inst_pe_1_6_6_n117) );
  INV_X1 npu_inst_pe_1_6_6_U7 ( .A(npu_inst_pe_1_6_6_n42), .ZN(
        npu_inst_pe_1_6_6_n119) );
  BUF_X1 npu_inst_pe_1_6_6_U6 ( .A(npu_inst_n11), .Z(npu_inst_pe_1_6_6_n2) );
  BUF_X1 npu_inst_pe_1_6_6_U5 ( .A(npu_inst_n11), .Z(npu_inst_pe_1_6_6_n1) );
  NOR2_X1 npu_inst_pe_1_6_6_U4 ( .A1(npu_inst_pe_1_6_6_int_q_weight_0_), .A2(
        npu_inst_pe_1_6_6_n1), .ZN(npu_inst_pe_1_6_6_n76) );
  NOR2_X1 npu_inst_pe_1_6_6_U3 ( .A1(npu_inst_pe_1_6_6_n27), .A2(
        npu_inst_pe_1_6_6_n1), .ZN(npu_inst_pe_1_6_6_n77) );
  FA_X1 npu_inst_pe_1_6_6_sub_77_U2_1 ( .A(npu_inst_pe_1_6_6_int_q_acc_1_), 
        .B(npu_inst_pe_1_6_6_n14), .CI(npu_inst_pe_1_6_6_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_6_6_sub_77_carry_2_), .S(npu_inst_pe_1_6_6_N66) );
  FA_X1 npu_inst_pe_1_6_6_add_79_U1_1 ( .A(npu_inst_pe_1_6_6_int_q_acc_1_), 
        .B(npu_inst_pe_1_6_6_int_data_1_), .CI(
        npu_inst_pe_1_6_6_add_79_carry_1_), .CO(
        npu_inst_pe_1_6_6_add_79_carry_2_), .S(npu_inst_pe_1_6_6_N74) );
  NAND3_X1 npu_inst_pe_1_6_6_U109 ( .A1(npu_inst_pe_1_6_6_n5), .A2(
        npu_inst_pe_1_6_6_n7), .A3(npu_inst_pe_1_6_6_n8), .ZN(
        npu_inst_pe_1_6_6_n44) );
  NAND3_X1 npu_inst_pe_1_6_6_U108 ( .A1(npu_inst_pe_1_6_6_n4), .A2(
        npu_inst_pe_1_6_6_n7), .A3(npu_inst_pe_1_6_6_n8), .ZN(
        npu_inst_pe_1_6_6_n40) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_6_6_n34), .CK(
        npu_inst_pe_1_6_6_net3051), .RN(npu_inst_pe_1_6_6_n9), .Q(
        npu_inst_pe_1_6_6_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_6_6_n35), .CK(
        npu_inst_pe_1_6_6_net3051), .RN(npu_inst_pe_1_6_6_n9), .Q(
        npu_inst_pe_1_6_6_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_6_6_n36), .CK(
        npu_inst_pe_1_6_6_net3051), .RN(npu_inst_pe_1_6_6_n9), .Q(
        npu_inst_pe_1_6_6_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_6_6_n98), .CK(
        npu_inst_pe_1_6_6_net3051), .RN(npu_inst_pe_1_6_6_n9), .Q(
        npu_inst_pe_1_6_6_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_6_6_n99), .CK(
        npu_inst_pe_1_6_6_net3051), .RN(npu_inst_pe_1_6_6_n9), .Q(
        npu_inst_pe_1_6_6_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_6_6_n100), 
        .CK(npu_inst_pe_1_6_6_net3051), .RN(npu_inst_pe_1_6_6_n9), .Q(
        npu_inst_pe_1_6_6_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_6_6_n33), .CK(
        npu_inst_pe_1_6_6_net3051), .RN(npu_inst_pe_1_6_6_n9), .Q(
        npu_inst_pe_1_6_6_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_6_6_n101), 
        .CK(npu_inst_pe_1_6_6_net3051), .RN(npu_inst_pe_1_6_6_n9), .Q(
        npu_inst_pe_1_6_6_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_weight_reg_0_ ( .D(npu_inst_n108), .CK(
        npu_inst_pe_1_6_6_net3057), .RN(npu_inst_pe_1_6_6_n9), .Q(
        npu_inst_pe_1_6_6_int_q_weight_0_), .QN(npu_inst_pe_1_6_6_n27) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_weight_reg_1_ ( .D(npu_inst_n114), .CK(
        npu_inst_pe_1_6_6_net3057), .RN(npu_inst_pe_1_6_6_n9), .Q(
        npu_inst_pe_1_6_6_int_q_weight_1_), .QN(npu_inst_pe_1_6_6_n26) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_6_6_n113), 
        .CK(npu_inst_pe_1_6_6_net3057), .RN(npu_inst_pe_1_6_6_n9), .Q(
        npu_inst_pe_1_6_6_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_6_6_n107), 
        .CK(npu_inst_pe_1_6_6_net3057), .RN(npu_inst_pe_1_6_6_n9), .Q(
        npu_inst_pe_1_6_6_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_6_6_n112), 
        .CK(npu_inst_pe_1_6_6_net3057), .RN(npu_inst_pe_1_6_6_n10), .Q(
        npu_inst_pe_1_6_6_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_6_6_n106), 
        .CK(npu_inst_pe_1_6_6_net3057), .RN(npu_inst_pe_1_6_6_n10), .Q(
        npu_inst_pe_1_6_6_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_6_6_n111), 
        .CK(npu_inst_pe_1_6_6_net3057), .RN(npu_inst_pe_1_6_6_n10), .Q(
        npu_inst_pe_1_6_6_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_6_6_n105), 
        .CK(npu_inst_pe_1_6_6_net3057), .RN(npu_inst_pe_1_6_6_n10), .Q(
        npu_inst_pe_1_6_6_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_6_6_n110), 
        .CK(npu_inst_pe_1_6_6_net3057), .RN(npu_inst_pe_1_6_6_n10), .Q(
        npu_inst_pe_1_6_6_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_6_6_n104), 
        .CK(npu_inst_pe_1_6_6_net3057), .RN(npu_inst_pe_1_6_6_n10), .Q(
        npu_inst_pe_1_6_6_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_6_6_n109), 
        .CK(npu_inst_pe_1_6_6_net3057), .RN(npu_inst_pe_1_6_6_n10), .Q(
        npu_inst_pe_1_6_6_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_6_6_n103), 
        .CK(npu_inst_pe_1_6_6_net3057), .RN(npu_inst_pe_1_6_6_n10), .Q(
        npu_inst_pe_1_6_6_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_6_6_n108), 
        .CK(npu_inst_pe_1_6_6_net3057), .RN(npu_inst_pe_1_6_6_n10), .Q(
        npu_inst_pe_1_6_6_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_6_6_n102), 
        .CK(npu_inst_pe_1_6_6_net3057), .RN(npu_inst_pe_1_6_6_n10), .Q(
        npu_inst_pe_1_6_6_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_6_6_n86), 
        .CK(npu_inst_pe_1_6_6_net3057), .RN(npu_inst_pe_1_6_6_n10), .Q(
        npu_inst_pe_1_6_6_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_6_6_n87), 
        .CK(npu_inst_pe_1_6_6_net3057), .RN(npu_inst_pe_1_6_6_n10), .Q(
        npu_inst_pe_1_6_6_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_6_6_n88), 
        .CK(npu_inst_pe_1_6_6_net3057), .RN(npu_inst_pe_1_6_6_n11), .Q(
        npu_inst_pe_1_6_6_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_6_6_n89), 
        .CK(npu_inst_pe_1_6_6_net3057), .RN(npu_inst_pe_1_6_6_n11), .Q(
        npu_inst_pe_1_6_6_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_6_6_n90), 
        .CK(npu_inst_pe_1_6_6_net3057), .RN(npu_inst_pe_1_6_6_n11), .Q(
        npu_inst_pe_1_6_6_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_6_6_n91), 
        .CK(npu_inst_pe_1_6_6_net3057), .RN(npu_inst_pe_1_6_6_n11), .Q(
        npu_inst_pe_1_6_6_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_6_6_n92), 
        .CK(npu_inst_pe_1_6_6_net3057), .RN(npu_inst_pe_1_6_6_n11), .Q(
        npu_inst_pe_1_6_6_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_6_6_n93), 
        .CK(npu_inst_pe_1_6_6_net3057), .RN(npu_inst_pe_1_6_6_n11), .Q(
        npu_inst_pe_1_6_6_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_6_6_n94), 
        .CK(npu_inst_pe_1_6_6_net3057), .RN(npu_inst_pe_1_6_6_n11), .Q(
        npu_inst_pe_1_6_6_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_6_6_n95), 
        .CK(npu_inst_pe_1_6_6_net3057), .RN(npu_inst_pe_1_6_6_n11), .Q(
        npu_inst_pe_1_6_6_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_6_6_n96), 
        .CK(npu_inst_pe_1_6_6_net3057), .RN(npu_inst_pe_1_6_6_n11), .Q(
        npu_inst_pe_1_6_6_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_6_6_n97), 
        .CK(npu_inst_pe_1_6_6_net3057), .RN(npu_inst_pe_1_6_6_n11), .Q(
        npu_inst_pe_1_6_6_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_6_6_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_6_6_N84), .SE(1'b0), .GCK(npu_inst_pe_1_6_6_net3051) );
  CLKGATETST_X1 npu_inst_pe_1_6_6_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n61), .SE(1'b0), .GCK(npu_inst_pe_1_6_6_net3057) );
  MUX2_X1 npu_inst_pe_1_6_7_U162 ( .A(npu_inst_pe_1_6_7_n32), .B(
        npu_inst_pe_1_6_7_n29), .S(npu_inst_pe_1_6_7_n8), .Z(
        npu_inst_pe_1_6_7_N93) );
  MUX2_X1 npu_inst_pe_1_6_7_U161 ( .A(npu_inst_pe_1_6_7_n31), .B(
        npu_inst_pe_1_6_7_n30), .S(npu_inst_pe_1_6_7_n6), .Z(
        npu_inst_pe_1_6_7_n32) );
  MUX2_X1 npu_inst_pe_1_6_7_U160 ( .A(npu_inst_pe_1_6_7_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_6_7_int_q_reg_v_1__0_), .S(npu_inst_pe_1_6_7_n4), .Z(
        npu_inst_pe_1_6_7_n31) );
  MUX2_X1 npu_inst_pe_1_6_7_U159 ( .A(npu_inst_pe_1_6_7_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_6_7_int_q_reg_v_3__0_), .S(npu_inst_pe_1_6_7_n4), .Z(
        npu_inst_pe_1_6_7_n30) );
  MUX2_X1 npu_inst_pe_1_6_7_U158 ( .A(npu_inst_pe_1_6_7_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_6_7_int_q_reg_v_5__0_), .S(npu_inst_pe_1_6_7_n4), .Z(
        npu_inst_pe_1_6_7_n29) );
  MUX2_X1 npu_inst_pe_1_6_7_U157 ( .A(npu_inst_pe_1_6_7_n28), .B(
        npu_inst_pe_1_6_7_n23), .S(npu_inst_pe_1_6_7_n8), .Z(
        npu_inst_pe_1_6_7_N94) );
  MUX2_X1 npu_inst_pe_1_6_7_U156 ( .A(npu_inst_pe_1_6_7_n25), .B(
        npu_inst_pe_1_6_7_n24), .S(npu_inst_pe_1_6_7_n6), .Z(
        npu_inst_pe_1_6_7_n28) );
  MUX2_X1 npu_inst_pe_1_6_7_U155 ( .A(npu_inst_pe_1_6_7_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_6_7_int_q_reg_v_1__1_), .S(npu_inst_pe_1_6_7_n4), .Z(
        npu_inst_pe_1_6_7_n25) );
  MUX2_X1 npu_inst_pe_1_6_7_U154 ( .A(npu_inst_pe_1_6_7_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_6_7_int_q_reg_v_3__1_), .S(npu_inst_pe_1_6_7_n4), .Z(
        npu_inst_pe_1_6_7_n24) );
  MUX2_X1 npu_inst_pe_1_6_7_U153 ( .A(npu_inst_pe_1_6_7_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_6_7_int_q_reg_v_5__1_), .S(npu_inst_pe_1_6_7_n4), .Z(
        npu_inst_pe_1_6_7_n23) );
  MUX2_X1 npu_inst_pe_1_6_7_U152 ( .A(npu_inst_pe_1_6_7_n22), .B(
        npu_inst_pe_1_6_7_n19), .S(npu_inst_pe_1_6_7_n8), .Z(
        npu_inst_int_data_x_6__7__1_) );
  MUX2_X1 npu_inst_pe_1_6_7_U151 ( .A(npu_inst_pe_1_6_7_n21), .B(
        npu_inst_pe_1_6_7_n20), .S(npu_inst_pe_1_6_7_n6), .Z(
        npu_inst_pe_1_6_7_n22) );
  MUX2_X1 npu_inst_pe_1_6_7_U150 ( .A(npu_inst_pe_1_6_7_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_6_7_int_q_reg_h_1__1_), .S(npu_inst_pe_1_6_7_n4), .Z(
        npu_inst_pe_1_6_7_n21) );
  MUX2_X1 npu_inst_pe_1_6_7_U149 ( .A(npu_inst_pe_1_6_7_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_6_7_int_q_reg_h_3__1_), .S(npu_inst_pe_1_6_7_n4), .Z(
        npu_inst_pe_1_6_7_n20) );
  MUX2_X1 npu_inst_pe_1_6_7_U148 ( .A(npu_inst_pe_1_6_7_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_6_7_int_q_reg_h_5__1_), .S(npu_inst_pe_1_6_7_n4), .Z(
        npu_inst_pe_1_6_7_n19) );
  MUX2_X1 npu_inst_pe_1_6_7_U147 ( .A(npu_inst_pe_1_6_7_n18), .B(
        npu_inst_pe_1_6_7_n15), .S(npu_inst_pe_1_6_7_n8), .Z(
        npu_inst_int_data_x_6__7__0_) );
  MUX2_X1 npu_inst_pe_1_6_7_U146 ( .A(npu_inst_pe_1_6_7_n17), .B(
        npu_inst_pe_1_6_7_n16), .S(npu_inst_pe_1_6_7_n6), .Z(
        npu_inst_pe_1_6_7_n18) );
  MUX2_X1 npu_inst_pe_1_6_7_U145 ( .A(npu_inst_pe_1_6_7_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_6_7_int_q_reg_h_1__0_), .S(npu_inst_pe_1_6_7_n4), .Z(
        npu_inst_pe_1_6_7_n17) );
  MUX2_X1 npu_inst_pe_1_6_7_U144 ( .A(npu_inst_pe_1_6_7_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_6_7_int_q_reg_h_3__0_), .S(npu_inst_pe_1_6_7_n4), .Z(
        npu_inst_pe_1_6_7_n16) );
  MUX2_X1 npu_inst_pe_1_6_7_U143 ( .A(npu_inst_pe_1_6_7_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_6_7_int_q_reg_h_5__0_), .S(npu_inst_pe_1_6_7_n4), .Z(
        npu_inst_pe_1_6_7_n15) );
  XOR2_X1 npu_inst_pe_1_6_7_U142 ( .A(npu_inst_pe_1_6_7_int_data_0_), .B(
        npu_inst_pe_1_6_7_int_q_acc_0_), .Z(npu_inst_pe_1_6_7_N73) );
  AND2_X1 npu_inst_pe_1_6_7_U141 ( .A1(npu_inst_pe_1_6_7_int_q_acc_0_), .A2(
        npu_inst_pe_1_6_7_int_data_0_), .ZN(npu_inst_pe_1_6_7_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_6_7_U140 ( .A(npu_inst_pe_1_6_7_int_q_acc_0_), .B(
        npu_inst_pe_1_6_7_n13), .ZN(npu_inst_pe_1_6_7_N65) );
  OR2_X1 npu_inst_pe_1_6_7_U139 ( .A1(npu_inst_pe_1_6_7_n13), .A2(
        npu_inst_pe_1_6_7_int_q_acc_0_), .ZN(npu_inst_pe_1_6_7_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_6_7_U138 ( .A(npu_inst_pe_1_6_7_int_q_acc_2_), .B(
        npu_inst_pe_1_6_7_add_79_carry_2_), .Z(npu_inst_pe_1_6_7_N75) );
  AND2_X1 npu_inst_pe_1_6_7_U137 ( .A1(npu_inst_pe_1_6_7_add_79_carry_2_), 
        .A2(npu_inst_pe_1_6_7_int_q_acc_2_), .ZN(
        npu_inst_pe_1_6_7_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_6_7_U136 ( .A(npu_inst_pe_1_6_7_int_q_acc_3_), .B(
        npu_inst_pe_1_6_7_add_79_carry_3_), .Z(npu_inst_pe_1_6_7_N76) );
  AND2_X1 npu_inst_pe_1_6_7_U135 ( .A1(npu_inst_pe_1_6_7_add_79_carry_3_), 
        .A2(npu_inst_pe_1_6_7_int_q_acc_3_), .ZN(
        npu_inst_pe_1_6_7_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_6_7_U134 ( .A(npu_inst_pe_1_6_7_int_q_acc_4_), .B(
        npu_inst_pe_1_6_7_add_79_carry_4_), .Z(npu_inst_pe_1_6_7_N77) );
  AND2_X1 npu_inst_pe_1_6_7_U133 ( .A1(npu_inst_pe_1_6_7_add_79_carry_4_), 
        .A2(npu_inst_pe_1_6_7_int_q_acc_4_), .ZN(
        npu_inst_pe_1_6_7_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_6_7_U132 ( .A(npu_inst_pe_1_6_7_int_q_acc_5_), .B(
        npu_inst_pe_1_6_7_add_79_carry_5_), .Z(npu_inst_pe_1_6_7_N78) );
  AND2_X1 npu_inst_pe_1_6_7_U131 ( .A1(npu_inst_pe_1_6_7_add_79_carry_5_), 
        .A2(npu_inst_pe_1_6_7_int_q_acc_5_), .ZN(
        npu_inst_pe_1_6_7_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_6_7_U130 ( .A(npu_inst_pe_1_6_7_int_q_acc_6_), .B(
        npu_inst_pe_1_6_7_add_79_carry_6_), .Z(npu_inst_pe_1_6_7_N79) );
  AND2_X1 npu_inst_pe_1_6_7_U129 ( .A1(npu_inst_pe_1_6_7_add_79_carry_6_), 
        .A2(npu_inst_pe_1_6_7_int_q_acc_6_), .ZN(
        npu_inst_pe_1_6_7_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_6_7_U128 ( .A(npu_inst_pe_1_6_7_int_q_acc_7_), .B(
        npu_inst_pe_1_6_7_add_79_carry_7_), .Z(npu_inst_pe_1_6_7_N80) );
  XNOR2_X1 npu_inst_pe_1_6_7_U127 ( .A(npu_inst_pe_1_6_7_sub_77_carry_2_), .B(
        npu_inst_pe_1_6_7_int_q_acc_2_), .ZN(npu_inst_pe_1_6_7_N67) );
  OR2_X1 npu_inst_pe_1_6_7_U126 ( .A1(npu_inst_pe_1_6_7_int_q_acc_2_), .A2(
        npu_inst_pe_1_6_7_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_6_7_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_6_7_U125 ( .A(npu_inst_pe_1_6_7_sub_77_carry_3_), .B(
        npu_inst_pe_1_6_7_int_q_acc_3_), .ZN(npu_inst_pe_1_6_7_N68) );
  OR2_X1 npu_inst_pe_1_6_7_U124 ( .A1(npu_inst_pe_1_6_7_int_q_acc_3_), .A2(
        npu_inst_pe_1_6_7_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_6_7_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_6_7_U123 ( .A(npu_inst_pe_1_6_7_sub_77_carry_4_), .B(
        npu_inst_pe_1_6_7_int_q_acc_4_), .ZN(npu_inst_pe_1_6_7_N69) );
  OR2_X1 npu_inst_pe_1_6_7_U122 ( .A1(npu_inst_pe_1_6_7_int_q_acc_4_), .A2(
        npu_inst_pe_1_6_7_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_6_7_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_6_7_U121 ( .A(npu_inst_pe_1_6_7_sub_77_carry_5_), .B(
        npu_inst_pe_1_6_7_int_q_acc_5_), .ZN(npu_inst_pe_1_6_7_N70) );
  OR2_X1 npu_inst_pe_1_6_7_U120 ( .A1(npu_inst_pe_1_6_7_int_q_acc_5_), .A2(
        npu_inst_pe_1_6_7_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_6_7_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_6_7_U119 ( .A(npu_inst_pe_1_6_7_sub_77_carry_6_), .B(
        npu_inst_pe_1_6_7_int_q_acc_6_), .ZN(npu_inst_pe_1_6_7_N71) );
  OR2_X1 npu_inst_pe_1_6_7_U118 ( .A1(npu_inst_pe_1_6_7_int_q_acc_6_), .A2(
        npu_inst_pe_1_6_7_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_6_7_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_6_7_U117 ( .A(npu_inst_pe_1_6_7_int_q_acc_7_), .B(
        npu_inst_pe_1_6_7_sub_77_carry_7_), .ZN(npu_inst_pe_1_6_7_N72) );
  INV_X1 npu_inst_pe_1_6_7_U116 ( .A(npu_inst_n75), .ZN(npu_inst_pe_1_6_7_n7)
         );
  INV_X1 npu_inst_pe_1_6_7_U115 ( .A(npu_inst_pe_1_6_7_n7), .ZN(
        npu_inst_pe_1_6_7_n6) );
  INV_X1 npu_inst_pe_1_6_7_U114 ( .A(npu_inst_n53), .ZN(npu_inst_pe_1_6_7_n3)
         );
  AOI22_X1 npu_inst_pe_1_6_7_U113 ( .A1(npu_inst_int_data_y_7__7__0_), .A2(
        npu_inst_pe_1_6_7_n58), .B1(npu_inst_pe_1_6_7_n114), .B2(
        npu_inst_pe_1_6_7_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_6_7_n57) );
  INV_X1 npu_inst_pe_1_6_7_U112 ( .A(npu_inst_pe_1_6_7_n57), .ZN(
        npu_inst_pe_1_6_7_n108) );
  AOI22_X1 npu_inst_pe_1_6_7_U111 ( .A1(npu_inst_int_data_y_7__7__0_), .A2(
        npu_inst_pe_1_6_7_n54), .B1(npu_inst_pe_1_6_7_n115), .B2(
        npu_inst_pe_1_6_7_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_6_7_n53) );
  INV_X1 npu_inst_pe_1_6_7_U110 ( .A(npu_inst_pe_1_6_7_n53), .ZN(
        npu_inst_pe_1_6_7_n109) );
  AOI22_X1 npu_inst_pe_1_6_7_U107 ( .A1(npu_inst_int_data_y_7__7__0_), .A2(
        npu_inst_pe_1_6_7_n50), .B1(npu_inst_pe_1_6_7_n116), .B2(
        npu_inst_pe_1_6_7_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_6_7_n49) );
  INV_X1 npu_inst_pe_1_6_7_U106 ( .A(npu_inst_pe_1_6_7_n49), .ZN(
        npu_inst_pe_1_6_7_n110) );
  AOI22_X1 npu_inst_pe_1_6_7_U105 ( .A1(npu_inst_int_data_y_7__7__0_), .A2(
        npu_inst_pe_1_6_7_n46), .B1(npu_inst_pe_1_6_7_n117), .B2(
        npu_inst_pe_1_6_7_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_6_7_n45) );
  INV_X1 npu_inst_pe_1_6_7_U104 ( .A(npu_inst_pe_1_6_7_n45), .ZN(
        npu_inst_pe_1_6_7_n111) );
  AOI22_X1 npu_inst_pe_1_6_7_U103 ( .A1(npu_inst_int_data_y_7__7__0_), .A2(
        npu_inst_pe_1_6_7_n42), .B1(npu_inst_pe_1_6_7_n119), .B2(
        npu_inst_pe_1_6_7_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_6_7_n41) );
  INV_X1 npu_inst_pe_1_6_7_U102 ( .A(npu_inst_pe_1_6_7_n41), .ZN(
        npu_inst_pe_1_6_7_n112) );
  AOI22_X1 npu_inst_pe_1_6_7_U101 ( .A1(npu_inst_int_data_y_7__7__1_), .A2(
        npu_inst_pe_1_6_7_n58), .B1(npu_inst_pe_1_6_7_n114), .B2(
        npu_inst_pe_1_6_7_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_6_7_n59) );
  INV_X1 npu_inst_pe_1_6_7_U100 ( .A(npu_inst_pe_1_6_7_n59), .ZN(
        npu_inst_pe_1_6_7_n102) );
  AOI22_X1 npu_inst_pe_1_6_7_U99 ( .A1(npu_inst_int_data_y_7__7__1_), .A2(
        npu_inst_pe_1_6_7_n54), .B1(npu_inst_pe_1_6_7_n115), .B2(
        npu_inst_pe_1_6_7_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_6_7_n55) );
  INV_X1 npu_inst_pe_1_6_7_U98 ( .A(npu_inst_pe_1_6_7_n55), .ZN(
        npu_inst_pe_1_6_7_n103) );
  AOI22_X1 npu_inst_pe_1_6_7_U97 ( .A1(npu_inst_int_data_y_7__7__1_), .A2(
        npu_inst_pe_1_6_7_n50), .B1(npu_inst_pe_1_6_7_n116), .B2(
        npu_inst_pe_1_6_7_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_6_7_n51) );
  INV_X1 npu_inst_pe_1_6_7_U96 ( .A(npu_inst_pe_1_6_7_n51), .ZN(
        npu_inst_pe_1_6_7_n104) );
  AOI22_X1 npu_inst_pe_1_6_7_U95 ( .A1(npu_inst_int_data_y_7__7__1_), .A2(
        npu_inst_pe_1_6_7_n46), .B1(npu_inst_pe_1_6_7_n117), .B2(
        npu_inst_pe_1_6_7_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_6_7_n47) );
  INV_X1 npu_inst_pe_1_6_7_U94 ( .A(npu_inst_pe_1_6_7_n47), .ZN(
        npu_inst_pe_1_6_7_n105) );
  AOI22_X1 npu_inst_pe_1_6_7_U93 ( .A1(npu_inst_int_data_y_7__7__1_), .A2(
        npu_inst_pe_1_6_7_n42), .B1(npu_inst_pe_1_6_7_n119), .B2(
        npu_inst_pe_1_6_7_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_6_7_n43) );
  INV_X1 npu_inst_pe_1_6_7_U92 ( .A(npu_inst_pe_1_6_7_n43), .ZN(
        npu_inst_pe_1_6_7_n106) );
  AOI22_X1 npu_inst_pe_1_6_7_U91 ( .A1(npu_inst_pe_1_6_7_n38), .A2(
        npu_inst_int_data_y_7__7__1_), .B1(npu_inst_pe_1_6_7_n118), .B2(
        npu_inst_pe_1_6_7_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_6_7_n39) );
  INV_X1 npu_inst_pe_1_6_7_U90 ( .A(npu_inst_pe_1_6_7_n39), .ZN(
        npu_inst_pe_1_6_7_n107) );
  AOI22_X1 npu_inst_pe_1_6_7_U89 ( .A1(npu_inst_pe_1_6_7_n38), .A2(
        npu_inst_int_data_y_7__7__0_), .B1(npu_inst_pe_1_6_7_n118), .B2(
        npu_inst_pe_1_6_7_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_6_7_n37) );
  INV_X1 npu_inst_pe_1_6_7_U88 ( .A(npu_inst_pe_1_6_7_n37), .ZN(
        npu_inst_pe_1_6_7_n113) );
  AND2_X1 npu_inst_pe_1_6_7_U87 ( .A1(npu_inst_pe_1_6_7_N93), .A2(npu_inst_n53), .ZN(npu_inst_int_data_y_6__7__0_) );
  AND2_X1 npu_inst_pe_1_6_7_U86 ( .A1(npu_inst_n53), .A2(npu_inst_pe_1_6_7_N94), .ZN(npu_inst_int_data_y_6__7__1_) );
  NOR3_X1 npu_inst_pe_1_6_7_U85 ( .A1(npu_inst_pe_1_6_7_n26), .A2(npu_inst_n53), .A3(npu_inst_int_ckg[8]), .ZN(npu_inst_pe_1_6_7_n85) );
  OR2_X1 npu_inst_pe_1_6_7_U84 ( .A1(npu_inst_pe_1_6_7_n85), .A2(
        npu_inst_pe_1_6_7_n2), .ZN(npu_inst_pe_1_6_7_N84) );
  AND2_X1 npu_inst_pe_1_6_7_U83 ( .A1(npu_inst_pe_1_6_7_int_q_acc_0_), .A2(
        npu_inst_pe_1_6_7_n1), .ZN(npu_inst_int_data_res_6__7__0_) );
  AND2_X1 npu_inst_pe_1_6_7_U82 ( .A1(npu_inst_pe_1_6_7_n2), .A2(
        npu_inst_pe_1_6_7_int_q_acc_7_), .ZN(npu_inst_int_data_res_6__7__7_)
         );
  AND2_X1 npu_inst_pe_1_6_7_U81 ( .A1(npu_inst_pe_1_6_7_int_q_acc_1_), .A2(
        npu_inst_pe_1_6_7_n1), .ZN(npu_inst_int_data_res_6__7__1_) );
  AND2_X1 npu_inst_pe_1_6_7_U80 ( .A1(npu_inst_pe_1_6_7_int_q_acc_2_), .A2(
        npu_inst_pe_1_6_7_n1), .ZN(npu_inst_int_data_res_6__7__2_) );
  AND2_X1 npu_inst_pe_1_6_7_U79 ( .A1(npu_inst_pe_1_6_7_int_q_acc_3_), .A2(
        npu_inst_pe_1_6_7_n2), .ZN(npu_inst_int_data_res_6__7__3_) );
  AND2_X1 npu_inst_pe_1_6_7_U78 ( .A1(npu_inst_pe_1_6_7_int_q_acc_4_), .A2(
        npu_inst_pe_1_6_7_n2), .ZN(npu_inst_int_data_res_6__7__4_) );
  AND2_X1 npu_inst_pe_1_6_7_U77 ( .A1(npu_inst_pe_1_6_7_int_q_acc_5_), .A2(
        npu_inst_pe_1_6_7_n2), .ZN(npu_inst_int_data_res_6__7__5_) );
  AND2_X1 npu_inst_pe_1_6_7_U76 ( .A1(npu_inst_pe_1_6_7_int_q_acc_6_), .A2(
        npu_inst_pe_1_6_7_n2), .ZN(npu_inst_int_data_res_6__7__6_) );
  AOI222_X1 npu_inst_pe_1_6_7_U75 ( .A1(npu_inst_int_data_res_7__7__0_), .A2(
        npu_inst_pe_1_6_7_n1), .B1(npu_inst_pe_1_6_7_N73), .B2(
        npu_inst_pe_1_6_7_n76), .C1(npu_inst_pe_1_6_7_N65), .C2(
        npu_inst_pe_1_6_7_n77), .ZN(npu_inst_pe_1_6_7_n84) );
  INV_X1 npu_inst_pe_1_6_7_U74 ( .A(npu_inst_pe_1_6_7_n84), .ZN(
        npu_inst_pe_1_6_7_n101) );
  AOI222_X1 npu_inst_pe_1_6_7_U73 ( .A1(npu_inst_int_data_res_7__7__7_), .A2(
        npu_inst_pe_1_6_7_n1), .B1(npu_inst_pe_1_6_7_N80), .B2(
        npu_inst_pe_1_6_7_n76), .C1(npu_inst_pe_1_6_7_N72), .C2(
        npu_inst_pe_1_6_7_n77), .ZN(npu_inst_pe_1_6_7_n75) );
  INV_X1 npu_inst_pe_1_6_7_U72 ( .A(npu_inst_pe_1_6_7_n75), .ZN(
        npu_inst_pe_1_6_7_n33) );
  AOI222_X1 npu_inst_pe_1_6_7_U71 ( .A1(npu_inst_int_data_res_7__7__1_), .A2(
        npu_inst_pe_1_6_7_n1), .B1(npu_inst_pe_1_6_7_N74), .B2(
        npu_inst_pe_1_6_7_n76), .C1(npu_inst_pe_1_6_7_N66), .C2(
        npu_inst_pe_1_6_7_n77), .ZN(npu_inst_pe_1_6_7_n83) );
  INV_X1 npu_inst_pe_1_6_7_U70 ( .A(npu_inst_pe_1_6_7_n83), .ZN(
        npu_inst_pe_1_6_7_n100) );
  AOI222_X1 npu_inst_pe_1_6_7_U69 ( .A1(npu_inst_int_data_res_7__7__2_), .A2(
        npu_inst_pe_1_6_7_n1), .B1(npu_inst_pe_1_6_7_N75), .B2(
        npu_inst_pe_1_6_7_n76), .C1(npu_inst_pe_1_6_7_N67), .C2(
        npu_inst_pe_1_6_7_n77), .ZN(npu_inst_pe_1_6_7_n82) );
  INV_X1 npu_inst_pe_1_6_7_U68 ( .A(npu_inst_pe_1_6_7_n82), .ZN(
        npu_inst_pe_1_6_7_n99) );
  AOI222_X1 npu_inst_pe_1_6_7_U67 ( .A1(npu_inst_int_data_res_7__7__3_), .A2(
        npu_inst_pe_1_6_7_n1), .B1(npu_inst_pe_1_6_7_N76), .B2(
        npu_inst_pe_1_6_7_n76), .C1(npu_inst_pe_1_6_7_N68), .C2(
        npu_inst_pe_1_6_7_n77), .ZN(npu_inst_pe_1_6_7_n81) );
  INV_X1 npu_inst_pe_1_6_7_U66 ( .A(npu_inst_pe_1_6_7_n81), .ZN(
        npu_inst_pe_1_6_7_n98) );
  AOI222_X1 npu_inst_pe_1_6_7_U65 ( .A1(npu_inst_int_data_res_7__7__4_), .A2(
        npu_inst_pe_1_6_7_n1), .B1(npu_inst_pe_1_6_7_N77), .B2(
        npu_inst_pe_1_6_7_n76), .C1(npu_inst_pe_1_6_7_N69), .C2(
        npu_inst_pe_1_6_7_n77), .ZN(npu_inst_pe_1_6_7_n80) );
  INV_X1 npu_inst_pe_1_6_7_U64 ( .A(npu_inst_pe_1_6_7_n80), .ZN(
        npu_inst_pe_1_6_7_n36) );
  AOI222_X1 npu_inst_pe_1_6_7_U63 ( .A1(npu_inst_int_data_res_7__7__5_), .A2(
        npu_inst_pe_1_6_7_n1), .B1(npu_inst_pe_1_6_7_N78), .B2(
        npu_inst_pe_1_6_7_n76), .C1(npu_inst_pe_1_6_7_N70), .C2(
        npu_inst_pe_1_6_7_n77), .ZN(npu_inst_pe_1_6_7_n79) );
  INV_X1 npu_inst_pe_1_6_7_U62 ( .A(npu_inst_pe_1_6_7_n79), .ZN(
        npu_inst_pe_1_6_7_n35) );
  AOI222_X1 npu_inst_pe_1_6_7_U61 ( .A1(npu_inst_int_data_res_7__7__6_), .A2(
        npu_inst_pe_1_6_7_n1), .B1(npu_inst_pe_1_6_7_N79), .B2(
        npu_inst_pe_1_6_7_n76), .C1(npu_inst_pe_1_6_7_N71), .C2(
        npu_inst_pe_1_6_7_n77), .ZN(npu_inst_pe_1_6_7_n78) );
  INV_X1 npu_inst_pe_1_6_7_U60 ( .A(npu_inst_pe_1_6_7_n78), .ZN(
        npu_inst_pe_1_6_7_n34) );
  INV_X1 npu_inst_pe_1_6_7_U59 ( .A(npu_inst_pe_1_6_7_int_data_1_), .ZN(
        npu_inst_pe_1_6_7_n14) );
  AND2_X1 npu_inst_pe_1_6_7_U58 ( .A1(npu_inst_int_data_x_6__7__1_), .A2(
        npu_inst_pe_1_6_7_int_q_weight_1_), .ZN(npu_inst_pe_1_6_7_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_6_7_U57 ( .A1(npu_inst_int_data_x_6__7__0_), .A2(
        npu_inst_pe_1_6_7_int_q_weight_1_), .ZN(npu_inst_pe_1_6_7_int_data_0_)
         );
  NAND2_X1 npu_inst_pe_1_6_7_U56 ( .A1(npu_inst_pe_1_6_7_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_6_7_n60), .ZN(npu_inst_pe_1_6_7_n74) );
  OAI21_X1 npu_inst_pe_1_6_7_U55 ( .B1(npu_inst_pe_1_6_7_n63), .B2(
        npu_inst_pe_1_6_7_n60), .A(npu_inst_pe_1_6_7_n74), .ZN(
        npu_inst_pe_1_6_7_n97) );
  NAND2_X1 npu_inst_pe_1_6_7_U54 ( .A1(npu_inst_pe_1_6_7_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_6_7_n60), .ZN(npu_inst_pe_1_6_7_n73) );
  OAI21_X1 npu_inst_pe_1_6_7_U53 ( .B1(npu_inst_pe_1_6_7_n61), .B2(
        npu_inst_pe_1_6_7_n60), .A(npu_inst_pe_1_6_7_n73), .ZN(
        npu_inst_pe_1_6_7_n96) );
  NAND2_X1 npu_inst_pe_1_6_7_U52 ( .A1(npu_inst_pe_1_6_7_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_6_7_n56), .ZN(npu_inst_pe_1_6_7_n72) );
  OAI21_X1 npu_inst_pe_1_6_7_U51 ( .B1(npu_inst_pe_1_6_7_n63), .B2(
        npu_inst_pe_1_6_7_n56), .A(npu_inst_pe_1_6_7_n72), .ZN(
        npu_inst_pe_1_6_7_n95) );
  NAND2_X1 npu_inst_pe_1_6_7_U50 ( .A1(npu_inst_pe_1_6_7_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_6_7_n56), .ZN(npu_inst_pe_1_6_7_n71) );
  OAI21_X1 npu_inst_pe_1_6_7_U49 ( .B1(npu_inst_pe_1_6_7_n61), .B2(
        npu_inst_pe_1_6_7_n56), .A(npu_inst_pe_1_6_7_n71), .ZN(
        npu_inst_pe_1_6_7_n94) );
  NAND2_X1 npu_inst_pe_1_6_7_U48 ( .A1(npu_inst_pe_1_6_7_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_6_7_n52), .ZN(npu_inst_pe_1_6_7_n70) );
  OAI21_X1 npu_inst_pe_1_6_7_U47 ( .B1(npu_inst_pe_1_6_7_n63), .B2(
        npu_inst_pe_1_6_7_n52), .A(npu_inst_pe_1_6_7_n70), .ZN(
        npu_inst_pe_1_6_7_n93) );
  NAND2_X1 npu_inst_pe_1_6_7_U46 ( .A1(npu_inst_pe_1_6_7_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_6_7_n52), .ZN(npu_inst_pe_1_6_7_n69) );
  OAI21_X1 npu_inst_pe_1_6_7_U45 ( .B1(npu_inst_pe_1_6_7_n61), .B2(
        npu_inst_pe_1_6_7_n52), .A(npu_inst_pe_1_6_7_n69), .ZN(
        npu_inst_pe_1_6_7_n92) );
  NAND2_X1 npu_inst_pe_1_6_7_U44 ( .A1(npu_inst_pe_1_6_7_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_6_7_n48), .ZN(npu_inst_pe_1_6_7_n68) );
  OAI21_X1 npu_inst_pe_1_6_7_U43 ( .B1(npu_inst_pe_1_6_7_n63), .B2(
        npu_inst_pe_1_6_7_n48), .A(npu_inst_pe_1_6_7_n68), .ZN(
        npu_inst_pe_1_6_7_n91) );
  NAND2_X1 npu_inst_pe_1_6_7_U42 ( .A1(npu_inst_pe_1_6_7_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_6_7_n48), .ZN(npu_inst_pe_1_6_7_n67) );
  OAI21_X1 npu_inst_pe_1_6_7_U41 ( .B1(npu_inst_pe_1_6_7_n61), .B2(
        npu_inst_pe_1_6_7_n48), .A(npu_inst_pe_1_6_7_n67), .ZN(
        npu_inst_pe_1_6_7_n90) );
  NAND2_X1 npu_inst_pe_1_6_7_U40 ( .A1(npu_inst_pe_1_6_7_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_6_7_n44), .ZN(npu_inst_pe_1_6_7_n66) );
  OAI21_X1 npu_inst_pe_1_6_7_U39 ( .B1(npu_inst_pe_1_6_7_n63), .B2(
        npu_inst_pe_1_6_7_n44), .A(npu_inst_pe_1_6_7_n66), .ZN(
        npu_inst_pe_1_6_7_n89) );
  NAND2_X1 npu_inst_pe_1_6_7_U38 ( .A1(npu_inst_pe_1_6_7_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_6_7_n44), .ZN(npu_inst_pe_1_6_7_n65) );
  OAI21_X1 npu_inst_pe_1_6_7_U37 ( .B1(npu_inst_pe_1_6_7_n61), .B2(
        npu_inst_pe_1_6_7_n44), .A(npu_inst_pe_1_6_7_n65), .ZN(
        npu_inst_pe_1_6_7_n88) );
  NAND2_X1 npu_inst_pe_1_6_7_U36 ( .A1(npu_inst_pe_1_6_7_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_6_7_n40), .ZN(npu_inst_pe_1_6_7_n64) );
  OAI21_X1 npu_inst_pe_1_6_7_U35 ( .B1(npu_inst_pe_1_6_7_n63), .B2(
        npu_inst_pe_1_6_7_n40), .A(npu_inst_pe_1_6_7_n64), .ZN(
        npu_inst_pe_1_6_7_n87) );
  NAND2_X1 npu_inst_pe_1_6_7_U34 ( .A1(npu_inst_pe_1_6_7_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_6_7_n40), .ZN(npu_inst_pe_1_6_7_n62) );
  OAI21_X1 npu_inst_pe_1_6_7_U33 ( .B1(npu_inst_pe_1_6_7_n61), .B2(
        npu_inst_pe_1_6_7_n40), .A(npu_inst_pe_1_6_7_n62), .ZN(
        npu_inst_pe_1_6_7_n86) );
  INV_X1 npu_inst_pe_1_6_7_U32 ( .A(npu_inst_pe_1_6_7_int_data_0_), .ZN(
        npu_inst_pe_1_6_7_n13) );
  INV_X1 npu_inst_pe_1_6_7_U31 ( .A(npu_inst_n67), .ZN(npu_inst_pe_1_6_7_n5)
         );
  AOI22_X1 npu_inst_pe_1_6_7_U30 ( .A1(npu_inst_n53), .A2(
        npu_inst_int_data_y_7__7__1_), .B1(npu_inst_pe_1_6_7_n3), .B2(
        int_i_data_h_npu7[1]), .ZN(npu_inst_pe_1_6_7_n63) );
  AOI22_X1 npu_inst_pe_1_6_7_U29 ( .A1(npu_inst_n53), .A2(
        npu_inst_int_data_y_7__7__0_), .B1(npu_inst_pe_1_6_7_n3), .B2(
        int_i_data_h_npu7[0]), .ZN(npu_inst_pe_1_6_7_n61) );
  OR3_X1 npu_inst_pe_1_6_7_U28 ( .A1(npu_inst_pe_1_6_7_n6), .A2(
        npu_inst_pe_1_6_7_n8), .A3(npu_inst_pe_1_6_7_n5), .ZN(
        npu_inst_pe_1_6_7_n56) );
  OR3_X1 npu_inst_pe_1_6_7_U27 ( .A1(npu_inst_pe_1_6_7_n5), .A2(
        npu_inst_pe_1_6_7_n8), .A3(npu_inst_pe_1_6_7_n7), .ZN(
        npu_inst_pe_1_6_7_n48) );
  INV_X1 npu_inst_pe_1_6_7_U26 ( .A(npu_inst_pe_1_6_7_n5), .ZN(
        npu_inst_pe_1_6_7_n4) );
  INV_X1 npu_inst_pe_1_6_7_U25 ( .A(npu_inst_n122), .ZN(npu_inst_pe_1_6_7_n12)
         );
  OR3_X1 npu_inst_pe_1_6_7_U24 ( .A1(npu_inst_pe_1_6_7_n4), .A2(
        npu_inst_pe_1_6_7_n8), .A3(npu_inst_pe_1_6_7_n7), .ZN(
        npu_inst_pe_1_6_7_n52) );
  OR3_X1 npu_inst_pe_1_6_7_U23 ( .A1(npu_inst_pe_1_6_7_n6), .A2(
        npu_inst_pe_1_6_7_n8), .A3(npu_inst_pe_1_6_7_n4), .ZN(
        npu_inst_pe_1_6_7_n60) );
  NOR2_X1 npu_inst_pe_1_6_7_U22 ( .A1(npu_inst_pe_1_6_7_n60), .A2(
        npu_inst_pe_1_6_7_n3), .ZN(npu_inst_pe_1_6_7_n58) );
  NOR2_X1 npu_inst_pe_1_6_7_U21 ( .A1(npu_inst_pe_1_6_7_n56), .A2(
        npu_inst_pe_1_6_7_n3), .ZN(npu_inst_pe_1_6_7_n54) );
  NOR2_X1 npu_inst_pe_1_6_7_U20 ( .A1(npu_inst_pe_1_6_7_n52), .A2(
        npu_inst_pe_1_6_7_n3), .ZN(npu_inst_pe_1_6_7_n50) );
  NOR2_X1 npu_inst_pe_1_6_7_U19 ( .A1(npu_inst_pe_1_6_7_n48), .A2(
        npu_inst_pe_1_6_7_n3), .ZN(npu_inst_pe_1_6_7_n46) );
  NOR2_X1 npu_inst_pe_1_6_7_U18 ( .A1(npu_inst_pe_1_6_7_n40), .A2(
        npu_inst_pe_1_6_7_n3), .ZN(npu_inst_pe_1_6_7_n38) );
  NOR2_X1 npu_inst_pe_1_6_7_U17 ( .A1(npu_inst_pe_1_6_7_n44), .A2(
        npu_inst_pe_1_6_7_n3), .ZN(npu_inst_pe_1_6_7_n42) );
  BUF_X1 npu_inst_pe_1_6_7_U16 ( .A(npu_inst_n94), .Z(npu_inst_pe_1_6_7_n8) );
  BUF_X1 npu_inst_pe_1_6_7_U15 ( .A(npu_inst_pe_1_6_7_n12), .Z(
        npu_inst_pe_1_6_7_n11) );
  BUF_X1 npu_inst_pe_1_6_7_U14 ( .A(npu_inst_pe_1_6_7_n12), .Z(
        npu_inst_pe_1_6_7_n10) );
  BUF_X1 npu_inst_pe_1_6_7_U13 ( .A(npu_inst_pe_1_6_7_n12), .Z(
        npu_inst_pe_1_6_7_n9) );
  INV_X1 npu_inst_pe_1_6_7_U12 ( .A(npu_inst_pe_1_6_7_n38), .ZN(
        npu_inst_pe_1_6_7_n118) );
  INV_X1 npu_inst_pe_1_6_7_U11 ( .A(npu_inst_pe_1_6_7_n58), .ZN(
        npu_inst_pe_1_6_7_n114) );
  INV_X1 npu_inst_pe_1_6_7_U10 ( .A(npu_inst_pe_1_6_7_n54), .ZN(
        npu_inst_pe_1_6_7_n115) );
  INV_X1 npu_inst_pe_1_6_7_U9 ( .A(npu_inst_pe_1_6_7_n50), .ZN(
        npu_inst_pe_1_6_7_n116) );
  INV_X1 npu_inst_pe_1_6_7_U8 ( .A(npu_inst_pe_1_6_7_n46), .ZN(
        npu_inst_pe_1_6_7_n117) );
  INV_X1 npu_inst_pe_1_6_7_U7 ( .A(npu_inst_pe_1_6_7_n42), .ZN(
        npu_inst_pe_1_6_7_n119) );
  BUF_X1 npu_inst_pe_1_6_7_U6 ( .A(npu_inst_n11), .Z(npu_inst_pe_1_6_7_n2) );
  BUF_X1 npu_inst_pe_1_6_7_U5 ( .A(npu_inst_n11), .Z(npu_inst_pe_1_6_7_n1) );
  NOR2_X1 npu_inst_pe_1_6_7_U4 ( .A1(npu_inst_pe_1_6_7_int_q_weight_0_), .A2(
        npu_inst_pe_1_6_7_n1), .ZN(npu_inst_pe_1_6_7_n76) );
  NOR2_X1 npu_inst_pe_1_6_7_U3 ( .A1(npu_inst_pe_1_6_7_n27), .A2(
        npu_inst_pe_1_6_7_n1), .ZN(npu_inst_pe_1_6_7_n77) );
  FA_X1 npu_inst_pe_1_6_7_sub_77_U2_1 ( .A(npu_inst_pe_1_6_7_int_q_acc_1_), 
        .B(npu_inst_pe_1_6_7_n14), .CI(npu_inst_pe_1_6_7_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_6_7_sub_77_carry_2_), .S(npu_inst_pe_1_6_7_N66) );
  FA_X1 npu_inst_pe_1_6_7_add_79_U1_1 ( .A(npu_inst_pe_1_6_7_int_q_acc_1_), 
        .B(npu_inst_pe_1_6_7_int_data_1_), .CI(
        npu_inst_pe_1_6_7_add_79_carry_1_), .CO(
        npu_inst_pe_1_6_7_add_79_carry_2_), .S(npu_inst_pe_1_6_7_N74) );
  NAND3_X1 npu_inst_pe_1_6_7_U109 ( .A1(npu_inst_pe_1_6_7_n5), .A2(
        npu_inst_pe_1_6_7_n7), .A3(npu_inst_pe_1_6_7_n8), .ZN(
        npu_inst_pe_1_6_7_n44) );
  NAND3_X1 npu_inst_pe_1_6_7_U108 ( .A1(npu_inst_pe_1_6_7_n4), .A2(
        npu_inst_pe_1_6_7_n7), .A3(npu_inst_pe_1_6_7_n8), .ZN(
        npu_inst_pe_1_6_7_n40) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_6_7_n34), .CK(
        npu_inst_pe_1_6_7_net3028), .RN(npu_inst_pe_1_6_7_n9), .Q(
        npu_inst_pe_1_6_7_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_6_7_n35), .CK(
        npu_inst_pe_1_6_7_net3028), .RN(npu_inst_pe_1_6_7_n9), .Q(
        npu_inst_pe_1_6_7_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_6_7_n36), .CK(
        npu_inst_pe_1_6_7_net3028), .RN(npu_inst_pe_1_6_7_n9), .Q(
        npu_inst_pe_1_6_7_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_6_7_n98), .CK(
        npu_inst_pe_1_6_7_net3028), .RN(npu_inst_pe_1_6_7_n9), .Q(
        npu_inst_pe_1_6_7_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_6_7_n99), .CK(
        npu_inst_pe_1_6_7_net3028), .RN(npu_inst_pe_1_6_7_n9), .Q(
        npu_inst_pe_1_6_7_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_6_7_n100), 
        .CK(npu_inst_pe_1_6_7_net3028), .RN(npu_inst_pe_1_6_7_n9), .Q(
        npu_inst_pe_1_6_7_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_6_7_n33), .CK(
        npu_inst_pe_1_6_7_net3028), .RN(npu_inst_pe_1_6_7_n9), .Q(
        npu_inst_pe_1_6_7_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_6_7_n101), 
        .CK(npu_inst_pe_1_6_7_net3028), .RN(npu_inst_pe_1_6_7_n9), .Q(
        npu_inst_pe_1_6_7_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_weight_reg_0_ ( .D(npu_inst_n108), .CK(
        npu_inst_pe_1_6_7_net3034), .RN(npu_inst_pe_1_6_7_n9), .Q(
        npu_inst_pe_1_6_7_int_q_weight_0_), .QN(npu_inst_pe_1_6_7_n27) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_weight_reg_1_ ( .D(npu_inst_n114), .CK(
        npu_inst_pe_1_6_7_net3034), .RN(npu_inst_pe_1_6_7_n9), .Q(
        npu_inst_pe_1_6_7_int_q_weight_1_), .QN(npu_inst_pe_1_6_7_n26) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_6_7_n113), 
        .CK(npu_inst_pe_1_6_7_net3034), .RN(npu_inst_pe_1_6_7_n9), .Q(
        npu_inst_pe_1_6_7_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_6_7_n107), 
        .CK(npu_inst_pe_1_6_7_net3034), .RN(npu_inst_pe_1_6_7_n9), .Q(
        npu_inst_pe_1_6_7_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_6_7_n112), 
        .CK(npu_inst_pe_1_6_7_net3034), .RN(npu_inst_pe_1_6_7_n10), .Q(
        npu_inst_pe_1_6_7_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_6_7_n106), 
        .CK(npu_inst_pe_1_6_7_net3034), .RN(npu_inst_pe_1_6_7_n10), .Q(
        npu_inst_pe_1_6_7_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_6_7_n111), 
        .CK(npu_inst_pe_1_6_7_net3034), .RN(npu_inst_pe_1_6_7_n10), .Q(
        npu_inst_pe_1_6_7_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_6_7_n105), 
        .CK(npu_inst_pe_1_6_7_net3034), .RN(npu_inst_pe_1_6_7_n10), .Q(
        npu_inst_pe_1_6_7_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_6_7_n110), 
        .CK(npu_inst_pe_1_6_7_net3034), .RN(npu_inst_pe_1_6_7_n10), .Q(
        npu_inst_pe_1_6_7_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_6_7_n104), 
        .CK(npu_inst_pe_1_6_7_net3034), .RN(npu_inst_pe_1_6_7_n10), .Q(
        npu_inst_pe_1_6_7_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_6_7_n109), 
        .CK(npu_inst_pe_1_6_7_net3034), .RN(npu_inst_pe_1_6_7_n10), .Q(
        npu_inst_pe_1_6_7_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_6_7_n103), 
        .CK(npu_inst_pe_1_6_7_net3034), .RN(npu_inst_pe_1_6_7_n10), .Q(
        npu_inst_pe_1_6_7_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_6_7_n108), 
        .CK(npu_inst_pe_1_6_7_net3034), .RN(npu_inst_pe_1_6_7_n10), .Q(
        npu_inst_pe_1_6_7_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_6_7_n102), 
        .CK(npu_inst_pe_1_6_7_net3034), .RN(npu_inst_pe_1_6_7_n10), .Q(
        npu_inst_pe_1_6_7_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_6_7_n86), 
        .CK(npu_inst_pe_1_6_7_net3034), .RN(npu_inst_pe_1_6_7_n10), .Q(
        npu_inst_pe_1_6_7_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_6_7_n87), 
        .CK(npu_inst_pe_1_6_7_net3034), .RN(npu_inst_pe_1_6_7_n10), .Q(
        npu_inst_pe_1_6_7_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_6_7_n88), 
        .CK(npu_inst_pe_1_6_7_net3034), .RN(npu_inst_pe_1_6_7_n11), .Q(
        npu_inst_pe_1_6_7_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_6_7_n89), 
        .CK(npu_inst_pe_1_6_7_net3034), .RN(npu_inst_pe_1_6_7_n11), .Q(
        npu_inst_pe_1_6_7_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_6_7_n90), 
        .CK(npu_inst_pe_1_6_7_net3034), .RN(npu_inst_pe_1_6_7_n11), .Q(
        npu_inst_pe_1_6_7_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_6_7_n91), 
        .CK(npu_inst_pe_1_6_7_net3034), .RN(npu_inst_pe_1_6_7_n11), .Q(
        npu_inst_pe_1_6_7_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_6_7_n92), 
        .CK(npu_inst_pe_1_6_7_net3034), .RN(npu_inst_pe_1_6_7_n11), .Q(
        npu_inst_pe_1_6_7_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_6_7_n93), 
        .CK(npu_inst_pe_1_6_7_net3034), .RN(npu_inst_pe_1_6_7_n11), .Q(
        npu_inst_pe_1_6_7_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_6_7_n94), 
        .CK(npu_inst_pe_1_6_7_net3034), .RN(npu_inst_pe_1_6_7_n11), .Q(
        npu_inst_pe_1_6_7_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_6_7_n95), 
        .CK(npu_inst_pe_1_6_7_net3034), .RN(npu_inst_pe_1_6_7_n11), .Q(
        npu_inst_pe_1_6_7_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_6_7_n96), 
        .CK(npu_inst_pe_1_6_7_net3034), .RN(npu_inst_pe_1_6_7_n11), .Q(
        npu_inst_pe_1_6_7_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_6_7_n97), 
        .CK(npu_inst_pe_1_6_7_net3034), .RN(npu_inst_pe_1_6_7_n11), .Q(
        npu_inst_pe_1_6_7_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_6_7_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_6_7_N84), .SE(1'b0), .GCK(npu_inst_pe_1_6_7_net3028) );
  CLKGATETST_X1 npu_inst_pe_1_6_7_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n61), .SE(1'b0), .GCK(npu_inst_pe_1_6_7_net3034) );
  MUX2_X1 npu_inst_pe_1_7_0_U162 ( .A(npu_inst_pe_1_7_0_n32), .B(
        npu_inst_pe_1_7_0_n29), .S(npu_inst_pe_1_7_0_n8), .Z(
        npu_inst_pe_1_7_0_N93) );
  MUX2_X1 npu_inst_pe_1_7_0_U161 ( .A(npu_inst_pe_1_7_0_n31), .B(
        npu_inst_pe_1_7_0_n30), .S(npu_inst_pe_1_7_0_n6), .Z(
        npu_inst_pe_1_7_0_n32) );
  MUX2_X1 npu_inst_pe_1_7_0_U160 ( .A(npu_inst_pe_1_7_0_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_7_0_int_q_reg_v_1__0_), .S(npu_inst_pe_1_7_0_n4), .Z(
        npu_inst_pe_1_7_0_n31) );
  MUX2_X1 npu_inst_pe_1_7_0_U159 ( .A(npu_inst_pe_1_7_0_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_7_0_int_q_reg_v_3__0_), .S(npu_inst_pe_1_7_0_n4), .Z(
        npu_inst_pe_1_7_0_n30) );
  MUX2_X1 npu_inst_pe_1_7_0_U158 ( .A(npu_inst_pe_1_7_0_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_7_0_int_q_reg_v_5__0_), .S(npu_inst_pe_1_7_0_n4), .Z(
        npu_inst_pe_1_7_0_n29) );
  MUX2_X1 npu_inst_pe_1_7_0_U157 ( .A(npu_inst_pe_1_7_0_n28), .B(
        npu_inst_pe_1_7_0_n23), .S(npu_inst_pe_1_7_0_n8), .Z(
        npu_inst_pe_1_7_0_N94) );
  MUX2_X1 npu_inst_pe_1_7_0_U156 ( .A(npu_inst_pe_1_7_0_n25), .B(
        npu_inst_pe_1_7_0_n24), .S(npu_inst_pe_1_7_0_n6), .Z(
        npu_inst_pe_1_7_0_n28) );
  MUX2_X1 npu_inst_pe_1_7_0_U155 ( .A(npu_inst_pe_1_7_0_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_7_0_int_q_reg_v_1__1_), .S(npu_inst_pe_1_7_0_n4), .Z(
        npu_inst_pe_1_7_0_n25) );
  MUX2_X1 npu_inst_pe_1_7_0_U154 ( .A(npu_inst_pe_1_7_0_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_7_0_int_q_reg_v_3__1_), .S(npu_inst_pe_1_7_0_n4), .Z(
        npu_inst_pe_1_7_0_n24) );
  MUX2_X1 npu_inst_pe_1_7_0_U153 ( .A(npu_inst_pe_1_7_0_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_7_0_int_q_reg_v_5__1_), .S(npu_inst_pe_1_7_0_n4), .Z(
        npu_inst_pe_1_7_0_n23) );
  MUX2_X1 npu_inst_pe_1_7_0_U152 ( .A(npu_inst_pe_1_7_0_n22), .B(
        npu_inst_pe_1_7_0_n19), .S(npu_inst_pe_1_7_0_n8), .Z(
        npu_inst_pe_1_7_0_o_data_h_1_) );
  MUX2_X1 npu_inst_pe_1_7_0_U151 ( .A(npu_inst_pe_1_7_0_n21), .B(
        npu_inst_pe_1_7_0_n20), .S(npu_inst_pe_1_7_0_n6), .Z(
        npu_inst_pe_1_7_0_n22) );
  MUX2_X1 npu_inst_pe_1_7_0_U150 ( .A(npu_inst_pe_1_7_0_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_7_0_int_q_reg_h_1__1_), .S(npu_inst_pe_1_7_0_n4), .Z(
        npu_inst_pe_1_7_0_n21) );
  MUX2_X1 npu_inst_pe_1_7_0_U149 ( .A(npu_inst_pe_1_7_0_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_7_0_int_q_reg_h_3__1_), .S(npu_inst_pe_1_7_0_n4), .Z(
        npu_inst_pe_1_7_0_n20) );
  MUX2_X1 npu_inst_pe_1_7_0_U148 ( .A(npu_inst_pe_1_7_0_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_7_0_int_q_reg_h_5__1_), .S(npu_inst_pe_1_7_0_n4), .Z(
        npu_inst_pe_1_7_0_n19) );
  MUX2_X1 npu_inst_pe_1_7_0_U147 ( .A(npu_inst_pe_1_7_0_n18), .B(
        npu_inst_pe_1_7_0_n15), .S(npu_inst_pe_1_7_0_n8), .Z(
        npu_inst_pe_1_7_0_o_data_h_0_) );
  MUX2_X1 npu_inst_pe_1_7_0_U146 ( .A(npu_inst_pe_1_7_0_n17), .B(
        npu_inst_pe_1_7_0_n16), .S(npu_inst_pe_1_7_0_n6), .Z(
        npu_inst_pe_1_7_0_n18) );
  MUX2_X1 npu_inst_pe_1_7_0_U145 ( .A(npu_inst_pe_1_7_0_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_7_0_int_q_reg_h_1__0_), .S(npu_inst_pe_1_7_0_n4), .Z(
        npu_inst_pe_1_7_0_n17) );
  MUX2_X1 npu_inst_pe_1_7_0_U144 ( .A(npu_inst_pe_1_7_0_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_7_0_int_q_reg_h_3__0_), .S(npu_inst_pe_1_7_0_n4), .Z(
        npu_inst_pe_1_7_0_n16) );
  MUX2_X1 npu_inst_pe_1_7_0_U143 ( .A(npu_inst_pe_1_7_0_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_7_0_int_q_reg_h_5__0_), .S(npu_inst_pe_1_7_0_n4), .Z(
        npu_inst_pe_1_7_0_n15) );
  XOR2_X1 npu_inst_pe_1_7_0_U142 ( .A(npu_inst_pe_1_7_0_int_data_0_), .B(
        npu_inst_pe_1_7_0_int_q_acc_0_), .Z(npu_inst_pe_1_7_0_N73) );
  AND2_X1 npu_inst_pe_1_7_0_U141 ( .A1(npu_inst_pe_1_7_0_int_q_acc_0_), .A2(
        npu_inst_pe_1_7_0_int_data_0_), .ZN(npu_inst_pe_1_7_0_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_7_0_U140 ( .A(npu_inst_pe_1_7_0_int_q_acc_0_), .B(
        npu_inst_pe_1_7_0_n13), .ZN(npu_inst_pe_1_7_0_N65) );
  OR2_X1 npu_inst_pe_1_7_0_U139 ( .A1(npu_inst_pe_1_7_0_n13), .A2(
        npu_inst_pe_1_7_0_int_q_acc_0_), .ZN(npu_inst_pe_1_7_0_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_7_0_U138 ( .A(npu_inst_pe_1_7_0_int_q_acc_2_), .B(
        npu_inst_pe_1_7_0_add_79_carry_2_), .Z(npu_inst_pe_1_7_0_N75) );
  AND2_X1 npu_inst_pe_1_7_0_U137 ( .A1(npu_inst_pe_1_7_0_add_79_carry_2_), 
        .A2(npu_inst_pe_1_7_0_int_q_acc_2_), .ZN(
        npu_inst_pe_1_7_0_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_7_0_U136 ( .A(npu_inst_pe_1_7_0_int_q_acc_3_), .B(
        npu_inst_pe_1_7_0_add_79_carry_3_), .Z(npu_inst_pe_1_7_0_N76) );
  AND2_X1 npu_inst_pe_1_7_0_U135 ( .A1(npu_inst_pe_1_7_0_add_79_carry_3_), 
        .A2(npu_inst_pe_1_7_0_int_q_acc_3_), .ZN(
        npu_inst_pe_1_7_0_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_7_0_U134 ( .A(npu_inst_pe_1_7_0_int_q_acc_4_), .B(
        npu_inst_pe_1_7_0_add_79_carry_4_), .Z(npu_inst_pe_1_7_0_N77) );
  AND2_X1 npu_inst_pe_1_7_0_U133 ( .A1(npu_inst_pe_1_7_0_add_79_carry_4_), 
        .A2(npu_inst_pe_1_7_0_int_q_acc_4_), .ZN(
        npu_inst_pe_1_7_0_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_7_0_U132 ( .A(npu_inst_pe_1_7_0_int_q_acc_5_), .B(
        npu_inst_pe_1_7_0_add_79_carry_5_), .Z(npu_inst_pe_1_7_0_N78) );
  AND2_X1 npu_inst_pe_1_7_0_U131 ( .A1(npu_inst_pe_1_7_0_add_79_carry_5_), 
        .A2(npu_inst_pe_1_7_0_int_q_acc_5_), .ZN(
        npu_inst_pe_1_7_0_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_7_0_U130 ( .A(npu_inst_pe_1_7_0_int_q_acc_6_), .B(
        npu_inst_pe_1_7_0_add_79_carry_6_), .Z(npu_inst_pe_1_7_0_N79) );
  AND2_X1 npu_inst_pe_1_7_0_U129 ( .A1(npu_inst_pe_1_7_0_add_79_carry_6_), 
        .A2(npu_inst_pe_1_7_0_int_q_acc_6_), .ZN(
        npu_inst_pe_1_7_0_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_7_0_U128 ( .A(npu_inst_pe_1_7_0_int_q_acc_7_), .B(
        npu_inst_pe_1_7_0_add_79_carry_7_), .Z(npu_inst_pe_1_7_0_N80) );
  XNOR2_X1 npu_inst_pe_1_7_0_U127 ( .A(npu_inst_pe_1_7_0_sub_77_carry_2_), .B(
        npu_inst_pe_1_7_0_int_q_acc_2_), .ZN(npu_inst_pe_1_7_0_N67) );
  OR2_X1 npu_inst_pe_1_7_0_U126 ( .A1(npu_inst_pe_1_7_0_int_q_acc_2_), .A2(
        npu_inst_pe_1_7_0_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_7_0_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_7_0_U125 ( .A(npu_inst_pe_1_7_0_sub_77_carry_3_), .B(
        npu_inst_pe_1_7_0_int_q_acc_3_), .ZN(npu_inst_pe_1_7_0_N68) );
  OR2_X1 npu_inst_pe_1_7_0_U124 ( .A1(npu_inst_pe_1_7_0_int_q_acc_3_), .A2(
        npu_inst_pe_1_7_0_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_7_0_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_7_0_U123 ( .A(npu_inst_pe_1_7_0_sub_77_carry_4_), .B(
        npu_inst_pe_1_7_0_int_q_acc_4_), .ZN(npu_inst_pe_1_7_0_N69) );
  OR2_X1 npu_inst_pe_1_7_0_U122 ( .A1(npu_inst_pe_1_7_0_int_q_acc_4_), .A2(
        npu_inst_pe_1_7_0_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_7_0_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_7_0_U121 ( .A(npu_inst_pe_1_7_0_sub_77_carry_5_), .B(
        npu_inst_pe_1_7_0_int_q_acc_5_), .ZN(npu_inst_pe_1_7_0_N70) );
  OR2_X1 npu_inst_pe_1_7_0_U120 ( .A1(npu_inst_pe_1_7_0_int_q_acc_5_), .A2(
        npu_inst_pe_1_7_0_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_7_0_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_7_0_U119 ( .A(npu_inst_pe_1_7_0_sub_77_carry_6_), .B(
        npu_inst_pe_1_7_0_int_q_acc_6_), .ZN(npu_inst_pe_1_7_0_N71) );
  OR2_X1 npu_inst_pe_1_7_0_U118 ( .A1(npu_inst_pe_1_7_0_int_q_acc_6_), .A2(
        npu_inst_pe_1_7_0_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_7_0_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_7_0_U117 ( .A(npu_inst_pe_1_7_0_int_q_acc_7_), .B(
        npu_inst_pe_1_7_0_sub_77_carry_7_), .ZN(npu_inst_pe_1_7_0_N72) );
  INV_X1 npu_inst_pe_1_7_0_U116 ( .A(npu_inst_n75), .ZN(npu_inst_pe_1_7_0_n7)
         );
  INV_X1 npu_inst_pe_1_7_0_U115 ( .A(npu_inst_pe_1_7_0_n7), .ZN(
        npu_inst_pe_1_7_0_n6) );
  INV_X1 npu_inst_pe_1_7_0_U114 ( .A(npu_inst_n53), .ZN(npu_inst_pe_1_7_0_n3)
         );
  AOI22_X1 npu_inst_pe_1_7_0_U113 ( .A1(npu_inst_pe_1_7_0_n38), .A2(
        int_i_data_v_npu[15]), .B1(npu_inst_pe_1_7_0_n118), .B2(
        npu_inst_pe_1_7_0_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_7_0_n39) );
  INV_X1 npu_inst_pe_1_7_0_U112 ( .A(npu_inst_pe_1_7_0_n39), .ZN(
        npu_inst_pe_1_7_0_n112) );
  AOI22_X1 npu_inst_pe_1_7_0_U111 ( .A1(npu_inst_pe_1_7_0_n38), .A2(
        int_i_data_v_npu[14]), .B1(npu_inst_pe_1_7_0_n118), .B2(
        npu_inst_pe_1_7_0_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_7_0_n37) );
  INV_X1 npu_inst_pe_1_7_0_U110 ( .A(npu_inst_pe_1_7_0_n37), .ZN(
        npu_inst_pe_1_7_0_n113) );
  AOI22_X1 npu_inst_pe_1_7_0_U107 ( .A1(int_i_data_v_npu[15]), .A2(
        npu_inst_pe_1_7_0_n58), .B1(npu_inst_pe_1_7_0_n114), .B2(
        npu_inst_pe_1_7_0_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_7_0_n59) );
  INV_X1 npu_inst_pe_1_7_0_U106 ( .A(npu_inst_pe_1_7_0_n59), .ZN(
        npu_inst_pe_1_7_0_n102) );
  AOI22_X1 npu_inst_pe_1_7_0_U105 ( .A1(int_i_data_v_npu[14]), .A2(
        npu_inst_pe_1_7_0_n58), .B1(npu_inst_pe_1_7_0_n114), .B2(
        npu_inst_pe_1_7_0_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_7_0_n57) );
  INV_X1 npu_inst_pe_1_7_0_U104 ( .A(npu_inst_pe_1_7_0_n57), .ZN(
        npu_inst_pe_1_7_0_n103) );
  AOI22_X1 npu_inst_pe_1_7_0_U103 ( .A1(int_i_data_v_npu[15]), .A2(
        npu_inst_pe_1_7_0_n54), .B1(npu_inst_pe_1_7_0_n115), .B2(
        npu_inst_pe_1_7_0_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_7_0_n55) );
  INV_X1 npu_inst_pe_1_7_0_U102 ( .A(npu_inst_pe_1_7_0_n55), .ZN(
        npu_inst_pe_1_7_0_n104) );
  AOI22_X1 npu_inst_pe_1_7_0_U101 ( .A1(int_i_data_v_npu[14]), .A2(
        npu_inst_pe_1_7_0_n54), .B1(npu_inst_pe_1_7_0_n115), .B2(
        npu_inst_pe_1_7_0_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_7_0_n53) );
  INV_X1 npu_inst_pe_1_7_0_U100 ( .A(npu_inst_pe_1_7_0_n53), .ZN(
        npu_inst_pe_1_7_0_n105) );
  AOI22_X1 npu_inst_pe_1_7_0_U99 ( .A1(int_i_data_v_npu[15]), .A2(
        npu_inst_pe_1_7_0_n50), .B1(npu_inst_pe_1_7_0_n116), .B2(
        npu_inst_pe_1_7_0_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_7_0_n51) );
  INV_X1 npu_inst_pe_1_7_0_U98 ( .A(npu_inst_pe_1_7_0_n51), .ZN(
        npu_inst_pe_1_7_0_n106) );
  AOI22_X1 npu_inst_pe_1_7_0_U97 ( .A1(int_i_data_v_npu[14]), .A2(
        npu_inst_pe_1_7_0_n50), .B1(npu_inst_pe_1_7_0_n116), .B2(
        npu_inst_pe_1_7_0_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_7_0_n49) );
  INV_X1 npu_inst_pe_1_7_0_U96 ( .A(npu_inst_pe_1_7_0_n49), .ZN(
        npu_inst_pe_1_7_0_n107) );
  AOI22_X1 npu_inst_pe_1_7_0_U95 ( .A1(int_i_data_v_npu[15]), .A2(
        npu_inst_pe_1_7_0_n46), .B1(npu_inst_pe_1_7_0_n117), .B2(
        npu_inst_pe_1_7_0_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_7_0_n47) );
  INV_X1 npu_inst_pe_1_7_0_U94 ( .A(npu_inst_pe_1_7_0_n47), .ZN(
        npu_inst_pe_1_7_0_n108) );
  AOI22_X1 npu_inst_pe_1_7_0_U93 ( .A1(int_i_data_v_npu[14]), .A2(
        npu_inst_pe_1_7_0_n46), .B1(npu_inst_pe_1_7_0_n117), .B2(
        npu_inst_pe_1_7_0_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_7_0_n45) );
  INV_X1 npu_inst_pe_1_7_0_U92 ( .A(npu_inst_pe_1_7_0_n45), .ZN(
        npu_inst_pe_1_7_0_n109) );
  AOI22_X1 npu_inst_pe_1_7_0_U91 ( .A1(int_i_data_v_npu[15]), .A2(
        npu_inst_pe_1_7_0_n42), .B1(npu_inst_pe_1_7_0_n119), .B2(
        npu_inst_pe_1_7_0_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_7_0_n43) );
  INV_X1 npu_inst_pe_1_7_0_U90 ( .A(npu_inst_pe_1_7_0_n43), .ZN(
        npu_inst_pe_1_7_0_n110) );
  AOI22_X1 npu_inst_pe_1_7_0_U89 ( .A1(int_i_data_v_npu[14]), .A2(
        npu_inst_pe_1_7_0_n42), .B1(npu_inst_pe_1_7_0_n119), .B2(
        npu_inst_pe_1_7_0_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_7_0_n41) );
  INV_X1 npu_inst_pe_1_7_0_U88 ( .A(npu_inst_pe_1_7_0_n41), .ZN(
        npu_inst_pe_1_7_0_n111) );
  NAND2_X1 npu_inst_pe_1_7_0_U87 ( .A1(npu_inst_pe_1_7_0_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_7_0_n60), .ZN(npu_inst_pe_1_7_0_n74) );
  OAI21_X1 npu_inst_pe_1_7_0_U86 ( .B1(npu_inst_pe_1_7_0_n63), .B2(
        npu_inst_pe_1_7_0_n60), .A(npu_inst_pe_1_7_0_n74), .ZN(
        npu_inst_pe_1_7_0_n97) );
  NAND2_X1 npu_inst_pe_1_7_0_U85 ( .A1(npu_inst_pe_1_7_0_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_7_0_n60), .ZN(npu_inst_pe_1_7_0_n73) );
  OAI21_X1 npu_inst_pe_1_7_0_U84 ( .B1(npu_inst_pe_1_7_0_n61), .B2(
        npu_inst_pe_1_7_0_n60), .A(npu_inst_pe_1_7_0_n73), .ZN(
        npu_inst_pe_1_7_0_n96) );
  NAND2_X1 npu_inst_pe_1_7_0_U83 ( .A1(npu_inst_pe_1_7_0_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_7_0_n56), .ZN(npu_inst_pe_1_7_0_n72) );
  OAI21_X1 npu_inst_pe_1_7_0_U82 ( .B1(npu_inst_pe_1_7_0_n63), .B2(
        npu_inst_pe_1_7_0_n56), .A(npu_inst_pe_1_7_0_n72), .ZN(
        npu_inst_pe_1_7_0_n95) );
  NAND2_X1 npu_inst_pe_1_7_0_U81 ( .A1(npu_inst_pe_1_7_0_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_7_0_n56), .ZN(npu_inst_pe_1_7_0_n71) );
  OAI21_X1 npu_inst_pe_1_7_0_U80 ( .B1(npu_inst_pe_1_7_0_n61), .B2(
        npu_inst_pe_1_7_0_n56), .A(npu_inst_pe_1_7_0_n71), .ZN(
        npu_inst_pe_1_7_0_n94) );
  NAND2_X1 npu_inst_pe_1_7_0_U79 ( .A1(npu_inst_pe_1_7_0_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_7_0_n52), .ZN(npu_inst_pe_1_7_0_n70) );
  OAI21_X1 npu_inst_pe_1_7_0_U78 ( .B1(npu_inst_pe_1_7_0_n63), .B2(
        npu_inst_pe_1_7_0_n52), .A(npu_inst_pe_1_7_0_n70), .ZN(
        npu_inst_pe_1_7_0_n93) );
  NAND2_X1 npu_inst_pe_1_7_0_U77 ( .A1(npu_inst_pe_1_7_0_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_7_0_n52), .ZN(npu_inst_pe_1_7_0_n69) );
  OAI21_X1 npu_inst_pe_1_7_0_U76 ( .B1(npu_inst_pe_1_7_0_n61), .B2(
        npu_inst_pe_1_7_0_n52), .A(npu_inst_pe_1_7_0_n69), .ZN(
        npu_inst_pe_1_7_0_n92) );
  NAND2_X1 npu_inst_pe_1_7_0_U75 ( .A1(npu_inst_pe_1_7_0_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_7_0_n48), .ZN(npu_inst_pe_1_7_0_n68) );
  OAI21_X1 npu_inst_pe_1_7_0_U74 ( .B1(npu_inst_pe_1_7_0_n63), .B2(
        npu_inst_pe_1_7_0_n48), .A(npu_inst_pe_1_7_0_n68), .ZN(
        npu_inst_pe_1_7_0_n91) );
  NAND2_X1 npu_inst_pe_1_7_0_U73 ( .A1(npu_inst_pe_1_7_0_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_7_0_n48), .ZN(npu_inst_pe_1_7_0_n67) );
  OAI21_X1 npu_inst_pe_1_7_0_U72 ( .B1(npu_inst_pe_1_7_0_n61), .B2(
        npu_inst_pe_1_7_0_n48), .A(npu_inst_pe_1_7_0_n67), .ZN(
        npu_inst_pe_1_7_0_n90) );
  NAND2_X1 npu_inst_pe_1_7_0_U71 ( .A1(npu_inst_pe_1_7_0_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_7_0_n44), .ZN(npu_inst_pe_1_7_0_n66) );
  OAI21_X1 npu_inst_pe_1_7_0_U70 ( .B1(npu_inst_pe_1_7_0_n63), .B2(
        npu_inst_pe_1_7_0_n44), .A(npu_inst_pe_1_7_0_n66), .ZN(
        npu_inst_pe_1_7_0_n89) );
  NAND2_X1 npu_inst_pe_1_7_0_U69 ( .A1(npu_inst_pe_1_7_0_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_7_0_n44), .ZN(npu_inst_pe_1_7_0_n65) );
  OAI21_X1 npu_inst_pe_1_7_0_U68 ( .B1(npu_inst_pe_1_7_0_n61), .B2(
        npu_inst_pe_1_7_0_n44), .A(npu_inst_pe_1_7_0_n65), .ZN(
        npu_inst_pe_1_7_0_n88) );
  NAND2_X1 npu_inst_pe_1_7_0_U67 ( .A1(npu_inst_pe_1_7_0_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_7_0_n40), .ZN(npu_inst_pe_1_7_0_n64) );
  OAI21_X1 npu_inst_pe_1_7_0_U66 ( .B1(npu_inst_pe_1_7_0_n63), .B2(
        npu_inst_pe_1_7_0_n40), .A(npu_inst_pe_1_7_0_n64), .ZN(
        npu_inst_pe_1_7_0_n87) );
  NAND2_X1 npu_inst_pe_1_7_0_U65 ( .A1(npu_inst_pe_1_7_0_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_7_0_n40), .ZN(npu_inst_pe_1_7_0_n62) );
  OAI21_X1 npu_inst_pe_1_7_0_U64 ( .B1(npu_inst_pe_1_7_0_n61), .B2(
        npu_inst_pe_1_7_0_n40), .A(npu_inst_pe_1_7_0_n62), .ZN(
        npu_inst_pe_1_7_0_n86) );
  AND2_X1 npu_inst_pe_1_7_0_U63 ( .A1(npu_inst_pe_1_7_0_N93), .A2(npu_inst_n53), .ZN(npu_inst_int_data_y_7__0__0_) );
  AND2_X1 npu_inst_pe_1_7_0_U62 ( .A1(npu_inst_n53), .A2(npu_inst_pe_1_7_0_N94), .ZN(npu_inst_int_data_y_7__0__1_) );
  AOI22_X1 npu_inst_pe_1_7_0_U61 ( .A1(npu_inst_n53), .A2(int_i_data_v_npu[15]), .B1(npu_inst_pe_1_7_0_n3), .B2(npu_inst_int_data_x_7__1__1_), .ZN(
        npu_inst_pe_1_7_0_n63) );
  AOI22_X1 npu_inst_pe_1_7_0_U60 ( .A1(npu_inst_n53), .A2(int_i_data_v_npu[14]), .B1(npu_inst_pe_1_7_0_n3), .B2(npu_inst_int_data_x_7__1__0_), .ZN(
        npu_inst_pe_1_7_0_n61) );
  NOR3_X1 npu_inst_pe_1_7_0_U59 ( .A1(npu_inst_pe_1_7_0_n26), .A2(npu_inst_n53), .A3(npu_inst_int_ckg[7]), .ZN(npu_inst_pe_1_7_0_n85) );
  OR2_X1 npu_inst_pe_1_7_0_U58 ( .A1(npu_inst_pe_1_7_0_n85), .A2(
        npu_inst_pe_1_7_0_n2), .ZN(npu_inst_pe_1_7_0_N84) );
  AOI222_X1 npu_inst_pe_1_7_0_U57 ( .A1(1'b0), .A2(npu_inst_pe_1_7_0_n1), .B1(
        npu_inst_pe_1_7_0_N73), .B2(npu_inst_pe_1_7_0_n76), .C1(
        npu_inst_pe_1_7_0_N65), .C2(npu_inst_pe_1_7_0_n77), .ZN(
        npu_inst_pe_1_7_0_n84) );
  INV_X1 npu_inst_pe_1_7_0_U56 ( .A(npu_inst_pe_1_7_0_n84), .ZN(
        npu_inst_pe_1_7_0_n101) );
  AOI222_X1 npu_inst_pe_1_7_0_U55 ( .A1(1'b0), .A2(npu_inst_pe_1_7_0_n1), .B1(
        npu_inst_pe_1_7_0_N80), .B2(npu_inst_pe_1_7_0_n76), .C1(
        npu_inst_pe_1_7_0_N72), .C2(npu_inst_pe_1_7_0_n77), .ZN(
        npu_inst_pe_1_7_0_n75) );
  INV_X1 npu_inst_pe_1_7_0_U54 ( .A(npu_inst_pe_1_7_0_n75), .ZN(
        npu_inst_pe_1_7_0_n33) );
  AOI222_X1 npu_inst_pe_1_7_0_U53 ( .A1(1'b0), .A2(npu_inst_pe_1_7_0_n1), .B1(
        npu_inst_pe_1_7_0_N74), .B2(npu_inst_pe_1_7_0_n76), .C1(
        npu_inst_pe_1_7_0_N66), .C2(npu_inst_pe_1_7_0_n77), .ZN(
        npu_inst_pe_1_7_0_n83) );
  INV_X1 npu_inst_pe_1_7_0_U52 ( .A(npu_inst_pe_1_7_0_n83), .ZN(
        npu_inst_pe_1_7_0_n100) );
  AOI222_X1 npu_inst_pe_1_7_0_U51 ( .A1(1'b0), .A2(npu_inst_pe_1_7_0_n1), .B1(
        npu_inst_pe_1_7_0_N75), .B2(npu_inst_pe_1_7_0_n76), .C1(
        npu_inst_pe_1_7_0_N67), .C2(npu_inst_pe_1_7_0_n77), .ZN(
        npu_inst_pe_1_7_0_n82) );
  INV_X1 npu_inst_pe_1_7_0_U50 ( .A(npu_inst_pe_1_7_0_n82), .ZN(
        npu_inst_pe_1_7_0_n99) );
  AOI222_X1 npu_inst_pe_1_7_0_U49 ( .A1(1'b0), .A2(npu_inst_pe_1_7_0_n1), .B1(
        npu_inst_pe_1_7_0_N76), .B2(npu_inst_pe_1_7_0_n76), .C1(
        npu_inst_pe_1_7_0_N68), .C2(npu_inst_pe_1_7_0_n77), .ZN(
        npu_inst_pe_1_7_0_n81) );
  INV_X1 npu_inst_pe_1_7_0_U48 ( .A(npu_inst_pe_1_7_0_n81), .ZN(
        npu_inst_pe_1_7_0_n98) );
  AOI222_X1 npu_inst_pe_1_7_0_U47 ( .A1(1'b0), .A2(npu_inst_pe_1_7_0_n1), .B1(
        npu_inst_pe_1_7_0_N77), .B2(npu_inst_pe_1_7_0_n76), .C1(
        npu_inst_pe_1_7_0_N69), .C2(npu_inst_pe_1_7_0_n77), .ZN(
        npu_inst_pe_1_7_0_n80) );
  INV_X1 npu_inst_pe_1_7_0_U46 ( .A(npu_inst_pe_1_7_0_n80), .ZN(
        npu_inst_pe_1_7_0_n36) );
  AOI222_X1 npu_inst_pe_1_7_0_U45 ( .A1(1'b0), .A2(npu_inst_pe_1_7_0_n1), .B1(
        npu_inst_pe_1_7_0_N78), .B2(npu_inst_pe_1_7_0_n76), .C1(
        npu_inst_pe_1_7_0_N70), .C2(npu_inst_pe_1_7_0_n77), .ZN(
        npu_inst_pe_1_7_0_n79) );
  INV_X1 npu_inst_pe_1_7_0_U44 ( .A(npu_inst_pe_1_7_0_n79), .ZN(
        npu_inst_pe_1_7_0_n35) );
  AOI222_X1 npu_inst_pe_1_7_0_U43 ( .A1(1'b0), .A2(npu_inst_pe_1_7_0_n1), .B1(
        npu_inst_pe_1_7_0_N79), .B2(npu_inst_pe_1_7_0_n76), .C1(
        npu_inst_pe_1_7_0_N71), .C2(npu_inst_pe_1_7_0_n77), .ZN(
        npu_inst_pe_1_7_0_n78) );
  INV_X1 npu_inst_pe_1_7_0_U42 ( .A(npu_inst_pe_1_7_0_n78), .ZN(
        npu_inst_pe_1_7_0_n34) );
  AND2_X1 npu_inst_pe_1_7_0_U41 ( .A1(npu_inst_pe_1_7_0_int_q_acc_0_), .A2(
        npu_inst_pe_1_7_0_n1), .ZN(npu_inst_int_data_res_7__0__0_) );
  AND2_X1 npu_inst_pe_1_7_0_U40 ( .A1(npu_inst_pe_1_7_0_n2), .A2(
        npu_inst_pe_1_7_0_int_q_acc_7_), .ZN(npu_inst_int_data_res_7__0__7_)
         );
  AND2_X1 npu_inst_pe_1_7_0_U39 ( .A1(npu_inst_pe_1_7_0_int_q_acc_1_), .A2(
        npu_inst_pe_1_7_0_n1), .ZN(npu_inst_int_data_res_7__0__1_) );
  AND2_X1 npu_inst_pe_1_7_0_U38 ( .A1(npu_inst_pe_1_7_0_int_q_acc_2_), .A2(
        npu_inst_pe_1_7_0_n1), .ZN(npu_inst_int_data_res_7__0__2_) );
  AND2_X1 npu_inst_pe_1_7_0_U37 ( .A1(npu_inst_pe_1_7_0_int_q_acc_3_), .A2(
        npu_inst_pe_1_7_0_n2), .ZN(npu_inst_int_data_res_7__0__3_) );
  AND2_X1 npu_inst_pe_1_7_0_U36 ( .A1(npu_inst_pe_1_7_0_int_q_acc_4_), .A2(
        npu_inst_pe_1_7_0_n2), .ZN(npu_inst_int_data_res_7__0__4_) );
  AND2_X1 npu_inst_pe_1_7_0_U35 ( .A1(npu_inst_pe_1_7_0_int_q_acc_5_), .A2(
        npu_inst_pe_1_7_0_n2), .ZN(npu_inst_int_data_res_7__0__5_) );
  AND2_X1 npu_inst_pe_1_7_0_U34 ( .A1(npu_inst_pe_1_7_0_int_q_acc_6_), .A2(
        npu_inst_pe_1_7_0_n2), .ZN(npu_inst_int_data_res_7__0__6_) );
  INV_X1 npu_inst_pe_1_7_0_U33 ( .A(npu_inst_pe_1_7_0_int_data_1_), .ZN(
        npu_inst_pe_1_7_0_n14) );
  AND2_X1 npu_inst_pe_1_7_0_U32 ( .A1(npu_inst_pe_1_7_0_o_data_h_1_), .A2(
        npu_inst_pe_1_7_0_int_q_weight_1_), .ZN(npu_inst_pe_1_7_0_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_7_0_U31 ( .A1(npu_inst_pe_1_7_0_o_data_h_0_), .A2(
        npu_inst_pe_1_7_0_int_q_weight_1_), .ZN(npu_inst_pe_1_7_0_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_7_0_U30 ( .A(npu_inst_pe_1_7_0_int_data_0_), .ZN(
        npu_inst_pe_1_7_0_n13) );
  INV_X1 npu_inst_pe_1_7_0_U29 ( .A(npu_inst_n67), .ZN(npu_inst_pe_1_7_0_n5)
         );
  OR3_X1 npu_inst_pe_1_7_0_U28 ( .A1(npu_inst_pe_1_7_0_n6), .A2(
        npu_inst_pe_1_7_0_n8), .A3(npu_inst_pe_1_7_0_n5), .ZN(
        npu_inst_pe_1_7_0_n56) );
  OR3_X1 npu_inst_pe_1_7_0_U27 ( .A1(npu_inst_pe_1_7_0_n5), .A2(
        npu_inst_pe_1_7_0_n8), .A3(npu_inst_pe_1_7_0_n7), .ZN(
        npu_inst_pe_1_7_0_n48) );
  INV_X1 npu_inst_pe_1_7_0_U26 ( .A(npu_inst_pe_1_7_0_n5), .ZN(
        npu_inst_pe_1_7_0_n4) );
  INV_X1 npu_inst_pe_1_7_0_U25 ( .A(npu_inst_n122), .ZN(npu_inst_pe_1_7_0_n12)
         );
  OR3_X1 npu_inst_pe_1_7_0_U24 ( .A1(npu_inst_pe_1_7_0_n4), .A2(
        npu_inst_pe_1_7_0_n8), .A3(npu_inst_pe_1_7_0_n7), .ZN(
        npu_inst_pe_1_7_0_n52) );
  OR3_X1 npu_inst_pe_1_7_0_U23 ( .A1(npu_inst_pe_1_7_0_n6), .A2(
        npu_inst_pe_1_7_0_n8), .A3(npu_inst_pe_1_7_0_n4), .ZN(
        npu_inst_pe_1_7_0_n60) );
  NOR2_X1 npu_inst_pe_1_7_0_U22 ( .A1(npu_inst_pe_1_7_0_n60), .A2(
        npu_inst_pe_1_7_0_n3), .ZN(npu_inst_pe_1_7_0_n58) );
  NOR2_X1 npu_inst_pe_1_7_0_U21 ( .A1(npu_inst_pe_1_7_0_n56), .A2(
        npu_inst_pe_1_7_0_n3), .ZN(npu_inst_pe_1_7_0_n54) );
  NOR2_X1 npu_inst_pe_1_7_0_U20 ( .A1(npu_inst_pe_1_7_0_n52), .A2(
        npu_inst_pe_1_7_0_n3), .ZN(npu_inst_pe_1_7_0_n50) );
  NOR2_X1 npu_inst_pe_1_7_0_U19 ( .A1(npu_inst_pe_1_7_0_n48), .A2(
        npu_inst_pe_1_7_0_n3), .ZN(npu_inst_pe_1_7_0_n46) );
  NOR2_X1 npu_inst_pe_1_7_0_U18 ( .A1(npu_inst_pe_1_7_0_n40), .A2(
        npu_inst_pe_1_7_0_n3), .ZN(npu_inst_pe_1_7_0_n38) );
  NOR2_X1 npu_inst_pe_1_7_0_U17 ( .A1(npu_inst_pe_1_7_0_n44), .A2(
        npu_inst_pe_1_7_0_n3), .ZN(npu_inst_pe_1_7_0_n42) );
  BUF_X1 npu_inst_pe_1_7_0_U16 ( .A(npu_inst_n93), .Z(npu_inst_pe_1_7_0_n8) );
  BUF_X1 npu_inst_pe_1_7_0_U15 ( .A(npu_inst_pe_1_7_0_n12), .Z(
        npu_inst_pe_1_7_0_n11) );
  BUF_X1 npu_inst_pe_1_7_0_U14 ( .A(npu_inst_pe_1_7_0_n12), .Z(
        npu_inst_pe_1_7_0_n10) );
  BUF_X1 npu_inst_pe_1_7_0_U13 ( .A(npu_inst_pe_1_7_0_n12), .Z(
        npu_inst_pe_1_7_0_n9) );
  INV_X1 npu_inst_pe_1_7_0_U12 ( .A(npu_inst_pe_1_7_0_n38), .ZN(
        npu_inst_pe_1_7_0_n118) );
  INV_X1 npu_inst_pe_1_7_0_U11 ( .A(npu_inst_pe_1_7_0_n58), .ZN(
        npu_inst_pe_1_7_0_n114) );
  INV_X1 npu_inst_pe_1_7_0_U10 ( .A(npu_inst_pe_1_7_0_n54), .ZN(
        npu_inst_pe_1_7_0_n115) );
  INV_X1 npu_inst_pe_1_7_0_U9 ( .A(npu_inst_pe_1_7_0_n50), .ZN(
        npu_inst_pe_1_7_0_n116) );
  INV_X1 npu_inst_pe_1_7_0_U8 ( .A(npu_inst_pe_1_7_0_n46), .ZN(
        npu_inst_pe_1_7_0_n117) );
  INV_X1 npu_inst_pe_1_7_0_U7 ( .A(npu_inst_pe_1_7_0_n42), .ZN(
        npu_inst_pe_1_7_0_n119) );
  BUF_X1 npu_inst_pe_1_7_0_U6 ( .A(npu_inst_n10), .Z(npu_inst_pe_1_7_0_n2) );
  BUF_X1 npu_inst_pe_1_7_0_U5 ( .A(npu_inst_n10), .Z(npu_inst_pe_1_7_0_n1) );
  NOR2_X1 npu_inst_pe_1_7_0_U4 ( .A1(npu_inst_pe_1_7_0_int_q_weight_0_), .A2(
        npu_inst_pe_1_7_0_n1), .ZN(npu_inst_pe_1_7_0_n76) );
  NOR2_X1 npu_inst_pe_1_7_0_U3 ( .A1(npu_inst_pe_1_7_0_n27), .A2(
        npu_inst_pe_1_7_0_n1), .ZN(npu_inst_pe_1_7_0_n77) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_7_0_n111), 
        .CK(npu_inst_pe_1_7_0_net3011), .RN(npu_inst_pe_1_7_0_n12), .Q(
        npu_inst_pe_1_7_0_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_7_0_n110), 
        .CK(npu_inst_pe_1_7_0_net3011), .RN(npu_inst_pe_1_7_0_n12), .Q(
        npu_inst_pe_1_7_0_int_q_reg_v_4__1_) );
  FA_X1 npu_inst_pe_1_7_0_sub_77_U2_1 ( .A(npu_inst_pe_1_7_0_int_q_acc_1_), 
        .B(npu_inst_pe_1_7_0_n14), .CI(npu_inst_pe_1_7_0_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_7_0_sub_77_carry_2_), .S(npu_inst_pe_1_7_0_N66) );
  FA_X1 npu_inst_pe_1_7_0_add_79_U1_1 ( .A(npu_inst_pe_1_7_0_int_q_acc_1_), 
        .B(npu_inst_pe_1_7_0_int_data_1_), .CI(
        npu_inst_pe_1_7_0_add_79_carry_1_), .CO(
        npu_inst_pe_1_7_0_add_79_carry_2_), .S(npu_inst_pe_1_7_0_N74) );
  NAND3_X1 npu_inst_pe_1_7_0_U109 ( .A1(npu_inst_pe_1_7_0_n5), .A2(
        npu_inst_pe_1_7_0_n7), .A3(npu_inst_pe_1_7_0_n8), .ZN(
        npu_inst_pe_1_7_0_n44) );
  NAND3_X1 npu_inst_pe_1_7_0_U108 ( .A1(npu_inst_pe_1_7_0_n4), .A2(
        npu_inst_pe_1_7_0_n7), .A3(npu_inst_pe_1_7_0_n8), .ZN(
        npu_inst_pe_1_7_0_n40) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_7_0_n34), .CK(
        npu_inst_pe_1_7_0_net3005), .RN(npu_inst_pe_1_7_0_n9), .Q(
        npu_inst_pe_1_7_0_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_7_0_n35), .CK(
        npu_inst_pe_1_7_0_net3005), .RN(npu_inst_pe_1_7_0_n9), .Q(
        npu_inst_pe_1_7_0_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_7_0_n36), .CK(
        npu_inst_pe_1_7_0_net3005), .RN(npu_inst_pe_1_7_0_n9), .Q(
        npu_inst_pe_1_7_0_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_7_0_n98), .CK(
        npu_inst_pe_1_7_0_net3005), .RN(npu_inst_pe_1_7_0_n9), .Q(
        npu_inst_pe_1_7_0_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_7_0_n99), .CK(
        npu_inst_pe_1_7_0_net3005), .RN(npu_inst_pe_1_7_0_n9), .Q(
        npu_inst_pe_1_7_0_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_7_0_n100), 
        .CK(npu_inst_pe_1_7_0_net3005), .RN(npu_inst_pe_1_7_0_n9), .Q(
        npu_inst_pe_1_7_0_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_7_0_n33), .CK(
        npu_inst_pe_1_7_0_net3005), .RN(npu_inst_pe_1_7_0_n9), .Q(
        npu_inst_pe_1_7_0_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_7_0_n101), 
        .CK(npu_inst_pe_1_7_0_net3005), .RN(npu_inst_pe_1_7_0_n9), .Q(
        npu_inst_pe_1_7_0_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_weight_reg_0_ ( .D(npu_inst_n108), .CK(
        npu_inst_pe_1_7_0_net3011), .RN(npu_inst_pe_1_7_0_n9), .Q(
        npu_inst_pe_1_7_0_int_q_weight_0_), .QN(npu_inst_pe_1_7_0_n27) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_weight_reg_1_ ( .D(npu_inst_n114), .CK(
        npu_inst_pe_1_7_0_net3011), .RN(npu_inst_pe_1_7_0_n9), .Q(
        npu_inst_pe_1_7_0_int_q_weight_1_), .QN(npu_inst_pe_1_7_0_n26) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_7_0_n113), 
        .CK(npu_inst_pe_1_7_0_net3011), .RN(npu_inst_pe_1_7_0_n9), .Q(
        npu_inst_pe_1_7_0_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_7_0_n112), 
        .CK(npu_inst_pe_1_7_0_net3011), .RN(npu_inst_pe_1_7_0_n9), .Q(
        npu_inst_pe_1_7_0_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_7_0_n109), 
        .CK(npu_inst_pe_1_7_0_net3011), .RN(npu_inst_pe_1_7_0_n10), .Q(
        npu_inst_pe_1_7_0_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_7_0_n108), 
        .CK(npu_inst_pe_1_7_0_net3011), .RN(npu_inst_pe_1_7_0_n10), .Q(
        npu_inst_pe_1_7_0_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_7_0_n107), 
        .CK(npu_inst_pe_1_7_0_net3011), .RN(npu_inst_pe_1_7_0_n10), .Q(
        npu_inst_pe_1_7_0_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_7_0_n106), 
        .CK(npu_inst_pe_1_7_0_net3011), .RN(npu_inst_pe_1_7_0_n10), .Q(
        npu_inst_pe_1_7_0_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_7_0_n105), 
        .CK(npu_inst_pe_1_7_0_net3011), .RN(npu_inst_pe_1_7_0_n10), .Q(
        npu_inst_pe_1_7_0_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_7_0_n104), 
        .CK(npu_inst_pe_1_7_0_net3011), .RN(npu_inst_pe_1_7_0_n10), .Q(
        npu_inst_pe_1_7_0_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_7_0_n103), 
        .CK(npu_inst_pe_1_7_0_net3011), .RN(npu_inst_pe_1_7_0_n10), .Q(
        npu_inst_pe_1_7_0_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_7_0_n102), 
        .CK(npu_inst_pe_1_7_0_net3011), .RN(npu_inst_pe_1_7_0_n10), .Q(
        npu_inst_pe_1_7_0_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_7_0_n86), 
        .CK(npu_inst_pe_1_7_0_net3011), .RN(npu_inst_pe_1_7_0_n10), .Q(
        npu_inst_pe_1_7_0_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_7_0_n87), 
        .CK(npu_inst_pe_1_7_0_net3011), .RN(npu_inst_pe_1_7_0_n10), .Q(
        npu_inst_pe_1_7_0_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_7_0_n88), 
        .CK(npu_inst_pe_1_7_0_net3011), .RN(npu_inst_pe_1_7_0_n11), .Q(
        npu_inst_pe_1_7_0_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_7_0_n89), 
        .CK(npu_inst_pe_1_7_0_net3011), .RN(npu_inst_pe_1_7_0_n11), .Q(
        npu_inst_pe_1_7_0_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_7_0_n90), 
        .CK(npu_inst_pe_1_7_0_net3011), .RN(npu_inst_pe_1_7_0_n11), .Q(
        npu_inst_pe_1_7_0_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_7_0_n91), 
        .CK(npu_inst_pe_1_7_0_net3011), .RN(npu_inst_pe_1_7_0_n11), .Q(
        npu_inst_pe_1_7_0_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_7_0_n92), 
        .CK(npu_inst_pe_1_7_0_net3011), .RN(npu_inst_pe_1_7_0_n11), .Q(
        npu_inst_pe_1_7_0_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_7_0_n93), 
        .CK(npu_inst_pe_1_7_0_net3011), .RN(npu_inst_pe_1_7_0_n11), .Q(
        npu_inst_pe_1_7_0_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_7_0_n94), 
        .CK(npu_inst_pe_1_7_0_net3011), .RN(npu_inst_pe_1_7_0_n11), .Q(
        npu_inst_pe_1_7_0_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_7_0_n95), 
        .CK(npu_inst_pe_1_7_0_net3011), .RN(npu_inst_pe_1_7_0_n11), .Q(
        npu_inst_pe_1_7_0_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_7_0_n96), 
        .CK(npu_inst_pe_1_7_0_net3011), .RN(npu_inst_pe_1_7_0_n11), .Q(
        npu_inst_pe_1_7_0_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_7_0_n97), 
        .CK(npu_inst_pe_1_7_0_net3011), .RN(npu_inst_pe_1_7_0_n11), .Q(
        npu_inst_pe_1_7_0_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_7_0_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_7_0_N84), .SE(1'b0), .GCK(npu_inst_pe_1_7_0_net3005) );
  CLKGATETST_X1 npu_inst_pe_1_7_0_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n61), .SE(1'b0), .GCK(npu_inst_pe_1_7_0_net3011) );
  MUX2_X1 npu_inst_pe_1_7_1_U162 ( .A(npu_inst_pe_1_7_1_n32), .B(
        npu_inst_pe_1_7_1_n29), .S(npu_inst_pe_1_7_1_n8), .Z(
        npu_inst_pe_1_7_1_N93) );
  MUX2_X1 npu_inst_pe_1_7_1_U161 ( .A(npu_inst_pe_1_7_1_n31), .B(
        npu_inst_pe_1_7_1_n30), .S(npu_inst_pe_1_7_1_n6), .Z(
        npu_inst_pe_1_7_1_n32) );
  MUX2_X1 npu_inst_pe_1_7_1_U160 ( .A(npu_inst_pe_1_7_1_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_7_1_int_q_reg_v_1__0_), .S(npu_inst_pe_1_7_1_n4), .Z(
        npu_inst_pe_1_7_1_n31) );
  MUX2_X1 npu_inst_pe_1_7_1_U159 ( .A(npu_inst_pe_1_7_1_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_7_1_int_q_reg_v_3__0_), .S(npu_inst_pe_1_7_1_n4), .Z(
        npu_inst_pe_1_7_1_n30) );
  MUX2_X1 npu_inst_pe_1_7_1_U158 ( .A(npu_inst_pe_1_7_1_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_7_1_int_q_reg_v_5__0_), .S(npu_inst_pe_1_7_1_n4), .Z(
        npu_inst_pe_1_7_1_n29) );
  MUX2_X1 npu_inst_pe_1_7_1_U157 ( .A(npu_inst_pe_1_7_1_n28), .B(
        npu_inst_pe_1_7_1_n23), .S(npu_inst_pe_1_7_1_n8), .Z(
        npu_inst_pe_1_7_1_N94) );
  MUX2_X1 npu_inst_pe_1_7_1_U156 ( .A(npu_inst_pe_1_7_1_n25), .B(
        npu_inst_pe_1_7_1_n24), .S(npu_inst_pe_1_7_1_n6), .Z(
        npu_inst_pe_1_7_1_n28) );
  MUX2_X1 npu_inst_pe_1_7_1_U155 ( .A(npu_inst_pe_1_7_1_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_7_1_int_q_reg_v_1__1_), .S(npu_inst_pe_1_7_1_n4), .Z(
        npu_inst_pe_1_7_1_n25) );
  MUX2_X1 npu_inst_pe_1_7_1_U154 ( .A(npu_inst_pe_1_7_1_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_7_1_int_q_reg_v_3__1_), .S(npu_inst_pe_1_7_1_n4), .Z(
        npu_inst_pe_1_7_1_n24) );
  MUX2_X1 npu_inst_pe_1_7_1_U153 ( .A(npu_inst_pe_1_7_1_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_7_1_int_q_reg_v_5__1_), .S(npu_inst_pe_1_7_1_n4), .Z(
        npu_inst_pe_1_7_1_n23) );
  MUX2_X1 npu_inst_pe_1_7_1_U152 ( .A(npu_inst_pe_1_7_1_n22), .B(
        npu_inst_pe_1_7_1_n19), .S(npu_inst_pe_1_7_1_n8), .Z(
        npu_inst_int_data_x_7__1__1_) );
  MUX2_X1 npu_inst_pe_1_7_1_U151 ( .A(npu_inst_pe_1_7_1_n21), .B(
        npu_inst_pe_1_7_1_n20), .S(npu_inst_pe_1_7_1_n6), .Z(
        npu_inst_pe_1_7_1_n22) );
  MUX2_X1 npu_inst_pe_1_7_1_U150 ( .A(npu_inst_pe_1_7_1_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_7_1_int_q_reg_h_1__1_), .S(npu_inst_pe_1_7_1_n4), .Z(
        npu_inst_pe_1_7_1_n21) );
  MUX2_X1 npu_inst_pe_1_7_1_U149 ( .A(npu_inst_pe_1_7_1_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_7_1_int_q_reg_h_3__1_), .S(npu_inst_pe_1_7_1_n4), .Z(
        npu_inst_pe_1_7_1_n20) );
  MUX2_X1 npu_inst_pe_1_7_1_U148 ( .A(npu_inst_pe_1_7_1_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_7_1_int_q_reg_h_5__1_), .S(npu_inst_pe_1_7_1_n4), .Z(
        npu_inst_pe_1_7_1_n19) );
  MUX2_X1 npu_inst_pe_1_7_1_U147 ( .A(npu_inst_pe_1_7_1_n18), .B(
        npu_inst_pe_1_7_1_n15), .S(npu_inst_pe_1_7_1_n8), .Z(
        npu_inst_int_data_x_7__1__0_) );
  MUX2_X1 npu_inst_pe_1_7_1_U146 ( .A(npu_inst_pe_1_7_1_n17), .B(
        npu_inst_pe_1_7_1_n16), .S(npu_inst_pe_1_7_1_n6), .Z(
        npu_inst_pe_1_7_1_n18) );
  MUX2_X1 npu_inst_pe_1_7_1_U145 ( .A(npu_inst_pe_1_7_1_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_7_1_int_q_reg_h_1__0_), .S(npu_inst_pe_1_7_1_n4), .Z(
        npu_inst_pe_1_7_1_n17) );
  MUX2_X1 npu_inst_pe_1_7_1_U144 ( .A(npu_inst_pe_1_7_1_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_7_1_int_q_reg_h_3__0_), .S(npu_inst_pe_1_7_1_n4), .Z(
        npu_inst_pe_1_7_1_n16) );
  MUX2_X1 npu_inst_pe_1_7_1_U143 ( .A(npu_inst_pe_1_7_1_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_7_1_int_q_reg_h_5__0_), .S(npu_inst_pe_1_7_1_n4), .Z(
        npu_inst_pe_1_7_1_n15) );
  XOR2_X1 npu_inst_pe_1_7_1_U142 ( .A(npu_inst_pe_1_7_1_int_data_0_), .B(
        npu_inst_pe_1_7_1_int_q_acc_0_), .Z(npu_inst_pe_1_7_1_N73) );
  AND2_X1 npu_inst_pe_1_7_1_U141 ( .A1(npu_inst_pe_1_7_1_int_q_acc_0_), .A2(
        npu_inst_pe_1_7_1_int_data_0_), .ZN(npu_inst_pe_1_7_1_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_7_1_U140 ( .A(npu_inst_pe_1_7_1_int_q_acc_0_), .B(
        npu_inst_pe_1_7_1_n13), .ZN(npu_inst_pe_1_7_1_N65) );
  OR2_X1 npu_inst_pe_1_7_1_U139 ( .A1(npu_inst_pe_1_7_1_n13), .A2(
        npu_inst_pe_1_7_1_int_q_acc_0_), .ZN(npu_inst_pe_1_7_1_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_7_1_U138 ( .A(npu_inst_pe_1_7_1_int_q_acc_2_), .B(
        npu_inst_pe_1_7_1_add_79_carry_2_), .Z(npu_inst_pe_1_7_1_N75) );
  AND2_X1 npu_inst_pe_1_7_1_U137 ( .A1(npu_inst_pe_1_7_1_add_79_carry_2_), 
        .A2(npu_inst_pe_1_7_1_int_q_acc_2_), .ZN(
        npu_inst_pe_1_7_1_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_7_1_U136 ( .A(npu_inst_pe_1_7_1_int_q_acc_3_), .B(
        npu_inst_pe_1_7_1_add_79_carry_3_), .Z(npu_inst_pe_1_7_1_N76) );
  AND2_X1 npu_inst_pe_1_7_1_U135 ( .A1(npu_inst_pe_1_7_1_add_79_carry_3_), 
        .A2(npu_inst_pe_1_7_1_int_q_acc_3_), .ZN(
        npu_inst_pe_1_7_1_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_7_1_U134 ( .A(npu_inst_pe_1_7_1_int_q_acc_4_), .B(
        npu_inst_pe_1_7_1_add_79_carry_4_), .Z(npu_inst_pe_1_7_1_N77) );
  AND2_X1 npu_inst_pe_1_7_1_U133 ( .A1(npu_inst_pe_1_7_1_add_79_carry_4_), 
        .A2(npu_inst_pe_1_7_1_int_q_acc_4_), .ZN(
        npu_inst_pe_1_7_1_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_7_1_U132 ( .A(npu_inst_pe_1_7_1_int_q_acc_5_), .B(
        npu_inst_pe_1_7_1_add_79_carry_5_), .Z(npu_inst_pe_1_7_1_N78) );
  AND2_X1 npu_inst_pe_1_7_1_U131 ( .A1(npu_inst_pe_1_7_1_add_79_carry_5_), 
        .A2(npu_inst_pe_1_7_1_int_q_acc_5_), .ZN(
        npu_inst_pe_1_7_1_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_7_1_U130 ( .A(npu_inst_pe_1_7_1_int_q_acc_6_), .B(
        npu_inst_pe_1_7_1_add_79_carry_6_), .Z(npu_inst_pe_1_7_1_N79) );
  AND2_X1 npu_inst_pe_1_7_1_U129 ( .A1(npu_inst_pe_1_7_1_add_79_carry_6_), 
        .A2(npu_inst_pe_1_7_1_int_q_acc_6_), .ZN(
        npu_inst_pe_1_7_1_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_7_1_U128 ( .A(npu_inst_pe_1_7_1_int_q_acc_7_), .B(
        npu_inst_pe_1_7_1_add_79_carry_7_), .Z(npu_inst_pe_1_7_1_N80) );
  XNOR2_X1 npu_inst_pe_1_7_1_U127 ( .A(npu_inst_pe_1_7_1_sub_77_carry_2_), .B(
        npu_inst_pe_1_7_1_int_q_acc_2_), .ZN(npu_inst_pe_1_7_1_N67) );
  OR2_X1 npu_inst_pe_1_7_1_U126 ( .A1(npu_inst_pe_1_7_1_int_q_acc_2_), .A2(
        npu_inst_pe_1_7_1_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_7_1_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_7_1_U125 ( .A(npu_inst_pe_1_7_1_sub_77_carry_3_), .B(
        npu_inst_pe_1_7_1_int_q_acc_3_), .ZN(npu_inst_pe_1_7_1_N68) );
  OR2_X1 npu_inst_pe_1_7_1_U124 ( .A1(npu_inst_pe_1_7_1_int_q_acc_3_), .A2(
        npu_inst_pe_1_7_1_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_7_1_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_7_1_U123 ( .A(npu_inst_pe_1_7_1_sub_77_carry_4_), .B(
        npu_inst_pe_1_7_1_int_q_acc_4_), .ZN(npu_inst_pe_1_7_1_N69) );
  OR2_X1 npu_inst_pe_1_7_1_U122 ( .A1(npu_inst_pe_1_7_1_int_q_acc_4_), .A2(
        npu_inst_pe_1_7_1_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_7_1_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_7_1_U121 ( .A(npu_inst_pe_1_7_1_sub_77_carry_5_), .B(
        npu_inst_pe_1_7_1_int_q_acc_5_), .ZN(npu_inst_pe_1_7_1_N70) );
  OR2_X1 npu_inst_pe_1_7_1_U120 ( .A1(npu_inst_pe_1_7_1_int_q_acc_5_), .A2(
        npu_inst_pe_1_7_1_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_7_1_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_7_1_U119 ( .A(npu_inst_pe_1_7_1_sub_77_carry_6_), .B(
        npu_inst_pe_1_7_1_int_q_acc_6_), .ZN(npu_inst_pe_1_7_1_N71) );
  OR2_X1 npu_inst_pe_1_7_1_U118 ( .A1(npu_inst_pe_1_7_1_int_q_acc_6_), .A2(
        npu_inst_pe_1_7_1_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_7_1_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_7_1_U117 ( .A(npu_inst_pe_1_7_1_int_q_acc_7_), .B(
        npu_inst_pe_1_7_1_sub_77_carry_7_), .ZN(npu_inst_pe_1_7_1_N72) );
  INV_X1 npu_inst_pe_1_7_1_U116 ( .A(npu_inst_n75), .ZN(npu_inst_pe_1_7_1_n7)
         );
  INV_X1 npu_inst_pe_1_7_1_U115 ( .A(npu_inst_pe_1_7_1_n7), .ZN(
        npu_inst_pe_1_7_1_n6) );
  INV_X1 npu_inst_pe_1_7_1_U114 ( .A(npu_inst_n52), .ZN(npu_inst_pe_1_7_1_n3)
         );
  AOI22_X1 npu_inst_pe_1_7_1_U113 ( .A1(npu_inst_pe_1_7_1_n38), .A2(
        int_i_data_v_npu[13]), .B1(npu_inst_pe_1_7_1_n118), .B2(
        npu_inst_pe_1_7_1_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_7_1_n39) );
  INV_X1 npu_inst_pe_1_7_1_U112 ( .A(npu_inst_pe_1_7_1_n39), .ZN(
        npu_inst_pe_1_7_1_n112) );
  AOI22_X1 npu_inst_pe_1_7_1_U111 ( .A1(npu_inst_pe_1_7_1_n38), .A2(
        int_i_data_v_npu[12]), .B1(npu_inst_pe_1_7_1_n118), .B2(
        npu_inst_pe_1_7_1_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_7_1_n37) );
  INV_X1 npu_inst_pe_1_7_1_U110 ( .A(npu_inst_pe_1_7_1_n37), .ZN(
        npu_inst_pe_1_7_1_n113) );
  AOI22_X1 npu_inst_pe_1_7_1_U107 ( .A1(int_i_data_v_npu[13]), .A2(
        npu_inst_pe_1_7_1_n58), .B1(npu_inst_pe_1_7_1_n114), .B2(
        npu_inst_pe_1_7_1_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_7_1_n59) );
  INV_X1 npu_inst_pe_1_7_1_U106 ( .A(npu_inst_pe_1_7_1_n59), .ZN(
        npu_inst_pe_1_7_1_n102) );
  AOI22_X1 npu_inst_pe_1_7_1_U105 ( .A1(int_i_data_v_npu[12]), .A2(
        npu_inst_pe_1_7_1_n58), .B1(npu_inst_pe_1_7_1_n114), .B2(
        npu_inst_pe_1_7_1_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_7_1_n57) );
  INV_X1 npu_inst_pe_1_7_1_U104 ( .A(npu_inst_pe_1_7_1_n57), .ZN(
        npu_inst_pe_1_7_1_n103) );
  AOI22_X1 npu_inst_pe_1_7_1_U103 ( .A1(int_i_data_v_npu[13]), .A2(
        npu_inst_pe_1_7_1_n54), .B1(npu_inst_pe_1_7_1_n115), .B2(
        npu_inst_pe_1_7_1_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_7_1_n55) );
  INV_X1 npu_inst_pe_1_7_1_U102 ( .A(npu_inst_pe_1_7_1_n55), .ZN(
        npu_inst_pe_1_7_1_n104) );
  AOI22_X1 npu_inst_pe_1_7_1_U101 ( .A1(int_i_data_v_npu[12]), .A2(
        npu_inst_pe_1_7_1_n54), .B1(npu_inst_pe_1_7_1_n115), .B2(
        npu_inst_pe_1_7_1_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_7_1_n53) );
  INV_X1 npu_inst_pe_1_7_1_U100 ( .A(npu_inst_pe_1_7_1_n53), .ZN(
        npu_inst_pe_1_7_1_n105) );
  AOI22_X1 npu_inst_pe_1_7_1_U99 ( .A1(int_i_data_v_npu[13]), .A2(
        npu_inst_pe_1_7_1_n50), .B1(npu_inst_pe_1_7_1_n116), .B2(
        npu_inst_pe_1_7_1_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_7_1_n51) );
  INV_X1 npu_inst_pe_1_7_1_U98 ( .A(npu_inst_pe_1_7_1_n51), .ZN(
        npu_inst_pe_1_7_1_n106) );
  AOI22_X1 npu_inst_pe_1_7_1_U97 ( .A1(int_i_data_v_npu[12]), .A2(
        npu_inst_pe_1_7_1_n50), .B1(npu_inst_pe_1_7_1_n116), .B2(
        npu_inst_pe_1_7_1_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_7_1_n49) );
  INV_X1 npu_inst_pe_1_7_1_U96 ( .A(npu_inst_pe_1_7_1_n49), .ZN(
        npu_inst_pe_1_7_1_n107) );
  AOI22_X1 npu_inst_pe_1_7_1_U95 ( .A1(int_i_data_v_npu[13]), .A2(
        npu_inst_pe_1_7_1_n46), .B1(npu_inst_pe_1_7_1_n117), .B2(
        npu_inst_pe_1_7_1_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_7_1_n47) );
  INV_X1 npu_inst_pe_1_7_1_U94 ( .A(npu_inst_pe_1_7_1_n47), .ZN(
        npu_inst_pe_1_7_1_n108) );
  AOI22_X1 npu_inst_pe_1_7_1_U93 ( .A1(int_i_data_v_npu[12]), .A2(
        npu_inst_pe_1_7_1_n46), .B1(npu_inst_pe_1_7_1_n117), .B2(
        npu_inst_pe_1_7_1_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_7_1_n45) );
  INV_X1 npu_inst_pe_1_7_1_U92 ( .A(npu_inst_pe_1_7_1_n45), .ZN(
        npu_inst_pe_1_7_1_n109) );
  AOI22_X1 npu_inst_pe_1_7_1_U91 ( .A1(int_i_data_v_npu[13]), .A2(
        npu_inst_pe_1_7_1_n42), .B1(npu_inst_pe_1_7_1_n119), .B2(
        npu_inst_pe_1_7_1_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_7_1_n43) );
  INV_X1 npu_inst_pe_1_7_1_U90 ( .A(npu_inst_pe_1_7_1_n43), .ZN(
        npu_inst_pe_1_7_1_n110) );
  AOI22_X1 npu_inst_pe_1_7_1_U89 ( .A1(int_i_data_v_npu[12]), .A2(
        npu_inst_pe_1_7_1_n42), .B1(npu_inst_pe_1_7_1_n119), .B2(
        npu_inst_pe_1_7_1_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_7_1_n41) );
  INV_X1 npu_inst_pe_1_7_1_U88 ( .A(npu_inst_pe_1_7_1_n41), .ZN(
        npu_inst_pe_1_7_1_n111) );
  NAND2_X1 npu_inst_pe_1_7_1_U87 ( .A1(npu_inst_pe_1_7_1_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_7_1_n60), .ZN(npu_inst_pe_1_7_1_n74) );
  OAI21_X1 npu_inst_pe_1_7_1_U86 ( .B1(npu_inst_pe_1_7_1_n63), .B2(
        npu_inst_pe_1_7_1_n60), .A(npu_inst_pe_1_7_1_n74), .ZN(
        npu_inst_pe_1_7_1_n97) );
  NAND2_X1 npu_inst_pe_1_7_1_U85 ( .A1(npu_inst_pe_1_7_1_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_7_1_n60), .ZN(npu_inst_pe_1_7_1_n73) );
  OAI21_X1 npu_inst_pe_1_7_1_U84 ( .B1(npu_inst_pe_1_7_1_n61), .B2(
        npu_inst_pe_1_7_1_n60), .A(npu_inst_pe_1_7_1_n73), .ZN(
        npu_inst_pe_1_7_1_n96) );
  NAND2_X1 npu_inst_pe_1_7_1_U83 ( .A1(npu_inst_pe_1_7_1_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_7_1_n56), .ZN(npu_inst_pe_1_7_1_n72) );
  OAI21_X1 npu_inst_pe_1_7_1_U82 ( .B1(npu_inst_pe_1_7_1_n63), .B2(
        npu_inst_pe_1_7_1_n56), .A(npu_inst_pe_1_7_1_n72), .ZN(
        npu_inst_pe_1_7_1_n95) );
  NAND2_X1 npu_inst_pe_1_7_1_U81 ( .A1(npu_inst_pe_1_7_1_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_7_1_n56), .ZN(npu_inst_pe_1_7_1_n71) );
  OAI21_X1 npu_inst_pe_1_7_1_U80 ( .B1(npu_inst_pe_1_7_1_n61), .B2(
        npu_inst_pe_1_7_1_n56), .A(npu_inst_pe_1_7_1_n71), .ZN(
        npu_inst_pe_1_7_1_n94) );
  NAND2_X1 npu_inst_pe_1_7_1_U79 ( .A1(npu_inst_pe_1_7_1_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_7_1_n52), .ZN(npu_inst_pe_1_7_1_n70) );
  OAI21_X1 npu_inst_pe_1_7_1_U78 ( .B1(npu_inst_pe_1_7_1_n63), .B2(
        npu_inst_pe_1_7_1_n52), .A(npu_inst_pe_1_7_1_n70), .ZN(
        npu_inst_pe_1_7_1_n93) );
  NAND2_X1 npu_inst_pe_1_7_1_U77 ( .A1(npu_inst_pe_1_7_1_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_7_1_n52), .ZN(npu_inst_pe_1_7_1_n69) );
  OAI21_X1 npu_inst_pe_1_7_1_U76 ( .B1(npu_inst_pe_1_7_1_n61), .B2(
        npu_inst_pe_1_7_1_n52), .A(npu_inst_pe_1_7_1_n69), .ZN(
        npu_inst_pe_1_7_1_n92) );
  NAND2_X1 npu_inst_pe_1_7_1_U75 ( .A1(npu_inst_pe_1_7_1_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_7_1_n48), .ZN(npu_inst_pe_1_7_1_n68) );
  OAI21_X1 npu_inst_pe_1_7_1_U74 ( .B1(npu_inst_pe_1_7_1_n63), .B2(
        npu_inst_pe_1_7_1_n48), .A(npu_inst_pe_1_7_1_n68), .ZN(
        npu_inst_pe_1_7_1_n91) );
  NAND2_X1 npu_inst_pe_1_7_1_U73 ( .A1(npu_inst_pe_1_7_1_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_7_1_n48), .ZN(npu_inst_pe_1_7_1_n67) );
  OAI21_X1 npu_inst_pe_1_7_1_U72 ( .B1(npu_inst_pe_1_7_1_n61), .B2(
        npu_inst_pe_1_7_1_n48), .A(npu_inst_pe_1_7_1_n67), .ZN(
        npu_inst_pe_1_7_1_n90) );
  NAND2_X1 npu_inst_pe_1_7_1_U71 ( .A1(npu_inst_pe_1_7_1_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_7_1_n44), .ZN(npu_inst_pe_1_7_1_n66) );
  OAI21_X1 npu_inst_pe_1_7_1_U70 ( .B1(npu_inst_pe_1_7_1_n63), .B2(
        npu_inst_pe_1_7_1_n44), .A(npu_inst_pe_1_7_1_n66), .ZN(
        npu_inst_pe_1_7_1_n89) );
  NAND2_X1 npu_inst_pe_1_7_1_U69 ( .A1(npu_inst_pe_1_7_1_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_7_1_n44), .ZN(npu_inst_pe_1_7_1_n65) );
  OAI21_X1 npu_inst_pe_1_7_1_U68 ( .B1(npu_inst_pe_1_7_1_n61), .B2(
        npu_inst_pe_1_7_1_n44), .A(npu_inst_pe_1_7_1_n65), .ZN(
        npu_inst_pe_1_7_1_n88) );
  NAND2_X1 npu_inst_pe_1_7_1_U67 ( .A1(npu_inst_pe_1_7_1_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_7_1_n40), .ZN(npu_inst_pe_1_7_1_n64) );
  OAI21_X1 npu_inst_pe_1_7_1_U66 ( .B1(npu_inst_pe_1_7_1_n63), .B2(
        npu_inst_pe_1_7_1_n40), .A(npu_inst_pe_1_7_1_n64), .ZN(
        npu_inst_pe_1_7_1_n87) );
  NAND2_X1 npu_inst_pe_1_7_1_U65 ( .A1(npu_inst_pe_1_7_1_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_7_1_n40), .ZN(npu_inst_pe_1_7_1_n62) );
  OAI21_X1 npu_inst_pe_1_7_1_U64 ( .B1(npu_inst_pe_1_7_1_n61), .B2(
        npu_inst_pe_1_7_1_n40), .A(npu_inst_pe_1_7_1_n62), .ZN(
        npu_inst_pe_1_7_1_n86) );
  AND2_X1 npu_inst_pe_1_7_1_U63 ( .A1(npu_inst_pe_1_7_1_N93), .A2(npu_inst_n52), .ZN(npu_inst_int_data_y_7__1__0_) );
  AND2_X1 npu_inst_pe_1_7_1_U62 ( .A1(npu_inst_n52), .A2(npu_inst_pe_1_7_1_N94), .ZN(npu_inst_int_data_y_7__1__1_) );
  AOI22_X1 npu_inst_pe_1_7_1_U61 ( .A1(npu_inst_n52), .A2(int_i_data_v_npu[13]), .B1(npu_inst_pe_1_7_1_n3), .B2(npu_inst_int_data_x_7__2__1_), .ZN(
        npu_inst_pe_1_7_1_n63) );
  AOI22_X1 npu_inst_pe_1_7_1_U60 ( .A1(npu_inst_n52), .A2(int_i_data_v_npu[12]), .B1(npu_inst_pe_1_7_1_n3), .B2(npu_inst_int_data_x_7__2__0_), .ZN(
        npu_inst_pe_1_7_1_n61) );
  NOR3_X1 npu_inst_pe_1_7_1_U59 ( .A1(npu_inst_pe_1_7_1_n26), .A2(npu_inst_n52), .A3(npu_inst_int_ckg[6]), .ZN(npu_inst_pe_1_7_1_n85) );
  OR2_X1 npu_inst_pe_1_7_1_U58 ( .A1(npu_inst_pe_1_7_1_n85), .A2(
        npu_inst_pe_1_7_1_n2), .ZN(npu_inst_pe_1_7_1_N84) );
  AOI222_X1 npu_inst_pe_1_7_1_U57 ( .A1(1'b0), .A2(npu_inst_pe_1_7_1_n1), .B1(
        npu_inst_pe_1_7_1_N73), .B2(npu_inst_pe_1_7_1_n76), .C1(
        npu_inst_pe_1_7_1_N65), .C2(npu_inst_pe_1_7_1_n77), .ZN(
        npu_inst_pe_1_7_1_n84) );
  INV_X1 npu_inst_pe_1_7_1_U56 ( .A(npu_inst_pe_1_7_1_n84), .ZN(
        npu_inst_pe_1_7_1_n101) );
  AOI222_X1 npu_inst_pe_1_7_1_U55 ( .A1(1'b0), .A2(npu_inst_pe_1_7_1_n1), .B1(
        npu_inst_pe_1_7_1_N80), .B2(npu_inst_pe_1_7_1_n76), .C1(
        npu_inst_pe_1_7_1_N72), .C2(npu_inst_pe_1_7_1_n77), .ZN(
        npu_inst_pe_1_7_1_n75) );
  INV_X1 npu_inst_pe_1_7_1_U54 ( .A(npu_inst_pe_1_7_1_n75), .ZN(
        npu_inst_pe_1_7_1_n33) );
  AOI222_X1 npu_inst_pe_1_7_1_U53 ( .A1(1'b0), .A2(npu_inst_pe_1_7_1_n1), .B1(
        npu_inst_pe_1_7_1_N74), .B2(npu_inst_pe_1_7_1_n76), .C1(
        npu_inst_pe_1_7_1_N66), .C2(npu_inst_pe_1_7_1_n77), .ZN(
        npu_inst_pe_1_7_1_n83) );
  INV_X1 npu_inst_pe_1_7_1_U52 ( .A(npu_inst_pe_1_7_1_n83), .ZN(
        npu_inst_pe_1_7_1_n100) );
  AOI222_X1 npu_inst_pe_1_7_1_U51 ( .A1(1'b0), .A2(npu_inst_pe_1_7_1_n1), .B1(
        npu_inst_pe_1_7_1_N75), .B2(npu_inst_pe_1_7_1_n76), .C1(
        npu_inst_pe_1_7_1_N67), .C2(npu_inst_pe_1_7_1_n77), .ZN(
        npu_inst_pe_1_7_1_n82) );
  INV_X1 npu_inst_pe_1_7_1_U50 ( .A(npu_inst_pe_1_7_1_n82), .ZN(
        npu_inst_pe_1_7_1_n99) );
  AOI222_X1 npu_inst_pe_1_7_1_U49 ( .A1(1'b0), .A2(npu_inst_pe_1_7_1_n1), .B1(
        npu_inst_pe_1_7_1_N76), .B2(npu_inst_pe_1_7_1_n76), .C1(
        npu_inst_pe_1_7_1_N68), .C2(npu_inst_pe_1_7_1_n77), .ZN(
        npu_inst_pe_1_7_1_n81) );
  INV_X1 npu_inst_pe_1_7_1_U48 ( .A(npu_inst_pe_1_7_1_n81), .ZN(
        npu_inst_pe_1_7_1_n98) );
  AOI222_X1 npu_inst_pe_1_7_1_U47 ( .A1(1'b0), .A2(npu_inst_pe_1_7_1_n1), .B1(
        npu_inst_pe_1_7_1_N77), .B2(npu_inst_pe_1_7_1_n76), .C1(
        npu_inst_pe_1_7_1_N69), .C2(npu_inst_pe_1_7_1_n77), .ZN(
        npu_inst_pe_1_7_1_n80) );
  INV_X1 npu_inst_pe_1_7_1_U46 ( .A(npu_inst_pe_1_7_1_n80), .ZN(
        npu_inst_pe_1_7_1_n36) );
  AOI222_X1 npu_inst_pe_1_7_1_U45 ( .A1(1'b0), .A2(npu_inst_pe_1_7_1_n1), .B1(
        npu_inst_pe_1_7_1_N78), .B2(npu_inst_pe_1_7_1_n76), .C1(
        npu_inst_pe_1_7_1_N70), .C2(npu_inst_pe_1_7_1_n77), .ZN(
        npu_inst_pe_1_7_1_n79) );
  INV_X1 npu_inst_pe_1_7_1_U44 ( .A(npu_inst_pe_1_7_1_n79), .ZN(
        npu_inst_pe_1_7_1_n35) );
  AOI222_X1 npu_inst_pe_1_7_1_U43 ( .A1(1'b0), .A2(npu_inst_pe_1_7_1_n1), .B1(
        npu_inst_pe_1_7_1_N79), .B2(npu_inst_pe_1_7_1_n76), .C1(
        npu_inst_pe_1_7_1_N71), .C2(npu_inst_pe_1_7_1_n77), .ZN(
        npu_inst_pe_1_7_1_n78) );
  INV_X1 npu_inst_pe_1_7_1_U42 ( .A(npu_inst_pe_1_7_1_n78), .ZN(
        npu_inst_pe_1_7_1_n34) );
  AND2_X1 npu_inst_pe_1_7_1_U41 ( .A1(npu_inst_pe_1_7_1_int_q_acc_0_), .A2(
        npu_inst_pe_1_7_1_n1), .ZN(npu_inst_int_data_res_7__1__0_) );
  AND2_X1 npu_inst_pe_1_7_1_U40 ( .A1(npu_inst_pe_1_7_1_n2), .A2(
        npu_inst_pe_1_7_1_int_q_acc_7_), .ZN(npu_inst_int_data_res_7__1__7_)
         );
  AND2_X1 npu_inst_pe_1_7_1_U39 ( .A1(npu_inst_pe_1_7_1_int_q_acc_1_), .A2(
        npu_inst_pe_1_7_1_n1), .ZN(npu_inst_int_data_res_7__1__1_) );
  AND2_X1 npu_inst_pe_1_7_1_U38 ( .A1(npu_inst_pe_1_7_1_int_q_acc_2_), .A2(
        npu_inst_pe_1_7_1_n1), .ZN(npu_inst_int_data_res_7__1__2_) );
  AND2_X1 npu_inst_pe_1_7_1_U37 ( .A1(npu_inst_pe_1_7_1_int_q_acc_3_), .A2(
        npu_inst_pe_1_7_1_n2), .ZN(npu_inst_int_data_res_7__1__3_) );
  AND2_X1 npu_inst_pe_1_7_1_U36 ( .A1(npu_inst_pe_1_7_1_int_q_acc_4_), .A2(
        npu_inst_pe_1_7_1_n2), .ZN(npu_inst_int_data_res_7__1__4_) );
  AND2_X1 npu_inst_pe_1_7_1_U35 ( .A1(npu_inst_pe_1_7_1_int_q_acc_5_), .A2(
        npu_inst_pe_1_7_1_n2), .ZN(npu_inst_int_data_res_7__1__5_) );
  AND2_X1 npu_inst_pe_1_7_1_U34 ( .A1(npu_inst_pe_1_7_1_int_q_acc_6_), .A2(
        npu_inst_pe_1_7_1_n2), .ZN(npu_inst_int_data_res_7__1__6_) );
  INV_X1 npu_inst_pe_1_7_1_U33 ( .A(npu_inst_pe_1_7_1_int_data_1_), .ZN(
        npu_inst_pe_1_7_1_n14) );
  AND2_X1 npu_inst_pe_1_7_1_U32 ( .A1(npu_inst_int_data_x_7__1__1_), .A2(
        npu_inst_pe_1_7_1_int_q_weight_1_), .ZN(npu_inst_pe_1_7_1_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_7_1_U31 ( .A1(npu_inst_int_data_x_7__1__0_), .A2(
        npu_inst_pe_1_7_1_int_q_weight_1_), .ZN(npu_inst_pe_1_7_1_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_7_1_U30 ( .A(npu_inst_pe_1_7_1_int_data_0_), .ZN(
        npu_inst_pe_1_7_1_n13) );
  INV_X1 npu_inst_pe_1_7_1_U29 ( .A(npu_inst_n67), .ZN(npu_inst_pe_1_7_1_n5)
         );
  OR3_X1 npu_inst_pe_1_7_1_U28 ( .A1(npu_inst_pe_1_7_1_n6), .A2(
        npu_inst_pe_1_7_1_n8), .A3(npu_inst_pe_1_7_1_n5), .ZN(
        npu_inst_pe_1_7_1_n56) );
  OR3_X1 npu_inst_pe_1_7_1_U27 ( .A1(npu_inst_pe_1_7_1_n5), .A2(
        npu_inst_pe_1_7_1_n8), .A3(npu_inst_pe_1_7_1_n7), .ZN(
        npu_inst_pe_1_7_1_n48) );
  INV_X1 npu_inst_pe_1_7_1_U26 ( .A(npu_inst_pe_1_7_1_n5), .ZN(
        npu_inst_pe_1_7_1_n4) );
  INV_X1 npu_inst_pe_1_7_1_U25 ( .A(npu_inst_n122), .ZN(npu_inst_pe_1_7_1_n12)
         );
  OR3_X1 npu_inst_pe_1_7_1_U24 ( .A1(npu_inst_pe_1_7_1_n4), .A2(
        npu_inst_pe_1_7_1_n8), .A3(npu_inst_pe_1_7_1_n7), .ZN(
        npu_inst_pe_1_7_1_n52) );
  OR3_X1 npu_inst_pe_1_7_1_U23 ( .A1(npu_inst_pe_1_7_1_n6), .A2(
        npu_inst_pe_1_7_1_n8), .A3(npu_inst_pe_1_7_1_n4), .ZN(
        npu_inst_pe_1_7_1_n60) );
  NOR2_X1 npu_inst_pe_1_7_1_U22 ( .A1(npu_inst_pe_1_7_1_n60), .A2(
        npu_inst_pe_1_7_1_n3), .ZN(npu_inst_pe_1_7_1_n58) );
  NOR2_X1 npu_inst_pe_1_7_1_U21 ( .A1(npu_inst_pe_1_7_1_n56), .A2(
        npu_inst_pe_1_7_1_n3), .ZN(npu_inst_pe_1_7_1_n54) );
  NOR2_X1 npu_inst_pe_1_7_1_U20 ( .A1(npu_inst_pe_1_7_1_n52), .A2(
        npu_inst_pe_1_7_1_n3), .ZN(npu_inst_pe_1_7_1_n50) );
  NOR2_X1 npu_inst_pe_1_7_1_U19 ( .A1(npu_inst_pe_1_7_1_n48), .A2(
        npu_inst_pe_1_7_1_n3), .ZN(npu_inst_pe_1_7_1_n46) );
  NOR2_X1 npu_inst_pe_1_7_1_U18 ( .A1(npu_inst_pe_1_7_1_n40), .A2(
        npu_inst_pe_1_7_1_n3), .ZN(npu_inst_pe_1_7_1_n38) );
  NOR2_X1 npu_inst_pe_1_7_1_U17 ( .A1(npu_inst_pe_1_7_1_n44), .A2(
        npu_inst_pe_1_7_1_n3), .ZN(npu_inst_pe_1_7_1_n42) );
  BUF_X1 npu_inst_pe_1_7_1_U16 ( .A(npu_inst_n93), .Z(npu_inst_pe_1_7_1_n8) );
  BUF_X1 npu_inst_pe_1_7_1_U15 ( .A(npu_inst_pe_1_7_1_n12), .Z(
        npu_inst_pe_1_7_1_n11) );
  BUF_X1 npu_inst_pe_1_7_1_U14 ( .A(npu_inst_pe_1_7_1_n12), .Z(
        npu_inst_pe_1_7_1_n10) );
  BUF_X1 npu_inst_pe_1_7_1_U13 ( .A(npu_inst_pe_1_7_1_n12), .Z(
        npu_inst_pe_1_7_1_n9) );
  INV_X1 npu_inst_pe_1_7_1_U12 ( .A(npu_inst_pe_1_7_1_n38), .ZN(
        npu_inst_pe_1_7_1_n118) );
  INV_X1 npu_inst_pe_1_7_1_U11 ( .A(npu_inst_pe_1_7_1_n58), .ZN(
        npu_inst_pe_1_7_1_n114) );
  INV_X1 npu_inst_pe_1_7_1_U10 ( .A(npu_inst_pe_1_7_1_n54), .ZN(
        npu_inst_pe_1_7_1_n115) );
  INV_X1 npu_inst_pe_1_7_1_U9 ( .A(npu_inst_pe_1_7_1_n50), .ZN(
        npu_inst_pe_1_7_1_n116) );
  INV_X1 npu_inst_pe_1_7_1_U8 ( .A(npu_inst_pe_1_7_1_n46), .ZN(
        npu_inst_pe_1_7_1_n117) );
  INV_X1 npu_inst_pe_1_7_1_U7 ( .A(npu_inst_pe_1_7_1_n42), .ZN(
        npu_inst_pe_1_7_1_n119) );
  BUF_X1 npu_inst_pe_1_7_1_U6 ( .A(npu_inst_n10), .Z(npu_inst_pe_1_7_1_n2) );
  BUF_X1 npu_inst_pe_1_7_1_U5 ( .A(npu_inst_n10), .Z(npu_inst_pe_1_7_1_n1) );
  NOR2_X1 npu_inst_pe_1_7_1_U4 ( .A1(npu_inst_pe_1_7_1_int_q_weight_0_), .A2(
        npu_inst_pe_1_7_1_n1), .ZN(npu_inst_pe_1_7_1_n76) );
  NOR2_X1 npu_inst_pe_1_7_1_U3 ( .A1(npu_inst_pe_1_7_1_n27), .A2(
        npu_inst_pe_1_7_1_n1), .ZN(npu_inst_pe_1_7_1_n77) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_7_1_n111), 
        .CK(npu_inst_pe_1_7_1_net2988), .RN(npu_inst_pe_1_7_1_n12), .Q(
        npu_inst_pe_1_7_1_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_7_1_n110), 
        .CK(npu_inst_pe_1_7_1_net2988), .RN(npu_inst_pe_1_7_1_n12), .Q(
        npu_inst_pe_1_7_1_int_q_reg_v_4__1_) );
  FA_X1 npu_inst_pe_1_7_1_sub_77_U2_1 ( .A(npu_inst_pe_1_7_1_int_q_acc_1_), 
        .B(npu_inst_pe_1_7_1_n14), .CI(npu_inst_pe_1_7_1_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_7_1_sub_77_carry_2_), .S(npu_inst_pe_1_7_1_N66) );
  FA_X1 npu_inst_pe_1_7_1_add_79_U1_1 ( .A(npu_inst_pe_1_7_1_int_q_acc_1_), 
        .B(npu_inst_pe_1_7_1_int_data_1_), .CI(
        npu_inst_pe_1_7_1_add_79_carry_1_), .CO(
        npu_inst_pe_1_7_1_add_79_carry_2_), .S(npu_inst_pe_1_7_1_N74) );
  NAND3_X1 npu_inst_pe_1_7_1_U109 ( .A1(npu_inst_pe_1_7_1_n5), .A2(
        npu_inst_pe_1_7_1_n7), .A3(npu_inst_pe_1_7_1_n8), .ZN(
        npu_inst_pe_1_7_1_n44) );
  NAND3_X1 npu_inst_pe_1_7_1_U108 ( .A1(npu_inst_pe_1_7_1_n4), .A2(
        npu_inst_pe_1_7_1_n7), .A3(npu_inst_pe_1_7_1_n8), .ZN(
        npu_inst_pe_1_7_1_n40) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_7_1_n34), .CK(
        npu_inst_pe_1_7_1_net2982), .RN(npu_inst_pe_1_7_1_n9), .Q(
        npu_inst_pe_1_7_1_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_7_1_n35), .CK(
        npu_inst_pe_1_7_1_net2982), .RN(npu_inst_pe_1_7_1_n9), .Q(
        npu_inst_pe_1_7_1_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_7_1_n36), .CK(
        npu_inst_pe_1_7_1_net2982), .RN(npu_inst_pe_1_7_1_n9), .Q(
        npu_inst_pe_1_7_1_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_7_1_n98), .CK(
        npu_inst_pe_1_7_1_net2982), .RN(npu_inst_pe_1_7_1_n9), .Q(
        npu_inst_pe_1_7_1_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_7_1_n99), .CK(
        npu_inst_pe_1_7_1_net2982), .RN(npu_inst_pe_1_7_1_n9), .Q(
        npu_inst_pe_1_7_1_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_7_1_n100), 
        .CK(npu_inst_pe_1_7_1_net2982), .RN(npu_inst_pe_1_7_1_n9), .Q(
        npu_inst_pe_1_7_1_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_7_1_n33), .CK(
        npu_inst_pe_1_7_1_net2982), .RN(npu_inst_pe_1_7_1_n9), .Q(
        npu_inst_pe_1_7_1_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_7_1_n101), 
        .CK(npu_inst_pe_1_7_1_net2982), .RN(npu_inst_pe_1_7_1_n9), .Q(
        npu_inst_pe_1_7_1_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_weight_reg_0_ ( .D(npu_inst_n108), .CK(
        npu_inst_pe_1_7_1_net2988), .RN(npu_inst_pe_1_7_1_n9), .Q(
        npu_inst_pe_1_7_1_int_q_weight_0_), .QN(npu_inst_pe_1_7_1_n27) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_weight_reg_1_ ( .D(npu_inst_n114), .CK(
        npu_inst_pe_1_7_1_net2988), .RN(npu_inst_pe_1_7_1_n9), .Q(
        npu_inst_pe_1_7_1_int_q_weight_1_), .QN(npu_inst_pe_1_7_1_n26) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_7_1_n113), 
        .CK(npu_inst_pe_1_7_1_net2988), .RN(npu_inst_pe_1_7_1_n9), .Q(
        npu_inst_pe_1_7_1_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_7_1_n112), 
        .CK(npu_inst_pe_1_7_1_net2988), .RN(npu_inst_pe_1_7_1_n9), .Q(
        npu_inst_pe_1_7_1_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_7_1_n109), 
        .CK(npu_inst_pe_1_7_1_net2988), .RN(npu_inst_pe_1_7_1_n10), .Q(
        npu_inst_pe_1_7_1_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_7_1_n108), 
        .CK(npu_inst_pe_1_7_1_net2988), .RN(npu_inst_pe_1_7_1_n10), .Q(
        npu_inst_pe_1_7_1_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_7_1_n107), 
        .CK(npu_inst_pe_1_7_1_net2988), .RN(npu_inst_pe_1_7_1_n10), .Q(
        npu_inst_pe_1_7_1_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_7_1_n106), 
        .CK(npu_inst_pe_1_7_1_net2988), .RN(npu_inst_pe_1_7_1_n10), .Q(
        npu_inst_pe_1_7_1_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_7_1_n105), 
        .CK(npu_inst_pe_1_7_1_net2988), .RN(npu_inst_pe_1_7_1_n10), .Q(
        npu_inst_pe_1_7_1_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_7_1_n104), 
        .CK(npu_inst_pe_1_7_1_net2988), .RN(npu_inst_pe_1_7_1_n10), .Q(
        npu_inst_pe_1_7_1_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_7_1_n103), 
        .CK(npu_inst_pe_1_7_1_net2988), .RN(npu_inst_pe_1_7_1_n10), .Q(
        npu_inst_pe_1_7_1_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_7_1_n102), 
        .CK(npu_inst_pe_1_7_1_net2988), .RN(npu_inst_pe_1_7_1_n10), .Q(
        npu_inst_pe_1_7_1_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_7_1_n86), 
        .CK(npu_inst_pe_1_7_1_net2988), .RN(npu_inst_pe_1_7_1_n10), .Q(
        npu_inst_pe_1_7_1_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_7_1_n87), 
        .CK(npu_inst_pe_1_7_1_net2988), .RN(npu_inst_pe_1_7_1_n10), .Q(
        npu_inst_pe_1_7_1_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_7_1_n88), 
        .CK(npu_inst_pe_1_7_1_net2988), .RN(npu_inst_pe_1_7_1_n11), .Q(
        npu_inst_pe_1_7_1_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_7_1_n89), 
        .CK(npu_inst_pe_1_7_1_net2988), .RN(npu_inst_pe_1_7_1_n11), .Q(
        npu_inst_pe_1_7_1_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_7_1_n90), 
        .CK(npu_inst_pe_1_7_1_net2988), .RN(npu_inst_pe_1_7_1_n11), .Q(
        npu_inst_pe_1_7_1_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_7_1_n91), 
        .CK(npu_inst_pe_1_7_1_net2988), .RN(npu_inst_pe_1_7_1_n11), .Q(
        npu_inst_pe_1_7_1_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_7_1_n92), 
        .CK(npu_inst_pe_1_7_1_net2988), .RN(npu_inst_pe_1_7_1_n11), .Q(
        npu_inst_pe_1_7_1_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_7_1_n93), 
        .CK(npu_inst_pe_1_7_1_net2988), .RN(npu_inst_pe_1_7_1_n11), .Q(
        npu_inst_pe_1_7_1_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_7_1_n94), 
        .CK(npu_inst_pe_1_7_1_net2988), .RN(npu_inst_pe_1_7_1_n11), .Q(
        npu_inst_pe_1_7_1_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_7_1_n95), 
        .CK(npu_inst_pe_1_7_1_net2988), .RN(npu_inst_pe_1_7_1_n11), .Q(
        npu_inst_pe_1_7_1_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_7_1_n96), 
        .CK(npu_inst_pe_1_7_1_net2988), .RN(npu_inst_pe_1_7_1_n11), .Q(
        npu_inst_pe_1_7_1_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_7_1_n97), 
        .CK(npu_inst_pe_1_7_1_net2988), .RN(npu_inst_pe_1_7_1_n11), .Q(
        npu_inst_pe_1_7_1_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_7_1_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_7_1_N84), .SE(1'b0), .GCK(npu_inst_pe_1_7_1_net2982) );
  CLKGATETST_X1 npu_inst_pe_1_7_1_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n61), .SE(1'b0), .GCK(npu_inst_pe_1_7_1_net2988) );
  MUX2_X1 npu_inst_pe_1_7_2_U162 ( .A(npu_inst_pe_1_7_2_n32), .B(
        npu_inst_pe_1_7_2_n29), .S(npu_inst_pe_1_7_2_n8), .Z(
        npu_inst_pe_1_7_2_N93) );
  MUX2_X1 npu_inst_pe_1_7_2_U161 ( .A(npu_inst_pe_1_7_2_n31), .B(
        npu_inst_pe_1_7_2_n30), .S(npu_inst_pe_1_7_2_n6), .Z(
        npu_inst_pe_1_7_2_n32) );
  MUX2_X1 npu_inst_pe_1_7_2_U160 ( .A(npu_inst_pe_1_7_2_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_7_2_int_q_reg_v_1__0_), .S(npu_inst_pe_1_7_2_n4), .Z(
        npu_inst_pe_1_7_2_n31) );
  MUX2_X1 npu_inst_pe_1_7_2_U159 ( .A(npu_inst_pe_1_7_2_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_7_2_int_q_reg_v_3__0_), .S(npu_inst_pe_1_7_2_n4), .Z(
        npu_inst_pe_1_7_2_n30) );
  MUX2_X1 npu_inst_pe_1_7_2_U158 ( .A(npu_inst_pe_1_7_2_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_7_2_int_q_reg_v_5__0_), .S(npu_inst_pe_1_7_2_n4), .Z(
        npu_inst_pe_1_7_2_n29) );
  MUX2_X1 npu_inst_pe_1_7_2_U157 ( .A(npu_inst_pe_1_7_2_n28), .B(
        npu_inst_pe_1_7_2_n23), .S(npu_inst_pe_1_7_2_n8), .Z(
        npu_inst_pe_1_7_2_N94) );
  MUX2_X1 npu_inst_pe_1_7_2_U156 ( .A(npu_inst_pe_1_7_2_n25), .B(
        npu_inst_pe_1_7_2_n24), .S(npu_inst_pe_1_7_2_n6), .Z(
        npu_inst_pe_1_7_2_n28) );
  MUX2_X1 npu_inst_pe_1_7_2_U155 ( .A(npu_inst_pe_1_7_2_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_7_2_int_q_reg_v_1__1_), .S(npu_inst_pe_1_7_2_n4), .Z(
        npu_inst_pe_1_7_2_n25) );
  MUX2_X1 npu_inst_pe_1_7_2_U154 ( .A(npu_inst_pe_1_7_2_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_7_2_int_q_reg_v_3__1_), .S(npu_inst_pe_1_7_2_n4), .Z(
        npu_inst_pe_1_7_2_n24) );
  MUX2_X1 npu_inst_pe_1_7_2_U153 ( .A(npu_inst_pe_1_7_2_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_7_2_int_q_reg_v_5__1_), .S(npu_inst_pe_1_7_2_n4), .Z(
        npu_inst_pe_1_7_2_n23) );
  MUX2_X1 npu_inst_pe_1_7_2_U152 ( .A(npu_inst_pe_1_7_2_n22), .B(
        npu_inst_pe_1_7_2_n19), .S(npu_inst_pe_1_7_2_n8), .Z(
        npu_inst_int_data_x_7__2__1_) );
  MUX2_X1 npu_inst_pe_1_7_2_U151 ( .A(npu_inst_pe_1_7_2_n21), .B(
        npu_inst_pe_1_7_2_n20), .S(npu_inst_pe_1_7_2_n6), .Z(
        npu_inst_pe_1_7_2_n22) );
  MUX2_X1 npu_inst_pe_1_7_2_U150 ( .A(npu_inst_pe_1_7_2_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_7_2_int_q_reg_h_1__1_), .S(npu_inst_pe_1_7_2_n4), .Z(
        npu_inst_pe_1_7_2_n21) );
  MUX2_X1 npu_inst_pe_1_7_2_U149 ( .A(npu_inst_pe_1_7_2_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_7_2_int_q_reg_h_3__1_), .S(npu_inst_pe_1_7_2_n4), .Z(
        npu_inst_pe_1_7_2_n20) );
  MUX2_X1 npu_inst_pe_1_7_2_U148 ( .A(npu_inst_pe_1_7_2_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_7_2_int_q_reg_h_5__1_), .S(npu_inst_pe_1_7_2_n4), .Z(
        npu_inst_pe_1_7_2_n19) );
  MUX2_X1 npu_inst_pe_1_7_2_U147 ( .A(npu_inst_pe_1_7_2_n18), .B(
        npu_inst_pe_1_7_2_n15), .S(npu_inst_pe_1_7_2_n8), .Z(
        npu_inst_int_data_x_7__2__0_) );
  MUX2_X1 npu_inst_pe_1_7_2_U146 ( .A(npu_inst_pe_1_7_2_n17), .B(
        npu_inst_pe_1_7_2_n16), .S(npu_inst_pe_1_7_2_n6), .Z(
        npu_inst_pe_1_7_2_n18) );
  MUX2_X1 npu_inst_pe_1_7_2_U145 ( .A(npu_inst_pe_1_7_2_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_7_2_int_q_reg_h_1__0_), .S(npu_inst_pe_1_7_2_n4), .Z(
        npu_inst_pe_1_7_2_n17) );
  MUX2_X1 npu_inst_pe_1_7_2_U144 ( .A(npu_inst_pe_1_7_2_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_7_2_int_q_reg_h_3__0_), .S(npu_inst_pe_1_7_2_n4), .Z(
        npu_inst_pe_1_7_2_n16) );
  MUX2_X1 npu_inst_pe_1_7_2_U143 ( .A(npu_inst_pe_1_7_2_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_7_2_int_q_reg_h_5__0_), .S(npu_inst_pe_1_7_2_n4), .Z(
        npu_inst_pe_1_7_2_n15) );
  XOR2_X1 npu_inst_pe_1_7_2_U142 ( .A(npu_inst_pe_1_7_2_int_data_0_), .B(
        npu_inst_pe_1_7_2_int_q_acc_0_), .Z(npu_inst_pe_1_7_2_N73) );
  AND2_X1 npu_inst_pe_1_7_2_U141 ( .A1(npu_inst_pe_1_7_2_int_q_acc_0_), .A2(
        npu_inst_pe_1_7_2_int_data_0_), .ZN(npu_inst_pe_1_7_2_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_7_2_U140 ( .A(npu_inst_pe_1_7_2_int_q_acc_0_), .B(
        npu_inst_pe_1_7_2_n13), .ZN(npu_inst_pe_1_7_2_N65) );
  OR2_X1 npu_inst_pe_1_7_2_U139 ( .A1(npu_inst_pe_1_7_2_n13), .A2(
        npu_inst_pe_1_7_2_int_q_acc_0_), .ZN(npu_inst_pe_1_7_2_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_7_2_U138 ( .A(npu_inst_pe_1_7_2_int_q_acc_2_), .B(
        npu_inst_pe_1_7_2_add_79_carry_2_), .Z(npu_inst_pe_1_7_2_N75) );
  AND2_X1 npu_inst_pe_1_7_2_U137 ( .A1(npu_inst_pe_1_7_2_add_79_carry_2_), 
        .A2(npu_inst_pe_1_7_2_int_q_acc_2_), .ZN(
        npu_inst_pe_1_7_2_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_7_2_U136 ( .A(npu_inst_pe_1_7_2_int_q_acc_3_), .B(
        npu_inst_pe_1_7_2_add_79_carry_3_), .Z(npu_inst_pe_1_7_2_N76) );
  AND2_X1 npu_inst_pe_1_7_2_U135 ( .A1(npu_inst_pe_1_7_2_add_79_carry_3_), 
        .A2(npu_inst_pe_1_7_2_int_q_acc_3_), .ZN(
        npu_inst_pe_1_7_2_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_7_2_U134 ( .A(npu_inst_pe_1_7_2_int_q_acc_4_), .B(
        npu_inst_pe_1_7_2_add_79_carry_4_), .Z(npu_inst_pe_1_7_2_N77) );
  AND2_X1 npu_inst_pe_1_7_2_U133 ( .A1(npu_inst_pe_1_7_2_add_79_carry_4_), 
        .A2(npu_inst_pe_1_7_2_int_q_acc_4_), .ZN(
        npu_inst_pe_1_7_2_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_7_2_U132 ( .A(npu_inst_pe_1_7_2_int_q_acc_5_), .B(
        npu_inst_pe_1_7_2_add_79_carry_5_), .Z(npu_inst_pe_1_7_2_N78) );
  AND2_X1 npu_inst_pe_1_7_2_U131 ( .A1(npu_inst_pe_1_7_2_add_79_carry_5_), 
        .A2(npu_inst_pe_1_7_2_int_q_acc_5_), .ZN(
        npu_inst_pe_1_7_2_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_7_2_U130 ( .A(npu_inst_pe_1_7_2_int_q_acc_6_), .B(
        npu_inst_pe_1_7_2_add_79_carry_6_), .Z(npu_inst_pe_1_7_2_N79) );
  AND2_X1 npu_inst_pe_1_7_2_U129 ( .A1(npu_inst_pe_1_7_2_add_79_carry_6_), 
        .A2(npu_inst_pe_1_7_2_int_q_acc_6_), .ZN(
        npu_inst_pe_1_7_2_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_7_2_U128 ( .A(npu_inst_pe_1_7_2_int_q_acc_7_), .B(
        npu_inst_pe_1_7_2_add_79_carry_7_), .Z(npu_inst_pe_1_7_2_N80) );
  XNOR2_X1 npu_inst_pe_1_7_2_U127 ( .A(npu_inst_pe_1_7_2_sub_77_carry_2_), .B(
        npu_inst_pe_1_7_2_int_q_acc_2_), .ZN(npu_inst_pe_1_7_2_N67) );
  OR2_X1 npu_inst_pe_1_7_2_U126 ( .A1(npu_inst_pe_1_7_2_int_q_acc_2_), .A2(
        npu_inst_pe_1_7_2_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_7_2_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_7_2_U125 ( .A(npu_inst_pe_1_7_2_sub_77_carry_3_), .B(
        npu_inst_pe_1_7_2_int_q_acc_3_), .ZN(npu_inst_pe_1_7_2_N68) );
  OR2_X1 npu_inst_pe_1_7_2_U124 ( .A1(npu_inst_pe_1_7_2_int_q_acc_3_), .A2(
        npu_inst_pe_1_7_2_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_7_2_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_7_2_U123 ( .A(npu_inst_pe_1_7_2_sub_77_carry_4_), .B(
        npu_inst_pe_1_7_2_int_q_acc_4_), .ZN(npu_inst_pe_1_7_2_N69) );
  OR2_X1 npu_inst_pe_1_7_2_U122 ( .A1(npu_inst_pe_1_7_2_int_q_acc_4_), .A2(
        npu_inst_pe_1_7_2_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_7_2_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_7_2_U121 ( .A(npu_inst_pe_1_7_2_sub_77_carry_5_), .B(
        npu_inst_pe_1_7_2_int_q_acc_5_), .ZN(npu_inst_pe_1_7_2_N70) );
  OR2_X1 npu_inst_pe_1_7_2_U120 ( .A1(npu_inst_pe_1_7_2_int_q_acc_5_), .A2(
        npu_inst_pe_1_7_2_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_7_2_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_7_2_U119 ( .A(npu_inst_pe_1_7_2_sub_77_carry_6_), .B(
        npu_inst_pe_1_7_2_int_q_acc_6_), .ZN(npu_inst_pe_1_7_2_N71) );
  OR2_X1 npu_inst_pe_1_7_2_U118 ( .A1(npu_inst_pe_1_7_2_int_q_acc_6_), .A2(
        npu_inst_pe_1_7_2_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_7_2_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_7_2_U117 ( .A(npu_inst_pe_1_7_2_int_q_acc_7_), .B(
        npu_inst_pe_1_7_2_sub_77_carry_7_), .ZN(npu_inst_pe_1_7_2_N72) );
  INV_X1 npu_inst_pe_1_7_2_U116 ( .A(npu_inst_n75), .ZN(npu_inst_pe_1_7_2_n7)
         );
  INV_X1 npu_inst_pe_1_7_2_U115 ( .A(npu_inst_pe_1_7_2_n7), .ZN(
        npu_inst_pe_1_7_2_n6) );
  INV_X1 npu_inst_pe_1_7_2_U114 ( .A(npu_inst_n52), .ZN(npu_inst_pe_1_7_2_n3)
         );
  AOI22_X1 npu_inst_pe_1_7_2_U113 ( .A1(npu_inst_pe_1_7_2_n38), .A2(
        int_i_data_v_npu[11]), .B1(npu_inst_pe_1_7_2_n118), .B2(
        npu_inst_pe_1_7_2_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_7_2_n39) );
  INV_X1 npu_inst_pe_1_7_2_U112 ( .A(npu_inst_pe_1_7_2_n39), .ZN(
        npu_inst_pe_1_7_2_n112) );
  AOI22_X1 npu_inst_pe_1_7_2_U111 ( .A1(npu_inst_pe_1_7_2_n38), .A2(
        int_i_data_v_npu[10]), .B1(npu_inst_pe_1_7_2_n118), .B2(
        npu_inst_pe_1_7_2_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_7_2_n37) );
  INV_X1 npu_inst_pe_1_7_2_U110 ( .A(npu_inst_pe_1_7_2_n37), .ZN(
        npu_inst_pe_1_7_2_n113) );
  AOI22_X1 npu_inst_pe_1_7_2_U107 ( .A1(int_i_data_v_npu[11]), .A2(
        npu_inst_pe_1_7_2_n58), .B1(npu_inst_pe_1_7_2_n114), .B2(
        npu_inst_pe_1_7_2_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_7_2_n59) );
  INV_X1 npu_inst_pe_1_7_2_U106 ( .A(npu_inst_pe_1_7_2_n59), .ZN(
        npu_inst_pe_1_7_2_n102) );
  AOI22_X1 npu_inst_pe_1_7_2_U105 ( .A1(int_i_data_v_npu[10]), .A2(
        npu_inst_pe_1_7_2_n58), .B1(npu_inst_pe_1_7_2_n114), .B2(
        npu_inst_pe_1_7_2_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_7_2_n57) );
  INV_X1 npu_inst_pe_1_7_2_U104 ( .A(npu_inst_pe_1_7_2_n57), .ZN(
        npu_inst_pe_1_7_2_n103) );
  AOI22_X1 npu_inst_pe_1_7_2_U103 ( .A1(int_i_data_v_npu[11]), .A2(
        npu_inst_pe_1_7_2_n54), .B1(npu_inst_pe_1_7_2_n115), .B2(
        npu_inst_pe_1_7_2_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_7_2_n55) );
  INV_X1 npu_inst_pe_1_7_2_U102 ( .A(npu_inst_pe_1_7_2_n55), .ZN(
        npu_inst_pe_1_7_2_n104) );
  AOI22_X1 npu_inst_pe_1_7_2_U101 ( .A1(int_i_data_v_npu[10]), .A2(
        npu_inst_pe_1_7_2_n54), .B1(npu_inst_pe_1_7_2_n115), .B2(
        npu_inst_pe_1_7_2_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_7_2_n53) );
  INV_X1 npu_inst_pe_1_7_2_U100 ( .A(npu_inst_pe_1_7_2_n53), .ZN(
        npu_inst_pe_1_7_2_n105) );
  AOI22_X1 npu_inst_pe_1_7_2_U99 ( .A1(int_i_data_v_npu[11]), .A2(
        npu_inst_pe_1_7_2_n50), .B1(npu_inst_pe_1_7_2_n116), .B2(
        npu_inst_pe_1_7_2_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_7_2_n51) );
  INV_X1 npu_inst_pe_1_7_2_U98 ( .A(npu_inst_pe_1_7_2_n51), .ZN(
        npu_inst_pe_1_7_2_n106) );
  AOI22_X1 npu_inst_pe_1_7_2_U97 ( .A1(int_i_data_v_npu[10]), .A2(
        npu_inst_pe_1_7_2_n50), .B1(npu_inst_pe_1_7_2_n116), .B2(
        npu_inst_pe_1_7_2_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_7_2_n49) );
  INV_X1 npu_inst_pe_1_7_2_U96 ( .A(npu_inst_pe_1_7_2_n49), .ZN(
        npu_inst_pe_1_7_2_n107) );
  AOI22_X1 npu_inst_pe_1_7_2_U95 ( .A1(int_i_data_v_npu[11]), .A2(
        npu_inst_pe_1_7_2_n46), .B1(npu_inst_pe_1_7_2_n117), .B2(
        npu_inst_pe_1_7_2_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_7_2_n47) );
  INV_X1 npu_inst_pe_1_7_2_U94 ( .A(npu_inst_pe_1_7_2_n47), .ZN(
        npu_inst_pe_1_7_2_n108) );
  AOI22_X1 npu_inst_pe_1_7_2_U93 ( .A1(int_i_data_v_npu[10]), .A2(
        npu_inst_pe_1_7_2_n46), .B1(npu_inst_pe_1_7_2_n117), .B2(
        npu_inst_pe_1_7_2_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_7_2_n45) );
  INV_X1 npu_inst_pe_1_7_2_U92 ( .A(npu_inst_pe_1_7_2_n45), .ZN(
        npu_inst_pe_1_7_2_n109) );
  AOI22_X1 npu_inst_pe_1_7_2_U91 ( .A1(int_i_data_v_npu[11]), .A2(
        npu_inst_pe_1_7_2_n42), .B1(npu_inst_pe_1_7_2_n119), .B2(
        npu_inst_pe_1_7_2_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_7_2_n43) );
  INV_X1 npu_inst_pe_1_7_2_U90 ( .A(npu_inst_pe_1_7_2_n43), .ZN(
        npu_inst_pe_1_7_2_n110) );
  AOI22_X1 npu_inst_pe_1_7_2_U89 ( .A1(int_i_data_v_npu[10]), .A2(
        npu_inst_pe_1_7_2_n42), .B1(npu_inst_pe_1_7_2_n119), .B2(
        npu_inst_pe_1_7_2_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_7_2_n41) );
  INV_X1 npu_inst_pe_1_7_2_U88 ( .A(npu_inst_pe_1_7_2_n41), .ZN(
        npu_inst_pe_1_7_2_n111) );
  NAND2_X1 npu_inst_pe_1_7_2_U87 ( .A1(npu_inst_pe_1_7_2_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_7_2_n60), .ZN(npu_inst_pe_1_7_2_n74) );
  OAI21_X1 npu_inst_pe_1_7_2_U86 ( .B1(npu_inst_pe_1_7_2_n63), .B2(
        npu_inst_pe_1_7_2_n60), .A(npu_inst_pe_1_7_2_n74), .ZN(
        npu_inst_pe_1_7_2_n97) );
  NAND2_X1 npu_inst_pe_1_7_2_U85 ( .A1(npu_inst_pe_1_7_2_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_7_2_n60), .ZN(npu_inst_pe_1_7_2_n73) );
  OAI21_X1 npu_inst_pe_1_7_2_U84 ( .B1(npu_inst_pe_1_7_2_n61), .B2(
        npu_inst_pe_1_7_2_n60), .A(npu_inst_pe_1_7_2_n73), .ZN(
        npu_inst_pe_1_7_2_n96) );
  NAND2_X1 npu_inst_pe_1_7_2_U83 ( .A1(npu_inst_pe_1_7_2_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_7_2_n56), .ZN(npu_inst_pe_1_7_2_n72) );
  OAI21_X1 npu_inst_pe_1_7_2_U82 ( .B1(npu_inst_pe_1_7_2_n63), .B2(
        npu_inst_pe_1_7_2_n56), .A(npu_inst_pe_1_7_2_n72), .ZN(
        npu_inst_pe_1_7_2_n95) );
  NAND2_X1 npu_inst_pe_1_7_2_U81 ( .A1(npu_inst_pe_1_7_2_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_7_2_n56), .ZN(npu_inst_pe_1_7_2_n71) );
  OAI21_X1 npu_inst_pe_1_7_2_U80 ( .B1(npu_inst_pe_1_7_2_n61), .B2(
        npu_inst_pe_1_7_2_n56), .A(npu_inst_pe_1_7_2_n71), .ZN(
        npu_inst_pe_1_7_2_n94) );
  NAND2_X1 npu_inst_pe_1_7_2_U79 ( .A1(npu_inst_pe_1_7_2_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_7_2_n52), .ZN(npu_inst_pe_1_7_2_n70) );
  OAI21_X1 npu_inst_pe_1_7_2_U78 ( .B1(npu_inst_pe_1_7_2_n63), .B2(
        npu_inst_pe_1_7_2_n52), .A(npu_inst_pe_1_7_2_n70), .ZN(
        npu_inst_pe_1_7_2_n93) );
  NAND2_X1 npu_inst_pe_1_7_2_U77 ( .A1(npu_inst_pe_1_7_2_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_7_2_n52), .ZN(npu_inst_pe_1_7_2_n69) );
  OAI21_X1 npu_inst_pe_1_7_2_U76 ( .B1(npu_inst_pe_1_7_2_n61), .B2(
        npu_inst_pe_1_7_2_n52), .A(npu_inst_pe_1_7_2_n69), .ZN(
        npu_inst_pe_1_7_2_n92) );
  NAND2_X1 npu_inst_pe_1_7_2_U75 ( .A1(npu_inst_pe_1_7_2_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_7_2_n48), .ZN(npu_inst_pe_1_7_2_n68) );
  OAI21_X1 npu_inst_pe_1_7_2_U74 ( .B1(npu_inst_pe_1_7_2_n63), .B2(
        npu_inst_pe_1_7_2_n48), .A(npu_inst_pe_1_7_2_n68), .ZN(
        npu_inst_pe_1_7_2_n91) );
  NAND2_X1 npu_inst_pe_1_7_2_U73 ( .A1(npu_inst_pe_1_7_2_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_7_2_n48), .ZN(npu_inst_pe_1_7_2_n67) );
  OAI21_X1 npu_inst_pe_1_7_2_U72 ( .B1(npu_inst_pe_1_7_2_n61), .B2(
        npu_inst_pe_1_7_2_n48), .A(npu_inst_pe_1_7_2_n67), .ZN(
        npu_inst_pe_1_7_2_n90) );
  NAND2_X1 npu_inst_pe_1_7_2_U71 ( .A1(npu_inst_pe_1_7_2_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_7_2_n44), .ZN(npu_inst_pe_1_7_2_n66) );
  OAI21_X1 npu_inst_pe_1_7_2_U70 ( .B1(npu_inst_pe_1_7_2_n63), .B2(
        npu_inst_pe_1_7_2_n44), .A(npu_inst_pe_1_7_2_n66), .ZN(
        npu_inst_pe_1_7_2_n89) );
  NAND2_X1 npu_inst_pe_1_7_2_U69 ( .A1(npu_inst_pe_1_7_2_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_7_2_n44), .ZN(npu_inst_pe_1_7_2_n65) );
  OAI21_X1 npu_inst_pe_1_7_2_U68 ( .B1(npu_inst_pe_1_7_2_n61), .B2(
        npu_inst_pe_1_7_2_n44), .A(npu_inst_pe_1_7_2_n65), .ZN(
        npu_inst_pe_1_7_2_n88) );
  NAND2_X1 npu_inst_pe_1_7_2_U67 ( .A1(npu_inst_pe_1_7_2_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_7_2_n40), .ZN(npu_inst_pe_1_7_2_n64) );
  OAI21_X1 npu_inst_pe_1_7_2_U66 ( .B1(npu_inst_pe_1_7_2_n63), .B2(
        npu_inst_pe_1_7_2_n40), .A(npu_inst_pe_1_7_2_n64), .ZN(
        npu_inst_pe_1_7_2_n87) );
  NAND2_X1 npu_inst_pe_1_7_2_U65 ( .A1(npu_inst_pe_1_7_2_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_7_2_n40), .ZN(npu_inst_pe_1_7_2_n62) );
  OAI21_X1 npu_inst_pe_1_7_2_U64 ( .B1(npu_inst_pe_1_7_2_n61), .B2(
        npu_inst_pe_1_7_2_n40), .A(npu_inst_pe_1_7_2_n62), .ZN(
        npu_inst_pe_1_7_2_n86) );
  AND2_X1 npu_inst_pe_1_7_2_U63 ( .A1(npu_inst_pe_1_7_2_N93), .A2(npu_inst_n52), .ZN(npu_inst_int_data_y_7__2__0_) );
  AND2_X1 npu_inst_pe_1_7_2_U62 ( .A1(npu_inst_n52), .A2(npu_inst_pe_1_7_2_N94), .ZN(npu_inst_int_data_y_7__2__1_) );
  AOI22_X1 npu_inst_pe_1_7_2_U61 ( .A1(npu_inst_n52), .A2(int_i_data_v_npu[11]), .B1(npu_inst_pe_1_7_2_n3), .B2(npu_inst_int_data_x_7__3__1_), .ZN(
        npu_inst_pe_1_7_2_n63) );
  AOI22_X1 npu_inst_pe_1_7_2_U60 ( .A1(npu_inst_n52), .A2(int_i_data_v_npu[10]), .B1(npu_inst_pe_1_7_2_n3), .B2(npu_inst_int_data_x_7__3__0_), .ZN(
        npu_inst_pe_1_7_2_n61) );
  NOR3_X1 npu_inst_pe_1_7_2_U59 ( .A1(npu_inst_pe_1_7_2_n26), .A2(npu_inst_n52), .A3(npu_inst_int_ckg[5]), .ZN(npu_inst_pe_1_7_2_n85) );
  OR2_X1 npu_inst_pe_1_7_2_U58 ( .A1(npu_inst_pe_1_7_2_n85), .A2(
        npu_inst_pe_1_7_2_n2), .ZN(npu_inst_pe_1_7_2_N84) );
  AOI222_X1 npu_inst_pe_1_7_2_U57 ( .A1(1'b0), .A2(npu_inst_pe_1_7_2_n1), .B1(
        npu_inst_pe_1_7_2_N73), .B2(npu_inst_pe_1_7_2_n76), .C1(
        npu_inst_pe_1_7_2_N65), .C2(npu_inst_pe_1_7_2_n77), .ZN(
        npu_inst_pe_1_7_2_n84) );
  INV_X1 npu_inst_pe_1_7_2_U56 ( .A(npu_inst_pe_1_7_2_n84), .ZN(
        npu_inst_pe_1_7_2_n101) );
  AOI222_X1 npu_inst_pe_1_7_2_U55 ( .A1(1'b0), .A2(npu_inst_pe_1_7_2_n1), .B1(
        npu_inst_pe_1_7_2_N80), .B2(npu_inst_pe_1_7_2_n76), .C1(
        npu_inst_pe_1_7_2_N72), .C2(npu_inst_pe_1_7_2_n77), .ZN(
        npu_inst_pe_1_7_2_n75) );
  INV_X1 npu_inst_pe_1_7_2_U54 ( .A(npu_inst_pe_1_7_2_n75), .ZN(
        npu_inst_pe_1_7_2_n33) );
  AOI222_X1 npu_inst_pe_1_7_2_U53 ( .A1(1'b0), .A2(npu_inst_pe_1_7_2_n1), .B1(
        npu_inst_pe_1_7_2_N74), .B2(npu_inst_pe_1_7_2_n76), .C1(
        npu_inst_pe_1_7_2_N66), .C2(npu_inst_pe_1_7_2_n77), .ZN(
        npu_inst_pe_1_7_2_n83) );
  INV_X1 npu_inst_pe_1_7_2_U52 ( .A(npu_inst_pe_1_7_2_n83), .ZN(
        npu_inst_pe_1_7_2_n100) );
  AOI222_X1 npu_inst_pe_1_7_2_U51 ( .A1(1'b0), .A2(npu_inst_pe_1_7_2_n1), .B1(
        npu_inst_pe_1_7_2_N75), .B2(npu_inst_pe_1_7_2_n76), .C1(
        npu_inst_pe_1_7_2_N67), .C2(npu_inst_pe_1_7_2_n77), .ZN(
        npu_inst_pe_1_7_2_n82) );
  INV_X1 npu_inst_pe_1_7_2_U50 ( .A(npu_inst_pe_1_7_2_n82), .ZN(
        npu_inst_pe_1_7_2_n99) );
  AOI222_X1 npu_inst_pe_1_7_2_U49 ( .A1(1'b0), .A2(npu_inst_pe_1_7_2_n1), .B1(
        npu_inst_pe_1_7_2_N76), .B2(npu_inst_pe_1_7_2_n76), .C1(
        npu_inst_pe_1_7_2_N68), .C2(npu_inst_pe_1_7_2_n77), .ZN(
        npu_inst_pe_1_7_2_n81) );
  INV_X1 npu_inst_pe_1_7_2_U48 ( .A(npu_inst_pe_1_7_2_n81), .ZN(
        npu_inst_pe_1_7_2_n98) );
  AOI222_X1 npu_inst_pe_1_7_2_U47 ( .A1(1'b0), .A2(npu_inst_pe_1_7_2_n1), .B1(
        npu_inst_pe_1_7_2_N77), .B2(npu_inst_pe_1_7_2_n76), .C1(
        npu_inst_pe_1_7_2_N69), .C2(npu_inst_pe_1_7_2_n77), .ZN(
        npu_inst_pe_1_7_2_n80) );
  INV_X1 npu_inst_pe_1_7_2_U46 ( .A(npu_inst_pe_1_7_2_n80), .ZN(
        npu_inst_pe_1_7_2_n36) );
  AOI222_X1 npu_inst_pe_1_7_2_U45 ( .A1(1'b0), .A2(npu_inst_pe_1_7_2_n1), .B1(
        npu_inst_pe_1_7_2_N78), .B2(npu_inst_pe_1_7_2_n76), .C1(
        npu_inst_pe_1_7_2_N70), .C2(npu_inst_pe_1_7_2_n77), .ZN(
        npu_inst_pe_1_7_2_n79) );
  INV_X1 npu_inst_pe_1_7_2_U44 ( .A(npu_inst_pe_1_7_2_n79), .ZN(
        npu_inst_pe_1_7_2_n35) );
  AOI222_X1 npu_inst_pe_1_7_2_U43 ( .A1(1'b0), .A2(npu_inst_pe_1_7_2_n1), .B1(
        npu_inst_pe_1_7_2_N79), .B2(npu_inst_pe_1_7_2_n76), .C1(
        npu_inst_pe_1_7_2_N71), .C2(npu_inst_pe_1_7_2_n77), .ZN(
        npu_inst_pe_1_7_2_n78) );
  INV_X1 npu_inst_pe_1_7_2_U42 ( .A(npu_inst_pe_1_7_2_n78), .ZN(
        npu_inst_pe_1_7_2_n34) );
  AND2_X1 npu_inst_pe_1_7_2_U41 ( .A1(npu_inst_pe_1_7_2_int_q_acc_0_), .A2(
        npu_inst_pe_1_7_2_n1), .ZN(npu_inst_int_data_res_7__2__0_) );
  AND2_X1 npu_inst_pe_1_7_2_U40 ( .A1(npu_inst_pe_1_7_2_n2), .A2(
        npu_inst_pe_1_7_2_int_q_acc_7_), .ZN(npu_inst_int_data_res_7__2__7_)
         );
  AND2_X1 npu_inst_pe_1_7_2_U39 ( .A1(npu_inst_pe_1_7_2_int_q_acc_1_), .A2(
        npu_inst_pe_1_7_2_n1), .ZN(npu_inst_int_data_res_7__2__1_) );
  AND2_X1 npu_inst_pe_1_7_2_U38 ( .A1(npu_inst_pe_1_7_2_int_q_acc_2_), .A2(
        npu_inst_pe_1_7_2_n1), .ZN(npu_inst_int_data_res_7__2__2_) );
  AND2_X1 npu_inst_pe_1_7_2_U37 ( .A1(npu_inst_pe_1_7_2_int_q_acc_3_), .A2(
        npu_inst_pe_1_7_2_n2), .ZN(npu_inst_int_data_res_7__2__3_) );
  AND2_X1 npu_inst_pe_1_7_2_U36 ( .A1(npu_inst_pe_1_7_2_int_q_acc_4_), .A2(
        npu_inst_pe_1_7_2_n2), .ZN(npu_inst_int_data_res_7__2__4_) );
  AND2_X1 npu_inst_pe_1_7_2_U35 ( .A1(npu_inst_pe_1_7_2_int_q_acc_5_), .A2(
        npu_inst_pe_1_7_2_n2), .ZN(npu_inst_int_data_res_7__2__5_) );
  AND2_X1 npu_inst_pe_1_7_2_U34 ( .A1(npu_inst_pe_1_7_2_int_q_acc_6_), .A2(
        npu_inst_pe_1_7_2_n2), .ZN(npu_inst_int_data_res_7__2__6_) );
  INV_X1 npu_inst_pe_1_7_2_U33 ( .A(npu_inst_pe_1_7_2_int_data_1_), .ZN(
        npu_inst_pe_1_7_2_n14) );
  AND2_X1 npu_inst_pe_1_7_2_U32 ( .A1(npu_inst_int_data_x_7__2__1_), .A2(
        npu_inst_pe_1_7_2_int_q_weight_1_), .ZN(npu_inst_pe_1_7_2_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_7_2_U31 ( .A1(npu_inst_int_data_x_7__2__0_), .A2(
        npu_inst_pe_1_7_2_int_q_weight_1_), .ZN(npu_inst_pe_1_7_2_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_7_2_U30 ( .A(npu_inst_pe_1_7_2_int_data_0_), .ZN(
        npu_inst_pe_1_7_2_n13) );
  INV_X1 npu_inst_pe_1_7_2_U29 ( .A(npu_inst_n67), .ZN(npu_inst_pe_1_7_2_n5)
         );
  OR3_X1 npu_inst_pe_1_7_2_U28 ( .A1(npu_inst_pe_1_7_2_n6), .A2(
        npu_inst_pe_1_7_2_n8), .A3(npu_inst_pe_1_7_2_n5), .ZN(
        npu_inst_pe_1_7_2_n56) );
  OR3_X1 npu_inst_pe_1_7_2_U27 ( .A1(npu_inst_pe_1_7_2_n5), .A2(
        npu_inst_pe_1_7_2_n8), .A3(npu_inst_pe_1_7_2_n7), .ZN(
        npu_inst_pe_1_7_2_n48) );
  INV_X1 npu_inst_pe_1_7_2_U26 ( .A(npu_inst_pe_1_7_2_n5), .ZN(
        npu_inst_pe_1_7_2_n4) );
  INV_X1 npu_inst_pe_1_7_2_U25 ( .A(npu_inst_n122), .ZN(npu_inst_pe_1_7_2_n12)
         );
  OR3_X1 npu_inst_pe_1_7_2_U24 ( .A1(npu_inst_pe_1_7_2_n4), .A2(
        npu_inst_pe_1_7_2_n8), .A3(npu_inst_pe_1_7_2_n7), .ZN(
        npu_inst_pe_1_7_2_n52) );
  OR3_X1 npu_inst_pe_1_7_2_U23 ( .A1(npu_inst_pe_1_7_2_n6), .A2(
        npu_inst_pe_1_7_2_n8), .A3(npu_inst_pe_1_7_2_n4), .ZN(
        npu_inst_pe_1_7_2_n60) );
  NOR2_X1 npu_inst_pe_1_7_2_U22 ( .A1(npu_inst_pe_1_7_2_n60), .A2(
        npu_inst_pe_1_7_2_n3), .ZN(npu_inst_pe_1_7_2_n58) );
  NOR2_X1 npu_inst_pe_1_7_2_U21 ( .A1(npu_inst_pe_1_7_2_n56), .A2(
        npu_inst_pe_1_7_2_n3), .ZN(npu_inst_pe_1_7_2_n54) );
  NOR2_X1 npu_inst_pe_1_7_2_U20 ( .A1(npu_inst_pe_1_7_2_n52), .A2(
        npu_inst_pe_1_7_2_n3), .ZN(npu_inst_pe_1_7_2_n50) );
  NOR2_X1 npu_inst_pe_1_7_2_U19 ( .A1(npu_inst_pe_1_7_2_n48), .A2(
        npu_inst_pe_1_7_2_n3), .ZN(npu_inst_pe_1_7_2_n46) );
  NOR2_X1 npu_inst_pe_1_7_2_U18 ( .A1(npu_inst_pe_1_7_2_n40), .A2(
        npu_inst_pe_1_7_2_n3), .ZN(npu_inst_pe_1_7_2_n38) );
  NOR2_X1 npu_inst_pe_1_7_2_U17 ( .A1(npu_inst_pe_1_7_2_n44), .A2(
        npu_inst_pe_1_7_2_n3), .ZN(npu_inst_pe_1_7_2_n42) );
  BUF_X1 npu_inst_pe_1_7_2_U16 ( .A(npu_inst_n93), .Z(npu_inst_pe_1_7_2_n8) );
  BUF_X1 npu_inst_pe_1_7_2_U15 ( .A(npu_inst_pe_1_7_2_n12), .Z(
        npu_inst_pe_1_7_2_n11) );
  BUF_X1 npu_inst_pe_1_7_2_U14 ( .A(npu_inst_pe_1_7_2_n12), .Z(
        npu_inst_pe_1_7_2_n10) );
  BUF_X1 npu_inst_pe_1_7_2_U13 ( .A(npu_inst_pe_1_7_2_n12), .Z(
        npu_inst_pe_1_7_2_n9) );
  INV_X1 npu_inst_pe_1_7_2_U12 ( .A(npu_inst_pe_1_7_2_n38), .ZN(
        npu_inst_pe_1_7_2_n118) );
  INV_X1 npu_inst_pe_1_7_2_U11 ( .A(npu_inst_pe_1_7_2_n58), .ZN(
        npu_inst_pe_1_7_2_n114) );
  INV_X1 npu_inst_pe_1_7_2_U10 ( .A(npu_inst_pe_1_7_2_n54), .ZN(
        npu_inst_pe_1_7_2_n115) );
  INV_X1 npu_inst_pe_1_7_2_U9 ( .A(npu_inst_pe_1_7_2_n50), .ZN(
        npu_inst_pe_1_7_2_n116) );
  INV_X1 npu_inst_pe_1_7_2_U8 ( .A(npu_inst_pe_1_7_2_n46), .ZN(
        npu_inst_pe_1_7_2_n117) );
  INV_X1 npu_inst_pe_1_7_2_U7 ( .A(npu_inst_pe_1_7_2_n42), .ZN(
        npu_inst_pe_1_7_2_n119) );
  BUF_X1 npu_inst_pe_1_7_2_U6 ( .A(npu_inst_n9), .Z(npu_inst_pe_1_7_2_n2) );
  BUF_X1 npu_inst_pe_1_7_2_U5 ( .A(npu_inst_n9), .Z(npu_inst_pe_1_7_2_n1) );
  NOR2_X1 npu_inst_pe_1_7_2_U4 ( .A1(npu_inst_pe_1_7_2_int_q_weight_0_), .A2(
        npu_inst_pe_1_7_2_n1), .ZN(npu_inst_pe_1_7_2_n76) );
  NOR2_X1 npu_inst_pe_1_7_2_U3 ( .A1(npu_inst_pe_1_7_2_n27), .A2(
        npu_inst_pe_1_7_2_n1), .ZN(npu_inst_pe_1_7_2_n77) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_7_2_n111), 
        .CK(npu_inst_pe_1_7_2_net2965), .RN(npu_inst_pe_1_7_2_n12), .Q(
        npu_inst_pe_1_7_2_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_7_2_n110), 
        .CK(npu_inst_pe_1_7_2_net2965), .RN(npu_inst_pe_1_7_2_n12), .Q(
        npu_inst_pe_1_7_2_int_q_reg_v_4__1_) );
  FA_X1 npu_inst_pe_1_7_2_sub_77_U2_1 ( .A(npu_inst_pe_1_7_2_int_q_acc_1_), 
        .B(npu_inst_pe_1_7_2_n14), .CI(npu_inst_pe_1_7_2_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_7_2_sub_77_carry_2_), .S(npu_inst_pe_1_7_2_N66) );
  FA_X1 npu_inst_pe_1_7_2_add_79_U1_1 ( .A(npu_inst_pe_1_7_2_int_q_acc_1_), 
        .B(npu_inst_pe_1_7_2_int_data_1_), .CI(
        npu_inst_pe_1_7_2_add_79_carry_1_), .CO(
        npu_inst_pe_1_7_2_add_79_carry_2_), .S(npu_inst_pe_1_7_2_N74) );
  NAND3_X1 npu_inst_pe_1_7_2_U109 ( .A1(npu_inst_pe_1_7_2_n5), .A2(
        npu_inst_pe_1_7_2_n7), .A3(npu_inst_pe_1_7_2_n8), .ZN(
        npu_inst_pe_1_7_2_n44) );
  NAND3_X1 npu_inst_pe_1_7_2_U108 ( .A1(npu_inst_pe_1_7_2_n4), .A2(
        npu_inst_pe_1_7_2_n7), .A3(npu_inst_pe_1_7_2_n8), .ZN(
        npu_inst_pe_1_7_2_n40) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_7_2_n34), .CK(
        npu_inst_pe_1_7_2_net2959), .RN(npu_inst_pe_1_7_2_n9), .Q(
        npu_inst_pe_1_7_2_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_7_2_n35), .CK(
        npu_inst_pe_1_7_2_net2959), .RN(npu_inst_pe_1_7_2_n9), .Q(
        npu_inst_pe_1_7_2_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_7_2_n36), .CK(
        npu_inst_pe_1_7_2_net2959), .RN(npu_inst_pe_1_7_2_n9), .Q(
        npu_inst_pe_1_7_2_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_7_2_n98), .CK(
        npu_inst_pe_1_7_2_net2959), .RN(npu_inst_pe_1_7_2_n9), .Q(
        npu_inst_pe_1_7_2_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_7_2_n99), .CK(
        npu_inst_pe_1_7_2_net2959), .RN(npu_inst_pe_1_7_2_n9), .Q(
        npu_inst_pe_1_7_2_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_7_2_n100), 
        .CK(npu_inst_pe_1_7_2_net2959), .RN(npu_inst_pe_1_7_2_n9), .Q(
        npu_inst_pe_1_7_2_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_7_2_n33), .CK(
        npu_inst_pe_1_7_2_net2959), .RN(npu_inst_pe_1_7_2_n9), .Q(
        npu_inst_pe_1_7_2_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_7_2_n101), 
        .CK(npu_inst_pe_1_7_2_net2959), .RN(npu_inst_pe_1_7_2_n9), .Q(
        npu_inst_pe_1_7_2_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_weight_reg_0_ ( .D(npu_inst_n108), .CK(
        npu_inst_pe_1_7_2_net2965), .RN(npu_inst_pe_1_7_2_n9), .Q(
        npu_inst_pe_1_7_2_int_q_weight_0_), .QN(npu_inst_pe_1_7_2_n27) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_weight_reg_1_ ( .D(npu_inst_n114), .CK(
        npu_inst_pe_1_7_2_net2965), .RN(npu_inst_pe_1_7_2_n9), .Q(
        npu_inst_pe_1_7_2_int_q_weight_1_), .QN(npu_inst_pe_1_7_2_n26) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_7_2_n113), 
        .CK(npu_inst_pe_1_7_2_net2965), .RN(npu_inst_pe_1_7_2_n9), .Q(
        npu_inst_pe_1_7_2_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_7_2_n112), 
        .CK(npu_inst_pe_1_7_2_net2965), .RN(npu_inst_pe_1_7_2_n9), .Q(
        npu_inst_pe_1_7_2_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_7_2_n109), 
        .CK(npu_inst_pe_1_7_2_net2965), .RN(npu_inst_pe_1_7_2_n10), .Q(
        npu_inst_pe_1_7_2_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_7_2_n108), 
        .CK(npu_inst_pe_1_7_2_net2965), .RN(npu_inst_pe_1_7_2_n10), .Q(
        npu_inst_pe_1_7_2_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_7_2_n107), 
        .CK(npu_inst_pe_1_7_2_net2965), .RN(npu_inst_pe_1_7_2_n10), .Q(
        npu_inst_pe_1_7_2_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_7_2_n106), 
        .CK(npu_inst_pe_1_7_2_net2965), .RN(npu_inst_pe_1_7_2_n10), .Q(
        npu_inst_pe_1_7_2_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_7_2_n105), 
        .CK(npu_inst_pe_1_7_2_net2965), .RN(npu_inst_pe_1_7_2_n10), .Q(
        npu_inst_pe_1_7_2_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_7_2_n104), 
        .CK(npu_inst_pe_1_7_2_net2965), .RN(npu_inst_pe_1_7_2_n10), .Q(
        npu_inst_pe_1_7_2_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_7_2_n103), 
        .CK(npu_inst_pe_1_7_2_net2965), .RN(npu_inst_pe_1_7_2_n10), .Q(
        npu_inst_pe_1_7_2_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_7_2_n102), 
        .CK(npu_inst_pe_1_7_2_net2965), .RN(npu_inst_pe_1_7_2_n10), .Q(
        npu_inst_pe_1_7_2_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_7_2_n86), 
        .CK(npu_inst_pe_1_7_2_net2965), .RN(npu_inst_pe_1_7_2_n10), .Q(
        npu_inst_pe_1_7_2_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_7_2_n87), 
        .CK(npu_inst_pe_1_7_2_net2965), .RN(npu_inst_pe_1_7_2_n10), .Q(
        npu_inst_pe_1_7_2_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_7_2_n88), 
        .CK(npu_inst_pe_1_7_2_net2965), .RN(npu_inst_pe_1_7_2_n11), .Q(
        npu_inst_pe_1_7_2_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_7_2_n89), 
        .CK(npu_inst_pe_1_7_2_net2965), .RN(npu_inst_pe_1_7_2_n11), .Q(
        npu_inst_pe_1_7_2_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_7_2_n90), 
        .CK(npu_inst_pe_1_7_2_net2965), .RN(npu_inst_pe_1_7_2_n11), .Q(
        npu_inst_pe_1_7_2_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_7_2_n91), 
        .CK(npu_inst_pe_1_7_2_net2965), .RN(npu_inst_pe_1_7_2_n11), .Q(
        npu_inst_pe_1_7_2_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_7_2_n92), 
        .CK(npu_inst_pe_1_7_2_net2965), .RN(npu_inst_pe_1_7_2_n11), .Q(
        npu_inst_pe_1_7_2_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_7_2_n93), 
        .CK(npu_inst_pe_1_7_2_net2965), .RN(npu_inst_pe_1_7_2_n11), .Q(
        npu_inst_pe_1_7_2_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_7_2_n94), 
        .CK(npu_inst_pe_1_7_2_net2965), .RN(npu_inst_pe_1_7_2_n11), .Q(
        npu_inst_pe_1_7_2_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_7_2_n95), 
        .CK(npu_inst_pe_1_7_2_net2965), .RN(npu_inst_pe_1_7_2_n11), .Q(
        npu_inst_pe_1_7_2_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_7_2_n96), 
        .CK(npu_inst_pe_1_7_2_net2965), .RN(npu_inst_pe_1_7_2_n11), .Q(
        npu_inst_pe_1_7_2_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_7_2_n97), 
        .CK(npu_inst_pe_1_7_2_net2965), .RN(npu_inst_pe_1_7_2_n11), .Q(
        npu_inst_pe_1_7_2_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_7_2_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_7_2_N84), .SE(1'b0), .GCK(npu_inst_pe_1_7_2_net2959) );
  CLKGATETST_X1 npu_inst_pe_1_7_2_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n61), .SE(1'b0), .GCK(npu_inst_pe_1_7_2_net2965) );
  MUX2_X1 npu_inst_pe_1_7_3_U162 ( .A(npu_inst_pe_1_7_3_n32), .B(
        npu_inst_pe_1_7_3_n29), .S(npu_inst_pe_1_7_3_n8), .Z(
        npu_inst_pe_1_7_3_N93) );
  MUX2_X1 npu_inst_pe_1_7_3_U161 ( .A(npu_inst_pe_1_7_3_n31), .B(
        npu_inst_pe_1_7_3_n30), .S(npu_inst_pe_1_7_3_n6), .Z(
        npu_inst_pe_1_7_3_n32) );
  MUX2_X1 npu_inst_pe_1_7_3_U160 ( .A(npu_inst_pe_1_7_3_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_7_3_int_q_reg_v_1__0_), .S(npu_inst_pe_1_7_3_n4), .Z(
        npu_inst_pe_1_7_3_n31) );
  MUX2_X1 npu_inst_pe_1_7_3_U159 ( .A(npu_inst_pe_1_7_3_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_7_3_int_q_reg_v_3__0_), .S(npu_inst_pe_1_7_3_n4), .Z(
        npu_inst_pe_1_7_3_n30) );
  MUX2_X1 npu_inst_pe_1_7_3_U158 ( .A(npu_inst_pe_1_7_3_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_7_3_int_q_reg_v_5__0_), .S(npu_inst_pe_1_7_3_n4), .Z(
        npu_inst_pe_1_7_3_n29) );
  MUX2_X1 npu_inst_pe_1_7_3_U157 ( .A(npu_inst_pe_1_7_3_n28), .B(
        npu_inst_pe_1_7_3_n23), .S(npu_inst_pe_1_7_3_n8), .Z(
        npu_inst_pe_1_7_3_N94) );
  MUX2_X1 npu_inst_pe_1_7_3_U156 ( .A(npu_inst_pe_1_7_3_n25), .B(
        npu_inst_pe_1_7_3_n24), .S(npu_inst_pe_1_7_3_n6), .Z(
        npu_inst_pe_1_7_3_n28) );
  MUX2_X1 npu_inst_pe_1_7_3_U155 ( .A(npu_inst_pe_1_7_3_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_7_3_int_q_reg_v_1__1_), .S(npu_inst_pe_1_7_3_n4), .Z(
        npu_inst_pe_1_7_3_n25) );
  MUX2_X1 npu_inst_pe_1_7_3_U154 ( .A(npu_inst_pe_1_7_3_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_7_3_int_q_reg_v_3__1_), .S(npu_inst_pe_1_7_3_n4), .Z(
        npu_inst_pe_1_7_3_n24) );
  MUX2_X1 npu_inst_pe_1_7_3_U153 ( .A(npu_inst_pe_1_7_3_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_7_3_int_q_reg_v_5__1_), .S(npu_inst_pe_1_7_3_n4), .Z(
        npu_inst_pe_1_7_3_n23) );
  MUX2_X1 npu_inst_pe_1_7_3_U152 ( .A(npu_inst_pe_1_7_3_n22), .B(
        npu_inst_pe_1_7_3_n19), .S(npu_inst_pe_1_7_3_n8), .Z(
        npu_inst_int_data_x_7__3__1_) );
  MUX2_X1 npu_inst_pe_1_7_3_U151 ( .A(npu_inst_pe_1_7_3_n21), .B(
        npu_inst_pe_1_7_3_n20), .S(npu_inst_pe_1_7_3_n6), .Z(
        npu_inst_pe_1_7_3_n22) );
  MUX2_X1 npu_inst_pe_1_7_3_U150 ( .A(npu_inst_pe_1_7_3_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_7_3_int_q_reg_h_1__1_), .S(npu_inst_pe_1_7_3_n4), .Z(
        npu_inst_pe_1_7_3_n21) );
  MUX2_X1 npu_inst_pe_1_7_3_U149 ( .A(npu_inst_pe_1_7_3_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_7_3_int_q_reg_h_3__1_), .S(npu_inst_pe_1_7_3_n4), .Z(
        npu_inst_pe_1_7_3_n20) );
  MUX2_X1 npu_inst_pe_1_7_3_U148 ( .A(npu_inst_pe_1_7_3_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_7_3_int_q_reg_h_5__1_), .S(npu_inst_pe_1_7_3_n4), .Z(
        npu_inst_pe_1_7_3_n19) );
  MUX2_X1 npu_inst_pe_1_7_3_U147 ( .A(npu_inst_pe_1_7_3_n18), .B(
        npu_inst_pe_1_7_3_n15), .S(npu_inst_pe_1_7_3_n8), .Z(
        npu_inst_int_data_x_7__3__0_) );
  MUX2_X1 npu_inst_pe_1_7_3_U146 ( .A(npu_inst_pe_1_7_3_n17), .B(
        npu_inst_pe_1_7_3_n16), .S(npu_inst_pe_1_7_3_n6), .Z(
        npu_inst_pe_1_7_3_n18) );
  MUX2_X1 npu_inst_pe_1_7_3_U145 ( .A(npu_inst_pe_1_7_3_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_7_3_int_q_reg_h_1__0_), .S(npu_inst_pe_1_7_3_n4), .Z(
        npu_inst_pe_1_7_3_n17) );
  MUX2_X1 npu_inst_pe_1_7_3_U144 ( .A(npu_inst_pe_1_7_3_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_7_3_int_q_reg_h_3__0_), .S(npu_inst_pe_1_7_3_n4), .Z(
        npu_inst_pe_1_7_3_n16) );
  MUX2_X1 npu_inst_pe_1_7_3_U143 ( .A(npu_inst_pe_1_7_3_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_7_3_int_q_reg_h_5__0_), .S(npu_inst_pe_1_7_3_n4), .Z(
        npu_inst_pe_1_7_3_n15) );
  XOR2_X1 npu_inst_pe_1_7_3_U142 ( .A(npu_inst_pe_1_7_3_int_data_0_), .B(
        npu_inst_pe_1_7_3_int_q_acc_0_), .Z(npu_inst_pe_1_7_3_N73) );
  AND2_X1 npu_inst_pe_1_7_3_U141 ( .A1(npu_inst_pe_1_7_3_int_q_acc_0_), .A2(
        npu_inst_pe_1_7_3_int_data_0_), .ZN(npu_inst_pe_1_7_3_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_7_3_U140 ( .A(npu_inst_pe_1_7_3_int_q_acc_0_), .B(
        npu_inst_pe_1_7_3_n13), .ZN(npu_inst_pe_1_7_3_N65) );
  OR2_X1 npu_inst_pe_1_7_3_U139 ( .A1(npu_inst_pe_1_7_3_n13), .A2(
        npu_inst_pe_1_7_3_int_q_acc_0_), .ZN(npu_inst_pe_1_7_3_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_7_3_U138 ( .A(npu_inst_pe_1_7_3_int_q_acc_2_), .B(
        npu_inst_pe_1_7_3_add_79_carry_2_), .Z(npu_inst_pe_1_7_3_N75) );
  AND2_X1 npu_inst_pe_1_7_3_U137 ( .A1(npu_inst_pe_1_7_3_add_79_carry_2_), 
        .A2(npu_inst_pe_1_7_3_int_q_acc_2_), .ZN(
        npu_inst_pe_1_7_3_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_7_3_U136 ( .A(npu_inst_pe_1_7_3_int_q_acc_3_), .B(
        npu_inst_pe_1_7_3_add_79_carry_3_), .Z(npu_inst_pe_1_7_3_N76) );
  AND2_X1 npu_inst_pe_1_7_3_U135 ( .A1(npu_inst_pe_1_7_3_add_79_carry_3_), 
        .A2(npu_inst_pe_1_7_3_int_q_acc_3_), .ZN(
        npu_inst_pe_1_7_3_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_7_3_U134 ( .A(npu_inst_pe_1_7_3_int_q_acc_4_), .B(
        npu_inst_pe_1_7_3_add_79_carry_4_), .Z(npu_inst_pe_1_7_3_N77) );
  AND2_X1 npu_inst_pe_1_7_3_U133 ( .A1(npu_inst_pe_1_7_3_add_79_carry_4_), 
        .A2(npu_inst_pe_1_7_3_int_q_acc_4_), .ZN(
        npu_inst_pe_1_7_3_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_7_3_U132 ( .A(npu_inst_pe_1_7_3_int_q_acc_5_), .B(
        npu_inst_pe_1_7_3_add_79_carry_5_), .Z(npu_inst_pe_1_7_3_N78) );
  AND2_X1 npu_inst_pe_1_7_3_U131 ( .A1(npu_inst_pe_1_7_3_add_79_carry_5_), 
        .A2(npu_inst_pe_1_7_3_int_q_acc_5_), .ZN(
        npu_inst_pe_1_7_3_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_7_3_U130 ( .A(npu_inst_pe_1_7_3_int_q_acc_6_), .B(
        npu_inst_pe_1_7_3_add_79_carry_6_), .Z(npu_inst_pe_1_7_3_N79) );
  AND2_X1 npu_inst_pe_1_7_3_U129 ( .A1(npu_inst_pe_1_7_3_add_79_carry_6_), 
        .A2(npu_inst_pe_1_7_3_int_q_acc_6_), .ZN(
        npu_inst_pe_1_7_3_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_7_3_U128 ( .A(npu_inst_pe_1_7_3_int_q_acc_7_), .B(
        npu_inst_pe_1_7_3_add_79_carry_7_), .Z(npu_inst_pe_1_7_3_N80) );
  XNOR2_X1 npu_inst_pe_1_7_3_U127 ( .A(npu_inst_pe_1_7_3_sub_77_carry_2_), .B(
        npu_inst_pe_1_7_3_int_q_acc_2_), .ZN(npu_inst_pe_1_7_3_N67) );
  OR2_X1 npu_inst_pe_1_7_3_U126 ( .A1(npu_inst_pe_1_7_3_int_q_acc_2_), .A2(
        npu_inst_pe_1_7_3_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_7_3_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_7_3_U125 ( .A(npu_inst_pe_1_7_3_sub_77_carry_3_), .B(
        npu_inst_pe_1_7_3_int_q_acc_3_), .ZN(npu_inst_pe_1_7_3_N68) );
  OR2_X1 npu_inst_pe_1_7_3_U124 ( .A1(npu_inst_pe_1_7_3_int_q_acc_3_), .A2(
        npu_inst_pe_1_7_3_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_7_3_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_7_3_U123 ( .A(npu_inst_pe_1_7_3_sub_77_carry_4_), .B(
        npu_inst_pe_1_7_3_int_q_acc_4_), .ZN(npu_inst_pe_1_7_3_N69) );
  OR2_X1 npu_inst_pe_1_7_3_U122 ( .A1(npu_inst_pe_1_7_3_int_q_acc_4_), .A2(
        npu_inst_pe_1_7_3_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_7_3_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_7_3_U121 ( .A(npu_inst_pe_1_7_3_sub_77_carry_5_), .B(
        npu_inst_pe_1_7_3_int_q_acc_5_), .ZN(npu_inst_pe_1_7_3_N70) );
  OR2_X1 npu_inst_pe_1_7_3_U120 ( .A1(npu_inst_pe_1_7_3_int_q_acc_5_), .A2(
        npu_inst_pe_1_7_3_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_7_3_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_7_3_U119 ( .A(npu_inst_pe_1_7_3_sub_77_carry_6_), .B(
        npu_inst_pe_1_7_3_int_q_acc_6_), .ZN(npu_inst_pe_1_7_3_N71) );
  OR2_X1 npu_inst_pe_1_7_3_U118 ( .A1(npu_inst_pe_1_7_3_int_q_acc_6_), .A2(
        npu_inst_pe_1_7_3_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_7_3_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_7_3_U117 ( .A(npu_inst_pe_1_7_3_int_q_acc_7_), .B(
        npu_inst_pe_1_7_3_sub_77_carry_7_), .ZN(npu_inst_pe_1_7_3_N72) );
  INV_X1 npu_inst_pe_1_7_3_U116 ( .A(npu_inst_n75), .ZN(npu_inst_pe_1_7_3_n7)
         );
  INV_X1 npu_inst_pe_1_7_3_U115 ( .A(npu_inst_pe_1_7_3_n7), .ZN(
        npu_inst_pe_1_7_3_n6) );
  INV_X1 npu_inst_pe_1_7_3_U114 ( .A(npu_inst_n52), .ZN(npu_inst_pe_1_7_3_n3)
         );
  AOI22_X1 npu_inst_pe_1_7_3_U113 ( .A1(npu_inst_pe_1_7_3_n38), .A2(
        int_i_data_v_npu[9]), .B1(npu_inst_pe_1_7_3_n118), .B2(
        npu_inst_pe_1_7_3_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_7_3_n39) );
  INV_X1 npu_inst_pe_1_7_3_U112 ( .A(npu_inst_pe_1_7_3_n39), .ZN(
        npu_inst_pe_1_7_3_n112) );
  AOI22_X1 npu_inst_pe_1_7_3_U111 ( .A1(npu_inst_pe_1_7_3_n38), .A2(
        int_i_data_v_npu[8]), .B1(npu_inst_pe_1_7_3_n118), .B2(
        npu_inst_pe_1_7_3_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_7_3_n37) );
  INV_X1 npu_inst_pe_1_7_3_U110 ( .A(npu_inst_pe_1_7_3_n37), .ZN(
        npu_inst_pe_1_7_3_n113) );
  AOI22_X1 npu_inst_pe_1_7_3_U107 ( .A1(int_i_data_v_npu[9]), .A2(
        npu_inst_pe_1_7_3_n58), .B1(npu_inst_pe_1_7_3_n114), .B2(
        npu_inst_pe_1_7_3_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_7_3_n59) );
  INV_X1 npu_inst_pe_1_7_3_U106 ( .A(npu_inst_pe_1_7_3_n59), .ZN(
        npu_inst_pe_1_7_3_n102) );
  AOI22_X1 npu_inst_pe_1_7_3_U105 ( .A1(int_i_data_v_npu[8]), .A2(
        npu_inst_pe_1_7_3_n58), .B1(npu_inst_pe_1_7_3_n114), .B2(
        npu_inst_pe_1_7_3_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_7_3_n57) );
  INV_X1 npu_inst_pe_1_7_3_U104 ( .A(npu_inst_pe_1_7_3_n57), .ZN(
        npu_inst_pe_1_7_3_n103) );
  AOI22_X1 npu_inst_pe_1_7_3_U103 ( .A1(int_i_data_v_npu[9]), .A2(
        npu_inst_pe_1_7_3_n54), .B1(npu_inst_pe_1_7_3_n115), .B2(
        npu_inst_pe_1_7_3_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_7_3_n55) );
  INV_X1 npu_inst_pe_1_7_3_U102 ( .A(npu_inst_pe_1_7_3_n55), .ZN(
        npu_inst_pe_1_7_3_n104) );
  AOI22_X1 npu_inst_pe_1_7_3_U101 ( .A1(int_i_data_v_npu[8]), .A2(
        npu_inst_pe_1_7_3_n54), .B1(npu_inst_pe_1_7_3_n115), .B2(
        npu_inst_pe_1_7_3_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_7_3_n53) );
  INV_X1 npu_inst_pe_1_7_3_U100 ( .A(npu_inst_pe_1_7_3_n53), .ZN(
        npu_inst_pe_1_7_3_n105) );
  AOI22_X1 npu_inst_pe_1_7_3_U99 ( .A1(int_i_data_v_npu[9]), .A2(
        npu_inst_pe_1_7_3_n50), .B1(npu_inst_pe_1_7_3_n116), .B2(
        npu_inst_pe_1_7_3_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_7_3_n51) );
  INV_X1 npu_inst_pe_1_7_3_U98 ( .A(npu_inst_pe_1_7_3_n51), .ZN(
        npu_inst_pe_1_7_3_n106) );
  AOI22_X1 npu_inst_pe_1_7_3_U97 ( .A1(int_i_data_v_npu[8]), .A2(
        npu_inst_pe_1_7_3_n50), .B1(npu_inst_pe_1_7_3_n116), .B2(
        npu_inst_pe_1_7_3_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_7_3_n49) );
  INV_X1 npu_inst_pe_1_7_3_U96 ( .A(npu_inst_pe_1_7_3_n49), .ZN(
        npu_inst_pe_1_7_3_n107) );
  AOI22_X1 npu_inst_pe_1_7_3_U95 ( .A1(int_i_data_v_npu[9]), .A2(
        npu_inst_pe_1_7_3_n46), .B1(npu_inst_pe_1_7_3_n117), .B2(
        npu_inst_pe_1_7_3_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_7_3_n47) );
  INV_X1 npu_inst_pe_1_7_3_U94 ( .A(npu_inst_pe_1_7_3_n47), .ZN(
        npu_inst_pe_1_7_3_n108) );
  AOI22_X1 npu_inst_pe_1_7_3_U93 ( .A1(int_i_data_v_npu[8]), .A2(
        npu_inst_pe_1_7_3_n46), .B1(npu_inst_pe_1_7_3_n117), .B2(
        npu_inst_pe_1_7_3_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_7_3_n45) );
  INV_X1 npu_inst_pe_1_7_3_U92 ( .A(npu_inst_pe_1_7_3_n45), .ZN(
        npu_inst_pe_1_7_3_n109) );
  AOI22_X1 npu_inst_pe_1_7_3_U91 ( .A1(int_i_data_v_npu[9]), .A2(
        npu_inst_pe_1_7_3_n42), .B1(npu_inst_pe_1_7_3_n119), .B2(
        npu_inst_pe_1_7_3_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_7_3_n43) );
  INV_X1 npu_inst_pe_1_7_3_U90 ( .A(npu_inst_pe_1_7_3_n43), .ZN(
        npu_inst_pe_1_7_3_n110) );
  AOI22_X1 npu_inst_pe_1_7_3_U89 ( .A1(int_i_data_v_npu[8]), .A2(
        npu_inst_pe_1_7_3_n42), .B1(npu_inst_pe_1_7_3_n119), .B2(
        npu_inst_pe_1_7_3_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_7_3_n41) );
  INV_X1 npu_inst_pe_1_7_3_U88 ( .A(npu_inst_pe_1_7_3_n41), .ZN(
        npu_inst_pe_1_7_3_n111) );
  NAND2_X1 npu_inst_pe_1_7_3_U87 ( .A1(npu_inst_pe_1_7_3_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_7_3_n60), .ZN(npu_inst_pe_1_7_3_n74) );
  OAI21_X1 npu_inst_pe_1_7_3_U86 ( .B1(npu_inst_pe_1_7_3_n63), .B2(
        npu_inst_pe_1_7_3_n60), .A(npu_inst_pe_1_7_3_n74), .ZN(
        npu_inst_pe_1_7_3_n97) );
  NAND2_X1 npu_inst_pe_1_7_3_U85 ( .A1(npu_inst_pe_1_7_3_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_7_3_n60), .ZN(npu_inst_pe_1_7_3_n73) );
  OAI21_X1 npu_inst_pe_1_7_3_U84 ( .B1(npu_inst_pe_1_7_3_n61), .B2(
        npu_inst_pe_1_7_3_n60), .A(npu_inst_pe_1_7_3_n73), .ZN(
        npu_inst_pe_1_7_3_n96) );
  NAND2_X1 npu_inst_pe_1_7_3_U83 ( .A1(npu_inst_pe_1_7_3_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_7_3_n56), .ZN(npu_inst_pe_1_7_3_n72) );
  OAI21_X1 npu_inst_pe_1_7_3_U82 ( .B1(npu_inst_pe_1_7_3_n63), .B2(
        npu_inst_pe_1_7_3_n56), .A(npu_inst_pe_1_7_3_n72), .ZN(
        npu_inst_pe_1_7_3_n95) );
  NAND2_X1 npu_inst_pe_1_7_3_U81 ( .A1(npu_inst_pe_1_7_3_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_7_3_n56), .ZN(npu_inst_pe_1_7_3_n71) );
  OAI21_X1 npu_inst_pe_1_7_3_U80 ( .B1(npu_inst_pe_1_7_3_n61), .B2(
        npu_inst_pe_1_7_3_n56), .A(npu_inst_pe_1_7_3_n71), .ZN(
        npu_inst_pe_1_7_3_n94) );
  NAND2_X1 npu_inst_pe_1_7_3_U79 ( .A1(npu_inst_pe_1_7_3_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_7_3_n52), .ZN(npu_inst_pe_1_7_3_n70) );
  OAI21_X1 npu_inst_pe_1_7_3_U78 ( .B1(npu_inst_pe_1_7_3_n63), .B2(
        npu_inst_pe_1_7_3_n52), .A(npu_inst_pe_1_7_3_n70), .ZN(
        npu_inst_pe_1_7_3_n93) );
  NAND2_X1 npu_inst_pe_1_7_3_U77 ( .A1(npu_inst_pe_1_7_3_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_7_3_n52), .ZN(npu_inst_pe_1_7_3_n69) );
  OAI21_X1 npu_inst_pe_1_7_3_U76 ( .B1(npu_inst_pe_1_7_3_n61), .B2(
        npu_inst_pe_1_7_3_n52), .A(npu_inst_pe_1_7_3_n69), .ZN(
        npu_inst_pe_1_7_3_n92) );
  NAND2_X1 npu_inst_pe_1_7_3_U75 ( .A1(npu_inst_pe_1_7_3_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_7_3_n48), .ZN(npu_inst_pe_1_7_3_n68) );
  OAI21_X1 npu_inst_pe_1_7_3_U74 ( .B1(npu_inst_pe_1_7_3_n63), .B2(
        npu_inst_pe_1_7_3_n48), .A(npu_inst_pe_1_7_3_n68), .ZN(
        npu_inst_pe_1_7_3_n91) );
  NAND2_X1 npu_inst_pe_1_7_3_U73 ( .A1(npu_inst_pe_1_7_3_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_7_3_n48), .ZN(npu_inst_pe_1_7_3_n67) );
  OAI21_X1 npu_inst_pe_1_7_3_U72 ( .B1(npu_inst_pe_1_7_3_n61), .B2(
        npu_inst_pe_1_7_3_n48), .A(npu_inst_pe_1_7_3_n67), .ZN(
        npu_inst_pe_1_7_3_n90) );
  NAND2_X1 npu_inst_pe_1_7_3_U71 ( .A1(npu_inst_pe_1_7_3_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_7_3_n44), .ZN(npu_inst_pe_1_7_3_n66) );
  OAI21_X1 npu_inst_pe_1_7_3_U70 ( .B1(npu_inst_pe_1_7_3_n63), .B2(
        npu_inst_pe_1_7_3_n44), .A(npu_inst_pe_1_7_3_n66), .ZN(
        npu_inst_pe_1_7_3_n89) );
  NAND2_X1 npu_inst_pe_1_7_3_U69 ( .A1(npu_inst_pe_1_7_3_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_7_3_n44), .ZN(npu_inst_pe_1_7_3_n65) );
  OAI21_X1 npu_inst_pe_1_7_3_U68 ( .B1(npu_inst_pe_1_7_3_n61), .B2(
        npu_inst_pe_1_7_3_n44), .A(npu_inst_pe_1_7_3_n65), .ZN(
        npu_inst_pe_1_7_3_n88) );
  NAND2_X1 npu_inst_pe_1_7_3_U67 ( .A1(npu_inst_pe_1_7_3_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_7_3_n40), .ZN(npu_inst_pe_1_7_3_n64) );
  OAI21_X1 npu_inst_pe_1_7_3_U66 ( .B1(npu_inst_pe_1_7_3_n63), .B2(
        npu_inst_pe_1_7_3_n40), .A(npu_inst_pe_1_7_3_n64), .ZN(
        npu_inst_pe_1_7_3_n87) );
  NAND2_X1 npu_inst_pe_1_7_3_U65 ( .A1(npu_inst_pe_1_7_3_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_7_3_n40), .ZN(npu_inst_pe_1_7_3_n62) );
  OAI21_X1 npu_inst_pe_1_7_3_U64 ( .B1(npu_inst_pe_1_7_3_n61), .B2(
        npu_inst_pe_1_7_3_n40), .A(npu_inst_pe_1_7_3_n62), .ZN(
        npu_inst_pe_1_7_3_n86) );
  AND2_X1 npu_inst_pe_1_7_3_U63 ( .A1(npu_inst_pe_1_7_3_N93), .A2(npu_inst_n52), .ZN(npu_inst_int_data_y_7__3__0_) );
  AND2_X1 npu_inst_pe_1_7_3_U62 ( .A1(npu_inst_n52), .A2(npu_inst_pe_1_7_3_N94), .ZN(npu_inst_int_data_y_7__3__1_) );
  AOI22_X1 npu_inst_pe_1_7_3_U61 ( .A1(npu_inst_n52), .A2(int_i_data_v_npu[9]), 
        .B1(npu_inst_pe_1_7_3_n3), .B2(npu_inst_int_data_x_7__4__1_), .ZN(
        npu_inst_pe_1_7_3_n63) );
  AOI22_X1 npu_inst_pe_1_7_3_U60 ( .A1(npu_inst_n52), .A2(int_i_data_v_npu[8]), 
        .B1(npu_inst_pe_1_7_3_n3), .B2(npu_inst_int_data_x_7__4__0_), .ZN(
        npu_inst_pe_1_7_3_n61) );
  NOR3_X1 npu_inst_pe_1_7_3_U59 ( .A1(npu_inst_pe_1_7_3_n26), .A2(npu_inst_n52), .A3(npu_inst_int_ckg[4]), .ZN(npu_inst_pe_1_7_3_n85) );
  OR2_X1 npu_inst_pe_1_7_3_U58 ( .A1(npu_inst_pe_1_7_3_n85), .A2(
        npu_inst_pe_1_7_3_n2), .ZN(npu_inst_pe_1_7_3_N84) );
  AOI222_X1 npu_inst_pe_1_7_3_U57 ( .A1(1'b0), .A2(npu_inst_pe_1_7_3_n1), .B1(
        npu_inst_pe_1_7_3_N73), .B2(npu_inst_pe_1_7_3_n76), .C1(
        npu_inst_pe_1_7_3_N65), .C2(npu_inst_pe_1_7_3_n77), .ZN(
        npu_inst_pe_1_7_3_n84) );
  INV_X1 npu_inst_pe_1_7_3_U56 ( .A(npu_inst_pe_1_7_3_n84), .ZN(
        npu_inst_pe_1_7_3_n101) );
  AOI222_X1 npu_inst_pe_1_7_3_U55 ( .A1(1'b0), .A2(npu_inst_pe_1_7_3_n1), .B1(
        npu_inst_pe_1_7_3_N80), .B2(npu_inst_pe_1_7_3_n76), .C1(
        npu_inst_pe_1_7_3_N72), .C2(npu_inst_pe_1_7_3_n77), .ZN(
        npu_inst_pe_1_7_3_n75) );
  INV_X1 npu_inst_pe_1_7_3_U54 ( .A(npu_inst_pe_1_7_3_n75), .ZN(
        npu_inst_pe_1_7_3_n33) );
  AOI222_X1 npu_inst_pe_1_7_3_U53 ( .A1(1'b0), .A2(npu_inst_pe_1_7_3_n1), .B1(
        npu_inst_pe_1_7_3_N74), .B2(npu_inst_pe_1_7_3_n76), .C1(
        npu_inst_pe_1_7_3_N66), .C2(npu_inst_pe_1_7_3_n77), .ZN(
        npu_inst_pe_1_7_3_n83) );
  INV_X1 npu_inst_pe_1_7_3_U52 ( .A(npu_inst_pe_1_7_3_n83), .ZN(
        npu_inst_pe_1_7_3_n100) );
  AOI222_X1 npu_inst_pe_1_7_3_U51 ( .A1(1'b0), .A2(npu_inst_pe_1_7_3_n1), .B1(
        npu_inst_pe_1_7_3_N75), .B2(npu_inst_pe_1_7_3_n76), .C1(
        npu_inst_pe_1_7_3_N67), .C2(npu_inst_pe_1_7_3_n77), .ZN(
        npu_inst_pe_1_7_3_n82) );
  INV_X1 npu_inst_pe_1_7_3_U50 ( .A(npu_inst_pe_1_7_3_n82), .ZN(
        npu_inst_pe_1_7_3_n99) );
  AOI222_X1 npu_inst_pe_1_7_3_U49 ( .A1(1'b0), .A2(npu_inst_pe_1_7_3_n1), .B1(
        npu_inst_pe_1_7_3_N76), .B2(npu_inst_pe_1_7_3_n76), .C1(
        npu_inst_pe_1_7_3_N68), .C2(npu_inst_pe_1_7_3_n77), .ZN(
        npu_inst_pe_1_7_3_n81) );
  INV_X1 npu_inst_pe_1_7_3_U48 ( .A(npu_inst_pe_1_7_3_n81), .ZN(
        npu_inst_pe_1_7_3_n98) );
  AOI222_X1 npu_inst_pe_1_7_3_U47 ( .A1(1'b0), .A2(npu_inst_pe_1_7_3_n1), .B1(
        npu_inst_pe_1_7_3_N77), .B2(npu_inst_pe_1_7_3_n76), .C1(
        npu_inst_pe_1_7_3_N69), .C2(npu_inst_pe_1_7_3_n77), .ZN(
        npu_inst_pe_1_7_3_n80) );
  INV_X1 npu_inst_pe_1_7_3_U46 ( .A(npu_inst_pe_1_7_3_n80), .ZN(
        npu_inst_pe_1_7_3_n36) );
  AOI222_X1 npu_inst_pe_1_7_3_U45 ( .A1(1'b0), .A2(npu_inst_pe_1_7_3_n1), .B1(
        npu_inst_pe_1_7_3_N78), .B2(npu_inst_pe_1_7_3_n76), .C1(
        npu_inst_pe_1_7_3_N70), .C2(npu_inst_pe_1_7_3_n77), .ZN(
        npu_inst_pe_1_7_3_n79) );
  INV_X1 npu_inst_pe_1_7_3_U44 ( .A(npu_inst_pe_1_7_3_n79), .ZN(
        npu_inst_pe_1_7_3_n35) );
  AOI222_X1 npu_inst_pe_1_7_3_U43 ( .A1(1'b0), .A2(npu_inst_pe_1_7_3_n1), .B1(
        npu_inst_pe_1_7_3_N79), .B2(npu_inst_pe_1_7_3_n76), .C1(
        npu_inst_pe_1_7_3_N71), .C2(npu_inst_pe_1_7_3_n77), .ZN(
        npu_inst_pe_1_7_3_n78) );
  INV_X1 npu_inst_pe_1_7_3_U42 ( .A(npu_inst_pe_1_7_3_n78), .ZN(
        npu_inst_pe_1_7_3_n34) );
  AND2_X1 npu_inst_pe_1_7_3_U41 ( .A1(npu_inst_pe_1_7_3_int_q_acc_0_), .A2(
        npu_inst_pe_1_7_3_n1), .ZN(npu_inst_int_data_res_7__3__0_) );
  AND2_X1 npu_inst_pe_1_7_3_U40 ( .A1(npu_inst_pe_1_7_3_n2), .A2(
        npu_inst_pe_1_7_3_int_q_acc_7_), .ZN(npu_inst_int_data_res_7__3__7_)
         );
  AND2_X1 npu_inst_pe_1_7_3_U39 ( .A1(npu_inst_pe_1_7_3_int_q_acc_1_), .A2(
        npu_inst_pe_1_7_3_n1), .ZN(npu_inst_int_data_res_7__3__1_) );
  AND2_X1 npu_inst_pe_1_7_3_U38 ( .A1(npu_inst_pe_1_7_3_int_q_acc_2_), .A2(
        npu_inst_pe_1_7_3_n1), .ZN(npu_inst_int_data_res_7__3__2_) );
  AND2_X1 npu_inst_pe_1_7_3_U37 ( .A1(npu_inst_pe_1_7_3_int_q_acc_3_), .A2(
        npu_inst_pe_1_7_3_n2), .ZN(npu_inst_int_data_res_7__3__3_) );
  AND2_X1 npu_inst_pe_1_7_3_U36 ( .A1(npu_inst_pe_1_7_3_int_q_acc_4_), .A2(
        npu_inst_pe_1_7_3_n2), .ZN(npu_inst_int_data_res_7__3__4_) );
  AND2_X1 npu_inst_pe_1_7_3_U35 ( .A1(npu_inst_pe_1_7_3_int_q_acc_5_), .A2(
        npu_inst_pe_1_7_3_n2), .ZN(npu_inst_int_data_res_7__3__5_) );
  AND2_X1 npu_inst_pe_1_7_3_U34 ( .A1(npu_inst_pe_1_7_3_int_q_acc_6_), .A2(
        npu_inst_pe_1_7_3_n2), .ZN(npu_inst_int_data_res_7__3__6_) );
  INV_X1 npu_inst_pe_1_7_3_U33 ( .A(npu_inst_pe_1_7_3_int_data_1_), .ZN(
        npu_inst_pe_1_7_3_n14) );
  AND2_X1 npu_inst_pe_1_7_3_U32 ( .A1(npu_inst_int_data_x_7__3__1_), .A2(
        npu_inst_pe_1_7_3_int_q_weight_1_), .ZN(npu_inst_pe_1_7_3_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_7_3_U31 ( .A1(npu_inst_int_data_x_7__3__0_), .A2(
        npu_inst_pe_1_7_3_int_q_weight_1_), .ZN(npu_inst_pe_1_7_3_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_7_3_U30 ( .A(npu_inst_pe_1_7_3_int_data_0_), .ZN(
        npu_inst_pe_1_7_3_n13) );
  INV_X1 npu_inst_pe_1_7_3_U29 ( .A(npu_inst_n67), .ZN(npu_inst_pe_1_7_3_n5)
         );
  OR3_X1 npu_inst_pe_1_7_3_U28 ( .A1(npu_inst_pe_1_7_3_n6), .A2(
        npu_inst_pe_1_7_3_n8), .A3(npu_inst_pe_1_7_3_n5), .ZN(
        npu_inst_pe_1_7_3_n56) );
  OR3_X1 npu_inst_pe_1_7_3_U27 ( .A1(npu_inst_pe_1_7_3_n5), .A2(
        npu_inst_pe_1_7_3_n8), .A3(npu_inst_pe_1_7_3_n7), .ZN(
        npu_inst_pe_1_7_3_n48) );
  INV_X1 npu_inst_pe_1_7_3_U26 ( .A(npu_inst_pe_1_7_3_n5), .ZN(
        npu_inst_pe_1_7_3_n4) );
  INV_X1 npu_inst_pe_1_7_3_U25 ( .A(npu_inst_n122), .ZN(npu_inst_pe_1_7_3_n12)
         );
  OR3_X1 npu_inst_pe_1_7_3_U24 ( .A1(npu_inst_pe_1_7_3_n4), .A2(
        npu_inst_pe_1_7_3_n8), .A3(npu_inst_pe_1_7_3_n7), .ZN(
        npu_inst_pe_1_7_3_n52) );
  OR3_X1 npu_inst_pe_1_7_3_U23 ( .A1(npu_inst_pe_1_7_3_n6), .A2(
        npu_inst_pe_1_7_3_n8), .A3(npu_inst_pe_1_7_3_n4), .ZN(
        npu_inst_pe_1_7_3_n60) );
  NOR2_X1 npu_inst_pe_1_7_3_U22 ( .A1(npu_inst_pe_1_7_3_n60), .A2(
        npu_inst_pe_1_7_3_n3), .ZN(npu_inst_pe_1_7_3_n58) );
  NOR2_X1 npu_inst_pe_1_7_3_U21 ( .A1(npu_inst_pe_1_7_3_n56), .A2(
        npu_inst_pe_1_7_3_n3), .ZN(npu_inst_pe_1_7_3_n54) );
  NOR2_X1 npu_inst_pe_1_7_3_U20 ( .A1(npu_inst_pe_1_7_3_n52), .A2(
        npu_inst_pe_1_7_3_n3), .ZN(npu_inst_pe_1_7_3_n50) );
  NOR2_X1 npu_inst_pe_1_7_3_U19 ( .A1(npu_inst_pe_1_7_3_n48), .A2(
        npu_inst_pe_1_7_3_n3), .ZN(npu_inst_pe_1_7_3_n46) );
  NOR2_X1 npu_inst_pe_1_7_3_U18 ( .A1(npu_inst_pe_1_7_3_n40), .A2(
        npu_inst_pe_1_7_3_n3), .ZN(npu_inst_pe_1_7_3_n38) );
  NOR2_X1 npu_inst_pe_1_7_3_U17 ( .A1(npu_inst_pe_1_7_3_n44), .A2(
        npu_inst_pe_1_7_3_n3), .ZN(npu_inst_pe_1_7_3_n42) );
  BUF_X1 npu_inst_pe_1_7_3_U16 ( .A(npu_inst_n93), .Z(npu_inst_pe_1_7_3_n8) );
  BUF_X1 npu_inst_pe_1_7_3_U15 ( .A(npu_inst_pe_1_7_3_n12), .Z(
        npu_inst_pe_1_7_3_n11) );
  BUF_X1 npu_inst_pe_1_7_3_U14 ( .A(npu_inst_pe_1_7_3_n12), .Z(
        npu_inst_pe_1_7_3_n10) );
  BUF_X1 npu_inst_pe_1_7_3_U13 ( .A(npu_inst_pe_1_7_3_n12), .Z(
        npu_inst_pe_1_7_3_n9) );
  INV_X1 npu_inst_pe_1_7_3_U12 ( .A(npu_inst_pe_1_7_3_n38), .ZN(
        npu_inst_pe_1_7_3_n118) );
  INV_X1 npu_inst_pe_1_7_3_U11 ( .A(npu_inst_pe_1_7_3_n58), .ZN(
        npu_inst_pe_1_7_3_n114) );
  INV_X1 npu_inst_pe_1_7_3_U10 ( .A(npu_inst_pe_1_7_3_n54), .ZN(
        npu_inst_pe_1_7_3_n115) );
  INV_X1 npu_inst_pe_1_7_3_U9 ( .A(npu_inst_pe_1_7_3_n50), .ZN(
        npu_inst_pe_1_7_3_n116) );
  INV_X1 npu_inst_pe_1_7_3_U8 ( .A(npu_inst_pe_1_7_3_n46), .ZN(
        npu_inst_pe_1_7_3_n117) );
  INV_X1 npu_inst_pe_1_7_3_U7 ( .A(npu_inst_pe_1_7_3_n42), .ZN(
        npu_inst_pe_1_7_3_n119) );
  BUF_X1 npu_inst_pe_1_7_3_U6 ( .A(npu_inst_n9), .Z(npu_inst_pe_1_7_3_n2) );
  BUF_X1 npu_inst_pe_1_7_3_U5 ( .A(npu_inst_n9), .Z(npu_inst_pe_1_7_3_n1) );
  NOR2_X1 npu_inst_pe_1_7_3_U4 ( .A1(npu_inst_pe_1_7_3_int_q_weight_0_), .A2(
        npu_inst_pe_1_7_3_n1), .ZN(npu_inst_pe_1_7_3_n76) );
  NOR2_X1 npu_inst_pe_1_7_3_U3 ( .A1(npu_inst_pe_1_7_3_n27), .A2(
        npu_inst_pe_1_7_3_n1), .ZN(npu_inst_pe_1_7_3_n77) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_7_3_n111), 
        .CK(npu_inst_pe_1_7_3_net2942), .RN(npu_inst_pe_1_7_3_n12), .Q(
        npu_inst_pe_1_7_3_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_7_3_n110), 
        .CK(npu_inst_pe_1_7_3_net2942), .RN(npu_inst_pe_1_7_3_n12), .Q(
        npu_inst_pe_1_7_3_int_q_reg_v_4__1_) );
  FA_X1 npu_inst_pe_1_7_3_sub_77_U2_1 ( .A(npu_inst_pe_1_7_3_int_q_acc_1_), 
        .B(npu_inst_pe_1_7_3_n14), .CI(npu_inst_pe_1_7_3_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_7_3_sub_77_carry_2_), .S(npu_inst_pe_1_7_3_N66) );
  FA_X1 npu_inst_pe_1_7_3_add_79_U1_1 ( .A(npu_inst_pe_1_7_3_int_q_acc_1_), 
        .B(npu_inst_pe_1_7_3_int_data_1_), .CI(
        npu_inst_pe_1_7_3_add_79_carry_1_), .CO(
        npu_inst_pe_1_7_3_add_79_carry_2_), .S(npu_inst_pe_1_7_3_N74) );
  NAND3_X1 npu_inst_pe_1_7_3_U109 ( .A1(npu_inst_pe_1_7_3_n5), .A2(
        npu_inst_pe_1_7_3_n7), .A3(npu_inst_pe_1_7_3_n8), .ZN(
        npu_inst_pe_1_7_3_n44) );
  NAND3_X1 npu_inst_pe_1_7_3_U108 ( .A1(npu_inst_pe_1_7_3_n4), .A2(
        npu_inst_pe_1_7_3_n7), .A3(npu_inst_pe_1_7_3_n8), .ZN(
        npu_inst_pe_1_7_3_n40) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_7_3_n34), .CK(
        npu_inst_pe_1_7_3_net2936), .RN(npu_inst_pe_1_7_3_n9), .Q(
        npu_inst_pe_1_7_3_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_7_3_n35), .CK(
        npu_inst_pe_1_7_3_net2936), .RN(npu_inst_pe_1_7_3_n9), .Q(
        npu_inst_pe_1_7_3_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_7_3_n36), .CK(
        npu_inst_pe_1_7_3_net2936), .RN(npu_inst_pe_1_7_3_n9), .Q(
        npu_inst_pe_1_7_3_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_7_3_n98), .CK(
        npu_inst_pe_1_7_3_net2936), .RN(npu_inst_pe_1_7_3_n9), .Q(
        npu_inst_pe_1_7_3_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_7_3_n99), .CK(
        npu_inst_pe_1_7_3_net2936), .RN(npu_inst_pe_1_7_3_n9), .Q(
        npu_inst_pe_1_7_3_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_7_3_n100), 
        .CK(npu_inst_pe_1_7_3_net2936), .RN(npu_inst_pe_1_7_3_n9), .Q(
        npu_inst_pe_1_7_3_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_7_3_n33), .CK(
        npu_inst_pe_1_7_3_net2936), .RN(npu_inst_pe_1_7_3_n9), .Q(
        npu_inst_pe_1_7_3_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_7_3_n101), 
        .CK(npu_inst_pe_1_7_3_net2936), .RN(npu_inst_pe_1_7_3_n9), .Q(
        npu_inst_pe_1_7_3_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_weight_reg_0_ ( .D(npu_inst_n108), .CK(
        npu_inst_pe_1_7_3_net2942), .RN(npu_inst_pe_1_7_3_n9), .Q(
        npu_inst_pe_1_7_3_int_q_weight_0_), .QN(npu_inst_pe_1_7_3_n27) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_weight_reg_1_ ( .D(npu_inst_n114), .CK(
        npu_inst_pe_1_7_3_net2942), .RN(npu_inst_pe_1_7_3_n9), .Q(
        npu_inst_pe_1_7_3_int_q_weight_1_), .QN(npu_inst_pe_1_7_3_n26) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_7_3_n113), 
        .CK(npu_inst_pe_1_7_3_net2942), .RN(npu_inst_pe_1_7_3_n9), .Q(
        npu_inst_pe_1_7_3_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_7_3_n112), 
        .CK(npu_inst_pe_1_7_3_net2942), .RN(npu_inst_pe_1_7_3_n9), .Q(
        npu_inst_pe_1_7_3_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_7_3_n109), 
        .CK(npu_inst_pe_1_7_3_net2942), .RN(npu_inst_pe_1_7_3_n10), .Q(
        npu_inst_pe_1_7_3_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_7_3_n108), 
        .CK(npu_inst_pe_1_7_3_net2942), .RN(npu_inst_pe_1_7_3_n10), .Q(
        npu_inst_pe_1_7_3_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_7_3_n107), 
        .CK(npu_inst_pe_1_7_3_net2942), .RN(npu_inst_pe_1_7_3_n10), .Q(
        npu_inst_pe_1_7_3_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_7_3_n106), 
        .CK(npu_inst_pe_1_7_3_net2942), .RN(npu_inst_pe_1_7_3_n10), .Q(
        npu_inst_pe_1_7_3_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_7_3_n105), 
        .CK(npu_inst_pe_1_7_3_net2942), .RN(npu_inst_pe_1_7_3_n10), .Q(
        npu_inst_pe_1_7_3_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_7_3_n104), 
        .CK(npu_inst_pe_1_7_3_net2942), .RN(npu_inst_pe_1_7_3_n10), .Q(
        npu_inst_pe_1_7_3_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_7_3_n103), 
        .CK(npu_inst_pe_1_7_3_net2942), .RN(npu_inst_pe_1_7_3_n10), .Q(
        npu_inst_pe_1_7_3_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_7_3_n102), 
        .CK(npu_inst_pe_1_7_3_net2942), .RN(npu_inst_pe_1_7_3_n10), .Q(
        npu_inst_pe_1_7_3_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_7_3_n86), 
        .CK(npu_inst_pe_1_7_3_net2942), .RN(npu_inst_pe_1_7_3_n10), .Q(
        npu_inst_pe_1_7_3_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_7_3_n87), 
        .CK(npu_inst_pe_1_7_3_net2942), .RN(npu_inst_pe_1_7_3_n10), .Q(
        npu_inst_pe_1_7_3_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_7_3_n88), 
        .CK(npu_inst_pe_1_7_3_net2942), .RN(npu_inst_pe_1_7_3_n11), .Q(
        npu_inst_pe_1_7_3_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_7_3_n89), 
        .CK(npu_inst_pe_1_7_3_net2942), .RN(npu_inst_pe_1_7_3_n11), .Q(
        npu_inst_pe_1_7_3_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_7_3_n90), 
        .CK(npu_inst_pe_1_7_3_net2942), .RN(npu_inst_pe_1_7_3_n11), .Q(
        npu_inst_pe_1_7_3_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_7_3_n91), 
        .CK(npu_inst_pe_1_7_3_net2942), .RN(npu_inst_pe_1_7_3_n11), .Q(
        npu_inst_pe_1_7_3_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_7_3_n92), 
        .CK(npu_inst_pe_1_7_3_net2942), .RN(npu_inst_pe_1_7_3_n11), .Q(
        npu_inst_pe_1_7_3_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_7_3_n93), 
        .CK(npu_inst_pe_1_7_3_net2942), .RN(npu_inst_pe_1_7_3_n11), .Q(
        npu_inst_pe_1_7_3_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_7_3_n94), 
        .CK(npu_inst_pe_1_7_3_net2942), .RN(npu_inst_pe_1_7_3_n11), .Q(
        npu_inst_pe_1_7_3_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_7_3_n95), 
        .CK(npu_inst_pe_1_7_3_net2942), .RN(npu_inst_pe_1_7_3_n11), .Q(
        npu_inst_pe_1_7_3_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_7_3_n96), 
        .CK(npu_inst_pe_1_7_3_net2942), .RN(npu_inst_pe_1_7_3_n11), .Q(
        npu_inst_pe_1_7_3_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_7_3_n97), 
        .CK(npu_inst_pe_1_7_3_net2942), .RN(npu_inst_pe_1_7_3_n11), .Q(
        npu_inst_pe_1_7_3_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_7_3_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_7_3_N84), .SE(1'b0), .GCK(npu_inst_pe_1_7_3_net2936) );
  CLKGATETST_X1 npu_inst_pe_1_7_3_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n61), .SE(1'b0), .GCK(npu_inst_pe_1_7_3_net2942) );
  MUX2_X1 npu_inst_pe_1_7_4_U162 ( .A(npu_inst_pe_1_7_4_n32), .B(
        npu_inst_pe_1_7_4_n29), .S(npu_inst_pe_1_7_4_n8), .Z(
        npu_inst_pe_1_7_4_N93) );
  MUX2_X1 npu_inst_pe_1_7_4_U161 ( .A(npu_inst_pe_1_7_4_n31), .B(
        npu_inst_pe_1_7_4_n30), .S(npu_inst_pe_1_7_4_n6), .Z(
        npu_inst_pe_1_7_4_n32) );
  MUX2_X1 npu_inst_pe_1_7_4_U160 ( .A(npu_inst_pe_1_7_4_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_7_4_int_q_reg_v_1__0_), .S(npu_inst_pe_1_7_4_n4), .Z(
        npu_inst_pe_1_7_4_n31) );
  MUX2_X1 npu_inst_pe_1_7_4_U159 ( .A(npu_inst_pe_1_7_4_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_7_4_int_q_reg_v_3__0_), .S(npu_inst_pe_1_7_4_n4), .Z(
        npu_inst_pe_1_7_4_n30) );
  MUX2_X1 npu_inst_pe_1_7_4_U158 ( .A(npu_inst_pe_1_7_4_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_7_4_int_q_reg_v_5__0_), .S(npu_inst_pe_1_7_4_n4), .Z(
        npu_inst_pe_1_7_4_n29) );
  MUX2_X1 npu_inst_pe_1_7_4_U157 ( .A(npu_inst_pe_1_7_4_n28), .B(
        npu_inst_pe_1_7_4_n23), .S(npu_inst_pe_1_7_4_n8), .Z(
        npu_inst_pe_1_7_4_N94) );
  MUX2_X1 npu_inst_pe_1_7_4_U156 ( .A(npu_inst_pe_1_7_4_n25), .B(
        npu_inst_pe_1_7_4_n24), .S(npu_inst_pe_1_7_4_n6), .Z(
        npu_inst_pe_1_7_4_n28) );
  MUX2_X1 npu_inst_pe_1_7_4_U155 ( .A(npu_inst_pe_1_7_4_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_7_4_int_q_reg_v_1__1_), .S(npu_inst_pe_1_7_4_n4), .Z(
        npu_inst_pe_1_7_4_n25) );
  MUX2_X1 npu_inst_pe_1_7_4_U154 ( .A(npu_inst_pe_1_7_4_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_7_4_int_q_reg_v_3__1_), .S(npu_inst_pe_1_7_4_n4), .Z(
        npu_inst_pe_1_7_4_n24) );
  MUX2_X1 npu_inst_pe_1_7_4_U153 ( .A(npu_inst_pe_1_7_4_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_7_4_int_q_reg_v_5__1_), .S(npu_inst_pe_1_7_4_n4), .Z(
        npu_inst_pe_1_7_4_n23) );
  MUX2_X1 npu_inst_pe_1_7_4_U152 ( .A(npu_inst_pe_1_7_4_n22), .B(
        npu_inst_pe_1_7_4_n19), .S(npu_inst_pe_1_7_4_n8), .Z(
        npu_inst_int_data_x_7__4__1_) );
  MUX2_X1 npu_inst_pe_1_7_4_U151 ( .A(npu_inst_pe_1_7_4_n21), .B(
        npu_inst_pe_1_7_4_n20), .S(npu_inst_pe_1_7_4_n6), .Z(
        npu_inst_pe_1_7_4_n22) );
  MUX2_X1 npu_inst_pe_1_7_4_U150 ( .A(npu_inst_pe_1_7_4_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_7_4_int_q_reg_h_1__1_), .S(npu_inst_pe_1_7_4_n4), .Z(
        npu_inst_pe_1_7_4_n21) );
  MUX2_X1 npu_inst_pe_1_7_4_U149 ( .A(npu_inst_pe_1_7_4_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_7_4_int_q_reg_h_3__1_), .S(npu_inst_pe_1_7_4_n4), .Z(
        npu_inst_pe_1_7_4_n20) );
  MUX2_X1 npu_inst_pe_1_7_4_U148 ( .A(npu_inst_pe_1_7_4_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_7_4_int_q_reg_h_5__1_), .S(npu_inst_pe_1_7_4_n4), .Z(
        npu_inst_pe_1_7_4_n19) );
  MUX2_X1 npu_inst_pe_1_7_4_U147 ( .A(npu_inst_pe_1_7_4_n18), .B(
        npu_inst_pe_1_7_4_n15), .S(npu_inst_pe_1_7_4_n8), .Z(
        npu_inst_int_data_x_7__4__0_) );
  MUX2_X1 npu_inst_pe_1_7_4_U146 ( .A(npu_inst_pe_1_7_4_n17), .B(
        npu_inst_pe_1_7_4_n16), .S(npu_inst_pe_1_7_4_n6), .Z(
        npu_inst_pe_1_7_4_n18) );
  MUX2_X1 npu_inst_pe_1_7_4_U145 ( .A(npu_inst_pe_1_7_4_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_7_4_int_q_reg_h_1__0_), .S(npu_inst_pe_1_7_4_n4), .Z(
        npu_inst_pe_1_7_4_n17) );
  MUX2_X1 npu_inst_pe_1_7_4_U144 ( .A(npu_inst_pe_1_7_4_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_7_4_int_q_reg_h_3__0_), .S(npu_inst_pe_1_7_4_n4), .Z(
        npu_inst_pe_1_7_4_n16) );
  MUX2_X1 npu_inst_pe_1_7_4_U143 ( .A(npu_inst_pe_1_7_4_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_7_4_int_q_reg_h_5__0_), .S(npu_inst_pe_1_7_4_n4), .Z(
        npu_inst_pe_1_7_4_n15) );
  XOR2_X1 npu_inst_pe_1_7_4_U142 ( .A(npu_inst_pe_1_7_4_int_data_0_), .B(
        npu_inst_pe_1_7_4_int_q_acc_0_), .Z(npu_inst_pe_1_7_4_N73) );
  AND2_X1 npu_inst_pe_1_7_4_U141 ( .A1(npu_inst_pe_1_7_4_int_q_acc_0_), .A2(
        npu_inst_pe_1_7_4_int_data_0_), .ZN(npu_inst_pe_1_7_4_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_7_4_U140 ( .A(npu_inst_pe_1_7_4_int_q_acc_0_), .B(
        npu_inst_pe_1_7_4_n13), .ZN(npu_inst_pe_1_7_4_N65) );
  OR2_X1 npu_inst_pe_1_7_4_U139 ( .A1(npu_inst_pe_1_7_4_n13), .A2(
        npu_inst_pe_1_7_4_int_q_acc_0_), .ZN(npu_inst_pe_1_7_4_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_7_4_U138 ( .A(npu_inst_pe_1_7_4_int_q_acc_2_), .B(
        npu_inst_pe_1_7_4_add_79_carry_2_), .Z(npu_inst_pe_1_7_4_N75) );
  AND2_X1 npu_inst_pe_1_7_4_U137 ( .A1(npu_inst_pe_1_7_4_add_79_carry_2_), 
        .A2(npu_inst_pe_1_7_4_int_q_acc_2_), .ZN(
        npu_inst_pe_1_7_4_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_7_4_U136 ( .A(npu_inst_pe_1_7_4_int_q_acc_3_), .B(
        npu_inst_pe_1_7_4_add_79_carry_3_), .Z(npu_inst_pe_1_7_4_N76) );
  AND2_X1 npu_inst_pe_1_7_4_U135 ( .A1(npu_inst_pe_1_7_4_add_79_carry_3_), 
        .A2(npu_inst_pe_1_7_4_int_q_acc_3_), .ZN(
        npu_inst_pe_1_7_4_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_7_4_U134 ( .A(npu_inst_pe_1_7_4_int_q_acc_4_), .B(
        npu_inst_pe_1_7_4_add_79_carry_4_), .Z(npu_inst_pe_1_7_4_N77) );
  AND2_X1 npu_inst_pe_1_7_4_U133 ( .A1(npu_inst_pe_1_7_4_add_79_carry_4_), 
        .A2(npu_inst_pe_1_7_4_int_q_acc_4_), .ZN(
        npu_inst_pe_1_7_4_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_7_4_U132 ( .A(npu_inst_pe_1_7_4_int_q_acc_5_), .B(
        npu_inst_pe_1_7_4_add_79_carry_5_), .Z(npu_inst_pe_1_7_4_N78) );
  AND2_X1 npu_inst_pe_1_7_4_U131 ( .A1(npu_inst_pe_1_7_4_add_79_carry_5_), 
        .A2(npu_inst_pe_1_7_4_int_q_acc_5_), .ZN(
        npu_inst_pe_1_7_4_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_7_4_U130 ( .A(npu_inst_pe_1_7_4_int_q_acc_6_), .B(
        npu_inst_pe_1_7_4_add_79_carry_6_), .Z(npu_inst_pe_1_7_4_N79) );
  AND2_X1 npu_inst_pe_1_7_4_U129 ( .A1(npu_inst_pe_1_7_4_add_79_carry_6_), 
        .A2(npu_inst_pe_1_7_4_int_q_acc_6_), .ZN(
        npu_inst_pe_1_7_4_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_7_4_U128 ( .A(npu_inst_pe_1_7_4_int_q_acc_7_), .B(
        npu_inst_pe_1_7_4_add_79_carry_7_), .Z(npu_inst_pe_1_7_4_N80) );
  XNOR2_X1 npu_inst_pe_1_7_4_U127 ( .A(npu_inst_pe_1_7_4_sub_77_carry_2_), .B(
        npu_inst_pe_1_7_4_int_q_acc_2_), .ZN(npu_inst_pe_1_7_4_N67) );
  OR2_X1 npu_inst_pe_1_7_4_U126 ( .A1(npu_inst_pe_1_7_4_int_q_acc_2_), .A2(
        npu_inst_pe_1_7_4_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_7_4_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_7_4_U125 ( .A(npu_inst_pe_1_7_4_sub_77_carry_3_), .B(
        npu_inst_pe_1_7_4_int_q_acc_3_), .ZN(npu_inst_pe_1_7_4_N68) );
  OR2_X1 npu_inst_pe_1_7_4_U124 ( .A1(npu_inst_pe_1_7_4_int_q_acc_3_), .A2(
        npu_inst_pe_1_7_4_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_7_4_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_7_4_U123 ( .A(npu_inst_pe_1_7_4_sub_77_carry_4_), .B(
        npu_inst_pe_1_7_4_int_q_acc_4_), .ZN(npu_inst_pe_1_7_4_N69) );
  OR2_X1 npu_inst_pe_1_7_4_U122 ( .A1(npu_inst_pe_1_7_4_int_q_acc_4_), .A2(
        npu_inst_pe_1_7_4_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_7_4_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_7_4_U121 ( .A(npu_inst_pe_1_7_4_sub_77_carry_5_), .B(
        npu_inst_pe_1_7_4_int_q_acc_5_), .ZN(npu_inst_pe_1_7_4_N70) );
  OR2_X1 npu_inst_pe_1_7_4_U120 ( .A1(npu_inst_pe_1_7_4_int_q_acc_5_), .A2(
        npu_inst_pe_1_7_4_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_7_4_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_7_4_U119 ( .A(npu_inst_pe_1_7_4_sub_77_carry_6_), .B(
        npu_inst_pe_1_7_4_int_q_acc_6_), .ZN(npu_inst_pe_1_7_4_N71) );
  OR2_X1 npu_inst_pe_1_7_4_U118 ( .A1(npu_inst_pe_1_7_4_int_q_acc_6_), .A2(
        npu_inst_pe_1_7_4_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_7_4_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_7_4_U117 ( .A(npu_inst_pe_1_7_4_int_q_acc_7_), .B(
        npu_inst_pe_1_7_4_sub_77_carry_7_), .ZN(npu_inst_pe_1_7_4_N72) );
  INV_X1 npu_inst_pe_1_7_4_U116 ( .A(npu_inst_n75), .ZN(npu_inst_pe_1_7_4_n7)
         );
  INV_X1 npu_inst_pe_1_7_4_U115 ( .A(npu_inst_pe_1_7_4_n7), .ZN(
        npu_inst_pe_1_7_4_n6) );
  INV_X1 npu_inst_pe_1_7_4_U114 ( .A(npu_inst_n52), .ZN(npu_inst_pe_1_7_4_n3)
         );
  AOI22_X1 npu_inst_pe_1_7_4_U113 ( .A1(npu_inst_pe_1_7_4_n38), .A2(
        int_i_data_v_npu[7]), .B1(npu_inst_pe_1_7_4_n118), .B2(
        npu_inst_pe_1_7_4_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_7_4_n39) );
  INV_X1 npu_inst_pe_1_7_4_U112 ( .A(npu_inst_pe_1_7_4_n39), .ZN(
        npu_inst_pe_1_7_4_n112) );
  AOI22_X1 npu_inst_pe_1_7_4_U111 ( .A1(npu_inst_pe_1_7_4_n38), .A2(
        int_i_data_v_npu[6]), .B1(npu_inst_pe_1_7_4_n118), .B2(
        npu_inst_pe_1_7_4_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_7_4_n37) );
  INV_X1 npu_inst_pe_1_7_4_U110 ( .A(npu_inst_pe_1_7_4_n37), .ZN(
        npu_inst_pe_1_7_4_n113) );
  AOI22_X1 npu_inst_pe_1_7_4_U107 ( .A1(int_i_data_v_npu[7]), .A2(
        npu_inst_pe_1_7_4_n58), .B1(npu_inst_pe_1_7_4_n114), .B2(
        npu_inst_pe_1_7_4_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_7_4_n59) );
  INV_X1 npu_inst_pe_1_7_4_U106 ( .A(npu_inst_pe_1_7_4_n59), .ZN(
        npu_inst_pe_1_7_4_n102) );
  AOI22_X1 npu_inst_pe_1_7_4_U105 ( .A1(int_i_data_v_npu[6]), .A2(
        npu_inst_pe_1_7_4_n58), .B1(npu_inst_pe_1_7_4_n114), .B2(
        npu_inst_pe_1_7_4_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_7_4_n57) );
  INV_X1 npu_inst_pe_1_7_4_U104 ( .A(npu_inst_pe_1_7_4_n57), .ZN(
        npu_inst_pe_1_7_4_n103) );
  AOI22_X1 npu_inst_pe_1_7_4_U103 ( .A1(int_i_data_v_npu[7]), .A2(
        npu_inst_pe_1_7_4_n54), .B1(npu_inst_pe_1_7_4_n115), .B2(
        npu_inst_pe_1_7_4_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_7_4_n55) );
  INV_X1 npu_inst_pe_1_7_4_U102 ( .A(npu_inst_pe_1_7_4_n55), .ZN(
        npu_inst_pe_1_7_4_n104) );
  AOI22_X1 npu_inst_pe_1_7_4_U101 ( .A1(int_i_data_v_npu[6]), .A2(
        npu_inst_pe_1_7_4_n54), .B1(npu_inst_pe_1_7_4_n115), .B2(
        npu_inst_pe_1_7_4_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_7_4_n53) );
  INV_X1 npu_inst_pe_1_7_4_U100 ( .A(npu_inst_pe_1_7_4_n53), .ZN(
        npu_inst_pe_1_7_4_n105) );
  AOI22_X1 npu_inst_pe_1_7_4_U99 ( .A1(int_i_data_v_npu[7]), .A2(
        npu_inst_pe_1_7_4_n50), .B1(npu_inst_pe_1_7_4_n116), .B2(
        npu_inst_pe_1_7_4_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_7_4_n51) );
  INV_X1 npu_inst_pe_1_7_4_U98 ( .A(npu_inst_pe_1_7_4_n51), .ZN(
        npu_inst_pe_1_7_4_n106) );
  AOI22_X1 npu_inst_pe_1_7_4_U97 ( .A1(int_i_data_v_npu[6]), .A2(
        npu_inst_pe_1_7_4_n50), .B1(npu_inst_pe_1_7_4_n116), .B2(
        npu_inst_pe_1_7_4_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_7_4_n49) );
  INV_X1 npu_inst_pe_1_7_4_U96 ( .A(npu_inst_pe_1_7_4_n49), .ZN(
        npu_inst_pe_1_7_4_n107) );
  AOI22_X1 npu_inst_pe_1_7_4_U95 ( .A1(int_i_data_v_npu[7]), .A2(
        npu_inst_pe_1_7_4_n46), .B1(npu_inst_pe_1_7_4_n117), .B2(
        npu_inst_pe_1_7_4_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_7_4_n47) );
  INV_X1 npu_inst_pe_1_7_4_U94 ( .A(npu_inst_pe_1_7_4_n47), .ZN(
        npu_inst_pe_1_7_4_n108) );
  AOI22_X1 npu_inst_pe_1_7_4_U93 ( .A1(int_i_data_v_npu[6]), .A2(
        npu_inst_pe_1_7_4_n46), .B1(npu_inst_pe_1_7_4_n117), .B2(
        npu_inst_pe_1_7_4_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_7_4_n45) );
  INV_X1 npu_inst_pe_1_7_4_U92 ( .A(npu_inst_pe_1_7_4_n45), .ZN(
        npu_inst_pe_1_7_4_n109) );
  AOI22_X1 npu_inst_pe_1_7_4_U91 ( .A1(int_i_data_v_npu[7]), .A2(
        npu_inst_pe_1_7_4_n42), .B1(npu_inst_pe_1_7_4_n119), .B2(
        npu_inst_pe_1_7_4_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_7_4_n43) );
  INV_X1 npu_inst_pe_1_7_4_U90 ( .A(npu_inst_pe_1_7_4_n43), .ZN(
        npu_inst_pe_1_7_4_n110) );
  AOI22_X1 npu_inst_pe_1_7_4_U89 ( .A1(int_i_data_v_npu[6]), .A2(
        npu_inst_pe_1_7_4_n42), .B1(npu_inst_pe_1_7_4_n119), .B2(
        npu_inst_pe_1_7_4_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_7_4_n41) );
  INV_X1 npu_inst_pe_1_7_4_U88 ( .A(npu_inst_pe_1_7_4_n41), .ZN(
        npu_inst_pe_1_7_4_n111) );
  NAND2_X1 npu_inst_pe_1_7_4_U87 ( .A1(npu_inst_pe_1_7_4_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_7_4_n60), .ZN(npu_inst_pe_1_7_4_n74) );
  OAI21_X1 npu_inst_pe_1_7_4_U86 ( .B1(npu_inst_pe_1_7_4_n63), .B2(
        npu_inst_pe_1_7_4_n60), .A(npu_inst_pe_1_7_4_n74), .ZN(
        npu_inst_pe_1_7_4_n97) );
  NAND2_X1 npu_inst_pe_1_7_4_U85 ( .A1(npu_inst_pe_1_7_4_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_7_4_n60), .ZN(npu_inst_pe_1_7_4_n73) );
  OAI21_X1 npu_inst_pe_1_7_4_U84 ( .B1(npu_inst_pe_1_7_4_n61), .B2(
        npu_inst_pe_1_7_4_n60), .A(npu_inst_pe_1_7_4_n73), .ZN(
        npu_inst_pe_1_7_4_n96) );
  NAND2_X1 npu_inst_pe_1_7_4_U83 ( .A1(npu_inst_pe_1_7_4_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_7_4_n56), .ZN(npu_inst_pe_1_7_4_n72) );
  OAI21_X1 npu_inst_pe_1_7_4_U82 ( .B1(npu_inst_pe_1_7_4_n63), .B2(
        npu_inst_pe_1_7_4_n56), .A(npu_inst_pe_1_7_4_n72), .ZN(
        npu_inst_pe_1_7_4_n95) );
  NAND2_X1 npu_inst_pe_1_7_4_U81 ( .A1(npu_inst_pe_1_7_4_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_7_4_n56), .ZN(npu_inst_pe_1_7_4_n71) );
  OAI21_X1 npu_inst_pe_1_7_4_U80 ( .B1(npu_inst_pe_1_7_4_n61), .B2(
        npu_inst_pe_1_7_4_n56), .A(npu_inst_pe_1_7_4_n71), .ZN(
        npu_inst_pe_1_7_4_n94) );
  NAND2_X1 npu_inst_pe_1_7_4_U79 ( .A1(npu_inst_pe_1_7_4_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_7_4_n52), .ZN(npu_inst_pe_1_7_4_n70) );
  OAI21_X1 npu_inst_pe_1_7_4_U78 ( .B1(npu_inst_pe_1_7_4_n63), .B2(
        npu_inst_pe_1_7_4_n52), .A(npu_inst_pe_1_7_4_n70), .ZN(
        npu_inst_pe_1_7_4_n93) );
  NAND2_X1 npu_inst_pe_1_7_4_U77 ( .A1(npu_inst_pe_1_7_4_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_7_4_n52), .ZN(npu_inst_pe_1_7_4_n69) );
  OAI21_X1 npu_inst_pe_1_7_4_U76 ( .B1(npu_inst_pe_1_7_4_n61), .B2(
        npu_inst_pe_1_7_4_n52), .A(npu_inst_pe_1_7_4_n69), .ZN(
        npu_inst_pe_1_7_4_n92) );
  NAND2_X1 npu_inst_pe_1_7_4_U75 ( .A1(npu_inst_pe_1_7_4_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_7_4_n48), .ZN(npu_inst_pe_1_7_4_n68) );
  OAI21_X1 npu_inst_pe_1_7_4_U74 ( .B1(npu_inst_pe_1_7_4_n63), .B2(
        npu_inst_pe_1_7_4_n48), .A(npu_inst_pe_1_7_4_n68), .ZN(
        npu_inst_pe_1_7_4_n91) );
  NAND2_X1 npu_inst_pe_1_7_4_U73 ( .A1(npu_inst_pe_1_7_4_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_7_4_n48), .ZN(npu_inst_pe_1_7_4_n67) );
  OAI21_X1 npu_inst_pe_1_7_4_U72 ( .B1(npu_inst_pe_1_7_4_n61), .B2(
        npu_inst_pe_1_7_4_n48), .A(npu_inst_pe_1_7_4_n67), .ZN(
        npu_inst_pe_1_7_4_n90) );
  NAND2_X1 npu_inst_pe_1_7_4_U71 ( .A1(npu_inst_pe_1_7_4_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_7_4_n44), .ZN(npu_inst_pe_1_7_4_n66) );
  OAI21_X1 npu_inst_pe_1_7_4_U70 ( .B1(npu_inst_pe_1_7_4_n63), .B2(
        npu_inst_pe_1_7_4_n44), .A(npu_inst_pe_1_7_4_n66), .ZN(
        npu_inst_pe_1_7_4_n89) );
  NAND2_X1 npu_inst_pe_1_7_4_U69 ( .A1(npu_inst_pe_1_7_4_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_7_4_n44), .ZN(npu_inst_pe_1_7_4_n65) );
  OAI21_X1 npu_inst_pe_1_7_4_U68 ( .B1(npu_inst_pe_1_7_4_n61), .B2(
        npu_inst_pe_1_7_4_n44), .A(npu_inst_pe_1_7_4_n65), .ZN(
        npu_inst_pe_1_7_4_n88) );
  NAND2_X1 npu_inst_pe_1_7_4_U67 ( .A1(npu_inst_pe_1_7_4_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_7_4_n40), .ZN(npu_inst_pe_1_7_4_n64) );
  OAI21_X1 npu_inst_pe_1_7_4_U66 ( .B1(npu_inst_pe_1_7_4_n63), .B2(
        npu_inst_pe_1_7_4_n40), .A(npu_inst_pe_1_7_4_n64), .ZN(
        npu_inst_pe_1_7_4_n87) );
  NAND2_X1 npu_inst_pe_1_7_4_U65 ( .A1(npu_inst_pe_1_7_4_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_7_4_n40), .ZN(npu_inst_pe_1_7_4_n62) );
  OAI21_X1 npu_inst_pe_1_7_4_U64 ( .B1(npu_inst_pe_1_7_4_n61), .B2(
        npu_inst_pe_1_7_4_n40), .A(npu_inst_pe_1_7_4_n62), .ZN(
        npu_inst_pe_1_7_4_n86) );
  AND2_X1 npu_inst_pe_1_7_4_U63 ( .A1(npu_inst_pe_1_7_4_N93), .A2(npu_inst_n52), .ZN(npu_inst_int_data_y_7__4__0_) );
  AND2_X1 npu_inst_pe_1_7_4_U62 ( .A1(npu_inst_n52), .A2(npu_inst_pe_1_7_4_N94), .ZN(npu_inst_int_data_y_7__4__1_) );
  AOI22_X1 npu_inst_pe_1_7_4_U61 ( .A1(npu_inst_n52), .A2(int_i_data_v_npu[7]), 
        .B1(npu_inst_pe_1_7_4_n3), .B2(npu_inst_int_data_x_7__5__1_), .ZN(
        npu_inst_pe_1_7_4_n63) );
  AOI22_X1 npu_inst_pe_1_7_4_U60 ( .A1(npu_inst_n52), .A2(int_i_data_v_npu[6]), 
        .B1(npu_inst_pe_1_7_4_n3), .B2(npu_inst_int_data_x_7__5__0_), .ZN(
        npu_inst_pe_1_7_4_n61) );
  NOR3_X1 npu_inst_pe_1_7_4_U59 ( .A1(npu_inst_pe_1_7_4_n26), .A2(npu_inst_n52), .A3(npu_inst_int_ckg[3]), .ZN(npu_inst_pe_1_7_4_n85) );
  OR2_X1 npu_inst_pe_1_7_4_U58 ( .A1(npu_inst_pe_1_7_4_n85), .A2(
        npu_inst_pe_1_7_4_n2), .ZN(npu_inst_pe_1_7_4_N84) );
  AOI222_X1 npu_inst_pe_1_7_4_U57 ( .A1(1'b0), .A2(npu_inst_pe_1_7_4_n1), .B1(
        npu_inst_pe_1_7_4_N73), .B2(npu_inst_pe_1_7_4_n76), .C1(
        npu_inst_pe_1_7_4_N65), .C2(npu_inst_pe_1_7_4_n77), .ZN(
        npu_inst_pe_1_7_4_n84) );
  INV_X1 npu_inst_pe_1_7_4_U56 ( .A(npu_inst_pe_1_7_4_n84), .ZN(
        npu_inst_pe_1_7_4_n101) );
  AOI222_X1 npu_inst_pe_1_7_4_U55 ( .A1(1'b0), .A2(npu_inst_pe_1_7_4_n1), .B1(
        npu_inst_pe_1_7_4_N80), .B2(npu_inst_pe_1_7_4_n76), .C1(
        npu_inst_pe_1_7_4_N72), .C2(npu_inst_pe_1_7_4_n77), .ZN(
        npu_inst_pe_1_7_4_n75) );
  INV_X1 npu_inst_pe_1_7_4_U54 ( .A(npu_inst_pe_1_7_4_n75), .ZN(
        npu_inst_pe_1_7_4_n33) );
  AOI222_X1 npu_inst_pe_1_7_4_U53 ( .A1(1'b0), .A2(npu_inst_pe_1_7_4_n1), .B1(
        npu_inst_pe_1_7_4_N74), .B2(npu_inst_pe_1_7_4_n76), .C1(
        npu_inst_pe_1_7_4_N66), .C2(npu_inst_pe_1_7_4_n77), .ZN(
        npu_inst_pe_1_7_4_n83) );
  INV_X1 npu_inst_pe_1_7_4_U52 ( .A(npu_inst_pe_1_7_4_n83), .ZN(
        npu_inst_pe_1_7_4_n100) );
  AOI222_X1 npu_inst_pe_1_7_4_U51 ( .A1(1'b0), .A2(npu_inst_pe_1_7_4_n1), .B1(
        npu_inst_pe_1_7_4_N75), .B2(npu_inst_pe_1_7_4_n76), .C1(
        npu_inst_pe_1_7_4_N67), .C2(npu_inst_pe_1_7_4_n77), .ZN(
        npu_inst_pe_1_7_4_n82) );
  INV_X1 npu_inst_pe_1_7_4_U50 ( .A(npu_inst_pe_1_7_4_n82), .ZN(
        npu_inst_pe_1_7_4_n99) );
  AOI222_X1 npu_inst_pe_1_7_4_U49 ( .A1(1'b0), .A2(npu_inst_pe_1_7_4_n1), .B1(
        npu_inst_pe_1_7_4_N76), .B2(npu_inst_pe_1_7_4_n76), .C1(
        npu_inst_pe_1_7_4_N68), .C2(npu_inst_pe_1_7_4_n77), .ZN(
        npu_inst_pe_1_7_4_n81) );
  INV_X1 npu_inst_pe_1_7_4_U48 ( .A(npu_inst_pe_1_7_4_n81), .ZN(
        npu_inst_pe_1_7_4_n98) );
  AOI222_X1 npu_inst_pe_1_7_4_U47 ( .A1(1'b0), .A2(npu_inst_pe_1_7_4_n1), .B1(
        npu_inst_pe_1_7_4_N77), .B2(npu_inst_pe_1_7_4_n76), .C1(
        npu_inst_pe_1_7_4_N69), .C2(npu_inst_pe_1_7_4_n77), .ZN(
        npu_inst_pe_1_7_4_n80) );
  INV_X1 npu_inst_pe_1_7_4_U46 ( .A(npu_inst_pe_1_7_4_n80), .ZN(
        npu_inst_pe_1_7_4_n36) );
  AOI222_X1 npu_inst_pe_1_7_4_U45 ( .A1(1'b0), .A2(npu_inst_pe_1_7_4_n1), .B1(
        npu_inst_pe_1_7_4_N78), .B2(npu_inst_pe_1_7_4_n76), .C1(
        npu_inst_pe_1_7_4_N70), .C2(npu_inst_pe_1_7_4_n77), .ZN(
        npu_inst_pe_1_7_4_n79) );
  INV_X1 npu_inst_pe_1_7_4_U44 ( .A(npu_inst_pe_1_7_4_n79), .ZN(
        npu_inst_pe_1_7_4_n35) );
  AOI222_X1 npu_inst_pe_1_7_4_U43 ( .A1(1'b0), .A2(npu_inst_pe_1_7_4_n1), .B1(
        npu_inst_pe_1_7_4_N79), .B2(npu_inst_pe_1_7_4_n76), .C1(
        npu_inst_pe_1_7_4_N71), .C2(npu_inst_pe_1_7_4_n77), .ZN(
        npu_inst_pe_1_7_4_n78) );
  INV_X1 npu_inst_pe_1_7_4_U42 ( .A(npu_inst_pe_1_7_4_n78), .ZN(
        npu_inst_pe_1_7_4_n34) );
  AND2_X1 npu_inst_pe_1_7_4_U41 ( .A1(npu_inst_pe_1_7_4_int_q_acc_0_), .A2(
        npu_inst_pe_1_7_4_n1), .ZN(npu_inst_int_data_res_7__4__0_) );
  AND2_X1 npu_inst_pe_1_7_4_U40 ( .A1(npu_inst_pe_1_7_4_n2), .A2(
        npu_inst_pe_1_7_4_int_q_acc_7_), .ZN(npu_inst_int_data_res_7__4__7_)
         );
  AND2_X1 npu_inst_pe_1_7_4_U39 ( .A1(npu_inst_pe_1_7_4_int_q_acc_1_), .A2(
        npu_inst_pe_1_7_4_n1), .ZN(npu_inst_int_data_res_7__4__1_) );
  AND2_X1 npu_inst_pe_1_7_4_U38 ( .A1(npu_inst_pe_1_7_4_int_q_acc_2_), .A2(
        npu_inst_pe_1_7_4_n1), .ZN(npu_inst_int_data_res_7__4__2_) );
  AND2_X1 npu_inst_pe_1_7_4_U37 ( .A1(npu_inst_pe_1_7_4_int_q_acc_3_), .A2(
        npu_inst_pe_1_7_4_n2), .ZN(npu_inst_int_data_res_7__4__3_) );
  AND2_X1 npu_inst_pe_1_7_4_U36 ( .A1(npu_inst_pe_1_7_4_int_q_acc_4_), .A2(
        npu_inst_pe_1_7_4_n2), .ZN(npu_inst_int_data_res_7__4__4_) );
  AND2_X1 npu_inst_pe_1_7_4_U35 ( .A1(npu_inst_pe_1_7_4_int_q_acc_5_), .A2(
        npu_inst_pe_1_7_4_n2), .ZN(npu_inst_int_data_res_7__4__5_) );
  AND2_X1 npu_inst_pe_1_7_4_U34 ( .A1(npu_inst_pe_1_7_4_int_q_acc_6_), .A2(
        npu_inst_pe_1_7_4_n2), .ZN(npu_inst_int_data_res_7__4__6_) );
  INV_X1 npu_inst_pe_1_7_4_U33 ( .A(npu_inst_pe_1_7_4_int_data_1_), .ZN(
        npu_inst_pe_1_7_4_n14) );
  AND2_X1 npu_inst_pe_1_7_4_U32 ( .A1(npu_inst_int_data_x_7__4__1_), .A2(
        npu_inst_pe_1_7_4_int_q_weight_1_), .ZN(npu_inst_pe_1_7_4_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_7_4_U31 ( .A1(npu_inst_int_data_x_7__4__0_), .A2(
        npu_inst_pe_1_7_4_int_q_weight_1_), .ZN(npu_inst_pe_1_7_4_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_7_4_U30 ( .A(npu_inst_pe_1_7_4_int_data_0_), .ZN(
        npu_inst_pe_1_7_4_n13) );
  INV_X1 npu_inst_pe_1_7_4_U29 ( .A(npu_inst_n67), .ZN(npu_inst_pe_1_7_4_n5)
         );
  OR3_X1 npu_inst_pe_1_7_4_U28 ( .A1(npu_inst_pe_1_7_4_n6), .A2(
        npu_inst_pe_1_7_4_n8), .A3(npu_inst_pe_1_7_4_n5), .ZN(
        npu_inst_pe_1_7_4_n56) );
  OR3_X1 npu_inst_pe_1_7_4_U27 ( .A1(npu_inst_pe_1_7_4_n5), .A2(
        npu_inst_pe_1_7_4_n8), .A3(npu_inst_pe_1_7_4_n7), .ZN(
        npu_inst_pe_1_7_4_n48) );
  INV_X1 npu_inst_pe_1_7_4_U26 ( .A(npu_inst_pe_1_7_4_n5), .ZN(
        npu_inst_pe_1_7_4_n4) );
  INV_X1 npu_inst_pe_1_7_4_U25 ( .A(npu_inst_n122), .ZN(npu_inst_pe_1_7_4_n12)
         );
  OR3_X1 npu_inst_pe_1_7_4_U24 ( .A1(npu_inst_pe_1_7_4_n4), .A2(
        npu_inst_pe_1_7_4_n8), .A3(npu_inst_pe_1_7_4_n7), .ZN(
        npu_inst_pe_1_7_4_n52) );
  OR3_X1 npu_inst_pe_1_7_4_U23 ( .A1(npu_inst_pe_1_7_4_n6), .A2(
        npu_inst_pe_1_7_4_n8), .A3(npu_inst_pe_1_7_4_n4), .ZN(
        npu_inst_pe_1_7_4_n60) );
  NOR2_X1 npu_inst_pe_1_7_4_U22 ( .A1(npu_inst_pe_1_7_4_n60), .A2(
        npu_inst_pe_1_7_4_n3), .ZN(npu_inst_pe_1_7_4_n58) );
  NOR2_X1 npu_inst_pe_1_7_4_U21 ( .A1(npu_inst_pe_1_7_4_n56), .A2(
        npu_inst_pe_1_7_4_n3), .ZN(npu_inst_pe_1_7_4_n54) );
  NOR2_X1 npu_inst_pe_1_7_4_U20 ( .A1(npu_inst_pe_1_7_4_n52), .A2(
        npu_inst_pe_1_7_4_n3), .ZN(npu_inst_pe_1_7_4_n50) );
  NOR2_X1 npu_inst_pe_1_7_4_U19 ( .A1(npu_inst_pe_1_7_4_n48), .A2(
        npu_inst_pe_1_7_4_n3), .ZN(npu_inst_pe_1_7_4_n46) );
  NOR2_X1 npu_inst_pe_1_7_4_U18 ( .A1(npu_inst_pe_1_7_4_n40), .A2(
        npu_inst_pe_1_7_4_n3), .ZN(npu_inst_pe_1_7_4_n38) );
  NOR2_X1 npu_inst_pe_1_7_4_U17 ( .A1(npu_inst_pe_1_7_4_n44), .A2(
        npu_inst_pe_1_7_4_n3), .ZN(npu_inst_pe_1_7_4_n42) );
  BUF_X1 npu_inst_pe_1_7_4_U16 ( .A(npu_inst_n92), .Z(npu_inst_pe_1_7_4_n8) );
  BUF_X1 npu_inst_pe_1_7_4_U15 ( .A(npu_inst_pe_1_7_4_n12), .Z(
        npu_inst_pe_1_7_4_n11) );
  BUF_X1 npu_inst_pe_1_7_4_U14 ( .A(npu_inst_pe_1_7_4_n12), .Z(
        npu_inst_pe_1_7_4_n10) );
  BUF_X1 npu_inst_pe_1_7_4_U13 ( .A(npu_inst_pe_1_7_4_n12), .Z(
        npu_inst_pe_1_7_4_n9) );
  INV_X1 npu_inst_pe_1_7_4_U12 ( .A(npu_inst_pe_1_7_4_n38), .ZN(
        npu_inst_pe_1_7_4_n118) );
  INV_X1 npu_inst_pe_1_7_4_U11 ( .A(npu_inst_pe_1_7_4_n58), .ZN(
        npu_inst_pe_1_7_4_n114) );
  INV_X1 npu_inst_pe_1_7_4_U10 ( .A(npu_inst_pe_1_7_4_n54), .ZN(
        npu_inst_pe_1_7_4_n115) );
  INV_X1 npu_inst_pe_1_7_4_U9 ( .A(npu_inst_pe_1_7_4_n50), .ZN(
        npu_inst_pe_1_7_4_n116) );
  INV_X1 npu_inst_pe_1_7_4_U8 ( .A(npu_inst_pe_1_7_4_n46), .ZN(
        npu_inst_pe_1_7_4_n117) );
  INV_X1 npu_inst_pe_1_7_4_U7 ( .A(npu_inst_pe_1_7_4_n42), .ZN(
        npu_inst_pe_1_7_4_n119) );
  BUF_X1 npu_inst_pe_1_7_4_U6 ( .A(npu_inst_n8), .Z(npu_inst_pe_1_7_4_n2) );
  BUF_X1 npu_inst_pe_1_7_4_U5 ( .A(npu_inst_n8), .Z(npu_inst_pe_1_7_4_n1) );
  NOR2_X1 npu_inst_pe_1_7_4_U4 ( .A1(npu_inst_pe_1_7_4_int_q_weight_0_), .A2(
        npu_inst_pe_1_7_4_n1), .ZN(npu_inst_pe_1_7_4_n76) );
  NOR2_X1 npu_inst_pe_1_7_4_U3 ( .A1(npu_inst_pe_1_7_4_n27), .A2(
        npu_inst_pe_1_7_4_n1), .ZN(npu_inst_pe_1_7_4_n77) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_7_4_n111), 
        .CK(npu_inst_pe_1_7_4_net2919), .RN(npu_inst_pe_1_7_4_n12), .Q(
        npu_inst_pe_1_7_4_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_7_4_n110), 
        .CK(npu_inst_pe_1_7_4_net2919), .RN(npu_inst_pe_1_7_4_n12), .Q(
        npu_inst_pe_1_7_4_int_q_reg_v_4__1_) );
  FA_X1 npu_inst_pe_1_7_4_sub_77_U2_1 ( .A(npu_inst_pe_1_7_4_int_q_acc_1_), 
        .B(npu_inst_pe_1_7_4_n14), .CI(npu_inst_pe_1_7_4_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_7_4_sub_77_carry_2_), .S(npu_inst_pe_1_7_4_N66) );
  FA_X1 npu_inst_pe_1_7_4_add_79_U1_1 ( .A(npu_inst_pe_1_7_4_int_q_acc_1_), 
        .B(npu_inst_pe_1_7_4_int_data_1_), .CI(
        npu_inst_pe_1_7_4_add_79_carry_1_), .CO(
        npu_inst_pe_1_7_4_add_79_carry_2_), .S(npu_inst_pe_1_7_4_N74) );
  NAND3_X1 npu_inst_pe_1_7_4_U109 ( .A1(npu_inst_pe_1_7_4_n5), .A2(
        npu_inst_pe_1_7_4_n7), .A3(npu_inst_pe_1_7_4_n8), .ZN(
        npu_inst_pe_1_7_4_n44) );
  NAND3_X1 npu_inst_pe_1_7_4_U108 ( .A1(npu_inst_pe_1_7_4_n4), .A2(
        npu_inst_pe_1_7_4_n7), .A3(npu_inst_pe_1_7_4_n8), .ZN(
        npu_inst_pe_1_7_4_n40) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_7_4_n34), .CK(
        npu_inst_pe_1_7_4_net2913), .RN(npu_inst_pe_1_7_4_n9), .Q(
        npu_inst_pe_1_7_4_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_7_4_n35), .CK(
        npu_inst_pe_1_7_4_net2913), .RN(npu_inst_pe_1_7_4_n9), .Q(
        npu_inst_pe_1_7_4_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_7_4_n36), .CK(
        npu_inst_pe_1_7_4_net2913), .RN(npu_inst_pe_1_7_4_n9), .Q(
        npu_inst_pe_1_7_4_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_7_4_n98), .CK(
        npu_inst_pe_1_7_4_net2913), .RN(npu_inst_pe_1_7_4_n9), .Q(
        npu_inst_pe_1_7_4_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_7_4_n99), .CK(
        npu_inst_pe_1_7_4_net2913), .RN(npu_inst_pe_1_7_4_n9), .Q(
        npu_inst_pe_1_7_4_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_7_4_n100), 
        .CK(npu_inst_pe_1_7_4_net2913), .RN(npu_inst_pe_1_7_4_n9), .Q(
        npu_inst_pe_1_7_4_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_7_4_n33), .CK(
        npu_inst_pe_1_7_4_net2913), .RN(npu_inst_pe_1_7_4_n9), .Q(
        npu_inst_pe_1_7_4_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_7_4_n101), 
        .CK(npu_inst_pe_1_7_4_net2913), .RN(npu_inst_pe_1_7_4_n9), .Q(
        npu_inst_pe_1_7_4_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_weight_reg_0_ ( .D(npu_inst_n108), .CK(
        npu_inst_pe_1_7_4_net2919), .RN(npu_inst_pe_1_7_4_n9), .Q(
        npu_inst_pe_1_7_4_int_q_weight_0_), .QN(npu_inst_pe_1_7_4_n27) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_weight_reg_1_ ( .D(npu_inst_n114), .CK(
        npu_inst_pe_1_7_4_net2919), .RN(npu_inst_pe_1_7_4_n9), .Q(
        npu_inst_pe_1_7_4_int_q_weight_1_), .QN(npu_inst_pe_1_7_4_n26) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_7_4_n113), 
        .CK(npu_inst_pe_1_7_4_net2919), .RN(npu_inst_pe_1_7_4_n9), .Q(
        npu_inst_pe_1_7_4_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_7_4_n112), 
        .CK(npu_inst_pe_1_7_4_net2919), .RN(npu_inst_pe_1_7_4_n9), .Q(
        npu_inst_pe_1_7_4_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_7_4_n109), 
        .CK(npu_inst_pe_1_7_4_net2919), .RN(npu_inst_pe_1_7_4_n10), .Q(
        npu_inst_pe_1_7_4_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_7_4_n108), 
        .CK(npu_inst_pe_1_7_4_net2919), .RN(npu_inst_pe_1_7_4_n10), .Q(
        npu_inst_pe_1_7_4_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_7_4_n107), 
        .CK(npu_inst_pe_1_7_4_net2919), .RN(npu_inst_pe_1_7_4_n10), .Q(
        npu_inst_pe_1_7_4_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_7_4_n106), 
        .CK(npu_inst_pe_1_7_4_net2919), .RN(npu_inst_pe_1_7_4_n10), .Q(
        npu_inst_pe_1_7_4_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_7_4_n105), 
        .CK(npu_inst_pe_1_7_4_net2919), .RN(npu_inst_pe_1_7_4_n10), .Q(
        npu_inst_pe_1_7_4_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_7_4_n104), 
        .CK(npu_inst_pe_1_7_4_net2919), .RN(npu_inst_pe_1_7_4_n10), .Q(
        npu_inst_pe_1_7_4_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_7_4_n103), 
        .CK(npu_inst_pe_1_7_4_net2919), .RN(npu_inst_pe_1_7_4_n10), .Q(
        npu_inst_pe_1_7_4_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_7_4_n102), 
        .CK(npu_inst_pe_1_7_4_net2919), .RN(npu_inst_pe_1_7_4_n10), .Q(
        npu_inst_pe_1_7_4_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_7_4_n86), 
        .CK(npu_inst_pe_1_7_4_net2919), .RN(npu_inst_pe_1_7_4_n10), .Q(
        npu_inst_pe_1_7_4_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_7_4_n87), 
        .CK(npu_inst_pe_1_7_4_net2919), .RN(npu_inst_pe_1_7_4_n10), .Q(
        npu_inst_pe_1_7_4_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_7_4_n88), 
        .CK(npu_inst_pe_1_7_4_net2919), .RN(npu_inst_pe_1_7_4_n11), .Q(
        npu_inst_pe_1_7_4_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_7_4_n89), 
        .CK(npu_inst_pe_1_7_4_net2919), .RN(npu_inst_pe_1_7_4_n11), .Q(
        npu_inst_pe_1_7_4_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_7_4_n90), 
        .CK(npu_inst_pe_1_7_4_net2919), .RN(npu_inst_pe_1_7_4_n11), .Q(
        npu_inst_pe_1_7_4_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_7_4_n91), 
        .CK(npu_inst_pe_1_7_4_net2919), .RN(npu_inst_pe_1_7_4_n11), .Q(
        npu_inst_pe_1_7_4_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_7_4_n92), 
        .CK(npu_inst_pe_1_7_4_net2919), .RN(npu_inst_pe_1_7_4_n11), .Q(
        npu_inst_pe_1_7_4_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_7_4_n93), 
        .CK(npu_inst_pe_1_7_4_net2919), .RN(npu_inst_pe_1_7_4_n11), .Q(
        npu_inst_pe_1_7_4_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_7_4_n94), 
        .CK(npu_inst_pe_1_7_4_net2919), .RN(npu_inst_pe_1_7_4_n11), .Q(
        npu_inst_pe_1_7_4_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_7_4_n95), 
        .CK(npu_inst_pe_1_7_4_net2919), .RN(npu_inst_pe_1_7_4_n11), .Q(
        npu_inst_pe_1_7_4_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_7_4_n96), 
        .CK(npu_inst_pe_1_7_4_net2919), .RN(npu_inst_pe_1_7_4_n11), .Q(
        npu_inst_pe_1_7_4_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_7_4_n97), 
        .CK(npu_inst_pe_1_7_4_net2919), .RN(npu_inst_pe_1_7_4_n11), .Q(
        npu_inst_pe_1_7_4_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_7_4_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_7_4_N84), .SE(1'b0), .GCK(npu_inst_pe_1_7_4_net2913) );
  CLKGATETST_X1 npu_inst_pe_1_7_4_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n61), .SE(1'b0), .GCK(npu_inst_pe_1_7_4_net2919) );
  MUX2_X1 npu_inst_pe_1_7_5_U162 ( .A(npu_inst_pe_1_7_5_n32), .B(
        npu_inst_pe_1_7_5_n29), .S(npu_inst_pe_1_7_5_n8), .Z(
        npu_inst_pe_1_7_5_N93) );
  MUX2_X1 npu_inst_pe_1_7_5_U161 ( .A(npu_inst_pe_1_7_5_n31), .B(
        npu_inst_pe_1_7_5_n30), .S(npu_inst_pe_1_7_5_n6), .Z(
        npu_inst_pe_1_7_5_n32) );
  MUX2_X1 npu_inst_pe_1_7_5_U160 ( .A(npu_inst_pe_1_7_5_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_7_5_int_q_reg_v_1__0_), .S(npu_inst_pe_1_7_5_n4), .Z(
        npu_inst_pe_1_7_5_n31) );
  MUX2_X1 npu_inst_pe_1_7_5_U159 ( .A(npu_inst_pe_1_7_5_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_7_5_int_q_reg_v_3__0_), .S(npu_inst_pe_1_7_5_n4), .Z(
        npu_inst_pe_1_7_5_n30) );
  MUX2_X1 npu_inst_pe_1_7_5_U158 ( .A(npu_inst_pe_1_7_5_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_7_5_int_q_reg_v_5__0_), .S(npu_inst_pe_1_7_5_n4), .Z(
        npu_inst_pe_1_7_5_n29) );
  MUX2_X1 npu_inst_pe_1_7_5_U157 ( .A(npu_inst_pe_1_7_5_n28), .B(
        npu_inst_pe_1_7_5_n23), .S(npu_inst_pe_1_7_5_n8), .Z(
        npu_inst_pe_1_7_5_N94) );
  MUX2_X1 npu_inst_pe_1_7_5_U156 ( .A(npu_inst_pe_1_7_5_n25), .B(
        npu_inst_pe_1_7_5_n24), .S(npu_inst_pe_1_7_5_n6), .Z(
        npu_inst_pe_1_7_5_n28) );
  MUX2_X1 npu_inst_pe_1_7_5_U155 ( .A(npu_inst_pe_1_7_5_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_7_5_int_q_reg_v_1__1_), .S(npu_inst_pe_1_7_5_n4), .Z(
        npu_inst_pe_1_7_5_n25) );
  MUX2_X1 npu_inst_pe_1_7_5_U154 ( .A(npu_inst_pe_1_7_5_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_7_5_int_q_reg_v_3__1_), .S(npu_inst_pe_1_7_5_n4), .Z(
        npu_inst_pe_1_7_5_n24) );
  MUX2_X1 npu_inst_pe_1_7_5_U153 ( .A(npu_inst_pe_1_7_5_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_7_5_int_q_reg_v_5__1_), .S(npu_inst_pe_1_7_5_n4), .Z(
        npu_inst_pe_1_7_5_n23) );
  MUX2_X1 npu_inst_pe_1_7_5_U152 ( .A(npu_inst_pe_1_7_5_n22), .B(
        npu_inst_pe_1_7_5_n19), .S(npu_inst_pe_1_7_5_n8), .Z(
        npu_inst_int_data_x_7__5__1_) );
  MUX2_X1 npu_inst_pe_1_7_5_U151 ( .A(npu_inst_pe_1_7_5_n21), .B(
        npu_inst_pe_1_7_5_n20), .S(npu_inst_pe_1_7_5_n6), .Z(
        npu_inst_pe_1_7_5_n22) );
  MUX2_X1 npu_inst_pe_1_7_5_U150 ( .A(npu_inst_pe_1_7_5_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_7_5_int_q_reg_h_1__1_), .S(npu_inst_pe_1_7_5_n4), .Z(
        npu_inst_pe_1_7_5_n21) );
  MUX2_X1 npu_inst_pe_1_7_5_U149 ( .A(npu_inst_pe_1_7_5_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_7_5_int_q_reg_h_3__1_), .S(npu_inst_pe_1_7_5_n4), .Z(
        npu_inst_pe_1_7_5_n20) );
  MUX2_X1 npu_inst_pe_1_7_5_U148 ( .A(npu_inst_pe_1_7_5_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_7_5_int_q_reg_h_5__1_), .S(npu_inst_pe_1_7_5_n4), .Z(
        npu_inst_pe_1_7_5_n19) );
  MUX2_X1 npu_inst_pe_1_7_5_U147 ( .A(npu_inst_pe_1_7_5_n18), .B(
        npu_inst_pe_1_7_5_n15), .S(npu_inst_pe_1_7_5_n8), .Z(
        npu_inst_int_data_x_7__5__0_) );
  MUX2_X1 npu_inst_pe_1_7_5_U146 ( .A(npu_inst_pe_1_7_5_n17), .B(
        npu_inst_pe_1_7_5_n16), .S(npu_inst_pe_1_7_5_n6), .Z(
        npu_inst_pe_1_7_5_n18) );
  MUX2_X1 npu_inst_pe_1_7_5_U145 ( .A(npu_inst_pe_1_7_5_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_7_5_int_q_reg_h_1__0_), .S(npu_inst_pe_1_7_5_n4), .Z(
        npu_inst_pe_1_7_5_n17) );
  MUX2_X1 npu_inst_pe_1_7_5_U144 ( .A(npu_inst_pe_1_7_5_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_7_5_int_q_reg_h_3__0_), .S(npu_inst_pe_1_7_5_n4), .Z(
        npu_inst_pe_1_7_5_n16) );
  MUX2_X1 npu_inst_pe_1_7_5_U143 ( .A(npu_inst_pe_1_7_5_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_7_5_int_q_reg_h_5__0_), .S(npu_inst_pe_1_7_5_n4), .Z(
        npu_inst_pe_1_7_5_n15) );
  XOR2_X1 npu_inst_pe_1_7_5_U142 ( .A(npu_inst_pe_1_7_5_int_data_0_), .B(
        npu_inst_pe_1_7_5_int_q_acc_0_), .Z(npu_inst_pe_1_7_5_N73) );
  AND2_X1 npu_inst_pe_1_7_5_U141 ( .A1(npu_inst_pe_1_7_5_int_q_acc_0_), .A2(
        npu_inst_pe_1_7_5_int_data_0_), .ZN(npu_inst_pe_1_7_5_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_7_5_U140 ( .A(npu_inst_pe_1_7_5_int_q_acc_0_), .B(
        npu_inst_pe_1_7_5_n13), .ZN(npu_inst_pe_1_7_5_N65) );
  OR2_X1 npu_inst_pe_1_7_5_U139 ( .A1(npu_inst_pe_1_7_5_n13), .A2(
        npu_inst_pe_1_7_5_int_q_acc_0_), .ZN(npu_inst_pe_1_7_5_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_7_5_U138 ( .A(npu_inst_pe_1_7_5_int_q_acc_2_), .B(
        npu_inst_pe_1_7_5_add_79_carry_2_), .Z(npu_inst_pe_1_7_5_N75) );
  AND2_X1 npu_inst_pe_1_7_5_U137 ( .A1(npu_inst_pe_1_7_5_add_79_carry_2_), 
        .A2(npu_inst_pe_1_7_5_int_q_acc_2_), .ZN(
        npu_inst_pe_1_7_5_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_7_5_U136 ( .A(npu_inst_pe_1_7_5_int_q_acc_3_), .B(
        npu_inst_pe_1_7_5_add_79_carry_3_), .Z(npu_inst_pe_1_7_5_N76) );
  AND2_X1 npu_inst_pe_1_7_5_U135 ( .A1(npu_inst_pe_1_7_5_add_79_carry_3_), 
        .A2(npu_inst_pe_1_7_5_int_q_acc_3_), .ZN(
        npu_inst_pe_1_7_5_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_7_5_U134 ( .A(npu_inst_pe_1_7_5_int_q_acc_4_), .B(
        npu_inst_pe_1_7_5_add_79_carry_4_), .Z(npu_inst_pe_1_7_5_N77) );
  AND2_X1 npu_inst_pe_1_7_5_U133 ( .A1(npu_inst_pe_1_7_5_add_79_carry_4_), 
        .A2(npu_inst_pe_1_7_5_int_q_acc_4_), .ZN(
        npu_inst_pe_1_7_5_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_7_5_U132 ( .A(npu_inst_pe_1_7_5_int_q_acc_5_), .B(
        npu_inst_pe_1_7_5_add_79_carry_5_), .Z(npu_inst_pe_1_7_5_N78) );
  AND2_X1 npu_inst_pe_1_7_5_U131 ( .A1(npu_inst_pe_1_7_5_add_79_carry_5_), 
        .A2(npu_inst_pe_1_7_5_int_q_acc_5_), .ZN(
        npu_inst_pe_1_7_5_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_7_5_U130 ( .A(npu_inst_pe_1_7_5_int_q_acc_6_), .B(
        npu_inst_pe_1_7_5_add_79_carry_6_), .Z(npu_inst_pe_1_7_5_N79) );
  AND2_X1 npu_inst_pe_1_7_5_U129 ( .A1(npu_inst_pe_1_7_5_add_79_carry_6_), 
        .A2(npu_inst_pe_1_7_5_int_q_acc_6_), .ZN(
        npu_inst_pe_1_7_5_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_7_5_U128 ( .A(npu_inst_pe_1_7_5_int_q_acc_7_), .B(
        npu_inst_pe_1_7_5_add_79_carry_7_), .Z(npu_inst_pe_1_7_5_N80) );
  XNOR2_X1 npu_inst_pe_1_7_5_U127 ( .A(npu_inst_pe_1_7_5_sub_77_carry_2_), .B(
        npu_inst_pe_1_7_5_int_q_acc_2_), .ZN(npu_inst_pe_1_7_5_N67) );
  OR2_X1 npu_inst_pe_1_7_5_U126 ( .A1(npu_inst_pe_1_7_5_int_q_acc_2_), .A2(
        npu_inst_pe_1_7_5_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_7_5_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_7_5_U125 ( .A(npu_inst_pe_1_7_5_sub_77_carry_3_), .B(
        npu_inst_pe_1_7_5_int_q_acc_3_), .ZN(npu_inst_pe_1_7_5_N68) );
  OR2_X1 npu_inst_pe_1_7_5_U124 ( .A1(npu_inst_pe_1_7_5_int_q_acc_3_), .A2(
        npu_inst_pe_1_7_5_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_7_5_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_7_5_U123 ( .A(npu_inst_pe_1_7_5_sub_77_carry_4_), .B(
        npu_inst_pe_1_7_5_int_q_acc_4_), .ZN(npu_inst_pe_1_7_5_N69) );
  OR2_X1 npu_inst_pe_1_7_5_U122 ( .A1(npu_inst_pe_1_7_5_int_q_acc_4_), .A2(
        npu_inst_pe_1_7_5_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_7_5_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_7_5_U121 ( .A(npu_inst_pe_1_7_5_sub_77_carry_5_), .B(
        npu_inst_pe_1_7_5_int_q_acc_5_), .ZN(npu_inst_pe_1_7_5_N70) );
  OR2_X1 npu_inst_pe_1_7_5_U120 ( .A1(npu_inst_pe_1_7_5_int_q_acc_5_), .A2(
        npu_inst_pe_1_7_5_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_7_5_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_7_5_U119 ( .A(npu_inst_pe_1_7_5_sub_77_carry_6_), .B(
        npu_inst_pe_1_7_5_int_q_acc_6_), .ZN(npu_inst_pe_1_7_5_N71) );
  OR2_X1 npu_inst_pe_1_7_5_U118 ( .A1(npu_inst_pe_1_7_5_int_q_acc_6_), .A2(
        npu_inst_pe_1_7_5_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_7_5_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_7_5_U117 ( .A(npu_inst_pe_1_7_5_int_q_acc_7_), .B(
        npu_inst_pe_1_7_5_sub_77_carry_7_), .ZN(npu_inst_pe_1_7_5_N72) );
  INV_X1 npu_inst_pe_1_7_5_U116 ( .A(npu_inst_n75), .ZN(npu_inst_pe_1_7_5_n7)
         );
  INV_X1 npu_inst_pe_1_7_5_U115 ( .A(npu_inst_pe_1_7_5_n7), .ZN(
        npu_inst_pe_1_7_5_n6) );
  INV_X1 npu_inst_pe_1_7_5_U114 ( .A(npu_inst_n52), .ZN(npu_inst_pe_1_7_5_n3)
         );
  AOI22_X1 npu_inst_pe_1_7_5_U113 ( .A1(npu_inst_pe_1_7_5_n38), .A2(
        int_i_data_v_npu[5]), .B1(npu_inst_pe_1_7_5_n118), .B2(
        npu_inst_pe_1_7_5_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_7_5_n39) );
  INV_X1 npu_inst_pe_1_7_5_U112 ( .A(npu_inst_pe_1_7_5_n39), .ZN(
        npu_inst_pe_1_7_5_n112) );
  AOI22_X1 npu_inst_pe_1_7_5_U111 ( .A1(npu_inst_pe_1_7_5_n38), .A2(
        int_i_data_v_npu[4]), .B1(npu_inst_pe_1_7_5_n118), .B2(
        npu_inst_pe_1_7_5_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_7_5_n37) );
  INV_X1 npu_inst_pe_1_7_5_U110 ( .A(npu_inst_pe_1_7_5_n37), .ZN(
        npu_inst_pe_1_7_5_n113) );
  AOI22_X1 npu_inst_pe_1_7_5_U107 ( .A1(int_i_data_v_npu[5]), .A2(
        npu_inst_pe_1_7_5_n58), .B1(npu_inst_pe_1_7_5_n114), .B2(
        npu_inst_pe_1_7_5_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_7_5_n59) );
  INV_X1 npu_inst_pe_1_7_5_U106 ( .A(npu_inst_pe_1_7_5_n59), .ZN(
        npu_inst_pe_1_7_5_n102) );
  AOI22_X1 npu_inst_pe_1_7_5_U105 ( .A1(int_i_data_v_npu[4]), .A2(
        npu_inst_pe_1_7_5_n58), .B1(npu_inst_pe_1_7_5_n114), .B2(
        npu_inst_pe_1_7_5_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_7_5_n57) );
  INV_X1 npu_inst_pe_1_7_5_U104 ( .A(npu_inst_pe_1_7_5_n57), .ZN(
        npu_inst_pe_1_7_5_n103) );
  AOI22_X1 npu_inst_pe_1_7_5_U103 ( .A1(int_i_data_v_npu[5]), .A2(
        npu_inst_pe_1_7_5_n54), .B1(npu_inst_pe_1_7_5_n115), .B2(
        npu_inst_pe_1_7_5_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_7_5_n55) );
  INV_X1 npu_inst_pe_1_7_5_U102 ( .A(npu_inst_pe_1_7_5_n55), .ZN(
        npu_inst_pe_1_7_5_n104) );
  AOI22_X1 npu_inst_pe_1_7_5_U101 ( .A1(int_i_data_v_npu[4]), .A2(
        npu_inst_pe_1_7_5_n54), .B1(npu_inst_pe_1_7_5_n115), .B2(
        npu_inst_pe_1_7_5_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_7_5_n53) );
  INV_X1 npu_inst_pe_1_7_5_U100 ( .A(npu_inst_pe_1_7_5_n53), .ZN(
        npu_inst_pe_1_7_5_n105) );
  AOI22_X1 npu_inst_pe_1_7_5_U99 ( .A1(int_i_data_v_npu[5]), .A2(
        npu_inst_pe_1_7_5_n50), .B1(npu_inst_pe_1_7_5_n116), .B2(
        npu_inst_pe_1_7_5_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_7_5_n51) );
  INV_X1 npu_inst_pe_1_7_5_U98 ( .A(npu_inst_pe_1_7_5_n51), .ZN(
        npu_inst_pe_1_7_5_n106) );
  AOI22_X1 npu_inst_pe_1_7_5_U97 ( .A1(int_i_data_v_npu[4]), .A2(
        npu_inst_pe_1_7_5_n50), .B1(npu_inst_pe_1_7_5_n116), .B2(
        npu_inst_pe_1_7_5_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_7_5_n49) );
  INV_X1 npu_inst_pe_1_7_5_U96 ( .A(npu_inst_pe_1_7_5_n49), .ZN(
        npu_inst_pe_1_7_5_n107) );
  AOI22_X1 npu_inst_pe_1_7_5_U95 ( .A1(int_i_data_v_npu[5]), .A2(
        npu_inst_pe_1_7_5_n46), .B1(npu_inst_pe_1_7_5_n117), .B2(
        npu_inst_pe_1_7_5_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_7_5_n47) );
  INV_X1 npu_inst_pe_1_7_5_U94 ( .A(npu_inst_pe_1_7_5_n47), .ZN(
        npu_inst_pe_1_7_5_n108) );
  AOI22_X1 npu_inst_pe_1_7_5_U93 ( .A1(int_i_data_v_npu[4]), .A2(
        npu_inst_pe_1_7_5_n46), .B1(npu_inst_pe_1_7_5_n117), .B2(
        npu_inst_pe_1_7_5_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_7_5_n45) );
  INV_X1 npu_inst_pe_1_7_5_U92 ( .A(npu_inst_pe_1_7_5_n45), .ZN(
        npu_inst_pe_1_7_5_n109) );
  AOI22_X1 npu_inst_pe_1_7_5_U91 ( .A1(int_i_data_v_npu[5]), .A2(
        npu_inst_pe_1_7_5_n42), .B1(npu_inst_pe_1_7_5_n119), .B2(
        npu_inst_pe_1_7_5_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_7_5_n43) );
  INV_X1 npu_inst_pe_1_7_5_U90 ( .A(npu_inst_pe_1_7_5_n43), .ZN(
        npu_inst_pe_1_7_5_n110) );
  AOI22_X1 npu_inst_pe_1_7_5_U89 ( .A1(int_i_data_v_npu[4]), .A2(
        npu_inst_pe_1_7_5_n42), .B1(npu_inst_pe_1_7_5_n119), .B2(
        npu_inst_pe_1_7_5_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_7_5_n41) );
  INV_X1 npu_inst_pe_1_7_5_U88 ( .A(npu_inst_pe_1_7_5_n41), .ZN(
        npu_inst_pe_1_7_5_n111) );
  NAND2_X1 npu_inst_pe_1_7_5_U87 ( .A1(npu_inst_pe_1_7_5_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_7_5_n60), .ZN(npu_inst_pe_1_7_5_n74) );
  OAI21_X1 npu_inst_pe_1_7_5_U86 ( .B1(npu_inst_pe_1_7_5_n63), .B2(
        npu_inst_pe_1_7_5_n60), .A(npu_inst_pe_1_7_5_n74), .ZN(
        npu_inst_pe_1_7_5_n97) );
  NAND2_X1 npu_inst_pe_1_7_5_U85 ( .A1(npu_inst_pe_1_7_5_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_7_5_n60), .ZN(npu_inst_pe_1_7_5_n73) );
  OAI21_X1 npu_inst_pe_1_7_5_U84 ( .B1(npu_inst_pe_1_7_5_n61), .B2(
        npu_inst_pe_1_7_5_n60), .A(npu_inst_pe_1_7_5_n73), .ZN(
        npu_inst_pe_1_7_5_n96) );
  NAND2_X1 npu_inst_pe_1_7_5_U83 ( .A1(npu_inst_pe_1_7_5_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_7_5_n56), .ZN(npu_inst_pe_1_7_5_n72) );
  OAI21_X1 npu_inst_pe_1_7_5_U82 ( .B1(npu_inst_pe_1_7_5_n63), .B2(
        npu_inst_pe_1_7_5_n56), .A(npu_inst_pe_1_7_5_n72), .ZN(
        npu_inst_pe_1_7_5_n95) );
  NAND2_X1 npu_inst_pe_1_7_5_U81 ( .A1(npu_inst_pe_1_7_5_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_7_5_n56), .ZN(npu_inst_pe_1_7_5_n71) );
  OAI21_X1 npu_inst_pe_1_7_5_U80 ( .B1(npu_inst_pe_1_7_5_n61), .B2(
        npu_inst_pe_1_7_5_n56), .A(npu_inst_pe_1_7_5_n71), .ZN(
        npu_inst_pe_1_7_5_n94) );
  NAND2_X1 npu_inst_pe_1_7_5_U79 ( .A1(npu_inst_pe_1_7_5_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_7_5_n52), .ZN(npu_inst_pe_1_7_5_n70) );
  OAI21_X1 npu_inst_pe_1_7_5_U78 ( .B1(npu_inst_pe_1_7_5_n63), .B2(
        npu_inst_pe_1_7_5_n52), .A(npu_inst_pe_1_7_5_n70), .ZN(
        npu_inst_pe_1_7_5_n93) );
  NAND2_X1 npu_inst_pe_1_7_5_U77 ( .A1(npu_inst_pe_1_7_5_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_7_5_n52), .ZN(npu_inst_pe_1_7_5_n69) );
  OAI21_X1 npu_inst_pe_1_7_5_U76 ( .B1(npu_inst_pe_1_7_5_n61), .B2(
        npu_inst_pe_1_7_5_n52), .A(npu_inst_pe_1_7_5_n69), .ZN(
        npu_inst_pe_1_7_5_n92) );
  NAND2_X1 npu_inst_pe_1_7_5_U75 ( .A1(npu_inst_pe_1_7_5_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_7_5_n48), .ZN(npu_inst_pe_1_7_5_n68) );
  OAI21_X1 npu_inst_pe_1_7_5_U74 ( .B1(npu_inst_pe_1_7_5_n63), .B2(
        npu_inst_pe_1_7_5_n48), .A(npu_inst_pe_1_7_5_n68), .ZN(
        npu_inst_pe_1_7_5_n91) );
  NAND2_X1 npu_inst_pe_1_7_5_U73 ( .A1(npu_inst_pe_1_7_5_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_7_5_n48), .ZN(npu_inst_pe_1_7_5_n67) );
  OAI21_X1 npu_inst_pe_1_7_5_U72 ( .B1(npu_inst_pe_1_7_5_n61), .B2(
        npu_inst_pe_1_7_5_n48), .A(npu_inst_pe_1_7_5_n67), .ZN(
        npu_inst_pe_1_7_5_n90) );
  NAND2_X1 npu_inst_pe_1_7_5_U71 ( .A1(npu_inst_pe_1_7_5_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_7_5_n44), .ZN(npu_inst_pe_1_7_5_n66) );
  OAI21_X1 npu_inst_pe_1_7_5_U70 ( .B1(npu_inst_pe_1_7_5_n63), .B2(
        npu_inst_pe_1_7_5_n44), .A(npu_inst_pe_1_7_5_n66), .ZN(
        npu_inst_pe_1_7_5_n89) );
  NAND2_X1 npu_inst_pe_1_7_5_U69 ( .A1(npu_inst_pe_1_7_5_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_7_5_n44), .ZN(npu_inst_pe_1_7_5_n65) );
  OAI21_X1 npu_inst_pe_1_7_5_U68 ( .B1(npu_inst_pe_1_7_5_n61), .B2(
        npu_inst_pe_1_7_5_n44), .A(npu_inst_pe_1_7_5_n65), .ZN(
        npu_inst_pe_1_7_5_n88) );
  NAND2_X1 npu_inst_pe_1_7_5_U67 ( .A1(npu_inst_pe_1_7_5_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_7_5_n40), .ZN(npu_inst_pe_1_7_5_n64) );
  OAI21_X1 npu_inst_pe_1_7_5_U66 ( .B1(npu_inst_pe_1_7_5_n63), .B2(
        npu_inst_pe_1_7_5_n40), .A(npu_inst_pe_1_7_5_n64), .ZN(
        npu_inst_pe_1_7_5_n87) );
  NAND2_X1 npu_inst_pe_1_7_5_U65 ( .A1(npu_inst_pe_1_7_5_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_7_5_n40), .ZN(npu_inst_pe_1_7_5_n62) );
  OAI21_X1 npu_inst_pe_1_7_5_U64 ( .B1(npu_inst_pe_1_7_5_n61), .B2(
        npu_inst_pe_1_7_5_n40), .A(npu_inst_pe_1_7_5_n62), .ZN(
        npu_inst_pe_1_7_5_n86) );
  AND2_X1 npu_inst_pe_1_7_5_U63 ( .A1(npu_inst_pe_1_7_5_N93), .A2(npu_inst_n52), .ZN(npu_inst_int_data_y_7__5__0_) );
  AND2_X1 npu_inst_pe_1_7_5_U62 ( .A1(npu_inst_n52), .A2(npu_inst_pe_1_7_5_N94), .ZN(npu_inst_int_data_y_7__5__1_) );
  AOI22_X1 npu_inst_pe_1_7_5_U61 ( .A1(npu_inst_n52), .A2(int_i_data_v_npu[5]), 
        .B1(npu_inst_pe_1_7_5_n3), .B2(npu_inst_int_data_x_7__6__1_), .ZN(
        npu_inst_pe_1_7_5_n63) );
  AOI22_X1 npu_inst_pe_1_7_5_U60 ( .A1(npu_inst_n52), .A2(int_i_data_v_npu[4]), 
        .B1(npu_inst_pe_1_7_5_n3), .B2(npu_inst_int_data_x_7__6__0_), .ZN(
        npu_inst_pe_1_7_5_n61) );
  NOR3_X1 npu_inst_pe_1_7_5_U59 ( .A1(npu_inst_pe_1_7_5_n26), .A2(npu_inst_n52), .A3(npu_inst_int_ckg[2]), .ZN(npu_inst_pe_1_7_5_n85) );
  OR2_X1 npu_inst_pe_1_7_5_U58 ( .A1(npu_inst_pe_1_7_5_n85), .A2(
        npu_inst_pe_1_7_5_n2), .ZN(npu_inst_pe_1_7_5_N84) );
  AOI222_X1 npu_inst_pe_1_7_5_U57 ( .A1(1'b0), .A2(npu_inst_pe_1_7_5_n1), .B1(
        npu_inst_pe_1_7_5_N73), .B2(npu_inst_pe_1_7_5_n76), .C1(
        npu_inst_pe_1_7_5_N65), .C2(npu_inst_pe_1_7_5_n77), .ZN(
        npu_inst_pe_1_7_5_n84) );
  INV_X1 npu_inst_pe_1_7_5_U56 ( .A(npu_inst_pe_1_7_5_n84), .ZN(
        npu_inst_pe_1_7_5_n101) );
  AOI222_X1 npu_inst_pe_1_7_5_U55 ( .A1(1'b0), .A2(npu_inst_pe_1_7_5_n1), .B1(
        npu_inst_pe_1_7_5_N80), .B2(npu_inst_pe_1_7_5_n76), .C1(
        npu_inst_pe_1_7_5_N72), .C2(npu_inst_pe_1_7_5_n77), .ZN(
        npu_inst_pe_1_7_5_n75) );
  INV_X1 npu_inst_pe_1_7_5_U54 ( .A(npu_inst_pe_1_7_5_n75), .ZN(
        npu_inst_pe_1_7_5_n33) );
  AOI222_X1 npu_inst_pe_1_7_5_U53 ( .A1(1'b0), .A2(npu_inst_pe_1_7_5_n1), .B1(
        npu_inst_pe_1_7_5_N74), .B2(npu_inst_pe_1_7_5_n76), .C1(
        npu_inst_pe_1_7_5_N66), .C2(npu_inst_pe_1_7_5_n77), .ZN(
        npu_inst_pe_1_7_5_n83) );
  INV_X1 npu_inst_pe_1_7_5_U52 ( .A(npu_inst_pe_1_7_5_n83), .ZN(
        npu_inst_pe_1_7_5_n100) );
  AOI222_X1 npu_inst_pe_1_7_5_U51 ( .A1(1'b0), .A2(npu_inst_pe_1_7_5_n1), .B1(
        npu_inst_pe_1_7_5_N75), .B2(npu_inst_pe_1_7_5_n76), .C1(
        npu_inst_pe_1_7_5_N67), .C2(npu_inst_pe_1_7_5_n77), .ZN(
        npu_inst_pe_1_7_5_n82) );
  INV_X1 npu_inst_pe_1_7_5_U50 ( .A(npu_inst_pe_1_7_5_n82), .ZN(
        npu_inst_pe_1_7_5_n99) );
  AOI222_X1 npu_inst_pe_1_7_5_U49 ( .A1(1'b0), .A2(npu_inst_pe_1_7_5_n1), .B1(
        npu_inst_pe_1_7_5_N76), .B2(npu_inst_pe_1_7_5_n76), .C1(
        npu_inst_pe_1_7_5_N68), .C2(npu_inst_pe_1_7_5_n77), .ZN(
        npu_inst_pe_1_7_5_n81) );
  INV_X1 npu_inst_pe_1_7_5_U48 ( .A(npu_inst_pe_1_7_5_n81), .ZN(
        npu_inst_pe_1_7_5_n98) );
  AOI222_X1 npu_inst_pe_1_7_5_U47 ( .A1(1'b0), .A2(npu_inst_pe_1_7_5_n1), .B1(
        npu_inst_pe_1_7_5_N77), .B2(npu_inst_pe_1_7_5_n76), .C1(
        npu_inst_pe_1_7_5_N69), .C2(npu_inst_pe_1_7_5_n77), .ZN(
        npu_inst_pe_1_7_5_n80) );
  INV_X1 npu_inst_pe_1_7_5_U46 ( .A(npu_inst_pe_1_7_5_n80), .ZN(
        npu_inst_pe_1_7_5_n36) );
  AOI222_X1 npu_inst_pe_1_7_5_U45 ( .A1(1'b0), .A2(npu_inst_pe_1_7_5_n1), .B1(
        npu_inst_pe_1_7_5_N78), .B2(npu_inst_pe_1_7_5_n76), .C1(
        npu_inst_pe_1_7_5_N70), .C2(npu_inst_pe_1_7_5_n77), .ZN(
        npu_inst_pe_1_7_5_n79) );
  INV_X1 npu_inst_pe_1_7_5_U44 ( .A(npu_inst_pe_1_7_5_n79), .ZN(
        npu_inst_pe_1_7_5_n35) );
  AOI222_X1 npu_inst_pe_1_7_5_U43 ( .A1(1'b0), .A2(npu_inst_pe_1_7_5_n1), .B1(
        npu_inst_pe_1_7_5_N79), .B2(npu_inst_pe_1_7_5_n76), .C1(
        npu_inst_pe_1_7_5_N71), .C2(npu_inst_pe_1_7_5_n77), .ZN(
        npu_inst_pe_1_7_5_n78) );
  INV_X1 npu_inst_pe_1_7_5_U42 ( .A(npu_inst_pe_1_7_5_n78), .ZN(
        npu_inst_pe_1_7_5_n34) );
  AND2_X1 npu_inst_pe_1_7_5_U41 ( .A1(npu_inst_pe_1_7_5_int_q_acc_0_), .A2(
        npu_inst_pe_1_7_5_n1), .ZN(npu_inst_int_data_res_7__5__0_) );
  AND2_X1 npu_inst_pe_1_7_5_U40 ( .A1(npu_inst_pe_1_7_5_n2), .A2(
        npu_inst_pe_1_7_5_int_q_acc_7_), .ZN(npu_inst_int_data_res_7__5__7_)
         );
  AND2_X1 npu_inst_pe_1_7_5_U39 ( .A1(npu_inst_pe_1_7_5_int_q_acc_1_), .A2(
        npu_inst_pe_1_7_5_n1), .ZN(npu_inst_int_data_res_7__5__1_) );
  AND2_X1 npu_inst_pe_1_7_5_U38 ( .A1(npu_inst_pe_1_7_5_int_q_acc_2_), .A2(
        npu_inst_pe_1_7_5_n1), .ZN(npu_inst_int_data_res_7__5__2_) );
  AND2_X1 npu_inst_pe_1_7_5_U37 ( .A1(npu_inst_pe_1_7_5_int_q_acc_3_), .A2(
        npu_inst_pe_1_7_5_n2), .ZN(npu_inst_int_data_res_7__5__3_) );
  AND2_X1 npu_inst_pe_1_7_5_U36 ( .A1(npu_inst_pe_1_7_5_int_q_acc_4_), .A2(
        npu_inst_pe_1_7_5_n2), .ZN(npu_inst_int_data_res_7__5__4_) );
  AND2_X1 npu_inst_pe_1_7_5_U35 ( .A1(npu_inst_pe_1_7_5_int_q_acc_5_), .A2(
        npu_inst_pe_1_7_5_n2), .ZN(npu_inst_int_data_res_7__5__5_) );
  AND2_X1 npu_inst_pe_1_7_5_U34 ( .A1(npu_inst_pe_1_7_5_int_q_acc_6_), .A2(
        npu_inst_pe_1_7_5_n2), .ZN(npu_inst_int_data_res_7__5__6_) );
  INV_X1 npu_inst_pe_1_7_5_U33 ( .A(npu_inst_pe_1_7_5_int_data_1_), .ZN(
        npu_inst_pe_1_7_5_n14) );
  AND2_X1 npu_inst_pe_1_7_5_U32 ( .A1(npu_inst_int_data_x_7__5__1_), .A2(
        npu_inst_pe_1_7_5_int_q_weight_1_), .ZN(npu_inst_pe_1_7_5_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_7_5_U31 ( .A1(npu_inst_int_data_x_7__5__0_), .A2(
        npu_inst_pe_1_7_5_int_q_weight_1_), .ZN(npu_inst_pe_1_7_5_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_7_5_U30 ( .A(npu_inst_pe_1_7_5_int_data_0_), .ZN(
        npu_inst_pe_1_7_5_n13) );
  INV_X1 npu_inst_pe_1_7_5_U29 ( .A(npu_inst_n67), .ZN(npu_inst_pe_1_7_5_n5)
         );
  OR3_X1 npu_inst_pe_1_7_5_U28 ( .A1(npu_inst_pe_1_7_5_n6), .A2(
        npu_inst_pe_1_7_5_n8), .A3(npu_inst_pe_1_7_5_n5), .ZN(
        npu_inst_pe_1_7_5_n56) );
  OR3_X1 npu_inst_pe_1_7_5_U27 ( .A1(npu_inst_pe_1_7_5_n5), .A2(
        npu_inst_pe_1_7_5_n8), .A3(npu_inst_pe_1_7_5_n7), .ZN(
        npu_inst_pe_1_7_5_n48) );
  INV_X1 npu_inst_pe_1_7_5_U26 ( .A(npu_inst_pe_1_7_5_n5), .ZN(
        npu_inst_pe_1_7_5_n4) );
  INV_X1 npu_inst_pe_1_7_5_U25 ( .A(npu_inst_n122), .ZN(npu_inst_pe_1_7_5_n12)
         );
  OR3_X1 npu_inst_pe_1_7_5_U24 ( .A1(npu_inst_pe_1_7_5_n4), .A2(
        npu_inst_pe_1_7_5_n8), .A3(npu_inst_pe_1_7_5_n7), .ZN(
        npu_inst_pe_1_7_5_n52) );
  OR3_X1 npu_inst_pe_1_7_5_U23 ( .A1(npu_inst_pe_1_7_5_n6), .A2(
        npu_inst_pe_1_7_5_n8), .A3(npu_inst_pe_1_7_5_n4), .ZN(
        npu_inst_pe_1_7_5_n60) );
  NOR2_X1 npu_inst_pe_1_7_5_U22 ( .A1(npu_inst_pe_1_7_5_n60), .A2(
        npu_inst_pe_1_7_5_n3), .ZN(npu_inst_pe_1_7_5_n58) );
  NOR2_X1 npu_inst_pe_1_7_5_U21 ( .A1(npu_inst_pe_1_7_5_n56), .A2(
        npu_inst_pe_1_7_5_n3), .ZN(npu_inst_pe_1_7_5_n54) );
  NOR2_X1 npu_inst_pe_1_7_5_U20 ( .A1(npu_inst_pe_1_7_5_n52), .A2(
        npu_inst_pe_1_7_5_n3), .ZN(npu_inst_pe_1_7_5_n50) );
  NOR2_X1 npu_inst_pe_1_7_5_U19 ( .A1(npu_inst_pe_1_7_5_n48), .A2(
        npu_inst_pe_1_7_5_n3), .ZN(npu_inst_pe_1_7_5_n46) );
  NOR2_X1 npu_inst_pe_1_7_5_U18 ( .A1(npu_inst_pe_1_7_5_n40), .A2(
        npu_inst_pe_1_7_5_n3), .ZN(npu_inst_pe_1_7_5_n38) );
  NOR2_X1 npu_inst_pe_1_7_5_U17 ( .A1(npu_inst_pe_1_7_5_n44), .A2(
        npu_inst_pe_1_7_5_n3), .ZN(npu_inst_pe_1_7_5_n42) );
  BUF_X1 npu_inst_pe_1_7_5_U16 ( .A(npu_inst_n92), .Z(npu_inst_pe_1_7_5_n8) );
  BUF_X1 npu_inst_pe_1_7_5_U15 ( .A(npu_inst_pe_1_7_5_n12), .Z(
        npu_inst_pe_1_7_5_n11) );
  BUF_X1 npu_inst_pe_1_7_5_U14 ( .A(npu_inst_pe_1_7_5_n12), .Z(
        npu_inst_pe_1_7_5_n10) );
  BUF_X1 npu_inst_pe_1_7_5_U13 ( .A(npu_inst_pe_1_7_5_n12), .Z(
        npu_inst_pe_1_7_5_n9) );
  INV_X1 npu_inst_pe_1_7_5_U12 ( .A(npu_inst_pe_1_7_5_n38), .ZN(
        npu_inst_pe_1_7_5_n118) );
  INV_X1 npu_inst_pe_1_7_5_U11 ( .A(npu_inst_pe_1_7_5_n58), .ZN(
        npu_inst_pe_1_7_5_n114) );
  INV_X1 npu_inst_pe_1_7_5_U10 ( .A(npu_inst_pe_1_7_5_n54), .ZN(
        npu_inst_pe_1_7_5_n115) );
  INV_X1 npu_inst_pe_1_7_5_U9 ( .A(npu_inst_pe_1_7_5_n50), .ZN(
        npu_inst_pe_1_7_5_n116) );
  INV_X1 npu_inst_pe_1_7_5_U8 ( .A(npu_inst_pe_1_7_5_n46), .ZN(
        npu_inst_pe_1_7_5_n117) );
  INV_X1 npu_inst_pe_1_7_5_U7 ( .A(npu_inst_pe_1_7_5_n42), .ZN(
        npu_inst_pe_1_7_5_n119) );
  BUF_X1 npu_inst_pe_1_7_5_U6 ( .A(npu_inst_n8), .Z(npu_inst_pe_1_7_5_n2) );
  BUF_X1 npu_inst_pe_1_7_5_U5 ( .A(npu_inst_n8), .Z(npu_inst_pe_1_7_5_n1) );
  NOR2_X1 npu_inst_pe_1_7_5_U4 ( .A1(npu_inst_pe_1_7_5_int_q_weight_0_), .A2(
        npu_inst_pe_1_7_5_n1), .ZN(npu_inst_pe_1_7_5_n76) );
  NOR2_X1 npu_inst_pe_1_7_5_U3 ( .A1(npu_inst_pe_1_7_5_n27), .A2(
        npu_inst_pe_1_7_5_n1), .ZN(npu_inst_pe_1_7_5_n77) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_7_5_n111), 
        .CK(npu_inst_pe_1_7_5_net2896), .RN(npu_inst_pe_1_7_5_n12), .Q(
        npu_inst_pe_1_7_5_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_7_5_n110), 
        .CK(npu_inst_pe_1_7_5_net2896), .RN(npu_inst_pe_1_7_5_n12), .Q(
        npu_inst_pe_1_7_5_int_q_reg_v_4__1_) );
  FA_X1 npu_inst_pe_1_7_5_sub_77_U2_1 ( .A(npu_inst_pe_1_7_5_int_q_acc_1_), 
        .B(npu_inst_pe_1_7_5_n14), .CI(npu_inst_pe_1_7_5_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_7_5_sub_77_carry_2_), .S(npu_inst_pe_1_7_5_N66) );
  FA_X1 npu_inst_pe_1_7_5_add_79_U1_1 ( .A(npu_inst_pe_1_7_5_int_q_acc_1_), 
        .B(npu_inst_pe_1_7_5_int_data_1_), .CI(
        npu_inst_pe_1_7_5_add_79_carry_1_), .CO(
        npu_inst_pe_1_7_5_add_79_carry_2_), .S(npu_inst_pe_1_7_5_N74) );
  NAND3_X1 npu_inst_pe_1_7_5_U109 ( .A1(npu_inst_pe_1_7_5_n5), .A2(
        npu_inst_pe_1_7_5_n7), .A3(npu_inst_pe_1_7_5_n8), .ZN(
        npu_inst_pe_1_7_5_n44) );
  NAND3_X1 npu_inst_pe_1_7_5_U108 ( .A1(npu_inst_pe_1_7_5_n4), .A2(
        npu_inst_pe_1_7_5_n7), .A3(npu_inst_pe_1_7_5_n8), .ZN(
        npu_inst_pe_1_7_5_n40) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_7_5_n34), .CK(
        npu_inst_pe_1_7_5_net2890), .RN(npu_inst_pe_1_7_5_n9), .Q(
        npu_inst_pe_1_7_5_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_7_5_n35), .CK(
        npu_inst_pe_1_7_5_net2890), .RN(npu_inst_pe_1_7_5_n9), .Q(
        npu_inst_pe_1_7_5_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_7_5_n36), .CK(
        npu_inst_pe_1_7_5_net2890), .RN(npu_inst_pe_1_7_5_n9), .Q(
        npu_inst_pe_1_7_5_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_7_5_n98), .CK(
        npu_inst_pe_1_7_5_net2890), .RN(npu_inst_pe_1_7_5_n9), .Q(
        npu_inst_pe_1_7_5_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_7_5_n99), .CK(
        npu_inst_pe_1_7_5_net2890), .RN(npu_inst_pe_1_7_5_n9), .Q(
        npu_inst_pe_1_7_5_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_7_5_n100), 
        .CK(npu_inst_pe_1_7_5_net2890), .RN(npu_inst_pe_1_7_5_n9), .Q(
        npu_inst_pe_1_7_5_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_7_5_n33), .CK(
        npu_inst_pe_1_7_5_net2890), .RN(npu_inst_pe_1_7_5_n9), .Q(
        npu_inst_pe_1_7_5_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_7_5_n101), 
        .CK(npu_inst_pe_1_7_5_net2890), .RN(npu_inst_pe_1_7_5_n9), .Q(
        npu_inst_pe_1_7_5_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_weight_reg_0_ ( .D(npu_inst_n108), .CK(
        npu_inst_pe_1_7_5_net2896), .RN(npu_inst_pe_1_7_5_n9), .Q(
        npu_inst_pe_1_7_5_int_q_weight_0_), .QN(npu_inst_pe_1_7_5_n27) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_weight_reg_1_ ( .D(npu_inst_n114), .CK(
        npu_inst_pe_1_7_5_net2896), .RN(npu_inst_pe_1_7_5_n9), .Q(
        npu_inst_pe_1_7_5_int_q_weight_1_), .QN(npu_inst_pe_1_7_5_n26) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_7_5_n113), 
        .CK(npu_inst_pe_1_7_5_net2896), .RN(npu_inst_pe_1_7_5_n9), .Q(
        npu_inst_pe_1_7_5_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_7_5_n112), 
        .CK(npu_inst_pe_1_7_5_net2896), .RN(npu_inst_pe_1_7_5_n9), .Q(
        npu_inst_pe_1_7_5_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_7_5_n109), 
        .CK(npu_inst_pe_1_7_5_net2896), .RN(npu_inst_pe_1_7_5_n10), .Q(
        npu_inst_pe_1_7_5_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_7_5_n108), 
        .CK(npu_inst_pe_1_7_5_net2896), .RN(npu_inst_pe_1_7_5_n10), .Q(
        npu_inst_pe_1_7_5_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_7_5_n107), 
        .CK(npu_inst_pe_1_7_5_net2896), .RN(npu_inst_pe_1_7_5_n10), .Q(
        npu_inst_pe_1_7_5_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_7_5_n106), 
        .CK(npu_inst_pe_1_7_5_net2896), .RN(npu_inst_pe_1_7_5_n10), .Q(
        npu_inst_pe_1_7_5_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_7_5_n105), 
        .CK(npu_inst_pe_1_7_5_net2896), .RN(npu_inst_pe_1_7_5_n10), .Q(
        npu_inst_pe_1_7_5_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_7_5_n104), 
        .CK(npu_inst_pe_1_7_5_net2896), .RN(npu_inst_pe_1_7_5_n10), .Q(
        npu_inst_pe_1_7_5_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_7_5_n103), 
        .CK(npu_inst_pe_1_7_5_net2896), .RN(npu_inst_pe_1_7_5_n10), .Q(
        npu_inst_pe_1_7_5_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_7_5_n102), 
        .CK(npu_inst_pe_1_7_5_net2896), .RN(npu_inst_pe_1_7_5_n10), .Q(
        npu_inst_pe_1_7_5_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_7_5_n86), 
        .CK(npu_inst_pe_1_7_5_net2896), .RN(npu_inst_pe_1_7_5_n10), .Q(
        npu_inst_pe_1_7_5_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_7_5_n87), 
        .CK(npu_inst_pe_1_7_5_net2896), .RN(npu_inst_pe_1_7_5_n10), .Q(
        npu_inst_pe_1_7_5_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_7_5_n88), 
        .CK(npu_inst_pe_1_7_5_net2896), .RN(npu_inst_pe_1_7_5_n11), .Q(
        npu_inst_pe_1_7_5_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_7_5_n89), 
        .CK(npu_inst_pe_1_7_5_net2896), .RN(npu_inst_pe_1_7_5_n11), .Q(
        npu_inst_pe_1_7_5_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_7_5_n90), 
        .CK(npu_inst_pe_1_7_5_net2896), .RN(npu_inst_pe_1_7_5_n11), .Q(
        npu_inst_pe_1_7_5_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_7_5_n91), 
        .CK(npu_inst_pe_1_7_5_net2896), .RN(npu_inst_pe_1_7_5_n11), .Q(
        npu_inst_pe_1_7_5_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_7_5_n92), 
        .CK(npu_inst_pe_1_7_5_net2896), .RN(npu_inst_pe_1_7_5_n11), .Q(
        npu_inst_pe_1_7_5_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_7_5_n93), 
        .CK(npu_inst_pe_1_7_5_net2896), .RN(npu_inst_pe_1_7_5_n11), .Q(
        npu_inst_pe_1_7_5_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_7_5_n94), 
        .CK(npu_inst_pe_1_7_5_net2896), .RN(npu_inst_pe_1_7_5_n11), .Q(
        npu_inst_pe_1_7_5_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_7_5_n95), 
        .CK(npu_inst_pe_1_7_5_net2896), .RN(npu_inst_pe_1_7_5_n11), .Q(
        npu_inst_pe_1_7_5_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_7_5_n96), 
        .CK(npu_inst_pe_1_7_5_net2896), .RN(npu_inst_pe_1_7_5_n11), .Q(
        npu_inst_pe_1_7_5_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_7_5_n97), 
        .CK(npu_inst_pe_1_7_5_net2896), .RN(npu_inst_pe_1_7_5_n11), .Q(
        npu_inst_pe_1_7_5_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_7_5_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_7_5_N84), .SE(1'b0), .GCK(npu_inst_pe_1_7_5_net2890) );
  CLKGATETST_X1 npu_inst_pe_1_7_5_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n61), .SE(1'b0), .GCK(npu_inst_pe_1_7_5_net2896) );
  MUX2_X1 npu_inst_pe_1_7_6_U162 ( .A(npu_inst_pe_1_7_6_n32), .B(
        npu_inst_pe_1_7_6_n29), .S(npu_inst_pe_1_7_6_n8), .Z(
        npu_inst_pe_1_7_6_N93) );
  MUX2_X1 npu_inst_pe_1_7_6_U161 ( .A(npu_inst_pe_1_7_6_n31), .B(
        npu_inst_pe_1_7_6_n30), .S(npu_inst_pe_1_7_6_n6), .Z(
        npu_inst_pe_1_7_6_n32) );
  MUX2_X1 npu_inst_pe_1_7_6_U160 ( .A(npu_inst_pe_1_7_6_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_7_6_int_q_reg_v_1__0_), .S(npu_inst_pe_1_7_6_n4), .Z(
        npu_inst_pe_1_7_6_n31) );
  MUX2_X1 npu_inst_pe_1_7_6_U159 ( .A(npu_inst_pe_1_7_6_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_7_6_int_q_reg_v_3__0_), .S(npu_inst_pe_1_7_6_n4), .Z(
        npu_inst_pe_1_7_6_n30) );
  MUX2_X1 npu_inst_pe_1_7_6_U158 ( .A(npu_inst_pe_1_7_6_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_7_6_int_q_reg_v_5__0_), .S(npu_inst_pe_1_7_6_n4), .Z(
        npu_inst_pe_1_7_6_n29) );
  MUX2_X1 npu_inst_pe_1_7_6_U157 ( .A(npu_inst_pe_1_7_6_n28), .B(
        npu_inst_pe_1_7_6_n23), .S(npu_inst_pe_1_7_6_n8), .Z(
        npu_inst_pe_1_7_6_N94) );
  MUX2_X1 npu_inst_pe_1_7_6_U156 ( .A(npu_inst_pe_1_7_6_n25), .B(
        npu_inst_pe_1_7_6_n24), .S(npu_inst_pe_1_7_6_n6), .Z(
        npu_inst_pe_1_7_6_n28) );
  MUX2_X1 npu_inst_pe_1_7_6_U155 ( .A(npu_inst_pe_1_7_6_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_7_6_int_q_reg_v_1__1_), .S(npu_inst_pe_1_7_6_n4), .Z(
        npu_inst_pe_1_7_6_n25) );
  MUX2_X1 npu_inst_pe_1_7_6_U154 ( .A(npu_inst_pe_1_7_6_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_7_6_int_q_reg_v_3__1_), .S(npu_inst_pe_1_7_6_n4), .Z(
        npu_inst_pe_1_7_6_n24) );
  MUX2_X1 npu_inst_pe_1_7_6_U153 ( .A(npu_inst_pe_1_7_6_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_7_6_int_q_reg_v_5__1_), .S(npu_inst_pe_1_7_6_n4), .Z(
        npu_inst_pe_1_7_6_n23) );
  MUX2_X1 npu_inst_pe_1_7_6_U152 ( .A(npu_inst_pe_1_7_6_n22), .B(
        npu_inst_pe_1_7_6_n19), .S(npu_inst_pe_1_7_6_n8), .Z(
        npu_inst_int_data_x_7__6__1_) );
  MUX2_X1 npu_inst_pe_1_7_6_U151 ( .A(npu_inst_pe_1_7_6_n21), .B(
        npu_inst_pe_1_7_6_n20), .S(npu_inst_pe_1_7_6_n6), .Z(
        npu_inst_pe_1_7_6_n22) );
  MUX2_X1 npu_inst_pe_1_7_6_U150 ( .A(npu_inst_pe_1_7_6_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_7_6_int_q_reg_h_1__1_), .S(npu_inst_pe_1_7_6_n4), .Z(
        npu_inst_pe_1_7_6_n21) );
  MUX2_X1 npu_inst_pe_1_7_6_U149 ( .A(npu_inst_pe_1_7_6_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_7_6_int_q_reg_h_3__1_), .S(npu_inst_pe_1_7_6_n4), .Z(
        npu_inst_pe_1_7_6_n20) );
  MUX2_X1 npu_inst_pe_1_7_6_U148 ( .A(npu_inst_pe_1_7_6_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_7_6_int_q_reg_h_5__1_), .S(npu_inst_pe_1_7_6_n4), .Z(
        npu_inst_pe_1_7_6_n19) );
  MUX2_X1 npu_inst_pe_1_7_6_U147 ( .A(npu_inst_pe_1_7_6_n18), .B(
        npu_inst_pe_1_7_6_n15), .S(npu_inst_pe_1_7_6_n8), .Z(
        npu_inst_int_data_x_7__6__0_) );
  MUX2_X1 npu_inst_pe_1_7_6_U146 ( .A(npu_inst_pe_1_7_6_n17), .B(
        npu_inst_pe_1_7_6_n16), .S(npu_inst_pe_1_7_6_n6), .Z(
        npu_inst_pe_1_7_6_n18) );
  MUX2_X1 npu_inst_pe_1_7_6_U145 ( .A(npu_inst_pe_1_7_6_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_7_6_int_q_reg_h_1__0_), .S(npu_inst_pe_1_7_6_n4), .Z(
        npu_inst_pe_1_7_6_n17) );
  MUX2_X1 npu_inst_pe_1_7_6_U144 ( .A(npu_inst_pe_1_7_6_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_7_6_int_q_reg_h_3__0_), .S(npu_inst_pe_1_7_6_n4), .Z(
        npu_inst_pe_1_7_6_n16) );
  MUX2_X1 npu_inst_pe_1_7_6_U143 ( .A(npu_inst_pe_1_7_6_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_7_6_int_q_reg_h_5__0_), .S(npu_inst_pe_1_7_6_n4), .Z(
        npu_inst_pe_1_7_6_n15) );
  XOR2_X1 npu_inst_pe_1_7_6_U142 ( .A(npu_inst_pe_1_7_6_int_data_0_), .B(
        npu_inst_pe_1_7_6_int_q_acc_0_), .Z(npu_inst_pe_1_7_6_N73) );
  AND2_X1 npu_inst_pe_1_7_6_U141 ( .A1(npu_inst_pe_1_7_6_int_q_acc_0_), .A2(
        npu_inst_pe_1_7_6_int_data_0_), .ZN(npu_inst_pe_1_7_6_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_7_6_U140 ( .A(npu_inst_pe_1_7_6_int_q_acc_0_), .B(
        npu_inst_pe_1_7_6_n13), .ZN(npu_inst_pe_1_7_6_N65) );
  OR2_X1 npu_inst_pe_1_7_6_U139 ( .A1(npu_inst_pe_1_7_6_n13), .A2(
        npu_inst_pe_1_7_6_int_q_acc_0_), .ZN(npu_inst_pe_1_7_6_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_7_6_U138 ( .A(npu_inst_pe_1_7_6_int_q_acc_2_), .B(
        npu_inst_pe_1_7_6_add_79_carry_2_), .Z(npu_inst_pe_1_7_6_N75) );
  AND2_X1 npu_inst_pe_1_7_6_U137 ( .A1(npu_inst_pe_1_7_6_add_79_carry_2_), 
        .A2(npu_inst_pe_1_7_6_int_q_acc_2_), .ZN(
        npu_inst_pe_1_7_6_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_7_6_U136 ( .A(npu_inst_pe_1_7_6_int_q_acc_3_), .B(
        npu_inst_pe_1_7_6_add_79_carry_3_), .Z(npu_inst_pe_1_7_6_N76) );
  AND2_X1 npu_inst_pe_1_7_6_U135 ( .A1(npu_inst_pe_1_7_6_add_79_carry_3_), 
        .A2(npu_inst_pe_1_7_6_int_q_acc_3_), .ZN(
        npu_inst_pe_1_7_6_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_7_6_U134 ( .A(npu_inst_pe_1_7_6_int_q_acc_4_), .B(
        npu_inst_pe_1_7_6_add_79_carry_4_), .Z(npu_inst_pe_1_7_6_N77) );
  AND2_X1 npu_inst_pe_1_7_6_U133 ( .A1(npu_inst_pe_1_7_6_add_79_carry_4_), 
        .A2(npu_inst_pe_1_7_6_int_q_acc_4_), .ZN(
        npu_inst_pe_1_7_6_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_7_6_U132 ( .A(npu_inst_pe_1_7_6_int_q_acc_5_), .B(
        npu_inst_pe_1_7_6_add_79_carry_5_), .Z(npu_inst_pe_1_7_6_N78) );
  AND2_X1 npu_inst_pe_1_7_6_U131 ( .A1(npu_inst_pe_1_7_6_add_79_carry_5_), 
        .A2(npu_inst_pe_1_7_6_int_q_acc_5_), .ZN(
        npu_inst_pe_1_7_6_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_7_6_U130 ( .A(npu_inst_pe_1_7_6_int_q_acc_6_), .B(
        npu_inst_pe_1_7_6_add_79_carry_6_), .Z(npu_inst_pe_1_7_6_N79) );
  AND2_X1 npu_inst_pe_1_7_6_U129 ( .A1(npu_inst_pe_1_7_6_add_79_carry_6_), 
        .A2(npu_inst_pe_1_7_6_int_q_acc_6_), .ZN(
        npu_inst_pe_1_7_6_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_7_6_U128 ( .A(npu_inst_pe_1_7_6_int_q_acc_7_), .B(
        npu_inst_pe_1_7_6_add_79_carry_7_), .Z(npu_inst_pe_1_7_6_N80) );
  XNOR2_X1 npu_inst_pe_1_7_6_U127 ( .A(npu_inst_pe_1_7_6_sub_77_carry_2_), .B(
        npu_inst_pe_1_7_6_int_q_acc_2_), .ZN(npu_inst_pe_1_7_6_N67) );
  OR2_X1 npu_inst_pe_1_7_6_U126 ( .A1(npu_inst_pe_1_7_6_int_q_acc_2_), .A2(
        npu_inst_pe_1_7_6_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_7_6_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_7_6_U125 ( .A(npu_inst_pe_1_7_6_sub_77_carry_3_), .B(
        npu_inst_pe_1_7_6_int_q_acc_3_), .ZN(npu_inst_pe_1_7_6_N68) );
  OR2_X1 npu_inst_pe_1_7_6_U124 ( .A1(npu_inst_pe_1_7_6_int_q_acc_3_), .A2(
        npu_inst_pe_1_7_6_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_7_6_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_7_6_U123 ( .A(npu_inst_pe_1_7_6_sub_77_carry_4_), .B(
        npu_inst_pe_1_7_6_int_q_acc_4_), .ZN(npu_inst_pe_1_7_6_N69) );
  OR2_X1 npu_inst_pe_1_7_6_U122 ( .A1(npu_inst_pe_1_7_6_int_q_acc_4_), .A2(
        npu_inst_pe_1_7_6_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_7_6_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_7_6_U121 ( .A(npu_inst_pe_1_7_6_sub_77_carry_5_), .B(
        npu_inst_pe_1_7_6_int_q_acc_5_), .ZN(npu_inst_pe_1_7_6_N70) );
  OR2_X1 npu_inst_pe_1_7_6_U120 ( .A1(npu_inst_pe_1_7_6_int_q_acc_5_), .A2(
        npu_inst_pe_1_7_6_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_7_6_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_7_6_U119 ( .A(npu_inst_pe_1_7_6_sub_77_carry_6_), .B(
        npu_inst_pe_1_7_6_int_q_acc_6_), .ZN(npu_inst_pe_1_7_6_N71) );
  OR2_X1 npu_inst_pe_1_7_6_U118 ( .A1(npu_inst_pe_1_7_6_int_q_acc_6_), .A2(
        npu_inst_pe_1_7_6_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_7_6_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_7_6_U117 ( .A(npu_inst_pe_1_7_6_int_q_acc_7_), .B(
        npu_inst_pe_1_7_6_sub_77_carry_7_), .ZN(npu_inst_pe_1_7_6_N72) );
  INV_X1 npu_inst_pe_1_7_6_U116 ( .A(npu_inst_n75), .ZN(npu_inst_pe_1_7_6_n7)
         );
  INV_X1 npu_inst_pe_1_7_6_U115 ( .A(npu_inst_pe_1_7_6_n7), .ZN(
        npu_inst_pe_1_7_6_n6) );
  INV_X1 npu_inst_pe_1_7_6_U114 ( .A(npu_inst_n52), .ZN(npu_inst_pe_1_7_6_n3)
         );
  AOI22_X1 npu_inst_pe_1_7_6_U113 ( .A1(npu_inst_pe_1_7_6_n38), .A2(
        int_i_data_v_npu[3]), .B1(npu_inst_pe_1_7_6_n118), .B2(
        npu_inst_pe_1_7_6_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_7_6_n39) );
  INV_X1 npu_inst_pe_1_7_6_U112 ( .A(npu_inst_pe_1_7_6_n39), .ZN(
        npu_inst_pe_1_7_6_n112) );
  AOI22_X1 npu_inst_pe_1_7_6_U111 ( .A1(npu_inst_pe_1_7_6_n38), .A2(
        int_i_data_v_npu[2]), .B1(npu_inst_pe_1_7_6_n118), .B2(
        npu_inst_pe_1_7_6_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_7_6_n37) );
  INV_X1 npu_inst_pe_1_7_6_U110 ( .A(npu_inst_pe_1_7_6_n37), .ZN(
        npu_inst_pe_1_7_6_n113) );
  AOI22_X1 npu_inst_pe_1_7_6_U107 ( .A1(int_i_data_v_npu[3]), .A2(
        npu_inst_pe_1_7_6_n58), .B1(npu_inst_pe_1_7_6_n114), .B2(
        npu_inst_pe_1_7_6_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_7_6_n59) );
  INV_X1 npu_inst_pe_1_7_6_U106 ( .A(npu_inst_pe_1_7_6_n59), .ZN(
        npu_inst_pe_1_7_6_n102) );
  AOI22_X1 npu_inst_pe_1_7_6_U105 ( .A1(int_i_data_v_npu[2]), .A2(
        npu_inst_pe_1_7_6_n58), .B1(npu_inst_pe_1_7_6_n114), .B2(
        npu_inst_pe_1_7_6_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_7_6_n57) );
  INV_X1 npu_inst_pe_1_7_6_U104 ( .A(npu_inst_pe_1_7_6_n57), .ZN(
        npu_inst_pe_1_7_6_n103) );
  AOI22_X1 npu_inst_pe_1_7_6_U103 ( .A1(int_i_data_v_npu[3]), .A2(
        npu_inst_pe_1_7_6_n54), .B1(npu_inst_pe_1_7_6_n115), .B2(
        npu_inst_pe_1_7_6_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_7_6_n55) );
  INV_X1 npu_inst_pe_1_7_6_U102 ( .A(npu_inst_pe_1_7_6_n55), .ZN(
        npu_inst_pe_1_7_6_n104) );
  AOI22_X1 npu_inst_pe_1_7_6_U101 ( .A1(int_i_data_v_npu[2]), .A2(
        npu_inst_pe_1_7_6_n54), .B1(npu_inst_pe_1_7_6_n115), .B2(
        npu_inst_pe_1_7_6_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_7_6_n53) );
  INV_X1 npu_inst_pe_1_7_6_U100 ( .A(npu_inst_pe_1_7_6_n53), .ZN(
        npu_inst_pe_1_7_6_n105) );
  AOI22_X1 npu_inst_pe_1_7_6_U99 ( .A1(int_i_data_v_npu[3]), .A2(
        npu_inst_pe_1_7_6_n50), .B1(npu_inst_pe_1_7_6_n116), .B2(
        npu_inst_pe_1_7_6_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_7_6_n51) );
  INV_X1 npu_inst_pe_1_7_6_U98 ( .A(npu_inst_pe_1_7_6_n51), .ZN(
        npu_inst_pe_1_7_6_n106) );
  AOI22_X1 npu_inst_pe_1_7_6_U97 ( .A1(int_i_data_v_npu[2]), .A2(
        npu_inst_pe_1_7_6_n50), .B1(npu_inst_pe_1_7_6_n116), .B2(
        npu_inst_pe_1_7_6_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_7_6_n49) );
  INV_X1 npu_inst_pe_1_7_6_U96 ( .A(npu_inst_pe_1_7_6_n49), .ZN(
        npu_inst_pe_1_7_6_n107) );
  AOI22_X1 npu_inst_pe_1_7_6_U95 ( .A1(int_i_data_v_npu[3]), .A2(
        npu_inst_pe_1_7_6_n46), .B1(npu_inst_pe_1_7_6_n117), .B2(
        npu_inst_pe_1_7_6_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_7_6_n47) );
  INV_X1 npu_inst_pe_1_7_6_U94 ( .A(npu_inst_pe_1_7_6_n47), .ZN(
        npu_inst_pe_1_7_6_n108) );
  AOI22_X1 npu_inst_pe_1_7_6_U93 ( .A1(int_i_data_v_npu[2]), .A2(
        npu_inst_pe_1_7_6_n46), .B1(npu_inst_pe_1_7_6_n117), .B2(
        npu_inst_pe_1_7_6_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_7_6_n45) );
  INV_X1 npu_inst_pe_1_7_6_U92 ( .A(npu_inst_pe_1_7_6_n45), .ZN(
        npu_inst_pe_1_7_6_n109) );
  AOI22_X1 npu_inst_pe_1_7_6_U91 ( .A1(int_i_data_v_npu[3]), .A2(
        npu_inst_pe_1_7_6_n42), .B1(npu_inst_pe_1_7_6_n119), .B2(
        npu_inst_pe_1_7_6_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_7_6_n43) );
  INV_X1 npu_inst_pe_1_7_6_U90 ( .A(npu_inst_pe_1_7_6_n43), .ZN(
        npu_inst_pe_1_7_6_n110) );
  AOI22_X1 npu_inst_pe_1_7_6_U89 ( .A1(int_i_data_v_npu[2]), .A2(
        npu_inst_pe_1_7_6_n42), .B1(npu_inst_pe_1_7_6_n119), .B2(
        npu_inst_pe_1_7_6_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_7_6_n41) );
  INV_X1 npu_inst_pe_1_7_6_U88 ( .A(npu_inst_pe_1_7_6_n41), .ZN(
        npu_inst_pe_1_7_6_n111) );
  NAND2_X1 npu_inst_pe_1_7_6_U87 ( .A1(npu_inst_pe_1_7_6_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_7_6_n60), .ZN(npu_inst_pe_1_7_6_n74) );
  OAI21_X1 npu_inst_pe_1_7_6_U86 ( .B1(npu_inst_pe_1_7_6_n63), .B2(
        npu_inst_pe_1_7_6_n60), .A(npu_inst_pe_1_7_6_n74), .ZN(
        npu_inst_pe_1_7_6_n97) );
  NAND2_X1 npu_inst_pe_1_7_6_U85 ( .A1(npu_inst_pe_1_7_6_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_7_6_n60), .ZN(npu_inst_pe_1_7_6_n73) );
  OAI21_X1 npu_inst_pe_1_7_6_U84 ( .B1(npu_inst_pe_1_7_6_n61), .B2(
        npu_inst_pe_1_7_6_n60), .A(npu_inst_pe_1_7_6_n73), .ZN(
        npu_inst_pe_1_7_6_n96) );
  NAND2_X1 npu_inst_pe_1_7_6_U83 ( .A1(npu_inst_pe_1_7_6_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_7_6_n56), .ZN(npu_inst_pe_1_7_6_n72) );
  OAI21_X1 npu_inst_pe_1_7_6_U82 ( .B1(npu_inst_pe_1_7_6_n63), .B2(
        npu_inst_pe_1_7_6_n56), .A(npu_inst_pe_1_7_6_n72), .ZN(
        npu_inst_pe_1_7_6_n95) );
  NAND2_X1 npu_inst_pe_1_7_6_U81 ( .A1(npu_inst_pe_1_7_6_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_7_6_n56), .ZN(npu_inst_pe_1_7_6_n71) );
  OAI21_X1 npu_inst_pe_1_7_6_U80 ( .B1(npu_inst_pe_1_7_6_n61), .B2(
        npu_inst_pe_1_7_6_n56), .A(npu_inst_pe_1_7_6_n71), .ZN(
        npu_inst_pe_1_7_6_n94) );
  NAND2_X1 npu_inst_pe_1_7_6_U79 ( .A1(npu_inst_pe_1_7_6_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_7_6_n52), .ZN(npu_inst_pe_1_7_6_n70) );
  OAI21_X1 npu_inst_pe_1_7_6_U78 ( .B1(npu_inst_pe_1_7_6_n63), .B2(
        npu_inst_pe_1_7_6_n52), .A(npu_inst_pe_1_7_6_n70), .ZN(
        npu_inst_pe_1_7_6_n93) );
  NAND2_X1 npu_inst_pe_1_7_6_U77 ( .A1(npu_inst_pe_1_7_6_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_7_6_n52), .ZN(npu_inst_pe_1_7_6_n69) );
  OAI21_X1 npu_inst_pe_1_7_6_U76 ( .B1(npu_inst_pe_1_7_6_n61), .B2(
        npu_inst_pe_1_7_6_n52), .A(npu_inst_pe_1_7_6_n69), .ZN(
        npu_inst_pe_1_7_6_n92) );
  NAND2_X1 npu_inst_pe_1_7_6_U75 ( .A1(npu_inst_pe_1_7_6_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_7_6_n48), .ZN(npu_inst_pe_1_7_6_n68) );
  OAI21_X1 npu_inst_pe_1_7_6_U74 ( .B1(npu_inst_pe_1_7_6_n63), .B2(
        npu_inst_pe_1_7_6_n48), .A(npu_inst_pe_1_7_6_n68), .ZN(
        npu_inst_pe_1_7_6_n91) );
  NAND2_X1 npu_inst_pe_1_7_6_U73 ( .A1(npu_inst_pe_1_7_6_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_7_6_n48), .ZN(npu_inst_pe_1_7_6_n67) );
  OAI21_X1 npu_inst_pe_1_7_6_U72 ( .B1(npu_inst_pe_1_7_6_n61), .B2(
        npu_inst_pe_1_7_6_n48), .A(npu_inst_pe_1_7_6_n67), .ZN(
        npu_inst_pe_1_7_6_n90) );
  NAND2_X1 npu_inst_pe_1_7_6_U71 ( .A1(npu_inst_pe_1_7_6_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_7_6_n44), .ZN(npu_inst_pe_1_7_6_n66) );
  OAI21_X1 npu_inst_pe_1_7_6_U70 ( .B1(npu_inst_pe_1_7_6_n63), .B2(
        npu_inst_pe_1_7_6_n44), .A(npu_inst_pe_1_7_6_n66), .ZN(
        npu_inst_pe_1_7_6_n89) );
  NAND2_X1 npu_inst_pe_1_7_6_U69 ( .A1(npu_inst_pe_1_7_6_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_7_6_n44), .ZN(npu_inst_pe_1_7_6_n65) );
  OAI21_X1 npu_inst_pe_1_7_6_U68 ( .B1(npu_inst_pe_1_7_6_n61), .B2(
        npu_inst_pe_1_7_6_n44), .A(npu_inst_pe_1_7_6_n65), .ZN(
        npu_inst_pe_1_7_6_n88) );
  NAND2_X1 npu_inst_pe_1_7_6_U67 ( .A1(npu_inst_pe_1_7_6_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_7_6_n40), .ZN(npu_inst_pe_1_7_6_n64) );
  OAI21_X1 npu_inst_pe_1_7_6_U66 ( .B1(npu_inst_pe_1_7_6_n63), .B2(
        npu_inst_pe_1_7_6_n40), .A(npu_inst_pe_1_7_6_n64), .ZN(
        npu_inst_pe_1_7_6_n87) );
  NAND2_X1 npu_inst_pe_1_7_6_U65 ( .A1(npu_inst_pe_1_7_6_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_7_6_n40), .ZN(npu_inst_pe_1_7_6_n62) );
  OAI21_X1 npu_inst_pe_1_7_6_U64 ( .B1(npu_inst_pe_1_7_6_n61), .B2(
        npu_inst_pe_1_7_6_n40), .A(npu_inst_pe_1_7_6_n62), .ZN(
        npu_inst_pe_1_7_6_n86) );
  AND2_X1 npu_inst_pe_1_7_6_U63 ( .A1(npu_inst_pe_1_7_6_N93), .A2(npu_inst_n52), .ZN(npu_inst_int_data_y_7__6__0_) );
  AND2_X1 npu_inst_pe_1_7_6_U62 ( .A1(npu_inst_n52), .A2(npu_inst_pe_1_7_6_N94), .ZN(npu_inst_int_data_y_7__6__1_) );
  AOI22_X1 npu_inst_pe_1_7_6_U61 ( .A1(npu_inst_n52), .A2(int_i_data_v_npu[3]), 
        .B1(npu_inst_pe_1_7_6_n3), .B2(npu_inst_int_data_x_7__7__1_), .ZN(
        npu_inst_pe_1_7_6_n63) );
  AOI22_X1 npu_inst_pe_1_7_6_U60 ( .A1(npu_inst_n52), .A2(int_i_data_v_npu[2]), 
        .B1(npu_inst_pe_1_7_6_n3), .B2(npu_inst_int_data_x_7__7__0_), .ZN(
        npu_inst_pe_1_7_6_n61) );
  NOR3_X1 npu_inst_pe_1_7_6_U59 ( .A1(npu_inst_pe_1_7_6_n26), .A2(npu_inst_n52), .A3(npu_inst_int_ckg[1]), .ZN(npu_inst_pe_1_7_6_n85) );
  OR2_X1 npu_inst_pe_1_7_6_U58 ( .A1(npu_inst_pe_1_7_6_n85), .A2(
        npu_inst_pe_1_7_6_n2), .ZN(npu_inst_pe_1_7_6_N84) );
  AOI222_X1 npu_inst_pe_1_7_6_U57 ( .A1(1'b0), .A2(npu_inst_pe_1_7_6_n1), .B1(
        npu_inst_pe_1_7_6_N73), .B2(npu_inst_pe_1_7_6_n76), .C1(
        npu_inst_pe_1_7_6_N65), .C2(npu_inst_pe_1_7_6_n77), .ZN(
        npu_inst_pe_1_7_6_n84) );
  INV_X1 npu_inst_pe_1_7_6_U56 ( .A(npu_inst_pe_1_7_6_n84), .ZN(
        npu_inst_pe_1_7_6_n101) );
  AOI222_X1 npu_inst_pe_1_7_6_U55 ( .A1(1'b0), .A2(npu_inst_pe_1_7_6_n1), .B1(
        npu_inst_pe_1_7_6_N80), .B2(npu_inst_pe_1_7_6_n76), .C1(
        npu_inst_pe_1_7_6_N72), .C2(npu_inst_pe_1_7_6_n77), .ZN(
        npu_inst_pe_1_7_6_n75) );
  INV_X1 npu_inst_pe_1_7_6_U54 ( .A(npu_inst_pe_1_7_6_n75), .ZN(
        npu_inst_pe_1_7_6_n33) );
  AOI222_X1 npu_inst_pe_1_7_6_U53 ( .A1(1'b0), .A2(npu_inst_pe_1_7_6_n1), .B1(
        npu_inst_pe_1_7_6_N74), .B2(npu_inst_pe_1_7_6_n76), .C1(
        npu_inst_pe_1_7_6_N66), .C2(npu_inst_pe_1_7_6_n77), .ZN(
        npu_inst_pe_1_7_6_n83) );
  INV_X1 npu_inst_pe_1_7_6_U52 ( .A(npu_inst_pe_1_7_6_n83), .ZN(
        npu_inst_pe_1_7_6_n100) );
  AOI222_X1 npu_inst_pe_1_7_6_U51 ( .A1(1'b0), .A2(npu_inst_pe_1_7_6_n1), .B1(
        npu_inst_pe_1_7_6_N75), .B2(npu_inst_pe_1_7_6_n76), .C1(
        npu_inst_pe_1_7_6_N67), .C2(npu_inst_pe_1_7_6_n77), .ZN(
        npu_inst_pe_1_7_6_n82) );
  INV_X1 npu_inst_pe_1_7_6_U50 ( .A(npu_inst_pe_1_7_6_n82), .ZN(
        npu_inst_pe_1_7_6_n99) );
  AOI222_X1 npu_inst_pe_1_7_6_U49 ( .A1(1'b0), .A2(npu_inst_pe_1_7_6_n1), .B1(
        npu_inst_pe_1_7_6_N76), .B2(npu_inst_pe_1_7_6_n76), .C1(
        npu_inst_pe_1_7_6_N68), .C2(npu_inst_pe_1_7_6_n77), .ZN(
        npu_inst_pe_1_7_6_n81) );
  INV_X1 npu_inst_pe_1_7_6_U48 ( .A(npu_inst_pe_1_7_6_n81), .ZN(
        npu_inst_pe_1_7_6_n98) );
  AOI222_X1 npu_inst_pe_1_7_6_U47 ( .A1(1'b0), .A2(npu_inst_pe_1_7_6_n1), .B1(
        npu_inst_pe_1_7_6_N77), .B2(npu_inst_pe_1_7_6_n76), .C1(
        npu_inst_pe_1_7_6_N69), .C2(npu_inst_pe_1_7_6_n77), .ZN(
        npu_inst_pe_1_7_6_n80) );
  INV_X1 npu_inst_pe_1_7_6_U46 ( .A(npu_inst_pe_1_7_6_n80), .ZN(
        npu_inst_pe_1_7_6_n36) );
  AOI222_X1 npu_inst_pe_1_7_6_U45 ( .A1(1'b0), .A2(npu_inst_pe_1_7_6_n1), .B1(
        npu_inst_pe_1_7_6_N78), .B2(npu_inst_pe_1_7_6_n76), .C1(
        npu_inst_pe_1_7_6_N70), .C2(npu_inst_pe_1_7_6_n77), .ZN(
        npu_inst_pe_1_7_6_n79) );
  INV_X1 npu_inst_pe_1_7_6_U44 ( .A(npu_inst_pe_1_7_6_n79), .ZN(
        npu_inst_pe_1_7_6_n35) );
  AOI222_X1 npu_inst_pe_1_7_6_U43 ( .A1(1'b0), .A2(npu_inst_pe_1_7_6_n1), .B1(
        npu_inst_pe_1_7_6_N79), .B2(npu_inst_pe_1_7_6_n76), .C1(
        npu_inst_pe_1_7_6_N71), .C2(npu_inst_pe_1_7_6_n77), .ZN(
        npu_inst_pe_1_7_6_n78) );
  INV_X1 npu_inst_pe_1_7_6_U42 ( .A(npu_inst_pe_1_7_6_n78), .ZN(
        npu_inst_pe_1_7_6_n34) );
  AND2_X1 npu_inst_pe_1_7_6_U41 ( .A1(npu_inst_pe_1_7_6_int_q_acc_0_), .A2(
        npu_inst_pe_1_7_6_n1), .ZN(npu_inst_int_data_res_7__6__0_) );
  AND2_X1 npu_inst_pe_1_7_6_U40 ( .A1(npu_inst_pe_1_7_6_n2), .A2(
        npu_inst_pe_1_7_6_int_q_acc_7_), .ZN(npu_inst_int_data_res_7__6__7_)
         );
  AND2_X1 npu_inst_pe_1_7_6_U39 ( .A1(npu_inst_pe_1_7_6_int_q_acc_1_), .A2(
        npu_inst_pe_1_7_6_n1), .ZN(npu_inst_int_data_res_7__6__1_) );
  AND2_X1 npu_inst_pe_1_7_6_U38 ( .A1(npu_inst_pe_1_7_6_int_q_acc_2_), .A2(
        npu_inst_pe_1_7_6_n1), .ZN(npu_inst_int_data_res_7__6__2_) );
  AND2_X1 npu_inst_pe_1_7_6_U37 ( .A1(npu_inst_pe_1_7_6_int_q_acc_3_), .A2(
        npu_inst_pe_1_7_6_n2), .ZN(npu_inst_int_data_res_7__6__3_) );
  AND2_X1 npu_inst_pe_1_7_6_U36 ( .A1(npu_inst_pe_1_7_6_int_q_acc_4_), .A2(
        npu_inst_pe_1_7_6_n2), .ZN(npu_inst_int_data_res_7__6__4_) );
  AND2_X1 npu_inst_pe_1_7_6_U35 ( .A1(npu_inst_pe_1_7_6_int_q_acc_5_), .A2(
        npu_inst_pe_1_7_6_n2), .ZN(npu_inst_int_data_res_7__6__5_) );
  AND2_X1 npu_inst_pe_1_7_6_U34 ( .A1(npu_inst_pe_1_7_6_int_q_acc_6_), .A2(
        npu_inst_pe_1_7_6_n2), .ZN(npu_inst_int_data_res_7__6__6_) );
  INV_X1 npu_inst_pe_1_7_6_U33 ( .A(npu_inst_pe_1_7_6_int_data_1_), .ZN(
        npu_inst_pe_1_7_6_n14) );
  AND2_X1 npu_inst_pe_1_7_6_U32 ( .A1(npu_inst_int_data_x_7__6__1_), .A2(
        npu_inst_pe_1_7_6_int_q_weight_1_), .ZN(npu_inst_pe_1_7_6_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_7_6_U31 ( .A1(npu_inst_int_data_x_7__6__0_), .A2(
        npu_inst_pe_1_7_6_int_q_weight_1_), .ZN(npu_inst_pe_1_7_6_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_7_6_U30 ( .A(npu_inst_pe_1_7_6_int_data_0_), .ZN(
        npu_inst_pe_1_7_6_n13) );
  INV_X1 npu_inst_pe_1_7_6_U29 ( .A(npu_inst_n67), .ZN(npu_inst_pe_1_7_6_n5)
         );
  OR3_X1 npu_inst_pe_1_7_6_U28 ( .A1(npu_inst_pe_1_7_6_n6), .A2(
        npu_inst_pe_1_7_6_n8), .A3(npu_inst_pe_1_7_6_n5), .ZN(
        npu_inst_pe_1_7_6_n56) );
  OR3_X1 npu_inst_pe_1_7_6_U27 ( .A1(npu_inst_pe_1_7_6_n5), .A2(
        npu_inst_pe_1_7_6_n8), .A3(npu_inst_pe_1_7_6_n7), .ZN(
        npu_inst_pe_1_7_6_n48) );
  INV_X1 npu_inst_pe_1_7_6_U26 ( .A(npu_inst_pe_1_7_6_n5), .ZN(
        npu_inst_pe_1_7_6_n4) );
  INV_X1 npu_inst_pe_1_7_6_U25 ( .A(npu_inst_n122), .ZN(npu_inst_pe_1_7_6_n12)
         );
  OR3_X1 npu_inst_pe_1_7_6_U24 ( .A1(npu_inst_pe_1_7_6_n4), .A2(
        npu_inst_pe_1_7_6_n8), .A3(npu_inst_pe_1_7_6_n7), .ZN(
        npu_inst_pe_1_7_6_n52) );
  OR3_X1 npu_inst_pe_1_7_6_U23 ( .A1(npu_inst_pe_1_7_6_n6), .A2(
        npu_inst_pe_1_7_6_n8), .A3(npu_inst_pe_1_7_6_n4), .ZN(
        npu_inst_pe_1_7_6_n60) );
  NOR2_X1 npu_inst_pe_1_7_6_U22 ( .A1(npu_inst_pe_1_7_6_n60), .A2(
        npu_inst_pe_1_7_6_n3), .ZN(npu_inst_pe_1_7_6_n58) );
  NOR2_X1 npu_inst_pe_1_7_6_U21 ( .A1(npu_inst_pe_1_7_6_n56), .A2(
        npu_inst_pe_1_7_6_n3), .ZN(npu_inst_pe_1_7_6_n54) );
  NOR2_X1 npu_inst_pe_1_7_6_U20 ( .A1(npu_inst_pe_1_7_6_n52), .A2(
        npu_inst_pe_1_7_6_n3), .ZN(npu_inst_pe_1_7_6_n50) );
  NOR2_X1 npu_inst_pe_1_7_6_U19 ( .A1(npu_inst_pe_1_7_6_n48), .A2(
        npu_inst_pe_1_7_6_n3), .ZN(npu_inst_pe_1_7_6_n46) );
  NOR2_X1 npu_inst_pe_1_7_6_U18 ( .A1(npu_inst_pe_1_7_6_n40), .A2(
        npu_inst_pe_1_7_6_n3), .ZN(npu_inst_pe_1_7_6_n38) );
  NOR2_X1 npu_inst_pe_1_7_6_U17 ( .A1(npu_inst_pe_1_7_6_n44), .A2(
        npu_inst_pe_1_7_6_n3), .ZN(npu_inst_pe_1_7_6_n42) );
  BUF_X1 npu_inst_pe_1_7_6_U16 ( .A(npu_inst_n92), .Z(npu_inst_pe_1_7_6_n8) );
  BUF_X1 npu_inst_pe_1_7_6_U15 ( .A(npu_inst_pe_1_7_6_n12), .Z(
        npu_inst_pe_1_7_6_n11) );
  BUF_X1 npu_inst_pe_1_7_6_U14 ( .A(npu_inst_pe_1_7_6_n12), .Z(
        npu_inst_pe_1_7_6_n10) );
  BUF_X1 npu_inst_pe_1_7_6_U13 ( .A(npu_inst_pe_1_7_6_n12), .Z(
        npu_inst_pe_1_7_6_n9) );
  INV_X1 npu_inst_pe_1_7_6_U12 ( .A(npu_inst_pe_1_7_6_n38), .ZN(
        npu_inst_pe_1_7_6_n118) );
  INV_X1 npu_inst_pe_1_7_6_U11 ( .A(npu_inst_pe_1_7_6_n58), .ZN(
        npu_inst_pe_1_7_6_n114) );
  INV_X1 npu_inst_pe_1_7_6_U10 ( .A(npu_inst_pe_1_7_6_n54), .ZN(
        npu_inst_pe_1_7_6_n115) );
  INV_X1 npu_inst_pe_1_7_6_U9 ( .A(npu_inst_pe_1_7_6_n50), .ZN(
        npu_inst_pe_1_7_6_n116) );
  INV_X1 npu_inst_pe_1_7_6_U8 ( .A(npu_inst_pe_1_7_6_n46), .ZN(
        npu_inst_pe_1_7_6_n117) );
  INV_X1 npu_inst_pe_1_7_6_U7 ( .A(npu_inst_pe_1_7_6_n42), .ZN(
        npu_inst_pe_1_7_6_n119) );
  BUF_X1 npu_inst_pe_1_7_6_U6 ( .A(npu_inst_n7), .Z(npu_inst_pe_1_7_6_n2) );
  BUF_X1 npu_inst_pe_1_7_6_U5 ( .A(npu_inst_n7), .Z(npu_inst_pe_1_7_6_n1) );
  NOR2_X1 npu_inst_pe_1_7_6_U4 ( .A1(npu_inst_pe_1_7_6_int_q_weight_0_), .A2(
        npu_inst_pe_1_7_6_n1), .ZN(npu_inst_pe_1_7_6_n76) );
  NOR2_X1 npu_inst_pe_1_7_6_U3 ( .A1(npu_inst_pe_1_7_6_n27), .A2(
        npu_inst_pe_1_7_6_n1), .ZN(npu_inst_pe_1_7_6_n77) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_7_6_n111), 
        .CK(npu_inst_pe_1_7_6_net2873), .RN(npu_inst_pe_1_7_6_n12), .Q(
        npu_inst_pe_1_7_6_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_7_6_n110), 
        .CK(npu_inst_pe_1_7_6_net2873), .RN(npu_inst_pe_1_7_6_n12), .Q(
        npu_inst_pe_1_7_6_int_q_reg_v_4__1_) );
  FA_X1 npu_inst_pe_1_7_6_sub_77_U2_1 ( .A(npu_inst_pe_1_7_6_int_q_acc_1_), 
        .B(npu_inst_pe_1_7_6_n14), .CI(npu_inst_pe_1_7_6_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_7_6_sub_77_carry_2_), .S(npu_inst_pe_1_7_6_N66) );
  FA_X1 npu_inst_pe_1_7_6_add_79_U1_1 ( .A(npu_inst_pe_1_7_6_int_q_acc_1_), 
        .B(npu_inst_pe_1_7_6_int_data_1_), .CI(
        npu_inst_pe_1_7_6_add_79_carry_1_), .CO(
        npu_inst_pe_1_7_6_add_79_carry_2_), .S(npu_inst_pe_1_7_6_N74) );
  NAND3_X1 npu_inst_pe_1_7_6_U109 ( .A1(npu_inst_pe_1_7_6_n5), .A2(
        npu_inst_pe_1_7_6_n7), .A3(npu_inst_pe_1_7_6_n8), .ZN(
        npu_inst_pe_1_7_6_n44) );
  NAND3_X1 npu_inst_pe_1_7_6_U108 ( .A1(npu_inst_pe_1_7_6_n4), .A2(
        npu_inst_pe_1_7_6_n7), .A3(npu_inst_pe_1_7_6_n8), .ZN(
        npu_inst_pe_1_7_6_n40) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_7_6_n34), .CK(
        npu_inst_pe_1_7_6_net2867), .RN(npu_inst_pe_1_7_6_n9), .Q(
        npu_inst_pe_1_7_6_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_7_6_n35), .CK(
        npu_inst_pe_1_7_6_net2867), .RN(npu_inst_pe_1_7_6_n9), .Q(
        npu_inst_pe_1_7_6_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_7_6_n36), .CK(
        npu_inst_pe_1_7_6_net2867), .RN(npu_inst_pe_1_7_6_n9), .Q(
        npu_inst_pe_1_7_6_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_7_6_n98), .CK(
        npu_inst_pe_1_7_6_net2867), .RN(npu_inst_pe_1_7_6_n9), .Q(
        npu_inst_pe_1_7_6_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_7_6_n99), .CK(
        npu_inst_pe_1_7_6_net2867), .RN(npu_inst_pe_1_7_6_n9), .Q(
        npu_inst_pe_1_7_6_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_7_6_n100), 
        .CK(npu_inst_pe_1_7_6_net2867), .RN(npu_inst_pe_1_7_6_n9), .Q(
        npu_inst_pe_1_7_6_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_7_6_n33), .CK(
        npu_inst_pe_1_7_6_net2867), .RN(npu_inst_pe_1_7_6_n9), .Q(
        npu_inst_pe_1_7_6_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_7_6_n101), 
        .CK(npu_inst_pe_1_7_6_net2867), .RN(npu_inst_pe_1_7_6_n9), .Q(
        npu_inst_pe_1_7_6_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_weight_reg_0_ ( .D(npu_inst_n108), .CK(
        npu_inst_pe_1_7_6_net2873), .RN(npu_inst_pe_1_7_6_n9), .Q(
        npu_inst_pe_1_7_6_int_q_weight_0_), .QN(npu_inst_pe_1_7_6_n27) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_weight_reg_1_ ( .D(npu_inst_n114), .CK(
        npu_inst_pe_1_7_6_net2873), .RN(npu_inst_pe_1_7_6_n9), .Q(
        npu_inst_pe_1_7_6_int_q_weight_1_), .QN(npu_inst_pe_1_7_6_n26) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_7_6_n113), 
        .CK(npu_inst_pe_1_7_6_net2873), .RN(npu_inst_pe_1_7_6_n9), .Q(
        npu_inst_pe_1_7_6_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_7_6_n112), 
        .CK(npu_inst_pe_1_7_6_net2873), .RN(npu_inst_pe_1_7_6_n9), .Q(
        npu_inst_pe_1_7_6_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_7_6_n109), 
        .CK(npu_inst_pe_1_7_6_net2873), .RN(npu_inst_pe_1_7_6_n10), .Q(
        npu_inst_pe_1_7_6_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_7_6_n108), 
        .CK(npu_inst_pe_1_7_6_net2873), .RN(npu_inst_pe_1_7_6_n10), .Q(
        npu_inst_pe_1_7_6_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_7_6_n107), 
        .CK(npu_inst_pe_1_7_6_net2873), .RN(npu_inst_pe_1_7_6_n10), .Q(
        npu_inst_pe_1_7_6_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_7_6_n106), 
        .CK(npu_inst_pe_1_7_6_net2873), .RN(npu_inst_pe_1_7_6_n10), .Q(
        npu_inst_pe_1_7_6_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_7_6_n105), 
        .CK(npu_inst_pe_1_7_6_net2873), .RN(npu_inst_pe_1_7_6_n10), .Q(
        npu_inst_pe_1_7_6_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_7_6_n104), 
        .CK(npu_inst_pe_1_7_6_net2873), .RN(npu_inst_pe_1_7_6_n10), .Q(
        npu_inst_pe_1_7_6_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_7_6_n103), 
        .CK(npu_inst_pe_1_7_6_net2873), .RN(npu_inst_pe_1_7_6_n10), .Q(
        npu_inst_pe_1_7_6_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_7_6_n102), 
        .CK(npu_inst_pe_1_7_6_net2873), .RN(npu_inst_pe_1_7_6_n10), .Q(
        npu_inst_pe_1_7_6_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_7_6_n86), 
        .CK(npu_inst_pe_1_7_6_net2873), .RN(npu_inst_pe_1_7_6_n10), .Q(
        npu_inst_pe_1_7_6_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_7_6_n87), 
        .CK(npu_inst_pe_1_7_6_net2873), .RN(npu_inst_pe_1_7_6_n10), .Q(
        npu_inst_pe_1_7_6_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_7_6_n88), 
        .CK(npu_inst_pe_1_7_6_net2873), .RN(npu_inst_pe_1_7_6_n11), .Q(
        npu_inst_pe_1_7_6_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_7_6_n89), 
        .CK(npu_inst_pe_1_7_6_net2873), .RN(npu_inst_pe_1_7_6_n11), .Q(
        npu_inst_pe_1_7_6_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_7_6_n90), 
        .CK(npu_inst_pe_1_7_6_net2873), .RN(npu_inst_pe_1_7_6_n11), .Q(
        npu_inst_pe_1_7_6_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_7_6_n91), 
        .CK(npu_inst_pe_1_7_6_net2873), .RN(npu_inst_pe_1_7_6_n11), .Q(
        npu_inst_pe_1_7_6_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_7_6_n92), 
        .CK(npu_inst_pe_1_7_6_net2873), .RN(npu_inst_pe_1_7_6_n11), .Q(
        npu_inst_pe_1_7_6_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_7_6_n93), 
        .CK(npu_inst_pe_1_7_6_net2873), .RN(npu_inst_pe_1_7_6_n11), .Q(
        npu_inst_pe_1_7_6_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_7_6_n94), 
        .CK(npu_inst_pe_1_7_6_net2873), .RN(npu_inst_pe_1_7_6_n11), .Q(
        npu_inst_pe_1_7_6_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_7_6_n95), 
        .CK(npu_inst_pe_1_7_6_net2873), .RN(npu_inst_pe_1_7_6_n11), .Q(
        npu_inst_pe_1_7_6_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_7_6_n96), 
        .CK(npu_inst_pe_1_7_6_net2873), .RN(npu_inst_pe_1_7_6_n11), .Q(
        npu_inst_pe_1_7_6_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_7_6_n97), 
        .CK(npu_inst_pe_1_7_6_net2873), .RN(npu_inst_pe_1_7_6_n11), .Q(
        npu_inst_pe_1_7_6_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_7_6_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_7_6_N84), .SE(1'b0), .GCK(npu_inst_pe_1_7_6_net2867) );
  CLKGATETST_X1 npu_inst_pe_1_7_6_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n61), .SE(1'b0), .GCK(npu_inst_pe_1_7_6_net2873) );
  MUX2_X1 npu_inst_pe_1_7_7_U162 ( .A(npu_inst_pe_1_7_7_n32), .B(
        npu_inst_pe_1_7_7_n29), .S(npu_inst_pe_1_7_7_n8), .Z(
        npu_inst_pe_1_7_7_N93) );
  MUX2_X1 npu_inst_pe_1_7_7_U161 ( .A(npu_inst_pe_1_7_7_n31), .B(
        npu_inst_pe_1_7_7_n30), .S(npu_inst_pe_1_7_7_n6), .Z(
        npu_inst_pe_1_7_7_n32) );
  MUX2_X1 npu_inst_pe_1_7_7_U160 ( .A(npu_inst_pe_1_7_7_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_7_7_int_q_reg_v_1__0_), .S(npu_inst_pe_1_7_7_n4), .Z(
        npu_inst_pe_1_7_7_n31) );
  MUX2_X1 npu_inst_pe_1_7_7_U159 ( .A(npu_inst_pe_1_7_7_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_7_7_int_q_reg_v_3__0_), .S(npu_inst_pe_1_7_7_n4), .Z(
        npu_inst_pe_1_7_7_n30) );
  MUX2_X1 npu_inst_pe_1_7_7_U158 ( .A(npu_inst_pe_1_7_7_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_7_7_int_q_reg_v_5__0_), .S(npu_inst_pe_1_7_7_n4), .Z(
        npu_inst_pe_1_7_7_n29) );
  MUX2_X1 npu_inst_pe_1_7_7_U157 ( .A(npu_inst_pe_1_7_7_n28), .B(
        npu_inst_pe_1_7_7_n23), .S(npu_inst_pe_1_7_7_n8), .Z(
        npu_inst_pe_1_7_7_N94) );
  MUX2_X1 npu_inst_pe_1_7_7_U156 ( .A(npu_inst_pe_1_7_7_n25), .B(
        npu_inst_pe_1_7_7_n24), .S(npu_inst_pe_1_7_7_n6), .Z(
        npu_inst_pe_1_7_7_n28) );
  MUX2_X1 npu_inst_pe_1_7_7_U155 ( .A(npu_inst_pe_1_7_7_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_7_7_int_q_reg_v_1__1_), .S(npu_inst_pe_1_7_7_n4), .Z(
        npu_inst_pe_1_7_7_n25) );
  MUX2_X1 npu_inst_pe_1_7_7_U154 ( .A(npu_inst_pe_1_7_7_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_7_7_int_q_reg_v_3__1_), .S(npu_inst_pe_1_7_7_n4), .Z(
        npu_inst_pe_1_7_7_n24) );
  MUX2_X1 npu_inst_pe_1_7_7_U153 ( .A(npu_inst_pe_1_7_7_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_7_7_int_q_reg_v_5__1_), .S(npu_inst_pe_1_7_7_n4), .Z(
        npu_inst_pe_1_7_7_n23) );
  MUX2_X1 npu_inst_pe_1_7_7_U152 ( .A(npu_inst_pe_1_7_7_n22), .B(
        npu_inst_pe_1_7_7_n19), .S(npu_inst_pe_1_7_7_n8), .Z(
        npu_inst_int_data_x_7__7__1_) );
  MUX2_X1 npu_inst_pe_1_7_7_U151 ( .A(npu_inst_pe_1_7_7_n21), .B(
        npu_inst_pe_1_7_7_n20), .S(npu_inst_pe_1_7_7_n6), .Z(
        npu_inst_pe_1_7_7_n22) );
  MUX2_X1 npu_inst_pe_1_7_7_U150 ( .A(npu_inst_pe_1_7_7_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_7_7_int_q_reg_h_1__1_), .S(npu_inst_pe_1_7_7_n4), .Z(
        npu_inst_pe_1_7_7_n21) );
  MUX2_X1 npu_inst_pe_1_7_7_U149 ( .A(npu_inst_pe_1_7_7_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_7_7_int_q_reg_h_3__1_), .S(npu_inst_pe_1_7_7_n4), .Z(
        npu_inst_pe_1_7_7_n20) );
  MUX2_X1 npu_inst_pe_1_7_7_U148 ( .A(npu_inst_pe_1_7_7_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_7_7_int_q_reg_h_5__1_), .S(npu_inst_pe_1_7_7_n4), .Z(
        npu_inst_pe_1_7_7_n19) );
  MUX2_X1 npu_inst_pe_1_7_7_U147 ( .A(npu_inst_pe_1_7_7_n18), .B(
        npu_inst_pe_1_7_7_n15), .S(npu_inst_pe_1_7_7_n8), .Z(
        npu_inst_int_data_x_7__7__0_) );
  MUX2_X1 npu_inst_pe_1_7_7_U146 ( .A(npu_inst_pe_1_7_7_n17), .B(
        npu_inst_pe_1_7_7_n16), .S(npu_inst_pe_1_7_7_n6), .Z(
        npu_inst_pe_1_7_7_n18) );
  MUX2_X1 npu_inst_pe_1_7_7_U145 ( .A(npu_inst_pe_1_7_7_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_7_7_int_q_reg_h_1__0_), .S(npu_inst_pe_1_7_7_n4), .Z(
        npu_inst_pe_1_7_7_n17) );
  MUX2_X1 npu_inst_pe_1_7_7_U144 ( .A(npu_inst_pe_1_7_7_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_7_7_int_q_reg_h_3__0_), .S(npu_inst_pe_1_7_7_n4), .Z(
        npu_inst_pe_1_7_7_n16) );
  MUX2_X1 npu_inst_pe_1_7_7_U143 ( .A(npu_inst_pe_1_7_7_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_7_7_int_q_reg_h_5__0_), .S(npu_inst_pe_1_7_7_n4), .Z(
        npu_inst_pe_1_7_7_n15) );
  XOR2_X1 npu_inst_pe_1_7_7_U142 ( .A(npu_inst_pe_1_7_7_int_data_0_), .B(
        npu_inst_pe_1_7_7_int_q_acc_0_), .Z(npu_inst_pe_1_7_7_N73) );
  AND2_X1 npu_inst_pe_1_7_7_U141 ( .A1(npu_inst_pe_1_7_7_int_q_acc_0_), .A2(
        npu_inst_pe_1_7_7_int_data_0_), .ZN(npu_inst_pe_1_7_7_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_7_7_U140 ( .A(npu_inst_pe_1_7_7_int_q_acc_0_), .B(
        npu_inst_pe_1_7_7_n13), .ZN(npu_inst_pe_1_7_7_N65) );
  OR2_X1 npu_inst_pe_1_7_7_U139 ( .A1(npu_inst_pe_1_7_7_n13), .A2(
        npu_inst_pe_1_7_7_int_q_acc_0_), .ZN(npu_inst_pe_1_7_7_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_7_7_U138 ( .A(npu_inst_pe_1_7_7_int_q_acc_2_), .B(
        npu_inst_pe_1_7_7_add_79_carry_2_), .Z(npu_inst_pe_1_7_7_N75) );
  AND2_X1 npu_inst_pe_1_7_7_U137 ( .A1(npu_inst_pe_1_7_7_add_79_carry_2_), 
        .A2(npu_inst_pe_1_7_7_int_q_acc_2_), .ZN(
        npu_inst_pe_1_7_7_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_7_7_U136 ( .A(npu_inst_pe_1_7_7_int_q_acc_3_), .B(
        npu_inst_pe_1_7_7_add_79_carry_3_), .Z(npu_inst_pe_1_7_7_N76) );
  AND2_X1 npu_inst_pe_1_7_7_U135 ( .A1(npu_inst_pe_1_7_7_add_79_carry_3_), 
        .A2(npu_inst_pe_1_7_7_int_q_acc_3_), .ZN(
        npu_inst_pe_1_7_7_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_7_7_U134 ( .A(npu_inst_pe_1_7_7_int_q_acc_4_), .B(
        npu_inst_pe_1_7_7_add_79_carry_4_), .Z(npu_inst_pe_1_7_7_N77) );
  AND2_X1 npu_inst_pe_1_7_7_U133 ( .A1(npu_inst_pe_1_7_7_add_79_carry_4_), 
        .A2(npu_inst_pe_1_7_7_int_q_acc_4_), .ZN(
        npu_inst_pe_1_7_7_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_7_7_U132 ( .A(npu_inst_pe_1_7_7_int_q_acc_5_), .B(
        npu_inst_pe_1_7_7_add_79_carry_5_), .Z(npu_inst_pe_1_7_7_N78) );
  AND2_X1 npu_inst_pe_1_7_7_U131 ( .A1(npu_inst_pe_1_7_7_add_79_carry_5_), 
        .A2(npu_inst_pe_1_7_7_int_q_acc_5_), .ZN(
        npu_inst_pe_1_7_7_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_7_7_U130 ( .A(npu_inst_pe_1_7_7_int_q_acc_6_), .B(
        npu_inst_pe_1_7_7_add_79_carry_6_), .Z(npu_inst_pe_1_7_7_N79) );
  AND2_X1 npu_inst_pe_1_7_7_U129 ( .A1(npu_inst_pe_1_7_7_add_79_carry_6_), 
        .A2(npu_inst_pe_1_7_7_int_q_acc_6_), .ZN(
        npu_inst_pe_1_7_7_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_7_7_U128 ( .A(npu_inst_pe_1_7_7_int_q_acc_7_), .B(
        npu_inst_pe_1_7_7_add_79_carry_7_), .Z(npu_inst_pe_1_7_7_N80) );
  XNOR2_X1 npu_inst_pe_1_7_7_U127 ( .A(npu_inst_pe_1_7_7_sub_77_carry_2_), .B(
        npu_inst_pe_1_7_7_int_q_acc_2_), .ZN(npu_inst_pe_1_7_7_N67) );
  OR2_X1 npu_inst_pe_1_7_7_U126 ( .A1(npu_inst_pe_1_7_7_int_q_acc_2_), .A2(
        npu_inst_pe_1_7_7_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_7_7_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_7_7_U125 ( .A(npu_inst_pe_1_7_7_sub_77_carry_3_), .B(
        npu_inst_pe_1_7_7_int_q_acc_3_), .ZN(npu_inst_pe_1_7_7_N68) );
  OR2_X1 npu_inst_pe_1_7_7_U124 ( .A1(npu_inst_pe_1_7_7_int_q_acc_3_), .A2(
        npu_inst_pe_1_7_7_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_7_7_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_7_7_U123 ( .A(npu_inst_pe_1_7_7_sub_77_carry_4_), .B(
        npu_inst_pe_1_7_7_int_q_acc_4_), .ZN(npu_inst_pe_1_7_7_N69) );
  OR2_X1 npu_inst_pe_1_7_7_U122 ( .A1(npu_inst_pe_1_7_7_int_q_acc_4_), .A2(
        npu_inst_pe_1_7_7_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_7_7_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_7_7_U121 ( .A(npu_inst_pe_1_7_7_sub_77_carry_5_), .B(
        npu_inst_pe_1_7_7_int_q_acc_5_), .ZN(npu_inst_pe_1_7_7_N70) );
  OR2_X1 npu_inst_pe_1_7_7_U120 ( .A1(npu_inst_pe_1_7_7_int_q_acc_5_), .A2(
        npu_inst_pe_1_7_7_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_7_7_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_7_7_U119 ( .A(npu_inst_pe_1_7_7_sub_77_carry_6_), .B(
        npu_inst_pe_1_7_7_int_q_acc_6_), .ZN(npu_inst_pe_1_7_7_N71) );
  OR2_X1 npu_inst_pe_1_7_7_U118 ( .A1(npu_inst_pe_1_7_7_int_q_acc_6_), .A2(
        npu_inst_pe_1_7_7_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_7_7_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_7_7_U117 ( .A(npu_inst_pe_1_7_7_int_q_acc_7_), .B(
        npu_inst_pe_1_7_7_sub_77_carry_7_), .ZN(npu_inst_pe_1_7_7_N72) );
  INV_X1 npu_inst_pe_1_7_7_U116 ( .A(npu_inst_n75), .ZN(npu_inst_pe_1_7_7_n7)
         );
  INV_X1 npu_inst_pe_1_7_7_U115 ( .A(npu_inst_pe_1_7_7_n7), .ZN(
        npu_inst_pe_1_7_7_n6) );
  INV_X1 npu_inst_pe_1_7_7_U114 ( .A(npu_inst_n52), .ZN(npu_inst_pe_1_7_7_n3)
         );
  AOI22_X1 npu_inst_pe_1_7_7_U113 ( .A1(npu_inst_pe_1_7_7_n38), .A2(
        int_i_data_v_npu[1]), .B1(npu_inst_pe_1_7_7_n118), .B2(
        npu_inst_pe_1_7_7_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_7_7_n39) );
  INV_X1 npu_inst_pe_1_7_7_U112 ( .A(npu_inst_pe_1_7_7_n39), .ZN(
        npu_inst_pe_1_7_7_n112) );
  AOI22_X1 npu_inst_pe_1_7_7_U111 ( .A1(npu_inst_pe_1_7_7_n38), .A2(
        int_i_data_v_npu[0]), .B1(npu_inst_pe_1_7_7_n118), .B2(
        npu_inst_pe_1_7_7_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_7_7_n37) );
  INV_X1 npu_inst_pe_1_7_7_U110 ( .A(npu_inst_pe_1_7_7_n37), .ZN(
        npu_inst_pe_1_7_7_n113) );
  AOI22_X1 npu_inst_pe_1_7_7_U107 ( .A1(int_i_data_v_npu[1]), .A2(
        npu_inst_pe_1_7_7_n58), .B1(npu_inst_pe_1_7_7_n114), .B2(
        npu_inst_pe_1_7_7_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_7_7_n59) );
  INV_X1 npu_inst_pe_1_7_7_U106 ( .A(npu_inst_pe_1_7_7_n59), .ZN(
        npu_inst_pe_1_7_7_n102) );
  AOI22_X1 npu_inst_pe_1_7_7_U105 ( .A1(int_i_data_v_npu[0]), .A2(
        npu_inst_pe_1_7_7_n58), .B1(npu_inst_pe_1_7_7_n114), .B2(
        npu_inst_pe_1_7_7_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_7_7_n57) );
  INV_X1 npu_inst_pe_1_7_7_U104 ( .A(npu_inst_pe_1_7_7_n57), .ZN(
        npu_inst_pe_1_7_7_n103) );
  AOI22_X1 npu_inst_pe_1_7_7_U103 ( .A1(int_i_data_v_npu[1]), .A2(
        npu_inst_pe_1_7_7_n54), .B1(npu_inst_pe_1_7_7_n115), .B2(
        npu_inst_pe_1_7_7_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_7_7_n55) );
  INV_X1 npu_inst_pe_1_7_7_U102 ( .A(npu_inst_pe_1_7_7_n55), .ZN(
        npu_inst_pe_1_7_7_n104) );
  AOI22_X1 npu_inst_pe_1_7_7_U101 ( .A1(int_i_data_v_npu[0]), .A2(
        npu_inst_pe_1_7_7_n54), .B1(npu_inst_pe_1_7_7_n115), .B2(
        npu_inst_pe_1_7_7_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_7_7_n53) );
  INV_X1 npu_inst_pe_1_7_7_U100 ( .A(npu_inst_pe_1_7_7_n53), .ZN(
        npu_inst_pe_1_7_7_n105) );
  AOI22_X1 npu_inst_pe_1_7_7_U99 ( .A1(int_i_data_v_npu[1]), .A2(
        npu_inst_pe_1_7_7_n50), .B1(npu_inst_pe_1_7_7_n116), .B2(
        npu_inst_pe_1_7_7_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_7_7_n51) );
  INV_X1 npu_inst_pe_1_7_7_U98 ( .A(npu_inst_pe_1_7_7_n51), .ZN(
        npu_inst_pe_1_7_7_n106) );
  AOI22_X1 npu_inst_pe_1_7_7_U97 ( .A1(int_i_data_v_npu[0]), .A2(
        npu_inst_pe_1_7_7_n50), .B1(npu_inst_pe_1_7_7_n116), .B2(
        npu_inst_pe_1_7_7_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_7_7_n49) );
  INV_X1 npu_inst_pe_1_7_7_U96 ( .A(npu_inst_pe_1_7_7_n49), .ZN(
        npu_inst_pe_1_7_7_n107) );
  AOI22_X1 npu_inst_pe_1_7_7_U95 ( .A1(int_i_data_v_npu[1]), .A2(
        npu_inst_pe_1_7_7_n46), .B1(npu_inst_pe_1_7_7_n117), .B2(
        npu_inst_pe_1_7_7_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_7_7_n47) );
  INV_X1 npu_inst_pe_1_7_7_U94 ( .A(npu_inst_pe_1_7_7_n47), .ZN(
        npu_inst_pe_1_7_7_n108) );
  AOI22_X1 npu_inst_pe_1_7_7_U93 ( .A1(int_i_data_v_npu[0]), .A2(
        npu_inst_pe_1_7_7_n46), .B1(npu_inst_pe_1_7_7_n117), .B2(
        npu_inst_pe_1_7_7_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_7_7_n45) );
  INV_X1 npu_inst_pe_1_7_7_U92 ( .A(npu_inst_pe_1_7_7_n45), .ZN(
        npu_inst_pe_1_7_7_n109) );
  AOI22_X1 npu_inst_pe_1_7_7_U91 ( .A1(int_i_data_v_npu[1]), .A2(
        npu_inst_pe_1_7_7_n42), .B1(npu_inst_pe_1_7_7_n119), .B2(
        npu_inst_pe_1_7_7_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_7_7_n43) );
  INV_X1 npu_inst_pe_1_7_7_U90 ( .A(npu_inst_pe_1_7_7_n43), .ZN(
        npu_inst_pe_1_7_7_n110) );
  AOI22_X1 npu_inst_pe_1_7_7_U89 ( .A1(int_i_data_v_npu[0]), .A2(
        npu_inst_pe_1_7_7_n42), .B1(npu_inst_pe_1_7_7_n119), .B2(
        npu_inst_pe_1_7_7_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_7_7_n41) );
  INV_X1 npu_inst_pe_1_7_7_U88 ( .A(npu_inst_pe_1_7_7_n41), .ZN(
        npu_inst_pe_1_7_7_n111) );
  AND2_X1 npu_inst_pe_1_7_7_U87 ( .A1(npu_inst_pe_1_7_7_N93), .A2(npu_inst_n52), .ZN(npu_inst_int_data_y_7__7__0_) );
  AND2_X1 npu_inst_pe_1_7_7_U86 ( .A1(npu_inst_n52), .A2(npu_inst_pe_1_7_7_N94), .ZN(npu_inst_int_data_y_7__7__1_) );
  NOR3_X1 npu_inst_pe_1_7_7_U85 ( .A1(npu_inst_pe_1_7_7_n26), .A2(npu_inst_n52), .A3(npu_inst_int_ckg[0]), .ZN(npu_inst_pe_1_7_7_n85) );
  OR2_X1 npu_inst_pe_1_7_7_U84 ( .A1(npu_inst_pe_1_7_7_n85), .A2(
        npu_inst_pe_1_7_7_n2), .ZN(npu_inst_pe_1_7_7_N84) );
  AOI222_X1 npu_inst_pe_1_7_7_U83 ( .A1(1'b0), .A2(npu_inst_pe_1_7_7_n1), .B1(
        npu_inst_pe_1_7_7_N73), .B2(npu_inst_pe_1_7_7_n76), .C1(
        npu_inst_pe_1_7_7_N65), .C2(npu_inst_pe_1_7_7_n77), .ZN(
        npu_inst_pe_1_7_7_n84) );
  INV_X1 npu_inst_pe_1_7_7_U82 ( .A(npu_inst_pe_1_7_7_n84), .ZN(
        npu_inst_pe_1_7_7_n101) );
  AOI222_X1 npu_inst_pe_1_7_7_U81 ( .A1(1'b0), .A2(npu_inst_pe_1_7_7_n1), .B1(
        npu_inst_pe_1_7_7_N80), .B2(npu_inst_pe_1_7_7_n76), .C1(
        npu_inst_pe_1_7_7_N72), .C2(npu_inst_pe_1_7_7_n77), .ZN(
        npu_inst_pe_1_7_7_n75) );
  INV_X1 npu_inst_pe_1_7_7_U80 ( .A(npu_inst_pe_1_7_7_n75), .ZN(
        npu_inst_pe_1_7_7_n33) );
  AOI222_X1 npu_inst_pe_1_7_7_U79 ( .A1(1'b0), .A2(npu_inst_pe_1_7_7_n1), .B1(
        npu_inst_pe_1_7_7_N74), .B2(npu_inst_pe_1_7_7_n76), .C1(
        npu_inst_pe_1_7_7_N66), .C2(npu_inst_pe_1_7_7_n77), .ZN(
        npu_inst_pe_1_7_7_n83) );
  INV_X1 npu_inst_pe_1_7_7_U78 ( .A(npu_inst_pe_1_7_7_n83), .ZN(
        npu_inst_pe_1_7_7_n100) );
  AOI222_X1 npu_inst_pe_1_7_7_U77 ( .A1(1'b0), .A2(npu_inst_pe_1_7_7_n1), .B1(
        npu_inst_pe_1_7_7_N75), .B2(npu_inst_pe_1_7_7_n76), .C1(
        npu_inst_pe_1_7_7_N67), .C2(npu_inst_pe_1_7_7_n77), .ZN(
        npu_inst_pe_1_7_7_n82) );
  INV_X1 npu_inst_pe_1_7_7_U76 ( .A(npu_inst_pe_1_7_7_n82), .ZN(
        npu_inst_pe_1_7_7_n99) );
  AOI222_X1 npu_inst_pe_1_7_7_U75 ( .A1(1'b0), .A2(npu_inst_pe_1_7_7_n1), .B1(
        npu_inst_pe_1_7_7_N76), .B2(npu_inst_pe_1_7_7_n76), .C1(
        npu_inst_pe_1_7_7_N68), .C2(npu_inst_pe_1_7_7_n77), .ZN(
        npu_inst_pe_1_7_7_n81) );
  INV_X1 npu_inst_pe_1_7_7_U74 ( .A(npu_inst_pe_1_7_7_n81), .ZN(
        npu_inst_pe_1_7_7_n98) );
  AOI222_X1 npu_inst_pe_1_7_7_U73 ( .A1(1'b0), .A2(npu_inst_pe_1_7_7_n1), .B1(
        npu_inst_pe_1_7_7_N77), .B2(npu_inst_pe_1_7_7_n76), .C1(
        npu_inst_pe_1_7_7_N69), .C2(npu_inst_pe_1_7_7_n77), .ZN(
        npu_inst_pe_1_7_7_n80) );
  INV_X1 npu_inst_pe_1_7_7_U72 ( .A(npu_inst_pe_1_7_7_n80), .ZN(
        npu_inst_pe_1_7_7_n36) );
  AOI222_X1 npu_inst_pe_1_7_7_U71 ( .A1(1'b0), .A2(npu_inst_pe_1_7_7_n1), .B1(
        npu_inst_pe_1_7_7_N78), .B2(npu_inst_pe_1_7_7_n76), .C1(
        npu_inst_pe_1_7_7_N70), .C2(npu_inst_pe_1_7_7_n77), .ZN(
        npu_inst_pe_1_7_7_n79) );
  INV_X1 npu_inst_pe_1_7_7_U70 ( .A(npu_inst_pe_1_7_7_n79), .ZN(
        npu_inst_pe_1_7_7_n35) );
  AOI222_X1 npu_inst_pe_1_7_7_U69 ( .A1(1'b0), .A2(npu_inst_pe_1_7_7_n1), .B1(
        npu_inst_pe_1_7_7_N79), .B2(npu_inst_pe_1_7_7_n76), .C1(
        npu_inst_pe_1_7_7_N71), .C2(npu_inst_pe_1_7_7_n77), .ZN(
        npu_inst_pe_1_7_7_n78) );
  INV_X1 npu_inst_pe_1_7_7_U68 ( .A(npu_inst_pe_1_7_7_n78), .ZN(
        npu_inst_pe_1_7_7_n34) );
  AND2_X1 npu_inst_pe_1_7_7_U67 ( .A1(npu_inst_pe_1_7_7_int_q_acc_0_), .A2(
        npu_inst_pe_1_7_7_n1), .ZN(npu_inst_int_data_res_7__7__0_) );
  AND2_X1 npu_inst_pe_1_7_7_U66 ( .A1(npu_inst_pe_1_7_7_n2), .A2(
        npu_inst_pe_1_7_7_int_q_acc_7_), .ZN(npu_inst_int_data_res_7__7__7_)
         );
  AND2_X1 npu_inst_pe_1_7_7_U65 ( .A1(npu_inst_pe_1_7_7_int_q_acc_1_), .A2(
        npu_inst_pe_1_7_7_n1), .ZN(npu_inst_int_data_res_7__7__1_) );
  AND2_X1 npu_inst_pe_1_7_7_U64 ( .A1(npu_inst_pe_1_7_7_int_q_acc_2_), .A2(
        npu_inst_pe_1_7_7_n1), .ZN(npu_inst_int_data_res_7__7__2_) );
  AND2_X1 npu_inst_pe_1_7_7_U63 ( .A1(npu_inst_pe_1_7_7_int_q_acc_3_), .A2(
        npu_inst_pe_1_7_7_n2), .ZN(npu_inst_int_data_res_7__7__3_) );
  AND2_X1 npu_inst_pe_1_7_7_U62 ( .A1(npu_inst_pe_1_7_7_int_q_acc_4_), .A2(
        npu_inst_pe_1_7_7_n2), .ZN(npu_inst_int_data_res_7__7__4_) );
  AND2_X1 npu_inst_pe_1_7_7_U61 ( .A1(npu_inst_pe_1_7_7_int_q_acc_5_), .A2(
        npu_inst_pe_1_7_7_n2), .ZN(npu_inst_int_data_res_7__7__5_) );
  AND2_X1 npu_inst_pe_1_7_7_U60 ( .A1(npu_inst_pe_1_7_7_int_q_acc_6_), .A2(
        npu_inst_pe_1_7_7_n2), .ZN(npu_inst_int_data_res_7__7__6_) );
  INV_X1 npu_inst_pe_1_7_7_U59 ( .A(npu_inst_pe_1_7_7_int_data_1_), .ZN(
        npu_inst_pe_1_7_7_n14) );
  AND2_X1 npu_inst_pe_1_7_7_U58 ( .A1(npu_inst_int_data_x_7__7__1_), .A2(
        npu_inst_pe_1_7_7_int_q_weight_1_), .ZN(npu_inst_pe_1_7_7_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_7_7_U57 ( .A1(npu_inst_int_data_x_7__7__0_), .A2(
        npu_inst_pe_1_7_7_int_q_weight_1_), .ZN(npu_inst_pe_1_7_7_int_data_0_)
         );
  NAND2_X1 npu_inst_pe_1_7_7_U56 ( .A1(npu_inst_pe_1_7_7_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_7_7_n60), .ZN(npu_inst_pe_1_7_7_n74) );
  OAI21_X1 npu_inst_pe_1_7_7_U55 ( .B1(npu_inst_pe_1_7_7_n63), .B2(
        npu_inst_pe_1_7_7_n60), .A(npu_inst_pe_1_7_7_n74), .ZN(
        npu_inst_pe_1_7_7_n97) );
  NAND2_X1 npu_inst_pe_1_7_7_U54 ( .A1(npu_inst_pe_1_7_7_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_7_7_n60), .ZN(npu_inst_pe_1_7_7_n73) );
  OAI21_X1 npu_inst_pe_1_7_7_U53 ( .B1(npu_inst_pe_1_7_7_n61), .B2(
        npu_inst_pe_1_7_7_n60), .A(npu_inst_pe_1_7_7_n73), .ZN(
        npu_inst_pe_1_7_7_n96) );
  NAND2_X1 npu_inst_pe_1_7_7_U52 ( .A1(npu_inst_pe_1_7_7_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_7_7_n56), .ZN(npu_inst_pe_1_7_7_n72) );
  OAI21_X1 npu_inst_pe_1_7_7_U51 ( .B1(npu_inst_pe_1_7_7_n63), .B2(
        npu_inst_pe_1_7_7_n56), .A(npu_inst_pe_1_7_7_n72), .ZN(
        npu_inst_pe_1_7_7_n95) );
  NAND2_X1 npu_inst_pe_1_7_7_U50 ( .A1(npu_inst_pe_1_7_7_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_7_7_n56), .ZN(npu_inst_pe_1_7_7_n71) );
  OAI21_X1 npu_inst_pe_1_7_7_U49 ( .B1(npu_inst_pe_1_7_7_n61), .B2(
        npu_inst_pe_1_7_7_n56), .A(npu_inst_pe_1_7_7_n71), .ZN(
        npu_inst_pe_1_7_7_n94) );
  NAND2_X1 npu_inst_pe_1_7_7_U48 ( .A1(npu_inst_pe_1_7_7_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_7_7_n52), .ZN(npu_inst_pe_1_7_7_n70) );
  OAI21_X1 npu_inst_pe_1_7_7_U47 ( .B1(npu_inst_pe_1_7_7_n63), .B2(
        npu_inst_pe_1_7_7_n52), .A(npu_inst_pe_1_7_7_n70), .ZN(
        npu_inst_pe_1_7_7_n93) );
  NAND2_X1 npu_inst_pe_1_7_7_U46 ( .A1(npu_inst_pe_1_7_7_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_7_7_n52), .ZN(npu_inst_pe_1_7_7_n69) );
  OAI21_X1 npu_inst_pe_1_7_7_U45 ( .B1(npu_inst_pe_1_7_7_n61), .B2(
        npu_inst_pe_1_7_7_n52), .A(npu_inst_pe_1_7_7_n69), .ZN(
        npu_inst_pe_1_7_7_n92) );
  NAND2_X1 npu_inst_pe_1_7_7_U44 ( .A1(npu_inst_pe_1_7_7_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_7_7_n48), .ZN(npu_inst_pe_1_7_7_n68) );
  OAI21_X1 npu_inst_pe_1_7_7_U43 ( .B1(npu_inst_pe_1_7_7_n63), .B2(
        npu_inst_pe_1_7_7_n48), .A(npu_inst_pe_1_7_7_n68), .ZN(
        npu_inst_pe_1_7_7_n91) );
  NAND2_X1 npu_inst_pe_1_7_7_U42 ( .A1(npu_inst_pe_1_7_7_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_7_7_n48), .ZN(npu_inst_pe_1_7_7_n67) );
  OAI21_X1 npu_inst_pe_1_7_7_U41 ( .B1(npu_inst_pe_1_7_7_n61), .B2(
        npu_inst_pe_1_7_7_n48), .A(npu_inst_pe_1_7_7_n67), .ZN(
        npu_inst_pe_1_7_7_n90) );
  NAND2_X1 npu_inst_pe_1_7_7_U40 ( .A1(npu_inst_pe_1_7_7_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_7_7_n44), .ZN(npu_inst_pe_1_7_7_n66) );
  OAI21_X1 npu_inst_pe_1_7_7_U39 ( .B1(npu_inst_pe_1_7_7_n63), .B2(
        npu_inst_pe_1_7_7_n44), .A(npu_inst_pe_1_7_7_n66), .ZN(
        npu_inst_pe_1_7_7_n89) );
  NAND2_X1 npu_inst_pe_1_7_7_U38 ( .A1(npu_inst_pe_1_7_7_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_7_7_n44), .ZN(npu_inst_pe_1_7_7_n65) );
  OAI21_X1 npu_inst_pe_1_7_7_U37 ( .B1(npu_inst_pe_1_7_7_n61), .B2(
        npu_inst_pe_1_7_7_n44), .A(npu_inst_pe_1_7_7_n65), .ZN(
        npu_inst_pe_1_7_7_n88) );
  NAND2_X1 npu_inst_pe_1_7_7_U36 ( .A1(npu_inst_pe_1_7_7_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_7_7_n40), .ZN(npu_inst_pe_1_7_7_n64) );
  OAI21_X1 npu_inst_pe_1_7_7_U35 ( .B1(npu_inst_pe_1_7_7_n63), .B2(
        npu_inst_pe_1_7_7_n40), .A(npu_inst_pe_1_7_7_n64), .ZN(
        npu_inst_pe_1_7_7_n87) );
  NAND2_X1 npu_inst_pe_1_7_7_U34 ( .A1(npu_inst_pe_1_7_7_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_7_7_n40), .ZN(npu_inst_pe_1_7_7_n62) );
  OAI21_X1 npu_inst_pe_1_7_7_U33 ( .B1(npu_inst_pe_1_7_7_n61), .B2(
        npu_inst_pe_1_7_7_n40), .A(npu_inst_pe_1_7_7_n62), .ZN(
        npu_inst_pe_1_7_7_n86) );
  AOI22_X1 npu_inst_pe_1_7_7_U32 ( .A1(npu_inst_n52), .A2(int_i_data_v_npu[1]), 
        .B1(npu_inst_pe_1_7_7_n3), .B2(int_i_data_h_npu8[1]), .ZN(
        npu_inst_pe_1_7_7_n63) );
  AOI22_X1 npu_inst_pe_1_7_7_U31 ( .A1(npu_inst_n52), .A2(int_i_data_v_npu[0]), 
        .B1(npu_inst_pe_1_7_7_n3), .B2(int_i_data_h_npu8[0]), .ZN(
        npu_inst_pe_1_7_7_n61) );
  INV_X1 npu_inst_pe_1_7_7_U30 ( .A(npu_inst_pe_1_7_7_int_data_0_), .ZN(
        npu_inst_pe_1_7_7_n13) );
  INV_X1 npu_inst_pe_1_7_7_U29 ( .A(npu_inst_n67), .ZN(npu_inst_pe_1_7_7_n5)
         );
  OR3_X1 npu_inst_pe_1_7_7_U28 ( .A1(npu_inst_pe_1_7_7_n6), .A2(
        npu_inst_pe_1_7_7_n8), .A3(npu_inst_pe_1_7_7_n5), .ZN(
        npu_inst_pe_1_7_7_n56) );
  OR3_X1 npu_inst_pe_1_7_7_U27 ( .A1(npu_inst_pe_1_7_7_n5), .A2(
        npu_inst_pe_1_7_7_n8), .A3(npu_inst_pe_1_7_7_n7), .ZN(
        npu_inst_pe_1_7_7_n48) );
  INV_X1 npu_inst_pe_1_7_7_U26 ( .A(npu_inst_pe_1_7_7_n5), .ZN(
        npu_inst_pe_1_7_7_n4) );
  INV_X1 npu_inst_pe_1_7_7_U25 ( .A(npu_inst_n122), .ZN(npu_inst_pe_1_7_7_n12)
         );
  OR3_X1 npu_inst_pe_1_7_7_U24 ( .A1(npu_inst_pe_1_7_7_n4), .A2(
        npu_inst_pe_1_7_7_n8), .A3(npu_inst_pe_1_7_7_n7), .ZN(
        npu_inst_pe_1_7_7_n52) );
  OR3_X1 npu_inst_pe_1_7_7_U23 ( .A1(npu_inst_pe_1_7_7_n6), .A2(
        npu_inst_pe_1_7_7_n8), .A3(npu_inst_pe_1_7_7_n4), .ZN(
        npu_inst_pe_1_7_7_n60) );
  NOR2_X1 npu_inst_pe_1_7_7_U22 ( .A1(npu_inst_pe_1_7_7_n60), .A2(
        npu_inst_pe_1_7_7_n3), .ZN(npu_inst_pe_1_7_7_n58) );
  NOR2_X1 npu_inst_pe_1_7_7_U21 ( .A1(npu_inst_pe_1_7_7_n56), .A2(
        npu_inst_pe_1_7_7_n3), .ZN(npu_inst_pe_1_7_7_n54) );
  NOR2_X1 npu_inst_pe_1_7_7_U20 ( .A1(npu_inst_pe_1_7_7_n52), .A2(
        npu_inst_pe_1_7_7_n3), .ZN(npu_inst_pe_1_7_7_n50) );
  NOR2_X1 npu_inst_pe_1_7_7_U19 ( .A1(npu_inst_pe_1_7_7_n48), .A2(
        npu_inst_pe_1_7_7_n3), .ZN(npu_inst_pe_1_7_7_n46) );
  NOR2_X1 npu_inst_pe_1_7_7_U18 ( .A1(npu_inst_pe_1_7_7_n40), .A2(
        npu_inst_pe_1_7_7_n3), .ZN(npu_inst_pe_1_7_7_n38) );
  NOR2_X1 npu_inst_pe_1_7_7_U17 ( .A1(npu_inst_pe_1_7_7_n44), .A2(
        npu_inst_pe_1_7_7_n3), .ZN(npu_inst_pe_1_7_7_n42) );
  BUF_X1 npu_inst_pe_1_7_7_U16 ( .A(npu_inst_n92), .Z(npu_inst_pe_1_7_7_n8) );
  BUF_X1 npu_inst_pe_1_7_7_U15 ( .A(npu_inst_pe_1_7_7_n12), .Z(
        npu_inst_pe_1_7_7_n11) );
  BUF_X1 npu_inst_pe_1_7_7_U14 ( .A(npu_inst_pe_1_7_7_n12), .Z(
        npu_inst_pe_1_7_7_n10) );
  BUF_X1 npu_inst_pe_1_7_7_U13 ( .A(npu_inst_pe_1_7_7_n12), .Z(
        npu_inst_pe_1_7_7_n9) );
  INV_X1 npu_inst_pe_1_7_7_U12 ( .A(npu_inst_pe_1_7_7_n38), .ZN(
        npu_inst_pe_1_7_7_n118) );
  INV_X1 npu_inst_pe_1_7_7_U11 ( .A(npu_inst_pe_1_7_7_n58), .ZN(
        npu_inst_pe_1_7_7_n114) );
  INV_X1 npu_inst_pe_1_7_7_U10 ( .A(npu_inst_pe_1_7_7_n54), .ZN(
        npu_inst_pe_1_7_7_n115) );
  INV_X1 npu_inst_pe_1_7_7_U9 ( .A(npu_inst_pe_1_7_7_n50), .ZN(
        npu_inst_pe_1_7_7_n116) );
  INV_X1 npu_inst_pe_1_7_7_U8 ( .A(npu_inst_pe_1_7_7_n46), .ZN(
        npu_inst_pe_1_7_7_n117) );
  INV_X1 npu_inst_pe_1_7_7_U7 ( .A(npu_inst_pe_1_7_7_n42), .ZN(
        npu_inst_pe_1_7_7_n119) );
  BUF_X1 npu_inst_pe_1_7_7_U6 ( .A(npu_inst_n7), .Z(npu_inst_pe_1_7_7_n2) );
  BUF_X1 npu_inst_pe_1_7_7_U5 ( .A(npu_inst_n7), .Z(npu_inst_pe_1_7_7_n1) );
  NOR2_X1 npu_inst_pe_1_7_7_U4 ( .A1(npu_inst_pe_1_7_7_int_q_weight_0_), .A2(
        npu_inst_pe_1_7_7_n1), .ZN(npu_inst_pe_1_7_7_n76) );
  NOR2_X1 npu_inst_pe_1_7_7_U3 ( .A1(npu_inst_pe_1_7_7_n27), .A2(
        npu_inst_pe_1_7_7_n1), .ZN(npu_inst_pe_1_7_7_n77) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_7_7_n111), 
        .CK(npu_inst_pe_1_7_7_net2850), .RN(npu_inst_pe_1_7_7_n12), .Q(
        npu_inst_pe_1_7_7_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_7_7_n110), 
        .CK(npu_inst_pe_1_7_7_net2850), .RN(npu_inst_pe_1_7_7_n12), .Q(
        npu_inst_pe_1_7_7_int_q_reg_v_4__1_) );
  FA_X1 npu_inst_pe_1_7_7_sub_77_U2_1 ( .A(npu_inst_pe_1_7_7_int_q_acc_1_), 
        .B(npu_inst_pe_1_7_7_n14), .CI(npu_inst_pe_1_7_7_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_7_7_sub_77_carry_2_), .S(npu_inst_pe_1_7_7_N66) );
  FA_X1 npu_inst_pe_1_7_7_add_79_U1_1 ( .A(npu_inst_pe_1_7_7_int_q_acc_1_), 
        .B(npu_inst_pe_1_7_7_int_data_1_), .CI(
        npu_inst_pe_1_7_7_add_79_carry_1_), .CO(
        npu_inst_pe_1_7_7_add_79_carry_2_), .S(npu_inst_pe_1_7_7_N74) );
  NAND3_X1 npu_inst_pe_1_7_7_U109 ( .A1(npu_inst_pe_1_7_7_n5), .A2(
        npu_inst_pe_1_7_7_n7), .A3(npu_inst_pe_1_7_7_n8), .ZN(
        npu_inst_pe_1_7_7_n44) );
  NAND3_X1 npu_inst_pe_1_7_7_U108 ( .A1(npu_inst_pe_1_7_7_n4), .A2(
        npu_inst_pe_1_7_7_n7), .A3(npu_inst_pe_1_7_7_n8), .ZN(
        npu_inst_pe_1_7_7_n40) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_7_7_n34), .CK(
        npu_inst_pe_1_7_7_net2844), .RN(npu_inst_pe_1_7_7_n9), .Q(
        npu_inst_pe_1_7_7_int_q_acc_6_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_7_7_n35), .CK(
        npu_inst_pe_1_7_7_net2844), .RN(npu_inst_pe_1_7_7_n9), .Q(
        npu_inst_pe_1_7_7_int_q_acc_5_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_7_7_n36), .CK(
        npu_inst_pe_1_7_7_net2844), .RN(npu_inst_pe_1_7_7_n9), .Q(
        npu_inst_pe_1_7_7_int_q_acc_4_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_7_7_n98), .CK(
        npu_inst_pe_1_7_7_net2844), .RN(npu_inst_pe_1_7_7_n9), .Q(
        npu_inst_pe_1_7_7_int_q_acc_3_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_7_7_n99), .CK(
        npu_inst_pe_1_7_7_net2844), .RN(npu_inst_pe_1_7_7_n9), .Q(
        npu_inst_pe_1_7_7_int_q_acc_2_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_7_7_n100), 
        .CK(npu_inst_pe_1_7_7_net2844), .RN(npu_inst_pe_1_7_7_n9), .Q(
        npu_inst_pe_1_7_7_int_q_acc_1_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_7_7_n33), .CK(
        npu_inst_pe_1_7_7_net2844), .RN(npu_inst_pe_1_7_7_n9), .Q(
        npu_inst_pe_1_7_7_int_q_acc_7_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_7_7_n101), 
        .CK(npu_inst_pe_1_7_7_net2844), .RN(npu_inst_pe_1_7_7_n9), .Q(
        npu_inst_pe_1_7_7_int_q_acc_0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_weight_reg_0_ ( .D(npu_inst_n108), .CK(
        npu_inst_pe_1_7_7_net2850), .RN(npu_inst_pe_1_7_7_n9), .Q(
        npu_inst_pe_1_7_7_int_q_weight_0_), .QN(npu_inst_pe_1_7_7_n27) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_weight_reg_1_ ( .D(npu_inst_n114), .CK(
        npu_inst_pe_1_7_7_net2850), .RN(npu_inst_pe_1_7_7_n9), .Q(
        npu_inst_pe_1_7_7_int_q_weight_1_), .QN(npu_inst_pe_1_7_7_n26) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_7_7_n113), 
        .CK(npu_inst_pe_1_7_7_net2850), .RN(npu_inst_pe_1_7_7_n9), .Q(
        npu_inst_pe_1_7_7_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_7_7_n112), 
        .CK(npu_inst_pe_1_7_7_net2850), .RN(npu_inst_pe_1_7_7_n9), .Q(
        npu_inst_pe_1_7_7_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_7_7_n109), 
        .CK(npu_inst_pe_1_7_7_net2850), .RN(npu_inst_pe_1_7_7_n10), .Q(
        npu_inst_pe_1_7_7_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_7_7_n108), 
        .CK(npu_inst_pe_1_7_7_net2850), .RN(npu_inst_pe_1_7_7_n10), .Q(
        npu_inst_pe_1_7_7_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_7_7_n107), 
        .CK(npu_inst_pe_1_7_7_net2850), .RN(npu_inst_pe_1_7_7_n10), .Q(
        npu_inst_pe_1_7_7_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_7_7_n106), 
        .CK(npu_inst_pe_1_7_7_net2850), .RN(npu_inst_pe_1_7_7_n10), .Q(
        npu_inst_pe_1_7_7_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_7_7_n105), 
        .CK(npu_inst_pe_1_7_7_net2850), .RN(npu_inst_pe_1_7_7_n10), .Q(
        npu_inst_pe_1_7_7_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_7_7_n104), 
        .CK(npu_inst_pe_1_7_7_net2850), .RN(npu_inst_pe_1_7_7_n10), .Q(
        npu_inst_pe_1_7_7_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_7_7_n103), 
        .CK(npu_inst_pe_1_7_7_net2850), .RN(npu_inst_pe_1_7_7_n10), .Q(
        npu_inst_pe_1_7_7_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_7_7_n102), 
        .CK(npu_inst_pe_1_7_7_net2850), .RN(npu_inst_pe_1_7_7_n10), .Q(
        npu_inst_pe_1_7_7_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_7_7_n86), 
        .CK(npu_inst_pe_1_7_7_net2850), .RN(npu_inst_pe_1_7_7_n10), .Q(
        npu_inst_pe_1_7_7_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_7_7_n87), 
        .CK(npu_inst_pe_1_7_7_net2850), .RN(npu_inst_pe_1_7_7_n10), .Q(
        npu_inst_pe_1_7_7_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_7_7_n88), 
        .CK(npu_inst_pe_1_7_7_net2850), .RN(npu_inst_pe_1_7_7_n11), .Q(
        npu_inst_pe_1_7_7_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_7_7_n89), 
        .CK(npu_inst_pe_1_7_7_net2850), .RN(npu_inst_pe_1_7_7_n11), .Q(
        npu_inst_pe_1_7_7_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_7_7_n90), 
        .CK(npu_inst_pe_1_7_7_net2850), .RN(npu_inst_pe_1_7_7_n11), .Q(
        npu_inst_pe_1_7_7_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_7_7_n91), 
        .CK(npu_inst_pe_1_7_7_net2850), .RN(npu_inst_pe_1_7_7_n11), .Q(
        npu_inst_pe_1_7_7_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_7_7_n92), 
        .CK(npu_inst_pe_1_7_7_net2850), .RN(npu_inst_pe_1_7_7_n11), .Q(
        npu_inst_pe_1_7_7_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_7_7_n93), 
        .CK(npu_inst_pe_1_7_7_net2850), .RN(npu_inst_pe_1_7_7_n11), .Q(
        npu_inst_pe_1_7_7_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_7_7_n94), 
        .CK(npu_inst_pe_1_7_7_net2850), .RN(npu_inst_pe_1_7_7_n11), .Q(
        npu_inst_pe_1_7_7_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_7_7_n95), 
        .CK(npu_inst_pe_1_7_7_net2850), .RN(npu_inst_pe_1_7_7_n11), .Q(
        npu_inst_pe_1_7_7_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_7_7_n96), 
        .CK(npu_inst_pe_1_7_7_net2850), .RN(npu_inst_pe_1_7_7_n11), .Q(
        npu_inst_pe_1_7_7_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_7_7_n97), 
        .CK(npu_inst_pe_1_7_7_net2850), .RN(npu_inst_pe_1_7_7_n11), .Q(
        npu_inst_pe_1_7_7_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_7_7_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_7_7_N84), .SE(1'b0), .GCK(npu_inst_pe_1_7_7_net2844) );
  CLKGATETST_X1 npu_inst_pe_1_7_7_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n61), .SE(1'b0), .GCK(npu_inst_pe_1_7_7_net2850) );
  INV_X1 ckg_ctrl8b_inst_U34 ( .A(ps_int_s_tc_tileh), .ZN(ckg_ctrl8b_inst_n10)
         );
  NOR2_X1 ckg_ctrl8b_inst_U33 ( .A1(arv_ckg[2]), .A2(ckg_ctrl8b_inst_n11), 
        .ZN(int_ckg_rmask[4]) );
  NOR2_X1 ckg_ctrl8b_inst_U32 ( .A1(arv_ckg[2]), .A2(ckg_ctrl8b_inst_n10), 
        .ZN(int_ckg_cmask[4]) );
  NAND2_X1 ckg_ctrl8b_inst_U31 ( .A1(ps_int_s_tc_tileh), .A2(
        ckg_ctrl8b_inst_n14), .ZN(ckg_ctrl8b_inst_n19) );
  INV_X1 ckg_ctrl8b_inst_U30 ( .A(arv_ckg[1]), .ZN(ckg_ctrl8b_inst_n8) );
  NAND2_X1 ckg_ctrl8b_inst_U29 ( .A1(ps_int_s_tc_tilev), .A2(
        ckg_ctrl8b_inst_n14), .ZN(ckg_ctrl8b_inst_n13) );
  INV_X1 ckg_ctrl8b_inst_U28 ( .A(arv_ckg[0]), .ZN(ckg_ctrl8b_inst_n9) );
  INV_X1 ckg_ctrl8b_inst_U27 ( .A(arv_ckg[2]), .ZN(ckg_ctrl8b_inst_n5) );
  OAI21_X1 ckg_ctrl8b_inst_U26 ( .B1(arv_ckg[1]), .B2(arv_ckg[0]), .A(
        arv_ckg[2]), .ZN(ckg_ctrl8b_inst_n14) );
  INV_X1 ckg_ctrl8b_inst_U25 ( .A(arv_npu[0]), .ZN(ckg_ctrl8b_inst_n3) );
  OAI22_X1 ckg_ctrl8b_inst_U24 ( .A1(ps_int_s_tc_tilev), .A2(
        ckg_ctrl8b_inst_n3), .B1(ckg_ctrl8b_inst_n9), .B2(ckg_ctrl8b_inst_n11), 
        .ZN(int_arv_res[0]) );
  INV_X1 ckg_ctrl8b_inst_U23 ( .A(arv_npu[1]), .ZN(ckg_ctrl8b_inst_n2) );
  OAI22_X1 ckg_ctrl8b_inst_U22 ( .A1(ps_int_s_tc_tilev), .A2(
        ckg_ctrl8b_inst_n2), .B1(ckg_ctrl8b_inst_n8), .B2(ckg_ctrl8b_inst_n11), 
        .ZN(int_arv_res[1]) );
  INV_X1 ckg_ctrl8b_inst_U21 ( .A(arv_npu[2]), .ZN(ckg_ctrl8b_inst_n1) );
  OAI22_X1 ckg_ctrl8b_inst_U20 ( .A1(ps_int_s_tc_tilev), .A2(
        ckg_ctrl8b_inst_n1), .B1(ckg_ctrl8b_inst_n5), .B2(ckg_ctrl8b_inst_n11), 
        .ZN(int_arv_res[2]) );
  OAI21_X1 ckg_ctrl8b_inst_U19 ( .B1(arv_ckg[1]), .B2(ckg_ctrl8b_inst_n11), 
        .A(ckg_ctrl8b_inst_n13), .ZN(int_ckg_rmask[6]) );
  OAI21_X1 ckg_ctrl8b_inst_U18 ( .B1(arv_ckg[1]), .B2(ckg_ctrl8b_inst_n10), 
        .A(ckg_ctrl8b_inst_n19), .ZN(int_ckg_cmask[6]) );
  INV_X1 ckg_ctrl8b_inst_U17 ( .A(ps_int_s_tc_tilev), .ZN(ckg_ctrl8b_inst_n11)
         );
  NAND2_X1 ckg_ctrl8b_inst_U16 ( .A1(ckg_ctrl8b_inst_n8), .A2(
        ckg_ctrl8b_inst_n5), .ZN(ckg_ctrl8b_inst_n16) );
  INV_X1 ckg_ctrl8b_inst_U15 ( .A(ckg_ctrl8b_inst_n16), .ZN(ckg_ctrl8b_inst_n4) );
  AOI21_X1 ckg_ctrl8b_inst_U14 ( .B1(ckg_ctrl8b_inst_n5), .B2(
        ckg_ctrl8b_inst_n9), .A(ckg_ctrl8b_inst_n4), .ZN(ckg_ctrl8b_inst_n15)
         );
  NOR3_X1 ckg_ctrl8b_inst_U13 ( .A1(ckg_ctrl8b_inst_n17), .A2(
        ckg_ctrl8b_inst_n11), .A3(ckg_ctrl8b_inst_n18), .ZN(int_ckg_rmask[1])
         );
  NOR2_X1 ckg_ctrl8b_inst_U12 ( .A1(ckg_ctrl8b_inst_n11), .A2(
        ckg_ctrl8b_inst_n16), .ZN(int_ckg_rmask[2]) );
  NOR2_X1 ckg_ctrl8b_inst_U11 ( .A1(ckg_ctrl8b_inst_n15), .A2(
        ckg_ctrl8b_inst_n11), .ZN(int_ckg_rmask[3]) );
  NOR2_X1 ckg_ctrl8b_inst_U10 ( .A1(ckg_ctrl8b_inst_n12), .A2(
        ckg_ctrl8b_inst_n11), .ZN(int_ckg_rmask[7]) );
  INV_X1 ckg_ctrl8b_inst_U9 ( .A(ckg_ctrl8b_inst_n13), .ZN(int_ckg_rmask[5])
         );
  NOR3_X1 ckg_ctrl8b_inst_U8 ( .A1(ckg_ctrl8b_inst_n10), .A2(
        ckg_ctrl8b_inst_n17), .A3(ckg_ctrl8b_inst_n18), .ZN(int_ckg_cmask[1])
         );
  NOR2_X1 ckg_ctrl8b_inst_U7 ( .A1(ckg_ctrl8b_inst_n16), .A2(
        ckg_ctrl8b_inst_n10), .ZN(int_ckg_cmask[2]) );
  NOR2_X1 ckg_ctrl8b_inst_U6 ( .A1(ckg_ctrl8b_inst_n15), .A2(
        ckg_ctrl8b_inst_n10), .ZN(int_ckg_cmask[3]) );
  NOR2_X1 ckg_ctrl8b_inst_U5 ( .A1(ckg_ctrl8b_inst_n12), .A2(
        ckg_ctrl8b_inst_n10), .ZN(int_ckg_cmask[7]) );
  INV_X1 ckg_ctrl8b_inst_U4 ( .A(ckg_ctrl8b_inst_n19), .ZN(int_ckg_cmask[5])
         );
  OAI22_X1 ckg_ctrl8b_inst_U3 ( .A1(ckg_ctrl8b_inst_n8), .A2(
        ckg_ctrl8b_inst_n9), .B1(ckg_ctrl8b_inst_n5), .B2(ckg_ctrl8b_inst_n20), 
        .ZN(ckg_ctrl8b_inst_n17) );
  AND2_X1 ckg_ctrl8b_inst_U2 ( .A1(ckg_ctrl8b_inst_n18), .A2(
        ckg_ctrl8b_inst_n17), .ZN(ckg_ctrl8b_inst_n12) );
  XOR2_X1 ckg_ctrl8b_inst_U36 ( .A(ckg_ctrl8b_inst_n9), .B(arv_ckg[1]), .Z(
        ckg_ctrl8b_inst_n20) );
  XOR2_X1 ckg_ctrl8b_inst_U35 ( .A(ckg_ctrl8b_inst_n5), .B(ckg_ctrl8b_inst_n20), .Z(ckg_ctrl8b_inst_n18) );
  INV_X1 hmode_cnt_inst_U14 ( .A(n10), .ZN(hmode_cnt_inst_n12) );
  AOI21_X1 hmode_cnt_inst_U13 ( .B1(hmode_cnt_inst_n10), .B2(hmode_cnt_inst_n7), .A(hmode_cnt_inst_N10), .ZN(hmode_cnt_inst_n8) );
  NAND4_X1 hmode_cnt_inst_U12 ( .A1(hmode_cnt_inst_n10), .A2(int_hmode_cnt[1]), 
        .A3(int_hmode_cnt[0]), .A4(hmode_cnt_inst_n5), .ZN(hmode_cnt_inst_n9)
         );
  OAI21_X1 hmode_cnt_inst_U11 ( .B1(hmode_cnt_inst_n8), .B2(hmode_cnt_inst_n5), 
        .A(hmode_cnt_inst_n9), .ZN(hmode_cnt_inst_N12) );
  XNOR2_X1 hmode_cnt_inst_U10 ( .A(int_hmode_cnt[0]), .B(int_hmode_cnt[1]), 
        .ZN(hmode_cnt_inst_n11) );
  AND2_X1 hmode_cnt_inst_U9 ( .A1(hmode_cnt_inst_n10), .A2(hmode_cnt_inst_n6), 
        .ZN(hmode_cnt_inst_N10) );
  NOR2_X1 hmode_cnt_inst_U8 ( .A1(s_tc_hmode), .A2(1'b0), .ZN(
        hmode_cnt_inst_n10) );
  XOR2_X1 hmode_cnt_inst_U7 ( .A(int_hmode_cnt[1]), .B(arv_k[1]), .Z(
        hmode_cnt_inst_n4) );
  XOR2_X1 hmode_cnt_inst_U6 ( .A(int_hmode_cnt[0]), .B(arv_k[0]), .Z(
        hmode_cnt_inst_n2) );
  XOR2_X1 hmode_cnt_inst_U5 ( .A(hmode_cnt_inst_q_2_), .B(arv_k[2]), .Z(
        hmode_cnt_inst_n1) );
  NOR3_X1 hmode_cnt_inst_U4 ( .A1(hmode_cnt_inst_n1), .A2(hmode_cnt_inst_n2), 
        .A3(hmode_cnt_inst_n4), .ZN(s_tc_hmode) );
  DFFR_X1 hmode_cnt_inst_cnt_out_reg_2_ ( .D(hmode_cnt_inst_N12), .CK(
        hmode_cnt_inst_net2826), .RN(hmode_cnt_inst_n12), .Q(
        hmode_cnt_inst_q_2_), .QN(hmode_cnt_inst_n5) );
  SDFFR_X1 hmode_cnt_inst_cnt_out_reg_1_ ( .D(hmode_cnt_inst_n10), .SI(1'b0), 
        .SE(hmode_cnt_inst_n11), .CK(hmode_cnt_inst_net2826), .RN(
        hmode_cnt_inst_n12), .Q(int_hmode_cnt[1]), .QN(hmode_cnt_inst_n7) );
  DFFR_X1 hmode_cnt_inst_cnt_out_reg_0_ ( .D(hmode_cnt_inst_N10), .CK(
        hmode_cnt_inst_net2826), .RN(hmode_cnt_inst_n12), .Q(int_hmode_cnt[0]), 
        .QN(hmode_cnt_inst_n6) );
  CLKGATETST_X1 hmode_cnt_inst_clk_gate_cnt_out_reg_latch ( .CK(ck), .E(
        int_en_hmode), .SE(1'b0), .GCK(hmode_cnt_inst_net2826) );
  INV_X1 vmode_cnt_inst_U14 ( .A(n10), .ZN(vmode_cnt_inst_n12) );
  AOI21_X1 vmode_cnt_inst_U13 ( .B1(vmode_cnt_inst_n10), .B2(vmode_cnt_inst_n7), .A(vmode_cnt_inst_N10), .ZN(vmode_cnt_inst_n8) );
  NAND4_X1 vmode_cnt_inst_U12 ( .A1(vmode_cnt_inst_n10), .A2(
        vmode_cnt_inst_q_1_), .A3(vmode_cnt_inst_q_0_), .A4(vmode_cnt_inst_n5), 
        .ZN(vmode_cnt_inst_n9) );
  OAI21_X1 vmode_cnt_inst_U11 ( .B1(vmode_cnt_inst_n8), .B2(vmode_cnt_inst_n5), 
        .A(vmode_cnt_inst_n9), .ZN(vmode_cnt_inst_N12) );
  XNOR2_X1 vmode_cnt_inst_U10 ( .A(vmode_cnt_inst_q_0_), .B(
        vmode_cnt_inst_q_1_), .ZN(vmode_cnt_inst_n11) );
  AND2_X1 vmode_cnt_inst_U9 ( .A1(vmode_cnt_inst_n10), .A2(vmode_cnt_inst_n6), 
        .ZN(vmode_cnt_inst_N10) );
  NOR2_X1 vmode_cnt_inst_U8 ( .A1(s_tc_vmode), .A2(1'b0), .ZN(
        vmode_cnt_inst_n10) );
  XOR2_X1 vmode_cnt_inst_U7 ( .A(vmode_cnt_inst_q_1_), .B(arv_k[1]), .Z(
        vmode_cnt_inst_n4) );
  XOR2_X1 vmode_cnt_inst_U6 ( .A(vmode_cnt_inst_q_0_), .B(arv_k[0]), .Z(
        vmode_cnt_inst_n2) );
  XOR2_X1 vmode_cnt_inst_U5 ( .A(vmode_cnt_inst_q_2_), .B(arv_k[2]), .Z(
        vmode_cnt_inst_n1) );
  NOR3_X1 vmode_cnt_inst_U4 ( .A1(vmode_cnt_inst_n1), .A2(vmode_cnt_inst_n2), 
        .A3(vmode_cnt_inst_n4), .ZN(s_tc_vmode) );
  DFFR_X1 vmode_cnt_inst_cnt_out_reg_2_ ( .D(vmode_cnt_inst_N12), .CK(
        vmode_cnt_inst_net2808), .RN(vmode_cnt_inst_n12), .Q(
        vmode_cnt_inst_q_2_), .QN(vmode_cnt_inst_n5) );
  SDFFR_X1 vmode_cnt_inst_cnt_out_reg_1_ ( .D(vmode_cnt_inst_n10), .SI(1'b0), 
        .SE(vmode_cnt_inst_n11), .CK(vmode_cnt_inst_net2808), .RN(
        vmode_cnt_inst_n12), .Q(vmode_cnt_inst_q_1_), .QN(vmode_cnt_inst_n7)
         );
  DFFR_X1 vmode_cnt_inst_cnt_out_reg_0_ ( .D(vmode_cnt_inst_N10), .CK(
        vmode_cnt_inst_net2808), .RN(vmode_cnt_inst_n12), .Q(
        vmode_cnt_inst_q_0_), .QN(vmode_cnt_inst_n6) );
  CLKGATETST_X1 vmode_cnt_inst_clk_gate_cnt_out_reg_latch ( .CK(ck), .E(
        int_en_vmode), .SE(1'b0), .GCK(vmode_cnt_inst_net2808) );
  INV_X1 res_cnt_inst_U14 ( .A(n10), .ZN(res_cnt_inst_n2) );
  XNOR2_X1 res_cnt_inst_U13 ( .A(res_cnt_inst_q_0_), .B(res_cnt_inst_q_1_), 
        .ZN(res_cnt_inst_n11) );
  AOI21_X1 res_cnt_inst_U12 ( .B1(res_cnt_inst_n10), .B2(res_cnt_inst_n7), .A(
        res_cnt_inst_N10), .ZN(res_cnt_inst_n8) );
  NAND4_X1 res_cnt_inst_U11 ( .A1(res_cnt_inst_n10), .A2(res_cnt_inst_q_1_), 
        .A3(res_cnt_inst_q_0_), .A4(res_cnt_inst_n5), .ZN(res_cnt_inst_n9) );
  OAI21_X1 res_cnt_inst_U10 ( .B1(res_cnt_inst_n8), .B2(res_cnt_inst_n5), .A(
        res_cnt_inst_n9), .ZN(res_cnt_inst_N12) );
  AND2_X1 res_cnt_inst_U9 ( .A1(res_cnt_inst_n10), .A2(res_cnt_inst_n1), .ZN(
        res_cnt_inst_N10) );
  XNOR2_X1 res_cnt_inst_U8 ( .A(res_cnt_inst_q_2_), .B(int_arv_res[2]), .ZN(
        res_cnt_inst_n12) );
  XNOR2_X1 res_cnt_inst_U7 ( .A(res_cnt_inst_q_1_), .B(int_arv_res[1]), .ZN(
        res_cnt_inst_n14) );
  XNOR2_X1 res_cnt_inst_U6 ( .A(res_cnt_inst_q_0_), .B(int_arv_res[0]), .ZN(
        res_cnt_inst_n13) );
  AND3_X1 res_cnt_inst_U5 ( .A1(res_cnt_inst_n12), .A2(res_cnt_inst_n13), .A3(
        res_cnt_inst_n14), .ZN(s_tc_res) );
  NOR2_X1 res_cnt_inst_U4 ( .A1(s_tc_res), .A2(1'b0), .ZN(res_cnt_inst_n10) );
  DFFR_X1 res_cnt_inst_cnt_out_reg_2_ ( .D(res_cnt_inst_N12), .CK(
        res_cnt_inst_net2790), .RN(res_cnt_inst_n2), .Q(res_cnt_inst_q_2_), 
        .QN(res_cnt_inst_n5) );
  SDFFR_X1 res_cnt_inst_cnt_out_reg_1_ ( .D(res_cnt_inst_n10), .SI(1'b0), .SE(
        res_cnt_inst_n11), .CK(res_cnt_inst_net2790), .RN(res_cnt_inst_n2), 
        .Q(res_cnt_inst_q_1_), .QN(res_cnt_inst_n7) );
  DFFR_X1 res_cnt_inst_cnt_out_reg_0_ ( .D(res_cnt_inst_N10), .CK(
        res_cnt_inst_net2790), .RN(res_cnt_inst_n2), .Q(res_cnt_inst_q_0_), 
        .QN(res_cnt_inst_n1) );
  CLKGATETST_X1 res_cnt_inst_clk_gate_cnt_out_reg_latch ( .CK(ck), .E(
        ctrl_wr_pipe), .SE(1'b0), .GCK(res_cnt_inst_net2790) );
  INV_X1 ifmaps_cnt_inst_U14 ( .A(n10), .ZN(ifmaps_cnt_inst_n12) );
  AND2_X1 ifmaps_cnt_inst_U13 ( .A1(ifmaps_cnt_inst_n10), .A2(
        ifmaps_cnt_inst_n6), .ZN(ifmaps_cnt_inst_N10) );
  XNOR2_X1 ifmaps_cnt_inst_U12 ( .A(int_ifmaps_ptr[0]), .B(int_ifmaps_ptr[1]), 
        .ZN(ifmaps_cnt_inst_n11) );
  AOI21_X1 ifmaps_cnt_inst_U11 ( .B1(ifmaps_cnt_inst_n10), .B2(
        ifmaps_cnt_inst_n7), .A(ifmaps_cnt_inst_N10), .ZN(ifmaps_cnt_inst_n8)
         );
  NAND4_X1 ifmaps_cnt_inst_U10 ( .A1(ifmaps_cnt_inst_n10), .A2(
        int_ifmaps_ptr[1]), .A3(int_ifmaps_ptr[0]), .A4(ifmaps_cnt_inst_n5), 
        .ZN(ifmaps_cnt_inst_n9) );
  OAI21_X1 ifmaps_cnt_inst_U9 ( .B1(ifmaps_cnt_inst_n8), .B2(
        ifmaps_cnt_inst_n5), .A(ifmaps_cnt_inst_n9), .ZN(ifmaps_cnt_inst_N12)
         );
  NOR2_X1 ifmaps_cnt_inst_U8 ( .A1(s_tc_ifmaps), .A2(1'b0), .ZN(
        ifmaps_cnt_inst_n10) );
  XOR2_X1 ifmaps_cnt_inst_U7 ( .A(int_ifmaps_ptr[1]), .B(arv_ifmaps[1]), .Z(
        ifmaps_cnt_inst_n4) );
  XOR2_X1 ifmaps_cnt_inst_U6 ( .A(int_ifmaps_ptr[0]), .B(arv_ifmaps[0]), .Z(
        ifmaps_cnt_inst_n2) );
  XOR2_X1 ifmaps_cnt_inst_U5 ( .A(int_ifmaps_ptr[2]), .B(arv_ifmaps[2]), .Z(
        ifmaps_cnt_inst_n1) );
  NOR3_X1 ifmaps_cnt_inst_U4 ( .A1(ifmaps_cnt_inst_n1), .A2(ifmaps_cnt_inst_n2), .A3(ifmaps_cnt_inst_n4), .ZN(s_tc_ifmaps) );
  DFFR_X1 ifmaps_cnt_inst_cnt_out_reg_2_ ( .D(ifmaps_cnt_inst_N12), .CK(
        ifmaps_cnt_inst_net2772), .RN(ifmaps_cnt_inst_n12), .Q(
        int_ifmaps_ptr[2]), .QN(ifmaps_cnt_inst_n5) );
  SDFFR_X1 ifmaps_cnt_inst_cnt_out_reg_1_ ( .D(ifmaps_cnt_inst_n10), .SI(1'b0), 
        .SE(ifmaps_cnt_inst_n11), .CK(ifmaps_cnt_inst_net2772), .RN(
        ifmaps_cnt_inst_n12), .Q(int_ifmaps_ptr[1]), .QN(ifmaps_cnt_inst_n7)
         );
  DFFR_X1 ifmaps_cnt_inst_cnt_out_reg_0_ ( .D(ifmaps_cnt_inst_N10), .CK(
        ifmaps_cnt_inst_net2772), .RN(ifmaps_cnt_inst_n12), .Q(
        int_ifmaps_ptr[0]), .QN(ifmaps_cnt_inst_n6) );
  CLKGATETST_X1 ifmaps_cnt_inst_clk_gate_cnt_out_reg_latch ( .CK(ck), .E(
        ctrl_en_npu), .SE(1'b0), .GCK(ifmaps_cnt_inst_net2772) );
  INV_X1 npu_cnt_inst_U14 ( .A(n10), .ZN(npu_cnt_inst_n12) );
  AOI21_X1 npu_cnt_inst_U13 ( .B1(npu_cnt_inst_n10), .B2(npu_cnt_inst_n7), .A(
        npu_cnt_inst_N10), .ZN(npu_cnt_inst_n8) );
  NAND4_X1 npu_cnt_inst_U12 ( .A1(npu_cnt_inst_n10), .A2(int_npu_ptr[1]), .A3(
        int_npu_ptr[0]), .A4(npu_cnt_inst_n5), .ZN(npu_cnt_inst_n9) );
  OAI21_X1 npu_cnt_inst_U11 ( .B1(npu_cnt_inst_n8), .B2(npu_cnt_inst_n5), .A(
        npu_cnt_inst_n9), .ZN(npu_cnt_inst_N12) );
  XNOR2_X1 npu_cnt_inst_U10 ( .A(int_npu_ptr[0]), .B(int_npu_ptr[1]), .ZN(
        npu_cnt_inst_n11) );
  AND2_X1 npu_cnt_inst_U9 ( .A1(npu_cnt_inst_n10), .A2(npu_cnt_inst_n6), .ZN(
        npu_cnt_inst_N10) );
  NOR2_X1 npu_cnt_inst_U8 ( .A1(s_tc_npu_ptr), .A2(1'b0), .ZN(npu_cnt_inst_n10) );
  XOR2_X1 npu_cnt_inst_U7 ( .A(int_npu_ptr[1]), .B(arv_npu[1]), .Z(
        npu_cnt_inst_n4) );
  XOR2_X1 npu_cnt_inst_U6 ( .A(int_npu_ptr[0]), .B(arv_npu[0]), .Z(
        npu_cnt_inst_n2) );
  XOR2_X1 npu_cnt_inst_U5 ( .A(int_npu_ptr[2]), .B(arv_npu[2]), .Z(
        npu_cnt_inst_n1) );
  NOR3_X1 npu_cnt_inst_U4 ( .A1(npu_cnt_inst_n1), .A2(npu_cnt_inst_n2), .A3(
        npu_cnt_inst_n4), .ZN(s_tc_npu_ptr) );
  DFFR_X1 npu_cnt_inst_cnt_out_reg_2_ ( .D(npu_cnt_inst_N12), .CK(
        npu_cnt_inst_net2754), .RN(npu_cnt_inst_n12), .Q(int_npu_ptr[2]), .QN(
        npu_cnt_inst_n5) );
  SDFFR_X1 npu_cnt_inst_cnt_out_reg_1_ ( .D(npu_cnt_inst_n10), .SI(1'b0), .SE(
        npu_cnt_inst_n11), .CK(npu_cnt_inst_net2754), .RN(npu_cnt_inst_n12), 
        .Q(int_npu_ptr[1]), .QN(npu_cnt_inst_n7) );
  DFFR_X1 npu_cnt_inst_cnt_out_reg_0_ ( .D(npu_cnt_inst_N10), .CK(
        npu_cnt_inst_net2754), .RN(npu_cnt_inst_n12), .Q(int_npu_ptr[0]), .QN(
        npu_cnt_inst_n6) );
  CLKGATETST_X1 npu_cnt_inst_clk_gate_cnt_out_reg_latch ( .CK(ck), .E(
        int_en_npu_ptr), .SE(1'b0), .GCK(npu_cnt_inst_net2754) );
  INV_X1 tilev_cnt_inst_U16 ( .A(n9), .ZN(tilev_cnt_inst_n3) );
  INV_X1 tilev_cnt_inst_U15 ( .A(arv_tile[0]), .ZN(tilev_cnt_inst_n8) );
  NOR2_X1 tilev_cnt_inst_U14 ( .A1(1'b0), .A2(tilev_cnt_inst_q_0_), .ZN(
        tilev_cnt_inst_n13) );
  OAI211_X1 tilev_cnt_inst_U13 ( .C1(arv_tile[0]), .C2(tilev_cnt_inst_n12), 
        .A(int_en_tilev_ptr), .B(tilev_cnt_inst_n13), .ZN(tilev_cnt_inst_n11)
         );
  OAI21_X1 tilev_cnt_inst_U12 ( .B1(int_en_tilev_ptr), .B2(tilev_cnt_inst_n2), 
        .A(tilev_cnt_inst_n11), .ZN(tilev_cnt_inst_n17) );
  OAI21_X1 tilev_cnt_inst_U11 ( .B1(tilev_cnt_inst_n8), .B2(arv_tile[1]), .A(
        tilev_cnt_inst_n1), .ZN(tilev_cnt_inst_n9) );
  AND2_X1 tilev_cnt_inst_U10 ( .A1(int_en_tilev_ptr), .A2(tilev_cnt_inst_q_0_), 
        .ZN(tilev_cnt_inst_n5) );
  XNOR2_X1 tilev_cnt_inst_U9 ( .A(tilev_cnt_inst_n2), .B(arv_tile[0]), .ZN(
        tilev_cnt_inst_n14) );
  NOR2_X1 tilev_cnt_inst_U8 ( .A1(tilev_cnt_inst_n12), .A2(tilev_cnt_inst_n14), 
        .ZN(int_d_tc[2]) );
  INV_X1 tilev_cnt_inst_U7 ( .A(tilev_cnt_inst_n9), .ZN(tilev_cnt_inst_n6) );
  AOI21_X1 tilev_cnt_inst_U6 ( .B1(arv_tile[1]), .B2(tilev_cnt_inst_n8), .A(
        tilev_cnt_inst_q_0_), .ZN(tilev_cnt_inst_n7) );
  AOI22_X1 tilev_cnt_inst_U5 ( .A1(tilev_cnt_inst_n5), .A2(tilev_cnt_inst_n6), 
        .B1(tilev_cnt_inst_n7), .B2(tilev_cnt_inst_q_1_), .ZN(
        tilev_cnt_inst_n4) );
  OAI22_X1 tilev_cnt_inst_U4 ( .A1(int_en_tilev_ptr), .A2(tilev_cnt_inst_n1), 
        .B1(1'b0), .B2(tilev_cnt_inst_n4), .ZN(tilev_cnt_inst_n15) );
  XNOR2_X1 tilev_cnt_inst_U3 ( .A(arv_tile[1]), .B(tilev_cnt_inst_n1), .ZN(
        tilev_cnt_inst_n12) );
  DFFR_X1 tilev_cnt_inst_cnt_out_reg_1_ ( .D(tilev_cnt_inst_n15), .CK(ck), 
        .RN(tilev_cnt_inst_n3), .Q(tilev_cnt_inst_q_1_), .QN(tilev_cnt_inst_n1) );
  DFFR_X1 tilev_cnt_inst_cnt_out_reg_0_ ( .D(tilev_cnt_inst_n17), .CK(ck), 
        .RN(tilev_cnt_inst_n3), .Q(tilev_cnt_inst_q_0_), .QN(tilev_cnt_inst_n2) );
  INV_X1 tileh_cnt_inst_U16 ( .A(n10), .ZN(tileh_cnt_inst_n1) );
  INV_X1 tileh_cnt_inst_U15 ( .A(arv_tile[0]), .ZN(tileh_cnt_inst_n8) );
  XNOR2_X1 tileh_cnt_inst_U14 ( .A(tileh_cnt_inst_n2), .B(arv_tile[0]), .ZN(
        tileh_cnt_inst_n17) );
  NOR2_X1 tileh_cnt_inst_U13 ( .A1(tileh_cnt_inst_n19), .A2(tileh_cnt_inst_n17), .ZN(int_d_tc[1]) );
  OAI21_X1 tileh_cnt_inst_U12 ( .B1(tileh_cnt_inst_n8), .B2(arv_tile[1]), .A(
        tileh_cnt_inst_n6), .ZN(tileh_cnt_inst_n21) );
  XNOR2_X1 tileh_cnt_inst_U11 ( .A(arv_tile[1]), .B(tileh_cnt_inst_n6), .ZN(
        tileh_cnt_inst_n19) );
  AND2_X1 tileh_cnt_inst_U10 ( .A1(n15), .A2(i_data_ev_odd_n), .ZN(
        tileh_cnt_inst_n23) );
  NOR2_X1 tileh_cnt_inst_U9 ( .A1(1'b0), .A2(i_data_ev_odd_n), .ZN(
        tileh_cnt_inst_n18) );
  OAI211_X1 tileh_cnt_inst_U8 ( .C1(arv_tile[0]), .C2(tileh_cnt_inst_n19), .A(
        n15), .B(tileh_cnt_inst_n18), .ZN(tileh_cnt_inst_n20) );
  OAI21_X1 tileh_cnt_inst_U7 ( .B1(n15), .B2(tileh_cnt_inst_n2), .A(
        tileh_cnt_inst_n20), .ZN(tileh_cnt_inst_n10) );
  INV_X1 tileh_cnt_inst_U6 ( .A(tileh_cnt_inst_n21), .ZN(tileh_cnt_inst_n3) );
  AOI21_X1 tileh_cnt_inst_U5 ( .B1(arv_tile[1]), .B2(tileh_cnt_inst_n8), .A(
        i_data_ev_odd_n), .ZN(tileh_cnt_inst_n22) );
  AOI22_X1 tileh_cnt_inst_U4 ( .A1(tileh_cnt_inst_n23), .A2(tileh_cnt_inst_n3), 
        .B1(tileh_cnt_inst_n22), .B2(tileh_cnt_inst_q_1_), .ZN(
        tileh_cnt_inst_n24) );
  OAI22_X1 tileh_cnt_inst_U3 ( .A1(n15), .A2(tileh_cnt_inst_n6), .B1(1'b0), 
        .B2(tileh_cnt_inst_n24), .ZN(tileh_cnt_inst_n16) );
  DFFR_X1 tileh_cnt_inst_cnt_out_reg_1_ ( .D(tileh_cnt_inst_n16), .CK(ck), 
        .RN(tileh_cnt_inst_n1), .Q(tileh_cnt_inst_q_1_), .QN(tileh_cnt_inst_n6) );
  DFFR_X1 tileh_cnt_inst_cnt_out_reg_0_ ( .D(tileh_cnt_inst_n10), .CK(ck), 
        .RN(tileh_cnt_inst_n1), .Q(i_data_ev_odd_n), .QN(tileh_cnt_inst_n2) );
  INV_X1 ofmaps_cnt_inst_U17 ( .A(n10), .ZN(ofmaps_cnt_inst_n2) );
  XNOR2_X1 ofmaps_cnt_inst_U16 ( .A(ofmaps_cnt_inst_q_0_), .B(
        ofmaps_cnt_inst_q_1_), .ZN(ofmaps_cnt_inst_n15) );
  AND2_X1 ofmaps_cnt_inst_U15 ( .A1(ofmaps_cnt_inst_n13), .A2(
        ofmaps_cnt_inst_n1), .ZN(ofmaps_cnt_inst_N11) );
  XNOR2_X1 ofmaps_cnt_inst_U14 ( .A(ofmaps_cnt_inst_q_3_), .B(arv_ofmaps[3]), 
        .ZN(ofmaps_cnt_inst_n18) );
  XNOR2_X1 ofmaps_cnt_inst_U13 ( .A(ofmaps_cnt_inst_q_2_), .B(arv_ofmaps[2]), 
        .ZN(ofmaps_cnt_inst_n17) );
  AND4_X1 ofmaps_cnt_inst_U12 ( .A1(ofmaps_cnt_inst_n16), .A2(
        ofmaps_cnt_inst_n17), .A3(ofmaps_cnt_inst_n18), .A4(
        ofmaps_cnt_inst_n19), .ZN(int_d_tc[0]) );
  XNOR2_X1 ofmaps_cnt_inst_U11 ( .A(ofmaps_cnt_inst_q_0_), .B(arv_ofmaps[0]), 
        .ZN(ofmaps_cnt_inst_n19) );
  INV_X1 ofmaps_cnt_inst_U10 ( .A(ofmaps_cnt_inst_n14), .ZN(ofmaps_cnt_inst_n4) );
  AOI21_X1 ofmaps_cnt_inst_U9 ( .B1(ofmaps_cnt_inst_n13), .B2(
        ofmaps_cnt_inst_n8), .A(ofmaps_cnt_inst_n4), .ZN(ofmaps_cnt_inst_n10)
         );
  OR3_X1 ofmaps_cnt_inst_U8 ( .A1(ofmaps_cnt_inst_n8), .A2(
        ofmaps_cnt_inst_q_3_), .A3(ofmaps_cnt_inst_n12), .ZN(
        ofmaps_cnt_inst_n11) );
  OAI21_X1 ofmaps_cnt_inst_U7 ( .B1(ofmaps_cnt_inst_n10), .B2(
        ofmaps_cnt_inst_n5), .A(ofmaps_cnt_inst_n11), .ZN(ofmaps_cnt_inst_N14)
         );
  OAI22_X1 ofmaps_cnt_inst_U6 ( .A1(ofmaps_cnt_inst_n14), .A2(
        ofmaps_cnt_inst_n8), .B1(ofmaps_cnt_inst_q_2_), .B2(
        ofmaps_cnt_inst_n12), .ZN(ofmaps_cnt_inst_N13) );
  AOI21_X1 ofmaps_cnt_inst_U5 ( .B1(ofmaps_cnt_inst_n9), .B2(
        ofmaps_cnt_inst_n13), .A(ofmaps_cnt_inst_N11), .ZN(ofmaps_cnt_inst_n14) );
  NOR2_X1 ofmaps_cnt_inst_U4 ( .A1(int_d_tc[0]), .A2(1'b0), .ZN(
        ofmaps_cnt_inst_n13) );
  XOR2_X1 ofmaps_cnt_inst_U20 ( .A(ofmaps_cnt_inst_n9), .B(arv_ofmaps[1]), .Z(
        ofmaps_cnt_inst_n16) );
  NAND3_X1 ofmaps_cnt_inst_U19 ( .A1(ofmaps_cnt_inst_q_1_), .A2(
        ofmaps_cnt_inst_q_0_), .A3(ofmaps_cnt_inst_n13), .ZN(
        ofmaps_cnt_inst_n12) );
  DFFR_X1 ofmaps_cnt_inst_cnt_out_reg_3_ ( .D(ofmaps_cnt_inst_N14), .CK(
        ofmaps_cnt_inst_net2736), .RN(ofmaps_cnt_inst_n2), .Q(
        ofmaps_cnt_inst_q_3_), .QN(ofmaps_cnt_inst_n5) );
  DFFR_X1 ofmaps_cnt_inst_cnt_out_reg_2_ ( .D(ofmaps_cnt_inst_N13), .CK(
        ofmaps_cnt_inst_net2736), .RN(ofmaps_cnt_inst_n2), .Q(
        ofmaps_cnt_inst_q_2_), .QN(ofmaps_cnt_inst_n8) );
  SDFFR_X1 ofmaps_cnt_inst_cnt_out_reg_1_ ( .D(ofmaps_cnt_inst_n13), .SI(1'b0), 
        .SE(ofmaps_cnt_inst_n15), .CK(ofmaps_cnt_inst_net2736), .RN(
        ofmaps_cnt_inst_n2), .Q(ofmaps_cnt_inst_q_1_), .QN(ofmaps_cnt_inst_n9)
         );
  DFFR_X1 ofmaps_cnt_inst_cnt_out_reg_0_ ( .D(ofmaps_cnt_inst_N11), .CK(
        ofmaps_cnt_inst_net2736), .RN(ofmaps_cnt_inst_n2), .Q(
        ofmaps_cnt_inst_q_0_), .QN(ofmaps_cnt_inst_n1) );
  CLKGATETST_X1 ofmaps_cnt_inst_clk_gate_cnt_out_reg_latch ( .CK(ck), .E(
        int_rst_i_data_addr), .SE(1'b0), .GCK(ofmaps_cnt_inst_net2736) );
  AOI21_X1 i_data_addr_gen_inst_U42 ( .B1(ctrl_ldh_v_n), .B2(
        int_inc_i_data_odd), .A(int_rst_i_data_addr), .ZN(
        i_data_addr_gen_inst_n30) );
  INV_X1 i_data_addr_gen_inst_U41 ( .A(i_data_addr_gen_inst_n30), .ZN(
        i_data_addr_gen_inst_n26) );
  AOI21_X1 i_data_addr_gen_inst_U40 ( .B1(ctrl_ldh_v_n), .B2(
        int_inc_i_data_even), .A(int_rst_i_data_addr), .ZN(
        i_data_addr_gen_inst_n31) );
  INV_X1 i_data_addr_gen_inst_U39 ( .A(i_data_addr_gen_inst_n31), .ZN(
        i_data_addr_gen_inst_n25) );
  AND2_X1 i_data_addr_gen_inst_U38 ( .A1(i_data_addr_gen_inst_N58), .A2(
        i_data_addr_gen_inst_n29), .ZN(i_data_addr_gen_inst_N68) );
  AND2_X1 i_data_addr_gen_inst_U37 ( .A1(i_data_addr_gen_inst_N67), .A2(
        i_data_addr_gen_inst_n29), .ZN(i_data_addr_gen_inst_N77) );
  INV_X1 i_data_addr_gen_inst_U36 ( .A(n9), .ZN(i_data_addr_gen_inst_n24) );
  AND2_X1 i_data_addr_gen_inst_U35 ( .A1(i_data_addr_gen_inst_N59), .A2(
        i_data_addr_gen_inst_n29), .ZN(i_data_addr_gen_inst_N69) );
  AND2_X1 i_data_addr_gen_inst_U34 ( .A1(i_data_addr_gen_inst_N60), .A2(
        i_data_addr_gen_inst_n29), .ZN(i_data_addr_gen_inst_N70) );
  AND2_X1 i_data_addr_gen_inst_U33 ( .A1(i_data_addr_gen_inst_N61), .A2(
        i_data_addr_gen_inst_n29), .ZN(i_data_addr_gen_inst_N71) );
  AND2_X1 i_data_addr_gen_inst_U32 ( .A1(i_data_addr_gen_inst_N62), .A2(
        i_data_addr_gen_inst_n29), .ZN(i_data_addr_gen_inst_N72) );
  AND2_X1 i_data_addr_gen_inst_U31 ( .A1(i_data_addr_gen_inst_N63), .A2(
        i_data_addr_gen_inst_n29), .ZN(i_data_addr_gen_inst_N73) );
  AND2_X1 i_data_addr_gen_inst_U30 ( .A1(i_data_addr_gen_inst_N64), .A2(
        i_data_addr_gen_inst_n29), .ZN(i_data_addr_gen_inst_N74) );
  AND2_X1 i_data_addr_gen_inst_U29 ( .A1(i_data_addr_gen_inst_N65), .A2(
        i_data_addr_gen_inst_n29), .ZN(i_data_addr_gen_inst_N75) );
  AND2_X1 i_data_addr_gen_inst_U28 ( .A1(i_data_addr_gen_inst_N66), .A2(
        i_data_addr_gen_inst_n29), .ZN(i_data_addr_gen_inst_N76) );
  NOR2_X1 i_data_addr_gen_inst_U27 ( .A1(int_inc_i_data_odd), .A2(
        int_inc_i_data_even), .ZN(i_data_addr_gen_inst_n29) );
  BUF_X1 i_data_addr_gen_inst_U26 ( .A(i_data_addr_gen_inst_n24), .Z(
        i_data_addr_gen_inst_n23) );
  INV_X1 i_data_addr_gen_inst_U25 ( .A(int_rst_i_data_addr), .ZN(
        i_data_addr_gen_inst_n27) );
  SDFFR_X1 i_data_addr_gen_inst_int_data_even_base_addr_reg_9_ ( .D(1'b0), 
        .SI(i_data_addr_gen_inst_n27), .SE(i_data_addr_gen_inst_N17), .CK(
        i_data_addr_gen_inst_net2708), .RN(i_data_addr_gen_inst_n24), .Q(
        i_data_addr_gen_inst_int_data_even_base_addr[9]) );
  SDFFR_X1 i_data_addr_gen_inst_int_data_odd_base_addr_reg_9_ ( .D(1'b0), .SI(
        i_data_addr_gen_inst_n27), .SE(i_data_addr_gen_inst_N39), .CK(
        i_data_addr_gen_inst_net2714), .RN(i_data_addr_gen_inst_n24), .Q(
        i_data_addr_gen_inst_int_data_odd_base_addr[9]) );
  SDFFR_X1 i_data_addr_gen_inst_int_data_even_base_addr_reg_0_ ( .D(1'b0), 
        .SI(i_data_addr_gen_inst_n27), .SE(i_data_addr_gen_inst_N8), .CK(
        i_data_addr_gen_inst_net2708), .RN(i_data_addr_gen_inst_n24), .Q(
        i_data_addr_gen_inst_int_data_even_base_addr[0]) );
  SDFFR_X1 i_data_addr_gen_inst_int_data_even_base_addr_reg_1_ ( .D(1'b0), 
        .SI(i_data_addr_gen_inst_n27), .SE(i_data_addr_gen_inst_N9), .CK(
        i_data_addr_gen_inst_net2708), .RN(i_data_addr_gen_inst_n24), .Q(
        i_data_addr_gen_inst_int_data_even_base_addr[1]) );
  SDFFR_X1 i_data_addr_gen_inst_int_data_even_base_addr_reg_2_ ( .D(1'b0), 
        .SI(i_data_addr_gen_inst_n27), .SE(i_data_addr_gen_inst_N10), .CK(
        i_data_addr_gen_inst_net2708), .RN(i_data_addr_gen_inst_n24), .Q(
        i_data_addr_gen_inst_int_data_even_base_addr[2]) );
  SDFFR_X1 i_data_addr_gen_inst_int_data_even_base_addr_reg_3_ ( .D(1'b0), 
        .SI(i_data_addr_gen_inst_n27), .SE(i_data_addr_gen_inst_N11), .CK(
        i_data_addr_gen_inst_net2708), .RN(i_data_addr_gen_inst_n24), .Q(
        i_data_addr_gen_inst_int_data_even_base_addr[3]) );
  SDFFR_X1 i_data_addr_gen_inst_int_data_even_base_addr_reg_4_ ( .D(1'b0), 
        .SI(i_data_addr_gen_inst_n27), .SE(i_data_addr_gen_inst_N12), .CK(
        i_data_addr_gen_inst_net2708), .RN(i_data_addr_gen_inst_n24), .Q(
        i_data_addr_gen_inst_int_data_even_base_addr[4]) );
  SDFFR_X1 i_data_addr_gen_inst_int_data_even_base_addr_reg_5_ ( .D(1'b0), 
        .SI(i_data_addr_gen_inst_n27), .SE(i_data_addr_gen_inst_N13), .CK(
        i_data_addr_gen_inst_net2708), .RN(i_data_addr_gen_inst_n24), .Q(
        i_data_addr_gen_inst_int_data_even_base_addr[5]) );
  SDFFR_X1 i_data_addr_gen_inst_int_data_even_base_addr_reg_6_ ( .D(1'b0), 
        .SI(i_data_addr_gen_inst_n27), .SE(i_data_addr_gen_inst_N14), .CK(
        i_data_addr_gen_inst_net2708), .RN(i_data_addr_gen_inst_n24), .Q(
        i_data_addr_gen_inst_int_data_even_base_addr[6]) );
  SDFFR_X1 i_data_addr_gen_inst_int_data_even_base_addr_reg_7_ ( .D(1'b0), 
        .SI(i_data_addr_gen_inst_n27), .SE(i_data_addr_gen_inst_N15), .CK(
        i_data_addr_gen_inst_net2708), .RN(i_data_addr_gen_inst_n24), .Q(
        i_data_addr_gen_inst_int_data_even_base_addr[7]) );
  SDFFR_X1 i_data_addr_gen_inst_int_data_even_base_addr_reg_8_ ( .D(1'b0), 
        .SI(i_data_addr_gen_inst_n27), .SE(i_data_addr_gen_inst_N16), .CK(
        i_data_addr_gen_inst_net2708), .RN(i_data_addr_gen_inst_n24), .Q(
        i_data_addr_gen_inst_int_data_even_base_addr[8]) );
  SDFFR_X1 i_data_addr_gen_inst_int_data_odd_base_addr_reg_0_ ( .D(1'b0), .SI(
        i_data_addr_gen_inst_n27), .SE(i_data_addr_gen_inst_N30), .CK(
        i_data_addr_gen_inst_net2714), .RN(i_data_addr_gen_inst_n24), .Q(
        i_data_addr_gen_inst_int_data_odd_base_addr[0]) );
  SDFFR_X1 i_data_addr_gen_inst_int_data_odd_base_addr_reg_1_ ( .D(1'b0), .SI(
        i_data_addr_gen_inst_n27), .SE(i_data_addr_gen_inst_N31), .CK(
        i_data_addr_gen_inst_net2714), .RN(i_data_addr_gen_inst_n24), .Q(
        i_data_addr_gen_inst_int_data_odd_base_addr[1]) );
  SDFFR_X1 i_data_addr_gen_inst_int_data_odd_base_addr_reg_2_ ( .D(1'b0), .SI(
        i_data_addr_gen_inst_n27), .SE(i_data_addr_gen_inst_N32), .CK(
        i_data_addr_gen_inst_net2714), .RN(i_data_addr_gen_inst_n24), .Q(
        i_data_addr_gen_inst_int_data_odd_base_addr[2]) );
  SDFFR_X1 i_data_addr_gen_inst_int_data_odd_base_addr_reg_3_ ( .D(1'b0), .SI(
        i_data_addr_gen_inst_n27), .SE(i_data_addr_gen_inst_N33), .CK(
        i_data_addr_gen_inst_net2714), .RN(i_data_addr_gen_inst_n24), .Q(
        i_data_addr_gen_inst_int_data_odd_base_addr[3]) );
  SDFFR_X1 i_data_addr_gen_inst_int_data_odd_base_addr_reg_4_ ( .D(1'b0), .SI(
        i_data_addr_gen_inst_n27), .SE(i_data_addr_gen_inst_N34), .CK(
        i_data_addr_gen_inst_net2714), .RN(i_data_addr_gen_inst_n24), .Q(
        i_data_addr_gen_inst_int_data_odd_base_addr[4]) );
  SDFFR_X1 i_data_addr_gen_inst_int_data_odd_base_addr_reg_5_ ( .D(1'b0), .SI(
        i_data_addr_gen_inst_n27), .SE(i_data_addr_gen_inst_N35), .CK(
        i_data_addr_gen_inst_net2714), .RN(i_data_addr_gen_inst_n24), .Q(
        i_data_addr_gen_inst_int_data_odd_base_addr[5]) );
  SDFFR_X1 i_data_addr_gen_inst_int_data_odd_base_addr_reg_6_ ( .D(1'b0), .SI(
        i_data_addr_gen_inst_n27), .SE(i_data_addr_gen_inst_N36), .CK(
        i_data_addr_gen_inst_net2714), .RN(i_data_addr_gen_inst_n24), .Q(
        i_data_addr_gen_inst_int_data_odd_base_addr[6]) );
  SDFFR_X1 i_data_addr_gen_inst_int_data_odd_base_addr_reg_7_ ( .D(1'b0), .SI(
        i_data_addr_gen_inst_n27), .SE(i_data_addr_gen_inst_N37), .CK(
        i_data_addr_gen_inst_net2714), .RN(i_data_addr_gen_inst_n24), .Q(
        i_data_addr_gen_inst_int_data_odd_base_addr[7]) );
  SDFFR_X1 i_data_addr_gen_inst_int_data_odd_base_addr_reg_8_ ( .D(1'b0), .SI(
        i_data_addr_gen_inst_n27), .SE(i_data_addr_gen_inst_N38), .CK(
        i_data_addr_gen_inst_net2714), .RN(i_data_addr_gen_inst_n24), .Q(
        i_data_addr_gen_inst_int_data_odd_base_addr[8]) );
  DFFR_X1 i_data_addr_gen_inst_int_data_offs_addr_reg_9_ ( .D(
        i_data_addr_gen_inst_N77), .CK(i_data_addr_gen_inst_net2719), .RN(
        i_data_addr_gen_inst_n23), .Q(
        i_data_addr_gen_inst_int_data_offs_addr_9_) );
  DFFR_X1 i_data_addr_gen_inst_int_data_offs_addr_reg_8_ ( .D(
        i_data_addr_gen_inst_N76), .CK(i_data_addr_gen_inst_net2719), .RN(
        i_data_addr_gen_inst_n23), .Q(
        i_data_addr_gen_inst_int_data_offs_addr_8_) );
  DFFR_X1 i_data_addr_gen_inst_int_data_offs_addr_reg_7_ ( .D(
        i_data_addr_gen_inst_N75), .CK(i_data_addr_gen_inst_net2719), .RN(
        i_data_addr_gen_inst_n23), .Q(
        i_data_addr_gen_inst_int_data_offs_addr_7_) );
  DFFR_X1 i_data_addr_gen_inst_int_data_offs_addr_reg_6_ ( .D(
        i_data_addr_gen_inst_N74), .CK(i_data_addr_gen_inst_net2719), .RN(
        i_data_addr_gen_inst_n23), .Q(
        i_data_addr_gen_inst_int_data_offs_addr_6_) );
  DFFR_X1 i_data_addr_gen_inst_int_data_offs_addr_reg_5_ ( .D(
        i_data_addr_gen_inst_N73), .CK(i_data_addr_gen_inst_net2719), .RN(
        i_data_addr_gen_inst_n23), .Q(
        i_data_addr_gen_inst_int_data_offs_addr_5_) );
  DFFR_X1 i_data_addr_gen_inst_int_data_offs_addr_reg_4_ ( .D(
        i_data_addr_gen_inst_N72), .CK(i_data_addr_gen_inst_net2719), .RN(
        i_data_addr_gen_inst_n23), .Q(
        i_data_addr_gen_inst_int_data_offs_addr_4_) );
  DFFR_X1 i_data_addr_gen_inst_int_data_offs_addr_reg_3_ ( .D(
        i_data_addr_gen_inst_N71), .CK(i_data_addr_gen_inst_net2719), .RN(
        i_data_addr_gen_inst_n23), .Q(
        i_data_addr_gen_inst_int_data_offs_addr_3_) );
  DFFR_X1 i_data_addr_gen_inst_int_data_offs_addr_reg_2_ ( .D(
        i_data_addr_gen_inst_N70), .CK(i_data_addr_gen_inst_net2719), .RN(
        i_data_addr_gen_inst_n23), .Q(
        i_data_addr_gen_inst_int_data_offs_addr_2_) );
  DFFR_X1 i_data_addr_gen_inst_int_data_offs_addr_reg_1_ ( .D(
        i_data_addr_gen_inst_N69), .CK(i_data_addr_gen_inst_net2719), .RN(
        i_data_addr_gen_inst_n23), .Q(
        i_data_addr_gen_inst_int_data_offs_addr_1_) );
  DFFR_X1 i_data_addr_gen_inst_int_data_offs_addr_reg_0_ ( .D(
        i_data_addr_gen_inst_N68), .CK(i_data_addr_gen_inst_net2719), .RN(
        i_data_addr_gen_inst_n23), .Q(
        i_data_addr_gen_inst_int_data_offs_addr_0_) );
  CLKGATETST_X1 i_data_addr_gen_inst_clk_gate_int_data_even_base_addr_reg_latch ( 
        .CK(ck), .E(i_data_addr_gen_inst_n25), .SE(1'b0), .GCK(
        i_data_addr_gen_inst_net2708) );
  CLKGATETST_X1 i_data_addr_gen_inst_clk_gate_int_data_odd_base_addr_reg_latch ( 
        .CK(ck), .E(i_data_addr_gen_inst_n26), .SE(1'b0), .GCK(
        i_data_addr_gen_inst_net2714) );
  CLKGATETST_X1 i_data_addr_gen_inst_clk_gate_int_data_offs_addr_reg_latch ( 
        .CK(ck), .E(ctrl_ldh_v_n), .SE(1'b0), .GCK(
        i_data_addr_gen_inst_net2719) );
  XOR2_X1 i_data_addr_gen_inst_add_78_U2 ( .A(
        i_data_addr_gen_inst_add_78_carry[9]), .B(
        i_data_addr_gen_inst_int_data_offs_addr_9_), .Z(
        i_data_addr_gen_inst_N67) );
  INV_X1 i_data_addr_gen_inst_add_78_U1 ( .A(
        i_data_addr_gen_inst_int_data_offs_addr_0_), .ZN(
        i_data_addr_gen_inst_N58) );
  HA_X1 i_data_addr_gen_inst_add_78_U1_1_1 ( .A(
        i_data_addr_gen_inst_int_data_offs_addr_1_), .B(
        i_data_addr_gen_inst_int_data_offs_addr_0_), .CO(
        i_data_addr_gen_inst_add_78_carry[2]), .S(i_data_addr_gen_inst_N59) );
  HA_X1 i_data_addr_gen_inst_add_78_U1_1_2 ( .A(
        i_data_addr_gen_inst_int_data_offs_addr_2_), .B(
        i_data_addr_gen_inst_add_78_carry[2]), .CO(
        i_data_addr_gen_inst_add_78_carry[3]), .S(i_data_addr_gen_inst_N60) );
  HA_X1 i_data_addr_gen_inst_add_78_U1_1_3 ( .A(
        i_data_addr_gen_inst_int_data_offs_addr_3_), .B(
        i_data_addr_gen_inst_add_78_carry[3]), .CO(
        i_data_addr_gen_inst_add_78_carry[4]), .S(i_data_addr_gen_inst_N61) );
  HA_X1 i_data_addr_gen_inst_add_78_U1_1_4 ( .A(
        i_data_addr_gen_inst_int_data_offs_addr_4_), .B(
        i_data_addr_gen_inst_add_78_carry[4]), .CO(
        i_data_addr_gen_inst_add_78_carry[5]), .S(i_data_addr_gen_inst_N62) );
  HA_X1 i_data_addr_gen_inst_add_78_U1_1_5 ( .A(
        i_data_addr_gen_inst_int_data_offs_addr_5_), .B(
        i_data_addr_gen_inst_add_78_carry[5]), .CO(
        i_data_addr_gen_inst_add_78_carry[6]), .S(i_data_addr_gen_inst_N63) );
  HA_X1 i_data_addr_gen_inst_add_78_U1_1_6 ( .A(
        i_data_addr_gen_inst_int_data_offs_addr_6_), .B(
        i_data_addr_gen_inst_add_78_carry[6]), .CO(
        i_data_addr_gen_inst_add_78_carry[7]), .S(i_data_addr_gen_inst_N64) );
  HA_X1 i_data_addr_gen_inst_add_78_U1_1_7 ( .A(
        i_data_addr_gen_inst_int_data_offs_addr_7_), .B(
        i_data_addr_gen_inst_add_78_carry[7]), .CO(
        i_data_addr_gen_inst_add_78_carry[8]), .S(i_data_addr_gen_inst_N65) );
  HA_X1 i_data_addr_gen_inst_add_78_U1_1_8 ( .A(
        i_data_addr_gen_inst_int_data_offs_addr_8_), .B(
        i_data_addr_gen_inst_add_78_carry[8]), .CO(
        i_data_addr_gen_inst_add_78_carry[9]), .S(i_data_addr_gen_inst_N66) );
  XOR2_X1 i_data_addr_gen_inst_add_62_U2 ( .A(
        i_data_addr_gen_inst_add_62_carry[9]), .B(i_data_odd_addr[9]), .Z(
        i_data_addr_gen_inst_N39) );
  INV_X1 i_data_addr_gen_inst_add_62_U1 ( .A(i_data_odd_addr[0]), .ZN(
        i_data_addr_gen_inst_N30) );
  HA_X1 i_data_addr_gen_inst_add_62_U1_1_1 ( .A(i_data_odd_addr[1]), .B(
        i_data_odd_addr[0]), .CO(i_data_addr_gen_inst_add_62_carry[2]), .S(
        i_data_addr_gen_inst_N31) );
  HA_X1 i_data_addr_gen_inst_add_62_U1_1_2 ( .A(i_data_odd_addr[2]), .B(
        i_data_addr_gen_inst_add_62_carry[2]), .CO(
        i_data_addr_gen_inst_add_62_carry[3]), .S(i_data_addr_gen_inst_N32) );
  HA_X1 i_data_addr_gen_inst_add_62_U1_1_3 ( .A(i_data_odd_addr[3]), .B(
        i_data_addr_gen_inst_add_62_carry[3]), .CO(
        i_data_addr_gen_inst_add_62_carry[4]), .S(i_data_addr_gen_inst_N33) );
  HA_X1 i_data_addr_gen_inst_add_62_U1_1_4 ( .A(i_data_odd_addr[4]), .B(
        i_data_addr_gen_inst_add_62_carry[4]), .CO(
        i_data_addr_gen_inst_add_62_carry[5]), .S(i_data_addr_gen_inst_N34) );
  HA_X1 i_data_addr_gen_inst_add_62_U1_1_5 ( .A(i_data_odd_addr[5]), .B(
        i_data_addr_gen_inst_add_62_carry[5]), .CO(
        i_data_addr_gen_inst_add_62_carry[6]), .S(i_data_addr_gen_inst_N35) );
  HA_X1 i_data_addr_gen_inst_add_62_U1_1_6 ( .A(i_data_odd_addr[6]), .B(
        i_data_addr_gen_inst_add_62_carry[6]), .CO(
        i_data_addr_gen_inst_add_62_carry[7]), .S(i_data_addr_gen_inst_N36) );
  HA_X1 i_data_addr_gen_inst_add_62_U1_1_7 ( .A(i_data_odd_addr[7]), .B(
        i_data_addr_gen_inst_add_62_carry[7]), .CO(
        i_data_addr_gen_inst_add_62_carry[8]), .S(i_data_addr_gen_inst_N37) );
  HA_X1 i_data_addr_gen_inst_add_62_U1_1_8 ( .A(i_data_odd_addr[8]), .B(
        i_data_addr_gen_inst_add_62_carry[8]), .CO(
        i_data_addr_gen_inst_add_62_carry[9]), .S(i_data_addr_gen_inst_N38) );
  XOR2_X1 i_data_addr_gen_inst_add_46_U2 ( .A(
        i_data_addr_gen_inst_add_46_carry[9]), .B(i_data_even_addr[9]), .Z(
        i_data_addr_gen_inst_N17) );
  INV_X1 i_data_addr_gen_inst_add_46_U1 ( .A(i_data_even_addr[0]), .ZN(
        i_data_addr_gen_inst_N8) );
  HA_X1 i_data_addr_gen_inst_add_46_U1_1_1 ( .A(i_data_even_addr[1]), .B(
        i_data_even_addr[0]), .CO(i_data_addr_gen_inst_add_46_carry[2]), .S(
        i_data_addr_gen_inst_N9) );
  HA_X1 i_data_addr_gen_inst_add_46_U1_1_2 ( .A(i_data_even_addr[2]), .B(
        i_data_addr_gen_inst_add_46_carry[2]), .CO(
        i_data_addr_gen_inst_add_46_carry[3]), .S(i_data_addr_gen_inst_N10) );
  HA_X1 i_data_addr_gen_inst_add_46_U1_1_3 ( .A(i_data_even_addr[3]), .B(
        i_data_addr_gen_inst_add_46_carry[3]), .CO(
        i_data_addr_gen_inst_add_46_carry[4]), .S(i_data_addr_gen_inst_N11) );
  HA_X1 i_data_addr_gen_inst_add_46_U1_1_4 ( .A(i_data_even_addr[4]), .B(
        i_data_addr_gen_inst_add_46_carry[4]), .CO(
        i_data_addr_gen_inst_add_46_carry[5]), .S(i_data_addr_gen_inst_N12) );
  HA_X1 i_data_addr_gen_inst_add_46_U1_1_5 ( .A(i_data_even_addr[5]), .B(
        i_data_addr_gen_inst_add_46_carry[5]), .CO(
        i_data_addr_gen_inst_add_46_carry[6]), .S(i_data_addr_gen_inst_N13) );
  HA_X1 i_data_addr_gen_inst_add_46_U1_1_6 ( .A(i_data_even_addr[6]), .B(
        i_data_addr_gen_inst_add_46_carry[6]), .CO(
        i_data_addr_gen_inst_add_46_carry[7]), .S(i_data_addr_gen_inst_N14) );
  HA_X1 i_data_addr_gen_inst_add_46_U1_1_7 ( .A(i_data_even_addr[7]), .B(
        i_data_addr_gen_inst_add_46_carry[7]), .CO(
        i_data_addr_gen_inst_add_46_carry[8]), .S(i_data_addr_gen_inst_N15) );
  HA_X1 i_data_addr_gen_inst_add_46_U1_1_8 ( .A(i_data_even_addr[8]), .B(
        i_data_addr_gen_inst_add_46_carry[8]), .CO(
        i_data_addr_gen_inst_add_46_carry[9]), .S(i_data_addr_gen_inst_N16) );
  XOR2_X1 i_data_addr_gen_inst_add_33_U2 ( .A(
        i_data_addr_gen_inst_int_data_offs_addr_0_), .B(
        i_data_addr_gen_inst_int_data_odd_base_addr[0]), .Z(i_data_odd_addr[0]) );
  AND2_X1 i_data_addr_gen_inst_add_33_U1 ( .A1(
        i_data_addr_gen_inst_int_data_offs_addr_0_), .A2(
        i_data_addr_gen_inst_int_data_odd_base_addr[0]), .ZN(
        i_data_addr_gen_inst_add_33_n1) );
  FA_X1 i_data_addr_gen_inst_add_33_U1_1 ( .A(
        i_data_addr_gen_inst_int_data_odd_base_addr[1]), .B(
        i_data_addr_gen_inst_int_data_offs_addr_1_), .CI(
        i_data_addr_gen_inst_add_33_n1), .CO(
        i_data_addr_gen_inst_add_33_carry[2]), .S(i_data_odd_addr[1]) );
  FA_X1 i_data_addr_gen_inst_add_33_U1_2 ( .A(
        i_data_addr_gen_inst_int_data_odd_base_addr[2]), .B(
        i_data_addr_gen_inst_int_data_offs_addr_2_), .CI(
        i_data_addr_gen_inst_add_33_carry[2]), .CO(
        i_data_addr_gen_inst_add_33_carry[3]), .S(i_data_odd_addr[2]) );
  FA_X1 i_data_addr_gen_inst_add_33_U1_3 ( .A(
        i_data_addr_gen_inst_int_data_odd_base_addr[3]), .B(
        i_data_addr_gen_inst_int_data_offs_addr_3_), .CI(
        i_data_addr_gen_inst_add_33_carry[3]), .CO(
        i_data_addr_gen_inst_add_33_carry[4]), .S(i_data_odd_addr[3]) );
  FA_X1 i_data_addr_gen_inst_add_33_U1_4 ( .A(
        i_data_addr_gen_inst_int_data_odd_base_addr[4]), .B(
        i_data_addr_gen_inst_int_data_offs_addr_4_), .CI(
        i_data_addr_gen_inst_add_33_carry[4]), .CO(
        i_data_addr_gen_inst_add_33_carry[5]), .S(i_data_odd_addr[4]) );
  FA_X1 i_data_addr_gen_inst_add_33_U1_5 ( .A(
        i_data_addr_gen_inst_int_data_odd_base_addr[5]), .B(
        i_data_addr_gen_inst_int_data_offs_addr_5_), .CI(
        i_data_addr_gen_inst_add_33_carry[5]), .CO(
        i_data_addr_gen_inst_add_33_carry[6]), .S(i_data_odd_addr[5]) );
  FA_X1 i_data_addr_gen_inst_add_33_U1_6 ( .A(
        i_data_addr_gen_inst_int_data_odd_base_addr[6]), .B(
        i_data_addr_gen_inst_int_data_offs_addr_6_), .CI(
        i_data_addr_gen_inst_add_33_carry[6]), .CO(
        i_data_addr_gen_inst_add_33_carry[7]), .S(i_data_odd_addr[6]) );
  FA_X1 i_data_addr_gen_inst_add_33_U1_7 ( .A(
        i_data_addr_gen_inst_int_data_odd_base_addr[7]), .B(
        i_data_addr_gen_inst_int_data_offs_addr_7_), .CI(
        i_data_addr_gen_inst_add_33_carry[7]), .CO(
        i_data_addr_gen_inst_add_33_carry[8]), .S(i_data_odd_addr[7]) );
  FA_X1 i_data_addr_gen_inst_add_33_U1_8 ( .A(
        i_data_addr_gen_inst_int_data_odd_base_addr[8]), .B(
        i_data_addr_gen_inst_int_data_offs_addr_8_), .CI(
        i_data_addr_gen_inst_add_33_carry[8]), .CO(
        i_data_addr_gen_inst_add_33_carry[9]), .S(i_data_odd_addr[8]) );
  FA_X1 i_data_addr_gen_inst_add_33_U1_9 ( .A(
        i_data_addr_gen_inst_int_data_odd_base_addr[9]), .B(
        i_data_addr_gen_inst_int_data_offs_addr_9_), .CI(
        i_data_addr_gen_inst_add_33_carry[9]), .S(i_data_odd_addr[9]) );
  XOR2_X1 i_data_addr_gen_inst_add_32_U2 ( .A(
        i_data_addr_gen_inst_int_data_offs_addr_0_), .B(
        i_data_addr_gen_inst_int_data_even_base_addr[0]), .Z(
        i_data_even_addr[0]) );
  AND2_X1 i_data_addr_gen_inst_add_32_U1 ( .A1(
        i_data_addr_gen_inst_int_data_offs_addr_0_), .A2(
        i_data_addr_gen_inst_int_data_even_base_addr[0]), .ZN(
        i_data_addr_gen_inst_add_32_n1) );
  FA_X1 i_data_addr_gen_inst_add_32_U1_1 ( .A(
        i_data_addr_gen_inst_int_data_even_base_addr[1]), .B(
        i_data_addr_gen_inst_int_data_offs_addr_1_), .CI(
        i_data_addr_gen_inst_add_32_n1), .CO(
        i_data_addr_gen_inst_add_32_carry[2]), .S(i_data_even_addr[1]) );
  FA_X1 i_data_addr_gen_inst_add_32_U1_2 ( .A(
        i_data_addr_gen_inst_int_data_even_base_addr[2]), .B(
        i_data_addr_gen_inst_int_data_offs_addr_2_), .CI(
        i_data_addr_gen_inst_add_32_carry[2]), .CO(
        i_data_addr_gen_inst_add_32_carry[3]), .S(i_data_even_addr[2]) );
  FA_X1 i_data_addr_gen_inst_add_32_U1_3 ( .A(
        i_data_addr_gen_inst_int_data_even_base_addr[3]), .B(
        i_data_addr_gen_inst_int_data_offs_addr_3_), .CI(
        i_data_addr_gen_inst_add_32_carry[3]), .CO(
        i_data_addr_gen_inst_add_32_carry[4]), .S(i_data_even_addr[3]) );
  FA_X1 i_data_addr_gen_inst_add_32_U1_4 ( .A(
        i_data_addr_gen_inst_int_data_even_base_addr[4]), .B(
        i_data_addr_gen_inst_int_data_offs_addr_4_), .CI(
        i_data_addr_gen_inst_add_32_carry[4]), .CO(
        i_data_addr_gen_inst_add_32_carry[5]), .S(i_data_even_addr[4]) );
  FA_X1 i_data_addr_gen_inst_add_32_U1_5 ( .A(
        i_data_addr_gen_inst_int_data_even_base_addr[5]), .B(
        i_data_addr_gen_inst_int_data_offs_addr_5_), .CI(
        i_data_addr_gen_inst_add_32_carry[5]), .CO(
        i_data_addr_gen_inst_add_32_carry[6]), .S(i_data_even_addr[5]) );
  FA_X1 i_data_addr_gen_inst_add_32_U1_6 ( .A(
        i_data_addr_gen_inst_int_data_even_base_addr[6]), .B(
        i_data_addr_gen_inst_int_data_offs_addr_6_), .CI(
        i_data_addr_gen_inst_add_32_carry[6]), .CO(
        i_data_addr_gen_inst_add_32_carry[7]), .S(i_data_even_addr[6]) );
  FA_X1 i_data_addr_gen_inst_add_32_U1_7 ( .A(
        i_data_addr_gen_inst_int_data_even_base_addr[7]), .B(
        i_data_addr_gen_inst_int_data_offs_addr_7_), .CI(
        i_data_addr_gen_inst_add_32_carry[7]), .CO(
        i_data_addr_gen_inst_add_32_carry[8]), .S(i_data_even_addr[7]) );
  FA_X1 i_data_addr_gen_inst_add_32_U1_8 ( .A(
        i_data_addr_gen_inst_int_data_even_base_addr[8]), .B(
        i_data_addr_gen_inst_int_data_offs_addr_8_), .CI(
        i_data_addr_gen_inst_add_32_carry[8]), .CO(
        i_data_addr_gen_inst_add_32_carry[9]), .S(i_data_even_addr[8]) );
  FA_X1 i_data_addr_gen_inst_add_32_U1_9 ( .A(
        i_data_addr_gen_inst_int_data_even_base_addr[9]), .B(
        i_data_addr_gen_inst_int_data_offs_addr_9_), .CI(
        i_data_addr_gen_inst_add_32_carry[9]), .S(i_data_even_addr[9]) );
  CLKBUF_X1 i_weight_addr_gen_inst_U41 ( .A(i_weight_addr_gen_inst_n37), .Z(
        i_weight_addr_gen_inst_n36) );
  CLKBUF_X1 i_weight_addr_gen_inst_U40 ( .A(i_weight_addr_gen_inst_n37), .Z(
        i_weight_addr_gen_inst_n35) );
  CLKBUF_X1 i_weight_addr_gen_inst_U39 ( .A(i_weight_addr_gen_inst_n37), .Z(
        i_weight_addr_gen_inst_n34) );
  OR2_X1 i_weight_addr_gen_inst_U38 ( .A1(ctrl_en_hmode), .A2(s_tc_res), .ZN(
        i_weight_addr_gen_inst_N38) );
  INV_X1 i_weight_addr_gen_inst_U37 ( .A(s_tc_res), .ZN(
        i_weight_addr_gen_inst_n38) );
  INV_X2 i_weight_addr_gen_inst_U3 ( .A(n9), .ZN(i_weight_addr_gen_inst_n37)
         );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_4_ ( .D(i_weight_addr[4]), 
        .CK(i_weight_addr_gen_inst_net2685), .RN(i_weight_addr_gen_inst_n37), 
        .Q(i_weight_addr_gen_inst_int_base_addr[4]) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_3_ ( .D(i_weight_addr[3]), 
        .CK(i_weight_addr_gen_inst_net2685), .RN(i_weight_addr_gen_inst_n37), 
        .Q(i_weight_addr_gen_inst_int_base_addr[3]) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_2_ ( .D(i_weight_addr[2]), 
        .CK(i_weight_addr_gen_inst_net2685), .RN(i_weight_addr_gen_inst_n37), 
        .Q(i_weight_addr_gen_inst_int_base_addr[2]) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_1_ ( .D(i_weight_addr[1]), 
        .CK(i_weight_addr_gen_inst_net2685), .RN(i_weight_addr_gen_inst_n37), 
        .Q(i_weight_addr_gen_inst_int_base_addr[1]) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_0_ ( .D(i_weight_addr[0]), 
        .CK(i_weight_addr_gen_inst_net2685), .RN(i_weight_addr_gen_inst_n37), 
        .Q(i_weight_addr_gen_inst_int_base_addr[0]) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_31_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n38), .SE(i_weight_addr_gen_inst_N37), .CK(
        i_weight_addr_gen_inst_net2691), .RN(i_weight_addr_gen_inst_n37), .Q(
        i_weight_addr_gen_inst_int_offs_addr_31_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_30_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n38), .SE(i_weight_addr_gen_inst_N36), .CK(
        i_weight_addr_gen_inst_net2691), .RN(i_weight_addr_gen_inst_n37), .Q(
        i_weight_addr_gen_inst_int_offs_addr_30_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_29_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n38), .SE(i_weight_addr_gen_inst_N35), .CK(
        i_weight_addr_gen_inst_net2691), .RN(i_weight_addr_gen_inst_n37), .Q(
        i_weight_addr_gen_inst_int_offs_addr_29_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_28_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n38), .SE(i_weight_addr_gen_inst_N34), .CK(
        i_weight_addr_gen_inst_net2691), .RN(i_weight_addr_gen_inst_n37), .Q(
        i_weight_addr_gen_inst_int_offs_addr_28_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_27_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n38), .SE(i_weight_addr_gen_inst_N33), .CK(
        i_weight_addr_gen_inst_net2691), .RN(i_weight_addr_gen_inst_n37), .Q(
        i_weight_addr_gen_inst_int_offs_addr_27_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_26_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n38), .SE(i_weight_addr_gen_inst_N32), .CK(
        i_weight_addr_gen_inst_net2691), .RN(i_weight_addr_gen_inst_n37), .Q(
        i_weight_addr_gen_inst_int_offs_addr_26_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_25_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n38), .SE(i_weight_addr_gen_inst_N31), .CK(
        i_weight_addr_gen_inst_net2691), .RN(i_weight_addr_gen_inst_n37), .Q(
        i_weight_addr_gen_inst_int_offs_addr_25_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_24_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n38), .SE(i_weight_addr_gen_inst_N30), .CK(
        i_weight_addr_gen_inst_net2691), .RN(i_weight_addr_gen_inst_n37), .Q(
        i_weight_addr_gen_inst_int_offs_addr_24_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_23_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n38), .SE(i_weight_addr_gen_inst_N29), .CK(
        i_weight_addr_gen_inst_net2691), .RN(i_weight_addr_gen_inst_n37), .Q(
        i_weight_addr_gen_inst_int_offs_addr_23_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_22_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n38), .SE(i_weight_addr_gen_inst_N28), .CK(
        i_weight_addr_gen_inst_net2691), .RN(i_weight_addr_gen_inst_n37), .Q(
        i_weight_addr_gen_inst_int_offs_addr_22_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_21_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n38), .SE(i_weight_addr_gen_inst_N27), .CK(
        i_weight_addr_gen_inst_net2691), .RN(i_weight_addr_gen_inst_n37), .Q(
        i_weight_addr_gen_inst_int_offs_addr_21_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_20_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n38), .SE(i_weight_addr_gen_inst_N26), .CK(
        i_weight_addr_gen_inst_net2691), .RN(i_weight_addr_gen_inst_n37), .Q(
        i_weight_addr_gen_inst_int_offs_addr_20_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_19_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n38), .SE(i_weight_addr_gen_inst_N25), .CK(
        i_weight_addr_gen_inst_net2691), .RN(i_weight_addr_gen_inst_n37), .Q(
        i_weight_addr_gen_inst_int_offs_addr_19_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_18_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n38), .SE(i_weight_addr_gen_inst_N24), .CK(
        i_weight_addr_gen_inst_net2691), .RN(i_weight_addr_gen_inst_n37), .Q(
        i_weight_addr_gen_inst_int_offs_addr_18_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_17_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n38), .SE(i_weight_addr_gen_inst_N23), .CK(
        i_weight_addr_gen_inst_net2691), .RN(i_weight_addr_gen_inst_n37), .Q(
        i_weight_addr_gen_inst_int_offs_addr_17_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_16_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n38), .SE(i_weight_addr_gen_inst_N22), .CK(
        i_weight_addr_gen_inst_net2691), .RN(i_weight_addr_gen_inst_n37), .Q(
        i_weight_addr_gen_inst_int_offs_addr_16_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_15_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n38), .SE(i_weight_addr_gen_inst_N21), .CK(
        i_weight_addr_gen_inst_net2691), .RN(i_weight_addr_gen_inst_n37), .Q(
        i_weight_addr_gen_inst_int_offs_addr_15_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_14_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n38), .SE(i_weight_addr_gen_inst_N20), .CK(
        i_weight_addr_gen_inst_net2691), .RN(i_weight_addr_gen_inst_n37), .Q(
        i_weight_addr_gen_inst_int_offs_addr_14_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_13_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n38), .SE(i_weight_addr_gen_inst_N19), .CK(
        i_weight_addr_gen_inst_net2691), .RN(i_weight_addr_gen_inst_n37), .Q(
        i_weight_addr_gen_inst_int_offs_addr_13_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_12_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n38), .SE(i_weight_addr_gen_inst_N18), .CK(
        i_weight_addr_gen_inst_net2691), .RN(i_weight_addr_gen_inst_n37), .Q(
        i_weight_addr_gen_inst_int_offs_addr_12_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_0_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n38), .SE(i_weight_addr_gen_inst_N6), .CK(
        i_weight_addr_gen_inst_net2691), .RN(i_weight_addr_gen_inst_n37), .Q(
        i_weight_addr_gen_inst_int_offs_addr_0_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_1_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n38), .SE(i_weight_addr_gen_inst_N7), .CK(
        i_weight_addr_gen_inst_net2691), .RN(i_weight_addr_gen_inst_n37), .Q(
        i_weight_addr_gen_inst_int_offs_addr_1_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_2_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n38), .SE(i_weight_addr_gen_inst_N8), .CK(
        i_weight_addr_gen_inst_net2691), .RN(i_weight_addr_gen_inst_n37), .Q(
        i_weight_addr_gen_inst_int_offs_addr_2_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_3_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n38), .SE(i_weight_addr_gen_inst_N9), .CK(
        i_weight_addr_gen_inst_net2691), .RN(i_weight_addr_gen_inst_n37), .Q(
        i_weight_addr_gen_inst_int_offs_addr_3_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_4_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n38), .SE(i_weight_addr_gen_inst_N10), .CK(
        i_weight_addr_gen_inst_net2691), .RN(i_weight_addr_gen_inst_n37), .Q(
        i_weight_addr_gen_inst_int_offs_addr_4_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_5_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n38), .SE(i_weight_addr_gen_inst_N11), .CK(
        i_weight_addr_gen_inst_net2691), .RN(i_weight_addr_gen_inst_n37), .Q(
        i_weight_addr_gen_inst_int_offs_addr_5_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_6_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n38), .SE(i_weight_addr_gen_inst_N12), .CK(
        i_weight_addr_gen_inst_net2691), .RN(i_weight_addr_gen_inst_n37), .Q(
        i_weight_addr_gen_inst_int_offs_addr_6_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_7_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n38), .SE(i_weight_addr_gen_inst_N13), .CK(
        i_weight_addr_gen_inst_net2691), .RN(i_weight_addr_gen_inst_n37), .Q(
        i_weight_addr_gen_inst_int_offs_addr_7_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_8_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n38), .SE(i_weight_addr_gen_inst_N14), .CK(
        i_weight_addr_gen_inst_net2691), .RN(i_weight_addr_gen_inst_n37), .Q(
        i_weight_addr_gen_inst_int_offs_addr_8_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_9_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n38), .SE(i_weight_addr_gen_inst_N15), .CK(
        i_weight_addr_gen_inst_net2691), .RN(i_weight_addr_gen_inst_n37), .Q(
        i_weight_addr_gen_inst_int_offs_addr_9_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_10_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n38), .SE(i_weight_addr_gen_inst_N16), .CK(
        i_weight_addr_gen_inst_net2691), .RN(i_weight_addr_gen_inst_n37), .Q(
        i_weight_addr_gen_inst_int_offs_addr_10_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_11_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n38), .SE(i_weight_addr_gen_inst_N17), .CK(
        i_weight_addr_gen_inst_net2691), .RN(i_weight_addr_gen_inst_n37), .Q(
        i_weight_addr_gen_inst_int_offs_addr_11_) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_31_ ( .D(i_weight_addr[31]), 
        .CK(i_weight_addr_gen_inst_net2685), .RN(i_weight_addr_gen_inst_n34), 
        .Q(i_weight_addr_gen_inst_int_base_addr[31]) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_30_ ( .D(i_weight_addr[30]), 
        .CK(i_weight_addr_gen_inst_net2685), .RN(i_weight_addr_gen_inst_n34), 
        .Q(i_weight_addr_gen_inst_int_base_addr[30]) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_29_ ( .D(i_weight_addr[29]), 
        .CK(i_weight_addr_gen_inst_net2685), .RN(i_weight_addr_gen_inst_n34), 
        .Q(i_weight_addr_gen_inst_int_base_addr[29]) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_28_ ( .D(i_weight_addr[28]), 
        .CK(i_weight_addr_gen_inst_net2685), .RN(i_weight_addr_gen_inst_n34), 
        .Q(i_weight_addr_gen_inst_int_base_addr[28]) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_27_ ( .D(i_weight_addr[27]), 
        .CK(i_weight_addr_gen_inst_net2685), .RN(i_weight_addr_gen_inst_n34), 
        .Q(i_weight_addr_gen_inst_int_base_addr[27]) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_26_ ( .D(i_weight_addr[26]), 
        .CK(i_weight_addr_gen_inst_net2685), .RN(i_weight_addr_gen_inst_n34), 
        .Q(i_weight_addr_gen_inst_int_base_addr[26]) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_25_ ( .D(i_weight_addr[25]), 
        .CK(i_weight_addr_gen_inst_net2685), .RN(i_weight_addr_gen_inst_n34), 
        .Q(i_weight_addr_gen_inst_int_base_addr[25]) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_24_ ( .D(i_weight_addr[24]), 
        .CK(i_weight_addr_gen_inst_net2685), .RN(i_weight_addr_gen_inst_n34), 
        .Q(i_weight_addr_gen_inst_int_base_addr[24]) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_23_ ( .D(i_weight_addr[23]), 
        .CK(i_weight_addr_gen_inst_net2685), .RN(i_weight_addr_gen_inst_n34), 
        .Q(i_weight_addr_gen_inst_int_base_addr[23]) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_22_ ( .D(i_weight_addr[22]), 
        .CK(i_weight_addr_gen_inst_net2685), .RN(i_weight_addr_gen_inst_n34), 
        .Q(i_weight_addr_gen_inst_int_base_addr[22]) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_21_ ( .D(i_weight_addr[21]), 
        .CK(i_weight_addr_gen_inst_net2685), .RN(i_weight_addr_gen_inst_n34), 
        .Q(i_weight_addr_gen_inst_int_base_addr[21]) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_20_ ( .D(i_weight_addr[20]), 
        .CK(i_weight_addr_gen_inst_net2685), .RN(i_weight_addr_gen_inst_n34), 
        .Q(i_weight_addr_gen_inst_int_base_addr[20]) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_19_ ( .D(i_weight_addr[19]), 
        .CK(i_weight_addr_gen_inst_net2685), .RN(i_weight_addr_gen_inst_n35), 
        .Q(i_weight_addr_gen_inst_int_base_addr[19]) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_18_ ( .D(i_weight_addr[18]), 
        .CK(i_weight_addr_gen_inst_net2685), .RN(i_weight_addr_gen_inst_n35), 
        .Q(i_weight_addr_gen_inst_int_base_addr[18]) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_17_ ( .D(i_weight_addr[17]), 
        .CK(i_weight_addr_gen_inst_net2685), .RN(i_weight_addr_gen_inst_n35), 
        .Q(i_weight_addr_gen_inst_int_base_addr[17]) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_16_ ( .D(i_weight_addr[16]), 
        .CK(i_weight_addr_gen_inst_net2685), .RN(i_weight_addr_gen_inst_n35), 
        .Q(i_weight_addr_gen_inst_int_base_addr[16]) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_15_ ( .D(i_weight_addr[15]), 
        .CK(i_weight_addr_gen_inst_net2685), .RN(i_weight_addr_gen_inst_n35), 
        .Q(i_weight_addr_gen_inst_int_base_addr[15]) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_14_ ( .D(i_weight_addr[14]), 
        .CK(i_weight_addr_gen_inst_net2685), .RN(i_weight_addr_gen_inst_n35), 
        .Q(i_weight_addr_gen_inst_int_base_addr[14]) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_13_ ( .D(i_weight_addr[13]), 
        .CK(i_weight_addr_gen_inst_net2685), .RN(i_weight_addr_gen_inst_n35), 
        .Q(i_weight_addr_gen_inst_int_base_addr[13]) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_12_ ( .D(i_weight_addr[12]), 
        .CK(i_weight_addr_gen_inst_net2685), .RN(i_weight_addr_gen_inst_n35), 
        .Q(i_weight_addr_gen_inst_int_base_addr[12]) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_11_ ( .D(i_weight_addr[11]), 
        .CK(i_weight_addr_gen_inst_net2685), .RN(i_weight_addr_gen_inst_n35), 
        .Q(i_weight_addr_gen_inst_int_base_addr[11]) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_10_ ( .D(i_weight_addr[10]), 
        .CK(i_weight_addr_gen_inst_net2685), .RN(i_weight_addr_gen_inst_n35), 
        .Q(i_weight_addr_gen_inst_int_base_addr[10]) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_9_ ( .D(i_weight_addr[9]), 
        .CK(i_weight_addr_gen_inst_net2685), .RN(i_weight_addr_gen_inst_n35), 
        .Q(i_weight_addr_gen_inst_int_base_addr[9]) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_8_ ( .D(i_weight_addr[8]), 
        .CK(i_weight_addr_gen_inst_net2685), .RN(i_weight_addr_gen_inst_n35), 
        .Q(i_weight_addr_gen_inst_int_base_addr[8]) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_7_ ( .D(i_weight_addr[7]), 
        .CK(i_weight_addr_gen_inst_net2685), .RN(i_weight_addr_gen_inst_n36), 
        .Q(i_weight_addr_gen_inst_int_base_addr[7]) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_6_ ( .D(i_weight_addr[6]), 
        .CK(i_weight_addr_gen_inst_net2685), .RN(i_weight_addr_gen_inst_n36), 
        .Q(i_weight_addr_gen_inst_int_base_addr[6]) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_5_ ( .D(i_weight_addr[5]), 
        .CK(i_weight_addr_gen_inst_net2685), .RN(i_weight_addr_gen_inst_n36), 
        .Q(i_weight_addr_gen_inst_int_base_addr[5]) );
  CLKGATETST_X1 i_weight_addr_gen_inst_clk_gate_int_base_addr_reg_latch ( .CK(
        ck), .E(int_inc_i_w_addr), .SE(1'b0), .GCK(
        i_weight_addr_gen_inst_net2685) );
  CLKGATETST_X1 i_weight_addr_gen_inst_clk_gate_int_offs_addr_reg_latch ( .CK(
        ck), .E(i_weight_addr_gen_inst_N38), .SE(1'b0), .GCK(
        i_weight_addr_gen_inst_net2691) );
  XOR2_X1 i_weight_addr_gen_inst_add_49_U2 ( .A(
        i_weight_addr_gen_inst_add_49_carry[31]), .B(
        i_weight_addr_gen_inst_int_offs_addr_31_), .Z(
        i_weight_addr_gen_inst_N37) );
  INV_X1 i_weight_addr_gen_inst_add_49_U1 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_0_), .ZN(
        i_weight_addr_gen_inst_N6) );
  HA_X1 i_weight_addr_gen_inst_add_49_U1_1_1 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_1_), .B(
        i_weight_addr_gen_inst_int_offs_addr_0_), .CO(
        i_weight_addr_gen_inst_add_49_carry[2]), .S(i_weight_addr_gen_inst_N7)
         );
  HA_X1 i_weight_addr_gen_inst_add_49_U1_1_2 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_2_), .B(
        i_weight_addr_gen_inst_add_49_carry[2]), .CO(
        i_weight_addr_gen_inst_add_49_carry[3]), .S(i_weight_addr_gen_inst_N8)
         );
  HA_X1 i_weight_addr_gen_inst_add_49_U1_1_3 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_3_), .B(
        i_weight_addr_gen_inst_add_49_carry[3]), .CO(
        i_weight_addr_gen_inst_add_49_carry[4]), .S(i_weight_addr_gen_inst_N9)
         );
  HA_X1 i_weight_addr_gen_inst_add_49_U1_1_4 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_4_), .B(
        i_weight_addr_gen_inst_add_49_carry[4]), .CO(
        i_weight_addr_gen_inst_add_49_carry[5]), .S(i_weight_addr_gen_inst_N10) );
  HA_X1 i_weight_addr_gen_inst_add_49_U1_1_5 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_5_), .B(
        i_weight_addr_gen_inst_add_49_carry[5]), .CO(
        i_weight_addr_gen_inst_add_49_carry[6]), .S(i_weight_addr_gen_inst_N11) );
  HA_X1 i_weight_addr_gen_inst_add_49_U1_1_6 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_6_), .B(
        i_weight_addr_gen_inst_add_49_carry[6]), .CO(
        i_weight_addr_gen_inst_add_49_carry[7]), .S(i_weight_addr_gen_inst_N12) );
  HA_X1 i_weight_addr_gen_inst_add_49_U1_1_7 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_7_), .B(
        i_weight_addr_gen_inst_add_49_carry[7]), .CO(
        i_weight_addr_gen_inst_add_49_carry[8]), .S(i_weight_addr_gen_inst_N13) );
  HA_X1 i_weight_addr_gen_inst_add_49_U1_1_8 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_8_), .B(
        i_weight_addr_gen_inst_add_49_carry[8]), .CO(
        i_weight_addr_gen_inst_add_49_carry[9]), .S(i_weight_addr_gen_inst_N14) );
  HA_X1 i_weight_addr_gen_inst_add_49_U1_1_9 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_9_), .B(
        i_weight_addr_gen_inst_add_49_carry[9]), .CO(
        i_weight_addr_gen_inst_add_49_carry[10]), .S(
        i_weight_addr_gen_inst_N15) );
  HA_X1 i_weight_addr_gen_inst_add_49_U1_1_10 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_10_), .B(
        i_weight_addr_gen_inst_add_49_carry[10]), .CO(
        i_weight_addr_gen_inst_add_49_carry[11]), .S(
        i_weight_addr_gen_inst_N16) );
  HA_X1 i_weight_addr_gen_inst_add_49_U1_1_11 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_11_), .B(
        i_weight_addr_gen_inst_add_49_carry[11]), .CO(
        i_weight_addr_gen_inst_add_49_carry[12]), .S(
        i_weight_addr_gen_inst_N17) );
  HA_X1 i_weight_addr_gen_inst_add_49_U1_1_12 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_12_), .B(
        i_weight_addr_gen_inst_add_49_carry[12]), .CO(
        i_weight_addr_gen_inst_add_49_carry[13]), .S(
        i_weight_addr_gen_inst_N18) );
  HA_X1 i_weight_addr_gen_inst_add_49_U1_1_13 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_13_), .B(
        i_weight_addr_gen_inst_add_49_carry[13]), .CO(
        i_weight_addr_gen_inst_add_49_carry[14]), .S(
        i_weight_addr_gen_inst_N19) );
  HA_X1 i_weight_addr_gen_inst_add_49_U1_1_14 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_14_), .B(
        i_weight_addr_gen_inst_add_49_carry[14]), .CO(
        i_weight_addr_gen_inst_add_49_carry[15]), .S(
        i_weight_addr_gen_inst_N20) );
  HA_X1 i_weight_addr_gen_inst_add_49_U1_1_15 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_15_), .B(
        i_weight_addr_gen_inst_add_49_carry[15]), .CO(
        i_weight_addr_gen_inst_add_49_carry[16]), .S(
        i_weight_addr_gen_inst_N21) );
  HA_X1 i_weight_addr_gen_inst_add_49_U1_1_16 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_16_), .B(
        i_weight_addr_gen_inst_add_49_carry[16]), .CO(
        i_weight_addr_gen_inst_add_49_carry[17]), .S(
        i_weight_addr_gen_inst_N22) );
  HA_X1 i_weight_addr_gen_inst_add_49_U1_1_17 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_17_), .B(
        i_weight_addr_gen_inst_add_49_carry[17]), .CO(
        i_weight_addr_gen_inst_add_49_carry[18]), .S(
        i_weight_addr_gen_inst_N23) );
  HA_X1 i_weight_addr_gen_inst_add_49_U1_1_18 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_18_), .B(
        i_weight_addr_gen_inst_add_49_carry[18]), .CO(
        i_weight_addr_gen_inst_add_49_carry[19]), .S(
        i_weight_addr_gen_inst_N24) );
  HA_X1 i_weight_addr_gen_inst_add_49_U1_1_19 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_19_), .B(
        i_weight_addr_gen_inst_add_49_carry[19]), .CO(
        i_weight_addr_gen_inst_add_49_carry[20]), .S(
        i_weight_addr_gen_inst_N25) );
  HA_X1 i_weight_addr_gen_inst_add_49_U1_1_20 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_20_), .B(
        i_weight_addr_gen_inst_add_49_carry[20]), .CO(
        i_weight_addr_gen_inst_add_49_carry[21]), .S(
        i_weight_addr_gen_inst_N26) );
  HA_X1 i_weight_addr_gen_inst_add_49_U1_1_21 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_21_), .B(
        i_weight_addr_gen_inst_add_49_carry[21]), .CO(
        i_weight_addr_gen_inst_add_49_carry[22]), .S(
        i_weight_addr_gen_inst_N27) );
  HA_X1 i_weight_addr_gen_inst_add_49_U1_1_22 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_22_), .B(
        i_weight_addr_gen_inst_add_49_carry[22]), .CO(
        i_weight_addr_gen_inst_add_49_carry[23]), .S(
        i_weight_addr_gen_inst_N28) );
  HA_X1 i_weight_addr_gen_inst_add_49_U1_1_23 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_23_), .B(
        i_weight_addr_gen_inst_add_49_carry[23]), .CO(
        i_weight_addr_gen_inst_add_49_carry[24]), .S(
        i_weight_addr_gen_inst_N29) );
  HA_X1 i_weight_addr_gen_inst_add_49_U1_1_24 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_24_), .B(
        i_weight_addr_gen_inst_add_49_carry[24]), .CO(
        i_weight_addr_gen_inst_add_49_carry[25]), .S(
        i_weight_addr_gen_inst_N30) );
  HA_X1 i_weight_addr_gen_inst_add_49_U1_1_25 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_25_), .B(
        i_weight_addr_gen_inst_add_49_carry[25]), .CO(
        i_weight_addr_gen_inst_add_49_carry[26]), .S(
        i_weight_addr_gen_inst_N31) );
  HA_X1 i_weight_addr_gen_inst_add_49_U1_1_26 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_26_), .B(
        i_weight_addr_gen_inst_add_49_carry[26]), .CO(
        i_weight_addr_gen_inst_add_49_carry[27]), .S(
        i_weight_addr_gen_inst_N32) );
  HA_X1 i_weight_addr_gen_inst_add_49_U1_1_27 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_27_), .B(
        i_weight_addr_gen_inst_add_49_carry[27]), .CO(
        i_weight_addr_gen_inst_add_49_carry[28]), .S(
        i_weight_addr_gen_inst_N33) );
  HA_X1 i_weight_addr_gen_inst_add_49_U1_1_28 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_28_), .B(
        i_weight_addr_gen_inst_add_49_carry[28]), .CO(
        i_weight_addr_gen_inst_add_49_carry[29]), .S(
        i_weight_addr_gen_inst_N34) );
  HA_X1 i_weight_addr_gen_inst_add_49_U1_1_29 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_29_), .B(
        i_weight_addr_gen_inst_add_49_carry[29]), .CO(
        i_weight_addr_gen_inst_add_49_carry[30]), .S(
        i_weight_addr_gen_inst_N35) );
  HA_X1 i_weight_addr_gen_inst_add_49_U1_1_30 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_30_), .B(
        i_weight_addr_gen_inst_add_49_carry[30]), .CO(
        i_weight_addr_gen_inst_add_49_carry[31]), .S(
        i_weight_addr_gen_inst_N36) );
  XOR2_X1 i_weight_addr_gen_inst_add_26_U2 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_0_), .B(
        i_weight_addr_gen_inst_int_base_addr[0]), .Z(i_weight_addr[0]) );
  AND2_X1 i_weight_addr_gen_inst_add_26_U1 ( .A1(
        i_weight_addr_gen_inst_int_offs_addr_0_), .A2(
        i_weight_addr_gen_inst_int_base_addr[0]), .ZN(
        i_weight_addr_gen_inst_add_26_n1) );
  FA_X1 i_weight_addr_gen_inst_add_26_U1_1 ( .A(
        i_weight_addr_gen_inst_int_base_addr[1]), .B(
        i_weight_addr_gen_inst_int_offs_addr_1_), .CI(
        i_weight_addr_gen_inst_add_26_n1), .CO(
        i_weight_addr_gen_inst_add_26_carry[2]), .S(i_weight_addr[1]) );
  FA_X1 i_weight_addr_gen_inst_add_26_U1_2 ( .A(
        i_weight_addr_gen_inst_int_base_addr[2]), .B(
        i_weight_addr_gen_inst_int_offs_addr_2_), .CI(
        i_weight_addr_gen_inst_add_26_carry[2]), .CO(
        i_weight_addr_gen_inst_add_26_carry[3]), .S(i_weight_addr[2]) );
  FA_X1 i_weight_addr_gen_inst_add_26_U1_3 ( .A(
        i_weight_addr_gen_inst_int_base_addr[3]), .B(
        i_weight_addr_gen_inst_int_offs_addr_3_), .CI(
        i_weight_addr_gen_inst_add_26_carry[3]), .CO(
        i_weight_addr_gen_inst_add_26_carry[4]), .S(i_weight_addr[3]) );
  FA_X1 i_weight_addr_gen_inst_add_26_U1_4 ( .A(
        i_weight_addr_gen_inst_int_base_addr[4]), .B(
        i_weight_addr_gen_inst_int_offs_addr_4_), .CI(
        i_weight_addr_gen_inst_add_26_carry[4]), .CO(
        i_weight_addr_gen_inst_add_26_carry[5]), .S(i_weight_addr[4]) );
  FA_X1 i_weight_addr_gen_inst_add_26_U1_5 ( .A(
        i_weight_addr_gen_inst_int_base_addr[5]), .B(
        i_weight_addr_gen_inst_int_offs_addr_5_), .CI(
        i_weight_addr_gen_inst_add_26_carry[5]), .CO(
        i_weight_addr_gen_inst_add_26_carry[6]), .S(i_weight_addr[5]) );
  FA_X1 i_weight_addr_gen_inst_add_26_U1_6 ( .A(
        i_weight_addr_gen_inst_int_base_addr[6]), .B(
        i_weight_addr_gen_inst_int_offs_addr_6_), .CI(
        i_weight_addr_gen_inst_add_26_carry[6]), .CO(
        i_weight_addr_gen_inst_add_26_carry[7]), .S(i_weight_addr[6]) );
  FA_X1 i_weight_addr_gen_inst_add_26_U1_7 ( .A(
        i_weight_addr_gen_inst_int_base_addr[7]), .B(
        i_weight_addr_gen_inst_int_offs_addr_7_), .CI(
        i_weight_addr_gen_inst_add_26_carry[7]), .CO(
        i_weight_addr_gen_inst_add_26_carry[8]), .S(i_weight_addr[7]) );
  FA_X1 i_weight_addr_gen_inst_add_26_U1_8 ( .A(
        i_weight_addr_gen_inst_int_base_addr[8]), .B(
        i_weight_addr_gen_inst_int_offs_addr_8_), .CI(
        i_weight_addr_gen_inst_add_26_carry[8]), .CO(
        i_weight_addr_gen_inst_add_26_carry[9]), .S(i_weight_addr[8]) );
  FA_X1 i_weight_addr_gen_inst_add_26_U1_9 ( .A(
        i_weight_addr_gen_inst_int_base_addr[9]), .B(
        i_weight_addr_gen_inst_int_offs_addr_9_), .CI(
        i_weight_addr_gen_inst_add_26_carry[9]), .CO(
        i_weight_addr_gen_inst_add_26_carry[10]), .S(i_weight_addr[9]) );
  FA_X1 i_weight_addr_gen_inst_add_26_U1_10 ( .A(
        i_weight_addr_gen_inst_int_base_addr[10]), .B(
        i_weight_addr_gen_inst_int_offs_addr_10_), .CI(
        i_weight_addr_gen_inst_add_26_carry[10]), .CO(
        i_weight_addr_gen_inst_add_26_carry[11]), .S(i_weight_addr[10]) );
  FA_X1 i_weight_addr_gen_inst_add_26_U1_11 ( .A(
        i_weight_addr_gen_inst_int_base_addr[11]), .B(
        i_weight_addr_gen_inst_int_offs_addr_11_), .CI(
        i_weight_addr_gen_inst_add_26_carry[11]), .CO(
        i_weight_addr_gen_inst_add_26_carry[12]), .S(i_weight_addr[11]) );
  FA_X1 i_weight_addr_gen_inst_add_26_U1_12 ( .A(
        i_weight_addr_gen_inst_int_base_addr[12]), .B(
        i_weight_addr_gen_inst_int_offs_addr_12_), .CI(
        i_weight_addr_gen_inst_add_26_carry[12]), .CO(
        i_weight_addr_gen_inst_add_26_carry[13]), .S(i_weight_addr[12]) );
  FA_X1 i_weight_addr_gen_inst_add_26_U1_13 ( .A(
        i_weight_addr_gen_inst_int_base_addr[13]), .B(
        i_weight_addr_gen_inst_int_offs_addr_13_), .CI(
        i_weight_addr_gen_inst_add_26_carry[13]), .CO(
        i_weight_addr_gen_inst_add_26_carry[14]), .S(i_weight_addr[13]) );
  FA_X1 i_weight_addr_gen_inst_add_26_U1_14 ( .A(
        i_weight_addr_gen_inst_int_base_addr[14]), .B(
        i_weight_addr_gen_inst_int_offs_addr_14_), .CI(
        i_weight_addr_gen_inst_add_26_carry[14]), .CO(
        i_weight_addr_gen_inst_add_26_carry[15]), .S(i_weight_addr[14]) );
  FA_X1 i_weight_addr_gen_inst_add_26_U1_15 ( .A(
        i_weight_addr_gen_inst_int_base_addr[15]), .B(
        i_weight_addr_gen_inst_int_offs_addr_15_), .CI(
        i_weight_addr_gen_inst_add_26_carry[15]), .CO(
        i_weight_addr_gen_inst_add_26_carry[16]), .S(i_weight_addr[15]) );
  FA_X1 i_weight_addr_gen_inst_add_26_U1_16 ( .A(
        i_weight_addr_gen_inst_int_base_addr[16]), .B(
        i_weight_addr_gen_inst_int_offs_addr_16_), .CI(
        i_weight_addr_gen_inst_add_26_carry[16]), .CO(
        i_weight_addr_gen_inst_add_26_carry[17]), .S(i_weight_addr[16]) );
  FA_X1 i_weight_addr_gen_inst_add_26_U1_17 ( .A(
        i_weight_addr_gen_inst_int_base_addr[17]), .B(
        i_weight_addr_gen_inst_int_offs_addr_17_), .CI(
        i_weight_addr_gen_inst_add_26_carry[17]), .CO(
        i_weight_addr_gen_inst_add_26_carry[18]), .S(i_weight_addr[17]) );
  FA_X1 i_weight_addr_gen_inst_add_26_U1_18 ( .A(
        i_weight_addr_gen_inst_int_base_addr[18]), .B(
        i_weight_addr_gen_inst_int_offs_addr_18_), .CI(
        i_weight_addr_gen_inst_add_26_carry[18]), .CO(
        i_weight_addr_gen_inst_add_26_carry[19]), .S(i_weight_addr[18]) );
  FA_X1 i_weight_addr_gen_inst_add_26_U1_19 ( .A(
        i_weight_addr_gen_inst_int_base_addr[19]), .B(
        i_weight_addr_gen_inst_int_offs_addr_19_), .CI(
        i_weight_addr_gen_inst_add_26_carry[19]), .CO(
        i_weight_addr_gen_inst_add_26_carry[20]), .S(i_weight_addr[19]) );
  FA_X1 i_weight_addr_gen_inst_add_26_U1_20 ( .A(
        i_weight_addr_gen_inst_int_base_addr[20]), .B(
        i_weight_addr_gen_inst_int_offs_addr_20_), .CI(
        i_weight_addr_gen_inst_add_26_carry[20]), .CO(
        i_weight_addr_gen_inst_add_26_carry[21]), .S(i_weight_addr[20]) );
  FA_X1 i_weight_addr_gen_inst_add_26_U1_21 ( .A(
        i_weight_addr_gen_inst_int_base_addr[21]), .B(
        i_weight_addr_gen_inst_int_offs_addr_21_), .CI(
        i_weight_addr_gen_inst_add_26_carry[21]), .CO(
        i_weight_addr_gen_inst_add_26_carry[22]), .S(i_weight_addr[21]) );
  FA_X1 i_weight_addr_gen_inst_add_26_U1_22 ( .A(
        i_weight_addr_gen_inst_int_base_addr[22]), .B(
        i_weight_addr_gen_inst_int_offs_addr_22_), .CI(
        i_weight_addr_gen_inst_add_26_carry[22]), .CO(
        i_weight_addr_gen_inst_add_26_carry[23]), .S(i_weight_addr[22]) );
  FA_X1 i_weight_addr_gen_inst_add_26_U1_23 ( .A(
        i_weight_addr_gen_inst_int_base_addr[23]), .B(
        i_weight_addr_gen_inst_int_offs_addr_23_), .CI(
        i_weight_addr_gen_inst_add_26_carry[23]), .CO(
        i_weight_addr_gen_inst_add_26_carry[24]), .S(i_weight_addr[23]) );
  FA_X1 i_weight_addr_gen_inst_add_26_U1_24 ( .A(
        i_weight_addr_gen_inst_int_base_addr[24]), .B(
        i_weight_addr_gen_inst_int_offs_addr_24_), .CI(
        i_weight_addr_gen_inst_add_26_carry[24]), .CO(
        i_weight_addr_gen_inst_add_26_carry[25]), .S(i_weight_addr[24]) );
  FA_X1 i_weight_addr_gen_inst_add_26_U1_25 ( .A(
        i_weight_addr_gen_inst_int_base_addr[25]), .B(
        i_weight_addr_gen_inst_int_offs_addr_25_), .CI(
        i_weight_addr_gen_inst_add_26_carry[25]), .CO(
        i_weight_addr_gen_inst_add_26_carry[26]), .S(i_weight_addr[25]) );
  FA_X1 i_weight_addr_gen_inst_add_26_U1_26 ( .A(
        i_weight_addr_gen_inst_int_base_addr[26]), .B(
        i_weight_addr_gen_inst_int_offs_addr_26_), .CI(
        i_weight_addr_gen_inst_add_26_carry[26]), .CO(
        i_weight_addr_gen_inst_add_26_carry[27]), .S(i_weight_addr[26]) );
  FA_X1 i_weight_addr_gen_inst_add_26_U1_27 ( .A(
        i_weight_addr_gen_inst_int_base_addr[27]), .B(
        i_weight_addr_gen_inst_int_offs_addr_27_), .CI(
        i_weight_addr_gen_inst_add_26_carry[27]), .CO(
        i_weight_addr_gen_inst_add_26_carry[28]), .S(i_weight_addr[27]) );
  FA_X1 i_weight_addr_gen_inst_add_26_U1_28 ( .A(
        i_weight_addr_gen_inst_int_base_addr[28]), .B(
        i_weight_addr_gen_inst_int_offs_addr_28_), .CI(
        i_weight_addr_gen_inst_add_26_carry[28]), .CO(
        i_weight_addr_gen_inst_add_26_carry[29]), .S(i_weight_addr[28]) );
  FA_X1 i_weight_addr_gen_inst_add_26_U1_29 ( .A(
        i_weight_addr_gen_inst_int_base_addr[29]), .B(
        i_weight_addr_gen_inst_int_offs_addr_29_), .CI(
        i_weight_addr_gen_inst_add_26_carry[29]), .CO(
        i_weight_addr_gen_inst_add_26_carry[30]), .S(i_weight_addr[29]) );
  FA_X1 i_weight_addr_gen_inst_add_26_U1_30 ( .A(
        i_weight_addr_gen_inst_int_base_addr[30]), .B(
        i_weight_addr_gen_inst_int_offs_addr_30_), .CI(
        i_weight_addr_gen_inst_add_26_carry[30]), .CO(
        i_weight_addr_gen_inst_add_26_carry[31]), .S(i_weight_addr[30]) );
  FA_X1 i_weight_addr_gen_inst_add_26_U1_31 ( .A(
        i_weight_addr_gen_inst_int_base_addr[31]), .B(
        i_weight_addr_gen_inst_int_offs_addr_31_), .CI(
        i_weight_addr_gen_inst_add_26_carry[31]), .S(i_weight_addr[31]) );
  CLKGATETST_X1 clk_gate_int_i_data_v_npu_reg_latch ( .CK(ck), .E(ctrl_ldh_v_n), .SE(1'b0), .GCK(net2652) );
  CLKGATETST_X1 clk_gate_int_q_tc_reg_latch ( .CK(ck), .E(s_tc_res), .SE(1'b0), 
        .GCK(net2658) );
  CLKGATETST_X1 clk_gate_int_o_data_odd_addr_reg_latch ( .CK(ck), .E(N28), 
        .SE(1'b0), .GCK(net2663) );
  CLKGATETST_X1 clk_gate_int_o_data_even_addr_reg_latch ( .CK(ck), .E(N27), 
        .SE(1'b0), .GCK(net2668) );
  XOR2_X1 add_428_U2 ( .A(add_428_carry[9]), .B(o_data_even_addr[9]), .Z(N26)
         );
  INV_X1 add_428_U1 ( .A(o_data_even_addr[0]), .ZN(N17) );
  HA_X1 add_428_U1_1_1 ( .A(o_data_even_addr[1]), .B(o_data_even_addr[0]), 
        .CO(add_428_carry[2]), .S(N18) );
  HA_X1 add_428_U1_1_2 ( .A(o_data_even_addr[2]), .B(add_428_carry[2]), .CO(
        add_428_carry[3]), .S(N19) );
  HA_X1 add_428_U1_1_3 ( .A(o_data_even_addr[3]), .B(add_428_carry[3]), .CO(
        add_428_carry[4]), .S(N20) );
  HA_X1 add_428_U1_1_4 ( .A(o_data_even_addr[4]), .B(add_428_carry[4]), .CO(
        add_428_carry[5]), .S(N21) );
  HA_X1 add_428_U1_1_5 ( .A(o_data_even_addr[5]), .B(add_428_carry[5]), .CO(
        add_428_carry[6]), .S(N22) );
  HA_X1 add_428_U1_1_6 ( .A(o_data_even_addr[6]), .B(add_428_carry[6]), .CO(
        add_428_carry[7]), .S(N23) );
  HA_X1 add_428_U1_1_7 ( .A(o_data_even_addr[7]), .B(add_428_carry[7]), .CO(
        add_428_carry[8]), .S(N24) );
  HA_X1 add_428_U1_1_8 ( .A(o_data_even_addr[8]), .B(add_428_carry[8]), .CO(
        add_428_carry[9]), .S(N25) );
  XOR2_X1 add_426_U2 ( .A(add_426_carry[9]), .B(o_data_odd_addr[9]), .Z(N16)
         );
  INV_X1 add_426_U1 ( .A(o_data_odd_addr[0]), .ZN(N7) );
  HA_X1 add_426_U1_1_1 ( .A(o_data_odd_addr[1]), .B(o_data_odd_addr[0]), .CO(
        add_426_carry[2]), .S(N8) );
  HA_X1 add_426_U1_1_2 ( .A(o_data_odd_addr[2]), .B(add_426_carry[2]), .CO(
        add_426_carry[3]), .S(N9) );
  HA_X1 add_426_U1_1_3 ( .A(o_data_odd_addr[3]), .B(add_426_carry[3]), .CO(
        add_426_carry[4]), .S(N10) );
  HA_X1 add_426_U1_1_4 ( .A(o_data_odd_addr[4]), .B(add_426_carry[4]), .CO(
        add_426_carry[5]), .S(N11) );
  HA_X1 add_426_U1_1_5 ( .A(o_data_odd_addr[5]), .B(add_426_carry[5]), .CO(
        add_426_carry[6]), .S(N12) );
  HA_X1 add_426_U1_1_6 ( .A(o_data_odd_addr[6]), .B(add_426_carry[6]), .CO(
        add_426_carry[7]), .S(N13) );
  HA_X1 add_426_U1_1_7 ( .A(o_data_odd_addr[7]), .B(add_426_carry[7]), .CO(
        add_426_carry[8]), .S(N14) );
  HA_X1 add_426_U1_1_8 ( .A(o_data_odd_addr[8]), .B(add_426_carry[8]), .CO(
        add_426_carry[9]), .S(N15) );
endmodule

