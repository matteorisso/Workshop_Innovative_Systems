library verilog;
use verilog.vl_types.all;
entity test_sv_unit is
end test_sv_unit;
