library ieee;
use ieee.std_logic_1164.all;
use work.fixed_pkg.all;

entity RALU is
generic ( 	qi : natural:= 8;
				qf : natural:= 8 );			
    port (
	 
          AD : in sfixed(qi-1 downto -qf);
          OT : out sfixed(qi-1 downto -qf)
         );
end entity;

architecture behavioral of RALU is

begin

OT <=  "0000000000000111" when (AD > "0000000001100110") and (AD <= "0000000010000000") else 
       "0000000000001100" when (AD > "0000000010000000") and (AD <= "0000000010011001") else
       "0000000000010100" when (AD > "0000000010011001") and (AD <= "0000000010110011") else         
       "0000000000011101" when (AD > "0000000010110011") and (AD <= "0000000011001100") else       
       "0000000000101000" when (AD > "0000000011001100") and (AD <= "0000000011100110") else       
       "0000000000110110" when (AD > "0000000011100110") and (AD <= "0000000100011001") else      
       "0000000000101110" when (AD > "0000000100011001") and (AD <= "0000000100110011") else     
       "0000000000100111" when (AD > "0000000100110011") and (AD <= "0000000101001100") else        
       "0000000000100000" when (AD > "0000000101001100") and (AD <= "0000000101100110") else  
       "0000000000011010" when (AD > "0000000101100110") and (AD <= "0000000110000000") else      
       "0000000000010101" when (AD > "0000000110000000") and (AD <= "0000000110011001") else         
       "0000000000010010" when (AD > "0000000110011001") and (AD <= "0000000110110011") else   
       "0000000000001111" when (AD > "0000000110110011") and (AD <= "0000000111001100") else    
       "0000000000001100" when (AD > "0000000111001100") and (AD <= "0000000111100110") else      
       "0000000000001100" when (AD > "0000000111001100") and (AD <= "0000000111100110") else 
       "0000000000001001" when (AD > "0000000111100110") and (AD <= "0000001000000000") else 
       "0000000000000000"; 
 
end architecture; 